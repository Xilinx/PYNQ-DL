`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner="Xilinx"
`protect key_method="rsa"
`protect key_keyname="xilinxt_2017_05"
`protect key_block
BwcgdCG4trl440t2KEmRpuf6QWQ/1MWxHn1PJvcEQxshsu/1eQBlUvlysaB8VF3OzORoNbb5ZvyY
R+TtbOoqPHdbUQ16Ay3Y09W5312NJg3ULW0gFCOySXWIMP9ur5hqOBwf7wa0OnF4NMMWMp5e5g6u
D9re48GSrAOCz4UMQvt/YsZTeqp1P1jnCOBoscRTzBPLcrpIQAXoUaByeZOcpDKaM8XHbSXFsZD8
3p/AyiI5a1KJ8r6fAEkOtjIKZIEU1l62ZxFuG1dcMlTmdpce1fKnbfwD2ZTqOVfiIOg9hZA/qvVn
Zizngh+z2AeyU9opRZjypg87Ut+2h5vSMcIDoQ==

`protect control xilinx_enable_probing="false"
`protect control xilinx_enable_bitstream="true"
`protect control xilinx_enable_netlist_export="false"
`protect control xilinx_enable_modification="false"
`protect control xilinx_configuration_visible="false"
`protect rights_digest_method="sha256"
`protect end_toolblock="EA/0gL5DSj+qIyeb6TyITkqBV2GDWgivWUra9t8PKCA="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1818016)
`protect data_block
Hg5KTSInq2NkvmerKPTvVsTIvVpXGAZxVQGKvS9w+IoZt3Ok+9sRI3IrOvNbvIE06fTNXeq5MXR3
8v1291mhrdwxZ+1iqHvtoz4nLDHQht7Q5ZxGivEpfuq+dGhdRBiUDGsBA0j1qrCrI4/ASym5dk9Y
KWHa5NEzJwKdohhU2q6M60AkphDL4Wa/6Zkp6STJlRMJo5peIRPzwqz8JvSYCOrmlr6q+apI6n59
7+P0A9/bDeoLkGxHe4chIJyycjlWr5cXpEIMUdkQOIjpfT+3gri83ha0H56w4XolADLRj7do1muF
BAVwYUpcOW2IGlQdgYJ3sLgohhhLZLqbwHZ8ADhUGzQLtA8NzvPGQvTRJ07fet3Spq0NJhtq0ori
DZ+NhPBqdD2j1RrH0ePbhrqIHv/OtcBql83+uzkK9SX6l32UoxGcFt77owc/gggpQEACsPKlqh9I
pNlGmQsR6n+VSe62QZWHVuD9gou+1RAbPBDeejRo8KQe4nJPzOJkT2hPUqixUsacgW/ldStBlChl
oo+dfTnKOTyTpEgZSppZCkkevaZp214SEDb2C6OBpNimkDSCxHUaa17RegIs8ocJk3+f5wdaeV4M
6mN99NMUPC2VSFJtIUtj1/MqAbogKKrhn9xARZMOTNLSHUoMKI5o6mkNMC1ygfAMnSzrYDktCh1V
WYpgZA73juyB7RDbMxzan3KhYZudpaZIekVw+VKWia7DAoFMyZ6mB9eBRRFVunZ9O28paXV4xnNy
w/4UafftW5YcZPnd7uTpiC3QH1X5lzINq8iM24CFCYuZiUBYonSkX+Khp6SopfernmZwQQ2SgXSg
y98dcrn1jw5Ngw1DIfjS3D+0/nYRe2KebjQqWINjPyaJ1w7expIGiIM/oL/ZfX+Fc2YsrS1s9eeQ
R562DqeZTXj+haX9HECM1dYAQVOPvqxCGapyFgwEIUG6Bl+zekquY0Y7TPCZ9l2Lu0aOl/wDj0mS
q6mBTfqAY9DifRv3qLxCP7azSU1iQXFfyVdunOXgJ2Gwwb8JyF2hJdiyj6BHPZ12HSZT5QdfzhuV
rL9eCekJN4b3zovVTEzgWND4JklyS5TNw2YNP+/phqxuPvblXLTYL+0B+gchEjkIKwc6bub7ZCSA
Xq/UL6vEOlvrMxPLhsWEwAJ1Gq1T/SsTvZCL4ONBNi3stu3pG1cU7EGqq25+LMAeCZgcA0csHWSo
FqLgl5Emqaa4CrRMtpGO8L2hopnjY08+boEnNjfQmEXHUjU58lbApBeLHJ9cYFnf03cys0cp0DQy
MHBsAMp+b8JT9CqGkYpVJfttTU1KcgklDdi8E/nypZVZHu2Y78K3GGGkkxGwETnaTEVxzZ3QphP6
UGB4L95fpu09CYCU0WBB3RV8AQUQCTyFlA4oTIV3s+zkinyW88pPkf7g9Wtf/0pRLRurK0IEXY6K
RBJeMhbMmM3zoMZ5diTb8126Sdr9pZkDlbiSljQ/kXbv6gLuZiQsatDePN3ktjN4XwieB6QtReGp
sN3PumHJwvNuxSFHbTtCdVZ/cgS9U5Lx94xtEIoHi5vilY4jo0U7Lh15y/amCWeI7HGpy30XfhjP
zPzGmfeJCb4LeJ4OXRl91+yyunocMOcFBOnYAwdn4QZeEaZ/+w7tEKIMx/sSi6zn4PWT6mnBPIuE
bjFLgYkQrghs5QiZ6/nqHB4ZJxePQUjJGeymfUIfYo3xM/l5zRsP54Z/ilh/E3nqPPiaQ12q8KcI
ybWDh4SAWoALflwCMNVbDLaNYMFh4rWB4VkpUGlI731WiK0tHKu/FXh0cjrUgII52SptKpC1AcKU
05ZrWCh0zDb4lG8gPjVBxt5vZ4vG7tUkElEPUvLjx6PrsQ9/KNZrViW4arYUJtEqOVA1HTIXYA9L
q99ElnGunGlHEkLo39fQ43TGVvJOvu0jCO24DZeZpsdNa98K98z7wKymI43Dyr2P7tnX769sc1Fj
cFqwktTIAPtG0m/nNwx5w2NbD70PbgtVHxTTprTok+RtCpLK1H48M7Fh1rsd1M+GaGlkICsonD9s
R51t/JIqQ6+LYniGxshW8mapPNwohdMLYsCwadz8E3rNpsFTrnkRKMM5CE/bnUdVLZ4+viJD6pZ1
iMLi9nHg4CYKGBoYU5Z9L+agzrEv++RpLN/Tv1D6x9UtELDdIIUuaU1CGReKnGs0B7P684Qb74TW
R+SEorHt03PNMZdEA/8DXwelVT0sMoGIeS6hGHwLp31+sb8hXqBDjpC3P2Mjscgl3h50Q997JSiM
Urs+l2NaShrjPQaxtdSkiLuS3hGkRtKtz0wuNcKgMULLaxDOc+3IKGOk8PnGBdo2iuZC9kCn8PJc
7F77t4bNv7Zzvpwmj4fcecM6wbOf5uWkNTdTSsYR/qzvtynq0xljRiVxnYdWdt/A8oXpDfloXfsS
1nl/R+vO0NoRM1frTVSkl+g+aTHkUgQ1D/eeahHTWPef0CTJTqNhiTbPFnSeME9GBQlnHcDlmHZ9
3oPywLp9Y0tunDQNWDNQT69zrGqhNG+QFKKUPeNkxdKugqtFyo7oXyx8FKvApdvomY2j/B+4lurO
O04/i4cBAXn88fy9IB7H+MGnE99lE+6Jtmr6H4imHWAzAgXs9PCy6AJQfC2C4sOllEmMf5jaCVvB
Bz1pUIhQJSZQPpEPv+HDoj3mTtbiEhGg4i+5MqGKe1Rr4EvJHLvfw6WYOe5g1qsKeqMN36HjTUf9
evuFEJihJ0tK1sdy/bAtomPCKv++xvsJGbZvwRpuFRh+yF7CpS+xdQB9WCP8t0Q0SBK5723R1FOg
teVEY2jVZh8ox/oWdd5UYYdgHTnyfH6i0CxwogyZVuaO+kprzQIsi7bki/Ft4NOO5lJ6X2kBjCF1
hZbPObrWv8ag5qf+YzDGDzsRIWux8Krz2DkNOabcuNzFZJIbEegv10Sf/moQ7SWKowTC+wH9wQ+m
CUvWS0sNE8yGjz2jwzERkxdEsbSs9jZFaOwTc6HBBJJCk8HAwM12V6fIzQ/ISPeMAbakj3CgdhqG
D3aQJYiacyrLsLD/Gucg9znCj8TtksJ5sXNXcv9ytfSYrhWTnbzH5p4Rb+pe731cskNQjQlYlriO
X/l/OhXj4LBXuj3sadNLdCBuHmJCity6Tzx49TCSTM38wRfF+OLcZSTppXOUPdktWaIeh1hWtJFv
qQtfM+67jBN8QjGZnemlmU+qBBGhuJgvHtQzBVTGusMRXUXhaVnv9Uvv7PmVNBwxDztPYrUT2QPY
s6naRdtmH3aldqMh+x3eEsexgTJzaJN0ykNRIYrx72oTwPtsyZBrkJFJ3XUIREGxliXxKB6DAmMx
/pPJfJdJyOQ5e5b2wvC429Zb2r6vWljI0gyPstK/CGxVVeRqxYShGG/xLiK33QZB/ls7RNLJkFcp
rj4q+4R/wqHKekm0SiuoDoDC/lc15DG4I/Ho+qCRh6Q3lJ4UrIM2wkYGu9VYbdWArXPcrbcwgaYN
K6GY2JvEDxWC6oJHC8YOOxztjNMJdt+EiXH1C5O5MAAdGcBmekuyRYdMQOM2XS3P104dN3ZV6ylt
Jd7PL0fCykqIi+93+L/Iatani4cLBCS+irnpIT9g6ik1/XV/YjJXuS3QIu967HR3qlp58vUFeTzd
2/TLew15L1BfQuRvK74fJJh1GOUvpmNKzIOs9VBQ9kFej+9FI1vT6MCywp5joR49icAHVqtti5pN
TiCBzs7ecchHLhhfKTtmPaQtKvBTDZfQhbSrsLlCLeCWMXDLZaHhxQL+UWpniNgKh3dJONiS/IIu
Y9Y7dC1Kv3gMjpTEs9qohui383EBtCSQO9jEJMlshxPApnLICSKmnHPdDQYZeFTJ4byiFwWygcUe
4Ot8orrFbzFvOgwEeAdu7qWECmCN3FjBX5qn44vG+P2Y57d/tG3Fx1D9JAY7O9QAGXzUHcoXnZm1
27Dc6ntHLoD/4LX7p5Bulgp5nrrQaeXJgiXyhTGqMpVLIcrv1qhmikOcfDG3F/s+wjNA3AUzYV+v
hcfU5vL/YErpVMiE8uNF5XXJZfEBzlZd9mFzV1LvsY0Poy72uAubRTjyaTfCm+lZluCw04wcoevv
kn0ODlItDQq+Iq+umR7kdbQNI2B7w3wtfo3uU0wwGt66/8pWfQIt63tQcNy2pXKBIA8gTfPNTqbU
6cUBh/vbcyukmzwYfWzLZrzb5ceaQbbIgNdDG+Z4cLbMXt9PhjXSVJUltzjWGKr59DqN2TrG9sdS
aMQ/IOKKHgFMgSaR8xQqMPkVpB6wG8a0IZ0M//81SCT/+Z/IbkHGDibaxNB2wGXJ4cnh01DbrCQF
O1Ui8Mry9xVNyrw21EU46wUYAWcn9oqEEXbjes62L3c3eiDRpn5YtvQLV7XU1tLaLDLLqTO0/w4R
ighsfgY2NlMiB9Q/mmn3sS4vV6fSStDSA9kKlDKwSi5P9zYR72v2cjKN0pIX1Zlw2ffSzJB8qOi3
oIojRdQTuzvZPg3Vp04MSTa8Ji808yN8V0eKDNhmS1LKZVs1ilyrcwWy2UoSazhhoZjz3/LRp/0F
sdrmwJi+nvQDhcdce8Fh/gvoRNSHdElDmXo6piY/AJBLI/hTlgyzPgHh3fx5+x2Qxv1frVQRQahY
tyg6pdMH6dM6ZJLK9m2CkaKfZHETuiM63wB5sDVXwsX1OqUdrkudaCGouXQVooBpo5sBn8zAXEtr
Xbuwbcoj6zFR/3+1OgFYpIjaPhASM6p4MvYdsen5roxOL1kL2FuXqr/0o3rHpsTrNCiYDWX8P8gD
MaprD5Gz7DcoFV81BX6GyHg/R260PVDn2kMoE+tjZeXhk6A58sYBGnBHVIeaozUFHWPHMUyZwruV
bgbL2clIubC/VLTgQTtFWzS4dW/cnEnSHFCKSkjfK0HBMpE9VzfSUG34Nu6Ne8h+iZEhogrDeKZR
ywZP2sIN3aAnoRKFwliJUTQ3dHYkunfkhfPIJ95gooZlsiNbrqKHitduqs/k01LQnTIgfc7Jr/Vv
bVsKNTpNNDBExrE6Fb+aY75w5tNTo6N/5A+GQFibSlWtAHP2Rnt6Tdd2LZ4snt8ifK43EdY823YN
oGBVS4A1EefKwme5u02ToC1M89QfEzO1lxwuPCTOMFrPWfsgnySSuHAnfd6k46xAJQhSkpOHaRbJ
KeVi7sjQY2Xg5q+GF6L03CnxruJlR6Rd/X0FcJep5Zw/w3aLJGkDUN1t2kBMCXW3+bl7cTNaxgHO
1D8al57NahDca/wPJ7TnsZnFvQ1fDLj/jKIZHKGv9oh2PkstAInixT58FJVBTzapndeP5bt5yx8K
Ym6NxNmHLM7De5B/04lHDdL4bS3cnHKaNahrR53CTz9PJ0k6TRuaml6TEkEcdcoBRAnPxXk9a0jC
59rJyoXILdjo7g9wHK6P4gq/00Bbl07GizDtN9cJvFHz0xQWcHyHP5OMNkI7iwsgy3stkO6cEgDz
5pTdlsRdok3mZyrhfjNjytwfF/lruesFsRnhkyJGteRTpMKSVXLgjk6od/0Vj1tU8XRZeRxQwtN1
mXv90209yb76xB9A0HwVI9NOMJmBytG1AQYAHB2q76g9v0sfijT7vLRIClrhEonVItewc2Cre+nB
2IV1CxOKQUKb1YxWAaYIkX6YVufxtCJjfKnGgU3ux8HSsCfDA5nQR5+dUPfh03eN4dIIHcyFAwL/
FFQiuQFxQBEnsWWFiSb4jw5+KGIadKirF5v89XT/ByNPGNeTFUM/OG2YnSGbmMCxEHma30sCkzFe
mfObbUKc7VX++NeO4djfLgSUZ9EC/U1EDLP36uhl460oI9X4cArl0wQrRjWDnKFK9isghrPrFKYX
nucQZLI69EkZ4RiwaDK7YN6Y2qVCduCaZLZZPCBxxRSOCuMrQ2JPUh9nVXpy/7HjxB7WXcLNtBfG
CoXw4n45cdZ41L+wIHGxNzPqpOOFIFuW/SnxVWtBmsTbzEEadti/T5oSRqhm72fnoQZwbnTeyKC1
cZ9MNcm7P6iS+YcatcLwrDKeM6TV5hTw1suWb4dEbkXIzLNe6vyN3IsITdVbb9SECtO6lCZAqp2A
97cqH040F1VlZUm3FMPl2DBytx12PRNbrAmpqeT/OPr/GAmUIdqHh5qCdORuKJJqDiyQ1X7k8Scp
rBW+rYQMAODZPaJlFlPKH6agrT2XqGx5Ce9sGA4hANDjI8ogy6Ues6sEZyTi9KMbjiVm2fUTNsor
tcMavCFY78O9Sx++qbTHWdI8j5R2UwH2SLFVZ01EIgw/YAeN+3Hje9fa8zRYWiudIn6CftDgkQ/g
Cglklvr6liTJsb0+uePf+6GVMaLgWOpG6JndjT8dmHK/VLmmEpgHCafuTKD4nmdU82KFzWpOVb4w
VW3CH8jNEXPNCL70DaxsV/P6gKn8zF5PSkI1exaKgx4PRwexRe1d+VvGwQDqN7Ee6vnKIuLc1P4b
1j7ZdoXT52gY/jwzqymjLT0CuqMv0UP233yWKbJ+eJcWsnVNp+dkLvFrl5GrcZcA71sDVPKC3Phx
wDkXGPCDbuzwkcVeksZLNF/hQNvhJ7PAJ4CkABXdZ2QxLTEcmMkdorUNwCeUgLCR0L1ANToCmXoR
nrKZyuzCWoZ+vZXWTi+DatER9aVAtGFSRg2aH6obvlfsfCd2G5OZhkaR14hcCwcBIq9+hlf4Npwj
+oGxD2rAVEhVq5ks3O1KIGJT+GXbyvUymvSEBY+o+PI3Fs16T3pjjnWCcxviioyYsLHeTkNSG7kn
8/oGZLYvdIGhr3Y+jUQFLl5jSBeVx0yTVgwICLZ1vBcerlATucz2Xuq4DfRjkPPb1x91QADNNkGd
m1A5JzW2K+GFuAD7pC++0Bgpsfv4ri5w4cCSCvFE3cHoAfL4jxB6uRAJkhmAHPS5uHNwstHq2OI9
UyL9xH50E+M+qURjo7KpspxfvqRsKhcCcemL+pHnzVHdUJh4pA2sskEywOw0mKOlfRc1YofIF7RF
F4DAJWAqVmBXZABHaBpbOCwSdC1mFisPNmgSMmwdTYdY1o++5jvoeXjXpQJiCEzd9bSzsO2DI920
BlYxRJOPnh1F438VvKm61D9IySyalAiCLTxIO1ig2jxcT8ENmeUWQyOULUpSTKpO9KY9b/fyqnGh
GayGNpWHpC3pC2e+V0HP67dMm5REiBQ59McaaomRuTxoEns+xECxbOZa9fEohuxqZsKTxFXUxgOm
i4OwiLExofGwMgJ4pgu8jC4ZswnDjRINPJLA4M271aaMxs+Jh3itsUC/+A+rlqu/WkHljHgK/b6O
oHEXhRW+jbitRExDSot09oefOmh2K6GbUxH2hYEhea1iRC3/bfnb8YXcJ4G4BasO0+oIqSGJC/2w
2RMHbIr8pJwO0V6MVFdSvpQnGkc5Y+xcYW9mQhf3tCLAhFJ6svSu03sy5+Mfz7vf5G1se3zhmlmz
hwVEqym1iAjiQhFFKivc+kQQ6XP/MZu1TJok/kqEqYdZ4/zLsQXjZSG1Kp4v+OGojrhRKgV57gQS
eVaOUZW3KKDNMullNzv/vBsgYQMXWVyqEw1NixLnO/Vi+FSCvDy87eag8f2Jwfvh5osodf3Ycggk
ja4/ySHy3RyVFwxJB8j4s9jTDKzs8j+UlVfyOYFCK7ESqOOoBo3e/IfMx2VA+8bG0vPz0N/0APnt
k26Ja3lxOcKRu2q3T0k9KopkkCGtfUhxuhGUBe+Z0k02sfaxVkarm4JY8pq6Gc3Jfdyi0xdusqIs
fuk03HoZx9r4fH70Mj08vaI2dqVB8V5bz6MxHFysoOvwYUn/QKa0CFFx4zN4I6n3k3rsojY4QINR
ZKw49qrXR2NOPjxl3VhsNv0/Dc2KCOLJ86ljQDpwMd85+XlNiRx1zKmUVk0XmitmDKgKSuTKgFsx
U9RhZCIBXJfXZGV4SGMOgEzRC8QTUTKtntbxLVU+FygQGrkXgqc+/YYznteZtacQbeRpkOmCSFZN
y11V7NDc86STLp+XXD4gL/RVAEZ1mm5/qm3TSaOH8QE3rwPRhc1J2dOuUgCCwCwuvq6NDYeJyVtt
TmqVunKFN3rPjC3vpkkv75WtOOJJKeLm0dJkVuUZSDSKN52xpDgKEX4sEAEQeuYlVatoUtCmOm2d
skANsuWScB02ZGixLHMsE0Vx3600HUgqhvT34Oo8UkvdQb4JFU/sx/JFGh1LLZgF4fq49mLCV4/C
T8Dl5010NovR84Q5AVs4F5XlAifuxD6cQjQml9NYamvfiSybR9EoYxE+YtYznXC18zH7r7famK1z
V9Uuu3VS/2lT6lRgSsYxtdTqtLIPBeYyQKLuPHirRSVX4qN/INke/MecIc9sW+KYcrzssCa8D77r
eEZZm1vdsT6DEUbuEQ7GuD8q3xIBstg30AIVrVEk45uzg8A/fvrWW0efqKBqEScKq1+nfA76QtTa
O7+YnpzNo32avmi8tqHuLIYA/2+gWXjZAW/W/vNvoF4gX1PNCNESBFqGJX+74t6WB8KA9LOAGub/
CuZTpJQbA5aILg9Wy48sg3QJtY1wTP4swIrfRKzgj75+uKhCr+BK9A8I8nbHsOp7QBO5udgpntmF
7heabwIvO/ogmKQdsZfJ9Ra2Z4CmZGfUaki87q3yHqHL0HgNLoWACVaFwYO+yuBHbP1Zk1vBHb96
6dMfU0JY6He+AP9s/de7iifz+lmH9xga2ADanF8blu/ZqXLpMg7T7p4ep/9EYwl9cFvELDDJbcI1
SDpNQbvZQXezbHxWOJalLE8A96EUL64nPAXNJZ7dc+JdfESsd2tkllnsrXsLwChU7xDmOj5lGcLm
GhLucITYBk0TYQrCPqdSfjabfzWKeJp9hhwTcrpcczKl4CWJoXGFRvalKEg+HWivnF8wWkRdTYZq
+O5XKVK9/fYipBptJ3MfkTw+XhFCgyXaUeHibu7X9Es58IaCNoKdji8uBhr9PPDfw2vKIoobH/rx
pKdiB9SYd8IfTSr6c/eoHvMPtz+hdzNf9DTg/f7iQSgtB8XMdtRSB0Ml4Pss+Zq2nndagM9asnw2
U0MgEAt5H0o6PK15eKaoPf5VT/j2PE9medbrxE5rTiQ3stXRp05/BI5dDPUDE4QrPz5dJuHfXIrJ
Kos+mKjesmTdfOx5WfzU6eGS9T4L/fm1we9let9dR+jhUR2zfDtsGCWNyqxO/JDisOKOa7Lwi72j
jy7/4mQAfkgO94DGotMdsNz8oBjxnF9Mn07tinYlwa7VV3KD9t5nKoYOLLDg64msUEUWOxFdO6wy
6gIKlI93sBXVpklrL+oIJxBAfZDoQO3VPnWf3sQOVeMRMbIqRjAzCrBXR8ExIxo3676dolchK1Xp
56rZjwa/jMxCm0VxOBcOOL919aG+48JfDd2LbqeIkVJAitMKRKRjAO91MJRckcAyIh2QHjK1kAvW
foYfLcQIgsEX2ZkhxMEhSFHUuGaIATTVTI4vVha9EuOG/K+dI+FztOFUcL8dE7CrWCHOJochignK
zfX6hPrkHRPT5V2uhFRM3o01GIr9c1TlXf4iQO0A3GsTTjqBWyEQRQHGitSz0UklSc8G7CYUXDjs
A50Q4x3nLy81CR/RuTjXxek9ka0QvvwkDpMccHyZizzHRQxi+c+62XTRiui8vgZFunzL4MDtkliO
MFetbQGNR5zTo0RGGB6BuxiKBOVOY+W/rbP2VVIkDmF1hpSW8UxqwRCwzqEQImSjr+W5DJGCCYEP
yvAU+E+emIVZa7we80SnSsHhiz6vH3/0U6KWCf6HXhKsyM4IoyKTSvhwP2N0BQRP57JPMJd6P8vV
qmbgPyKWHLGu3c7XyYiZq4FvfaJlkzep6ZToOPi9ga7+/lEORh+91seASkk+QabupvFOM3EgWf51
4muX4gn8khlGVr44vkfWKcKGuqEZTuWbOzB3OS5KA44EZ91bc0qhpBEBa/xPqRH/XmFeQK93ZGvO
LYOzV/5eqwBKo76ktXm2vCB3NCoyH//o6bKbrXSdWSBF9jT00GrTwz0e9cwrmwtI04QfKTVhrAWY
sUCuyt1uvtOxSJKvZmS+XiwKI/7AUfQ42xJCU162xgiOWVmtRxz6VurLv0MYbFNlDHvwHtjt9jN9
RfSm4FzqOi5FnxXKuLAnSl2vlWhcbfsS6HJTYmmkXLsESThyNfzcoTKmrdJ73am/g9LBnkUgLqsV
ebJfWYGqdTttGNU02+lj9S5L3wTNDZ0GTV/AHKOrIWCq5wmEZhyd53VTbFy5e/0y+Xka2i8OIagc
OMfVI+31CmYZB1dtMF8lbBuXkOPyeUo/m+kZR7FPM71K06bMCzYw81XMFzRwHsyw/M0GUc0eWTh4
HE4rtPL1dxb2mF5C0zizxlh2G7nOnCeIBVb5cAQtifqoiQpuR15lsj4ex4eTyDGwZTjhMJRjK88y
rkL1wecUkOoy3Kog5FyN749wnmngTMP+ude5rnmwrA1xCTkQ3f1JXSLlAjzALVrqlpIP/IaRJ1Qr
Y4IhgXq1l8CrqeFMhS48BPdeAUP4uOqYpn8g9lVOe9DjIM2cNx9iiVDj43QyLNoU425zc14tLU7h
Uza+Mjwso4dt9HLWVmYzHHpuS3F/8MZqbdL2Sr3m1FlMW8z9T9xA1QhI3J6cTkwUylEkiDdeZYon
l8KwkGEwXwqM92QZSlkuczt+qSMyOmqklc0SvB+/dHB58W7A2VhVgXDuWvnXXg8NlTKmengwuKMf
X1TuIYBI4LyfwKWmIa3imGBtxCccwhfmE415XEz+1DVx/sqhaddOxW6l7pKM1SqbHWHD299ivmyX
x6aim5IsNltPjGLgn5YoxMJFpuxy2nf092H8f691Q7aGGLummz9ey3a3uCO4gC0FvCJEqjBL9xBr
Sl1DK2AlI6B9yptn9vJn0kMgXw82c3JxOHkCcbsnr8k4Mwsf0Ux3tfwKrTqWJIAsluz8qes75+kG
M93OEAkA6yIbhZYl0+aOsWDd52f2Dk4DqQZOvAtUVZkoHg3/224sng69fPW9atkCTStsK8GG62XU
R8nZ+W7b+YeUPq94ZTO2jTEgvMtvuiFZsAkPWcsEJz0gO8pjVVKuZJQ1StyMZCK/JQWSNGsY+4gg
ueCuvMa5cQAq/HUEeFvZsUCGxRlmEXk7FuIlnIoR05gXbjNhP1SkbwBk0TfihnL1+ZGZIq+81pV8
NzH2sDDyzooWpcyURHefMbSvT8YH5Jvf57oFis5TGyDY182p6ufHt98zLRAkib5uqmopUKEiD39O
xMsH0C/VyJCLQMVreHx5CXNINfrujkx5hW/utoPgvd5ywYaB68frLUgOU3px9f46So+xjH76qvff
EaidHBMIwJH7t82MzuRcSUH1zMT51AAxzphu46JTz1MdfI4RIqDgoW7VU/O40Rx0N9oApznXoaMm
b/RlMjCYV4ys7Irb7cFZj0ztCcALizWzQY4+3SW7tL6fyH3DKIvcbPP70CrD4mttpkNwnJ1hMYHT
2hE9Fuv8PjaF8q/8sDOmrrGPP5zAOdammE3XS8JdtxzNVKJX9z8TNRsdc3S1kRgbQaWx9QGrF/UD
y2qWT3ziM40X7MR+4OZF/DQK7qYYydOnzhOIwJo3crhfHaeF6rTUj2EJX0DHsGMYPSauzew0mpMv
3yPmDax4WlzJXPp9XCZ3CxzOJZy+EfcJOnnFLGUICbsjpMkoxvis59yNb58jNSaoeLWLliYvb4dr
mIA2ESkzDdNOrbYHnZlC1gWNqFKKFS/adCDsQvLA3WivxbS8K0cOl0v1FfE85W2zaJCzIOODNliF
zDyjlQlAxeb0kNPpIRfouPymOPRvE4Q9iMExFmO/iB2f9WH7lFtQE/rqfzFTE+4lZSdxkTC+re3b
yMZelYR89uaudVu6z4jpALy+F0TiIIfNqmwqUfTIFmHwDWuq8tIQ7k5W/5bRKuwdeknIYgBDYUHn
VtnOLdkbIA98k5ZUlNhc9lir0y2307kUKwUXTHmORCOmrZ3w959J4seSB2Ieu5hHSQ/au+9uk7I0
xEPCH1+VonKU2kUoP953mIi39Hcrpf/dKRH66Z645EXzilIQk8K2RQXw9wU3Iba46zRkhzozjdGZ
0jc9m6f5k6UQaU7t0EFgDbrtGPXA2aBBYVU3pKM7ZoWHp2aPbjeYWvt6I29UHczppEUpnn2pnV/h
0Q543pkuNt+/+KS0QM797c9xumcdI6TpcI37X+kE4+X+UuLlmqjH37ni1NN+0BYXGW6KfKrJf4W8
kqLjCnhK8VBidaQcHD6DZRkOCctuv2tDsmpYdIKMCeIxbHtSuA4Zilv9/Xga5Oh/1w7s4nvTsug+
0Ej2OZnnO7lmoS5LYaUoVlPOwi7gpHOXszUviKRPLvaVIH7eIUM885dIxdYm8LJEh4kUa9ZJ2tjm
Kt2GF08Qq8wLcR6Ifwy2VZjZDgpxIqPllmukPyZYlv66Tb1uLTnNs/NxCYGbtUpxzH5+LRZ1OSuL
VCAJ7OUOVl4Zt1vEk8HU21KCqIxeD9ls4ShBvbYGtOmjqRBFMU42fSp2PkBOuP/RDabgi/+2t8He
kLRnZnvUroeBJxc1Nzu9KiEAgTx56Ptmb3ZK5Aa72F2RFLdyIfbQrxNu4+OhHNQPIn5GF2/oc4Kc
OuN0TRIecB35X97CmyK6CckQHiWibcRSGiQlqVAuGjt82f/oql72T1Cu/FxcbzHHAOCl6OEI4b7v
ub72VJzZNKUzak0lBH90+9j/OjxrpLkv4UQ7HLpi3iBkanV2SSfXvYSTVcbu9sC6kLlmST6502/R
41AVUt+kxSLyjB+FFGqgNNadvsE9zmt5pWj+t+ckIQbfUHmhFRqNesisCqofiHZ3QgO6nKO87G9V
imShkG1Q4nCtzeClI/A+TKAbXmwfkg9+13ovE5qGZ90eE7CYW/Lehch0QqVcNos4sBdmAoKUlt+x
xDfgO4EIeJwujvfbEf7lnGp1OCTAUAWuPE6AI5/klJLOKkqvT4JYCjXV0CamWLdrmEzccSQhZid0
RXTS5AhpVATQqgHAy8DQlw1xc0whWvP0DFmY8DzUsYys3c9xTz7Ym1w80sLFQJ8P7sjTFYXBpE55
HHzjBr0d7EvJCoXaPiIlPGCsJf3+T3tYVy59BPb5R08BuJB7BleiZnv9v7H9EkVUTWjuKY6ED+qq
Xpo3u0Cx9Cpb85zKDpxEQCyRu6TXPq43igD/aTgj1txPqOpK4cGCY6xG/TrJs2wMyc9V7inBielc
jQJMvS/ZSStdO0oM5wOILCJ+kgVuId+9ffPH0v7aw8Iyt5xKCM/kyfL4D0ZaZ8MVXMT/R2jhXosB
gvbLvao2Kr+h/z0+dEhCsDddvEox6bU24jK6He6cF2zL3P5evvnyt0J5BGKi/OChcwuG0pSF7X3h
QmPmoyrgcqs5vUG6eDGVD/imzrGP1T+vvEUCvtwJEuxLdOXM9bAPpaUXVUOiwH0Uz9WXJTrYXjck
wwrBwV96dMzO5IU+ftFEDIBdgrkjvvs9MvF+93emPJTMs4CDigLQBESAlUdAltp4fEgx5moUjfba
JaUgNMPZ5yivaV5hRwFsAqOLzcAnD96yCNYzA9NXXpgOrdsbma3GN51DnXjDI7bO23wW7nj4C87y
y0DSCnUVsMZJaQtyQfZf3mZJ+ml6eBh4cyRbVoavTVbUCpiFOA9DrCmGZQaxYUHeceEdlLvugPp4
EbWeIHnp7GufC/HSFhev4aOF6tKY8i2StPZlpOLvvtfXM8+E6k1obKRNrEp++u1dWFibB+YI1Foo
x/KyPt5VxwqoPn3IEjuPtJlTJ2dholV0pmC0vHVUR0Uvi6Uo+7+yEUOHaixeEHY9jWLFEmXeLmbN
o9JqgknvyIa7EbyNM+rVqzKzmbW7S+14jkXoHvT6CVQVCHQf4YWRbhCOU4uVfCNa83LTFwFfBnF1
yaGW/mXAzbT9lNuN/vVVlUKLUYbu231jjEeekngTkE17/5d62hWwc1Gb5dcAjb10IXD1t3GMDRIw
op2eOkVgkM6KlRHLfCCEWAeX6XK44hUgx1z8UHXb46DvgQ0ozB+0Y9H+zM9q1ye86VI9Zej4Dd0A
xRfv9J+6Y+tEofUYoUsbwGAByYTsETXci+exjAJLL/i/6ybwJNMx15Rt0C+xppB78dMB6dNetdCn
dpxQbeNU5P/iigJq4WVpIji3Pha1tbNhWmRoaOH1ISMkBHOG6ltPTFQIOcJ6i+IGh+yzCAUfLwc6
rFhkzMmpIiw2Q5kWbxiZTllZQFhJw4TNfyHICpp56Hjkadg+HLfq37OQmVns57omp3+DiXyKLZHS
0WAey/9uxByvJ1ZC5uY+lwg4PTd9rfuUDrK95dMTkzqsbr3E7sFBYU4KzhQb/Xc0h4p9WBcWP2vA
VPmEcV4L8ADdyMRWQFJzeH6DsJcya6Kn4LzPCKIx9uHJJWeBTqjHb4109b6pW9g2Lxxms51x5pbB
Z7RRxzHPfaKteM7NiPINVsHsJwzFJr4R4QUXzPP7E4bNWzul6tF8/xSVCbD6mqPPahxv+G4TXCAJ
zvNP0Np+MSiY+s0rQwqhdvIeX+dsHG7QjUsfXkfBGPjS+ULBv+W6FT2p2ZDMsxGyrXZrANqeGO+r
GG/FPAMNzXQrXJJ4VpufiZ67tp4Ci+mR5/CzSi+SGMkW8rixTL62ASu/F9yUMBacDLxoyskOvT3U
8dehQlGX/87mHH/icPDGHlYPOnmei6Na+BSy5TqVkp6WEPpltXF++Cw+x6Ngy+O7PGnuVbKKa/f9
bkvu3jvFoNii6989H9LMTla5V9Lqj8Xf7qiYCcOfAFjaD30/CRCEggCIdnBSo3YoKsTEJrn3PQYG
3DqNmYzty/vR+BuyCFjJdZ7/y+y1TGo5Ughnk1JLp3rIJRkoC7jnCNhLb2GYs+yZz4dv1tYeGSf+
pHmm9dG++bT1OdCztI/Z+oy33DeGncWacI1dxiWJ5cRL9zM1MKlOK8ZGS9I87XrTSW5IIHfidPDC
Qa7QW9HxWQAvukCBHY+/9uC0uHJEbquHZxn1pr0sLi97pRuBzdpjOfgBIlhBnmmIdOVbW4onhFDe
06P+R0gSVvlj2AZIqfKUQalhUpmhRokY0kBPAABlqN16xtbTQJHIYKpwefQVn59/JP9RRWEGhgOg
xEaN2hDaSJH6SpECncghlxSrYu5AwXo0fOWvYoMhTl+WhCGZj5xbwnSm3LK5o6eCmozzLhXs0zhA
mq29EylBPIljLkLD8lFJESUgd9TSmcyv7xhGPLtAB5RCpn3NDmT/OqjSPdJvoFGYeDxtovP8JZy3
FDMu7MT7ZYOWulwfEHKIILh9vuVLyDuTn5YM6iWsHazWOjfst0R+Nae6SYzKfz/FQemjDSsL6H/p
4m5EBa4o3fXLrEDrKWoh4BXNsLMK/FU+BwXw/RW0cyWz0i3j6TmXGv3tQIc7qaiL/FOxW3cEQH8L
gHbHFzmflr8xY4RYjgO9Skb+2D2NYk+jkO8mvp8j3yQQ1DyXUkqHXLPjUFe0SclX3DtPoKF8PZL0
YLlQOh2zOP1OTsDKQSGy49mzdelKqBeZ89/59etNkU+66OMCCjG6FjG/NQc4uq5kYZX/3mcpf9aF
4rQ7hawj6cMl+7MPsyJr1+ogjypDThvotEYbm/OW0UDRB0HzIUEeFOqTS7c+S7v5DFhsKMPgfTKV
kqsS9+NKJerXG36JsWzeXbOuFloijLgz9RvI4yeTfyVxx04WfQvW5Kir6hvi+arYNEazm0YypoSo
xiJbh9j6YcQaQTxVIg50bZ4W0AAJpsabVvAWKEN/z22XMezJPYxo6HB7J/PYfjYjMvhR48hliW0g
uezLPlFPAMK0dmJBMUsf3q247PO2Vrpuh9AqbH1ETofcV0UJqtWYS/09qDObaT8zK5w6nre32cgS
FKd16DRlQg3lwCl/vTRALhpV4JKXF8tfnx0xlmxznJRjaQAoRKAxYdpXmx5Kn9iHdkmqy8PfR0Nc
iXUipDz6HSmIpYAqL8KPDi5u6oWNZmMm+aWraQ0z/WZZhoLFso6VPjHJZJdc18j6gZOpAxKleEdt
M+NTqa1sI2lgrMjqcWKj2Cq7kfFtjROfT1ugzEDlBjzzR/IBx77zgQyCEfMbpNkXP6JeoxtY42yH
UNNhMreboKSXuEsfflvl+mbX21KO8nYRCidRLF6BF1lGolfnk4eMrHyUy2AfBkX7FKECU82mN73R
jjlCcbalKAWKAFtJRhlqEpOVoS+OQMcjWROKbnOWwz+ZOk7Z+yO4YPDgp5LQlQNxr+hNcgJoXpYN
q6pJPZvjhkwTqfzCMTS3wM+jgI+ALco0SbuYGb7Yu/DoNIAyN31o24FY1cYMRvePliUi/ZG9DtM7
uPs2UQCMGH5fNIYtx1QEPirGyjVHbb93JYhQeNHs7WEOGWsWfzTSeifQyt+dDx6IzS1CYCaQclfY
tkLXb1FROPS+BLmWqTxPboSec8NyrAQpagJmW53/QGnFHHOgwT3/yYdz+r00HvCLMMavi9V4PjKU
OxxKDDmgFXS+xM4KhPsbxgcznPEuNKHJTs0vlWThB5GKXlYaD+WEMyXtVNJJGboepZLn0KVLP+dm
RU7fBDA8mgu+XfXfy/hYlKkMx2BrGKwy7TrEusKPl6ek813a3kbWR3k6Ysp9R9WqPe2kG38tzdnX
NzFyTd7kdtjGzlIimX7+RmzC9e6oed/3eIX3jmgg0Ii/uS8RVv44WB16MM2c8nv4lyDx28vWfmU/
Q4+8sMO7juPzli/ZGh/QQA3kzzJ3lgeZwSobLZn9C66VdNnKdgGuaVh2QvUKJ63Quv3kQkzgR0Or
l1U5UfbhtfcbM6UNZ1Br4lXr6dTNLMXcYTsFwzugnhVhXMDWRRqWrMWLKpGHewxqG0rTuRS7JuNB
wahI/sizoaFwVMjxLOlpMl7Mm6RQou8fAYzlB7AwEWdgH8vzscclKzWePAwMKS8tSragiUP4ftnq
mQj5OVI9vvvCxbrSF3uKdYjbZx9EsOl1sF0wkJ318Ps6mcRiGQdeweZ0fUrVcgb6WLaz4l42tv9Y
CQj+gGZX+tLS8ZknTeAX7c79w2TgfdSovVwAqEtgY0GiZWK+PjmWb5idMIbZYeGOid9R4vmHzx9K
RHfkV4jWNC1cTHfTG/iHKYkcgdPrV0jcvHuYMcGGW87VfduOwy14NV8hL3L1VnJRrY8g2gTo126Y
tDfv9lbmOoyweDJ44tlv3vjj+lTmiS1oC84cABZ48M3T3MQiAoiaZ2qjKA5iwDA1bkhcjxLSV4Qa
H2Yuu+YdYwiCdJ8oHbrQ9gE+PFNKye4nj6v1iNP6k5u4SK9mgymEBd7f83YIZ5+OXde7seNVHe15
EW8jsWANCm0gCK195yboifnivoaIWux9Lc6+XMgKlccI6VLDfT/mLH5QEj/zjtMk1ONxixOTdjTD
Q9ffJOvP37yE0d9INLQLdpTucpYkYQRPaq0ZDzFlA8PvzxYs4KlDQ/xLx0bEVF3LSrpbiLGnWDbf
xmtSOLuKq8sP4s1HQNQRvSPA+TAHJDCpSPxRcLUQOpz5nNrhVPjNP+i6+EtEG2zlhUngJaO5JUzK
Jrf7Oz9fXZbrXC3mzF2ewvzb58lfs9xNjSh4c6Xbh6hEwh13JhCO32v9KOyW/ms5Q9/zJiwMpUBM
YjcYLIDeTLSKYZyv4kyzFewC0ErMMvlMzHj8Q5zskAWETKsCHWt0RifHOOUAHqlt7ErtsZtKl2qJ
v3SlhCP1n5arwshvQhQx1lQrUNPiWlkxXfByxWZv2IaZuXzk25Yb8VgeRDKUhDoc9ijKsHSRKkQ2
RhfO53fBBkY1SLlBOEfGaXwo4ZCdkXmcCIFBl940R9onnuN4+8zJpTUk2M1bCjHZosa4pXiBsuB7
tATUg5+1KSbV7d+BgiXHGkoYmAB9ddeRzScvg/yWbZq2vKXgW2S0lyZSv2mCkF6vXWf5u7jJDG7T
exmmdztyXdL/UBR2DVTYSSNZSaGQ7igVPxq2nXHozWy3PJDSdOpNAjrpHYxa/N3Ssk9vtOr1yH6K
8lmiV/2hrkBqjFx1xEiS+YhayYCCkmEzG2KBoTdJFA13ZxDKai6yMFYEtTpFRzvQqo+wRBUHFoiH
z/YzCw486KSzuH3FS8vpcrudV1Hf5lGNC3IsZmL7pEIvSH47N4YWIMEY04lKr4I/t5xPeho7PuLg
2VGNOrep/wVvXC/tjEN6QIOrH7JhGGLNGaYAnjvGlw2sN+zmxibZe/ahQRHZZRZq8Pnlg8Sdn5bS
0qJTRhzS9S+dCMB/blWFnJBv/LTFU2bekdtJPgReURtoqrNy+TNtkoEBsY9RC9yNDawwy/o9VYSU
i14AROZ9imIf/ORvAIgNmxRlHIhyvnMOhBnrIRzzIkEExX/8B2YEke1pTRPVLxlNDLFH0oy5VwEN
/TZvHjMfyd8N/BSHaBqdnCq1yuHLoJ+9FguRnhNyOOW0iFlztCS55nJXNOMLmNyFYG6siNrT3Oqz
z7W5yjrUUCxU/6WprLysUMLaMTxPsbFfp8TiGxz8KAhj3/XGO32far5ebe5+gFmIDQnWkqZZ8k+w
qjSA9cNjTfPIoNjTnemlezh6yDX8IjYSCaLUasB994XSmgvuwQ0wi2wKVhFdrQ9D7s44iHCaGw27
DbYgirAu+doXbDrx01tFnOjrq2btA91mBkhFeR16z/eAfTWsnzrXZ7zLuQ22BNukhHG7tn7iuhiO
a5KQcbEANSrpc6hiyaYr1cOkPj6C3DpyMWqlJRBP16OGqmKwHadrBRtamF0HXH60G+thZHl51Ce1
Vcuv//Fh1m1aua5bJj6PYXxMlMJpaFJ8JUce+DLBmoVycQTDJoVUDu5S77rFrEKkwACH1hRekgI1
vMgdPBAlBKWC91tFX7pvD6hTDE+u6Wt/ubW2/M2rHhO6c1ByD7LTAHHFJ5ylz+b6Tj8rEegcCDQZ
rq+GaKcQqZFZumg84l8e3ckPmJmeOAEH5QQBgzF4TGbZpwmc9NWrVsUwUUWPXjkmuq++YZj6BGLu
PftFvdiVF4JNgiDkzP9DdJd1AlP40t8SAH80xWKABPmpJNj4699owVLwW830ZHJL1nuxtVchMg/O
Kxx3cf2WhYv3spUxt+jwukCDLjkwXicuZ24vk6qXkhNoePVFlL71ZdyOZCNxpe/tdCQQ3hwwA89d
IgVxQUsBzcNDNTk382THF6l7UdUupNfK5+k/NEHzau4OGMh07exvC2UCX1nRFtgegoSMYxjC4JY4
XDeOIDgX/KaHXZ3j/Y3G/rPkCzDUMMq769kK84sFoKzvEh2t0U9dgOyiLsEpo7OuLh2rDpggRCTM
DyzBzxj5EOoVwR67l1sDDXitfVNG4S+ZGep0EtcqYTsW8Wv2beigqXA2jwVVcZX9Cwwu/tKq97av
+iy6ry057cN81+EJXr8EuUhfQHbBelq09GSaQdKWifBD0orFtKhZvm3YzKUmS8KPUNJJ7sn3gW2r
bS9wIdWY8KwiUfteuRf1zfyOYTebvKHZjuzlzpx+KaXZEJ2kVAhaY75URn6y+CQG+HRg1IE7+o76
6tim/dl/VORoodJF7r12Hdfy/EnesfeMZ2TeqouYQpxm6e1fvwN953b0/mubnhX6lYujEfiTRaDv
7fD65+GH9v5HLAceCWZZqEJwgmBiInE/Vo99tt5yW2glxvKAgROwd0Aq+KYMZ/89EgI+EHSF2sZO
9i2AaRTNcNCkJQibWQWUKJqElOXIWOX1rR98v8Hgqo0k5hjyuaehAZS3klc8A7+dPUfSI6iIGPpw
GhE8ioyO3N2EjoCEV0HoajYSGdWfrrTAPWt/VZ32hiUAszWg0cQJZzeZNW611NXyuz/uECYKigud
yn7P2tjh7SqmcudOMpJo/qKJaY0lVEbwoyzmMt71CDyRo5ZDDHXDOBnP18uK/g9BhedP7xmyE49s
YHWtrcwDB8k0IZ93qx6C+TcbzlFccA+5QD8S4nzBAP28efrBVRj45sOBYDLzaOso3ltYetb17+Gn
RtyO9MNeD8p1miDpSzV6+8rpVEXFuvoxblpfRRoWhe4ARuAOpn8XvPchOOnpKqK4XcYh2RA/G0iV
goIfry1GD9cZfqXf3GaMq+nayjLYrPmDegsiOakY7899aZZsTUzn5qMpfsPgW+YW7tFAiMYKc/UX
bJY3k1ON4ZZfgrtWl5/fQC/TvQsBi/Am+nlwCDqZnsSmWk5Dc1XuCuBSLbUROJIjheSzr1dkjWaj
Njt13Kg/Co9Wsl95a6e0P85AqHsXxszNVPdNzbXwTjbrDjdjrDcyDj+3mvhhRou8xAmfj5NQDV6X
fDDf+re+NwD03GWMYYs6OsDty4940KHlbpqfRY+cr0zeX2ZLSN6JjLZhAQAR0JfS+ReJrUvmBdSl
5GXij9f9Ig/2AaNDm5pgjJpz2lHddkft64nF00tzdO/HwLAYmihb4DhgtmQZXnfKvBfcZ/QYhAPP
jNrmt0eZk5cDlNwFIVuaEGUjHBy32L9NrBRZKTKavR1IetTASoPqs4pKESL2SWim7sSpmrF9OHc6
D0VWvnxt59NMqnMK5n2babq+M+0LA2sSDpHSRmuRG6gESEnrh1blslXr7hoWGP15YWcIl2gwBEsr
C/2C2D0XCWRT53IbRhWXxuSl0HEAtelAyCEPlxIxXQbsjAE/abnD9+R5O6aXEa7b/d0iNnYy05u+
YUCAGOsaNcktLLd5caN7YscT4sVNEpEFIDqsEa/cDdSwxu4inmg8V3H4FZFxxR23RwClFSETieoI
TNHIGAOWSS9Z2uQCQW41kbyi8t7d06jA39v5j8eIQuFv969jMxew0ZTgpYTM9Akz1zAbSCZ6ipmf
nuXOszEqLU6PudcUqUMRBJMzCjxQUDvZXuGnLgHZ1jpn/lprCJJQmV4jLX2AI1gR7w8Cafhs+4Mb
rbUjtNiEVRO8lYZxfPJsUY4jq3SP8g66Etk1lEqBVEgLiOlu05Y/p4LH9CyNKo5QwOMca5xcQV1J
Mj6TmoOEwwunl7Rae8xKxsl0EpAXSCWzXTYcCYdxsCSFIQKSG2ECvfPO+nqtJYm5ar9AKFYBRrx1
xcavY8xMdYQI9jA4vA7aiFQervARBPrI6n5gj4tDeSdYi50MpAVotCXMbQztwjhFzndnYrrVsmy0
F0d58BgQOb4YmMMozjR7DCAXfl61oBUlYxAic9TcID1OBjzs4vMj4W0KcOX1sTMkdGuOEFoVQ6IY
Jm1LQHfCQO55vujUJ4P9BElCgRRuacDq0x2tFNuMtWj9wLQmxIGJxRD+fT5jyCceC3//PR+Dtk4Z
/qWwXI+m0LyqDTjdSrIj3fLN4k9RA00wRPVwCvO9NWmvoh7pjRhNT4+ScvgK5HvWxoUNjANHmRy0
THva7VJb3Lspxvak7Yrk+7BIKwa0+YBiyf3RmzdlL5NpoNJKqauv3HSu8IKWJq1cRdHVjp6tXS5s
u1YqqWL8UgJNeLgGyc2GJvsDkxzHDSJ/fW8iUzLGmAmFMY5h5+U2dBDfKby2p8CJ9jmmQ9gYY6ss
cLMpbhLXiq8RLhN95IX4lOnYfV2t11JZw+ePAjMIEZMPCR7GEVUv3g+rS2k4WgGNWDJl8kYnLVXC
DRymOhm3nlqYW2rnL6Hvg19c2AaBh2/M4cfFaPVcjojQ7ef9LIybN13/iZCA08Rt1d2X8BaZfL+h
q4cJeNTPSycTTWQsnnLdGORQ7m10QHhqTSnwk1F0Vt8bO+zM2wL1RPULA4ISA/SdtWnPc51RLsRI
t72lQ3sSpcomz/G5PaoV1RIypEPkqOinsBCnP95Q/PZdUAkPEGL5NA8oB2hJD5wn7Y8fRKN/HpFW
n6FNScJh+E89Wr0dvUjHyl9r9iuu3S1CDqXGKjH9mB0QMt9+myjfhpCKyxGgxhCcxAQiEmP6OgmY
hxOlAITa+V11z5Q15OtyqtFnibTdBxZ/2I8tDX5/6MEf/EiaNLb9a/bIbKqBELSH9f/Qv1tqYKWg
Ny8PPuu8Qx5XIot1eFOyT2HyKm6UB+Ab81KmX4Q4tNpWDYUhy1Ej0QMG370iXWlZJ6koSrdXnAS2
38KQvdI6hqg2hFy5sCCyZz7scy6EfJr/5eiWTPtYgQEYo7j3uiBbNb/PxdunM38/hGX5ep6VB5Ms
EigUeUZDyGDGlF4LPTZj7jdodMqtVk5rzguamR28VWCXecQVoULygyWFNTf+loihTdf91rK4dY6Z
ZvBfdQWubiVjAi8OyhM03ZhNlYXh37Iarr14/XNqCVDwouTMCrGDEuZTElyFp9O3a/QT5yUppRjq
bYxZ5d1nSOadZl3q2IX2p4ZaVjf5W+LKKotUGfYEynh9MNJGg5sXAQARdmD9iUjyg7jmxcJ+6hIe
FDYocHzQSEzh7oSh3LcPWNdw5JwlSz+YuPmtf1mXnOLDpZvSAJNqa+Yv1pgM0SyIX1Gusll2AqQz
vGdRVEsDt3vLPKArd3fylkAu9f3FdLcxV21d8E+v2igjBqPXyRie7H39IcaYLz5+npyYMIU08e39
SlGxS6pFnHfA+iXTf01Zxzdh72Iw+eLSRDoY0M4w9oe0lbLUcrWn0WAMECMgywIwBz3mxjSSEfbP
G8BFhcqpxg/pIq+ZD//Ctcor46+2e6fXiveGdnlw+Mi6tWv2Qf4RZn1Q15lwYN7rA8Fi8SPCAkGz
l7K/hklEyC4AWZvSUQ8WxWOYZ98NFeoLR+bGbGeLf+I55q9ZH7rGE2qF4xeE49M4y/SCG2Yw5MrQ
szuC88X6eMrJzfGOpEe2fzyURk/qBzN3eFUO2U7L76rbNDmakut4UAG13fYkb4LhqmQaMWhct+W9
CeJG0f8El/anoCZp5y2xk9i2ZkVNDVzgusdMsp6nCldUB47QfDVsbtnVxJYWmt5TX/5CbZ5JLsEK
qwow5o2UAMM7T78GN0ybKA8xbYFNmLTEFuMyGkaJRIPrj5O1LstdcRGLOlgquFt1MsEgJCuAqaw6
SrEyDb2/RzhZrbvWNlhq2WeliWljv9U1wMwIXvPdALalJjAHnWVI184DA358hYWRIMWieVyptc8K
EcTX3pNGwyucxP46wrMq4BF4puqEgylFYqfmJ6rOxGBUuyv7JE8YM7soYQfkMeuFLeZY3hih2pnw
cpE+GjLW1lViImDl+qCY+YFrfocdpsYxnU9da2NmCHqBTV6l0uWM7eYQTz4/vaJvWEaRQceEDJDS
sXCindPbfi3HTKhudUO9uT30TDAgDPnOHSRvxvqQCTdqw1c3ckYwTwQxzMeb3cePb56gS9rmQ/94
Lfe79OQOwC+eRp/17t0312IIAbauC41RrAmDWtn7OwrhqW2DuUN7fwnwAB7FbIR/N5ySHtUSYco8
qCkO4WzYv26oXhjzxyDJxtCjmVJzBZlQtJJSpswXNS8mrGgO1Q++iMVlWw6601skkS677ENX8F5B
bDn2l5CXZNk8UH0KkUCEiPpRPHAKvC3KNpau0XhYjTkmsusNa7WJnRKzkDZpimwj2LS2Sqw1UXO7
6g/mGCtV7o5EGXbkZe9NiqPeOJkYDABGaEaPQvAGCREcx5Uqoc5c/873JQlN6lwYPmGEEeC+wF1v
u0jzvEbSf/UPKPP68iPsTb6Ms0F4gdZO28lSOElGRGvVkDkgObriBwZPwew+r+LuNX1X0a1NolBu
7VaDByAfxbVBpq2lyFNGmTSDhgE4FkJbvhDGgHdDajI6O5RR1Me2KG8FyJjflrl1SNH/bbtn5CPl
9ah2KNqrTUO8m2bbN8/DSv+9j1w5WnPuZRIUf7m3HvEXD6hDGdyspTAYDdf1SO/vcwAxFUEmh6Sf
/cxFOBWOWgVjKLYJQYd6i+Q4vZcaQHhHhnFfJnPl8mUFi6RUl/j0FvXwVs9ENSN8LHnu+HBqdIb9
6sAlfukMm3U/95dANJfyV3SKD8Zt0BvPCaqUI0QWBkcQJq3itXFHKQ4zF/IuYqs3r5dLeLEiCMCZ
O1vq36jElcLeA59C+3/qgOxcw/AVvuePpR2dq/L44/BhZHIaF74EU3ExdJKnY1pT9NPE0a20gp1u
LYG2jH/ldiFUNRm6leOUSSoC8v1iSbkqWTjgmfQYt0WC9PfLkm36FMm5D7rfCy+Oc23nKsf5WuSd
F3lDbncxdOm8Q1L3hXz3kzngs8j1L1S/evUMWuCEgU+1ppDXLJPDmQCXcRUpk4gbUPk7vJl6GPOg
nbeREC3rf+lu6ckzB2qrSUm3wVGjpjWdy2/Vnml+5sarDTw2U4rwTcPjAnayWCPYzD9AB4hQVR9x
BWKbO4aWtU6eZwyK1PgGoDRVLSre6JZHw0Dzm9RXs8yyAWz7FXeY58mZ74r+K7Y6hfWboV3RR/Xj
e07ggBIgxI9ysc7qYNI2ilTD1V1bJsdYMwXtkBHv6WeQ2ZSFox8FLqoLQBT9vt/McKugHWn4iBWD
sNJM9S7AZIvmJJflFEsV1ne/lYvZ8WR3kq9A3E8tWLsJlEo5MViwFfwmGhzUKZL7Z/q/o/578iez
qF1x/mt6wbckkLZm0U8Y4nFBRGHnh43gVrn6VaD4pGvvZ+CuRH5vSZsnphBOGo0WDGgna6oC6Y/Q
U5HTFSgCWh9aQk56WwXjv03QAmBqEfJjai4K46T5ucQxbiUq/RF85QnT7TYsFHQY+ZxPKSsUFnJ6
k08PCNF6ZD9wXPVLQNKV7Vy/6pg9i30eJi0HYkiyVxzjkifA017QU8h26pK2bJVFlg5u8UKXfYsd
r5laF1smACcqqDP2OuRb0Cmqi4/chXxhJ64zl73K7Uf2hJGD/tevjNVrJbrAJBlBvyiLVIO/eshY
I0XTM3RSdR5qmNvB6JE77wMpdo0Hue/rS9AwQd9AABm4YirWoMacF8K931X3uuq2J69IQhzCu3+d
oHQlBuuh0J8M2GKFPn3Tqf2b7V1miEfYFQ0eXpJMXM6Xq7KhlmyWCYLhcgl2YuY4UMiNqYQlFNr1
62pxSDWIxFccGZIHnZHR+46floJyvhtoL8SeArCGRCgxe+LigPpGRmeg1NHzFMCs8Zn+pl9TSOW7
UHoxeEVVFV01+TXrgPtwGezrsQMjaj8pbktQ70amZgs5ExTpAOY1dd7pOJKOO6kl9psbyN9EajQw
ZspkkUA2o0fRch8++vh0XIRE8m/nUhnBuscnhxHQty0TlxPbeYvWmRwgtAGUzR1GMTzYodofpQkL
chEP3aodA/RPY9ETpKP5kH7fwu4mwzOgwcN9ioCg5vNXd5QOSpa2LGIWhklx0MJXsuD3Y7PJ3bdt
6uDKGRdQEd2olYLpPfgTYCRuwQJop8l+DYjvuZ2yvp7FgmPYs9QuYY6y2kYkhmJO5RnYjP/G81i+
+AJOkjLyr1c/EzrIeqIkBavrvxsetnTbPlb5WhMmZ6w0cx/vcHsb2Sc4RTEkHfwCMSAj8sc//mrE
H/LKLEpqByfw7RrtexY5FnXLa+NIvSYpy24jkJRy8MYDHzQwM90kyG07u0E7VD0XFOrYotpj9PdD
xzM75d+N2PvX8z/wL2FPqRzIzjOjW8W+rs8t+/dje4hPedPZlrzTsR7GAxEjI9YjBgwRpTNX/OjM
yRq9YNQaNppbzfypO0b/5Bu0MBUPhHYQlEnTQ3Jh7dyOE61svppwC4caquv7rxYNXtOw0KgBhqeY
Y9hX4oVFGUjjZscDIZ95yZQ4CsIWMf3SpWeOERYtxdjL8VVbJJEQ34QMJo3JRq1ee+NQg9dKCg5m
bIwvDBT/fALSUZVNjzXrwFC3JkFX3QjC/FYfs1TeLxTq5mq2MeuIDKOlvRooecJu+2hHX9KykBRd
giQnWqSYJ+CVgB37Nlt8ySq8o8QqHRtP4VVVKkV/X8pDukCUyuis3QAI2qvKnWJQFiZr82W5e7ja
7tkrcWIsdG98YdLphl1lBQHZCo/8Oj80wRZd2b10g+oGV4Ae8BwwXlGb4GOK++WQj3RsxBL0VVqn
+ZHSKiJygxweIOE0wwexaVuGc7+ll2CBokJyHmMqzynOAo5N2N9NsYC1hoIqKlkInDwd7xzCwIPr
hWIcgrf8HbSSYQa4dlK0ysx7QeoCyVvu8zuzpXdowAaUiqE8ObmikCru1BQfqBjAI08mH0tkArGw
l3a8+esF4tJjc2L4hdCv+4d0BalUNPbMTUyDzHD1VIhWwcfXtnmY9eMIyzEzgNmLYzwjpY3AQtba
P3fpsl+T6JB8fAyVI3lwP65Bd24/RVaNjaL1qYKbHv0VfHM42A+IQfMXmqvkJ+uuH+MxiOQ/5bHI
BeAA5VTg+uY1R6C39sFvSwVZBk+4LQWhwczqx7mhbQ/j521kCugPRz8IedWIsTQIuEKt2FDNAQ79
C+6YK575DNsKlQaQXohcMO4xp5X8fiwrALARDjVU60NlbWGQrhbxzCH5RuIDmYY4GKPq2JX2J74d
QbFHY4LRBm5vj9yF+8NUJVExlOzkv48AnlFP7Zt/yQkPjzOGNsE68tZDh74dIVZWezBpoh+dkNGR
38t4hlPvGWoN+ZJGhGZaN57x5GMVtQZiWCYBUSGlscUM6377xqE2hwItEWf49Myrq3OBPuHRbbCT
2+bH8sFANF0esOJ6Pqw90gW6NPQoTjxTTUowIoORvBUmTYb5WjN6D1f7Nb9WiWCdgc347t68hL4k
Fp3D18qx/d6khKbUWZfJjBOdO2JbNhVV10p/bFbpPy3njf6PWwgnjpoMhA9aDQLKqjSvkiHl4iLp
M3ruTmKCl5oPp5VeK8lqC/EFFc/msyL2qATboNo0pzkhwQdr+ESlhxXzmGgddvdIrJIcOgbrmEr5
Le0YKcFlP7oX+SMDTR6motgSchEg3nNUwVgdV8qO6+q7nMJJ5UrLD8wGi/G1bR1V9rqerKJR4vdr
1LIY1MV1HHxnts4p7H/fXAPeqwZMvdrUyK5W0PHIClint+r/8jNCKWOpuyVbWg/zYgPe8Djm5mME
UN4kPnDc8AOHiKl2Qow/YPhEEoEjAcoiWsExhSM9bL+FJ4hDo9Ku2ZaM7PR/FdFjewzoCsRew0dj
K2rNUVU4CuIB2fCit4Ppd1QnOCubbasFNSj6hvtTtrthTH8wUPhr/TSPCoCiyqahZH7HIxVvRVJc
NHJOdFpQe1bDBasB0q0XvYN+134QYpfPx7vu8Lpq5+s5YIIblcQ1EPumCpnIMTeo2Ht8BWbQuUc2
8AbmT39hJWe0YaQs9XxhKJR/vG35r0eXWm0vQgwjUB1C5UKWS3OmMPCdK5IfvDjXRh+E+QzlLTU2
SXjJePRD6di1G1hBxOFhZAqoQ1cnjLP88+2c9JBqBa/ky0R79i1K76HUbuFXRJPJXkHfHvs9DiD3
iTXfWlnLBD+eRyk5EUq/IwrSEcUPKxnUumvi44jdEt4aND8esyq4CYy8E4iRyDx2pepwOyqv+FnU
18Y4Lf2I6sFDu73eM9LgoaDxmnmCOG998ahGh7MYypyR36rKK8JfhZMz/AiAJKM9PdDZq9wcUx3f
rIlpAEjn1ckPnvSerR6oRmvUYqL3hJ5wJ4X8cenojMmZyqje5P4P1Bu7BwBvzYq4imtfUjOGJyE+
hZeSW4ITNnjD1qyWEBgDJYmE84zOY9o8Fo7cBgECTVg7sz84qwFEej1/bt8ZhKXrz35CSUyqAlCK
mTVAcogkN+LECp0y3WQlrD/qScSx4y8Fzwie504iZwtNfxDynCnpmqEIr5SF2qf/NKzDN/oE7ir2
2XzURlLul7eg+OakZl3ef73PYrDr+YbqXx+V6aTPZTvYL8RqP2wKB6grrachUGEb0KrNntEA5S/P
QzepGnQNPK31RTOZ/Hj/uiXcIo8jhbbzqKCoVeyXMKpDmU6WfkpjF49VqxtpmRFX9yqKltQf3n5Q
zd+EfbVz+v8Pwcve6DKRKC3r/0GEpSEMrNFZbtF6dkh7nEoIQ8DhzLfFqBdMWuuGQmk5yHYZ7zT6
o9rI0gPHxZp6DDnP/wIBykR3dwJ/Bgz67hC4QqAzec779jAiHeLxdXIPCXhxqwIzIFsO1RdLrB0L
6tEu579LL+tI3K75fTCtA8kPSBz4buhsVajMlg6FioFiqzAJEKFEIBl2841tFYsaw+emfZ+Ou/6k
u7TMtk4UQnbT62SL/U4E8YEbemZf7FQfRjTWIrcPCbIPaPnpK9rKFCFg+QgyHB7NyDN1XuAAqhOC
zzoQjiw3ZybzXDyql7eqzqH82rfS8y5MKXS2AhAyhysFqYp4kofWmmE8VUZvuDUfb7o0ThdKBBGM
ZGvq/dS/OwtKcWRjyc60gdyqlV69fLi+oFx5c48yGknwCOlAz+qslXHrlUoMfmdNw8pE4rgvpwZE
2yzal/NySFo+8hjLtFaq7aNhI2AcxPWDrZBAA6ivNYPdIARiOMd7Evtr+ymxxUhfjRV5Fdux/eWv
i60f3nmsdyzNyXbTeTyrEzS+dEWs5wbPEn541lYJB36+CKZrOlq9aHYd5XiZXhdjgDC7cq0nEsIN
4f5F0CZ8c2xyZGNzJ8T8cEEdT9d7545dhJqZF9hGA02V5hXApS8gLsKBsHi5g5VHHMaj2co77paq
GnRAOrGOY+eM5Mf1EC6yz3g3th9AsI3OMHIdDonNf2cPlGaX37uZKS3DigSjEFOzN1Wu5+oWROI5
o0fJnPOiv6nCLZCTi7N8bhZhHZwasQtHaj6TC98vWFR1vUQXxnOt62w+1FVlTGObdUXLAYHUXHs3
Bw4snSa9lTqergbtBufgd+Nf86Y3eBkdmyhz3wLkZ7cv6dk/nTTEv0ISGMFjDNcqKnA1aF3S+gpf
tUy+ut0oJiEW24Q9TVonLLzu0XQjPS6D3EzfrmJABbCl5PrrrfslfShksidLE+sSHVj245156DjH
1U4LKSdwTxD5i/W1sstDPxwHTr8Ydz6T9C+0Zj5T0lKQ8WDIG7R1GhLpwAHq2sSQsXHjGluJGKHB
fSCIv9iwwNo1xYmaYzngJlKXLv9qk5lCXbqBvWFBNHIrEsigGYSfSzIz4kj99WtQr2KCAuMlbez3
l83YiNjHx//XHVor8RZvyey47A3X1fJki37RdHZToB6YK0l5tUvnxci78+9sa0bVYN9o1zEjA8bj
z+kgAWafhSToiIg6vdC+pUBcSHBoulelpd8LW+qRBRpiSF/CG4X3Zfi1351o+90pKzVe2j5JaFpm
fJBNkgR+cuy4TUm5umcvx0JspCBpvsm6qGRwG7vy9pOm/NCu3FclYg/TUhFk4BJRKhgo6PfxPRqr
17KXbRSvZuKN8sTxIkAM8PKKIgCfGH/pQDbZcbRaORD0l0adGauZtCpVWn0DTjIYd6DR8JBmVExu
VuteKC/D6Agk0hYj2H1WQ7J1AAxrd+PF9wNIiZ34MJ2mi7TbFGqW0a0qdJ9fLAqsw8pTN7AHNtYB
QGCXZ/9nMUp8NH7fIL/35z/kRABB8Bx8fwQmYTfscRkX4ffeHmdnfAO/UjrvY63+7aEToKcQ5kgY
E8DtQzpHS2dzZsnO446OibZK9FSJi6/Ot7PZ/qtXX8+JPAX7GMRkn8atAZf2rD0MbIu7qcCbnnJq
pJmSksHkflKYJvC6ysI8hDp/ytPsBcXTa4fis+uZPqxH78fSobKyvUnEDvdxL0vV09Tt1GL6w72G
c7B0QSBRpvscuFrppJlxBMT/rDuDmfylZlgfEoDfYIGHg7DOhZ1vJjvImd0/Y/oCev8bJEqXfRHt
B/HeMhKbubjmuWatHfGLqCglv1lpbhL6SXIgVTSYJMxTNjznJkJhbmCM1PNQ/aMJVSpe6DW2FMGg
0M2DImcpA2RuX1PpO3OYjDWTKrcjMT7RQGkUxAoNeUIu1yBhRQ+HWwlPozoNMkCAfIRn732KRuWA
cIHwlPusQDFQfOdsamreHSlwSr+BSSiOfKfLsXIuCXHuJDgcoehfy+syUAAdsvaG9FD5RZV3Of+F
Kkk8Ot0+cBnNgsuuBFegJBVhgeE7Miqs41RbAoImAiGE84e2ny5aSOI0FNb7f5sSwrPIDFQHeCr/
7uX8eMS/EBA8KWLYyPb7YyIo6DMrElFbad3TQpbmMXl004523eDfnvHQDX64ew9TU2oH2y2/v6rZ
6ExEu2FQUyqG4GwysX1iIH/bNWg9T8Ifbm66uSRyEnQhd5y8gqGkRVSLwCo2EaLlSFcgPGZJMxKN
01QB0UCljJOZ3RwgxnqBvO8VLvuqdbEg0Xmzdjfi05NAQ1EFIE3HbU/YekemY4K7y84kQZUb/F9I
LgXAMTX3eogukyPOYJCNlDD4vWOT4JhZJ82eMK3NkUcBexhUpQSbNAqB7U78d3Rj+7F5/1QE3YYj
G+71IRB3wD3mMoMqeAZjb67f3adnzFaWD0JeD0caRsWWlJD0C76t/bslRo2ghhwCqbUWqfG1isgP
nj45yEXOOWpeLh23Hyin8Im1yCm78uJda+B72j4TPEpHpx+5Pzw8P5K1wpi+I/KeYyPClg0c1M73
scCu4gn7sTbxcnyZ/2AAFCqviZetP54y4WF+tJpWsXyCyRCyhkrFuLPESwBKSrKFpxPorm1ySt7R
lTXzbSDwREUMhUNuoyp1ZAEaxYzNLBaQb07md46kVZ0e+tcEgLX/7JZaPRLXdpAxC7+ZEgkukGPc
1jjByfBKQfyIgVe0g1892k3Oz/YA3BKB5cGmcMQV8eJ/xVf+yVpjn1BHMz6Q0mSyuWS8CPKr21gs
o9mBUJrJphiXUs1gnrtltLo6XQR5mqSQBaT4Mt8dPCS6tEdYtNba8ZPSvvZen/Rnx9roKyfw4Uuj
OG2Hc/ZBatzIaL8L4J6f69ayKNPngPRlDlgR0Ykfv0EluFi1h/TbLUdal3L9oyMLj8M+asYLnmz5
P1gW1AyLYEpXAlI1D0D3daEZQCkyyS6xTpjGe/J8qaHJ2Rf/4HuIDyVi28kcp+z1rUFAPq1Zc/Na
AnKKBYRM51ngh/nc4V06D/cJb8ygPP+D5NlVHQPT8FSaicQqVOOecvsmsMMlxloS3nlAv5G+g4TI
r/r6gKO/+PLOCQkz49cMYL19TlD7RSjg0S9F1Izl0CQcw+Pm8VMsg5Wt2gFCvZVrh0sEhRxMS4y5
49mIMYw7tYPGqQ79BTDLlka5X0LEgSh4pwigli+TnZTRY3d1tlaiDQAqA6Qcc2PsEpRPKWcoL9A7
PZ7E8+3x/gQkbSnVlacjJVbgbN62MfI0UdPX7GElkEGlNhm4vViInpbeD0SlxJfr/aPrPLtGntpe
Wy6S3JPNoixRvyN00TYYZzYxSx4f1OMnJQKhstyGq3kmKY5hvrAo8K9aFJkNKYZKareCVUfihsdg
0jNo2JLiVQ8OloK3dOxmA52DG3tH+AogCmtTbeUCqbzNMMykirY6rYQDgnChC97AM/jJOp3a8jty
ZIhlNUYrXO9vBFiB++cokm4htDzsuxLBffDMFvp7whqAkCMJ1l/1v9ZV1AFIGwqq4Dn6MdAB8tM5
7Q7iKKT2K1OsVXZl7FtYRtH5jjW5gY0de3HMAUT4qeOB6rd5EAT1VoSv3ZFCYMZcSfQJpkcs6gcI
bOQFM9vSTImqyF7FHmpd/oae4lIi6z0fxkJLS9uQh4nRR3gO5GkDlG/ox/aLG8AxEJXP3rlN1tq4
Lo9l5L/F00lc8wUEanBFlLBaMnaHzwiEp/qD78kI4FIiMx4FsDoEq6Tz/waT+Sgkhk+HITabbK5Z
7w/Cw3RNtUjaLqvGox8NDhxaRBmzVQMHgrdRbxKmFgKYjLIAfmv64t5zHX04/+zm/YLtJRtlYp//
O7bOJyQe6JrISrA+2WwVSmq2SDzd6iyR0+OmfiRojp74vQopJAzdQ3t1fEBB2KnElD0fVYAwywqn
y36LYub1qTprx2nza2zGFf6exMY+U28F2cQW33GXl7UXcTBYXThvPTX58lYZbJTmX6TJ6T7DDROt
ZFOO6AZDUqLUG5TmmuAbf6R/JgFl86vBo7aghxaJ/Zio3WyA8cnmUfotsoKmA3kW/qHXNF46f/jG
L+6fsPtIsLAyeheZkAoHtIzjrp+iebrGEGNa8Q8h2qajvRsT/5hxJtr+SwPGQXDnq3IMq9AzrL6+
p1eAocmDyIOn0ptVr6ee7cOC7ZVfjujwF/LjduFM97erGgBEj4UfrQvQZ4OdLbWnLqxDs15euN4v
q28ac5R8fIhYtboUkONIDULErQVnrNHGCxYVOT7n/GurkZmKqk3r3Jo60St+NK7U+iQwsEZi0TEc
YJXfcuV9Fr3o0mGcW+P8n0a7LZMlDhrgbBT74jfj/VxBiyXtk0gWqbzLJjdVWW4D48cieuMDpx+V
64m74IK89YPpJLajJ/A1CdVoUt9pdiBMKcknXtraYbcocX1EI4upgZryJQ4ntuclaJNn0wMqMhcD
f5cr3+tfaRpGG+DeWkfIWUkIrw5llrsS7IDj/9X6vB0evKI4Mh3OiKSQvMwDiUh2hZnhDFHhxZVI
7YDBNqegzyikpoIoGGakgrmbqPx6dBnXSjcHY5BNSWG1eKwu+fUtuzhwn7auI+DtaxaSn3TkSkC4
T4gLFa4Ad8hjzn930K6lVXVV05X/OU6NeKmgNEaaRezYL9D4Fb9ukiB2gH03Zd5JPkssEKJ8pGKw
kPe/SGeuPWUcIXrtT4n8aOlAS49H5Lct4jn3ea+BYWrwznDGuTU607V+oqBHwaxwWz5vhdAnKoII
aOXEwvRZ1ElgVnsAinyT0G0Iyhg/S1jM41eGNqj+7MjWm4jBsNTiKZ4VLXLTtfuRiKheszc0G0PS
Hhf8P10ImYYV04GRwxy1RAScBxhwzQDohmzq3NzGM/BpPL4OXg98mIPFTJicjmIGW6C6fcYyxmmQ
vJi3nHuwg+ljUWZLrt7eBwh6/KFYMMmNLa0PYmr5ArQPMfHCe5ZLiMFknXFcJ2Orl/Z6JfBgnv1h
K/UtVc1x9Wq5G6eAwe+/n8vUvpHeyNKzGDYjtU2DU6TIpO6KLuaooSkaCNTfQ+Mb88M7T76k+Wb/
JsYiTK1t6OFq1M9PX4xpDhi1GWas8UdQ0Pb0WzVZzACTFBFIeggvzoPmQuM6pfmTAq+95wKETqV+
1hEUHmrBq6JUHgZitf1Yz4XhZhmDFUqxz9KRzhsQyjtX7PmmlQbqlP6Fhp1EfzcZa5JWk25YWsSO
wWQ1uTnbedWQhsYLZFsqpB8SjTWVBCm6AAc3U94smmwb0cNcxKBnZDv+Im84wvYSnZXPg86zBFKp
KrwT07TWsodZqQThoA4jrD4LbGLli1E32+XoCiWk+Q9JdFERoJhSzBGKtejkHtLwHCmOebLkayRV
ZK6/6ktJ5247k3lFGtKrRjptw/eYd1O4Og8uRvKBpWUlrJjxYGbEX4WKcjUfbERUx7EO6yvyQpSB
3dYVpI7OP2Q6qnM9R7LHME3086cdXCMsD8yXi0z4fJ1t3fz4OL2VTAgA5nYMFVrBTaBn+/Dd+EzG
8x4RYVCtRmSQ1wAfmrYmsYW+DNjuFEsfkDDM5knDn0C/u7EWgcR7W/6KhjKZfiZPFrI6sL84xebu
yASPRPur9MWTSXMijQCu3Bzf57kB3qSqzkvsWyP+syYRD4LcZI+urc72rxOb3/RE/JR3g3eKjGen
22Vv839M3i0YDxjjIOMQ/4Q0nwqW88ZuqnO0CP/ZiiCjBBpUeBzi54XwF2FsAOD5ig8A6UgkYb3J
bjAfnLrtBdcxZPueHfbI4eG9G3Wqk7Ns4R59UCODra75xC1mRjSBmAFszciWYmmBF6KnZRUueqNp
eGy0g0+SxF7Z0WcEFd89AEbwPj/B1kw5TwgvmgAiym2HkDqAovvSZ7WcXVpwA6uvRWj4A0w5wkn1
4MQH+oxo8KZJn/SuaUhMhfe30VINej/Ucsfnc+XoJ2z719mlj3qtpjJwDj8ry7AaiMOCEqNgvKnF
zGlP3/EQj4bBJ9I1JJgbJqyGwBuTSmuHpXWYOQhuYb5/W1/Vut3wOM7OXJvUh4jt1RQd62cDjril
a0bb/7vKYMUTWm2+nLJmFtdiOoWPPSdfNwm5e8yWP9yFPsEgF9VkkZ2M9yv6rYd3OAF0t9CqGHTs
OICa4/vygh34Pk2HjFyS8smL2SyxfwWoC483LvrOXAuOpbY+0vyI2Z3U/GlfZNT0OsvN9xbTUXpI
3d1/sPILfVTu9DRB/MoN2aegM8fr0NlM4YaAdhYE3sfy+CccdG5qlg6syLEyGthDrUtAPbVrseJA
Skx+kwVw3VyTrhKOnPYUesQojphIzf5Bi69tE57MHCsd8hmlWTRoIuZPGKqqPkzPKoa6GYQi2mCS
YGtCl0QDUF0AMWJvO2BNsEuLJtmgeeKV/ZwtL5jnvU7yPFitMU83sQaZ0YTIAyrq3kZPSwVLiNep
fYSKk/xikqn1cTzzitIEtTkZlYnh737YYANG1CmSoncvWwn8b5O4C9UlRmSU4QCfTa1v2WA8FVrV
+h7e/jVgj4MNPEjd0ONfuUposki4Ua2ki2s3OVCOH+fEd3HaLTOfamx8bdLP2B6FpLX5b3nwrpgQ
/on9o3WIeHKJSWeCBf8LsuEdjMP7OSxW0Pd6nO43luztBuJfVndn7xHYtz3fKK+b4Y6udhfHAoLg
JSvgZ6P33balboynFcDyjIEi0Ym8xpTDW+7tZdNxTDumOPqmJOVcge56dXDPLKS95TqN9cH9fDAg
RmpAMQZZRCxqIK0J5K/UW5FwA8bpV6M1liNgCgAXk9fzQH2M5UbQsgCYg6bP02ynlVgw7fFaanYI
s9O3ILww+orufmrrHg95IO2vXHozooBMgF3t73Zg/qP48DObO6yDQ+jSBzMljK6SP3C/ZEH2N6NN
g6UW4wvpwriDLZI8LgHKTSi+WB6/Hxfw8EFy2axOe4cECzBEZrS54pF1mLf87Itj/aHrtRsK1RMG
ABxfpSyHBmKURUNKzdtFTa4V7eDEzLicP7qTTKRPAwhx41xdeRG+8CK6VJevvD6CQlMppPUr4kCl
Gy3KFY0BA4whVAELbQdPUm+tf9OymTcIoOp37wZuxC3HJZUvvn2gr+k8epY+HU8+sRbtMrDUWTtx
SLZYilr53NN/KulDAu/aEPtHHOzCqCLo/OrT9b9YKtOJT6kbTZB+458t6uL7uXOy1N5Zqs9SyoO5
a4xx57NB5QgI2xUHrv7tx5iVsh380biHBcu5P6TWpNO5OgTFLpFqj/bYGPLzb2TXoUdHRcpKzuXy
7nMLUMfff1jMlU/EdrBD+p4Hcwhik0Iqb/o6cA7PKJKeH0PK5ve2/2PvffEKYLQrSPe7fw8xRLqp
2SMtrS8tjj1n3qcvhImfo872EQyJEl1F/IELgt7Dzy8mpjYb85oCF9An4QHQZI6WENi9CPpfI6kn
QIB7vKbojOH2odrzbAC37fb02sOlb4IMdBBSxHJ23JLprg5if2TmQCIjxd7cdNLsfitDvjWGqrNG
e2S6Lk04VVFneAnb4lXwLXSPoZL4Klf0n1ZF8HF0CMN9JDQsjA1vVg7Qds5Ae4AhJaLhmBoUQsLZ
qBCkNGDyxdTUZP+dCPYt1oDQE9lWETIJ6Ou0Nr2jAmsqq4DpbakgUo7moAecTI1Iob9fG1FhMArU
p0Of61QKVzLHN6bygcNxBUykUFf1plhew0PYYGD9KkZS41Uu7Pw1ncYUsCK7q56r//z/cmztp+iR
+mqhQJgiDjbfH7qGiFDUacC0Pde+S/hRC/0dCpL5Rez6BjtrxG4WQ1lExGVgMEVA9OyK7MIVohAJ
3PEdx67OfltiJNmpJ2n1d1hOSZf5oKmis8P+boU3L5622WqfB+L70cuGw+bbaUf/Gh+MYEKgMoHt
wYDbVfYVnhXctM/wR18uB5JjztZRmD5nYdYKN5PU3X12yPkqZP5D0u/+Zn0JKBk4MD5+50I+l9lQ
uH4KY5panmYWgD88pcC/9rpToBum1pf1qBaXA4ppiWgf0oI/MSxcu7yFLaUs+6V4ZBfK+IFZXPJi
eNpHJ9Tcg2ICWiLs3dzWR6Vb4LBckoeJ4j9ehlcfmK89S3roKJcu9W9nf+WB06thnnfwNXGVy6Gv
inog5FMXm1cG+b7VXjJYH/urQwH2FXS9wmqWikkFYk9bRkv1n18AGJMnRjo8kBYv4w45HHhehbA1
7lhOmjVl3ZkjVo5svDud8JYbwWwH6a98o62GfH9z0rckdDS8i/Ev6BMf/3Fqj8iO3+PpAahrnCHX
iWeisZFyU5pP23o5H8Sjf8RcZJTZOUiOREbI5aL/sIV6Zv3xm0mI9V+uj7+ZsT7dPnZc/44BEkLr
5QzBElpt/VcakIe0wXxcJ4s60h5uFJ+Q7qP9bF2KrflTppv+6bpKCwsDb8z3tx21zfG9BJm3iv+I
JZkkhzRXFnhmsqOStnxhW3FC2+0HNM01Ku4g8OLW4zMzm7Q83NppGX+qZ1dHjOXQKjBzNkWR2D6i
379BG9zCLqtQcBshXB/+llocEHf4SOgUuqYAYcEDgx4q+29bvIqzh7WdJp8nNqMl6BzcIm4BAaus
FbVllKDbCGDT/zxkhk940Dm0/n+zjKJMArfiETAPuCjCu4iRDQvhtZhpyhtwltK7Nl+5Hqg4qrXC
oWEAluDbkF6xyaU3E1GTr3vqBhv0PmZHrotTn4Ag2sGaYFmRtoRKGn7EV7Agnth7UUnlLcmY8RYk
wL4gMpBFr44tq4sS+7XRcyhOnlfTlCTDhCmPNgBpNMbMEd8u4cfaZZ9vGdj1Ehjv1uo7PyiR5jIC
Ke4N9MH75V8HLAYHhWrAcq4yC6eJd0YCKUUONQs2J5QS95xYkvALJTa7ouSV61CNBVfGByd/TtLf
AxF6/JE2N9vknsElcsrpzCLASugnkWSIPHjFUvU4S2HP0JgvTgA9uQaHOXtXBx6868D1KfE4MiAy
JCjQ8JT1pgYKAm6fMTl+Zke//MYGiFiJq0Mr7r92Q+wVgDAr8/k0aZu5PbOf1yJeaAija4jK37Af
LW4ozMgM5tzBBWowyhp+AkvuWp6Oe8HyPDi+klEsyudHK9IxlqFa9AqB7kgR2wOj340zwddBA3IY
Qw6/MBMSmvWlG+WrGCw0q7auyX4U40fZpovZkN4N4TplSb6Krlsyv5ch81JvSPyTF9BkFen62UIm
+D74F9ZG5EYply8hAanUEDa6F4eT2ldggWE/LszbsVP5fkOeyrY+pQpzEbRQRResVFMVu9TPM4pA
xalutqx0ix9ahUUb05XroY0ZQwQMlkArteJCHpuaJR/zHAhkayxbCRx6viRckVEaCHmOQkQdI5jQ
DNAVRChDld+IVNw/o1/Zw66NyaVbcBxRctvevFFayVlr5rCBGjaYFxsX3ZD9m6IVDnpqdP7QZVL6
Z5yNGExZn2bdPUT11yp/Y42mvwTzxw8OZsGFx4w759AEOeQ3UQz2b0T76mn0U/HjKayeYsI2nW5p
9pHcMRFysAD4pP9Ps4GPracIJ+Bgba05fOyb7mkBT451Obaznc5AS52pscnzBAVvLwfzi+7aE2KI
bvTQAUlesgDz3CiQ4eU8hlzwZ0QPbRcsg/aQuPOZAuvV6zlB74AoICbtjDWgp9jg5AocBqC/EzQW
7+RPlSYf7icgDe0lY0yPJCIcv5PoIIVASsOnF6lGezhX9Lu7uasT4No4rEWq7+iQueYvONOE7tgR
9S816H7sA/7gN6dY8VS3GQYSHTjDsnMgvmyC/9NLbryCKddzFUwMUoZ7J01hu4rSVqIP2qp6Q5eJ
SiYoiLQja7NJqbgwYdx5zAv5Vg5M8GMGEDZpCYjGrpl6AgqVRLpGgRW5l+w7cgFrEUofcIYs1ZwK
jmPNmXyWA4AISwJzhxNAkucCm9/jppAji3Bh3Z656ZdzlplDZOfU8UMYPPPSVwn0SHfcwffmBeFi
yF2KY4l5ENqafX9GSSAyCtyFVrT+jX+LNlLQyS7Vs3QDXkKgzzwhThupHIE3phh/WvjPQHolYI1h
abRP2OkWVd7KxAD2D0umV4WVDTRlQ+I7uWtWTZBxu/ly5xKXgUmX9Nhpel8IcX/e2OWILH/q4kVy
4HMgnfevDVf7qH49cSlDvIKObK8ZC2phM233inwUxuT4QOSjkyNzHT6fgwtjFmLgTC8FV1dvFWaN
J2UwfICW6Nns/6j1TD+TF7AAMbCxraw8ZKk+hT8Fs9DFb5PMaexoiYTOEFBVnlBBY7c5tVgJUWr1
atV1p8soIl9YJpjf2pWRC3li4IFoOvJp961eRySOGywwAixDromgr74UCyYmP5gk+LNbENQRCJ4r
QnZaxNV2O2fr6CfdSiR5m+Z5CLwH6Sh9mMmCWxqw7glraFl6CmIsIwsMnG8d0wh4Fui45R/8bXdB
ndcuTZ7kOIh2RXBJXJccPgZjGTXfsbxC3PbiuaSNC+R4X3ntfFgrPj86WgPyhYTU/rnHD+SwcbrG
bH6PkQXpFF3f5H1YejELyLcnmyv9t5UUA76uSbydorqC3dhwly5/CStecUO4+ENJ/FDjYSQPSRu3
wWT/OU/p6yf9ZiMUicmy/HUUQW3oURC6KqS5dogAmgVYj6wMaVKfjwYdV83doz3XxXA5wJ3gYwqR
eU81/qzFpS5JXi27lFl9bAOUED/RSGTS4P231mpHqs89Whk5HyI48bm4JyPtWX+7Y4rYBzkwbA+E
Rh6zfGFr+wyfjXoHuZXaNSf78r8JlWTAKEB91ZEu+71V2waUDjRRFlf0IWxbacsLyK/EUwm2+2hp
dQo+ghmX06e7W/oNG007fgwP9BmxCxgih3E2QFVrSwejpSTRBfLH7CfvfF1x96oGgbokp/p7rj5o
1m5wQGtrrKoBy50Jsbok+7HPrz7DXzc0AX0NQWDleeFjDYXEg3DTsSD0kv0L3vPl/BNggRfmqE8n
fTwJjdMQhZd9ENuPCw9wxspJNAIqXsM2ZKA/d1HxcPvlP2AmbvK/w9U37MP71PnqGfd1to4RMTyD
lNWMFgt0S4/n5eWxWWj7ib4WZ16242hrnTNUbWT3NZ8TO76TkICYHWGo8oxWS6j5QLsyB0Bo8gfX
Cp3ePqDREXJVjuiiEusYw4lI4DbN54bYY4My6tyA2xGQXcOTCplO/S68cWlj7HVzcKfxk3MbLYaG
ER7P3x/wTS1G7LpSH7KvoIhA9m05u+/Mx5rRnYhB+zwBa3xhNhUAg73ntnDZAiHvxHTuwfMTDmea
0dUb9qBRzhvMz2Nj85F/UL9wt3o2VtOcUwA4uQ/+trGpcioJkk0IlN0u6tpmo4bdaC09dUB6B5it
qezLhNoG3tBnIFiPEJs8FbBBt9pTyDlijhSmK3nK4TfN0KOYVVcWdofhVi8dSOHA69mmYj4btOjO
CJw7bVkOX1JmWajEB3QZL67D9zoV09Sc2KVAYHg+nEUSGWra56SZJfydqHhibZRt3DWIHc4MTI+N
QHvRxoIoQ0xMrVtt1CLYxumeLSkGbt+9m2/1lKMjxMzblQ20q9y+Nfhr6gzxmy3uxAglO1Ttcr7Y
j6MA2II3i65a4ejTQ8a3Q1AnoIgzH0dYSklDwRGG3vtvAjHCQAzeTsf5vHvjHARdeE9KCsXT+/h6
lcvpfTw1C90DinNtutU70EADqo+olvVB+jWu0+6leOibx931gwBDf4dUAmYxvUnq5xBrLVxf2rnU
wKCDTMQAvBsY4xATutO3CjVkfPBu/DAEYGSVhmfG2lqafsNbRuYRJJUetSZkRF1aBWghs+lrMgJF
Ubb4z7VMz9JIBIGiWtanKDlyItrVQoFoGYUVjg1Ew82PoO/GAe6BekGhNGdJKgoavu22ZAPnKE10
rw1EvBEkOTpZsN7wwaKPt7i1XP8IADTFWcuf4bDZTX/haQ2qtD8DOYS8iYMugPcIJTpRhm94V7nC
DwboMqwirCwd8QApIVVVTCFaPoGVKXjTW99O71dosxJ4zA4SKZFA3es6eKEJkXEw9M4ke4rcJQkx
LZ0WTNOfg5Z/L45EHpJ/ly4QBBSS4J//hxOUGGXm9TIW6/QQ/kccgP/v2/h8lJbcgLdWMmuVF/Ij
TaZ9DZ50DjaonqUg9rpYPpuDIfv3TO0wO3EjlOBIxU8jUyjCFXyKwY3WNT1Rlo68M5Rcupp9eYu3
6qGVNvTAN6cK+oldeU5kXqjCLc9kub+FAnH4nRyeYi2iknCGw+decYfT7987Zaqz9J4t9wI2q80Z
U+fvE4Z+U+x49PtBA3JcWomFnVZq6N9Z3PXiNmcolt7UFjF2SWP0Jv8EFIRUaLuj3I6lvXiuAhV9
Pi7HMlu+g4G+CIYf5DNPEnNYz92BPM3gRB2u4ts3etAz27aON2hl8LYAzVAf/JzKaLC3mDz0msj2
znwuSQ2yeDapYnK8xD6cFWOxWiXvWtksFMMnWpmdAbyTuJ6g6xcltobN9Dezo30JZe4/hfvzETAS
PdsyI5cLqleXTeHWpW460X0vwiRoatH2JlHzO12wDHu6nrOc2Rqa3RSD/m0HhnWCCQbyPqrpQ6YY
fNPsdXKYDUSiItiInyNef5ZIFoveot339dQ2Vju7hm4+k3jy646J1aBfLatqniE4CHVgdXAi6SUW
5nI2mRetNxPybmKZwARD9S3lgieKPQhUfPHxexM2i0h6V6Xli7X9f1agySPCQTwxkhLK+Hh9jsce
ToS7aVQwTV14SEmjaqpDHCQA9cMH0g5X6/Kgy3t2lOQ6y10Q63uMGzeeqlZQq6LL2aaDM06dwgh1
+3Zxp1lPFLtEVr0xd9GbKXlzlJwiCno47KZSdN0RNc+nF1jmYPN99XUYXijjTTW0MWh9HHLlSmwj
Jkjb+qSt2PgwBPlg37P1c7Nl9G5IoFK6iKtHXWSEPdLihEyrOdK0eY1f3XiRqhw++m88yimwE9vr
QftPqd1RvN+TUmeMLnpglBncjXewbpKftb73CrVXsa0XKMCtRquxCmFhWh/psQZ3QQ26qHx9BNsg
cSjjjmYmfKWFiAdFNIBe8E1h6FxrMZjE48txFD/ihaXkMLlEH6t5PIfioMAMsFUecwkn1wE5URKy
IqVlNMkp6ywzt04ZWXteKamEqDTeQ8Ow7D3ovl2vZCuBcVu7DVBZ8EhtBw1q4lCSWQ9j5TqCOfHn
BZB/6TtKPIeXhAlyjepThnZq05oZ+ARnn17n+KO2S3K/ydMg2fzl7z/F2+19fyYbzZCGpJ7sfw3z
3JYHtgEKKFb9tLk4wGKK0EyGrhGvpmDfDsk99v30OdGK0+xhM9kJIrPXw46vGoquyGHs/vydp9jy
h4F4GspevI1axjkMtAkifN7wS1+7V8Vbr5hKQsumyt4vRRlct7PO/A2Y2u1Df1MzU9qjScymvMoJ
anZmKNkPnURl5FUli9z6EUQpDF1ca1AzO/jv2R5D9wrj0TyLYwO82suDtmfIM9GDb+4C4QKZEuV7
SvHpleNN7SR6Dn1/NDKiet2M6Ba7kJKuVzx5tGF0twR8fygGvWH78U+LX6a1AbuV+kejJ4iAcwju
TkxZE/+rG28CwHtHlm2ezjB/Sl1n/3iOKVcX1YmBmEL4Y85d3MqbXeM3kzM1WmqR5IBz7zqDlno4
Lz0I71VQOHkUJa+myrJA8PQeItyuFLk6+B1QFlCagWxmUmUxXo7oZa9eOtGl9GjfAjeW9TGkCOYt
7oEbVmkWw2ciXSaqdBGtg83n3E1tVN93+BqgW3RNgsi3abpMdp+usSJaUHyeSj4+mCgp7RSFGd7c
aet4PicKxoogbQG+nyQj8X5IowT0JjRnr3e0weSwuG6523iSwLCACz+3jLo2lqvBtqeXiQxyR9e9
ySYlAldwH98VBz8Pk1MTIJ1K4DtDXUsm07e53iXRIpHtmW2CtuCh1V/lPOHHiNIuuP2piJIgXe58
Yrit0Hmkvvq/UC4XDrvWT5B10L/WqITeLE8HcjfnIaiyM2bntyhelv5933KL2T7wXhy2ILwd+8yw
HYA8gM0CsM+OQ6HEZnwp2xaBaLaLgR9gTMAaiJZ7msTDgvAn4U/u8byULiZBOTuplXF0cFKyNy58
UFZ1bBweGMbX2Qfz04H6bABsqEOKCO8rzYldwu9pfSK0s/Bzu0obiiV23OAze13qmdGZeDvV4w5T
o1Y9LbNkP410WxwpcbOnLRP+Busq+EXbXPU+Pw5u6d1BknIVfMKmGCg9vQGB+nZI7bihuBviYYq3
zlhhcMo9M6hcJ8fdGB5DUn7Eeqi1Jsjh90moaRS7oVj1MCBLKgIf0UEua3ZnsBQx6bswKwaAmN0X
WxQVfbLhy0ahVHOd4oNTnaUBf78WeGOTWwQw7FPoTr+5gbwi2Mu1cE4LDxNFkPb6ZUX5937CtAop
4fYpN4ef4DTx2+oKCblxNrCZHwvg+i9RvCtNVMPiCAUUXYh9t3032qc6cpMclGu9+YRbgflIcfDL
1jbAfMFsN7F+ROtBhGtggjp9NUzOuOgpbtsikWnetKDJMKhbI+FqjmetaimDtv9yYkJ8EXQyEDat
10WwCQU2a+MJqehgtDn1GO+6q8KvQqWUKuELOYsO3yNQHgmRZBUeSXRY7cBXHU5kpfxNjDCIupSG
tlNV3QYXA+SZg44ExUPO9CnsSvAKjUlcHZhG93XierPMX14vr377eZ2k8tR3dW5Zin6J6RkuRoS1
2mg5EzdPpKt3VsOXONxgkjXXbpUO+AW0n563QOYH9BPGRBXFLXC5whJ+bx7VUgNCMCsBNjjjUw12
oWdYg4XvezuCDbiC/MSKZd5a7aNE36/lzSVftmXu1QBXQgx+lDpPXPqark2q+aZho1iDRoUFQJCf
X9hBInglhY3Yap+ZPeZQctr9A6AY4QzmymRzJR9wrG+bVOWMHRgghQbNSVBgFrKAh++sawQKdvGv
JTRjh3M9y9W0AGXG3dXvZtQtnWmtnc6UH3UVqY8y7JJb6BvZ2PqkBAkIlGMrKnIgHXqArXhbobM6
v7/iRuZWZOAyrj9x++GNtnrMyPx98vBuQgg+eMIqCa4SwEhHYVjNtrrDoICihYxsy4NYQ9JKZIDM
vR1sB0xvLEcaeYsytMbaL+M7sedKRT9Kmr8XNagzUuLlc7pepjLdB6Fhg4FSIu88ed0pwxIC0KTo
fMCCfrU7e4oJtdOcE+W7vSiOreMS/j4RRQUfBNwywxR6JTzurYopP4/9jKrGKzdfr0kHuXnYlGhc
YR4daoWPSByj6/9UgRu4KrhAjd8iNw/7sxqF0NdBPLl+KI9rtmUzOn6U5Z9KslRhUChXmbMRcMto
cIjAKlI0LEX6HAgaFtQFQDCKJD1Liv0mOLR30zXCae3fkJwDwi2Hpxi4x0YtekT5gSvti0cUUEps
qaDdj2R8vlyOLonb07IyXDAb6JLQmUZIcEsH6ghmk7yPRZcpKHwYEosbP0f7MI8OKCCinR2GND1m
uj/ie2brCx3Cldcnq3px7djxInKsQeV90a31s/x+7AwQKU8XGZvdO0mKP3EOwbgPMEWg7duJVpBy
aMDTRG7l8Std4tGRvaMVS2okvPvCKDleTR0zl/ajUQmsDRvGlP6SZQzl5N8tOn29riMxGmHzhld1
yUA4QhtVmuHH5gbx//hfJII1PcGaYqSe0CXjJEl2NyYJacTrn0XOb/gF0crfZo+NHQXfNmVbzqej
KlTHZPamkAlGneTGyexNXM2yGN9t/MsuCudyA2D7v1vyixY6afDBQAEPLwywmZ7JnBzl3bAVQ9f9
bK4s66sSlGO2h88pLytUAe42m2iScjTgbJ0De0J/LR0tyGJmlBNioGJumJDgc3wZ+6417ScBF9uy
qRlX08nb5XLTDdQOx6eEZ7UNZgASIBsorGz09/WDVeSEUi15LZXh1bvGm9dxKkvqCLgSgWzbpT+i
1UOrfb6wcN+ijZEKz5pjamC411/WqM7k+n5rWRYxJ7qPVcwOwe5OYsdNKA8oaGZVzJ7JR92mT86U
OUm8kJGdrMam43f45VjSVB73Jo8xQcRcYlVm6sMzmVVmD9EDtKFXv7S+A7FPOPlufVx0HKo0CtTO
jMEIjnHMxMACDLRDbZinozJiQlsZci1V3LrMigM58HFEjbd/+77I9fWXuUJEjMh6VcDh11Of6JtW
QLKtiHOzUahPIaC5pMN2+sXZSBtq8J66bbKTd+GX8Ft9GKYbTSFaMRXuEOp6mGFx0e1MzO3WFReG
w8AN3HVx5O8Ndw5x5dO9187B1rnGTZ1xnOQsVp9UovBG9PBf+sL9Gxr6PQm+2m+9iAxIL+Bp8/qx
pNhTxrKaV6AgrcZvvbvCa5qWWd1JAAaarZCIIFYnkCxpWeDFtBq9WiJyBiXdulG2HjiD+tKlQuO4
HOZwfmLjYE+K//zvrLfBwoTFI+9zyyTrxMUCz0rHAkYi8NinGCQsqmgmsJkhzICuk+l9wVlo3ROq
PAd9MLpFZIgAAk/duu78lQitBFH9YuUHQxGRF1xUPh2SFk18ivoctg0ANG4bYfU+a3pGatSz3PiH
Q8Qo7yQOQkKdnoP7PhajOkS2Ht3JeV+SkBdaiycyOLnaaDQUOiPZ/Afy1xjJhL4dcSlsBz/OQmk3
ZwP9FGeI4z3D+GuvLNfCYk25BMOfFfImj29PWkoUvAA3YkVJxWey7eJlOxJf93diExrKUeuQlR7z
zTizpHsTZODONt/d75JMw3CqfvVdcdib64vHRBhwzeGTa2CBunKJpJYm3APEp66zFFC4OWP4lptl
R00JxXmZS0YNqlREVkOgpvwJwORnxyWv20CnAnK0DAz1iUKgToVaWVHGuSmF0mkGtAts/NJEojuN
qv/AItHwR0I1v1vhyK2a7EPtLZhUYMTs/60rhEYliO5xXmnfuwCBhKdPIxC4L7FQ9F0wnrPqZvBt
5KGVR5dvAxGWW+VFiHtOdG4NJhaFr6NHTeSyIUuyVA3zEtthNPatLnVhTz4N95uefZ05cyZ3VwJP
uFQ5yvqDtGnn0NfZ6vrNTjKINdYwM/FKi5N3PXuLT4Gi+Xir7ohiQYe61nY+DZjLWWYijSC0gwo1
YYthaT/tizlhh2gTfIQnd2a8eBv13dO//6WIn45m6XxOJKLbNknlJMMw+u7+o4SVDfy6H9c93qwN
sS+D5DYtnQFhQ8wu1cY1+W9iQVuxlCHjWaZffM/h6fgQgsivredXTY4vbCxSvjzTYCnP11NnH6FJ
5W/YXFjR2sCG+zStRZvlQDcY4TcW6j1phHDbFT2FoCK3JVVRjiUMhmHwaXd4FD3ugFTEClaWL35K
FFewl9hSIgIPRdxexg/Vth85/gc13vKOWUpL1m05cKyBOp5RCAxo3DTmS7lx/UcyJNpQ2ORUwSIF
uBCyobIOsxPrtG0PW4i+z+mIMhXjQYl+es/cuh87J02ZqGiIo5Jcf7fiaiawHBiFmMw2UocWcZOg
2beVWZf2cGl/Po7NY9Zp9O396++VeLlVV0gIqdhf8hgsRtpg7IBaW+oz+jxsYLeaFcjLCyGPLprc
9+PpMv4MDD3Bbr9Akww1dB24FJ1Nrw/MzshJHUEbsL87OuJLy1EM69lyVhuaX3SUsER5oNcHphMA
Ii92S0phLSgzOFNvOuP5Y12qGEF0RnIkKa9YK4kesqc6Jrfg3KcHiMPmmSNChqeyzcparsnuFOvl
NoyxTKdEolHq5qfljaMTnyyvLny2nsOCrCJPZo2cqZTMM//Jfbs1g5qRh6eDE8PN+mp5exo/oKIc
O59WnQP+ev9rtzaWQYempHl5mFDwZ0TGZMkCQCk8CdBkfVwnjbLt5+BuueL9OjPSRO7dURrxMxZs
hVyHS+kydJ5KNwJaGHy+cRYRn7F7BcpAhPP3omqjFkS9MQ7A+x/lFDNkfJNIUxFhVNe75F1zB99X
92OKa5APN5hkYh7oWYkuDScDbD9pJEbyX3mWWxIsdzXe1ctSHq8Ba8SZPE3jzMHet47WclF69M2M
R9PQ4RBk8gwnm5kh/qIOWdy4ql2yTyOtCkZGCS7mxAhz1xUwt6o3uc06MI02rd/BpNSicMip1RNt
NFe9yRZGe5CxuMgxlGeW69tZ6Ta73eIV4jTJoz2S2gCT+taDxoEx+SI0kZfrSog8zhFGCJFrQuH4
a8PAeP28sBskKPbfNgjVQzrZUOQo/OSyHEkt35H/l84rdyrOk8axU+yGGkW9aZjHYXYr/EeUW5rS
9ZuUaN8SVRL0mMrpslywNYj3G9nSWTohFYp+9MD48grDn9MiHP2IV+3jSZzVhdeZdFDGdehYSZJo
WZ9J3whnkWMMf6m2AJG7FX0+oYeAkyeEaQm9JzDWlzlf/85kGKi2lySY+jq1NzH2li0ghZLl9ri/
Ok5xhF5SmiyFsxeuxSHusz+7AIXdc9OJ1UDsXwTdd0F9Jg/M/hihL4jABsFr2YmSpYXo/eDehQdB
TBt1W00PJzhs2DUoJFu1fH6FlpmvBTk+O28u0i8s4b7B1t5VnK+g+9ndqDDhaPSBnOzrQp93xVLM
9vmRnkGayr0Pro75Xs+7WdOrmJ8tMdPhEfzqppbFDMsd9x+4+A8a/pF1pxT6c8OgsDpbgPs+8k/O
xe9bhKTJkrROc/v7mop9U4/B29BFcouV8Gil4KDFseO8bXjmfTz+aGYidfleWtmxCW6+HdYZbVY7
qWI1T3V5Nna2iyiyVWPzCH6MceS6j8jhyizIyyAbBit4Z0AGpFrXHzQjVz6fDjf2hsJTk57q+gBU
3EyAcuD11wRPC1soaIlHxFluSYLEb7JzdmnCM4BZO+H1TLH7dTf0hJMjh9+OJCvtCVLcaeCaKzcF
syx7B+Trvv+73dZ3UtWffhQV+0Gcq/YYAE6DTt8hAKaMtY3PmI35mqDKzRkYQVmgZ2A8F9UDTTmZ
m88YF3JOP98ohyl6T4MeJhkF61YccJ8abSWN6UlCso8zb5FTvqPEwAUTo45yACklmXTdmcHfbDum
WpihhDpSzsT88SoK/Foi1qilpP8ObaCn3pJVnPwm31WfBkeibDeVjNN0zb+CXEMhrlzrnD0Ox82K
vLsV2wchnYrXfvYQypfxXMuYlzl8Jpe5lUvQSsFTB5mvFvX0Ub8Cox2zPYYYRuYr/k/hILQJswrh
pyZVGEKAM2h2cVeV2NZTy/naj7RgYsG2OYb2Dlceuqkvjf0qUVnaQvIgxehW6pgVACPwH0skmiKH
63jXfQaP51EZqTxd22G7y8uPk/UuEOPeg5jVGr133wNQXUK4Pg+iKYr6XRjPCMd6ov6r886/nUGG
k+nVJMNqKHFJ0aE5Eo29pPzWW+ZfxWJ6tGlBtGNhozJRSHvVdXF5piAr4B6+5BcEEOxxjAYt1QbQ
u54OhGd10uk0oK/iAKaF4mIYsBl+QZ4dwJJ0Bhdoxu2pflmRBqzgivrpLeLi1x4ReVkoCSgjWWLF
TFDefYGIXRMNKoNBKGHUyoH3ZlG+7XqnteztRUPCTp0aql+rkC+TmDf8MBcEA76GCIx15NShwqd1
oOaqQCYKxjV2f819pSS5BS2RjQp878AjCZ81oWYHWyUseLBuiGa7mU5UBLk4/d0UpaHJ/l5Nkl9Y
i7Qqu6FpFHl6rxqOPInGSX6kNF321tM1pf4fLxGBW6uqkOZtgiJjXA/4D5m/pPthEHkXeQw7fyT6
gtXLyBJoohsc/qM8mXrWxNQ5pUDflmQ2qZN/SsPzG99urvX6NnKIz1vU78gjfDchdzHzc6ThJ3rF
hzoJhU4T01Ak/aPrLi8wYzOhWA5f9z/1PMmp7gNoO196wO4kOo4KOmjQPJzmAcBBj2tC3j//lJr+
6XPQtRx9ezKjYMSCBHe0odbcM6SsNYac6+J1Oprzya4fGHxyG1Em1rDbdYMZRsXRRkveshBEzvOc
1QqyQ17Z+UfbmqxihG5Gym1EWmZ46G55bj7sLTd+BfMWAteV3RYGI/doZV7bxHpI2r4v4A2oUL18
wVD7moaaviuUqCO1GalyyTvkGhU1fnVepNtEDg2rawfp9Z9JyjNrcZdCryGKlQSAvEx8eJ7WxDnY
NhJciRlDWtf4ZAmaVzyvxrARdTGg4BeR8NMtYgmcwsKL/6BdWURO2N9OdU9pJ5kbLsh+k8IpFn7L
HIfgWNXz4K4cPFhXmBtIp0XdE79lIzouSB3jXWbxVq57doVSbPzZqoQY6oNvH99ZSqfGPj6KOygs
E7S02OcXN6rwDYdYgPDie026Q9Xoh89YcM276ZgWFZaHN4t7qHn8Nd8h8ncf8rB4x2MySun0Tu/g
RlLodGbhbi9akFpFpORfYLAIFKs8kwmvUqBt+t+j4e8HfHI3a1Ay/IDqy9MuoIsDjJVvpMOYvM+k
ZnYB508Q687LNKkoaNv7fQ8It2BCG444xJ+e6CRkcbgCmjqxLxUubLSp4aCK2sifii4/6j9dNBg+
MdwBxlntsYtAU93CKmtsz46KtFuvKMThEHSt7dhO1W218ySJyM7VgLhOMJJiMR1X8p4Yosr177W6
uQ4tBhzq3l8QJHkx+gC1YwLcZTf8n7/aiebLSWvINRL4IKPjKLlZCYV+rVpmtVGtjQv7TYsWugcM
1VuhjCNkF6wVW75gQpt1jtBmE4MV2or3LPZGvY3zS+jL2zqYHe7BtFDEB864NOdT1+CbJYkgfHbw
OxEFKrIXpelFqkX775GxjlDb4NqmQCmYlUPoUPqg5+Ucj3NTVT5ap/UbhhqIL7xXfjIOubhOuIRx
bnS+x7U3cZljgTntpKWfUl0RmNtyBS0xBg6FgwcchLETvlGN6J2q7WgZW401jFjTjXRYtxZ3h6Rs
4C1SOrSGjXvwcMWKkVN9DMhrlzzjbwHuvq/5unibRIQ+9lUzk18wkh7ygGLHHFOHmm/Tz2Rk8W+s
Kdp5GuQnitv9dyp6CiP2Xj29OuuTrljdmomXXYWNaFnIiFr6bWlSYVCKzWb6PNKA3eEhwJVe7wge
uzJqnop5JndwQSNSRVBAIhFTMyivgJT2Q9WYdqR3UG36AP3ehsuNSNpmc0rlCc5QCbb5ZAQwr4aL
VosPb1aOAMjqzWvKRsot6HVbsjHR49O1XcW7wRTp4rPzCFNvziSB0PphB53DgesXfZbaJh24wHuz
XfwouYMgpFXe+9laAbMIV39bMUh9/VrljOsPNE0Ah37v3W883RMhHzxRRwM2LjPFg7hJXs+HDzN2
NotoquWJ3QQMOWlfiMLruAHOOL5QrFEG9KgNgIrzyz0E2Do4UmG+atQdWyb7wCb42TzybkbNJnHQ
EManjdpCKHO3Q8XTbc/fgxCYCwHyX+Dxgf6ixCRpacX1L+RF7MP75UqQ6UPur/PNZci21qc7lxmC
uaetxsBbclF0+4eryG5Ly8o4XsuJW1Y6oKg+sVtMCZLn1vXDXUSNfVNHMXn/N5A2x1csgSbqS1Sb
yxVUgYcTZAZVQ8QEG/Cpfm4YnjkiOTpufdZp1CgpMwVxacU/YHAwPfQS1dyjdcUTiu+LdxHkMjF6
nf/jjEQUj5idqrUEvuR3V15RJrdDOO1YL2i4Z5HN93+rCnM7wNDOnkSMNX43wkiraFjMJ1IZARA2
G1JcQ70nxWBmR34i38kL9w3E/N3h0pSmfXjPSp1tbQgJdeknCoWFUoA5C2CJeamQvdiNkb0dVcCh
qzXqk7W2SHS5V2n3VmO9Cukh1Rbvf1HpQdhxu26IQa5HemIheqe0yb/m163UYrimEcboWt9ycjmi
GHWdnySAbV5GAgyx8mSg+BZA/Ro6MfFNrdEE0xZc7MdzgvgVCL90v3HuxBFlzcY4c6/Nl0OxQ3P2
qhiqIfAqzCbfoLSRhxpXYJeYWQVWXpbJv/cr7+/kWEHKZUtV6/XYfHc8HjgMEVH+tXxoXLAK7y1y
5HnQwOHVgwbkB0AOgMUv5a3GvjrZAJZSyS2eHcm+GxTifc7lr/xZpjoXWVJgMqahS94PSW+6+KI7
2MbT0OAk/BtLzYyDyN4AC1TzHJAg2kG2MD+9M/5al9PjCTIdjIwuxQ/Tyyok4BV9SjJfR1f0zbOx
WyyhRzyX/cnvJ9bFr4BXmHrTEnF1/qvZcVoKjt5EeTeVsg6h1cfAy4WZC+J8mWOMgoTGzAFbAHEl
wztvSwp/jyY1don/PvNqvVzWILbkCbnLLHVLchFHa6cZUvyYkWG9APkY7i/q6TLpZX4DOkIcMwlT
0yiIuqyfBW0Ajy3GWG6fJtJJAkZY8Mtlczz7T1Hrb+sCnSHu4x2CZuH6gtVh+Mj562IgytedGYTY
BN4cE5pbcFBvZJoyh0OqBOnp37x7qeXWilJc1WCqexrf6D9ROM6ROazUEFDoTVBtiLFKcW29Yhtm
kOn80zO4r7urwfuTaBjSyNKo8YQkmRvDCa21P7IQH7hIaVZEFlFfA7oMUzrqm5+nLSym330jvAbJ
UCxOZ60dJybSxogA1m5LjLPtwP+dVvm1AuKsZxDsb4+O6a2q6ksjWTYOZRyouDUiX0n0sxVWGSw0
I5wNE0tW9LPJ2QdUzW76ct0culBTI0lpGDrLTVSqLxkm9XDwBgjIFPCOPW18dLfvRU+mrSspvBgC
re5rRdrGPRXo9eADAOYNDABsHwpPKDrt0cJTl0u4Boyq+FdpgllXcEiGCU8LA/cH5mK0xoEbrsAz
g+E0pWORUUQ5uy5Yxtzb4+Yjnr8jd95UntvgD/KEG+nbMnRVkvmYiHl780vxXOCyg6mJs6oOnnLb
w2j5wCCYgLrAXNRdzc6MmlpOSl8xvQC9Fow+a86tyCSuhIAVy9xBF1Iu/tZquKpmsUMeR8tZWoGr
oQ2ILWO2LwAPgU01A8yy3GCTCCRKZzT+o1M17SLRDg+fNw7LRVoWvI0rBA6kcID45h/+efpVgDjj
/D+0XMZZJxzlVf9PPoaVsPQ/Sg2qnL77g3UrSrsy8W1Vtl44PTXuX3Lqe3JV2AXTSMPEpQvecuDV
7wSU3uwh3WjfvayQvvzs7dv7iWWg490Oc/TVrNx4PAIZTwc7ZFlQy797mgher1uFp98CMk5TybtD
x08GJuCRCN9Hzmx7cmHN1zaXV3weFgfB7+56UZNFyaybOetbnXLnbJLahIFvtmVwFXqBeCWQaF5b
lBSTG8GoaBBTXs81A4c8xj652I2atmBmeLNT0iuYqQIGuOtFWKTHS/Mu0c+CXEtSacoI8FO1rbJ3
sSUW2HtP4t1okggPpEJjOmjxfXyXmds2gAgcYRlzCSQJn2cVxdovz5K8MQ5bGOongvT/qif1xTrf
XzKPryBk1gCOd67Vmb8epvXaRfDZZnWP6GOnwRObULfp1OzmFPdMbEG1R+ennEW7u07ugG1WR8vq
Wqp5xO5v8QCnLWRCyx2yHhIj1/F/QqR4YRVZoU2732FZxa0MzLw7IAvZXiwXgEZVo+xWsOzjMxKb
bvwf4JhGXSAVK5DCwWZPRLVAUuUr7dMmbD5fRyNhFQ+x8VzbVT6EIpJTNM2SyN+MJR6C3WA+JFjC
Q9cz8Z3EdbJgKe5PaGZxqGZCrLPgTzgt5q/WYRAtGAaE9Vx4qKl6oU8jRflAVXuPgtv/WDZQFmg0
nYt5Q+WydhOlYtS18TYXKCB8ebSMbdsK0YcaViF73ecB1Ls2f+DOYd7knFyrtklYruNEuEiwl6SK
5tc1bHebjRjmkTloLQ/5lAXQPNQnv3AoQwIk6DjgIm7bneQfg7Alg6ffC7Y0DjAZ2ze67GG9Xz4Q
K4M/4q0wu+pT7ZKVcGuDUYPIiyvA+/4UwZkIJDy0EAi5DpfV2FJdUXH+I3OzVLEIfxfDxqKbQ5ZZ
Jb0t4klyMn0btyUllX704IoXS/ttC8MDFOoatr4BiOvTjd0a6WvHvk/o8VZEnsMvuQ0DunJfgVsD
uFfIOIjELnCH7BwtXlqTn1ZdGIMQ+6LBdpb/yEeeIBFrFWKmPYoTdl3V7ddeMjqINX3lDOGnmCG/
OAOMi7uNqw0EYeVaf1B8URB6n+goHJi4qccmgEtpaFLdbnUSIlijtRi2CsQcVr6g2DTYYopENEnn
CFRpZzhKgas4/o28X+kPUGZif8QhbOKVsKTl1FwPxHsOQcAu8gfvL7BbenaCEbJYlPfBxhKfdQP3
q/XgkQQ+ev47pf437tRKMvYvsbCJ82eS/JszKFMWc/YD408sBoKCcEKG0MEzrc51bQw7wa/uINPg
jTZnRTkT9lLFtuXa7qJHrBdDMFrcWL4MAUwA2gpkahRu0qAW7TA1nX8dzYQ84gh7mRx1USayAn/k
kNIyDxg4zIpoPZRRaK4o7SZVgIe691/zPCzrCOS30WixMScs+GBWNXN4mOuMCsPebZvyNTu1QeWA
/CNXEhs6X96iomXS+reRwpVtZL5tSDHM+n0poHv6QfoPM9wTf8hnOvxkvzwW4uRSwAZvYWe87J9I
BncY1UmTktJCW/MoXos1UJwJ+O3r7UeQh+KWwCwbsOXiPcyebT+U5VtizqUM6+CajBFnBVXJB48e
jhkT+bgMfBr6xYPtwmZX4tBgg7naVQuedepSb0ZMs2FGcqgXyIpTSBFFfLbdpmVqhzuHK/qAhLfX
xG3rb6MPo7HoM2UXooIrum4wOuU1sYIxB62OMPFEZKeK0RGUa4p6a1ShVm/2HZwK9QpBQomxyqbX
LibW5mdr3d4pvF1dwDYPuSqt29O8Abi0unAXmP/+we+y2I1vbZQrjQgShyuE4ZwLTte6rRJmsATh
nbbKBgd1m7epuhBvn82vt8kxDzEnLNG5XhQyL7IzsNziO2En1eqF9uR/dVP1bRrPUpWEL0jlVWBT
ZMo9CTotnTJJzxddGin0QBaiBmz+XenpaJRFyn5RjOS/VuMk/VvIO0gJ6pj5MY8O5LYijPdtQfpb
8FUoJ2lkNE/t4H8knpgajlYRHul1dr8WarnOCNMEEUmSYPbud5juQ8zy2fQl7jbvt4Aq/JSlnxvh
bjg7/CD6ZJ5xXsV03BhgqRXs953zLIdqjahfxEMWG/sZHceyWM/cvem1wv7qr6GjWB+2nF8ZFLXi
mvENXeZSstiy2c3EhmIqcGtDTqCIVY2vimqtyqg5sGU7ge9zLeE6k0BrNl+likeA2HSLoFyF47lO
TlGx2nlRmMskFpNSpZHNLtd6hHmO/tjgXzOSHV61ULCvCSfLpYYFrR2zUsU5NqN5mfyrMrJGmXZm
wBCYBczhHLGGcFLO2ApX/GuS4qVZj264nGo17BuN6fGpZCcztF83/LH4xeb+wBVFudBPABTQS0kw
QnUB4Ub+QUjRo9EJMeA86IDMACQgiwYeBRk2DXNtWU/HEA8vNPoDkrDB5VDh5JAqebpAKkDQg0Hm
LGs/boOYUvMiRfZY33pwUEFFl6vYJrYGk1oQ2UA92Yf8mAPYMLissJ6TvR/ktEa5VXzQYKQTvb6L
4X3nslXrGQsky5/Rl0eHsntDADVMQ4aoMeE5ICZF9/g7ZpcV9SRaeKbMEfMT26uKUSUMeJfK/4f+
3ipTUdhHjvsWduhOi0hkVsdy0DG1bICMRUPRr3KPz1HVLXKarN9UjMnxruD3givkM6z68++vVlyE
VhsWGVjsMJYLVkp5y1GLHWDRZS/4SYPtZfSvt0M5o3gq8eLqkHTVU0bSoAc9e5SRHgaj/Efo7tQL
RZ9643sEBobHuer/sUsVew8jOxq4uE64wUVzJ8SYfuPTI1v89U1SISYdL9lIlnaHHkyKtsbtQ3vz
RKJcZMErc37SygCHKHclLl+s6pLlbB+oaDjb4iRYQGY3GsAMBRFQjPAJ6unODDl7D6MrHxzXg4Ox
ejmm+sWr0jrf1+NddVV2RWE6I2Z9UhkmO5P8dzMvVYDlpzWIodmZzrmY+7IVnDYC/DqzmyESANN+
JT8eR1Ys8I5FHnYJOUCBQa6FnMBUO+uC3Uk2Y4xEXRNCZvL9nNH1n89DWS5iTDmbRgxFt3VZwfNP
SoGpKFzIpYXRWCX1YKRrg5YlDEy6hl0Rr0WeTgs/JUi6SPsRKNyXwso04gCZXm7aD0P1bQs8CTTo
vAyylT8+3nHmdXgpXTZsObxinnG91w03d8/mTBTL5xW7ITYyavtqfPOV3nrmTPCSWclf4V+36RnB
NtWuzDIOUvDeTneYwasRJcc9AenG2XaXpNBZFscgLd2nVhYn/LlJyY3vwQkWheWZRVeA/8usuAzj
hid/vaP/rn+i7ECZyWeaetOnKe1J858wXTg+jyIhyl1GokHE4Ebz17NkzDIfd4zLvPh+QDc5RD+b
vWpo/fuxLS/ykf0Yh+LvfrgfhZWLd2LlpaKQ+0YFrIg5whFfc/KDMl3baN+it6iwD7csxqoau/cN
0iIz8fIYNB89T/tY/oItsczibZXXE6FIwEbutMT1g2MNOBrEikfawmOC6L37wyNS376fc+e6BdIp
11n/2AZuGj2ChqkrjBhUP7cH1Lr+SBrqV8wfaWYnX1hog674BXcasvGosf2qR9tn4fnnRUxRCHRb
JnH1dZfX4QhDMsg/b0TVDWPgJpq5qRcaKWHK94MGI7OuPOLk+i0V/0TAvHMWSdkE9pl8IgESQHw+
gU/swypT39XkTkU78Bg1CjkGXqol866ZkPgg0vJ0MPHNPOOvRy3OsXN4/yfFuNlK/ldb14ZhvzX4
YAlJKd95rtria8VZCf8rsi71lWaRxRv30WXagdOFDF93YMlfZ4m6ncINu7hHdGjB4sB8W0iVqPKI
RarEXYVY1zLGNltFcdBO5kytxilW4sL5ab3i6kJwvqNqAFRQpzbnehrta0YveIcN9eZp/AZloDw0
Ud63LO6pidlK4b7rmdy1DC/Y1+ooU39TpDFPY+W0h8HBiPy8xmFTwze+h42k5BCPwuEZTYL3itUH
t6mxlVRY99G9Xhz7/PVENbEHBoA93tdO4bqmfcCa9C4+ftn17r7MLiIMNR+v1QrtaRwNm+R89sNR
DiKe0jhL9cfEXFk9pRPfKJbIZdUepz6DKAX0rsu27AULshgz8FvQYeerQrl/XCoZdURqzUTlZA51
HluTXHeKpaGViGvxnAPpk4Ayo1xUED/ojcgZ/2Oaku6T+q7iRKbLx/ZyZRq2hvShoMSUgExwhtkH
2bhVNHktyW1E9pkr3cRmqoviOce8aFz4/fLsiYlO24yik87GFolScthJvzu2oQWJQuISstZYcIh3
8sZNuXQPWNyocWeJgsgJXjHgIiAA1Ln2MK8hSw6RbK0DelxbMJanQHaMa+ILaj/m/gWV1AqWoEFn
bgTdlTHxatDPv4LpMSCdIZFP/uoxCM4w8PBEMGlsbuZ5VmJtnjqZPZj7GEZbXR+wx1K8prV27zrF
TwZU+r5PChijLVd07mGaaNlp6jMbgToJmsUno2TT+z+2b3TwirJSqMZkHs/RXcO6cAKk74DumEca
EdvjWnntMd55PSQB/+aO5W2bEkNAGPo1OeWS/Hna5XmpuD190zVQGZyFMOXd1260MHiu1NaqF7Sn
k+ACnW8icsF56e6+rWXZlJ18IOLi+0wXnc+N/llevOGklmYd952uSoINAmo6R2nB5W27KKSHtahO
4zrWU6/a5DMCJb3lcgs/LIf9rwHJszQaoHZDh3aNe/zX2TXTTQ4gTX3F1YSktwz4y+WBfPPrq08K
KfwQ4ok0ksasuObBGDdzXk0gHLJf49WyPScYjZZQXI9jPUB3JpR4FTA5lImf0ospHWAP8xrIXquo
o4i9UyDyX890c9DTduN4ZV7z1xbFanwwOT24CW4xHVwE1Yxx/0zItvLrGi71OCg2AiyqjQEiXjwH
huHo80Pawc+Km14/NRsl/nEUwFAn67iFnqdUWdi3P8nYEK/iqttJ/4Lrwe14VJuFh0nNKSz1qCkK
Wk+soWWBRy+7/UwSKNpt7ckERMK4/WRDF3YFhZV5FOmzdrY16VzhlmClCfjjxFHqgKsds0UymU6Z
rN5ZPKuJ4gIgSKjl0ow04ItGekmTDF4vIoUP427HZuMZzasSZ9znAoqw5cCE1JSO+g5vKOZKKiID
FocDqM6mZaxg5W1sy2e1+xv1EWTi19AK5JvlFUmRbOH2v8/l2MzXP6l5F9jCgHMslmLw019HGqd+
PqPZTlZ5CQg28FfFoLTOAsAIMGFh/2XeOtyJzg1L7hPiBx5SPT6dtHjJCBbXNkQ3BNoHSB7yR2zh
LxXxy0TxdcnONS0UcHYgDK5jNE8tBKjhpHchQlhR6l1tKuQ0iG7ZYPi2NCiQoLziyjQpKD29Lhkh
nP+Qlx5ufECa7dZ28qZH36oIQ3Iz8yKr9bZCDpTRp6s5qy+bAueOxuzdt+2q8OOfT21erPmmwwfl
06AO4IypHuiCQ6orgdwY3cq66+uPIb8hfBme+9sSjUTU3+ZVsfpuErlZ8MEkezKmTBI70wSkkUVS
+zGWVefTs6IrHGnX39F4EiIR/Gw3HPVUeZUYfSxW17ePfxtiFCpoAI8/8q7htgXrEEjllFdEVJm+
3aYEb/UocrEFVUCLufdwScRYNLG7mtJZP2ZaWY7Xhw9DXvAv4pADLnKru9FPp7gjhNg3khR3leZx
UBbNh2s1XE5QyZE6ZDvIX3DLAnWknZWcIs4Sawv8Xyz0cwl7ckLXvO/807aSqsxBZDCN7qvk90bG
KACXM6BlzQdemE+4n1k7emNUMR/tAz1OBDcxVHhCcYWxwec7xCH1PhvNVXlrQYFzGWdxa/mKYdXf
/wWRVI91N4kl8vRkrxABA71Y104ttIGltHs2KQ9Njbe+L3e75Xs2HISvtj01OgD5QWHRm2/1Ge6E
A23HmxtBGzuPvpmIGjY4aYD87gls+oZZq3CbJZfdmmqEgdRdTVJkJbpeJ1BbjbwYd4E5f7owpJSp
+rJsmleKvLsaU8Sj8Jf7EK5YiFH2pDkGRYrXe+LK0nlRaaqTtoYrBnFo6ejiQcgLqTKXfOYgJDZn
YnMKOX99sueZrm73yZISuBImSdwI8RyXXqKY7GfCsRYv0E8A4zmbM5CL9KAqfeQrZilHYFMOoTwZ
oaj47u724aBzCdvBLV5+EyeVekNtn6ZGpDWiqy1zOgE6Mn3n7GDKi/Ed+5bn8wGg446oD7rTBfga
cxRs09Fnialx2b2UliNDUR4OOKpXRCbbTI6WeDunmveqF/H/IZu+aqPwIxBDKyFAUVk6se5SZODu
WXQiu0UIkknUiOYDtCT1VzCfmW8aJHVktiKkiiYaKkZ3s7cmBqliTAJPx31lNvoO4boWG+KW3+yh
Fd9rGEjZwe+xBMicgmHWy+5WPAglsEIOoFN5KcYnF0SjuE9tbzePOy8i6YZITLfKh41dHnXX/4PD
sOkywQyMOxgsnsxuYormQP8DoF5yJFuPB0FPRB2WdtrmVD145zMkyA00aM8fR5R4Yb9awFGhqsLx
BKsKHwJXunSNqsx9G8CJd0OFdmkYUrYE6gt88KVHa5WuCispB2XcTLP3EKup1ANBA7Nk4F+It9t9
wwWH6iwA7ZlsKBXvI2iZvrdYQrM4cN1CVHWVVTbTmeOv2YMVaSape+YCn59h0VHvcRbUVV1prAzr
I3QRRXOSvlP51eIQGrZ77jX6uzT3HJylTgfQQYcXgadkl3rsjXgM6AHP+yG0zeO6NhA8LTfUMb++
+7RoV+0flt4fnSGsrUA6ItMMMtTUDVt4ZmUKjB/jyIpqkDRICvbbBguNgZoJXSX5JKnt1Z4+kQqZ
P+qLs6eM072t2sHN0gX5B8y73LG+/8fo5hOuNvijiwN329r0a4fJenmwouxj7Mg/fdPbq4moqnDK
/6Z4Si2vXStU/aklI9pApifMXP1cdg6UGX/fU5pr3nRBdxm6YxmOrsQYE/N8IYAtIjSEeEN5+/QB
YLP+fJPNFrcmFaj1pxKr58Xo+xw0Fp/WXcnEipI7ZKMBp60+18KyFAqUzgKNIPfzArmDta86Un0F
8KjxW3XEBeTk4NyO61RZguxEmELK8wHyplRqJG8eiuzkitds+5b1Jjs6PHXH2hpyFetJC2SIvAw8
s8C6juiN+oY5jfFoXGj19x9kTC/PEoDYPLwRTmcME8OgV520jl/VjUs/yaRzK7bkP1isxNt2eJyJ
TkeXBqno8PsKO4leV8bCpzVxmZC//sXohLl2v5qGMOJSpKE3EvoDGoFnxDbp4rC43ibMddh+5EXW
yF9z0eX/YRjvUPC+GjUwoQp0RbeNYG9uNrvcI0BaErV70fuV9xh/R2eHXFeLzdof7VJF5/gwJihG
Dx6GOn/4efjXIq5lDy7AmtKXriKQl9KVDmZMylvjCpA/SS1pAdqAliAXWA+K42cz2Qe0A/DjDom4
fdfwZ5ThRtswPxKZQ7oVwejTtIpMDH+LJ3VF0q6V7Ee8v9WFHjkecHWK2k8kBt4mZ/cpP2bGFFzO
M6LBJt/Gn59Zi+RzAczhtrHx/8jOapa1w69HiGhhPYiD4G+V9ohhR7AdNBprBOJR8CWUvSKxtBxl
D/DPBT5LIHRaRcYOi7z6Lti9ML4e7/ytOpqtbffBfzuv3XzeVuU3dWP/Y2UKzXDK/dl+CiNLJphl
WQgoXn1DNbWmwcwvLYuTkbx6MWksOfzbk/HrLWRJstrNTY6bEUEE5O2IsMuNMfNY3W1tilWosUv6
liK+6sDRhF14Fnc6X/KY1dCrdznkungsRpr6pBfaUSnT8II/0K3nKU2rxZH6c8+qO7hkLjMzXS3s
QYOwvd8VfrAZzJqRUti6GWMlk+ByOsQxDLIHBrTPF0okr5sFK7IuK1rxpjTk+WbfYm6OOP8E4KMe
0Fn85Dan9KhiRXUQN2j3HgAKkwDSIcL9WmBvHraj9Ckk6oP2jZUEeBdNkFx/6vJJ2X0VxFmQpgJr
34lZz5zdWdEeK3bOinzytjFwIzZtIePiUuCw/moBRCSyq8OAa1V5iFLAcI8U6LwiYxAEbI7cKkEV
il9YYh8ygt3QsjfZG7qRsYl76utURKdh/NtT9xhCitf5sw4FnBuJibWFVMNiLfjWUs1kzcNZy+uH
LCdHnaipoeOM80fFiU1VZaTENVPap5uU72MN32UZsZ9eMyCokPU7iwiWvK6lXmj6Ga1duL9sJ0+K
d8uRrsJ8L/d5gX7wDWGiusUMu5hi2pcvlFVKBnqE7FBDJISIX01YtT8p84Vk95+U/OOEI3KCEMXo
8M630zayFwFNXLSc14lOM6cSy61uxRoMuQAQDgzZeezwXodZQEk4xjP0yrQeEUw9nS5fiMCp5759
odU2feEADV3zArcYfo65PhlfJm7V8Mg3awWb20C7bhyMEUrJ4U/7wwDKJLyGwojcCEKQKoIus4RC
9sr6YqCSrFSvsy4OamgaVRUmhU+oyI6ExohOpVnEkR/GWZLPnRFZnL3oH995TdSBvlRXkhPTMplk
LyiOHwupLT1txYgqlCdjm0HRFynrvG8gTktsma2oH1h3vzlywv+nPpIiAaevJY/kOSoRMKbvCDBm
V8YO2qUZ6+y5seUyGHkvLTO2DEzw4CqVr7b9tgb3O9OCCpZp4hfAnw8F1GlnQKcmHmGQFhTI8mAw
kGNgDFQ4p8SHDjZeIpgGxco2EO9qLbEQwexw7jkr5WtG7+BdEQR/DzzrffuZ6prP+KCqeFxE/G6O
dYnYbaqB1MRjEnPDRlXdGfywm6x3m6mQAN4qbSLZVm2ndrIYGHAeBlgZMhg3zxo43IFIFAgtu5tz
ktyPhS683b20naiDhjJm/2vWAVvYfOYcD/up/VTYympJP+/zoT0poNeCF1Q1JcR66kcKAyAtgY2w
5kxirnslAtd54CUkhVikeQs0tE6gLN2ULYa6qBbVrpGXT3ZiKqCkKVZjoSoWnrU+GwliwkLiQrfR
tEPe9Clc1FHV03OhOz/EDXKgU4fHT0iUuPN+7lXFJMd3oN3+HD+RrcNCLtUhGorqJJ4GkP4bK/Mg
aUZ6vRyxf9leMnsj1Z5xPeFH70OvrFpkgTADGegyetL0Z7mHLWmbSYv4oXoL1UXvbLD04sFJmVN9
TjnAAG9UedSBokpyZrVBrqLU7oHK4ocZ0bqXQlyal2keSyOh+Dl52obDS8Fdm+duKUeFEUByArxk
x/6hqrbRmFrYRsmCEVsOrjrnXkgofZLu0txbx9pEOjbzoFCDMCOX7ZlXxajR5bLaNRfKsjI4B7fU
IXqBQu6l53aM/solfIbZOayHGNoDVN9zxYnRJXlJfFJRmAdzKiSxHZN4dY5IlZRTSuebtBNEXODO
WmRluL0Jb6/Hb25WG0RqFBaB7Nf07DIPGA38WeSPuYdcogC+AZp+3VDQE/iGuPyC3WjakmEW8l/N
5ASireyf5Ihs683PGvGxuBKI3/VkYvsyhmhVJ8Jo/tU8KFVQ5nUhzZ5hsQ1xXsxbrPtDHBvmsMoC
NK2BNpBTrSG1LPI7RVTfL2hVJe4wViz3+8jBdrFxr/87GJzGcUMhtkYShN7xSTiswCKRIG1w5XWV
ks45ZAiL7zj4rDyuGvCgyE4u+a/5av4coIppL1GWrnqBR9mAhLE3VWYtGwhofmEJHsMUZpC3wWGH
mdWHL6+mZeKvCS2AfKfVsMriVZWzFKxUHqhaIy17565gM+L/HBl9CieEaE8c9+1iX3Nd+Sw7WXJc
TT2e+evZ99i5jcRatyssKeZtHX1m6y9xua9LTC8NlxPk4pNwYX/XYVemSDhzi/5JIE+I2KDcmUYi
xrKGRxBJ2RYO0RufC3VMhfzX0E4v+CygPOL0qsIdXcK77QnoraZHarx2LZOw1OPvwBXU4Nmwr/+M
FrdTBXVrS64xUfSXQkcUrZuu4estgWvnDDXS/9l8LqixWHi/QHC0w718Fm0LbKGa5wJqOYQJYVxT
YrfrHznYYK6CImteSO1lTEeXpbSLd61sw1UDUV/0Qt2dpAuLsRGR3Cwbmu/OjxW2kUvMjil+f8Xv
TJFHVIqWtDAK1Oxused/tlCw098evBAXBPLInySN++iz9kG4LENnlqA40Y9XjBzNOhe4VgRpcqrM
NN910SF+BUAbzcfSLayak1sm/efB6aJ7IdMtaWwSZyd7Gz493NFdTrAnt1kl+EeiCWQAZne09Vaj
ivDMRvM5wju0hDiO/TbEGp7i10umBZHwNtOAZqwpTnUVfGyHxNu0DJnLBZoPGqRS1BGWF/3q6d1B
ARwu29RnGvbIAb6ygTNA7GEQmuS2Yww0kO5KOWStVuYkl3VRN0I08yrEoblLR7+VzaYdXVfwv26r
uVUEEqXKh/jlTDf0LkwCUkYrnCFRG1lGPrVfn5UehUNA9IOz5I+V8RZqQiPEgPtQ4hMFgOTOC+gX
V5ZxudakMCpL5uY4J4noMvOuJrh8pma9YNRS8DV8XogHXVUF8gDctbBgsgBKFPp8XzwrlR4vWPbC
nK16Z3PFbpK9f08rChua8GuZ+WNNwwYOqpFP9pCQFc56MsEPcUgy7mHvqvLUu600j67ZNZcodcAI
DfZn56Mx3UNZzi1CIJupwfJGfFM73osCJBsx02XF6CymRQQzkRWLZwfHIw1HP+k9XyODPjjNV7fD
xDI8PlWCCM/IWnm1lyuHoFiKcGKqnJLMTaMpNzOIiJnNxSK3xHdZLBK2xt8DzU47dg9rQ54ZuKIM
rygjjGs+H0jvEVGEgYmPpjNcIhznWQUxXrsZDBfwEDnWL/vl7cwzpVvoPaCZUpy7D/nW5HE7RLEN
Mb9T0jrjuVc00wmaeVinuWtYEyo5pJU1TtOaih2TSraKW95+wamBsCebv1OZnGFsVwHWMsgqzg6e
8ItF5zY2n/yfme/hmnzFaQlUbWmmNZQ5U106VflEDUMOxRAsfwM+FrTJDnI/sMhJnYwz3Fao7x0X
tfRa1hW8O8PsHG7H8MZk4L419dg/Ct/j5d1XEQF/Mbec2GE0LegC734a3cifMWyIP0cX+Z0b5m0W
++sGBEahkDnZQpvrcU7QIiIhgQwQCsPGJcb/Bhvojw2s5KZ9FbK47n/Rx6THvKQ6IEpuQn3QJruk
fK6IL+KSZoStbl7iP7d/cxOFKCRj9vgGT/jPS1Ngte9KcTGFrYlx7jXmFQA3rPplRo7aom3UGIjQ
8E3LOp4Xcia9JtXQZDtee65dxYzKYZoIh+CE5xCqt9TdAUpVDgawFyI5lLHf5wzg/6xmt7j1c7l7
Ags/Jl434Ugqa3eLAcUvVRqVPktyff23PNz9pE+43nh2XreoaPyXTojZ+EV3cGFNRc9hrTdRZNgo
1CAjUj9HPHPWR2KoAKMI6JluZUUMOGSAscG9WYaPh4MSVBzj/wTCmch9vIpRFtjAgV8jp528o27S
fC5+PvVA4rhB5NkB3KY16SmzlCtvd+F0TeTCpYVGGeCi2c0fdtaPltTnGR+3u1aYbE2PjO8E/s+N
lv/3VFL0zg17BpRs/92usSYgmQD/AtQ9eju7j7b8QnFjyRd8jwK5evz1hrrF9cwTbe39E0qeeZLD
wUCpxtRWxWTBLftB3e2VODJqgQlHMKpj9rwA7IprZt6+l6vuX1NWquA6y5faxRBBGjAupxqP1pAv
SyN68bj/jvZ9YCQugBb9VyrIMaj4hPO+xcrtHWsudIRhDIR3beVHnAq0flKvbTt6GlmDjPMKnPYm
ozuvsOtAeR3U8hleCNBnr9WQF03XjiWmgGD6r0KlM4qwSfaSWJjDQgmxpVgPNUWDTewixNnq3ooU
9Daae+e6jThl8sZNSE/7st+T+6FEjVqidO+/2zQJPxlr3Gkc+rSvmhoPSerP2cEz3+U1D1n03R4C
F9/uECdm7odp+vOoaogQZOzgoNR+FAAMS5esEv3GWPlQ3GNIk648NdiVhEG0KrppuqzVU06W3EnV
Hw0RKjzQ3ZFFsDrT8C/2+6dhq6B1A0ouuHL9+qUnarbIJ+MuC3TCZe8YivFuKIxM/b5TDWz6QHhK
7ETfKIYXKoQovtVRvHWa7HF2vnnqWCR2i1B81XlClok272UJAQjXpwi4/dcdv+CgERN/UqFnVdC1
2Bx4G7VOuLc+kWDz6nmUtVKR6ANg/FFmrW4F+jHwBHy+woXweOQhsJ2S9tWFQKbfuuf9JXJsBRQp
mETV4MIE2psmNbDwGIMV76f/8hci5IK0hGPV9KWTbXlvKEABg4kD/o2mw1J+6lW2iG/ILeMeWDwY
NrDbdzxDuv9kMuQNeDY0xfECRt9bc4aNZlTbA1E/fznS4hWDFK6TVmza3NINZ3OzIgIUzOfohuSF
7iJTZn+ZJ/wziluAlx1ew14sWFQ9T+ouhJlBX3D/MXtnXjloc6uCB9M2Dwy9yllgQOOEhV81ZZuT
8WAP5yN3FedCN1KoFz+HbIwQ5gxXdul9jtoKNc825AIohgdnyUw2M1CL13PhVl1w1QgXXHtQK6tE
ofOfYiem6qec4YVmfOClbc+gz4UYqTDDg9ulKtH8B/9JSrSvOSqT5Y3Xzeexb5TSfDpk4kiPnhg1
aPZx1I3dPyR+uAIcdSY+ArkxjkrlROFcWkLDqR7EY1DAddrVRtzQhdQm5WrIwm2chDgqgG/XA7fH
FZfkK+8WrbQuTQRZv81rXPfFE/bn2E4cT5vlBdoxsLZHNjgs+rcWV8AcLi5QgflZPM3rmRmX3iaT
BIakxk2CcKBQdvF+zJCfBfr5LHb6Lx49kgcq4xlMr9Lo8Ct4DXAzI/45n/XwVINSZzWLPC1+qCFe
1k4X7OYPGQ8GkRKWbmr5MmWatxTFT5kc56xnNc7YwEVSDF0AbViKd3RlnkHsyhHEAGXCcSQpKoaS
nu+nhpidg7MvGOPV9ngscqzGJt8e7t8dX7u73qh4+F6hJ2aW19gN7/W7ekIWoFkXx4lF5mKVbVLN
UN6BI/zZSOTz4TUnDdvy8HdUHMbTGu3Ac5JN5suemUTumc/auXR90CxCmkAaDRDa595B5/RHribj
eQOVrf87n242oDoB5yYWJkZwXW0OgxmJC4qXbsLfT1TDeFb0vXUMxHv78nONjCcll+pu8uZj2NdI
oyraZmikHKp+/xEfyLyRHvzpHr6+RMzAW5CLjTbphSFrtNh5x6HT+KGIhzX+GQLD284crcRsLKu/
lb3GLUigmLMDmFxDCC5475zbJpiX8t1gS8Sg6L6T020hwgkVI76hojQrPicjQSOdSfsTaqATk4pR
DExVU3SSUbIWF8pI33YgKObTDKro5k29sCT7LI7IZc9eZIYDYwqtLIQIRBr9ceBQ7ijoYRa6GHQB
xsZZH+Qd5MH8IZsdDkniW3eCcUFqd05KmQGZefAg60cWhG+BHPuXubscBByMp3K0jMFgUuaDCiPG
PqiTGtKOUgj4OAIDAdQOFcHa6CT33+SfMgnnd8fyQOmBxMQH2FlVsQvmTYKQBu6XmOKyDA5025sK
nOYeQ8ZEhBGmTxSCia5vFFfJKOgZ73sUHDYxAdNWaCUoGr8XYBHMkOWECIdyZN1XsHTiPr/K9LXO
P1Aru9WrzDGcmXl003Bj+Upz9b6uVxnTRNBJbt1Wc/r2hN4wPWHBhGWM+XEurb0PWjhOEUpC9i0h
ZbgtKl0eSN0/802O4xCaKAXRKAevQhZpgNLxYOiAJNMbTU8tw0Cx8YWElzc7o+AoJzGHtjWsRs1k
43Krge9NW9jJ4R3myHz52bzxm9aZBd6q/sYOnD11/YlnJIRAPL7Z2LP7Riqvd7dnJ0wGOf0YmcL5
8sLSQ32gSmjeelMJFOLmoSb8noh7XaOGtCi3sB78LPqTAJWx0Ns9azDXe1mTgnW6TtsEH7IHQhQw
KMSI9rF5Mik4QMPs2ePM4ARRxU7bP7AEGaKZdzmXVQgjacdcpWbshdtZasvUqQhEG5HxWgELAz47
w3Jpn+VEMcrxWhhcjBeGZit1rNqFEYEYiDA7B/UWNibJU6xxu6XE7N6rqddMiJn7/zxuLhIk87bY
tm1hN3jXOyr/TIYPA/5+UQ8CkA3/MuxcI/LeJXUFda3YTY6zmHRiunM+4jdoNexNEwibadwV8Uwb
cWLAgjABeLeiFHxEGBLfJ8qXlfWnHsCLDi+N73/VhzI422MgumB4VsDrgzGt/ywd9UdJGqrzL9RQ
vYn55PSeDKRrTwQG/V9eZ4iFX22peOk1/wzLogmq5olYf5wBAb32Zw8mTYAnjCaVPTN96lPqsKcf
wwanRUiufezZ6frt8//dYC4sxuDjwWVFl0nIZ6E33fJLeNjZDbE+kiJzjIUFMO1gsjYuFeR5DrgX
2B8UJe/3AFyzY0qHvhIb7Y/j/s5JlsT/un8IsyxyHy2tpZGFMVGpGnDuLlkUM88jpSPXFTTwu1Lq
y0y2kliYHIHfaONOinNpraZWSKwpuJSZzKZaaFlj4uzkM0+r1Il3OkPR/3pdXzJ1H73XZlWWrQGB
Z7ZQR00ZVGrYr37P1VZwCyV7cL71B8SJXxAuInSqVsKKFK2Q3Opx+xGJTTx2d4l5rTHId9S4sCNa
iWZJXzI82FMaLIp2AiYif/3vTjJUddU/msTbUFFnzEQvF3IJI57KTc8WI7HlCjpZP1vhjeR8IDE+
A73OqiZvWGDHXPGBg0attMPXsUl9wFHxnJIhNLkLlVYoFeYX6zYXu/guvof12kfLGhlpKmdaV1Xe
o75XAUWfGmDDwxZbpiEVqpeFCC3zljiymKn4Pas8V+tCrsq4+jZw34S/VPSL0n5mVjw4pv6kOuyf
RJ5uMkfvrTW91yiXJS4OiFTBTTQOX0YBQrcZTqet6cMu5N36StMeXFH8BApRAnfgnl9I6chxSMVW
Efaz0q49kVKVRdst0KvyInL7xTT6E8Jt7u0VHEdGBf9WajA3PeMigbKDfNLRc8x6DGFxDWFleOcI
E6M3p1t5wxhxVa5C4nayvkrnV6yrUxWo+4ZwzXWyXL0516JAOZwV6eFZ5BiUIr9mqk3c1szH2gvv
xbRwweSuufXOzMnRJpSTDM6iAEFJzWZ5VphlTE2nTYbCSlNEg6NVlbGN14jQJMOzSfCMfXXiJVc/
I0NKoZqj6LYt2A7PAHkuP365zn6zfPWrlqCd2HzcaS7FYMM/5U+Y88g6UppmxPKb4W6DJozPKT7k
Xj88+ghrIvD4IR7GUYWrFj1ZPLlIdWzGzA9cVshrTljO9XxPdMedvIUZM+8DmcFWSDy7qEPitG0g
oxi7yKUKBrpLHCcpoyngom3qOnXTSDX37LDMzsAfXzmWMxGeUyi1Li4PqrOLrSZYrV5jfRQWxt5E
zlTHi5krQVdOCW9eKc5HvzE+DwccA2lB8BRncBQK1/9a5qomtzZ12GSA/oq92G57XmYouyF5J9B8
gF8FyGjFGN21VgBiFD+BmrDWZBaDhGYD2zV2y+2J082p0z+vAFpZUZoxnMsFWzm9m9egFtDXKTgR
4T/+lw6ngGDyjau47kk1tubA56qPasAkDhW3S1dGCGiY8b5lcvIZ6dutOOLzig4lhlTKNKJMUrQ6
E1wgmM+vjokrz/YQwSKyFrhQH37W9iDH3HDqgnn3BPOGMkdLqXIg/BewJwWppAL62K4864tWTxvB
ahEZ96bpXl59RitdzNi0moQjB69dUAgE0AFjHGk4CjgL6CF7PppxLCCVNeR9nUhjW3ZDJJByajWh
YP4juDReoz+eU15MJuTTe8EIna3E7f5xz2sC/hAk2DXfASHKzj5Bytpmt+IA3Vv5+OE0fAMiARbN
0rcMSTxxUtvTRUbFPfaLNz8AcERdRDaalEexnsqo9cPBPJvDjJhA5QpMBhsLgfJ8V9p8wXBlCkPC
/RQusrmeOT7u6EqiFjWIuFEsnmrWWGn1x5hkPNlnxWgPsdoa0ts5kVOnDAwj4abi5dfKaC9lOuO3
m9i3KzcOBJNX1OcPRbl6HooS2U68U3bVbKOenrhSkV/WJ76yS/YfutzpyZ1kQFgMTW+tpZYS3AVH
IMkEq8TETRclQaiC363i4w0XSggAgVIHJwbbsJ1fgpSfzEaZm0qb5qlJPZhyBGEKsX9pZ31C7Jpo
5SdSgfVjr2lue3cALpZC2RfFoKOuvIsNUJRUV1wx+PmGvJqY/z/5bpuNJAyGkU9YlIwyGDQiEm7Z
uY7G4dtrYKOKwckHh6BUWQx8XeFlyT70Uv+N4jOQuh9NZY59AbaNRUxVIKKF01nPhv+kJ6Mfoob2
Q3eKYnBs6y//XCUuabFRB8wjg9xUnP4p5ZAr8RQJpcuo25ZOSom95HYZ4/s+WOwu7ZwbREqokEBo
OAVBzR8465SpTaiZBW9rZTAi0AFQzS8FyJKgfSuw0kCq6uYp1bzjSFciciQG+COYIdThSA+voaTv
8mC4h0zZeJ6Ss1GXdBioLcFVLxrDdoPXEVMuYmlLGiBar6GMEtCDZ4Iki3WhBNAIGH+hah6ZzKpM
7Kcn2H1Ataf4tQ43ZX9tsnfemiaP1qqp8ancNVkUvAzbqgUp1rV23ymGSDsLBqIHcvKyr+94fFvu
739f7Dbia/EPz98JWZeQ3caCpDbUidHVvB0wpYuRvZbk9+3gBKll+jtzBulh3+B8kjOBQlvuWc38
Gl2kLgxi0kaRSbdf1JEhrYAOF/2ohQlCukD6A+YrPFsYdS9KiGaHCSjTVzn5WG8HzrKaQyTxc6Uh
yoFmK49orPw8DAG84rvKrWDK4uvsNupfdJ1kxuDcwidMTP7S2UkMp3zVf5oftJsB/32PepU4we66
9MVCfAFeJfU8vTD+lIPoQYXUfNqjlM0OcRdm/w7x505sO6LWHKAQtH2ebCQw3wCVVgLyou6EYweX
wosFBwCWgWdo2zbw3bI1rlRySQB1uJUHsteup68G3ZQNOUCLqHwMD2pSjABrIOrjeCuj+1dl2nFE
j3Rs/Y4ZabOiYtranAnzGIKj1sCxfRc8K6SGyniQIPZPq+i2Q8sEOwuLqXqC6GwKjVo0LWR+D9CK
M7VtwHq7J4ga446xJKVcGGLFqefW7/a/30rNcru4Nghvzspg9s/ZdPe6vsZCUOEmS3+e9pdSjqhf
jsOtAFV0/Npw93VtnVqo+xJc7YKxGTGDmzb3o5Mi04CI6zjj3E4amxQtVf1KCzutOJI/E9FzOYbM
IaGrDyNcOr7/ctUw8vvh6VG2k4iy3M3kJCFhFHH23w96YhZB+5TIsrUVHdLgyC+zWg32yqXARcFq
B+Q2/ZEfYPQ1psB8Fgt/ZUbwO8lihX3bR+LuTfOUt1pHxkVPJ1GbBF8LXFrE8GEGgzcR6oVlKLe3
dmtHgPiTlLZFZHm+1Ps/QtugX5aOuEH8WEe8TCxg2LGOCQdEO6OGCZEedtNgP3HQUpP7T1ATMgjs
/sN/47c0IXkvqZucIR2nj652VfVniDwrorIl+jYz2JHLDSiigQBZ73GQv3ZIeY+SoGJlBQYYBhL8
xY0DU7CGpyjh4+RYr8O09TyRziYg65Ix+R/bSz0wPs9eNJ2K2FZgCbjMZQajoUF6v5OM5B4UzF9C
J1TQL0gNY+Ap5QCuJKdfubk3cGpFals0Ni0tANkdxGLVlPT/1lXJSqaBL4UhcbG120bQCPdZkmHY
TFwndD/lPJy5J/oXY6uo8MG8+XzV+7c3c7nDxkR31Sh6ROeRRXVkatbeLPCP6Iz5kSnJG00O+Gvh
UWKXnp5I+kojlJreNtHT6Gl1tTd+q4GHduX9iS/00mpzx2E8iU1WC9CiYA1J74duX0ZS7tlH6eqI
La2zIyIFOB4KX8aXM9ih38zS5+zepp0ADHjLa6muBtwTSN4Po8uNamzyXn3lT/lQZ/+AeqLF6y0b
pdAuUMib2j2n6OoWM7b3IAFNJP2zMDsixLIPXkHGpi5u4y8JJh9LnagKvMa6w4iGyQB6Cq+vhUCe
7Yj0oYtnzpgLSh7OdHaQnDNxMmct47mn484BHLR8Fcii1tyWznqBDRMEgnAQSwOJSKrxdLjjGEv7
Bbp+7ZPsj0DoSPmfdPHQEHibbWkLQNpHHNDw3gqbLIu0xkBO7L/nNexEHGGHlvSQD/nRbXfURH3M
cJftVhnoM7xvF/1sTBIwt+dY0sUm+HqGEXf89gQ1SHi/VpkiLkLRswKi1Yfg1AnJz6EOEcUkdvyh
aWK16hu2c0iTq0obXU9w0N5fifJod9b2xZFzV/+dQDm6ypNsuIn7ByZsZxJuJlaOUfTHzca/qXn4
6W0ohcSl/tTR7qDpCgmXMhGU45rhqYNJYXukrlZANWzOhtB2lExF5aclbyBsChMOZGEJyWJOvGNz
5NuVJlpbPkIiKJOxjtOwVmw+Bd+UgDlZxlUihmH4RT91CNUhWgnPELpK9paB+uVR+zdTfa8OEYgb
zLVxwaSfvjPLGZpy9VezbmDrx7E9bH/dKavgS2Igx+yU2u2zXpHZZhEc4fE0Xwg6gZlbe6R4xMmD
HedSA2PvpvzePR22yeQMQ2ec5lJ3+m4am/FrkcwXI3/hmSzXWcmTFzIvsYH4uRGPqmrw9mDqIBd7
xxBFskXsUVB5VGZKVEcikJS5pfpftx4ct+teavSec34nUUOcFZBW7sdk2W2GcTFoYnW9C+HfDqRR
zIYmLz4VBqyTncypDmLA43yT0iWO8afrDJWNMrQsq/wTkBTUA+EZ9al/qO/pFCNlis1N7nmb6chN
tH3f5/UfuN/UWMxW2n82gm6ykLYKWDKcOrtaZmrvMjs/LUHaMeHT0flY+aXbJ4IiOQjJ8G+8ptPI
kiwrhLK4aGKBkW3T390kZ4KoYAxJ3N5JlppWMjFFNoKOnJauGG9LC6QBLrNZmDRzRirhkiUu14Bv
sL14yXQKKv2Q0WWX3l4BskH5NO6GB3+jLlW2S7ne+3JYFTHNJYFPOi70Gaze4p7Le/HV6x+xg7PW
uC6VsbxWbKgeKBJtJmDBDBY2gk4Qud/bB8YUXOhCd4Jo7oGn4U7TnISWuWpYE9GCo3EO1aZQ3Hvy
RCHwcpBQlmeU9r7agS3VciD3lC8SFAKbzs11K2MDxUKJwNDU+GC47r35JSLLb0MgtKfeLC22vfyb
drCGR7hd9OHjKo3N8ZyN1WdnKVpTF170kqE3qW0pdl0jZNdd96PVDEu+g8Oa9BVsMzPg1rHX9pdy
h2Qw5MmBYe/CjZHJsu3KZ/NmCh8NzyG1ffpsPtlMez5DWRbfPecvH4hhnZEmmpWYbOi21YfmzT/n
35qMvVtlrGNwnMBpVLySdiAFWAKUeaSQeI8ZJj7gsrh7gU54MoFaUFHwHt2IRFW05DXrm0v5R20q
Xl1xCEXK5YllypaUGi6I2MGJL/wZxpOxtnFMh983qeHiTTp7CmNwytSuvnXgF8i+KEeaVWEEMAf7
LFnH1t2yQC2z4G6yt8E4HknmoTRndct3MyvuxybD+F4WMc4vY/ajHopKeIKIde3EZzZUvBKxcBoa
97VfQKNCuzC9B9MKfdSAUx4OpMO2fAfshLh3bt2NKBo8QVBHfg/hYp56xbz8UJvHi8PsKBIjZxm7
lw/adWVLs0k/pmr70STz8gV1Jcue9LdfH0XyHfAGRQuov3K70DWB0OwnMQdzmcW0fHj3ipP/zPGn
PVNEF3VqJUAzJx0jh2kZ37jBiUO/xVblssFe8cjClE3BfZHDb6/vpaKC71tqEcU0sjC1qD+FQ295
7qr7AuzM+1G2F4aa3KDEenSz3tasG4G0DDlv7MMWBrlU3/O1BVYN0YVdZXFpSOhpsufUrJYdKPLk
4RqV5/7qtZTXE1E1gJfGCb1MRm75vA6yzK+4OhANEZk+j3IQgjrOn0phYCTazmJItUBX934p09Us
RxZliKCFdRPkYd5w49pCpfyCKWsrklX+Yzbw+lJ5w/FTAwIc7tUzo3cT/IRPCdk6HgLcicy+kicg
VYeV45USNfX5Xd5cQdKTnsuJ46bnJg5dgeDFU4RaIfdUpoJ1hYWrdHxhuoxjlMf7Mlz7nw7pSiqw
NCE/gJCMs7r5jBoRsxdDrow4oJOAfhFdVALwxAafNgQNFGxxlEXK3TIt4KGZ+0xs/+C/w9COdnJd
JpeRbxqC9XVha6r6JDQNOu+MU+lgCW+tQjY8ZDFs+1D8tjW6NIGNmRj1IOpQaXq6sKK3l0EutGFY
qlts/z1638StNzw4I93xDQWSxusGOLBAzBG0ApkQqt9loUOiRK6SWXz5ypSAKlWJ9ZFm6e2DKEkh
vocnGaHzi7dYYe2ur9KiSi2eRKGmPd4Fd95GJknsgkvJUdlH4S/d/L2HiiUw/543aUSdfTBbAwa7
ssA81/fBnHAEhmoHOBLuf2rsoIdhBwGNbHHPtph98MgTerg3iruDFS/TpGKpKUUmi7Klp9betJnk
frHcjZVcBUdJw+TLiVRednwpzoabNZDNm1Uk3u65bEJeEae+lUukT7CouazZHUzIl8DYyEug/XW3
j/2rZ+PEHcuoQ3rZKjNzA3fk53SRkDQmo9K6oTJlGmZrspelrYgh7dkuopnBSlei5/kS1j7DLetG
yEwbz3qlT4cNe3ou2kuZ5mCkx0zBli/io7vesU4anIt4J+cTqIbQOrIcdnH+N2DIrps8tOvdj688
y7xtci+8FeFOswgS70ktV/Gethw2j2O4jRYRtJ3/KSFqL9GPSNUHkRsee+b7rKz03Df8Drbdx34y
GM+RuyNtAUqYrdRBt8sqbbhu94BX6B8j8cSDTud8psI95FPFfwK/94pej/1tXbh743jAl2hizEbG
vCkfg/vAT0h0elEIJVQwamSngJ8gXclCYEQyg3okH+ezNVbIlNrsbZqCP1as3fdEnAZp+CMmxvW6
JZDSFfNUueLoKUE/NtdOCkGuuaPXMIGBNQy+XAAelesKrAA3WO2Hrpa8ILghX3VTsRBch3MUxQ0i
sSWQ0iP8DSZegu0NbS7hZHNNqHewbuvPUfa3C+aoKhUKEKPsGkrRb40aX+jCg+r9hRwXVrQ8eXhW
rbRmXd5i5qhdGBqX80RJ1jw6pTiQG55lKmdW05GQXdrH6Ks2+IcxqGuJ690H6J4ZaAiPGD9AHQvd
lb9YSPEZcaZTWY81LOIYl47SU8r3+rBK0ZBl6s+UJOlMYkLimzIOgL8Th24Yh5dsJKqneXh8b4Ae
6pVZRjziCUIYVahDSIkwKMiogHBwyGV5CHdQgzp208vpIEBx39Ob+s2p2qIgASIwT4vxRHDW/Q8W
lOsSKWahdEkGaz9agjmbz7uPktNL3Rb7/6LAxdMy7lYHVudM9YuRXtgnV8a7QAsfUcPeg33+z2aX
i039X6i8tpSOcWNNRQwOVFJA5W0P1XL6Bs2sZiR0bxKNwD9PbC8D7k6Oav58KhcgN9JPe3rgXLNE
mae1b/3PAWPanPPJXnVLJcDh1c/c+4G4ReYUMtBkkpDBKpaXy9WQLvCg6TC3L3GyohbwZ+m0rjMN
N90nf6iTz5dcBS5s6S9RAxmOvNEnKdIevWQYSHRHv1j3BKj8rLmJtiu9yNkUFLJzngw33cgvO1ME
edWIhFexTSr/esKCibG8mP8lNN+wTtx1MgDtPJqOUPe76oDgrA2Jf8BJVCDkigmDabZ5xGn/zp8G
ZI5CdZOGkVU/N/0dTxRsojdd3eVdTTSth8+dLN/iFS4LmS5r3nETclQlll4DtlDA03vpNjD/LKVF
7RLo0h4X+UmonEo103jI9YxFOc04DHTLThZelu09Z22S6Y7Pr4XQUzYhsSSq5wgl57iotJQT3Xf0
6ahOKmlTWOInLxpIf/EeqXCXMFh+9JsMp5g8+1eiTSDOaaygRlNZ2HiNMbTnRwHBsdzskSwhhiJz
yIHwW/0LXnCTgqQgn6lddx7yqN1YTuD6kSbBz8ZG57thPOXtjcthqRjHao/wYQjIGQronzKegWjj
AKTKIV+1pT8/lXQoBWqXU8xPGJeRbFSK7nAUTBED44XA0fTLyvmEd7AbO0INGIelOWWoyxGPEAi/
e/DWisRZx54dJpDcwSUWRO9GwPvzVWlZySfQnZHPBHOS2WMOU2EqHN2V6ocxNo2//35NY3XGlfHY
/UEt1hcTCduX4FrA02yX4OUR+FDqpKbLSms6NsBeXarc1HVyYmsBVlPQJy7xK69t0TzZoNxntzVf
87gns31N3cW0mVysfkHYLy+BkLIBMCujkJoS82vtbyWiSTyK6dZ5RKMllEJJNN9wYNcoOGa+NuD9
dCIBavLY/Vrmq4ejrB3GwRRuefVxTz6lOO3yfuXOugoYZOS/UMMv2o2s48OGxg4bcl39E17JOoI4
f9a0ErQNPG0q0N/ozkB2N1ofE3QIJbccezERbgBsaMqXMfUYxTT39RcSc21rhGCb8zJlvU2qG2a2
iKkqGwik4gw0nTJ3mgxBg60fcEFzKc9w2ROyJvz+nsd/bw/34ehvrhs9JBiadVhx+wROjfLjmAIw
OSE5eq3sBJeWmO41R5HsDaq1G75cxCpxTJDAOFwgtEDjgJjFpwm3zcvfcDO7K5qcGmmEUd4Kzknc
tEsd2GqOGu8ElNLiDF44+6pnyukm5GLiMTXnjdZ3tVpT2EjfLTRS2WtKD4C/PRn4cdUVJAJtX+Tt
xPv6+2T9r+x0dMiXMtrnvqnZgiwM2nQPurnYOpfZ8bRfnip/58TgNZJSLjfZFPft/6L8MtyXicqS
VHpw/4G76pL4gNxZQJIfGqVTkvm7gTx6ZFmYdn7Z8hg6e0F6438xb3rvQTaG/Q4qLdJFC/2v2USJ
+u4kNLvCuiaKg2oMO1Wc1HXo0d8f04g/WTpZP2PMyh99T5aZrKOmP+mQmS9Zf468a4MFOOfYIqHk
hPQUe+hfBR6Ld224WrVpEEmYF48yWZByCop5vf04LCsiaYC9AHD1cjdiXUGarqcEiSkSWkKxIVbt
WVgSvLGAuBV4lAA2XdulPaDEowHUx/PHQcD+R1nhbwspxcSj7XAYknHRvjChVssQynW6Iug8V97K
LGDS3NshYcUa5zf0NjAwZopmFynGfp1PH7yqc+8Bq8e6n07YHtf/YYjYZ05u08N6NCZ5D+n3/BN6
uSGDGYvjsYoMJOg1RswD+ZP2TbAasCBsW7Bnuolok5VNAFSYbGOxMSWD0MuY0TRHvnpkCeQx4R72
9pQweE5NSRvAzTZcVAjcsFENGiJ5OLqTrQxkWNZZ5b1g3mbghijHD/AGOdcT3jqJq/MumAchWmB3
me9XjlRh4tkA4L5OrizINxMZBIN2qrhduVHChThGCZbes7FDSC/4k4Gq8/laNbFks7VfoqGU//bq
Y5Fj/usoDSiXS6NXzZfyKIoSiBKZ/ZyARRnvbfy2Fd+z6jpJ+v2VSxoybBHBf2Pt5rAm8+wqKRzQ
BMrX8xL6baRvqzWOy8WWIyU94GUINKxeGmdJr3Vo4QpiF0AIfLlUTPxj7Z6/xKutVc7xHbb9ddb+
wZy9lL0BDdQdKs+9u604lNlOxeyXiBHMPQzZ5wq7dIk1THZFfJ9E8iHv1A8f26nw2+j9jWM4nCCp
KnMRqVm+okoDQSBb6nXVjYQdFq8vXW2qeCC5+VjtgwRffO7LBBLP/30EzhqKcVX2wOXsxctOvfGd
7zbHFddnST9Nfdo2vB593ZQgcv2TxufWem5sNVZmxE+kWYfNnbOIIVy6kx1SV+qLrmUh9gHQlAB3
gBV8kvjWNjpLTnnwe/4c5ZwQgbEzDdlxH+cV6+wxaYSH+Pso3rFLYh+RoTxWq1mFtBYrmcNp9iuB
6aASe1fGNnsRADDr7n21xpYCnZ+IdT2+DjGJRJD6QL692HLBDNADseJTU4b88mpf4RSHJ1DzIJiK
kccBU3aZAaH01wVGxsmi7CSzx2z/7b9vsqx6Lfj9dgRCEIjmZfGAFlFJsvyval5oUS7ypbxP1TPh
ristNSM+sC6F30eOvqBEmBKRfLHJ2nLQMrQGrRZEKGgIppFGR6mnvMg7VaSf79cUhiH7ALjYAMNw
K1ksdnZQv2I/MlnoAWqUN1fZGvJSOu3GCoLanQbvsArQvvp5CX1SGQHTq5BaWAWJpXsQMqOW57ad
eEEvIzPQ2Pp7dirQXkctjIxRpQfIb8zx2QpCMJDKYi+PurFbzIqUF22Cswds1j/KIYapLWxfExwK
vJFlqfHhPVXP1oW3z+Jis2LSpIYhshLD8L/cC25v7W6Jrgbdl/5WOwrsSUx+hTZ149Pe33HJX1Ay
ZqqSsMkZLSLZr/+jjiVAMdlSRCuUFc5KJX4EsOQKtqfkS96xGEjwkw5Fl/mtbaf2HZS5R1xwdwPo
U7fEFpLqNC2OapnTE6Y/IU3e1Ek/j5UMtvIvMxb0TKhMYL+OCfLqrou8zxiD4/YOfAf5S3XlVbXW
A3NCHNVaQDlUlJOJN98gN900G7W4hQwdjajmLKycf8Yj8Z3WOykjAQhz4qvL8RLx/JpgXAzeSk0p
826+1IB3SSNSDdK1Rkgmc0Fi1AKYgGgsW+M+Rn5adwBVc2dvjtVnFm8hbjmuAqrAplQuG9prYHav
3BAlkE8wVgZ6ZhRfYaUz0Wgh2QWmdtMMNltt9yFNvic4gEBFVTld5pjtaWKBaboeZq+pExcZCuHS
bBhxruFoeY84PA9lKxfb4mBlcgw7ruSrgY7BGeUqmGH+s6BsvtnbY/13Yo83+6fszYA/NlA0Lndw
vPIo2IhpHuD6y71wDFHv0ZKS4mtSRBk1tkAfX29ADIXmtNlCTLdKZF8WcSfhdDfHu1cC8HOAfQcT
kZopSh5bQdVwuT/8xjVZrjLGqkq9QkFzDDRJ5hILYQzaVBFShY9GEt/w4lL3oLsZHXhDI+3Qdcjf
2TM83MV3ofjeEbi3DW0bxDwlmahGTq4TGLuambCO37U1JKyWAhAJEHKrAaWDCCqEXLbPYJ5NJApO
ZaD+qIo6g8bntjhPZJIb/2BwIULWJRExDY0TxTWWxQc4u15nT+2kTqEJnSsXJQNSjsVeKyvK16th
VgRpWJ/Np59iR0t4+OEmcGoeyH+GfZrYchjB7GMZdqq6FMmirzpdx7aXW9a3HWeAVEbNa9udHFr6
61DqWdvuSgEq5rbDOKIUjcpF8wZnNt1f9Dt98dijKSyTU1m6LG/QfHP+eSVbAJ7v3ToZGTvdmNGS
vtRZMy4ExiUNMYqe7oLlRWUoafBTAgjF1ti4lKfIOdb0NcYVJ+j1NAN6GUdKo0dLhvx38XPXOERE
1CID58Ghdg+Uhf5XOQ7V/piYb9oyR015QXjbRaNZ5mqLpz8CX/P/VxIGGeY0PiUlVv3XmKJFTsRb
/Qpvimn0aAES0bFoBRgWATkEwbe2aGYiyDTba7PqJXgRG/laQZ2kx/FLZm14+qwonOMuGDEACXTu
EV+vl2QQUte0EY6YBasStBWy+M/aw/CA/MtZowedSFb3uJjhVmPbtToniuRInLc8889VMH9BotGZ
xOPp+7a1YtTLUIsQ9LMmvHZxivBp2uA9GhZJLLrMyIKC2+u51cKWstUSJkSlFUvYuv1POTuFfcSv
wc+i6t6eUTdo0+fuNkKIpEvf4FL1Kc3Ff/ASHstl+nPq02RRk04pSCvqJ55FaPD/6Ij3t+O/xf0k
2kwUES5vWaVhKYw1nNsmuDjA0W4n9Ro79OBCPjySpY8rtQLW0O9rkLckBRe1AsBbt9kvJ+gnvQyv
aMueAxivCzPJSccaGIp3E+2HEIrb6w7hYvJlPPvm+3gG7DduuueuSCslYKkT0BudkaS+77I/ZiQd
LK0tBCDoJT1ODcJiOtBDY0heZCVccH+RrXXCVkewvtEU3D2Ky8pmRAMdC1mNqcJEo60FdDvuWDYZ
QvF1aKTajFRD9CrQhQ9Pqzc+QV9Vf2ZH4zlFvsL2Ma1MMMeOw8NMuWnyTOAV1RqV4b4TRpIjUboC
N72z8QWXfIVfGNVq3oRNDdap1TEb9yR/yyFrjH5iPezG0GXaDaG/ak/kBX8xVa7merWkAhpbrlJZ
V6/2h71BD6ZJ5S/yhVhfvclzvzQT29cAGcIw9F4XhoQpzdfsIdN2d0cWEItWTGGBJnSYFmGzri2M
oxTnCBJznCAGm+mcWxnaf2+dxY+wJZuYwMLdBICmsV21krAv1w57ibGdJknnCWKRdPtjDBWuiXZU
8qAAYKcqxtYD5OdqfJC/FMGio4/KOJbxatkhSXakSibq2o7/GtdXxAjQkE9SkJIeaskcSKUVudwn
8jlF/5vn08vwafrL09d1ZEy+tHUdQw3i55DysK/Z4xnzI7PoLwz5uKeljxApuBtv00//dKdBF/+o
g3hDYTUIg0pCLVrVVbs6pgac4yxToQj53GPdy3raqZhLHncFJE9dISWihHAavY9mga7YT9Dmricf
2kKlrcRKeLjbx8wAbkpClArRglS0iksa5L2bzzxLo+WUm3Ggb8XA3xOVi8m6odRqBEvINl/s9tAG
drzya6HU+NfLAzhbcr7ac8B22UQ7eT+ZHQaBGENn+Qr9tmqjUbtwMroNQLLMkmPIUEwP7QK0zcTH
5MSxcG6yZMlABDMuhQE9Fuh6EH9l1Te/UmPC3hKiE+oCKE5kbMzw31mIiRR7hwqdRG2O8cADrWkJ
m05W2UVQwZ4HuX+ypw6pMjua1o7r2gbr7tsAAyvW6JJlGr4cUFT8i6+DgrjCgX92fb/yAKU8t1/O
+UNT3WN6o4jziX9ZMUdZnNtRMFRcs0nC44YXDv8f7UxU752EiDe+buWlQiYukj8nueeX9SvXPTxP
jrbaKr90w3OzAQUktZkxrrnj5kRVXjIWmnqoIKLkhCCxMpgNwZZuE9keqhiwpQCYf4GpYuro04HM
R+8K6kqIyqbxYJ6bpPqLLsz4I93RB1Sll2fCDPxWqa4kiBYBkfw6rZRVZ84rDNbXI+25UFdWOEBQ
w3aEcrd+U/5V6qscX4HjjLvl1wjohlavAuxYGBb5dCuGqYZYA3fYdOROKwSPnvPGOyXi7WJKYEDG
A8TQVNvnBwnL3OXUOqYcU4oFfOPHAUs3xcfhQzbPBJLdUZLrbh8Udt3gBH4AsgqX4SMtwwoEtoa0
s9vv0lMBjTZd7YHd8M8jXlGS9cVCyVAohfBafGhIQjSSbCLqf+3RhLeeR7i6dEXnnCBBXBgA8bHl
52qQZDem4KEdOnbEjg0CKD+aHkBWD8fgNuvXcTuGMZ8mzY+6M8x/m1Mcj0+G0+DNHxDoB7o9q1Mz
kjj+OxeY4YIl83mRmi+tl+P0kVyROsniyrT5pN+sky1rPQkhpV77b+DpCmPSLq5or9/aDYBtF+Pe
or1aF4Zg8+pLw8aO7S5Fkf3QwyYX0oLEaOWCjFJdry8EPYwA1vaXlIXeE8njSlcWlGzXx8Hy11u2
9Qobm1GJ3nuGIv2z9sj2UrS5zPqhk8ApEQ6X3nYGWBpsXrreK++qWRrtNGzONaLfvJlOG4YLUQQp
xY6T4j0WTivNOpV+y0BhK9DcKoP5ijl7i7nrTKbdkNM5GPtu8GC5OJgPFA1a1RdpkKwFTtV5gH6q
8plITIjvKBNIw4R6DW1U1CliKmjowJNmb+fl7B2vvlpqsyPTOdAj6VRhnbwk2m0bGghn/ZB6mN1K
AsOMGcu7BHIwfLboNLNuSEzGcISPgGBhM9/Yj2D3E4K183Cp7ex50AjbF1U+aEHX3HUNASAZaSyj
21kvti5ah2wtK9oIkeHorEklWElxUPMtJiFU9QFZgRt6dL75Lprw1O0QYbTOCGgzW4UAYOl9ducX
xxH1AUli5RCfetiMeHElPr6DlNHT7MSTYTJmHLsv4ezWpG59BCyIfWd/MWH0OFvQnt0oe9517ucl
xVQIn8pQI0KrHmdWNMJsHGkgWRiXUR3s0n4vH8FAQEoulzrfTkS8CHznerii1Vi6fUpuleUGjVVf
iq6JA6hRFC/TqRYc8ySeshtHLZflLeP5Z8XvVzUFz59QQeewJVQYZuOjm8jYND3HD4mpFtmLIq6m
Ww6gK2FJy4DzbR0jmlIJ03mNMZekz/ulzg76MLNVIkHvyTeRY1lPqzNYX2Qht0KIWz+n+CO4U7TN
NecbW6KWkm1/iPEGPM4fzAf1FjDsOyinnEsd/iSuXpUqJiInb2l21Ui3UZRIWnoCuYZv5uGrp2mE
Thge9I5kj0u4kmr/lwzJnuUmXDP67Vp1JwkR3vVvtLGhPNUy4EHOvjr1SZmAthbWzVPwLC5X8CiV
OIUKEgCxF2rJTnwDA36s+7+h+ye6d0zMMhthOPrbwnjy9WFDDAl27vI7wGZ0BlWO3dpX7hxhfzDc
2F0Rko9xNeGJhqYy36HrD2tA/0mEIJYZ750j0YgcmubjQWNIG3SsulXIK8XrJpk1ZG6BMonMX7gL
kUet4sdwvn/wFxyirY1hFMBZ32aeVZboGDBCfzTWTNyyncLIjnhE7HvWz92T9Wi1OymcMOGZer/U
YFruVYQyEDlAPwDe63vg/XQLfl8AVQIL3M7xAV1FUJA+oaSdqgrpN5ZLa7FOIh1+UNSqv4w+5eCO
bdMAr9XiJbYNaleq5Uv+WDMDhGBPACdROVY7HYN+v/GWjavwIzYXZDbKyUdtI3rvFyRTFpsjOr4D
eznw2cegtZfLQ+zBdjodpgD7oawWyLUzuP4ASwklbqMgypnKTQK16tC5jbcIKmuoRtJmMa64WQpW
mRHGjIdVBNi6EZQbjklagSlVIBY2f31jnQCRLlpdiFGD2SNKG4Bo9CX+Nh3lOenlQHD4/zZuPpFX
jUk7UnRkIsVuItHawINSeyqjzrBfvNQS5/ZIXg4vTK7uZRDTgXR/5PRtafKFVCL1nSJGfbzMU6n7
avsqOqSqj4lW7aBEDH0HDoFB7PWy+9qxbdM2NeENo0k71QoADVU4XlA48bCxHRdl6KX2AHJJMpHy
v/pU6KIAUhshL4uDFcWwpLpZ/cx2Z/j5wiChdl0HZba5ZnXeqVQTS1wGnoAPndpxggWqeqBpCKfy
JutSD+7ci+mw9TZSrYSRzGU2R4tObiFDzSICCK73OR4pZjPT5E750rVRWmjtyB6Dx3AreB2pGrQ8
7/sLn2q7Mrq40ydYS6ahZ0AS61cTfm0rC2PqMMuFx3gfSqXTTIBvv/ou0NoZqsCxSXz24Kp4y2ki
TeGQ0exR2lBm2HRJoUK7Y2k2ayDBNpOS3gtvPDdeTpPRxUfOmeoHghetW8Dp1ZpGSu46g+mGqEFt
yU6/ZmQ5alL2uvzRQi1WeozuSfIhatjOJeoOBAYe+5yrZkvzvJ9MxtaExr3x75ogvLE4+LbmNzS9
rJbG6FnAS+kXBiz9BZrmMLoB8bnGk162bUZsb6BZ0CX3OjBpDdcxXtFmB4hjjWE6utjG6i3ZF/Fq
hTjjHjgqulMCbOgQDco5V1aXN8H+dgCbcV4++p2FaMifAPkQYzEq6BbG2/FMWqqLS5hDn4HzEuIJ
rX9fclAAsABspv6A4ZXP70Ymfu2FZxsGIF64oOOZ5Fj+A9xEFRtfzoCiPFw2DWHcWYfPSl1f0NQx
yoOzXk+/jRUe4Wn06A9YG6IYyZdc91MrPv08v/1b/RDwVmrAeVnTtuEqn7RrmKt6U9H3X6xR2XOu
jCvOuIMcXikakKpU6npkcI0a78g3gI52kRH5+++GiAMSMsjrRkYazsJIQ1qBuo0SUA9zY0eDYNtm
0Ze+iim89kIzg7ckReaKPHJwBDHWmKauMRZL5dashgzHZstpTLAEMXtfn5cH5QOmENmgH6EqNMeq
DLRPf3QjlqfRAasK9xR/j4TUoOTtorhhCA8RJ5uURU5MgMVp9svmybEuGlsTHfK7Ijx8J6Pi5eT7
21cCwbAlNqS3huRo8hC099x2bKb3e5vhGRBfWZdthQDDETqlLmWZ63XG0ADl/ZeWv4ysoWh6QaFQ
YRwFdShavmgq1WaBwOGwo66vQWD6GHJ4nPuQ5ImcM6cDsUPEY2ncn+8qbrp5fAl7Jm3DLYQ/TfiP
rI7NkCvKiqb4alK+KU4eQ6FXWfk2CKW7p1v37hSJDQ74h6FkMHmw1lbfcqvQO9inOQE+DKOv93zi
QKLe9HeYw8WZqeVmU+zmmktE9nKdXRFty2SQY/Hzz63Y7sgwYjXFPbz2+PY+G89EaS41jjJ+NcXe
Hw8FrKrYBr/ZxQr/4Q4teyTUP8Gkqj2T18av35HPmylv9Yq6qTj4x2OFD8Tb4PvNFyKwPda9ZfUa
3XEGZLpHIWM31Olcl4qO8wEYJzBx5f0O1rqr8meefEIGTYC2vQyEWq3mo9KZzQdx6hsqMzgPSc7T
RaGt09s/mjnJSvyN2ALIl88hag1WQEzf5y9h8fLyu4VQPY8N7lc9iccyEj31VhogTWGLZw1aiygQ
6s+84zOwoKLpHkRZKHVViMWdhk+DjhYbdEIOh0obc5hm26g90jkuPQd5NsMntH8niVNXCMFW0odJ
fzRnEzcBf+ukUpGZVlG/d453du8xKruaomf+8W/qT2jqC+r5y+eYH7URQDdCVncZ0qkV1LKTDK2t
IjdruEvFHM+Pk1TabNjllpAH9wEZ8Uzl0qNlV5AX173pSDTGs96/JtZbENDqkW57sc4YCfZM6PaX
hLFpnXWMC+sa+gX6azzVzuJpWR9Z+0VsGAfJkhPc/ZkotQO+gCij6rl7RypPONGExYnTBT5l5DpM
yqy8xotZNssua3RZrfJ7YIZWBc72YlT6AknfZiX80x7t6ZZbeRkAMaC1YKypAEPZAITr0+/jLUjv
dvnXmXUgznrfZrRFTTh8FRaN9GzbV45sxDH0RSDS4hcAjjtlViUhhJVAvld7mhkd/bJDWXI0spH2
j6jldVjXtlUNg4NY+O77gDkFjkHXCpDR7IiBHYhZ9tq4figsxG1PJL5oOvFMRpLsMW7l2UNIc8/i
FVhChEy7AAPgVubVAvo7UXA9f0WuCUxs4+oysL5z8D1zz10v3eoZgGQZZ/v5H3lUSXbC/I7thUL3
j+u/plALNfRIZwHlyc17oh1al3+phY09YEKqo3swsqp4AnH68Kx/oXhjKT/bB61rDRLo0WFUPMQ5
1uxWZDTCeAt+OiylYnrfUzHeg8tjc+YCo76OEcWjB2V4y8bFXX5eothu9EeN0lyA+99WsqtrLIu1
KzwnA/yEouOr3+0fYM0Ru9mLuojC9kYz7x+zfZZoKd44+c6mXgRiR19+byjaXdgiRRvKcP3W8C5p
sA264KKY4hgHFWF6VFo1OF0dm8AsfDgbVdDsDBZ5IXwpwUdeX/QO7jwICJ8E36zmv1VUjVMzSIvY
rtGrLEUIkIUKT384dEC/6m4+Rvx2dzhGv9dWMeu441yHEDyVkIrKgJWmzbWsZc4xvb0J0mhlrGsq
xndAk7QXG3Wm+wPEGCWGHQmBRj9hflsJzWcTvMiX7vYSXaGCzgkzHo6syYdyL4+AB9CpSDXuaP8a
MY2niX8Ae82Pj7syxzJaiEys5MUB+WozSLD4YrBiamVpCU3oiZhY6Cvlby9emO9iWMR2nhWDzoNH
vgumXk5cwLkb6G5DdgBcnC67E2bxEkFK3qT9BqR9WnWigAhtAB4e8kjWEDLfZR61eiDh1DY69PIy
kGXZ6ayEeYxSTEWeh8nY94W6Id5K+txBpcV7CZ6u+k6KVUuaV6D8MDCiko/c9eBECCyK1bIGWmhj
DcSVg8wSrvmKBtPGigax9ogshVwUzWeDjVHF1BJ45jPCTEp17ZGyaMNjxOiFEkyfPRWuTWgfz4ID
cAbiLMBGfIoCrnZgYwGDk2P7wphrQ5nLTZSPxPxdio4PUfBEhI6cbGtfhNdS8a6Yunu0avYmenbT
cz57Bhu0HagtAhDii7lHe9B1IyEEq0mfLlVT0doShuk/iXDYBgh5vN/8/NN4RisQhycRCQ9NVhfO
UxFdRIhNBaRAw5pC4JzoJm7+Q5I1wFa6VhN88tnAwFk4kIeAS+dbGVm3rwCSjThTsgWMi9VdUzcD
RnTG10ii/ORwU9oGSPPunaSJSlpZg9N5TDKpgHT283oHtyIPzIl5eJ1wd9KZ66dyDAqtN4TSuehB
DW7GFPXxeQCYy+doXZDcl+TVvZGo8sBxZOPlSrntgA3IbB0odIICx1XNGW/MBGhwwJ6Jg4CyXSXC
DUl7YXdVvF/9CPxkxUSQLyXcUrUg/Q8SAQ7VXtB+UPuJNqBbADr75cREWlkmvsqYOQzKjVnWC7or
l5UX65siDmH+QwJDrL8HaI4WpSkCjrGRjobi8aBkOnpGgEYNtWM6EhvW8+OeW2HmXMg0Z3c1VRtz
GgdDdg6AILZAdwiybuhGpl1MQ6Zw1SuRx1xsD0TfVYXAPxEQWsxYBVyHIsIuK3cvs1UJum/Qmr+Z
eBPSZCSSai87vEC4iw/64pndQU3Wgf7XOP7RTqcFlLKhciE2QksrM+Svu4WQtxM4Yd10tbmKgVB9
k0eIaUAXwcR8P2esjm61qLs4awdHbqv8OqiSuwQon7+pwLYWmdqodBVSwTl45Hl9lHBi5/boLmpt
4MAlXG+4slupLPeD6GUVOz/VQcuSAjx8XLKPHcqp0VD+zUiWMDaoFxRf7bZjzv9gMGuaYUQT5iI7
8vzYdKKsvHUbEzNneleymXIAK3QxlnAOtJUSwVXbP0Gtod4ymQQPecEwkL2cGgXvcjhvL6YGiR4P
i7JIHc1Ov/NrsWwoVqtfwZDEPFsu0bPlnfbbqdodUv1m0S6Omer4y79d/2EPcfeZVol69cxVBfn8
BrWKkUjr4CTyY0o6N7Q0pmDMjmlD2Dt+s2T3XzXYTsTVhH590F2KydPSItJl1MBEjL9eZ2oNVk7W
U0MjqNEGlE/xVKeINPQlDAwqenruhKW138C/pDxZMPBeBvtIatpVXdJsN5PjwMPQwl4QdPTOwSjU
xfE9bp+rYx6SaBH2zmRXS3Lu1QH1iXYo/581XNdcmxJKHmrPwpmbubCYGwzVF0RkEWvJLRLbf76v
i9Gv19/VkpRhoQE+0b0KXmSDt1ZPL1nl9Gp5yiahVGpzwHuZKILO8u46LOdEEjzPRy6ukgruSfsY
S+TFVR3+oriIGV4EVP1w3r86yTB/RVGPgA5QpK8VHuaZ/VhovXVWPH+cejJoarEp3KpUdAx+GMPT
sTvNIgIgUr+1xam+ZlVBD7IVqBxfFykcVWazlu5JGzzIWMy7onzcXZPNC7Yspk9ZPYQ4DznuZ9r9
GsjkWqyOB7tpNFO9FKkidIgzDT4SIq0Iy+LWpIqdJWqYCPEiEBBblryonMqRl36vTpsdHUsc42sP
QY7LcF0xXeIVXzlFb9X3eUOvbU4fwlZsvRpIraeluIpDLyRbQNSzSLu5K/TbkN6hPrBBFzOBZAE7
TFJkMclshXnrKu2Yf98l41duBCaPbqif+Hkz19w2nC55lT7a88PMXjMXcvJvj1SEnLX2WtML3Wz2
6srkphn8GR006yWW2DxjMH8/cpoAHFlFCR1WiTGVhMCoU0UrzyLZx6Bn6pGaH8R2uKI0FV40wwty
IV3M5n3U7LiEJJ8/PIGdRoT7K3ygYiuVA6LqPAzvFoy+XTZFfoE720LntHskrb/IOV2hEtlnSDKB
MwISAnYXJ7e9aXhaN3dQBCq2YVz4uhru+yGc/vwt/ElYX3+69Ok9u5CqFSUZBECt+JS6M7M1Rcx+
9dl0t/GhndZ98mPi1oVoywwfCft9wRfVX6YqFK+ftkn6597odhPb697hW/IZSroKft+IufeA0lyz
9EuFgJBw0d1fK30itvw/lSAuIJgDyGG4mGF+IIflBeoPvm+6JUCZYjjiUwTcRrbdl6ohps7etaaw
c8z1kT+oZJagHiCEov0nXvHYSH2QcmI3leBhuiNEOZsGrra/BDnaCU49Nau9h7vahYiagjZhIUgq
Zd1+Al0/E7Yu5iQxYmJ5T81sjiuaz2Zja7IK2q9qa3c5y/nrFUZR5oadLE9OnSZEvulagQiLXi32
SoHR5RiNFYZ4bESmbQyTMGXGTTz4sTSWKgkpnbcAo5D/ZuFsckTOB9onHuOtbqwCjLvqNVm1ixdd
yY03SmVkpxd3PntbhXKh81jMZByfHXxkoXAo8/0I6QOEz59e5hyMWqHpF4yq31VMeVtJLCLyw41V
EvdHSfMEVMxQDVv1NZ8FJSn0qjEFkNPITguQGSR6XTSMImYjUQP8fRCbc8hdYUHISkyfiFhYHG2I
god5xS1niELNxHDwqWgwnlyCXTGmtxzrm3UiK6xjRetOehJKrcyB/AURkH5/9O1a/Qc+fUxFRsMR
8JKO2fCjCC9qe1B3VWvALTA+/U0vpnkVIXF+5rX2uRlK++XEILa85SNEPIoX4qrvk0pkN/B1pUaG
d0GRIMdyalaNVkg8o2S0ufpOjVmVirnUUI4yagN7jRIeIrI1y2Jt0YMsFfPY7qJ1/FfT8474ga0m
F7PcafhtfLDQbqYtG4oA61YFIaW5eHCgZupHZZDWVbQnJsMMq0bJD5EP1S6Tx92RCxy+Uv4n784/
T8oSdjPjBDk5fDQhdHSWsedldAWJr0E+ggvVjGuQALDeCWkBR5fjrEQQM0D45k45dPxbKLvtR8JS
AYbSHDtDypaEzLcK3miEE5MM9YuFMrT7SpQduHiYKyfEo4kL+iDJQKoDqcwEqMzPm9pxs9TFaloY
i353jo5ZndcgjRX5Ykq7aSm4gT4HOrT7vcO9nxXp2L2YDvj3W8Xnjy4MVcSxEkx3ZqSvLn/k/Mr3
bJc+N83SBZFt+G6rEIf8UNOG5t5nYJ6MwknB870RMEB7rOEL7fIFes8BbEYcXCmKkunT1OhzR3a/
llaJdageOfW6LRG+VMOWnnCMJJCt5l4gqfqCry/b6extGDXukkBYca05s2zUj9WVCFALd93+MAbn
LXM82zgCXpr/Y7ZZVMTW1RnO2OeOfbBj6lEr7npGyriCLulQLEH1hxlidb+rbfiFUIckR24PuoN7
iiAv/Upx8sfphREWmWHbVbHFaFBRrDiMIPnMUMxRb5Z2FD8dHkvyHG4Uu36cC6XOZktTDm5a7+Yq
aLqJ1dyXUcDXKxZLhrV08kdBZE8/UnwRNIr+zlqEUYgUvp3vQUcD88HIHAbgD4V+t1cnXdiX3goj
ml4JnWF4mXVTNM+diGHisRySE+XGxpONx5+yrabRzZIp9TmvVlTzqaSaulL/Aszd/W0E0snQZmXF
qdAI0lImP09pkyTiU3CCTeCVmALfX4Kt4IYbxocu7jlRn5wteCBpvYb+J8pQcrCuFyu+1+/i6xnR
ZYgYdUaQWiyh8+heobAsx9SJqltzVwh+lWMA6aOsPWVXgTQDTJoGSGY4Ua44K1j+IaVEpr0NTBm0
rtANpUGW+gSOa9lwOHjh50r8Ts0Kil8SIr0VRbfJyfBuyVGMdYHLAZjW64kMOeMfl4iRqZc5C/f1
BI7T97VHOkajhRa+w3UkNlUYzd2lQrBLTpWhMM83rB4Rpx77xMiOoTvwoQ3dyWmZcGzfm1/Fn/Pp
cdmZ20Ft1/2Awm7V02UpmoT43uJcglkbXReFTQUhCfXwNVdupluO5vIAZkdK3gSG2lGB/UtPBfHG
JQnoI0NFTbzt7n+PDGtL/CweV5CmrRiJVaSV/dE1x/l1iRTL5xv/zFzf9QW9NK+1bXacVT94ObkL
sr0RNpeEkiYwIGFzl89timkhjQmu/6rnreQZYPWzLGGgoJUQKTvOI3+YBMPeB+FHzJYo36PiAzKU
Vm8sU5pl7zutrBQHyLTpsPsey5GWo61J6PjMg+VW+V2tReoCEUA0yXHwKOyR2yfcrNHNzBAVSXM1
FeEjKuCILkea5PxeMC4B1ftDqaYt3zdic8hjlmzuDYaFBM18muWjyRCubkkwHasZOozC295sXAoF
HLWYay1AkHbVMQsoCGDkosa1p+Uk3J/IhzxD/ZvWzHGlHoLu5HNuccmdSPO9emo4Q7CpyaUGJ5Jz
p3k8RFW8vftb2HhYxVfGrI2Lq0jQGrUbZ+scKcfbi3cCl9zj8lkjRrXoDi7MtavgggXPH5s5348X
nxPY0pQ7nW1gWbBol+x2TkyajWqBTnJqHFGG0Z53vZ/46eVih3AK1m4f+G3Mr2TLIc70iCfMJxeD
iVEmj1+SFOf4vLusJ+hOqHzdhbyfEYDwu3ugJyipbQZuWLyKsR3SeEevORm+2eJ03jo0Ks9eHci+
hYVOoZ4pPE7US+TtQHycebo2d6/0BX38Y/pTa5O1WI9LGHsoQfjQKGcbP/2d1Z6zobJoR6HNHY3u
LCEsZZm9P3A7uP184U7G6xkF4L7ojdKEocZZMMqsVS7s2kEECZcE+dfVlsaDS1OIC1UwEJMqQvQI
z5GyK/roZlh7HSXUT5x0Xo2yU0W5aQ+VHuB4e1irrWaXzCE7i+UKEI1Fr4nrbNbhgSry1AnYTjLS
SmWnkPn/914tQZbVZkMO4w7VrcVLlvVA0xmnxUSu8cSC6vq1eXOBIqRDSICKAIOrFVdJXbMBShl2
/FLQI/TKvn/rfW0pjk6Vls9l1Vt/zbwyY/a0ES50psePufA04nLkhpXF1paUFvEh5ND9RZOSIB+W
foRW/GNO2TAucsgFm+7eW+atKUVi+K9Nr3P5wc6ReeguhQZHapaX0pq2A/sl0QNkYTH+DnC3gtvy
LY2aZXrtLmKHyREFoM84+SpxQPom8su2Pj6zbFqYeKFQ69hbv3L2JGqVQwpSsB4eE5epCHefyjAC
6k6lgG0eOEX+1bnZiebycQD8nGqfsb9ZIR+s7CjecwQP04Rg3hdp3klkZQuyRy6c64jsXIn1d9hq
+H5dutvfzGb/nKIscyZyJscvp1sMCvBn/nOPx6ffrN9z/SG4ICvTy0MpvqdM6Zg8ksJH540aHCTE
a/g0aMzIiUEout7fpQpfTnvct2IgRKnjPXuXY54SM4joMkMFvk2EgDvVHEtP3v6N7nVL0sy7IW5+
Lxp/lUOwcNEII+ifi+pcWz54/Ua12X6+J67EZoN/S3R6966lokJDWcch1LoBH62vdsULWg/I2ngl
WSQbr48suDD+SnlUDhOlVF9gbiI9P7DEobyqaz7DCZ7r4gSVrhpTomFK4Z3ByM/pUE4OsNc0dEww
RTBpycvkroaTBCU2pW5AckUrznOGkTD/1HuepMEgbnmHWqjyGwfFuL2QeWUxeDidwbr1aR+2lN7n
ovGmERRCtr9AJ3ki1eFk14E5mBtvDTVR6mjDOj93lhHpvEU4t0SIs+n/msjQYlx0spbJQsVbk/d2
qcDTHU7V1CQ6Rb2/1HkAgvD4JhUcTk78m9Z93H600SWNS5KGqHl8JIDyWuEqzr4JGQpO2C3id2FK
EcCqaNrsZEdIgaT/xOKVdMGPtQxU7/g6ccueWau0zEFoMDrXGTxvZ7knX/mNQ0YbRDQRukOZrpT3
e9YGE1HOuXXd533mt51BY3D/rOXNRkHa9Uzbo6bZz8+2Xgeae0tBt1e7KJwvMT5IosxWDG6xADVp
A2k06Gv/1QxMekcT2pPH2h+6TlG2LkNBt/NHif91vRQMLELMsBOkUDv2blJtXQwnVZpt7qv9K+0g
eJUPE6222yhhmBpcApHKVCDQRIrXiJagqoBBsU8Jyb8WmQPjC07AsGS05VmPl1LR5FRiSSksMtF5
SL1Q1yu9rcesmZY5OtNTRgiQei70omCqPvPGKU/fARl4dv2rpRZOqtVRDUkCp3wULRchof7YYnaZ
EmtwveBcB/H7aFUsByImtfrWemVf0PTfh07vBkHIp+5yP9hpdlP2lsMdcuPQb2ZzF70X7PZeUa/y
oczQ7ItnPxAsFFIGC7u4VBftlBx1DxFB++h4g9cj52LhW6uJ+4R/bVfUtv5EHTp043LwN12kpIcQ
YrjKyEnYStgCQg4equ+WfHNBxeG156KiffQJo5m5ELRL1SvuXQSDIeTFN4W0zEYn3c3xPtMkPmTY
XZC/Txk4OnO+rk3zKkiwUoF0m1/2Jq/8kNnGUagI07IRUU8J1n3dJQKzFWhI5SQ/781DzMDKS8is
hHtVfOP43gt4oxClY7LBr1D9cfQtA6WwrwHSm0LZM9Prue4ccfuX3W5LmJNCR0W7abTGtIwpLw3J
XZp5ERZP7BGEh1Ru/Wu8YsMoiQSXt3Hj0Yo9FP81KBUnTsR1YubNdVLEjVL0OAgg9LmCnpe62OQ+
o2Uaafx9UmYxza3QFOSVABLNrAizVYcmqVYBl4FVEGiIIYKQXSLV2Jw4GDptzjazsgsgfNpwCmQO
NgZ4iQX5u7XP+MgM8NE4qYhoQdsZySecN6yFdhble7QfNTiTicATW6gjKxVYF7a8PKKc2WY72yXe
US70c4hM7JoQ3uikog8p4RW89hD/oUbFpROSzQqioV7ErneaFylfvADgnmHIUyUj4y4i7jrTsOIN
HAQkou1gZvHCAV1xHgeNFBakG/UKOGcmTeNZ1rbgwxogF7IP5fJpFEYwh0wxUpBK2jqw+Qplup1s
AHhB8384nUNzmqMPTkJ6r1TPvKRPou10BWP0J76vDrJ4/RFoozBXHjR4/7t+T5nY7+o041GTqCTN
fWqJ5RE6zRow1Da+xzuIj8Ur2jvCjQ7Z+jWgapSLPeQ/McvFYmgruZi4tqlItlCAw4C+Keb/qiXy
O9E495rsjdYiz0bVChSeQ7HHGAGEA1bd8X8ROeSKUm7dYcVt6TLa8edKvAsRRoQPxGeWjw4ABEtB
scv+h8h4AvGNwGYUhg1q/gcr88RRMUmo9JFLv8YV3eidN/dEvw9nZhX4dfh0BnEs+ZzUD2gBbKnr
q2WpI8nXiiIDjYb7BYcKAg3XaAAjdE4JJzRg6xyWN4RQu2lKdYLynVxGOVgciDTXSllexxvtTAMW
yUSQXaAIy2yPrKPz4pfUyTU7Y5P6AnqCFiuXx6+lCdTuxAapzLTXyLkSdhYhlSgepYMKvyL1MUJN
qur/eP5kx70dMUyUDkEKHDxkRd9OPGTNuppolDekfh+r/pyZJPiDJNuW2R7tsM+VdUaRjZNvjHnG
v/qof0eTUlt4tMlbzLE/m26F2pR9vQd0PPstl/Z4WEd7cNdwhoucjVpYLMhegJW0xCrECGFOU2Ik
Skk+c6jDLGTwZWG0+sdjAzj35cNDxA9+NV8fUod6+MCU3f420Y3zLBUx5tLZNClN4ICgWMubGjh+
1q8Dzg1/dw10r0pXfy/OO0UWz9wNdkLrW1qArdb4+CIj/OIiZ7v10Bed5R0wQpsA5PFdhC4PV0M/
oAi4vItzJ8sm3L7VpBuotEWmIznc8D5cpLFVGpHur73YtwuD01hXViCyGQYOXHX4L5K9a3qqqhhS
muRdimrsGM/OQtyI/vS1KQDXLxs611YR1ddXKfJfxGzFGSNOnRTgUMOqLIMXA6QM8ihg3/DQah0X
/qcSGONchLxqcRF8wGB7b+HMeOGYFb9PnP+mLNZmw05A5z3NPZJakpV51bV/Sb5vHlPIEIFsT2UJ
EfGW+p/PkD4V9Ki+wSjbqVdmQdC0lDrC6tqXFG1xBaIdy1tw7UOOZwuOZnUXdxSy9ZIMLj3PVpTY
XIG/VsqJxEOB8a6a8Aw6GzFEKiwidzQJHMqCtnULJ6BKyyVoP3PlYWrItSsMHO0YhfeKtFYmtKdZ
CEbs16AaCg1VbdSZuasszXEbRWQrkwIBPNxNcGDHnV3dsiskCtXc7lK/nZk1mWWdv+W7FBRMlSfU
Xgl32W+Vxhc9SChsEd35Bi0kvuOObsGsesTFbldKOlensJPwkvImQ43Xr4y8thjPtJnIGIb4LOQ/
L9FSli97A8MXkhMsXN9hlYuWlL51TSOmcMbU3W0USA6gtBi+7+UtHt+eWoANQtVAbDBxUUSQTZ6b
8Uq5t9CF2ibVy/8zf7f3GLiCVz2qbuT4n0y+4Mb9R68w+FGH35vryHCxuQfLv2IkFtG+zMDsBx1y
ENDHn4IAEv4ehFXXxJB9CfMoDmwmLn7z38aZ7+hSLTxtkqFHqJBFyZoc2TEODoFQj2K4c3rNoVXJ
wSAJkLxzqJ3S4JycKTXEhrUpCfiLRzHhIdjcaTaxVWlq1ziB20CmO3xpwINVHZc3ngG2iyjeIjsr
dBv2eieRkUhzgL2tp4zk67AfnSgOV+d71wyMaxP/bBmPMKQzPcCVo2ccDtkJhKcQr1RMVpfScWR/
70bPT6Q5LU1X+YW9M2olPsJmhcnr//3VVLzQD6wfXCY51qQ5TFgi2z+AVTKgcxD8xTCUMxl0QkGc
ZDbB73nJCjCVJvdSR34wsj/HM35DCduqm6xeuordOab92ATZuVW6z76tZP61zUz4wBj6rgoTerb3
XIVvYUML9fSDSudHR0g3wRqI2Rpu9tJVqEXwE11mUXPMH9HAQd1bXU3bTeQqGUIj6OPCJyXX3Rz/
YpqKDWgZZU732IP2QN1KSqiBKlxawtYH8tLCkKgJRrZ5XOFfZj++aqNky/aR92kAwm86ow9GVPMO
KlzsAvWJDjJGqHLsQW2QVHCsteV+WaxWkrk6yJQfbjoSn8hP8cSnpQI/oRUmUfm/o6UvR45gkawt
/NzCOCgnFRuPghKqxmHQ/hXpN184BPkSl8eX5sA0//h4p+YQHtC4qm2ejV7bMNFzmAND2wbPjTcb
p3spuPS/HDiDEvlIIaZmWRNS0VqtSF3FZ5fCl5Bqd/6ftsbsR/hePYaYGrIASlt4VoWsxCxwb9kb
nweMGUk1WsYgBbOCrnpZe5kWs4CcNR8XM6ynVDwvLtXYTMBszyJnr7GQ4N0YZeK9aWHs3rs7O0mQ
F3QXkvn/MM12kVqijr3ZVweD67PswDJNeXJal5ftxKzmbtKOcs4U/U3zAw+q7qW2QBJh6lrDOT/Q
1KbQg1MdL6uCyHTxHRYYViS+M98VsREcHA3lEAklREO1nxs4ZUSIDR0odPtaWGP9IoCkwOBJvH+W
Ztt0pB42llp5lUzUHRnSk0T0Weid9HMZEPPM8g8/2NIRZmFxaOj6kVM1bl5lTRpSiXzwZCokeBi3
Kh5doSQiJPWX9Ab7eHBnF3T2xYBLD9Phx0H4rUG7W+m866DCgrYlfukpFs9JW9dkGlpvu2nEuE3h
N6tXiBQ21mPd1rOvTPUcqQ0tyspRccxXdIHgqWodJT5ToFqUczKFSQzyH+J4xDvwAFbFFz4PDb+n
pEPrsTnAG8BVw8K4bCYMi02itAk3tlM0Bmdy1CxBuz0hyenUF8hcBhMKY8EnPSHi/0s7d7iUM2i0
qpvU+rsUSj2Ql27A1IGRZb7EoMmNTCtX+VgE3L45ExY7hGNEVJNFFqYp9IHDLqkyQpsThBtGcPYM
p1THn2WKnl8bYeXdg2bX6p8fFZo/wf0pWHTmIZslj4Y6OI8QwbUg94vMNllae4uzPjz6mi3WusFv
P3TIqQkZsFWWzfogehvsTtgKiSi5uaJ1rlb4oZYpdVEZwEpJZ6wRFLwPlsa44bZpGhUv5237/UK2
vrMfIJVSrumm5zgsp4BeS6EbuJyX/GNI8bmbS6/nytua22qNrrSjzlEq6YWpB5xO59aKYq/i/0zr
NlIQPL+h38p1mjNVTQCNFNWIrbWRQtSKzGy0JRu5Bpc+D9PiSNEMruJaXQVb7HrbTCgEWcKgrVzN
EYL3QNo6wb1g+j9Aov0kY1vG3J7b/DvlEZAf1ytzhHMY3LdHO0YbYD5RUTv4Zvflr7DMq7+yPiSG
ef6pzbJvydtZqICfRKvkPt8UFIlVwU7HrKZ/mt/v5gTYXNPTDzTjV9Fcn5tm9UhqP75JCVUmWOZL
3AZuiNPaacWPBXTKpG4bpOpOqc8r+1g/1P24VbNnMeJ8W9UPTsR+qiNUHTx+RIxfo0oouhQrZfAu
G6hVfxj089H7R9wAe026Yxv6QAb1m+VQIbaxvEhrLyFaGw50xjR9xScjHH60twjGOA429MCXTg2L
xEALU7oMrfpp1DvN1f9lvK9pQGk5g9oJyc6h7+8c19Sd+oLJjSx4NcBDy3DPR6/p/pTBWaZDELvs
iSdJ6U/kwTVcjdKAaFMLG9YfTGwk5OYBh0km+B3OQqFnkgRU6fKrp47XTxzEiwcoiyPP94QtFLp0
WduGfqFFbAo3zVzmBndJbsORLSmTG4fwdN4XsO/fLTAB9Lp48VwxaTbgKiuFIU7yQyWw9Xo7q17P
xiEA7iGB44yeaR3vfTtCUtlUb7jnXT5S+Tc2UI/vMlICpxU49rOnjxAaS4GPb3eSSHJpsBAorAIz
NDfLzGe5XThvSJGyV59ezbvnW0GasUpJnhhmzkoGYdBP2hxGTbKpql+GDsLy4pC968LcGGtW7D4B
hAZSs/VRS43lMYt5JduX002ZX2VT+5DqSufqCEj1rG7RHsueI+KGLjD4cXeftcMKMGAuVOB4/bge
ybG/c3dazrOyFCAW7ru8TsnhxCh88hmviJTZ8v5JWx5dyuOi5tiFM734k/9g65Pz30O7C+S/3F/v
vDeb0lmkyGbwKkela/h8EgDvotqMP406zoG1cNsKHV0AxaYvn7hlz/Z7aTQveNLqRThrScnVR7Tc
jCpu/adQxVWhFL9jlm6kI59gLIs/K9bJhgjlOE/kJsVsAcLKWvn0YEW874C3xooooVfymVCRx9R5
BhlUGdCbz2ek76DvJTCqjIio7UMF/Q96d451uM4izvhwLV2cS9Ak4EkXbRo4/j4pgoRU0znzQbdd
cauf+3e40FL1y1AOnIDXlQzjqkg92YH/pjYp1jVtFaoFZvAXncytxnzugfOTONE5jWKH1vuiA4Vv
ZXYGb6V67bjxVi4U0fPgEHrtHJdA/kELJLeg/ybBPMs2AGuienMZ9GWvKVS6twAtX9maY4D5W2lO
WGO1tNe/bnv+3BN4Ss0h9dZPCDkMW7vmQJH95EmnHSrxj74hiHLo8K0x371B7YtIU08tuxcy/3Ox
kuGUnHJaZ2W3/Qj7wyrq2uSW9835HZ7zoPOlzSkwoBvr0MfxuoTNUzgipmzveBtpoG39eHjuO74v
eTHz8is9XWEdLu9W0dP4HUqVhImf/bH2ti1EstEsfNwNqeq+y2rhdn/r2650D1SIpD5YxkuPyUWp
4aOL0mczo02q7jVhgUh7U1KwxMgm8v6kwjzV/03I8oe46KlMJgWNWInupaBAeTArG/17uZYMvqCw
01GwuW5nv1cPPFkBpi/tz3xwU2lySXEjfdffltLlFPAID2Q6NiFb8FWgmJdXYYy/mvUj1lri43h0
J5tlqLyzgBOkIDUW4i3FJNHLGfmfhC1AryliGbYB0m+EmFvqWnpN3WFckH4opfwNa/J1uFKZCFRP
pWg19scQFXuLm2zg/7qMatDUR3q81foikZwcyNpMVjEs3h5vmx58OZzA/3GKXSWmeqniMPs/g+68
U4aC8NW0WK+ovA4efmNUtbKqAqQT8M2WKMxVlztKuERQLe+IcZwbBfcj9HYNjzIuC7ZBdaMIMY+H
L38Laz3oXX3a/WCtIvf8owFVzL7t5WLkBF0eKHaeo5b/pCmGZzYANud5OVjVUlxkwbk+Uw+v7Lbd
wcikR2Z+rYQJ00ltRtP8ul+60J6ug+TKZGrRbCO/USZIZ2TF58M3J97NzOwB8nNh6EZVmbnN2LM8
y72D4LI8ardMZ8m0bSFZrRIuSGqgE3ME92elXFl9B2e9ytzbgRqtusLni7+kNfyDc6T2kp8wHASD
24IVv1SH1pi9jco2QN1XA1JAlD2rXyZtYOI4M/AivexTykYqmNyOfl3NpoAauLFWs/QuChClj5Ja
TLq/W68B8u6JWCROZaFDJ3gAaiF5TuE4rKk25+iNV+TaULwmbAAfdgQbN3tyJffHRXVVXcRXA/lp
KmOrj/D7yPp9h+hTNkjbMV2kRgTp5LZGReLlhcfcNcNaWAZOgWpiLbyFJBrh9fWhE8ikNFQnJSDk
uTYDuEsO8fcvzLSfWQQuaxnMaw68yfAV+dnPLWlPjV47R8rRv6WuPDFbOzOXgQlGnskTIf0XM2gS
f1mDssuZMXMtGzrNDKTJkXBY8d71NoK2+39UQ/XzAGtIdoPnfL42MLpgOHsPDGwJcuqMfYysNx8q
QRgW5X9bvc2p9Ls6NH2yLUzQKT9SZaCgqlcsFp2aJUX3kEEDrGVt1VxeroTnAtVg66mv2kEBfI8z
4kw4pEblaH8kNWzOWgGxs6ivtYierKSRP+dADUsiO4bWhBpTtV2E8Vvcocx8ccdbZzk2vQCWu0up
rADN4vljQM0nepW4NwMzt6+GqLPh/p+vsEWfjNy753G7Fe1+nGu+nJh1pHaD75gdDlY7Z6vSm12A
a/uY3QDg4bNf1DOYe2+qwUU/vSjO9hoZIRkted70jkQfCNz35vLXSV4/FKgcCc7nHRoVnofG+8rf
UXDNmlNd/iRhFixaqUpGrrheOZyYGA/D4WU3IWT6fAIMm/9A2oqrGkhtrnTtlrZvaiN3qqq05ayG
qyRhNv4ab3nmLfaT1D8ly8o6KKpeMSLGBpZBNCcDth2PIighGNui+iks1HM5Xh88O3Cs3+ZDKXsL
8YBmFp8ONHVvYKT2PM7sg37HNiGEyF60ASNorHfyfpYQ+e0Ml8N2LabKD7P4aepMxBU60QKzitxw
KKq/WFY+9cb1Yxh2aODfTBv9b3U5ejunXzIEukMT69IN4Zvpt0m1vNYurYd7BleXihHY/omL9kPM
I9pxNSluSyPbNarjv3N9YWoT0Zcw3lv9MBIDb7zsS+saNIBaeACiOsY+xWHIml/e7+UQkNHdx+eM
HaVeKbNzUGLPGuV7TBMKq/sUili+7Fid4BcdEDQ5rEb25tY8L68vI+JDrLh5/WlfoepZSxfXCVnq
MmsNZu639ZHNC+n/7DB26WG+wBQ0uQqWhpKpySegRxLd9JKBH7MVHARFz6eEssJjSvKYmSuwixkZ
7n7m0gROfOhsSNDxXPrOcMJru0mSwuV419VHaGNw+D2SimOZt1A8XIiwRrS+JcS6kbfrGjvwAVvu
dcSNvAc/ZfJ39N68hfINJL1kFelkBaAufkta0TrVL9QiH8SqqQ3YyVlTnYgw/OUaJfiRwSOnKWKU
fiGeSzJ/7TPBwUfnD9fLoj966DPxE+oS2e1jFP4R9EHt/yxfS94Lw9uPXFZ3Sq0p7/1ZJLrVRSN/
uN7He8uZz7R/KypsPcG2aB/0o2fRGp7JhMBvIMji9rzrFMBsWOiona+xh02aPWQzwIxgfkl+fAeW
eSyYK5yOvYTX//wvw6/TGKadzt9iAnx/2SJJ0X6sy5P0fyNHEgJdCbpuM6uPtM11f1/APUvVn5CI
US1uM8zjlEmq2p+XX5KusDJD7VAl1eo+c3bVCilRPfj8SttxCbSWhrIKCRHABrrkuRqRJ1VrUT4U
zHJDN8vsQ5Etp2usWSqw7ADdgqiECvK3xeDxDUukmC9EWGu05JRLKjapaTpsmJe6brGsrHBsFIKx
1f1r/LgCXbg9sZ5Sp/aj019ew4ZLKh67u9rptd5GQKCGRF8OwoWiGZdlv1GkyZmkl9u6zFA7/MlC
pFp56dmPNt/mGuBDs7cGiIDhcYwH7tiNn4AYTZH0CluiiWL1qfVSyQFB/RcrRrX7GZ5zd+SN/OvA
LcAxYKxLgZu3qDB5Q9bet8/3gCR3y2eBg2LodwGWYA435ANAnrpIkxRkJdo1FsKATQ2kYnoZELfU
O97+GvVqt1/7uUd2+t4c/sksEy0cUMI81FHcw/D7B27eXgxGGe1fM/Yv+dSy8WPsYk+pYF9j0BLm
Miel0zYuRkdCe/E+5BCWnMKr/xydK0lUwDsmWOBm5ZoY0/AUiGCKg+XMHYU0t7hwc+QkzgvtUDmD
RGiHemrxvlFCONSL/2FLhdf8ukKpp7ggjrJ7BNf2ECJ5MjvApliE2VjMQRWrVVe8Yuuqe5RBsYh3
oE/MQn8WP7SR1UIku4YwiZ37zBLI4QhlY+ngUwtQPPxe/L6dfcLCnW4QI9vduMlJbuZFKFn4FN4+
pLI3w29inRGy9xij5vH72QAxVqiGbCtlMDLZOokKU/FGHamNWqpdoKf63U+M9170U5zZ6tP40wtg
NN4Ap4hKpQMFojpK5tmNugsn60djmkEpHnFMzPLtsOfwcYr83eUS8alzu/bYkbo8jjkxkBxZ5QFk
AQxoX6Vuxd42yMB5SDcV0wbcNP0GUvgV4C81MmVCBdmYbHPIJ6Du9s+XtKqQbjB7wI4XXjlnJbMa
ZQfXOzIQb5oq9j5GAXh4YoevtkAbfsVJmNk7eWvBhhby0pcv2lcYRbf0mc2ZDDjrnfrlQM5mwMDK
C0U5CPYRjC4sAdKtFGR6QJzJekJo0WbyfUNlmAf9AZ6EMRPtKs/tvH0vADsW+UteSMx/NJLiwyMu
0p65HaJT5T6I/iLYi6ZaTbJf1idwieUSGPdmP0lOgktlgD+hSlOaRMVykCJMHfvGDwTX9WyVjHkU
U+o6a/ydumIrd+fQjFzllVwO7NlAAC3Ol3U+3mT6v3+unmXdkvGN6jnVP24vo3IVKJ+MbzRm6nmh
t51fAY1mYWQsafm279EG4Fq+r3/XqVn1UXYHV6CPJCsns5oj0KMKL3Kg4mWVofSmPHq4Xv1UI3+f
0cN5cbVs+NCD+T8rG5zuWL/j9Rx4RrdQ6OmCYN972ssTe7A469bNG8V7EcjhBxGDeZrJiZ8hUVl1
4tTQmZ8HA23Rc6nAzukTomO1xzoHk6/xvSIpb1sr1Ei+AXnSC2oup4u2poisZsqfrQ5+WHjm/U/h
eYMD1OXAfk8eLi0pOMEmW10kXFglj6VGofFquEV+yiKM0ABblolLsRfr5QF39QyhkXgjAy2yXMhp
RWg+po4zPAelSDG3JBNPXB7y4UxrUtqsGBatVNgFMRiyUzddKdn3LxnG2nHDohBWcpPk8RVYPVHK
779nWq/XRTcFmGqhrxytk7v/xizVq44vgGp859WllcOIXnLGnzvYpYHx6EcOLMZDTR8tt/JycDix
XQsd3PHhXmEBvdWPKqAC+PXUGtqFW0x3wseYzdovlpibcaxOAYKbjPw+ayXjoTbiKMFRsr2h4cya
zBd6Qc+kAWfq5091kJUuDuiCp7NXbDGjp3F/cUkslFoDc03KwXCGgyL/mxp+kMJNgiWRYlUW1jaz
MVELnsyquoGv0SPE2Uqpj8N8Mq+IUxmreRNL//U428Xo/5MKI9j5Zs2qcBaio11F4ZTjSg6n1cCO
LWhb9gSQ+m9YIvRfL8uCoOysz2BtQeMzOIAPOUH2eqk7fia7rY8vrr+GoAXl8Sk3sTMrKZ6QaamP
slewZdykfKhVUDHu/MI4GaP2r/C0/7vtbQ3cvx1iRVAPa7XOr5aNLiQM2gqbylksf/XTBTExw+Px
36dpdkn/LkjTffjzSBhBEPPRpYFnOweiI7R10ZjCvWswTv21X3amTLKeY4QtFc4Y3P1/Kjj0VytN
y52c5SaPHpgOFw1r0Xpk5bOy25doomsPwTTPIIRaM+DQ+imW4rgBNSTRqUC0oGA9heW894e7mo6P
/b8g5WDVzRTdJpsYW1Jhvzcw+JHkBNmTKSzqn5lPFRJlts/1WsbuQEO+cDuumAdRH8SKvhrWf1HV
BFsz9pI4vqO5RrbumYwN3zZKLssZqCRMK9/hu0qYZamXdu6pQM/ghHW3zFflQFf12kaY/X5B9TFb
j9L2gGIFsU66LcQJO08mHzIly2AUpnIGNoT+DB5ne6ASFT+c38TzFscniIKcchYlsQKgBzzF34Ig
+O11pZklzxSEIH/IYEfZW0ymB5ZUUhMTW5QSoC1WnKsS2Wg26vN+rq+Bc29hi1o0DXO/lZp7u8eN
eO5AwzH0weW0GXZfjFwhjUUws7Fko4JRxXaahIglFvJtyMXz+rDoo0L6cl+SyAWo++HXiYkWAZQz
LHfgbrQEUiLycf/yOyCxYy743+coLloHj2KphQ10EOu620GrcIfq/yZAl5lXFuhZP0K2aEXUY3SJ
Ot/XzK0LMg1MxEURf0y05OMC55ZX5aRrtACEyM6tg1HMvu786A2ux4GmNtV5eOTwk1JOB97xMe2+
tBf5KGfjl/rCDyMkpvjUUw4dVNGXv5Ko3ltBoM7wopMPpSEa6Dl15RRmevRlGWSC8JH/405HcF4j
ayq+JfgVPeEUvQZYC21p2+UWc7foYIpydwBOodU8AzWOWkJFtDhbkWiNBFkE5JQctOAfWy/yUPGF
63R8NbBopS7P+4Y5vapJyh8fMM/m42Gn8DkM9QBRcwmSV71Js3MXIbsJh6ZQrODA5VQpc3oeOX9/
n7Xj8SAqYubFK0w9Rc62WtW+W6jnUgnXj0ofj6yTlEFBPNMOlYWmlSU3tfy6TfVLTgKnFkhdOYQ2
lIbk2JUvSbVLMwyHe3HzjTD9pxi42lsRJKVUtAknaTlUwYB+fB9HgnYcdIepxPT9Go7H55g3EF7I
kDDUyV6uHOKVnLKOofP/LrRClpY4Qd4TAgPj4btijX4P3rbQ5GegUcyzphR4sT8JlU8n9s4CzeaQ
KtvuB6B5eAF3ny2aA7T1n0oNVNyHpOA84f8b1QduRVUXwX48Gji18caJnTQx8gagmhdlpS8Ix8YA
zlPkVX3lIZdRhRj4mvhJiQtwUUojArWSB+d2FXpbK78jTA5bZtEYODjyf3JNrTT16n0kP5F9naZH
tKl7ZUfkYrasGdoQbITmK6deLzNtG5bHLE4kEvLTGfl0OJp8zt3YPVDZ9Bf1YbUhM4qmMd45xVwq
9mxQ9NG5pc6lm/kBMcORyPXIufN1ZgMj1BSKAFc1ve9BK+YscpoGZew/LbLL81Z+QysuuxO9wive
bpNgzEzYRe5OJ83csx1lmYIw+JDTYW6uX+i/9XnshtVRKJEPHtoqzIhYVyCkmfZ/cbqhj6g/AuWm
2iMSh1Q20iSkAG37PZ19ipT9EsYJJN3eJ99Pmh139q3MHBS+H/cr/iYRACsUjPElD46cXGP2ley5
HnA4uTxj5l3T1iq/Woz7uvFCGHO7IJ38/o2pzUTW3A5DdN/gLRgvU6w3f/v6AUJaj4fcD80QjQOH
y4RTmAIZBSysazkbnTegfVM3auLXnQcTJ9LgQmiYkql1BMAvpUvGTIx3axC43aq2KyHKdezg0nEf
aDv53rY+pPUOkotnchiFOB5WC8eU+6a6OdopWAPcfVREQHq8rfw9FWn1Irx7suVIBm1atDXjF3ta
m9M9jG0qt0ELDwZORMdNYt7to14XT1M0vnrD86W0I3r0MgU+vm7M7yjdMyiz+LzGxVSvz9SgrS25
Mbc3SNBBbKohCyzNexUew/GW0FUDs0jE9Gag6V7Q3wO+o3v6ZPlO0Xrc90JgM44OSeS9SZlJPBI9
v6+FSw9vaUoh7jdyTCkQop8stj66GmWxP1wZXaW39X+B5uTueunMGF3YMGVcEoARUJwlmfbHy/tA
c2N4ywjK666fDTAPnD1UTsKeFWS/nAmS3mNdinE1OiRmZj0zkDdy06pXBphJiUEfX7ufv5uQK9N/
IQmyTeZ59+6Paju36cBQf7TXYcnjB+M+zRKbHOLmW6fbgdwasy3mjbIoGe4066I+Co5mVbb8WYpV
qwQ2nRTHVN0av0HmVoU6ar5j6tZaJKBSp83xpeiBdewwdoxzqe7b/nJK2Kh1L9hamxGV7xWPnlVF
xVIXf/3EfNzd+PLExEzCus+cHqEuunPxZHxcf+V9OGL9UQstB1O7pKguwaog50ygfZIYYML9Fjjw
a0XcZCGenlYYJje2FRPkxjebnSV+rhGF5ToHEgPwI/CYa8t3x39laUac+EsHPNsTETkImhs5lCQD
B7zY5873Xq93/uO6YNOTEKhXD1v77TUc1+hOFT5QocMN4e6mjNeY3nuamd+fD6Q1xTpV+RSHUEv9
75qvPEYDbccfQsH+iSLXZOn/VEJbu2WMUChz+ee/nd+NzcmjGYlRQs3wVdVLzrfZlQxJPHnnlIi9
LuEZ+eNdNLaT6h3SZDq7S5JiE8Qz+N2pvYoZ8j+fC94xBAorF8JKO4/MOccaDia07eQ8x871geQM
BL/SVuVfLD8jedZ8H8NW4paLVkedautUYx3sDHaouR14vuhbTeYbJhLocUssiGX/CYfBUgDk7KqK
/ZpsH7zf9e8CvXLsw/bpImalv+jxyPi1sbcfOP53np+WiGtA9Dm+csUZ2y5wHKk/SBaboWiXg0Ec
v6u+W3Ka+qWJ8gs2+Os60g8bc2qTlBZrhzvl0UwC8JLKMVBhHZtvXQI5g6UDWeCTZzLO8ZLvWqKf
zdv1MKiNMrairBD7n39Jwk7Qlp7DMbSXstBxTGsw9PKAm8+zswnO8yFCauq4LJtcT3IWGNwipxtb
7Jy6YFpRaAaMCue21wkakujOippm+uMURGaOMW5nGYLr/PLf2jU67z/9yKQIzhFMIkeBtnmDG4QI
v3RDuTVrm+ygfbZCEQP0/qLrmp1MdCO/zPzz7me2HZE5t5WjLs40AllD1We/No1DqCEFG3wUVADu
6ja472mFIRIRHd6odY73u37Xv0qL1QmwYkq41gLvWY0DcJyPhAi05LixlucjL/RJHPuCU310RbTF
pvAQPcpwAMYsOz0v222jaLtc+NefNQK7JoX6QW2bLHLABhtIWLSW0zTQwRIn9g3L0npHe7C95yat
fkDrCNAkutdkx/BvnHSaPtcNMkaNIqyRmAtZ3Zt+I2DKFeSc3uLKdZKD8WeUIv9v75VoIDQjgnqK
/oAFGy4HE8CiIQ+otN00fj9O7sq3mgrbTtX9RW3wC64biqD62KYtW94xuJjrgO7CqLAnIhGoxCpt
LMhlFAQb6qT4fi2doeXKiQ7EQBtLiYUMbAwsXSGOtDF2nCOAcbJFG7EFYcb2R8jV2fbj65rvX+6K
SinJw+SURyuHZ/gV+YPAPVHAMKCpbqZq/Ts8gpw//XQzxeQ0XVEWHQQXCaGP4ZDD90xR5j9bi/jT
DKhvMtAGzpwL/99IcXDDh26vx29noCqh/uvtmkL1W55D22UKD1/UpPLEj4IHz+LFK0udgWoYb5NQ
Q3LSTs/v6O3T4jmhXROIBwfLuC+X81lk+yGEndgwp3wKHqoeciTI5Iid7+wnnJuQXXJjmKKGNK0S
zkFaKVdk8uFZXP/28ZoTmrY7fc2rEbcmQURiRpA6YdiOETfGGChMAvO2nwyFT/RBcxcs0LoZeY7i
RDmakuB8Qrobt7gQJgBGpnRHyI+UrizDbXDqmR3wY+EJDLzvPs+K/xzbY9JE+Fz5oB7B56uvtg9w
ocPYMtxuqwuXg+rXsTR5I568rIGgbg4dqkyx++5cP7s2MBerUvbjDE9/e2WSsihdpFtTUSsFE6PU
nmx2UkASfpiQo1RiUaHthVzEC1T1NCFF9Me9nsselBXCBvIkwBT8bBAChlzrD+08HnxOw4CVN9Db
CGzs7unr/9Ob5TfILzJQH3D87jrCP+teSxW0X5EjHgEwdzzyLZmg4vFqiWDTXW84Ttfv4PAohNgi
zNwUoJyAFxcStRaU7cwU7aRjNYezVtrLVDm3QSUmpB7IfPfg2RNoh3mzizRVMEaYsvAXax2qS7qk
BM1baqTpGfiDP8CnSHUSlTkMB1E5Wnt/39UXLRBV4irM9HLJ+kIbt0RicNqd3GiAgWclFBcPI8OE
Il2ITYVgJPvOPPyP/r6XvJ0SkwCbQ/W+Cs+vAdItcu9rkjvOozrl2OPi1ZsAlJg97lCXNFP3WtPn
kRbJk5I0UXVn4WwG70/Ij+IS47MzENN7lkaxmbFq1v9BgeSCqwfY2reGPXdJnVWNiAHWzBA704Qa
4guoQVohaBFmFrkIm6fSPZ8OU/BqmJBitk+REzrVRXvNWeIgDMq7RwM7Fmhp0yFdaJOLHc+ZOuyN
5BNgzYKhOzTS3OtewwXZ/VfAvIJOIDVTizjB5D3tuCdB768k3N3ZkinydBrMmWpubNNT86u+EHXO
nn5hHFtOhpwVTBEGBBJpsYE0gZF8z/2AvDr0mxNuNc3z77M2pG6ynkm+DuYoJX19rXOm36yw3scr
YKM5b6i942vJ2eNE4V1JzILtcOAGNhl/AdW9vEpVzz/aGcST9YGq7HNDn6NVI9ACMXpKGbi7yBU7
SUMLwZ1J1xVwJnP2KUB91fxU2EUNPPAQ4FyF22G9kG4REd/DXREtRoYzARIZWRQShZuzfN8WVj4X
pCPMTkEyqvjMnuhQDFp/zlI42fbw6EzagRD8t/fZQ75Pbu9TW6xc8rRORbyfCMqsnzNRCoHhUMHR
6KaEISZLJi7ykNK7Kf1fcZbWM02pR9+nJo/XEC7dMLxyhfz70q7QoRBNbXfYfw6eAeAYhbILhXWc
JOP74ErM1Am1um69kqPOyPKQ0EVtVOaWeql1TBCUnlfzTNTctNWD22q3lnFUUafIfZn3fGv4WPaM
Ach/U8WxMh0xwByGsMTv7i3CtYvM46nWbIRPo1xFDqq4e2yIGspP7t9pS3WxomXfc9yOIRZLSjIV
Z91/aMMe2NloUKT1TBnNFc+JnTCLUnU/yxlBFqmim/pkGWFFHo+fR0GujNB73hg51/hAePRfitoI
K6CO6vFnQ3G2GU43WVQMJREqJWIjIlZ3KGbyXt4Vbii1QWUKiJ+yOTpkgC4yUrQMwkB8CVXnSIfe
u5MYQcA/XreIQO82AcBW/kapp23nnIyerAnZyq90PPkb6mOXC9HxuIMAd4qRuw5j/amEvrifQFzX
uk5lD5TfcMoyRERuXBfg8j0PIlEgh+/DPZ+7y7lc/DDtMKJ7c1GZVrWG74APr7Zi+E0JrYK7qWRq
YEtd54e5W7mBvL2pTJtSx2zVs3/auSNFtjqtXyKmkms6RrJ5UxNWt3pZkuQ4BTMScKWEZ1Qy9upO
PxG0sFGOM4tv2cf9Y8g+JHIf253ETFIn6RQGJYCJ7yriHhTn41DDTkuN4tGgcWCsJmJqkOlJcLSa
CGp+4s+he2longMQNkmXKtax65pxvwSkgp4QSLH6PrA9Mm0Cd5Oy4a3slM0YgHAkC5pHl4MRDM3a
7qQgf8VAgeOjjygNo5KChC6LDkkYmT45pl8go53Bs8yURabdhP9e8U2DlGTTMbPadbTeefK+P5Jb
OPvg7LLYhbCUBwksKl4Y3VEbJ11ow98MdoR/90RDyQ0cJNqA/uQ1bHX9/fZB0fq1MQ8qEYKnWWJQ
SVFo/Q7VCiLF8EuE0BBaGSUf1yp5cEBgxJzB47t9wS3IlXa8DBJblS9XqLZNyteUfvLT1qD/z6Tz
PuVqlGrhpT0YQ7ff97YHg3ubfxrFOWE77K/LXw9czjc8q9UJjjsDCFu0FmPnO40ADwGli1RG9aJz
s6MLuItTEUjr/X/A0kjKK1HCU9WYgJZvAwi1f0jfy88HjN+Qzriv0/2/l9eDgj0Rojo/CiDV2bYQ
xAYzSmxTvtr757DrwWuvwrDqitKwmceO9l7AZXoy7xgPAAJZeHxIhjDnmuNZ8FJBMBcOkd8X8TUV
TL4iEimV9XmUXo3k/TLXtEbBjyFJKCIf8cWyhIXFS2M0g/Ijcnq5hYlo0YZbBBD2FK24QjYVNWSb
jOuDKg9GAXq2Ay0j2s39w27aaHyzJRX+CgklhwQHV6GPbaf3iyJPGV+GRH94bbs6zEf5A4yYj4eU
n5mFF6BfFjWuyf/cMx/qcSLCa6+aUD7OdWWgYtOU33PN1loH6HCbvQ0PGaixjXlOjirkwNBCy5pT
nWw3Fq4Gij1IZc9EZEkwow2DeNK5G1LrCTPPHlmUIExrZdQ/GsvlqIRMeZ6z5QWb8zjfOtgwPP4n
CJXc1jZUat/G5cq0rvip9XbizvyUiz+O7V5t9eLX3S5VWL/NsjoEhjfz+x4OTOvQno4R00YD+nuQ
usnpfK6OzvVTVL3yXjG4rQLsRgDUZAYEqGUApUroQeGDXeCAxliF3ZJ+MYOE4Ki5PLClba090xtx
8DZROa1ZnErUeadYDI1OHrXP6KU2ewFFtTd/o0f7cPaPNXhXIgcHU80AItiyLeoY9Ay+G6lOYXM2
LUIbYcXzspACA7UNATsgTdQOuMs14TOs0hnlVL/t0ShjLtYmYvGaglUI92FhwT4PLf++N2l6UhIn
pH0x2L+xdBKA+VJazhiILst6Mn+wXlg6eepqRrLW6HBlC+c66O5fOP0jMO7CbiRSdq5cjPgtKDQy
s86PN6s92yKdtE4oIYOvPwmm8ZvlvpryMEoIrDtaeRKaAfo5vhWKqM1/RmHGH/Y7NSKjfm8ttd0S
re/V4jCU7gFlwLTCzKGTol5eGl5kRA/MI+TFtbuH5yQzMbLovKToOQDiqLldA6EzrsSWZum3JHca
ZUWD8ubs1jqOiEj5CO6FpzZBm6fw266++pcIbMkSGGrsUKfmWuUvR6TiFSeeKrwo0Oz/ooHL6UWj
P9bDqZAEp3DsdQecvBYE2AXzESDJsrNFcf1HwQIsTv7ckK3RVAFzU299MzMAVCr1f6duRkQZmdM0
bv5oejzAglsaOquGIgkJcVy5UPRFF0OQ1XsQCGwZ7lM2TKhvYR7/yWfRfzmDfVdX+JnxxgF7iR0u
kiJtHr8fn2E13YJHGqfQy2uhmiw3DsEvHuag9fcF7IjI5V6thrwl+DBEmikY1//bxH1hJRbL4S0F
i7LOwz5dXQL07ZQ1UcHk+S2GXIyg/844w0WuRtQIfq3wXlj54q6M6iCrfTq9gteIQv/C4BZwbrL0
CSW1iDZuZYgstW910PPFiVYFfvSzJqNlbTj31luwGaO4xK9T86FgtEDCc+oRNoLD8WA7rKMNXWcR
v49+G0LgjYtcRldA1HCUqs1F2AwcyUjZv+7HTzXfNG/tZe7oxM6gXRd/OuUObDudaaz5xmuhSAEV
VgICPNzBsnr4ZBQD5jrYjWOTT5ZEb9MxkMYBdRIyq41mH1xEbzk2RBg8+LI53SAzpVljk/BO/GJ5
ruXhMnkGNXpzvfdcZXo6Hb/zY7MtbJEiaicNx2FZH/Tlrv4CQZgKkRsK8rNrBXe15PhRE+tILclu
aRR6AzDi+pNZgoeNEj3fUchtDs2z6dlnkscrwzmhS9TKbLwnvdrMfbNRA3LG1QiiBR8letHLQUXM
Ot+tyS9Ar6qJC1UUS28zNEtJxpSH6wn/TgvcPPraAVrIIIrdMu6hiwVyYL9BlOMsA5lGHcd61+73
oiAXFXehhyJqixJA2riAeAFOsIWWmm92Tv63bP7GlqGGfj6oOispP6gLVqGRaHHbZjf0VFQod8oM
LMYsutwjO44lvny7xI0ROdPYIDFCoC2URZbawXFWozzC+bcqolJVoqcy8ylRvi5PHdzjmbfs07V6
oGiZ0LBzmeyBvj0S1y00L9ykgWk92qp8oWl4YzpgFoOyAhaUO1gsOWHDtGsHIKV5LG8ebWw4mBIY
W1gs2M40sb1ELry6zNS51i58g5H+5p71NvQ72+i+KY77BkZcQuvI0jWAI5l9umV1fnJtdnaFww//
PbwuDH8hy+5ZIAmUpF8qEG6S/ZSd4QpRIg5OUuaotgwLlP/F00hOVQH29cJLiFJTDVdtC4CHO5hZ
ClLYD7no8QB21pCdkYTtNkI2/k9olU15XxmuNFr5r1LG9DBfZlbaBh7xR20zT/IguAd6EA112wb9
jsXV0cTdyZj1zvzwTF1wy8x5bLM47hVoyow6f8yndwHJgYF7dQA+rpk0JLq1AjvN2hn5CeU6mySt
grZq2eCqMw5bxf8UCroy3ycHr5frbbo3eG+RS0Wt1FqR1AoccQITVuM+7fbqlYjoFAtnMCJ2YFoR
wG9wD4b4lszPd3tZfBGx6Lg5qWMCJrFpp76ikVJV7XnaaVyJQZn3coDv5WecUVuz0tLXlzNikHmi
JkYZb5mXvpK8fS7MQdNOus82ixlTrWBvl+w65qKM0DJJCoSu8zGGWgpn90MsXzAMTQLbsZZuI2ia
rAX7N3XbHaVMny7nCJ7C+2/aVHwigsSEyE5OLxEsSoX8L+yPNtby0N4LQn8hGSBJ0Im0MZ6Tb0q6
bsg2tiHQAODD7uW+7fqOS3urvHkr4VJTNAuh+nKmrRnERHFXXm3sinYf4OzY5c/UxQtuqJ6c7b+/
FAFd/X5Wh3YA5vrh2rew/C8BRuyPBjox8STiZu/1T3JZKctvpdDo+Zyimx6OcCInl8KodbXlSbTZ
MifoKF0QIs3Ajl5cyqcv73iqyS48km6fxvZxlgQRhej3iGSTrvoWqa1W4yNLqBRVoIBvJ6i0h+Ac
YS1atLk3IaBn5lMftVWcA+RCFfn7jLh4MQMiO9gZMi+XhxCYQ1Ut3WG/cg9wDBOoI0jINCpsr1f6
tNrKK1US7j21xWWjooUSe7Zi9/LN/eGlS36CZyyqGEtIp9VZw3C4I7YrrLVkOKJPPf1nrE+e0Vw4
gueS5EPTFauZCDOnzwaV5NHz/7nMMqKSQKgIgszTuTy+11o91Hb1WJ03IPGUzSzIhKZp1Wy6p0FI
34EnNLX/w9Jbqo4BRVf0nx8tGMKsJuG0vXg0d3P2dsO4kQt2uhrPilWqe44Zc2f3uCl3BnhMQ9TQ
OWVyWyI26o7QVsd5J7+CsjF8mmnO1TpXTVeOXLoDZ89lmwNtQSkvS32O2JuBiKyJ9moTuLP0mb5m
tid7uu8Gw+munW60GYCvpZkTiVm5duqjGYzJ3LrEladO8dzSGEpHNaCtJAh8Rks4/76U3jniIilj
KU5JFMee1WnMv4ZrHhf4vkmVfCiERQnBXptVCWbw9uLD1aOTD58Ac4MKLEd7d7NItBvLjMOtNBq5
0dWwWD6TVacBxAVFhWitxcRVFjzqYKBScNIbXXctrKQ2zoBHBYtMk1Mg+6PeIEKmsNXE6d8BQJMB
MYzTTe/6BGRxAU6FNsbgDe5jE+j5UiPqf18YKVLb3FFIhkWmRf/50ezz5ZgA+0eXhVHi/Tb/2ov2
TTc2L14LeIKeY+8GEovURg+ozYpxU07xOcESmIb+pbYHNUFt8hN/OsWg4E7lqI3tdnpzpNOSWRfZ
yAV5krjl8F2VImHoCQiWoH2YKxNoVgr259lv2x6rsUsF2AvXDE8MJ6+wld3n5LYhMpKNRgOIx+UX
HkmRo9Mri0fYwNjRovg0VJguMrzWoOAJz5u3sXvsGPYj1GWF0EaFxWHJdsuGZqXgTSlAYfcYOcN6
5gzGxN2ketaUrr4WOlXhgQU2fXlh9wDz3otHpmkcI4aAAw4FtC6lNwF6+UVu06HOO+9TRMotqtp4
6WMpO8YQyIOSlwXa0999HWUsZyRZlrotfJSZmIzA4Q+uVQUrPqIR/aMh1MpcBR7O1WuFyt5QX9dD
dwWbiTA0XOeFb9mXdrWnQ0S3FF6CI/N23SwrzddtI94tCqgXDNK03AAFgTg7oLuZkuxoDn+R33PK
py4lVo4sC6k2gUlhYDEow+h49MjDaKnRfbwhGApWv40HCEcr+1cM8NKAtIVLjDNXjKdptChnwpFm
YktriWN8zQ39XMXfeh8C+PakJWP34E40T8YhaMvkVDjgXRUy4EISqng9frGemWaVTNrxD/j7Bu0J
/KpmjywPjC9IAb67+e2EF8wYXCFp8LbDE266vlnZjczEtozFFDf3qK9pFaceuCLirAx/OQuyZI9R
426vi8XRhf75F8d8i47UnZYpjZiqIfPpEulNlET6XpBxPVOV/E57VUgGmKVgri2BmceclPDoZeRA
CydHPPpe/EtyeE3y6mNtQEizgQR3S09e/Rrj7E0jHymNv9QHVwV2ErY600uilekBZwhJHwuZFYU8
rETtjUx9sGDxtTtrEsczlgZugH62Dec13C9thTQ9zpHLzeMu6tbG9t4Vc9NiPZ2o2LOYRTvOISl+
xTTUZF5UKXkI/WEAG7G4+WG7ERKjqmGZxLF+4EOlpgrLgQfMLAnkZDtNv10m2fnaW/JUPnF12bER
JdZyPzp3+9MDjiWAJDNGC3yd0mlR7/PkSSz1888y09K/SM/D/EBzlOx6Kmor+zfttwK+6lit59Ag
dfzlnnzlZjHHz4d9fPfF3NuSWRrX0FEr2sJN9cQtqOwV5cT5BmCzAX4bIWsB86Q0aYGooQ9NJ7z0
oZn8koUUDdKsmy4+X3OMCvfKWFADxwLwDnemPNbcgwRSARcm9O8xbNse+ZqhmuCHNXOBEqKrP6RG
IuBiEaLkXjZAaXadvMi61blclfH+78OjqlIgi9wFT1ECn4XESXgEY4o5yM+DWO77GQDzg+DsTAx4
FUVZuuYWWUtnL6RKrIAJyeJxhv4iKtHpnj1Kiwb8c5fgtqpFRrkXFna/oMN6IAkzgS/PVDT1/5N3
J6R2JXXzeIW9hd8NX1+Q/MceoJI7i1zbf6WsU7zQa1DjMfGsL+aeABditwl0qFc9508mbDurQBYX
HIoQCbdrpzExfrUYWOPWjSGRo4NhHzrKTHm+PC9Dh0aoczVthZjxjeVp9TPM/vmU1wQZTyLTrHZM
ebVi1EWeNTy8wJ/+HLib4vEAAEqy4e9AlYa59oe6zq6I5H7IUUh5ye8wHFtT5KblPIXGB5hMAL/A
m7FgOFAf5n5csSGVo+Ch5dwy+3pal511F1gQaLeWBLDGS6uJlFAsklqHY13+wVoOSw2J9QxdCx1f
F5GyXrbdbR8YPSruRylfsyl0Ds7mwhG3Uuysh7VvZ50GYtLhzBQnPlGf5JC8fng305ppVsn2FAxO
nw6AWHCT/E7xAeboN5iNZzy6T38F7q/KazcVpC362GF5JC95n6chJC6SZb3uItBNADGpoBdAP+j9
9OURVMfjYvxFKSxbyi5VLInz39XmCAGuN/+3HyTi2aUJenZBwBl56s19kuoui0Wj2x125w16BP3x
tS6UizbGMDVuIrt6VfuPH2rlq4gnjUv0ZCpM8kGUnmOf5qsNdRganE4dTLNS45MAbRRJU3M1pRUZ
MnGe1ayOA8Ktkrqqupn+xD8H6a1AuW+LCTRHFRMYiPblkqAZiFV1QDc2FUJeCUJXhxHsvzX16rHa
IZQVjVx5P2w9BlROQpSA5tfQ4m/r6dgvkr/ffgULLqdGWQgPGLmg/O2E/hszRL9KsrlXTYhDjMJ0
HoLMKAcK2MWe0JP5pdYvsb26Jr+V2ONoUm2nX9ITIzcsHkZE7X6cfI2ZVUtt25k3wlPJx3obl56m
SdINL3csmzNQgKdLM5o69U3UxdEWtF4crvky0WVz5DyckJ7XN+SmhZMP2w55wKX3vsW2zoaiWBOZ
0TmnAjg4abg1I7ep1XZKRpB/i5F379zCfBXq71m/e0sUFCure1wMI0c4EEWv/ged8BLzemIE97dl
+iQ+vswhV+nLgVqgKahC4f8sUPmiOHfjzyXr+hMYp9DXu7HNLQszBYvojVdIpvnjpCWALSZ7ejdw
RwWtX645fk4SpuQRpXFh4i3TmXeKF0Vw34bznZP/Ec0SMjhBBjmgfzUMg/iexdriKTtseauumGnw
h4uGQRSFIDsnC4UCWLC7IKjTWR23y6aM9AP3sUxTv24L+7mhtSc2B9qjnEXixbPXw7RZzz00/v/B
gCe6cRkbprunJ7MhknsZ5J472IBsrQ2T2QLAhEyJmimVqQWlU2xjwswyOCtyE3VKg7E9syllI+Nh
UoFGmpfQVDQdS37md8VNPGub14jZdBkApJ3PCO6mGx8IiUm2lddeyXTHZRulFzAHNqqNbe1xS7pG
Vve2LCjmxJR9Sf3830O2+ecmExuX8cKV9jhtgTUW6jfBNOe0mM5dPJMuws0rjWt8i4Bvf8LJNEXX
vUwozHuauGK1m+DiC+QBn1Gn7swnbSBl28Datlu5h6TkBtY0ckDXAH2LzDRZ/HNuuzd57El9tLM9
7RytHYCM3M63Tg8iTiaugTM5tP1eS7Ry/jF6L58bUOTPfgeTwP7IWG3af+/Vgxojdr6+QPrq4srI
wdwomSkNjCB+b/A3691ePcOOSHKB9Lpt+Yr4nOFtDvbQtUqk68xMfNNYafKEK+VFtidLh4uCL5/a
qlERcmm0cw8bJDEbyM5Wd8N3HMPGM+AOVg5jusOkRPsG8AqECEmcv7f9wvqBRbNUOgNZdl/0zzck
iV556aTmptPDjaLpVZPK1+egtmU5AltwGz0WK7d2qf8MkmTcYDwfnzDMuQ96P/bdQAzu6oUeaY27
szj3EgF6HK78YsgfwGWdsPiFenXt/YbjlhkmT5/l8Wb+ZMXiUv+BQXPnhKHIdxohsvOfWJAkYjod
actkPPXrnx84aw3tIj5JZisTpljIp+DxkVdhQHziClzYZ6GN/lVlWQwjmD0wN0CZhxvYe6l0Mjyu
FDrp/7wGupPYpnbbjrfKg6KbZ0frtTrk4qxjOUZc4uUG/zNcw2Z5TuejJV1C/Vg4Ai3XSeJg+0AJ
6jfeAw8YQvDxy5eKITy9ZK8cNVEM+b4SSxzkmKNiSmT6q/7so5DgVkj2tbM3lk4uUkQaLdS1CEs/
ro00KgbpJumD4LkP4wQ+82zjktJhtZ/5KsjvGX6hhmTcpEoQQxUR86PV2c5N1jcXZ0/LcU5CnWjG
nURRdjENZqRNSEhjWX6j8jNLf6tIG2MOOiEWbv6aRiWcDBB46lFI47ldzw4PPw/gOLhu4n9r8FRP
g+TWhVoWSjQCA5OisYbu2FHWn9VpaQO4a5GajOXsnH8Kf2OAFlqXwmTmmAC/W8aVAwwWWvKtYOMh
rG+ChRI7ZDfChA919RsbMUTY6iKUko4u2qd7r1r6M8KzrkRXyVxlTrVVJVWMovxyiqidewdg1WyX
rz0E7Dll9/VJj3fgl3DP6IRCL4Z7NsBLfW+VuF7e77bJGxWGSgi4qpnXvU/5lQMTID8TtuNnZwss
6z4F+Gc2CpANJbd32PoHB50BqHLZXjpBkw7Sjzhh0u8ulwHD0m17J1r8Ca59jNLI+cwfTRwoI0Gf
jYrgMTNC+XzZpZ8KNMYwI1A9c32Xbgs1dR6pxgiKM5j1jiQFVjNK1OyUqjTBHQha76hlrTAB20iB
4BtdkmIByORQK5fOgsY/6e8GV6KJCG7jZKBVcQfpxGeiYupHgDYm7gl7I6vpH3D6qxkCrHR7yTXv
QzkVZ3KedNZsxou1TO75lEW+8Z78u75Fdy3AEVwSOmXluBFaFaKFxxjsaR3DivUIOS3hOGzUYXnz
wxeoMbEOdeqe9kVNYYnIIpUWDQqQrigxP7zn/45eBHYx2oBDyvlSfVX5i2DCFMQCG/fKXybWUuZA
766ExxoUsKnD5tzm6CtabiL9NkcLxl7rGQFRqJ6+tvP2zyKVInp4kcQq+iSfS+2eZmCRovAHg8nt
kry9r/Gc+8rPQkROtpjKvoIDLx3F6/tsRfqx4k1JnsAlh10cJT5/YyWnjJ1ivgodkraQOmm0AlwR
mPSakQlRlQDAHgJzDWvoOT59yYBvHhM1IrA1+MHZt73+XqCAtJG2hg1MDmY0PCO+IsHkP0NDpFNu
jrBi4zgMqagXH3aNzeN60dG4GN19JFYGeh5fEPaDohzVIPD2L8Nx5q4p6qEw0pkkhClA2BSUVzwa
/p9lusfiMvT0DMnKU6FgoeruJQAN3oKEos36X1xCRXF+z17l1AwH4Xkw9oeHMa9/WbupiXyh63jk
vw9hGljX+iZV3pNAqzc5PSxYEVNgMhoMuh4t+J9qpLWUOxwElWmHNGHjdzgjAndtgdMuk268GuhY
OYvrjvwYrTqTDVQWMwSXr2P3jtxJYpNhiU3XorSove0yE5aKpuYWJuDA8FQAFPwKFatbhpxY1fkp
lg7xP9RTc9zyfVo0SyM5j0PsJgQr3X2+r3GeI/tEcCbB1ifus84VyyU3iuq5Xs01pnho1pGFVIls
N0xySVgTZB/pkQ+MfRr4Dpz5/h8gYv7jXH7qWDvX3lJ0DmYol1jG2nW3Mhu6vWurMKNw0kx11JGn
TUt1agcNJ/Lo6/Gjf4TDoyz8Y3K+53yOruH4e8z8b+RHHA9y7zH/Eoy83E5caALeeUqgiznCpqam
VKMWwRGRSjyztSP6aBxLKw/wsXTSzQR6dNLBtLZjc4qFQeIWnp8HfHHwOG3+sVvgGUQRH27ApeR8
Xyx7enZxalvGGLWIyi6eosiY0abm8V96ZqeY+gzNS8dPAM8yT5qYHTOfCMs4CgBHCoussMSXfpWp
wSSapWcuqBoJFIznLim7MFSk/V25KMNqAuZiG9rpXimk/W/4m5pXmzHOqplSZCuLnqpFq/X3ygKs
qRxCa6MdRbGFMFkNk7bO2ae1IXROGcsBURtSWeaYmpG7uzXAXJnK+TZ3vgnU2O/EaL/zs9io9hap
2uA44s6BjaZXgmlFmFlkY/WAXF/K6R1Az1uzyU9GahehI5xic35NiljmE1dhDc9+6oEZTngL7h5R
c6tKSUj2DKPYBc1Ik+MVjMLMYHwswO4da7tayWpmaYpm4Es4CYRlqhX9uszylIcPX/bOEvMKR1u9
glkAJZ/eHtJJboSTGdV3A84A4GM1kvOo3PqXVGUUsQqAXYbV9jjTRWOB7IQ+kqG7BusagN+uvTBe
lDYrYStVUxP+dM3gf3s0SfmLwzCPn7QLmrEiKY5frOHs3SkJGKX330vunizrfiKIJJ4oW8SDUsRp
WVR+OIb8qJkg0nlAgFks6ajib2hmtGgNMNUzmbo+luHfTyhvQeCysqxPV0XDziZaszJ9+hhxkCl7
OrS7Wv6z/4QJ1/pEBIkGTshsgj5+Ap77xDhu4jM1mjkLgO0ZF9HfhpvQViqLB5mbaNvBCnU6zgQU
rSABqrHrxq87hIVAMgB7s4FnAFHdkD/udSssiBri2S5Vmjrax6dHuSM4/CgMBrMXTS6Qvq+tAUB3
74OBwDzx27UCrCS/jWraTl8PGS/+JXAuqsQMGv5O1uwn/yyR2iTB8L22DA4b/UXh7ag2zaThvG8n
sDYQloONFyvYxSkCMH/+5gxItuqBm1VOVtEqwj4+QZfhYMZcfV8SZDCU4XSfLcurwv0DGE2ZpyE+
lN7/dET8+QKflctNVQFyaqY4JpKfrKlBwJp3M/blNeUV6ql9e67UJbQShoNH1xkdSC0rszSRtfGx
a1p+DHF7jGGVdr4ZX39UPNU2gR4PgDy//WFl8htENdBekCoQSYdSY7HckedcTXACw3fuGoN/ikCV
KHFC6GDA55SszajWJfyJbx4xSsgVneBwnyyBXf67ijxOKhuK4IA3idJTAhG3CFhdlYuvvP1KP7SS
2Hl6mPILod6CHJKH8fR/Pjb7gfMXLdco3Rw4W5aXJ/OJY3fCdUywS+e7JFJYBe53yt5lalQRA42u
Mua2uEQywQzOBQ12wAKy7i0AM3xTH+XjNBOT1oVUvvQWrqBrrstSD9X83zHdKPJg8ttoeixFcEQS
7xktdjrn/1zVQSfOXvYTjks5oy6Dul8de9LV7g31lOdnKsZKliiqXY/8z1U5vMrq5ZghgcxGOR9/
I6Z6VwIaoBw6EnNlB5tsD69dNF4Paex7WMZYMzGAx4TrjnCVEHR5eUa4is8KY+BmrXjZsnfrHeUi
tIk33voW7J38FbXuPn8KQjkkjNrgWpdIzicnIFo7nJSpTJ5O756DhNF51NMTXnmJOjZEdrtS32B0
wBfzaStdzAvLHbabiVkRKS/jNNowZCw0UW9cAhlXhXRWkHW8itSbU4A4Z/kszhToEkExtbyxOXI4
ArmQ4B7DwGzvipWHLzmjJIaDn2FDzDINfzGpcQ6ypnrpYpM11rcj5S09V2sGHPRgCHh2RojgM2hb
FcNVo4x1SV+k1wM+nhizNhDgQHjKlhuI0mClvEiKD8dmiCytHgXp6pUYwEgKoHLNC+M66uk84g/G
HXMcodDcHc5I4qntz80ClGMzxbroB10RW7ZGviB9f6LI/YD3jCxtCE605VD0waa8tvSdzqyhGDyj
Qn+tAtT8xFuT3x/DjrPot7/OXB+NocL6LmAZF3uZWVlXH+LK4WyyZwaGxy8iJC7kHRzHvwhQi8zY
sVmxUHZtnhH4xl9RLQbCXqSLYXZrf1g0DE7Xq06oRm0eeIdP76iYzMvwtbWupt8lXDY6Kx9ENgga
WWXfVuvUuUcC23ASw21WccqIvfdDQH1gq+zR7xgfWKbmsB2p2/gh3vMt23oCmD1VRUG8b1bih6/t
2Z0rXxdqmdonTrST5vmTiugPba0tPvuN9lAr7mGV+qNtDBSIqcsb0LgBSvgIvI+5o0UloH7YKLJn
XmIAX5MkT7rr4W9Y3N/LSO69TzffXkNtD0/hp+2xNZini6qFy/VQx1lW5sdpffvUy6IUQ91s6+wN
idGIHNvPbb8RB81pykBGh/WBICn9X39V/58ZA5XkCuw2KC6WF91eIn2nJdsngQTA3XW7KluVreZU
c8rRCaEkB7DCheltdJrsoj15El6UL39nDb7+/OYlNdPI+8484FlK+O9ihJjaCm0wkwReXxWgB5o/
D6HACdmDiLixkt4ZmGCMajEFH83LgKjosBt+WmfQHluTqJSgUp/h6kqS+WbOlBPGXoCb9Mbobcq2
pNMfAWlL7V3vgiiMKhzJ3C5mTIkiIWSlhiPZmz5p8nDDyzuMx+5jblsv/01TDq8IydrVF4tXZPQ9
+4aYhczcNMktmwdq5oDZ5pLIHfZPsgyLHP9czWcGQIUoJk2e/a1HyZaAQFH5lSYY8klmt6Ma/FSV
7QenyXUi/AJDlWjZh+G0Bllp2wbnMmhePwODHbaJvtoJOstOpTa8Zx6K8mYA5g+z/ise9DtyWuHd
ZATe2Nj1kHc1qfKMSrKyhHuO4w/8uZCAb56y9YqUb4tHoinTnyAwoOIfbg83/cy/pRW2qckZNpce
NZJCPb9o3mr/2ZbyRgzOOZu7UVuKPEil5ZdPMqIeH6LV3hC7wKww3JUfMbaI6In1ncubUn15KRiG
zzibinDeJTxVmdPpXpItPmYKYu7T+IFIyQUexSrLbsAPb1Jq3zE9V+vQNrFnhQvdLtHkblVouIeB
GM6oIOJw9iP//tqUO5Ou75Q1rdbxjfWW6kUR/BNNEbIpuW/FHNyffqZSSzryQsDycsglXZb0tWdn
k0mdpDpYhs4HFcQHkmVIw/3TcM5AwBnaQMUXROsbGILXX1N6uCde5dVBfiVcGL1oYKqGoADcuHBE
Z+oYltvlQJwrVU9sXKBpE6/r0b3YTZlPySEecSyAJCh3IKgwhCWyfi7E5EPFpZF0E0sBFu60CZ2T
HwzR419KLZ5GatO1R0yp824/3qlAXNf3l68Gvjx/ss6PCbY3Mti1N4ygSibe1DICP4ZK/MXJTFKU
vz5SDbW8ic6Zq+LRSWm0Ycrbw05Z0FGrWKHvwaxUiQC7F+gcRaXBTMbU3rehw9a0+l2E4HVMvte3
roHq1S11Cr4mKxOBXZohSJ6/IYpjdyNiWulXKHnk/IoL5sgwBvwxHG7oV/jlNoGstDXneacDINSu
y8W+Gxd/FoSOO2QpJUR6yQAfLR9M4JlV8HNhNdb0K8nMoauvGwv/+e510X/UKGftGFTxFxAC0Lk5
WirFHXgcgFaZWjdmfbmrttLzXoRd8HHT2koBFK8srXf0akYNu5KrRIZHbXjDYkgfcaQ8DV3BeLYI
VW8nF0RRE2PdWr0El3zRYasNSsTsUqzdxQZgPm3fTQJXhk2mbZXfGZDhksP2MoQdeBVczkJ02zWu
mAAKmH07Nf9V5QwMtbpwLwyWYW4DEHpO8spaMksLFgMNTyolZGq7X7+mcnWUv9uYeTA9QIkJlmaP
xPIK5HwFYleapi+n28M1d/KekqY21NXtHh0+Kr3jPIr7kv5S5mTKmox1EDDA/3KEgJMg4GjJAIZ2
uJJRwrdsCrraGvetbGwPLwp91ZWca5w/mMAOeiljCk/pyF7Az10XZJ6r7zCyhPrrgf1O/jICP53Y
VLd5zQeppbPaGzukbIB6EwnmlPAAJjBVxBlO3gHjrt92RW6hnPy4G7p8IR0PrYeFrt4fiYOPEhW4
pPqHwnZmBXXAOvw227AvWmUbCqN316zKOvn2rDUajKE3zked7de8a5NwKXH2oVXoWHx4l+sDFAuZ
oOEGyBkNQGs7b6OmqcdI+JE6TBdQ7kTX4jH3JrTInpVYbOb1u36dQcXFkXz3mUhj1lctOnZe16Gw
61eFRLprdJgjdn3N9jrHAb3o36lqNz782VsaAd7R+bk8w8gUQPSZHA8Pmm/Gw5BWOP1713ojxtI4
RUkL4V0y1zPomnReOI4YB4pZCxoosHbTAXBu19c1Ag+dVV+3iVQUQT2vxsvJrXsoedGksESk+qPC
zl+/EQaBJKZ8/XZSO8f0gKQl9nEOPvFSAjsI/x1ilW/m+Xl/lSSq3n5IslvTv2qB7084TUvMllZt
nAlYbOBZ4BSdWZaotni/m1PhR4YtjRjalQ81Jp0pSAVg3XHlFVse01jGQ/pNVCrX4GLf7+tRXbSR
txoZ/FWNQvSROiuQx52aIfgZx3XnTBJXIQzKtw3voWwCat9lV6dYkpDznko0UEwzihlND91a0F+9
WRR2naKXK78xwylGiS9J+OVfKMy4uMFTkWwwqGCtcTOo1u1lxtYUDfgO1zq7nuZQn+PNUgeMhFlb
QIpthRMMc1l99CFVzWdo47TCAEjdiZhRiqZib/nNarxfm9pItFWnBGqWhAquqEhG+jyja74DZPST
CpjjT6DXtxnPIL5ttRqK1aBgSUJw6XkKPt3EosGXPluncWbi45WIL5rJSnKc4Gz+upjfAZACvqaG
DBK/GBAPozHpic9Em4hR44lR5CgBb22e4MUDPfaEFP7W9l8nyf/UmUo7U0KRFpLgn/+ZEOiB1wSo
fLE/WpSHl1rdKaHf4tQEbGJXsxS1C7WvLYslnQF7CGphlEI3NmqE7y+C5NKzwEyQ49s2TQDOmZT6
QOWF8BquXQDBAKvacONvkoi/1HZbkD1zU4fAPQjcNJ70WNrdsMy5+1wAi+z9kT/p2JXHjixMerkx
tjdC0iIUuXDQSRNHGKFl9Y/okTozW6PHAZZnR7gYbKVlxhItbwiNfljgV5LwcgJBUMsYuBRVpY3z
2DX7u5gCZA8qnhK0zagnYGor3LQFmCoyNStyPXzKaUEGcOKyDcEMeDLQUMr1GVNhR2fX0OC/4h15
lz+WuJ8/W2Utz1zKjEcQT/Ya0Sfc05U4PT6xBH2q5rLpGAFYJhOciJtt9fyXvDQCq1aPzS4CUNFx
Rah0a3Dco7q/gv/kLc/64507EcdJKmmtFhxM1YLvSlQZGh26vZ4BaA7lwsM8ZSmB5VQ6ui35jXDJ
CSfsgZHCF7hGVUoYMru1vglUftynRR8p9TaI9Si4AnrvdgLWwEeApqW1zaiiySIO0IXZKXHHh/uC
KPmOF0AD2jZ4lLnJdxkdrOY8qTtlXIYHqyopWWI6OR+bD58GfFEgew1IsHbNWXMqi8LVudTtd/Rv
0tdi/QamHoU4fmlJ+pQtVzSNdlJbezgMEvibNq+4swPE0cCkkGLHXJNlYX2uLDkDpHlb3xQuIVc9
SXNda+Y8g3VRL49QPNa7Gsgu44me8bXrASxCCyIVOLNimKWgFJ5SlyPsj9zr5DlqW3nGFp8Cm5KP
Kk1E1e57IWlEcnnLY7qufDQg/+EWcxrG1zDwn3QlxQopKZGbupxvp83Y/rfHUKfaKfiDBVr0+uKB
X+uF3KeecSxHS7F0pUKwi0hdhmH5Vizm3IFo7mPoN0ozY6QK0JMxd/GkSm+YLR8kd8OsfAx12cK5
oY4iDuxa9RzHb+i2+AuK77/u2gXzB/6hgIm7x9Ge2bJoQI7KYlCqckdozJx74tjK9ElluaA9oP/D
xT8fvcTA7DTgudfNBSxZzjoNRWpFxlcORL/9CGP3cciUAchoVY5VxiRtfqnBdJupsSP3N4GfgrD/
YK85+1mt4182xzna8XSNIZChyPPOHg/5N3HWTkU6ZVjKSZjO7NOpgAo+PbSwVkMo2krTNLYlhY7M
iB4IF1B3kmCyvliWWFfC1ZdJjjmFyBBEzy8gMljStcBNAZdHv4yLf+TY9qfSCJkrCXJfTzgGSSxu
rKrmtHf4F2ACtAjmDCvMfdXVv0/VR5i55F024x1oLHFVfy5hNBtm5Tn4GBGrPqL8MGID3a7GOk22
ebTvzaGrPFULnFAhW6OGQz7HvsVkaptN/KIz1HIZCrB2rh4o3p+SncUzze8cXnKic/Ilyt+cvbz9
//vjxazFYcNLqjI64Yh2XFgx55/IEVGKwAW68tVF0FpmV3DgVa4TC7ppqYIshZ+PDWZwuhilFEbQ
V6m38a0d9I368Ypn8pSC/2HdFxg2FOqEVlV7j7jKq672R3TPCm2+9KKJwqOXABTjsiV8Jfs5X66J
YN6j7czGMdbBexuEHrs3d8MB5ZlIhrs7WiNLXjO4EONbPuvYQl1g1nmdkfi+DiW+vi435/15Uw+C
Hs5LTdgPzD3qSHapmSOTGtI7UZ45xxsLGC7prlfx+6o0WSaGweEtoVno+2yBBRsv8F4Shn1j4Owz
rRPu8u79lFkXwFijoGVWJKYDz4BJZbJgtxHVtvo7+T09FCGtVdiFn9f9PiBmxOiJG5Kz6Fn9eVO1
t7Gk2sKWw91FQPICubXLbGoKptiIq7HScgBktrWJV3o5RuulGt95SgHjkT3Pr8GljTzVtlSXupXW
H5PYhP+AvnnlDLbk4mzqqyJ4u/UXl5naXZeZnxnPkJmmb/Mcda7ep7LFlhq3ULbyu6FNm0yK0OM5
T09fa2F3LHs/gyItdXe/wQI80+TRIqWcdht4S+Oq+IfcCDaNVCgJfNdNi+DmxDKCtVpHP2kLPR01
WGl+5qGKdAxxZH3vesBuwSy8dCxcCw+HgyfzkDz8vGXLkeCY7d9LVUTddCvs44dLRCPh+lHvqNG8
7BuB7RHpgyiC6Y8V0SfLGltarITmI2PF4SOG/XbA5AFVEUoZ9Tr0A7b+mSjMLhfG6ILPFz49K25b
S6mJPTDYTolRrZi+G3YZcPCVK+h8afdGYUdAwFaq9MRcSTSPb2YO1UwypeeR/58Ct6MlMGqWw0ec
fIJMecWVRI/zrNnIu6lTLjtfKg1yvRtjmxQZaLbeAuypJXYbpCVn5HGDtx3wmpC6iOLC04tk6T0i
vv7B2F3tjoDZfxv/hgjkZ0iqS881rga7EYYKp0pzrQZpOfDWFF2ST2PwIAXeP4RZm4xrDf5tnAKI
KtWAEqktELb9HEhOaTAjYnc3H9esv0Y1lbgqaTL3XGL+fV0LTAxwqCOPQj6tBgytjh55US1W+axI
UTsQ6JeVo0iGfAr78qRC9wEXsjdJ6PmUjmIQ7MZsXVx9a3ScjTxxPDcQB6lQeJoFAriQ/TYkC+Ui
EKZTkF/6ekUnXI2Bfl7miZLoRVxcFmeCaHUceqakxvSxm0Eq0qvCqZ0dJHQRqF63+AxVG1x4amTH
nKuqni2XGwjjegxz0PZro5f7d+gQ545RjaST4NTL2cvpu3NS4AnblwyD4VVo/BVsKx7RppVK4co4
983+wmVwTTvfYEBWermg7HQUIO5BVT90lMy7QL9PKcqh6GNKF6HPeAGucO68eABG+w2X09+Nioul
h68/F+IzOXiSehU4hX+lq0krOKFOjJyQUUfOD18lrebNbb9LCmkpOIHI8JzbdFYl7jA4rn74OBVN
0S7rm3+9e/ab6FBmQZVHexJZiEValLRyqT7NkR8PALtYCdfGyDX91HieiwPrkgAHbpvmndn1Cm7r
mH0uBIZTXcfHv0diDD3ztl/k0VpHL/XRfntEIHFJJfZ1y+9wg09BKeOHjrAEcLoQTWFV4LokWzkL
SQEvxW+DcAnxpsxpFPK5M75HAflC9TIB5V017B4Jef0YT6CK4koxAzulh3NmrKP00Oz4mBR2bktW
3Gjqd7b9zY353LJR6nNdT+P+wwm8a9r0FkDVY803fOTGrxFDiG4p3jGfqDN1NegaXMXmCkRtTYDE
d5t8zr5GIl51Hby46JGBUvBA4FScNVE+rXYUbtACdIv69eQpAErFM+xbYhB780w5s5CI+cw6/MM/
N3gMDsRXoVZV515eed60F3RGfS66LPkQCwfk1mOvUf29PYmnUpSHqIZObV3AAFqYlexNrG3fLK2T
mHVB3CmJ2Yvqr5msEBrQp4aI/MO6UzA5pVcsPCPd5FjANgsr96MgipumVqbzOVCcK+KzyY6e5rwo
pRofaCR1Aga4XlULsvsg/VoQwzvAUPqJ54KIU6yY9WkWC8k7s6JdkRRqHf2LZzvZAaNwQj1Az16h
VzFxeknzyJUeoLY7Q4tFMMqo4KDZaZwlXqtLIr4NC48EmwET5wgZMYrM2FX1OGS5Mxq7XQBnRbmn
W17+P35OdooJHtpEggVIv4DQXF766jkLJSQ+l1J20+n8qN/lH5aTnHi5E87LXj5S8iPN8Lrtsru1
GfBGsL5LMOa1DgC3OWFfD1QJpJ+1qOW7sgIu3r6VzbVBbw/5ucJR82MSLNcDQIEUlSajKX1sE7xS
RaUMsmRu/84ipab0nA83JwOR79ehxYAA6ckIxAeAXraLBcYdeYx+5x+DWNFHlrl6Fxgak1QnyvT8
HztyHKjhabN2KQfYhQ6PYyPNikhZ/xbS0JDn5RtDe1UB14slZxUxr+CQCnrPduJVIO9B+3oTNhMo
203unuiYkPXX7po9ORhCHFI+77ek4q+UbXxubb086XOUzhoqEK6RMf4QxPdbJifQ4IbMBDyVhj7x
Ibafw9ONxjm7Z/uP1m3kbDpCYlVX3IMGXLlNsmRCn2yiicwh+dlfFpoxAu1J+wosPOG2VqOZdVdT
zKBHMrzWFQei0i2o8ISbGWGX/NHuatRjIPAhyIDgnsQfXMieRvkDrSxhndZtQlr8PDGwLOs5CAwc
Q1vJf1ybYgYWFOxUHiVbgOQPgxqrdCgRWEWugRTlzcBLl4/qiwtp7rDhRESNwbQg+h/D/nz0juLq
6PtqmqmAwc9JEE0WOOS8i3kfU9K7foyimzdHTnINK4CuqNE2q5gB/iiFMa1XVwE+D/GIk9B7lbZ7
L9PcR5o6rlkxHNV6YB9BPz7eXOPoD+m0lejxIWpldPbVDEyYAcWqo/XxzILA6ZpWbTxdvuKKdLiK
hmjYhpHDQFrA3Lsva4vu0iyCItYeBq96bIFc6Vymm5SlE30rMp8xkO2O7dxUZAVMJ87mMci1szi3
qp9+ugWYOn2/jZgpNc9l9Qc+HnrRMZKcHJUT9D+7CzZ6EAqBD+sqoKlY9oK39a4zOS+k2/HbgRdL
Q1Um03aqaV88A1KO+5k9OlEdIvoWzYAAJpIgYx3QyqUb5hB0DiJ6htIpivQvN7LiDToEvIUhmig+
Z9ETaxY0ESfAeTkF66snrXf/+cb+K44y26E8kTYKQyMya/+ws/+wJZwv88dtKYfNheNngBmXOK7P
pun9Qm4Vhu5Xc4JmzfiRuGAhar+7uLrNh7Dz7xoH2tblf56yyM13MIldfexupmKEqjlTU5Js4V0o
5B3Qezcvl474r52JYMBUBuDMn+sutpS9MVqhGTD8Iqc/A6FfY3upzsw8jM8E809Rtlh1Z25y1jMh
QhgBkn+2x5iWQZQ76Y3lrIQNVVtZnD6irqxlvybJqeQxXQghJ+YdKB7nx2x/QJ6/xEhNXkZT7CLj
1w3crJY3Ksx9CYwjPoc06TpNko5ZznByc8VhL+KchetSfnqvI0HgR1ivWJyZflUt0k79/M6YNgIv
FrA+jUuqH/4aOLQLUrU73PNTBoGFRPYplqzdSGp0OuU+OWIPoF6ZgWsi6VHkq9NyKcVoWkhLyGDT
sqd1UQfIbsH+1L5EgwYRtopydWY7i4cfx28L3tbxT2h9TOO9CVMSs5wmua10J6bCrveByTEGQuSa
YXZ2uU4tNxKBzq02A2drvE9WUi+QfCPH+zpzuiWpG84hyvaXrH1fOBh+P5iWfzsNC22yRSS23l9/
ZjQF+UM8DPNifs12D9cbOu4nufyDkBpsMg4Med0PElq6ntSPUamGvlefILXUNnq+rp5CV9411xVT
eW0lQwiNXc56V2hyqt4OJh2I9z8Nd6PaAUkfvr61THsxCLv9ehuw0+2My8YvEP+JorqrGpry7hhc
Obnl/BM3yYgRwRUwItQj7JXh65iyxXWbAjle6+54+zyKMaYmKJRyi2tyRqVfg0N/h4vNqMFPMQKH
DUH9LjWq2AFBVeoqFkq2XvTjiyleiIVa/31C0Jq0wL4CQH9PwJdRw4FjMotkd6hsowJtd/E+zCPz
TRRYBlNBNX3h5TwAi8+eouA2ci85/N0mWJ26SlTi7t4iX9RPZM2XQ9zDwMDA5h3LTBm8gqkQowU0
oKai5+qkeH+8ZugVtJoOJwwGrK/7XdK2lres+lktuXMcHyPI1Q8Vzg0m4+jGf1JqQOl4APIexMNv
aApv7hy9ewwmkRc/c1rVdiwpxmOHMeogWFz6G4KZSpBPw6ycHT7QRjtmoAXXUC5YEGsZUgtyZt0g
ArgTN2icgRH86NUbcpqKW6u33WQ6PBKWKSjd9UVE2OjwFdFqx4HYUL7A0AaEdzNSXRGs53jYrRmr
nkKEyTn8J4hhERPv2ELy4oRasTNnHVz4/CiZtUr8+ZN88EH8uysmlXTKdAv8petfxsXGrnFY8ket
q2FvGeCKogXqiDeaQOsVHNehULwY8S3PLjo++IkwmWhOsFYppZ29dHFc0MVHOD2DWInVo4mM3VZi
tNOylOBvsrTxch45NzbTS/SiV1q230z6+1E4+0JyhIxbZBPpqrlyIRdvY2esmkr+3jv50hJToqRk
q0vcUOYXyFNz8qdU9iiQB0KpioYoPniQS9zxexk3TXeUhaVi9YNZG/5boRJK/JIJTSgsEHVOoobU
wWtA9ueldxlY6UN30hq50id10cFcg7xIRTZcRNVQZGqibFgt9wpd1o4GvUkYJqkBHpxW9qaN6W3A
h+7jw0lgZI9vkYTU6PHLytRJtHvV/5qZ6pguJ8ji6EmJ69kewp16KKiGy1fSEPB5Fx0y9I0Hdort
zPFWpXCx79Fb+mNIyx+UeBACTVOoLiKtaSWi1dqPKg4lgCZIqI4ESDl1TCSn2BvV3YM5YdS4uHuC
ISLUU8hlSjd7kVts1UG58V1vlbGRatooTLzC6C8tr9VUz1u7Q2Ru/WwZj0dBhpyDU0ugjCq2mqbw
HG0of5z2XDA3gBjyjbv0fXZW9YaJ36JRikHycI9DLkuk5+EYlIv7nkZSVHmYq2zklc+Dqk7y2xti
0GB0KYc4HzD+dIikyjf5dSyDiYbWo51dOjVfDreh75yOSrITAnoieuuDvqtdyw8kVUp+ylXsAWiG
DdqPaXqBQ5VomJputqXrulYIBH3DT2H08lo8R4kaMZOcXRAmzkahyd7vyWQbC0wJ8TgjO0fETMea
6Rd6HsQHaQ1XGwBVa+qNgMbkWDNTrGiCyxT77tlfP+R/HIokoT29CHCl3hDAp0ODWBWjpDck7K3B
hy4MmAVp3MbcbYcKvZ4o/L2q4gmd0AbQKKx1HrQNrV1NT0O+4BEGLrqo4M+Eaj1bsQ0R3VACnbfu
2QJOekzAqg+5CVo0ci6Hr4nMYyC4AuWLaocitDAOdrxyMsjn+2lW32DvyzMYv+z7/4XAmfeuqHUw
AWObt8+cUKUUVEms+2Tnac5f0BxvTi0SPfVN4Jd/H3gixpcRqdykaK2SNbSYJLkJjA+jJ9FvyANy
P72k22LVgF+ZHli1poYQ8ge/8VfCXoUk+OSH/Gfmc6a0CosvuVJIgXE8lAfDA77ZPdm/DxsHUyRo
byV4zYY3dlBLTFj4JAiQA69W+UPz4cRkl4pJelP0gM91XLash/35EH7YFwkDT+tGHYOCjDPOmkkm
T+q5J8Or7vUQG7CSlAhQlQtIQxz3zj+0CZGBSKKRooNisK+jtydjhoSRc0ORUfuQCNjOnUm+IqLc
eqyV9FTEpSI1g6FCwScxHVDrPiyue9T6ZDp7dt5ARIgU9BXK+WIVrVYRw4bu5an1faGLc91P93J6
N058u4ztEHT5OhJ6u3Lf8BAPrY8GAwkOX+ZmWbvFSyBE8AEWXXasa931d4Ygi4uVUaNBFqPwltW1
CpqyVTlBniWLw9a8MiFsOqbsToZOEFcR5Cd+jn97VOaWhCkeJG2AMQaQSmYYjtObRrD1uaZHzH+D
VUhzRv5gDQPupZxZ1HjrXqSPh5onQiV6jC1HEHTwfltEuTZhdKWXH0OYi6Z3Xi3IT0S6xe3Xsw0r
Sd3zFcUYzAWM1yuMKdYNPBa+gG/McQzRww0KKw/IY91tXuQHML3td+kUZfMZVyGoIbVxT4yVWTyn
f2RPwrp0tPAS3S8auMe9/Kl8mGAQAPaYPPGs68noNMRwbJ3JVdQNvvr3jyDG6GKLtCBWfkJoyVUg
0cJH8VkEGJde2USn6Rhu6ej2+omDL6XR8M4sq6FI0mDNaxdLRYJd87li9UXbgnzbPv9ul/rvpZV6
nzkaA+QadPIixA53+tvunIDWskn/QahNuWnCl3Mk+YI5l6VKWACXZc+zFInPxz15WMXEWbqylyzR
mRexFBDoeT4zyJpqvKDZrucRqBZ5bPNdx3eBNRxxxpAOhpB4FYEafVfOVGEOx2+zR+Yae06elwGa
VCc7j3EDhJOc2DWtBZskXU3+lKi+mZ7FqWUJfAA1GF5ZwNhAHektM/wMyLSuOHUs8ZweEW+b8m8S
zaieDRIPww2NVRtRDVUvjxcNhoY6H2M6XgC2jmsWdTHaE7cCOENM26pvToi/Nrj3GxgWeL1UFYYi
WB16FV07N7zE10WIaaTVwl1SDCfZjHPZj+gxkoOC+/CMZGDMXJMSA7fW8cxDyQvuq4hvCzUhin4+
0gywOlqHYxd5PFykIu0+rgO0tVjvrI0AwiCvPSHpkkssz0FOA55ZJi7ZLEVlnlRO/qwErJOVbbKh
YVg92NOZY/Cd6zhPq99bNzztRLOtTJ36jVkFjZNGEfSmEI3gScaswiHCHTzr/wZ7BN3tTaVdp7nb
sB0rwgDQaoaEC6pPWPnXWsjpHK1zX+wn1OAFkM72esLpBr0foWNGauWPvBytx+QJ3YFyU2yPdCDK
jUYoeyVXzYDhYFV5QfXtP6LGIkDUUAjCyR3tSVDeBZrU0mIKxPwqpmmJVBTLwYhwBMs8piyXpYUL
MYSbD8RY49zMvhZQXZTYPQ9WW9flFWGRSLZKfCeIts/ZiwjIgyMfsWPwMoeews2QFu9NT35UzhIb
tBRr6qns8dAE08IITFXyssgfm6/2v2QE+nRkibQ7lUH5KF7LYQwMFcZ5QtxDWihKSz9JmzyySkX3
SR3fZwu09UAZSv01YgcWSAUEZDh5hFEeeYTwlcU/LlgXyfaCNH3ZXmxybP/oV6yZf0X6s0vP0deX
AW9g1wi9+aHxWNjFvCmOUcT+MmWAWX8MwVci8HEGFEmC6ZbWCLBekq7tT6NNTq3Hm7rbanvO/oER
bOk6UYcQYUjNX6RGT+rrN0PBZWKbxnSmKbp25MGv1tr3oVXDbkZkvpNG/+nCw4slmRXVsgvqwnK5
1OQnzbLTbaUvIYn8plvF5n8hYUJ+XsUR3QX0kTxNSud4jaUGA8DtpoI8tW8eNDE5GHKQkEBENDbl
Ic/WRX5CiPQLFxnpYOTPJTb0TeTkPiA29y18IvdCaRI+W89xBY/BXZgsT8Lq5ZGnl+q/GA0O8EFO
is/+X2/i0ohP70gL+v3E0ss4eZ75laA38SLYdLM7CsYau1orcC+6BRV1upi4w7qTlJo9fA8favON
optMlYntjH7YlrWD3H1+CRUZLhvA+QcC6FB9zO0IxQ7Ah+y6Crx3Gbes0TVWGa3j4frzUQ16joBY
2GhQoPnh6chxh9xSHge0U6um2aIpDU1jdzN3DzWmNFvTe9JzuhdRvs0UazsJcHABXJtHbLCXXmGB
2so6m6asnFBZNHsx/5E9rt5MJqHf56e8zUX8Ca/D6LAGw0ltWixMwER95yhSLJOiefyrzrcaVyK/
wH1xTtjO8h4qLz5FMrqfiWC2pn8aNfm9r9ZYu8smeYZMwmh6l34ZmKt+kvQTUjJ6vlfQB5A0RxdR
aIYGbQsUQEvVtP+8LUw7r6nY/rokvYF99Dl8YgDxye1UYbMaZsaREkOHWBkBdHwSz47lxMr7LGnL
HmT0ln1B70ZN2VC5jQA8QSpUa6uSt2fFJKN73gQEXDOjTD3WeSbhQOrhDHWrw56ME/u2LbuNmIUv
9UjTXik23fPAoest1i+EIeFqkGMLPD4goQfNnRqtKg9jd8+Yx5QcaLJ1+djjfJNHkdt9BjoGtPkS
pVQCs0lZY8ymTdHGNIF5O4TP6SzCfDFxdsRbqKNUpJyrhCXNdF1FcvGadeC2u3fQMgOr9EfbbvAc
ilE/XAtNNnuoneYUTfhOXTRST3hcI0wZm0ESUdvr8DXPM8LymO+afVldAGicOd+Fq6hM0hCgn/Qs
crpdZ2RXHJ8LoxiFFVhSUMUjyJKUfA+6v9IKZzxS2phdK4DMeXkK6pnTHUcdeMZtRllWHou/xPYI
CEvXda0KYlAD/4pFvSa7qbZCkrAkm9TA60qRWVmYRtTokI6N3F1MC7HXTmBHrM5yBhOSPIC+417+
cx54Agrqt99LdX5TssWTT1BqO04ngrmLbLRklh7/blInBv/CGZvX9NU7ezBuLT1NFHWHG+0xDMnZ
gpMa3D2drlv4taimQXcDrCQ2wFyq6aFn2vAWEmbYtwT+SJQlUskFviz0o9VJBfjQZaif9XWISg3w
QvZWlcMZvFHmCdaJII5dBqBL4guWdYAB3WMhKRA8M11hBYJcq71jzN/k8GRBn4q5U5V0uttOebd7
8XTLAyn+uT7B1hz105xL/JhVu71m6xJfQd/3uHxc6Z0pn1begk9YYLlamsuoJZWEyINCM2tZD0gG
UTUksctjKj6Q045QSj7GBlT/12+DbngnZJKbXiwIihiQsYsrJELQlOH6Fo75GaSS+DFAKJzy1GD4
nSKXyezmUpPG+pqu8Z0aUKNGgmM7WZbw6ec+sIF0U2EkRPGgxwsDRoYaVVhksbZCs7Dl1mjKaxm3
8G8EHporOrnFWI0fY7oz98Uz4fiu30+IjVbZG6DunXKzRIgLjH9/ZnMqUJuQK4sYVC8YeJUJtJtV
rhr4uxbt2kHau2dS75xE/62sfkIZwbrE+Bj6ZJyZ7ZvgcEizQyR3Kv85VhamyC7SwFM4fMLLkFSM
FMjPQsfMLVu8iIdS1Xpliu+jy0cqE2EF1z7s2rfh88iAFOzaMUq+bM1apLdTEUtJUwgaOatdi66D
PqRQ3uTUSLF07gQMps2wC7OaUaT8f9QEj1pKN92ZSM2Ph2h3vBMeMtXONMkkMgGCF4bkgTHplzM2
8TdMWXjLGN07TzQCjPGDjEUxv0Wpew4EXhvckzthvwEihOXLR9C4D1D9GKe0SyNq+O0HJ7ZaBxsk
p0Iqxr0IBuzSETYVeKCmkcmA6LZUllY+jGjqWIyrIJdla2Xv6FfqJHmXhj5zouHsHbkDk9uaStIO
lmi/Fr+Oo1eodaoax11DPc88JWmOPcYiNQRuUtku4xPCfkWiChJ/BruWdaGYQnBQWb2DzGo4jV+E
/KEFo1cxRyaT78m826fd9sGxrWQymL51zvTxXT4v7IDT1tabupK6o/kVBSdWZqFLAZitgu/MC2QY
GQkMlyIm4oM80eFMrBUVZkZJWhyLXm82toOeTseqVkPby4AkuxxRL6eyBQwY3sX5f10DwIhkG4En
ThKwuWNi/LQleWPieVhF2UMkCUpXLBm/PXvvyYL8w/tqfE9/+p5q/wHZylgZHv+gBPmLCJSE5Y+X
926zrP+Fpp8wsbNNcSeqTXKoEsgl6XzcbgwfLnGn37x5PB1Yxn47hsWSUDLmdajMSN+81+74XEnb
AdFcUgyAgQ5RZSogTIKcYcEr6cNmmx80nXkeW/WPyPFPRqbi34TI1Vqzgu4i0I5gz7k6DiT/DADB
hWA5z/Tnbd9BuKzSxXcyEUdj9l9yqLKSsznqeAuo9Sd/FSwpMrsNycdkI/RliBmClTgkyHPZPRNe
R9u4g1XL+zKvBk+aw6TmFPvZmz0YJzRJrwyNkVOSPF0dNULaKuhBiCA6bE/ARqT/wtzxzeELg1QF
NcgyVZ+WrGjol3nc7+ChJeuo1ef8W28Z3YjPd6YByAi7lapHCA0cSILfByZSeYqpoSNa+UamtBu8
/nwo4ctHApZ8pwoDSQgyuzYsYAxJeNuTe5wtYO6CBAwITOSVDlKK+5mwuM2LeBV6hxXd7lVwfDaQ
RArIIt/HT7fCyF4hHz2nafXMmTbh8WryzBgbceA8Ivgaig/Z9N7FBFqoWDRCgCCIgEME7wvDqzm8
xh7qHVjLbI1zW6cXX4/Iy2bfoNdZg1y9e9jhu7g5dB6J2wtZYHWJHOD2S0yrqa4ODVSMqMBeuhPu
nfTh7KbHkcbYoUCw3WZY2TA8QgFmMRknpKy+vr3ZfYfsSh91B9mUyLp4XHBKIZkiyizXp7BxlwH+
5P2tn0+5xxTykjevlijxY5sklC26bqTvsvBHh4SyBPS36T8LE75diTNEP314v2HvBY6++9eItIj9
3Bm07i7kAS7HDBK/cdGlpjS83KPAPdTmIZvS+utZ1T/Osd5Papq7c7Mv2y/8UKYIO+QTSR7BQRTo
V/Cpi+/3VDsEhWL0xvbOlAiTvuJ6Mdxz6uG1m2KE/ZSZo6G96WexZnnt8ptYAvliFPJUIhdZLg3i
qN4e2f9IAQ3ec6k47FRMej5An4jW22yvVYYwz4GCdwifaq/YjWbA90cNZKIUHbcc2Hkbtsok3zyI
ylh2SLpFA0cA8y6PuC710//tYNKrrv+aS4hXcUUn14HNrhvc/26SYujBr/wDAlNOgK+wsCGEPjUn
KegY4bDkRuVyZ9JVmBblXcPIia38WEmHlj8m18vBHhxN9m+8mLE4x49WfttNfBFyS1g9eRx9rBPO
cCexzmtlTmd0vmKQTQjKznlXWVhSXT0q/Y9h2wHHf3Jq6U5xRLQkcJXsnooO11eJevLryqToVUnh
JdQML4UgufFBRZEkqtWd3gJzP+M/nlNMnZPI+N+3Y6spcG6rVmhoWxYso3njG+VJUKNam7+0Cnyr
8ZnFcPrDg8cjiEPax0F7F9q5Miic3eRkCf2AcKbmVMCYIXQ+0RZu1rry6mpkv57BjyOzOknOo+Ty
4XGlxXyJMsym+b5LCBGxpFjV5VNzk8SQEeHCbB1yqyMlsqAKI9Dryow9oh+8dEwkTd3Wdulf06N0
2ds/toS4h4HeRzb4R/C+EtriYB3p6cgCcmadgNV343qInAkPUXVXllVVSrEJDjF4JMDinJJElrHm
yRQh2ocU5Awph/nauTxKezHZkPv31LHmYqlDGnQqG0T4zYHhqYteQSlR8MNRQJMhLjdkxvNzpJQ0
A7tZS7Mmdr5oHJYJZboX11YXx9Y4hxSeKWShYplnSTSaD1rBUdRn4uo6ccLBraajs/obHaq5n0eE
3xz5W/KuUpVekI9xuHYPGamSvvolEa6+0mpKJbvC0ek3Uhep/mYncmzdkhGAC2HuoEAqy7gy3wqq
EjrX4AVxFfZf13n3ANA6HN7Uj3GMMCoD1AxRT5KU/V1eyvEFLPrTaFX3d90iZeih3USGNLjg32lk
XeotKnbMRRy7ZVIy1OnGzt2QdPnP9HZtqDtmjR2jEIxHEPFWdnCahAmC9s0CYolM8NTxJr/nq+Pq
fTfpRBk4YiTZ6Pf5nhZOKt17E+APKbwHhSOuoanaMWo+Eohh4weadB3X2JZfgZzqAAgJhODPeoV6
o5E3VpCQTOChHcejrB7VwMjC5+vy29MihH1yxb6QwFsnZCrF5u7TAJPMmS1b13AQjQDxDtk9JVmL
24bm1r69j3zxdePImiUxYIJy8dQTKLlhKwJ1WTu1Y48tChMHj+OqrPs+SkIt3PGv5V2DK4l4EcdH
XXNcs7pVg1JEAdi/TaCeg8+WArzsOH/PrRwqDZ5BLJcguQKOG2t27ePuFJIe80Ekb7MTsIrPs332
gJh6l8USVqEuHs3ZT/kiKBe9T7MqCiZiO0mrn6mjAo4G+rD45lLwOOFVAQ6yCwI11z5S4JD153Dx
5hQHAmI2zlb3Pij6cXOVUyD85KWAtW+YMCFJ2um/cNce+0aJS+Teb8vgrDyruXlTXKfj3P0g3PQP
FcRPEXxKrrp1FzWGQ1UF/j86eb45UQJfzeYbPn1Xa2kVWKCm9G5SEvIoBrgfV4Tra60pVRrG5CuZ
662S/X/aBWqTxlR9Ccm1NI70NELJQhtMiVkY/GIUAIRVJ8JuqF5y/tgFdawSlWWOcvMBSgguotXp
BtGaktWYdH1/C6t1SOf6rlyiaDJw2C3wgAW0xD9wrGgjz0ZtLW2ILxlKa4rAC3G5Grd9fWJClbNf
tPOPSLv8BfRQa8PsWw9rnwsw/YlhsA2TZ9hS2kRfRat+A2GndOG8l1rEnl0DbTqcPL7jbSo5YSOV
nfElW+77DncB9f4KT8uC9581cTDglVF+asq3/1NAfBLcGdZO3eBqPwEKpEZwX0/bdM1s5FCr2XCv
Tdq/sLpd3WfiBU/o9YzgevkCL+ieZkTcCSkWz6YW96Oa+Sd5By5mijzl9nfjUGu9mDBGHvKBXZlC
hLgYRaR1x0gpOXYtFu4GTZzRnjY+l5yPOWANagPR5eJyrl7Nx6IhMQaa2gdM6zlq8pMGBfFIJNSb
2DC2I33//XvLh/AeSBB4wi89ibyUBqPnRqhmn4bSum3wkeGjiqj7l6wWFvC4AZuQCnGLuGsevaCI
sOPLrjevt6LFAX658cj/zZl8GNfgGDknog37yGcmT0P2F+U5BAt6IoAZIoxRps4gBwKCERZDftWi
v8/d2l42FmoKE9M+GL+JlhSaocTS0UAvkJ9cVKSTDlQGewmUqdqgzi+PU6HPI95DSs4mvOD5q4VZ
X8MVQFUsbKRMX+zhnX7Qy2aP2C16KecABhFXVZvV0E7Mt8ICVXTolkJ0F0tp7B1mhcvDssp7FqiZ
UwttJtjvwZ7hRfyZQW+qSuis/S7IqJt35YvLwbqv5JGRx0enZWDjNK0+o+0UYZ+aQ2BROIzSkFeL
pFqnd1MbVSXHBkitAulmCT18TRjf1eNOHwB26yftxslPK2b+3WHXU/qiVFIkzNpDA++T0Egd6Cu4
hF3TbZZz/cijjys5fzQUEJOVkh/jPosiHaAzz08eVzNAaTJ3G2ySuBW3pafBg3+PyfWVq3Ey/qOJ
SP28Is+HJgdKJx0eIpw682LbF5Csp06nI0qQaHG2HXr/YUY/4suBUbSIpwTayK0nLotEcq8dDDUH
dHq8OUedlGbx9CyA2Q0cudqrCWArGnaxus1iuZTruXJuvhEMFD/6r9aEIXEDo59QOaFWs9qiv5c1
Yos3u5WqvfEP0qCfQ9LgLg6ZMzkc7eUCnewPREkFvHhUIolbWZzvKV3J/uiS7/eGMFGVNyfYLnH1
dIecPlrvxCf+AYUQ9LolEn4l2KEuTgM/8NmOuWnXU45pTQvAOxeSxMULKRm8d1aH7JsYj796QBvX
8D6VVlS8tOXXb8/QW0JwW6tuvesRC7x8y5zxIrloq6yU4XFSTnJ9Ktc/n7zmO8pVdQJY7yfZDDZw
1U2rlN5BN3+JxJk67zM8xjYpdtcwBbrhlqS4KwnfdCMs6gqYcjM9cPCGeOSXng9jOsTfyXP45S47
Lajc3PZOvwNKU4B43LIeHWkctJRA5g7qlNJzNz1Lb7ywh27Bbfb67/o6rg1kNCPTOnvlRah5O35Y
0hjy4GtlO0VmxhbEdqWY4qjOY3sJNJtsUatsY3MOFvwipA6pZoHrdR6Q1XA/fQWM+Lv2SC1sLZQp
rfhWVBPgsraKohp8k8R2jl9VebxkNgY4Epi+JoDlWP0c6KIdbk7ZV1W9aJGyZ4jJdXx1g2OYT/hz
MlhWtD1s8H9DxLGeoPAcBsr68OPmMJYMA3Z2iUGE+4sFCGVpa+XiADYfMKZjdBwUL9YMDYTLXqPg
+J/7ImIZRdpTq17VaG/0l+1l0TlRL/hitivR0CCauZplZzhuRtj6fkx2UD/PxreyXz2O6f4uupt5
uF5kMfJFJbWxUlu8H1ciqycvx4O4cOxkxg8FzSdAxQonFNomlgwDHcN7d7pgvZ4pss+YRiEXP1Ao
jIYrCjYkKMbdA3o4JuvRLkmuxfkp9+L5+Yz/B9/EZW5y7BQszkXLqeltQgPEB4zL13lFHH6rQ6bJ
DBMx3Faf9Q8opwKYKLQzZMsEwb5L95MZj0eSONFzK0U3rPlmtHDL9alocannHVwA1oV1k7QqXxpD
70BTu/nvpK0IvH9lBPeWeYL4FIlYgXa89og0wfFA/yRkx0UeXi8rkcj3yzMFGprQ+XeVA8y2/ZVt
BYC2c7URMBEgKGZjUl4HhHz4X7J6WL+5R/L85a/BmosbpqS87CE2uS9faw4fS1VCnSY7SrlzkpVS
qpBcuwrNvLwVcJod4d3xm1jOUnLvNA7aFpO/qCfc8UDLVDNMjXoHw9+ZikgFlRJAr7XW9TiPHcNt
nhCHS6fxRj7mRc/Y0mGap8OL+3d1oQhDxjs9HbuA+ZdEGUxoNlpvBbtzpn1W39uvQqW7f/oVIuOr
TYJnGWJLLjT2GrJH1ZG/8q3Plv90oR7XQTE0syjFldoKmWCn5KFj0O9VUnCSs9ey2JtY7XTOFAPQ
hsmEHZwZUUYeHOXTLr1HGg8H7T2gNVyY509UWa85Rlejq1LGYkfEyuEYGtZgswKDMXGVJGUuSSgP
HcpvRwylG3kyCVVYMe4QLiQyHiCaAIA5OiqKlLW9jwpf8xJOqRvBrgnmmimnyIe6u9ciSidzy+T0
iMpp5UnweY0x8YUemj5X0ay+WvYXrVLpwnwEc51w1zDc8hJq4nbZqC/fe2V/Ge88Al5PdB9jdykM
2jKbx8gnDBlz4cVkdO1zTjRw9PM/Q27wtul1EQEaDc2NtNh1DgdRQfxmgnZLtdCj7Vsy98wdQgjy
a/pschgsyz18lqvady8xr1jcMn/LGpAlo50jaIuD7kD/33B8pgD2yHg1JXF2c/252Zzs5z+Uvz3Y
aP2tGLVEF8Ptxhk6Oe6Xznc9tFINxRdkbiBj6IT1U5h3LKvq7MDg+GmHwncEudnIGSgQGPu0eumk
V4mIUpwYVszt958s3R1wSCwE5MWLeJGuyVSqnx9sGUZmewl55BkMLGBcyP2fngzEcwabPAmCcKez
pdC/I/T8Q4FbikVZvj4ly2Qg8mFXOzxAcmHq6A/YCO7jHOopQ31uUL2W6LEzLHX6wU37QAhyh7aj
8kw8Kv2Gk/LrCV8/145QpCuBER2/dM7WVHnsi2WUkAFxVOa7hf/xnotkYGQgHYTOR7UciULcn5K+
oloRuKrfDhI7Pm5OfZl63+N29KbjPMLN4e0r8/ktChLWzZ65GrewDTJBW33LnnoNk+Ei7gBVdPDP
e5MdnhVqZmFZQKa6tV8eHBXqsglB81qnJ67Xg6Vn1qRoQYeGLlJaV9GPMN0HbzJXkxJcrvhXzxdw
f2WEASuZMBQVAkenPCnj1RHXVORg8QI3FBab1+EWL80SwXuPLkRi5TH5foXADUlpDKfeVU2r7Xch
ndmxdJKt68oaTe98vBH6pSorqk2Sg69BqD0oJreNm7cp4Zy+NwdzYJbTpJIf6VUnNMNxO1aWA5PQ
9xGZvGYc5YgnrY6ZtbTELC0bNGCqEX4Z5hfBWV5+R0d6EuAz8bFsx7Wk7XndwpbCJm8Wf3VW92bM
H5DuqGtRx+cU/RCciS5njmqvjH72f4BDzg8KeRYPQHkC7N058Y9yi/McurE+iCXxqe8ZrkypvRCI
8K4wx0hibnC0evb2NBrovDEHweYgO5PZ/UDiL/D6zjuTn1KjJeb9VBBr44H4/Vi2mI+qLwHltmdm
foH+oluwK42sxMw5wkN9CnV/cBoD0zvlWPsaY9ou++mOcqGSRqDTJd6WJWxDPQm2arGANMMnl5FM
7b0+biMawE2PSrXX3noYbo0S0mjL3XZCzOS81rkFZBZXXOVqk9Ao9/lPQVs59Pww1Lc8+Ux7wC91
RtR7ozoZOtQsb2/muA9IPzjCK88aBZmvYGf1PyBv7ScsmdMuqeZOzmWg3HwSY91XYulb9LWSN61n
vA0isWnkPN7OsazdjiFQLZVeCs8uMtscpiVDe0p+mJWLgMK2DuJkXWFpIjWITlULC6w9GYlwFQKn
KjJU7Irg19mcR5MGRrp53vFXhvjVjEM7vbHkeQJcgFJHEP1jtCLPoxLRV1Xgvvth373PmzQMmkmp
PKlOkodZPQbUedh2WN40QctOFkrbD3IMKjp0SZc3h2nOWpUlgptX96/T7sKvkAuvsCQqzq8lqE25
KqpM5hatg3cpuu/rrqL9QEd8CuITFg4iNHR2gGIoCjXwQLus+xBjAixTNWVFzQUcNny9+sgI+hJ9
fvFE8ciwxU8tRUZqtP36X0cxe9EQM5ovFvL+gAbJxrNMghKZVNGmph9MHHMRCUuAnKHvPGutMxsd
dEYoLpKC+NacJFyrhZKAaJYjgIZuSKSu2Nq5XF/V0aHaTDVKw6yHBxuIUvfnxvVsH+l4RuHIn5L9
0CRtZatp2crPMjLkJsOW5Sli9JoH7dboupZIJZkOD1rfPw2XD3JNfKHujCh1zuDYlFkB8SrYfPKF
jn7IhdzCPXR5Y6+pDoAEq3u+t4PwJLGLXlSl+qZJ86Ha81jMRPZn7s+dYsyOy2OR564mnkVlvQWi
933I13UXh0EDssyrbobpi5JWIpGF2D+D0/yyZ/NVwcsTkgBk5Zjo6vyIB4P8fXESB/SlDyOJ6RYf
SvBm72HCNOpv1RH+ZKStKZ5ebnoqkkWRWCdp1BxbwaQIKDG3SoFch628QM+wiwCvatWbw3bhVJLZ
QKeXSBvhCydCP8VrtElA7vZEYHnXWElknoROjTfyaGQieIiWI8Qehg83yWkswZ3o6I3dE4XWkhBB
OQrPnjFZwgAIhTQrhTnD6dg1uNSMUqgdwrbJK5CXD7PNxeXU/JY+yvJJHsBvgmnrqBlpebpiZeRc
cish9bXGsO2kGyTkrGjWgEeLKq9MY7gKVIxAbc50w0V/zBs62TLG445+EsnTT1gwnCWPEfFn2nkG
RRonQQWqfejpHNRLdTaBaeE+/RgTe37b6ozI872fq8zJ3Kkblmgo5saOoinA+I9XyxVKTMVSVRoI
yL22BT6c9k5H6258AHyX4vTzF7dMs7nOcDYaEEowkLLkkwKjrEIv0lxvvRFHIyyAagjW5zVmMby8
YwDqj4q/btESjJy02NSq1TElDoU5iXfYU2ryhGB6qRhxADaEtpVzsEEGPPPPdqD5r5t6WSPMN/EP
j/vCQwydinf8MfJX7ArsMy0sz/rXcKIfbd4UkCf0UoiAqH4oM8vFrEQplc9MicTMMlG1lS1v0MZr
lMs70HN4C8zVZnkRLoc0IhAxcZrgieoVZJBsGbCXyjZfTG4Xr6/9LMw0k8XYbOyxC7pb0orqoH/t
QmL9814jtd0BjUq3mUvyjsUQkBfntmnkdQ0IRjIRoa1ZkgE8PEyPYIcWp/hNLE1hOPMzi7jPpKaH
RtNbBTNhA8OOsImWxjfDSJpJ8URYUmZNfLFna/U3gTmU+EN2HDOZHvWFuTX14e0PT15/AVlBMmnn
yt7L2BDnejJcEDBhC5hNG24mdxQ7VRjbPx885BQ3lZAJGVJ4jRR9YzCV9kzeeKN6WnUkVlOAubXn
3jUTtgdLhhejAjXq5IstJDAaBYDvm3VhsPnpjHDEl/9DJ+tY5S0ngomoWrpiKdEMW4/t1Uay/q0O
741J39Cl6DMz7fqarJ/AZr6mTMO7knCwGx+XYiJnHZyGkoXIhgY9q9kfloQ/R2CCgm0l/woyIWUH
XcbmWDrmOyCl5Xznjr+wIYvKL7rI0n0loyfUZtEL9v+c9QymR1Je+PnrMXe1Q8ejOWUh2MjldC/a
ppOlCIEKMyxDIz9WBRVORUEqBnD8Vo9kJ4tNsEAxX8KZZ1Um4G4XTaS2OAVmvwAEVDddPtNsnl1s
jfkxNEBwxpxlbkqIhmOMTvwxk3wxDFMWgFN9S7XUTFFGh/RAjbqsXRaQMhmGnKMAmLCGR8LfcWcj
OeRJ220AzfGOQHdvywXEhp8iYX3S66jSycvaUFzDWdLNNdbxsa8mbDcd4INkoCbTwLof+K4GAlwi
EshLp41IYyDvfPPj68I9kSaOd9FUybntFTgXB6L4sKkRHGVWMP6ZYpN8MAsc1emwFPovvKmql21i
46e/t89ZBX88IDd0SeufVSqAJHh0gXGO1hRZV5UDBLq87z1+ukKojD9un4wJbhVq2xQRQ/sLk5t3
HTqh+HM+J9rR3qjsgbn1zO3t44I+f+YdSefVRO2/+J6wtDq/PIabYqHr/olzAxhv1suo6nvWct8Q
n+aRAl0+bI9bznx2T+Gf/3txPuD2o2IuRSLtAIme3o4wPMqDUQJ76E6y5GuCYiVmouzyvYi4CMeo
KjT+ogzwGmytj76uCzDrWMdbx2ddoG+8u6w6aa+aDIufPrXfPC+FF8EWhtSfKUI620kmkL+yWoCt
9rPOMNfz4GIg9NAbcXMrISTBAUaNyjK7UmlOihSYezFgWMJjFoMDd4VkDUwsjOmJ+jfEezpGqz24
Ixsu2X2QeF9NGWq6CvfNlbSngycnbAKzVkTAmAn6QugNaB6jU52f6vWnd40+XYkeoqaTEuH7SBWa
Fb3wYla8oDX5cK7LkdMROg2+28EHdABPVsaoytEIG67px7AHwIrO/exOExKGpJJ9+bl0d23ay5Y9
HWac9+gymweIC69OQp0jk6sEXmOSHz6YcoFfObP05hxKEkbMKMFXy55aeqsArZNwGssCwzvP2DDG
yG7K8Gy1T5e/yS2fn+TYUTycbvQJuerAe2nvnIe0GfaWwxMC55yFlGkGOWZaY2fiON8vbSrfRHQV
1BC2rriR6wM1+uYnxgRqqGI7QKDVNWWt/25m81msiQ9Qx5pugkZy6e4q9HyhpBySMZ2ju08xxX6s
YB0nE8BbFcIQzUNyOKl676jdZEWB6wnv5O6To5D3SY900bIPM2hhicRMBtb1fEObOgtiCi9ii7/I
J+/J6gq6tlS24LbNxHPwVn2rurhfSdqgkPn9FUlaXpcU8gxTTH3n+9PFFvnEBaRrhRhJ7JpoiYmB
ozeenyu9wMJtivZ2zL1u+3d/JjAifIWB4fnISxNEqLmRfIZqX9zT1zxxito9+A7LRdXBmCji9r16
4uAU9+mbX//1Nx5LrSMfYWiCeBLU/gK9yIrbQtGVF4YtbMlKTwfjDdCjB7cZKOlIzdobvzkl4fcB
bHa+DyRThomOhTbuHwLcAHTv6O1zA/cmMIFy016EfieDoGPtoNykZcAA/dqkxnkbtKqf6hFLVpHe
h3FozKlkbqU5aNh79GY7DAG2L5GEIJXwtNDlOtFAAhKzk2diGYbx8Y1zsJeM+X5eZhASN0eA9rvK
EkB9ohtT+f6/6nEhpnLHGaAaVAyxJSa1kl7AvCBEh1PwkEBXlKMg9sPUKhwnCABvDx60SxdNUPTg
DflRsLQ8kZiq/3oQUNIyZS/ZOoIuFbow+G4JlxOFQT9etK2KT9nZqbATgROrQlAQzOD5XmULRq/H
8xGdBHNudoR9cpVRSnVXi0bI3ZlTO1oQQwoDuDB9ZpdRvIlIyChmCntezUr4AlzcPAndKZrauTRT
HuSDTseZi93RrX+n53rZ8BXz4uBWVLBbdc+HClrHLtTjagcKVsdxIIXIYZ7OkeB/FAUNOKOQWkYe
nywhss7Q+JPoidcsBcagiJVAFeda4+TLRBUoKmj/pffbrDLDMogxPcOUfwFjLaBW0T/7ORBRgvFU
4JtO3goTkUUrfbrUXw0yTyfKige1WFqZPah9/HMQ0NwcMgwxfX57bgEGWpowgKNntFrlxIvUFFMC
/B/MzcIOHgutmSQlYMvEcLYYPOj7y+zTtImC9uwprLBDUxsaPWPjSzejXcUsabMjqoS5eQ30CY2E
vGZ2beEZwsuhyB6YHIBzlnPuFJesDS1AK916yQpQhfHaaRe5H1rqzCBC+YDBepwtrGawLLCYCfcR
I5XprkgM21Tk20BSUSoq9GOtfvla0SlDZsdhuN9BP/7+wxeUYe3STugqZeQbfyiD1Jv/ggjbywTg
pMxWes6bggzXYCt6ytHVulzsqh9/u4qWBiD74xXF+eZBre3s2BWjhSKLYzIwaWwd353/wksbGROu
tpU0KYWFe9foPmsiYnXL7zWwIEhJCGeeKVtLMgK9fUomrC+0j7YkPtYjLrZ/oHvsdB9SmcYtAsgx
k7aE4+Y466U0TynDrperYUB21K8SQJLKwsBJl+HLdNLKl7Y4cWYDyp166aqsM4paAf0ZE8GqSaT4
+ko0iFb40GrQw1M5oJfFoiFHpRYsAWIwCIJogX59P3VEl253tNkKbxxYnVnAwvBDIkZBFBbwFkNr
C3/clwVrrawm9A6jrXgusjfgV7JAf3mMvAR8vMZxRZbZEi/gD4L2fOUgKSDIcorv5tNUBYCeDkib
oG5uXobcykL7zIjlAcUCkerFBASL/za0qmonARnf1swuXuUdMMq8pDkGKWQiv0X4ba5Qye1btYZa
e8xu+B/4ZPorpATUh2XTuZeWX+2wwTk0PceZ7ev1mTwRX2txAhBAPpXlPYAV91KokO+ebMR4I6Wl
9TLiNiH3qKfxUJRbAk5/GF1hjVBg7r6GgjqKJ2Guhm1VxYjf9imfJY8kEwuo6CUHcqXrRP/ym1lf
c7ZnnZbws83+SrNm8L5N/pPTW8jofLtMCqrIH/mp9KIuE4aQN3NBseb+O3eqCcTxeOQCjrvQ+j4i
WJ4/E1xTP0G+E1REtaZhuIFAUXAYd2VD/KMe2eJzto1f2ta6u00MKUbBeF85B5RSOcpMLEnxYs2a
/fAuPcgUDyNSXhCPhNc0io6yCPpcgOCF8HcPh+iz4eIFRSr3QVKdbxOXWDQwWxS5h5xygBTaGiXy
dzQCJSgvhL/Mfa4k6CwWoYafBIXXXA8Ku8EEtxivBujZYKbxHMOL0qfnwZ8sxgwJFESrQEzULCMj
d0h8XgNo9jD1VZSmgPWg12y8eHQ9RqOdajxO2vDr1oQZEginWCNH+urjJM5le2nPq5VJSgsWbbvv
vPDZwNRTOaG5ISWXx2dy5CevaBUtbU0J8kOFYz0n5x2jhM1ZhZIxMZkKeA/ps/lyvnI6dmHmww7L
rfV23PpoxC8dBe+gTU8H2mVKnA5zTi1Sll8mauvN5Bwo7JbHDUVsUh1yqmP6t1JeK56zsFgaRGN2
wqAI73G+YWggt942RdRPSL89Z2w61TDA0l0jmhz49u9hoH0JkSpG/2saOLgAreSzqs5+/ZkSEIZ1
SnIpMqqCkrlgGUI8c8MV4GUfhM1uvMaKKaujCHi9vpdot7llzpSpK+HV9t1/zRuz1jezhz2UVPLQ
pOpKqnnfhkFOUqCnlwJIJbJQl2Y/bjAwv7VEQEo/46I8SK7dMjr0iXXRADMSVLp83FhAILmrsBEz
k89N7IAdbREbpqQ25OnYrdevCqHIWm8hN/AaxlYvL9RugDUk3HqZ2XgrjAKtwAihyIOdan3KyBmH
8R2JbLHTSKxF79/uv7bJW07wqNUVnIrq7NAlWZaM50gX9jF/jXHT/Xc1gi2QrOv1EBlzQ4iHgOvs
688l/4EuPUlJG1lGFefE4FZq0zf/2vTLxFpoVRZtjL6R4I/xcg4exOkOGtuvYr+aYLzWsiymlJoG
7noWkjtPu1NcWfxSoEMRasGSOYXAnUlWJeKUJpof83E0Unpk4CNuU/Yawuu11w43QkkhbD2ej57J
I6HN6PVBqrPKfm31pe1KYGBDUAFKZTrvqlgv1qq2KGON+TIfub9HqGqtykECIM6yQmljoxrKtyqY
f5XauPFsZDFm+hxDJkvxD0jBYnyZ+pGS3dUPcBFqXl2kxNPp9ycfb5WtsEVK5GSi0Dn8Ro8bVuDM
yNCu/Lnhz+Mro8XMqGt6dKm49jdZ6ld21jtY/zOa6JG9T5cehQeZK4yw6fpIf9WGyXSO8H3WpY+V
TA+Lc1cMvxfQ8qnJc+fm1W66okyuYem8x74k3gx9289KUxl1QGBei5X2ivGL9umPFdV7Ikyh9oOr
TOxZ/wpw1jRGmVIZFOzkKDViVVkx3UAXXxR2FKdgN+PvvkOve9P3PxXKJcU5cmZxkiselG02EU1x
pYAkU1atI6ZjmtVEKlFemfA56X/frWhHTUwYnDvabxHIRJGKP7oDWU3xZK81+DwtLRicsL8AVgfu
nSJJpDepC8DTJvICjjfAXAUcjXi/q5bGU0hblMITb074fj7cNl9QOREQvj+vti2WCDrDHhXoZbOV
vYjv5I+Z3dryprYFUBShcH7YIYBq/AXe/VTPduY/hFturSxmuksUPBX23pLw3ph7Qlf2ws4d6oWS
Gj3I23rnCp3lajTWpEzbnzqUW99w2Wkum9LCHcCf9wRKercm6dLr5N9b3otbml7vG8s1Brv8dn9y
UBXMrrLjD/yinZKJ4qF7vbh58w8SDLiTSznwFRBg/VV11V2udJrx0Uxnoa/2GLZALTe5eSeAqrr4
Hm6uHb+SF+m3XDMGW9HDBeYBTGb3g6yEF2a2Huhqt7rn637SDQ4rGtu+X4Oqz5duacdB1q/bxrV9
2bRUMMfrJc6lfNuOxMjH/U/3RNARsMds56FFM/LWkJOJ6NoaFcLh2FxrqYAt2cRhf78HXjmPhvi2
+Ew4tEfhSq3qzHd1aJAOpXlkOUaE2lGHmaSkulRmWKG+kpGli5UjRvjU3bfskiV0myR7W07ygJqp
pdHVqf4mYY2bHMKpUFYIobYc1/o7wJtRrdO2yjApGrZFW+WslJhXeZkfY0jptMh14AAQM4fviZtp
UaUTWpkeXNubjDhG7wLIBmVSgoYAVr3VXqnQgFS79By54gB84reQZISqb+3XLgVwWQdSm5wOwlXS
u7noY7PT05kISccy5eFO+7x4KBwhKiakDqnm7NshpKtgi3Nh128cpw43bKNK36EfLJHEvGQoaqF9
6GQnQQ4BfqG6QU4pP2zn69dRnGxknjCAW4EIxMr7zOZmlpYC9TRDmXJfXfuFatrqJXdQtfDgoYqA
2h5bzx2AlKHWMWlt9bRwRnIJgG7ZJMVNPt1Jradj8k3y8lNVC6xQ0jzNKIzJ5nt6U/jXrmccN/7k
XHiPhCMS5rn3WR2FzdZG9FgYyVK2vcNECNEtwAxxRZIlUoVBYti3PF1yAgunIj7nhb7uFOy/QsLI
tdC1hLkab1UgZXx1AoN2Ewi0MYGrIFSy4xY05VoISYNl0pnkC98ymUHm5sExg0C5VkQT3ktUccz0
C9bGfP0l21qu5WeOfHTn73gZWfjt71STNBDBrcemycbXz7i85LETbznuAyMibKnKykbfLJG3JF47
WThfEK/gy90N7MnNa8uwy0MbAss9b8gLGYvzFV0MUezJXEA20tGayF7RmUKKrG42Xk8zfIu6vYRe
U7papsRuZznUwwsc1XlFpdLnJ5MiSKhq2/a57MRRx8z2pCIJOmApYmyX58DmL4ex2KRPGNDWUmd2
zlHpFJ21PQe8EsFx6495SGv54RuoWfhB39ePCzK3mlbd8xWyIM8cNyisrASp6imx4WqmFUkzvrO2
cBRW2/CyTX9watcwLXZZ0BF2JcECOnFy+/1VL3TqvqZ9rNpl4qt/urpkeQG1ZOFFASGiKh+01mVG
HvJapGcGujb/sd999kokcpsYwfl+dm+FqZZqzO+BEgDXrFd5VUAhW6df3YMisKfuscrYCPDqAXgZ
SQ4tcZlL2rYri3BJt7gKmeKN6Pb7eKJb7wnvJA5Pb0VA/Hyet6dHAlMvu1A/p2CWmBsyK0BlMw0c
8lmy32VHBwRAThUInbSHp3HFcAyVVOopF7Ucp8a2LFOP2VADtNAx70lylvdRdadDAJN7gd1/+ZJA
kfu+eYh0szsTUUzlBL8Gh+KEMXPL5Ac4U6YH6VNycx/Na7iO8KEuZO933rE9Z6Pcm1+0dnsoByG8
e3odME8QHQ2R2JPpC7aqptR7jYWdTQDRX649Loz+FUqlb154jLYM43golFSwqAWbw0POf9AxRbvp
AXfU6CrY/aFAdDt9kBTmsieBNhYar6CMSmWbP0zByDCqIDM0u8/O8XgPPxC2cTT9xsfCTfWkZyLj
aHlqxpKJ1D8ekUxh0vGDU0mf2fhGo813H7yBALKGP1FEOql12PbEqXYp/hYfrBqYl4rMMInSiQYI
Zpd70BbAuXqufPUvpSWoA/cc1YWuKwz1Wy6dOBamahZXv3jgiu74ngD0x4BKtFtSHu4zPi4qmKPz
Ip85+M6+4E7KEYePdOnYAZbIu6w0VZt3QAj6sYm9QOcgr47kEqUswfcuza8GPY11Jzo0LCSRyWCS
Znwau5l9LAB17otc1CkzBqVvdPd/4TSgMhIBLry4tu0KhZzBQc4mt0D5Tit7IQ8RCl3V+C2WJg8b
IGlS/ngWfa+5TTUDEGPNEmh7OLk7NBR1f8aciL47d4YJKmhsHDsmfRYMGqe/GsdO7TS6vpZgi5SW
zmBEQ4nRbTJwvK0RfbmeWx1tB66JXVqxwHj3JkvzRV0JdS3dcf8G+tCrPAHqJu6gw5+ApFqxMdhX
Us4DCfUHUGxNkbI7T6ye2BNs8JfPnDAwQcZDe27FtRjX95Z0YIQcWCdjKg6BNp75dR4nFMWxPOQ/
z3DyCkgxOMRuNzQ4leVQjow8xAuBX2NuDaKioiq0fXI2u0z2E+nFLgEOZiFwBLMouiXGd3WmeqwW
KYLjtS69qAN8ap9xsK0faBgaJ3N/VcV0ilohSyjEF8rnjtdH2p36asGDrVD0xAHcEfESbKe27sUl
0IoVkhHFIJFDPgaK3Y+sWo5DDiRbhn7Aw1hvQFIaKbeoGWsGkPeEY9q/8Ars4bSl2Ed6JChfzf9o
seid93XHWOihRaeyZFnzIpyWjxBjAaTz9cvE6F9+dauSfFtBxz9eelT9Su2G/TnXKS7T2BpOwT93
eU8HjoxEFD66YMEMzdPHLEOiRtRwUNFaH74xHVOzSeAXdriJJD44dDQB4xbOhODYgM5SWI9DbIvo
J2Mqg6N+igZxvbTL2dvQ0bybuaruQGOSgqheJhjB6gftIsa9R6xeCtN8GEbZ9ZYgoeyANbetCk+f
f5ty5CpzCKKSdO+mAt+yp3UoujBPS8NmBtCWNCBBMTLvQXpLQbiBMKe2D9ly+aglpyLRRxaRDNOm
XnleGl+UHQIxUZHIivYCJsddJK8kac059aJnsuqk7JHNTYCDQOHOob+1EYKp7WPLz2Bk25qggYIR
VF83N11Lex+0TRQIGWrfqBH95IaXiWPmIZJglAE0HmMzmUXzwl4XLNkJB3HBVXCU1nX/9Kn3udNH
441+ut8gTOh1lLaykdnK2UDyzMHZL2Fa3ac7X/JZgyUna3DSeKMIDetTWNDaVqbwLdxNuH5opXhW
JzZM+2xp2O6vjePlU1bW3GtQesLJi9pHf5fzUDC82VLJCWZSW+gCjzOnwIIgN++TxJk9FwucbBM0
SClAoIg3EVOlF14JYaElBOMUo2AKtWOIj9RdlGUTygEKqLa9QCYXfi3j6PmtOs9Q9vJ74087d/Rc
/YF6ilh8yq2YLe6mAV9xUD69E0dbtkpOadMOYVSCS0gU4EwGUPDBQn4wG9HR9ob5zXJztPB6zYUB
yoN24SjxTs0BkevZZeZhfXSz+OcwS1HJYwNWCuiPsLfCJlaL1NVKNMEpGqHdk8vLc7NfLa0gBiBp
HubdEGmGwVrOFG+y112ZpG6POUQik43RYKc8VdPQvv1od+n7jkmcqQqMX2AYx2pz8g7tmQ0bAtG8
a2qVzRQzEeVwDa7hJfybgEHh3hElvJys9HO6pnczDpz7tPWXK7hiVQ9Zky5bJ4RCpHxS8PHFX0A1
DK9yupvvPCpGFEKQXlbTwbC8xfLezOfXTift1FnsK0ibDUqHS7cPVt/G/7/fzIAcbKtDgp4OAYjg
PWGOpQpW5cwUudVCLKNMaf2IEiQBTSosV1INbQdokzVIya8yP7A/fZFSv2EdwYzUhPskhLoCeTIq
a4P9NC63TXp03ltZKGv2WVnOX561ITgcN08vE/OZ82gSXBdwbAYo8PxfIRFxksFZVCNHjDjcKIl4
ZaKPxArK/aRbBrGamWemByH4Y9gzX9jMZib1WD23qFhD5hlVXpl69OkxiVaCf1MNbtcjJIIGr2LZ
14imVYAqLf7fzHoxe61NEz2+GKr1c/yFzAT3XJhU4WWfsHTbJhrRAj23LjvCZhEHxL1iP4igi99V
GDnka+13Q1+WOrKzdP6641yGBORkjqHnPa2RVcHYbOySf6UVLldurIaesM1+vTThYQcBw/G8jaOX
GnLGkF+/rAOkQMA8R50L4w8ce00PexbZsUko13C7GxUxGFQFrDULZ8SG88CEsu002Dg2j7c943uX
TY3cdjVJGL0msTUkFQiABvqJJGI5r8ZLYMNppODXLbStb0Rug9/3Q0V1TDQuwXwfRZzdInHfir8h
lay6vybWa0qxR66kB5yYRNnRwGJ7s0DdbCTosb3LtOn8N4zoB1PEdftsHiK9rm1nq+ksWiWHpKra
R8XoRq7xgDTd+HjMkDZ+GsWI5j5cbGMWEIspV24/JTclWTAHMG8fwelUUB2YNdpypjLDPbe0yKyR
XCsLabIS+MhpKLwlzPnuJI6M67qJwpxeWpzDIPMZvl2UMtNZivW66cBRokHoM7jWpFQ3ZXyQtf3d
+MOARLCqJ0Ya2/LDjIx4fz6X0Fl4QjkdEcc79OpP4/ay8cy/UAcquizb0uLSVHD9grdeXzdxz1pF
3x4p9iFAhx3UoW+QQ1HE2fG/jgvW6v1JpabuYmWqpznL7aQj8qt0WFJZ0abVjvctkigJ4K/5Oy1q
RWB2xmv9E/iUAQv7EsbZmJ/HY8K0e1nNrqJ8t107nX+TLQJzwkP5TEGPG/S4EZjPaNaE3jbqTsha
J2QJcYhv+KVINy4OBK7RUJEwt1kGjHgqXT4xsD0eCC7p8V90eROOMEFxIx0bE+LF1TmjhwrJ8Hlh
0xJgi3f5TQOmEP2dbAq/Dj+n1Jq+nRhLk1KxvmYKZ1OLKVEm+9LwDMR0msROo8PFYQrUAnNITQxF
kLI//CIt7xcwj4OafrrpF6PWSZVKym0fBT8c24aq1F6JqGvtxy8J6DDF/hSU4t2IE/PAT5J+IzYG
Zv1Ir/cozpr8xbVaOoy4l5n21GC0MzJjjsksW7nsHzFjg6a2admiQMmGRuuc48VxDeCD1L0l/wES
V+ZsEB2fXDbXxwhH7ol19F5FfK9IM/mwTVV3w8FG+6A461vDqAlbXIBc5381Pg0lVV3orrn8EiUq
XA/1l58FsyMhFwz7yb+uCYGpJA0WwNuacgdHVV3TBlwPejIRguLXHUhoNVk6Jk4SZjHsLRwKtBVx
WowaWHxcqO5RI5DQdWwEoSYytqvZGHait47Y1v2hxoIYYCEwgEfadDQYJiCFtbsJ4qgDpun/h1le
cX9pFbmtRPuyDtkec8iv18P7xDaGJFHOxqd2s7jolowcnuA4ounCEtvTrJ/YckLQeQYh2tHo6yvg
9hqTVFazWbdsCLhOtx8bkC3k81aHe/rUlkvcHw6lJRk36+o/BQXd2s0KRVt4Nq7Zamhig8Wj+fRr
z7Z5p8ZokX22iEb6ckK6eyGvsSef1TqGCQI+5PQFgGfFK7cIn+0ugp5u+fMpE+sdjein+w60uxa9
7oPUDXQ9RwGkmcXDwMIIeBBIvRrwNWMAB3KsrXHuvI0cx2I5J6OlRGRWrPNmw/8mbURJlnhxMB/L
aNhNzOyTs9NCq5s5pkhmK/OJauNGDRoZBG0UOzXeqkHBUjb/JVZX5BbYHcFsUrjmDxag0diy9LF0
PQi2vVGpkJI7QMBW/dJBMzDXnRC4xRfj2QKaNc99owh4F0TKeEKScZdUyhyTS/SS47zxzFhjQDAN
9LfZQ5qHkyh59qNn6GUjAolez2ZS1oc1fXNU8SNgiUUQfkoQNa32umpRj2G5yFZ6tt81fx8dYkAI
WkhRR3RLDWcnS6rOd9nGmitEeQ3r+xQKa07KZ6GZ1UlZOvqmnTr2Q/w+A36jtAXIcyyRYv8bmpu9
/I72q+f4wqBUC2ryRe3yzBR7ojzrASYffsJtwxbsGmO4T8h8+NyH+RU7d51uzAaY7Tij8OSzIugC
RHuylPZmgPBTGAc2SXaYG6Lgpva293oppqPTKt9AJzdmVZMSu3PIBvlRXwjDJoCqwjuBbNRU1LHM
em4BwYIX8WSJyoeGcFO1n22t9R+Lt1La3uWvIHTB+5r1qjWExI1KrLxvl+N/T3FvnWeD3fLN38w0
6N/d0EoP0bJnlVJwPSRkfhAzp9h8zonqx+7vbkYtgAUn4N5YeurEIrFlA6vrb99wTk11YiHsnHsG
iwUO+xKJO6cYkud0DP5W7oA38rbZidcFeF1nQwIRgAUxuIckBwSY9hYVY7dvjklwWqzEUziBTbZq
uW2bW7/GIYKATyyVEDr0cE7H5ppeXpX8+SgGmqcEWp1jtLTBPnmB6l1xfrWT2VcSrT4UeJnvSfJs
69hD10VQgkRj54fo8WkSZKH45ukyl0YktIAUE+uiPGPtZVgQ70YF8meqrIt8oyZuzOgRtD83phUO
rWNlVVMU6ddvRx0nsyxXuK/fC64IyoSIGrPOURJarHOkQtcwmaHcMFLo9P0aWmRSdoolui5awmNF
6+n3zr7EPjPGTDPY/x+i3eQd/pXMBzG9hOCwNLHiduqyntuwhHSU03F8EFCint85ky8IRrx1cSYU
C1OMuJqFp0Mnmf6FxdWIEA1BUrVgr8WaIgWkY9R7h/v+4zIlZ6uuMPOle5GpZh/mca6fRjDmnC8h
4RsgJT/C8SJCql7i0IFnBu6Gs5X9oeL2GK8c0ZchSRkP6WcWXQR31YORdEsRp5+5T32xYGxsRlIO
cvzF5zjky4ZcKo+IPoCyKnyks8R8tX16Q3R5z7Skr5fiCEGT2LZPXDQCrIBHoSFAVIfl5nN5EXZE
3dMQTcYBKJc7Jd3K0SZylXA3GMQUWo52pOsYtT5FhKe+HD1JC0e6cQOBgzp3RRTkA6fzGZtxpGvY
LppLgv1DQXfIi0dJUIsmEpXUyfLmuOMPWBXQot3VU3AnQrbi/xmzUwT5gHkn9dAWRuzRye+A6SFJ
rgSovhWgWiCGv6Z52/nKDN+iNIcTVcC6q337YHvRvFyPXI5oLf0hvYTmVktzpsvyMQz5cUMmOJjs
dGSz6wnqMZZ7wyTWc85eTuOzpxYASnGdiQDSHnKsDotCyKEUY1K1cjE18U5T8ukLQZA4rKoc8wnE
LWNe5Z1Nb1WoNAlKfLLzFqfhEAaxv7yFGpU66FrMBtNNzGs/ums+mXxDxGVwal9jEPuD0zFp2uCG
oelrQZthKqieCYZS1lFwYo5h3+Xg0rW2M+jGHzUbPtRvYxixHdPDCv3CHFQ3qh7YdDC8MiHWouiV
WPv+wZcUlHrvlxCzY+YMNK6N/RQ4NsYZGY38VQLaSa7hhF8Y2/V66pZC+Q2c+AOS1dq9yhtpaaAI
dWvceJdHmmJQWK5DilNykjD/xU1tn4oa6n78rNtN5hLCWps+ZiCSpybRb3j5/bobGOb+6hzCsrY6
SYJJT2HRSuxjp2IDI29RQ2wp/6s0mk36YTDmHpfajIdUBlJFNDSAVLmrs8t2o3pEJcytJ+lcGkpd
HlifLPJtME5MfNZkXNQOsn5jMwhwJECLmomsYJ8pm6NTL5H+QlREj/EWPkUUGyLqeqazKUH7HqyY
YE+0zdZ7HZugb9YtLPP7wnHsOmudB3e9miTyL5FHw0KsL6DTawuoS7IbQ39ig33QVUPk8Cu5Wqmu
aTlLAFfafC0Frh95AnCdDShag9Co0YBqtq8RbO8E38SexJATGiTOHMuJCzaFnlXU8PBv2yqfQ4r6
MRZ/K7qyw1MAV/IP8cJKE16yfydRRQmao7Ebmxx+IuZ21B/oyHrjfrZPPgC8IIBXXi0cPXxC0QR5
4kKHgTZosIHEzylTuNNxOup3LgeQ4oinGS+gIUNcsdrlmCYGZ/wQ8HdthDjwxAI1tE0PlxTdGQKV
81t/apUwKlWT6V8NtM0VFPDoRZlvlYM6S/ZXSjQNYmWJ5SJUAFGWsuk+Zn1+uP8RiR54ajMjmdmm
qqWDBbu1qOg/OK39m8dQwlf6WO5da231or3wWscu4vSdMcwhQWWQxB9CScC3mrkOdprvXXiSBY0O
bMj2mQbRrCJdntIcsJJ9C1CsGr/Q1XbP1a4LwoCGXu1zyV34UK46UJuDKC11RQN69kRyrJTl/ROl
XcdYefCk8v+g0WCsCuGwtpwsXzK1JMwMQr9rYwYptTkNe2GZrXBx1Anq7YSnlzkOYgnZVWeDW9kX
x6v2R+bSCxmUuZWPTwTjYlk+Vb3sKqDXzmtLHGD9pKp7aMT3hsVXaQMZSu1CphYiKDVOgFvttg2T
XPs+RWjx4zeKVGJbVIb88MOyYoWeNbugaX+oQC20+EP2JzY5+E76zpnaP+zGZrHr6BXCHRohjmZt
iC/3B0HS3GjiG+yfeHfd51ZebP5UjOwFBridPipLUoLH5j9dIW4bjX06Jhjti8hkhMa/Ddf+IHFp
6s9KJ4jk0RhknwLJxrte+V0U2pLW+zJ5tsPTAxIG1uPtva7G5IGAflKqsmodL+psJ01HromJLRvK
OPA5hfomwCktcCWvN+AjMkBKj6XLduBTMFB7qRRcnmfnPlEAMmN4VbM/xMoiaZEUDgPQxcpxopJS
iYpBCzUgpT+2IVI7166Kdw6DGvLlZsHTBM2ewL0ripU9cLja/6EH08XBSyrE3p+b4otaUj4gi56r
+RV3Gh99o8QlefYJ0OiqKYdCv3fKkAE4u+9cnOuEuoKnFLoOT8f4tTqTdmATi83iEKkGjSGoTH/r
6CuZlybEgfn9NciyRENZLuYG6B/8MSg1tuw8EsvZuUb9f11E6WUHXhHQpn+aOfHSkLHhpHRYl+ZD
aX9HTo6e2PA2jZ+zqryneKa2DQdEdpe777/MWOiSVVnKkeBXm/fi6+ifQD++HbfbYzMzkOLZFo7N
WK0N7p2QUu3NUSuqQXlV93TtRspvvZttpav2t5fGghnlpJ5hbrxtgL76Ju16uA+/daa/daJU3BTH
bz6VYGfxDFC+V9ExN6D7g8xfntgj2FMoHD5eFlafIh/FfvtPXKIaIZ15ISrlWGCiPrcjc8h+1j+b
k2CErmJ8e5QcqlWDc6AyyJy6MgHmhveGoUscdpuU5bUjRWc6Ldj0HUSIhLcNXRbCaozXrhEsauQu
+2AdCAYcEbrJ4rH+e/A7H93GMy6vWTMJW1BHYK608O1DMkDqvgRmoYVJr+IoSirY67lb2MkTOGKN
2NVJy+JL7HDiFkBUxuIcMfhUtJqgQLqqPNcL6VAxUoALYBQ34t3kZqpXJfYDQlzkCnmk4AD3a2qW
dmaPjLDVyUDrIOFpxlXRZDURw8ghkCBT4GmnCfmufOYi8Gs0P0chqRAidpYGzpz3oXqPEVZf6Qza
Ayi9ji0V/UhmvrK3Jsz/d43Yt4GhpPbgAMBvDhuVZCsqROKyR2q1GdnuXBSLTDhJT4vTZsP6sqNc
2woROKQ4dpT6XC4PiFpEeuRpO0Lwb6hoPCjmXeRTHTK9Bi/66eG9ZuUYc7aaLU439/LuVWoOD99g
yPB6vQkYWwF4qdqKvJI5GbzV07+aVOqfOE/rfUwIc/OTWYBicPeasY7UyaFqqou1nH7SE/f35lGz
MR0KK22ucSUyEOV6yxUwCMtX5VlqU56EDJNzvEyDrnhbPG5DgVn94U7nbIGTKQxtnKC6VOGSM9WT
9plkA7dmWPTSQihcS91HEobiFR6hzw6+2nVp2sqf0TsXj23C+/LrF/65A1CnPps31w6zWjC2cO6u
rmBGVBCgn7SO7Kxa+kn38q/0wXyH8B0ksZt1cWusm3i2Wt4sCxLxIW2M3FLJcGGF9J3B4fUdGkC3
gF2PVjRm9jmmCBL3APkxos92stGJTBEu63czC2tXcfSch79EoRw2YZXWneUA4oFTAeaHkyPinp3w
CZLeZKbH91J07EVaFZc9b5KKHyQsDGQswyY/Fa/I8RLzJNT41VsV2t7XQw7n9glf8IKi/sv1o+GH
uwDbn+F3gUJTD6rOE7pA2biUxFRlSpdG3y9ahbckO4LfY+3EpxCJN79Z1QNf+kSopJeKwbSgAFRE
8LuIRrR0C8zgtBJwtLT8ZWpo4PqT/akiwGIGFp6p0JwWa5TsVQiHPw/GjAfUsc0s20LgaztNyVtZ
ZDtZZhkeBNAsajUFmPNag4jW327yrO+8vwhGvx3oMV1ndzMvOJbh/t33CsYVDXQscPyuzfIxSKSY
eCIlbcjX6KusCNMpHD1H58DotHIpVydUBBBDWgDKBvM0/1IS5aSiGs1EOfSOjFLVbxKC4+wsT5Ro
IHRwc0d5s55hNKaBUpE/kU9hEQ3pErL7MrZgq3pguJ0mdytizDTfE9QROjePRsBnvWKfOGkPmPj6
usRLZV4Mz4CxKZWNW5LPsd8HqH9P3010RlKvcKoWEpFXu5/aYgZPE8hemUaYR87yHeJbIswWBctB
d9aONuzOb0RoTpZPlBYPFgtalG8NjY1oepags4G3WlOemb5j/7m1JI1fBa/iZfT+0Imz0Q35ZY2B
x0tWt9MhUys07UMoTszNGNhDfthfdNdzfT9Ea3msFhLro0esysf53E3WcPJKG+XlrqglguHtUuGi
SS80Ea4/3smt2MTKXRioVeL2sSbK2iWGGQVcHdn9dKd4SMulT/oJ1gC6MtIhfR5WUQ/cmfekX1Bl
1USidphJ62yhDcKEfkZ8KY3R5e5LB9MsHFPJuxPqTAuNYI/ROpZBepatYrNHHxN/bImzdQpq72mA
MDIyQ7pErh656dGbHk6+Jbw0+QjcqkVgCfwD18Y0/61SN+fCmH2XS5gBe2Tw0XPSlETB6Y+pJ6y9
baJkbBT5pS3cZkrsNTzGXPkA9LG6opTi11biGVIicnvXdSKMMgvklrfjAwSRy6M3lg8cr5NAn8GL
ftzy8s2yxDJ0qTkwCC6YkGIZHXwkGUaPRQYOVj3NZjGM6vdHFf7S2MhreZXDY29yYS4EaYngIgFz
mjPDI5khRS5fea3A5Hgh3KMLSFImE3Pg/IaBGMFx8QhGxKHxfoptWlTtGeKQqV+KbqsFMxF0Ch02
krOhdtHwMWns40K1m3igEffJlRCqgQU4CnHYeHXIilO0Zo7LQSniBnqryoHxJ3TrN8FDmVuumla4
mof0Uq+RYx9pMswpZJXLwPEdLiGNWJ/+5ic0sLrfmSPZPUYBDEKzkKWLo/t33WwQw9lgCWYF/GyK
XbLsP0PA1ulESVQnuK6ktEEkGCTZ+DJiGZZ7NYbspb5CzZzQ4t06JZIwwGf+K/dQIodDQS+6tOXk
YaQdup7UXsEKY7Me5JWEN2yPWwlfTc+4lYxs26t4ZmAkwR7BLtkp+KdLE5piqaA6CR8x1mWuEuYr
5lBOm+Y5mOSlAQo4dUvlhT4ud+DGIPZck7cSqfiT4BtfDTdwQ5+rSIFBSmnX3vnSp6lsqH5fPo4y
v9qPZoik/7x/Tq9G88VzAaNDVkmdj9RDTqOuGEdZtXQVROSHMjog9HpzsIrxz/MF5b4g/iVnhLYC
GTGuVWqPrm+yVCVlXYz9JnVwDJj6AeYVMKAc43+xNwEKMdVxiqssxmc/g1tYCf+ISt1RVe07GVjM
OGcpcKEAvBlDfEV0CMUm4oX1laSsLVsmF48E7WzxY7QldWNrZNAl1VXHc28MnA0yIYN7M5wyzGJ9
pR4txVoPoWW1hwIE5XLm5B+pK8ZnRWfHKwFbi7l84HzUPkHf02PvusJpREqWOgc8fruCipj6S2Rt
ZwYoSPX2IKtFMIw0Uq12H19DPLyg9HnKbE1UkZRsmu51URRqV+HHORjd7VllHWz+J6dL1x477Pic
hLDlTkk6+7bwvJkL9f7B0kXpi+rvh5Xhn9d7Hzs9Vfj+ANj4y7Lo+TKMIJvLmiGfHw30UlDsVeqr
PLN6pJ+CEGorU5tsa2BsySMN4rSFAsSXp0jF1kQhMiyniMs/YkU/O2nmsKVNG6jSN7lFyV5GTDDb
sDTSIPpz65+73AW5vQeElIFDc0GPsiaQgMghJgArSw6LNbGDlZ9p0M/kklQjVrX0rg7ot8PQlBIu
ZaRwByhUjflC/UUdlNxgfGSXcZX4c/CCSoVN6QXqTeddRHfM0COHrKZZWaw7q39eY2Qtcsa/c8w+
Atx3FHuxaABc+ceafL+o2ma7rPGsDS7QKDVzoCae3nglM+CdZ0J6Fi2PJrADBntqQxpSCN3rzYzL
/raROgNKwJawoTkjvjvxjGSN1+hLEjlLgNlMqjLgkBPyG8oWGkYCn4pK43SLj7NJBOEfRWLrdn5z
YV/wxiF3qGySim1bl/fMjDpSJ9M/rav7DXKiauWLKwUjFqCq1n5viuHzjP5rYu7gkCvQGM5swQU9
1gI7nQ5FjWmxAJbVqZz44Dqvp+N2OltMWo8uvxlNq66wIktYB49NR1CFRcKk1MxYq8QFLcO+ax+n
VeN1YWWwM+UT7e/W11bjApPEZ0UXs59JHS19B/ttp5lB1Qh0yzmG2LiJcL75mIacy9DGUcZ7wfXD
puTR8Vw6ps3yx9yxhqoLBtQeU5iTw6ZpQU0oXHYOi1x/yFxGouG2G4nVybCw72NFeSut6WYnq8Tg
WpqV617BEylvp+SMkmPAr/1//csQ0uipP3GFFCWVk4S/Ag9npqfngFpJ9XxuFhu4DoIHMgm0YwwE
y5qLgFZ77e11pNhhIUuw3r2ZY4JrmD40dhA7urtOyr5955LbvDwyBulu/ulmBmoIEqkP9P/qpI20
B+bFEep6a8sZ00utpckg4gq4A1I1J07S7F+WCWCmOY+lGgXSnh5sVwFRydu2RedHh1xlRM4PeBdj
TvygEIOSLIarJYmfJ1sLoO1+4jM5Yy4DZaeI5t2uwaB1QiSfsTPhF/SLtvK1WG/qYys5Lfdpj889
f1JUZAic9P86RZBIhmS68f3BW+pYgEoaDFu3PI2AXVHMYrM8W+oQCOaYPR8j26IecnLhqOFzySc6
tcKsUEeBbVWJyQPvzncoFBrGZFxjZsjYkuPtyPaRCirjqXtD2/gpUsrL7u9TLMx5SN33QiToqdrX
nypglfpxV1VUf95oklLMwqpgSZ49VmJoLgVFFOLVybpbwh22Re5vPAEO5R8XrR10sydJ7OlMF2db
c6vUdKKCn0UW44uaEn9tw57mbmGE+AsSGSaxWTpTMYx/47iossAtmvtEhhp7AAHXgwNXV9EqniGl
PTu2tW9zZJzCwHDxJPctcNVhxMY2zBTjByyKl+qUoKIYmKqs5WDlLcIel8XEO/QpIrjUFPOF3SLy
zzSgVJvZM/TalZczkbvxgFKaZHjoISxmp8ZINJDc4lzWvriXnZ9o8Ryf56H1821VDz/xJhrXKrdn
3ttfTrhjIwTY+2s48XwAiqrm8/yqLpvX2YoAW5fV6f5DoCwikL9qTNZVfzTvzIbCIPvn7L7dP6Pe
YagbsIVIafwNcy/0S17l41FACAjdzabD0hvywEaVwxBgpSkzvyBzlw+5giXjSWrbxqVMi44DnEaR
9m/BuX2prj6DQwCXQeCe6dxRW/nZv1WPqmspWTvzJaABNSB4BynXxysQ3kelwlaa7DfR5zRCDQbD
hPrBxFcPbg3IHCkXLgHCVB4UScRYxdyGSV+IL51W4Sx5Sj51Pwg7k217vyfAcwjLVjZ0EI7WcEk/
Kvl2BALdlpagxWaeB51MRhhkVlzcQjD22PBqyxCQ14WMDZPq2UksB5Y30ULSnAUYLxnUU3L6t44V
zZ4FBwmcrsrZcB/a3s1UVUtQOqfXtGNrB/mSBA378gm1u5WWtF2WYQT+v7aPHiPgpeVzk/OqFK0f
KzEwIafV1Ym/aXltIUxd/trxGLIthAh7qANhJlWoh3lcln3TucF5RC4HToA7W2RREOrB+OdoN0F3
Hid31Yc3ED4W4SnDnMrVa/yDtZbUQBWh2gC1XU4u/r7+lzyeoiCV+mHGMm8odI9y/DBv8Er/Z53B
pTZAFIQog7yambx0YCyAE3lIBkXK2JNmbf0PbwGqw1oT7Vp04KCRPB0LCnpgW3CuS99r5jWprjMT
bpBUUb73TutuD/mAHiU3xCBje/94/EUURxE3U5N5QaWW/fNt4d14zd17837cJJaQsI9vEAVsCTQ0
qyeztbnJ9TNPpq3H9Q4A6XrT28G7SBWOcdRzhwLx25V1m4EZwGmD6qmfn8XbS3+63DjQn+VF5+t0
YQ7NY6R9x9IhaVkEjri80MKcpCMUcRiuVdIDHNDAIlCUDWHqvkPYgs77+Ba6hsq/xxXzokYY4oyO
cDWim9FL56NwAVSZH19Nx1QlD9CSRw0KvG2gH3POsd+ad038wVfB07tDy9blp/ad+3oFUVUtuUdS
co/ERFM+MdJZGGPKJD727Q4vRYg0i4/t3sqRmtRaWcieTE10uA5RnYYSuXjB6QOtUEnLQUB/BJwn
Sfnk7KVYIe3Ufx31xu1f66vwby6C5QD1Z6QKmpWdyX+jrd+vRMNTQLrS1S53U+/6QIce9Qa+CXqA
gzLzBtad+HdB3wLgoxoRgkm3HHkP3m+J0e0dqw/bFaZe5+l1SclPPjqBFbudYSBip6nkyJNFPd4t
AdbM0dlgUf5c0gHWOQlCEcgyWYWYydNYPtsHXv/mZazQWJqYC6sHbgr82Y6xhMNjVRBH2V7BRPpD
msFwx8VbOeGm+kExo0TjKpaURvjvXtkTmj9Yk4SYmF8WSxpfjxK6sA/KSkr4P1pSdBu70SL8A6VS
M/B3OYSZ7sR+R0qLD9JioSBSX68sRjFbDCcssRC1C9qf/5kRiHTVmFnNiRi6krHKtgMrq7qhT/UP
+AolGokOXFCBwUmcBzBlb2Ek6RB2tQT/s8Il1pdpBbbwUn3BXZZpFTXcp1n4UMZIUkmL6agNhcC3
Lr4hHmrug+Q95ag9mmk7GsMCQxy4arJNedagCpc1qzChOoM4+nhLisjfRWZZ33z30bygGuZ4FC7u
NCkH6AwEK+ZGqaDquQmU0QlRruIBzeqjJF83D4yXrIG61VRSrCxH1XZNAAuVPqJsXFga94oBhXqY
vBOoMt0XRpVFNqEcskF/A948pbAt+Nc9LQySMz1qL4IQJ4VyOY56/GfFJs8HZGfoyk83kkb7eu3O
mxS5Y4uojKrjjJX/1bTpHoqCY7WAMuiVTQym9f+dlLvbDcbxLsGheYB0L4XSAj8HnfgMIL9vBkAQ
wkprDkzApGqCsONNlBGSnsYaVSlC7EW65O2U3kqlYwBW0UeWTeuDLDlWP8Pp3TVAbRItknU9g+O/
9j9Fy2gn+X9rF9yGj9nJaETi8hSVxMp4S2jcycFrCi1uCiwsQtugJgbYtrpiFqrOAZcDUuXABaJL
/GMu914nXnlHAEHowZE1ZaKbyKJ9odya5nFnGtprbC9jcUFsQwuZvSfVzIhYVrzQ7TxcVh0cCDfs
5BfdO0p5CgFGo02rqKyhE3Iq41CqrSvSQ4yMph2XYaTLr5dh3L3lajzwc52bq/7HQuPWlUBc1tpk
FNvIYjq7jcUJ6pRR6TuDAso7zZxRJGPZb/2YAGvEnwnSeObhRmgUbCEKn/ZHkFXbejrLwGqTrgjI
VXmuM4e1VNsD3Z4ZkhZQIxkVUwjN37/Kx/NCUnRcBgqt5IA5dKjRqvB6MDYEQfl+e3spyhoAysTa
bKOLH/dmrLVTIZnpxQvTwWVgfaklUKMuFq2Xncu24wWBwlOSCcFXsXeidXdJlHxk59DPcQ2E3Rb+
O/Cd0Nk8c8zZ36TEnwhgnyDFJcmrmifCcuzeVz27idEd+KrUddIFnbtOwkr19F2T2OvhDAHIMRc5
dGAglvHphwORpZSFd7UkNCVHiJEhVgxL7yruBMolOydrPZShGkUfYiYz2h4m9nB6n3Mg97shdlRm
pzcbmx4Js1DW6gkalg/w5SEyiP6pJyQ6jzHb1eojLUDP7hZK3cDjiHEimUzcj/+40RTHtlaaVKpA
9UlyM0i3SIJzabvXUH3TUc7hr20kJ+1XyCGwnZF4dkbYzQBgkGgxi5CYlJC7GH7OmKBeO7Hw24Jm
GKDlKk6HktN3EbCe8R2LFw22toFimJTc4FNPEj2wbIOMdK1lOj3h2QFEP/166IbU+kIhbRaI5l8G
x6zAHsjGy6m9OYL9aYI26AHoolUZTTJNmHDAX8QMzCEdDn5E4Mps2CIpxwUMCOkMlnyYhYzxZvLD
nVqgbM1j5E6vepsKQom2p95v+1J/CtGplxnimCx59NfR03Xq2L1IZ38Zr5KTofRe3hGgQelf48I5
V8wLZpfKSZJJWjq8/PLuxNe4OQFThZm50WUqQVIniBAqmcKSWRoLhJ6cIku+ieBKCI8EciKLmdFV
p531/f+OM4s3ebYxmw0kPBswPOpZEbkgJN5Z38l8JbSbKXOXvaVHu4MkFLdIbyeaByivaqbO0otB
5JtM8jA+Te4W1j70aDnQ0938kmKLyHFmFuUR8xKdkiNzJwj2SMgUbZQpnL0Pu26LUj2vt+qtyk12
twtYf+Dcwg5BxFF2hr6YcJ+pk3ArfxUIHaZeXHp1EGjNVnS32ak2KisB7QPjngZ07JEfaLMcO0t5
9HT46e8N0Fu2DMdUgrxp8rWRitxQQfntqur/IZU+3qOmVsK3+AH27pT7fQ6CwguY8nPJ+KrfZh5c
syO1SWFtsNIaQizucRiVPEtiV70vkr74H6r1HSxi/BVPk5oKBPy9hL535s2QqQar7jB0HHjXFN5O
zmOFSJekoaHGWeIQhQcUQgVTtAd2xY7nWkjxugTy1UYzcS57XkErbms1VtL33g/bfMtWHVQgz8mY
mzqBUGPZrtX6xDnwWwSzk6nRW7InHDRy1pHWS9qsWIRBxWtfOLg6GYJNBFEWDozRiQ4uaG/FDDWt
M9Bwy09z0/GNUBwNzq6JQKoF5CaREvOhTdJ+w3RB5r0xFxNyzgfYleJie/C/bZYI4j8hvuHgLaek
A4fl1ycdCGx6ZUIrbNwyPWu5KAuIK/u5giJEpCGZ2tQGqQOT2eS/4VSfOihqupd/YV6BmBjEwveL
nAAt3b6/4L4zsSSUlQEz6+LITS8hc8aCbSNAOIJg0ULAEAKfe7/4dcGAVMW3zgkhFi9Xfq7dslle
dGjXWCrfyivstG5x3/U+1v75mEitF0nTaWzid9iKZVp5y16G+oQyIzm2RsMz8a32cSAI6DEkfnre
7lb8xxbrcq483yEhEj7ZCTcYskebQWu8FQvTTCVllj+1QrawO+zBHNRIEDXQ7CiwQgLAVSPK7TM3
Edj8RO9lg3BkUqsFEK5EZ1iKedDy6w1LM8BTGK9sI3/vioEx3AjEuazL87xOSO2x5pMAH9aMI/+c
aKABtqKOtFrCCyrXfiNwYcevbp4U0dyn0vnv+OoFuTTQaX1I5LmWWXC4NjooJyxjmtUH9AKSE43r
ucGj5jgx3MFBX5pzlO/lvXlLpxGLM1z+z40AVjzif6Mc9AjL1Cg8Wk6KjEsvdUfOxwWlSeDdSxH8
BnEgd7txFbdIak7N3Fd4eYnWPOJs+U5HyWVBbZa3+IHaqd+8BnS742Yy0Bguc5Y5K5bw9+wmVQ/U
mmuKqJd11ua2VgMjAafUkM/DyFm2IVpySGdaykk6uyMHzCHgqoXMXR0HB7IBAoBPVImtoO2pdNJm
AbF5UeohfxwHU8SSBphZQlj1NvyLOCjh0fEcVAbK7IbHuPGxreOn/hUJyMrb7ODZZkt6lgB1h7od
4yS46XE7qwcYNZz7lCkW46dvAnm5T2d0cuCbonIB0nDlkSfNkZgTnSEufIOqoAQ3GmiL3gkq7ZCF
eA/8uwSpSAFRNDrzOoaMvTqhBDmBPiB4WTuWkujbym88mTtJ/15Eqj5QrU4WyER5VXaYJwJxDxhB
pGapQKGSBXdtkwPRKGA5AnsmpltVsOdjutP4n6Mo1QodloroBSIjCGr5oJ2bW/IiiiwojKBNtoEV
lLWyePSth1RIowgyjxP8gbgVumrYUpHbOuc/JtI7FDNKNQ08Zh93EdJ9XvyYv4KgwhsABX+IfRmh
a5lXTSBPUMU8Z+zkC/qbv9VmhPL5TjQzm2gGpSsfZwbamn8qS7tPehjtyG3RL/RvgHu+9TlvdVgs
SDrF5UbbdrwOkFyvzqW4WIJok/G3ySNI8uDVIhUL6hWRNqBpEl3/bdZbKW/AcqriU77PWzrKbwjK
EKy6N8pGD9fxtuNMvxbqNJ3i6IJfPW8SvDCE2X3c/+MpdPsgxwuC+t2W2yLqD1KyHGg2V+nFR6GY
GM/nqkvnDJ8eJHdj+YAK2bCyInQZf/+9p89Dt3kBil5ByIUm+KNNEyaVKMXgtqLxAXmxbURldD1A
WydgDUEQ+GfTqpAaRqWDptPX5W3H1RCN/tuiCGkTd34jtgE4dDGTKTS20JqBIx/VoY8oBphHAU/s
tDvAJIdUVqDGH+mlXUzfeyOwNs20fRS096DjcK6qJUgDahK+nbrcI9L716Dr6+RYaiUvO0Zh5ycm
KAIj9vX6ClEPMtw7Jw/VxJdWKDHIoL0ZeBKhfNxgMqPn7TVSf9VI7/Oxs6iskyOAtvKY7eFRj/00
/QR5ZnPQvDe6jWYAfRRUCL+p1xJAxV4VLfWFoPH7TyXZ23G4Ek+huwXN8WR61iHdXPByMwXuiqND
y0QZyGyeA5gxpHfALrFcdGyO0B29gS5gllX+TKWDEY0hmGx4+TNvxU7FKLSs59RZLmxxBq5A8RiJ
jQDKbpZB6QWeUoleH2u7w9adyzeWqB6RGXhlRr5UJaJAsgzwiPUjjfhTSC7ienHU+ey4jxeWEpLU
XV8RB4w6cat4F264Ke3+HU5t7RFyWBRNx/VzIywmVCFnWGhOZssR/jtnn5tnnV/nHdFpp/aszbNz
lSQOSTWZRgtP/PGoe4olCx9mM4+tSMZlemOYAVdJpCqOE3hf7YRjT0QPHXPG4sFYKM64vcG3NeF8
ey3kFOXJwkpNWp0KS58qmyfZOWP+uESZf5fw6O7kDbTZpCMzPb3iVnuY2Ou+MO+6CaFPCLFPwqpV
PL9RIqUaNPDztonvLEpbBNkr1C6fkISkRiQ9B270u+je7nyZncA0ybvl7gdREJSF/XnU6U0TxF4J
ITlxw7pzzTqidj0AS+CeJBOtI2e0paPgRhsE82Z54OYiH8oEAwoeGfLDiwuGsce5jo374tax9Bd8
lkm9LqGsZfuzsFdRk+xWxEGM7ouClaVrV5rDycbWjgt0BdWll5mKoD5lJ2OSSRBg0bX3C1XTojcL
ncQm4ps+LavBkiQgaZDiEYdOEp6jf4rL2JiP6CdZbPigsm/4X+B41yqgGAW8bmsZlfxyCyPJrDjO
zRNHO7Ad0cAToPwIOhP+FTZXz1Q4hrqsQGXIUOIFRnZqHrllhjBmJG6CjbNBZpx9da4hjNFH3RmV
mlo/Y1mkMpfV397GZI99KxIrQInZjI3fo+tT8tspGtDiXPmzd9vmmixLF9Eo9ZYx5SoLJeJgghei
rQVlAG44UFHBPlpL7xjfmD9GdZcj5A9Tjs8V6co+Xeg4YH+fu7r1TujRJ4ur6akKAAtatD2/DFMK
3g8rl9+vUsszHz2mpnFUKSVEEJdI8Nu5rL854jJ/DtEPq8ImOHv/VEKKv2V1G2ZjJhMiXT+hOvKb
oEsFXUG5zaBXlgZrc08JGqzmzu4PFUQX6rGJzajUxqqo6cuXVxOCDmImf+f3LYS0zTXqG5Fd0N2+
0UcQGK/18z0Hwp7aOzAnsu5PFAoxQWUVWPWkn7NBO8tL6kjoPdaFLElt2H5o/ogmCaCRKALEnHfP
e0dLepMOPuiyG/adOVNfhGoCK1agWHzNKGeZ3M6EQRzqm4W5JDcJ7llE2qLQH/TXNhzNtMAQtrNh
FDpBlAVa2de5honawCTVt5HSBLGSiwbxyF2k8xUiPT3CHbOUFmSmG1mkc6RzPbLKEB/U+sWKEN3+
s31u1lvvZL2delQZBJ4ysOSLkVd9Cfcf7UEHh8xowjaS79D+tr3P9s/vNJbGm+OfZnaTgYDFUOWm
ohccS5zagN8MtDP2lqWPr7qqgG7DxOdCjl+BhbKnyoia3PMzYnG5IU3iVS44pQCjtGWY2hPuWErL
bNkzNQVTTvbTIfZONa9aeyqP4fINitwLoujk6LQ/biGhV7U19IrtKGFtm5RVQ3IZM2f3KTvVlnvD
WJ0nZODvog0g86EpKnaKRlnHKTSSxEPRCDHZXNtj52xX/RLP88qsuTUoC/h78WGHzpJy1mS3roB4
6CqZo0j4pV5xDqMNADsOs8ueIAk6TfoN6Ojz/iQWfFDQ2Ywk5oDhskdgFb3RVU2dHN8yVN/wQ/QK
cp6uoDVtUbpeMhjnBTAL0XASJk4aYg3AjsytJyyLsIuX4SNFO8vhiOmqS5oGwBfPkuWluU01Embl
N4Ns0MSHRvj9UW8oxE0sUkCqYwOG0ixVI4IjIQU0Gje1aGheWUjsEYresRDWa8ViQ/uQuCXuBAN5
za/mw6XBxN+VHi8NTqiTYCS3tnOoPES8zx9kW6GFelNerBhpH2GyP7caOO6VIFzJ+548TyHz+i+6
EpHkxxbfLsn4YOPRs2Ldxz+kDud8Q4UPtVeJaCGJnHjqG15uPO52cdn5qNGGIbBaWF6OjpqsOwcr
q150dKYiSSS1ot3PhtmAyXsWrIOD/Z0UgB4FeGPgDwa04QW9Y4dthdyUip+SxUPQXe2s+oOZp749
uKgv9cmONBC1sTazwoU3ebCgylIYt6uXSfBO0EBagOJPwZFbc2kx/2W/ATSdNEuglHdrSUGGW0ot
SR8jwIrE7zSOJmSnYRiyXseZa3Ej7ZU4T6hD6y3tc0WbcEvQfaG4rwOWZ0dKUz2ssTPUgUGkliLN
ORpIIPReV0cdRc+oIzog6dqgJWiVHodXTL58C+VsHZ8XsuFBXmHNggKR8E6/5uInUi0RRzU4BmWC
KJa7Wh0a9Yzm9OIaNkahpHOce42kFr4UXxpJMlarRpCPUfVUC0gjUpfj26mCAdE/HQP8u/Ly7olI
kicTIgD5De0l0u/rd9QxtXf4Fls/2leo+CAwKIFmLTMzFK9ORo0Ny/4QplsGF6Ki3FgFLgcXr7Cq
2qGbMxTJk/z/iA6yQMp7XKgVx7LipUXCNF4B++6vqOBkZP7w+mLdupFk6khNNmScrjHVVaxyqnep
bd5D6vHM+WV5aU7qdLXcODMEm4AZ3PuR8kj7IceiR54/qWinvP06guhlbnji8xhh8nSKspUcOCsq
FVJLwym0OEPV/Xwgq2S1YFkg2M1sVQaxBQrf+vrPFa/mBk9unnnwnyEscDc1O9ir33cEKuyjfj73
o20GdejaUMpZwT0AuTLf004c3sjFKSwNXvYGxIFPgaaJU5vIyN1MdiuQsr3SypG4tQQ6wBhmFzRs
e0DoLUoVS/V/DC5772KnWTy3fv5LoV2RHQmLLDoDLSAxl3RVgoeYx55ziwEEajHdafOh3nCzd8hZ
/7EY/sHIqoxFGRPzom+LO1BiX75wVyEpG7hyJHLHX3MZsURSB8CFwmNK25oRVK9fpxD2IN0ne118
7Yn4XMx/xBk+vEGRSBY5Q4IXFcDXuFzLZGN071ezoxwnbSklbbnSpcrCTQgfmJda9xNeYlxZuWQA
LWWPBHfri3BJrMPf6EidCRFXbPUGcyO0Nn3OW+oQWIjzClSH3JrVM6e7furGBhhF7UlIqtDVznbV
Efpt3vfFU2uvJYjccDAbGIbvi6qMqDkav4SX9KiRnRNc1AhkWXpEpn35eTZamzaDn8Ca3JD1nvj+
clrfnKOfSHp4gXIzlBTPeNk67l6EV6Jz0GC9DqYKwOtMJzifiFM4SPh/Cz2R0ZsgkHyRutsY9sqS
SqaWub9Fm7kRYcA3aD5nfNwPZXQyO7IsCT6+Ad8/L9aGU50ZVo2Wj7b7RnWjsPfWvmav9rvTubXJ
WwheRmGwG4jd8nH3b6rIJVBUBxneE84v4xCNZjv2swyeUBX0p05VmHIB9kDgRHFS6kgyJT6jtmXL
yfSYB9V4TVNOvscId0+vX1o9VKw4op9JVrw4riaUdI0kH1pQC4qmI6CAkHC6qmiTKp9DGzYgIQ0k
DBne7aBZ5SuBvc+mMBHB/gTAOdo4shLUE6Eebvb9+T27QxogQwHLtS7ZaWu7r5CHq9ywvJ/PgA0S
mlImeA6M7XAnTpvEXkoRKaJH9AdjVkuLl0fxpczFfAogu0YFppQqugCT+Rpu8ODyaKC3s3sF51JW
1Y2r0lQRJVXejM+S3Mzc4g4fJR2CyfU9n81AwG1ZcyU4rt3omD0HkIRYPGuKLcczrKCU/uxujGw2
M2OfespQdjbCLbA0fgQErttFif/iBs8i4UM/YRaKfhho3AFh+NuRsDkS5jSqizovbPkuYnVNgx3n
lIkV36z3SbtnnO4Q2NdZu2nT8Q9n9x87ygFe9a6lkv7jIKSOXz4ZmS+F2S4PeVdK+AF5FkQdz1jj
fQHOEGTUsPm3Lje/WSMZy9VIkVAGQlxanN9Q9c4p2DJ6pI91Zmp+Uvt5D8gFNxn1r4zMcsFH9Ker
jna5lcmqehWGQ8g/c6CXWBzomDgwO9EHus8hs1GOMt2koivEutvGVqIQkSCe1rG2qDIwAtTdQfaN
D+040ZOT2f7TRDaeCnH9p8z570NpOHVmK3LCIjCc52Qe48uEZxAGN1EzpVrb+WowSasmEscCwZGA
pE+3b5G8bJGY+OhLW93sQE+SRNknW5idRCRvie8eihR+/m24U1EBKESwOBkZoLHepsOUG4iF4mTb
15HG4l015Dc5Ye3dgy3apn94CV+w7HvGuMHO6/r47ELhY5cLHTgWLtHUQfT/M18/BdbcgrFrzdTu
oHDtqwnCYbcQeCqxi36k9A3nC33VFmtZU8KLgF31y0iNHWdDK2pHk+uAfXKgPbQcm3ZVgqy8pSRQ
xkXPEIXyF1FPbXkAZ53pjd2FtEwfNghb5qlHsA+t/QQwomPMdhv1Zg6tpNOuyBm39Cn5UopsjRvK
GLb+EqeAlt9mwU6l77+D8dqGB+plyuzjPD0U8WSK/TI9YBDT8CvSYKkF53GOfPVoZ9Q1MRoR8bFZ
cz2VbpOG88DsCQloCBl9QzlbBRplfwV8rPD79Cc/d20bTwFfd3tB9Sne2trVtuPKN9Ev7aw9lwqN
t2cOToIatMePROrK+ueg4TZcHOZfKr9dFjkVc8ZhPsr3pYhsJZLu1NKuX3q01FVDV3Km9qW3Zxr4
HzB3LNYp7Mk64WH2MYpBGLq6FQEqKwLYBOzb0K1m9HZwu6l8KUlVjy/5qzSEf9G+xU9f0+hjNvmh
wu153vTRFhUzH9zx7qRrCLsHBIp1v9EUlZRM5xVTjE1eSDBcXtRGT3TnOTpEFgdshmAmOWKp4Zvn
X69EM1pBYcnYsd8562NPpNn1tBPUkau+zVRcjMVgerXaKjSwWlRjsa2b8sKM7h/9HaOIZ3r16uTw
ejDczpXfBybWH9hWREau5JaHOY3oegPi+cd2MAyfKsMadcfP6O2Wh2LJAn50aTZTYqznjmJjuMZB
Ar/Mdu2Mlctwx4ZChLaEI+mqajp07R7olC96J2BnR6Zmag67CPqYPEONPq1AYzxXTlLae6WcTDdG
lZOu2vrenTolvnIZ0g5xFRQ/qXSsv8Cl3CCZ1pve1iSMByaIiYHnoTXk7WqExw9aBka22FwwkmlV
o2spIv/cZiWtVruOhiNBjUVukbbGAeLEvXfgS5XYP9tUSTLJG6l1AQ1Xjgh8rk07iYSzfc+DUdfW
fOs7kDO5DehiaadDF/fMTNjX2USp0GEWTvTyi5p3HI1PvW9wGuHpTmzfcHJ2c7OqUSAmbveGZJB1
HxaM2HxjZQEHkN56Y3vRjjWU2ziTnoCFfB8AskWse7dSo28cr3NG7yVdQBsV4NQvTs1ooAGXVYk5
KjmNceB9UJzeLXYjS9d9yobnIVRPNmMxhiJrEhKavV45VQu1c7TphI/gZCbsEMdreei+XZXd3eui
lIAtM+xFwRUz53Q9gJ12hs3TPWHSC+yYkxhdrBfYJWM3ADcIxEXXlIJDLtA0yiUVrNXqUiYXUya6
FpCP50eIbyQH+Lp6kdzhOMCAikQLz9uXig9qcACm/al8d7gIYxryEd9NwxXsXU9Lnifz621Ufsfn
/pJMZR+owA8TePhOEwtWl9nG8v984fpjTSCQ3odl/iUduqF7nRpSctSJdOl+eKtTHovmU2L2ZNRU
vhRsgUub0JGDJWywwJfRoOyiPMTQpS7/mDWggXKYKjAe+Oc/eq3hTI/V4AdAf/FLAkja6EWhId2r
HvYtVYcZSpAhrHv0wXE8qzX9j6kxmq3vzQWlR+m4fjjbJs/8txxd0RL/ybHvt7Q3unrQTntZHCO0
fjZ2mQd3RfqXNNBMaqx3ZLB2MCMCcykzx+jDUedEcv1vmUEZq71GiUL/DEqUK7SJplIUDKYmAmBf
Y1agOq6ovDO1uofxLSMP+HWSRsmPtXdS6M8QqjWa+oNe1cmjI+1roTpvdMMrywwrKtszBRoKaPY3
O+OOyF4a88k0aU0UtGvVA+WFymykkwU16gtyfW13zYqIZPkNnk77RE8iTM+LNyTNY1YLEdH4GWEB
kdITVaHU+u4plJbf9H54YS0A9HfYOYbqEQMobFJboiMoO/kH30xV0OwxIdxsNURCzAl1w6A+jCEC
hSUHPv0cmFT3aGPo8Cn/RLE/H93Lfah7hPCak+/hGijNaAP8ICg/zEiXqChsjTxgbqUcO0VLf9pQ
CCy5RjL1o+T7oQmMLXYgZWcgoBS50OKrnGWFANYLP3Ls88qrBV6PHWvVjQUKcevY5VHo2WwdTlzn
QMwo5tIgMWUPg7RjSpuwX62hfSs1+hgfP8l67h+LZEJLV1Yb15YSEH7OUF1y8zijhR4fxVo6F//z
cctlDtF/Kh8495U+FbK9evf3VaNFk0G+mq/dhF8zq+sqz2pi6+QnxMdUjP1Quxg2H2RsR7keaIuV
Fv7sOgAxlXMYsDJEuUy2scxzTwcU0iZv7Vi25YwDUBPr1Jo5MnCsCq9Z9u4FdeRcS11CJgminiDR
AeVhn6Ek6j5//V5/J0GRafAcqhOtFP7mfAQ4Ebt9bVr1F8pbhpzfEkDQvqDvUMKCgKPN3rNXwTAv
tQoP3SGnTMfHZlXSzqFu1yRI1Q1sZ73c48ocN1T1mKPgXJG20d3FhW85N927+5dR4RRT0V3Z6eHH
PPNo74UphFJ3gMGQM7jifRzvTfNk99wh/9CXx+F8X0hapMrac8sh1unlJgp2IdBtO+V7z0WCmL2h
kpYGapJTcGwFBuuBxOKXYnXP39I5VUy32+Lo+o+JHEa/klr5JZWdcDLNvveU3D6xRMlW9rP4+rOL
iVQHA1dpmQoO9Rbyq9xeRKb1Pq8+U0d0GfAhJuLyTz2xYOvwjPO/nLU8m9pNkTd8rQeV1Ryr9DzS
xhVp51PP6ha9eXvALw6oCV5EPColUnAebJL/lbh+cvLBouVwjzJo4fy1jnq6n8Cc2sE7dIlPeYxF
adjbOQ5gzQ4uaUOnxKNbdauHDYR7I+4AnonONZhrLJnP/pJtXfycKF2/jylNhMoKc8l4dq1lTrP/
riUR+lbRXrCK+ERyP09VkCeJwtMiGJuMjwKNh7Ljmxpd4EJy2+4Aea1sQyadTiIbt9cEEoahR3We
Ed5I9aYG7N1FHGMw5KHsSz9SpomMFjEdg3ADPN7bokyUExPcIlPoyKhHNBTl/AXDATTHNeMlum9D
dW5fkL5T7O1tRZGucVp1KGy2M1AQ/xwqclPAYjwvhTUqoKCr4M9gWR076NfbXOy39zBRdUXUj2NK
I992qdwhbK5gFFwVdbvnNt/bdHCfW+8fayZjpbCw5YaOzMB064Gk7VP7nDSKZ3MvZn33nMjeEYfk
z5Ud4sg0t3swuZw/ujCxexkjqhTpk0l3wak2hJt8zDS/jOJWjsMJomdFgOn2dqRdzcf0Oqd4r6a8
m8dzU4Y4Yp34pe/BlFz9Q71po3Z2iLjMR0GJTaWNer9yp5WY2w/6t++EZFPbGBvsfklFV1ridA9j
U+WlIqBAeOQtVMDlnmVRioDFuOGFKhwRXNAHkRffcwviCcXMIHsiiPXlqM0dJOos/g5EbafIYv8Z
jJMwVcGzvMB7umNkeNQ3FzCIY/AvWlkPRIDouZb5ANkwHLyVPjpF8EGlgYSFBUyF9+Q6uTNZwO7K
8e0IhEkKcot06tHcmmLQWPcEU9J5ccDxXkvLfT1iil/eaawfWn/faN/DBb+nIivqmO0xMnX3gq8B
/1+ffmGiY3RK+Xvoh2vVVDfYS0/oqSqpvMAtfC7JioSghZYzoD0B3Ip1c5l86lSC6vB9TUMRnXHf
zepqIzN1cdQoFhSdpOd5IhDcfOrDMEwdfDugQDJC/4UEKghQyZhIbHPplfVC/UC2sKjbifpTp0tA
JYmRDzm12dLCXP+nfzgvtmT9Ej1Sbn6oN58+d+9Ji0mgWobSS1omUDmkp8UaZvaR5ye4gYPCu96A
/cYjd9zbw7HIl/Zi1hVc7HCz6JqVWwO/VIURbMZPk0p2PHuGm1WfsczriIFQlmVNv0ZEICk/zIC+
2AI5hVWFg7iAgKellkUNA5pRYjFWkJ4f7J1PIr4psoBX+s9/lujcrzJoC0G6g9jVN+0npsTm9xTr
MMxpyAK8hgY0R3pMDwyfe0CxRwYOHkcLMuyJzXdfxbpI9xLsHSP4NEjvKfmIiMpFISZhlM0w3G8L
RsycKnIYDSFFVNh+wE8vB78MY7HCilQfajK9CamqnTGoI4j7gPMOm9ScHcOIImE6Omrc0X0V4ck4
wtzNqgIga6HuYikJlX+QtPiM48DRCraHiDizOaVoE1tcccntT3WznZD7+M0Wr7if3L/ql/8ccxaE
viu7A/cklSkv4MMu67PiUyphqSunVUg7bKr9eQ2MMD/VelucQAozA57i3nCne4EC4lw25+gMpnPo
N70tqlLTOkNQlcvu86mYKSW7zD0rLCAJLIUeXzoxBZTrVdNPJ+MrPsCqU5f173eytAoG9DMPkVqF
iTHn9ExEB1tvV1tinoj1po1rfYYj3E3x82YBgoyPqn6JH0LZ8TuD/E94eT/pByG++dTZOhpWRVf/
ZG4UL71vHxa5zo3A5hVUzaMwCCzluOWrXbi0bIiEZkZ/6y+QP0s5v6xEqQ6yKLjTWCyaBxycSOqD
QQACc1FxQTLM197jzlQoM7gqdN1ViM0SK+S4YPSLIKXqSfq7CN/+porNB8zqkdvvQh4velnztkVW
GwP2Hp/ybsfVvpyI59hMOWgn8NyYG/G0f5DNN/ZyBlvqI+muVaz4MBBtRsp1DFdBFpQk71zEx8rE
tZUNyGuc18cueHJVkRdigB1YiUP8/qWUJg5Pp3nedK4xD9vIBVO1JPAT9MXxPJEgFLetEO0/O5Yj
7FuFN2l4s/w10mnYAEvEAh4dCVXEzW1/VqcBeORcrdOnU34Q/aIPQQrHzBTbsXHeXKFuIFm9OW3b
Uxd87JTL1HOb62gWqWE3XjoMPh4Z0nrwOJdxqm8KhpVUs2p4mhk/EaeWlI5d3+NyOX7mVUYpwQ4a
JvTljeTA3Iq6R+GddgIANU/unax3FujTpLpcDm16QQWtw4HO5M1H4p08UbI/T+inzNDeRLjjWfND
/mwyZqDw4BfDhLFgDshkYFP5oxpjG9B/DptnrvhIMVmty50Q+fCrU8FFopOWimrGrvZSONOnN8P6
6XjHcrfEb6Udy3aWwhwptLuYE18DqC90yaZ3EwMhvTeQ/2sS877eIyf5iVfHPv9Dk5Gl30rh+gxe
Zznq15qfK6kV643jD0/X37k9vccFnyUAkxRXMdcs3wDaYNukkEdSZxDkz0gq+UBVxA/nFoOKPy91
izo0lM3o6WziiRAjTo9HiWe1u3EOvEt/1ShSzdU/sSgKY02WAJL8LyAvILgQDp4R7Sq6p73/uyL8
9hwtEBI2Y4ch7AsQTLZclYXxRuBwX6c5K0sagQLI8DR6MkwqMBIZPmZlSkXMDH9Q+3YvoOjv8iI0
4r//HAGhyesIBpxw9pVwI06aNHwX84nptQUoQH76qk+mXpG68YQGOQYj//UuJRVHpZy9KyfhT1vz
BlUxUgJ+7cSv0agLNjsf2U1xljG5owDFsi8qKj69bscpq49FH2eMRp7LrShncJcl5AI8YMd8bkYs
RTN/1Ea4faYyGruWtLebh1IBklK1rLO8Ec/B/3EdKTguyu7RV8l044opvy3KlC//rv++AUcocMIq
Zc4f5KlK1ZO96Cmf5bgzrNF7kG2MWrE4nEXvEFXfYdiJgeo+GjMhSPHbJ9BADbw2IyCWORQ1AIGO
ZcrG03HBk5O5Cly3aCI6y38eUKsieDhWBAnq4F3Y3XVtKWIdlaVwBeu+iywT00a43fRmATzmowNp
ZuOLxHLlGKj38xRbg5RAFmgj7JvpRR7fKq+Nj9y3D1moFcwbuHeqvR0WbVVt1Kahs7KCbzjtImqv
w8u8CE+LARCWtH08Zn80p4nqfSmiU4EYVuH1GL0YcAHB9Qn+DVoFr293dkK4YpvTnaDoAVYqYuKd
VxSck5rFEJ2C5NxnXGXQVSfHJwoel0ZqBk3h0AqQELAAbnjxZXXaL9Kd7uqzJ5b8MRXGE2Gg8kwx
WaoQMYcXHNUimGHnZ81V2GTwu6dI4iZxs0jkyMZLQaFCmFf63VZIYvChtV1uiGg/yrbzJp/OvqBi
Lkw8ttBfn1LdZAAyd+J8kRBjjIDJ79XAKaRIEc6vm3SsRtDM9C3Pb0ITeFzvvvIPPDlwiPVEEvDB
6RA4yQUty7Slu8k0U5ltL3exgvlU+6f4fywnQFVm4ZaKFmyAEZaAiCyveNJapuzC1Ic87M6WKrpL
Ur45xKtYvHsAhSDcqBgS1ZyVcp87xwZ8l804NzAnniRlbYu48IoRght93wLnMMvz8cVNMt5fsovE
CbIAT+BR5kUEUz9X/KSLtlvzNG1XbtBZxJTI7AVxU+B6kxxfYemYL9qe18le2djczZ6Uv1sgcTrX
U6nJ+0U2pO8DK41qmnFt/jInWIOlP0FJp10ECbS87WrtA8l5AMZKhnuOjLahkPMId9VV5z1is21z
f8lJdnZv1ae8DgmXsw3lbkSM4owAYHaPhXxSyZ6/AYpn0boxugVAEpVlKnaIG0yRh0gkHBvEAbmb
6SXh9+AOkhDJQAn1kJ2p4ly77R8gawOSV9+nGiIXB74gXuaJwcZlFKpJ1Bu3OUUTG0eewWV1kGhF
yGAozqHCxhwnH7j2TrmXkE0Lb7s8LNTqqWNozjN4fEuY7VZjEnVWgn72i5elhQ2gTYUoP8ZTW7bQ
WN+W/1+XXKXbrWV818T+aS85YhE7AvPYHUlP4wgEz4OpvwmYg00DGy+WozUoRECjdJo1+40J2Ci/
b0qTqwQDZfFUnl3Pf7CdEbrKvXQzNFUr8grm+/p63GhiYlQN5EanoUX/Fh31e+FBC64Y8R7iNPLd
bCGFfSXQbo9SoTkrNhn3+FQ7Wo7BlHB+h9Vb5aUif1MkLxQn/njbPhk/OyGfIa0UUx0yPBdMt+nS
Y8uIJtkShR3+cT4ZDTafXaZm7oBes+TGpx0lKLCDLs22zFNA0pGN90oAyA1qLxG+2YtYhCnk40Rx
Bx0jDD+7pn1t9sLBDnSG+gSV3d9fIHulB4SgTNdKtHK0SrcI8z1PY47NhGjfaHNyUI/bPjUOGBHu
YSppNK+IRaBDb8w7h7kIDMUHNbPs7vmulfkW2OzwoMUpPt6FsIpSsIYNiv2lZ3Bzflwef2v7GQx0
emnfaDPR9nmjieKoQ47JKYzvarRnzOMkuXLgJ3mtKNWmilwA3no8VnmkXyzGi6s2O3qWNo2lav+1
2rQWbYPPV0CAGvWg59d78qCYZv22fhVWNSp6jRTdGEMIcgE+t/QiG5fPDEFYOiJEEcm5dxucIIwd
sC495vncY1vRNJsiNNX+k1V0XsfS3VwlACnVitUadXJbyIQv5apckmr/kq+Gpt74C3l1Pfv7IsKL
Pu4UMqYHd1yVml9lWSHsq1I8uLcJnGOqSvnl/AO9hSMfH0xHxT7piUku7h7FPHqvnpazd0gr8XTT
K/lAqYwb1r+X6jxG+soncr4xrYfpKtyctvqri4yey+poyE/tU1DgkTWxtuSqjIvNqSO9+oB3WyS4
OhvOzjKdpAAwJyCrh1gJ4tbp+oTAHNH4uRyoXWVzuP93qyeeFwHnfybcXgpRiyg9U7QZwCtmFPwN
95JmdUFQMIIPUlv7VJDWbLqhRx1Mw7N+7xKAjsJp6dp+/yS7J4Lzz8VwPDmdSloagcCww9RS5yyx
eg9bYCEMlkKAqptjNq4fIk+tM53OHrYc8Y3aGopo4DZkS8XTJSxWMuqKGk/qfX5V0OqYgDw4nnsX
PpEsR+Ofu1xVN4Rs8wmSbs3ABTJ2AJ9dqYOVHfax7Wl3sVXZuL2Ux8K1gXBBoMvSRDy5iAhk2hN8
gqX8FIEZlXfxOVY75RS/7MGqzrSbYZ10atoAN8ZNdveXWPMQrtg4TsVtg4nZy+JAnGgOhegTQb6M
x79qPs/2Gc0e1Thy7T9AcdF7hFP+mWsNRYLodjk2D1qIYwbPjfYDeGMIy+I7551osgKLLP4nMe3b
n8hbQYQ6LhxAWm3RIVs+sqqet84vuT7AOeRI4oepRURwZzjp6w6ri3sXeuXbeWKfUrgKuMnkV0jV
P3cYk8kncanDYsblRR8kCWg/g+kAAWLiEbf76zNXQ+hfHb8E/x3Km9IgLZ88q6UrICGsmBcl9C25
gb6eDog1hAVVa/IdWxfrhNyjOfwvuhZPCAFuHxvDLDBPLRnsEwjbZx6s/ODDsotxSLv8r1rS+BdU
NP1T+jE3zTCUdbmA21XtL1QBSlSm8sqBA/+tCadPzL5oj2FTXCi5+EUNnhzUxsMqDc77KQhgFNPp
caEMxWDFs75sGpshBmEn9xFW1v8KAILX5XfRjEfjP9ET8us7aljazGtEYCB7zQEgr5z26Xyv57tk
EvrRa+9tb4yMc4b2Ft4cNpBZwDx7hzUU71WPqaNTjMU4hogqoQ7z/V2iPoTcAObp4cFv+lFeTg1t
AWljQwWexGYfS0Lx6xV66nNnyupsFL6xb0RgzR14UwKZm94+kyyzSc6oqJAcn1HMp+YwMComG2lu
gWBSjCiignmIu8PZx1UhGMjfmrsFZg6llqG2Mq7WzjdS49gHCGl0H9FErgstRRoSKPF5oTbhonpY
eDsL8VjSysvFqDEdxcEf2IAP5BbQtFwBaKiRAuTuLUOR5wLGWzpGwo/RNmxStZE6vLS3IK9zUkQJ
T3lRScoXjZJ1cyg6gtcrZ8TgoISpE1K4QfS9qFLkHfyyEbwzU1ZMdHOdJZhxfcVewJLAdY60ordt
RbyDEmxSusGPuiWqDyAzjn7sDwTn9t9j+DZonvKuwy6o/sKzYAtd5wf+t6hXUVe/4405sb6yrBHU
+6OgyJCsW3+f+0mC+KbXOz6rUmXtdkSJxetBvje5rvlf2DuwZzDeh1YiUMrJoUKlhpyUIkSgp7u1
c+y3bOdX8K9OF6ybNQcIornlEdUymGlO4ffkcwDdHSYJMQPakJ7FM0hnmDA4ZTJwVnalKFAGsC7x
V9cyMmFMlyjPq0hszoi7NPt5sZgX0lMqQWxPC2dWBxN2Bj78UXUNtu4mhY2XzmxrBbiGuAyuQ1H7
zIwtR4HYwHFBBKT2JfVMXbQtQ1xbIOPI9y0qAb4dCBYf0x1FtOyf6Z9JGoaemfmbXklUydUaQkdw
RiEloAAptxwHAC4fex6in+04KH+aX/YNUGndAyaEs0iRAqp0VVBC4YtzDDzOyT6I1sVOQ8nIGm7Y
jcNBq8h+aF43EXqxvnB83cKWp1NNCcL/s7Kss3QWsQqShIetyP3CvtLM/mEBoA4AcdZGb3Ur8aCz
Hmqbq46gtGpnosZ7irRGWAdYdM0Q0Z0SM5yu1k2/F1ESNMPDrOJ9TPhECgzodd1OD7cKNUqGAhNd
g5hTGtIf5SHM5QsNyeC1UOb6G4St0Mt9F5wt6Fmh5mp19+1WPPJHu+adF7H7a2T2GWr9qG9FmtFt
kYRLahwFoGJrUFXJqMAugUzS5hkaWnndXlBvmvyl/hZvrUsCh4kozpu1+VP/f94/5tupcL8Cq4Dt
+VTpd+LDDZFmzUVT1d0vWqXiZ2e+nd2svG8DUmaiMA2fsj03mNPyxX1+1FMtsOKbX+abRbv+TfHb
00TAPpFwV54OVuxA1U4KEu7lX3PaVdHjrCEDtcQI/JckSxboFcSCmI29OTuv+yA1RX5ofkvJ1Cfm
1Rxy2BEBG0x6ttvz3kNG8mgpOynIGsS/q14fhCodj0DWXAMyXTeWgSf8vco9U9l7Cuwah+WZOp6k
NMqfgpz9wxh4rbEYvuu2CLPWvZZmuENYkaE5vx+SgRi2zTC6pAEUEtpMuAh5YPxFCHRUlyKZj5c4
WgqS2BmnhenPkM3U9vHBICQsC2+7qJaDnaaGXoUiHRrvXD/GUKcwImZHP3W7EMlDL/1aV6blPC8M
ktwwKZ/kUEeaxrGJjC+3kXu+WwZfTzv3EADLyC/H478I+q1zuTxsfO1LkJAtfNWC74DNNGgiKLpv
TgIVPzC8lFVxquH4AFkObe3mjC0PJubOU0OkKpcUvTmzUJ3AGRfMc0vyejO1qg5chHGbt6R229uX
Z2l6LwYkVCIdeuL/c5i0PGjAZCmOetDZdODGViRux+Odo9TT9bSPHXuZfrMucfO4CNc4Vz3YdyKY
V54952IA9wR++W7jHrdpEltpJ4Rw4x1YXcGQw66/uS09FPzcmfon6fKyMuxJTWCAVYjttrFA2JqE
llgzNh4Yo57Pcq9yGwXXYWJPldtINYzLOtN1O2na9CQS5XgCJ82KIDtRkaaQkju8JD9SuMob9qR1
Jnp65kvKmtJ+magmZQGIjhXMltqDABSMcjA2DufSsF8dG6xkjOens6G5X1ntx56bNbRpRSpezuwo
ON30SG/x+ShtJaHUniamrgnFLuaHPSbkmFD8QtGC3lDXCjjqQZei3g+Yi0l1S3uyAgMR+H2Ru84n
v6qpcFx2CFrebDbHMq0+lgQI+wBk++uIhxnEpymnlSjGa8Eo/kMi8nB2WB0D0KpJQ3jRiN3jlgJC
JMLiuOLAIITBD7r5U7luytu6quCXqQap4MwdXNVKuyg7vhPY/AuWmc6SBLo35fAVqj3YfiWAsIBR
j3Ggi7nvZkww4ThESx8v0ZTHMtUL9cHGfTOj1wgrkhwzdndbaz+FyWKtGE4QeuAaNKMeslddUQnq
bgjXRTku2SUik/HvBKucl1LwP2s7wStk8oYm/XniQOiLf88i8OF3tfekP6eAfcwT88rUz/meTgOn
C8i+0BI/FGXluevEWnW2/1TFvZFI35eSawc3XK9KH04OrVeVIt8qvn1mD4F9lwgz0uwTir/T3iu+
dph7u8bw5cNLmIPlKJfejxAaD4jsMFMz2B/O7H5LDScH/d0DrZNiJ+LovJjY/ZUd3xT4jIKUO+BC
mG3dTCTVb1643RVT3n6n/siXro4NA75Kz8iUtfdsYtCrq2qO2TLQKxAFDD743igWuW1rQe9OLogN
SxVVitwrM7R3XDDjxlAXqRnhb8NNOUJ1Vy2z0jdNf/KioKwTmio+ayN8TZ3tzhNMBrArtUSZYWrt
35grlDnzmhJ3s3Ap1PYQNKjnUUMXt/uR+YLaUKjexKT2ibzXiOMPGQnTziFMJT1NReOOnqqcifX+
05UYB5KmcwGY52zeTvnscGzpQgsjHmoz1qe/d/16mJ4mdNK99TEUwRTXQvbUg/naQbxiAoj3Q5E7
hX4+z0/Pr32f4myJAB8k3ot+wjg1CQunLDyuVrFjkjpl4XIin/7WMCN1eUQrPBJmpOfBBmmwdbCk
UPlpjTKv/8+DBKokyldFqlgu85cRFTpzDakEPbsrMri6HkaVvYxoclgLCDXON4s/SFyJsFVMTXsr
Rbj/1GJrIqAloVsWu/feKHXmVR66CXV3Mcg/dWMLFkFtfmbfz/ii7LSEe9SwsBSwr1KLq2Ldd8bO
uTKxNHioFE5btW0eEG9lce1416p+lF+rARnvXFdVZrtNHrgCsGD5C/5MxVyYVIt7V9Giaoe8pGBe
aSlINW+OY68FcV07LK4u7Dsx1/tHPZfay/o1KgKACnagdVZQNu1z9tw7m0Cl1OO+XgYRBTAce6IM
tVmUSUFFU8kKDDLgesy/oq3KWe0fJpQiYoqfvhLBb3f0sfE1Mfs5dm/RuB+x5XSrT6MygeZ+eTYV
MqgK2+ikOc+JtdyI0EfdveQFVnx0DT+mIJGAlY1LqB5+PRIa2W3u27Nkg8DJ3ySYNCLn0Hb7d/IG
HTjjAMbiOA40enRFPVdzE5YcXVCrWOg/y8mGRkgysmHRXSEb0IcuKgr5h4deRuKwRf0GKMZfFypH
9l6dMtQu/JWHDWNdbueWTtLT9u23Gxgl+nUxG9Fc7qWY49671lVLq1cBz256brd7hHezH+V8GY4t
MtrYiMLm0BuycgtvGVzWIrSuaNPN1sjDoHu3SpfKMvzLbJXeLElDSNVNQNNpYDgEcO8q/EQ6yFdd
u3y2wJjf6S3X11hj5kuYgD336byAaDqNPeTYHj8pLnc4Edzvnkq5ze3nEPs1SHRcQmtGngVoyI8a
2P0SaGXQBUBi7iRvZWyswJNWBYO6cDplyS7w+PkBH4HC/Ks9S712l+bKAlNzU+OEUAQDYCJjlHx/
MH9W2M9hYnH1+JmBulRQdsrWpewvMd9xHAV8enFiERFrl6MMzjwSvuR8eEcWvTtVTSxxWj5g08Fv
vO4bBT3X/7kz50w6bSzEsDRHtQR9JeR5+WdLEjs3ru2kjma0hly/QnXD5/uLdEjWkidaDDU9GhKl
QGQySb14Ss/9j/3tefDRSelHLtto+qvpRpZvZzuqrV5IJMZwky8IV5S2if4kOXNGOWxcSeXtwPWN
o+dC2VZ+hBmtMDTth0Sia1deBMRGM5KPYBVMyj4mnZVIQBpijfszBUJa0nbcKi/9cov1BA73DdDp
MjgGgXAKl20pKd2OKPXVT6gJ7FPo//4R+Nh7gSddnO9P+nYGCHuGDefoh7ecV1Np3G3uMqdsmkEI
pVppTa6nWv911Z3H8Hrsqa+A54wq4I3GBBEmtzcbS0Od/zJzWEFV/opcV/xhJ1ey/nIg6hnoUSHg
c0XGGyB+gThab03AccjUX63ZqOL+qmtsNrO2mokSA+3LKJbIpNM01AHw3R14Rjjt4XIHfax+F33C
FHIjECwbiBu/hKWkwp7lkrOM5a5mlSQwr9YoB40FHa7c1lqJg37/XrFGqmYt/R2YDzCR3ALCscqt
t26ggI+bAwOgkt7rDlqAu51gRQanSY4jaQDYatA7gIgUmN0st1WbQtGcbpuwR0tocAV3PZo+Ogpn
GlPNrHYMr4AoqqmUZ1q5jCV0srXCDebyHXD4aEqmARyd6CLZM14SKK5BrvBlcEbXHrxD5k6zEGPE
DWBVXbSz/0oOgHJ0FgL1Q9Fwh5QTtw9ra8MHXX2BUnZVjYZE2IvDKVWzkUUwRRtp76Ob6NsiLOui
KP6ariOdnkE83QjkN91nd7KtpK4yyxQBkOdnbOqCh6zo1iQbaKI1XmQr7KpfZ3sxBse0c0AGdeSW
BOXHX1teCO15zx7w1RaDVJmmfVIzQ1qlxF/2cdaqBDPJJdCvB3eQpauPJT9DxUUzjKNKaGaaqRYR
dELrpfLTzbABoJvDYCI2lKHRDNp8gQtwl8ofkygY6BgUSjHdq9JCDfuxQ3EzKxO/7MAAfL3Z7Wn8
ew4HBFWGkmTDM4ci5rqLeVNXV9s2aaGWHGa6ydj10AuQfmDetSs7JEBK0Gpdp3+3ae2jYAFvr3nk
YnshZXPQ49kJPWB3wXNelxYA0ntSk56wK9XKEw8AvMl561aDubZdLZzqcafRb+7+SlP9Y8RH6ZuT
pR7kxAvU6h+asyDBe9aCywGW+GUTfusk3MrCMz4g24W103vap8l+OSB/VgEiNtLZCpGB6QO+ZhdN
rXyNRNhwmjERUx4ySKMktjPHEcd/2jrxxJc9TRj7rpQSsXp9sq4mcsSAJMMKerNRokEzY/rU4pZv
hlEb12zD3PEsD+H9y9S1nHPBRaWQ8dnUnZY44iKa4vCtleNaz1XyZWyk8ziSoXnNJFgRzjFzv44i
ZhwifIVTU/A5yBiAA/g4FzFwvFkA7Oi9ndembPK8f29NK/9lvw/8KawknZvdz8CMeoKknjlEJoMI
fwAenRzWzPppsUXmprgPnTH1F4l6krc2euCxZaX3jII88fibOTulqxj4gxrSQ5l2cqscOxJkIVIM
blxZNL06zFgBhE832AfjDwBsJR/BICxmESkpt6j75rqkwGvQcBMv5bCrKZ7rHFxtSH5WOZZ1UIWv
IQgMdjwweyCqP44ZUDMfY9OYhIZs/Ec6/uMFqCWvyugoQzbvgxEaKfAUIHWsZyIkIML83b8KUDnZ
oofSwWvb/hoH3wb8jp5Hr73hdXO9PWp9UX++MJXobfa0GENNhbH0Xzi/i3GfVLmNTJJ52nRyEByj
LbiA1yt2qV1aJg4R0GCz889Twau04iPVWDxXa/tKMDv6WbTJxUo7ZxDSGX0xoAizUaBqpjNxo9hU
ItLvvqzr2lBVgnnaW1Kl+u5VlmNcKtqnvg7H46/tJuc3y1o3rddUvAkKwrTLMfp3fc/kxN4XMOe/
dapGg4J8x/cDgxmfLg58a29qFMdwcYF7Rp8F5evA9eJOpeI3VZA2Zh1CkdUlSVXZrQ63fToIocDV
y0IMIACG1P1bVTvE0xo2jApIU+BjkP1+cOOZAdHHgr44Lgy0oatnIglQ8qSMF7B0eRcUAiitHt7F
1MvCHcOLcuI+Ir1o6fn5uXVpRVvt42tUPwF33sTFn1Cp5tHWXkKbNHgiXSiYvTnmJ7Q7AOjFfkEg
qm/11rfMKP4XFFbMb1GzMgZOzPHsUKpKINiwmaTlgbYWoBBX+2FaB0M9NleLyNyTfCoVWOGfIiYW
BiZ3cq2zFVHpmFkaWvsCHDb3L6Gbc6tWp5oC2yMEadF6VihgqnHb8IFwsWBGvLOcravgp9oVrX8L
OsnTrc1WHPu/SwRPImWXmcb8JoqaLqZepPXk0S8afIhuMdG114NpqMooK7pb0dBjF/vCG8f2j1sG
pMAUQgULFcDOjJYHj38+I2PBN72SISi+NQP0BuO3fAWivOc0nAqNg2ehBl7gEmEH37vSXbbweh/J
L9boA+kQdg2J8D70WOxN6IO94EbR4MmYAtsjZRfKVZSv6K6ArKBLCNTNZ0Phev5O2vHvKTlruK8y
rFPYfRk4gaXlFk/pJDKqbl4jehPCImyVuVExdHm3s3CQArB1ELz4t8KPnj0eSxo14IoCUkGn+vZ0
E1wdc2wUpYjrryVhqGLPWwokQfnhLEdod26MxIlI+71d4JmXjYeDNS5H/259SOIzwK4C4j0KTDFg
vZj0DwJOPL5pvi1qfX3duG51AxIiiC4+Ud4w7x9PKvNahfK6OdCb9uhSJnh2eYPBc85bpgmjT3Vf
xMo/ClH+/RiQSLVbHCuqaIQYMcIuehyxyJt+CDkCf6VJfWlvH820Sj3S0oVJT4yeHiy8tLa1hkQu
k6+EhpQOG8toqS0Q2a7GOytkKDqhZZ95EnZQkm/qQGEyRZsHxdyiy5pdySbz7QQD9ksraQGEuC41
QxeK8SkPJrnUbEsTRo2SVwKIX6mbQt5czjW1dLeWeKsA0EggsHrqRgs/ZY8FQjd4xjnDhvIDITfZ
KuuPN89hyavV5To88ZFU8MOGcDdyRSRjggaNtcSaiIZbCm+vaB8PT51jVzB/FSdazq9rhbYpmqdg
aAqJNzXM+q86rHO8p/SYZoc/wF6oPsIfstb9XSVpeCdv3hYntIHYkf+IgIfBK+5tWbGJhmu89b8H
M/CjboSiKo+ewOFnZFFh60PpuOcDaurFEnwHIv8h7XCrrURpHJsWViP871kbeQQPiyABgD98S4Mp
awmLEM8Oj1eQUeWC9B7FDNelTkbGlrrocvafi5Cp0/vDu+w76s3lYltB13I5eA+4jFR66kuAEd/k
t5u46WvJZhykoYNQ+8Fc0YBdg+IJ1/xWSn2cNSxUNHv/qNxng+poyfQtKIz3Jh9w5MbemqOikrGs
HcMHLDLcx0e3/gy0LpGC5oE9LWmnHgGODUvJ3ToRkvfO3AyuzqKNhGt5azbuW27rk8JiOLmZrIFk
7w9WtS+ggX8ZTCwnpD/5vYdPxysnXrOhLab+u+ok0UOjhZ8YHFcZtOy2I1UZweCcLvDU5m1lPrL/
UQKyqi0IUk2fq2POGtH3sq87eOtj9UvV9TZxy/WAclRacu+f23quOqbANXUqBvvaVws2UFLdF/e6
j7wk82fyfiO2O0Ucd8CT6/+9q2FpABRBzlENYV+2dLBWmzzZKW60KMyizj/08gq/uIbrnWGNnN52
vxZ3OL8lYFJSp996btVpzhGjyByoi/OqVEuhWiA5PlyUD0vq1uFoBUkosjM5pDFmA7vHMMMMUfYN
lMbP6nMQDUtihwLy7acVyERRjF+imcOP6IvakwB/aKdMSUpCpJQK5rSNsOyWHUNxdJWmOvvPju3T
rwavV2odRp2aAq2l+MC46VdSBHyL3Y5jrDl9HdAoAziLkNpwki/mAJSyOIahQwsnAsU4uf4dDkSO
Mn6vpWAmzrK0PKjlBSSYOxX5MSjyVytZk0NkvPh4k8EAc19HPuFC3RGKcS/faKACFssHi8bLt57R
rMM5ki25Tt/A1MzVfmpH1mTTRlp1cnwm4Sk/Pe6yezFjq+Qe9xC5E5Cmyae4XLLFHOVLTCHe0Vku
eEJ9Z4GR3PX98cRmbrZj70PvVB4ZEfAE6ElUemB+/I8ti6dWcYA3qaILKuyB0Be7a5QtvHmNYBnJ
taUJgWIQm+yWDOy6NFjm+L6ts5WiYUO/mZJVfJrPRT+FZ5GjIO/AaDdw7jNvMn865NN1LjBDnUlg
rlIh6AGZvrlu42kjMhgGJTU4JSeboR0baSKkcpyn6j9FyQgiwle6GjQuYpjXOYrf+1RSvNutqZDw
kJnMr4EuBgXRtZBCmtIhk4JRN8N/AMknJliyIyaiCYPctLNCgicoTuLYYrX/gThwhJwSiMI9d7lH
u+o77zY6o4fygKfRLVRmRhw2wf1g01sJ4utDk9m9heGFWIkwnLPO18zk21Um2Mx9dTX9YwbgooAi
bac8igaCq8JuQBaBf9gNMh2RhEDou7Lo1cnGfl+7Az4ZGocK/mYdUJ46imFK2SA8/ZFmGJVtw0iI
4nBfrcNNsQ6P6FvKLj1Q436EpDxOWInsxZ90gSIu0k4YoUU/bLRQlxE5RO0MBnMGsekDdXLBdbf/
CEag2jCknj4edxqKADDT+Hoc5CF5JzUFsqLUtmMaqnyg6TC4e0uZV7ae7agxC1rQtyWosH+BYFym
hKEHvTcqBjePL8rYQnn7Ck86Pvu7E/Bu8jaW7OgJj/0idVUQRy+EvHRIwZ8QiIQ2/Uw6iYFcqbP0
ydNL+KAccJ4t+7EOyF50fR6SdvGGnoJoTbRSRMPhviDurt8OIZSDV/z86wphtOOI6wOUTfHk8rj8
PrD9h52oPbd5IcKj37W5N7vGNpjX9fJUlGSQ+MAE67vT8SYNVOTt2rKkwK0cJmpySSNUT8rNUWy6
zwXgLgmVIUqCGRUlIvvmV8JukzlyIr2mCyB7AcAp4yJQaJkrwsvSoGC/tJhVXoV0C29J8JcRgmal
dHnjE9kkgAQAWYJe7gEKSb8F1rG/EMKL6Wp3gCxjZ/6nVhEDx02UvLlQwJ2Os7Y7GmtouEIBkbkx
jJHCOs73Y40kI8nQSB9T1/Ueppd6xZPH+eoiewyY7DbVezAdJ8aAHhnHdNd4lZheh9eDVPayZcRG
B9jq6Kls3MZgq/DVjuRwM+UKxSeFRRkHvF3nrxqTuUk8/O+gD+wWkTUP+/cBs8dsf5LECSmBU57p
fOjwg/QeB+chrOHZRlXWeZpcNdvpv9zZpAwHDXO928e4PotJ1TlXZwgVSXNHZyT4s7rl009YyvvP
y8dCeyY60RbqhWCI3QtkSiJSHjRlhAfDOuDC8CKlPZRjsgtsqNqg1gahtpdANIvs9/KkoL65B+Kx
HrBgu7t4MKPWpcPhoFXzcZgDXpAMbGEWVMPAJc9UZR+TMAdpDqGD/qKl1g9a/Dx9qU2ojxgsp2J3
HpN+NzLZ1US7KHknG3GyQfSuZGL/pL0AQ+iPMOLqYm6tTcLnamP/uLHHr7WAfNYpSVQ0cUWBR9gP
UcDVF2T9mTROGpcfT9zZSf72jS/7LrZuZFGE5geKKL4cX0V4GeXsx4bm7jSUFEQ4FM34uvBWDEBt
6YvvgMamgPRfhy7Ibs8Wjbkm3HRw7Cp+qDX8r/i3sQLDbWJU5Px8KGWio58o9w3tXPKp3xDWkag5
HCsVRgEf+NF+XDpS5xid8/yd0lsG+y37MmpghhzYpJIaA5hv5ql505wrlIAoSJIkgZ6JIKI+38NY
Q0ZMRZ2mwpX0tqf22gU9Bn6HLguPCMZ47/hDZgceAUcPrsfB1TD8tjBFjcHZwkxeECZft2vpA9IZ
Pq44Vq05QBqJxk7LzDU5UsXoLJUqFfGN9c0fVnnHUPv5XiV/MK92ZVIOMQsSvhLwtGGi3TYmJOau
f1IC20+luSOyXRkdeI4rgsMD370opfdT249YGXBKM8CGzVMVKZ5ZZDTK71AhmX2+1hehAZ7IieVK
v9dkF+yenmzN3mCixRPvGPKzMou5k+u4dvxU0G34eriGN9GLzWiaO8So/G7cSemUxlyu4utHotmz
xu30rt1YspcL5k2ip+3+OWVA1cccGvCmzYXPs0WEFUUDHF+wDcpZ6iffASOFJ3jGbBQUgerF4Ag6
SihDmmxDbsMsVDO6XqB9cIf825VpwxpfXcU68Au3wbqsw4ZHsaBceOZfnUL5wxwbRyORmqBPkK98
g0gMtG+XGN7VeVnl8aOjTzEoj2qZrvQayCXhpVXggjPXz429HJgiE4LgvJ4z77Yk5KNwCZPeidFR
ZS3oMTkW5eaV+4dcoKUhhKjyM6oOQXt0CD5CGfTuC6JF1WjxK1rhcJgVGqQhRcw9zKsWdcjDTd/K
vaewmyKSwgx+TirXFWmZIsX8ma9fxI9kIKkbWgUf5gEa7BPy1qXn8G/9QHQg+zHFj+y3vMZAPzFX
1wi0j+aqJ+TpexzGyqAnvUYi1Xys9zrMuzhIeEr8it7VeQ6JbI8qx8gIhGqI79SHx+ZZ0C5DQliA
sTxdV0rTofgHfa8+qaV/KZj1nI623YBhHaCggGD7KL4MMkLTNPzDXb3WTQBwBGorbXxk7kXbo+2u
KeuGuwq0K3bqLueyqlJ629AlrequJn85WonSSB8rDMHXlaERaw0OM7LEIq3w1sb7xVbgmFmR2h+U
NaJLaSvJJDpotpDheNKAZyXHi15l9pkfraOlAXc5ZG1hcn9etJMJop5vDXFQUE3P5WmwnyzumEUl
B+xG8IZvyYG0l1MLKkC0jnCwPiR8iadHCZ5ZhxXaKvhRzhHOqHN98WCscr+aojgKvFSKi/WwqXcB
03NAkOh3aQ/HnBhwMM+BIH13ixyoc7rvNnZJo8zFTv7Ygr4ZL0EK0AZpYguMXWO3Ij6w17xelMdu
P2P301q1y6oB/lCKuZkD/3KDCoRyuDm8v5IW1N3XsCqqld4fk3P1BYmWeaZ+F8rE0cMVzbRStcKn
Dy7a89E+hHnqPMRspVKPhQJCxLUVIvphVazIeLFTuG5g1EhA2jZZTg3YKwDGkbAOQyWlRZE7wTQo
DL4CFF5+iTD87X15L09fzOGKNmqkTc1PVFVh0Qr9J2G6PcFU2hz0TOBrIllQWdVZWKCdbb9eZ7VS
EgPi3PVKtUHaB/86WIZJl5qv2apUR/AFBPjJz3b7Ew5oMScNtnz0fwvN0dzdWC5mlAEE2V6gOcM3
rfVHV+qSMYZLYrVzRVDPHB2ZbCDsZn6EiHWBid9Ki9+XFPr6SQBUJk19JvtyaB2RHDs/vNebXeeg
KWuy0jgpgpzWZIoaj60j4W9xO9j0Sa5k/XGqrHzBVIiOI1iJxZMSY9XBLR81gdSFGBeCVcntWYzz
erM1qC7crZdrLtCKES+LxPNfl/9rBvqq8tG4vlG4AR03IzdsCyf75D57cszKDX4+ABgD9xHGTQSN
McbknmaXS2k6ZpDWXvkCNqU+0PFFvABzhxEh4Hab45TuuNm6k0MfHo6FdOkbBFkj0ZGpzEZeIAPr
WVhpWo7lhPGflBIqj3MS/KaalYBoORwRWMFuH9OuGY6vMwyaRGRktA5+NyehuOJaRPZydKxcY3eU
A9hOlrkrIeEqhKSbnypNiONpvORhIgxHE/nxuv40TAJtfVSzpxlifmMMLs0ILNGbYyJ7XjPZzTVB
jUquncqNzWAkOBiitIwEi+bHwMI4ht2qO56Ag3EQYR4dx0iJC7CrAa8NZ0CJuw2sHf1QVARVQfI/
1VnBAq/Ew5Ire1FE48A5NNJN/PAwWFmBF8IExMt0OFqWXuAwTqYp1bRg5KH9Dvy9PYRtBnRhAWvl
3WH7kiEmSR8Ksj+9oWzqlIOTI8ImBxM/7m+pMxKx8H2hqyVjIE6uctjZVO6CVczMQ7i22rgcXmCI
wIKMYcrAIF7Hc1LKRotRKZwrsPlm+HsQb18++ocpUkoVKCfUczdhWQoYdFMQNRgSJ46JURekt7Mw
etCCSqy6XPamk7LOos4Jj8Vmhdo7gl/8FB74xIXvlzKKVysc59YsAOhqrcd6swcHoJzTjVEpLUJ5
l4B7qMH4VyTn6yUsVuzAMZ3kHCZlm4S9vxjiJP5Nr9MDe8L74j7YI3CgzLJtzqj+yGFr6FDUBcuo
kHQc4EDlxrylFUW7crsQYgtdS/ZO4A0d+4GM7hcYQsrU6L4U0H0LpUW5M3cJgcKoDrCFZ1vm/O2G
/VeWOn9+2cKSNnr7NS+Hi2I85q0UyYZLkq19k6lpHyedHEcLtpek/YmpJbgCtX0d50TdGI5Ue1f6
MWIuFtddbJt33q62T+xUGFOVPsLjAzEOdhOAIX76uwQuOVHbXsVY2AqzDkPfHkhRzfT1oHH5AAiw
WdAFEGxhNsBF3QrzNuGxYjXy/npA+N7RfICARtEHyT6GRTD7u+ro0S/zuNmqGYzAVcFrjQiGhcwz
TIAFMa2x8Wf4blgEu3VZh6UwMNLyOPaxcN4FEfxOIlnAgcHppFyY/MCMQ1/c16jz8sjDrXOJ2ELS
5TEG1GN3TEBr8xX6WFnOpVatXYOxdwk84YOwbtZYQnkSBKi7LTX+kluh94QNV1O5jBDikRE/gxW2
fcqQm9V0eC7ffmzlSjKEkX56bRC15P7XK9DjGxdVajAiV120l7aX82QJx790IRWk47CWURLZS8l2
VxHekzQc1bLaHv7gYMXaU9WdIPUlyCfumLcPwaBx5flVXQuLoqsUbyTCf6EqxlsWiIS+eVCHEUGU
JHr8cyZki4kbOchEkBGz2G5SEaeJhNIm3DoPiUXQpIskF217no5UehKgQ5fP7rJSqt14uKT4wsme
SgqWiEH70A+O/NTE+ajs8Rtk+4Bd2hvEOAifUNkFdiXYYf9YvIX6j+uymJEUvn6yMdnkweOFCcKQ
UL6KH77+kTR4S6NRIDtG/dUtW9QIIU7bYY6AjMFMZ4SdKgH5w1GzPbUGe6OB2cvraEQqg0UF6FFb
jxJ9/94yftHGgtTw1sYIdWXgx6NA0gxP/4zA7QtS6kKGcJ6j56s5oHzBf4DtaidybAZ+H+E1p2JN
0cyN/rW/tz+KL+rg6g8M82y5el70OHuMbpwzn8smE6Wsthyd3D63gwI0OI+kAFXs8dPRte/ufVDw
sm5gyM+toNVe2vnlcOooIvRiQcdIflWGLQnBnar+wCLYvxHCh3kS4fcpTu6r0aFKYkvh59wZiJVj
RBmu7By4/Eak5eNF3oYlAczAAhD+uUiErUyT0E6Xg3spSQe04HyCROp6OHVbIXQe9cCb8UcSSj5h
1qeVJ7YIKTP1tNo/+L6MQaZde/GyGF7oBkpoFFM0aUeHFrRbnQVrIHt0Va3DUVvaB9AXwyEEECHR
qcPyHHhhnVUQQylcpBGADEfr9webtjcayynYFAqMJHALadm9fOJbiYzb4vjTMZYVostDPELkuBS/
lpH0ZCUP+ioWS0piS1g1eHHGaIh2rAKVehFXV0cViZR6apLmzPx5RVW42ydNf6DymGTzen/YHxlJ
tVLMt/XYRl9H7d7vI/cb1oJwK1j1xOwxabrVIme8ovxklE3f6DIWHDFcbPp9Ye4olE1Fu/FYiVzf
UjG/4rH62i/IKMqqQDLrU5zyKGNJtw3OMFwbkwRyiiiNWpOjfYMYtGp9XRAThMrfxASvnnCoykF5
QRdQevgN5vDn1rXsqFP1w2pHdyuyrXZlfTSGTegUsxNANgDsshYvn07ylKZZDfjVOiAbWDmAfdp+
hHzKBdjELzEZ+XUBQsYMf4KRY/KSV/Ai8q/0YSSoicaBoLzzlfEQd6jKxqngo5247uME2nhfCxJV
MPdGpDs3+YOiZAQWRVVfWBEyYWiPf0u4L64frsfM2mXjrsO6sLQ0JOCIWblM6nz2hDvb6qddswmU
NFaHD6jiTqU6Z8eR9oEyozMqIfyLUbuWdPH4BkJhJ2sV8ARHEwrFqgaSlCrgRkqiRQ4NfoefV38m
ex23nfA1a609TvNWRIar0PlPWQRgXA8I7+BOupXLVDg2difHcZYx9zYxKMzjrYT4h136Uk8S3yR/
ZFAGxnaqzJnT+GjwNMjSEMRwZBzvU2uaB+2m7piOrEzqiCUyACX/df9A4YlZ6z+Y2xHsc8y1A0OM
4SPsMci5cGY+1kjfuR3lwgSpK0YbPBVAZ2a/67et3wcWefd8ZD3c6KYGWWVmKRwGPnLYs/DHGPmh
XVQLuQsGUjzB8l12SrnGxyaYLn+CfNTp0q+U3L2LVsieYTwMJkKaCojgRTtasSQWm080vnlpMZDw
k6HIQcx3jzmRMB/jk85SANDrcwS5rfu5aBj4tprZUNqgpY/eD0sktfnRhD6T/fLZVOnoyev9DvjM
NzlOMNV6LBuGl/UP4F4s1UllSkxWuEQl8hCjg0/v9oRLlT7ZWsCDz+92RGxMfXtvubKxXz+lQn28
ZjIZlalULlG0uvJji7rAIh3/Ol+NPjoELPHdUAR9f9sJndd1SIi+TN9ca2sJn4l1DvUHRpYbM7UF
5Tj9X8oAyGFERXo8TnRB8TVzqbSLv3GBj0vdaD4UkhfsVGC8KZxwq0c7VPLlUY55T7oLMcIHr0B1
3Qlg8TJPl3RPlWsbtjBB47tR3mJe+T6x45ad7mzRS86EyK6xbUfWcrT9bIz20CDw1BSxDYKq4k5X
if8rHeIYeSpTofrdP7EOlnZux6qWw4v6ueLOuLi7WhyelI4oeDQNODtorA3MQRTcRRlqV9t+rMKl
e1vAkUgP5tVZ8Vf0DxUEDSzQrCDXjcrTB9BMyzg5rlNdynfBXMinC7JkWz4ex2UVhVLpIE9QfxuL
1jmvhwPkpo8gAE7d4xoUTJywNEBsFndqs24AxW+oOoV9iA2vKETbmqUc2OyQSkFvk8m7xu0m9/V/
0doSKeXU7CAtk//USMXCqYks1om21Y7PJaqPY3mxqMQJdsT2HHHEIv9i5SmY9qFv/wd43Pfb0G0l
+ET28TVQqiBmHXpGMs53HZlkItiExR3nMnqi7g9b1DVpbiU7Om9SAjwmWGFXy8YldbDTW9Her4jL
JklzwGw8HNkz4Bh8t9LoFpZ1qvorHwUtR5zTkscIyWar3o/UeK1m8THFNDrwLjH+NFsArQZYgPKN
o4CuVrF73WL9fqu//kXqR5a3GU42saPOjw6z6DYaicvuGa4/pQ4eMmg8ztg9pRY4X+ZlyF8eI5aF
lvBTP/Na8pHurcJCJ9w1Arj4gS+JLHSD7p6oDRwau+i0WvABh6ecNHvzjB7bzixJg+25XpjamwSO
kFQQ52bE39tb73gdTNbiOva21exH/3EfZ+vPXq3+OxpZCNF1iuKR/Vz2/PrWqmwBqV5TOSFQDtcj
22VSVsKGf+gwWN31G9t5Ekz/8aiFlm3UA6yKjEUXuRmRNo4G/D9iqJmI9JiA8PxN1/4sdAkT0VDg
yuJYAk0H8I7NHmXSoeJdXB+PB424Hp1F1HsnNCrkMVNa55oa7LstJNHj8UEU2VPALjAxV8m4iosX
QuKVWs0rjvCf97P00lfNVEDyWuY6pjRjhJKZxBJzKo8zWPKVnYwjpjTEtWY0j0axKYKouXNwaVJG
aWRyRQsnRYIn0iSDwVydK8Dj1kG+lURYfQmppGpLnJlbiA5jPhGfUF5nDPlcOoJYtxagpBPJB3oW
mPmXXGyipvKKMeYuUgUrDzlsClFAv0iSQm5ZCPVNp9fccHvDzPfloMon57RiO0awajCaCzZsdTX7
G+EVSf5zrGsUUCGEPSCVB/Dn1e6nsvboYZjMTkyG5RoiOZ2qtHG9AjONnmfadm3P0MKYQY8Sv0Xw
4RPXYf74K3/VTXwvPTDykRKsdye1MshQOOJYfbx0yMlGxVG87a8xAp1sy59m3L4o/oYOYcTYX6F3
CbD2GpzL6S98Rdw14DgJd0TL+esL+sIGeL6DxlP35QmTMcFSvKmnvdqcWaq2IsKPvu6Kdv3eYEo7
vam/ey0vi5Rw+1aGl8MerDW1BTqXiFMPznJzpSvo8NTRZCDbsy/ecCM9NyZqiBw6UVvkSdVCYM8P
PNY+Glatay4UujAX/UGnioX59WPGYvYOIlNV08YZsZqYCZHxSe3cbly/rsvSAj/k535ZVD+ibI1r
S3vNmEXGnGbUYipjdwRpRrPJaodY8/DGjjplE4soVmgFuw4Nc3jc+m+AgDbDlnoM2fIng+MkwxVV
fodfX3Ya6o7LeWrzmYAkFRayTvE3I7kUSVFmxmUinhmOxXcLlHVV7nyQw1f+YIfs3tZglZfeiKe+
D0VHwZJTU54N8xDrGirnDJuvrZhkQ2VMPexdHXPMCqz6ec07+JrnzQ2UNJayb6GjK2I3yD9CGH+Q
25wuMcUIbaoiIn7oTNpGTVali0l0KG5Apg+ZcXX4ol2mle26Z5pq+WhUaO3qzy8J3v7ZBA05NSfX
jUqXOEhUjcmSTQx4QQcGx1TuoFyRdvcnDgRthpB34nEBABb0A1gbUqCOaZBlx/dxbrPAGzddfjO1
41eDk52mVF6B7jKhz95jlH3nPbRm3WE3TLYcp5sFBFqmIwu34slRqYVkJap/YToxJruFXD8IHofZ
baSF0emdN+yXZm5ysuBaQsP0rqWLiDSqm8M0qT6PKyx5dwYPTKyvVWE6GwZKVvJqaxOE5ZgknqeA
trJCkkMBgSD9pnVg7vBewDbq8REST9zxQjnT7wGE78XVqGyd566wUI5SCWQag+6qisplCOIBchAQ
9ABnOzo10oTRMUlGDlQErwD16kA1HDoZncMQkqKwx1thNit132AChEoilUseEJpOGmas6EWV+hcf
xLDb1MtwW8yUvnNCDXYPJvVT/onKYjX6GH0O72OOvixCyGm6CA9iPZ3ebXSey4tPR6b6LpmGN7HG
0ej/Cp3vJ1Eyjs/jOztjVpkRoWiepG1mGbvC8Ouxu6ZpSfHCSF1fcxcMqosDk0LzCNaLCrlneQYO
tO3k9C2Zhj7svsb1zCW7TtaxaunWQg1v+aCgUvzh4PPqCkzrYGFlkc9bNbzdso8CTEKlHyMvhb5Z
XrGFECIfU7EEBLs5plAgwt3mcCJdhhKlPOPs/xoR70vShBKxAypnEIoSkUwdC3ScZ3vmEvun1bpD
vBKtl4wwVx0fKLQQxAMRROSHfjUjkkNkKZISuqtgNnWX0MtIkjCFC01/d65HtRjrwAziY/xtvWXu
Ly7Vuxe+QyJZU853Lpsfn+1iRYsviZaKABv+5xoaWRERuiFYFHqX096UDCaJLMCTwNKa1/IgqEYx
T8+X1LOVOFA3p2999ApzWIaMB7K/4SVoczhl/HTbeQcAgppJm3D5bBtbPuMD/rgrNYooGUmMuc0J
GjhvA9Tr7hyByliMc7sGgaM5Z4l3wEuu6XaP4QWCv8joQnYQPg5QMyOtCtKQjT1sjbjiD13Lg2nA
hSHE/KTIu/51GoCXw6b9i2fvUlivQ2M3EcksRJnXAI8/IUtLsbVieKdcQycZ4ogyEZAeuRVEFXIj
Oqwv71Q8WnasTQfAPT5NKIQCbm9hhn3u9np1WXIiNw+ZniDxw5dlUX08lwfcG3vlrI8kONeHX8dt
KpE7JZodjfn5X4EDt79C2GuEXlkKUnMCUqLY+gGsiietsUa4pK8XMISbWG3oIS+aLajXur3RgSok
C1/xKi7iVXDA84dj11k7opkuIUOz9F0LZfBjkH2wQsbTFBv+czI24zvYXUs/z5HwX7RP016z+Dr6
7AE1KDJMW2p3lEKbdawHNrs/Fw4KT5ZdWAUc3L4XdLPedmzDRlxxpNpQM6WnkEamg/mI0Y2gKXB7
qJTUXxp5ZsrTWaz/Hv6wOT5duaWVwwqtCR8ZkirNS0VK5c1KPf3BOWgxfo6heUDb2bkCKjjkGTAC
jtX1508K4dIHIbrNdUMqJnZngpRlfGoz0FhWH8Qu+tvimg2cL+9R1S+5G2gI7pyQXpbFApIHNDD9
Xjr/MsszAbVpVGmFlFHkh2R+G30H0T0aTMUtBReA+oiUf42gS767g4L8ktzwV4mGQCZfZ83RW65g
tstWtwKnaKrWcDkRex7Meu0qe/COA157eY54+dkLZbKGjt/vFqWRkMsv4Yp1I7/cqSkeQryVNkeI
H17mLirL7s3PK/Nk7a9d4XRQ4znxrVWJKmwP2RslNj61XAx5FETKo5m48AWRAkiVCLgzlPa9giN0
GSvMI2+Hk3OSILwF8uCl22LMuHL+x2YqRnPjUVCHssB7vXAHNvNaZvgvXwzzbHDmTdhwQThi4TmH
vDihjJm8XH7OLdhhR3l5+4baEittQtNLV7AOOw/uwnxfKKm2z+aURryIBHaGu326bV6vnAQOiXwl
zmeR5bNIgYP+qYJuvtIev9tkvUEgfzbyaSup72v9axD7xoZwh/BbVlZWroSRL8nb5v4Hz20ipEH7
QCp/wyhQbQQ+9DjFaOfOytf6bsSFcwgSbt7HlM40AzV8K1oQ+jrlvBYGeyY3B3C0UTCRMUHgxcTF
y7F+45T5ZtEioZ6s3YpSFazuIRBLei2CgVjSvAm1z06TeDnDCQ3a+6U9rAdNGvNLIxgHAyphRq2i
nA6I+aWXd6U9KXDHXj/BgGHZaxsBpLZ5Bo1BeS+xRNEVPwFGYCTWlrobbAvUHRp+cY1sMT/3o7+Q
XOIONo452RciQuJC8yJu4Jay0NmRc/fwZPtOlUI/yBLkO1X7sPRafOx6E79EsHkWgOjJ8An/kr1z
vRmnSzVg97ROpHsUmTx3q7ClRnTxHOQF4ITpD+3mIcey99XsDaThzG5P6skveRwPxJlDgWsLgI14
T37PMGbyHIRVxK7NpKci2/gwCaz6zh2ZzUpqpB0AOXRtlkOmY8LQcOsVxv57FSZTuEWUKCpW5uTd
1BCFOceixBaAZ5cqjgOJHLQLzwkgCGILFc/HWGJh6NBcq0P8GeRbAeMpQUV4i9WxXkZbttkKul11
v+kWlISLBac6Y1MzR/Y/6QUXG77C1pjm9b8zIXZaF7X7ov293fKj7S3K/wMGd3z/XhC4aAClvxNk
002NK6PBph0Z5n6nHNNz4FPhCRY3lhvo48Akc3Trc13ZaGdH32PeFJ6MDoTzb/uqsed5CKM7dCQI
ngY+RNBiaxM0MYPsThpxML+kGVLulLXTY8KO4Oze5kjxKKHv4ANNBxgdt2VYc4e1AV9Tx0Uzd/iM
qIFvN4z9Zb36dLMeeWWmIK2T+DOx8VCbJaV8XK4Q3spICscxgwBMBSswEwK67/y+pYyJqZpxnScn
FqMHEBvjJtdguH/iQPXTl9//trqJV+EE2S2teIwxzVjQYDalBpN0kKZbWOgbLGhpVGckooYH0imt
TypFs7UpdNk8ZPzaZbMN9ZON1wYygG9l79Z3VxFcVDVL1CF4Uth3YBTQBmIQV502NoED7oyUwwa9
ueVUKG7nQanXDFxbn0PBsSV/uvPMAWd55Se2wNu3CFrnbfbekf6dFopDezs5MOxwn7Ma99bSjhDM
0TaE+EjztW33jH2hvi14Z2ZyuI3KqpHxw0jpw+WNSth1c8dj5aVYXPKcpXfpf+cM/dbsvjNAZ1Z0
3EBBSnzqo34wJFICsma3n9TEE39CkEwXXT9/g8l8qyMeHsZZalptZsN/n/rJnnJEOPUiPjmazq76
KD9XAXPQJY+v1g7ZaPu/FBQP0fN3OpsaidMErscs/raC4RYFacXccxYfHD5fIFjU4llgLeK+E/1k
jJETged4NlNdkw54u8+Gg/GGNaUO5hj+t8V5Dx57l1CjCOHaKwOcXHmat0c2ZzDtAlJtE3luOm21
wXnKKsrAj47ZasNYbiJ8dPwS7nBU4oSbfBE98rpeT4kc/zy/ecbW63U9E/L2ht1mJVlq9I2Nz+PR
ciaay5JNtfZrXg1X2JM6sVIyqDy6NvJ+unZ+DsUEPCMbf7wLhd3SjTHz5XlXOaz99PhYKWpdA41s
HQ3yU2Xwas779DIbhLX2u6Hg3TQYE7ZiD0o8zllvafQCOgPFAqJJozQ+bc0zDJS0a9yagqTpzINi
nSSd6G5+kVjoCq1sHbIUV3zTS5aJV+SrVWKRc0mS9N1YmewylmGpnyEGFEieljUDcvQ+i/0SsNJ4
aUT+io1JDhqztPhk4KYtm1eJ9DRdonYdFKM1n5QzJd0fENWhhvkTtfY1vy6AD1+M/EP3ZW+WsMvg
V39Gghk0lo+G/3XIsWA1oWsDHdB8rSlGD48Ie2eUXdgwQC9j4eeT4H/jA6ztnZMkhzQT6GFCwV0W
N1/AKeFSkXZI/Np2LLo5D0JcWbC+rX11SQKdjMivHEUeSQI8vTaXR1UyFc0UPTkAUYJAtI7nGCeF
aJfEQh9H+TGoLB3b8XQispQv1JTSzP1bDy8B4i7YuY+L4rThJNMXrD0OX7PKQAYlRUxsUXN8BdWs
Ow+1uy46ALEoF6SH88zCnFsV5G9EyWYdBlSeRdn2us2HiNwu1PPU31SOwie6wtf4Lv0wuUc2UkCP
n8fFYTeDEjqbJJKWaJar/Zh5sThDWMW7WEcK6X+KjGbyo//Z0PpUfsGYXVYmoJY7pdF/m8TrH16b
wix4vdiDH4QYplvZQpO8Y0V19y/ngngKq1dYNUCyFiMnlnvNfVYZqNEDzcpWnFrbTkel9ZtaePQt
LBjzvjsxh/kcspCVWVQGFo31MVCpROD9DvlB1eNX72GhIOeGaXpx3oNsdnVixcwCDjSklt9yyFL2
a6jgkX4lH5A7RAd4WiZRk+KPLGvXCSS34w7cfTE1xbeJwqiIGt4u7XE2IPlAsZXrdPZ8gI39rf6/
Yrd5o9v7CIYsKRPFOArSmWgfwt6QyeB9cxK2I1U9QauIIB0zIFUYWX4XtkUSAvPoBj8fwXyZ1nx7
K0K0WX7WQMHoQP2b94UcWMCIeLxYyJb5OfuC3r3S3rO7olXQyWe+TA7MuV86Rm91q34LTkxwt96h
Ac77c0F32bt2wszkkTET/RBND58XrTT5FRGEcOWHL0EKWWM4fkvqDvAmh9NWgk3cZYjGiCBL/54r
pN79QMFHnlKUW2ora4IK4CaqappCjolllbSaHY3cPN/x/YGBy4kmrpE8J4KMNWOgZljLEYhnSBqR
0comVVBIyNzvIQtxaVBE200DP4RNerz0nTgBPNeXNLHltUd8WkbiYaS1ksgXLz1hcZFhJpymVqbZ
jTotcIk9sapr0I1wwe+6ZvNSIeZcuUEvMuKfpRLvfHbFwMciZeawTUXlXagoB1AIGj4/iSGC1deY
apYso6Z/6J+SP+sa0QI9Xx2rvASlErvYu512S57k/uwhRGtOE+VILXWrZLcxSA5tRR32twgyMO+X
mbG1rnFzv2j7jqdrUomDgm/X4aWM1k7QYJBJp46hXQZ83DBUmiPkEpXCBgpbEhxyUvsrm4PdAmrN
+0vpiWGB6RRWuHBnFSh2+lu2uBRhJSlj/PJIXwtLNfGNsUHTHDyxMtysobCwVVjVw27NXxL9A4a5
JPYYv4Ln9IbETky+gSI8xnShF0uWtGpVIg3ZCX2Kfmgrc0D1XfD6NaQdBeMsw6hIOaucaUsl0HeF
WVmMjAcH/LWN+ul+g/+qW0sKHYoerxnzXUUc+29M6O0M1XejOuI7BozV1ql761J7ZL9P9PoH+msX
Lfo1AAYEYIA0bU2ua9c0ezZCHMzolioK2Hu5oOuig2cL/lmLYIoVp2LJrrvd9iVo8pxC889xt7n2
CI0nDjZZmq6nia0qeWzzUFGOelb3sekx21LevudIe5wKaLiYNAq8dFIiZbPvv/fLQVukfi+Tvshs
th/3mPvJe6oFQ8IJ0gAYdmnuFag6zIhONbiAnmgm6LZ5zGIroz0c1pHCD/SjCih8Lft8SeNwXtzt
cyu2tiDLWa6pWqePPbEm1RSJlsjnPxgyiPIrnNMYTBiYd8LwTD68dOYlFuSDMCBLraOcR1p7+tco
3TlfAuWZxaIt0LmfWy1zQTTfM6pfTeDo3GFDisgcpuiK1X0UC6ugAyFtnu98BDtG7kcoQJGvL4Mf
8kJfQxUuywRcdg63PqY3I5ORLyb1oWqwcVKCNzs6sfyldbDhLGtpAmnM+MEahQvps+4hvMcSlnUo
9Afqc9XyZKwvwi648T7eyW7uPCTeEkAV2xHD+fvxyZ1RaArT7Pxt+NXUjwnZuL5/VRjyRLuUV8pW
o+aHF4T+pizq2n5rcFlnP6P0AJqrzXFGKpFSiC5hMLtez2sDF0vdbM7qHZ56pIYro03SJ410CIgG
YubzuiAhStpxiKE3u/OXGRC3ZYEp8yzjSpqRoCZub1hHghaIhp94/jnc4L3r4VmdgI2lp3ZF+UE2
UrP+lQXQ7cZ2T5zjaEj+sV8P3OkuBmy3VQleIz5Eb5IS+7yy0T1xIua+85h7sdN7+moLKLK9WjYD
oYgPcteOCe2lj8bTArr+sqoS4KCjsr3xHfcMZniQvAcgMqh1/r5MWjHaBnrcIG1npKBqTZ5Eryts
gnz+7UKjly6vffDGGxNJs3xaybw0KXLj6fMLdQVorQ4BvIeXNo9Xexf+usvO3xB7n/lFX9JDImQS
LZRu1ueMWR6086WSI9/dBkp7F9f76ytKNuwhLKVC8981AtpdDrmoKx0RzfUMA7YwsvS2Jp9uLto0
aiwE8etediEpNKxsOdJR0RK+JowZpsE2Jaj3ZQARx2TOi2b4IkoMlDwvIGRHcJ2PrIukMXuiRgGg
0R6JvS0o0KOUqikhRS9eF5tlGzxmFuFY6U0qJd5VofVsNJOQ6eNTQ1Dv9SxYoa6MArWx9flUacH2
u2Wp7AOJMj0Ro0hADi8FKHYIQA1rG/bQYP16+bTM+FQ9s9pFXTcTnFkNJ9phDKVPCZaWe16dog3E
h8pv7cFtUwIsON9nsbHTX72cc5Cn1STvLqzoiHYYGZ9PjQcOGaHUZ/H1JZGXu3uFXuqMYAKcmexL
KQNdbhKboYY2+40LnjyIp8bJ9izT5pAO2ADOM2O9umncaJo8zS+iRVlwb9XDmDES6MQo7rndDxUS
iAWxdJZDF4SzVWMMVCVSmxfP0XGQTF8h30OSNCKs3e1X1PPHub7iW8qrfXF4XSQ4tCmf+eRjiUvs
29oEGzxfpwHChVASeA1jhTelGfXdiEdPic4P3IF3djdbaJZx4yGltCahqtTosYkWIg5km9AYx3mJ
fU8rFqcEI01pR9sgZIlUAbluIPUvlMkwHN9hRvN3T7w2o+t0imKeirqmFXS0h17Fm/LKu4fiHByg
CVZcI1p4ukp5tzt4Nc/Xw1xcMkOEAiFIbWFGr2uav67jJAj3BM2tbL1+l9XxOYgqnWPcFZCXQohU
h5GyF64hl+NAQJP8OWkCHZP/2bqlTgNSBWaBzKBotmo18f4UONVRUl16G3Xy+Bf9Kz3uZL16Mepy
F75S98nmaj/RSo03TSbXSu//78QB7jBHHPd9hYijeNDIzeftP0c6ANugkSl4a0Vmr6tU3P8nJUdL
rm1tUJsD9PlS8Yj3OI8MPrLerveBK5tDbmYcns/lG2WGYONDIUAYn/UKtIPi4V5d3uObth+0SPOd
9n8DJzR7ifIoqXraPgEEridIomDJNUd0qZUdcYjof4NJ+Le7EXScxG+Fbu3UP209JN+Irt/s9YUb
nltXzgxIIEcZjygqGowP0MpBznXxctrLrVqDtRRxp2LYZNsWkhud1HwufNEDKic2deOcx3AQlXj6
E+0WotNpWFX/5YwyK9ce1XzrQCZ7oTI/JkUjSL6qOxNsdPROaX0HvnXG2V0foQ6dZP+QwTGLTc7P
IocSJlOAmKY1MmNvpEMG531gjHXQxgDB+oN5qp35OCp5XyzKSuDr0GrhNQbcNv8/BICX4IQY4SZE
0W2+v5Sc6Iu0EGgtd6LJ3h3pPjBd8E2yroo304FiybvGN1xXkLBwrmXAiMsLuLM79qrfKSnQe3sj
kuDc5uo3AJDkxUnbq8cWExiXDEyxzcUhqpnwlwVKMUtBdU/0wXteZgD0ym4NsfVuI2jIOONVicX5
BeIUmS5wWW/4b86c3t9kNAtilkRFkKTcWXnZb3tionHHTttJvoizzj52X6xiMwwrK/P8FckWI5q1
AXyV5IGU2+nU1T3Nh+Bubl3utoLX+SFMBBnyZ61DfRwjppVfcsjySGQotGi6jwcycdvbwIH98KxN
xiO5+5b0ZVLeMxVliAtelv7sNTzoAmV0v6vEI1amX9a+8fTCm0yuO6lUU872w7XU+LtSNalxwYNy
MJpSr/IDVsYp208qeULNrGiKViFn1BIHe0nuy6flSwRpS7tqxTuiXGjTeDqADN/m2ICgNhgtZoCR
08QG2xeGzHZRaPZXivf7INRMp75DznMKBCUjp/OPfuexNwpNbhzCtAGCaLLV8FvVuj938ffj7zya
KJQ3M8v2+OlehXYe561OqMo6kUE3fLndyE/Uzca0Xgf/w3gAw7aWZFY0ZPjfgthkJdkx9HMvO0FM
JZW/qxJI5Hg6Qvj33zbsfFF8ZCSgXmAjihXmWosb14INCJ5AT5B+g0MwK72h9uTwMUoWbfFHWVIv
eX+yb4CjGjeYbND/er1QV6grCTJCjHcYydp81kvxVoKgnwmanSA5hKal5EDjMU6YQ2mKTU5EP/+i
1qUf3YCrBEN3L4r3N8Ex8gu21Lb+2z3uaeGq09pmvAl8Z+kvJONd7zxbATB203aw8bRjRxtiS/T2
00pOPcKpiY0+/Xrvwfys7hA7fhU3w17Xm1Ag6aVv10m+2blFqZ4OQCaPIyUxvu98c2C2F0IQJXuy
taIv7FyvOiMZlaDNqCfWezY4HBNCNuRrwLzEfAxXzysfThLiFyF/3Y1b/5MpJgttaI1nd2vx+XtH
i0VSY9p36h/XwSAc7pYpo/TjJsVoLYqhrij+hZLij2MAUzRDUN87cHIYyS79scMVnrlGJPsNId3d
8HCgKlzeqn/csYZLzoaAN2EGGx6x/KuH/HGKaGABePQuMUlkhnxzi44TPlyuITC+XDP2xtURKmGF
6psOgnRVJn7kNAXz3yOsLMQUc3UFKlfbiy0NDuMB61p4zi3HNKXvF0AU/FCBt/Pd8YXyDsiqP+46
YTTBGkWu5LeQAlA7o+VBDs/sMAmC4xvb3hw3vZBZ9XHAh6hFM6R+BjQkOpZGQRdm19JhaNA1+/w0
TH3mCPlvy9z467MpEbuaA/NSSIwz13WY4GyUfXtcDfpZ6aBZTeg8GtLRov4Nk5yAn40mlWEATxn4
vfiJRvFD5O4HPLNVs6/s15zVcwpPwsuv0qswXMcCjsg9mlilNLEV/5pGCinbyq/z/8XfNwZz/HGg
85OOEoCUMVns+cn8w8iP2zj3fvrZiRQFa7C+LNC+rSqMAJfYiENE4I20Dt9jARtdcanpoW51idTo
7QKP/ZeqVDtd3v0erjfCOvWQnpzrC5//gs9++5e/m0BnDB3x3lHMs0ytthJ822bqxfOSkQkzimR0
XGhLsjoYGm0uWWcwP2crps41b6QZdh1Jxrf3yf/OTCkPzx8sNg5CjfNWpBTIbfQjw9eX02IHqD4D
AXuABuWZZ7PUdseX2zqL9cbKI3cqYzeLMS6NpKXSc7kQrHQ4NmizIiLxPtyHTG2k6+tLxf923/h6
hLAWKvCWbvfXLLP3cw7NcCDIYSg6rThIXr52KZr5OcC1lyBdfeQGg8CDB91qD/WUhsxt3MNP/O3X
JnwC+4aWV9WFD1ontHwcm27WSe97ye3maFHuiHIDXIsE2StWIiMy8krYNrTX3iSnTqXQzFEoBhys
SQIVoCpFnLgftrC/0eSoVWnHsP/beqL+2eG7S1F70iXkWpZgJ2/OWipHxxXBOb6NOE6bgWkz8INC
hGr1WzgS7tL05q5uiGavr8LZTsuX4Xw6RWJEmwyprSpxalJIBoV/QNYVrCQiDcZZ1vf89P3fxxkv
QEHqFiZZ6//c39e+aBEzfzjI3q7Uw7WiZqZS6QTcd+s0GEMDQYb0lQBB7ZXFE4BlHPSpu7YmnoOz
L1Jyq2WnlUh3D88qkovgPxApdZC1FrFYOCLSYSItvWdXXINrVG4eod05rAWeCm9CU4iqw7/yRSD+
2hD5073zt9JOi86gZ6MnCUnmp7GlhywCgDYXMtbNPNooCgWopf5bVZ8l6KPNZ4hOvMvQJVHTSp3T
6Ymwr+u+IKE5Sc6RN9ZrsAMkfENZqgZN7yi8FjRKeCpOYvNdmB437iC/zzky0kfE8kjEnekMjf5/
qSGI/SEVwHCHSEfhsIVMT8HV2Is/r04byKNms8ni5W9Heu2FPdcedhEdPOA97uYq4r0ns0b+YiYr
qRrZU1/pVYJUK3ov4NIftruIXGzpdFCCRTxKBPKn5OtfygaBKZEmWmRvLUbddkcfjV9HS1K8Z3kb
8+B+g0MXpLaGUgmN0Xrw/AVoBjDLabYFeeAaWnBiAcOdrYaUj9xCD8yoS6Cf/ytvnp8EeyAn8uYn
teHgXSBTnnXBJRviaag+TuJ6x/bK6MT5Bihq3rP551/zdOeDfGBRpYTZXDIsHWHs+YeFvXYbakXA
mjVfBX+s62sb7jRzZtMvvwRel4dYnTD+IqhXhWHqCXXmB0JnWJrHgjzfblqYNRJuigxb+TGynrav
BUHgscSrvNyGT9AyueUVU5f1+FcpVLO2QdxvmEp4DF/6Jx1KoMNV9niwTlMVH+VOQgklxWC1QUgv
TqGqKNdBwOz+cozfmNV6VSJ3HI/N4aoB42n4EdNbBdOxYuD0ZBr+APy6kS/mKq9r2kiessLyQxn7
9A9T/4HmBYCExD3QScOGsFXU+cv7xJmybIreW3rMLSHSOIjmc+1BDzO8tzuDjTTMkGzSbLj03glh
Abx6VN6plIq5f+duXIaBmLZPMgN0+FrbbsKEyYSu06ONeqCGt8SIYx7AMIMCg8T7Ivftq+0JMcCc
4MeQWj9qOaKAb1BbnZ1JyMylXzAv3acmZSs4lJHSQlidayJ/1e9+TK5sseL95m1fur6u8D5f/N+p
V31W3LmKmOtwMMDsYgVd8nUnpU5ePGnALu1Sad4DKf9mtDBxXV1bZrtCHL5Pu6x7j9eSjGmqoxCZ
cLXkqOKB98tZswb2XG3jDQIx2Z3azumvOgOtrb4fMITTMj5yb9sJA2ofCL9NVLE8JrOJLtMREMNK
1Yo684svW6soiwpdYxoBtC1QDiLDsYasTFjumuXnULkcfWXEMEBPTuASqE9orUm4gRpXoUl+jQny
hHWL66xfPHzyPYIarFRZc3lc1pxuHVDYjVzW7A7kOitJcTeWelGDf2pjflZZEOP8+IvEypRIygf+
08b0E+7UZSO7YUzke7h+P2qYlBneCj7GAM1JIN7BOjIV3gpMXoiYuOp3eLl635n+jj6+vrfY5aoV
6Ee6uuS7VEqmvBRTlxALUW/kMGQDpH+z8PucDEdP3b2T7LP3yj6spLzmmqVIN3GyDhRxMAnCgADf
eJD0vTHJEJQsjMQsMb3/XiX52gNw3lr38o2BWutEHUcneuPdJiK4AzsQLRofFhKWvbmIbE+wWAUM
KFjgaOPxdZ6Rdkeu8i/9xaA3ztvThCua76g35kSjOaIb1RpDADcnPIh+TReTQbz3MDlglnUVMrXz
6t0nq5LYcksxCN5uqFilukcYC4pjqzGgbB5hy5B4l0geBsV6H3yUQp8S0Y6RX5iMyB2C2jlwcquR
FsM8hN/haZIvbI/FNFbhMumn5tkPomc2XhbhZ3zQRxVtT26i6RPX4LbpOzIN7XsfpYnvpy43K4l7
Y/IXIBRT2H0g7OrffZXlvYCCZ8SIoBtTqgJpc5fBONWOPKC4F7sXQjOYUnscrQhOJRu6/3ArbdtM
eDc5lOi8MbeesQoOjrlZRh5aMaDYk785oqoBClxfZwnf/QJuv1pU39kFTZisEsa99W3vBa2jP9Hc
L+VVb+I7EtajdN81Tkj0kSphBhztWYcEpYCsO+GbqeCI9QMt1KEhMuPb78JbVbKN5E4qgps8n0Ui
Fg31/fX67OkCve0DRRkjTki2sSKvWxE3UJ5uNPtBH5OaQ+RMBTe3C/OP4+kRrvUXz2h1O2GGx8fL
7h8xRGa5HQ9e7gK3+i03ZLpCchRpLx+xLrXN3556yYWzkVqU4st8WaEMlSmKB53JJIepheF7m6sR
/UPyWk6wFhzuglgFDTJh4V9HX5Y0/2Van+S1EiREwfhut3ObNg/6HFvPsBBKDteTdlwwr4Rnj05t
0InP7RB9N/0K1KQFvVLfkW+V0SFrXkzv+YQIEOykV+mUifBqlMcNFyGvCHVeGSYlgUObY3Rxv9C1
5Gt8SQl+BxQVKgwhVEJ4PzQtWNHnlZ7lJENv72GlJ4o/ZmwpiFHGVGq3l4jo0RvVnCk7CrXZjUj/
MFXxvKRuYRBzUNm6kYntDmZrl/kJysNDT4UQGd3fWxZ3pkEbgOzthYSVsFxSOoCUF4zAfhZlDTfC
7J5huJfUif/DGmq7r2UnpKl2mVNlqNC2CDSGJ/w5U4+QBaZ81t/m5U6plYQ3rnR+eKNxNIj18UFR
fUT7Nmdn+gbMYrwn93GEG9SvwP1QsYXHX+0J5huyZp82mOs5/7ONr+pzw7L+SX06GqrYU6CgduN8
FV5TalAQTTOohlg8xJdeJNxqoI4o0Hwali8IzeM794oQ097fXThbU9TbI7vS3jSVbq1csy+q8ZV0
gyhBG27T14vbXlEt+jm1e6aKakfUTfVgo4CE/+1Zj7e4qP4fCTvEaZz845y7uWuYSDe6PASYU0sr
MZZgWokIKwur/Ybt7wFL3YbLkArAOa0uTruXInKnHXYvUmxkPnRoJXn0oUEKglMUyH+aNtjl+cZM
6a+5Ja9+C6KqMqV42Z9BvACftyDpRyc74tnkOcx11iFJeNG59OnfutpsnN7CMl2ohchAOTUQffd1
imDVEUzAuSCl3HSPwH8we+Z5m38n7xJ9ETw7ftNKNPeOh7OLtGtoKz+M/r9kQa7stN4IELdztcsz
DA4D2JS1yZ4+YjYoYSUzCtMxTxTc/MY6dRsPd5CrB2QUy2r/ebIAq4cBlankoCb3NNm0YnwHp161
AdFTRtESShSPVVGVvRwlQ1PwshEViOo74vgh46N6yVn9EO0ObtVB/Zjuy7kvqT7/jCuLj/W27p0z
+tTgYxVFHrB7QbmRhdzQxbxnYUIUZHjC7b2QZVGVhG49W2ZxsAa1qld3Qotri7At8YG3ukGJJme+
/ImcjPC/gJq0MCpqRc0B1ZsCIxoKjzVuomWgzvHNDF+/IUvLGf+pFM1Q1DruzsmtfCaebJb42pzq
5xs3axaZIDs/Wc91mrOgJDhsBCpWZnmf8+31HhH8EqWerKDybVolR0NxbCa0sWBIVe9RJKTc7ooR
87kmbotpd61LJXT5RKMiBZvgBqdKFX++AxfHSquBRakiqIrQdMZh0qp+CINfKmR6aL5ij/txlKix
PNSrowjcroAZCOu7Ei8V36yuNNSv5JmBhX1l/aoTDaq0LRvw07Xiag/9DxMGHxVjz9RclOdAKE84
Vhh22ShSJMX7fSg/6P+qweDf8DZeX0FQiW2Bsh61BkrmBDKGvg/ObM/5RDeJBS984bm0epC4Artq
z0410pWgwkBDR515nTfCvzlrC2Bgl7VBU1qfzM+wg2z4iq+OtBQaXYlQdiNNghpknOY8f13h8vHO
d/sMsNlFSeA68vCn877PLzeV8vQ+GKhZL5IOQboGDcoEeyGdmDpXjq2ilKLxNLMGsbXXSIyjkqaW
8VBrQOO9peZyWNQm/2LQUIFQcyn67oz8s/VpYnqXn2S/zoqbXxgSdIqHa8xwo+f5Yn6n5aWMdLOP
wVZ9C3dcWV36kJGWSRh427eaCEQ3WXASyZU08r13MOh4U1y/pa664hmLqjUo81VJN7KeuUWYMWc0
sD2gkeUTjLBuV3oO4ZSRRI4/5ULKdFnpdR2+yMzS47bixkI4td6pG3sXT8+zSM154gMCzCG64eE2
dX0NBKFuIh0D+hM7pPDbBntepoSnxz7MqivcNCQYYcDDhritb4qQrozkZ0g4Fa/CwUzvgrd7/o5j
UhwtNupyHcMA8g7eoiQhAEq7hhh5dLEbq5t9nmvXLid9qUxApUk7CfuayRsevF3UeKOFoL7KRjlx
QPt14gEQFwVu3Ao9vSVdM3d++EKz/gVYPi8eQWj0nt1p9euyr2ybczCakfNvYn33VisjTCj7cDeF
Ati2oIiFCe4oml2TXZxKsOHQUh+DKvBWlSpv+HW0ed5Tq66Q0vfrxKBghcRPO6M1kwPq9Ex9aSAF
mCshdW9jW7x1THthZEWLyFiuGCkCAwkXRBtz5hfBezmcdmB6IUvm/yirLZzW+T+xdaN7WHho4yyF
XEejgRPeG1XBFAE537kjwN2RleFJVzyp37NHJ5PvqFaMF1wa8o5888Vl6A4GNxPGKmlbljqGI3F0
nvyZfRuiPAa+X5wKKuG5LuEoI2MF9MDcRHqqkZWOeDvssvX8fUlK+Jo+mggff9LGCYBPambPcW+u
izjnJkmX5mIOCULPe4U8PJymIEy8gWsuLXXFqDroXJ2QgeYR0F7irI+acXf4fmrYzqGECWaUYAWb
65X/2tCw3X5my5C0SaUa/Qe0w88wenrpK/44U3kxJk5AGm6WCQ1gjYJlySi6sfdC1evcdP9z3p5t
1URcj68w4ApIOlFBs6KohKvbl8SJ3LD53xvTpsoZHgHaqjdGil3MJzIWLgJjZ5mKb5jN44a4/L7N
4uwvuy7reHWJ2NCziImOoG1ULPnak7wF90ts+DLmSMPc/USV6qcV1EpADPHaAk8pyDsdm1wIBz48
MkOGCtkx0QN7oRaZJyuZabkw5XJ6wBrBKD2h6yLr4l+TT0GIfxIMQuCS7iLonC7+cfal7PQAt89g
aYANDoWea8OoX2VJ7ZpXPUPxBA0W1qBMoxPGv2rjVpGEAX+gBsEZqq9p/18+1eqhWMeTZ8CJQvEA
tIzmp1NcpMoHnn+k16jUIZ4KDlid9xpgwuwV7ZfCgg294NHDVbqAktCCxPmLB90S6xPJRSaXWEgO
cDi/Q0v2eviYLwj64EKMb8F9+yoXqOTnb05t2e2MOsMBzQqrax/cUZyplR5SoeJ8nAnV0hpWmS5+
IoafJi6swQnnqylLCDc9pQPyfIFX8kiN0IHo+GzxhjRYhiH980hLc3uWIfkbBJa8q51SfyRjN3Ow
mn9GYYQnU+DLox0gsEVkkdp2CeOLafcf6G5Vu9QWzqtqKX0Vb8oGClsPQJ4lXeSoE2P2r4Z5MnMw
Zp8WPmp6T56y78GHFefiv68DJqbYIexLf+4/Bb7qxLeGni4VnOMa3UYI4e40DR1Arriiwkzpmv2e
YvgsvcnBFSBMQavs5JJ8xIDeQSvCzTab8HI8YGqBfilyNl982ZjM9pV7bKoXoWyKt3nOcy0vGJsD
jKw7Xwykefe8rNDTOIu/Pn+Ffjdvi/P+FRANGjcj9HtAtAdPl4+fInl9t0wXgQsOkDPsLdWAJr6Z
hbERDxDAv/CHmWktXJQpcfcmD6UVfDdSJ6SP5/qlGAGXmO56uhtPNuqiCeEX1BF1DSPzfgc3lLc6
diKyRgHJV5JGfoDM7GdyA6AEGnlvMigOBDUuvuBvgkbpgRA3c5UO6gIyUwaO7NRO9wg4IzUSuTev
zxBg4yLD86FglPhv33Eg7w3v9JZEuR1Z75nM8/fzjm0EarXgGXpsm6Cz+2DnJSNTZHZiXLJa/uCs
jyLIoZKkK8JoDzsmgLl/5S9gw02o3e8pDl81uR9WA4z3ZuVgZQcE3KoZx4cUeMvDWEM+bbffMV6Y
RN8JBjC5jS+ml9+Fdd5oqPBeozeVPX4c2bKHrf+FaR6HI+TaJtENE5sqyHoAKpnU44JUXNmKhWPY
FZX/hWasudYLWF3XLZffYwWuFGrrY8dGB2qBG7LIY+6YLCURFpza2Hl5iSI0Q2r7mReTuRS1GSsm
oKUNRYH1HFuqHjhJfRfhKHp+FAmqa1gD7em33xxC1N3cgYRifgkF5BoM/P+0cVpxy8sC9afBQ/5m
y2maLvPFlG1RQS6H0xj1UZcJvvYVJDllYp9ZQV+AIkAad8AhxYxizK1Xnok8udQZdnJkzu2qnnDL
Os6yzEgM6d2gn0vGbjzoYmlYQywWWRhV+FvPgW5kBD71XoJbRFWphnEdwaG0jjOq3Sxvihg/AId5
/RCfJ3xsHpd/tUNAee5FO1+ejqovXZWLz9Gsw9qkhG05JBCFW4v7XvJRq4cHg6OdO8jDyR+UO4KH
5U53OJfKjJLyDCRkk13WQDbTUiEr4WUQ71k0l7WbbFCB3hpGJvzcXhX3ZWy3OmDtGTEKAwO7vX3X
Z+kfYVzcIaNymRay7DCBFnNI8QNr8QglYG70sbxMl9bRaf5ZNY0k3Xyxof5fwC0hdOT2aFB38k0g
cHROxKEFIn+3v71vKJVs9jg90XVawUseM7OE4CTjMXQD4dG/GRJsHE+2e9i/VC483io/3mMm6YzE
agmiUJ7fYSAJpUJgFs+JJxLjL2UuNqfr/dOotu2Yp/KLCdK3GXG4Pd96yaiIWCfACb3WKNC5M07L
dhzC+1t9UHBLDpDwBXBa5nEK5C8dGavw0cQebZVhFu+iHVf4JcGbLR+x/hlNjtaxY5RHSCutz6Eo
m3MwUUt/KizvdaFcwDTxBj/2FZgE6tzWt/kMV2h0oNRIgF1AxRnwo1IulDk0afAbyEfvdxejEdWv
M8CpJqzEURkqtpnlzLijiwAYgta9Jg1MqmwU2qwP9C1cKiz+Z2HHAkaInRHxviRVsFyGE3xcUT/i
gWc/ktkPO6jg066P7m20qU28WCeiVx2J+FBtjt8IyYa15mJZwrbdI4639rl4Jb/BmW0R1pz5QGuV
OYRQSDeAHrriSW5k0BkgU2Adt/0f0Ia7dwClAmwQlUmAjdy2D8KmW/fGK2iNSXsoHUNh13ZdE7nM
OfQue4lWhO5umHAEfYj7Pno+usRZicrO1PowZS4xefBs73rPxvQWp+dkiFK/1c0MID56kjWETinF
yTHmxyVVTsf9TxhKtgH5IYoUN5edl+LaJWoTA+Pj2WUB6CJAcdMONJb9a53RSdsfr6e3F4iQ82VO
CBUOsGbCRAVchf7qNP+Mp1rJnqdJikfuyZHDWvvC8YSrAqcG5IHHJHzTVAwhliEvLMHC50EoiXGs
U8zcPZUqQsH/3Ns27Or/f3WqYOPYkUPHzb34OLdkueFLIGHaxniipJm55B3xyuq09l94Uz4bkiw0
AzrfnV9wJYlmw++G5/tDBlKIOr5kmKxnxUqu5Ynut3ZZYldLFrmeMI8iX7u05ZSSehgBTzwEVu9Y
CcVVSXpn5liSShyUFmzk795vyOx9vV8xA05RSydwoEe1LZzR5Nzf6i6Eogpk+0lykC73wGy+db1u
4+wg99m5/IpLnN6W4IWP1TXPReMXdhQqEvSLavx0i8RAk2Ws1oF+DH9dz9+dWB1x3EWofjPRCanM
ZyjJRXQ4ZK0PmHzy7vnSyRzef2QqtQIjmhCWtIZsIw6HBG2sDcuhbMSlHZsb1qBeUckDCcXfDat9
TIzRbDyk0shnqtlUUSGZuQJnLcUwje82Yy/srsRAw7/k3/pXp8NgTiSXcbjIZ7JJx6ClnVBxfQ0K
GVSayRtqXmpIvqVYuY7AvWyqtvfj5nRdpOXvWRrNbjjwJuewWplIvn3oeKT2weQV3Rp2G+dZfMLY
OXWg9DxHc3iRmZDnrg+DS9zXeXZ3XYv6okjtsQwLaDqSzg/EVnvxg5DGd7BS/TXJmCukmoZXUp+O
FF2So3hOJnfH+TLXA/tbBIq9CDlteAOf36LtjfXsJ75PPtGjduG+mAj0rcWH6yPeJcmAun8Dkrr1
WrUZC0CR0MfPI7A4QSTR5NSKWC1pDDdYEfT1sanNyhDdpVjASMzLk1XzKj77ZJQUCs5t4e89BMD7
LUvZ698I+IShu5FQ8i4zOVyI32NrJYWOj8/cKuAwozl4vyNZZcwbYvAiIb/zs3Movi/J765iWyFQ
ehziMSXptK/nTaDfuZHT4LrPFQIXLg4PInljyTPc9sOrSlyhIDyQwQTZ2tEJbKD9qq2HoeDb0IHI
JyhTPvQvmLEtYIx6wc3xA3Iv36+1EHcbAdi4NUa115SJXcFvtYkWL33+n9Wrb2aymT2MKifCwqSW
V3jjLEPPuRMFrQg53kw7YIsZS0b/rXs3Y9K5y53VCOWo0Xvgtf0ViHD/yTvP/paNeAAGnB7JbKgm
Z1qFmz4CBho+s3xoCi+KTohULHeD1vv5g2jAwVN+XTRVyID2IkdLdRtGaTI1qkbwW7TCswIs0saF
hAz+HpjGQyToo1Sl39w76wWSGh+H9JUlEpKSQ1446xd9z/LN8726LmRPtL9+osPgAyoe3vUp+oz2
ycd3l8osfngPaeOqbvLRqRrttLOrh1R7xxXZqOip06k/bYdeXWwgaZAOuXJH8jtdaeIYl1FmbRWb
vQDLMt6xQCZ9fMB4F+tJfXfnfEwAOvFuYtZ8Eh5KXC+YdcOpj2UoiE9uoj9IfGyxOQjlEb8vCIbw
GrHfMtzsj2F+AP4zk2fvdY0GpSysqzvZphny/iYVk681/z6K0IRjiYk3wmgAHOacz5iG8coc+Bqx
KBMc8hPBeG5CRSgtrwk35kO8w0zU6NofjVOASELfcbRao/Phg3pFiSM+w6DFdkeZVLCgSsiaTl0E
lwj7X6pJMNukXUxil197C/vcQGvj7+2na7bbTTBjFY2PajFOge2wVNMsPSkTdvTUkCPr6iI2h5Gf
mEtFeIqZjRLE7svhELoWqPhPESbiUz/f7nN+yiT3qi5Gwjh026j5biu+MrdDrSXWmm1XS30H35GH
6mkutml8wV9wMyhEPywgjAqVl1L5L3k4M1fKliKhGJ9NCz9qekcQ02trP3dx9XLU4HR9gPobhJr8
JjcoL635psG/ap1Yika5qQ28gJW8iAG5sSDUBjH+m8zz3WgnMDlam9wLqWNGiPrKgiL8qYUT9J11
RY4rd/mGMJyGVyZQ7k4TINcHOIYBdfqkEA3uk4anCQkvR8W+YtFvZkx7YDrUCTAAjkq79usBzXHN
tjGKrjGZ1qe48ClsIZwEbX3s4wF2qrWL2L2eGaGgQMZgkF1lkUVwOM61qzlsy5uoHu5dybUQtBMt
5JIuVhzxWMyKK10o4LSSlXM56kF+fEGt36Awd26Vo+wmtumNhbAyAbdwzipDB5KVXvu7THdhtKwz
4ZdI61MdERPjFJJ/cXizmA4AditUvu0xj+KVnO5zYKqwC1h0AZz0aS+wf8ecPTfDuZtSFMxIWy5K
Ng+ItHpPS8x5f1J+5sdEDLH6bUglelgdQM6+8IjcK4o6cqIqox+hNNDWuU1R0XxxIu8077XaCErw
Po+g2hTeDPwdqKF0F///ZIzfC47HHYVmoBu/ZKc2zQWm4HLkpu9kr5pS/8q5ohrgdnQU7NNl2Xl/
llfIeW8vqecpsKj5jDeWXVahqwVdpNO7hHytkJMoWExxylN2ideqaKRN1mav6AO9mLC0C4HNIkqq
nlQ6ZQkYbqjyMOVbhS5qxOGExb/fqxbGgvyBhmZFfJzMcKcDHhh9fvTh6/Ks/vEb8Ub5GCwqtBBh
1mkxrLja7dRbsnW+MoyGtQwub25skxTL2dvXI9jvOh9KYPf/o/wOeN6zDWQD6hSqGc7ee2rW/tJt
w3XiKhEnBAaxYOzh84ohfdnsk6KeYeZ9DUL1ImtahditpUhrfA2ZtwKIzz+wvTEnDWyhfB+fzqep
za2KAg9dCzxIX3mhb7RJMBQFLLV0pXnWuS81Y2VMiKNZGU7UWYEiMOPaZubglVGIHhvNUwO0akg9
9wM+t8ldXR1m/T7FYwKX8xIi50Py5k9RVmPOaOLYBB/VJyrIJlZHtrf/N/Spu+1dlMD9MSr0tXX5
zCyuGLsa0LtQgTK4DXy6U+0HrxeL2AQM59HN9GmYt2ENNFBMhJU/DC8uHL3Xr1rLBn7CZlbD3fqx
CCd7jGEdRqOsnD+kmWfZd/IeOeL80BktQIFr5iulbiZ/hE1dsGuaJZeKfipJWvGo0tEnHuLCmI1j
OXsZHKAkIIijwKWAg8zUfGBs1dRFw2t6UYV4VMZLr4/3BmF5k5aYzsPbjcZ1lkFJ4WkyPY1gkys8
hDrIhZBPz/2bb7OG+NolcpdWCR5GPAgm2Mr/l8EPO8gPQeLIrhN1uM6IFaTkwdRZDrOMfVt8+P9A
oxZ3i/d5oc7UW1uxT5BTxoGITqVNKyRaewy3oEoNPI4Ti6LUtfZVSzmKYYAlu7t5HF1Vru335rgh
BcY5XE/2onGHhaS7dNEb1k19fR0W/hZP0aDgqpYKN6D9mNdQGMXnK3SxUP/NgU/9WpOT3G0GmhW1
rFV/Gncmx9NDT/PwdZxWGRuk+odqDGHYY343jUxwRPJa+c2lwZfMC6lwC3a7gwpL/xODbm2BZmgD
3w3tCQtVCTWAsd/yQZhtgIm0TTSfkQM4ua34D68KagOPA9k3Ibzb2DzyymyJEIIFq8XR57DoaGbG
HwtaskEgo3TQhXOZEmSRCYQt7zZ1hmm8fUo6OcdBYWUAVWUMnW/yfj7DapDuVK/leqcJ3VUF/KwS
BGSHLXk7DM3TwcyDZksBmQXHXKrtHWrMfFBCfaWV49gjhOGppX7yfUhwFQLGmrgItacVqj7VYWzR
vbUCLLYYAyurs3N11dpGoiO3C+D73Tc5Dr5RwXaK7QmMuvkD6l2t/uFoaZEBbhS2LL4pjLkqQAYz
lVC16+gekDL2PB4l1XaqVMQ1kjw/LuWhakM4bTzkabGYYMZUNgep0NYcrOiojnNgi4RevFeVcp9q
wPwKdL+QUPnvHy9jAuz6wjYwBxGYvNoMJcBGzYxiwlN6mMhs4GzKhVc7vsaXwXw+fbOu3QxHQgsf
J0au2R5tY5S9UALZV0kmyNSRb6kRqkTfv3kdYyaC4PeUkmqA/PoVBY0SpMBVnMNo6Rp4pHmalcKF
MAa+goiruVFPLrvFQSX1wOcm7WQFJ0O15bTwbtey/RWhO4wWjACZ9lN4C3Emqfj4TFJc3a5UCP2w
BPbFQ1FYvh4LqzLJmQwv64hzQ5O0+OoVcKs2OjtY7QE9BrvWNlYJCfpaYDBfYFCfhCyHTr5om/0/
H1XmUsS8CsXjxVb87hBpCm5lovYSMNfOBQ2v6ZVWxw2vgMb8wU0eJbhMknQFXWhSBf8+kMxSwkFM
QD+BXG/5Z9I1sC7NySA6J9x+z4e1AKcX6boQJNlWBCwiqjs0IAoIzYlDx0sSkZSVYkqEFlorQBHT
Igwriup+/GMlMRb4EG8DmP3ISz4wMlukZBG4HvNDaAek16oMI79Cnu5HYepAAmQnfADlfbO6OEIz
xlWJTwQxBvUF6p4Xd5smMATU7zyvDbqkYi7xxehtwQozw8BFqvjCM06YNYrPVXjsRz+V5b0cPOr3
OuRs3UjsU8kbFp3Rj2Z5wenId3FaKNqDGAzcfoogvRHFzugUKxKb8KND9/zND/xFfqKVhTuM710a
FjEgu/3u5mCOjWE/KmrbAcbblbUnL1k0BsurWGMGYQMEnEGXTBJiTuENUJp63g+Dx/EFFhqUM66+
OVKck+9hD8XmmrzV8+svFGcEY1CWdKAACz30FvwO+aykacySh43sJSbF6C+B8Guo9Ur2w4XjgEKJ
v8cT/aGpwWVgqDGw0KOrI4xZ6Svrw54UsIQCZUaFbW7STAJawERMQ78dehdzph6ll83H2m9ybcvF
AFknw8JPv7bdxngzGh7UZg4+9+oBxSuznIVIcseVVyftVcg9LDT8xeo6v7L4f5mZCCDyKLbf4Qp6
GpzBB1lxCcj2AY9Kdd/Xpn8yG74DQNUYLfWrtsQXRnE9Y7dF2y922H6lbvztNcx///N8yDpBFLHp
AtSPjxFF+Tbm+FxdbuZis9p8SBTyQCD0U0ABzfGaMLWkzmrX1yIETDkRHYSUCfA6gPBUZ04E77eo
hPuQc9j6xJ2km/B8kDnRjE8y4Q6aJVrmKcMtfpOGwIEEGRQG8D1WquXLvhL+GTwU1a1m0uPR1Npj
2qTa+qo7v15u312wVQ7MpK0BVaxjfeg2m/1kNLuUG1HwiPCMz50aB4xYxOIYvezjT8c5oqIS96I6
87+Jsx+3aXCMJ1Lo+TEquuxaE62hw3cG/7X3QQBCjC6cXuIBwgU8BiEMQkrh3q6CxdO0aUEMSFRB
NnoC+V7pG6Qj8ol5FG7gf+PPBmtlsDvP6lCVnmFCdO1UQ2ZWOEP/ZQB2bBOkq8WajPlHFoCpwW/i
ZJWyxQh78JAJZJNyjug2Q+bbe8yec2xRl0U/Bql6m0MtSNaUS92/iRuPsC3HRKx5OgMHA8foQ1sp
QGMMTmNjlEwhcDYM72GBTE745tTII5RTvuFzlnkg41MOlwPa6bqx55E7FjA95CEGbGjnBIhGcnYy
k6lCs0dm+sLd95OfeA7mzW3swcL/m/TZHlY3dBd8hCecPLvwi/slgS/xVW0So3xH6q/1HFUmc82i
MxBdAl1+WaG/kQ8Hi0X0jG5oYkAYIqUFVqVqkXY1dVdau9Ar8gfQmaxDhOAYZ7Np4g2V2elLwBrL
OazO6KqJOBfn8CSclEx2Vgc5Avqh1pzmjFNESH1hG/I80emTLgtKw5u+zn7K1LxaAsBE5Jq7ljvF
eys0HQ7duAiUZ1FxQvhLxnTfwiHUQziDSMf8BKn5QENTiOZ7Ehqumme0ribO0MsRhyPFzCudFIj7
NGWzPYs6vTJirSioRbbFJhv5JUJ94OQbJx2HDoxqGbHL/I2MauTS5byuaat4MTsehSl7DZL3zApe
vFbTqUt8X26K4vDXem2pDmpkfnvP5xmGZCMs/3xImi/FTgkOdlMhx0VIhmjyRaTy2H1ywnjZ34pE
unqQ5k7CVEdibba9y5vnm5sbfgKgITY07gAlId6K+pXvEFHiydXDq7qjB7EXHUCQdFpWeyZcNwIM
r05H43o+x41ajYBoB/Q0K1q3/NYm+D9Iow1kbv/jVcn14aupD0PALMTyRTV7W+MC8Fx+sa8xor+W
744IWczMHdXuIGvyWmNnEH0PgXZ/aOk46Y2DaYQN0tl4Xs36K+IVVjM25FYIjK5wv4SsiJDeyaFt
7eLjEDT076gzt5FxsUAGFgaGbxy262UsBq4J+HUIEUUKr6q9JQXxa4BfoJt7uakoI0qob24+P15z
Ah3EBwXE9nvDTjyXizPmlIuqwkzp4FjCtvpx8XbneVt5Hk1BZU+AJecPg/D+Ei/FxzsLlgPdyRk3
tsTQ8T8eSdpn4RqdvZb7rLjdVlUp4OvQqyzhVCGhGKt+gP3K5dePHaFZDjTGnCTsU7Mif2rG6Q14
UmKf0CJTfAHwBbgg3N7b2Vqqyqg2aIQXflIuaXwcXo9vKEsuvimgItkM1NeHkwV984OJO9j5EGzX
Go379FV9EYqrXX5If6AzJN3kx62Q+IhyC1afzPqtbh/wH3iXj5x7eZkaB7686AX9yLsM57BXnLUP
eyQ5T4Dz5S8YQvSXriKaX4nkWrh4WNgWt/YKRNKzYnPuo+PqFShbUB6QK58cIRDCFJwO8GeEQWn1
JQA3qpO/nSIqhCXJuwOxuHf9SSthzwGVaN8apMbos5Jh+SgRzY1mj6J893rGaokntBpS8ovz5A+H
vUV74fspHz0zWJw7bD5y7KVg9EBxaA6YR9rNQTAA9sBgNuXj5dv06lsKbrZdYsMoepN1N1r32SRW
Dt2nStvHe3gHR7xh0b3PffJqH6tNgcY+hdg2yg762iUmgTapA/KrmC4iGD5+OawsfU5QaFwwdIQ9
1UM09QzYIrGrtizbm4gHiojBG3wH+2bKX8ZACASonTaL2FXjfKMtnkPKjy2UtT9QBZVpMhYGdQ4L
8dZ2L8xc2ot/MCyavvWPzfL6atxrE3d6jt6sQRKIMJcEJ9t6SrtwsR1Rhbm9sPa50xg/oLpuguAQ
dGTiekDca61jFUsxmO1IHDKf9oTI4xlsaZMig2Rr56YlZdV3GMH1Db7vcddQw9rz2qS+Cu+ZsBj6
qiR5vGaG5ctvHNaZ03dsJr3at1oMAmfT07KgyCR/AuPqe4QM1H6TS1kCqm2CE+woATxfPphv2nkl
8EOdJFluq+yAdldNtWEZVpD5cYLN4XdCVVcR7QARhtHXtHZRv9Yv8MIo0Jp+jcWO6sDVHZlZ4Ohh
w5gU53e570bizg+rdhLv5l0dILmcmdmNjwo0GWfCfteVVprpE6eO/SAVEBh1dqvi8gOKXcNK6Qgi
tvJiHaWWjBhe/fQfxTYObzg0JJJPwmnjBRb0TGQyxljFxdXSInYCaWi5HMWc0dZDyJ16nyEy71Yv
u3oMYVbxzSktGnBG6Z1VCN+cliwaIZTriwOF4JE4Ffl9t6IQAx9nBoToG1qsO5Khzt/tELyDZHAi
kd16QjSApMZvcV7Zg8BjHy4F7zEYSRgVpS0E/DAmOHxxi3QmkM9u0xdDYxLPt3GjAlc6kvDUH/iN
Xl5iwEwLvoL3FZf5bsK2+zQhygSTd2Rfb6RzKfuf2fVA4I6sb6QPx+r4iQ5+tZV3VLAlHQS6sh0l
WXf879EOwf/hYeA5g11m0KxALofSDb/O/jfLp5CTgU16KAIRgy2+LRz2AT4T7a5vFGzMIlHyY2nR
PuZUOLS4bjjxwYG900+D9dTMZDGlh53rRYWEedF1Ss2c3gBHnYyHF/V8C3YqiIQAcrIArTkP/3Kz
JncVvE2EnLHF/qSnsdLqa8nl3TLMt2nTvfrGv47dxtOSxNOWI/SAu3eMKHyApTtfa6bbmykll5ND
UsslqthvjbIu8/f/lNQmkRePXv7MVHr20KR1igzPApu34vGTAGsPWcbQuA6JiUpuAEptTZr2dMdh
gFJpHUUdBQkJEG7zBe+FAyFZFIE/j+YHXi5Xg2wGTjmX3bKae5gskUvGJoM0y7tQa1zlcvB3XyG0
AIYPMDLYjYyA84wWxAwiQzIWWR/P3WiDn2MsaJUQP5lL+N8tREplZRgOLkgS4lOgp4Z26mIOAK2B
n5OxhzVjheHJmrMEC0o8igMjs3hqOPPMTnhGUVG6N/x0OYHJo0lGJWuZXiceFmwosZU/x5Wwt9Ae
8GQM7W2p1iUhO4xxL1G5E//Pa4ApP4LxTnRB6bFNemmukVOAfcMlCOzorRnDA6Mc9EczfGxlPBgV
nhmhqhEItxHjiJzoWk39yaGfLCXgPe1FsiNegf2p2tg52zCFHhNmcG0PUi81fFjgb3I3Fqr+uSY9
YT0/rJwWBlxTF9Me85xU9ruxTJDXnyYIGK33YFnQwwH6bMpU0RpwwnDrgfI1LjMLMsITumE6hrvU
qm6iWo/ghx++gcGuxfRgrrmiAyKuYmX4VzMdYbvvCE26f+vd1UYDt1IvCdpHE6NRIDPZe6aIDruC
zaSFJblvcyuWBg/cEDD8KVwJuaUv6A/h1ZapacNjdBjiN/1HEp5n43BsRB3bdIem9DoJ1UDFf34M
OjTGDLuohsG1S8rwFHKBJokMFllN83C+q7vGvXQaGkzf9VOTIRx6lEjbhFrQjLNgIqTfuvKqe6Po
GlqRSTX22yC1nGyPE4FXXVEpXddLy4Le3Ndp2EYzTHnoOIBUeS7MBw6Hcd4IStIsfQ7x0vdFcYm8
4DfBuE3iwWIHOB+I30MGEGCK9KNprsckjmExa3lR/2Bez6BNnA5KgXqzDfm1V8scz92oUFA3+gpe
GOWdmCy7uyli8F+LdWIZmfoKXO0C/hAxFD7gaHU45QeNgmw2NV1v7VouB92PvNII83ZSYauiRZrt
e1/5m+kkTHQv9aZh7IEKqWrpxWpABEqFQATE4U8jAR0OBkUnukremmyyUoyCrJSWz/GMjRIfgiX3
vlFCnD+l3vmXUObN4YX9kHJTvyPIe+JAsPEbWsrMijSfkvZAuUGwZNWC9M/HQ76kQlq9BEUq7YZq
R3GY/3e9/KW62pCAtlRbje6uh6Ga7uBwqiiYFJF8OKl942zfrhl6ZYcpzhbT8wlBgu9Vuq0b96oe
126KEbDlLOQxehGP0zUB0Mf1lZfofQynJJpjMNUQ/c5SFhTWPxRXjdSYGPSi6dkM9G/3sZHTDv5A
rQ6NBbMoZBQMiGDOK2U2KxaIHhSqxhz08jy0H51YtEYidmoQJxCXlHEJp40irRbp7HpqBsKEIB6F
g4CCuf+eIKlP/ud8+qg3z8hSIOTCsTxdjibmYa29EuIiv1JQc4wZqYPSRm8wqcbH4A+gSjoAZq0D
BNJmQiUr6llvjiC8U9xrqFPRYcytKXk89QebNFa2BKHj9qepMd/utIi7zPYYkT9VLEhVQtKEvP+c
YJT/0mQQrOmGQCVxuPCsFPO7S3qeMhYm+/hoLaO825pQuhXUzwXD5+cMWsy1+e8k3YuFdI1K10A2
AWhqDdqhnvZCdXMLXhxgysgSK6p3lTM626eciVRDd98rZ5ijHvT46UaZ9JvzRRzwL0UJnspUPR2+
l3jEk+g9Y9b9+X0JoXQa3+YM6KUZaaUOQpM0itejQ1meuRehc27bZosTwXAIG2GwjSR530Q4oLh5
OLcJcQ+f7uaAS7LaOnxAUi7UNvDrojaABIzRy+HxiX+zwaxAE+Vg/mOZ0+p/eVpF3KkPeYXmDvCI
t8xPSNEVy0YhDG+iU4dW5JGceNNmvtXcBmHfME+q3KaZHvpvAIxiCbpFZZS2cuU+VIds5l30h0uW
/yIrglDWXhB6YVR0dx2nlYThPDYtfOi3Yg8j7XFbieOfZG5YJoxHxIn/mmrYcYnLT3DIcAeisjMS
qBl5P9BHyxTaZwNSDhQG33Fh5AmmYc2f0/+/ZufKHCyWLkBLvad5wY87TiDB2Wa8MaNbV2385hjM
Mx9Le+9i32FaLsMnF1QnA71AoX0EDxdFd67Gk5v82BBpqQ71DpiW7F3d+LdlNNk0TAZgTF0HhUIw
Y9YCQRd0kupZf34Fo6akklcxSDHJvVB/xypmrknNBMFPdnhizQta6BllXYF8My/nyr6+fmxR2FVy
CU67gLYEDv7/7ww/bbOi8H0KKxMa+bfvoz+h0Ni1EyYFjsY2P/TcchkggzpcVw1wUAh9usU5mpys
oTFr3/cHB9VDQmyIrtIUqrI3T8db7MrYJbfhRYgt0zf7tvnr4CtAdaYOJwcXvxuhj+UqDUl/cLv8
qij42KXfY2l8tti3XvHgSN745xOL+Elz3sdDaOWWcvY/hFdQEV05VZ99zlC0azSnAhJ+VBD6y78X
OLtxmyBNeyatKe9ZhoXH33PE30IxFyODbYZH1ecJcwqogh81Fj5kLx9Ls/mw1FoxfedGWL8bND8s
k25m7duBjJu0ZwUywgPl8yBjbsDp/Q0RToh2iDZtukpRId+viSWNHmNo0790SsE9MGRpoyIDsqVC
pZ6xjW+wZygPIWkC7j6WlvON2TuTX95cTB6enHU3bNuckhdBgAvfxTKXDIOZNhi7IcnbbhnMWn20
spfZ8MBWSNxVH6A+vkF7QKSeKj781/4KPvzwHCyz2IUXmEhF+bhjUbNx2OYM3FsF3Rl3ClUtjm0I
fGwFn3odxymLO6PPydc3cXwHzWsqa6ZdCRJoHNyrMfFyrtajGaxRs654WKZJEHJSrtJ7Kiq81QQ6
O4aksaNFl2GfbpwaWXYo7In+KUhWB7W2yCR4zS9Gc91/z/XvDr6vWRVXRoMMCdXXY5WoHNgf5Od3
KzWfEWepC1U3oUwHEPdWlTMIkx4aHQxr9IM0hVBxGFMZHTktihODYwywYby+nfw+rgLsYe4DdEpO
lpJ3JhEQFrP9iquv9ICRXRPB1W4E8C0d6FGdKUjESfZhj4TrugMTTrFCBsgYh4oaRm/HCXX7Vj4T
WD5AC42aE2YBHTeRxSdM6mn/qFshHwq4dnj0qHGcYCSxDH4xzzkF04A53+WVEL4O9tYMP9PiBAy5
/Qm7dSTeWisnjjgSnkLiCAovVEml3HOXRLFaWyBoASKxu9FcIZXQnj9Bx3AiacfZltVwtm551jEg
ljqr/b6NflVKzwvAA9Onp9Gvp0+L0ZJFIW9PVfW8bMYjubvUJn8AQ6nwT/KujhFNoDIgJi7p1DcG
fCksFoTIg22PBgDE3OOVHUfIK4wf8lqCv/wAiLDdqNihZ/XamVlmcpDpZif2LToTcA43zY6Fjgph
GOY3Z+5rDkh3HLibtv/7yiwtP6Bl/IhHLAPO7X+3eAKSfkxsAI8QZ+TyYqWIuo0Z+hInHhjP/NFj
ykqI919kCpAo9JVY4AqUoCwSs96uI9Zb4/KLbWX8QVqYNgQNHSEuFrtTe1C5ISlFf50BCC1PcacW
xFSr24hAEMCG4mnYjtS6l4aS9Y1LcJZFV3277OZr+efY6z4Loy/2/cnFgbqmwimCTIPaNe2F0QMc
aIq6OB6TSRNr5qNfs0yqfWxsT8sbATovRHMO1nncLaMFzASkK+V2zVQ7tTo+2W4t+n+hnxhPv+sO
oFZsD1CJoNpxPOFpsnxfSNtkbIrOmFXnHCaEm8+COLsR6lvs5BTfXgkS8eA5o9mtoUnVlfzgptY+
eOlOx10w83HBrTGqZ4x2mpizzTWEDVGI0cicSm+YpBHKArPibYvMvAhw/xUWr+sXKwoV5ZYqOXYf
Gs1dTEral7jIH/ICTGQHv+7qWHzLyl71UNZBZ7P+zVCkVK3fcD+IC0Dmzl7OCrH7hQ/V0wlxG3Xo
l5oYTuPo9E6bA+0Ual/XFTnsA5QirXs9tUZPIMDHnlM9twh72bG1syIyNgm5Cgk64JIHhu7VZ30E
lhc4f5rHhLfG4ATqI1uUE1Kj2htH5AcccNjDRxYjTMv/8dSo7980d/Jevfq7vjI4/su9HDAer+Aj
ZvQl94qDugaz1RK9s1eb4avgU7mcayIC4gsGCG2lU3pjw8zPSqh3RrjEu4uMNHK9iIEbBqLbqFu1
B+NfuwgVRKlueMvHTklQihime6yLrWVoAWGJ7ufSoB4Rs6U85DRqNUFjlFU89BAIuETZBdArDEEM
OSYDCZT41VWdoJE7IcKL27ZVA9emFJL667CVJ2H3OXu4P2FlYNJkBMWr2YdFaaddQdA/I0ncNvAX
/QwI0jLKSRHWUkM1w1QsMn78ORhe2oDICcNl4H9OTixxEHlJzh6qPWEUrDzMw0Rm/i86f23179y8
+hillx98bflwtjoLoxFIX5o8wVSNUjUpf7DSzWnWJj71TV76uggnPftDiFF+/SOpDZdiuddZ6nTt
Zi0UkhIpALHq/UQO8JSUjsJF9wGqiM6PabVZ2OfGCRPjS4VLDgx01DgFgIgUzpYES+KLsn9T/w7f
xbTUjWlf+08j5R855risN0Apwfmah5VucfbxUYiR9dHqBse6xLd1JXG8x7EQuDmPaNL1GVV6Xn9N
QEn6oDWE8dkdKI2VSGd5+YwhIUOv591Mh/a+6aGeT7KYEv+Nq+pB+NzWIK0+EV4zc3T88KykQn5j
yglF9ww3Ly+An8WhEpJ85KYXB70UD/Smo4aBPw32kuS2X8KyqNqDpEJRuLfYS6wddqh3aI44t8Y9
ZCcQzWnNO11O5FhmQv5Yd5BG2LHGR8zw68jxjORgdlyhM4kv+GPU8l5IaittkLnn38njRTYrIUuG
Jkq+qhqDzPpeAZCEafdOsMv9DzkBx5+UQ1pDx4ySVsQHmfswkTc4nk4XdDYFNIVQt8MZyj8PeJvc
8sng1pME6IXgEYjUNK0u7qFtu1E+jnUeAVjdDK4nmnCCWXCkwLSRmoQYt5EiZhqxg76gdvpCkuax
X1T6GW224T7NG2vTK+VXi23G53tJF0+Tny7RQ0/OcKL4zvIVWZj0TwbN5PNudNJ1PSWDn8fXgx6i
QT93JnvD+gAi052HaVhT2Ms5O0aVbl1HsiyET+3UFvzpnPaPq0ZqlF/T6x3v5ibC++K5WHfTVmi5
LjqcVN5ElDTJhlvGwAN2aKPrVOj+ZnM8IPCwZCTncrdNakoxD7gByZ1eBdUMQ+3Sb9IA3i3xiEWp
Bxw1L3O1Y60hHNncwSXR7pWiQggd2wWAkRMk7rg0OehZ0PjW/OzYFv5CwA4/JhX1lUy+0Yo60Suz
3Ji3hCu9VFL1+mDBRRZf2MBGpMRGdrXDjR9BPm99iaN+7H/bPq1rox7wn64JDe1rPsxM30PtVOJm
CO2Efbhb5krpVUqnKpEcPV5Sah9VEYVKfNoPm9LRGNwSYn36PwY8eOv33TQb6QgCHxoo7SClmBZL
NFfrlNy+FhlmnDHEWtqorB7x/rou/+OlUbKDcR3rJVThOMxjpPIVUEUA6sAwIHpFg/c42E/HDa7s
HvMC/AwwmJfZ9+APf1rjeT53oaB2BvPQ2pKbebPW31JNhRK8ZrHFQd0oqC/QNGJcQuqnTHwBgqkx
1P1SskAqSXOAlJP8hLNw9EaeZeML+ITWKJdnDapubojfGuf1GhZWYwdEbvki9mzlRVmxiJtoYvyi
RYHev9cq4XuuYcODlap9pj/58tW32Pfg1mRvtK+1i3tLdrDeQku6SMHB3gv2MjO4rgl65hbGrTNx
Wj7qoX9uCriLz26CQc+Cibbs51EE13hDrrfDAELvvRUVeqCf4CDOvJCUpi3HG1oSbIiHhkGfOvmO
MVEMvFOSfT1/zzDCIVu9PdKaZ2nELdMaWbKsfRPT1uvv/CRi8dFWo94SIVWwKdMW/f8w+w6LzrD+
geL5BhxZ7MP4j+clGkqa4HaUYFiBpq640jZX1QvLpWGdiLNajgNMpHJOPPYxqR2UMu629rKro1uf
BZizfWqw01QTTsmbU0FobpmwTHEyFlRUqR1/l1VHs9sipBxqlYehs3Xj1CxLtDEWNlPRdjXbVfig
2GchJrahzerv179Dfgct4m4wuyz6QNpeB/Sua5uFAz81GYSMhgbYiC+dppv+g1JpJjn/1b3iFKPS
JHe+fJCSLc7+3dbd5/vVC1pfcXPqGgQtzJNdwcTsCmGs2PNSJIxUuzup9960xfdWhvXz1Eeii+nd
WQBRkc85PnfAxljotrbrVwgq/Ekp1WgF6zRamCGKglrGJ5MH33/pKKXG8sCoRnemtw3ogfXRygxR
MwynjXUpaq4OqHqzLMyFO3oCvOL19eGc+aF6gykuglpR3XWgJ8G2scBvQPJ1zyyDKZTXdVV7KGZr
tFHkNhPDLuk3lEnb2CVoLSLfoawxpYnHjgaP9P0cs4DJje6em586z5z/aSJxG8TCpXqUSaM2JcR3
HwvShrJu94myoXsIrKhBLCgDK8USIOg1rzG2S/Pcio+1ltcTj9f0rcUU7meN3oOExxmM0XbEJuH7
DyQztzjTBHeONRnU6NoQhSYAjxFsZgyrOavs2W4j4JEs2UxSFWWNYQDU+k1VWwN25PJarLpnE7T7
98cJk4gfa3e0xT3rxriKI0gig13wxLc+JeJ4GQpQBTIiCqgl7cMc6ZehGP0qVamiwHyn4W53DDAp
X1td5ddljD46onjHMkUqXzPl/KoD7wGjhTm7LKA66AJsuRBGTlj59fGhlPt0qoWZGrOhNrJHRhey
H7Kd8DRhzx2bEDZV2VnNKjNevROt3nTD3+TiTwPQA3pWNam6qPVYgbiMI15YT8G+puI1vZYM5uFi
KDohF4IhggvKcks0XXNcoWwsRIIRhXFFQq1+rHmmGoSC4byzdewM9R2cvu3yWZo+IKw24B9W8PmI
PpK5jraeiGg18HI820J50NvHNJYJ2TUZjFL4JrYuDgT0OAeHtldV6GSjvQUB0NS0CBwtWMnHrlxJ
OTsRV6Y+uYCWzJvfDYDiouoK9VltpMzhvSBTgiCe8DRmlX62xbyakpUaF7b4mebwx2WQRG5Sddgr
GAMBrTPbgUj6GeQRS48bWaT2Cv1GYW8rG6Nu7rUJvib8ikCSK+G8Uw0OrWkSAoHKep0jFJr4zBNe
YPoGAPIixqrwl6s+ofr0XubfSAPuitURkddJj8R8x4Tp1ZLZ/JfZl4maf14NlozXWy4d5xr61iVb
CGPi4JT39863LXo5wxzUb08NYPsQyEU0mnNnaDC6eXFhIXB0LQlsMkQl8ujfjSbrQNOOGdw0hFvI
SWSwjicl3CtLU9jCfEHLQanSsQw5bLJkH0Sv503dXJjyiUPowyhps8ifjoJ4tS6GN2LTjNMRPMnW
6rBNEk0ixJUIZ+ZMUpismpFzk+1KfrhXD0+9HZ4joHOdt3vLjc9TpQ2nryfyL/u5jm3I5ImXdaRk
tA2PFPNLcpbGjtqqYCFc+dHoMrkEABAxBkuq/9kQ53MqOccBTlSgqZG+Ux27xEFHOEvNjrF3aIWd
xe8z/zEeTkSxj8VG8feCJstuX8ToJ9IXwrM8hbdp8GRKEUt2DLkVLK8vjgzYNNCl2fMObtrfFyT7
6NEdC4yr/sRFMdxXv0E9+0HT6rrG7eMrldvRPi6oHisYz4EQiuiOMuccLiN/MSrHiRtZDr8Iqiw/
5U+q1//3uFK7KL13G4wmDJa+2CqsIK79PM5kNau0EIDCWqrSELwP3PPU5adHvL/33w/Zq7l614E7
Kie/zG4Ktgr950Y7yqvpZCNpbD36mpV057GInDkaWgGenVDz7DoPlz6TgtelQQ2hsETv4IOWcWlj
MpHBzZrGYGvVq9gR0cbFLELBDRGx0x1O22YRHTMdHCILlLjE9To15rIbFx7dL+6/5p7kb4pp/VVr
vy9iS3LbGrhFoVDuxnLSd+3fxzJqTBdaQ06Xm/55Ggu808o4Bm8VWtmFyBuEgaXRTaAUdo2CRdFG
pyMgplOAK1c3+g1ibOiLrUj229vIEgKH2wanPLWakK50MsUApG1wivKfeeSpqycIADo7qnDeKqS9
onf5D8JJZPT/XZBB2KUNadqkgQQ6838WqUhPdyedu4BSx8/6tudfq+wZINGCxAosbUtX5MjkaUj0
L7QXlQyumh5v64P2BBLIXJ6Ji0OxAyIr2wJT9gpeQ9+qwGnHZ0Jnb9qzRoaRwwXONn5/JjD88QU8
J0GKDOF++td0Z33oGHPDajOkp0NbmWdDMjhGr5dGXzLNMAzMJPQVsLgbrUdR8MIm69jeW00TYIRw
/5JlFPQDvWHGwDtEJFnPBfEeVdGYpTbwzxgkK+YDh5lhWWPwQuLXdv24RMhudYVK8bTMTnuLiPqn
A7av9/AvD8i1wT30GRuNLuinWLXH/zlUG0b/prIpnn9pVH70/+E+YTK4aLznYeFfeFqxUjw02jvS
Y99ol7WGj/M3nzVIRV9zm7TEKUIiIBLm5gUPKOhEq1JMk9k4Dg+FiPjpaZKp1UtNBwys5rzSDUx+
Vidl7EAxbj6oDByt57r7C1z231bcqgG3gu0oAYDEr4FACz6qKOSrqztBDFeCtLqV79G1+nYhykhN
WTH/nB0hetu6j3vVMj/vzRvxCzWJwbfu+PjlFvdMUk7IXVaKg46v1C2brp+hkzViv3QkPfZ41yAZ
DmVR13XgSqWy8HsNytZ1w+3WlXjZZjGj8xmpQpI72X9SaG53qZ03hH9R7u90y0crvr/OQG8M4JNE
IPojXE12Z7wknYej2Lq2Rteoh5ZeJ43e0eTuNUk9EPS0ONb6M8U2sLwbgdUns52O1gUjfnf6CNEv
JLDNg1Veh1YbhJRx1Oi/00aD5QMnG/SCtOjcF0ZaLT6IZO2l0INHQ+WreIHW8nCGJZ05f0HZpDNX
VeIglU/TQCFDaWd9Nvcr+5tL4M92AQa0UdMIj/OCgdXyxL8i8u2CtU5EqtJacfh6auiigEPuyAid
6ZRMXjExzfwtpryxbq5BUMlIRoSWz9ouREsfGQU6SwsKUAjPiNwEW6/CMUcLLKacfKIa8r2WsNF6
RiMt3PtmiejHP4Xt5/sShT1xXLUfv0+Sbfp2aRMLZKcdpwFEwAmS7BwXXF+RqWKe2FWCTWE6frym
D2+Rop9ikwBzASXINefGK4cFOczen+cCQrpBrVBN5/fzt8ip+/B45ZnOSlMBXKVywmP+xmTIuEWw
zvCX82+5ZN162/sI2DYeOCeuVKjzh5cfLWiiXOSUZoLLjE3OJSzbpCAmhM2rIWUHFhnkalY+0xXn
YqXcrGmGvWATiEzeRTh7JIjqsEk8xUYM7mXV9zqogho2yympqvq9EfYTzvk1eqlUWuRdxXdaFtz2
8YuJ1QdECkRCa42Lu3ViO9gOLzsK31T6sS3W1V7EA/P1eQUq5P3bOWQeEj9g7uF9mEq6LBArGhJR
6KRrWBstR+W9dYpVCfWEx9OIggSRX8p227W9u/GEv4AKc8NNjXeRAIn/UFAx48RnBBvGef389DVn
oHhRG1dX1iWh6tqz8PQh5T0FVnnw+lJqW9rlm6DLCilJrf4x4b1o0gR0BQXV8Z95dXzQ3cGtg+Zw
5v8BoRu5bQR/K9OFhSYDDqdYl6SWO90dQGZ/TM77QVDhLLwcOci2suE5j7S53Z7hFPGhPwvFZESK
y2hPHItmH76ZXt3zjgUaewfmmhSanomFGrzsoAU8so3QueKmFzJ1IF+Erq4ezkiQhSd4g7KIbnWw
W6+lUMpwuROCoPIqGccFgZu1MSsauIcXNXWEogGXwoWt9GCpSmrcXA3wPa2+3W2Q7u3DUoa1k3Ku
EjIlecXnD4npYyTGk58gP0FeIKr5yGl8flX77brhpYUnqZSgqAtW+u289zGTGdVlVWjboU3rL7+H
qjjA9hIlymTPWS0bO395wN6647T5ToYfnfg2I+q7DQEqnkBXYretluA9PYNFAFZFX9bo1JRGvCH7
3C7SVMkG4EJ33jh3qc1isL71sC9EmAIOO8C6tkMLamQtZpMiGdnhwWJqJ41SwLJH0Zc0Q0CoFRVJ
fAtftRdVr8nXTrVLj63U2YF39iWfw8i53eWA/3jeicbJyOFClc8YsuCO52NpqrLqloa/SpYqRaw5
DscxuGV7bkPIULOsJF2fuXiDtdt7HIj9g9yljfy5rpmllI+OUw9B8H1mh2tPkxEkE053SCWRbRK3
OCP6XwxqwyKZ6k0XNbzNrUrhETOGZjV5TdWXnVHxybSukjUyvQ9lqMOc7gimYiYAsKzdRib9xGug
vGBMPS2xBYWXNbadt++6rMVTj2Ho07zINmS4flC4ScFz5zooNCM42ulQglh/yrfn9GKuFNsTXBgP
7YSz0io3AUpwZpiSW9o2c8RpVlqkL+3kTYWIedKbab2k2RfAZZNmnY+Aumhd3BwUi2MEDeOWnIQP
lzaDyfEFCtdjuzswKe1VG0uvaVrIJUw+ZuBD0HRW7oxonfsUnx5I9j2Tgysh6Pw2ypPk3vBKPuMy
aEh55K7YQPzI8QEMFpj5n1+v8NaePRgT0qc8LJc4Jp835bZfJZ2XtdniPFggWTaYvO7SP6PxuL3o
klkk2h/2so4M/djp2He4TY8V47bV+uzyNREAyblY/W16E7eMA9mIgGaC3pPqR4/1to4ENb+Kyxdf
j+ZTQdS4MbQkUIu9Ju8KNMe4DGSLGLXu5gwasr5Ok3hkcYvoRCrNvmHWFCmokUB+ovxFDZ4iQI8+
5c4ay2AuyjmiOAlFGT1boVokpU/8CP+PadHGjhvBKcd0j3Sn1W3+IqNQ5sRqAjoL8yQqt75tkbem
pJXl/GK07YQ+oEQkfeom64jS+EfWIJJ1Tozc7V9EO8V8RJu2mQmgeh1+QtfSJ8Fpd0XyLc/IvG9j
iKInv19ZenlnkN/HmInOorDTpAriTpnzNIMhR142RSuPu93DZoUhd/lid4aNuRO8BqX37pIxEVdU
Est6rmnbHqNUlPDHkingR5+Gze/o8dOGvHCUqEbEr38rIyOyrpNEramePsTrEWVrkdhOvrGn8Nrh
kABN2MgttwFfuZKQpIiF64ufSEV96+0syhirIOio4wA0rQE2D5/pg3kAp3A7Jh+eNVA+sEAHr5bf
y9jyxa3A1NW3o3tA/4OOgG22/yfBFKSBFZMMouN/ukoVcgOPidERUynj931nY8ED+7EtJSIbAB8r
51TvN9vwk1DNbaKiW7oAZOQKATb9Nn+59X7EOOWoE0ZuD9RwaYlqXaKXa20FA7q8lXvaD8FFFfC7
Xs03mFf8Rvp5L9as75A9u+vdFmVN6+WoTr3cIFHIyq1kiecuqy1G/kw2xx3mFFSz3Foix9Yic2x3
CEkGMhHsgjbTV6sWYqUNBndty8rLLRrQOIDItcD2nNRK0lXAJ83xy6lbZFf0KGpmcxw0sUdul1l4
lkUt0o13kmHeOP1W23hsTbhX7BaIqXUGUIUOy7Y0irwsL+7IV/qxRTKPSMkm/0M0YRXPQb/m7O48
bVhJTEmRqaNRg7EH7hW8S3hsONI91Vg3loAOz/IMqUwdXpRClmYttMeI5gNLOKibgbY3gEgGgF16
UtRNVWhMoESPYTnpA3vinhdqZ1ruNGC3ZhXLAwEgw/1aErMaVEJQL/S0VEk7spNPWVhWkBEQtCrr
r0jU+6zAPs0SxvGj2vhjoY4sUDRaaAxApBWVcvDZ7AohPE+JCrFwqHLY948eIUEfYnJPHXC7t8C+
ShEeAnzxwCLWIoGMTRbDa4CLtfzf5N9n43yZt4By7nehljS7751Tp31EQizZ2KCc9MLvDjbSttyX
9PHwh9gfTO0tXjZl2WeegARUGUrXasRootMmNekVmO5+FTY6iF2addwPYQJWu4OHshzqpbwXFG5C
+YMuIkvUqn+aTYAeKug5LsW33odqyLU/vFozTdyB6C9T3Np7AaTJ92/W6sThdzxalnhu6IS6Zuk5
L/YaHBZLD59BjAHITJiFf6Ed2JQIASBuY35R3vNKXBKq72GM4LRj2fLB0UawdIui4XjOPcs8JTab
sseY/agceTkIKXdUe7f/7MAfqV+1ojdhaW9juqEllTibmf6ijHNy1N4ZJA3DaBx7q0+brctJqRb/
8HRb1sgUp750cT5j2xDL5M1zNb/3naIWdfciz4d4RXNhl0vxXlh1nvmyk2PIsfaKLgnHD2xCyic9
dBZKeCeYJqjsUt3/J5BEwSePWOhddnrya/gZmVyTjSK5+DiCpVjDd1QO3sfjWoURnkk8vfMN3vlh
JExeFmUKeHU0KVM7nAlvRyOtYocvvN8iYUvCJ+tr37LAouocHeFDv8AMEAaOpjg4fCLHcGSp1jll
sRfvVjimzMjroAtvDM2wOCeZlNQ+XaH9TBJcCr+1eXup6eTZezCDu38NjxGBEqjF7sS6Tr6KJqcP
gZPI34PB1RQg0lS1Of/aljvmJAwngFQCOM/ZgYmv7AdIfV4KjOIrzpPnKBGEyJmeXKiteaK2bavj
Qe0OQ/kcK07pyZJaEw9BJHrpypnEAA8iR9m1T18QZttgzSbajmlKBlPCqhzeTsqiPzZoK6RVAduB
YwoSQv4M5kk2rAmQ+reCgygRgu/EFomApxlad8+VKvfkeytVIS/rWU+UC0LqVysGYVrBTZBJfD3e
9aCH79i5JK2joIS4d6VFFRmW+L/6yX63zE72nWXGTzjGd/izTtE5AKk/Jr1M+tvlm28OThPmqb7L
LHx0FSB2c1WlZX/agRKLsKysbJhR4Msu0Q0y/bzLmVGPJBlQJ1bGJwW2ga1wtBtEIZG+eC3sQ+Ka
TfseykdLVj9mv3YR0q6MAqlZIvoDYYY2CCCnqQfrwiuiXRPPBH8AseJgqM8HiNYOAc5NUNSUzSYy
gwo+LytNMqP0ADqNL7hLuW3uWrBMcm12ewgn4jqi2egO2S4QYP+6xGc9FPkoC7l4hgTXCSiFpznX
UEiHx/L+aGI5aPLUQQAt80z6xOz0gKDgwq3Ug8gTyLk/dtINtAw1FL51ZTbaUtdJFGIjNdzzMvIJ
43LUL1mm2VBpO6CpzcKywn0hFnJ5T72Jwen+jgrqW4+UPVm28pcqzEsVDpibV4a2j3fr2jp3QOrC
Y62BZlTr187Xgt9XsydE4DMfFh9J6kwBgPjDb/P4Zr0COiZWVZZDQhUC7Y45HAam/re9KL25yFfs
mOhG1qbJaC2jDGxUbs8AQNDvP2atWVUhdwW90qJwwIFM/lFWO33erAWaJFFKGliejaPStKvSaD3c
p/xYPoazSn5Oi5nopSsv4s44QESisdSo3fa12xQmXLmdrw4zQ99pZF2g3vzgTzTCH9G5av3e0aNK
rckb8zMGP9t3ZDsFHjhPNoEq56evLaY2l8R2bRNwdhulLPto/ZvgwTbBfoM+x+/UEtdY0a8dbtCP
shS3LmWYiDpPFScXBo1C2s314+DqVWIqfgCHNaZGmLOGoxOnUxFayjNrVYYlOYc/3dQ+EU9FrF+0
LFmZ/mrLeKeewSfcBwrMdpq7DRug+XBQnrLBQjPscjJamd4E7NxnwVP4rum1/0LX+hp2IUq2H0HG
pjPaJrfTQXoeu9l81weM1+AZUfHEKqAnhl9wKd64ohgu8vXvfCGnbeLbVN2hcf+gDojSgDZOUrGF
EMffU64XuPmfo5fhe7gnQwMsyuonXlUD3JxP1trL58HjwjNpaaKbmi+TXDw5hYR/uCPC2iOhw0du
9cW5TFCY77NU6Cocuf8rR8IvoIsNc1RVZO2yuexHvaQamZ56lk6aa69x/OrHV7AlmSiYhEyCtlu0
cDIIsLhm7Z0rTIc7Rdl01b7R4UR6i0og5+X0PVUEecKuvnTgvhMCuPq0CI/MHiwdr3gLif4htQfZ
WjJbePBM50U6YvJsFvURVVz0pMiixW3XP9IuUDSzkxs0UIcVv/pfz/RmGUsmCmoclRTvlyDtXpI7
t/5uXrjE5MGx1WJGLSJ1Z6bF9wyoxYXIg0zm3AdAWaenV7SSDDGoPUSi++QCXEZOZtmDKdDf2q7J
KdpkzlxpXEZgR64r1+KWHUPhqN/CwkaS0JMFpD18aWeSNSiBvOFNIj73Ayr0+BIy5MU1nE3LilKQ
f/JKXBEVbvhTENDXvjvOPtVwZPTKGsnhCHa9PE1XYO2AMxxCj5mFkKR8bHiGX/uGGwrHNmN405K2
WlQKi4UPsiNguZ1xG/IWZ+xWRZX0mBc9EzrJ+re+sayUz6g2JgHt2KvgOEdn1szCD5YO47HTkjjX
tOr0gQkPhTfbcXytBDW7H2suu4PVy+BL5c+VsJ5aGdsIoMQGUHS7zv09CC0AgrZ8KU4QEoZwdklL
wuGEDUH+AKAhkMJJr+c+nL/U8o8Gs3y04soQwUPS0gsWaZ0cJDVL2hPfU3eu7JjJDHs2S+xS9lFI
noY2Bcc1qWLUYWhOJEHkEjlcDt8twdmgm/BIwQgEreLZV4saCNBPtfRwkYHHXMm4QDLVHdbrZBJh
HqwGlbVntoJ7iT50uHswxILNXN9oaQcMNQy4QsKFKe/n8HKx3e/bKCGAKnQPp4NahNJs9Y1uIdZ5
FIkK3O9lQJFDh1hyT4LDq6X8qfu1+REyO+i9k8rVV6Un5e94Alk/D0Ih6/iNyALK6E4LjD6fZGGM
fEBAMKso05JI9pwciFC8U/PsbYNPPF+JPuDNd1xgrpH1n01bcMi4OLnvnar9OcLilsEabImt8pKs
CX+XH7EHxXBXQt/GD5AhjG62i4UQpe1/E1yuW9OQMRxVCt8MoWHzD22LQMRa0EUC6tdvj8ivoxWJ
dg/66cAGmqQoVUjXc8aH3ADQfgRL+JGgnxb7qeplW/exFsd5yb+ZOw2cXsV0AEsWpb7soqCWEtrA
fENokgQ4gDpPWPQHHYkcpDyVyKBleuk5eOYm482248CdZbscrWLRi8ikjgnkZ4sQHG/Ske4dtHGf
D8ePz3GfJyx7cGmVqwV14Pks/2w6vaGxxltdefeqJWwD+Pw2uIgNgJJO3Y0THkkDmz0ViddR0Ht5
uJoRLhmFNRePCoEcpv7KYoG3TGDeYBfGbwyTXnizEt8icuqpuD8llkwCcDJxdcRGMufvsnPm9Blh
Z7tPQ6SA5AU6YEB06lPjNPRQe8EfC7HpO91bFSGh1hjVaMbH/LNj11evUQBwz+MxaqRGjnf5ERUN
snYC1DQ71DjqjZgLBvr8V2/UbTSDbefVV8rRczW2KsPW/0T4NVkgReLvYk4WuF006jEbuTqMfcMo
EvaJDM525xJeOhNLfVFdIUbPIhDFb0rPDgCaV8vuMjXksT8Ayh5GOAhtKFrgEjDhBcmfEwILRC9w
v9SB9aKPZcc/YxhlvV7dZpxj9hrp8HsX/VUK5bfCG0lwTzPuvpqvfFLlwBvm+c4TiTF6zlPo0phk
N0WJYPTqvXmh8tTGbLCRHe3TgwGuk32KiV8d7iO4sl3fFk35I2vqiHADE7Nvv+kwpRtxEWBPSSkv
nrwVyHhcjmPIsVrIJ+fUqI/k3eenNiWhsDQmh4AQWtmvwXL5ecaDsG5NtubRO0/csDUW0yVD5wLf
YkiTpcz8Ns0SNslW41ECX5+kb6UM+4ojr5bnBObNCfchvTiQsinAXQWh8br0BgGlSvzcsArGAbbQ
Wk3yCzfTwO/9iHUleruPBiAleVsWaWWdJ2DLemjOx/fSvw7NGSG0uNl6NpZDn/OUoJH6SMVIVxTz
H+LPkBRDMVLmtUD+uJxC6CB2uXDLo4w/eIeHYF/DfGkjvPAt+mqr90/EHei1ZREuN8QTerTPORZy
+RbMpSlbqtq5knJj2dOPdiab9K560fzM3rJ5f/5L1XChRllncvghylrYNAjPttOl4bJrXlQhuEff
0nufdG1FCR+RAF8c/IR+l920V5aC0Y/3zuFXvJEJWJCJcBBvoK/VGa/HIgsB5qJ82FS2lENacZYF
Z1Mra14e63MFyzVBgIdAafjb+QBFKWYZxmHjsSf3hpd8/DoK5yxaMcPuIbMHw2N8s8kXhc9ecvQi
G8i5sOIlGOYg3DsJOM7WhALld3CjS0X/ASXd07XrI2piXy+gREH7fx3idJZzh5YK5piQ5OkcgugP
8VdE8Cqwt4bXL2/KYGUolZt1fQlF+nV9vT++7KnWd402y9Rd0Mh7UgKt7T53efavBu7w0PCxylPE
fk6XC8AZ3lqM390rl9oz8/Q2R4xMA7HmsEwnftPLbQBReU7Q6kF27A0JbFm/ppIoGGDKRLG1vphK
F3EIoOYaj9paAFrcNphsiIoStU6v9UbHh/645CmwlKFXoxo4qQ6o9kP4ovv+EbsJBXvhwyx4/MrS
+xEXmAI0gclfUEDpCsEZs2x239SmrbCpyKHwrLjqq2jZhYGnEvhu+ggFXMy97GQdcCMPhStyUWsJ
27Z/aK21lA2luB0L+aE3cKn6skL3FTVvlaIOoGrXhoen5gvENrTDv9dVU+HlBY9WjizLh3wFGCJz
bM9kzgz6dFZKSizCibqCiBgRY9VZyoXZICKNKfuIO6IM/1MqwQXVWVFFmd9Hayk+18J9PqAW2dMa
flrWC31zz/IZvlPkHFJV8HByBlRbrCD6eTReB+5S+hg848tPysFhmHlnA2EVn035fJcjzKCldiVg
TpPnLSrrUP2sRX86ZhlikxQdI65NtcuPRBJCn1q31padwurLKIUxnFuJJuw+Brrzmu/7BZ6GUT4O
WcB17izo6jdA8iyY6qYFRkitxOhuaJ+fhbtkQJDg+M63n4zjF3XyIjofeiXvncfZy7kuAiyP24Md
c1l+IsEiW7i5s1DHPqpzB9PQeod/tz9nC2GJ2lF1C5JxP56qJswBW8hszzFxc9xurj1gFOQLaUyN
zJjKnmKfao3Eh4/NwMJtO8n2GQwn1TISZPDkMujy7czuHHXMm3eR0YGejIHKUGWMfarmXwhpEOlm
X3rAT+X0PZRvKPgWM4fLUvwq/Dc9hV4i/rShMeOi6cNY35U03reOLrDTf0qD0XrH6RdzaYs/xVsb
+UJZIx+LKD7e4EGwAQr7FRrCG36/xDZt8/goxGeCLQX927XDDhEANlQPD65eXhVFAkWBlrLhcK+c
fSt+Glkhd/TZegnYPSDbiWz9DzqB8bInEnOHoQvQ8Y3Wr/UQrji0w79NXjAD3tYLwKB1eGb4BtVV
9pQcltdj4jBF0q9Qx751JXTdNR7KSwNUR1QVGFnNqSjLlcWu+FG7PJMVmjUhWSEnX9FRovhGAAEt
YhsHwZjCgDxv2sTdp+BT81jgfBJSpViIVbfO1nHD3ZmjE3PPhKzIKmxWgRn459OJp2cUDUZTqGqk
cuLrX6Ku0CQUEwuBcVJx6VcqSCx/hG58AuQsQbNNFeDp/0oWfCcCyBsuiCWF0ep/QaBDCrFJKNWQ
JZTXGExkrfN9hNYUobIUFB/DZjbgYkkLcXBS2JfCoZetwWhi1AyENudkmWOC4oR52J0excdojXhu
Npg11s+usmJkKKbWVdp98FG28VJapp/QoHLu0qpMQQBYu6sJ9D4dzROwXybLMmls02pALExWePak
mXldr5jXaeXh5BH5m+4+ueqD5Jt1LIj77P9fEu70kkkZtFjgZL0ly/ilPjEWazKmc9R2nRWSAlyv
wGpfJVHbpqBtzT2Yoy6CtTFRRz+crtxD2RqTKCYI0WZCFJU5oyl5afjy7G30qxmYAkID0oxvpaTQ
VM0WS4gfMf45GEW/YNE+bvvuT1vRaNbOI0XLNT+yEHksUzlTL4c7l048teaBA8zCA0ihBGlRQ5tv
o642rgaRJWEI6fC/2XtVVScL4lmYIzFNTmTznNUuIzAdGX3ZLgawhBnGBj5bkIDvZiwXDoY+4x2Q
ZZMYGIlZOGz3MMGTCo5gkscDcDfLlUfeyTCfzplLZOI8t+IFKhZ5WE6pOTF+7ubrEAMqoje4O+m7
GO1n9bXH1K542PXNSEs7JDZp1yKiNsbpywIuT9nEVJQuDBHBl/D1sDCTk0WZgxtQ+ixZSaQLeTQf
GVloDuoCbvfYHsQpydsxkQaCk0Ypl9kP8SmxRyPn0II6ArmqVXN3mstZSTYEm2cwS3sUWJ9b5Yub
pQWN4gMAPbpdJx/d72AE9ohA8aq/fE91CFAZ2DH7w+edVYF3/HUat75W98pOB+poed3LapFrlt8L
Iw4fF4/cHL/lSC6mGuRRfjHpoHQxzRcAZVG8/Q4GQuR5/y5gA3HkqCvFZfIPkRsfN31kMVGqjySY
VVrfOt9U5zMAoo3K9RC/nuE15d79gYBHdIOFn5OjUn5NP+SAoaUVeO/KxEzu4DC6q2h1JWktDV/g
t7+fcKl9sVqpeOZjYiqdFYX0RAB6CVSnDmH6R2hzW0cuQGRzCVMGEADp4brPURLiSqNxYkXyTG8w
i3xwje/17qkZBu8+qxDQpCdKYMRcNMLfd0cxjtVYJRMNTSJd0d6wYbfK+VobaX/GWJwu0NaqCriZ
Wvgmi0yrbLe4Y4BYNQK3Au89HQKiuC7zdA0FFBAmsHKTPM1n1CF43QbxHKwSnqXz05oBp3VkXEKC
v5tlmBWZFNT6CWLOZ83MlVx01fzCclI9HG40x7w4FM1VIg/2/QuQyq2txPG+Thw93pg0iiy/3jT4
V3yH5/BCHb45I/N6yyQdE2yLdTjc84acQe3qfccTrnpl1Zryc2MyDb0GI/kuodkNJheTu3ytGj1j
pnuyu9Z5wpBxxl8hsPvMWpuHGoSbH5r1sfxwzchzPEA6iXcrjUjM1Wr3l5JN2UtPwJgYj67WyWVG
E7x45NG014ZKb8T7wlgDgtNA30yTkmBuCefGx2XnMA0a20pbbPCEO0uqLYz9FW81LzGzO/k+wqzv
3nvqnx/OSMi6aJvaIVyFwpQUvl7MUkRhxroWXzuJxVgRojGKihus1juRok1L7IPC7G6AiLPiwEVP
GXTQaxC12dX5W6NiAkoMSCCCbLSWqbYCLyoHMVLQFLaBxuPAACedNfem0cXWBt5Wx590MjC1OVQp
2CwPT08Q8xzDm+jmSY7y6kLc+4yCz4OjdO9u5Az4Fop9C3Wwf1i7MDTxGCf7D/vJ7IiMFDKej328
xVoUnNjoh3c/mtOBwixPN9js14HfcnEHDTccw+NcwcTW+ZBvijqHt610lDaKr6+fz3N4tKmQu6EK
EQGTyfWAmM0qI8cr+QB2ftCglxVja3WCkq5YYiPjcjZ4bIANvgR55rV5baIX6NLFQARUzdmn8JBr
SeSLm2CwjkFf3kkPcMIkxf1SZaHXYwqLY8egJZbxHDwVPfA3V3HEot/wgwz1/IKeVkMoEuIQ7tf+
IwNuhBPT2EJH2wb80z53sChPR6WuquKx8O98ugSmnw2oUWSW635H4azdQKaOm6nhU8jVijHPPXzZ
DPogWGAR3OXpgU+nSNGl6jFqXAGPFSrMhZkXx2RK2kP8vpqnjS+fae1ONUwTzFq82FF1uwvq4Kkw
Gvi5Pa5io7KYcqHmCZLdjD4iRc3rM3vVx8rOgnBz/QJrE3KM1mMWgoENLFv/XGK44poz90wDUzpu
igVX63LYZMJor6uOVus0qY6o1xU2rpqkPKaftZgNJimqUGUS5da3AILyYktuquK38bpjxRn8tbR/
xNf26QlMFzzbUpGs/J85XMPSCW3EtsLqQfluT3YsxuCznoxZ52yf5g+1OLYdJyS7kTXEJuM8KirF
nxeRI525hNvnOSrYd8rp+V5Xq2QtJ9OmDIdVB7mjGjGP3C7LgRsDiK/Y6qlSd0dy+TWBdJEcp4Cs
AB3B+Kxq5vcegAtDoYWVo//uLmAJ1BgvEOTxzBYCoDeNm0ZEobUAVMUEIyXswb/3amCZS4pgeYNa
ivYx8Cvs5ASUDzCQLCDyN4UkPkV86yMCERn6s9fK3B6ueINJslYMCUKnnI9EXiCXQss4wA/W+dNd
NbGr3EqJNB43qCPHQgnmPqiCFObMJrBKBbxHFjmraNQrvBp3VJKpfLo3KY//qabbvNcowDoTEvSj
hgxzLWaSWaA6Ln3ogA95bTw+eAbxoQuZK4cIOi/2o9m73Yqx+E5dY0bOsTW4u8DCVvem/mzKoobC
dwgc6y43k8PkbBZHhw2e9eLnfnofQk0ymBnG6hXZUJv7vaLyiYiDWU9CgBvfZm8/8AIidmceRz0I
s05JtASUtY3/4bb4n6uf39neo7TE3euf3QFOvZ+5XqXqQLTf+DB/lb5WdhK+xj8DOTttekezFl24
FTLRIa3L4S5DFzC8kqps4ElE7+WqxpJPffEZatsnK5anyJ3lNbmHGVeO0NWSnK9YrwwngatOKFwB
qfIYBWbfA64MpIT4ohQTfsXfBAiKyR6q/OqPcssrpEllTm9fFQLrJbFH/WbzFVqLjAhTPzuXTfgl
Y/Kwu8D76Yr+BMlQDObXVDlRWib6tlsQJoyNq2If10VvqZT1v9BLxET5/0vRpRSR8Z2GPB0ITxlL
7KCTdZPxG3SFJ2VAuzdwNgnxB8E6R9/Ed3I+A+IeZU+TG3RH96i9s/dTEt0CZoaBTvBoAnJd2YAk
YdyHKk1zmHqAwke3c5YqWqQZG65dTNJIdYB3G8q+JyUZZVdqP6eDW7HRAbo/ev9U6eqINJ+hRH8e
gK38g18R21JSTvGDWuy3peJlb+3KLhAyGg2fnewe67oShiqq5tce+3Wm4SAUHUdhQCPRy+IpvR6e
qAMRSgSL5nc2dm0F8TY7H7wQB/kGA6OeVoYCrDMvqGBNfTLBFHHI42qGKwrwc58Chw6krMiLgWOp
xajHh5WIXIB+R8UxaIZtZi61XH8D8Jv67RB+1uzi81PjSRS+hBIVJkrgUQZoI8lZ6gHO9PU7nmf8
ul0M0wPbVhD0quHksDC0u9vjnkM41CJeJattNVAl1LpW7rqG6O2MKAueccMGavC32oaMTptFk1zv
EuzWMZ1urhDyg7oFtWZg/byTAi15gd/Kd6dypmA36A4cDQ6gVudCBF//p0VBhjOJYbODMXVur4Js
c5NNJhqCXAR2Ylv9D43W9RALHIrBG59ySF/8UIVmEz2ufSZdwX/tvmRf8HjdteQXlEley7VvAltQ
QRJ/kLdgZNPrQtKZf3Ud75wPEOSxDiE5M9n2Aoy3UX8isO79DhjdB5YsU0u7kX5HmHzlkspSBxSZ
hUOamNVwXmI0eAyKNP+zQpIYJL0WWeSAfRwUx/8oSGJtAC6TOtWAVMriA3QNufbXfyaL2WBbP5vr
fNs0A8loQLRzTQOJWcNMm660zkDfl3prbOviAHU3wCB291KKSnqxDYkYmF40xDyJtbF1tjCHe4Mc
SQtLGIrMz8VKk5w1omZDL+Gsxn7GbvUFo4E56jdKN0rUYrAdKMUPwlRTwIbuGns/LuLBcvkfObJZ
GPhiPSJjzEaQQu/35d+zdBiV2gqMauzoIA9tQs2IcnCUFyQXqmd7Fl3LRE5xvH4+FSv1K0CWTE0I
fNU0/mlHSk1yHPYtDCrDl855pwiSOIBxlywnhoO4OBjJkIeANQ6fG+dV2XgwDS08/a/9VQxHVPYA
6Z785JSKoZ09ssmYLzCWkueMDxV7bin3VJo7Xah8I3oxD/+JmT3uEoMwYS01l6wWLU0jJGc8WQ1f
CXw6gs5pE/nLr4DkA/iBzQLaZIWTm7uGgZvuhD7x/sXkW4C37WBxoQQEqc4wLq/wDUWAwVQhcLPh
pFrACTPrxJbGSQlWdZ9zw3vkjSdqTwUKUDcNPMmtJeE0IF58vBoDBvefjR/v16pWKE+7kj8je3Rv
LeHnXUL/bvTnYt37T5Mlf9pAG10QsYutWaA6jrqc7k6BauiTgWtrVVCneHKUW43ehMLzB48bVH+y
aaf6CqEn564oLs378MzSN+fPwuhRkbJfBbIrt/Lwu//tFw749iWhnOG6UwFYXhTVS7ylPRj6kCBB
PUAMJC416TCB3YNJDiikNPBbWkvSKeT7em1HI/u7yq7IytIFY80Gnh3awRs0pFTCyJp3mmkCV5eC
x3WEaXhfPX7yCf3Y4CJBhzRvQbQi+c2ZVGP7Dx8WmDc7UH7sB2+m1Q5sJubbag08AZN/z02VFCN/
6b5DhqkZSUBfUsatwBnp1427q8pAVNQ2zZdw3vFE6pcGMZD7SEMg0/PZeTXzq53Yar+PPARyh366
A9s6jkTB6n7Cp1Abe/ovgP8khOYqB0d5qPysZ0HOHf2+uY4+5Unj4cak9z3MkB8W+p48RI29XXox
wcajSzLwnVkJM+zmNA/jc3WzWYMcsTMxXb7S6UdYdQQONaqFBeHIbvE0WbLnP3ilqgld+Cd1w86j
HOxvuGPpy+pQ50Vr5MUI6cZgSkkWuc5JXQCo7P1kHAqlmDeYwK8WmZ8mQsD0oOP2CVca0V/sMR4n
r8a8lP0smhAT/RkmXFDYtbOiQneH1jZgCW3Lxf3dbqZN/AS02VCghw+8BNKES4A0Gy5xDv9KG9SW
ULJQMTn2RapSSzGVkm2YroPv3+oHSa6XiGT861ahRHXAi2NX1PXUYuGcpwRbz+t9TiI8prZ5NVSA
aku55k3lDvZOPD2pFd+PnwA9jpUHByw725z+OKHlwyImXel6yON+CIJ++6V1zINiBx3VhXRzksnV
UsfcjIh5HMbIL5vb9opoovrvgt/IEx3mwSnsSFjUlmNF3jVTTCEVssA04BrKJSQ5JIPXNxUvNGFo
GZBNtLug2UhukMpqVViIwstUIaYV93cj4qY2eBz8MCYowoVZXRTJrqzcrKf4o2ayZcxBjyylTzFt
A8JU1q6MIitXwop2ET0UHWT8TeQroe2iENDYilkz+BypDPkOmfnc8FgOIbmqLOAEOn9CDf9numUr
UDoQIVj0hA7nkpymJu1HjgENRN41MKau72kgGULLEuIHlTItjVcWdYuvdP41cKeu+yXS11WN5yrQ
tx1ZAmJeuwCDhSI+cIgLMFQxUxUYQez/20T0FIuVIlXvV8TCbiuvEsm2Uj2d8Lc4y12/EQ2hdeHi
wCyIk2zpd6uiQzTWiXG04IGAGYevMgXL2JJIRMUFxgLS1QkDEINhqD065tWFlvvPzGy8uJ4bgb3k
CnApYJr2P5y3fFarOSp85MI/mDHyk85NdqC6uRuePTtD3xXnNGzTmq/AC/zObUYApwypZDs0TeY7
VZU0lwwjquj72a5gwBeJD90nec151kq83hOpGf8u1MPFQQnyucvI3nM9DBmrtjd9EyeP/udy5+8r
BXSk4twEsSLbUGLlNnaQKulFnYBoRqgVhBRaObrQL0arEJxa7BqBndlQ8S2VbUXQLXCZGCcgBmZQ
v8uHMZroZ+Ne/MYKoUQA0+oiqgyXQIZyRuAfDrSzMX8sym4FITFNZE8saSkg1iI/tT5K7fPaOyJx
cLXFJQnjCrY0Jds9JWo6tDkKLtsdet0iBSXh1hyujZGpy91P69bYUl4qrNsdPgvEHFtRJWL02G3S
a679/nUNpUEGYoDqtIsT9WzT6fdpMLntLhRnIWawSNqte2zQX4iKSpa3CHNePpNM0oPz51M6Eo8s
Teb5lB5GDSyQgcApm+/2MmDNJy7gNzcJGW9W8T1lKOdRYGJkRo3MUG+k6LDSLpPcPkx/HI6Gvda/
Ul9j8v12+vxyKFt8udCqP44lMPHO8paxt9yOxkG8zpgUW8Qrz5jGHKY5N48P5WfBJ/GwVe01DlEc
j/4uZhKvm3JEuZ9WwBW+y6jAgpriTySUktCXuZCA1eKMGOajyRkIiajvqpqnPMyA5/oaoEwrqZFd
YP43suIJ86E1AtiGIgGU3YNj958R7R3lGBi6XbmMMA3+ktXry/yMC9BoaGIfhrmEH7nbFjB3frZ8
rgbLh7NxxdnsmS5gjbMOyPLwWgdk4C6uc4O8X7p3V7Ac6BIktsvf0NcSU0E0J80ObElsHFihCT2T
Y1wvFEJl7sx37n57KwIM5LOXCmG79F8E8nMWdzcAqsc46sXjlr1qSGsDEIAI4xeN9pyoBnVjoBnU
KkVXM6yTLnXuh38PVfu8guU+VmrAAdsCd2AAkAx7oYqpnBpwRlU8aAtE5eeMaHoU4SFMF1bdYBx8
vik4snfhRFm56hIzovWOuldi4Z/c1kOTv0K+ZvUTxdAeXdS5cWHGHqmNeeEHhdRCOc0vJxpkC6BQ
cWdBac3qml4D9FPpDGnr+IjcYTSupElv+k9JB80UokPC1byIo7ofPYlYXQ8hWFUqHOkNUcEGlRNe
Et06Kiw9eRbmJOrcHtMAeRfFoVI4ZJHvMao6XPiCZ/4rI/W0OQ7HmZ6TZI674FKyOGFaEL4fpeP1
7cJvbts7Ndqwj0sozVx4fsqIyBTfxKJapu2Y91fhVDwKEqgYwlXx/92+snjFQ200C5uvpU9Lw5l3
ogpVwwL5b+OAng62e0Z5gKi+ZOvTRTjf9NtDTNZILf3rZ32OApajwzktE+HrnXpe2UP8VA5AAz2S
ghygQ2D8djrNfZj2t20yO0qNytNEUu/aL+zWi9OAZqsqTSrX86bfcoD/dmTT2adDm8OsPWrnr0WD
sLGyDO3Mm3rL2nnXgthLwYjfW9NQd/8KPjB7AGO6RqZX/BpNVVSQgU/cC9AvK1SMYM27FcM5Y6Sj
hQf1fSKr91vm4uNTi7Ofv/H6+YFCeYIYXZhhN259HvdgAeXE5fuycnTWaYz8RfoCoht4bc9MJFUJ
NwIoIwrUGlKrTq6kd2+57i39plD8RrGYi0JavjP6yTwNEGF0dlqBLAljYQvx9Q3EBg/NHpCXI2pf
aEQWOBvp6Kdzc7PT8pkxZmswMqvvMIu7LRd/8eXFVxjVBL/BMX3QVRcB5LdQZx188ryYUT8Gyqbo
R41mYPiBxB5Z9SmpALD9XJ91+w8NVzPHzkjhQBDl8nSw7Hwbhk0e/To9BTdq8kSVz7niih6vWLj8
dLoveLNEKlY76xkjAQbqfduXHtHnNcu2MAPSfQ6+QvN2hk+m1p5A/mDyhdmF+yw+LmtKPUNAit6B
z8nDi7eau6l12ZwWJTrkDiRTMcgRcTLJh1GK8Q1wY12CTXCKoNDwBxmPmdaNLar7p4HgLRyuU0sf
RPOoSV4ufcaObviUWt7d5W3p9oYOhg6mlRCCll23dBDeyWFY/zn0xKEBKwYBphW+nG0d+xQLw0RT
bx536sFWTpzC0fkeU1tQ1zd2En1OC2RRjvAX9EYcB78fpT35OGaSzTgwZqB+qT5A1RjzV6NGpqNH
atP88sIV0+Zlo/XzmcYrNOJpwtEr+QqRYM/rffdEsYERSb5YHWANyeyzwyUZonY48WghtcjKYBcM
VEvdvbDOmRtj7mpxY27xeT80e7rypzAnKpJgIhf4yBAjlgTVMHV8WSJUfvSzrJsbygD5eHlfiRby
lqCLDL6JxsB+rGflLsk0c3420N84DuYT6At9dlsOqxW4xUzaTav3sI0DRvr2I9fRz0m39YUCxwKU
Z+5fqHzFB5sEW3Uef7cDHtz3JMSuExGT3Qc9tUkDBKW2qgUnwG9LB0xnsNo7MuARXjVRM3sIVMY9
XyzkUMPP2+r0f2shXGooxPa2x7j+MEblyffmax7n2JwZqapInmwbeSiQKMqDhgYxtETlSztLxsEN
D0qgAzTIvjjKyoY0rzvL0DjWCTnwf6Dlbz9+NoIEKrBWUzmZzMVcludEUuIGI6e5C6MqHYVZOHFi
LcaUHNgDE4LtLN+9iQm9r9DlOvZtpB/aRXl4aSGSG8MyH1Mp/nqfgfItKqkfKLHH7OAgwphkqgzl
0pltdvkOFunuVZg5b3EgODXhyOdra+2Li9Dw0RnYZKLPAZS48SbeNOAXakI8TqM2n1zSNZ01y13/
Iz7ImnjJ1vFQMVUXHpm5sWFyaWpqiQCL7y+HeHmueWAVQ+0/eOPzFULL04CQQ/v6tgB7VNMs4XwN
CtFnUx86038GOD74RdsW0X2+nAslZNZ+oFyZo8d26zBIdDM6jq7XrbwU5YgG2eNRwSqh2J2H4QCI
fTOk0NoVreYc51XwZv+89cFHkQm8dSpK9Lxp3lpfUscPAipAnGHsiQddwH4NukXrzny08S8QAQq7
KK66sTanFsHfxhAEHTKjERKUn2w5s6JymrlNGNUYPjrYwI7/QYjNiT+DITxhrZXeqRc+5zO7wt8K
1+NLYCY0w8urorywFXTCzjnqqzLzS9swz6osn2Y/upMa+GLbMefIl7VqY3xRQBtdDTiX34T43+8G
jbmEWyHyejq80L4Fn5F1ysmjmdc0xHAULRRJIE1KY7afWjKdEk5iWLEBgTTAZeXlZUM6zcRVayXh
LskruiycZFjZtZ59WbaJjlN+LUzzQAwoStvIIWpuA2hHmp5rxcicmQvi86dZzEoBeedJPuuqqdGU
j7s4ddpjrdAaSH7D3f9D6NBlNan9dTAUYTH6TRLiJ2GjHCHvwG0GX1ndOGeLV0CZ/QTZsdPMAkB5
DMryvC6kCW0AVTUj4dMqJDGEBq1D/rYs+q/IjvloZ1GdNsAPbw/bivqw+NuanWC78JlG8C9wblT0
bKx4OOnKSJFmZJgg1RP3DBxQ6f45kLYDnc/IVHRtDSYs/cUiFUpLQ51lHE3JuJwkRFx50wZxHhNz
YSayA6KbWtLHbLk5r10AZslOa58PQBE5WcL4UmmLaIVLHZt/3QTgdtMWjH/gzLCFJ+T140G3VXj/
zIpCRDIcgmzCrKMqxP73sO75wtsZQmnztDWGfFxppC15JsjfyVuQ3cJPFr072R+KEW+ITB8NdWNX
R/x2yfAliYcajh1kHs+t/ds4XitTtqW5UjtzAKloPaI4YhcsXvyboNXt1DEOSkh4mEbViqies3RV
Ajh1OVyPX+kpG52rE9yRK84Hh+MxjmkWsOOp63wwgeJGNAQOhByNkaLd494czYlhaJCVYwJXHmL4
Md8TJHyKU0C/AriZWUVEq3pEUaE8v/tLDPJGN51nIY9tN3fh5C0nOtz89SEEPNK5mKGDcyZ17Vnv
akNm9AX3aqkvwQOWH1gtq8JXZisrYF6VDMcj2Z6AzAEsrDfu2dgNsf0ME9wh/kM7pwegxHePIm0A
SNSr0Di+wDbvVUtEtsz7OU7TzV6akDNvjNJe5NboeYyyJ/fAJcKEpVR1K0CTRIL0h0RpD+aSavEN
Y1r5Tbx9iHx4SjvrN4XJhYwuuyRDRm8Pzo5eTOB05/zcQ9+srPtDcYKj93dJ/WKsE7R4D0b9xWyK
Javtb6EYitwczd3oJ75ZszvdeDZOl8669qvLXqrrp/jXRcn7y+OE4RzmnCtWuiRZ0Q+sE7Rn7jle
HQBQS2oIW+oDtFsOGzmNVDYgv3faGDu+T4yU+RCjGGaC3z4ilPPCqjXnuJscxy0aAnejg5ZzNfcx
b+yx53fjnB3jgRdKvTqduMR2vXo0CuqVCTxNqGLaAsS+iMJ/e4dGR2/AaoKbhR0rfU9jOfCR0jdg
TZoNd1pEfbHWuWTN8ijqalO1ZYjbs3TnDQgT4QFhmzjMO6Rrj7w1QsZxOIi67NkaeFLAaM/bpN/E
VcgEtKF0BAJryI149RuGwWp0KbNWh+a2y37B2/BzY1B9e2KPAB0AgO12ojDR9UbyRd2OJVWAjZ3T
TP7DuWG4LHwtFv/L3bbX89stMoKhy2yUVR2Ef3NZgHlylR+NKeJrBkdweacP8dQdkVfdtfVFK5wz
VtEUzFoTGZlXPGIgr2TN7wP5iHcFcj7cD9FAVliV5UgBo1PfZT6tX8aWmWwm9wP+n7h23wcotMui
HVTnsa8UkBFXSCGHbLB3StqGJgyRzkxMNAZgZdMcoOdNmSZ/m2U770y7LNze3QehB1QydqZwGcXD
hW8mAcoXh7sI1AwLaqrb9Ox2lV1Y9cSspadM7HLBFg2OUzrN24pLCSgsFVJwxxj6AXB7OwVa6Jw9
wnLRZq81Jce6VD7I4Au9VMGvVA1dAVsV3Vv062LhlupW607K460RJSuK3cPDf4AifhZlF/TQ2n8r
//GRpNSnpheXTemR0N1Gihh8ZrSSA/IwhLWtePohtXlci5k2sZepVGm0pRmCWmVVjagl1DmyY3Pt
trJjlSpUtjSmFt/gWZ3tLzPclcW3IT2eo0sYEK/pSC0poQ+xaDuWqenTl7gbMsG6XAMCZfaP7I/w
5mMxJ7NusfTOBCbgXntvSZxecBBHTrhcJ/RH2SJw43vNdt5VDHeN02PJt0sIcN7e5txSivV3mMSE
NcTeXwt8ekBAE5whplgiQQn2j8NsIrjPVcGNeyG/w+4HgvKbyp9JoDNY7pnn33N7yX9sKkjB0KEB
2bWrxG2/V0mUzzK1/fKpsw8t25TR1LuXvi1RfSQyoU+zcefG88Cwd/dJi05C7Db6PGyhkXghlhNz
St2/Lv48SKBxDKBJ5oRfiNwiaO+kS9u1BubF+DvP8o3jNppNlmI6m4GaoQc8dM99hxnndifb0VqN
1BXVLJbZaUEdX/VZrE6DSfJALCladEuooJxTthW03dXqKKDL9yHx02yJSyCSpn9wn1H1bYUv7Dw4
hW2NovfjNBmQkqZJmNtu3vGPvA72uXmCJ5V/02NVaUNx4ZfnFD9/1I/v41iZ1rTReTjhTuoUcfcn
DHdR0Co990b+pSX1emxqNbQfqaDkSm91M32Y/zeggUbB240iuusl5JIqGfS7+HFZzNbgIzh7IyO/
3n04/EnlVhTOfbbS25o5kHRm/UraagB6l59HsSpwa77DSGa5cISWVfC4FYVZzmS5Qo8n6jfZpmZ5
hdWvJqX+VE/ppMLbmd/+j4Za5vFQmMp4vYzSl3M9WUV7Psj5Yy6oHvu49CNcTZ14X7fFU+cV8DYe
6szwe/RofM8buE8swyo7OBrRiUTukO/5VUYyMW0J8dHVpncoDjrfYzOSpi1twJvIi1Pc3Rr3lRUL
/BFXcjBv3ygRkuzdWvvXvYhNivrmxIy8a19TCvh7H2kRSabLQv+QNCEiTZdQpQfVbEaIhsBEQiD/
IV3PEI/wZ3o9WWdkjCMi40Xi84FG+kRFzjRhxmy6sbE7NbNtYuuVSQ1T14K61KXMw9SlRtvc5l40
k5mvaeElz4nqGRw2IYlHE4JFxyiT3+o01VrL7vUnW8pe7HuD0hBF0KSMEYpjhDtdaaB1QGWLEJtO
ViZueaMVdkD02yhAX26Yg8v0HM3zK7jPzSR7dC3RNzpdzNcFVoatTZTFkX8a7VX4vUM0qlSI67E5
8iFtlG7w7knnZGasgZqtltQTgxtEcqWSJCMdn3d8E6KwtGIywnvPzbemDl8pjpkxXog84ug0sTAO
92THCyyJjHOzr3nnEY/DZLTWYEjtRWis9wgFHNmB5H4JLOVdvI7+8zpN2FZLhdWrWAxq8wej5M//
3x27PQCbV2RGhNU46dj4RyNQ79hVXVUvp9tdqZV03IMu3IJNPRgKaQMBKPoR324OarpLWJ23y+dU
1LK/KvH+r/ArJ/gUOS+pzouJBOK7+kS8yAE7vvKM5LDht9ppSEzMxIAcXU/BFmOROWWKk3AVnVxI
Z/s8QGwbAYZDwfxZ+wqRIxw+Ftxip67kcyyzaB02Y80OEiQqaOejWgSE+V29zgzYaLMw+c4ZQzKe
IMCIO2ti4gRj1c0lC2DpGgZCZ29rFcOxc/fRhqO3xjm1cDQ/TwNJ5Qyvk9dOAICX9vXdA3nytrgs
xErhsSWgslgEXRQfuX+VQ/kRlx39PwR1Tx4H/IodBmBh/9PwIJa771U0PpkxGTMGWn2Yu0TJhpyE
oFIBGIyZ+IB2X22vBCF19WrZvTH8+Yf1uKa0N2KV776HpttflU/ul+/MSmTr9NAkab0fFidJ4XpS
y6gGX0+gXWv9QJm4SZtiJVVsT3dT1Npmh5s2vazfzVgHMDHRTIMR6zFRM29kq8TNtsTxdl0u6zd0
SrJddAR+osL6WeFn1DMfFPvt1O9H8TjHOJkfMj/Q80FF0FIO/I9ofGBKg/0NWBzHLlp3Zv/DirFS
cG/GW87/mLFugDT8dil+bTHs3sIXM67FwXWlHHkVePzQAo7QEncySvitHuhyf76s8EjysP0mYjGW
VUtHapMUxwASx+lu8PA88ivr3f0e+4lmlQW0dk+rAFRLM+M/Zd1HuhhYtZCziisCAMPfz3P1V6np
gN5PdIS9wUT6sU+M4I7a9Vk5ccCQcNcqtB/OEyqBc+GwvAv1QYHWnsfWs9bKXI4JczKLkrw7fZxD
32ZOW/09dmJQNdGHvnGPxU8Rpp5z6FyE9Terwl1Lc0uw6BSQJlQnVKuipfPt/G9drsHsaimqKAoa
KF67GSR1484GMZh4FIAWghVEqSveFPpRT2WhMIqN4tA1ee/l4hgoWSHXypBik56O3oJtE07MZJIX
679zwxnpfk0md0QJw6lj6ORnfRglEsqBursr3qE17wWgz0z1rPEfIwsDxNPS6IK3/9b+VIaGv6zg
mRAlpAzH0jh1ek4kRQM4Iya8mZ5Qlh5yX+/QBPdYZGid825sD/h/1QZf7sxU4c6s6lN1iOZ8ahhL
Awpt1LVzzMaBKtj7aN9DjNnsXE7OS4gm7e6MyUnF6sYi7sgUfh6jVR+9nTj9kz9SJ2Ls4AB6Bawr
vX+TThRHgFwRwaxw0B7pmt4rlxGQ4wca72srbxPZzpJmowDKaIVTmNhkiMc1vkIeyNDvBlznZBGP
Z7n+jx8OQ7RE6Yp8r3AT0+5q55qNiT+9JJrX31n4JNcXwvGd/nQCJQNSkGCTA2RFAHuAN9cyYkP8
mUn/VtzPIXNrWqpgZBlmJ/0BI+/XchlXfPpY8nUiTRvb5eC354fSlRmr2oMXC1hi6vgE1nq6bsgD
5yj3py9k4EQu17xb98bBJvE4FqusLPC3CEARi++hM1lve+tlB5xLJVNLWQeU22TS53DkKWlivXkW
B1U0qUINalHr7SZ/5F9LXnRvuGlQiigWAGPHqfwx0bDm+vhwyAJASvkpYCxkKl/cWaq+ABBiv5w9
jwXL52W6AoKMmrD8sdQPCFUTflia5P6vm7H4l/eglAPvr4JK+T5Q/rZZ9U17/Itrs/BQ0otbuHu+
D+6E0Sf4Kf/geD7AJx9Ee21NfhegkZCdg8hMWe1ARNsijLm+itdmDsp6wUCTMLPwNrqDqBLX6RR9
TGmwMInWT5hxjguFpduha/WXJSDUw2IpetR0OMDqwf2w40YxAh0m+9MAJDdWEgJPt0Q8ZEa2o4gc
Az9dyVDDQeP+bNQ91XPqV1NpKhJrZRkcrvXUpqYxgs8Lxt16+FkNIItDIClB5PMoWoxUa/6HjAL9
6EbxlqPdFX/pg+/ZXH4XA3J4Ye55FIXhIBdgwK8ko7eWE48FIuNyAjYiSAMMsWCspf9OaEUHLdEI
TnDdUxMGg5dsWO8EuvkxEj95Pu+5nP68Ix7fXtc4ysMY364QLRdoYjFsv/0czlJRrr/gihAbV6eW
/FVxBtLS2eksur2YeRF5rsAQS3SkCu4Ix9MRUWKIurAFxBd2mYv3S4g8bpa3qLFeg3PR2mq8Pwf6
6DaSrkNVR6t059qqiSJLaVFWPGmSGTNEGKnLF3RI0AqXf0n2Wchr1gkz5pdqEAMVOqw3KeKCSG4M
uxGNEznBHOO0b/fSLuyNrYBKzokZmOiVD6gZeDGz7F+EhSzMFB7u/WbrGsn4iu/l4ssTAcNKfGRq
AcEe2euzBWYquwAZSlDukrTvDkeRXuXpRHuYEm7J1797+rLO9ZFhywTc6U7jy43OGw6jr51hZvU8
oOdXjHMuBB76poegTD3mGHqpoMg+ly4Axw/faBK+OEqoWGiRi8lP/ZuMyGjDeKyXJPi5TpMKzU6D
/BDIGhJLsfXZ3sXmumI7mb6+rIm31luEZlMjWHOieiWjMz825aHWZeiy1QsDHA8lE8+FqmxZ1Ogj
S6tAjsWPvRWyku7d2FWlTz5Xfb1COBqWTAr4q1I5iqJT3hTWkzkMSfWMSnWz3GIwONyhooIvBZMT
b6hwiq6OArjKTB4WUmNy2bMyryo3B5+RA4K1m/CT3LGGRr6XTcua00t15H7RLMeP4/P5wq6D3+Ty
/qxLG3UPzKROkDFzER4jP4/BueyUsEqKzHqRwxMSxdNTovT5I5yn/93qDHm9vuO2RmUdDWo+PzP6
MLra+lB7htKIaZL+77JS/bG21+6lXT72Df+qWXYTD/U77Qh0KYieNsPK+bkmZBoJ5WjXKFzDseRI
Z57zRE6Kff+rOJBQUNFKC9rQkd8v/EWpAE9owSQ3pvvLqRH0SJlZLEsFBDEv0WJNy028qFYdqdq6
aZSo1SPWXJGSDkOqwKgdxRiJJHQAulhc49e+V08IskkJamRQgabB5ckLViwpgdIfCv/9VZbF+sdC
266B5qnP5lgZ785X0m65Qd9cK8+bJqGzaXi5DGIpyYkZXVvb9H8rAmP1wtc+Z0pU6xHWBlwBspOe
22BqIttFtYXzPcKaAjuhO/UrNBBUS7yGoq5GD0iyU71uMs1FNLeuIl/dTrsaOvh/Ciy3bL8slu1R
YJ+lLuHsBEA+r8OnWEV3YWngCeWNfSpcgiOImCQ68XijQ/BSgvxS80A4vBdCkb6cZ8tDc+ZDXFyp
ahCe86vRfR4+gpzSR19uEjZiCJhdncx5+i8k12+N3y4ArhjwbcsAtPp5qqNyYepckisMig7uXI7T
B54VVV6y93r4p/ez9pAZZkpHI9PWnT5UdiLMY3ZzDJNOvVWojpHGvFSxWAxYyWoa3qrmSyN+04+v
36KLRlmZ9ON8mNoS/w3OZG4hMcx2xEMgLplKyAplkLAgPhW4vZPm5VJxr0LiNQjm9pNoGuFsfYv2
+sIAU6b7JFXL5XCYr0ebiGDiCPtEYOA9syCdZvfLzWsP7Kc/Y48YZG7AFVfs4/zWiq9AUYiu78g5
bXwqT0zSn8BnikZsXpJFbCvQFWWx+sqRvVxIMjZDlDyyhhH0OExNx73/w+Uakn22IfhV3Ef7BJdN
l3lAtySaA4YoXEIrUViffGO8jarfTwWHm5FveDEaMuGl2uJygU+G/SNVXK891KE4zu3seonA+yFR
V/u+tOdqOhkDkIZxEz4qoM6uRYYyq/D28Nvo7q9gAQiEfJgFbUpohV+Rc4LYOYHXCkvqNtqXmTvk
RonRkAFv3Wzo/ls+z33GSt2U5V85dkZKmpBGF7ngFNu6XFZlj+4EA1bEZdEgPLTOt2FFbpAJGLQO
Lj49z+BQwVpokmCMQ6qR8x+i48Inb697OjzHRrel70a9paolR3OAnMYTqZxyktIKb1dFdRlp5EcC
mrk2s9wQHpWA8xkkkoBnaEZyCEkwBBPpjmkjpl1+2rEKCPSVHDG7ynU0KiUhedv0DRZmnrpJqdMs
uU7/hvIWWiKmaLXm9DntDK/g4qQ9IfHGSrcfNxKuBZ9kWK7ph0cFrGmCAnK6HQLQvBb81b+cD4Sa
HK1rqGVFO9nLOWZJTthu2wHiXGb3XvUbGgcEDraFkV7j+ZWlxQ7hVE2e9+Lg92x3AItUkPg+Pb/H
PPuKHXN071aiXREIPQ+ms8MPkqxZbD1qJftVex8zmBtwNBqmJNf6cQVnSPJ/Lx6C2OXbwdGhdK7+
ojb1wK7hUVH+Yz7eeWfW/zCo4e541mfRNcQ3nEYcuogSAtyTnqATxOcSHlycmWB8INB/WxaSTi21
OGOpUnA/SAhLtgau+zUlOQSpNx+PfHcnRd5DdrFy9P8na85wxa3+H0kfthxSe81Qkv4M1AZP/y5a
U5s2oaJxFveM7v+x8inSiRgstCktdEvwo5MuCdieFgkDPezA3ZYw57dQcLsW9fB0X9JfrbV/tjUk
2x4mpgPnrD0+hesxhmowPRRrwRYqUnySFNWosRXTxCS9S/ThGcSFRKX9icoEf9Gnm4x4DTx7LAGY
1zHsyOa8ZcRLQ2RDX4vVHoC/c/BIEjlx2YK9rnNpbgvNUdoYuYtFtfrtvYBCO/gKUmGoKjDd4TnF
0OUoxdGCctmWaRtmLC6Hc8HigWE8U7deq34fPFSJTaethdH0CKGynYIWSUmPIOtTNGkwDER4zoWB
ogXxTdMXbcYhhAm9Jju3tqq0hlv1tYfmarUoVOkrlACk1860fPKbVXSmE/9Iwb2OGblSNhi2WWyB
Yc4f7DrsMdmLIyh5uGKooTVd9q4UVCTe9t3mC5a3AxGUw46PbqBbh/RLjKU6zovxBOibPsX0XnCz
KxMzl2C7e0k01BN0pH1/31M0GmY88uYk/VHIHOPsXlAqeYG/owRbNQyoKiw9mhSwqKfDRdS7n9ur
jrBZPT/l/W4gwvUc5zNE4e9FjuCAtk2PVlKR1uenEM6wgjvEWcoTtQAoAO0+pqcuVW0qZ9ZRyw1P
KjIatpCDBeVSFkLIy8oBPDyMMkztP/CR2RzoTqLN3F0vQALtCZ/1KX+hjE0+4oaAVMv3iQ4V/5ni
+8L3jscBnnipoJDMlj3JAoDouPgQkGlFBgxTf8acEdcL7kLJTRmce59m5pwKszdNqtJUQH+HOOOT
iyc7IrMQq9KijW0bOerXDSwwijJUrMyydPTZB2nae6/a7lHCp2fV0/IJqzTnk2ycXr7PTIGhkvF6
ucWPAI/jgDfRKyt4OQbXQm4lU7PeZf3EKK0VfORnh9gN720/i+nWxhpMn9eaVA4RzVL0QPODmiCI
y4WB94Jga7jNfct0fyXPpJsllj4eMGkMajJOyTgc6HARHCPNmJp6lnaaK8mx4+AjAJVPm1EIrzer
lJi+Kl44PfIlD+uCTktrPrFPHREC8jWIekGx0YOmF0niF/8s1ptZGFqU4B6jcy9DDRY6lCfYd5Ub
ZrFYWMhdCDDvyYu3g6mVGVQoW9t9PuhKtXkNv8nOVZ3s54uo4DwfGqInbzvQ5MkMhMDJ3whsKtcL
JnPMHAZ38niV2ucHGFj06qRni14lzIiXZbBP2rvVeP+Gsv7GkLGWB6+PcoWd9KzmPjVZNaOaxcWv
7t79ooVAtXn/TDB0DYE+4bgij79ZYdn0PnmrayyEn3XxGRxtFn8kGX9AAHSg7ITFq7I5OYk8ZVqV
X0Ol1x0ElypQNns/XZYmUS4pp10tOWhfDg52ZjbG1Z0qjJ4bSrNWleKybrHPyHu66aaKBssdZTYf
GYLKGL32yTXz8Mihg0SxM2qYZ+C+VXuuiysUpKsmiyq7vhdxXUIjvWSNqiCrm1GyGFO8E5svpMLy
EVVyw0kPKYv4uxUy+QO5cGDlLrgzvjhloZpC5cIySMCHx5AcV6kLAtkurG+qS6wX2mZLc2NxPJQf
p2z48IA24dTuHsh1Ag+ZIBHC4vyTJcIc3HPQVyvCJeh+FMG1pCAYVqkBKfSA8t7znGY2RhH3uNxy
ozDMROGuiAvZMGfVigH0zuaoJdDgUVIpxTOUKVxPK9Mwhhy35tuLXf3AI35JCYe28vTYwmrDivTI
wfx6AMo8I1J0wYSEJysq6VYOkqf7661xAy0U1CSiFS+dg5qGhrqFVWxJtbTr+8vNonpXgZ0AveXi
8HGihdkVDbdjlSDWS1jMFdNzdFfj/ovnLOxcK0sAlGyr1naDmaDMVxurr+csbtjFI+B5xTpDrUeS
GkhsxTrNi5C589BlPUu787KrrlLHUM48SQwt3uE5Uo236E/cSwW2N9QYNNNo9vNrcY2UvKXdYCdS
W4Dv2SL9I0YXYNwO9T++Rgs8yASF7E2MVWg3ZmDyXyIwZlJ2vgy4vfuZVZ3Czed0HrzETAOd8uX4
s/OH4O4WZZi3Ox8Y5TBJW5QPcJ02kX7ep43/0pY/2TU7FTUa4d9ZhW8ACaFuW1e1WN5Q48fl/WSc
tnXtgWvtNigPYEJ5NSR4UHZTRZk1/3t6E8JY564vx2kLcfg28vVCrEYUr4HHBKvrR9JxG8a6fs9E
Uu9UrfOy4eRaO1O+VPhOo9wQDLJr+3Qh8b0QXbLCxyB3tWFVJ0UIJsk0C+xQylhBr/+GA52QUgi9
iGfXVCzB5QH9XOzt3WB2np7JERDXSmfJso1FmcBtk+PDMi/4jrVgFgWB1J9tFYR6MleJnySFUCmz
lI4w19LYdsMeiZNCuDcHOXfpZqlagZucZu5z7qlBdn2BqdA+qyOqyItz5kUsfdA43z6Xw0SITAuF
amLAn1jtcGV6tRmsdrnG0+oR+q9iqgM7on51SmVpUPEmEZ6PdBAc5IpMXvrVgN0ENYEyiVqjhVab
sOJTlzeyZk8NA+eDc/qEO65hqKwW5Oq80EALGVJPofSMSXq9z7KtvCyqdhI7wuYKXkX+WAvcIcvB
p+c0DCWhqfhX16KB2IR7gCEh0c4J39pkvVZKpzb1cBRoKgN5fpbcMr9ZiNJa4ZFdvLQhz41+DM64
Q4qjSzj0j57GeEWYZZQ7tmU3dZ+cVMsOwmR9IdyxEDkBc8M32Q7GweC+w0uTk1Wdc9T/Qasewdmb
ayYba+fRQ5e5ZnnlCg/+4IkX8uBV4TVHX8zwieellFEsqFQvxVUREFon+mxMl+LIn/YJywlZThfY
cEoK5tD/MQv6WI8ABgnzCy+bEX3iwQp50IgtrcpVkUJlhkiPEjFyKYTnaZSjP469BKe1Zme40AtK
xwp3brliIoAyZskqeObmbrhtrPc8u4Z1BJa9toy6CRNTBg/whfHdH2SiWIU81x1TWx5fNPKrXO/k
mTlas/kxwy8vJMBkNOnLNz5+J0o2gUxU2d8etfO21xH59P2M020Bb4QmZvpY+EIb8ZmyfpUVRlf3
6FYZ5JBPiMNqUPnvLQaRBQXTq+GNrViwDOHamHZ9XlJR4fLNQdBXOtfS+QNIa7bNCO3VrIAc06yO
1cw+Kty2cKfu1KS/gcXJYmi2KmwPnuP+xCEjCYNQGLKJqU849046iVkDDkwWvO2mm2vnpauEULmf
pRG8djrxPRggu5ttVS4YyD6hXZGyI/g++vw3ebmwDRPWp57uBzNu6b9Wd25bvHn5dtkkbKov26xL
jIwmhiqd4+aQt1ACddSXkTjcqhi89Y7BM3lbUI6K4W67vACeR4iGzUQq3H0rEi9t29IpiN2QfQda
57E7tgHjmWDUQJcXAdmvu2IuxqIjnbaJV6A+N3VtcXUHN+JY2HTEGSRNYRNbTViwcweo9hleGfEN
AE0iX5JxZ8JD36g74UrUReTW8bm2Wrq9jm1y4TPppz4l8VbnhMpZvDKF2/XnApPxVaDAZ7nftzvn
Uznc4Zuwq0wIs6fE8QLP6MaNVbwO6grDEkx+bDxpsTovzK03gcYb3b3+z177HhM5PImFmlxrwWP+
fp158Ldjd68cN5fJlNX2+CW2nxoLBspcGlaJmkoGX16cW7FVQI2trbs+jtlAhSs6gEW6aE8BSk+P
u0cxVrn6DusZEhKUwwwnkvHc8BeKQI6kaxtuGTH/BgdSZdcW2Oz/lyTkvCN8kj19Y/TLDMggmOmz
uSzdCWAh+ZHiAs7C7dMwh6yoPYIBJB/V5gDG/iivZuoutaNEqy3Qbryovf/fzGW2ggQrTqECBJ/m
jrLyqZjRm0BX6Iy/v0a73n0U7o+3J9mgK4vEPpriyXDe+4QUexvLPHLUSfrkbEPakVQF4rolfQ23
RqfFed9yvj2iPPVX1xReHxFxTZrwU6/n51lfFUxzlV/bN7e0DJHLcwE4YLD6pMiL2n+lJ+C64F6e
kpcq8XZ1Qm/DkUmzbo3aVrbyd0oPekSry7GSHv1+GR/eNIA8aY59ju2UKGTq7AxyzuQ/jMdY/isg
nQEMbFHsIwOba1HZtq9xzQl3ivcqsStnhabsy+QWA1SnpRea51MS20thdxw90iKhjpK+F5Q5kvcA
cRyXZPyR4OH6sHtaVXzzSM4BWQIAJ71H3Y1qEIAXuSKN4ocXbQeiQ1m6nf4n9hXJgBvTi21bO6Wr
OKTzD21ECFP49rR3NUUh3wDYHayrbxBarcAhGNlabEKRaKJg6RGuq9fz3Z1VWsu0IDZR72bJK6X8
BD0B8tdbJJlf497dHUfH3z2hDPPKIPM9N8Rsv8h5GvRmpIL0G7b2NjZeGP13aq6+yPe2Ob3OSSnQ
oV0iBwxRdoppKbvhOOroaQ5XdoaO4WM6yYjttx/58pTkKT42l6PBg/7i6+rceuSrNXhpcX3T7FPX
h6qVTAjuoJZ6UsJfVhpSupVUxj2uOiAL0FO/ECAZK8XhTdeQV/LXqibyPi5/4Cg+O3xt8TYx+2GF
TNeItIPl5MCwfF8plcOaAMs+bzktDBY73e9g3bW0wSlr+ifBqPt79Z0g94mKa/kkopsiDhCtVAhJ
ovIQPYhks8crX+4AAVmfOz5pzfpSRf0T5qD0HVv0tcxyXR8TzBkTFgTGy01JPyZMfTdZY4oClOj8
84iSNvlxkGPGZw9G/NQNysyoVr90Eb1Vi2zHxRelLbxgktQr9mqvvDBKs7ay+1uIYu6EQ313ewg7
sMecHPTU+8M8BkdA7wtRLujM3Q8XhBzcAUcgkw0JIcLv3x8faJCLEiy65hlUgl3lUAOSHLxBccMz
D6i85j+o5iBVVlSZtvbuLHs9CwhnSpKWIhpPN5bwbe9FYGgFPnxRvg1DJ8Eh3ns3Ll/YM6Jed4h3
LVfA3Z7gftDRzlSgHkwvRGDM3C5jQpeWR9slzKyF96+G+jinsrmNGC8kkKraVEP7pnrxMF8E/VMh
wi1ZPYLfwrN28SpWFRmfmCFgV0gKMjU3Cvpij+uKgwIMmu7jclzCqk7uezj5ojWVV8sHstbvD4c7
JURpqEZjNpQUdAUd837sKZuI0YaZyKS9C7DLDXdqYw3Vie4ziYS0WSFc5CQLOxfBzlkPxstxZLY9
tZoZxHrR8vbRt96FA4pCok2j/NHPEIvD5EPPPoNhnsMjAbqoQlXHeSNMsKPfmDr26LgL5xXKAVh4
aroiB3dXhmRFWHJceb85ksT4o7gKUDbAhDBVVgJpQsCnDYUgU1D+Y6Iu4EOeeMFKXbAZfaD8kq3+
kvMzFZ76VqyXVPdKyQ9eLsBFPYQGykILNYDJHK6ms0o3uIcdiaq1WexsJ/n1TkFfz51qynd/6gAK
EeoZ2hfo9iC/yATixug1h9oAX7sQUB3A6JRe+ID/+uCW0WYh1QOX6z4dFxLvU28Re7kdclytS3yf
13ps/yfq5jKgB4fisyaVWq+hVvz+gfVLPmFaIyCGuIQr2HX7eIelh6lGSulwKI1GBx0NEXwUIKQr
ddnh4kGRhgNCiWuShLMJ5jFi8YjI0T/2tqRT/lW2UKoeTAYS5CZGVdPht+XKKy7I97LUKDedAXSv
1pFsXCGHrjX5mZtVGSOd7WTN9NWHp2/h2sOA6tbuXYEQXwTXja7JH60VNYYtl0plB6822aFAjAHE
IkszjvupUi2uOFxjW9cLY/fsJvx9kj1yShWR08YnPna7T8RVCkTugX0B9iE1Ppy/MW4bhNZIxCNZ
bsc1XmejUSE7dSE1JwLEa7kDdOCcHtIIbb2RfwRWYCbTDMyomrgr3+ZS+ssxjH1wv11hezGb5bYw
LteL6R2yGnoPr5/0eayl+xQvEvWkf8hxAqHW8XOh6BsfQTxSW2si5i8Jj+6p/DFOAny92fuhxcIY
0Hj1SCdhx/MDPjO286juLPi8Lhzg3CLoXpsDXYMBXpxE8kEwXj0KSh1Vkd1FYK6Z6otfY8S8Rx04
UOdzJGcH37JC3La83e/TFeCJ4eDCZTPDCjJyZ4DFnRgTK8rIdHPr6e9nN2e0z+w4FontlAwvfyfh
QbQEVLhjezCwe3t++gBSHvMJM3Zy75X45iKSITWLI5q1pf0uWRWunh4YE1QzJvuqX2j1mFMit6XZ
Aidka2WWBz9B9edY+xe+5XnpeETfB7i66qYhq2F0PD9bBxeM/gRFN5KTHZpZix8335Eg4795HVYM
lgrkXltoEDqEiiKSXJtc8TPULysoNB+PsU73QSJNx4JECrlpHCZwMKBg4+uc4LAFE8NLsJI5pTLQ
ubM4X31m81evvw3UmuVswuWMo6M7LwXxog1I6W22L/EV991TRzqkUmARG4nyMn6tS6o7NN5bS12Q
N/UF19XFFlaWLyu24exR8+Ns1AH2CQRSgMN5P9V6u63QyH6MF4T0c08TdEtb+gR2y/QolnWesXzB
7Uw736XOhLWHory1RC54p3zCyk5O/5cKeYc63YKcSsijrPYM/0Ukd/TXC5TjkIMPnTx5WOOaF8ea
jJUfum/SbBKQiDUPNaJMSPm6YNlfHERvjx1F8enTSxqNAfaQdKxxIqBvJl+jUmDGUIJelaWEAu86
RrQSUH9HNRcLP8VPVqThzFiNZB05QDGok42lKooUdqKaFh8MswYRc4bee/7huOCL0G9wy1LoGyZR
Y2CJojR6mGtapMgEtPfH5SIWZ8mzIJqaI87HiupXyfv83+H+6fOQ0ZMGFNvkHF5su90fcRXdOOQG
XF1nMJ47YBdi+88GxTTvrTPRv9OePxkr00L2+wU5TRSQgUZ62lkZNKwbchkanvRb0Sck7cB/7SDG
Nnjq2gWJAF2ScjYf1j4/+RSskKmrigSq3Nzu2m6dLOLYZ3G3lJNpoEnmal1tP/atgfK0G/Msu8Ez
6ZuEOoYkYEAS/B7BFIs/0rqA8hPM+qXVhWqWs3jnfzO3S0N6PLlZzXAUA0d1SeUIIBxiDlC2Zwv8
doFTtsm7M6Q8MyHxqzY5wxny/o9EMABqhGPw74k8v2oF+AKU/VcaHfM9N3NRPtfXjT4WkA/C69g/
sMFuVxsnabVS1I+25Qv1m28UGjQqYvYd3khHMeh0KCWUz0UXXLPmE1RxCi5SgUj4Kw+Gn5QS7Nw4
FPqDDApiT668Ci8XXfGwnLxFoWoCumstO4Z2yv5m85cZ8rF+ovbv3rn3a5/Ul5YWDAmdwmFJvC8F
bT2WNgbcti2Qsiei08OHoLPmgrhj8okiMQjZObEEElPZF+6ZfCFRqJecFDYJGSxyef+NIMuaZLE6
5Gy3rojK4u92BNZCmGfYqGPZyKiiX6cO0jntuIHGcTlXEJUF5KZC9Ubuhq25rKcqxhlq81/tMmF9
8TeiLkK0SlOiOIYcxj2K4QiplmHj7oLaUw2h3LX5C72AGhECmwffnYP8C/yp8oWvEwFDLkN9gVAB
NtgQOK5KZzoGfUnx1a9Ii2hO1ZKMX3O57RgPiXshv1oUZXuTXE6I5C9oYkJ/dyagqXKhgmT/OfGr
rImLIwIJBF5JnRRXLqWuIpdgy3mRjw++RZGh0DMjZkm1ncVQI0XJ5E/YfMvvGiyyOJLD6AR8t3oC
4mNLHte95BFMPM+fBhKzSTf6ZZM+P+LpS/BwAA4ktRMXhMUCP61Bpiw3HGoFV0GAMLxnGta0UAYq
bHH7QPRg95OZhOCMviZPGKZXKuJCqQOppPr4tC/ZShisjy3xxM4YcS7+cWpzYIgcyeelLOAUHw5I
tpoCIg/iZbDLiNPaDds+tUHxZ9H+gc59IBS8UxBVfAiPoJHaoKLtAv4e/3eGmg/sN3hkdYhQsKXb
4vnDI/U6TnQO6e0RbNvQN8uER93A7Gi59FP+kDT9OyUdb7F4G/IOrnJW1e8TAAGFDilTdGarsh9I
5Ig7j6lWuXzVDD1ST7JXuddlqzUXvp/uXTqCT6/9Q3V5qhBYY+uktBMd0nPNuMo3lLmoTy8ENTus
NmhikOwnzTdhTEjviHevvnNWKW16E1mMKMkpTIbQ5QtA8pgIBtaPm277e3rtWAyF4dL1Q4lH5c+l
AAKKWXezDk5GNRYfoi5Vy/iqeCeZ5w1drA+NuaRovmBCIzw2jSfVQLPjDd86jDkuQBoNFVL7cgyG
jy8uVg8QXt9bSk4UJlkPcmKGyMKVfkjXya7rHh1ELYFffm4Wg4DZukSqbYmaiHZjQI/kd9qpoC7c
pPT+NNOaxWp6xvMqnhFpTn6rMUxvy1TtkHK8yvtMwwsyLASCUCndepH1Le3pTx8drE4foHyxImRd
EOdh9+VgeLBumcHH7KqQAKHsMEcnNBxQVzRNiu7p6CJyHSMu7UnEXC8yFPKULrSbg8VXy+AaZLp2
JjwO5lNehCXg+kME6u7qDqKnQMoCM9gkCTm3hJz59Ub62+L3iOvz5YlSKRyj4UG/lt1NVW1suGxp
OAP6VotXAje4NUQMfTayD4xJHsjO5rRfNczkBxWpQsvjB+wl3XvJZ+UhM8ANjCPN1hnlzz4E1Wbt
JW/0RewO2WVbzMLE+XR25eI112cTF/uIc1YO46Dk2WIsHaCnQCSVxqYa6MF1yjcEUychRHyB1jfg
eQ9tVrxyPqNSaRpmq+mFy8m5zWfsHkigbpRAB7U5Z4iyBJ7gXa3/tFULakPr0nUKOAHrGyxeYUOM
cbk3nXqv1nOuNwl2h2tLuuKq2dypBz3v5Y+GSi+bgPN98mSgXq8eA4MbW47uXVcq4BQjhJdjOvpL
LPpu7hxhPhye4R/2HKCUfBUjDZ/bvl5wyYqZZwd983X61+m7DrucEswxJV8RX4iXPxPZagRqwXxJ
PjvRG1XhjxsqA/5dbG7sLQBfPHPrAATMEBUX8RTLbfR3Sw73wWrNMGO18AxnCs57QpWx5rGA3gVj
A+bZSnSrpI/b/2BraGcEl9GRE6J2qOEhwSjputEReDhLu5efh2AM+jRkaSoKdyUKq00TRcn9+5Im
oaOUVPRwdS3QwEyFaZqpVyC5RM3GLKQuSDfl3xJVeaqaC1Vvxz9TsBplsJ+7y4sv/y0ofVZzIzqE
jGuNhomtxxEtzbfquB1+AvNmPLyGL70nUTed4yd6mg6m18ecKhR1BH6/QPFZpFw14+hgvGlkZ5GW
85WWSpORMK0eVqccsi9zq61gG4O5RIpyyaYxm/j7WGjNNnyaBFeqj85ozS2D4sPiTji2mPI9BpHd
cKMGHGUctSEokpTbBWBhU8EllBRqOJXGms8z3OUNer5ZLMGvjAd5vADvEoEKuivkTef5s/UaGmCH
KBDFDkdVbCC/DlBjs/cmkhbq7drDhjlA2/ZA49f9Fq3Ie2Z74KsMRDiktVryk953RZx1xuP+9IQr
WdBINSbDVurbzGYgHjPc2QcRger7PXgptIQ/E3rB2L3OvIL/P64yljjCQbJ1sNfrH1aAZeF2PNO1
Yeca2QFy8/JLK2Zadvy+1C6WFJMVFYMKpHQ0K19DNgn892Y/2OzKxXhxQVbaAcRnuR6opoWUfh9R
WugwhZdyF/4eBPn5W0qKucEEaIw3cWU9IXH7A5Pby9xpR0TlnsyJjtlBvaSmves0m3DfNzq+oR2q
juPRnLj24e5H2lqKrfxSTYbwpjcXMNQpe5Q0QJUvbX/i8X8Nqeh1/Y558uWjS39kW9fPuVMLRr2j
V26h+7aekNS1TUZxz7PIEM01UQP+j6IAepIGfyNNxusLgKVl4W2XaWtN1GGossZb996RUdgEElxS
NploNfZM8hgC3ZfXny9da4UCEXRbEgDwVBs4YCs8mk3TB2SUPU19WpGRKtiYpyvX4oIxNlXlmErb
/gsfT7zrqut5f/rYaoZsVYHjilrl65svcgt4Q2NOr+WBVf9cYdyncw1AaO5mnRoE3orodyd4iO45
zHHYMsKRMKqENv5lKxFAEXdxH1Qdo6EE8TQWUKH63+Lm96VMc0kAWnmSBj4kusj2PARvPirtInP1
P9r92r31BcLDTPHUZtoK01iS6QoY2j2hT3SUoF3o/AFkAe+l5z+91yS6TkkHX0niLcGcFOAykZab
0TA8MpxiriT9Ma8QDQeO2RyTedYHY8XGQ0BL1VzDigH1S6oa0O7y6EE69AhsDWpmme1ZuvPZ+fOQ
B2G6ND93pAJPOSeW878u9ZpQbb6VNma2EBkMAJIhNMw1KBNgNMssVEatSokJVUhP+J0i6BR8McWs
7+1BB+PWgnuUQD3jo4o2lIeOBKCnzzhoOir7Ce82W6bsIoEjSXyF0E/NChvOmaYUBs6GINHMVIkH
eAewOijEVjczj0asBx8c38ktdg80fibgY0523G2epqPZH0/1xb3g9QqUTXTJuNsAcpwa7WcwskmD
yyC2XMyddgadJxfEyDuSgLyRU+8zZ7v/FpAgtTPn5H9HbnnraNrmBl2wMC+2VWCKY0UZrPSlq3xd
NFOXO5Dav7AzJMhGGVjPzi1GtYrCy8GZSo+wb6xHd3sPEFznD4MXr6P4fGbCzf4uwbXOHQuY40Zc
7KKqKjTp9j60ysK7uM1hk0HswnfnW+g8ez3VDqkBQrkIk0kP/QFIoroA7xHtmsxgHDipdIiawZPv
Dhj/g63feirEaTykvCAId0IS6ap3GspZgwFJsiac3nyaoKCYZuOhhBwvQcun7cQ8l4BeolbKiT+R
aAL84boPsxBf+g5K/SmYtORhREBrZTSW/6OwruAUk7qzZ9EFC+ZOkDwPILRfXkKqzxFM1YcEaMoU
LM8/wuKnf1S031j2TGUmXUIZtz9IdKRjHQbhGLhALpdUew40UfySa/czC2rlCWoDUzgwK9i7lWek
L6N6Ao3300n6N0FgfPALZW3g/4CxcKVMyDqpFOI6TP62742iajUb/3yX5un3StC2VPjZqsTlk7dV
V06cJpNf7cPvqlEOL0UeSNn0v8ZhGLhsTlAv1mFwmy+Un2VIPs4xHl74poiJYKfIVP0lUpuTrORS
mY5ZGAa8270Gy/Z26knDa/5Lx476fPM91aL+mQ9IvXcUCBj5iWepJPMoCZeyx7dtg9AduoKx63KE
7JsOGINa4+3At/UgudDazX602zysBBGesXBkxHKISJZxpHjyu35ltWE+RpYAANdTD+FZ/AcqZEvN
IlTzw0J22TkuuapTYdpg/Xh5cDWkwMCUFz31G7wri82VyNptXzBKQ13nqkJJVxd5wNtjURZOXl+7
PmGG9PY78wIj/9ut1lbykOBa82K7zydJFvUYa53Q/SBQiDadVPUace1x9zdFqtOa1nClQNEGnplC
YYxRyz/aw/CAe9NnVA3JUpu0vF0HlWAXcH9zuJt7nBigFqaggMp0bTGOxAt6dxB1V2Qrd/MRcIlP
dyeR2iD1k5rYQOYBEAQVTe9/rofDr4qhDw1ZFi9PicVHRyOHI7jRGhNQMC2GI5R93+LOqwb37dis
IOd5zNnVkvwcT0CVppgsnf7SWhFM3aJHpkiD/doegYhvnvEe1u2CjYn+piXsg1wif+Hft5YutJUm
GBZPVqD44LPVwlW0Jx9nbXPmfgnoUNTYyniJdMb4EOYENUzw0qCHsD8K9Z6VaAcZj2iGjo0iILgx
JI0uDcCBBbSFEb/dx6f9R/obsLKT7sUEbNjRHl37URAhQH8XkHDjvSjoZAtIJdB6i7T6wArpBCCE
Ip88QamI/IQEKcNBOW+L436AwYtUdxlHjtaDQovXJv5BY3kc+iAa59P1tjqvqmFSZJm6UkMBgTAF
nl6i4sGrWv98KH08xRwsGHxZ/8P2F4BH02pB9h4/KVIqOISWdaDuTk/I8CdxzxQlq8Qc2I5sa/4O
7qXL+1Kx+awZoh56EK8LCjIE9N03LpHq628GYXJYf++uT/jEiOHw3DLLxn4ltlKbG7xlLW8E+vCO
1mzgZ5NebqdhydlIU9tOMY2Gh65ukYDoxFCGsXoRFrQacKFeGphb/0jZ8XNrnvHVeXVo/1tBNhMK
O2Me9g2YRAZfXNqtewkiyUD6+k4B3oyB2jgsDYDX10RCAMXNCq31Ar0F+Qrl4Zi3uFvCVCcPHSei
cLUTOIk2p/9gTxZP5jqpQenkd4FOIDxa9NLnka1ty3c5iEYCHgtqsCK7kD/A359p0OZv3Lgo+01B
EC/fi/Y/WOqbnlXRuKEFl/JTxDUBdpOzMbD6GdFGwMyUzFOiqJA2gVsXS5bJyKLXyaXtwaaGOGjs
1gXyJMf5/pwRNyRe0s4o1/Bn1sjeR2OQjAHmVkX72tKngnzXzMOl+tJD5MfimgRlYv9GY+FVMNVh
39wBBU2cMnugwQYE9qMS/Hk4zDyiDM2XP2zUUW8BBk0qUub0loDJ9i3gp3aZLeUb4iEeEISWCl3d
0a19SUUtyGyUhDMZgdFGNwxLPVAV0j7NT8GuRRF4bWvofF4D1NFUZHzDfe3c6H4/GY4joLl+X+yx
temm4W/nTe1QXbIJd/sqMv74nX+Kivqq7G5vox9oaXeXdCNu4ylRP5hiawv6iu9bvqPPPHvastCQ
6OzVrN8vwNK40bL6nPOCpgW9CyFgiR2xI8ZX4UCqK0SWz77/+Pva5ZQymy9LAEEJ5AAkDCykIhdD
RKPCQFQbsNeVXhIDGLYlj5oin3rXm2ySMOvDxA0tjgdOcxwi9KB5+CHa/3my5M2mvjeS5BHAElPf
PECWp5nv0peqojDaXCAbv145YPvdCV0nlmQIQ9SEztMIOg3ulBLtEqJ9YjF+ti9TuguaUkXp4USw
ZsNpJAotGMsKHZWmEskck/4/63Xtd2EV8yY86p1BwIGhhjIiKV8I1VH2x+RHvJ5fgWOTWKE4GlDE
GZV3hywIh+0CuMA6yWg+YgOOCreCsLYOljrcF+315CQ2eXrrDz6ZBeeVqsZRIevnY3NwKzojxGa0
tx5NxMGKxEq4YhsLs+KowKjQ7cWI+tyahgf/FSQyj6QTnn/dPUOJ03YqdhYg3PFmKJuP13lVPWpG
iRcayfZXyxoeU/KawNPpZi1mahFUOgvDm9y/c2VG61f46la4jy/JkCL850cRQfGs2Acxd8WeX8mb
5C0Ri1Agg2ivoejfaIax8Hgiwd9mFBnly4i54M+TamrkIkiGU/iN5LRFHjv804f144MGNudS2RsM
4xsRmcRib8+/3FU8mfeBj3TU8EqhJd/JhFB4Ii58b+nnaoWtijpywAUkFOxleJaVdE8SDmDTu714
ujhevvmsAz3Ye5YQ5yD2LgBAhTfU3nwtGlnHMZ8EYG/ttXGtY4A/daijpcWvpdbZIuMY31MlzoTI
6DgJyZfaWhpWE6z7bxux4moig2VHJxsehxL/zL6Z/tuRkwTVKRCow4M3TR0rBd6thmR349qhIbqb
BFHYYOahsvzN90dDkxEZONpnnnLg6+x59n6QahNxqr6vT+Fo27wPiEqc6BbffWwd9Tix2O2MJcjJ
YTaO09N4D53a3PmDQEJAQDdd0QfP+iegwmQN8riB+ZNOWAibJrNBVDCLgMNxESY8emKSGqzSDmIR
BjjqKFeHApDzSethK+F9MdjneSMBSKJ3cL76zcpPnJwMVUvRxoBHftaFh2qQ/g27BdbQnXlNn96O
B1EmrFZuBvVcdXLLwbrUUX1tc08IHCSVKXAQ49sEJHSePGfzhTFMcNM5lslzPUiSHLXuDAdBWqL/
Y3N/d+k2KTgFscVX5RCEh3n1fRN+zZYpDSAUbggdwvsfw6/n3PkcMolIeTME5Z/sq3OOklNAPb8G
qPk1OP/iRT47kXlCN69LOXtrbnH+arLvn2e3nM6jur1cux/5C/uFHPiP1BzCGOfx1gvSeS8R3UuF
3KMWfCVzzaLmCzA5ekNrt6b8fdux+t2i2Ej9f/Iy1lRvgvQ2nsqj6z5p8Y51OujBfRNwAZWK8/kK
M0OJ+RxJQBoJOMTev1XOmfYISt1PPWZv+EtUxmG+qRpW+ksERUotIsZA/imCV61ySkI2Sm8yBFPH
Af07ZBT6d7mhocLYsf5cTWzGBX7HJ1RBX5vBx0OHLCe76RIcON+xuZO2WiRN2xdNzywvmr5r3k6t
xrfddthks4drG9VH+quVe/mrr7IpUPIBdeGI6lgrA9ASCZn8XTino9Gd8bDndoosYnzP1GmGiT0q
kg6+erbFWM6NFJ8dS2ei9PTOUGZ1nbPNmK1IgMSWdWE6DngoNh2Yx9gWgqWiQriN74Opm1iuzFtE
vP4LjEHRuPxdncFnZ0w0S4bU+fxZAr/kQam4p3fWirCJaLz8VtSqfa4tiSagUH9iyCOlxEtiVjHc
TXYVUjPJ4fq5m2hUI2gonV0OZq4A6ZD1wVlb+riHiONk3NFsf6+SPUf7X+WHcPbQSnKokXmN3cE4
xBr9XTwh3im+kJaljf2Dy1kF/6rqJmmI3GYZ/EDETpXvRP4poDQxKG5H0ZyLsm+uxWEEA7SaLBs8
/ypFfQxqxTbBRtNreu0ENVDFYQp9d7ilWnvquAEvKKmG6CPhdTL9zSTgAjWVxwxoORFIfYjmiR3U
E9yg0a5S2RmH8su85WtwInFvrTceMDcDMv6mCnjlNcoGMlon3gTYR5Kqkg5QrZceq0DjhExOEVI7
WEeUo3uxD9GEVJFb8bG5zruZbsCg/dFrlBi2GCnjitEM3Fzp+P8wDXIXcqfn08vvFRBi267rFix/
11xYr4YRGlMMQ59V2dFdoFUj4F4YsfQ0qyBHbPP5W/WCzPE5weiNhTRSDcmkECuu2mFInZ021W0g
PemTZbUI9kocu2P970OGohXJPW8p+d0MM5fm5Y+3GbZKMmpJkEXxBTCGEXdjMLqj+ztnZmvKwOBb
MB7GIo3yvE9DSCLcOqo/EGwOezus9jhympBIabzdUpTgvK99bq9iORBagINCoFzoNJpKXgiHgT5M
DRKY/GML/zgpFpF3El5w1edeXhCr53pVve/mbxg3wf7MIvwPhEDUlbHoSgw1dVJ7+9ArvHmqJjvM
tMMzH4lihy4xgteoAtj3IcMVTbfG+PUi0rv+bRBFWgREFZ7owTXWVlfiFp1lz8bRWVHAa1XETIv6
g7xixyvWoMgXOiiMGNLozKsW0+zWjki5cFTvyYXdL+k8Nc65DBbiZx4OBgQcU8YbRLP/pW3Aerph
Fs3FVcV93E762Ry2yiW+bsMCLKsTNh1URAfd5vQH2n862l/eWNR2d5F5za3mwi1fyH052e2Xw+tF
ZfqsQTULyy489RYmNC4P6VeIeGGgVXL5OqtMeRlP5J6O2SoKcVsVr7zjbaBNdXyEEJHslDmTypib
Qyq3pRXe8viNuI+e2BTbbK0Q0GEYc7sS/2epRMPmJ8QipoUDn0FvuwSF4SXZRbIpzOBNkDiaWfUp
MQ1LBy0K8e8RIO3AmnLEUre4ThrTODCEQzoR91e3IemhD8fi+RnGo2NnpuVPyKcW0LmULctsneVr
q6uqykrdfGFMg5uAlK2azGmZxvlzpEbwW2IDhDoOoy3t/e5+LCcAiOopsSR4HZKmOi/yM5ROGs3v
gzkwbNHaUyy8wzPmz+udi3Sa0vwzU+MYnnEPeDkBrpRlJ5u7bMIyIsgdIUa0baJCVyACM9C8gXlS
+JwYL8qpq85wvgQOafa8/t9RpiHG7CtJXoFk/3wbhQ1/s8RHw6uy/9Xbt2akbUOjMPycX5U2HI2h
UEAGkTTUf8cIi2vwTvzJUr3Z5fE98J+ouGERkRNLyJlimlVi2ZjdZDalXfKHdZcQ+G94Hq7gY7q9
v/OYfDTPnIsVUK/LNYuefgLc4MXjNlgd959UaZIRzoDhwkntL0G9pbVmLjz//5P6aGLB1AFQEqu8
Rt78xfUCI4SnVMjTE1ULQwTRLrE6gXlR9EvWTwe+SxSl7cUoOEjvgY2swRI80sYWBN9N8YLGyWPR
pv/t9HsNuBclzVNrwIEefVpbXG1KczVGsQ8SkwFJ0AA4iXiXtcm5PcYWlOh0ACwgRn4d0Sjb3vOB
vLNyztCuIo1xc1CtoYi66GQhFW2udFY6OpL/RkFPSXcfOymD173A/1PdzgDWf0ov/77Jt9OX2+/b
4+GIhl1h1Ge8JZHs0DfgARhRAaMVT55HJFaepTZw1ZvKPhmme+D3lXhe1Jlyzl+mlme9nV87H0eb
doNJYguswgghtdj0P0PrIINzi9xkJATrttU7Rtto98kFtpYSLNSL+T0ssMOh2wU/4yr1JUtD9qtE
B6CmT1Qo0pb/Ct04u6KRPtl1ohvWDusLxAU2EWIHEFquoL7UDOV4T1sS5y3XuX/kc9CFe56xgHpy
YCqGLGcHM++1ah0lknvTO+BkO1Mf/eyPzaDdmMOKV/MW08Ah3YCKvZz4etCN06PEt5Mt+2Y04bKt
IqcObkIkG9lKLXQZI/wByUHFIRLXkqdANDj1lkbkgYAZi/QZOB7t8qIkeg70t3lqI+8+ezfVeb3C
UhbCjKzvSODxjpC/VPLtY+lsq5sGe9Kq6K01svR2QWB9GxrIZ4wNaMapH+4vUXZKmM+mfB6uvOMY
njS/Qjzbtqhq0eWfEO+Sc16tfkVzaZtMJmkF817D4TaQRMqNKIBf8AJwKAVAdnxs43BXTmxGUlyv
1mIbJok+/GdCTAYdKBNtl2nnt9p+ddeNPKOvD6IETuf2kCsWADKI8U5OKE1IfBguTuQ+HZUf4zCQ
F9mnB+cez5VJuH4IOhqjP26chF0M6ioxsI/ffVZtuOFAPaLhX7ebAOYh0lhk4YL1iTNlxOf13s7V
9vWGojsfKItdSmT1RR5GKIKQqKcKLDbspka9vRTHz7IRTXS28cfkePPra80MzPGsSTd9ufrV3hyT
d3rk2ouBoHdLPxRj7ivUIuIQgBYpwAjDxojGExHVh2uCtbH8+w0OcCDyvPDg6xKeQGyr00WmVC6q
6g3V+OT4iRwrdt/m3Lnt4GQ7D2lLPPXKwutwMD3dqqOWUcaHOkvNBeTt+8yuZKLSIsYJyoLEH7NK
GzwKI1am0w7cMe1GCU/2CTK7JqcIKVJT81phdNOIlr3/DQPi0KHjix6isOHEIc5OdVZgj8h2S5Bs
jIyHA8AlPs1gI3wAVvs4LrWIPaJk062ShwTCOsaBD2z7E6CoquW4AhIlQN6RqsKo0MYcE97ifWDX
Iz0m7DsWTFKeK+vnpX0YdTASN7thqutaPGgARzG0SKELkv5W3L331bMLqTyTDiYc39E+UfKNgv1V
HJrookYHsaBvSAZxTM1WHXbO4YY1yJn2K70T5emvWBUwUNLUkpcmgjGkkJKEUSp3fdRI/Jc0zbiz
Y2sh+dnIyW9n7YA9jjgPNRPpTNqt7mwqOPMwNp0P4z5dZb2XXIhfwJBk9ufHa3TDEWJRyeNRC2y6
Xys+nBhB9nlN/HZZRurxlza/Powz8mElLPabqtRAsfT/rPVJC7vNzv1/A8pZstjEgfq1glP8mV6Y
L5lZ3bZ7d1w2yOTYdJ22Lavp7+N5nmmyrQ4iWEh3LT/VbGzFm10NT8KROOOt7zm12C/XUUK74T7F
l7jYimRZl6A0nyVphAYncR15ZB5S9fkJZ4L5Gy8FDXCcEsF+6hpUIZzXBmZFBw2lXbG+JoMGIB5/
ge1HowKpYBpYbpfG9TAd/JEl3Lujhwy1objplylIN9UqAi0SrE8wgk9IBpPSoOLsDl7GJDwNuUUc
KkJlDIcZP6cVLW/rXR7Qdyj7TsWf8Es1ZuzAtMRNq2R+tGNbA8O7XAMGvpjskiefaZG3SUe2V6VB
EMmKAg5+S4JVikh8ncy7HBdLpDs0JVZ73HeEeK+7DLzAt4YYCzZamv+DIuzaC1hHUhZsnsrE3ZbV
xTI0eqVra4ZrmYJD2QgJUPN+p58oOxZ8zCv/oZkH/T9QlZNHv0KIM1t+b/HkQb+hZS9vqmPumwut
z3LLJ7oI939GYknwNKe8b3qhASdEds2tqGI+/LL4IG7NNyOgODUjO1yG5hGwJwZY9aLc29e3sx1N
prMbAKc/KxhRdQnyXV7fhT/LdFKsJiPo9Imtjl8u7qSCS489W9pz1B0RHNzvqY5YAaNAl191s6WU
XI/TYlcB19nuDVl8z0NTedEtZkgKusd3sBK1Nx+IrvP3/zqUGdqPCK04FkvqSDJWaPX4FVWsYOOC
CtQ5uo7KEvfb49ywxSZhJUwkdsViL0LOBXxZLnQpNieDyENrmpGZYcS59WBxlceqCcyRGgN+gJLT
zN1AgGPT7tbM1jHF8jkaMLE5EYBw48ZJLDeq4YdP3SpX4xmBrFS5iazaxPJQNLtfMbR3m2NvhhDK
ak8doUF/1u84C1d1yIbpayWUVyQRfxRyqR25IczclpEAzJuxOVgihSCPgC/FboaRbzr1O/QLLMkn
yJ30nj0sHVt2mSBa+hv6WFrIs54Wi9iH8zE0pJh8oVViZ+ddPTLupmSOaoE/gYN9gPRCJHFZGKkn
DD7tnVlTDYcop26ciX6fDEoRPBe7fVigahApyN69YD5ouvoaaDTbBimJLfKyVFZE66pAqQiEgvwt
Nerz6S7IhPJP12Qw6UzuOqyW1vQuYLDuNNyirWVkr4cegowsARLADKdlYuOt+tdzkTTywuj5mXqK
ng1ix1w3pOSCC5wDv1x4FOw7KZfK68k0sF1fOx7HKK9kb5Bb34DKwvFwuL0lHZNau257kPz90vp/
OUYgwlR3vU1c2HAPuL3Fkg7fZm9YLnRel0ZaYsP3ZBuaq6H2iXbI6T6YbzBgLKowXnzRuKhs3V3V
NDMFRdQUMluQPQjWrBNpk9cAA3vECmB0wx5AKeNTXUw0h32OBvnlYvOtKTks7fntehOHIR5lX3TA
J0tE6IxlGn5TEnYhP2pkaZ+eUjqdUwucfXwt92dwK3ARtpa0tNfkBK5WSCxDJunCrAv8H5hu9j8/
RUBGMsdFGd7yClxJy7MonJF8CC/xFIB6tjT6kukye59OEtfzDAGo0fXKDEVm1AcOR/gI110d2PME
HMrWnN41UiVWD9D+kONJNVsrchkVt1oCUFeFOAeqwMQa3dZrIhqwzApQnb90vcU6MNeuJXhSb6Gn
7LmhP3z8UtU8u+XImrBVDICFSMOwh7Vjuf20eBVIy626DdusKFPtD6V4UXmUJrLaxUnwRaocM+i8
0Vsu55NPOJ7Hli5LnKQA6biRYEaZWntdVUNMsf88syl5ui4Ac0ckQNXRRYY/Wnd/IEs1Ov60QLm5
lgJ/pNDgsSFkIS1Uk80G269zd8hT2KotLvH4gHmfCJ6/YEsp5jzYMVafVFli3FEBOit0T1+eNP2Q
vg87RkGJj1ZHqfZhW8WnafomzZJR1aW9nVSHeaNZd9YdgK31/Nd9NIIX+OMDYoEwVERo0QStsfkX
ijy04jzqyafUG1Q/DL9M6rhWqk4Uqzjx8GOH6IOYSj6RdUw3LhFSTrI/pmVk+Be0E4Qegl7Tsy7n
wKQzWodhADQGk5yPr5sJjQQ46WrzQJNEQm12okRRO5YAaLLL+8+q7wIuozq8x/QMDl0qokdCsXYc
SDDygvspjxgF7ZNtfRlCbI12WrVVmKnaU7UcjfvC2ropX6gihArjUcI1Q/yeqD3XnlftrHURLMsb
nDr7yKgErcwkm+TrD4z8dTtYgEw2Ofqpoc1loBG6joby5Cma5MEMQDfpiHd6EZ4ZTuhFJHlYF5m/
kBCe7RALtPiDrUycA7FXUmD2e5wJQBN8NHS7lZ3CpH3/bQt6dTynstwoPAl9XVf0tq5h39G3dqEV
A9GqYSk5ZGWOKjyePpJ3YssHuj0chWuc+F/Mboz/JeGsvrtp62Bpbd35HHsa+P0PHiDiGgvCl3mY
u5NuczQJLMatvEp8tC5+vT8AnGpG09Df0v1PlBWUaFY0eRsoFUYe36Ud9nddY8YA0T5XqF6okR4m
4SZUp5pvS5aWRW7ir/NLbCYaw1mYDXyMasA8ym/sjxbmnuObc6vRhQkte9vZsOIHXZM69Xfr8BUn
lzmP/BXxwslrYniKQ9r1VnKaMVqQ8V/0vCJYnrZDlaDg/FfIIqz8FDS322HqulPlLoZHTIEn8ff0
giumNPh0Z5fY1CoIHlZekrkBv8GCR2XBloE5To7nqf7sQ83WWPrburbc6FKop/GfwGir+9dXuyWZ
XLy3pooPR3ke3+Pl0B/15mCUCEginzEoz6N7SYFBKm3/Qq3UQG3VK27Olq/zfVRUFPOabngTmxDj
LnBheBNaGmACriYfygcc4/Ys/ahC2B8E4MTqu8E23e9ISVIov4Px4dhtWS0RQj4rFYKGbeYdtA4g
rK8ghGp+kpo3g3wCGqyPF+EySkKsnsCr3uxesgunQ4VKN6yUVDSs3XSR1VjwUB2i17RnVFL8AbTu
/mkfI0DJvUO5PiFx5WTkN11dYQAdHNAAUXmGabO1FtRPzoXI+aOy7xeaxG0yHDZkNRrt0dOSwRFX
Hu1O1mbLlzOka9wmco+tTHZDPsiB3+da4LaOHMq0wDytynbNlimYO39MTopj9uNZ8ndQ3YNWqdPk
cOrJC3h2KzSTIWCBUAdvHW2wmDsUhuDS01l82/a5GZhr3GQSwzsgv0BPJuNcQx/XThmJOqKSK9oT
V4Cwb6d/F8nlStSV95Qm1PyIC5Lkt3EarF8rrz5rFWWg5qNTIngTJVwDMu2OB6GncGvbqCTEhgM8
6lsnlVl2qcfxextLIZbDm4jiNeRcCqXP9jOujrYaau2dKzJnPgWF8ddosYB1MlLmGE+rbI5gyLQK
sYep5in/ey/Iq5IxyaGUqaOmmDSbD32ywKimg7rxmx2PeSBPjYAifEr1/L924f+WrXbE2HVJisN6
vEeLyo+wUKx5ggrA1/eixytGuI2K5uFLHsdPWBhymDgc6JhilOYYoGgcZuJ764PBDMG9imq9L75b
IOWlrTjA+81zF5hC6fcP6ohezoUEtNHviou10NzmujDQmsPnXJfK4BHj7RMmh/4FYTdZBx+zesy5
8zGCxoHX20vwx6zzvMkzElXGw7ENJPPWiNAjk2uQFS5E/aiYN6aWABxF6BYVpL9BBZJqf+7wArkH
kIj2VAfgy3ZMU6qTK0ZQVzjfa5FhqqU4EbACio9zGiy0A9LLYnWfXBCpE2VR015OS9Te+1aXwTfW
SkPSXjpETnLbh9OvhJa1DEgftcJJjQfuJCrLJqsk3euJHwYbLjPHeNFs3e35ChDdlXRyHBw8vw/a
nJklQ5iYpSKyvCe3ztzX2volmcRvyTk33DGN4JQZAnD7E3kov0TDNAgjhDwm7BcecEKBncUgm/tF
WCa4ngZQEDHa4qXldRi38MMeolnFvv6ij32ChLjCRH3VahCYhmJ9P5LQ6jLZH4ocC774PrZKhY3m
UHPw2oFaSN0fSvvca5EjOu3MeXZw//IBHX+vUNHOTxUlgnpnTFmXqkqcpBozgiX5QrDFfa7fjl20
f4ikfuoG5qiVdJn7QB0NesAEjntca22XdQ4OfXe2Rl9EQSImdz96jiVMQ9ulBzbADBKGTpxI/UaO
soUtzG9DKSboWGdwNrQ9Pu/JirR+X5e33VeptvmPzHcgSfKl3rJYrFmSLrkDy7mcx9PGygqq/aIW
m36TwIpcMzQSDkXL13l52y4Om2NCrZpjbZSZrRigcI3dGvpMOqpgl4DUysYkoj2qQDbGn6bQTbj1
G+Ilz2xi+Ol9TpQXVwDluElCzHS7rCbWUPjJBIQ5R14PStJUaD5ICyPgXBEd62s56/62+4cumbX+
db6NhUB4Cjrl0qkCl8guANUFnko1xO2Cs+X04LEYhJEVY96cCnp6LktooEAl8w08+lnLXtv+ZMue
oqtnwACYmrDACNQ5T7SvPAVkXrYB4ID0gwh4SMV/FCCrRBlyZM4iU1fP4jIbFLdHsufaqLKlelBn
FYsRC4d/qhq0TEzA/wyqN7S743nZnNAUuO0RYsgrXJswb19ImQJevxn7OEnqu/wLwOtt/fhPsn/l
B5CIQ0bUY99HIfAEKBcegzsDti4QqO6BpbOx6HI0Xhdm+DPz10iDn8Q4tWNFxJygn6qO8if56gP9
H6CV7msxUABVUGTo6ayxGvvNJ8JviWWRp1FeYxdNKGAeMzXypiAufVmW/mctAjIhlFWCobKrXfo4
5sWBI/Af+S1Ta46VZSG1LbZ4/bXTzP+DpMVG7itwrmUWnPS4BOJ8EJjgV2rd1u2nDfo9bv9qsFcB
EfrXVC+rjmYfZj/QZtebKBhiPGE/Q6kR1eY/JLFH2ou04tsx6W7lXareU3hmc9KpqigkzHoxTCsj
3DtKP6Zfmy1+ZKNZrTp7ZNwT+AnNug2qcVNW+ChjBElpS4x+qx+oZAYXJJ8r1ZlfWp0S/AT6km8h
dIdu6jioVF47QDWKyj6fNUj6OxNA20++mypfyTTYqS1Dm4RuVyFKeS4pIyhAGy4WiQ80C3BNgMkF
ubNj7Ze913HaPEaNmTlk3SblI8NxAeO4R2OuUxNOoenDODZV3L04FMQ99HcDIRgWXt/eEt6P5DoI
U1T3XDl8a55e3UeXd7H2Z5YAglYORmtTtR1zDdo9X4SIssG30/WqxO5n4TmpT+Fmh0UwD2VBevFV
hHCCFsWgzrpdBz9R2qNbjyuOi+Oa+pZAzF6q9oV+FOHNxcIj7i/Bslk6z4sC4s8En11SHmm3j/Tk
cuBWLxd4F7S77iU9X7hSr9JUPZFf5Z87neFLZJfR8LHE0BB8ovAKFuFgSEkxSMn5m75B9XXEOftK
JAelruIN0QzT0KVF+x02lGFFvjJMu88RvPd+gWWf3tfe/L/CraSAyRVf3DDyjejC0Je9FrMv1obX
JKrgDDVDD5HuLrBhNPudlwKN9ZGFWZyrwqYjyu0oL5GxC+ct7KmEQH9d1d5S70gjyY6MW4Hmn/P8
qAp0Nqt4ee/nGrHFcosJHYOG/A/OV2H4LyVoUOTGblS6Ky5xKaDYjEuOk/MaO4QufNafvGRLNG0Z
zOpcoEoSaexTINcd5ahbLtbfWaD+eIicTtWpH0T8irOG3pMDci/9r4Xtv3wZjAw5YoqL0F734fwi
GD4DuwTyliJkZUNkGQ5Rf19JTnHb8Lt4J8I8u8U/+BOXZziuYN7HV0c08I/s2+/ExjbqQHp5KoCU
Z2JxyKOfzCVy+hFSCXjHV9Actw5Vx0TADh4zBZR2pWPNOT9uLaUyqzQzdh/h0JVUWdoRP5AENuKB
FvrSIlnoStSOgAPmraSD+pQif2i+6iIs4cpLsHOkfgfR0YvozmmXw+z01RM/G0aqxX9OZHWOK7G3
gMh4qZC12AzIi2uAdWGoaeZq8WKSD/PY/qZ4zAbwj8r6plXaoC/0WkK6nCPq23+rcddmX6E0QtlB
+zeCS3QSn3Skde3ipR6S8817hnqPpS9snbDFZutFP6/CazrU4smEasTamTh+Sif95G5ErjBbmm6L
ljuep2zZCt6gAlQPrJH8g/4WNsxU7uw5S+Mwa9XYoHX4SEf5681an4xIbOwOULI55/HjH4yr6UcJ
AOygjHmUI7c56nXtwVw5m4Kmi71VonFJwDWSFG+GPDJmlBt7SXdqp0P+n6i0E0MsJpGPPsG+0vMJ
TDtdfnouum9417JLfRvQYn4HMciTwHYG+6R+3/07LDxmdeTOvAyVvOfMkS7haP5+82nPtryUnA6S
SokYKptkRFHFUTHbCyliTbRBpgAWWzC8TF3bvOUNkHrdwUByUALeMesjvIBOw3OEZw7RrXR7h0DT
bVO0+qAT28wMLdDl63yOSOY0NoUArtqg258zdJTauFTBtu7nlhqYVY2JtiW5hek9ca3kdzcSVoZL
zwvr2OX1rZnYHFTw8B4MJ3C7/tKV57GH7d8ox8zHKr5U9thxfWmjqXaz0qi95xBUtPwiZENQ/v2k
7VAmxHr6tBP8dfG+07I6ZhQPh+bGHC7Nklj0tvGdz4CE5t1dDxcEqgntfm1a63pOxjq+zgh5iO86
9Lz6/NJZ44AHXAvcQsNO0g50ioWMays62GGgfvCvMI8/kjSl9y134NnpXnOq+2Uu6XW47xat5Rsi
tBhD1XxyLnCPXmXUv0UrkCg6qwC60wrDDW6nKL5Az5WRUIPlCT4UipBmNTq6AXbZBrRQGgTzasMi
4/i2sXP2cHkxOW+E5O6KHmSqz7D6V56eXrMBUg3TkBVomI+renP234S8mQuWGqIYN8MRtLIbnyCg
mqcj4Ry0F+nBXBjb+LyH2SL8paXI1LCRMIH42ubfGQTmavJge+lm1KbdI6T3lQqppCPpFjeAzCgY
10Uh6De5defQGVKWCEaM8DX87910yy4AvywoFEj3FjTnwiDwO5CpG90nBug08APCIyPhU/p95oGd
IrTvJNBNzAVWtaKc3fIyox77GHFOmA9jJTpAVrlsK8q6WKJdz3f3lgYY3st7SAgtDIyEwkmaoQrV
17n5JRUcUmdq8sPrFnw5mzZptWr2IWGW71IydsDy3nUueSmr6t9xVo8L2aNKKioiLd5599kyLTV8
TehXHy7WJ6Snbvjgri0x7nF+0hWnx37s/yafo5s8Hpkf/VgWmVeA8Qd8rGLxJzjV5Ok1ViCssLAE
M/tNU3Air7pU2fiTmofbf0UD9jj5u+F8NTgPjQlrTNGe+/av3wLLupNuVGT2Koy3ekCB/MT+w3R7
U5rpK01ZRd3+30VAZjHrtPvL9Mcz0vlwQ1XRk5Qnq+tBOTUtRtMKKsY9CNoTXepnHLy/nCCrzx0Q
miJNkaUu0rnZMK/M47+sYYuwCMV4h4s4cddw64cEhEmtzJGNli5Kswpypud2GK1G65VHcvkB9e4e
MDN4ZObXnFU5W5jfdxx+JXm0rGouttR1CQWqFTk4vdJveQAVDeENc7M3RSJlOeMgU/iULcmNdi3y
8h/yd8R/5QG+GO7aahLc7o90t3DbxOomL5rThs1htaxR/r2SX42DYsIEhjExgxNqElJoHo9N30hO
0REqwgp7VRhACQ6/M9iAuTwzxOv43k9BXwyHERPkaGaYAVZFSPL5iEU7GvPJfP2EEDTD7TxdXC/L
ClaZUTEoZj7SXwH8A1C2FTYh5S6vTGJJ+8VhDCNnAf2v7Mf9q1+UvmbNH//byTNnAZAad8InbnYg
pApAS17B8zF2tpUtVNRr+70yeR8qUMhU3qParI1pygHavwTqWAm/YK/gpXshDPISvuIcqodX2xys
JLnidlbFk1Mc0bmGi9dtNmHoPGfTVVZUr5zs9Of1ETpmsgDy5FwuxsS/+4Y1oEJe7nf1/tlpcekA
2F28yPcGG0FHLOjOQXH6vYqYcdBzoOFHQ2+Tpnkje8/kvz0mrBDPni5zl6+/1MTUPtzikzu6HtOj
sZuvrsEcvKR8U4P0enospAU/MFBvZ/q0sBB6wMZbka+hrxtuYPf3ZAGueAwQMaV77SV0f/51WWYH
ELYAa4Vp/dLbZJYnGIwC5+IAFLJyK7asi5OTvisqobQa5W6HCHtBUDE5AVPRTO8ZKM7rv3pqXsli
I4Bun/5x4cUr2VMCYbVr314gsAbEXpfnev1DTuHFVrPKDnCz5PHbCDIAR57osERdbi3QETgO3xI+
VXKhYX8/6PfbfNGETciX3FKAfUQV5y7agjOgRo++pFnA0altA72+B51Uphv/hdX4rfI3lEcp7zh1
sQ+/jHkY6u4AFG450Mp+t0IwKqsSa5O5nwhUm68Cw3VyuWoXCQHmG50WwtYa04qE3L5Sm1YjvJxt
O5AtQIPXJ5O3Kbdh1TDqTjRClPW0lJiARi5j8kn9E3zp57wYkfTtv6EETYcLqzGD4zm08ZDq2Eh0
bgM+qXmRlXi8t/RlT4P3aJNhRfFLklMFGuPtuMs4uy6wxMJz5u/G2frKYeQWUtnddeaGIsWJIzTa
8IwGGahA5b+SgpO4WrkkZH3VCzNVe4ZoDNFNeeHgrEpDyfRUY7riXLns93q29YhW4EyiSLXoqwHp
OXFxaO9FtsgOgJ5vKp0fabI9R/cC+Y9NbevCRO+z7pWOtY5DtfEVrKwEXqVvMAYBhRNPHVjizfAl
PLnfwxWCpwgdvZhduBO5l/I33RXpzX45mfPDe0ngaT0lahDeOlWIFB9hrENG9UN+IG6WsHRzbTvx
CZQ7AU1ATT33McxHCeGz5XNkhFZbl5JW6v3YN/Wv7dWbXnCNy32AMR3ZWn2hl6P2Pq74tTNtJJzv
KmaHl+sW6iAa+PB9RU7rO+Lk4AyuWJwM2Knzg5mNSSktfz/qZgvqOwyfsl9on9E3neLiWd81cTb3
vsWydkAuInG3l8kJJateA//UOVZFS+yPEOcewUxXXvoys71CNh0+d+I29TET2ZioUty463t1dwER
4r+bi9ANGgMjpyJQmpXm3cmGFtdKsQPhgxkMh+8ZNkmXB44k6zlLcXqezJvsJKvIBIicZIkGLRz2
JIPNLX0GbOmUr0SxWp0ro7BXKAhGRoHtou52Kv9xDtrJc0uoP2jdlbeQAfIU3rdGJsioWuxrVWO+
oDqokf2ike19+66trGdKEvexX8CLo7Wcg5km8uGZjO5zzGV7Y+vlg23hhx4ZnFtralid52S8Bq3/
Hkb1EcCLvQuafmr0P5jzihKReEjRf7qeLibz7GD/xz6M1iRDGtrt4P4MTcTPfbVswzXjhIlmF8hx
2cD4xem22aRu4rOWxd83RA8TpIbOZjuM1t2gHFuaDcRiGico0zhBZ2W+w4OwIfczpkwvSsqvMQPv
1HKiOHLbQoChPUd3VV5FLYGmUj83Ds1l6mvJl59dHqtuI3O8q2in1Snw70FP1oXQH8YDKaY5HDKz
9eT20dMDMYsoeeTu40tEqx7nD1U2vgX7CFl/vX5Q8kGOx4qCvejhwB/J0ijOp8b0hNtawd5xLDM7
XlHjvO5/DtdfOlb0kwtR9HAdyISkdGVAxLluhGX6V0BTf3O4GtC1F/H7yLyDqEuCnH1nqzyJYhLh
33jbc6YvbhPU7TuD5FyhHJtfYuc3boIJFVNj+fXw51t4FmSWOld+6kkRAE6knwMPLCU0GjgrtK3R
gSJuom7IsJ5Hvizg7QHfdw5HbbMJtyhGrX7l5ppKvCa06VTE67iB3sPrOLiFO+RPAtB9XrXJz4Kg
fQxu17GjRTlyCxWxB7cZpj6DvLFwCrsI6sPrkuUtDfuoSs1LMigaL5p17rJN4r2o6HgxCwy9rtxu
w3szvnD+NSNHnMU1mQ8yFpwsqxCp6bhnB8mFQiSuUiu/KhXRiHRHDTJfwqq1J5Fb2rWGQRhkIJd4
RKD4EdvaHCotHori2zoZ9gsf5Q/muHVA8XEi13244MCMnHl7YAofItOsNQ4TVRg/bZIQMmLcV6y7
rynf6pAvDBZkX7VAgwWrEB7BgV+Qd8oMCwtWFKIvzXlWijrxipPcKZR7UEpBd+Q9S4tVM2FkENAL
MMC6C6akNzdIBwuzEuqVhQdyGrTToshVCWmboN8553isNFC4Vm+362pD3LZWCSYRlcyDb8pr0AKk
wAbGcQn2L8w76KHSca2R1lcQOkun26rzLcKk0ONDfdaLsRlzQWu9ezikJ0+xYY3V8OY5HSXr8JmL
fTd9IHSvdRApKs7MI2pWgGoSDkbjY37RGLvpefMhVQopqyP4Hn237cHL/WtgmYYfqSKoG/FaO3kO
2kfeaMbOl8dYeBrV4uCWaz+4R6FuA7Z3p1MR3L8n4iOq9GhcFHbDGfdRO0A8FNEUZS4EO0eLDlJz
BeACl19/de74ohsOUMMVEulkAi8kDu6w5DembciF65YStm1MYM1M4Z5QXNGBz6WQvCIh0s6K6Qsu
DciZejcKLTr3eqFsXhn6qeke2UeH8b0GR8Z83h7kWiJkTe8rhc/UtkdL/K5s1f5WcLAU5xShGSRv
cobyJsb6EB8coxOiNCrKdBNHyxZP1T5FR1+krbnu8YmAjv5yIJKiYIlPPTps5Vbxx8Yn6P9gUqLe
KEP+HFoVHiJ3JWgWmMhD9nff7aVXhRj2uGfyBqIqWnyYtV/cdfkDXMdbVoT4pu4Orz5tTugqnnUj
lrv4KnPz+zQ85iJAzQ2iGkrJIEYopzELv+D8rprShBP0SEUKhtHJ6CTNCN6/p1xCVXhSzPNgc5oN
ICacfal5zApbSVlY7K7j8Xx1ndcyk0UpYXOShBbWCVjhsbG5BvwwVjavMFS0gAqra+gfm4UH3wCa
0h+K4zpDEPv8bQoJThX4s4vEko+CEJb19SKQ5UoKhSB1Oh9M33kkTwLGEkXLHbpNGdyCJXrY+oIj
R5SCH3ZSMxEEdqWyLQqvo1q2Gziq8lRBNKPGJmlNTm9EtIrsHnn+VPQ4a5Uq7AjyDpvdN48xB6X+
7OlCNkiuLA7OqriHctvO712umh3oMXzk8p2+8Kxy80NyrIx75gCv6JcG/awyPRc32hiYKyprFNcJ
WTWzRAGEKF3LZ/SEZ6OhXFDVecPs3oa9+/MQTE4rxavk0gQZfAMyykhhzz/Pwu+u7AdYRg4v4G+K
hud2K4CRjuKeMy3wqGszH9MuWdrtMN56E5t5VNo5MKdUDh3jRfbSp0449xNkuIAtsbYbLoBRI/1H
WgY9g68Vpzyc7cGHWorwD2CoetSyb+RRkxJ8xS3+yP7V0YhuWtqRzqexeui8RA8hDECTGc3RPW0d
USt4Ar/2NpfEDu/besFAo1q6u5CIBjBxFLLMEiJwzpvlDc3mopdT3cNB7RreilnqXAMcqtGDG2r1
7gSSQB0TLVNjIwecY7ow/BWpyiCKT1n4Pch74sK5q5tsSNMdcMveKLwwDZgJca5alB7hprur/YGS
ijcxN8Ov63kCbOTN4bg4+fD4ceRhVQ+PMzFoEYBNPiouS051URBP+iCWPXkXYNH0te2cJ4Z7BVzO
OEyDDka8C6qBu0gyt8XiDZgugrh31vMWEUJDy4aufzvDKUENmE010CGbtQUFY/J/3xGurm1nSpQt
iD2GSIayoLmX04BuVdQFvn8G8VetYrq5zj0dldvdRqAp5jgPy9npB6SQmZRl7tK13qQ6DpD4B/cy
T1ZbfygB5qIX5G3LePlFaOs0vRdut3kCTy/N9j9bmkVpZP4zFMQgJnT15v4aj+66cdaHkpocsh8t
4oXGveHKFmWV5zsJuiZDvwRhlK5uDKheoJMqBtF2WzaH19UxwK1kpX5TVngUOy8iwcjdgEXBCZIG
b632/ireKLrQasWbC2Z3c7NnfMvI47DYz/fWeUdfnx4O99BjPIrG02eHDIb5xixLNRovGbtKkPmU
0VgXKGzK+VeDZj9VAkG606H9sDucS384+aqt2IOUnmZeYOaFxoU3F5oQ8po0GoZg5a9tAB93EF2O
VvEvuRsNGzJojxkcVseouYdaK074YtkTpEz3myOKRSd/dbNXaNqFvEEioOUBELeNjGAaN3ZOjn+U
1VXAl5uTadDRfBVmyn4vWaj7cLVI7QPbuLrA3dzZ5EUdY5MwH/Q4k1YFCxysgrs7zpEAfrK1lyd4
AYgroLCBqb2Q+ccIl05hQDmA7oK7Kvd+45SLZ68r1tGzNxTq453Yv6McKHcePXNa5CNQn6JkSAlH
OlzIQr/VCQGo0p6R/llTfRq+o/LeILxLJGoFKAiAaQOC/ouuVS4KgBKu6G7uhKKhzglTLxD/zi6q
/x+VDmu3BkzP+LLZJlYYVnLRBc8wHYoLc0k+3BZm9mUjB3phznZIr4qJQ19p4ngYlAO4KnicSwUc
VNABX8XySVUNeBUeQiH6d4Kzo59ka2dTi/O/lv9mbzNQvJW8f/NliYr+GGxcqeUXcTyL17CGpTVx
01LOCGPQ9T52G8D3HssNjzBUHa++nJ1nekkM/hF7JgTTZf1FmHzQtf6ytKRY49vezY7lP18NlyiU
Xzjo6shDl+BR3x3XhsQtQoQ0ubg9Av//ikkj0Umwd1RhC0HVsTGjkbMR8hW57DLOnX7NDRCAGngh
J0Vp0XXQA8mtxy52H8MWuoqAtXCDdTrCdnXwvzdUjHzZyOdxcO+G1ssZc+rMoX+KGr4N0r9bgdzS
CpDzZQPRT8qkW5FIkpMpTh4sjdtWXsQmkw28GHdGBsQuFCNm/B990jzQG36SezCPz2plxedncSbM
3P1i+zxFomhlbHoRdk9qopEKlZ/ZXX5pVdBB1ZXtT0ef4sdR8vVqxcEuRcMMmaa0vNDvK/sAsAq1
BjbVsFpXnsOdDZQI31HF0bTdzsl2R37BbJc6VqwVAkLE1MAkD2gdomxrZfh/4B7CaXtj6x+mQnkE
tBpzyUTiLgcwZUA8dp8E7rarEkZEzFMSkUcYE+7HWHv8lciB3dT4qlSQHFVo/0r7MNPmPVXwh0WP
mzADyShkTafgypsQw6XKwHk0P0ffKLh6fxbXzXBM7plSRBTWnEqMbU8cS/dq8n0g8uG10iWlqXDu
IWXfhi3oPwRDyxRnEY+Gq8MarkiKuA09KJPlxzUiFFMrc8AzmtLrlHU9c8TONodghMg+bBPeIu44
/Gkb+9F8Vt5JIeFHZXD6kdmvibr0jyCdYR1fVyPbr0yCQBclHj2VNx2KphWytUSutM5uLSOPSO3I
Xl/TJQg+/IZUhsPI1i+Ot55jyiD09EWU7yfzUfFI+ZLxZF7AWydEED4MfCz8+CghAdyqs4jHTvoE
ePhxljVsYj66vUVxlerrJ+vhq4Z19nEnFZh8oWICoocjppeElvB+0lJhUnQqyrGMJySlJnGK4gn6
OuyYfBSVUo+CBnC53919LZn2y8dAlqiLYEKzSEyzaEDG152qzZNcFZFj8zByRQe2PrZworONKMoo
UqYq83T17f+3UjLgXI99bdcypIXhosvgGgnPWcLtaO7xFHJelIE2hqGEKdX1lrFKEH/TYKod1I8N
44hIjDQOcmBVrSsOvBVai76Ds5IkpdUkPbyZoE1dKivCeHfHxV+50g2BruP3m+SwapRm8xFES3u3
Sw4BxxMXp1z7oaO6iaUW6SgP3//Qtz7IcOixhfJiQQkHeZYcmLYFXnSiasyJrVa0FJDaLMIL+/X+
E9VkUzm4P3vIJgqhyVEHhb2qCcCYrRPNhw/5oD5s2KYVuiJ7I6BA4p3XEw9ktotIcrBkwyxVYnXF
G2Jeel5hJaMFDEXcZs0u1F4c/MkZ6H/QQykMaKGYXcBMYMbmcFkVRJMper8uPzP7Lcjae9kkgbjp
yi+pVM8ZeIwkMPAhfyeeIR+CQxdyrpD30kTSehiMF9Smt4lpdmd3fgAQ2rkqR+BUTJeH320pxDTk
zrlgZ52VqgjHcNyngw16SJxHNdz+kMgYu/rDsABqCUVd94PVF1mZmbRM6ym2HAfOCCxYPD8Ms6Q4
MMbU7AQHCwwm1UyrvDbAa05O/n09dV+7NND1RVTDvziDH1JrXX3nskY9rrE8Rd8q/kGRAYqKoxJ8
Y/JmS6ZkyrrT7a7i+XAN0nN4o2G1pYB638+SujbTT8KaJZ44CsSMQBP12H+Fa6lhHBJWKPUPNqo4
Rde0fCzxM1nrG4syCShamG7uq+SOpj/hpDMRAKRv331T4RVruHE+m5Qq5pwnLoGy9pTn5p0VeMCf
wBFsvNXfUr0/lvLcEPM1NDtzv1k6sz5/djulDaWv0IUoCZC4PPt7/wXJi93tEQteWyqWLeVlkgnd
XlFzH68dFJGBYJJfOK3Lix5x2M5eMgF/n7M1qCCmSi3iXR8EBZlvVBqQT23tsHc301o+57BJYq7q
+pb86VuHqHQHVrZmEgBFx7BswHVAgpBeoYGJgoT0Q+ddGnqi25ptbRYu6LrV4tdsKr9Fw+UbyKdB
TiurVg7BFDzeIqTLQv32lNfj8KXJRtK5Hpektv+cYSme+Hfk8bW+P+gl0s2XIXX/kKQfz3NuE8uA
LXAx7s8fPy+V/uGGFBgebhVH3R4NUC/IDJsmJIzAvIioKuOQTpm/GOjWGmPb0Lil8Bab4kGCQN5N
lnFUf0MzUn0F/N8Rf8b+mBkivbrEo8RflBB4fzu7p6htJ47JqzP06t6csJ+KsW9vY8yjMy3essA6
OPVlGFGhSJuhr4zJHQ6mmKYXlDLBwEY6yh8RzNyyWd4i6OOWWqh1oPKEGtbXhPcGduksZtXKVnPe
arLYAqaKL//FtN04q0b5f/P9PQuGzgnL+rgorOIFNclIDvElK1wg+xIeFVVU17Z1gCu2nmG9SH3g
LaaYSbRikf6YDs0O1f9MHFgs3ovtwh2Wikrpx7se01QJIw6Ebe1Jt5uCI2uUE+08pghrikPHxnMv
/y6/K+2w1z+nYcBJbUpWkOOfVA9QoG9LVQwoQYjABmUuzFjPWQV9WXlqtanqQeiPzlIAGyDjl8/2
Ghar/GwxW61F0qZV3mTjPj5uN1pVDnd5a5iAZSGJQ52asB/LKsOY+2anGBqErqLojrXLtR3+RR2Y
kCBwn6w4V94lf9CB4kN9PTirLsvBtTKXq9mrGr1wYBLwk+drbYkrNcmDOZ9HAQ/x3RvlcNLGZUHZ
KOSrhYaxsfG9t/CNHBI+zwJHHk6WjbZVOfVAgD685566dL9ByeXA3gT3DZZqoAksLCyWIQe88qvX
+KHNmKPH7MiTLU5IAFWZbaDlERkUVTif/nIQR59FmVLmnQSzvWvQPPpiXZbHMqMs5ZuscHJCH4wS
thhdOQ+ZJNWNG74ZFoM5EG3l9YN+OaBjY2OcKCuEehCSnHQYprOwa3On5/5h56krCtfh+Riqpy0p
KszGrRr/HXIjWyW/umfEYDATAqqnAKDP6iBfBR1x1Qf5txZU7yIGITz7XpG6p0BYhZdWFjKOdi+K
DuiEWLMhdJhiAND2nt+KumLe3xEVpsd7w/en7fzahILFFizB2sc86SOWf67LlivjGSVDjcOwpl5z
dNhGw3W/jp6sFdonTclPu5yEqIewDHnxbBrLHChAckQ9l7oMj2JUqW7+73mo/6wEK0uh4EbVMLOC
BCCAK1jpVcTSo06yj//VphH14p7zlvcoOabyaskyYAu9qz2ASUfXHw+uj7r0HQwaObnjzI96Gdvz
ueotRszuSim8iJ2Ced9BDaJJHEyEDIqF+iweyhhwSZH2bQLHsgAYLVtFnCF1obHueZulHbjPvuRz
bCDVwEcHTGoG+Gt6PX91gp1P43Jw9GyDt+tKVtxNDsiT696Y3HVSC5LDym+p4cSRoF7UFhRK6wvV
totaYl4nLaDcyNtKLkYQTQ6UoAWQAOYyqmIeFm6GS0eRInO0EOp7Ley2k+t4HlRP/2cGMpjT3t+b
8gjzXFwIHcvfNwGalSz7RP9oQzmxgr9k1xkmpRha7Y1H3mh1gpF55gMfRgbPB6R8sJIfarCUz2py
1PiWP4mDuFl31XMDcz2NhEs4PllE0t97ShN0B9yHzj8WUuMZkXj5kIYM8kWhkv+wSNdPFffrSiZY
SL44/a7HzD78lFjtwM8nWi9o8plrJeN1S0r9vOt2XHpg+dbLoB/DEug/hwgAzZbcPfzQz1UvWhKv
4x8MNBb2k85zMuGXkMAURP0QCUUQNigh/Xx9dD+xqbH7WfbO1tjgSQkr30LAI8Vln+8UX3eDLTOX
OU2n604qCH1xrQ0c9V7yiIRnMb0VdvvFuppWa/R+FamEaqD1jIXgLcw6YF2F99xQK8tl7DpBHyS1
0OJZfI0vgAPwVHL1X4GLctv9Kz0FPvqtLL37xVVCcr7w4uXdHekrrVtWXVixNael7/Tt5H4ZAdou
ohIqc1cEyMe/orH1ddd0CEPF3v/4IJmP5DSDIaWETgoX3tzWQMPhVmYvdB7BR8gjhAdE+WCQdQpq
qrefE9jDdrmHBbVUSe8VtLrsSyzmaDDMdm2v7Zlvxd5L65qH6B+8dx0DQlhinwakJIIk2o+6KYuL
E4M7/SpaKxIxfDBSgON2XUZy1Rh7J2Q9LXUQefsmueTb9UW36snwQE3PKO8loIUL/dunCuvlz6uS
Mzm5RKMXbEMr9xSTbK7rAxtUCpbOrLHflL0+zUvX6J/RgDJOLqlkO/QyfQPLFcevBl4JKBd1pMTt
9nui4oRG6J1gUg1gnetd76MBH3tlLyBdeuD8YwQY7tiPj5wxGFf3mJzXtgDzTEZh7HqxTjta46q5
grzuqSt/Q139tVLyFLYZxFhDwdGhVGMu3Gx3luxsO0zpEmJCEWy91ijetFjMFmQwr8TsMCytGcWK
zaIpF6TlfLfBAXAaL74oAacf/I4uHNycBQNtTe8rvxvY2PJKhAzyfBKNJuVUsC+V4b/PDQmmG1Nd
3biqNhq8ovb4XsVs9z2GI16HPKek5CerIz9RAyj37DkBXWAx740UYPrghqbteKH4Ip7wMr1+pxp0
HLvRMisMKav/XuT+v7wuTkza6Sk1QHzWNZG0EvfnTQW+U+AfP/2Z8J9GXdjBLncS4XNw3nHqgYQY
KfsCMnnJ6FMxsn6gVvdJjMBYtbOIKsm9h47FGpsYkEGX62TqJNELi+niYwHYLfjuLqDvHZIc8qgg
HVQ4mWT5gSna5e3Ey9s2u9+UfTA+ffEKMmPO8Fvn1myCOiQxqNQQ8x3MAZ/X2P8kVCkextX9+qOZ
0QxI6V9dq0ti+JaSq6Yh+103ZyXIaP3v0mfKGoJJO+vn+sb1hpuoByvnVQnvM/FbSwG4Mud0iT/O
n3f7eW8LVJxRgUlwTxBnk1Yxpu60hKnLcSor29A0LaLxjKfl+KB8bSI49dw0LD8a4lIRtsYP7SVs
JGoumYD7FkLaJT7Q/ZgL8m48z8qMqb3hM0UEvfwdeFQkXSsemnxEtS+q1Cci65Zg5NoAUlMYvXNA
EZKSLyJbW8hQfuKRKoNjxFiymA/TmszZAxeXM8GNRiAWB0KGp45YjFbQlc3vRUH67hTrf2X8KSlu
cENe3ygD6XAzvPI09uvQ6JbUI1lQqNKd1EtRkM6Inm888CVCHIMad2EHeVEzD2p1ZnIM/dPVzApV
PwAU0YN6bdNIZKuGMG8KrA7rmC0+Zib9p2T34xxnJNmis31DULrIlfdmb8m0k4PQIBd4gFjoYrtt
jrz52QFHY4FrJwAHk+i330wogDbceYRr3HozxV7VfAiWtSCYqOHncXTWr4mmAqVsOPxIltsW6RdN
a6yBQ0ZzWpeJksu2hASVKK2ac26/Gbf8k5c1i/RPMwzudaJTzvhB/wzNs+UnjBW6frm7EO6IiQgU
ivpTJf2AdmtQSoTmR4YSFN4HqfK80VRQ8oVmvRKZ3+V/o9Dd/S/1Pv+yFEQBxe1Ez/ODhnC2WnxN
UAFDjLQZOX29fSCWUg0uLH6cum1xI6W5N+x00kKGvBtfCl8XkSoJrykJOIlDnQlc8diJ9VjNhgVE
vc89oYq1/ZRp7aKHGrvIt+VURnEBbHhU+2EvT3/dfmFsKdhhy6A/7eGL/ETEB3jTvnX3yUQijP3p
oGVuyimaw92XR7k7qu/FeIvbaLUjHBnmFqkLw/OszySgCdIXrAyOLUpF9y7UeMFQk0+/RdWdQHhW
Te8wHuPc7WIq/pEAOgkJPs2G/XJlUGPwoexStUSNi6U81896+cRwVAmg/ed95HWMCniMSt53ptPk
10zRt9ZVy2nsBtVYvPyi05pC8qQGOZFqVWY9Q5eLmDub3XSD6Z3QWNeLm5JMoTsvllCxPKcU4jp+
N64PU0/zSd4pJQU6MZKC9y+/yG/2JYHSBnfi7LdyW8w3hnj2L/TljNSmkXglkkjgNF5djWCaRPGe
+n4OhCUwZ1fTn/JIVYmKTmfosTyXd7yTM2VG/Dgiwgo1umAH8qocZvMZBu7d9HLFpB5a2BlYDgD3
HQg/yierfI3msN7N0QSrs6D35/FDZQcNC/oLp/cHAaG48hiB4mgk6NsL0oidfn9bKCfaAtsH5Zif
LaAVt7XOxY38QIbkUKUGoVfXK152pUlyCaoC5XKLtS2Wb9yPaG4mfDykgsTLYoufqTll6rtUGo5/
z0AhLNdD8EDgFnzGXGm1zaUI8fij3UOaY2aLk1mAbjKVujahjrdx4tgmk1J7NhNnIvKc7sDDJPUf
lWHiH3aNzzarzkhVMp0LidV77WmFB3t7e9QGDjEQJt29KWKTueq5Qp2XRM4ECcSK2iC6on8iN3Xi
u1SQBn+cXJeAnfKZT8XaFczEQHgUT1zkwvYPjF3znQpRWWBvdEqA+exAYsSiiU/5+hyyzOI0tnvz
2QC/GepHSGUbaKNubQjcVk4Ud+QS304F2Wil7KONcx2DtPqnLJpQGpR6kQ1A/nOugpC5VZ6bwO6m
UTbKgC2rrnX5Vu7NECxpSJywB7ppkXh9dPDt4eBNWiS1LguFFdMC8DDCpF/PGpOiM8/IzNX8G/ML
6ih8xa9fPPVE+5dMWGaSlfUNb4fBJ026HXLuxWBgaPDgrXjH3vMwcBKg+IO3bYnWwXQqK+89mFtU
NTJypqVXJIQnJYXWbN3JQkeSMfFi2EMJYSRmDEDN8OQr7tiOzbroKhHV4lg5rkwWdMp7TEaMWodm
GLmYbneEbnhPDuUb+xAsQsD7EuICQdrOoJaNbwZasGMFz9oFTPEWqLPKtNzLYMTIXfonuMJuiwnk
GzrX8hWAkLxLHkD0caJrmvx46QzxvbIhIy0gYllACVlaFo2Myh/uMGO2MlmSPIbsFbzlrCsg+oOG
mXOlxFkO6mSlm2S2TYEYK2KwvnzniYAc5T+Gm2O3KP/f9vKbN7omcHSRCd+4li4bcQBEFBL7NS/8
Gu9LsnY1DeEOL36Kc3DenPNKO4PdQESzwQWpT8xRmJOTn34Yd4WTua7465Iiwee45DuVSgtLc2Pf
RsbKr36pikObnJsCxnjS6co3cQFabr7dJ2TFLXaleHZUrfUJ8rz5KKW2eHkKlLHnOJHcxgOlHESe
fjHZyzuCBKbZ1Ww+BhHNck7Cu9yifTAHkdLXt51rLY/6rPJD5Lu9KQp34HbozeZ8wEz1mgRabyqd
wKCAz1Vghl/xohdZYOOlwYiylb9qy2O7SVUu/4G89b3kaVBI9V5EdDYKMcKuJI4NPyODhWobHFkl
LoOSlmSgiVd1J4MBogrLYLNQYqb+Ty/mEVqLfZWE0qsGrNMC6rbbLLKeV5ZU7ag+QBsOIyaH3uXg
XGSU+iUltivyhjA3ADFq+WcaRw9cw/g/5RxuTvHbNad74rMQykgpWjIGHRS3dO2ubmNpAw/4neDK
WthbzsXpEdfxtBvXvEetxZ7i5epGXSiWOPfIg+H9Oqqnt1RVzfBUC7BMyz/yf6+2vAL8Uh5R2p3M
08IdlYRxXaCf5FUrgp5wdHoX0ctYWznM8fWy7LvOrNiKOLKbokXdf4CkM106BBLCJ0hK1CrabIjy
y9FOCa5p6oNTKoN9ydqiHTbH9BKqPqRzeuSi7t/m6U053u6O2c64R05TY6ueK9S7Zx0z1A9GZUlu
ir6p0fUI8vPbs5mgYWFYYfUhWd4g6UpvaswF1X13lgpV2yPyTKrsrYR9o37h58wSq3TvTHQwLCSc
7RCZ3NEQpO0GuUXwkwZvWl52Krbt30S2yvfSB+oabeQduPpMKMR2iRNCTZKH2twlAlgqSP8XeKR7
8idqVMk/tbNh7EnxiZfdeDyGhbp/G7BN6jxqfEMXbyd4RAhV2Rry9c/Q091f/BUgpK+gNBJ5J/SV
0O1EVtzsH+fnHW7zB9GFZJunYCWOi+m1JSvtc/JoHOkCSDeggnqAf1Dg0L0CDw4ISrcR3XWsZZvg
LIq3ewuSilUKkxMazGEu9Z+MoCBvQDqfkc8AG51O9n5buA641zFYpIJJFnYv+CR6ecZcKxBUmp+/
0aO8gWHKrGFIZa3YyHGVXcAyjyBJ9Ri9G1Mgvobc5EWHz/e00SrHGeD9fD3H9rwrV7pdBwIxziY7
Px3Pdh0QRuYNUSbFVXOJDMqNeQ46bE20oFPju1a2KfYhtzaxd9UsnafdCDEOjVhb6vsP8qqNprLB
NHSK50qCEt/vTazUxChxSHq3gejPq0V+rnFpr4FnuxmXGC9fZH6k24AzrlXFq5hrTF8NLtK9bLMR
a8cqiJMNQplewNv0dC5PfEATk8aYLKOPFl7JpAtgJ/V496vOLpcKru5u47z2xiCnHJIT/7nrTLVx
QvmNhNKjbuU02MGEj2W1ly/r55MKeHYK4Ekd8CjJnjnaHgPNLsvJ/uDrcW/wtebZFVfGcEsGmiLB
z6kvIMGJaTvsJm6q8zqab40Wzxn319XdyHVcTvFaOYs0Uq6HK2pvbuWWS1kYNt0cg0Pvx/etrTBn
ImcjN+hm3F3yTrlNPy5TDXk++jrbmJkZAlWNHPAPqr/FCZnqrmjWEL3Q6jS7dUsEUWvAb8RGTMK2
4R6WQBbrn6hIQGeIWU2qSudausB37rBDAPKHSr2O3Edx4If7l7bCceXsxXxdgmj56h+2iX7kGmHs
zQUz+DBIQrnf3giaigLhPduOPk+UOisGYF521cPz7PILxG/rKTKQgQALqjm4lU9u2KrKX3rPqLax
hekPjL2nQunlD1dZNp2bRiROQ39cpe621fjz/HebTDdoO1RGdjP1/uZnFUW+U+QkGGxwSjeWB/+I
rcd6oKMJ4bKx+PEORaDi63SkkP5/k3tEHTD57j3KxybLKXoQyiZ6FyI4d76xQYK12yMIWfoVY79/
yCPkk2ghResF3J+n2BGAyfr9AnlnqINdLkboPAy8gPLsMp3WDAOskDk8x34Fv7xMc+FOcWZziiy3
Z/k4SsBYVD0iJK3qOzWTogessslescFMNwKZadFzmFI3eygY2GDqohkvEEon9mz53KjSbXsA1hBw
FN5eQKHrsXokYvmV84JEPNUfDHJKfiy7/7BOy7LgDrodDzGFHzjvN3SZPW7vDxb1uxA7C6xTfpmA
J/pqNVPbhEh3rp//xyN5al66RRmrdWRVndUNP1Cp1Uo0nRDLqC96bdvBrMTa4SAdmbcHa82yexap
ukXtrX1feYI8g4zzKOxFADYuQSBzsqXI7r6OYg2vNhyOBUShKufvXtTRMhtxfDUoEDZzP1zRfiR3
0qFDwhactyKSsXRVv1jf1lXpwMu5iHlDx/yPLPz/g4JFg0ZnEvZnoRGBBEFavlysGQYpwtkqJXE7
eGsc2MsZaeRp+ennzX2BfiE1T6sS6rTuUxcZ/m/TGVaftTb5XBzuuzKc1R3ddYL23bAZm+rup6LQ
beDWbSTAF/ii0Bo4b+GpeGVcvcGfFNvOjuwdTsVmkRYYUgZG+PDx7fUGPCeYTKuReVjwspvtc+3t
YnF0qoUS9QWE+FkhH4gM4UD7hVdrc+ToZGeghSB04ECN83gRB+bb9dHzTlCrUW+5PWC36eNevJXN
A3VbJd+9EHivt2Gaoh3s/wct1YYdo9Vf2YZMRkNRZmg9J+6LpP8p0zn0D0C2G73ZIFwMJyrQgSsK
/5BRUIOxpcU+6D1IJKsnjNiief8nQAOrZCJ1kIv1Y5CXStwiY/JLpEjC1vKwrl1x179i8Q8BFKac
1c+AkCdpBEHoAua5+WyIkOovlHTWjds8HwokQNVCXZVqRcrifV7tcSSrQNTOcPHblK2kNGcQpW4t
adAdlq9mFsA//4RvK14ly2GZpgPwlwk8GJLs3+hqqs7ebprmrUIk7bVIM1964NXs3Em8DDUM3ubv
/NJP6dvUXKkjT6otfUfnIYwIV1qlKpWhxTNSPnBTJS6p/YJFBFtnui7Abl8uNdngfxlcZuLyVZve
2vAwSGCvPxi9xAt7/ssO/d3cCmOp7CFmzOat7idIH6WrJSPCQowXwKg4B60BLw6otYCEHjqaOiL+
b/c2/JbT8+WZMCuxrlM0tQJqIJnZjQKjWcH5dtdodxr0lXqle//AHyzbdKdXuZHNJiBMaGP1v+jb
Mw5jsjurWR1mCxv0zyQzcw7ZI5zOlo6LIgYx/0dRug8kbfUFSjJ7p51SJopn/kdEgTXWOz+L0kxz
zUMA50EBdms7N5sJd6jtKd14++cx2voJe/fii+hdMXaojar8kmjFWBpXYm8OcVfyw0Mp4UFt67JG
8uYQcriqZk7Afxr34EJE+jA9M+6XGHTxWIumollIzn0y7PnLy/Z8rTXJMT6Mb6XCPISOz1rm7Qbb
Sz546eIudEim9/vjEEqbOG9gp1yteB7sshL1tnC5tDVNhKvYqljS30GvppeiGit7neYb7CD5yZ9D
99LeJMh7BXVRlLHIJJND91gHwbDe7cYz6XUyN2bjF8GnHiG5YSSwusKt7Qsgi+omWl8FEhHfT+Y7
ybigV/x4lfgJmgn3dei5z8TzdlLH+MqRHyuVrk+AX3nmfsEYRvWZI0kWp5jvgCpk+lYa90tpHgTX
Eki+Oj0+TH4cNMCMaw2qRVwLVljmeKJQ23ngK8y9nMCL9u8xDLITR3VFHr4jCXpUbmFvGRnS9KHn
oJWSTkKCVMkAkNCLu34vv8Ra0EDgo7xmI5IKv0LaBjsjJD4zcZj3OhOztdIq8vrnw5icEz4Q+ugB
ZXJZyzcRYuKcgFrVpaXSRL2xOcq31Jr4XR+earQltDRaox0Wejh3TWegDU6v7oAORc+oev7Kv2w1
GeDTLCM/ruUZWCh5JBfNwDar+ZCx6y3kuwaBa+UUPOuOXfGX8kytRbxg41oKWN91oT58OR95nQzq
JMmYdwCyEfOPv1TFrtnBZURzdeky+I3L9+eoBWWSmOnPpvg/t3Y5N5SEIcwfobw2y3NSJGr8RODl
+VBhikDAEjHjMMEmVHll67ulwnt5NC6PEWflePoHodV+7wp/+NJakKsiqK0xWoiqvbPRFDHMBsbN
aQ0gAnZaz+EjG/Y6KfQ2bJYj7425AJ9CsdCmNHafBoXdE2u/gFpPbVDVj3O4kHjLk/kt1yJ2Ka2U
ECJXmT1mKIPGucYDxbhtGDqzmHak9t4c4+I9iuxPX8iLNeF3bJXRxE7ES0X8dA1+xpEJCuYWkniD
6H/zCr1pI+jtskpUam+mWZj0Ei0530cq1nP9ITEpVlPeLDlA67z5arqmYBDo0Ohmar6oyWGm0yhy
VRdojOdFBXFqxA3SaRuBUyqdkJjviBO+6j2ptV12maqozdaeT+snOP+sXIDUYuRM+P4ibcwUqrx2
3Uc75oulSPH6ZV6mUyhjVDT+r3It5mPaMKTNlkCVrsLECoJ73ZE+J8/bO55PQKrMNkz1zdT0PQwM
F/rVvtvN5Pl8UeKoEOoghF91Bq+hx/yWgiwlFhLbx1Yp1cJS3kYJZ+qj0EK34o2gUd7bh3LNP1WH
KycHhvXGBwr0XYgxEfri9AK+HxkXkdRiIwv3o/GLSV4nOyj5u7bo8mv6H+rooNFqlbUf/TANL5dG
IMEDh1iuFX8zAE6Ld6tu0KiRihZiRbjCIKyCx0lfKoYRA7QBa1KLAtIcWFYZ6CwMld9fS83vn9BO
G3GJR6gz3+BTA8hJSS21npfKYMO+s5rkYFd9/YwTqo1O0kK0sgPVw1YL+yq4djz+SumINpNI5c/W
Ww7Em63+Jg15scJX6aqAcXMkHePcL3vqPxWakTSgcw2ErxOivNvkvs2AdAJLvmTS0AHNTRFYy+1f
lSwio9ThyFfOYkCJ6R3eop3tRSWUa2H5Wg6uCETKFq6vPxTxAYhk/0EE17hMlKrHG6wSeruCfn4D
dVDQ2rc7TeOB3T9jUOcasfM9NTUHJ84Wsz0jQZLgKfRY9tq/uoWiscS60t7JgWThfyNlonvUZdHt
7ZM6iV1Kag83zYf4+NFvDsy4m3OOPGIC9fwYjjlM3MtYToLuf23ePyvmUThbCMHpLEPI89f57p1i
K9EBGAlkFPSnX+hYwRBBh7lZZaYJ+t0G2cVWXkBhT+h9hDrLOFDoixk+5raEoS1AJiAm1TzmeGqF
2gwoO/mksm6Awe9jb9eItyePlnwdxZud+Br4Z/UnBWpwM8Wss7aYNDx5ewbpBYLIZ97Tm8RTTx49
NyvekZngxVSguVvPy+ecJNfn5jCGXHjOyesHaO5Szw0EoB4DvNuCnH6w3pPKIriUL3hCknAEb5H2
765/JdA3id42ViCPGWgDQVty9JQgYpOLYAhlc4bR8aC2XCGgzYJEqCtb+tuMM0qMAMRQExu5Vl8W
wWhlowh66J9hwM83c1+o7yog8R+NXi/6WJWxe8dJufxAnrUBipoM6YPSrTHiPQ4z0A8hfmNp7GH2
tzpEDDnXdXacsUSv9ZImVmrjoxDqScbfGeRYIGAGqLlXUnmg7F4DWT0QEoeaa2FxjogIs7FBvft8
NrrfwAMKcnbnv9ZWYDHOJACflLs22AIcjO+KaY/d3DW8P0L1p8N6wgGPrxOT6Hfyvr+Tel+0iU3R
yT3HgfhC6uRG1qDcs3eKGSUtfuRdPxrtHf3k3cqvQ2dzSMe+EV4gXDddvXmQZ6FQeJ8Sr/KzzwWP
XLugbKdruifNi5eszDQbAHOjR13qnlGsyz0YmG3fM+Yj2d1ab0rtO9/t7Av1cwHCR/RMAwOxH4q5
6AVFX5Mus78qBD21S6ePSskOu3PSJ4wU4ObxN7H8R4wK9idMt+HqlcthTY171ebpycRcGY+gBU6f
lIpcazZJYQ9MYH5o/47VpJMZ2zQqahCR1gP4Dbh1RVOl+zeYZZFzi//SySypp8fKNfDCack7FIsS
RJLmvX5oNhUdmGUhxONYP3Ue3nmsX8UdCgCV1o3rWgT36+iHjvPAZPPDam2MF4V+YREr4TxVjObZ
5WBMRUvXEHzl4uMIwnuePNkQl98sqYOVQOh4akiV7f402wW8fxMuAuoF93QEzWPTeUb/zma5ABpv
env14n0dlUf0dcCHPZhIUeDD1yM4Gyk8JN67cVzs0yJoOYRqZTpgb2aAjfOChQvsV+opevbfoKpR
WOg4IOxPFsxzoR5zPPUYrqD2ierIJ0RQt1ddVV2+/HtM6DtciHK8I+Y2NJWYFhf4+bviT6YiizUU
Uh5VJxd1KPszM3W8xFLgxjIIPgqC/UMWzL6OXR3ogdSFGbJS98AcaPlz8Vr1IWSpzWSPc42NdnHn
go8MHEQXw9LrCVVH+FVwhONhTB7kXFSWqV8mh6A9Be3Hk8+NH5PUiuPEhFJD5GrOefMXIPCL8Zm/
7w8HP3n2DT0uL51vxkIoW8jajf7yk5S8fOmPb7+6ldgOIJ/kyqI17QFUA7Gr7AMxukDEylvD59L6
GbCDpc90RBEFz4tb6Odq7GMTe7DTHaUbumRmqyD2XaPwqyD+2BtP3vmJoJKM09gaBa2/Usn/yonO
2rGnQ8CPUnX3hshJa6GO20sBZOVhWEqh8TS3wV87cY2kjBl5fSihJ2vS3DsvdjAJEs0iYf1KGC7/
qjryB/BQxsU7pEhMSDL5eBz6nkFO+6DvxM9nmMB+YuGmK7wc8BWrTb6+M1ODDPEVi+vUe+V7kty1
wjKqTepcEqX9dMhKxgKElhmsxwiwkztfIU1mNOaSj+/w9PLGg1seQxzqWYhABHVVaUhZj7kFv9k5
huhbpX9IYah1opIfe9wFJjSAG7dHCSyrbFLnIdE6jxhfbsA3AEQMkn2UV8jCu4VbPfFY/JxaaVLC
MvqzKQDbtvy5Q5Z6jE4iyI/HnILsdN5Dx95zePOsAD2CHV3nTNd54L5tOpWR5ZcAHCYDpTpS8gra
QSRF/w8O1cnGG02ur9EQ/eIUPL43fFmQvnURKSOF4jWxVO7xDPHvgBQUi8lFxDo+wPV79sjARyK7
GigIi6zI3P1h6W0J7+MiT/w92uVCV9EjzP4hxFaxfOl/+f3KRuRaRxA+FH41d5/c7Vz6R5jraNEk
Wieoj2FJ9SJ/DdIFlNdYdaWMy7w1imhJrzyyBtXQXoFru9mLTnNrC0t02J5LNa+El5wJ6ee9sJ7s
vLy3Ux7c9G3jpUSX+WcWHeSRZAlVSLmDaPYnFc4z+EwE+BJj4KLujPzgeWfx69sR1puaqA5+ULRn
uQp7XGWuLJbhKlhK3abWOflEURU5kiNYBxhr0Fyu99dMmKqXY5mR0x6fdn/QpAa+c0WW2sQeCWZr
i+KJo5QH39usZegPCf4k3Bzr1VQdiAtfzxRxHlF/qLvHPG8tEQ2A/XllQwp3aRvnn0lDa0kHQGBM
cHxmq8QlvLpO/m/kdmxhEIItA6GGNTorHvZgDeNxmyi8cg79QBaULELO83ya6n3mDlg1F5slIxSU
zI9LiDmTJnsCH0jUQ7m8I9mCxRukXjoGKS+pEkddJfrcXsP7WsUIZ8hNVfMy1Jgd9iPFkDAormlb
7PKfb1GsUitjNx7tQAo+FL6ueveNwwaCyfV58cIEtDDboPqtMiwbxpGPXu7rgZY8KJFUh0t0g2g4
f6NyHe7PsjoMDxoDeFcGm4Io9d4u/lp1/n1QWO9th5XimqcHo/kv/KVQ2KKOr/8KA9xBjpLJYK0m
IgbUfsNlg9HG75gT9iHXbeZG1/6cf+6taGWj/tnXpUSaMtUzzDnH9OBWore6WXcO0GcyYIIDkXRN
tx2VHshlHFXdWkKBVTVHZxR7UF8Qxt8LvH9kLUWvoRwWc1/megR6O/gLO6IDfAkeF8rG9BMu+UHK
HT0S7wFCPjsJpGvdHPgYO/3LicVM86mDbhmSCqQKF8bzhFzwQPFLVam7aoAFVm3gVW+Z7VwvCVET
AvxEHJOQbjPEL8TJaxqsAocQJFFmVNlbqibxm8LKeELrv6S4VHFAAFX4ZflAZOQ5zi95TmY7E9BI
8eKJ9dLfKpnEA/HrP+h+oGUJmjobvfuwgTeRNoXxLTzZ5ZMLusz+OItsrCcyU7F8HfbHk5vMs0Hr
ZmJW1vjPENgQWa8nVdm9S7LqNRguNrl6o1xuvqADRvSUIOVphhcrNhBLLQCdaWtsch9/d5QE1jXS
qG6JodTf9v4f5IXqzkf4x7oxk1WzK2SvRhgQEhrWO1GfQCirLrVIJIeX5BB97VPhmTENm4q8ZoXu
8C4DiFaDJ67sci/L0WWZgHeQddCaWDnicJNbnnOJutarGxcBVzAaBBwcOiyS0MTC3NvZB190VryR
9qLE5zFR1pvYXA4Ura1trCZ6GI/VJmpxAiNgvGtwvhkazFzsMW9/aSxVgIyfZMTe31clpJ6I+sGp
/Php1rvlQuHjU0SrfuU48L0XRshq4JiOScEKTSIvyTI/fghncbrtYkS3ZEX7vurk7XAzYPQMou1b
zV2lv0QOB0MPz+VJv6hcRM0cZr1Y6e2DLAEENYeJ0/C269uziZSexs9e1KCDtK2IwMRTmnFcmRib
MDtfDinoSoSoBfl9T3cyYrmfX2msFSLyS+tOFoR2hMZRG/3tFyJwXmopCTrkYaLaKWLlFrRBmFIU
omMEY8ljiNMbm+Y4vtlzWLajlV7ms5FlSTlUy2hPMIGFKojqgcFHp5TG6uxqtanWUwpj4Cjvwaie
sZjTC3043/QyqwYe5xCxluHssuqMkf82y2/48YzfaJELc20u/le6SIqdUIf1hI5EBllzTq6OAZTJ
XLsNE+cm43Y3mVRQRrXiX7vbv3/1g+WKxzYfPeFTAuq1TuGmt8bOB6Ho6p9RrFtfj/vqbkFoj342
E+ioRDr4xc1QdeYSK2oPz3LKMDKXgVgSM5hnQ+X5NGWblkctb/BmyxQIgtOiYOHvSx9yKWRPxaUH
a53hI6C6IM4t3JbIIwQ1yz8YbtS3hEiUlpjNYMZq40o+yhbLTeHdtQp+f+oj4sijgwKCAjQNiqnv
1K8+3d2hAExUBFS6edFHWTLZHCOdNhDT/lVzPFG2hjdk+gqOSs25/FU4gmSZ6LTvg7SMSO8SPn6g
P9X+j5PVQ8hOaul+kyzfiV2VqcEFIw0KrmvqbjytQQ4f3l7yc01+SjvnnkdqqJIJ2Q5REbIXZFV3
Zmam0LrvOqELbaGKxQONexwNyYEp/UmXx4ajEOt7JQpWo4vQa0OA7s8BnT9hA/ysIXQTMjRH8IsE
UmoefHpgrQUIcI/9v0u7svIds+Dq6KPI9/aRRfLtFZfyWsbN1q6bGPNrv768/FIY6R7m5J4jDOQE
2vG7BCp8BtVVzBl3K70LatQelHVVEwndgF1SDGSrK9KQPC0tU+Hp251HTwGNIhk0olIjpmD7Laiq
3JcM3AOnU23Uw1kTnywkkSzyqjel0J4QMeiNSZSdQm/4Y5TSvuJmkeP1CYFurbzfsGzskgN1PWYY
tjRnEKOm4A6Yh+I0zEGGfncXju/LmzGbRjDrf8CpEh8NJpVojZ9ycPaZhl6tycVUqS78Pb9iE6h2
hc4U4eFEm3JRTgjjj5h7RwrgDkGkwGtgoaKeaV7ORiIhZieYFxlfH99E9NLY8ZczrmbMrBMpTHzZ
JQ5R2+cx+gGy0O7k9zTyIkha65CyRVGVn17FiZDhosTFoe/T0B/RIvnqmsSEzrQX6DvE3ITLaAm9
56oAqWAN9qrPFGS548Noapp4VnOvcONgne9UHlmv0geuRN1rB3zb9HtQpbt+pv1EeVHyHkYAiItK
dXFfX9fPkEVCu9x11uYFQp2j9tekssPbHutEqYRzbhp3gAWht0AGMFkkOtLaXtCTQX6to9sb2fM0
p3zC3G19peicUPaUsthQznIiO4YgKgJIV6NXfrsYJj19SXeIUBQcV0AvISV0/SSiUTgXNOecxpUM
U08Xh2yqNyvsk/auxrTyo2GiH3Ty736fRJ2S5agSB9sKG54PNZIlB3Rwn0L/PyPtYSS88GLMtNuR
tvB2SlchxzTBfHdsE78x+uaEpweGnMesWriPkBufkjuOG/ocwZvYf5Upk/o008tnakRlz+elClAn
YapfUdnxFi6lkHgUkMkvTHImUTBzZScE07YhDGeUDU2mGU7CAkpMDFxVwgIPzklFUdU4OBlYL8o8
aEmRymChmSx0GHDS78fXpiP0xa/vKvnLb+swJ5ZhxIRG9JRf3t9K51fev2wevd/ML0dIhutJV48k
zYl94QUISWQGz4PFQdSQa6Oi5MO6rLgv3FcO7QjRzNEvqgO0Gfd47bDqlafVKi8Gaf8fDUYtGcMI
U+8q3t6R36anyg1Mj1RsKOSCsPLR2XzOfRf7TjxXr/95zqPlPhG9B7Gh8z98fkJXx0UQ/VsZGb3U
m2CwNgjylN8AcIptnTRhqDLqh2QIg2owKawfKNMLvmT6HSBj+GMPN/Miuh3JPzCh6KTScUUayqt0
qpLgia+leCAdOARgw/by3yGdgSxldJ5w8i3Z0GfEuCgazxQft7Rq6lLK3X44jcnuUq+CtumHQEv4
oswKk1EOtFT8xM0GCTI9blqP5yuPrhd2HrIHttl4iWYWZpe5G31tIcjg7kC/2V0W1ytZf04/9F1i
4Exmb0Q9MnjSm3cXV2+RoaovkvQSdWNeOjMqTKuHJ7OJn2vgTOgYDuqn4kshLKKiyySWJKU7y/+s
Mp1nPQ2zoFNKyQLuo5VffUpv0iOP11+yB/I7cIXH3yAoWyWhQGCcGanzYteLeFoN3oR5AoxBz4DJ
GY4vyvd+PGcZO9MFPlsAm2O5cYnSJal3pSlBuAcW8RK+eHGURrR3ydkM1OurmVvLLujdriJ26Kvw
4s+u0Nxi3IbyskivVsZ3YPTHph8ce1iUHSd4Gos0yI9Pby+cOI0/3iR/cVKFS4hrNsTsHsErz3Cc
Y8n+6JRtFzTiG5Oe0cBg1dVTgatRqmf1ioKG1A3sfI8crutd3w0uvYgwKXDUsGq0RRUu62Afa9hp
gYM4o5lZh9dZAFVB/UXgzc0s5+ZFgNPPm+ScXCf645LyQot9iFAOoJCdqLK6IEEqFvIV3PEVQCwq
q+APjA7cyHF3bzuxPmnbpuqdJCd2EHhHnLasNfqOt1XJg7cFUXMqkQ3A9zDTEDBNh3t4sCpFFgxu
qNYuPY8lQc8kq/ETuIvhv/fBx5xTus42NdAkp3i2XMK6Hja9rNsM/V4t6V07VXimL+LeN57SGPaS
S4AlTK8Ospr9AwilUzByBbJFFphLtWCsz5d4JueTIu4D03r0kmUxdvYw835lHbJdalfh1ZwZpv9q
axQkbzi0Y3ckL2HuAFskFSp/RiuAYP5HIVLop2nQiNr0UZC7NdK7nixXaEpGSlUVGcw1aoUX2D4a
UPIICQu+SzANgKipGgNBtVZd4P1KgrRObw2dWLU2Q68bFzdDBpDfM8mryKeMsPdFQgreGGAHqcqs
lUpNzL1Tp5cdH8G8cRqfosJDtFd78a45NUvNWcl6jHgh1sBmuFmcKws9aWwl7SnAARgrbCVwdC3L
uXNaqu5elc/gwrODuRDGu9pPZ0juqBa5N/GODJj+AVlIaQ8A0qpSRsQJ98DQLnneS/qFk+kesVvH
18OqUZu6QcnfxiJub6hJMTdwY/5iuXhGLfiAUxx388Th6b870ZqMHoyepQnampYRZtuW/bYGk1hs
td5jh9dBxBzu057W9hkodAbrnkSKytWpmIj9/y/kglQ3DOFUq2NmRL12I8GDEZfFASSwVKZddGQi
fWhLAacKnhBOl8eNhdOF4RFOLB86ysZEE1/V8Uzbq6EDfv3PnT47t3ecLxYGJdiH3Nb9R2bNNwol
GbKpXzLhIOUDSTuZFqiNKhc//b9A0cQwxPMIA1Y10yQ3onsYfU5+L8Jft8Qw4gwT6fp7ojIGEbrm
mpt7aVUD5USJ6D32sC2E1ECUIp8IMQ5bTjkuYbGf9RHAaXCNQquqAdgWOF52uku8LqDlmptSIynl
QTmwcCP0ULB5BMb2YJtqakubf1Gyfewbi1+pPwWrsfszuQ+GN8lflYg2bjNZarHQaNrknAcSUySQ
tNW3DujrVC3o5qBxsWUGqz+6ZkmShxJbGExPQ6Ndpm/6wvgebuIkrYWaZrmqYzQNQk9bR7iHsmPU
c8/9oE8enRvzyp9M8XiMsuGLrZX/oFT1DrPVGbOT9JTIK3FwNqe/Sy3cbaQdEEvpBvZZFUKKcml+
19hLkGZeVKstsFPNfDP+hUzhUjOalhUm3c6R9hea14zuQphcGR1Ig4fKmoLCAucT+5lDwOnwsXJX
+YEiqO1rce9w1YjjDvpR5Q8JWUL8oSmsbI5Oq6WXQaxAtKqVq8glUf8Boo6jd76eNZgrLzEmrR76
4kE8HOY1WfsFwUEMR7juuMz+P2hPTD0/IceaqfB398qHSGqS52+ZnpylFzoO+PjmAMKV6qW7/UFg
4Mzs6SuqkIuDuj1vmBDbreX+eXW0fP2/VPRNEFxmOUtL8G1xSiek5cNejnEJriGkOftHEdCfu4WK
+X1lhlj+W902lR93XGZRJHSdynNEwiIQEsxdS959IqRM9MjNqDzZ9ee1QNrhouDaIr1UA7DHReQX
Nex57FZcriClaK5U4I+Fh3rjqm70tbdTSZivD2BIw9xK/okgq8FxcKOtDPVy0xnGJgDPp6CaRJ45
QjMcB5J4XmfLFpsDGo50RP5rxu4L7u1oYQ+AAYEnj+w9OUv/MwemteHa4YyGtApY7w/hNh6zxOcy
szTRlOBVLHNfIghI8zuxlMUMDA1xwaYJ3zWFt99jXO2iAwmef+V2BqzQk+GqqEHUOoGTBYE3Tycu
ntWhVy4xsuGVHBLAJyi7yapkGXLHY3/pxXFvgVfpDh18lmmWDowdWyWP0LPk8NYK7ZhyvErtJAZr
xetzQIfnHdGm+hR1r/vJzEJg1ag7RYjvqmk8NE1CicaR5ywMgozxnL7uXmX+X+7KAue9eBTqXSrV
vVz0QhCak9yrBQSlNGpkuD7f3AA5G3dnrfqOBR5xkP2Ll+vR+sqhR4eLnGmklpwOvvfK8ZTC40/Y
YaqYe9ML5AXj0vegZNZdEZJlC/sZX+sZNithTXtGQCgoGlQ4EO783om5m2t6DO4HaUPoOaeNTf4J
r9gK5Fv+vBCOX5MYOeexvmIb7HFBhIerXylCG3DxMmIijF8LCnSj3C0wuMF2173Xf1Xhl5X3YY3c
i468AGuuySo+vJM7s/OKGyr3aJq9GdStdrHx11sBfPdVixMhgJry18XJdQj9jCR6dglH1OA6kXcd
3nDfOhMt1+cTuMjVLyRLfWqZsuL5tL2QqqR8HsVS4hYUN0iwtexglDpCR5OHldMlhr3NuFLHBRyG
XNOBnBHwMoPjPxAKNzdEVhR520uovnuqBcE38ZC7ozjWzALZAKlQRVwsoRaWWSEyiqTewCHs+I1l
qtpOeVh9U1G0d0O8JSktV8o06g1T7S/7pPkvPmTleuHfP5lP8+jpNb6AmXTEvbN/8sb8tMYFT0PM
jffpg3UFg6+Wq0QDa4UcPCo3Il3BtVUrNU3M8QfCM/nY2bF6Q5Tn0WIffrmDYSPKlhrjmumLMavw
JnRhP7a5hlyCUsX73E5D6Ggx0YoLOAHdxar9u3x729L9XrfU6OmIL3nmr7xvUUMgZS7B9/bw28dC
xsS8fZ8vkonLN6ATZygHE7YqxyX6fiA8m254BCPoz4Xw6+a/dM+F04pou17EY156Oq6AW3+K+PsI
/C5filDqt0YPmCglmHtuImuLJRlSYz/6CudX4bM1dmDFdP1orRAEAjK9t8eU1x4rCQumG0gOtW9v
aVvMRgNbzbwXoUqnNzP8+1Vb7Ge4F2ImjJ+y5IOlKe1OTiuWxttzzn9yMjmouo5nJxR57Fpsn4DW
d3wpoGXFiNYbuDtMqcDIvrgV5EjF88WtZfYgoP6zv8bAOj03gyMGS+8+LnJdtdJyW9VBAetmBbUd
aP9KLUVgyP2B0nRn9xRowk3+nkgeyeC5BUA66zXM6YPbcKeKfLbcZZ2IHattXLBYUeaM19IPxR5z
QTJt8R/nwTNgoxekRUm190Ag1Mqu+2efszgV0Qa9Vrls4lfUkOurJy0AwRpramXliEC1PS6gOgrb
UyIn1m4xwkq2edvII04fRsQMROpxk97KsUGHmsRN8r+fHhIDsHur0SY1IXXnd1TlWP/CKV5hq+dv
u6vezskxDUXuE50XS75XrbC+osMD9CjxrCqJ8xXcBJdZHLAuJJQCeCYjVCCKIEoEh240jEhLRbTT
aO3AV2RHnznaEWkPhusdj/AcjCRhv+gLGVYPE3GFlfFmbQCmxYMkTLhdtTjT/hM4Y7moU2s8ur8D
Neb2XxOJtfT461PLYQ7wht23MWJXQFkDwOIOuh3ofTx0SaaRY3tOzPtEC7FalyVHPCBQmE8O6LIK
NPpyjUcnOc3YkAIz30cA7Apl1ukWQTwzwi/8i6q2ruomk5AD8Ox2S9g0ddyNMs5wUwcVjRDK1rfT
PgbQMnPU9He66bXk8jqICpCEyqfU6uGQGGXKU3CtdBfeDvqeoRBAhadIwn0mNjfqx6D0Vkfd1iWI
QKj4BunP+FDokRKFOIWR27l0npRiXIUykIZ5JlRxDkpD+our6BJCmCkRCzTWj1udrEIL798mCggQ
soh2iuOFjh9iegLeE2wDAIKFiW4VkTDZXGoqeLgV1VykzurpW9ej81yLquEaKvfsG0LwfzYzYVo9
wYavQMdiuyo3qpXDKuPBf7zrHbMB63+uV24YlN6FJNaOmBf40IckQUX8jLmRadLesCBWVOwkgpKD
CfOfYj7nDW3F3U4GpyiTBIBmoyfb2QzalMvXj6CEFOulttRCqMhOfqxUXlPEp1MC2fSp9EM76JBw
oEoaWMdiU4vhN+ekukIgAgN5LJz09HK9/+bDXM/eH37rZBvhwpfNPEpW1bigSowZCSR52xQf1LD6
XvWq5wszqgKmgtHQ3dzjj7eMOFydSOTpludYOkoiVeDSEr0CeBQiNc69tEFYaUHMFxNhViz2PFRE
FarlutVZ6yYBmD/fpKVb5aYQTnKDst53e+xysXc+CLKBBTj4dhQE+2spy+X3yAdLK4k2PiknhbIK
8wOfSEiR3UM3KAO7e+YlvSstsjX5pYg9ZEJwc5qhGKf4QomQadJ9SOJWiAWpoqpP82Zsijafi4D7
bxFvSVqCDeJLH6w6gh+7+YAUAN5JQz4/uSezOUtPeavPhdwInzXyhcZ8eJDL+sCpW6w62oX5vCZ0
T2UM7ngF2SOVYmG+pq5QRzycObq6dZEpnwdAj4GgWcmKqtlcjjQ0pPmoPnKilxI+EdzSldAnX10U
dV3f9zm1weQRIml7RVlFqfRzmA6gKdwcxatSFDwNXRkhG3UShGRKyOBZH9+xZafAdjmrc/lmbkrX
KBXy8pHLEXkMtgj7AgI5511QZdnc4Gyo4Dj3eI97WsSSu6VZhyDieFXkEFMuMwarPl+pTSAurXhH
0fZnZ6lWokNpG8bQU3IkHvwNDtGVvTaEsyIQnNx12ydRfwIFbNf3e21go1LOaI/S79xEHYmHnTp9
Ewft6DqLs6m5KnmKJYQn4XtWTO+ilkHx1XxSviFrG/fMEcsHt6J3wOqkM7TWQYOEsODd3BHSUYCw
A0iZGezgV/FcKQY333zM6Wb3SUswbaEvsIhc9rxhqZMhZku+Nd4bRuMUpUzLbZmhdms8K4jib2br
hqDFhry5DEuo8DqM25yEN3duttQxy9phYGIUiONaxRCPZQ3UhsDKYlmuTL+GVnDjAtIZQJCpsfVF
LP/P26cB+xNprTo/2hEUnNXC67lHRryYheAcIrGkdBNZ1HuEpZCcWc8GAtPNUyVbjfRPm4F6R46n
XauzhDfkBkdg1lYcOuj/8uO/rN71Ef649dyzQWoWX4F0oIUAjvkI1v7aRUrv3JgyH2glb2uJHE0x
y4JB9wXMl+puy2lJOHfYDcl1FxQOetT+0/FEt3l5BJcCaFq2CYscXvrYJ5pf8HQiB3aKBWzFS7yT
BCiEBBfbeiWXqgjOdC9OUi1kUvsSP7vlPU7o/Z7ilXB+9CKrhk2k+6hn4Hf8bFexqj9EhxPHbr1g
xo0TOzDhwynjjZb8ay86+kgsRJVwUB5Fo/fCTe1pbvxhzwMxnWHDPPWnco5fQj2uC52b33GE47Lw
+ltOoJ8KG94Lkth68UXdhFST4Uk4LKIlC/pSIlHLkad78uPK7axbxx/NUfIf4KsnAzvd+f4Mfn1H
JzN3m6BHUKXCkE5kS7qsLt4riulo4jdQAnD1R6Gx78gx3F/lX1NoU6RXTF9vhnzFjUgfIqd1Uv0W
PDVYzd8UAfferSME6OP/dizBo2sGxiQv2yJK9cbngCe57zVJaYsE+QrcsiHHlbf93WA0spC5/+8t
i2b9bL2DR7H8B1YqPmnA8EeNsxiGNnELmOhokq0d5c/3W084ropx/3oO1MNOlFY/P64xNBIaZ5GQ
gmcPx0euXBJIgZ+Sr3Yzz4UQF71NbHBYYI7kz6az9ntwyzJcE829mY4SfUxrr/D8EyFf6SPW4ctd
X8P1xl/MFkPf2GckJ8YB8r/jpoPqdqfzOTMV/1RPpEfncWu+gCEXjoDYf4rmSZtcRLQRzv7A91re
lgJROyFxZDvUF/VruQYWCZJpTUMLX60N7KAd6OkFpIfoL7qQIhgdq4FnqaPh3CVqwawrITTWy8iy
uY8vapxqLOMmIhVvxZsVc5M58ZlY6RME2okXdtOBpfmV7W5VrS236R7O9F7Vz/WxqTk1KKDJndGf
411c4BpO4U/yZVeWU/xbGql2ySZunC8OZ7XFi+ayLGwhNtdXOdPi8W4R1UDMilFDKt0dI8efxLPY
fddl8cV6lm0v4Y6m5tnKtkvWuuBPq5XxAOHMmkcCpVRucYFccUupmVAclUA6L58cZi/e8URTwxSj
HLAcne/3wzaVcx0ZEvK3QgWsHazrQG4ef/EReXp53pyk2WTyK397QM+cjPxoc6xVC+9D3VQe+7nj
qKwX3NEzjDK7gunWP4CmcJ5aMgNbM4cODu8yQ7KjFgFhI9U/WNi94WKVFzsQZ2vpciWsEYKXAOBS
QMdbfivZzPHsnQGOVqHtNOFKHnjtTkZx3zKSh9DrGX7P3wrKrvLJcEXXt5jyGr9VKqqkrMwVTEO1
RkBELF0rdDv4G0ZqDktSzEq0h/PWhdXkczNAMUgqx8OkbS/kVG1fjU75Iphln9STzAPR8IEhfCyt
a/fnRDDRJd8aVG31x580n39uesnn+n1Gfemp+nAR8wDDx12Wbgk9d7VI9rzGrj6CKvTHRCxBR974
61uvSpv6AnuNM0hCylC1ayKmQv8yIoRnQoWqFPXgh2iJvV8pvR2j6vcsAnyM9Rz4vlCQYMFTRk6P
0kl+0chtTkuI3ucyDs2sNA0aoxFU9oy9CVkEKX160cEp2M/vnZrJgRb6227493mBcnAp5Vw2/p3x
KfZ7f1X8hEGiLSFsmcBmvDKNi+P8yMo6VQtabRXvl8mDBFOl9tzOz3RU+Fu+M+2ac7EmBPn3Vol4
ngW7t/H+hAvjeWVaCvSGZLPZvS1JfN6IVI0h/a/wnOsK3sUXJPLZ/QL2/N9x/p3INq2IvwbRe+pE
DeOkdI8VbqLHI2KkZAXrJ40FnUyUNRhNJ53X3ci6Xr/OOsCUdojg2sBQkTpB0ESve8EMKsMUnDal
7i3HjGhAg+qIZjCxfjncpI/VlMUCogaN98UZUxxs46mb25gBF8VbiPM4VBCxPa624xKVJTTTd91H
/VXx11rFA9XOxlL+U3vr8JUJB5mAnXCES9UYzHzxDjgMR3j4ZBvW+ycPYQ7g+LmpiBuZodSiH/Wd
xpZJS1Vz+ibihJIvujT091jW9VE2VbEn7Dee1O+DR3nIIuC7dMr4op3CTujVuY1Pnx3NRjS0ZY1v
e9sNBOSE7vS3q6BhN3V++7NxswtL1bwc/QACw/jnAakRbt5bGL2j3XfFC6FRYF3gMwdBQI7KuCx8
owllgKCiu0ikQIeP6ParQbcOs+iljNO2dkW9OO/KBDLRALq5JsJur3+ZCc30kuXhPdHwTnFJVKJC
u/H0BURcqQsjICaV/0zfkHM98E2V1kyFWYadh251P8ZlvuWr9VrDjbOoSDKhcvq/YBCo/l1HOR4G
pSTv0o/WYKImJ+0aJqoiRxlOJmyeDnBLKSESVqjaSl9UMCAOQGCJmNlhsWt5oKrBaUCpQZ/owWYe
VupfHAy5UKU4u0QLPgnub3lwCjCFehmOzwW7te9Djo1xGE3QYOR34V3pOORybXuoRtg8Xz/QtTZX
VBPBFMKp8BsHkjnTKRyiV8i4DIpnns4aH2mUWofvTTPZY1Xp6ez9v+zWXTFSa2m5VC6DU1lPyLca
6fx50h2EFMri7vsZ9ES3rFu+JeFC7RQcjWZtwAI/3jiomhDm6X9jGA34lyJuyJGOcaGF3NkexH/a
VRTfmXxqU7SQuhlZnSR7kDiYAeU99fz+eYtdXopLYjsG6J1KOv8os1uoNAg44rOodqy9aLdmUiQC
VCzxi9rfCFoikH2SiX+HQ/hpN75e1TSZaxjrcF7+N6Vq6pwapCNeiBaViUXuwuD7FbtitnXGW2GF
Ous3ZcDpqn1P7OHiHkTcSQkA1hLTIyqHQrJu+RZx93up7jgKId91+F9tt6xsKp/A5EaclP7J+zr4
OSTJVjeqE7AMQd5X0qxJIhCekktOzZzBNnycXsEr0cjrWLSUC+pGXD+Dobdb/r5z2nTZ0F+xMF/0
J3MzSesGTNJstxUJkEgqv60l6AvG03PHL3p8kXHh9P44BylgwA4UaFw07a6GJWG2OqXMteBhlsJv
yfoslAfslal2bz4ojndkCXl21w41fxR/E7z3zNrmtwwkuF30ERsOqPgk98JoW3aGpv4cnlICk3iY
1fkzTTsBSOo4FiQ7lP1Kip57iOKfoPfHr9lf9OBprVjRm8ZcMnwkdFq9Uuk/bCsCmfCqx2NyoJB8
At/c5gSRyCsAxRRriiYeg7K2m92xZOiJuikz+sbyZ6VzqidtIOVPNPQ4MElEAsG/ReD8o0nsS2F7
754govoRf/uu7KkvvfRBJzvf8BbOg8anvYy07diCvuEamaQetjt4rWexJbeEIzGhfjOZRHHfqBKO
UiV/j4BKjsJ3hzbSoW7QzzzrK0U2F/l8d5+thOBIjsnO8p4idE8NhYxkhy1kF0TzlRThvp/ArQ/0
5Z3bJx5+JY9pzZInOQOt0iU/MVuSc9cJsCdq7fBR9vKkn3KDQbQSefXd952TFyF9ovt/wns6HAlB
28HW5oCmBnWjBw5ts/R8iWpXOpa1V1GBD1rS7EURKiDoXlOGq/vURqhga1DJFTdcyCe5tXmUEbuz
3H7sx3eJzRQX4DznoR6SGruXg0fvusNw55sLyl+IMLas23pSslxYjAn0u7ZbdCS60pj7yoVwMhBl
eoFQkm+zFs98bSUB4+y2pPrJmqjFtShhwegPaaGJ3unyfONiO1y3a6gs9e528vAU/Ylu78PUAywx
aqMdcKXGPEzpAzr7urkfctaSIDi5gTCYeMeCFQ4cq7BvGQl04XDSP7I0Zos5eo1Mgc3HYiARV6wZ
VdMz0LoCBaKboRIbiIv+93/O22rqIbY8ApIL7dYSgGrA03wexyZ8Qz/N+cDi/JEx+U6ah9TR2M3P
0XyrjhLrUCXKOb8xPOCJ3aztmCbMxpMW3CvneUlzQ21sMSqkBEuqnm+2AciKGbS7nwS9W3VXnyyI
EIMWHGgcTPose/02WeX2DRLyespzwxhKiv52INAkHC5W/pF7JFVFZKAZtn4pX4bjbaw5+ArzzHS/
KlV+buxOQfMuJ/w+PS/zk4vuaGCHrj3z6Oj8JVeZP1nQJYFZxyTNYAR1ZSbQNcJTzI+iRInmMRFm
o1DGHr3nZjjzuRXquezVV2PHTldAdO/cFMNEBGYLg3EWuLnhWoFcOOieXivNkYdd5gM0Hp48z5HF
UVk6Yy5pCPJCAsPSBdLrohMtHX7GxSp76kVUQGRgnMC0d3as1RChr4ddofvgHkVzsgPyVCGXxeoV
vgi0FEZqoIxGKXlaysaxvdMYJITwaHHRZbC9a4V56CgzEwYrUPAaPM4Oqqo2oyOJpPcet9Xn3r22
UTq7EJrSXccjJ9tFz7HAzLadIFi/xVnIWa1cITQmMy4UZfL4mzvGmi7IBkXR5hRjMwLF7vBLvyjB
FGoaynHyKIpz9LVWyOtasSWJ06mtFEV3IFHxW/vwgUWfCj7Jlm7Z0CLQhu/qCWTMy5Z+ZFv6UyaB
0cMHF6Vdwe3T1yFwH4ZEJxkd1BvkDMl260f/stOh6ElE/Q+UtkLIZOGvKn2ZXlTeKRz7b9nLt0wl
yPPVVtlxeNwUUCGY+n1o9ui3WHFbl1RgbZSXbm3X/bdg9Ymr9UCt0lyWnpQI0BGMRuv4kRGMnn84
mkhrXZehe5wWChZf0AJRaWQaQz0OKklJsNgHmrVTHlyT/NLwayeSJHO0lBeitIRATac5xLvXc1oF
oDFrotGSczeWysY5Og7POA0nigf381UEQ4uJu0VMUvDHdtqQCBgwO6t91RuoIybLuSw6DaaVqnQG
B+j527fkvt0UVk7fS95ECDe41TocMDaq/57Jz2P2X9xukpTBuYYoQiBA1Nt4i3vGFfBT8AgPS04m
S/QC6pCaKzKY95vNxPL/3hnZUOMCoB3bmT5sEPOerASVxkKUtx/P4aaC0/O1nQV+YUPQi2F+uvLN
XRw6Y77pEgy2K4+126KpXU2kN7hGTZcHC/OYh4KTVz9l6sQT1lP9fQoxdyBykeZOo1m1Dqe4YJi4
Fj83r2R/w8ga5pugwVMS7gckC7Ai0td1QeBbPbzNzBmf9nVN4v1YsSoWRftBWyxfbLbjNXilLfWk
amqdZfMGOhFlgW8RH3adshcKpw9Whcz+b/au6syflnds6wwv6vAyr5zSApQNIGZ+XqOkbyv/msde
n4r90JblzkomKIi4ZJn+BwA0MEqHQRLn5gYVcoG1ACXiXfFgjj2OrZNfyq8/w+o0oAZ6EchePdMG
bfdrTftccVXY4wDqgfR85I7U/HpEZfpvHPCitwwdWYX6M5g9DXNgcNbQhIcO3BhPtyaiPMb9rr+H
yBjZ+C6IhataOfU0K1TyiTr63pAgoaJAixuo09qVNP18VJIFAEoxe9+e0eVzxDrlrbzVwP2Z1J8Z
Eya8LPw/lo5EW4qAVYFq6Jt4FoBRDczKrYg52Z73Y5zsRSZslUWsEaSkrOdQH2aTpZZkQTwYsoQe
mob/ToYNxrzNILo1EV6pYfi4G5ZkyA91JG/NqLc45C8A8F8t+i6mrhJz2gidLlj/BRUXm+2kuh+P
hPFNBSx3Rmad+8cYwSQj3/DxHcRFBywvdhEwimNn1LC31ezGLQ5IQKcs6+OL0FUnYkb8FTbRpHWk
1fSZwKoKZ0CWnP/GPq0WoVQGwa0ovZVMA1dsDsOAd/7cYx53V/zvD5zzDC9/h4Rm0aJhyH+LN0Hb
r4ZizIMmDY2eei4uuUCh+Dmtzec7oXEcZKr7rF8NyX1ltzGsiiM1H+Vrevjh6E8hF0J0qoUDoM+u
k7lGwTy1bIFXx6ZYQWmghoXar0FDQOOTwucLLdUPk7ZWKJ/ErtDdjMuT4sxxtGQsmtY0ibr6X0V3
RBfNuHFr8LZa43eUigD+1RGONFbEw4dPtfO+5lACAVjH+kXB0eATMUppJfWYV73m7W889tRX9PlY
CqbaiEB8JijhuTNUsRZVK1vuNztFoQadfyOJLe499UfpskRLF/rVhvGAfIIo3hZjGRQdBtYjjskP
JqYogcrbi/0rr/GH/V4j9DMkBHCQHns6svhAvO3GVvOpXICY3BIUJtEjBMVFojGyiKe7khN6Wpe5
Enb8uTkG4hNchyoJHhKIRGLlupkgIdziiIphaGIxNAuKgMXuO2S7U426CIwgHcCA19n5JfVLm/27
H2xl9sFeIQ87L9T3K1UL2MQuQ+Szw507tlYB1YbkEoX4HcRbOyhavs+4yb+qg/DVurZjbTCi+Sdk
88mbvesblFKD+d6Ih+T8i4IyFr+68Wz142RmS9q5wm82iQ1JLBrGU71xNUF8qFJvEMwjU3gLS0u9
Dk//bXLEVfkjrl+NVDm6Md7hqKag8s4zkC2qUi8kkBjZOVDRrFOgEAPj/hD/QCluwcbSXxTIU40n
aNCRFGY+TKTLbnWivDgM4R4jCoqH4pdq4d6HnJsFIPBKxIWZKL8BHeoXg6eK/Skkzx1l2hBPMGJq
IQSOOQIVjVsfpGSrISg2opjVqt40yMkSTHEA+xvFkKQWkUX4o/uNDA4H7ImXYQfM4w2ysft/VDK/
mlTqHdw2zCFQjEDgEDz/CP9ThEoQdo4/zaeZ/l+dF+YI8Qy00oOSYvc63vVjISIcyrJfTALhsy3K
3Kqz8tVfkpetubM2op2hTiCur0i9vwkrvgwBdehNse7l663WO6yv5OeDypjnh+/CihREpn1B4eP/
HoL+mmBpTI9VnradxYrJwiF6FaUNCOm1Q712P3EOJCF7GBu88VMZiBm5BN60JDyFNPWmXZ9oF/OK
e+pNxmwuUTrR+Knhj/vNkvlcLoGo7VqAzrPSLGWRe5qrVb99x681LbWYME2HLFSrouNG+iOU0J/S
HnvAZbN+SfUKu9Wx7KHm1jo3mq++dvyKt0UAMEFaKIVJZ1pIS4MsmtFfkDc6YQTpihuq/abxficY
I1JfKUpvLW7qfk6dRry9cgbg1giIQmGXloN9c7Nx6LUaNEZ65wuybH46xF7MtTcBYFdS/y4jTIEW
q/U5t9FFrxnze2xOMwSrPKTgI2HAi/F48LsfwO/hTOXx4ok6WWIfyJk3bqAVXYXK/CDT2tHRWr9D
D0Qm8hynNs8bBrI7XEVbKvdzjxGuZHWjT/ljC3DfaOZt1bBxfl82cIbM1IoA9GmUne4eGbmbl8Kq
2S9xABUcWXyxqXbwH6MyQc8tl0Fo95Os6KrfDoxlqImFt7/Eg3e13CudPWRP7TqJfNX81Mio/goM
VfEeFy8zg6c+6yyOBxZYmGurf87OzJb+QfLxSsRh+V/0aFiqk1HQVgkBQw8U7NdmOT3aDE88bBWf
rkieUrI8wESDLXenVcrSLrGFzrtytYC3O76PysgZZ7mQymHWmyN7S1rxBMcIC1u3rUzH4/KpCPna
vhWEL7bRO7pLmQ++epRv5sfz8XEUoxacou2ipY6KZoAYvI5AREcF73ExIFyA2Mlr1EvjcThjRGAB
28zt7aRJOovp55nV7NpEV2ak8G+zVlgn1qSbXeL/Ht9TjyZJYhOle1Lzc/15r+sz+T6oVXHPfPaU
+eQan7IhlsBabIRPk7t+jLSEY9T8+LKJmTo6yEjAlx7NQcsXNEdCg/n2/Cbgu7azPN7tRvH17d5h
k+pDEGXVJjFG9iQ9Lieq/aD34ILgd0S91vh3HKI+i/3yR+gTtMt43kCTUn7jB9/ZsbOwywQNJOVY
qoHdG1X+Vi8tE/uwHabemY0OFsoj5A/gnwYdbdkEO7I0iUZ0xjCraOHyasMv9xEGb6rjXKlXeDAC
vAvh4hYCJKV3Jw1m0YJjxpBAHPu8BFAp5vmNJc/W8KPJv4R/Yv7obKdMQM+D5PFw7idAvtob+BAO
yizZ9+AhGZt8cFdA6CSKfkehuqWniMnU5RAL8Q1ZkveY0o0cRRqsJ7Oei1KRnaeFIdpVh1bekeGt
o+lIx1lHa9ldfBg4fdJKPIVy2MwPvuWTckM7Ghd7Z+kiiaJX65ywNsdECp8BcC+3Y4VcKWpMvWO2
tErc6RAEXaTMfFVCC7rmIwajiFxcG+a0wwrtZWVVOlO+yOfEzeufKUtWtOHXdYQU+yw2DqmBMsK8
UHR42KI3ZEpuEoG753YRCZTIA40gGB2RxF9Bq8cHQgoRzvzZJmBwWVpSvO1TphYIt1g0gc4zU+QJ
zhVz1UIurscZKSN+cn5bdOb9u7D8D12zHkhp83RfVPY4yqVKxp2O63zMAC6jTbLNZDntfIDnkbO7
R/TtLsL8lBWacUDL2e6243WmoORGH15meqUghBDbsYvXUtH3/fUjOh1H8n1Vmx/nvACzqCeJSNAy
dQh4vtokg78AlegldfrWw3aJj5WC9s0lrEoegYyLfueprz/Tn3dEQCtPJ0UEEcJNE36SYVAkmvOL
WtDD7cnAo0+ZWYhE4mWbSU2wCSeDgsIT2oCg/uKV7u2D9e/6n0oCnTwAyJo5pFa7+ZiK/WNwzas/
g6YcFkbxTDmku7vJIu/8Ju7p7oEl6SSGrNgqsyKiHUdjy/XhmMDSY2Q4cTHNYTUuDEwvsMhOey2u
DmNEOLiWRciUTRFwU6P+6WmD1o7DoPs0ngwpHxKO9Hl3DiyHLGovY0GLEnWBuLoRhyNVWxAiU9aC
zl/emZm72P+vak5gdV7ataABJA6LNlSSCLZssqL/ZDv+2B3kz0WsSXyrgccQZfBGncr9Rnsx3CkR
e6lkqrQPs7RrrrsGhdgw5ayapWbRATTBd36GQivqVwPA56U4OHe0KI8xX/veHRriGGn2TqdrXeZw
mDTDMDLCT7wtrdSaiHwcY/+rAxq7nz2TCgHOlxAegdr6kFKcWbxmC+4zRshiMokjK3ztFG60bECI
kVjzGYRVoLnhQFTKhQUIRd/eKTK+2Ykrnl48vsRgv15O4dr6QIyn7EwH3HOWPxQH9NXFmvcMqOLE
dlKvZXVI/JDJCDBpI6N3YZaLTjNEGxPlkqLZUEZeOa6vrR8VysL13IybcgGyffJZK7NxSQuVcBW9
STXr5plkH9Ciw2sIf6eVXXPrzsQGkpn9YaGblx/I7joOUMaVCnP0YL6b8qhbVnewTh4DMnNB+o1E
V7kr+j25y4ZB9bYbzJP/Kye8MMz70aEonB4gEKJ8I+1FP4Q1SCw6U4AOulDwTGD7vTPWRpp/9NH+
vWxPMIczbjxClkIIQlx1+qJhDm1AK+Zihceaq2PHyrjd425XsAJPUkZ8YpR4wChTQDdxC2ajWkF1
+bMGyV/a70hEM69CrHCoicc284Yadv0i55DN/iVginNh/94wrmSLqxDs3milr2vcNqf8Y+a+6iat
7EgF0YzXooniZY+efcjJfLUGZELAKBMxUCkfWjt9wRpzGoqp5fLurAfGNodWX6HbvXDdbMSRPwXl
/pZN1vSM3irRB6SUW9iO7skwnb2LeHZg/ACEagSdkmrR5fbICRr0ZYnmjOZIg+HWDSpz0OYPb0AK
9CeiISVmknt10WFaEF29kLHCYHpcIq0Ti6INHfeA3l7p0PB1ffe8UYgaDuCuXhP+GLCM/wnS5zmY
LeJgHFbc5rCBXDNJnD4ZaB/y4kYY764RW0imbNbcUndBa/IfAo1HgZ36teY9gkrSOCH3QLM019RN
V9vx5UYvs9uIJz4TbNGZjnrtXqqhFh8F2nW+4uh9OQVf4+zhD54CBzQpqiwIl8BYVQJvtR2/B9BY
16TGcZkPnFIeZZgOLwt9DerbMLPfI+c4kRv9sCcc+1TOrIa5ENZBt7Ugh3CcFPcFtV0oGLrbayJO
Lpw6oUwH0clb/b0gakzTtnIX7GMS7RzpPE5w8C7oaYZdnwO4KVGu4XrJASsTEktRKDjdhKqCPv7Q
NEU5ECXe2Okp0caR1yq5HyGV9Tr6TblHkChOvpJTHbUYNJuN4XFPZ+m/y8TmFg6iXnEzb5pHoiBR
py3VM9vN9jOACrA2WEiWDLzE4ZgeKZQzqHPWMGJlImC2nn/ojF3N+eVm3S/GEzpQMqfJY3+t/P60
wHZSsArFAZY0eTqUWek1NvclLThBGjFJvVIj+kDjEt6PCp+ZNkNl4Yel4avqAnfcfuij/4NCNPSG
cEV1nEbH6Lbjn/v8me40PbpIKwQdAMRumwYC1wwtPyB7fS+b5l4RpIuxrkeiFk+0v+IhLZn50NG6
430fdJlWaS3GLHiaH6iyMKu73qW/zaDIAmocVrWxGDkTUUwblOG4mgl2cZs4eqOqEjL+wgD5mkgR
DHraDtnU9EejPwMwaUaG3Igqo3U9oCHjA1r6GhPKMdn8SVgYBSj/sN81pmXqueZmGPOuopA0OHoH
4Io0D+Nf5rJwCb5IdH6CCIW6bHtdNm5JE8F8H2EUTHn2x2gdHD2FxGQlgM/7CIlNWv2ceFinyJhq
LiVcMFutcvouc+K9WvneOH0y6/xCphjvQN8W3No03qoJJ7753Yl5pGLhrY3P75FNFQL6Kgj1p5DF
e0iJKyhW4RDM67DG60jA1IpbzZYbJ29X743YL3qmUNDzpMOGh+hWRb6WFRsg87QNFu+68hVvVK8Y
Z/1sRWDRyCg0kdQZ6V9uKOC6ZoZQ9MUU+Tf/OoqF8zRTC6h8rsgzn/vO94F9GRuUnzCp8qovD6yf
qoASWXRoOs78ta3SpYJ4jKnLzucn3u8S0tJ0JdqvqesoAMC+5Y4xezhRzyuDwP7o1yf/ye/uXt6M
v7wUXtuTuU4jYmD+uIk4jusLsx2tEBe6AqkrkWJ8MxWcIwxo//KBOC0jipvCMmqtijjUmjnpHpDg
XZ0EdwbNsIzlAoyqDTSuqQcMOrT/9ORyyBlGP4nVikVXhlQAwqDzbgVV2TE4IkyX+QELhopcTxMQ
OfuBt+gFhT+Vgo9yw0F+IPBqvRvSBova1ss+V1g4IAFkWysS+u/MuTqWLdoAoFp2ZKKWPD3JY45q
8siLuOMlvKsko7aW7ffnbdZx+ClNDeCA+GY7RefshNh3lqvbq7OUqqAdzzTiH3zczY4wF01KbPEl
InFGMYRR8SM+tRPIZy3ks5lFUh+GueFgHyFCfDbuogf1WA+X5IJRfZmRSMH6fUqmxQdLfsmFm5mc
+4Jdh5KR2XjQcPQtsPBvoOM5scn6zTQw46k0t+UhORBpNcgnoVOHEKQLplprwqzsHKNp5ehK8pH9
m3HJDXccJssPrEXDFGFPE5JOFfFXNKDCfxdjqlKTz2Ffd5/R2tDpdIIwH8N4zB3SlIDqzQkgpK6T
o0Jts8L3M1Ee7ObyqAj6zQSOHscdK2DhtpcWUK484SO9yx+Mu//uFKbyxvDRMU88UlDPOwp7S+yL
ShV5NStOjQ2Fmc6mBo7z0miWRuWWAt/9wjP39yjGiOpn7XonrmaDHqCYmqu8GLaSqzi+y2uNQYSH
ddckZeToANHvTk6QWkaJakFnNbrKPtxbevUo0vnoqmDjNqpXXDd/NIktkrLSerp1ZtmiFHaV6dMO
eXhAP4MTgACCGM2cFQriaPhzp6CAO99S443gnWpYJlbtNjJA1NhHelXJJEQNpRiJE+VR6ZB777+M
ZMST3tU6XAjKcjFEdIWbsDkCalggWH1KOOCyk+TlLWA7wteWQC2YzNFb/ZIOyNoWqU8PJp7Oe5Bt
R/9WjuVUAnP2oKPKkQgVe1bxXAUvWnaf6wnBzYixO8RkUbaWkLeXwvf4NZtv/dYHFM8Y3XWq9pts
X366yqAoOwfpuyE9sBt8DJWVpuj7CHRvBCEGPvj+vRc9BVR6xN+WBG8oTJycAVbH5mVsbytEHHaf
ZEJ7XSLmzsciCehS3UgDFQPtJ5SAFYIzLGC1BIR32Sk4vK2CfV5t8o9pPrCt1SGQGmrWsR8QPZug
yALuOGa5gu7yK1RE6Tb8kprkiOKb0IGd5UgOZlwZBZ/lQWl91IyNxoaOsI5ALBzrCY1lF2byt/e/
h5nMjPfRLx4zZfTaBvuYzunEPw2kT49u5AWqYxtSk664NLymK6SM9afSzCI9pL9BSPp7yU3Fxule
1VABk8lJEfCjEFGy2GP9MV0oRLRm2u0kEJqq9fAX2j7RWI7zUosShBwjx4TKsYeKBNrZiYvSTk04
xAi/bHu0mm+lLffFlvTple242gC9s47GeoggJMqR1XJiON4MHvGDMbwytHfKC1QlS1HfvUtpgfsf
rxwsaPk3J5LIzExpMJ/CeAa/x7v6M2bhSbGdV5CpoAxIKhVcWVNEpZvfHyItxli4gpHf5FC7R252
b2n2t/uBQ0mXJYXRhF/Pl/3w5F3YM8Kk4lZ7vQr/q2Ni8i2Zz/qInjgGJIR21Vo2tAe6/vUrlvRH
D/1owU42y5VF5WUjfpaGV+57BA9iKLKFXpvnQuokyLisqLNy0Uj2+cu/ye55hufCZJd2nYbKPe7s
oo/xb6lypDkevI9ye7baXLZ2zw+nKPRkMISVbcml8yn0xXA6A1xI//tASGd7S4AbbMplfYuSsXWp
6td182nc/aTtbH3Uab5VspnDVuSPWWIjqCtPho4OKwSappoQn20LZWQ2yIYRVTm1ciYG40AHfN0w
1iaxi4J6w5wFuNgIstd8PozmR/dEjtfrcRdD/V7fPF67F2xBuTaB8HZdOsFPd2r1miM1VeL1mSMo
cKV/2ZLdkNskyNiUXV18TDXSyajrxoRJdfkbUIsDmbVYwzWUU45hJk/RwMG65P0lQu4CsJQLwj6Q
LXOn9sQano2dKRgaWvTsbpKQazvKMmmgVLxaqPFb2+qhjmJOXM8vNCWBEBh8olKpcCeBQ+ULZ8Sm
RtgxTypGSwdXzhTOAGuDeyGPPdFJfZUVZAiMg3yb82hz68hW+T5sRRM0zL0hf+rvgimy/pmZxMXO
WX81/PGLRArJlecUqFcccZIyupkgN1t0QcfCoO3PwAelM83uJbRx970JH6nteYwqnktBbi66RjvQ
TAOmcdbw4CsVx0rf88CkEA/xnNG3ejygMGTYMCqCe/xpK1ctZtSRmNaWVEk5VHwqvBpz8GylXguh
6heKvkCiFyNr+nZ81bqu+KF7jd2m0MDpQbyba+irYbcir+MMMtu8NcSR63k/EEd9pt40bgWYJ/UO
dAkGubBB8OLFJzXj58b/el476SSx8EYI4LI6kj2CE+JfTexP1GgISxvEOFCBgCwX2E+0UesC7s8F
ZQAovUIe0q2oss7pUQrtJBbSTQToEz1ViUG5XJsDvBH+tvdr/0ETPQx0lLJOpMecb0CEuaM2yphs
DN1MvVewsMBILFYqbnVhEO2zOgdgvn3DPefXuNsaqVivfdMC5r4WszS/nCJPyuJ3hx5WEloo7cyP
PR97K+ZQ8+sY02ylp3C+PsyharCj5z8b8RygDnUaq3P53wthnB437s7uLUrZbuG4dMn3tBIfUCvD
49g3CSgdcl0wg8Ube0clMdiZZrs2aV4TVY/RlduP5cIYtLgFAnkjIJkzsA4fBSyy7Jc7gLzFOCjT
BigTN4vZtJSwyYTrN/kM3LgmaRmoR3UAGeIU1d2/b0a2RDd1/AnFY0+qofcnd4FKoNObOFkbZ2Ba
gujuLiWE9QajIESmJ/KBsuqytYPvLySKVwkXt+hi6ukNkbR8YStjRXqMVlgiVcqqA2sTGUAxiv+D
UDtO3Tttnc87YjnQz4UA5XclK7jf3YKmMYY1gOm2AskWjvFn9x3UfDXl7tfswKF7bpuV7RXgQmCn
bqmEatZBjnXMCssnnofJGEGK4OABI67BKIIH3PhtuuY/aXrECSB5Fm/c7kZeFlGQ4QXZbEsd3ehl
K63ulqYaoKpHTn66o2DOwYUD/0Niz5a3b0NQb+RuyeI/NoNIP77kKZ1NSJhmrWe/xNsPE6DZ5g+Y
rPyuX64PZbM9CJ+U/D4nMOaOE4z++DYT7nN8+Fj0/Gk+CbebBhyU0z9yoEECDqzIvoMS49wSETr7
sIzvDsUqSVTGRhBxcAzOiTg9QCxcW2H0vy3Q0Y1T/z2qeDyuNpmUPSeCWS5dtsnzI93u4L3whkHZ
AaVYA5uagP7HF2WCumQ+OJmCEkhdBuMstTCX8Hlov6m+Ud3PGS7jh5Njtng5NBh6gLeg6DrWEMn/
vYyGwRs3mvXcRx5swWH6Ornj6U69Rye0pjezqS4utbyzQCWH7rOmRgB9KctMNmLY2IPrZlbzDO+i
6QgTgxY7JUn2jezXm4G+qzTuBF4jDfihRc9hjiWLArwYI/EdCko2XujzYKFOQQnoADDuyFg4Y0ga
scodXesJjvt9v4peTVPapw4npoZwNJhKYM/yTsr2VoWRSkUX+7AA1AKP2nS8wYRwFa9/tzhBxso6
qrfRdBuGOQWrBenxf1d3lDZlehVrYJuT+aHgWDNPnNIqEVeAeAFmKoX3k5W1XdeOJRuXoNkVHHOF
RR3+ZHbycEMzfiBNdboDowqnagqcH+Slj/HKCgaNr7oUUkCk5i79wTu5o82XA4jXge18AylNsFUd
jTlaGR5VdKgkUpgoALhKLpszgznmFij3AkZU4hKKyBD83cre1MH5JW5pqCfQX0KEkjldlO9CLjsz
K0zqwCbI2YsjuO8pIqD3GATH2+9SYBZ5dnnUvKN2YsJ/1u6OBa3f5EUwVkhKGLXswPEcl7Fq1mAC
N8kpFHj7CzZwJX9uhuuWbdiJeJRiiawDntD3Xbo+9BcCVW2UsMPhym4p/OXqr8Y/jFrAweXzEgIH
7kYDXXXZrIekJF87vUUv9m7zFH3Qnq5iUjwpQlrP1vvDTpo+mL9pcerZGDRb5g62AtGkYmp/jAzz
2spOt5dq5/x+DynIo3Gbnau00d+OphrenCLlfjMcOh6JUrKrhqQ3i0yy6j7OtXJYIlQwYi/hlN8L
Es7Zw6e2h4ZK39d+HdTGxgYcjyoQkE4+b9Lst1D5cPChXjZFgBMrNlFd1xpCIcvoRwwi4EqC3MV/
Ha8SkYuq13rnBdRusFd6O7UPOhj81bUTxD/4PWG5qeNl2iFIAyUqfkNzB3aFDhhb96PC8gWZs9cK
21kZRF5Xgg7fUHc47kwEhI9ayWeBlSwNU72hmQuUlAX8Ngj4cJ8xCOOcBIPBbGF18DASR5qA05hE
7Tbsw4SeJhUf7aGWAly28cf19HiQCqPauTssk5exWCcK5KfwiPA6ezvN0wbCoTElo5R7EdDenJ53
9CwJdD/4HgYsfVi/9fBL3KwVIj8LHUyUz55gp2bb4S8bjTWai2HIl3UldzOyNdlhS3P8CNJFsg0z
ItS9hzhCrJ7dqfyJqoKgigeNOFf2kHJebSDG4hnL6c3bZ7bDbPbbrgYjPZqnBDO3LjulCReq/uq4
j9n1iFRfP+DWT1eqh3jxhXDqOpfLG1tnGVUihLZHyN/INvJVeumsZ/7o/tjTyFdemH18N9sUBRen
xWdcpUAiL2e6HfK3HEJW94WG0sZcoERDRMEtMFlqwu5ZsQM7F6lv8ORhXka9G3VaOGWCMp3orUh2
5tGVqZUPyQId4otqnztaCIWIy7lwj++7Ktann4FkaqBDL5WI+24mgkjksudZRgCKUkniYKl5XKqP
Xrv2wvoQ2Mm4gFR0TJ3wpKJ1d4TzXP4t3LZPKw3ZesvT2T1g69NI9q7A3VKWAJnXmPKGoryCtV3x
drM5yhSbHfjOexkaN2mIaJjMJR59BhMY1RfTZDhkPKXxyPAZnx4wRuuLjXdwbdKX2dqJDeUq5m9y
RsTwe/5hlTn3I10N9HVifNEzQWg5boWlASV8jhwDyGX0R/3Cdu6lOfd9EEJ137uhIzMTGBZqwgG7
421gihf0pFQ/z8yaaI5PrlS8NU1D4zRFsDBmG8eMk/V123Q/Jyr9ako1LAlZijLk1HIBC+48bjhy
4dLgUS4IrobJIKAjtBYW04Gr73Kx6i6c+R4JcVf8vni269XBTKy3vRHgv14ZjpJCYirU/W8isfeg
zT4yzOHP/0W6u4+siom2tDpAo2vhdtFO1m5PQlir0BN2V0LWj01GL2+f8B5q2B3X59mSuaiNhARz
oU9UDwIs4009hfLhVPDytGg6Pff64Ym+1y8Ht95YSXUXWGuu4mRO5jcatxiKKt9cPq//KgAohk1w
qjptWniqLGy2RvT7zF6Va/Ygnzj5bZLUAgPNHrxbKrTnS1z/dxw3thkVK/2Sm8LKkQTwmkYDvo6b
HWw/cJe0Mw/qpSBMjRhAx5d7zASMvMKvjAVeulwFHSQHRlaf7SB6yW6VL06lF1zZvEsM/EZyiBc5
J8HZ5qtkXPYAFTKkD6OFeCSifqygSco+lofAQF+5VNp8mpYK1Y+Qu7ZTWLtoS6TVEayJHLKzzrrO
ufX4F6pfHnSbTCYV7dAil/cmqZ6oWFdpeSi4lK+brdgkC/ZzlCcFweYvI6fhJjuphQq+XU7ojUEh
4girZyfefYhZIfJY2G0qqBshK9b954Ed8EwwO1Xq7phF198fJmzBJBkyPiUKD2cj/AncxZ/YzJLu
GiqHWH2Q4a+uC1bkjFtFbiffkrbdWZJDj5J0NKCFi/qHxRwhLIC+Z3pRGM/46T4dzHBnAVWMlNkH
CNsfEH3oRDlAW2HOLwJ8h+XUCPBl+MfLJMXmq7TPxRnwRBVHLyt4it/9LTFDcAR3TiOOvF6lWBC2
gBtZOZPnSsl0gLj2k57w9jfiD58obj+/YXo2djwC+EM1nJNrxLBaxgpXPYs/gKu4QluGsJU5y95L
ecuDeHIkpQELvR3P6tDb1pU6066VaBT5MT7pCpb0tUnHGt9by95MQsJd5yGN5J1NBb52HURiT9XD
d4IKm64O7zCFPlxpmCZSlrt5rpUcsmWxsaJd5DDOpionuAf0P387vsbS7FHaiQV8TX5yhP4P//m9
AwL8W+Pna0fLNPvJq6YociVZusPdJY15WuVjQBJh0EZ9xFGRIsjffqt1979we5hEdJwQuE/Hzn/2
nK6wFBMtaWSl7abjSpsRJuhqz7D3GHFamMoReH8mU8ekEwljbMsKguGBwgdkBxgWgbfCAPM9y2Hi
WKeC4bLoEW9w2PdD+JuAUwPLfB100YiIkByPyOvbGd+wwQfpyrpAGINiqnlGvmGS+hGvWZZPgJXr
sJ2mWwrWEHZyjWpVLuQ58LI/rjHdy4z5Dogx5iRdtikKPrQBuZZoL2vekmkCCvJGFU3t7XJsCokm
SidzIRqgkpWCUZItfLH658H1I12uj5N43y4sO1OCS3yHNI0BFp/46g+/Mi526WaKS2sU5RIaoUmI
NPn1lPLkRtfOlbF96Adu1ek5VQnZGHY+fKzK+kTOt8ZmXyXDBRDJ9WIxsYJSM4gigL6Rz9GjnPpR
Qf1PE87DJrFhAko9vEKRG4gVnmwwFA5WRFEiRxvYPNvlPW3kl6/Q5XkmHn9/OYj2tdj/UhpevdCb
2OQ709br+E7nqiJjok8NDBGfM7vpt7WcFGy12Dtr5oIzPirkWhD2kg7CMcPxm78Szf6layevy01t
SH/RWafnHSoBG7g6Ont72xllZLrnNHbPZbMCFJcelxbJ+B57TnVzEcikaUArlpjIrf+2KLL5ba6C
kuQtlMutEeVIdnNwfKzKXlUqdqWnHGcOGONedQmTWHOqV21RsDuWYxsG2MVLpK5KjrpnsQWoeU/k
7+LrmO954fhveqqEghe4xna4tKgRJJckRd0CAshQgCwWNoKcE+uy3W+N6iBWwwZlvfV1K+dAn5bx
Pq6spBmUb5ushyKjFSJ7+uFkf7b9XsZlvn4zQauRx2eZVOF6kUYmnXK/5aSqt2TfrRxxeIFw2vhA
ff3lXQ6g/zENYLFdzqVigQ8PiGnsSjkkU5Q3KNvTAT2zs6ANUDAqryixMBUBHUJiJYlGn5BvB+Fp
ZZnCSnKhuAyaFGI9fzUwcmcWB6N3LAvXD8FZMDjKflnFBAVHUqLMTjlX81gIFWXIoy+6TbfEy8oB
Iu97upYmzwF2cxxJsmeOa/4P53isddhT0qdDzFH+OnQbHejeIWqRQWBEk+dy45Ppa5EYXGOXmWRb
dZksNZGEhMqsDZ6BdEX+OnGpieHBMlPin5jy7p7DZ463itSXvwp0TEYSFz8pniYcYsvWbvQD86Gk
ebHhj3lsXq4uup5JF23ikgS/O/YyUDS6bjBBjEra/Y9fvWg6MVKqfjfA8a2D8LSGpthJDRsD9Fox
7hz7qCy/JuJk+WSvSz9bWWArtdev2FNtSPnbP/qaEdc3Ec4fYKP9dJqi4jXqcEGeaTRQIGL/OZLZ
QpU/Q++077hITNoUrisJEEcPp3bsqzGwVCYNU3qt1mDPJF8zPr8wneOULkTZwyhEOu2LufPaSk44
AcSyApKuFYeg/7gUhe3B1sBeJ4mVNKCNQKw3bxtC+PVLW8a9vgJwBy/+hR0ec2U2faAM+YqbA62Y
bJnCQ5nn93p6k745ir9wwuFEwPtBgAVNCX00T4aixIcS6ilAfVXA57fsnNoctTmizqvXPMAsF/7j
UvKEiGZPVRv+jw8ZI8s8+WCRnSybJ9IJQ/v7HIGlhbSisNE/BWn9Q970zMljiW2GQtOd5JGprI6t
arRR0EKVXXzfrkWYj4WyqQDHAouscfe0HXMn6VbMNVSPaCpFxmVPsvcKVWa6JbpxaylIb7Y/qt8h
MZ1dfo/j+G+1X++kHx2SxpiAqbI55mTXEpkP60H9rmPVDhQAUDETmsQUBc3E/GiG7asFLCIdGtm5
8+VOpdec3qSCvs54Zr8Y/XnCc9OseqDX2RKYQ7tBDB9eMA3KTYFAg3dhhxG/ha6efQiG6llkmTiM
ZtUUDKv4S0/bB4PhtuSU/tFxKd49alaw28bxdT+l6c7oILG3f7WPOz8pi77R2kPc5PKTvfAoDhou
NM0yjRzHMpbiQ/w6qJfIkHxSZLyC3b/POIz68ijSNHMOKMClGrPzQdNLcUAoFl9zx8RQrb/xK2kY
FKT7IH4Kb6VuKoSvZHRUTn+D0UFZsjK0jlHgTlkEhIs8StciiiLuoHwPs+fz6oRxjo7lZ5j2puqD
spBDCMM7lxi54VvjkLWSMuMKN4ukc25WZySu35iEV9EE7GaGjVoOWKpfPajBWctBaFhluubMi4Jh
4RAf4+g6fXVsuFOgA+VEfi1bB1p9nLtyB0NbeJ1gPJjM1LtcnNGlMXEG+xB8JTClmEVyjPGcb820
i738+lVtjs6xrV3HesWP0oNlW2EfTn6wpiU19m4o3CirTcXUTphepa4QFqF8jUqeUW8PWz1bphoa
P7BRoCAawDbqxSLg7Z78wgv0Qgh1UtoT5hkyXFC9Ldd5VjovRmMRDmAEz6jjcdAneCHH+DAARXxv
4LJKp2eMqwfj0f+ZqjSp2eGImX5o6Oa0Su14EkoEA6ZzziaENKWRUt8QXNbRtUlbPtohX3HKPIFZ
s+3IszGNbIeREzXgbGfCHn25mvO5uTmvrxmwEG3ouckb18150EinpPCn0JddPgDNdoIxh9/Ri+fX
cH1YikHjdj/7XaNx17PZltBMYF8oCBZnM/gajB8/Vqwi0Bh/75MX12rP+DAsPKTpBxXOU6OtZ1v/
jAvX+ujKBUB7Pkcqxwu5TZ8eKYpZ5a1W9RlW5wkuzt6CKCwbkPKHTsNtjT20YJrVqq28hWMGjiSG
l+tXJuog7fY1Nr0FQHMh5WG+KFTBUnpyTsh2zoeoEOzWcntgxw5d3Bl0oUdWdFniWMx6S5J9Y7RD
XJO4O+9x1xZmK1PTqbCR9GzGWkzeMe5f58mJ/qj5NbU+aAE896Ct6bo3diZ15PBw2C8bu0YXJyx4
GcqVs1IE/QoBiwV7S0eQwT5alVuOx4+mGSUEf4cgqSfzBTmMD65558D1uJFLJOdx8KAq8X5Ecx+i
ojds+iVfuOso9cGb+C614MEv0a6+jqXOc/PrRxXJ9Sft7F2j43a5BXooWwEePdqP0nj21qmhRc3L
RNoZzXgE8qbLTPetrOpz0S9Wn4yVotz2xHt57r2gNzMTIeWW/Pi2VaskSomrhC4Unb4e2uRuTB0c
CSJaCQU9J3KQKFeI+Z+NJCkHkHfsDVQQt00IorkqVtBZ9KJyMoxOvVuz+jzzc511AgGvOO1Z31CG
Fs7BKafGGT7F4wZkiVMqJfoTELxZnPbQS2C0QCTUMyKcmz7mKP2s5zMH+CZL86x1rvW9vOcNYAlO
MF5ZqLxubZUoKMCGhGFsYe7hDBJSmMDX7lK5RHb+VD8EpL5XI6boUcHokVrGJJdAlGU7YIxD/zZS
6G8lbye40jJ8qJHhYfiv++S76syOR+fIDNmyxy1Vu6rNzMOJzOpr7a1K18yuCigUFRdKXA648WYv
mY1I7DwTS9J4X72ow7Dr6PtXT8duf/2mpVAI9YU+BI69c6uLhG5SIoh5JYnwDnbHEBEur0IKMBl1
JyH4+sySHqCD21DgHWfdYETrD6W1yGYsWYMrGo6h04Jr6p1bcwlgIfxA0oGYzq3hnid8KM3iR4hq
Igq916b44dhmbJKptjOe92SMULxzskzRN4OOG813HnYdapWuX/v6frRKMpZcBdQU1KbnmYkbkxl0
a7f4W4p0gOK/ieUH5cvMgemwHbp7GPVx/nyxnCWbMs2Tuwdeo3J5TcDhq5JP33OvpQnQkZX/HBi6
oqdE5K2wqCW9BFlpGtvIDpDtXLbs3l89+eScZf2zJDFmbu2d4qy8+BLn1tiHZMPTMl9ff6oNLg25
7mcjbbXHy620sRJhJLh3wDrTphB1UXZ6fTO2ypmfJlFpdRe99AsxttlDYYoRIANYly8zOe/EklLW
pa2IbIYRsqaLU9e//Xe8LFvJs98zY+jpT3ykBkmbcqM3Ezkf87irIMQSxCd1ykeINV/czYWC12zR
XvnbTzxXMqnO7fQ9duHFT9ozx82159kmM+9dfPdHQDm2iYdJtYtzMxcfCw9vRqxM+kmln8Xr+L/g
M2YIdGrUJjTs/GaPn/TlhLkJr2Cc3SJ0IqHFbXIzUBAk7GjpAofknyQirTnei7hH9cd5JmKbVjhl
DJ9NANOHNQK3s6t5bPW+1h8pPgfWRFl8w6KN5e2h4Du42ETQY6M2e4lY73u6JsC+oeJzEuhFGheP
RV3C6hMSKI67xd2X3Mxbm+grurvICqeCUW6Fx4Zjx4BzZA6P5Y/GTq/p88JJECW3nAGJm9Yv1aG0
ToRkLJ5ymUYf9iBt8s4TkTjk97xwZHjZbgl4GSKSbPwMEnkr2afeIlKbzKmWgFevqBQcUwEwcYOs
jREYa3hWEcl1IY/Z3gNFzaOWGrfkiTilkT6Bt6Mk69CJp3mCJgP0JDizWnJOcBe7MLMw3PL8fu1/
JufhMBKAZbvuX/dMbgzu9knIQZRpzymxDs2FdzfujnEifpx4RS6EIe6dVwrGdaKYSjHQU07g/VSC
Fr5kowZFZUZ3FDczJxpXG6TymL6DiTvfxlLzbqSHrfoZU+mu7ITUC7wPYH5DCAgaOtD8hqhdErnh
3e61Ike/+hNRFzUtbJXaySKsTWCVng3tZy7ZcMhD90+mFUwF/T2LbJzqoNoEYjFKAWccLq8Ko9cK
g4p2/WplGPMsjz+P4KMPBiUhtRkoMpJqEmXU6wz3odqi+AEWFmOCLjkak2nd+uiiUVkcBKBvG8rL
lOqIGt+Dv7FZ28RNo/yTWvdWW5MQpKsUK3aPFJPipDNzOBbzNoIQw+oWyYX8bnzbdchEpEt12/+o
/uNi/ZoAvD9ZOHy9vbClA/+NXXAZuJCN5kcFTogmbbLFm/DlSN+0qALAekjI6jxc+QMGArRJZxzF
SP+SkZb3YXMTkO0PqR/J2DmW/5hZFWpLM7YwvAqCuZBnHLZ1DSh/wDClNU3kj4kcjtlW9sY0wWIQ
3llP0PDxRFLgTwq/kVxGDQQh0oH5+CwSoiq3a+scu1ITIkBlVJHRCxp7+ls4YF90ZDGttxuwOQv7
0LrDlFEdhaHZhLxBIO6Lb+ikCH0JMwAybC0xZOjkhdfbRnz6tgKTAPgfrfsp4ghiLwGjxFneYjfn
z3rHZkR+98yU7kzBz7TTgM21qcAx5vMm8R9wmmJC0lVkj/rgkqvpw3iT0uR7vJvJgC1ulEl10Mba
DtgfdEC7cw+06Js8s4vJw2SE9uXTrnLBKSw7NLZdLyo8PAmAkF7YUoPVIXu3qT65Z0c0EiiO1Zoe
F8PFvCY92pOe1Nz7A+U5yMDdAUflVZ4CtpVXatCWDH4B2oYm0/GNrNl1GwE+3hZtcC8N6jUjbpZQ
3nfJcMWNNznDAIijVQlv65j2DKO8MHaLm6Zl8mEm15XKELg3MMvgalFzAr5xn2cp+QIiucYdZz08
7cDH3EUveAKBbg9AjSSXg4cM5uIm2H9NTDmc6uD+VKPs/qC8bQeJ8RmaJHXJ5AuaaLxu3uxZbra9
Y93HRWAobIq4BgSW5nmMzepFe4xAhJ4yGzV4gRa/ZYVItfpkPmxf2U24bxwYNfC8tjee2+Ig6rTg
t/W75KmI5ZTSH1Xoalx63Ih6OUlnW82/oVR1cGw/WKCInrv+GgXYaznqxQLFcExcR5Kyy/IDkj34
vxecVTguDNxFU+IB+h+az2ttEB5XhS/0oOsSO07ZsyQPrLeC5X6VkoqpbzDpMpjG0DBB5C9BrO7Z
76+2QlYMligkHXzIY6hg28LMLnNYk5iTwvWfnj7zUmGVFucmxbkIUODygaQBLrstBwkLIatIZ8iL
9MBobpuaC8PQmcQ11KlbAZ70J9s8cIqL6x0+XUmvZTdOgk5bt0tG+sA+edcKP8QhJfrCfs8n6i20
i7X2THpmLlohNT0MWR/vGg7tO7eZXdvO+p4AuKBWFHl1f2gR5kZJLChkPuTFtDW5sV/b7y0uNRY+
Ga6ZnN2BHb1+2PbAoI7oidf9ZThjHjI8m8hmnA6z9S+ZuaL/dPDbKD+nWpOA+yNc56YWyUxFZcGT
/JpImbnvKh5cudziq/9byOJNKrmkKxzI+R7EeIogos0nn/rvF4IcMV0nXVUzaWfk2G4/YZzWIkew
ASWKDvs37OdWxrxH36jVJi2T5DNXjZnQdkApbET7AVGscMyn7mqXZPUY5aljnIcv+c5G2ESaOPkb
m1O8mGhkDRFLoKNOkm+jybiQrdHURoW8vPQs9ZKjQbBwhB/aFBWuh2cYGN7HpnSnbUk+dn7iBkhq
rbXMf0fFrKsQaMoYRHr5JA8e334SeHJmJjSTAV/Y36e6FiMh01ZZ4ZI3a7cQ+w/7KppJXMMSc9Jl
+ik/hUqbHG+lZm2JrQIGoXvJeNGLUNcoSJkQ8doZleldItU5/j+EF4cMwBVbXXhANr07e2WBzLIl
OAyXA5L1J28YjxPfoigKkURQaj+aFxHf3qkoUZsam0HSV86TnKg5qXjJphf5yeVotDOjzytjVdSr
MnkIZn3CCy+4TsZjMuSMLwEhqeAjNqCZ7mneXpF079kQt6pJbiOqbwc9LQGZj3dCR3iD9dNylz6T
SWEXUmXwXufr9JjS6HFYqAVDWQqjAUCffKf1ybElIDh5uzpIkYgyAqIUI9XPCLQf6QqRjY+yKMpY
0XgsKOhuOrw45OXMbXSs0D5OOxVKvyo3egTYQ2KDjplMQd+ufEb0t342FbmlM5ayaQvx8FWcua0H
kQv2z8sMYxb3EeoaIan8ct/6aVEDUtgHlCi2iKqPUaonlWDuEqW2XsOyWIq14sl6UA48DKnTKpWP
M/nLtgeHF/ylekU7Apnm0isE2IaEQtZuMJQBXod0Ru/l6WIb1MncLa44Sv6ggOWfIvwOTyT6yGGW
t9OxciighAJCfMV6jwWTG9Q7IC6qsvGiFIdzvUPXh7QrZTs5gb0xjZixzYiDtMnKGwUMgGnrGIUi
HdgzxVDzfKFaQsnanLlQkC2dCihdBgKOqPFBrPfyvH0Sr/7XcQbWinwPiLt2XQGGowWRlkPVfbdZ
GwABbQIX4DT2Zt0kfTMNUNVJ0utoys4ZiQATzPCdxohQ+45bp7pA/3R32hzQcqzKBijorVSF2RY4
BcjCFZ45Ldspe5OXvchKBnh5Qx+nwZxiN+y+s0UNjNz4rJGKC7t+gwr1oeOAo5vu7A1vvE5jOHIi
afRgMzkllhkQFh7ZXO/2gyoWJQ4d9vGbzIwkYMXuF0Mn1DvgLsAMOEdThNKf8JLqBCp14rAFgG6s
xGEPiW62dRC5GeRTUs8dKSTkjuWFsLmxradYfqCSp4l5nqd1QPJ3QaT3dl+Bk6BOodP47YhLJJ/5
XrFxqVx3rUrC5sQ2VzD1F7aXUwuc0t5/c1gswJjf7O7CM/eXcoZAae8O8/cg3Pp9Id2OMRB75jdM
i/DR52UViogBtuMwVjfGInOoyy4I+bColN+oHjNXr6mWyaUhkU9lVkkAwpBJCkNQPNL+AXHsiWpg
VJNPyZdCR/9NgEbXoeVz5XfCAxg0sdv24noLu0ZhuNLBulctLZdB+mxHYHgxqzUjmkzgZl+C2f6O
Hx37znClHZ6+K4bM6Z3qvZ55wzSo/rou7r01qP1s/50ECGYL9/stpg/l01RjTEOPi5c46ZqsU9rq
RMiHA6h0vPkp/5C5JDGyjPxQoiSdNABrxR/x6u2lDtxNPuk97eNinhxMU8yfYi/5sAzsUk7tREYx
4/JV27RzVih0Wb0AN3ECUAOS81O9BIRVeniDXz/Sunin+xNDK8VowA9LjQI8G89Opz43yttnaxDy
GgeNgXIMINorrcCyWLhoW5Yt0iARB3bS1u+nLA0MRSXljTtIDuVfz6sIYCp4cVV1g6w7tLSUXYIs
96fBxXcwT27tDUIkclkux2UBRzIfuNJK5OTsj03tl5F2S+5NUztCurCrCBOQFChcdSsBXdYA/fE1
Qd5dyg0SAFHeg1Jvul6Rok60CuCAOg7zKRUWaP7XppjI8PkqZEEKtO629gf9zWFj+HDN0JxIAHyv
dxc64thqNntLGLDsMr/4L91Bw+yLbrFokexu67lOZvhLVkgL0O1VeZXoCd4TbPN4Q+DW5oHcvVWc
lJ6fYlbqYxjhW9FMrkYae4LtTJYMDCrurMaKqiGvPnwNx7WcAWOgqdk0YDStHzFIqr2UgLgIQz+Z
+i9xH0HPpYkhTL6ziF2O7vov8utqdkdeSv56+oiBZG4qYc7WlOCEAOcghz/nEldnrM1VXMPXwClC
9sqkZG20Llq+0BU6gqAy17KZEkHUj4TzJvOspmi117mXlkHe81tA6oqKBC6prLB0OgSTUnUwtcSq
yb5vXmO004DmbKauA7w50fOW4k4LXPiHqryIXQOaqnIjuoy6syjYdJOeUabYuxl/ywyqCjdef4Dv
ri3oLQZ4bUILTB+9pHBxO8cN14CVZy/wzMfeFXGL1pJxueGJwg3y7v8gpgRoW7XuA5TtanWcgVN2
FCRmU4G7mNxwg+w+aJ47+qmmvu9uoF5KtEIyL31Nu6rHeMF8BOJrfBUS6jqfkNdO4SWYUNdDgTmI
enG2WbLedDTXQRiz5WDAAfqpRtuEWllXOCDdQZ1egojumc1LlcbPERK3uyfXOn3wfDS8Xbfo2z6R
F4tFEcpLl8jWp8vxlYMnPi9LBsoqq/CSlqb7cs7H0HlU11sJMrM1BSjIYBWxQwq6c3GV9c/Z48K+
ZkP/bBu08TgxDWQKo91MxzyjMhqh31sKjsCkFPXbDXjV6wnv4vdY3qH6mbQFkm9WfALrCBpZwbMB
fxN2x3pup/Ai/P2lNmqRSTN4g0WfOOIcBTE9GtYhRHqcOtwdemxZZoOX5gmcWU2Ala3JI1qeovQA
cSToZvgtBCkrf41jBo1xdpfgED2P3UE6kVz6Fy/1/cXPC2bVJgHkStssVKAf3FQ48xxFDhqCq6ve
PeRPx7RB7ZWmMBP0FvC8RfwDn8kZjB1OUVGbs/rygLxj/o/BgjDjNv2L1u4M0HvluIPdLTz1z10j
pXp6VcBRFn+UySqZ59zWgD3H2QJ2MfEnD72kRRMuMe7MKKQAm0YOFFTRsnPVZNM0jZTTbtRBtC6t
56P1z6Gt9ZUZSc3IvddHDcEwyqeXYmm753KMzFFcJ6acWj6sL7fUCl2Lp2qop8AGHoR52fqJqo8l
0vy5jCJRvfqOLrZ/cTD0h/888TOZ/zlbUTsXdyGHiv8f9min9YCGn0NZv95TvDJ+ZuoOQUqv9gJN
3pM98y3b0gfF8jv+5BvNLihEC9LcAP0fUH/y2vJY3ZR3zc9yomSy09H8HWnLgqJwizjg5mkuDYlL
3AAhv5QcWpFCSXdKB/teWdz0i7vmumKsJh1oHsy6VQc3MkoGi5CnDzFNDxm8m2cBGUx8/zeCQ0fG
lYVJxA3pZ2agAfNtzCXjzP1IO/4tRsBND1Cy4hv9qPjAth9BjZw4Mfq9+Y1gs18epVztRgfqv2g3
905L64AdCBC5KP5+gY+RAWzH4M8KGqJ5C3RP+0GoEHGJ1vVyPpIxzGNm/XGPXcLHvLgvpMqmsegh
DMmLL2JXEY9Uvb5RwZ149LzaGMXX2NLKW/jJd9fzCM5cQNzSutB6YfMnweyDTcy9x96I3hPzJfrX
T/flaOszNeypbdmwTXuTzNv9FC3TaQUd070Ay2p9eB35lBcFN2TnxndtRGsfVDqxMevQ72eJ1OGk
TlCfW6noCF9TgX7zfwOXhqJHEe+1LKYpSsmviNqO1w+3nvZiF7m1JL79nT353wJfabDE9rJbqTaf
Lg4G90EJ6XAtpijt/K1rZUDNQsA8HBVHpygIi8PRmRxdq/18RVEZo8vqI4RcQDAIRi7pXZImUU02
KXD0F625ja/zDNoKku/KwiN4iSdwYrVmpqDdGpxoEoBM++ReImR2ly2tyLDvcSedaEWcRSbSgyIX
vmKLZCim8Bk7Wj8YBz3P+g55ozmfqvuz+iBsD5ZkjTqCnZukLdzALI6ulrLoX5sHNX2qbOIVoEc7
rVEpyuAQmq9JHXfnQ8zXxwDU2mIBhNLHvRiO0lWRz0JiBrW8Bqjh4FTD0hZ66IBhSAG5eRDf74Ka
jv13C5WPVDXYkT40ixI4sPHzGElmVwdSgQ4OOO6JAIYmoRc6gyzG49A0gbAzmlar0aYfYVuJr75h
n/3SmhT8yeU9Dxc1Yrj27BmclY9Hm1lLvvLFrmVF5hUZhV88+zEeEgb6XwbL/n1U0S/sJ8Qb9qw1
OX0E2Kzeij66Eb4Kmg4swMbHsafx7abD897fSl9Qk5WPFApQAmZ0YZNtNQelp2IdpeP2Q50hsgZU
z1ugtXVVKWbjn67drgo0ql/5Nq3HwnBF5iuRh7UKXLl66WCDGM48DYkcIF9O4dHmQ0j84kvqbBlM
jURRmv2LAiymTt2q+eUT44nguRugf99y2U1dfD6pChrtlQsNIojv/Mcf2f0GtBrl4niLvVD3YRZV
AfAEdaqfYpDub5Jg/2VkaE6Alsz1P3TYJG53/WNXI45HYii2grpppMCHcYCHeFqkLipq39LCF5MY
alkMCG5DjSRPd20lWBx+LecziF089iSenLvxN2vfWNwF+CUiBYbKmjV6Wgnc9aEFP2az0++SAp0N
QJwxLqweXZOdxj0Rx4JGNIEup+eS0Zvc9DDPY6l/zfez71ydXLdSGVqq/eNxWJ/8Pg0l1YT7q0aC
gH/A/wLeCUzDTjUxuYJmw2ouVBimzqaGfbywLflK8dMZnOSRRjGjyvr38Tyw89aTE90Bbn6V4WVH
3OWAMk6asM1tJ6Ji/LZIkouvz8HhGji7DSQa1MO8dUcu5A4msYs1ehsWVedHPr/KbhsMKfYnOz/B
JhzgXyxSmC1G23aoIOpEuyL67wlfXCtu41M3itW57Xbi1zWZtVBWFrH62q4el8otRseTnr4eg7Cv
td/Muk2r62OUnu0XPI5xy8jBYUHpF4XlTc20hwHIbm2shDpZKltI7S51+6WQuqDXO/esu8WeXO5k
DeWXpG/JrvVilMLBMuDL78bpqVqOCZFtNN85uyyvyo+TEdjiMpoFdZzivAFwS6SHNu9vIFcFaOL8
VRbD61i/WL6Iq/ea4oUtTkYlxOjC52YpUGgrMGAVvyG0lJaTVz0G2UCW5KwAa8MQHrlx8Zt0mayE
XmLte0BY61PhjzlcOCOoJ4mAswVL9ZvAr+ZsZDE0c9vyyl4eAbitwj02jiEd4zk/lGKwVcvBEDc5
cNC/BwKQJ1GUhX0VZPe4MOCkHEIz7KkxjQIzq6jO2GfrW970fyGQwHdO0DjcvpYvDDXyH37EssCP
71BQliI4KGSiL4GuwJVasFkqaWMifbFrXXCchVW7muqM0YcFROlCkvARTtkuAljgzeWq5URojbnK
c+VDkrb2fVhP1DHA09wq3ytD+9BqmCyllkzT8ZegbLLDzWmqMYUMuHPrqjX7DqCXsSXHoL0VMvZH
Fj62QEj3wA9YmmwAAec6mahOhMXeB7T2Aa5ly4D6craucgx/961HvH+fY+2HlO9VxODjDJiWaEv2
d8Jxh4m766d/JpNT7ls/pSROLxD+40tPBXq80Zx+AAvUzZaba7uFHCG8HIVIEr5/t8UaCFo9SyLB
JPrkJVhuY8pxamHWCaZHn2twlVSpW5SXecgfFCpPx3nmc8PhpofvH0n954RGvlDRb1nHNW7HCqm+
hDu5mHT6i1tt7BAV3VTJaEKWALqwLet05WscN6fJvVQZkLFFCdEhxb2+TXRSggWFwMRC2PQOps/e
Cr0pGwQSbA5SDnQUwxJcqTjs8jj8edsQJSTQCWIEyDiKnnfz+kkE+QQmQhcrIlViSvu+CPn065Q3
464U48eH0m61mOQt5O1ozTB/sKAu/guLh/oGvTeG0bhAaMXJhemuY1f8mcM7it3Ch7yTRiAlFQrM
WvSWLC4E0o2dmCdcinwkssMr3+HWJMzLtByUnBKfK6OPm2jeKGUCYIw/uOirR+YDxhUMeuesQDPI
fcBfeCKEcBQBRU55xLIOivdzIZbA8htQVkSfAQjMVWedRv/ncOGrjkpcQkVwcV6SOiWeo6YBsKM1
VlGxE3MW6GsjcBMunYWfYDAmigaqxgoHd+UMHj+4jnUnMT9iCTBW1oDa9X0YUoonmi1TfRlIVI1u
BzgcuSbBNzcn0L5e9w/xIH1+dqcRmKL/bvwQDhbYsbSX8t5bMYkRq59si90IDEekhKTEmwbb4Bo9
lzhjV4UgUFDpNoOFBfVdkNSa85nS/86Zbp/y4Ih8ve3LA6KO+wUfV1vXQZPwLD9jx4Rlg4AhzN8h
YllPWuq7JuyHO8Sj21UFl+xGiYvLG32f/PidYHBxHUHVRYUVud4n8vxav5/LgAqGGIfMllWz6ahx
dKTBn6m5c5E1cwAgwiWJFd4SmsqMfKdey5QThRcsnD1wXHw/AZ8ksgEiUd7d0L7lPQywdTp5JJwD
PXPWrUksX2y+wZ1Gkg09Csk2cWrx1GvTxh42B4uJaztjbYvSmpczLpVTCy3pXQp92Aqk5rB799rr
4DUHH1h+woYxy9A5erAx5m2eEnmGGYZ4nHtYWvr+mqmoU4Cx2vd3MmWOHAxIAcg8sd8VQ2JQFTRF
yT2RCWIVY3KvFN72lTCj+Ilgtviuz3cbThYpyeojzqgS8/u0cEgyguXBnvq7KGwx9HFwJksav72d
PHFgXUUuLJXQJA/3kbuHPWKpiMGqncLX7fbV9X8Vno/Cg0rEvZZ8tW5AYsOnMse+0EoYK30uQxf6
pYi0PU8FJZDcTeNjy9pMxYA1eL+0x0hhu+5w9axUZBSwAPlrvFMgoUmFBCYc80yitrfitlgx1You
yYJxxvqT3IWUaBgx8QcaPFQjuXMcyyHgnN8AGP5+XNgLUVqXI/YygvHdBhAdrNxZqT5JYKlilsx8
v3z6LKxPEUIzHTTMOBsklrPd6iiKeaR2gGvVouLTCHJ9PzD3xK58/7Clgz8WVrDck4/b59MndrxF
0Vv1JWhz6+sDSAqCJxlQ0pyztrwPVTimHalMzNjPrQuaYAbYLv3w7MOC8j2PJ7986eCoDqleDKv3
zDVdDFVcwuMZ94utT0WMYef8Qk+brbT+Sht8Pc4RM3p7B210ahyrwXHVcce4U4KtsZpABMx4/LoG
A0gwNwq+M0S89Rn/WGPIBUBCsduSJrySsIZMdGOV1dCLvumZXG4wMy2STNeC11T0vCRwldLQzkNS
S5Am8Xs32MWIa/aQM/GWG9EKVEQFRFAL9vUti31DjzFMAU2H23mM/nVbnnrRTe9ZkYM6kqorxBso
IKew/MgdVCBwvnxvY0+fu5yje/ggqu41A2T0LfQHYFo0tVSjYozCFF/Qgs/Ps09BTBF62RbV8Oc5
eEhHhr3GQWp54J9jfjigGpHsksnmQiZ9ogSVmc+cC9yYztkMHAPsSYMGtn7i5D8//jcMdTLn6kTz
65wPzh0t84wJN8NaIOyznnvHsl+M0jIwXRaF2IDVCoaPxeVZt82uOl5mX7947BvuYjZZBzWfT46Z
jWGC8ovWmiROk4yJYl2nbq/QeSAKdZWvM9gg6ndQCdbtQkS3UkF/1uT7rc2HI0eNJJ3AzuVgZMhv
85qpshJFviexXhN11kE0GwwIHyQ8Hh7j29R+8wAe2qyVVPR8XvfeKLWXFtUO5WemonYv4B/a3S59
5X/ApcF0CFBQKW3AH2gGojiWUWMf70b9hJ0tPV0+2A9XpJ3HhDY4O2Ix8wD5045iBiqesKT/RW/9
CcVv7H68SdICaa9MzYUOKgJM6tLLfRlF7I6rQIb9dVYQJnhifovWW/89fY8QV1TepcZ0ViD2fkiZ
Iv7KJmhhua2aLeyoTOikGq0QrUVjgyjO2luRrax06a1pOTYPUuHYNh6gLr9UYjauETN10pIEXLgO
0aIHfmI2q5JXQY5bUWHmDb99VUACBmwprbh5MTq9RYi7HCc5Jz8JOzEs4ww760AFufa+u5yPR2sj
SpDTQlKFRluWKXysR0EL8e2eYWlKWGtQHyrzOxwhoK+e4f+1d0W5qsEwfTPhyiwWUuVGjlgB2/1i
OPKlxsokHtWa9+iWWNkSoBybt336lYcXOXQOzjxsc/WsgVDkX38eULa42ZOlWJPvIDC532uqeg1s
895/HQZ9puHgPQRLkuyyX2PXuRgXl/QsBPG9EsqwGEBPs2Sa4e1nEsxYyy23DYsY4cjLBjcgpzws
13V4BtrXI7Rx7a0qgVgMeMk3Cid/dP2Sph4/LPXfWAw4+QDm9wEBlBygIEWds3k3aA1Wi2jqOPZW
svxlFiXxeCvoHSsn1oCZ3ilmtBKB0514cDWSsZpcTMxfPaBKLkJaiPz9EfuNSJqGZrF5IcrhVbJW
/RJEOnxY27e4//X1Gmon3C9Kpv+M5nJe6L63dYL2l1ZBXwf2bTkf6gk5J//qSBXQMbevf5wtJJ2R
Qv0/tW2Z45fcQHXcR0R6QncoihZ8psOoAPsWD9yF4N7bI5i5k9kov7QyAGgeRgvKmQWlF/lHhE4G
mi6gajzrInF3JkyX+CB+b6rz8Gg0izbb0yVRwbA/XGJqnnXUad2lyWHPfmecnZw6EkwY8xOk+qZE
qlRfu8dAUMSfji+W96t/utHkAfscUt8s7aPWMoz8rSJZipznwmeGwq4lyU0WiQVu3Hw1BRhXIyVw
EyaDRQ7D5fN/WtHVxlOdmt5Rpppat9L8qvWifBrmCng/YgB3AQ6wms1oV4wRr7sL6qzR3M2p+y3b
3XFZ2AEDz6KkxMCBzJoNFR7TOoCARddoZ5ph/fZFWd4drBx96czftqpZLlmksfC5aS5vWex6fnNA
YuoiOlct6y7gqO2sllQYvQPOmEOHbXM+xsQuaadvZZy8E1fE7vWS0B20GH24pzylrKfIeopqg1q/
LQyv+Y5rsatcDm+M4QsUwipwGEwupZ/QercMbqRgQ2T9LKJFnYEGevaXL4nkdZku69QGMWy+p+d6
z4FCUuxq6l6QLnb9nZbuslmIoVF7LswtOfONSzwYTtXgMs5tCqgdX5XhBNYtbKZ3kULqmm0yQqB9
DOfhe4zJr94uJbZ3fJ80LvmFf+z1c6n34wlfgEHzX61w+vPAMkXy387/5P/XchiDMoE82PSi8fe/
dLW5e6A5q93zM9yNcqWlSr3JQy+jHWTBt0yeiFDAR1xxG454R18+PQK5lGZNX1x7KVB0Qwe0pHrr
eiUTtw/m3gE4a6F5yq4WmRflIf7/ogwa1tkrmZTDAPHeMv4u6aj9OqKTpbPmlwjt6dHRKll600q/
YaUcpELU5ZHFSEWXnSUoQuVKZ8vEJzQYJzBCVDiln09aMiU36EUGlrbXPIIhzJVIfx6R0kcJDFRL
+GLOPfBjPc5OwooLyYJXCpPIPub85fqjoD6gOeeJgncDf5iHnWdMjqhSrJbyiWM5zzzvRBl9os8I
4cOEuZ+wiZFhowtWmXFH3Lznsu8mw1VR0stoBwtsySW++DHR3xkXmUtvQ/LHv7BKBWnNzWIOuS0O
ervGzWmS/Jmta6J/bYZRzm9+yxTrIp+8dWpA7IyKGjYDgt81gl37uYOtBwSOzltFSySzy9fv6r2v
wyt+bvwP+TLC9NL/y/Qq37TR64CFp4Ww0FNKmRhlIoQXGIc5l4g1z2BH9ZHvZBGS/Sw+dTZLu9cu
MDW8sERVX0wT7pPOXsonDtaym210wVaYqqe4zpcXN4vTD3uZ45YxLXaXqQA/Dbi4l3a96pb0YvpJ
uVuApy0LU3X45ZN3RmAuyDxgP1/wqiLAdrwoDHsKtSnqYH9YjZac7PfGpuZdtB8oOqWuqjVkPQ5G
MqjJVpHiO0EGac7IQVrCzAckU2W2Oe/q7VY3Rh7gXoI5LfsjKkDfQwIURxsJc3R+QaQVgz25KdbL
jcJCnRnqCNKWWzUA4lkX2AmLXLECQqlWanHNReN6qbftYUcGfhuUKOPN+fDWIa4/6MypZyPCH0Iq
arD4bxvr2UIqoDf6KuBi1zpjn54FNNpEqwN2YlbXn28b21inptXRsZm7aTGO1wM+lzBaPtHrOdc4
FJvtN3wQi44k/t4odglEAsORu2fCSkbE5mODTwjl8+2pvGIs8wnx1H2Xn8ZeSmj1j9YfWimt0ogP
6jiSTbmRgLnH4O3wfC56ilxcn8XoPHgef2uTsmKOBGpYdMIlbvjmKLXJ1Fx0yxrlPjkwoDiKOFhR
OCDm5ZpKBfYcrrPx0sUmngBOON+dMVKbUv9mdYp6Ye5ox80hnkElxvCcxZ+xOFK3uVNc8JlaD+0D
Gq2HUroj8db3/EH4Hk2ThHo8qyWLpgFDyHpo0WgWr4lz/NkhOhOaB6vCYTJxIsjPYXc1ckSn+0os
j7/WpzL2ehrzPH7oyf6k+pIdtnlNmGLDxtg9AFerSC1OnNxrpv+vvLyRfOPKXaaaviIUPUDE48uV
kYAdCjdkbfyFSKLxjiTx3Fk/iHPbEft3zK2sGFNy4SaAkDmctJmGmUvwfxRamxpZEk+i8PlyzRWB
AU6SOHe/2iB2w/pRbNzzoPWK3gK5p2jpiiCl8ZA36sWcifY5dx8P2h3Ov86T+eHB+GcfRoqJ586u
YDnXoEb0U/+TNce/Tm5p2tnEIVL4CK5X3kIRwYOj/uB6mgQmItIuI7P3wLcH5h83hOEHYc99wAGZ
T8F5dAhd+CSesZUH6llKUnvy9f7DvVPdBHp6TcKnepU2vDNEUuUWjWUoHNSbSQhMrQbFFHRYRIbG
Wm7AKMERX5B8iKkxS7KrUCFuHZIk+okoVXmNR6GL139jHhDrv+Md8aGgXfctsGQcV4JGSk2AaF++
C1OmBJKgrmavl3Zd7NDmoVLlWUkphw3wTU4vF6bUHbA8FGhasaUJSAnwbDF1BUkNYEf/S+833ztf
Lw4nTucHylFszhNqGH/RKz7d1dFzvDXi2xvSwcq5LNVhrXYor3fE+EjRkE82DdigRSwY15W9hD8l
LeXmjZNKlrPGH+DHEsm3slizpBbpFLSHlNwFE0h1Pi7T6KpZktyTUo83cSDKYRgKc95e96GTqOoB
ErYfJBhW08iYClIeA6+nIuYJ9MunaSvZHw12me9fHILaXJquqZLormPuFS/JBhinR1VRcUVtN1Ir
zTzfuG/KTL6h1iTtbKr8eFt2XxiW+F8T+vjsTkFk98eE4NLLYICxg5n6t5c/gQfNuy7Y/uovYy4x
nL6FrJy1HbrZcPVK1IvZbIT2bY1dNnhEbwX/g0LThinBsvzcCfnZ7SzhT0NnZT2uGSSYYl2m4jSn
Z9GPerOHRRz9j28+1eursm1tslj2UjSkcj34Wn6+XoWYUd3RNR/ewAt66+pkUqVlf6DYQNCB9ZKN
RDMzF///GHY5lNzaWWeqUi0+X29suAeu4l3JTCiaAHOMFz2C7cjrw1xz59872nRh6Rbs6jj4/9Lu
K9poHdGjG23X1Ez5VGX24MyH0crhXbnZh6d7giElvG1LGfs0CcGuVrGPN/4YY7FBoEkpqM3ceVYU
lkgM49SOO4Da2CCXzMkvpWjdZSyFcotmU9TDXe+3BlCuM+G7yRnkde8m5TtMRuykwmz+VUY/SVPf
lI0nHBKZSFiLV1+BLUQ2ck3Diuv5kmf7EfL+ynJpzK9AWuYizEhXB+5BtZjtXqk4m71znb+Lj91C
RKMTPsw2X+hFTXCtpwUD+40aifhsTMhQMD1cUAWRqEVFUJzODEZXqtHMmNWlpbcb/Zq1Zun8oaF7
y5nb4XtgLxYadG2B8RxgxmBphZKydwIZb9blHK4zfvilMGk3k2a25YfB/1P3+g5t97HHL1coXdOe
su5nE2CYzSLnDJPV9oSxd3k3E9SVOlxz0sjzniPnzZvDUApjW03du0AiqXRfKmIu7IS3zLFMw/s/
seC3RdM3wjDpK+j78+ogo4hdphq4/624jndK4jPCliK9qehfemiYub/cyHGcNWDmTaHf+Qz/gbg6
iJBz04nOWKUDVxenXzx70C6TQMtUzk+a2Gae776iG6NJnslK/fQRkbBrbfMlwOTYYM3h3byv8MEH
7zcZVtXM/LNey/CCfYUN3l2rNWQ1uHvNKUaynPqJ7SpnS0uDwp87kEWcxgq1E3Z7QukFB3qLeXVL
kGZmh5pNC22bSdKWnbsIsH+Z6NQFpWQrz6JMwuNgK8shgLhuEQmVgd5zIkUigtIEdf7/pRTTONqg
6swvV7i4H/y9rzuTUMoFHRFRACxHiwIPca5Hn6m0rRwc10PWuFTj4ZaLwcrlbh45QmYI69K/e/2e
NKB374O91klWgHLqInAFYjlMo5AV39XFbAVNUEjaPMP0+0FSK9EReYuqAZGRkl4G+mR/h5l79XE9
TAHhXpGWgCgqIDd8aER9Mimq7fCuSqBvUkjyp0HpurAFZQ4O10duNa2ACtXMAYBoysCk+Q8i2jMl
hnyfRSnhKHivpcQaiCHt4FeBXm1bFW49ryuoy/bZmEvpkkDcDmZNwC8Cy5kVCtpMGP+v2fHzmG98
1kybGxg/KSqkovb9g7u76sSH8JV52mLP0gss9FcB6td+oDNjhOkxZ1I/cQ853SjQPYhjqrfeyRJK
3KHV0rKTVnlHnLsK2Ol5CQul/Xx0iAYNVOOFP/G843HgR9riju4qaHpf8yHuXX9mrgcDJECrohJ0
Zo29eBeQj4Rw5oIupGcgeIe0a5TP1RfX8qsScxsQRZ08jThezAbAr5bWy56dGEIAiXfypML8w4iy
aL8+E58NnPBHrQErX+9qgCAPj669z00vAPhAT5QLISd9TOxRhI6TrNJA0C9Mc8sPHb/NaRzRdNf5
rv72j0qmhmToNmZD5foERdX6iPRbiXsx0sG/I3/fEaef2+0iT1wIjW1zww/giAxzts6I8VJsg6XX
5cyV9HcpAx1xGQbU0RthLGLBjkICxCrlTd/sflN1LhMwxWRjWAPbePBXtRmeQn7bOwPs78osU9GY
kjBha4VWlGcJ9dto+vthQh9+e/XLSAQZzhekY2fYSvMPZjz5rFkpJFiQeClrCkYhDF3L9yMFZg6w
aBTV3mRtzejdt2pGW/QN7iOrLp4kWbxFR9kgv6pOzPOp5bQOKKLlc2Pc4zgXOgI5O7eKTkiYzJYQ
jyBTcZ1MMPm0ZEzE2BjepGjX+g4xdt8JzF1nMsN3Zcxz46Ke85F0jMkXaTkntSQHhx1J7uMeHmxs
Y7VHjn4PHFjsJtfOOwWj9wGppK7JcOEbOKFLsKU43sAyD5npz2TUD4rzoazB354Yoyl0kGYden6r
AfGIvLpJPrtmjgPVpTVEbpryxZvwUZmx4uZFji+flPsprkFhdSMfHG0gGBFJgvFEtTjd5bv2Bf6N
Er9fT9NdZ1N+xA/vgaeAFE48YVUqu7MIXl72B4zbplGEItnNU4HKNsckiqutSULMep0hV7kLOoFX
jc7i5+4FbUu3fc7svZCajahIxZxSYpRDH8Q8t7skI4X10aSbLSfgx6YeDARIpwahRARBXRNwrUHv
OdqKTsaVLOFGQy2PvTGrOGHO+XMThf4qNUUl0LHMtwtGj5wox9D602GO80CvLwMDSPeviND0A4cj
Gn9fqssWG2WMmgBc1maV1iCn7xnNkhMfKAXQ36JbNM1IsffBscYbxNq/UDsZ6+PADC2xFxkppnpo
mJwVgS1z9HGWBtl1SJ7f3OQqMNBPGeIPuyV/xsdcJGGq5pFm8ADRp89NZjz7k7KkBKdY+hWXI6/C
WpIDxdLIN0civZ9jGR+wccK45oPJLrLrvQef7nXEhGJNmoe9CmCpMhDZRWp1hDWbWJgKGZVUES2g
zp+dpiuE3+qOHc0X3oER9fly63SaVmK4amo3WSn0O9W5DXxiUtsjAr20WrtVGobb2wHmloarpyBI
D9qB5HnPGoHTYOU2cHoh4ZoftjyqcBesYt3qbZ3xfyPV13bAsYzM3UzSItf/pGg/gxBPsb8uaBr2
QT0KOsWRbLkUs+iEyZkUelKApkdu69V0lRNcsD1+oH14HyS4AynfcdwNFUHG62oJKUAwQrBUuj16
u4MTdvpSWGm6PhqfdRSbg4r9gXn4uDlmAcy2CbLIVCat98YcA/LcL5lgDUPOCbvDREIG3HcSDWrY
cxVU8NGs1/4XbXXXyYg+dMy+OMjy0h15pV5SWeRXaF9WysUroSSWr4XbH9SSXILMPk0XN3g/Bc/d
1VNIzO5s31bbIUqfIeiVxq1BnSmDAJNVViffWUmVLWt5JT1k+87TzOQtlDkT+6YrhADg6o1LkOPy
rPotWaZyk5szyfYu+T5supgCdlljFrKyyRIaeYiFqrvAREUyBd5hlVSYPn0lP31qsd4mXEWXIbv6
rIeWO5EBxE7c160HdOnHoxNVs5ikCIokbLNELkY5afS3qH0QDPR3Bit8sClL18NcUptKK/ioh7Ui
1DWFiwUm63CW8g3eXM77mPsDizfJ3F2YOI+N75CHJWGaPS1KgUG8PruBRp5xhqJnsou4/epF645W
O3RRLk+CWY1JLlYnY31LYTslZHsGrnwh7MrJPyMCDEcN+Xly9M+FCeMmT79Y0BR1Csx88WU5OEnI
G8+Ms5owIfqZE421FJWqmscgXgOWEnQ41zSceBQ1Xmf6zIrujXYBo/6tSpKaa8jrTw3/kcxD+2tC
CKvRO5nQLfzoVk69mw31mm4mzuh0859Qp5pu18RWZJMo1OcgBjehjSa086bU5NTiGvnH4u8L7elI
tXHzDL0DX4rES1XeV+GjY0dSprewrSaLu6w9IAT3U4rHbuYvnP4heVHrZxN5shyb9oJcZN5MbA20
3gLehB4Q5HMdBQuXaxGiZYtBeUzEdPUIkyHb8subAXJ3eaCg8o3Nlb607bcmV9u473OfyHszd2bb
SzpwySKM0UVy+eIDreOiJTk+a93kt07joSeOTwtvOK24K9SJ1BhTpGUNtVLJe2zNDHaHL5sn15zn
WgKW6C33CHFx/VJKbiYHAzEUXUiFrG8OjPeifhTOSGIvXSOM1oyRB4xY+6frU2lHyo5+xLuhuvia
VLfuU7mIGbx35Xe7Pt2dLfmHxHuI3LYw8RkZNL4k8R3a+3rSobl7D8D6jOH9j7qdUmiNZCfg93J5
AtYYWZoefjDWezOmKKuEToJ39ZXIUjByvraPewlqecF3MHXXUQvejy93JR9X6p0r4hLlpUC844IJ
8R/psACVXQD+SGMEB/hfRGB7qUg/NJOLcWd/gf09KidaMTnothUmpiHnE4rSZNSz1cvg8JSR0HMy
Q/t5LxJTEsvobniDpdbqKR5vWE2S6fRw9xccm2WeCZNq+PMmwkdaxlhHEx24L/dHFbH/5to+sJzu
blFyWIlCKAkMLkxMgLjPKSuOSnhLl58PNqlrgypI/6cyCt/BRBSbYfcwJQ5yNGKaeGZyEmRIWcOb
FhnZWMgmzb3R8bcLld2IcBeaqNOrZrslVmvy+gxpj5nu/RWS9pdftELzHGP2li7Ke3EEO+ny6NaH
RmLgzNrKkqTvK2m7haWUT93q2sr2qz01xKulrAJtE8Vq8goubU/UEHrqvDlZGgpHOM0y+2FLheaL
ftbyPxE29ue+859yIx6p9Gt9vU2EOcSokA7PGQk3yI2WsjQDm7oXY+VDRbfPC1ojdUoH6h53Eg2t
O8i4SMUFU5YaQN3X6dPI+GzgoDYGjOlniUZ7Jh/54yoXL0wmrF7WxP0K9DmuEghGsfdmCt84NcCl
R+qMXrf24MlBwS4EyiF8domTZ52mugc8PqYuho1nSVUeLJuRmlEWAbu4+VSm+eLLWGPSYaxgkqRN
RGPpeAtb0aunWDQUCm3K6qxiGBj9iDR2NKZUJNrKMANcpt30c/vhpwdZlQPgZh35eTY6hT+XPDZf
Kq5faEd5NR6uuf3A6zcelwRR9LLwaCiDLIrTvXayBCmE9uDSLRc4Fki0VHJkTek/QaoZesrshAcU
lk8MZmBptphkvUnY3nkVKrzBSOLCeVQYvfs3dfp88Uyk3UoZQc5NW9FwBhNA8/WBFunxC4z8X+mZ
txIo582w/559mFiq7X+R6IA757v7vD9QjCcGZhTW6lMfV01+PZ9Hi2GaXBIm3Y/YnRgQ7fnpNqJH
9pJehqCqabt2EhjsiYJZU/MFWDLl7SAvIH8/HXNTzmkLxun9r2eOIB/3EBmBegKkcybYvq3b4T4K
ir7J6A/IQ1e8aYWWMYrKP5TrjaqAkvxkls3hPMp0Ln3OgnoPeueJqW3WYvyDfyfW4RTByHO9t2ig
V6pdRtCaG+Mo/jaf3/afTZs9rhdbpT8V06HLGP3hKWftTCs1/IrSz5jzD9jCMaQVdLKSbO1gBzVb
g8v0ad+58G+FbV5Xk0ItsCdnLvnNzEZGJaOau0IXjNDVgTnoJxeWlQR/AKJGRf9EQNZl72rZsRAP
XuA+CnfoeClHPaIxI/RKTj9YwXm9UV09dD+0zd65AHFOeAZxpPHjp6lu97kvsP5sKI7lWgjOJV/1
DnloNASD0lsCjsDWSQduxqLF3+IkbyN2FwGmnJbdtud0cs/sHEvdHMIZBchloprAuQi9ikSEDpH0
2ELR7pzUzr3nLjv/TqVHTNlh1wL50JBI4v5UA4eOvZvdCrV9UpEXPyqGlYthp/QqKFC39fpEJduQ
Fp6NwE7Vh0Rp/MFnSs3jd2Q5t4CMMBrg8vwW2RXCQ8KXYfysOd9jadeQBTvR3fCokmKCTGLVe6ZN
dYKMHmW34++WDdXZiDlicYzr4T91bcighb52xsTxW6PZkZBm4naisyns69c49iHOl7JsLWXOw75q
OgYF01Ozzv0X+7Q0nLOdNKd1nIasox8Zs/X9EWtp5lx2u3sVBf+nhw6Sr6s/vpCH15U9YVh8Hvfc
GYgNsjgp+JbJpl8dYAz7nd4iYhvWZkuoQ36Ff3vNga8ZyGyWrGD5OeQ29UQSXfmFJB9aABlqGHh3
LV/d1p1B+kLJb3PMiOBUeETcyMrslkfCBnG6K4CfqOC2w4ziL5p2rPttDKkspsfSmiikF6qDyejI
rNBrD7eF9ttt4YydUwHUjryBLreJXJJ3oTbYVSWo+Nu4/nAe+iIqwUFIz+d97J4tufeDeGaANj+h
WWhUSATD583JM38ZcmeSRecAh0H9oa7AuCPmTOvN8gW5xZXOCiw5j/n+AnrYrb+DvPMr+TM9mq6X
oUR1s4BcYsbZq1G3Sa8WtDs+r7Da1N8Q1qutOQKLodDnJ7xkb1m193VzJCsJUEDUKnxGME1qy+lr
olMDkRAe53SPtYXXn/wvO9MZXu5VNZFLN+/5Ob/A/kXWRS5Y8o62DMk2/61t3DO/oCFgYlYG2PQj
hQfed97u9cS90MLX3E74DfgvniJOdwNRiJKhTvhNcNggiduTlsxz43Zhgk53z3EIdIG6ldSITNrg
u/FrNfQNvLyNQWzJnuQYFtjL2yaLEkoCml1UBC5VTcdCUTEOCu9E1J5HnbIJYzGOPBtu/Rp1VeYl
zaZc4tJCaeY+dGv0cOQznic3duepzzCFrsu7ZU0LLUHAXsS2Ouk8KaYqi9vtzG8zV2X0pU6nTkmy
/Tm9ejYKNabnhyV5PMvxwAQ0FfFgd2qZc7+qjQ3n0faTp/JpNILRvUgVucB90qNbU//3Z9scfNM1
Ptnru99ZjQApYG5DjhiHip/Mg4V5fWg07uj6D9aXrtv2m5tEn2uUurrkY4EkNLpr/NQR+TCd5PpF
rR5hs+MyVTnN10bu+AO6wbpUgyJYuMdpeMUhQ6YKgRckNzaAGoRhuOJm6ZkBPiywUXPoJE8BnbtR
qz/l6ZDeQtgWuW0ONWtQcNGDnznTZZDwaZw2eFTaYju93XpXEmAxK2KoWI38alvCvnAopH2/3aUs
1zlkC0iT4RvDYs8CSopeOf5nkMMfytomv8+1lUOLvtIs3eTXN4jCT7HdIjrl2KersJQeN+vNJCvQ
BTs/EteGql0OUyu7+YCBbnmLbEVT0BxuHIfAldiCpyC44B+G7xSfOAY/k47eeBbO8UjU5coK+1Hl
5GyiiKMTGyN5C4K/C9HharWVSODWAEahNU/QG0bwWiJvDQmlMc1niuN1GUxStrTnoViehzhJg7B6
+uD0hBMbIoiLshJFI4sGCUrRYfxz4jzIGoTsrEUmlosNyuI+hXNrLcLG1MtciVCYGQ8dsuE5eP5W
hl0nxLrQcm7aSubsFvptG0yNuN4KOBs4vQvS+awblfCgtjMNVNLBzBchjQEJtlaiG0cd6Jnah81l
tLEZSEG7ORm0rFkXM4v9UptnfajbHdQBeFkwv4a80Vf7m0yJC6XwRx90q7xBgS/R+LU0wpXP9AZ9
TOhojns9yK+7QkQHQt+CRERpvjH3DOUa9/Izo2xEyLxtPEm2q5ii5mtXMLLgi7AJ7EA/wxsF3GXw
bxYc2pI6oabpu0Qln/4UBrRG8RHiLheK1/0fHhnYWFofXs7jEVZSYpTVmSZfCYGWIxS6FZ0BcegI
dhMpoWEE1G15Q6a1w1EDj9NL/vY5tCI7BHoWpHWou4jakQNprx+6YRtk5nzoEv24JAKKmsSbTpQP
Cn1BwiM8hANJSpWVhqOozEY6/6ilPkSbONnYrnOhUZEEfYbvOmDUxbkX5HDmJ77+hyoTjb33qBZ9
yE8OIKtmr+8vp+rKVv8ivwWedZkhRiMfYJb/TzMd821YLqcSSQYP5LJGtDicicP+wsoVmVc6AvZ6
tHLlMV3DYEyns7xLhoBGgSo9QIkH6ZeCgkbSBnEWHvc++JH45PRQ8KTtKnKvMynzUAFRTyB7ti2k
z2QstUq1xL7HIg3J6tLfD3EqJLHdoK0GJm4Rt3j4kYvR4+ef7tJMZO878IIjBQhzVXeDRlXr375L
ngQH89tyKcH5Ph9Lw9O+ZgXWTWx3w2MpRSOSgRAGkZZhlCx6SfETUbCtxZAxeT8nHcsRUxDsGKxd
WsqPZ6ZRWop9HVoWhyxQAYtieikRsmXibESfS431pLW3/rm5fDz43cmLZstUOmIb9fsvx4WJMnUN
I5KaRn1U5PDSh2WWTfq42n3xP9TegXIL3ijLTCTw0ArMUUoG2lwRR6LYHcraExjX2MvKa+mzwkYu
+cMegJOF1GyPAf1JUU6zzSR9uGQ3guNZnoPPhdRefGlA4b4fU4ZrSMex4Prhx9t/w+vek5w6Z/8P
u05S7+r/B9vEAHnrPZgcOxBguzFGnaKkGBPyAzqX6ja5kEcpUXNv362/eZrtcJyP1vdS0Bect1MB
azcqBjG/4aCsPAK/dnQBSQNqeS1TbVw6tjUtbeJ7l6eFe0lmEURIRGvzJ7ugaXmLI4oeR4s98UIn
bph5RP6cwEf4uUgBgCTEDj7VFj/xPjxh+D72Gzj4cpdqNmJmFOz/bLd/t56xVUjbRN5rQXPNtJHA
mR5zYVR2iM3ALmAk58v4IdNzznyat4bqOe7dlG1wl65p55qMsWrGduuuoz65zkq48irx/4C3Dcj4
yR+pnTNtu2z+F38rTCKlE5zR92h3p0Y/AjM1dboieQR1X0WTtkxTR2JSuOxk/UfyfQSvvK0HmvHx
/AyNY5EJZVGUjKjb//CRGfzaaATCiKANH5g7jgCxXXCTL8OVUj6hOefGQ8rRArSYb4Luw+2KV6SP
ZX+hDtQ4V070nbAHjHQhRVFX6deHia8e3KPXpxMb/qufC+YIv2j7TYRSxq8MfIwy5eezd3RE/ZSC
HQ7wQq1JJaXAoGn7b+ZW4hsNs8RUaIed3+khglYGygxwCeQ5uJt0IaR4OjAIvGN7TiFTJcAi4Hmh
ZcTC68pL6LU5i8mh996zP7LOnvPf8FhSnU+81zKqWtVcXu15nvw+oZqi9ZN2usx8LvwtMl1mYsyy
sZOSbMqF2D7iCUJl1vjlZ75gjBEk9oRbl6uPMPNZlIV1x4dkbCOiKj9/L4UOXzEeYZWIdcwbGbak
Mk9jRsvb4rTb8tcFHl3ZTy6CFsp6v/Xa4xPw0BzYfTheNiazrZFYelNyG+yQESc/gQ+BC3AfNXDx
y06I4goecJeoCLXs1MCwMsXyUFWYi07KyJNrl9LUoNPHhEVEJ2J884p4MjliEBAEAlXZeySyPw8o
aZPmmMsXAFeh2AhcI2Du1MWljl0oOxyUas6EEH5RIqbYwWqstg41fMAO9wWnIwjzKa97PL9+IEcA
i7yCiKF0OcduWCfCyN1jRYzKOzggcqjgEnVwqN2U3M9NagJ+h8cuE+rF4DIqa1Bb17BZdnL87EW7
liEx+nwOWzAwCTpIoZAWmkm3ufL4kgGB1NEQfhjSU9xTgLVCuObOylZtSt9ZP2/n7sPRGKCSYQBj
CQpndfElqg38JdMF+xMGRFsDy7LJuxTz3FkDTLcosJ6qJLP4nKH3jCP7g/JEEysuhMW6LEXgere3
cxmHi/Huk/HesDbtiud037rtuzLMBEHpbePYvRNRccudw/a0YE0J5+Qe2d+UMH+8RuMVJzfBB31G
ibokl9vMMDITpIcet1EPUcQOapyWZT7Q6vPTunMqGC5JFLfG74I9NtaCBGp+YB/JLtgkxWM2ug2y
DO7ecRM1XQV856trJxykGWcKBYz2onmpoBTAQugIgHsoiF9eovWM3VCt3FeO5Q/xNh8XyRAmevDO
MuBlsgrUVpnKWN7S4EZm2wJDoy7Ddkvl8wUhytgxjtc0NQyFBEZU7nhjsfHt0iYs5f+smwQj5wvA
HaXcGo0VdVHFQObjNrhX713cSmHObWnjQoBRO/5jVO55Wgqwm/InuWiy1eFGOpEkNDsKJNAeJD1h
6Js6Tdpc2glWhQzVJ6E7IyvE0WyN2hBXMhHgap5x6MEznKJW4tOgdoLjeV5I/JItF+AoU7eWg5lT
l5HOr/ROsX4O4Pvq02LBjdvU7RHCbhX6iMRb6B60v37giziRyKhrBMDpcdF7VUtrruyJj833hrmu
DwMXEaTf6Ur7QYT0ZB+1nwvpWiEE2XziCjWtUsKWLiKqf9ubPxp2nyPUmKzEYB4yXipB2NZqh6mJ
CQD2Y2bfcK+jGGpdIRPCre6bNrUU8RG921IwuL2cB4VobrdPuHEPRIUmAZVxqkj9I/N+kuuzw0NH
2/OZtKPSdDf+bpqvyxLcDtXdP2glHVG5TXAbaKansrDu1xWdpmvrq6wD5ZI89kNfYKfUJF4J3gWE
uYPzlFboFZ/x7h0X3LIijz/0vA4gqm3UiSZJDoT9n0gqVZK1JuvAGGhQXpkgSf3cidZ37ZZruRU1
tDjP17ByoVKhWy8oY0ehnPhReV2dUEGHZ1pY304BFZVnN4o1SVIOY8Q1aAIi4W2ST5WeaapP3zi3
VZQcXVb5jzzDd9kdCgxOjpouyRsb/uOxeeod6aSuHOUg5CvU78e+yVq8EbhZzFksr3V+MV1RAe9U
UWVC/FFov0FLZ71FmLq6Zgem+ijN7ZKM2bB3ivWXu9iXEh5eZ4YmH6fB+2enGMYj82rzT6AO82HU
ucmnCU7r5LL63V8ze5DyZ9u+9ZHqcVKntAhf0bWH4uNeu9y8OTqSEABM5qdBFuwHd9t6qiH3MrFF
hCTamHiaQEzcKqH9ucIUJ2ZHOs4Ob/kkryajlbDr/c6y8ELQ6LA2gF+7dXr93QaZCAerUv6AFYQ4
H6GoxxuaUmrcaAuvB08h/Ne5MBwga1lOWMggNnOOkBfeXusOVFBlqY0rS4i+nchQAXc6U6JOWZN5
l+Kw1XR4dreZkfLlP2mq2ODiSZeAhVUKPqjPAGCP4Ijt+3AJa7Yp343chD4dDAysYeYpz3jsbj8y
PP/13F4DuIvgRq2KEnw9+U/p3fjsYrJuSkxHlwpdNlodXLQzMGk6UxrIrzXgxOhwXgpR/kIqR13c
td6AoKP7S2PUV/h6kCBg391lXrql5T3zGQ+Z5rBy/Z8nUJRAtxFbqBwupOcJOxZLkX+/bJcJ/egU
mILNTs4dgcG8EFsUBmHe8P0+hvkSj8Z0LPKCHhHc/4roYZSl6bO84e9BHF93FeIDE8h7Ge61uTHM
7nAqNvFJH7opYxk7Wo1xplz3n/mRy9NTkdGl+iS7IpAmvR/hbx1swr6foK/kS/djAic6JnrGALu5
37pIxIEsPiugkIyYqHg5sIwkfLnL38j+nYwyLZbPotK6MD5oobsw98jYKp2v8xAX4DOzhrK9yUVq
vxW87WkZX8Wc4QBC/07xaqUpZBVg7/L3OOKHN3iIsEPCVvSZwMBcwubLznatsBZNCZ3+cfwEEFsP
dcPM4cO8YocUPhFFYCzs2twsTQr+yQRY1+RPwp05Nrq6auYUkoLYR5qgC/mNProUf9mHDHgjcYDf
W3abv3YngkWYUvhcePkTuCRrzCdmv7Vcc3z2jnZ95SWLI7Hxzzu0TtrrPJsusgs5t2V0h05LgOml
fJskNrKLKJxsER2+SJ/60GEaGQ4CBW/OF0hiT2gpJGTzytbDXm5FG4EUvdV/A2PSXKZ+vjxWy5AT
H4TeVebgNiBk/2rM6fDS3Dx5wJhkwgk8M8flGIIz+l6eNp6KVVyGRuzLMvwDZkqGMFjL66ti8FBb
n4tOx3wzE5EuTrhnOfXixfGW5+uzuQ8ei9Lc7jKQwpbZsDfFROzN6YFc/xSPCxZpKSHmDM0GfG9n
vN5gPU0QnO6HDMchH9Jjj1ECRkhv/3i/mHohJsRFlOpo+Wi7b98/1H9N07sTdSwN74HM4k2F409e
MgyXnzrZHirgYy8ucHAce8AHmAqlY3fDL8tmzD3+F8bHpERhLUuf27S+StRCVZc6nE49Tj3QsYFm
n65FTPyzaT639iLWMdlqbB2A9Xf+O6HkBL4sFFJ0+ZBfPAItLKzC4fTzSFCCjVwiRcaMEIyd1deK
CoySHpJROHvhUAnWp6LqBtnHDdT7V/5Dx/kRYyQZp/gR3N/jatR0BfNCNXO7x2nx/SGq73Tp6Nnj
QwC28/6+EA+lkiWnRbPMBJw+DL9XSaArCyQjRXRWO2k9ics7vRTR9GqSNcbnQdzsZckVHVDEy247
8sNvgV3jNQQkE3f4lQZUljI7YTIW0IecUBTDHEBMxj+s0Vsfa6ZbssCS5DuuLcnATZOJ/s4+wEdZ
HI1DhQcZasQ/yNEvIlXyXmJuGXqZMCK9XzViyx5lPtb8ORuKeU3vh7vIMrxzmDgEq4SNh/TP9Ilw
ZCQMGnc7ImooDTheL5KDCqAEdzNe2jPviW+gIvA+xHR/E4qrGoWXm9bvj6Wsk/C/pt9SPxQv2Osa
bE7iftoycRWV+auqjozh2tBzuijhyctoMZBQmVevaeSTQ9S4quJI4+Bu6FvX2A8XUoWZvJ8K8T2j
9rNzwCYPZDn/hYgO1xPfxMTyUylbOtE/eVRpLb8+B9hDoCKYb+CAtQY7jQ+scPhwuTYCyD/e1J/c
zz+ATLSbX8nrzFcYq8j1PsR7AMLAtiSc6QAzU+MRxQfLyHbEEUDLPA3vVcZdunBotFepBSXNMFff
JRLBvJEMlc5v6/1XIRTY9Cg7Yjz9hIPvY2LfbfjU9u/oEYMMB8VLy+u2BR8/dAi3ypFR02iD2HVn
rta1tBzDI0ry1Ba7fg/CJoWmkTG067Y8AjqQ04w3e+blB+4OVFSER1Wk0iEZ6WfD0zw87k015S0K
LVtxf0oMToA6lzg90NFmFjt6LCBPFQW4bZasdBcvjTwNJj3Sdk59p3yGbhKQ9JKMC2Zk29TRqPpu
0Ov5wclzP2qm/BFtEsqVY+tfEDnSnbrw7p9t2Yq6yndxVQhKgyjN0ElfYr9ZXz3YHGK8znXv+P7a
SPhDNK1GhLawYQuWa1lq4bUEm1GH4DnEYXjIS8aI2dCmRidZXs6lw8Z88CIlIF00syiEIzmWxcJD
webDxlXvPudtvH39ssJtX/BybD41AfHEkCS6OxCrpKias2gvmqUMjUYfIddvnAxRkSRSyNujwfwQ
/fcz7uvxLfW1P7StejSB9TClRba1yIXv+1FB4IFPFCmsNmXnOlwkiHKMvGD3Dai/3UKKYaGPR826
dDPMmHIH/GMj3n/UQaIDqm5w6/j5tM3AZGNWxh4gby+afMVH0u0PKFQws3HsFBi1o6uNjektuH1V
69iwt7QtlteUql0nCGOpQ3lW2RYGzUmcq9DM04kfYVTah3ZHTtjWRNPXhhae6Tb9EzR1PGkEPiOw
9/d2LhAtuhdTSAJzJWJltufFyYQQnYAleJgZKukQ+xDZXG+IY/Xv9D/nECx4Wwjvrh64o3JesT0u
wuNNbWwxFCab2HaWT4Ytfk5nRtanyZf0KVjahI83cXfPGdWCgjb+P+dUp81IsWiRXdatdruKTIvT
x8z+Y4Ea35gyAcMJsPR051PFufnTD4WoCf4xjopmPfSctGzrC+3lSStPKslY2h9r7YwZ3c1IGu2d
GOEHXkY3jf/Gh+Cv8xxDb4b6JIk0MqPXhkhBeSvLS/uIqNP5z9OWGTCFqwbQBMv2zeJJyzSdqY1u
Wa3scrW8VgyyG8I+bQ/cWZEbHyiIKoixNaSfl8oAAmuRXdtrHBnK7KU740KSRRM+oNygcUCfcQ9H
vBCMgJCAAxuo89d5sB4h1v89EzFrPX8QzVK24kLpbUmHvMCwVzL03ZjBQkdO7x85/wpcyAcElc6O
VGaEpJN8phRRjhv/NaZgFvBTS96MeLST0ektAKBm+NUfz9LNnycaiSrUAahAwhBBpnqjEj6tqskh
9iR7pS0naeGmC78Lniem3pHUmavvObeNW3c0uAFb+wSmgPDpRn1+yhHvolpldj2Al0faP5Yz1lV0
5IYcSxGSr7kadcOTNmYfVsPH7KoBRUX9xqABY5GVem1oRHMKQp1nIIuorHAi6PMkYSsakeX3mS0b
bsrDn+NVRzgIitygeCiw99kYnGb+BE01ZI9IEBiV9YR5yHMu9s4rPr+9DJFVeRXm5r5OdC17RJvn
ZHlB1aAmJvZP7WbJovbhcUoPDAvSwFgBQKenB0RoUwJmNwTNMbegnLdzC9O1wJYlkS2bAqt6sONP
jHzDqCt3HDBwaY9lvv15R5eKxY7GKySrJI1d1Em9BLI4/qBYnTOGyDnyNdhG6woTQzXH7ke/lwWu
vnVsw1KxprCesZQpdqVqAwely/6euie4t/5iRrZa2hK7CXvbFVBa+IdHGu2IdCspUwe7tBNSm0yO
ff/LnZ77aryp/wGXJjhp+JYACgOqy2b2FRDGGdvhfUpyGnEN2ELNLjgmfDUjqOhZl2ujfBnquJ+B
MwSQ6uz0R86yXdBgp8sVsPvmItkuV31vorTMDTUjl72cPiOMXxgPmReYbw0hjh6hcZhQXoaFiC85
Wwv/eze0sqSqYFatDWfI2VX+u6hPtgB62OfNewZOd+JRnha0PJn02lk/sIfqIq+2QNHkjY+saYx3
rwizA85B8prlgDoJ7Q+E5qVPqK52+oejFkaXxtJv8lSYyIrrfkMOi81S4QlTVJelG9dDamc85Xmw
3OP9AasvFPZpZSoTHpxUt11e0JQaNQUtncfcaBPuXwNCynlX4lGUjbfuYwXXWVC2UW5fbKKzJ11s
+tITPWxfeyJDfaRva/4bY7h4d/6mBa1k5N8cwGYR3+kCRLT5hgix0X96tl+pmICFpxSN3xbFzwoC
8jQnpVnYt73xhp4elFYZBjtkDygbvgftJiAv/1zdhuVz05SyWXwIG6jyobnQ6iNGh37AMnN5e43F
Bz5BTuxvVxFNM4tZ7byfxiUbGIdWa+Y8bGlDPAvMCFFn1tc6R9AvE4iWM5zFEcpBvNWOxDtmGWKN
VIP0eTIXS6ZfmRefaw92M5GWVzGjkEHT5C8/Ul+JhMZ9qLJukQpTeVlER4xoad423QHsBZT2wZQb
7GIN/I+12e+S2jZ93KXpT3wI+Dd0SRbIqs8OABr2eAFHlgpKi5kp5QuNg2rypKo57kbCHe3VzB1o
Oo+WKu8GBzmc9QjhFQydffVGPaPAOt/xbdBDuPfXpR8rgDRsdRr7Xx1ZgDoYZAFR7QSP2b7ADzuZ
9HtkmdEkS11ys4pDKt3gQNjPzsgUrbGXzh5wkboRkcI1tZH66ouv8OSLfeB7hLg8GvdNH47IzGHz
C0o5y6l+XQEqFknf2Jg0OjMMS0lPTn+b0ytheUp/XDhnan3VHK1tD86IUcXow39kwlxqK/RienTF
gaXV/Q6UgC6SJf5GmPXdhiziLmnp+DMjI7r742WWH4AIxWzI+8UH7iGa6lo1E4umQAndnagfUQd/
UG+p0FIPKF5w3nnsMhZgL/WKqgzoixeCudXCEG8eGShtNyw2Ifax67OpFyptGhZtOib7mKj4cpgk
tcrYttC3PStmBy630I9YQyITcfD90uguUC5EFKiPhAMUaDeLPT9tB7/DpDKEwkBs/AIjYvHit0rA
RCAA2RAMCyrPNf3qA5jFGhMeyPHLI8n4umjKNM93glmw+ziZXjUbYCQyMBOZXMfzKJ8mgTXOQaIF
HjzuKftqrVBJFREosyGj+/MGSyXYZiOuoMmw2AUVMGpcnGzB0WhZ5Gw8EVUj+Vloq27IUpt0gyY5
wix4S7VhYwVtqk9qQA/aroej1cAs24vYIgAVeEup1hVloBtRWCW7/Ya3GnKwDES6FyZLPswXwXLv
EJvjVZnpT5xEIRRrjIXZdKcLFjRNcfy0LK1gxA/wqB9YGzXtMes7Fuh+rMDZ9GzgIo+uuJWMxtVu
1wSwWqT4d3ETs1sv82hqZml8Q8R9CDte3c+mpvMZx/ZNyL0HsdsG4FSkYvv42Gg9fnP0nvjhoz/x
LNScxpwdrmqfJoC1/eF8IBLneTmoaO5NUJR668gQa+s3QfuSJAYB2KT998bZGW9pwnANgE/fAXAj
HHZWh4RlTc1PcrZdMpXeZNAUFzkHbZV6lizfdGmNEUu96Yo+dsrdZzxD1JlejzBa5t9EYAtbGjns
6ZyRkDcIeZYp7UaKF2cmK/9VerW+EOY4h5X41EIAxqGCiTXkmb/1Qo/Jzyr7gJU9Pf4HZ3Yb9NfX
9cScci+u/ey/cV62XJtWjXUTtIftl5eIJsYDN2qn7av5iXi5I7z6PikMS03osMk7ir5QYQEyGBeZ
aPo+QZO0RpjO+L2RA3db2vZ1MwTkbREV3SW55tRClgl2yupXbNpxgXhjpAHuScBNui1n7o06NJj/
SBxjHgUQ7Dk3MwC/fN1ilBHanub8jDhEl+JRE1/9MJ+2xnJPLdY1/J/06nYWVrymttDaXy/iGSdf
PoLL/YK0D6EEN1GMuhmKasG0xfbH0+gOA04qWvHyyv+SnGPseiQqjIS1tnxQNlHRWSfy0MTwqr+O
MaAfG36yxfxK/UCwkjCKtgAF1OPaBkuu79bET6ky8dI/pjJ0CmMlKWVKpLzOBQNCdPDDLo3CU1/T
RO14HIYw8lqgd7H6+y5nCObgfumThlLJW41K0NU0FMnbOaIVfzujaRpGbTqQRf571CxQMoCGDFRZ
EvI39q6pSAxVgbB34FzWL846ijSHdV0ALYnHtvF/cy2XfWwD4XDZDxlOREpkP5Wn+7nuPfL1E6kg
z4p9VIJ70QhEqFDTvmeRXjjZ+v/4Gk3YIdJRUytuqsPOL6wM59AqMYfrn4QmNauHDpvEJc0PQyjG
hBaIF8zOzgDfMDgFAV17Q2Vn80QS1dY4WUvxAtfQkk1wrckLNHmgXVl6oxUSUnIXB19j9aJKHbTF
Jv7Wfjb9HvXvLOf+Uo0paJVrdr+LDVgkK3SL9LjvyzPJNI1/gGsrXezNnxR/b1Lmfg3fwcurqrWC
oPWru3QxqyUzYxReLtxiNVLsAD7rosIh5n2ANfxX1ujrAmJoApHfxAl1Zq3x/KSMld5GElhgC8Ap
C9+KLU5jAA7Uqa3cS1mGNHQRc8c8EZrN+kC+rTNZ0X98vBdlLldOYZwm3YSzgv767+gWlYlOMNYm
0zXGbKQHG66nzNYhcxFg4jiSLnWYGGtv77IlbscCBv9uiLuqWJYJ7SZdLLOriG8hoXXGlxFPfp4T
9OEJ9GoPG3Eu59bbuLH0lErIaXjWlCogWQHwF6LB3IXtWLs7eFK6T300KKTsDg06wLmexs1/8agL
exvR7mT/o7RgD8nG9eqUdtoDWFZX2HQYk6CTj+bRJc6+Yrrc6pGQdZ/pzgLYnkWl4YKVyyaxElXo
mSIwRF64vNgCaQSX4280lGnWXbPPuGkgYYtgCCuUBP87Rt2Cjr2SPQXklDA05KfQPWN1rv3+pTsa
q7dVl+GTGZjRG5ZoWQUDGhgkEQafNp4KCgAOYovHKjS2QwgE8YBIKNADrc5eGxRMmqbqHRLxO0Th
5UvXQtNHWdFeHXooa9L2lfNK4eNhHiW21iQjd03Wucf3wzMf5ZR3uc25De0QF1XvrQ5BGJYoIpEi
TEHqhHZA8lf4fuyEARSqxKnOSUBasaFN5sn4L78ZI5EAyhd5mQBB74Edxd8DQUHVUjdZgtvr6f0L
4dbTN2K1YeMcUeAXAXHpsRmhoeKXQl7vhvgB6HpUm4OhoySCOsJqeWzJfL1CMkIvSxgFZEbLXmdn
BbXbv0A0vIG78KfKWTcjSyN7Zw6a/tKz31Zkl2r2aAsO7U0bVU0ejYy6TkqyuTifxP3zvrhIG2bC
zmjfav3n9TKgOYuTWHWlCyELhohrxaWMLsvXvU0D5z6dpLkQ9gNHVaWUfLl3hHhQ4jYjSk5uEAo3
ZdbT5QFd1ZYBBeMVjoRfGIRl+k/0qoZZPRyylqOJ0Yo6dBMvhOgv/v2XMBp0odN6/uw8Z9AKyWuQ
GSbwWheA7ZFg4VhW/Z1++C3Dqs4zrLKf4d9+NDzAtgk1uJUCHUy3OG52Dx9Wd8F2pQl8p3axtCPH
h9e75UL+NF13JMBD9Kkv0z9oFuAPlAoMZW0No+cMBxUy65bAt0VPvgc13yH/eewyiboSTpv/IQo3
JrlTXFI+mH4hN6E5vuHFEF1UOPBHw0BNUlSkF5Ubveae13o0fH+MAu6IF1bFO1wKjJlvAtopf5wq
fiaAIgGQmLA8Ec2KhVxkQKYZlFVWlHJdyv9X587fnChS9fX7Odp0DYrsxRAOCHxACtsoZwaXAdSc
qZ8blfdUzPx67aqREi4La+naflmWxohzoOFoZYGZoCEtkZzCkI+TBre5kp40kJ+GjjtNgTRFNwj0
XvjH5e/Q+sb1O5uOtQAdloCyvx1qG80eHEGjtG8wNc3An8atGWDzvayP23clx8izT4jzd0jXV7ox
onEvIN8WCxThSzs5nVd+Eape+oBP6xX4Yx5qQtq5efgJ+IFOuvBfKdz2C1iIC661l59dZvBBVUYR
wuAXQ2WYNJoLY9B2WWwAgbTFZdjoVXISQq+zTa1jNcO/onWJmPTCZklcfmQS1TDNYJ5z4SPvhptl
KzaZtqrRIZXP2lxre04dmtHUuM1IyPxFtqVLBAD6dbTt620Wky73G74tsqL5OHZfKy+4WmcPrbSI
tkofKRGq17cv7L60sc44z3FPjSeSPDHoPRxCmdDgD5tX7nd2iWKBWVXb+jbSvPok7oOKGHvdtnc3
SoyVq6PMSmKMioTbCsfqaqRvlWSNbuT4+sz3NqSaySl7YKmuUvvfwimG+H5KSqw4ZBsEAXbnFV+X
lBm/H9VjpqexUA0nLLWLbnVTpuu2rBsqDR0gykpTKUkrC6axZFde1dh0ePw40RZkvsglHTL2SAyX
BemhJrbOZ6q8Vd+GUciDVZWLgm5BjBPICkfBV2Q9OTGjt0Pu5j13e+V5sf8jsjieN76PbbzUCQ7c
saQnm2UU5Ro5mOgULx6Yxh9czg7HPA9z8c8nm9FVJBuO3jMqlhK4j/VXFYGbdZFVX0LF74viaItm
GqSvHjyOZVvrYeEZUiSqTedIpPSiZWB/yNbT0Jrv7fiLf3wuuorD5PozMDlL47/RFBzCsvzJrm/C
AlSmxUqS77YbySJIdQQEEImBAPqIO85Bs0s9nC1qy1Lt2BW91oKlJzH7wE844aBaxeU+1AGryEm6
W7y8nHjd/WvMLKpvIxORVWGfLeyn5SLpvSEKePaLvP7PfTwVe3MKeJTt3pcvKHvemRIvAGzUIL8j
hfq9tGYFNsOn9P2d0s8JDJwYoC2QiVgcUElwpq1B3m4dikdtDNxWUWY47qV+PLCpEQ8MnGRKKHT2
fhNSrStFwmxs2r0C7sT7pc6XYttlb4vBxYsSdQL5KUI98Mj34B3dhPn1stZ/lOo1FHRJWwor1ytp
uSOGLhanJQ0tvemqG7F1M9+kCL8X5XBQ2+pu7MjjR6hUbQ61DpdpjheZZ0OiUfoGCRx3wqzRfSOl
DpXZ/qvW3U4Je445SLHlWRpv0WCuzbAE1i0iQhlzAPcOv+N8ogMkbK01DHZvMkaw7UH6nE1tnS3Z
ZOGcybe6f4uiyTrVQM4T4Gs5qj2OPoN1yH3f35gyjli70OQ/BY2Esmmi7JCJiyuk4k7adDJm/NBl
6kdcz5Z5sNmUvAxUNZvtGjOiFD/ASYLChX5PpbpXviHRApbWOV5Of8s+h6sOz4hqmOqsr7IRHJ73
6OA139ebrJ8llzCmDcbVsuP/ctpi+MGQm6HTgqN+Bkp8lVAnj1Vh8IgD5ObTmbieb9YOz5vSWGs5
WYat4f1KK1ILyaXhzdOT0PwXtiKz9txn/nj+H34M9Bi+/lH4xYuHQEv9D/E4yK0ViV0Vs48wq13Y
PZi4mJwI2iPcvOcCbQYNhTYlOK16VlHmid4SsWewJVbIf3TPXgCEslskH+ZrtPe35ei3OHGOfWyD
s8nMl8TFfIW53Fyb2YwHWeYWFj+/hQiy+p03TPa9aM4TB0mqR0njAfz5m4ZqK3g+3rW+Cfrt/Plj
rs4ALJXhLWmZETVRzHxA+OdigbTwTm9EOZVxIpBHUxDftWEeDx5PqXo8gJBqLGi468eiq9gTqAZb
qfnQr03qnvlr9C8Crthe0g2oktW4qabVbW9Yw/JKCyJuKckTnfmcg/JXDRzf+PkVi0e+nkK3zIJi
Hxnh6Dkwfp5+tk51m+XXGonFPUvyoqpexTF0WkfzT3L0yv+DAAXk+THZ7fvRztFwo8DhC4EYUYrB
3Hln6P1Z9YlaF5/1MnVZjwSH63s5kmF4KO8nO36sAQmvFHCXzmOZ7ItoSRN4G6iCQ5LdsOZKbFi5
Qu7QNVdFefLgBc5Q1PfFVi6DD04sJ/lLDPBa6m3GppgItNlfbaXNawxJXhscysrAdLp0DdRVHz44
Ylr+DX8Ju5Z7ubmLoGAVs8mhPug729IneaJr780NfRPPVrKsA8CpBCz/FteW6j6N5h/vKEORlLU8
mzJBQEEIGdHv25MiId27lm6Z/F47MSg1QMcE9UOHlm8WCAxkXcu7tRZQxstHS1WLu1LWE7e9PJCa
6LFYRTF5SOQv43+c4kaCM4xPvS5B9ftsrCzH3In0xb5vwwBNKh1TB8zsyal+ANQOlzKPD+sP+W8R
S0nuIv+s3melrcfzEypLQVt0jlUcardgk9V2H8hpNTO+0oTX28K5A+ExpPQTGjoGaoUNjQs2hx2x
py5UXMJ0VbKKrPfodIKxJq8thHKpJ8js1p/tG79eahLOvR7NejzrGXBWCXo33N3gUmQjQCxnEAp/
G2hb06+dFUlsUggJR90I04mfe8APW+ex8JIdkVcQ1a6TbqKEnZqMK/tzzcaiGMBwH4qsA0UMdMF5
OYoNz9yccoSahHVLp79ggsK0gApJ9iuWhYLkFzHSHU6nRHYKckQjkezkvB3BSexj8RbkLjpl5GxL
UymQP2jf6liO3RGU/z4JLYbp3Jfzgm/GR2bZpXRoHuhYnaSJyUGryW/SdrF422qd1lXwVBFkSMjg
a1tIOHt9WS3/XrO0tCnSQTZvonsMCJgRImAGaZgsSHFwbudlOEB94nLhhr47yHIosCCOajTREmaw
pEQZqYCR+p9NpB7Ud2YWbjbomDqAcbwK3NaOh6cH3aTZ7iwjZLTGOgXH8EGruJRmy1VTQ/qZwU+Q
rRZkU042KTDg9pRNzyH2OrWlIHcnNpg0+ElTmqCYHIGj6oLM/Qf//q//mastPFaYTvyWhqMzxh+f
jn6GTzIgoBCJlalsuQhT0OLOmCiosI9kU6S11GdZIHn0X3Ngpd9CU5RNAFFihKf2dJnAQLBYbvj7
dAR8zeizGTgRXWZUXADeyyY6noWqbgyB08q9AQ0eP6VQJpJ1pgxxDhqiiAq/2XztghXWdpwdL4U9
sTTH+Qx0H/7SsNCdns5DGB1nmTcE35HPvNSWlHF8JMQHiaKf0vHc2diAex2OlvU9jupLrcPAwZN2
B7L2bI3OT6GvdINnaumVr0LeciyEbICkuwn7Wuq4iF5cNrG8C3G12eZbqpXbqkNdG58KMyqg00lP
RdDLTCdvCjYzlyO2CsBsYvAPsg/ddauNfCndeAMVrNQ6nYuMr7NuSv8JQYsh3y56Oo8IOAPSGrWc
0VIZySEhKtsJj3OWudBh1lr+U+B87x0S6rziVdhE+4HV/YBF3T6/W5q5+YUDWMDxURnchI6ujh4I
G6Iz0iNolEKkd+JNlO1K2/4J/J8yjQ+AsFN0p7edIl5sTO+8yUAfclTtULF8O+TWmMcXJOctl/iG
RiQjz2ar0qDUheTPMKdOaSB90wCZmEZwgFv8qdrnpdlCZ7moo8eLTEDd49pHMEhRDz+GdQU41XdJ
GDPz+kmZUTHGpK6EyQja1qlesHuA4XcZ/FLdO9wQhnMBYplv6VEaC7rKYF0DG94RxNFCdAXYFJIo
OfcI15dTAyB2lYxhKWMZGkufyEcCpv4y9ylTqFHpW6fL0wqekJ5Bj1uEegj5f7G38PGnTxlylFMT
Ci3IzEirHGgI/DGfLuyTCcHRmgGYvD7ef4a3InoRq8I1QKJYjpV3XOZTJUYhCv/YaLFlHGZKrgM4
rtED4PCm79TReGECCc1ZYecJrq0YP0Tgkx65vSn8y3+VirBN1KOY8Y6eRHk1kwinqmQTvstCw5D9
r3YyA4720k4Id372ku74o0Bfe+++a4EvGlBON2PH4QtP+LbdVnfxA4b7lRXkJglHiXk9hGwZjIKh
ocEKvglGgZEh9/tG+c0GfU7f/y6pZZAGgx1XKEgDmHSJTzwDGHLJTuPO7+HqzspIzY5DVh/2Tosy
2x61Y5rEa3+Qx1TPLjge1BBqxgp808aRWj2bGOg8blD6g1Ez3zLJG1MSnS5588SyZRGwvVXb7LKk
ST5oCeFonJCWXVARcp2Tx/Dj4DxBWFfVqcht4Iwy1o+uH9u5kqBpr9+CzB/KAFJVmL5gDBfgYjz7
0ouL19pOvbpu6v/1yt7E01NNJvRir9l+mGsis7sDNzW5YBejRldVS97OuNhLhnoGWBiK4VKjGiyW
VDVf/fQHTuF59J3434+J4F+YTotOOHg+FE/W8/+tOhUyMBtY7+sfFFKLAp7ZX/9QHcSL1SKElw22
NQ0Fj7PJbMJvHEgw3MocqCUDi1OuWMkvQ6JAvZ/9zniF6Zh9b+FV4h1KMZGSEjpL+XxIAeBHOCoW
PrJxoGeR1KuRZIdMMmVVHilpJMEy6N9J59OIWohFmLHxvv6egCISZIWJSdZo8DKyWupeXqCDstve
0ZChgkwm4QVCa7ReFChgom5Mikyh6H4GizhA6W3SVEmYr9khD8f002sFwO00ATWvC0X+ByVRaASn
0+XQsTi90k9M+zF0Gg2YQa417O9QWtavXWujlzCf71SvJ5+r8xDzAinEPgtLeenWcq3R94TT5Gw7
EvHx5Zp8FqKe+bdrhTs2A3wk71KUZwQQaxq8mlDIrDP0nC8BW1uTqP1mywqfyCFf6iC5e0SvyX7w
6wF/biBgzk/dOLBg/f5Yic6eshqjxv8q7fJFwzF4Ocfkf9Rk4BKymGsOMVbWYIBaDGQ8kbhinW3u
0bvgtGck+OUE2Rw2p39Crm8aTZ3kMvudYvUQhKf7CPSlhkLszUEG1G0JD/3p2hR19V4g9SfaT3VP
EPx8ekGAaAFDW6ROEh5SKrkMsp1rCXa7VEY9sGqK93rDM8/X5VcB0OH597A+2cEIuHerLV4+Bz33
nfzqKn3ymzErAdW7F20CyQmDEfidTwXLr1psV4l3eS3OA9ZVQhIMRMU1yO1wW1+vpqD2B46BtfqZ
TdQDkY7xb48y6aNcOFLRXBhgUMP/F6ypIsniPkpx1qWd69RMpN5/dPgHrOlD37uLkdj5lwXNju1F
bSzlInFo4zqWTkkrpZsYA5OGVjt9pcRcW72DO555Gc4gsAtF6N4hPrvJM5gSca3W+ig8k4T+tzbP
e/Yt40PK6X1Rrlo3PktpLf90CZL/Z1SY6id7FBynuUd4r4NIQUELpHmtI4slvpp8OqCzV0PFDTNH
BBrG8nuzbnnXwqm4gVuqPNM8hZL5uT/NP9bGqSqA2kssOoNqzBwVLRDo6FwvDWyxl3FjZAVHaxjl
3BDPX/ZZB49oOHrXRU4hgRdZb+t5JOD0oITtLgvFT/RHI36oFb8F0yiBTjFN7Kkth7CeHaUVxOOX
7HVlWs3EmlfKwONGWDmNT6ejqH4vNFxrcKhYFVI3XW5b/5VsJ6QNogCyOqGy9nU+zMnB6CCEbSE7
9Vr27RiB74fGG8NXx8oktSOTo3578PNvVj+iDXlwBO/HIPWhtUPVVOTisiFWVeeL11tY1dZng6ju
56CIzzej1/2xJ2WNw5tVYoN2Gbi9KiDJnKffYy1QtjTBWzUheJZoCx/9TQ5WAkhrYqZ0myaG7rf/
bg0wld7vqwSEPdWcesCcCRI7OurhCAndm+vNe6LfhQzBt9T77eZ1Y6rdgT1KVxJBEdewwIG60jDx
RjyWbJuyO0qm9BurS8O2jfRmA8OdJAubccpsD28AIu4dY9dDwTTP9LQfFWoDJXB8Eh92Wmlr/eYz
fByQLy2EQRlSlb/qM3a9Bm9jbBufhGYZW7TRpePWJAdubrLUL8jTwCLgARGiaPoGvj92XgtkZwcy
uUiAjmv1KQrPkPOEqNFQsCeVvdhNCu4+LLNFoh3IAjRIKdlnq3Ys8x0CsmHTYJKLSp8btKbPn2IZ
mwyrgziSSQ3zoB4uIkjxmmsxS1bUSjXaHFMZ5qnSpuj8rFsE0ZqbLOdVSsGe+U/P4BCTGZoxLQ3V
jaxZUtREA7aMMOPWgPn3sU/1W+9W+fRwIlS3txAmmOGc6aCXZ4zvX4kzn81T1xD0EKIJuJAbexVY
CFNHM9eWt90T6bur7aE+oK2p97kugdLAC6G1L1kDE17LAM8U1EsMuj3+qx7/tOVFnmmLYKJmDZNE
vGk1iOwvkRDprPGcGv+kFCsAyEUXgKd5nFA6ajrJzmu0HLwTptDXVYaJLZmR84H1lllzK7XzdmA0
dg/aQnj+qIIYkNd8cMscnIZlRv/tn4NTDh5fKGUCfwbO4izeqZa2FH7fX7P52NusfD9sgZ/e+QCV
IXIKe9mGxn0wEUqU430xnrS6KEnWKlE8sIP99HifAReCcNmKI1YN6qfVtWNinJ6j9LP+FnCtaF9K
0LNCr9ndbzI2Sxu7FEQhuVqbR0gbMFVrcgcWqH6VPQx/pgO61aQEjQ0hBBH43S2mTJoAyNxvofbR
5TeRdhKbTsnl0fOrkkk/rwR0x5MAtIbI/UU3LMJwD9A6Hcds6sIQlIivC6Aaojd3VKEJ5Kwvo8hM
gx1nObGS7D8cbNYeeTm8JkXBmhz8cvqgMnfPVOxAwWEg+slqcCNVB9zV3IYja48UPjk/qzqvGyVn
1++SfWsKDDhrxNuIpGyaretbYiNcAfJhWLd3DHWWGbyBEHZo45XOsHQRgD5h/+agUpAxWflHauqr
LAmHMC+5AluZPk8wxZruAwu/0LuhxXLStSKtALC/U6B9EKqI58rWRSp3CZkzrok5resO5e9WgSH3
u6XQqsornUhjf37g4WaZ6PT/4+MQL3FZqGnU2KA1IATbiC+hteIGFMeJkOFSCKNZ7qUd1RXXFgX2
ivmGc9CWVuwhwlEGCutpzyUlj6XX2Ly41gexJI9DfI2B/lFyJbqzUs+l0FqBWJdvOSpp6HB+O/g7
Zr2nhEfMn1+BUFj+Ri2wepAGqzrbHUZOzbx/UTHK3ZvVfLIO1jzqSU084iQvulE1i3dRl3FcZijz
ZD1tP+5+jauhjWixjz524KEyF9Sh9fNlOe8kRAFOaomC4fllWoi6xPP9rRnqDMf8wpSzOHDdNwlV
6qFdRdPsakSYYW7QwU5bQz6oZEvxpKE6z5FgjPx580fn+NUNSgi/0IFwuG78KrFatSMpNPp9kMve
NHWzaSuRmS/4BeudhPb6kkeDNn5ybySCh+MCZz/YxD8KSA5xGiVZrRT3/gLn1xLiOknj5zs4uEWp
BZHLoEMJvRK8ffQdDkgSno0cCOv6CdMw/fcPYC9buI0mumdcbIC+dXbtIKbhQqe7UDPJH7nmQf42
ItMSuyZXlsV9iOHAscrlklRHEDDoPeDZzuHM3Vp3rHarGo2eg1dOZnqkhGPmD6/+AjrHHBmVj9BR
nDCcNe5sTvT0XF+SvXko2Ptq1FFEJgZE6SSKSGsD+WWDvH7GMmN5uUIUzqCIyxPMxO1f9gArFvt+
5GttJPYthNRPR4H11ZyDiYHCAi7Jhud838fVbC7M3TdJPWWpU0AZMTVrxXYhGq/5spYUuQpG+jAL
zFz6WL8WgiZke1U8xtSF3Kn2kwt6VHehRhy2VYtqIakKrHv2agFYsr9dDAnlNwpYXMqRf1jxowjf
cUIVszUL7vj671Su2/g1ppriCkE+6TWj7jtdYArOBIZqR6mzPt7KQkvP+5SlWKFoRt0T0sN4fEOG
DBt8qJ8I6yHX8iCl26LdCLYwJBoqG79ANQji92lGa0f6aSgCwMfuluyJswt0UqcXpGT+YvXFgZwz
Jw2pTtlABX/YStryKDuTkI2acriG3J63nF88eOsCAhvY54JDQSdXXt136fYxva+Ttu6US4RnVpNy
ZskvRBZBFmCFHFeePn02jumCZbkj8yahS4AdgYdqoZEvrX7UphY+NgFPVfSTe8likaa2UPxn554D
hfP+vLdZ22ZAFOExNemFT9ghzZNA4DMwAiVxytWNVNYYjAQICLGUcwBNT6lq+el+7/G4ALRvsLMb
QNDK8ydF3RZHQjl+2M7sakxt+K2ETGMuSt+wzfvRHhsoJ7Mlht/xKhW5wlVpgOwWKA7gnD3G+CGg
WJCBQz9c2vNTHFST2OWOgpi3W7GOEKlU7vGhh++soXfcbuZ3rZZXvL61PA98tfPqEVFERWYlzp/m
mR1RxB0a9Lfm8FT0QSPX5CHn6v60Ik248+U/M86XnZ/9w82LyHdi6oWY+7zJPo2kAjdyYPJOSIvb
cPMLEMLNCsQnwMGKkflAVhxlEVdwhCAOORs9erWpG/uyHAjU1g79VQLFA1IXvOBEl9+YJ+piWv/Q
NNqgi8t5ae4IQWVfhq8q/AoKAh4s5Vc6gWH27+iSHGFgBsSxcAa+NiG8bfuWiReilkGE3XQusA4N
PGwM84LtKurDZ4vo28p7myl7HSICC0Gw7M1/hfuBJlz18+zcY/yAoB5Xr0kUtQOmDj/A+mZNDXob
xVIS8AcuXdtTJS9gVhIylnqhZ4uOo7xjkEjMhEaiMcnB9owzxiAHvk98ZDcLgTxxBB/wrqwTKK+G
YYoplaKYmVybMw9gaFyeirVz/cGZGu6x8SOsNM3vV45Nr/hFX+XYsU7N8CX6CXPl14DFECOpNmFD
tW+3UfURiq2t51/lGl5h+3ugXLhlwB7k0v01LoM9taLAoXKHqUhKLgXXBKFn6+DYTefVQV4OXjOy
WAQd0MnFLsKgVQ28fxBq9Q7Ss2W/oBC0qzuDhOyXLYVptAYVn9XZQG/bUaXSzqeeWKuaUWy+Ed0/
KP8hBlbiR0w52zdRSr3XtzJsdHqGMAGbaDEgivq4p3RT+Ns3rXSJH8spSP7nd6gVQUiTobIlRQjB
QJaYwuOekVTrhcG35uQdYLxsIfSnt7MZGZp/txpFLpp0ZI1aPDfzhi0b9TEwbMbxaCdEnILUY0FP
BvbZAnC9vLngP4eEkSZkS/usagcsIxRsOl8rA1A8EP2madiDzmRp9rodcSP7xXDUMU1BzKq6J0no
1wcrKN3gdjIwfhhqBkUfE0yAKGg3NPlRrvKEu8E+SREXDH+uuQys6NykngUgD1alRglwXvi27yCA
mLC+g+FIM40jNiEURT18e8AdQTyppTDNdMpPiivGlVuNWjYXe57U0w6Y14Kg/+OQCq9N7xUsAwyW
JyXLeC9M6/W37MjEcZJb546cu7CBB+PVkjepUJdA0FpjfW5OPdJJD242rrTqZ2Nl9E2cn5WO1pOk
q99gs0R0MnEp+OaZumIrb4SPv/HqRhrdnPFeqRLR5Y1zZdfm+cJp9cKhphDZxl+TjafrXhJ3n7DQ
ALxStzzqjcoXiviuXVzt6BVTAZGPz8+NwZkvN94R7T6jr1PFdvbJy86wIzQAxSfDHrXWQayDDYap
RczQRKqp2ci0M6HLd3R10eiOxKqHgImB3qNJ62MDjY5TfMWBoyedxa3fRRaUL44DE4KX4zu+OVGw
Wef/hSOLQaRYU4hZfuWnzAzEykyzNuLOdIvbl0Q9L4J9NF40cKIekNgdth4D9pbCRqH0TnC/STFz
NqwD6BmYX2MgipVhM9CI+R3wsOBJrtWBWoKuXAmPnc4VOhaJ1zYodgRpNmRsdWzEgSUxeKiAoYdp
ITSMQdT9GkB5EPb6knMSA6+hLC4XcAWzQBawKmiVCnqLaWvNkemZWgdNTrshvvLRldHlVJXez+Lj
Xj6Hpb0+GxfpDvlNqF5QPe4dZtNNQxciIJ958cZ9oLFnp9PWPUZDLDJKlJba8nEKU6u4xcMEDjh1
BMZHrCGRl4OxvAKlxquLc2FwJ3ecrSKze1sMozQHIDozRxvACATDcyCSEP9s4JCt/1kA7A0Y8DLC
Xn7LN7ENvrhaOiupMhK3LdMAVOjQwMvPo8EwXaAWv0hjnQdLNLvs7wyvwGlVG6JjAFLVKE0LWWUo
twefTQFJJ5wbnWFulNGUUMJCTF4V2CFvlXMkL6qYNgA8cW7r9VQ7GEL6qbIyjdEZeY1duQ5WMeXK
Mer9V06ayLb/NhFmJb9eS8OsaTDtyFKZ0kD5+xkJZRD4S/Vccb3On/81zF0iVgN++Kv0sXnQG852
btNR5UEu41JiX8UWNfJJxoOE0t71bB29sv4aAejE1vJVBvlKbbZBXz3DG/XCtbypVRJZZhjwrA2i
4Qlq1NEbOuHYQHni5SP/ZLxWLEto6KLJtsiXQsjYrFcVxouAYuLrVqVJV8f0zXWeMUTCW60M8dSx
RXat+lRWz0bhMd2tqg8iXy9kCAkPnmy7i+kKaprIGjzlCNl8Nx7PktbFYbVIPiql1Iv26Zxbkkz8
4vgTTJbBXfDFKTl/9PlMrxYBVqN2aldU+eBlB2fmJ2/KHNVRGzxJ/cPxWkw1OSbq3a7l0mt2JD4O
kJxLiIcwTckyQepNtGd66Yqmrl21mo0HHzvvRVnPPmIPLSM7GjVyg/mZuEkUapO1/2F35ws1d/ix
u6SFvZKlJASDqbRZW669dH0E7cpUQHWSekv2B0Qywb1lcsha0PikzSmiPAqlCbv99rf8b6k0f4Qk
4Nl17vmSGeeAk2uC0VmiI7tZJNP3jvmia+VBBlM4DzC9B6dtsVbZ2v+HBoRS5thUMSRRr1iBlJU7
RhTMZ8SEAnUZysVuW41GmuSFsvbhMSGRFMEMu6ZegeetBqkm4jTfo5GAV5HpEqspBUjCg7cp7aAS
jDXGkuX5PutoKaQQBNx54KooVKYdXnY4C+HtxhEQxZ2LfAMIu/ktx3Qe1fozg0HKKL2cmCvklc5K
+KVmC09IUg46sYR5xARK1tVqtvLRt+Cjd8dSKvaKMIofYJAYxFk6aPgqr8mRJ16beYIhlvqpVXdc
a0NxCk1gQmMaOfbH89RsBIzCnNb4hSxfUpbJPKF240rBgRyMD7G8HdpqFdtpT6uD+CjaCnCUW92T
yNGYJU6SV3Pgp+M3g5IGlBHM/EjzfYya0JrN1jVhq1FATFzQJEAYoW95AOHjH2VrUQUU0/xjcPEt
bftaObRL+fDPXR0i8InQWmcl7yhjkZTLEBc+5i+sAh7EI/yzH2bqkYrGj29vOO41EbfypUIZWJuA
gnp53/d7jJOrsYt2Mj/V3HIxvaVQoUjfj5DJnAQUGnHW6sfI6iXQUACNXatPfU95YZbQhDShVHDh
4/i/bauTQWX6NxO/T8tuJi1KTGa/nLIjgw0kv8KuRNQH9CTaR7+n6FuI7auxh4DW2ItYb/Mupuv/
Rk3q62b+toaAC9Z94PkyOzgBqd60W3zPG+pDf+wdzIQdwGnH6TRVTXPzKrBYM2MmGcAAlhp4cKpi
mrZrLH1JBCMAe35dCENJ3Ev/MUQ+W2I0WLNqmsESaTJF+RPDovBYoU1MCRtHGmHo/kDki+YosTfR
3MEc+ahCcLvdO6sSccVPVOeA4aYhWkjscKI/ecrZLlbR+6W7/6K+zgNh8bMIr38A9Nfsg1I5RetP
+0ZWrL78lfvRLWtDAzGPH3aDDlseReR5ks096bKram2cIU6KsPQ/xXPYFvmtNRutCorZ+Y7PsUj6
+6fn6bu/BAJoc/J3TgF4jL7V6GzxYvHESMaVOOJ0b5ktV9gTjCUBXNUwKyI48WrRSIyXJ/m6jTwJ
BUgLMNRRH5kOpZCC86DoDE1aG4FU+c40KUoVU3J5KNxRZZ+5mnvk22zKxWgYk9GFL8vI+2l/2uKM
qUwc3N52FKGnYXMuZnDYoEK6Z75M+WNcVLqh9Rk679+iLgCZzyEfXm6EkJZQkgIDZhjpTqMDiyKg
PF9vX8wJUVSKdrg3Bwc/KD0upS2wkDPljGllyumfa3VrzWp5XQ9Yk0p2iY6C3agkbMf16tHWiWeI
AN3glZt93xNy+WkS7r9AZG9e6+O19B2iouulz5R7Mxdx7+KlTOc801ioM85k9XtaDxh63UeJviha
Nm8aYTm/g028OSD98EkG5O61P7Ceqmych/+bUqxb3piQMWlSbGxKk1d0kJ/8xKCKqEehS0bp/QK3
6XGmZkpf4HzQxz1+aV1Vl8rAP5ANjvvG883Le2+zk06dqgZJa02KKcr142wbgTvUd6soUTy8jZxb
gTiWlQeS9Qz8Ug2uwTs1ryG5XZUpPAuGM5Rl8jVSF3KHvqrEYyO2BywcZO8/aXe9WqGs6zwWTdPI
S9W1EYhOc86peZkqIszu/DnDAVTQRwMGlUyM0ZaZo72G1pg1ezP8DvkQ3eB5wj/ENm2smWs4/MNL
Wj8df7eA8L/hh/6Io0zd0RNQEQyTbtTsGxH6qjhpRHF4ZTT7uYUyzopKSJAzp6W/UzsIYw0xQmEi
a78OvCS9LPHh3oxVepuNwX2W4nNDzgPKyCF69oceVp3GZG7lKxMJ4J0ejLtrYprvI/bT9Jd7F4hV
MTYCU0EfjQfCh7oiMKi6OBC1AjqVjw6rj/jVg3M1ACN+juceNOT7c5ls8vOZQ8b2B/XAtX7W1N50
ktZ/n4q0galToTCbAWA2uyfhiKL1Mdi040Ah0nUzY48glMcGgsfgjQOFTpWjcrokCyYJuGhh1Gx/
2KmQgVHutv9NhJn2Pj+ErRCL955hn3MUkq3q2nclOobRMJla+GE80evaczOeRyUvsmkxNMC6+0zw
NrufBLolALF2RFTIfNT/JlXR3zhlfQkuodoleQscndHmGiEHMH0jCNrT1s9iq23VdieW47P4rmj6
yioBrw+mOYw7D32GQCYhL/Cw2QGrklssCVFjNt1pF6P1yLc72OryZi75kf46hrzebYdc52Wyg/Ne
8+blaDB/hb+mFnEKTcvH6S7kL3/AjFR7m8SMSLbZ4HACO0WM9oWwIijnFbEXWr45Nr0Q/h0vdr6/
xVbTnjxcI8mM7RNGE2DME7RuTLYcufTKQ8g8LZdRE9t0bBIYbHDLe4ufdQCEq6J/z9359ghUS7BM
PNdK/J+oWnpXCTedOQSNL0Ae/QVziLNRVazD1NrrG4llNjhgMJauGftjhko0Nrn1+Kg4XsXXDNpx
zo0wtZyc/7qFEc6UZyhv0kdHASiljAoQKG0qp22MLPTiGK1nmQJUtIyvlzLaV/Yw67K3TnyXznmM
ETwetGsnNHDjJ5GJi3+58cC+kYCisEgX1JXPW5x5hSs+NhvHA5k7pJC/83QUxfogPfotdhKgC0ug
26WMSbFUyKw9haspq+AJAlGgdHZtsYIj93LwJAgFmIQmBgEKC51d5pWMoyqln5tL1zsGGKWYJeAa
B0F/1LD583pqxzrHNcYzXCsJj5w5F+GoZAjMwy580tvk8G8IMocsQwfVoL5pKYU+SqDjsP4i0zRf
4wtTHAueNkzJByZDdtnyuXs8ahczpuvClRCETOUcH29XgBM/ukJnDFAfBoD2X2LUg5prHlftxT6F
VjZzjhKtomAqbGvEupgPQEJiqvVgUjcw/CJYZqgflEPcAYGS3edVeXvia7V/sWPcPOjDwUOAsOdF
Jo+dGC9PkRYffhqURG+ipLhfycPFLhyqUBIJnZna7RggvQln+MRWPamj/AOKvoachai8/MBxgRxW
kVlpwOEOdPmpTVeYfdaa1iBgpWWgedwGB8wceLaL6ChLkGZnOqHMLuFVLUDbg7FqbJGC/wD0olKt
9pkPcGAOxQ2b8PsQrFiHuz+QQehddguhXHwmq3D8pVVFxfg8lDnc5LElObLUUsKp0rB3SzTZ9vb/
sp0GoCprBliq5qKtR7kU6DID/oGuJEBFOloSH1jGuLMfish7pI7ZozVStv4r7qBmUhHn8M9BUCNN
bvLH+dbcXSzPxZ+4NKZSkwcsfKOVpOjYrCxbrFwbHbfmzCAKUToyoLB1TrZILI6uiLQttKaclSxA
3R1aX7ai+HW+I+0t0lAujOPeBn6wfOsvSY/0R4NsDdF68WhNrQBBt83WRQdGnnldVsIWDtWbej9+
q5jlATjo18/JTj+lVQhV9b8chYPt9S9ffY8Qn/7NVhzFL0uPX6fW3vEm/wSNEkuFGbm9qBuHIhi9
H63f2D7GKWe6O+CbquRa+hEe51/0l2d+p/DvRtyv5CbUeffbeiuKWAFgV67SQoNs0f9+d2GGw0C+
J5puqamJp5ogu8lqljW23Un95ErlGA4v3yDyhwL6c2M4j00swA444uOAtknIuYTFpJy0cFaS4qk8
ChUHkJaouHFHBa76Az+/NdVCPNXVijnvZKG1/RCLXSTSqe6eUNwXZmle3sPCgOItpY5NpD4geOMB
jKOF6T1pRELfo05f7ujmZZh017qVna32Ucp14Rt+iUD4/9GuyIpXiC6BF7f6ohBJx/7XD9Pi8we8
cHaXTw6dPA++9ZlbXo6kazrzfV8plg1fm6qhWLUMDJ/+PEK5Px0J77SKXNXuAPdTQel0lFDWvkLz
t/z7YolHXiyo8cN3SIc8di12+QdHwe3YwCNo52GNkisLD778F3SIDvuWM7rRTuSCPIKcZIsgZ6Bv
gCRCWNukYMP5m6oFfq97a/CNcTGwmCr2ybfvgxqC2mYkqlcCBfFpM+3b+kH489sgLQgglq0FFHrh
aKsnLoEYi9fhEoH+LqeAE8QQ70FR4GH9gzyIhbUxO0fR2P1U4oRxYY5Z+baCH9xSOtsg6v/60ZV0
YgaMh7JlaxYo3AT0W4lW8sAKBJQH75qhT6NrT1bUhlm+ncV42Uz6uJ5mg+pae7C092nxXMO8IWWx
CkhmySQTBYrsdNQb1qYRKfmJ5stR4Do2FGQwO5O16w1plFF7rrZ9WeeK3UTFanxbfazmVrjV9YC3
pQJKMkcFzX9ILB1gkAFAXSJjwfRPWTBF5wHcCVdtmXpwasDobkW1N8dma4Q5jBhg5Ej3VQSCCPsc
mwdIWuUrkWPZLhejtSuOmRZQFPRGfaKV6BwOOF3zv6o76CQwo1RCFmeSREH/B972hJhMgstNEhKd
yOSCcTi0c+sBscMoasfO/uIQYA9arrWq2gEzV5Gx3dBdx1eZINYOF1oeD57hm4Xawoqv4Ew6td3t
tSNB6FmIPA59SOvKukXb4VPG8VMx2tb16lKqvDXG0HQvvuiOzU7gXfUxkstB1XT/poFI5yvNgPPq
tDaJNFL8BTdL1REOxeQNwSQnW54YCh9JQJQ6dk9IwzlgJdRV5K4j4bvdnshVerb4CZ6HrQhMZW05
jMlOCCfAEQVp8FaqIbViddZxJy2oRokWW5gP1StWAkyazDYkSIwT+mpIES08BPYSzQKiTtsxjhVo
fgWk5mjqV+LPrV+KEF0H3dVVbCa2I9KlFcNQn10423Gcnd3ntXNPIIVUXLCebQDB4LailFVnkKlX
SZomDHKpm1ZENYAdLE+kb2F4FJ/UZFzI/ktB8Yq2+QcPi5054098fjTFxW7IrAR4i4M6A4b9RAyB
dwaNHxxP8VynC4s08qzpBJCtgixYZQpDbFZxZwbNEiycYyQ6p+wqGbLgSNima1GTjf9Y0fH6n9CJ
IUYzP1VB7H1WQzn4vx9o95DYveMikMUMNKD4yazf2uMApvoAf1VgdMl3EGw0QV6dj8dYmwCv2H/J
5rlkuBZwAQd/IUr9pDWxUqL7JpAajij9ADVS5qBppIPTjO/UENFE7YGDTMzsOwJnRObc6Dwi9YMr
buGxzXBF9mwec2QD8Xr0G1Cw/r003C6Z6NkDV8HAUqtHPo9HUwbKomY65aEtDX4yvwoMXwxe14hc
5mMaf2AyAG08U5UHUrl+l6wDYc1xTlglrIREMyAzTdbVmYRPeJV8PhPSUAdBPrV2QKVbTdm/IFBu
iLzP9wQcXiw/nObqxO3JQpAiSj+iqj+QA7p/av3EvGWquU9jrJTIU0+nJQosPOINmPImZqujnUpJ
/f/fW2uiLIn2qERtJPlpxhwyMoqhLBCu1UKYoopF3MbTxshX6UwEQ0+UZRPT5ZctU9uqF6uDR32T
ZCnCyGWRKMI72r1VjEUU40WWsv36bzw6HpEMoXowvIy/qZrt9xf/Y5NM8Q/WqHUuPW1WNnZklOxR
NgtCnMUXVKJRJs8CaQKI/cXkusz/39cl8LoXK+ZISFpxZu3SgVZLy+h6CdXTyvYvdgs+liQdAe1N
p7T7l/5/yndMdRNkkD3nb1swpN+YpkjGGFftQfHx46vK5qEpV5p95LCOrL3Bx5axkyfeujB7jlEW
GVEdWT7DDHXUbsXUDATRMqF6gQz+NCG5n3KL5RAzABkWZKqQYk8lBLDS4ihGUvsAmSG2xB01/0/G
wendfYA1HL4xt1tOTZUcH5jgb2VKB7ErZEkaklGYQuH8wL3npAXT2i23Pj7qd3IjjlZC1aHFXOD2
Nc80Sry8O9YnOJQpqjVIwHmXrDPGtSyKRjmOoL43vMmtt0OgUNUIVCNfjkZBra41WjeyBTTSGHTY
gRJAOeCyGNo/IFKmatocGFhxfhoi8KWMNXmal2/OQqOtEUUYauky/+hBFHerED/kyXdD4DGgtHXJ
CoI7iJXNrFyEO1mrI+4EFM2iAuuKMIPMMyVDrcOYsDlNCE4SwHY4an/NDRGgvawivw40ODQK6U08
uN3G/1JpBgyDp3mek1EfIqX6HjO6ii+T1EUyyo5TQz8agA7A19czFjrcx+RXa4+I2JQl4L81YNbs
97eKxDHEiazO/slKyHJC9F1i8BsY4L6G+x9C01bxcVcx+pTciWtxP3gQSK9898tqBBUzMeVYzeOd
Dq7WGcp8bskEXlAy/lr2fpjPRpcA+BzlGT6BoWKAE/0MM59PBYaXf+8tMGTDNp0RPVGdbY7p/jP/
5DFo8C6NY/dSvx36/kaWMCeApzvZB51bfveu1yMuBmwH09XurKjCY5cjjUOCAUvsnQp53yVViDBm
kTUknzc7r5bTgr9GFPHRQi+CFIxkoWj+pCzJwAypZ49B3IXAMDOyhH0oH8qltWZO/CmQKJL2NjEa
UJmY72gzhhlslmFQPm4hSly3nI4zaf0jg2hPyXiU5GBDYKWbqfNBBOV1zrsksDnUDz1wUZeHLOnG
u85IvxWMRtKM7dvlRhXw2wINT5iEFB+V97G/4+Rbl6bp1nS3Y3gkYWhzszmiEr3Hk/Wd3ol3559j
5OEc7NOdcPHNTXy4XbQ6C3SfiE/0Dcuk8rvtG6P/TJQyMFFU2fNBC5TINF9YW8C7d8we2ayRXDnf
L5Uxrj100qpvspXcpVU+eXGa9Hz9ClF+lTJlwpWzL0dgv1ZcYCDryW7DNG2lvRD2setoxQL7+HlN
NMZo6+4PaAVuj3H+oSSeA+VA4fjm3FthLmXUIe/AhE8I5MSQ7NrUrW6pJNJRU5KOK7vaTPJHv78e
uvHIUBt5TwE5f/ii8NCZ/s1odd6X8bYBS+v1Eru1/nxBN1uN8jUmpiAitKLMDUvEwr3k72Mo5hPa
70q6rOpBesls+usIrSdNEQldX5YhmLEgRnDiV8RbRyOZxzOjTrX8KDz6kcHTuPVaXj1LZ+puaLYH
tqxCI3H7qvNh4GQ8WM5Cx39hhdotH12OYK9JVCz9zYLk+f2LWRcBfGZgT27L0C3K/lYj3JNLd+YZ
MOOwkUr3NL+Tonc8QYeQsPg+uepyY5lAJz2ayd8ZR3xQQDK2kOQNu+23YX7aevALLfiwDb1ZSw73
ub6+ClXRuhyfS4RSm7J8heF3NTzaKvwIjhKL2RAzfG0uwia5+YeqxOoE4N+jqpbAbaQxBzaNEpBc
nq6Y2pusnx+JNrImCidMDejSFOLaaqT7EAny1liSshiLvjptwR8JPpixx7wS8pAR5fnuEzrgPFW5
ixjYNV3wmfEYXs16QZ4ZtAorexyBU/r6aGU6L1vOKxhkO+ylX5Sh/Jg8DZ9UuLSvBLHPzONUf6W5
e0Y7ey/ndj8/DS8FjRFyk/JYcT/P8sP0PrIj/AuuqrEhnPBErYEfi/RdWudi1UeZLxpzroRs/lI8
KC8s/nT+Zb7W8jizUg7KYvM69KnMVGjiUBRAxELUBgRvnYDAeMl11gppxCyIe51JrRAWwGBNO1L7
mEhSzYkqtQ00yhuUhG2p9McVEaF+O6MQbBfFyelvuQqqAfRNDCHa8dyhdqs072Wrq1N8Gv0bfLmd
KwGHLbhTdqxn3dZb1G949yYLJJNF4Lp5NqmJA+N4+84dtAShhu073jeQqBxMhafA+UxYaJ9FT7/N
9+BGNxHCOjKAppESih5DlwgBMCpgOTyXSkZ2NCx/WSbV0FhJvxQ1JpJyvisS63gdB73Bjltpib2W
vcfjh4X/+8Tcch6tzuA+8lzm0XYgrVwkdmj1keU6l8ElzAsv9QiIif2IssQoCY0Ur8uYAE8jwUFb
+sPc5WmD3YlOR/GH3doRM9q89cxAIqg2Rq4MqzTwKPRr+v++IBmKPpsaCmLGALOULLBR5Fkg2qM7
XdVOKiAyvw+0NF4JA0eiYcUKH5COOHAYrF7+LNQletxPfejK3HLFgO8hJd5NoA5eN9MFku/sLgj8
bjXQKOrEN8mFRxtJQvpFQPDBNdxeL80F7GITGHvYtUylQq5WLP14TcEU9JM77SdWS/LyD+Hl09Hd
d351FK08SMxxVuRk5tfAnuUOLoRN4iF4dCLx+seC9Z/IIbj+bRNBsnMXmqNeetcYFPJj7iyEZBcH
xrnBiJh0axnRniKEsUlDjGfbZoOUnhwRsuSbAevlRCttaXU82oS0EE/dU6mUIBrTwrv1350X/itq
8l8VtEeijX/i8jyNmB83VX2PWoHkvmahyEHOlD2OyvS/jSDQO+RL6jlR2O+Nc6uJK5RXrQIdkqmr
OnyKYx0F3VRFUcyHWBhuWCt0PmElUeXsd9FHWY/Ajqx1XRxJqdXPvgA92f8g0TIg5zV3vLUnjMPx
B0N/GcCMf/5xx9lqOcoyxpTvud3cw/gyH7xDaIXlr2I03bE7tzFCatsXrMYKak8Ry+6xH77IgBEi
QmnzH4OS2RcdYzl2vCAcVZFEYZ9gWNrWx+o7U58r0r5X191k2WzAUxaH0CICmRZ2hQ5cAdAP9RB1
E0lz3Z2ZRe6Z93GjgBKXtGwG6xpeMYro6AvEjpcWK1GE+WwPEbTtdei4vol4qZeZ21n7wXm6bnKQ
0Fvi4DX+okKfVkhroGPW79uBoizD2E6zpEClEsPRpS8dRkEmmGwXn5OC/ghjz619dONojW1ER6KG
K13fiyx+HLWkbS34NMn4ma+r8bE/6DOPBSczx1gcU80tvqvJmgL2GzM5PTqo9Wk4zs7KRkpI4CTs
4jQZ8pfikJ1z8ZbTkCtdWEq/c4MoKTyjTp5yY2mzJWvEu1NCpksUKHucsOqNF+hlD+8Q5TBt+umE
RP4fudtKafBBZcGPNr3Cpvv54q9y9Z4mXVYhfLqopzsgR0G/ZnHHnGWaTrnPvUSTVyTUU2LBsxbn
L+k4Nl0vhpWgSTKutTHojxYZRSKp9XnXO1VZvFdMGo9LZD7uXfABFBJ0IN7ksNq+9I/5fgvI1WN3
YJq+uXeKzuBTEOjyBoa638ius6E6Ut1cCcZFzC3UvNovrdHB6s3mcMUsYC+UkLa8IGEYOhtWIz6q
T291jnrIcaFjVtytYLiNMh10Pf5i/9j6s+jTX4YOZoBCaMPCW+hyayXdCO9sl92HWvI0emCd0I2E
mwFxhOGGuxbB0f4q5O7NFvJoRWp36ulP+7TWnKwHuN0mj4G7ez5XK8CYhfWGediUXdtal60IddUD
jnWuc8VTNvi8on7wwPIaRJk5YESuIZiIslzcQ1oa0icjNsxNG2cRlTcbdNugcDSiZIbeIMQNwQ0p
DWq4kVXQuBsu9EBl52LJqhcd9VD/Sb2qRRdjp/1s3LZxXco/JdswTCPGqpEcndQ1twpPpRBPD/Rd
/bqPV//ckAb+zSzcqFTo/lPgz2SKDuIsSB88rBbjeCPN2Wsrc5BxihvV5DVncdRXjYSmYk+awvMS
xVk4HpETN/46GWX+RRlgoG0RzhzktJKh7VQXieJ7JToypewkLlX6rHNjpXeZChACrU79AsEg9sFu
FDxyF50kMP4oGFLW+b5x6+y50KjtL4kBWjdlB4LqX7NKl6+lpDn2rui2Vqitz6xuXBkp7Z+l7wgE
h4MH2o/g7uCqhN29u11OBqd2c5dSiBkDBytv+l5ddN8eKzGE0nxb4/3Y8VfQvsAPkaExrHUFi0B4
pOEaUvt0qZxTtXTRZm65AzXBJQZxN8N+M/+n4BoV80aPsIWWieqJRAUCFlvm1PNaoVJ7zedGgDtD
7cUHEtCuxSBzlFUJed36JUbG/XKGWuVlZuQrRvHVk2Y8y3YOVHk4n03HwFhIZNOaULB0gXDJPcfE
EHe03Dsik2mEHrESEllXxznLyHJIHULMdlFbDZljYen1LuzkFxxloXDgESb4+gIX4z56wZJjGgBe
uJN9m+xNoE0Sg65we4rwSTr78u0VqMYZNnpK5Jm3RsZ9O9SbVces/UWnjZwQR+i5kVts3hOvqIYB
IiRxI/X/qiRl2HGUm5sRl8N8FqFrGk19A+n47rmZ1IS5anJqf4OMo9SXZlKkxTt/mv8FR6QFBDG/
3tAfX7NP1WAkiaMXEpeTn+er4rUOgSl3xA+956aL8lFIMNMBl77rJtcBt+Sd/cfms4VudRnozhe8
7ewzNBJdQggWurPsNTKyS8JjJ5CJ4WAuDkBRbENP3V8JOsx43f/XFlTRAnPWiAkhO5c/8NJOz6+m
FchNy6k+hRuxJbTfdky7yzvs6q0w2ds8FdqMN1K+0ccDTIAsaLJ5nAxyp9JN2ELZaojaQaHabSQm
r+JWqRxX+Tlu4PRJtt6eTh2XZZtOn7pupQSDDBw0elpJVR/sEX5Tu1leedC6grpV1GYew+TO0kv2
Tw1h2uOkpep1p6lfQ0pmSVP94P704CANTux5VbZkhmBBoW3KJddAsiYD9xoR8dq4x4glSsPuwKQq
emHjztcIh6262Nm9mtA3VNiF5PTP1TTbwgXpfIiEvhP7zTz4rGN+ELhA7VCHxBDXUk7ipVXc7vT+
e/FCw1YolhQvVmBFRdBVFFajiXS3AXdUfRKF4pSWdhxtkcXFTkhGVZQIQQ96+WGQ0d0Wxwg/UizP
W1BLMKVZG89w9c38qittJCAvJNc7jyPKwSNgG0Ba+RTzN3kegtTTk3X2VXIgghQqmVy8voNM7DcL
SvNCzKRI1W0QXzHRqvmKiljwJ+Qy0Td5kj9UiCqA6W3F9ddyM6pAXt0XdYe8BmeyivunLfYiVkbQ
2WeYWzuE1jYGdpYX0bhXcp6eneYlE+ToWb9HjMzeJNsgpcfa0MBN/TQjwK9cIaMFFfwZ8Ebqa0rl
dYwcTzrYvwwQRzlXOT7EM1MAKy1uZ9pS3RmlTTbQR+ztW78u0IR/IkFJj4EH59X6yKJ+FdzrhymC
dwySVMax39ivO831MsFYwZhHlqRfRCDisnbY6tYaiG2R8yh3FjDLaqlVnDGeC5KCeuvUl3WGpWFt
FTNwQvGYAHA9uVpDZ6t7UicOIRsenJfP3Abby8nwkHReOTSkazLzTnAO3dLHDbnIqqMbob2fatfS
2fiCOpAZe1vhnr0HotOailsJwJK7CjjNl3gsiHR8n37IL5K9DowNnkPqGJ2dgpsHiiYMcYcfrBH9
98phuvWXvMjJhiLNNty9NOQVeyCZ5WiRKjUHmdTWz6zESFQnkY4fBdB76W9iS6Ej/lVNRSzYYWwk
BbhAlrCDoH40ao25Fo6jWDdolUR/p6A0WSLTx6r8vwGPNpAxP8tE+EC4HOwt5TukZrvAy4UhZGwc
NxipHJziW45di6/oKlsQhECS/l7Vb+80WrygpeoPiWi5CldDcA83M37g6dUKYnzqfHDraa04kY49
Dy7T/4wmOJfFw/1zbTPbRp3pxMWE0WYWS94sI2Ol9P1b98OoXULRj/yLVcD8Y7BihEPzBkfN1bdV
0ILUyiWLLENGukDZDSEDgyvDNEewjD7ms0mhC7dLtJb2cyTiy7wolcUJyKnNsQSVSG3rNopaR4z3
ntoBRIah0cQ2LC6oboB1C6nlkmQoPzO+ECg5mESObqzBZZXY4nAt77VUf4EWRX3mkdMT+XgiYbjU
jzD57NpK/dBMk3zzaZjK/jecE1s4Q1MddyQwNq7IjTck91Soc+C7NFMCTkJ6te8FMUwJd4W38BMB
btzXLtjG8WkImyLelmLXbA0jqQc2VsxiD49KGZyRoMXVlQEN6j0gvgQcBqRcVoEqWtozMgsMprQL
rYzH8eVcPM8fj8wLwd0nhVETrMUkIDYHlLWuvCREor+c93DoFJmsUi0OM02sZ4U/iqwcz5xeAcG4
B8evPshNkld+dJcgj1BypUVzmXGO3mNdSLuJIzQRM+w9qFI+ayAZmvU7qzLcFNgffc0Ct8JF59/h
rAMc5qTLaLkWGgu4tahMvSOO5eLRsyYzEAnhUWQeTMoRjhDTFxrZ8WRzBafR2BjWFEPXnekkapol
b1nvmzfzbxGNkOJrng8/YFNtaSDavLsbCdx2THRqwdBemZ91gybhcMmSTtzpi0Ryl77unhis7bSV
FlbbUYbzyOLqzS047UkNXRzCtjDCueNsNfxbgH9NXbfbLTD9Ajd2F4oethwlw/HC/sgsG+VaKgxQ
V47Gu2fkdPUGTYysj8GI4xgnHPlFKe64R1gxZIL7gYM9ZJ7ep9w66pQzb04kbtYa3kBXlSS683d8
O6MnJnkm55DGCWe+13qrekqH96sm7VWrKDqiCTHVhqsf6kkHRJr9XydeLmaloI4yQcDUZiPDBM46
n5d/Dy1PTuY5HgbdNH0vBP7dMvv5MOKJXwxYz6IVXFopJfWqCKbYkXFQz7K7kLUzhPsI3KB2yXO2
JctJd/FC0aJ3yN81J8Wndbx9eJ67T1rbK5s1eouCOg8lTI3mYVk6aX1YbBbBCq4KEnJqpie2rY1z
0P5utomtn90aVFSenMWhyRiKMHb8kzYhFViuYkygCk4KEQbNde4JhhHEAWqsXw/OukxiEokFBeHI
0yKx3qNh23Bt3TRA55a5Ktzy1x6xZjRqTTEYOaT/xfF7WGcPB9gtqbnsXUrJWovBjmmkvuSrSf0n
qTcsDDCgVrvZuBAJMBu2GSqQRekSnChVWH3zGwMZuviWlTgigLM0fuLaWdaC5TDoaOXsm2gg7TR7
XGJUWayqOUFn2quhmpRS594cu6eIawRYUgOwqya0xWViQsGQzbGzy+KE+wzrxMU7g38FB5Wc9cW8
EWohWD1RbiU96cgW6znDeRP/ESktM8B9wfHodUCkz2um7JTuTuF4/lYfl4pAcdN3xXH0jLRaNO6X
VmKxVNKrpBIzwwDCN1eFoGVrH6ypNQkYSB/yXThIWo1iXexkozdnwszZYop7ni2TFxJrhUvw4UlM
aiNeSKtkIFrMN5ZlMcxK3yHFTmv9p2YS6SNvGvcD3kgqeZ8U/YIFuP0FM1sXo4Cnf7/JMvC/jvy1
R2UvMX/gMzq/yRv+dAhJLcOt9ZXDnijuw+UAJ7JDbkMK7WC3Uyfea5Q0aAkuaZK37yhHGYVxh08l
4ZYeSPbBdJ+T41C+f1DJ5GhLwN5ubyK1b6VSzvFnEATwXVXjoxrYFUJpdqj/AhjaEa7T/OqLiZ4z
0M2gIyKZVGzaKuntBlQ0dWB6T5u9B4OlAHNJJjU6v7jFL1hUOXqw4a/VhOeGooY9RdWkwe4zxSyL
z9DF4C9ZlHDLmVWFfuoerOGIxS6obxhIB/V3BcZ19xkyGWyt1g9ovY+FdugIhL75WDyT2pt5SbkN
FcfACISYqFj06VKbI5sqFyAvqPSGpXR5XWHm9Bbzy5M+cKGL3JcX6oqquXm13N5ap56joYZflnZS
/xXgY8kknoGK5L54gucaw70oFyv+6RNTmJkElh3YTQREF/hUkc9ViZ1nhFnlXCOJfFjT3bRwIvCt
dBPNL6PFYIHAZVw4aU5jBURlFa80Ii7WGqhgxkhDf0U2SlThyeN+fOhI/BRF4J6cEs/YeF7fg0Tx
C7DnAn3uTo65SrC8nZaKShgKa57VVMIX4TZ61iZ2cqpBNw2a/D345vUTM65QfYX3l7AS4dh24v7A
q2m2rAdMF/yT1n4giQ0bl3/DMcG0G+sBEkSTY4H51ZK1GKBbx1g3OSlk4TlBQjJC4ep0jzEtIhm9
WroyXV1OpPysLtbGHzV/CXgemiQDzz35gxDxOeeXGrdBUuWfsbYtV5Mc7p0OW9RyOlL1+l7XfoGl
yetv0L56ri9cvaqRHyYye9WzGr3MLdoUKBVs7qSzrTqm8Gvm/ZIihWP5P2QSKs1fOVp0OPrkOxDM
fPEbbi5nmfi5AddnpKWn0OAHx+te+50wQ7Qgd5ul+f/bvG9OHVKU/HTITmMakzQaapn0PNwKYtKc
2FhvOaH4X+TSDSZP+LMYe2LHTkLwsa2KFuXH1izvebD4uGmyrz8Ou/ASNCdSL71FGwQBnhkk4iQW
mXUNA0qBD7LRnwu+MQ5lYyTRueqrcn/qsfJN3FkAIFU1OmKEoXDNJCPX9Xsb85Myg86zt4FYdfBx
IsJYeW9vJgiAofuuq88UkfiKzM7MQZiZb9JxqtBHTkWprpgneglb4u6hSeU5LduVD1lr5o63PNnc
CKyQoZefvsqxEoFcX3/vBiHLUzku9d0xk2Iq183VUKpCQbsRIX4lkjTF7155Lpo8waci2qRQTBNw
ncB6lowm/jR8jXu/gI+H/kUQ88+WIqQBZ/dp+cf7ipbjsKE6wXYeEhmTyfmQ2jANcV5Ixat2FH/8
ShvBxYxRvkHO69k6LdhS5yesdK9clBlirb814eIw4klO3xPnkHj4yAjf2e4H2O+zbuhfmHAzi+x5
d11plLiSorSlFB3nUcL5ITMAcZG3wKIGxNkeL5Vl+FtXMX+PqkgvYuBdxh6yzV1EGQxaTJxG818V
AOQ7rV4mb8PYJVA4ZLhvZVQdX5OFbTfyowD238F5gLGjxOiL8Gx/NKW2gowywYq69Vfu3qFAt/86
0NCE8HRY63ze8laAkBcRvCZ2zjMvHhYkkd0eJafSo3y60vh7lzLLjvCxTxiFs8dm//8yoowuS+D5
3BLbTpwkFEgxClC22FzKzrZzWAYJ4jGG7Z5hD6IbVKp7+d7CzBPWJhD/37uyvP39NXg8Gh2WekMa
+NGV0yKB5mPG5dMyXt1SmQlCWYGvj7M94mtejqjl17Dpcvz7bASSO+U5rHcIEN7wrfVpLMVm4sA0
RVE/CH8mojtByNJD7Uv2YfNqujx4WYIkR3UyxZ5WY8F0svnTxa+Zz2oj1TkhzFcdNfUiO23daXNC
IBYCQ7V8cIIE8YIHoZ79P6DrWSqA5C6ygorXHM6uDvYIAXK+K05Z6c9QjOKGOFm4bBJI7gTV35GT
759aqKJo0cEj/f1zaPfQhxPmy5O7vCfKONTYjNis+Hbk0F03teLQiJ0FBh/osqluntBYtkepLDq2
JJ5W058YSzmgN2Ym4pp3ZDeFWCaEf9yz8boBF3rFSlvUo7KUlh5uCsFKEdEJdE/xhj5BBOiAfem3
Lzu5U0piEaCABDSHJmlI7MbyNdv7/S6zkpKs8a9Rkji7QuGsZMD3lp3rAg6UxjrgecZUBu8VTkYN
ldheCWjHW53ilhB9+T7HsfPG/9mLS3oqXsnAY9n9fTST8lKOSmeRU60I9eXSrbfKy6YS7vBKDoMO
pZKPqnPNPwl0N9N52vsapwbP/PnBWReYWE5P4rzLl+LajVOO2MlxqKKDvUeeXIIuvFbtFCtPCaHS
JDiXJC0PlmJXPRQfncCPxCPwYZofqWb4yVsVosI4VN0AbMZJKcHdeALk6d6URzJD2EpKjVIUsRmS
37u9dQxuoiUZhH8ao/uFlVhLklQ8ZYZJJMfFbPwiUYOtMMKVXK0vbXtxRGP07+BNWVxUNqKXBlGJ
3tsymnF6UuBflhOmf5gA13+W7qErR5DvkSS91CpSB9qq4qf81XVGt0QQDx5sl/8vXKtvnFampCyE
hxI8yBx6XSsIkcj5Ibgd9a09a/jx2coslnunBpgUbhOYOZaC20txy8ucR/5uDn8GH641HzG34rfG
OBuk03IA7ZC9tlVD+Vt2S5HCqx+k8iGkpWrv/dW/Io6YMQ1csL/Lg6AqWh2jZjDr5AUN4m20I1AM
8hxAFUoVI6cSI5cKfGpm7/bcUUuyhh9mLbdPLMjK6nuo0otmh7yeU7CVrxtWjXpL3cBnNdP4vK0u
Wn4F+e4tius8W/16/T/3/x790TKlyzGYea31JUa7+B7zLZRu5f/dbGdIIlzLJtsTEUuazmXQMAst
El9HOZLm1MzG9e3jqVu06CijvcDwRTsbiBuLV2S0YA1xaj1rKmfOKj/RxX/EdWZ+PTbfe5v1tBBo
3UJAQcnAKNlL3oQiQ2+iQZe/6w80CwUqNZa/OcJH/2nbqT/4C3hn0vYVW6tQS1XFIy3AMTAJC4CL
zK+dw8Xmb/ySVMq4XnfYl5ky+7Xzfs0GsCW2Po3b2Uo89T1bFL4SX6DtiKbmaoPkcDkNz8N9R9C0
6wtj6J28BEiOg5gD/gW+GNc7j+s8GFF4yIk6URpy7E8hb8rWFrjYoC5qKMUJQG9UFVEEY7Lt7dXW
1nhNXdPes8WrUL8GW9scAlYneAgG80xCsjkjEzUBbFAHsk/T961HlB8NjU8Rx79bqDvIJmZ2/V2t
YMPqhht8tkYimk/01x9S9znMOWwIIKcaplCblPirc9D46kZrFgqfbxohg7EDgsMwt2meHrZTkuM7
cYbDzQSrumd5bAR8ID5t/nvNlEDZEbf8ZP+Dr/BQJecN0RJaZBsjbz2DwSkiZzvkRF0A+7a7zSPE
k+5A5HBNLtkLA29afDZqAnQ7ZjFdwPxSFd84CkvZgnRwtN2VSdKT3OjeqeBnKFI4NZ8q78a72rNL
m4GC14PzySdr2ypbjZW2sDSkU+84IM4kG7DR3uCwZn6Et4UBK8LDMEl9lgb8SpoCLqwctONFE3Wn
0RROrMb/9SLuu4QEVN9ABuokM8hd/6E5Dq40+JlLNeI7N2aW1BHfSvBnV625/xTwT7+0FGl7pd8P
l4S9CZ4xJuxztlME2oDuTLgwslULVRUJyEdk/QYNayU4Thn7PEoeDOMKU/ZuE5qO1Nll919qxaQM
oGgCkMO2vmxzY1vvL+ttbr0YPZaj4RbAHRPbnRCMSykQ0SPBL4q36O4iH4c81WY2TMLL2oKIOkUl
griP0DKTkqpXxr71MfkPQrWGDAPVMjYLXO3Yd8PJajT9ifBGC3z7onsH28wZbMps7SgFkuTJbfVW
v+GNahjXViR1VVAYE2nCPvwBwAzC6gTbXzW4gHSIysMNazZQksppDmQMilbdOcA+t2O8k9ucbV6h
6yWa7/GjXHuGl0zhCdoNYz3TqAJKGoWUFSVyMzEkBrG7FprQPQQMvpP1P9xBl55JOmAPDTnmN7kb
oURg/cxZuonv8TtsWN+jXWfrswGDzWcClCwL9KN84AUzTYvRpsTk0Io9v3sQJyecofn+5xG720gm
MhUOpeyNbD4z5t/aKT6QDaV+TEDR5JccncxX2iisqO1zTyV6ef8nq/yAlu2ChFXkv5QMQZRJyMt1
yqMuMgWawVzgOLOdFN5TV0VchvJsrMdBMP8gRLd3MqdwapJpAJ8ur+yZ6BWDhb6bHLHReSom3iFk
QJUoQc32b4RrfBBLDdnSnY2LqKI8gJUzICzYeUdfq2oLB+fBZaYm3t/YlAtDd2ZPJBZHljMeQ2u6
OfRQ1ykK5VfVd3Rl4hc0r7X0tEXWPI2MhbWUPDFDrfAB514L8Nr8oJIfvRWnUoZhjAi4t55hU4Cb
y+8e/K8RjIT/gwEpmIS7bePlv5yz1GvK0NOmvUlE1nuOoTnSKXKpoDAMO5XaTu4RzB5WQ3Sl3BXk
U7/0oBBW7DiRX0DXZsCvyKcTy3MyDamYcY0FwHDHollxNoxZpLv3Q+77/xCoN4zgYcflYIkc27fJ
bUIqTA1Zpc6XA0UYl787R4mUHylRRLhEtAP85sOnIaT2Fn9L5z5Xhtx7WeowV5O06CriAVC5Jorx
Af4mEkUYcwOQfyJbc8aAJ3l7BIlxQ5Kt/tSw8kat4PaXEIgip/F7EB1oF/kRZTVlnhk8iuTi7ODW
RwJmM42yhuMYvGdjj8wZQGdhEOjOXJ6YbIfZkPU/3z72ZmgETOO0TDs4m1scWBB2XdQsKM9lyCAr
KGx+7XBGiORZ6+kwUTOY9d+qT4+mp8yFv7+fi7y4ANmdDaG2kzsoBG95EDYTg1MKqzHDPe3StoqP
SoaW9jMqNXpObXJ6KuJ0y3jZcYJagG4y2pmtT+vNvr5mBh/yfqppSdNYqH3RLnJLWVpC0YTaG95o
ZvHMVb9Hojy2IwBCLYz1t7Qfs99f2ImGiSN8dwrBu9E0VrX1slz2ByJBgATGli/nSXb/KeAp3kdP
4SM+rf51e/g5ktK1NFeInaFYKpjDIdQ343aI0mJVt2aAXFTuJkzadOUXTk8Wz/YMStdOujO+P2qn
xqmfduiCVUzl/e3/iJref5AVZcJjOad4HF9t9OABoXNVcPw1rk8zGjXoPuggW1Bcc+i6RG82WMpA
4h7pcSRowMmGtxfoK2v3fnHG/upw+QIbSuiJmQlctyOyRnnVQbdm3Ht5NUOlf35F7GlLvGyptNhb
PiFeiJfI2WfdC2fWPxwwoNm2/PVvFty521GylaacW7zWuN6YMqwVyJGU/H3jKI43/mRcLFmDIrYF
7v65sZJPqHD2gc47DzTNRg8gq0+7GrTBegHPtO5aTQMJMrylDINq/tWNTv+Cuf+qFmSEZWQnhpLH
Fcl335Wb1VbCKuVVoOQGhp4ZpLbsqDGG++lbvY9QluPFwN8IVAX5HyjN/01CYFaBOk8qg+Zjt5tT
2lzJGgvNAPazDJvhuKzNxHHlwE3P4RB2/YbkD7jl/niNj22ktCamdYgFnC46sEJ+qBLfBeCnZNhh
WqVjRa7cK68mWcwJqYz1EvRUZH8HaZaYI/27dV7PrbGhMRgjRZwr90qO728L2RmFybqRua4y6Uq+
QRlA12glj8MzHDx5PETSjVoPUaPcrDFhedPF2+1PkkTT+za6GePoITnGe35LZtteqb/owigXHdb1
XItYkrEvHmI6q7aFUd3sUw8c9LvlmAdC09UBJU8B7AGzojGxzo+IduZIAHdLW1njkf4yqJnSB+Oz
RTUHtim5kLGoqbx8Zr7msmekn9eI1nfr9lVMhuJJtaiXKarDBS93w3kPxY6NaVbVvyM8BVA7dvAt
BSzQ0sAgB7G8DP5grb1pWOmAOxq/zDCkPuWYaC9AZlMqWML7LA5nwojPSRC7/8IH/Lx8z+Eb6ICs
lKlMOZjHQmV24fxJnOZTWvDV00QQAKBgHx/oB+/9MXgktbsgt4pu7WrtpnnsNBrkEUZac+9nTPh4
V8fdOfH0irMIKlstyt/QhXZmWZoTVZb8407TtssI0cUAU72pm7rUwIczdrmq4wbtp0EzUzuBvysp
nN5fDLpwetSp1YTFCrxj468O50sq4H8oPGGQlh83pqJgSJxBVxftizN0HexsnIt1IA+Hiq1t27c5
IXcmnKR3kOjocvaaGq1mYLjk2LzLe+OwvEnAYvl+8nMdu/9QBjo62hH11qOuID7nFwIUh+lL2RUK
ssKSb3eqcTqcL9O0oUORlgh6PHyB9ykNWmMb4TaMGaPmjlwW5KYLpn8bSoSR8GsDXbTTDuooHFn3
fyIWx8GKKBY4+IP4M5Sgf0i2muc5zOGBMMJZ5AswOA24jyRWylfk5CEsEpiN2ZNZm5+5+H+TzVQ+
tVSEGD135LvUMmj3tvOLsxk5mrYCptm7JHhczkOYeSTSaDofr5YSVKk1UhdOPTGm2UunYXzaMMN4
pi6TjUFezk4dQan2xaqewvkzMaEb/0Auelj8/YmKk10B7madefxXphH8bmrJ1HGqtVtGpK3/93w5
SF2uDWTYCjP3WAg7omlLwK3/K/gAq8CRoFepV6vEWgf7WByG3xTY5Af8RHjsF/vgHa3UO/oSKu4q
TT2xQRs2JpkTBky/sa244qKWAWamNKV+p0ebTUPqd+I2kJUpsRq9CW2zIgJWJhZRXVFPtM7m2hUs
/Vb/kKAoHkqA1LLl4C3aAxM1bryIB5UBvpYAWTL9WRPFKs4wgxd7p+N3XgObuHM+R3Rp0o2cGaXh
16THnGFGHCdgIIJiHNtLRIorfBHvNIx56osPUhdCyB/RwjMN16/QAXB4El2n6bCojtrhtE90BAS1
Gp+CmhXjObkgnueVJmAccISkopgCD/u21NlW7XDY3lPKIo9Tmzk9XjaHhVymUyln2ogipFugfRdQ
vB6ksJELv9asHlA1WtM0DQejlRM6yXpB+av7X9nqVLx6eDiN/p7e845iB7GA75bu8WDIh0nbVBXp
i+dabyjybyUg9QaByQfzEnkNQFYPcLOA8L+LbuHP28xHleg6UoYH8pqjecZKnbUpkb2FbMyUrbQG
VY3iFKxk5vMmt9nS29ByjiRjxkFtkSC4uw9pyzbtXkCmbcof+N/fgpZb6Im4H/PW7tWwUARGVryC
cNv5sSnORfKVGTH1xvvk2pCZ1D2aAFq/HQP0wjcEr/CDOOktc3Trn9FZpUiEhBu054YuZa39I6C/
23C71dHNBfo7PIsVOHdFg7Qo2bqj2OudUrJki5VteOZMXlWdsiKnHjAXQKywvIrCOZtEUHPWOd6U
Q857hYVWAP2DDh7IZdI6MPJWLJ/qPtjoTVUqH4eZGX1cWa+9N001JaStMQgVRAptEc5KkQHXPhFA
TU2nNBpnlOZObZpkXMul5whzWFingIRDhoVWbaA7tKoNxDsCBf8BBRx68jINBvk3CO449Dm8HUQl
aFtzkBKKc9sjuRRFiYn9/mou4ud6ImR9yDrcde3uFSDJEzHLIuFYF04yEK/un312Mr/DwOtSyKw5
zoC5TtizHbcy2DUXobJgC5L/v+hjk7FL1GCcN+XeIn2veUh86FR5WN80J1M0+JYz6zpk7NQVq9Om
7hMT8D+4/TYacVkwoQQfuyI1Q8TxdcJ7Gq5ywWfoUuq0xTqc8NpTlrpBg7KByH1b3HdQ4uR1nMOC
cLoliNGZDM7dntAPL1Pni186IpZyBZkRz660KmTbPDXdFdpCjM6jqPXrNWRe0KZwA6LtqDQaOwcN
OycTXMSueomoKABTXT+R/UfKjiYCQ481YAd+cVaEBjKGbaVdlQi4LBLmbmVev0Ut3iIlF/TUPfxV
gmbxSpIOMB+yFd8qR1dbBcOvhXb+VcHzFpue+bwcb6EwYBaK0VvywMfyZfxCpemnp8dRT/Op1gkJ
1lGhXKyuf7DIiBMCZh6uCCIcsRAy44UQUsxiJgLqeuQK9nS9Ji3UqaWJebGNjbNXBlbMzDu5QTrl
ImXfUuu43Y4ud9b3N9Z/jWwQG1aab7SBioTuahKRk0ld8KsKwr0d4oN8tdIQXKEpSHL02RcwlGTg
dv6uNtk7wNvA4pGKxbobbDwG3+BFnLKM6iX5OqtHO/VmxVFmzgDBt6oRmThu3XHTkQQ9SkFBchIg
HCSOpywBdfsHXHaopgF0RiMaIFXsb4Z00OBBEU8unRaOwCzJnliD+R8mZAqodeb4OhE5/v5RfA+J
USUz1LiGU1G+7krKKntzQjpNeovvyR1V7X/UUoHflqMtUuOFmTeVKxtuyFz+ICzXfS9gFVXQqsO+
P27U6dMH9DSnIc0+pQ+9TB17ThVBWxyAfYapTNNtw8hiFOz+Q8CPwA3cpCCmy7oB09KZgvjWwSua
LH9hKEG3R75BfSlkN+1rEOUaZenX3HG2Xs9AqvRiHNiglw8GhaNkoWgX3kvOqTOpX3Mz2TUP6b9w
a9vaGnZXuHpj2oqcRaDd5HjuHJ2q2NYnuBcrkyprbR0UFYqL20tfv08N8FB2fReRlHhlu3l7AEUE
zrWF7ioVX7COGlXfPH17agYj86uLGo/xCN5ASZIDjUnuycEeDfE6tPpdRTVyj50HePZ3d9yAGul/
gdHlXGyfgIOtHgDCi3AeiU/okrVun6CTpi4725Cjf9ftgrcal0lXxO3ObBLigfxnPrSoJM1GoN0S
w4DtAe5wqNpjqPa3Ir/2KbV1T2YgfRsH4w6StEZj0W5qjQnTBQcPKuIJUwMNNbXIhx42UvGYkwwv
O9IQX92LeyWREBgA8MReRPCU9uJgGokdj3V77BTQCNMACB0Kq2ne5imQIKUNC8ZHp+V2yhwquJBq
rrtGujvwGsrJYLwKAKerAwbnXlhZaT/nh4+Td68WK8k2JE10pmrS9ZKCSJzhijSD1toO4643xZmt
Dj65R2czAbzYJwiiz0OLPexCmo9Nw/6smjs0WXyggN5TeuzozaVtfmYJhuVn5roi/MEScGmf5K56
P8auU86DZ6LNhep1RDi9lkPUCLYZEbkdYTrnnpGDFcw1gsVs1Jz3E1OQg/sbCN9fc+pwLovrJTvc
bl6azKR2cOhvI2X7LugBXEJZd2k2w6uI1C+sPksLO6JlKt/k/mgP801e601gJ1zo8D8IRkqsNCWs
hu6b2+A8zVf0PtCVom+Za8nzIKYtiQSdr4Sasi6ryHuZFUEB4qO7n707gnc8fZeiM0AAWdqs4r4f
XYnvYmBG/89jVLgnpmrQ+Y7nMZxlahaU4TNJHD2bB6JhksaQUCgn5FmMVIBVDv9XqSTscTX5F1cD
LCZwvqs4kaXRY29kgDCp1mHhjd1nWHtrmA7MvEdjJHp1xetkB3Q+/WuKHD2Om20U4z+RvlPnXq37
HCld8cYmYqngURhWEo7q0HbVZmy1w3bRsy1wXn1ZUap1CDpeI6o5pKRerrfatlFZpUH5u5lxr1bf
e+gtA+vioPIxlf36txV/FuG5ee7fv7JKPQ8PQsLx9ZKWjYDzitZiS3J1l3Y4qz6kY47BUyrsKHjj
q6Y+y8+QW58MNK1jxtwBAN1fU3mExLPH8b18w1hrqubLArcL4JteoHvNPziShjCaL7PWounPEKYM
iWIV/zhc1fKHaWtZYpeYKvcT9gqhPvlilpDzhjSE+R7O9WWUON3jAc/OQCcITbHS1R1Kg5Y4jYad
IcpZsP7xgkP3CRUh/92p+HFlUahfTgCgLfyUs1a84j+XDxZw1jQeRcxQ/gznFXMZF9pAQ1OoRJKp
hRuLSjhBg0PBPu+4vzbLiWC5uWrrVaGIPmEgXM0TzspHC9v3DUAzeDLW4xVBE1wMQfV5QXanM82X
nk9gXwdFx6L5od8/SHbXsRTOyFjjjjeTtFx6Lny8cgJWyw5ovSYcOQTwPjtWIet5rQob2wPfpLcU
t7gvL+/sQwmkQ6VgpE7XFgEpOaz6Z/+cD280N2I84pq+dDVn2iWFLFgKRp9OROGLnODmQsjsMl4Q
PdCZOqAr+cQOu/jFnG/j4lCKVf90N8MdKuXxfZJjsozN5tNoH7c5AsckurZ/BExspo172azL87Rq
pf6iG2f6hZJYSepMKUuNeBM1Xr2BUv1QOjMQLowz//Ez52EwubDKgGAKEvN2NE3WnYmsN22k5nQm
a5QFG4DitGztQXxlgJ8LMdeXJj2izrU6x/1+oIbfCu0/Gg2NrXPC/3657D8uDhIjy5J3NcUb+YXP
xLaAqiNMkTuRlyjAj+32AJknBRMwzZHM51WfYNUP/OFUljasCwXv9/4nqKWN6CdFCUGCtanYUvTH
QC2WZkVubDfSYCRa60b3p8QXCHhpd9g3/oKofWx+WqYtnkmzLG1jMHYVC0jpivFHxL9BpNagcyC4
SBXCGnBRTL2ylWqere9boHaGlLgnqkU4RZKS+uuuXd1CnnAmXQOl3RH0/JqrlcfPpbKPlgV1AVEd
PowjVa4VeASXwfGhgNSeEDB2Mh2+B1wl/VpI/ung4y04IFog8pxHGzobqQr1Jib2yxOlwCBYJXj4
erdr4AoBp77b4Y5VIrkxYWvVEnLFeOhLy0pBrgH+sCkDosWB1ck2AyW8x2x0hHPBrEabjtq3y0Kz
kaNpc0rwwtL7Naly6J5bsa7cH+nwcnXr5oooIhcK+CF3T93O4oyxUVLeYjJ6qp15xEmnvNs08TEI
yoNDia/FT96Fn44zJhS949ipiN4458GF2WMLvTWKWTFTzzX5iIB48wTOasdp3pSaUnOAOJXh6ta4
yJk49eSCvC8ASi4/6jEOHHwQbQ5jC0Bn4ivNfEpTcP1WyV58cCRKH25VY9eNymCBL9POiDBAvf/6
gPa9AlTZJqnRHJ+EO0UOrwLq8hwwgNBVoTOoGX/LhurPsSLT07PDgLveJFMzNeGRLYtSrQUTTTNP
qCLMpPKZ9NaBUtSy5YebtO7Ow83oQqVU5lJ/BkckklSdvdeoJHPFtq1VFP5HQNOvNECzInXhzm1i
H1hYO39n1bxTuM6G2f7xpv20eeKsE/Ia2kFXXdQm8veO08TztacKPvNAfHdSZMTpXDiu+3QLrCqh
tYl4/aDQ2mZF6BxtI7gbMJqQZup6Kh2LVb312/DWDdESnvtk078SoPClDXA7Vpjjj12QK2/pHvkX
ytF2SFHpFASTUvSNH5A2FM3RwG0/owO4lIf2IHZ0AhoAq7JlG+rNHM3C2irbbFnXvIXXIRCpfy4L
0Ezf0kGcDWJrlHA9JrT+houYpDNbpN2rtqDZqQ+V0HUme+xZRS3Esl80JAXKCMsuYVedZv5WL7ii
zjjHbwADEzJG0mPE+YdDKpqAwb592zkgTke7+Zw+CFXvLxBKiK4LfmKHd2015V8GPgKY6XWLF6q2
5vo8iiohRmsOn2OUFTgCMINJRePjwf+HLEIqTlPLWyHPN0+UoC+u54LCzFbm1ZF9X+csGSFqLmGy
vZPpx/avOBQp1nNIPNWXdQLzMWkjtTcH8wb02dDERBiWGor3mI/y9t9iEUskFeslK6M7mlHdheaA
C2w3bCgRINM9eREfbPHrvfotHIPp0JvIln/4VcYP1Ppd4MaRpDdI3ND4o7zx+hpb5k85XhdNwsjW
7wiYu/+crjqYaiVgccJdhoKMqIR99kQ9QiNrVhzqaedqk7y6O7f60GVzo3e47qwMHTwN5c9qi7as
9nlLzUr3pJITqrZZ4KLTLR7kFx5rjdWIfA42Jg8Bv9epLkVz15AlZNdwafRKfgPLoqOshrFOENGS
MWdFBuDfR9nDsY3kRiUIdQH9jIV5ovjYDI1zEQnCH3WLs7hSBV0+7rDIiQ+i4uBDDhF8MudxHZ64
t7znkQPsy1U4dzYucez+xfnTrb9lqHjmcyvdum/kijSt+nn6JfLCCUizJdiUg1TWUXrB40rAJIyL
YurhvtW8aFZ3j4Oh9/UON/kd5IKw+cd2H2v+dgLREttUCej774RAvmG/0gVdk/v4WemBrSwNdVH9
Ps1MVsZ3TZThQ3uuwM49NJYzGUkZQg9gkCl/yb88NQ6LX6i62cLYRU11PvyUQxK/dW6V/vPiJ6NK
Rp48havO7QrSgCGkUsXJZD9rH7Cm40WLqr8TFpNcC1ryRrM+mGjjMhFeTifX5QFX3ld6WxPKLKV4
uqR4oj9FerQyHxrzboc6P8/yr/9E3AhY1zr8N2QyGXLWFfa4PbJYTgFXeG3GbQxvTW60Dp7O7fp6
GbXv8BYALVt8y/dUAfvmt7l0iMadd6fbpO+wGPycAFX1pZYBfUh2lESWs+6Z/6OkQ+wL+BO79dDu
Io/hpmP6BluqZyIU4p+bmxMMJ8Fjq+OK/A3bcNMmE7MiBws3N1vPWAJ9WMI7oXWroueqhpmYumWc
+a9J916pEREZqmzwP9eHezC+99EvXFRtx8oPu5tJfyxTyuNhbwy7x8jB3sD11C+MBbq3+u4hLX+u
4BhjjHH4cjuaU7ofp5zEKvSGZYzw8n3/onC/BKQ1q6bUDV21guGFdcvF4t0IpoiOnBFwSW9AuRna
ucHSRkipCYx8BTl7ENaAjzSiHNereOV8j5z9POAdU5vPhN79CfD4hUiOwEXzypvwvuqBVddLTyxi
4UcMkC4xaixMj5nFiuStbEmuYWkN+KzY5gl6yZ7QyfZYYAEJ2mV7lNJCG3SDCCQ+a7+w5CLBkG0F
t61PIpmKMl1jHk2l7izBESj+eXktcxOlBlPGaHF7nIqdR94Cw/Un9YYV+u9hUKOI/XeL18/CP242
zFj3BHUy80lBvRQDXrPKLjHDk1Sqpg/nmRIryGRXuV5thl7QvCgiFjfgs4102/gWPVsKoSjdhbfx
uEpbIw9+S/Jw4zfbqY/4YiX0gWTQL/Qz28WwKESSwmsYJO+5H7woQsXsAj3W5nw6uvvfdUdvOWSS
pMhr55KxK94C4r9gc6adDjR5ihIduT2ZCmAj6iu5iPrJKABa842WI4xsPFV+tJN6rC9MzsR1jclS
bpQVQaClVcDQBRCbvelaqpRsRm6mt6M5whLS39gvl9KubgOQ0vsqEM+ccRSgq46mD3SilFnbmsbf
jrcI0b5aLhiTyZMTcG1OgB0ozdB6tAT3/a5QMuXEEGCV9VGbe57nYieYYkGvFaH1xCTUKfw2/V2k
r+MdwT706IwEC0GO87q943w/CiCGSJPvkiSxDl2wwbVWvcWxTXlafJgtnFRC9i4SxVSi9YllinY9
Iye7lNf97X5yg0eAT9i2UhgXj3X+NIohXYM2dN6+Kef3e/Js8fJQCv7K/kEJwP34GSDuUmChLPFn
bizNMjM0EoNWoIKzSDsd4Cx03Bb4nSx1YtOhUf/C6HePHzKabhxPfM+SC3AljLqRD3lsHqONI+dI
9HtLIwgukERDGRknW5KiS3bq0gQ7B9381YZKdpce29TKZNCZJuCOcXNuWf7IHcCZYfFfjQl3IXGo
wK8vIcr9BqCWt2T6kuJHqvzpTMydrj0bjXtJan/idRyoJyUq+oCo1+bQFGxQNG06mVLtBeUTT/Ls
gXbB1a0g4g8fhCGeHUi4lCfAto0gHvCex4HivwRlmalBp7Y3MtY/HIquv1Dg8Q4POQt5Ni6RmAeX
/XqmuTD1V9drt7E6tTmgbmIr34LABpzmx1PCRHBRPaDICmuJtZDlpO7KEcHEJJqmUvWH4w6t3LL4
Zr2XwyiJJpOZcVSFFlBve9aUru+CKWhaQAc9qMognVyHsY5FtBtpYi5A2h/oZdOG0is6GXsp0UCq
zTFpPT4c6jy7bab5fJPPf7z2OpCGJVT1ddgYZyOgoTj11jwCpHldbIsNsDONdyzrCZtGKVvbOo1F
8iRW2bi4RXMgAXCW3CgdDCfWwWYLFChbJwe7+3qM1PZWphC7NIJWDAqbBxLurYODGVsc+CMtakAT
JflEGXSwd1TKNuStKQLklWdFqF8DF38uYeqdCZT3V9cAO4z+ZGESVoIAfaaYXptesP8tEI+kPda8
iHlZ0w7vtTYibC/yqWRedUb48SZ3oclq87bYbvRnQTDhNafzNhAFvivosf3Tnnx4KJkJZ7QfYOvZ
/TxRqxOxBPiMvJtGfYQ937QU98AbemdUJRW1alqdI45mqaZ0TCxsEg6V47VHHHfaQ1TK4sRIs66C
kIBa4ylkXWciblW9bRAYs03wyLZ+rq7Nmx1+xHPdexzsqNEifCuL/eTQsNrykWhhKhs6N2nN+S8a
tMo4jelImLrzZi1uj690Lg+My8Kv58arqJhi/j00j/HzysPFLJm7q/4d8FCAJi1hPUGRLw4cEOII
K+wvgYj5hWC3jxgMEI/PtkSzU+zCPWSVQBNSPUTO4NorH29RSI+V9zBBP9xXjbck53TaU1qySBup
HjLss7vNZfq/NgVmvRCXX0NJuq9dg//r4Urdqpx5krznOdkQr5umtYbRICV1HJZJb3rn1K0BlVYE
0IoHCSaBvuZ6uTM0ViID9Jg2jZuEaeyjvEQNVmAWOsB/vVr2M81gXKHiwyoA+OiIMsF8QVFa93+2
uQkAdiXkliV9qx2Qk5lVLyiDFbtAhXQxWMr0F4/NGDHAf7wWxIS92uh39VUioeKtMwURsB92+nek
Y7ZTsojxjLwQHGsVZihhUjEU6XO5KAxGtEZb/Wn7O2UOiyeJTjd4lSmMkfM7NK+SNlY+CvRNtSQo
G/nVlSZ8EBJz+dKkqEm1uvcTokl9IXUp72xCypJHuBHbB8K+LvT/MQ/bJoAumVtPs8KuSSiO079B
bY9/S5zwTQurgLJnUL7EqsZyg7juOp4c9BOP4SAt3cNy2EIUOYlD49/HEpJzUlx+OViSC+ev35f5
kljVNWRU5uqyWjjr9T20ggxENyVX5+nBKnpXpBi6aKRMOJn1hoioD/130qMsY0AsMFH9AMc7ahhP
RoH+8DveXNLIwBU7dwnbAapOaeP282AEIwmvG0XHZoW++pVOMTA319xwPAe7wuEQSAs/pMOv0MuB
3VHjdNcewOMlvhJFgXpmegW/Tc/U8i5PUN0aQhmnbKbC2jj43rROjAobxoPmtn/iIbNYo1+J21/t
b1aWfriUYO+zCeWfIOagNI6vYsIwWUcf9ymRGwE8wLps072WqlSf3VGTDttfLvqh8XnPvWZFTelO
e8mivLiHH4BibPig+6esuXXE9vrt4Fy3JmqOVYKIZfQ+s6y4X4GVwUO3AlCYYtPWWwILJkfnJQlG
AeUKkYFJgcATf/QN2VuSJBjLRmDrRmSSXPMuJyogQ9sPjcgKSdewBLtLdCrGbcz1jXAY4RyK26FS
OguqHEnrL3P9wM93NREIeKwaJH9zZxN6hQktnsiv9FJLiIXLAHtvVdJ/p0ou86XWA44m39CDtICw
6oWKkSG/0VzQ1RY7Lvh4BCD7bXIGoLwAU91z448JA0QRfqqYY7JSWmAfA5vzfx+rAqAPFW8+STdP
yvbuKIvIi4ioaymZPHR5LrEmhoFXLBW5Cc07YdXGibKo+uDh021T2gIKd4MdvpEHF0fBBMdbr78m
TTck9/c4jYzvIk4rxavpbbtl6qjdjS0Vtv1F3haBOgxcJLzZRf4dfJ9kYdf/eHzeE2jUm3QsOMXA
5mGh1cVa1Dr4/yJ4vXErqFAtq9fbdigqRwu7ZRQDG7U8RMHHxuPe1BNrOKCsD1QbTa1/JaKUt5Pv
JTiU7F95Qz+d0QCCsnCyhqK/gmJB/4WUM50NRQM5qqyQVrwSJIn20mHGD1cl6lX40lR8nn3eEBhm
JEtObITLGyldZe65gFA3bnmpZky8L/fOxU6iltvSCwKi9vUpi0wJ4Wx1fTuJV6PFFZ6+zYLvJIiP
thGFo0FKJ6zcLKIico5plxt0cvDwN/fxCmnr9LLa/JWikEa214B4s9qdwj5fOTzbFWUEDteqMcor
MCFcQgm36gYUMmdZJKvh89OCSUttI0B2TDllnqsREUUh66Bj97025QwwQCw4L/YyZi9GaSNhT8Aa
6Kr56/u81h4MymwSnzXRteGKfZs/u9ZPSCZIboGZF/35vON8X7HUxDVeZiaJ+2fDmaX8exIACOBv
SdXSem/4fgBh/yoVBITCK8wvdgVIK753WG945umG+k5GEcbsk7+Q8FoyIX2oTa135F8JhPVJd/TF
C7zu0TDgrhCFM6/u3SaGiyR/f3io8CBSgVT+wadKbci0TXaEgibCNyWVOZ3XsC3rQulELQmYDEOb
3jlHCqpxeh89aog7RWHD/XCV9iLx42mdjmdRMV+cR5urm6oXpV5EimZGliWZCml5jM0VYSisv1vw
JnAID24YKLB3vWhsO44SW4Lk4B9UkjzBTiyHYHKSkbwphQmqwDJ23XzI5j3Ib6diynaq3afz6D2b
omPg5xwWphLBr7i3t5ZTLvEkTrq6Xnj5QlMA9OXKCzMP09AFFe991KPDa5aDh9/EegN8/bmrfh78
gxvxerlHJ06vHSq3Et0gSszQqRLC2qk5NszKbPkLkNiTiOvm+VR5mqDP3LFLFF66LNh0NMONLA4n
Gv34JqMHBTpD3JHdmGeaJU13BOjH++bh530YApUVAmaAHAypbs8Y2w8+uskK7SA0cZSG6Xa2QXo2
XFSG2Qd5zIXDF1D6859w38GCgpOd+3bH6T6hELNb2nnod50CBUlv0d049b5H1rI15CHDVNd+CtBf
Rj/N/UYNFn7Q5RrcQd1Nq9Wt9y9Mcv179X7gPsZse5kqh+2ViXhNRC4MCpVoWYzJ26+uM+vsxa2x
LzLtL1aUmFHjcF13h4W5D59YZftPFYeHA+17hoxq5r/wyMYsfdCGDEwAdwSX5d9TRLTgoZn22RtX
otjV8/xRK+Zj8LPUSYC0TymuSNLuXT8sXSffKPVZpi6WjLJe3Ckf1TuA6ScWIwcMbNDiA2yy08Sl
3yyCdmgXV8ajP/b4h6aaTDRsW6jrelciUg0GtPJ3tO9Mjd4y1I/tZWbLCybAOJm0l6eGvjQCj7sl
QNterqiDLT6aBxocv6NHVQ5rQEyczctsO+dnPvqeqUBgWyUU5qRtpcpbwz6ci4dEQiu7yW5pZ/5H
DhClE/1S6Yd4qgmIZajns1Ygkk+uUgiYebQlRMlVNfKBX+8viQGzakYk7hhvCf05ymshm4aXQsE8
d+xMpbOKvLKB8RMgGwq5d6sUt5CKQRgKxpGnuvUtncmyY96eNgLRyFvx7tlGoS97/1at/UWQH6kT
iraDJmVCXjGrVU7PK4/kZQUUF6AAmp0CxxqGeg2bxk+OgjWns9gjY+XyWYicUs8R+GdBFdpfLjUV
fnJAxLK4BTfw51zUHmaMNNAR5oTQ4wpGwgp9qEAQjFHPKPD7uPOC76dsmubP18RBqbKRyLgmHwp2
L2s9b0PZt7fD9Qxp457JDcUvE7Owml1FVwaCGEpCihPvViNSF4QsnS14pTzaqTOLy8TPtwb1rW29
bPcCdWEEQW2YVirL8/hjJQ5G9Jw5daGHAzYZbBrlyCCNPZOhVEho98uOHCv/j4t+/+6FYtr6k5p5
qzaFT1x+qt9+IsADQciaLe7UaoVH6d1k72PPDbz5GiK373VfRhiSe2O+Xck77EKBPjccrwUXSyDK
etXN7tyIrDSeQIH8ybtA//ybClbchS2QUFSm/6qYBRUS+g3oCUODPqGq7K+BCcWhsOVBMcp+Cs0U
oFk6oLcIemQ3k2Vnrv4xqDzZyMSI+9r432sZJ/K+Qf27m5XKnk8eu7KmlLcF3UdEvJ1LgO1Ty/KS
w2UCR6dd6BKNG8h9QMEeONQWTNbj39D/l8Q0JM3Wj7GlcOu6yTakdnE+7ufjrfAR5lRjqmj0Y4Ru
cMMb1/NuBhJjKU1qXyj1P0gNpT37iQcBgrBmz523nzkWmzJP8ndwDE2XZOzOnVx0aDQhLUia0S4d
kaIQm4KbFQNvQOkvn5r8rfC1+zxtppo+Z0KU00PBgjlvndzEvHhKA3tCjEc+EJmdB9+XlEEDEwEk
l7vB3FkgUNzrkWaZ+PERpZ9puCir0k6F43oMXGfN9vLd6czi3o1MQ3VHQibX2cyaJwRY98DPmt0p
d3lxdFC1ZjIoSYSF/ZFxEnaGbopTedZShYhmyhMohBwOtZmcI4qBKIC4PLDYn/dgijeZvlD9g/Ha
qQ1EZpr7gZJTlh8PCv3agkGhH/KnVDf2eEy8cSlxBg87cAJ1ZyyEpcGD2LCLyqVk6VMfPmU43X8W
5duYBar4GUA50Qu/A/avKq919/xrvybhK2J47jGlUJE4+uEjR6i1XgaaDL6qSwU8l0vG4MZgoHB+
GWJLiE9AQPw0z0Un1xvD4bTYaaMPPhNrxV5z2wIryE8HygLH5ezNuVMd3V1i1EJlsQIcddLcoNfV
ak/Bt0ThOwmzGff/rO2cmNJVD+2LlTM9/K1pPTdMNqRD1BGyB0mjHMNOk+hyu7nOR6zTWusaT+kC
I8Prkk6ChvcfxrWripaoY+l8gIa3bteN6rBtMzdYYLYSDwLB1hCBC5+38G2a0umhB3zA4UMVlF0L
nU3vU171AqboLfeRau2KjjaWjYZVOyY3o9qIMHKHAT7CNeghlq6V7rgwUGmzND/4OUlboII35LHW
puegND2RpO8DihWW1mNxXXCi9OntafXNlUvnjd6K67nFHImd46D0sRMJpmQwpcWgsknhTP0dkguA
zqUDUmi+RoRr2YHxxOzV/C2yKB8+YKWz1pJiV4homBhZksBvuHr93mBro1oMz5sew5VwSJFzUXnB
vCSoDA8MjlGZWvt/eCPOUPT5gjuQxRDxFwUFhiEO6z+witt0ymq8BCk5tJHWddJY62QAdJDEpMqF
y07+aaUsLGGIs/+CUFsK/i6FNpx1UUdZ/RWh0STqJuypCITLJmNmSOiA68ZZQD2w38IzRyzgsSQG
5taowxIxJSlXlrEGPLy/K1wJW4kjroXr+LMMoIJ3tEsB4UOJF9meQWnB0ZUYD4ASiA82720cDyPc
DpLAggQZe9MQ0sZ0YqZoFxOZfQEAClA7n7wJuTzFL+s1a4WKhrHYmIQAdTbkPRAxmsZ31EW5fE6I
VjN4RqPg13SHW/5TPBBt04VI/1XPOgYo6DlKoq50M3mQ1QwwxMLMeWykDPW39xCp1MQhFztcJMcd
uWeg5YVoLAKsKBvY/3eqLwYarkkRFSJe8TYffF0ggz45j2gTofrKMB1tV1noO6AomIVWoNRkbSVC
z/waKCoQWeqNU8HvRL5snlzOssxR0qg6WW8qsuyUVllF/JEjkm3A+9I83iAaUc7jqeblHyZ+antR
7h2il1ccTL5oHpwfb4D9pDYm5yAafNA7iGNfFuMojpDBplC1ldqXoEAnP7QZkpCCc4SbZyojA3YM
dIe7AguvwE2mBALOTcqnCt/LbwADhp7cW+Ix3eVy7hVLC7aHi29fb8d2Lha78CBqK//Ch95PsOQA
wCqrlPz49LGMUddCneSyae5Y6xfu4gpZtzIr74JQquWmMU+/HpHD4M4uYjryEkj+tFRqIrdX+AwK
lXJZ6BN8XSbVzFzZjLECnK93jWp0/Tt+S2oJQ5AKNCngr0X8QLg2jVmzNInvpnier7wwUn+OXZb2
6NMSCC/Yop4WTngEHbsPcIUNQ1TdwmpSkkQNgJaGuvSi63VoDDwSg33C0D74rw2Do2Us2Oue7wHH
idYtGxrHjtwXHNsNzwWeGZzR2HEcvIjDiXfUtc1/UvzO1XKWKev5YfsX36w0DNEQed+6OqLXvcoJ
lJ6f2ce8wGoGxjl1z5iT0du2bpOZ84FfAHzH2XuUofa+Uw78ffrMHx/4b7dP713REg+YscJmUKJb
5T+6NzYNoamgLWMQIfpGRSSCMcU6yb52DIaq4u0PtMwedU45fweEssALoWaaodx508GbY1x2DBZr
uZBeO4qf7p05Kca5m9WgEVR07JCz4M93JCxGGYUoO6dOXwVLfuNXpB1QJBsnAfUAmfaD+nGtZw4A
FpWPUGhXP0VqeiNjM9ysMmHa5mxFP6OXwgPgLiPT9OZ0c986OwGUMUbwhdPGZf3giIb011Pj2X81
3tcYzZW6SL7jKCGQ0v85bXqVYHkhMasfhvx3eURSSf/q+n/OzeiuRSGSYdQi+dQXxwsT385dkax/
4s6Ev5J2j5DzhH6awSyw17Ce1+PGOjUUxxKnzHycSRQc3ckZ4DrFWdsZ21wVZjaKchpVuZI4EoTd
sww1jO5TNXFDIbftJhmDMw5HE3cgNsM0WvlC/LE7g30h/isTtt3UdxoIzObi7Bbs69tfLNLQGLFS
chLGmeZxeLgMgal51hfH7XQxVaKwUBuZSOjTaz/n8bVdelU+osTUQ2CjVJEulUE3JdRN1c0HZDKa
yAkZ8wQ/1jUe6/ikgULhzgFdUT4MWeupO9jI0CfNR+SCnjV7FPVIkftdm/38yPjLhB+hP79lIJn+
FNmm10jc7M2R1WRCkYUrADxp+wWZhIhs1kKak2JUPL9HXanUo0hQ5AMKqc4BHWte4vVfs+PzhM0J
LEsd6doucvFHdV/Py9JQwvsUxwe/2MtUZ/rNZeJo96CZSb0vnXC47NZJMPTNLajCouGltOH2RUfm
QNXfOgLRkuFG4QKsmZbL2mG83dM2+DH2BzD7N0TRwMmHHbo813siygiukmcF4CVlexrUUJZEtJjI
0nYGmiR/7OPfseYWWaDFpcOxk+ty1t5kRvVqfftmyLoV73XBIC4siW2MIf7gXxjjNemHAIUeSt3/
oCVn+HOE2i2LkiR64ggnDFqrKe71Z3XAJqf9pgMOdEhg6k1v2K4tuAvcC+J1UMct/U1q6I5OoJ6w
WM49Zg5N1QMtO6YK4h6/IhaA/vPX1mU0FO5NPFumTGGIBF64bggVbR/o58K5t3wGTwx4r629W4x5
dCOubcoDzmZsGVA3+MylYnLJB7iskpmB0eG4j9jEaEVBRYu3iL5SGIY3jYDl2vxcoRJE5jFoXjWr
xcqEba4otrvhTAMN7DwQp4VT0L8SF3r3i6+2bUScSgaHuVuOg61DfEc7huKyZs+lDEF1/u6ZL++N
z0Cbnz/BM1lkSVCUJRr9TN4lhyoCHSyVm2vwVW1mq3K+Y8DpGXBfNU+UcgM6iH0G/LtTR/c/d1/x
BEiXn8yOep9xjif84oxl9AwEyS0PZVyd8Ekrmv1sttKFtkWykm3PL04JCpewfmRCWjGSQ7rzmGM4
BTGY3woIiCsKrGJTiMQGHIYC6R/4V0pV+HZmi9FRT9530EkmH0gjkz6THUZTBY7TzyLDNna4bPnJ
0eItiJyx/NS6CTZhRn7cOzxQVvqkuAb/hAQIGvXw+yWt4YbN8AG+ObbvBiPcwn/So8oV5qcAoi35
ypAnQ2ktzLqC4Q4XZxL3jkqvhdLbpx0PwCe+7WkM/QwJufQgW/DKFSTksIIMaXvhHGixWmljmrG0
ElmsyBlgsTxvYjcRCGF0XQ7swP9vWoU/y9F1E0+bK/98VOljG7D/UomiTk7+GAMzZ4p+sSORwrXS
AdRhzuVbMwXZ+CQwaLm7jDJHe/gjSspmi5ceYm2N7wZYMlargnb0JCA40TLP/MW+02+nx+en1AdA
QQSZmXP+IJ+JX1aFES3ZuUHHKLwrucIZPIM6YvqRK20Tj3ebBvLTufx3faFaBNAnT+5sdAoZ+GNT
p43J0IjedZn4lwGBOQkaPcXW0Sp/wC7FKiUh5iurbO+vxOzGGgi/D6lhTWSqozlDTLGp+QseWgxL
3bkQGETYNpDXD2TvqNXAFCIt5DqwL2E+V2mS6r8xaRFi1x8TpsCjpD7WIXa6obSflOExcpULGKoR
VmZdZg1x5jqr9X+uxz7+h0siWQf7r0y7H5aDZfEgbcDCZMFFPleiGySe5oGPO07s1d61lhQuM/v1
7lq5w09nIwkLnXhY5n9ZPthvovvwiTVo027tHUATTwFugX6FGTC06CfJ4F2qAJaxLoe0ORKR72Fn
R87NjrSJdRrK97N9JyodH7lLDS8nkhrgY8lkKyu0odHHdPpZYONUNYYVxWNQt2pyxLRbJfbo22gQ
ZcH11w2MVrabLLzgXp86J9rdijlNcDBB7lSc2oMtRedq22ZvOvK+8EovJUPC/23DyXDnKTRzhtJK
jfDdZ1PXNtA7UFP3Rp05g0MfaIZqn8FFGvFKAIbxAckPIKO+Gw6KGRWSUNjcwuolypvl4ubDIYAJ
nErOMP9cFIQfhoKZUevTQ6afJ1BwKkVJw2OImkD3I5FlOTujtlH6M0ALP8gmppcQ3ekdMT1nGuEZ
wway1j55Llb2a2fhMf8oZUhphTHzQskayJYmaXdQil/SkJr9fB1Rn93EXFpxgjK/ThZFwffZsVn/
4j+H00Si5YM7LYymYaViBiI4mf8Shk0yA5Dn0c7zNHp3lPkxMuDmEPrrQNoBghxHSb5nEPnUThcB
26MrZHRcUTeIvKvagSAdbQ8Bz9QgSaGVrgTczgCkQgQytfc2i00zYzHnyLUbU7CawNrMYqBrSR3s
X+NbwKFjp1sAVRSeATbZs3g2XN7hiHHsWZSOoFFHMoefSddE0c606hoRrUiIaihIqZXFA9/tBXlg
nts9LAeeIokbfueO8P0fcoWiffxp86p7HitstVqdT0GPiBAif49gW5uGoOgYunF6gadlpxvAgkCk
aof190yrpKCLZDf5jxE/v+vR6tdhtsmSP1itU4at1O4+7gMho4gs+/FSFlZNsdnKeQ92PGnQmXZS
jrHO4ymOWfmPRgmdTQCBk/lNtEIbkdxmgOKwW4j3PsN8p8eG/y5pqvSYKPpA00gA7hedOFbcf9kC
yUdOAckFMtNWTTt7KlYcPbXBhdi+1lcYc/9IGtZP4muV1ckq9N3xrUUjFvUY5gV//4060kINSTnf
ARX+xdLP8Wunfy72+tYBN6doNb/qtIclsIe4Df5MnxGXERUWos6cUaaTPibEO1Lz7tavhF29kcD0
oEnzJNKzegC/mVTmisnXNe9NXthWlaQr1wr0IMZz8EQQqp2zJ0LMmkGxaUAjElLIX0VGPl50NXvm
m1363yOXJ9p7ZDaEJovVSr+KcEx63sFzQK3COfMp2J7mmf0H4pvrYmib/Ai6+WCCo2Qznml5qb6n
uNfHd2DLR7RGWT1nkrZ3bVjFZ40GJ15mvwRI9pOPKowMpElrPGJ0+Ww6ktHYYtUJGhu8jFjD2ki+
vnbwEON1N0aktAjUPEJ2vHPWhsCi7kKm3NMliaEYvrUwof3evy2hjz0ZaHck230nCXvvvpFEgpeI
XWvLoqdyhZ/7xZ7+eETMYQsimgZs3LjedG7z3fYTMqJT5ZEyJIzPuJvSRKGgx5uA9UsX2OOp6ihJ
n1mm3a8HetK/0jKU0k34oc60i53d7r7pQq3y/Prpk2BUQ5zeMP9sHLIFUTfXqCD6rw1X5r5hkbUY
xf2Xk/ogDaoaK5gyZf5IjyF9NMX6ThKoyPHxQbtrFen08ziMHSln5fvY9G3nXwdJiX+dzr6l5wId
cC7tcIGhBgIqSyCmPGbOsZyhzGP0+VEuMlzhvCdryvBFJKhnbHW8saG/x3+dlsAP6OdjYQzg0Vhu
x5mljK+uweTkJi7YWCvRvyzH1GaqVcZJcXCtf70q4cp98Wk5Uu1N4W8iJqffR+MLQ4iXbamJnwCP
tXWADRAuA20IOJ+e52S5M3HvmSYwC4vXlmjTcBBeFTMZ2nIh5emmqfU6bgmtJoSeFFyI8HrfYQDe
MR/BTetBdVi4N56mID8+ypJdEQFvvGZWZ5SjIfWlv4//u0wm+LeQef9Id2xlbzg3J4H+OaPIhRP7
cW4bosn/Vhs6IWQiGPWAZLwvXhVbfnqVYjZ9dyLRTlFO44oO4q8hK6EjUtxWdu9GU+SilmAMYUKo
S1Fh5snhD3UywANBx3f+RKRcbASWFuIMOGXc24dUQkSgaXK9UCnjYkE+q/bXVMbFbN296l+l/Mh2
cYlB2XJ3NvLULZvgG3/b6MT2iLs6JtgHQMagPW4zqt6iFKh/kzP/NI5QTzEFmVKHgSWJmN9I79Px
X6/vy1UKNvJm8eX6JTDcRNPy5zzLOkCkaB14zqMHsV2EBhl5IDzaIwdLF4lLmb/LsM7eT5+b+Ywk
QXzgJvItH7yIEr13tRAaS6r2Tgyu+rovdjpFD+np+sVlvf3SZ9ddTOqsJlTftbF89CVJUcdxPjdJ
FK4VSTORT1+BJjk0kX3xdKEArXaa6zlxZ6MQJBtxnAWNOGhqEFUmEBEje/zgt6Dfl/0OXK4HR4Rk
UaALmE0+eSkStDQ6bAtWfB/1yR0IlILe5YGXcAGzsJ7lXlryLZPGb/90Gbpi5/TfX4nrTlsVt9i4
n+Ua1DIrgzDwFq3SCt8+JOMrw8ClJaE5o8f/q74xpziCvilXX+k+DUMa8KwouFveA4uPtGZgTSJj
E6PeFrgptGvNcF5wFb4jOcLKKujsiZlqiuLWbdMbG8tCOiWlAeOQUeD05/aEYxVijntIzSFz339b
cCYUzM+AXXXg8GJfOAbb9Z8Cf9MrTI9hp/ql4fEF5vIWM/isLjutsplfsRd/5ExooemQPCysCib+
wIAMmQn6nC8VJtq2WPNr17/dCpe6Ma3r7uWy/+KiyOJD4ZOjP0rSfH/9a+VsYZToyFDlXep2CWJw
AjP3d7NlG8Cvuxqr0Wwwkiqc0OvKpyf25JqwHrZVkpPrUtIMLXP6Pl+YuiK6FK2Taj3PGsP/bUt8
p89WuR4Rqp7wP2EbQcxbvH1t3j/nw5MQ2vE120CL2s4YbHSi3n2LTBdIFTo+u4XXPQ1D1y9h/UxL
wPa2o4Go6x5NlbVT0vI089aYMBWn6R2PdIHXl6xUfoMqlGUcwUxrBCmXiUtmsZZ1gXJ3GpYaN1dp
TLd43qduLpvSQJawr2RJXbyAOHzBAlOXgnTT9XQe8Yvld0pysZXdwuFLMk47e4ajFOV3WR74eWLZ
JniZ90ANgsi7cZo1Q8ro35QtvmB/wTkGekE0/008WnDAC6MGTCxLtSHJDVDj/6CNJ59XeyAggOY0
XDgZwuWFTHG5r4Fuz/zA2MorYdfsVV4nXcqeV5dMru0YIv7wjTRFNhwUSlLuku2CVBHhFJlB4fpg
vSGhXX/8jlAE7JQ1BAFns+xrlQwEj8ViQLOmtQXAj5h+rqGefBT0iE5vgljSBNoutLpWBp//e9H+
MbC+RutkfpjoqOcGk5xWCXebQkYmSIsIM+jhwU0WJN+oG4KTSyvTnaoacgYqrXClQGGO7S9w2kiy
KF7geM+RNvOeUnAr91CC+aKB7XBIbyy2+dNDqZqlkHUTQgSv/rAxWdgJ1Cw22ySfrCsEyNUjWoVe
YYXgx6rTHBg1Y+T22WlwXcssZDFl2L3zDBdfiHYcp7SWnnaUIFBoPRrZOg9Np8slm0wmoqYsEgAN
TUHLDo3lUqRDQxGQk9vShZqmeB9v/iPTC+7JviMSJvSmvtlzTld2WXgM4gm1kFq6zAvvI2suEIkV
+WUeejg0lGCwpfPlUaYD35o6h4c9T0xDn3uFauW4TxM8cufzzr1TifEy4iV2gJKORpsLFhYwADtg
rjE86FV6Myl2AUpEzDxHhi9OmLElrsmP1+Q0njjvpFyHB7qspe5bY5Xg/Eu7UdBlYCKfbeIJo5Ps
3XXisCraEtYtTD+RFnOrXE5V/systqbKDJLUJkH3+jELFg3q2MlFS80Ms6VmH8TcqcPb2dHa/HOQ
m1nfcKH5Bg4erPyzum1FZGQvAGBdGFFaZKyqN4rN3kbM6PiZuGabyvjILIupBV9bGtSaLjFuZ3bN
cXF3J27D4TVlTKSPRFVyerzdVOV12dNo7mk9wnzYD+oKyh+KVhd4wCRwOtl/l3gvfr7t++i1DNam
HRtVk/eHSr0wFA2eZcnCCc8KzRhFaEoAErGbbY+6w35Sy4DQSVMoiCc3V3LPn4969efi0Lq5c3Sp
K8azwuK8gZD4Uaa68EXga7/eYTBgGdBFuugrChc/pfoBLEyQHSt6xEpBj7B/z5+60EI3DeM8NoSw
hePVrVJcmLIPMutplVIhajqpYnJcotMczLdrzHo412iz223WHRxc9GUS/aFgpLn+oGDtqZJ51NcW
6oBom3lj+6noTyoicGvOrzQkyXJYPv9o3Sn6x41QQQtmTy/6I5nzcnfG4bpPAWPyka7kDEhiS5W4
3Orum662dlIK3YBq/OFbrT87GTGrEyf9Y7r2LFckGTzdlqb82phUpc5sMzYwl5ViJdepcQBvKThY
zJKCF9XZe9erp/VPT21DnB0e4gHJZWY4Jzc1VD08+FSl+3Cz7f/GQV82gF0Ambb4RqnqluPzGoii
21lSguPHBOs6r2kLxYYTvj5kVAq0NopZ2zgF8c83RubvU65Bl9r1FQK03RJzuAYidMDoWGjM7XkS
n67zD6ElHL4mEK9xbcAAnUB/N3LfvP5phD8sHDXuWcaWXx5QzdvOs1XE13WD+Sq6yNrOmFOUohnb
U2A91ALlnMDRVgZUSKsEXmLfsa5jHdAKnMdW1nm+lbRm9/piMhYlpvJlMBrRlOKHxoD+horXOjBn
15JKbHaMHVc3wZ/G4twyIZUDSMoYImxl6DHOepvNBYzjWRZdrfSe+2QCeWm6+A5FoZcRkmyYMxGE
DV+8ZaBeBZ93NweZ2758rGoMFf/BBKYpcgRsHu5hOA+Pv81gsFjKcnULkNy206wuzqmfbATWx2qK
fZOPqXeKEqOpy/ubgbMDY8VnoUdVkekcGAWradxHT5c89HF7x+hh/SKxSAZBVYUMhw21DM2CeFjh
qTpbUfFNh8zX9UuzYEfBS3b4BnGWo6Y3w2ZctYQ2sE9wMFHpQuhl1m2SClzJKd7BiDhQYMxpQa9I
CjwBbwFnN7JrJrpnYjLpPtErsOmcjcO+hYatZXko1e8FnHSwXM5JL8quow5JKxCNUAfGgzl+sXtq
xo+3kcUHRQqLx9bI4VrrnQ+g7+SgbFhM0J0/xsWMRWl8O3vowVDhOgi0L3gZAUc3YubsVkUWjYlR
RHTxPg/fer6gGvgJHVnBL9PZL0cAUPPHfRqyVjXSv2n4lurM10KxNmBoXIxjhlEgpyG0GvCQr4tR
tPe4uLVQyNdYagDaLKBNgQeWOLnvWOSKHFEKgsZtLRcnCXmFSoO4dKJxKWwKmu2cU0Sc1Tdtf/mV
vlFPSt1J3ndYxaxWRX15J0sHSMhVaW+q5z/5cv8awFfqDuVQdl4fNpodfJFioTPz4fT3RkZa57Aq
2kz4po6SAyNZiTy3/EibHxeVMo3nSGuoOe4n5xdha9n9fzlKRqYO1X3dUg4mMOJGEfcpKVSa7cpm
X5YeOpKytkwwYW1cJIxcArZwxHa1ZtPJzLxVjP10Su+JumKKBNfCvHMkNN+AVoIOkUKqKMMJ6Bkg
4SPGBnxZ/15Is9ebdHeZZpxK12K8DjhLYNfvk+M+nGZ3FZwlBqbxjCXJN0GyD9kB6UsYDK/0onnq
FJdGxG586nQPfK+KQZbV9SX/a2Z/5QJOmns1XEimedKEhRm5mei62zit7o+OEeb1VJrxqQhN6b0N
aCkF5wIMbD6Q9zwLrXN6pYAAVvu98O3JsWgxGrDda3/ryDRdPFA5jKyD7+M7vNyhhFSrY55TIN/7
M1YG0Z2OrAZuY18qAxDLGO/mbF+YKkKHJsEWvY81OBrKdhTfPX1HQxcWhoDZkg8ZW87qbDZIKuKc
Zt+DNCra1+IezpT5aY+pY+hLPBwbqthkaciZYds2oE+02kut+WnuHBAK3EBptnZ73li0BSMUJ97u
5U+PXcZq+/2UB8qor9UXdmk52H1bSBS10Z9wHpUcgPZzeQ7piVHfWjLRhSIb0YmHVN0Fh9AAj+O0
RM80MUiOoERg2beDPezta94ltEaxGD1Yx8G8u15BqWaKH3tXchK3vo7oPIwlmO9Yi86dKKHvzaTZ
K6SA+RVjktOuig43OxZfNMc2OFHqiFT1DqtEGNyItEHoDajjW45kpydcUdBkWtGZgD2pE94Xt4j5
qQcRGoTrWkZi4r8Z2bIxH2cbtsbYcqTxu+5XPwnmLxQBwtur0loQese6cQC0t6WIyEdZ+/1UJpDL
GZwnKP4Lc6NlkmEx7jB/i9tXTW7sgmQnf6eprhWxQuJHnHPlMWQHRoeGE73vpyC2plHtRNB9xeCR
FftGzyLgnnEtqG9LQwA7K24O2VDquDdqvM76wM8dsz6WxLmoMRF/14I7yjYzXFTKluUDNBM++QI5
M7M4umkBMNNgJvg1Rmais0vn50OQQCJD8/3kT7fnqgT0bLiBJBNSy4lgr9SFcQq0HfO5G2ywSjca
jzCvTU7ZjdjY4OmYQARnfsObBtDUV/Z7vR+WUBmMzVpfgyO/X5KHM+KKTKKijxn5WdgwRzcgwM50
jOP7eNT7pa3pba3zivD0Hbi38XKcKKgkNOft7hwJ1ArDrgqDlRorYZcBoFsbf2k3biAt+0A/P+nl
IgmmwY2oZT+lLjCGF9Dpc3iJSe+uhR1L6La0lZ0eHtUcM6TfhXIu5w/hlyhFoJO/ayTH3lLQNyK0
khTiPMjB9ctRZEhnXC/NLUmOoRyG8AHr13C8XZaQE0NukYrklxUVL6njWMKaPps713VXvBzf9Zjs
il7Jx9GRil+3igVBqE8/NZjEc2MfM0lZCM97ssvN2bwEI7JLRgGhA1trwU3MjdYpK4fXvLvztsJ9
P1mF0PO3jJXrTShEu+FIZaNc8k8VO77O9Dspba/37B3ZGaRlLOBAKbdpXmZbKOIKY8EOsHhRTFwX
q/OxHXZj8Nv5nv2cMl7ux4PrK5DNMJVKQHiHKLSlU023meGG5v9/oVb0c8sgVeVR+ePc1TwLlZWA
LVR8TbW8+iRwx2naRX0Lyl72nfxHD0ppfL536/F9CKhkEmqpI2ybwWR8vGWVRT0D5XTfhTS2AbS1
07PLlzfjhIAXm0eSZe0hbn7dLaOe8a1bYy3ujhY4juZcCeTxLMM/fZ7dGa1Msq2RClEAeUlR7Bpo
oPw1Kf72TcyxA+peGD81yax3uqxdqoyET/RxfeLRcinM0P1VBixShldNb+ksx3bzelQSfyOLpujN
L2sgCJW/ZujVJfy+r+qJfgptkARxOimNJjztB+o7L4l+1wpAYsv+DYblb8fdKNeZTVQ2SH2LfJSs
NgdyqTPR8wv5xhnzxSJoYQxoNJvxemhG+8OcBws+0pVIavSHnmziZrZhQ1bWFadeAw7ZqX0A4Nwk
Sbs6YA+JT1Y0PetRxfP1IgN/vB8lOUfc6+MUORf4Ac5RkKWQMZY6TnCi1aMVJ4/nDZPoLooWN8eJ
iMJFXjgyi3wG4ZeAuzfnLYmUlq/QB9lRnzrBRWlxTdIEzpNh+kpgqPK5+vBjj7AB0I9DXgiQiMBC
biDuJeQR1QYR67S8i0QQ/0bZTQfc2lYDBG0deKbx73uEDqGD+xqlJTAUHEsC55Ntk7XTkxpbD5My
OLxWgAa0ECMm6KcedO2W3qC7QTPU6QHfMoc4TT8U2Sk+opgOx5FMsjYKTmmn/tEyLin1xt0tT9vR
JdkG0j4+b6W9J+VHUoceX+JMvNjvJlGAx30cYBIyI9PYXQO4fkmsbkGFvpc9QNiKQUZCgu8Z8lGy
qIZpBFMRYV1IBbwOZBjLEp2pBaH3arlNknoEcviNQamundZ7d3xQLBL2VyRq8dZwD6zvp68HzpzH
uWyNuzwPA7kwPIVWrEelm3Auh5siSPzAoMOIxeYvlGTDdu5g8XxKzFNHSlmLDxqo4ijOpHvSdwu0
n/KaGphVV9j2IAjcx/kgqw6yERAxnsL5c4Xgu8MP/sMbk3gJFyaU/oHR4DihxslngSUb8fIRygsB
/OElH28hlLC/jl+8J7ADpOUUugqK3ugioZ7s0nUW8ZTdD4b2gnBdima80FngYg4mM6+xToWIBudn
4koikA9FFqgDExzdBgt3pbCT7VaAMQ4Vmb3ZWrY4VmF/vhg/0x+ckZpureJz8US6vV06KJzVeL+c
eu2q/+LCTKXT5DwUoYASUUW91Sx0Rl6LmsfEmiiqqmoZwmSU1cMBstXCEz7xmauK15y+J8K7h5Pl
XYE9iKkHBwXvwX4L2yDO+OxD1HORHY0wNvuUijbJ6D1eLVJmIbbtaec5YoUWVWWeQ3mv70s1ZSdj
eWTVJ4eQ+lVj8vUfWgWiJbTXEXcdQlfOpjKzCKWMCDUEiL+n4F6mprTxU6DDNNdUN3T0z/Pn/xJN
RbGA3kCA9Zgzpg/a1WXz5e4phlvp1zzBLeI0jjGyERav80592WHOQVEzDyTO1goGzHa78Hi2tnLX
6UBkQN3JL5+ScqbnF889uMsXYO4jiO7dehJ5hzeX7MxLaeYdLrdiwU1uKA3gCDFnsh1BD5P80dG3
L07Q5+jLBy77brZqugA1i2c1CTdWF1Mdk8m1kmZ+IH8GtN2LYepdjiZIE4ixtOyuFQsx37Q3hhsb
5hEGVSLqOTaLuALnlEwJ3ucOc3d9Z4LLvqM80B1bAnulYmrE+ue4EHjU2ib8H/VaHb1jE6giNaIX
moTc7U41eqE4BFgIPBDDrY5co+2osvEU57uNG4yEtRWDlrvJbQcaBN4I+aFIOBbKZgY13NULPmfU
0w/2z+amYkWeBD9oGtgJ3H1qNNFU08KzAtPYI72M0wocQRCvG+gEEhWQMECHKprv3eDvOqamdwgK
6uuL5PRxv7V91Zsxqo6IE2YvkRqRjaGf33qN/CgXdBahd9lJAiJjGBtiMl2coAci4hLy4j74p4YA
oHDpXjSyG0Hpxyxn1hoqHVAh22gZecKVLLpYfrxwl5XBSwh0ihUCYlWkzs8Db9FpQ/VcIAUvA+HV
pNCFnE9YSvsaxI+Wqkzu/NMhfS2JkEPETJ12vqttjThEaAaKsN+y6JDMlvDaJO/UA3qWgZ2p3nwV
4nndvgBD5QM53KwGAF0FWxVAeA9hfPkUiJk+OnffZFDJL9PuKgYBVKnHuTitGSbpmvr3p2Elwl5c
W3lQAO6fEDeE9Wd4Pg9I1XQ/PqO+UzNw64pym/CTy8j+fl1GyoiR+VGVn4Nd5fhI8K9MbYbKXLYv
iNWDPaUnpIR58QJ7EFmyt+JDxRRUP0q9TANJWIHv2DtpfBURmmjs+MtYoW3V1adSunGaxxS0cbup
vSc8EkwlT02kPVBB2P51HkqqbZo1ts01c7RkOYMbC+JfgBj/+7o3VLasgJgTflh7rot+1zc0Fm+e
L4+rUq5tNm6ozFV2/hSqoNoqyR7klNyFo/ciFx3WrNUvve7+T0wAc/gQ6Wqs9ZYXdzO8YCeSoOU2
N1zeK/xy3cEoUB5wSvOSw2wB/EAqMsk5Ir3cVrbExRbLDI+hOjkTHZ/JrKyJblg3sZL5vmcHfVtJ
IoXa1k1ZgMFbW0p1TZgFK+YwssMri5TtZDhVpQLZbEzaAJyZNW2XGGQs47Mn88psaEzGUwrZM9sO
qlwSaFP1ovdJoRKTa9hNhzzubczrVzxaUmsmJnYHKciO02dIYHf0yi+kwphPj3+IkNeVCUZhglMr
C9GwDtenG8l62FK1cpvjZI7UHHjNgclm1grAogHHEtY2hj1jkVV25v0vlc1K0lj1QRK0Q7UdLO9O
Psb3gSFwX0tbL20yx3/QSDgRFGqDTVqFlmBRlNju08jn9YOd0pW9KCmcOp+uoXz8iD9ihVfYAwri
4fy50pbGe1umhV3jxUmi737Zg7wAT1GX+lJgnAC23JaG1sT8HbaHce/bfCEzXJdY3O+z1XDU0hdr
Vqlv6bIEsoXEWuWk7vr1Haelko1ceVjj1PsO22wHCgIxq5J7oE/09JhYS6sAzRElDVnOk0RIbzZ5
oHrXA3gKDrLY9xTu9PfHfRNAIDdQq86tSt93qNDxFa+Pwl+wtzYsp0ng0VTykjQwhRAtRXgEIgJp
mADPtkGAWzhMTrNSILZ1LzMoECh2rZAhhhzqypwHNnrIuuDmnW4F9ft5icvKhHp9E1Cy3e8zHmcA
r4TzrBJr6jhDk05jlEnMudUjok6Ar8utw6NmJ70gUjgFjYICkQ597R90Y94rpN+s+Aux3aEno2pO
JB4vfVEGAnQqT/6WRVjZ544VshfclrNATceq835epBeQO4h9GGAQwBrVMlkFDfLVudb4owFauCR4
FEYihv+6oH1bDlL9n5gA84GtYHDsl1ZORQ61/icpiki2iA1DHCJjj9sBx/oNe9RNQZHCEnPJ/83B
gkZxZ4MYow4AjBNn2idZwsluC2pQ/oR1ihTnFmE3sjg4fDI9kgRfI4BBb6Sfpjr0SBiALdYnwm9s
A08ZR13ji4VeA+l1jE9HUoES2zv+0PA1avANXlRWoiAP4khsvpuhQ2vVXIYk062Br1GLH37uvn8J
qqKTRvw2xK+xfaRAo4Z+mX9ZPMgYFE22KE4VDwZCRw2Cx93NEzklVHgU/mdfmXzDpzgYPPezVkwh
4qhiB2bl5Jl/AabsGJLm2uKN8BuGhOKLYO9rc9tHxQIQj7shIPLRmhMtTbTjssY7HhAkZkWjE8oT
03vafLvYTgqWBQekhcb2sQNt+QyWmsBIqks8p2iZ1O3NMi2lhgzR1ES1BfLGaCdoA4MAxv2UIWv5
17oesWW9HmMyzCUwc8y1hdR6UNX2vhtebC0V3VTeTvmXyB3jeTfZVUfp6+H80oaUFboCWps+NIr3
TJsW1usEJ5zRln/iER4OKi6HFFfKljDZxYRkuGrEgy0m+3W6qcE5XrxmGhWJydukdGKaI9Ce5DdD
5HJRgcrk7KHlz1Z5M8LsdGwMPn0vVlRhA4f9RboTz4lY2xLVUEb3Owopm9kV3/NsxfHCO3FmDqji
NhOl99Gg3V3BYtQSgo4ae+VxyU0Rw5OCUeP6m+CZXAfIIFF5xlxinNk6e3PYcV7RIhF5q9x+Mawg
UOW3UXWKBAPBXEpok10Xq07w8sbu6edSzLfNliwX4G26b/LyI58Ipsf44QUXrs9lUeOuBv9rNBN7
LYKKALeEMlND9f0rDr5b3ake+PAq+z1mz0SwGzGy7CEC1f1MW/c/bMWCCvra7k4Qq679QXLvymdS
egZTeI2bGQI6uTQDPZMxTxkPWgCIU0HiMGhGqt/RnLw9qa3Htf4e4s6gbrFMX5UyO2yPlZfiwGOV
kPd6RB9S6pOImOBvwKCL78KaigthyzKUeNbEFZcp/0gzCsZmT+WZHmYsiNSQWKPHEQtKmaVX4cYb
2CLTMxSdlWkFSDDObbM3VnF7wryE7h5l7Z3yRUQuAgr8sTJgJnyaoF7/2/U3irEMEo+EwhZVzNT+
Purr+B8PUUPQGIV6/m1OVU05sewEFz6OqK/9bp02cR+St6zFgU/j7uaUmtt1ZOicgdrOoZBpgLv3
rkOFmeYannUd5LXi+SBzw0Y6vXVZPi8hDII4DowDjq2GdqUVxY4nwhUebJV9QwVYzcWX31mMAdVi
3GjceTgE/+wBPop/s4pULCwkM9YJAdH72ot8oSo9+ZzNkzBnGis7/EYgVTOLJxVws6AX0e0MhSN9
FXTkABYaxbiuMaFJsACgZbmqEPzuSkIrwA6AuZ4gwXQQGVfiULsWYc9loX4FEPSGLuaCSTnEA8kQ
Pn216q4Ua8hSRtL225XfcE7mHOdS5Dt4yQexZw+9ko9/jSyR2lUOxb40kGfO13gDmrWjUHG8G06Z
SvMD16CE2RzRsW3BUSQ8rZUj1rr4945Ud4Wlfexh68rvTy9XHiLJMZ+jjrpl+brQunOYUsoLCPU3
mqCS5aWMe4xPSCdxE4/Y7XvTizs0ekgV0lSBR39i6xekXeVxrvVuxcXUV3SbJ9wjqytMFQdU7d7+
5/p3zC8duOnF89OpsxdXNIOHh5QQGD3MMS/0Wzn0lybr+Kqv8HVbixxm4pBLkRyv2cajL4scXvo2
vWvCinsrqtjB2TzHIESbjIGjB2KA243tLZa8vCA5kjezk92EabhiPDDrBHiEu7AYeqHfaA/6Mipp
Lyv1un6W9MmpbXPDrlMIjzFWn+JVTiR9XJ6Bqb7jJKxi7rdMq0WSIoJoRYJo2tZTAc7/pJKMv86k
ahKCktOuvTcLiIO/oRIzdFIsHoCrwuIZh0JTAT2Uo1Lk6Xy7hsm3PcUogAekFu0p/Up6sSkpmf7J
VMVMkuP6XFRwYKEZOGomLvEN0EKwEKMmbOV2DM3lq1iFLbSJfnrPf+3jXwRcy3AoWqU1vhAk9Ry5
BG+Smx5xnv6bBYABJNuxK7q5HDygcLELiZO/TmRVh6E191osGKnbCIkISkuKPPGpxGiwTK9sd819
PR0PS/2H7zVTqH6QIYgj2IKKuNpVm+Kky3kN4bk/ir/S9rhFt5XqZMxVXEMesodc+D2OlkS/1tVC
HLK+Ww5AkemfqBrtK4nD9rNCi9DZnemMPbxy7dbQ+qlDk4vYxWGfVkL82XiI2ScJhkPLf+AdPPSC
R4YgvCqm/lpkGpHQk2ozZMBzuvtgpSTTTuBpfNfH21EPvWaCVGAJdbmrM7am6sAzq6ovqyPRG1Sc
85iiVDwXHTUG6FR7VTFZb3BuKOz2pLV0tNs7l/zvVQHAp3b3+whvg4t3iGqjyT6nYxL0CbvOXMFO
hIk2rrBq/gRYbwkF0kAmHSKkONCgrOIfMFIc/p6rs33WzgmphNDbOZnn+ugx1Ww9AzhVH838M6vk
hOPWZroY6wpfI/izNms0zQZJ+iF6KGE5RzQE4onzwYDWR/OvD4bi3syLATTXfawxhXrRYXYLfOLP
WM2G2mlVzkGaGjUtkMlfUnfmYsnU0/+N44MFY5VKf0+TOKohY62LbUBJujbaOkhiYWfu4R/EGdam
91n5mRqCSpSJdQEDlEjkWjsmoCF+LNxRXxZVSuwlVyzP8tzVRAn6YohXyisQ+6dDKvu/ePDKQa3H
ehyVTMN4yQbA/ZHDrwIox0ub9bsJGYeFuaS8nlDHvGAlLdGKjfuL/4y2Vz3tZuUKpO0oLoptnOlM
XStvQniWvxxDw/NBjZN7nN1l4ftl2rEIocLN3oG7iLEslo1hCScHvMNAG06JGJ5lp3xutJdpBD7p
qA9aIsLv62740KRLYgLvcsm9zrfniamdaazDnC9dvgFWnuWdHGoGTENSRpcOrSPjrYj6lTabnzMG
u08Y88rqJIDvvtUerbUYNrVPaE1xKzIjRRWm2kJwE7VxlPqa35+KVlj6/Kb4r/0kkuwbQ1gH7al4
k+c/I7ZYbVZDlomeF1mQWzaur6lte2jS/ZGIupKm09qXfuPUhz9dAFguaY6eRgN1zuq8czrKbS/2
5SV48CSsyfp0eaVi/vhizI+/q07ESgu/+59GjWglPCzroln7v+xkHAlc0+qh+GktsBBkHpSsjlcJ
up8tOv7NKLzkmTI7JRYaZbq/P1vx89DSTlMVCuFWuMye/RmlAZIq1Kbmw9fpmadK/VcIn0fFDDmE
OaF711gaVQOk3CNItdtzXhm1e8rFDd1aJ9KAhLl9O0yc3MUXchc2x7R269rv2sFWSc9xz0DRJxkj
D2vreYXAXY28Kk2tSK8g7zy0NJFlqJ1zDb6enwfT0dcF0u5fnhT6WKRw06cANizNd6DodJehxRZF
CCECTSfC6PVpi6glJK6ECt98y4forCKJVJggXrVv5p7IepGh/43sLBWc6pYYQUDcOnamKIJmTARj
UljgOrxlgt0R7vTShCw6aAF5ytG/YkbctRcs0iapWcJz+Ag0gBrCH6SYiqvR0Qr43DzebtyGArrK
ZqK1HfL+zbwpd/EKS7h4WDkRoBf4uK35AHiT5TIlTuCYro3WtlGGjjCwzOh0c+b8AMmKVe3yfU58
N64kAjDd/yY9T/OnOfsoMtdJoi4lp0vZvI7BcdwpcYtVpr4LzSzOIOvjsYnYRbk2SzARH3ssLq7r
eqqhyOVMRmcxWoLYfBptwxll/j/quvY9sr8aGHX42rOXopmq2EAej1YkXyJnqvVxCB6lGosmMfEU
BCyWicjMtAyDYBkJrJTh6LbchZhnBxYTHylyBQpM09rifkCIfbSQnBJ2mlpQNwELbISLENpXvRUU
eHw5s3yhGJteKEPpxzqgSZewnpEVVqp9M8LMtQFBFhUI8/bLheX6gBfB6Zlx9MztJNX8SnSKqvFL
mfll1WXhAyV9Qh83TAXQGUcju3A1brjl05B5Faj7emXR/f/atw4P874iCuVyKb9X6aNi1sxTm1e6
ZnREzbOLNWCnshKdaCy03v4D+U0yRoAuocvtoCdbGOBQLjcyVX7ieBX9kCXVsyy+VUpZaPYurc/v
a/ph44WaKevkoK/0oO7dUGqyNr24agwP+7+9BdyG6Bpr6uEROFC9gsJaEA+xghPwpnVcjA0KhQch
J5dAICXgeVja6BKUnFB9232q4hZl3lVhorFwcXtP5qS8+z93vIERGoL7bzpt52gULlxZliDzxGV0
hoyYunQNReAO3JfGkJppMJmTy2y4Zc8RuwUKj9Jzcus1G45vo1Ms/ZDP1baFH0u0CLlpkpIE4a0D
aAUFidFMEgaAzhGgAAtpLdfWX4Jt6+O0GoNt6xM3ePDB98Lru0vBN19kfmCU25i5hUAW6jHtDJi5
czbwDxC1KHdL9drm7MyxfRYHW5U5msUwAVdnfsNNQN6fil47R08y8oBvPBB/Nl6t+M+rvIgetYB8
JGm23Ujnv8owI7E76Jh4QlKDqPabWu58Z18dBKJrIyxTavI3Lz0z3xz8qPd7qM3N49YKeH2S8e2c
WPnP55s0kTfKCtAG3lKL8/Quu4txY2Vv9bj3YovbzTWU5sjcFklgpayw263gmu49sLqEktylQZ2N
axeRx8Q4hksvsl/PcnNaXmg8MLH+qUiZ/0nnT7ZNrrJN2lKQLjceRKgMRVZ3sTMjUkMX4/UzHJ+r
tOEz05wDmpXoSNYdwmYl29U3y/h46Fu5XndN3z2YOYOiCm361bEqJ69cMeVzMmJeABce+k8mpMxJ
67uVB0nrSNZTll5N9WEFwWsPwaY61W66QSaNHx1BaWyL7wrmc+5/R7K8dKKIDZLqvQ04gzpBKDoo
IYO/5D3tTP/TiIp7hGcdEkP9+jy+BPa+Gl51wMBtJAFGUOTJmRtNah+2fT7m5sW7aCVEA9cI5I7R
HSut38FMd72YUABzRnJQGj8Xd0kWDFslHxLQ6VXA/3Zl8zf2bfcdW1V07TLFuAcO0eHY/xQUh+gX
pQc88FuxwJd5AqJm6BX/hGcHY6UAYpqflRYS/IFNZdAlRCT1JbI2MHHEF9cLF1YSRIT63todpCVB
pUg+rrC13n0KtVD7ZccKnRQymrl27uZASlxa3YVwEa43GrWDsmmzPfD0xs/KaycIgxXrXMmOTt8v
RdMlfe811+pjNhzLRvs5ZZ6O6RO3koPmg9cSkWUOe+E28dYR9hD3PS/t09M0N1fM/6XOS0PKZsKX
BHnjpMrqUntHRzwEjtOIDqpNQM8nXA7Fxct7L4RBVlc74EeWHVUrJIxxwdTQWDPu9a+W6K9mOhcD
z+Gl8nAxo+Bn2QHg0zF1h53w6kTUXhym/6ssEyXjiPmRPepGKOnUfWcUo4jXRgR59ACvTQ5OmFI9
akGZVnsEopON1YOIfiFJwPlveSHm0YF5zHUM4PNmM2IlFzUlrFb2kWntXFFStkyoY3lSPjlpMt1R
8rfolhF+mrxyBFfBWwvEopl6sJO6jCYQkH089IX1+1TalsnCd4OtHg3KbguwDjtLOIsFU2dCduHJ
nsO7vSb7Md6qT/L31F/58pLRkHHz4Kn0qkyjXmf6k7qs/NlOBuiaSd86qYPUvhbdy0EBYldX7Bgr
K28Z+sSAwARJl7majQ2KClx7+DTX18HJUiFvvIynOFXWlCfQJOI8lzaH1ZxYSBGmhlcRxNOHIonc
fsdBANVwuNJyc3RshVkJF4d+zT+pCvBqkYLWGTm3GwuJldzy4Dp84CySPaMcUIUtlX87Q2N9dCgD
iok7g799z9o4KpGMr8zv+5/cipob+BtQg+vvg6gOjFmY9p4PEm4Qr/4DxcH70wWziqWGDE68FLjd
3lIBTfLzGpzh5c7u6Fb8923BknoArIkrTpYHmG4C77V9WIUS4t85yKkvUZAL5qI8GeNFXnRJRFkN
A8cOSHBcKG7ZjKNWRFk5EZA1g1VixtbUDLVNkBzFQI4ufuhqe/1rdK3FQGmoSWV34235B7zWbIS6
d2SKx1LigIWFmMxAbUN4kyHIWWBnsCaH/ROmTkAOKN02Oo++KdgR1D64bWCbtgMqxvekvJzxAQ/k
xVdEUHWr6QgHyLs+9zxRUDiJCON8h/iKpreteZj8yufj6Hz3nmPgojKq6zns9DYZGAyjYvUXRUh6
+Fcgb3DD5VDPo1IRL0+RL4PhvhFEX6fnhGmO/9XIaS/vZmhFCaep20R+7hoC4e3SXjzXxpavm9vu
jA/n5O0mQFeGLkwaDNxvlt/4w9O3Z584eht+6YWug7pegazNl6UwgX1EYGq3/C6TumAL5nWeRHAh
9Q5zB3MTKHcyd5eyuGxlfh79vr6yaweE9jXDklehYmfz7FrOn9msFqiMQsJGHM6IkxZLPPm5Fykt
EAQzF97AO3uAH45tP4ic4WTLMnMzQ136oC2CLtYwUKEZ0ZlrSXhnyzTt8XBT5i1bByPmBxKlnujN
vZGDax9xQL6q0QPQUSt13hMlHfyQzWxBJ3wi40SrbXVhjpiQL2y81eVJ9QzUbO0ozoClQLRzi+ef
nICt7ZKyBer0Oc4h2a+vGhp7h2EExiP+4i8mLpMse91LevV9CnhceIadVSSmP5Ey5Q1yrCPStA9w
Jt0PrGtiZm6UBM3OQOTtKliOUafSzJ8yD6e8ZmD9WyyTehOlGEdDexsTpfPHg1b802cGax5RhPMO
yIdougeik4S4vTJVVXF4T1lT5sA6kc1sCgklAHw6tDdQCmCfchbiAFuCtmG5cKblA1spgf4HtLwg
msfGVutiGvYqrt8MoPcqvyuX/yceAxW1enU/alYDQkaBO05YDnHaJofXtyN/mAtXuP/sStHF+vvk
o8HYXt9KPnwn6TJvsntV5m9b6iO+8Ly8njOhUiq9ggUx0bLdn7iuzRSoF+JcEnEHn0nmRrF4oPsd
gTOOkLL/AQtqE+eGvhHbj6Zj+t9PQZk29yEY6KFXtaMl/ZS+rUFGA98WrctKj3SrsZ8F4YfBxgjc
kh1SbsVzO8sbbmXRQM7upfONE0nbvhBrUEWAfmSbR736rav5VbRLCKJnVHiKSKjDOkei6My9sVZ1
/MevH71d+EBcWSscfEt4sB6eZaklxiPwfFSyiMad2nhF5TFpF5oZ//DJGyLo7icR07uD8Ez6F5QP
76EFCQhr1w/WtP+oGyTCyAyayqY10AFITH/4ezGCHQ/FAd+DfpCy/Y5wlQzX84zUtAuBfy3hRDdm
m/vrpNQ3AzuN5h9dIH3r32c8BzQoqt6E+sWH+kMuqKiMmsEAk2mlvDKmQWXZGXQc6C0pB4YTMe0+
7R4yQDDZOqAiNtXJnmTfSQ4OQTbuBPu7bjOdZT8BDNHxz3A3c08CgC8D7qrbb22JUUHyJWE7hSM1
D4STMIyHkKSnmzqx7JSH1ZwI0Yj2H7Lwj81Ov1RMKUf8T6xo3GMysdYTNd0zG8LJGbbBOSkfmebM
TPyb9Mmxh4oF8gmtXpMHwu0+Wr7oV46NGd4N6bze1FJljFVMDAV0b+qYZIt7m98IH3vS+0PMRpjo
dRZsDhc/c9Pt0ye2rI42JF7hWswtUPZ9IoB/nbQs7fqld1yYri0rXf3wcwmrZv7pOmQpeC4lwR03
ozuWub5SmegD7EB6bHndjb++XM2A9ZZ6caBosLar5nxtBfcZa0DzBYUcVpbGgRuxEYcyOAck7GBq
hUrJ1tz++JF2+UmBtUcJs1iarbruQ+sQUW6l8cvcgIOEeaIYVEEYAErhMRgTR729sMPP8NGZqhrp
qlNvKGEMglOz9o+HTxBFRaooEISNW8WZBtv+7NdkmnvhFfwAkrP+7JmUG6VpWkDXNTrgQdAdSlTP
SH0A4+bxHxI7xXpNpZoNSyEwejPJ9pErjxffqHS/5IHiMeSLcIZ2rDN1eJLgypB4xhqmI1HJnXgD
CrOxjA008odT2RB3xNDMJoN44trkYk3IYwe0ygQxf3qXxN7cO7wrv87Rac9puVO0T70R8uLVqSdq
NfQgzCKcKAmG6p76XCo29a1q3xEf/4sr/mvw42S81axy9qLqXXXwnNwDOkFIQx1V3hao5x45Xdcg
xztaTshYeECkkoaz81CcZFezocLs+L7CRxbehWNMXLhTG+A7oeLtGngdhvcAkxWbsUDjiOGm5oiX
E3JEEi0/avT3aZHdCzPO8jW6MZxNOc3VQn0Z5KfPXfC9DHgDsyZrwIEVhNCYN4mbs2L3qsUCSMB2
ao7oVjupjjJGmCBBO0hycyuUS0X+UVd+1ThS1c3m5sorslG/lmBw7ejwnXo01/kExOX9ilYmT1QA
wSczNHxrFkjMjeoUOo1tnheNDDiaQXLAy8QakC4vqDFyPStpYZajTywWuoIW54Dhmi1rLODepRR/
9bVjskoeuS/+NuFrosCYGlq5wFGHvD3STAc0UK5ZRu4zHSZZtb1vlpSdWijZx3kBJ7g9PPiFWFyO
QYpnfh/RFiFsbyoU4WHHe33rRtB5QZhS0ELTLVIsKI0TkkKcEs+FMAeCLg72uFcGFARERy4ExxCx
mpRDFsC3qhimyIKt3p+umvKCkpl0/HQK47MccwhA3c80aAC7xgvzJRShO7vcx8oQykaMQ/VFjGw4
l21zANVUttWL6bOR6jxf0hGgGkW53m0ak0oYjOn/9SKvi9xjNrY99O3wUSHu3p3+yMmRtdEmlRNr
cXeYOJVTz9kdHQtbSAqS1hiobZnWwwPZHvgrdQx+yXWR+qBCnGAktW2eNwcNtXdJgVhbqaxxV9Af
M6ZFzEUhZsZyQleIDI4eL+pxo7TCNtm6pwh522SMOuhwNI4VIR14NU+S2CszVWs4AVo2xHPCK93U
FCjj9+QTF4+imxIeJq3nQmmjn91UVKPNxM71ljgJfSEtWJnMENw9h/AAkRIgXg178+W4wMKY8uW6
axC5f8uXy/lVPT2jmRDuOtzRaFJ8sKd6DurKs6YbZl3+9zuvmbqwQiVzNbGgLMFeISA+yJ8i76Ng
4qZk5UeHkIjLQeOCOX19XCJfwSJ3G6JMMQE3jDpSednqbt4L9pVjIQiGhIjDlzNo0dgWRsiP+RpP
S9qHDLz2MtCrrgTe98ZI+V1fT8MgY9l+Vxj0kGh/8No932cUVrenS+wmRvFQA9VRhsSsj0svOF6e
1Anxe9wgUjA50H8tV/rT7sFif0XRaviQ7jlG9Z4m4ciNpgyz+tvtqLRoI2kHlmkOTEw1iGak2VMp
nQXExZmDkOF8uw91p7yUlXCSOCacIJ+WZt0UmOgs4LOSHZd1zLhuxnz7yDJis7E2cJlgzroV+3nE
daBX6GOA3Dy7+LM59n4EH263L4Hsa2g2kIWd0nDa4n0navexMg6/0eKoCOUqGFr36WhBA/8JOeB0
stFXQyC1a+AvchX0JbnsXDHSwK7jhK/ToYOc0l6mc8VlZrp6qBHZvEgGqac/JItj08w9OWRCtOc3
UIUOr4nIr3e7QdIM6L6fDHypV48ol6b4X5jmdZHtl6J+nWDBmk7+7vqhAwJ/Z5Zd0Uc8Xu/+TfZ/
yaPciIdyMj8Ukt9O/iy2oBb6MmmH3PN9/3azEIce3readdx+C1+fYuuCET6JZdk4IbPvXBxGl1q2
Z4Ua/pRHtyrVheni22cgmchFvqcDJ0uUWNFO8P91NVCp2tNxmd89XReg+nV7jSqg2J6uMczLHYIm
XNtLwJ7GB3PoldET0HQY+YW+epCjHGKdeLlV//TMB5D3nM0R8+aNEqSS735OBQsc5vIHr7TUyT/2
OJl7lgZ1/wDknse8K4pHPjtV4G4K1V93x3xt06Wc0nwOqKZaTcYHtL103rkekFYwYSwfmJgf5CGi
cXq9/yBIwAT6Cosqz+IsW+X2qXaMZm+Mrq3Nk4VoG11IzhmiDgX7lrB0RR5sOkm64qRKRYOX2iGj
sQA0ZLlJ5gvIbnmyocmZ7T7c6PzMp/9Bj7x6RVV3moodqTyDKd5zuIxrXK2ZnZViWnYyj9OAqgAq
M6t7JqayeCWttH3SQEekTNNEi01JwQLoHvsYvIJbxSCRH3OUxZshUmKszQ6jey8ZJO66roQf8dU8
bYUAECg5CRbBEn6BdyclfkmspfbltGTwBygP8V6Lp4QlgMDFAgeE90XyT7dZhsItl/t5g55rjuTY
AMZ1qsLWmOHFg9Ve8O/SrBjybaj9Y8sV2Gn6dM6s4RJvbgArwMJ8Gn0dDmsr2pfiatB76HMmOthb
NGp3R9ROnAQzuCfhjOaXUlcwtpt65fre8nHjoAhKkwJpL8pAm8JSWjW0I889k8u7uRNWflG58ijP
6NZNNjtiQPEh6koZKedjVS4guCI5ACVPXyq4omeh0X1haY7JVRHT9LZWqltYhiz9r60fvdqveXKV
C4kBCbggikphZhhse/MxgWxwcmMjQJ8SHJvDClczbzvYVeXOGecryMht5XzaME8u87ZNu8Oe6e2X
089iLNURGUwHTJB7SSjxPdwhqqTLjIv1KS3mCVPUM2INPZ1XeBkv3fK7+0EIn75jl3XUpyJx6TaW
jnUQGYplHZSJZHDptXSIdQ97kLchZ0Fwc5oa9KZHRMQdgMdKCzmfXZv4dcO2R1eq5z1WvzQoJhkI
kg99RFhkGo4Am0047eXxdaczFBhpFIhrjZl1YS8CI7fLhkDvoxY9X67hoawcn6GVSMjCEkrwKgsw
IegT6BOxRS33Q8d1ByVM0y3xZO7UEcPMby9+tDbprbBSiczN6yV5IRRQl7VFwZgo0QYh6GyBH72L
FcaYWUwz1sXiTbaIpo32mK6ckics0PDf+z2cduXBOM5Zfv6o65LckQ+sJ00i15zfkrB0cSgObhI9
SA0AURK/9hQWlaClrHbwGbLFijiRvITT/AD5mNPcUuGski58tfgDxU91elQdk3huyyq2a9GXIP4I
sOYpGsgQH6EzjaT3qIqHLLb95x2k3Vqnio6rYZLXoeHtMLXREpnhJIOIUkgfcmJuNRcQNo23n57u
YvZd2FOkEDwlvtddwYNrmFM2Jh9GEavFjmj0US0mUZ4dVYS4LOOZZA8rqM15Za9iZ9uAWjSsdj5L
pHJEMlf/rVxZ0E8JCa927EBOkj8gY0akOAGyccm4paY2z6/X5xZi39pScC6I4ZevbfxD3ezQZAb7
1oAbjXJ9seYddcn3oA2rgjcCBWEpsPh9Ab/KDX3AkmksZBmGtVUmK38WxCGWiJ3KPzoKG9nkfAUq
8MPD29rq9V9vauvoKyX9PrmSY5oCo3zaNqpXXKyYlN6ZlFkcZIi+1eGKEJ9QecJ+DDFnod9XtYU3
oVknSmUH1/RwAlQxVi5Rc4PqiGTVJe+I/8rrGOhpqOoAr/Ahw6Zl4hE3gSyUlTE5YbHgZRg6zqQT
yjNxeCBZPSe8A4jfkyfhu7ygl4qXgGZFTA7V0acff3wNRqZfZnyVG3MEhCMjnaBhYLONKcA7rAYA
ODF7lpe6lkxb9nOhftb36K1DR0UDTAmvurY1D9MMf1T/MolCYwubNTTIDwL8j7skOwFuvwobPMCE
CNvuoxWSHIJ5W1D283ZRvTRML5U61zh+o/SyygNc9tdq3us6hB8ZHTUNGptAY9KyKqkGNKtLbUYF
U6Of5YvLqsdxKwA73RgifHjnnw7L299hd1YUOuXwI05Am21cJrFCtbD/d+RGN/ten/XY75+QjZwg
0rAhq586A9loKc5gcdUeNUYO19jOYWG2cgPp79uE3zBGfaD/k1aKz8TntRN1lIttpiFal0JnV5iU
uZoVsSNWtJxzU3+jcO+fKkeBkxD8JsZPEy4jhcsfd5tgFuxNna/m3V9yWWBR/TVHxWNdyDXziJve
oUgT+LYI2410EWBY4zfCQoFcShx9F/58vrHsBGmMW2CguNpHx4Cs5JKYNAnQBbwxh3LKsdEHX2XK
3B4e3mY0xNe2S0TS+OrV9gHjPUfruY348hpbvFjxk7MKMnM01pkDBzT2+L419K9xrsp7+hnsALk6
oTGz+BE0YnpnIlB35uhBY7eFEX+EaR+MBaGE6DRHmXa4jsH40xoXmxof0eMVNfmocCUvXIWIfyVY
sDCxBl+QeCZLEHyKw66x3XHqNbNyGCUqsDB8i0Uw9TPi8cdNmWnGGyIh5Wnd5farOhQTJaqz2QOQ
ka3Ibns7CHUOD/ILyafkMPEHbnbPNIad1YMup09gJ088Oz0UA0FAsrygZLSoYHB8z5kZWpboTHI3
AYHwhooXDFywyzJWuZwsqmixNS73L1vpwETBI96553N4LQPwqrnmZch29aOIwGr0tfTJ2nY4ohJq
SnfgNOZZQwbj5W4w0HxACBaowT6duq9hcSkTMxGh05y0lA4kOzDgF/oHGxBXmsFoyjS5sVVnFT05
GkKRkdjlmQI0B1WR1d0q/MSYS2xi3DpkA5yAEByZ7uvYOO2yn1Tk67xlFK2V+cdpV446ORbXWbOq
NZQvEqQ+jiZkUi5WPsGi9fOEBbMGqQY7yEFzch/JzZOTe38qxmQ3XrrqVmBU4hqMryQPO7QYL/F1
wQu8HTHXeIltqrUhqg4yCP5U9eVAYtrELVZBzdl95CkoiqRqPd2GHSpNkLwSY5E00VVH0lGrneMA
I4mhDhQWh+ASdHjRpqWrC7Eg6+puhGnD5VTjp+lRKg5WGjMHazx9z8UD0GfM3OEN5fGmJH8Wt4/u
8UcyAPG62GH0P7hy9k2FjB1ZyxW3+CAODYrp+k9twc+hs8C/PG3quX6m7/0KnxXJb8AaDAaB0ODB
5mEQ9nbFt25NcXiQZD1FEVBgV4TG2DPAf82UIfD5M8sJfStBwWLPr46at8SE9GpMRFSmgl9jQc9N
OoyXNCFJhKsrMLycmPBaNV5G9Y27KVPqwrVJ1S6sYeOqZQisZWCccM3Qly9kHGRqB2W7S7gF6D6k
6FZovLLAAZGHzEtq85xYqsFp0suaFunp1QbouJ4LHIhYjIPz+YOH9FmZsOlYenb5vUZzLBiorXDF
KuNIeqi04lMR58ve9919xcqP7gYKQ23ziK9C8CJW3k7Uf4WsKnegB+A2F9uaMCVgXHj+6VT2sYuY
UeKJQJMQQKZtup5AWIZeF2g+TOPq7XeWQpvsKGwqHFdSpw1ucJp4GF+IwR8174wQthgVoxcqIjEm
1TP6qwOftyVIcFO7JRV8yvyMTG8hrctpXoakrgfwLQbOqtJEYMh4Q4UelM3lh/WW3sjcRikhaY36
AisRigoYoGgo3ampDfV5kK30COW3/Jykk/Ek2UAAdYTpPN3tAk1nQE/lA8sAZ2ek4TcvG6Aba+0/
hfwuhyuXP1RXgXiO+sHr9PyI8WQAwkkRR0SOduhw+pxNgZGU6LmsN2zKaDHHc3XfYLV4tusThurs
OKpFAtSHce2oUGMsYs+77tNPmw1p+VJSQNC0bdGKV2WUeVC6RiQZgZ8Y2WbcxN20AQtY3hJzUi1F
Q5W7wOcBYLoN3Dn17iZ1C4o14BTubzlY0eZGj8b8veuN3YM6HsbTeKLan7TdwGYTtjUK4CMZsT1H
MXnX4m+kd0AFObAfyYv/1D1VzpJhKVG6JRH1hBvDuHthvpqO09mgEqpLGRtJf2ravqFycm4yz9IV
o+yu6lsZnOS2xXKsYF+BkQwZQi4l/FiH/bo0z6U9OKljKUWQ+6HCUaZpFi8tahYAAgVWBdR10n3D
1YQ6RfkNIrwvpfH7wWQXUawSMKX1il+LTjDhp2sRvza7kOV9TiUQpzwEyZyBvM8VzgWqX3trobuO
m7S0l31jFUHfbeDLF9NFz4fdo0HyR56fh8oL3vxIYQ28WGoPjOvX4vqED3CyMGGgXD/4gNkVtW3P
M3Ba+utzv4tHueg/WNBHSlyPrDotCk1rzja/Bu4pHIKK6feIxWk8uN080uW8wFzSItrcDHmh26VR
1r0cgesfXrkb7NH8pJiC2jR2rnlu51KEJt/g18N13VAxSfF3TdvDHya2vICw6VOwZqMn2oHu3Pd9
Fw0UW61xlPUf2Ra8+dlYdCw9kSNTnig8YH3L0YqsWQpVEzB7lxiYRv9ytmzpBBSnYw6MwFgNHIsb
VENzsOyEnjlleMsQUUjbwKUyDwKCMK0OIiRAXj68puUaVmjlUlenHKd2D/1PUnYasl9d8QkD0FzS
g2fAv8RkL8ww775jDU6VWkv+8c15fW1Wzc1/GRXsYLUhkAOeUwScR0pIRRE5m/jWVjOuLK0Ssljm
6uU6m4cblkYFlPcDM29fqMVCaAooLJgNDNYb3YqKonZXUtddu7uAMTs4La18O0nBwZ3DWM9phGJ0
5Qlr+NzQTV7YUvUkCY7Lf/OhvJEGSRbcQUNrW9vqgyCjmcniCURdHxbjTMw/htCEOCSZ0z3SMqcP
U3T5GO1l9w1qnN9tuIfmTDkDh7KHBXTMhRnuSnJMg4CMt1YZg3+pMvIH4p/+7hHJBOFZIMb3UAeq
JrYH5SDSrv3deHKpVkXMasPgFsgeeS65H7STuswKpRNV4xgrUj/sR6D7DZHOMQ6JIwMUsgR4fn0z
Db23GK9Q20xD+amOdLQQqn3gf5NJuzZdicdDo7seqRy9ZAxlgpIS5Lo+k0ygcWEKS30hgHw9tUbn
POrbRcq4ndRyFdSuhdZh4VPTj5zSiE/wrxRU29kGpX1q3ApCNrE+rqO8NwPYWZwoynQYu0TJ2/RR
rzsCpanmJcX9YGKCHZ1W6xDRbD57mGnSZ0QYEuZ4CeWC+F9DOdiNxYtSwM+anSno2KENP3DZt89L
+1PWhQ5k3Fph+Yyk66uSHlstKLCjEp7QVCjmDS7ocAHQ/HFV+IWtj8fTKnKVPkjSHaZpkFaRed6Q
7YCLpx7gddbapO39/BrHcOXEt3SttoPa986Bl9VuOkCBT58P0QNJ2iRKrhVnQ0K0bsCjBILLh0/R
45krmmgXqQhKCs8IY1p0BVTeyOd0xuzN2eiG0y3zY4hBqiwr3TMdwsjHd9EGJM4ht1+Sld380wEf
NQ7JPzA6ijjDs0ekOn3C/Ik473hvv02Adpat5JGn6DWHmR/sQ0wptpst3rHlTVHOtXk2y0TdLCK5
FcwQuG9MzrsRgZPZKylOOsM4mqPlaYJ7/Ds3//nSdB4iF+sr7NlNejzmJHA5exIdfMjdnlLRM0DI
vw/+TdbRSUh5+fbcdhzWOVwdt4//biKPCXfHIODMAdlRP7fxW66g7WzqzGZd48vBplPlSdwJw4UI
moKg57ACzCZngvZ95FcaBNQxeFNlPPyL5n5Lo8yaU1OjtceXqzU29e5KYdv3X/BIOpPlmCIpIT08
+BZrt2mgk2X50yv55fb4LgYj5APxg6Xr3I/fLQKxgomQ3YphOMaPIPK7z2lI/GRYmnvwErP4YJYq
xh92/qg16BvvZdPcSpGKExDIlIjVaisNN9wt3O8v6i8jPqYNbJ9TaRjHH+fvrZvAXCSMTCQtlS2a
Vc0mU6NhsQLlVvT3uHPnc/vpi7bf5BO7shu2vY/wdMqm4h3UaVtYr+nSMBe8+xYdObeJOryXVJxF
Fh2DYpd9RjFf8wKRNRVBlAdAB4DFs6mpwhA3vOoN7uibm1OMH0CGdlsFNAMa18B7fuXtE06uCplI
tVkcBigXPxgPHsS01a3am2RBbd1hBxB8NkxweQglvUDgp+aKzNEsnrdj93LDwxdX77w+aOa9N18A
9jgvWW8u41fw6T73fV4LbriY4M3wEoKcSfffAfwFYtab/8Dowwc+kEtSIV8XZAPQTVy+QKoym0iP
KgbM5U7mM9DmwV2vWD6CS3leTj26nnHdl8KS0yjA172/kt/rZLoCxXfiiaqt05hP9xdw8rLw1h5b
Zf1px1rFr0EzGahcwFEr+jS/F0vtqAkdzPH4cWARvePyFQKDefwQinM9+yA2tkylOPOyC2dwMd9H
/+NoRi2o/mPFdhy6eqxG0g+tJs1F7tjdlVT3P/4NDCYEKF0M56nMcCfviEqh0g+XtoKZd7dP34im
OKR6mivn1J790Top2CpMKEIXyyLVhQ2FIZpItrvi6rCWC4lpPhWUPAt2uFL0s61W0oB6bErK35hD
8Ku9XE/+MOV8CwxXwJx1SLdnk3UeOehwWT7g1qEjLaqIZ+Svcwy7NgxoV7CqTNs6LBK7GWRITyVj
NJIQboAJbWkv0AuGznxvqvBncezo4PYkszANPeaLAnLWIC9SX4cFit+jmRxKAWKKvjrP6ibeioT+
6vx6rwRlCNzr/8Gc85b7+epeY/Pwx2hsOMkrGGBSn7d5d2kVoU4L3fmYwa4q2/AdZ3i5ci/ldNDI
LxCfENrzRmDpDVgjuYIkx3wgubf0EBModObW/9hY9RI759zSrADK6aX/T6Uxnyvz5zMGxo46T7MN
o1umqWY8fLOV58e7qJRybJ2wJ99sIBUXbZ99jZNJ9pqGIL/idIcqRexSFiEOPi5SrEKAOWL4HkAp
ggjr/pRENT1AFj5s5I3vEIKsYKnWcXP8Xrk3JZ4nWgiZntV1uAQpiRbzaCp39sg+69GPSKgq3sRl
czOKxP4ouZUf19axE5y9H3GEGzr2q03llpeOWdb2/24NeLjZy1BIHN4Tno7KKcWMBH0I722A2NV/
VszRhKG8QfXUm0zocg2BT//rCbm90xSreI+mNxT0/5YfWt+WiKHYN8mOqMUbZ5g1RAfP1IbX/i0P
fj5wIFcGphn6ohQRWaQxq6Mq6Hsj0tZGynvVlIT1gKzhoDtlxq01Mm3TPLSV9RxmquD+hWdyvsbx
QfuGnUroJzjUHTSYOMjbU897iINKGauiLBzBjSfSTYmkFq8IsI+DzNvBFl3dE0Lt/2NkJq5jllnV
gjobfON78J7n8HsA2A7GdFMCz3URi/di1Spf5MQ4Lz3D+8uKyIs3e9wiqib2ahm08vt9Gnxz4BDM
O9zu2ovx4HofvdOABVkZ2eMCMg1pMe0easSEUYXbCjcneLv9Bo9WzM2sZeH2JIJ1xAOUJ5hjH60X
KH2wjpmQ7A+brtkoyOinR4RsSUxWKM3Fp70qoxmsFbyNyaxoPBV3WIG+09/IDpXFDK+vpWPHOUzu
AeZis22zLvt8Bw2tcZs1UVK9iUG/6uCYbWv0wcHV6voamD/Ax8jCsTIgX4E743OXN8lq37CRmv3T
CVxI6lnnO1eNzPDfxNbsXiKWBWKorn+TgylfI8Fu3mryFKNk41HgCrO7o3NZkNIPnDnVdmUMYqnq
JJQL6/oxECgM6BXieQsFVkLNfW8deMdLGRgZpVvH6RGpDowQ4ZxvJercBeLrS6CZZBk87iaPRJ+f
uPWfnbXCAJZLpMgx5R/KDKJkFwB6Hxj6nlkCs9Ouqs9omQ5Ss4D7bLH6mZZBnt7uXBOPjk71r/e9
MLJZAMrdQNRum5foVRhI4MO3X9Ygibc+UDaEFZ5LfIuiRk5YU58+cO9bRu5uFsHpCeCBGvP4dMKX
qg0+rc+fKa3jirUthivJa47LTVjmYo4rbdKDIYAehidqp1xqoKCF/+ts+YxCkR3JTPije4/fNxTm
GkxpFFibWYg3F5AWXdBlAdkfVYw0pf7EgaeuhNFCggvhQk8Jun5LvFDlH5I56gnNakgoqTaVZrzw
nWD6B6OvnalRT5izCVfTyZkuivXP5s2bNRuI0BTkJYE6bo1qkZVgiTHY2mNntCy5BHR94wQ1bt4a
gZdQWjZDu1qTLh3iNO0V/Ma6IExSgvKZKFtuNvmOh0O6xLSCVPJOnzcdo4iVn/cL2IMYhOjfDoqV
fBTehX+N2WEK8k65lgJKMKYYWX41VXm2TJboN48LQ2WMsmaDomBhWp79AQMS/QTT3SO9rWOktFoL
PIPbFa08hJRmmmXh8vs4Bqy7Xpa2gwcOxB4P9mHp7h8YEPxQEoGvytKvkrctj3VosdfqzOBrdQ1H
xCLXDjEirNX2+GWskDPkQCtXK3APbPNBUKPWsTN7+KFO7lNGHY4sSV6SYZRhCW2fBGqQev/Zjszx
StKZqa0ETPlxQYRgXpGlwJ2j+wdaz3yTEpdWGgVzpA7JkRlT0/dIxhUn1BLIGiZvLSeURIIZwwUp
IVgWBwRxYJln1X/gXsuwvb+fNWsD8B9Lx3psIsTOilrTyQXV7NDZf7pARA1gZnyKLExYH6kYG2ui
j4KaneTrORfprM9OeRSwGTOl1CmXM/lCkW2W0e6y9TZPw8+K0BTsoDvY30KjvH+GKQtugE7065V7
XYQa6K93JOdZezjpgN7E1+ajFng1hHhqvXpSbM0aATZF9m8w9OVd6G7QkVP06VdQ7wkWEydyW4Jb
XmUMJKYlGa98P18ZkFRia4tMw4iytYd18Ry462meuGbf2eElxhwp6QmyOu6/pk+qGc5pKgk/fe5x
EeKLUYTrmFRdLqmjmLA2f9N79J7OVb12wjV/xcsUB2w+RaNQUehessr7uvdsyVHtj/1wBj0ZYH2Z
M62ZqEFNQafeRBVuOAifMJ8cJJ965QGwPFFQeME2gVgqrE0VCIKeH2ItwIdMB7VX2AxYcnhhuRnp
iuDk9z3IeGsyfIUKCZXQ1Gsc8uzo1mbbIcd9UZapfLqC/KJKfpQ45bUb6+5o1pbJEMwz7QMTgsKT
oodF6qJcQ8tNdwbGHoxTfaSvO8w1Jws0vuXCN5aRoXs1FHemsLgwOY5mk9bqw0FXWHUf7qZ0HChM
2EEab2raBch7jF0y4OX9Za2x7JTEtbjRk+4n/fUcTUlNDtq8jpb1FUVX/+J7HNPY5iNBCF6Q4Vmo
Yaj+E0ahvuhLSdW9LPHWsahaD+U6zM/zXU6oV9/U8jv2B+5xnI0/DwJj0F1Ejml6LKbdkVbFS4TD
DuB7j8vHrha5dMSvrBNTJbJruaW8OpE2W5nknLbBN/1lpLP1NOD3ggeRnFV9wchUNjJWaXQQW69c
nluY9H/v1E0YR/tVrZw9Z4tkgB5SPHI15cu1x94/ptloS/ZWq8JY70u3O3Do19T9e+TwkqSj/aaL
eEgmYeZTYMpTt3oKmqlPjuk12HS0D+n52xpoW1yBwxtiB1603AqRSS9U5iIJxncmxmMdM81FqX6B
s1orcAukSNaHozUHSh0bkcxfrg/SUxNxQjJ3rrIHJT/pgf11VFAKlRXj5qZxtHIf1nYkH84IUxK+
NTZs49TscGp/hEq9kuqcze/LshoM+bFxy/km7N+zxTKEp7WOO3EXIijwjuCldqyO8hCr11/oZuUg
5Nj6AnWkJCKrQ/iNHzyVibBVYbMEECzRS+OwRQr8G7I+7zFHl3/2MxSI3LxkbAktYTtCMqNb8I2K
XEEiwUKNDCUvnGmVbRniwHeSff736/HtbTqdqlPuxPZUnc3JDbnEaKSkfIebau3lumpZMZsrmRNp
3UyUdmNT4Fn9b3jRKgK0Tt6JD+uY+nH5cuUmYPbioYK7nN44fDs3hv5xRvP6EbNeuDTdwuuLkFPu
r1HU1uFRKh7AZzcdAT1C2tG9hmNDyO9JJMQCrI+oRnshzOBU29VZi3e6bFzjmhlHjpYrXwVZHK1y
jTIWch0y9OXeiRoXv8PKaHmU4OArQkVm1++rTjc+bp25+Y76enpYqEmPTZZgPsdudMJN4YotvsKe
lLFMGhsJHC86qWnoVQtzehFXZh1y5wl0HaCaufJWH8MmiGTjo8oSBdV6YDNo2mELO8W98bAAfv9I
DOquphe3yHYCGRi0qsWqgq77xPVui/Z+ximLEhuzTR6VxwcZV3Pm5BB7NBB5wUpjyZQCXnUaPL9g
H5uo2hIq0IRfj16G3eKOdHtItIE4cRnsYAl0703Ohx0eZ1W1KlnQHNYPjFCiNpeNxjeaMYE1NS4R
925dDlthLio4tNwQs8kL0m5SrZtBFQAXs7gUcpZBEezZf2IW18AoJ4IjLHaXjsF//2D5YK8FJWQN
hehJXXX+IAjr/LtN7VX11v/gEKHWNni6BS3tIVxebBTSiMB/xZ8WXNczmUVF9OUXJbbFHlJQuswk
v7kof/25vvwtAdTHcVrKOQcWp6il4/J7ffEZ+YmzP681CfFpoU1nR8uQTgk6aLFbwQGqi0YtX4Zm
VjOYdYm/yjovkycMZDf/3EwDU6vCCDJGfhXwdI+qe1IzRXvxRxx5y3OpHxqGNtlWBBnWBQEFkVuT
sfW+n/2wenZ75IZPmYuo8+NeKPTmArvDpCOSOYf5cceMC2aIGPBgjlddzKW/V2lg3e8I7sJ3jaM0
8s10hJtxiHhyCRIEydH+ZSUwCNcjjTGKA76JEmrE68srwYUNoPi0Ln5zbkzamJcpYfU2Z90L9JlM
QVKWTczoWQKDviaDfV5ZWclmVLWTvd0e8Jfw0uzaPoJ+VJbc95Fv/ABiTF9CEWByKluGm41HmM1F
wW8dNqn+D6nibNLGx7L22kCKpgwb2J+ihq/S1bBGFIwFv+zEPhV6vnB/TXanUnx2Ite93OV0EYQ7
xHAMP/Xr2qf7jKzESzs0oUc/T24Vl2hCxgyZ04VFLT8TORPTxhKrYr9wKLlK4S99Oni/SYZ26YYA
IhP3+wFveOWwAuB9xb8B4IEW0P6LkqxvQGJu2IosaRgSO0gU5LFYnAt0fcD+65XyUEEhedHOM+xQ
zBiphzo9T/NszUU2qLwToCmjmX4Bf+/GpuDP2XC8squyAM7BZ3dD7xwdUKUFFbKJH3UC7lQyADHW
p0XDTV9t0wPp+Y586AaGdX71cs+x4bpqFIhD4SeVdGVapbZ86KqROjr9FNEErwTXN4b+rqth1D0P
tEzjxeO9JJHxt3s1cAmPbhJ7GcvBg6aWV9jobIM4wff8dsQp5Bi0XDipUj5326ZwSfgbU013y6Hm
1esl3X+1acr0Nt+awbccaUggL3ppwFn4n/KWxePFWvvJOS/CjcUTUq3xNtBJCBSThMKK0fjQeoad
LTe3W0dK7xKjAiUbsrTrBVxZ1u8YJ++0tYf8mM0Ujl8ZBj/v1hobUwnPTFnDipavixrPK4LCdv2G
UFqb/gk29qEIjFTOEfPFJsU5Qh7z0sIsHy3fNH1QHafohLGqUlQ3bucHGU7wcr69OCPj/YEZZpz3
qp2DSCAJ8fxHw720S3cBwNIGyWCCh2bJioUOwHJwjb3syy7B/Ufm4XjIohQsnP+dV5Xu97SN5916
jMoIqeVcKNZRP4rS4MBNtEtADjjtTPa0OR5u5e5MISMkdKzABa3e+JETxPr5vfTb0E+Q9WervvWZ
S71xmEG9ymyhLgqiQq7339ats2lr0uF68yFkvvXpBXigaoUelYy4tLuP+//v1Li+R8zz8fQNkJ46
vXZYHm7E3eApMv2RKF8waTrjYKBd4RElAp+DwFsktrowrdgYwrJL8eeLj+23TGCrSVLYdGdeeeG9
yuAAjtJ+KugiSg78tNMQtExfh4x0NGhvPk703kYe5VdpuBnGI260jvkxcX7ouH6Hg9rJ5I7zEc9y
gaeGJx/IHnu7pfqyHu00HLovSSshlfa0ayMp5bPsolsuJg+dExuj+1dYnwI/AlZF8YgNlpsC2VE1
IEFp74BYDsP8328wNVPadm4d+NfJxu0H/IC4/Z9LAnwunYJ73eVpEWR/XUavAuvGX8NFOybCujJ+
MZX+6OFaBBQqKDdWz9lprSz/wR8ovo34Dm8u37pK4z7LEk1rrPpQfr1fBH9Ftx4cbPajNs7Gf2+f
le20gFVyowjOQvGewxq8a9+ePHoihr/8uaQaxLAkO3OW12R9OoJQaxUrWTwW9be5/V2k3xqHGmX4
833WFEfvxZOqnwnhPedVhc9VeyX2Uls9FL53Ghj0iMt5rGIDHuDda6DOxn/q8NjXWuamfqcPDLAT
RWAhGOQPqh0RXPtzjv6slbYx2LmFm89+NyIi9j8n6pswHuOvbjoKCi33ODouOQCUGmYxueB0VUxN
cVWKWHEaBkDwecz7815Cez1o0Q+B2iAWcCcsG+0Zs7KzC945NfXdzu/UvSzEAQWfNxWv9bmjV5Hf
9LlYguAlXX78sD5efrMgkGFhtE+oNv9MknC+nGdkX18qWoIjomTQHXQ40vj8eUTVBK6sARzZi8Na
FgSrAswX8iecfdIxDGmqqDv3Jd25RL7mlMWxHUww0P17MHuRA65ZPpOxvIAl9wmosBv6E446AbkJ
oNRk0tsiJ7VVByJ8bBr7e8kZi1Yob9aokaYcLQXdtRrI2KlE62GnyRIRRDdmY0SuQfcBqgA6y4Kn
SIqvA0KcNN2P00lwKEBzofTJZPJpVK/z9fW6DGCd3tM578r2MrC+fmZiz/Ge7zkRDdHTmjFnxYGJ
xKKex6guwvp5JeqUcD0kdD7xevw7s2al22m2XS+SrnoNFtCoy6ifZ/pUlbQgzDBgt17SY5gjFpAR
lZ+eAs0lovJz03TrXhYsK0D1/Iv5RUUPW3RZ/qzCcZbvuGqt+ZmodmjHNaKGbu45H1sW/I0EB5lk
5DJVJKjaBD5eRcTxBlMJEiHX2qbEQJvEzE4AWhaArRqAjzMnLALEB3jUBPChhD3935OfWDgj1+S7
RRX3wuWHGo34qiRd0n76h3ODODrskFD3j+nHiexZo7ECltrPGIbGl7tmEwNlhZJSvoOHYHcOzNXj
oos3zjcqDSQiSrw09UTuvw25apYBi/UqN3tOoSE81uliEt7ewrzi1wppv/vgeeYQVQoZSJ5IoEA+
ZLZXNZufRFmMJC2Vk1VNPh0+x7RQQyQV24xZvRab8YZvK+8aELDUWP5Y+H7/mrzn4PtPtDSJH7MG
4UvFQUDUqAmC4qyqSd7RdtZCb80SJq0rhu4ayBSNjWe+6AcCCzkVsIv6qMKeDMXFXwmScYr+VoJv
vsxFSDXyl3WZPI8jMb6LkDeeLucBC+e8qsqDb9gOPEhG2SRU586VhqT8lF4M9yMa9/vUwmQTl1fi
R6xJHL2ulCFosgLrQ35+tEYKBiHhuPcBeteuc/rle46St8+e3//iB0pA/G7A1eG87MHEUQ12DfE3
O4ymfsIMPYbeyklcRVuR75zJ5qrvWQ427xkPHkR9KKqAPpbjUXsHUEJ827iW6+rr8eqTZFmflpKP
D1OjN2P5dTarlVwunfn/R/EaoUomR+P2bISFZu6qAOpQCmVFJ4c25uv6d75UdhYPGdOSL1G1pNjZ
WJNxKBEDx/rwR2Po6VmQs4ER0YrK8yEMT0BawghVHLyMlWHMQfG0cflnIJEFWOpKsz727xfaidbU
uRujISnHLxr/ESgY4YTe1UnBHMf09yuSQSxAfpTSO2dFafiCZpvTZwGRSH+n0TW0NWRe0UfpUUuh
AUhGg05QOr7RLaX5R0Ef6kqOPucA5ehbvucbmLPmugoSBuanzKWoBhADZdwiuohNRYtlVhUL/ni8
R42i5HImH5VjyaFdrO2MbKC8o9rZ362fpP7A2/0N386hoPeFByhh+20y2FULRiGmNwqivuZLp45C
yed4RVSbZLDxU26QyX7cjlD8936c6ULksG+WTxpeUiPfCR1G0LfuB8kLre7+/x8eAXF5dZW8e5Rd
bhOAUqqhKAwJJaVH5flk54Z40E3MZudmWqAVumcGd2t46Oe1Bd+csU6ySQ7XHee6kiZVZ8EQZUQq
2rTZx/eTKJT6BkEq8HQ/DR68d0KGUGnhotPWGYx1nWX/9YpZ947WLYCkw/CGWrsza+NNFhw3fHFc
euadYyI8j3qsYZlzU8Mz6QH7gtGeuavXdn5bbF/WuPJUQjDrNU8hJZKQ6xpaa/aSq1BQ73vB4gxw
ykt+Na5L6lSc4TiAT15OE9f+LPFR4Zw6C7YgW6axgDTTwWAIVxQ4dbwLDctkVjUVhVODjOR+MxN8
ycty2z6jKTtxDySrpSytLFruVzJ5KWQvjY+jXhRizrbaWAxdmuUxsIIy7pCtPCCR+EfFaVm5Rm1Y
Jk9BK4SRU5G+ZwUhisEUq8uDeQzXJ8V2+UWOyNeXbfvNb3XcrgCxxAGTC0yhthh78jPRGvUwniBg
y2N42Es8hAW17tu/7Cdo0Mdy2T3HvhSYOs0+Ee423vzICRlOD20+RK81j4NAyoFBse1iY7L7Ey/D
In36bK71feq6kTu65yw7JSMcRuNpPMzx7zEh0ZXASuIVS7nPj9VOsCbVmJAhYMCL5akE8ryWWUNZ
i08XhQnerdA4CFn/Rv3bVFby8vneE0lHC33TjUT8Sve6X2hqKDpA5wXt3aQ+PWQdC3Fg0+cQVk64
6Ni+od4x3GpssVZcWaErRxPlYHDooIS7ZcC4CekA2+QbbK9R+Bd/3bedJ86GqReTO7kg6e4ZdDhX
GQqiDv7KRCr9lxOWoDH6mb/bNSezAhdYRBrKMCxizhqiGWmb32POwQTiJhOB0+TpNnPapSnSjRxt
kdB44fqj1hsYS3WYL9Ws2gRafUpjLtxaClke6aGfL9fO44P8HW1zi1d+6/iSZ2GgSD2+cgzpTPki
rzCdUUwpTjYfuTd8EVL7VBMq1PdJ6B20Cvbb1CVXZp2JeJxnIF2x9fE4a8BV9qRyz5nf5IR8Dm5z
cgOsk5Hh9SvmrLy7j4Y83+Hae9kPsc0NzNCyuip58c6tb77ua6hFJshupQK5qSEYHwdgW/mk/C41
HzplkYQDdYxudXScfLTcFrqMeuZosYU1FWkLCA4u51nVbJ55oaFgQDmFVAGdmMcc1JmWczc8WX1i
O+8OKdLcKg77LojGFVdjr7vX2Ai6Pn8KrhGufn/kPBn9lNUT8MUCLr8ZJ2h/JbnuGoTOrfrdoMYU
CIjqtIIlVPuqseXgkRZ8W00m7jlnXKNaBxwllbygrPV8YhrvbMFb0ZYXAXE3WZfLAJfMxPUTUVL2
v8OD4zRYJuu9cRJR3bUiaHmRkjZe5TFnFeGnvfDKCUvibEekVtOIevfFijyXtBdRK2VFCA9+ChA0
dEtBq3ruFiAJCqp5JxrQpEc7HurmhzyAyD8JuMRF4/ews1MvzSauO6fXaLpJ2oRCrUlM2ucId9Fn
By/Y9w2sgepxoSV8oDvZodRxXjjAOIP7pLapNR+/3SaeLBRjnXZ9CSf+m5CQtcRAtg6HNrgeVfYt
/vd9LMsRrQO2MZaJhpC9VJ1Tlesnm/BlQuq/QW2o0y1glyDlXygWV4OdO6bwYxtEZQZMSfE8voP/
/bIKVBr/De37OrKTdq8MhQ3M/fsv9gN6BvwFCqFF9k9/mN0tjVXdrxGI3Fv2wuJnRYbO+Cq2IDXe
6Zl1Pg41x641BPJiK8DjLcRGndnB27Dej5fcYrkTihl5tKY+6FNntyiuJPoA2bivBDX5pOh24m97
HEmcKJHfSILyrCtxNnMugPO+A89dAKgM9zC1VlEn/a0PrQ3YxXQFMoBcdZaI8kmbvJZ0CobW+i5s
4wlqD7mhfI2F68RuFqA3ciu/U+Gxw+KMpbhG/uU/MivY3I0G/xCMBBuAtJkX44HC/hBnxuQ+9RrB
scssmDUqJYM90JHIc8bCewVR6dSxIuSFg5opDh4lOlS8HfQMEykoT0PATgHqwsOQzioUieSCoT+N
ZpyyA3cLIAeSKrR8VqnoQIfL4ePfkM4fcFkCXRFVDH3d4TJ74jYB4rGEoqXzbqPq2k5csHctGcED
jP6glCF4HKqHkOZ7xCz7Ug2HdqbuJd2WMyXlFwz2bLWnRA57a3gy5lJH+RR+XrpO4tApTsyFGVlY
/0VuiqRm8MfB8Z5akvdjmyfFC+c1NI0HjGsQtTpRFzJW80OI1MT9nLAcQ93m9hDwQppxZ6keNw/k
7IWVntX/5921iy6vPlQUDGhkN/ptiW0z59k4AdVNXt/fdazZNv7zAZBBNnr7k+PrvJW7Yw3JwfEo
tP9qLrdqSMjZYAw7Z+Rx4yRQgC7O0K/ZBpGnEi07miezGYAkfbk93dF1fvvbcFGtfACtabWbfH6R
B4ZZg9OiaGA0VU1D8C9zNGjvJjyhmN87h6jSzZ8dU50kKRqEjYzCz7ixQe06GQGW9wfxIRSvM6qI
Q7AX2EJV7pJ6yo+R4veityA/KSrojd9G0lzvu/iDylh3UOwKyLGPupnk/ldomlfQTpDlUpMQr6Qv
bWsoLGLcjG6dldeSqViD3fZ1CeAuWg44et7GrFLKVZNBNu2hlvlN43xmIHc4qm5j3Yp6NEn+tO+Y
0RSod3a7q0teQa4cXRE37Ix9UlDxq7r0gnEfGywK3AZA2uae40fEypkfgN3yUHJloZ3LULKAonv2
Rw9iXFx8aD8CNPCFGMfzLUgk704jaBBCsHdBelKwztWjcowMTFgn2pgPEYxGbMhPYMCpoHuyYYZl
Soa5YOeMq1zwdh/MKDwg8uQPJBIOd3Rxrr3/oQUvqf1GX5POs18r2Fq8Zb2FB6Ty+VNLzD8H5AYb
iODA20erLPjRXi4hfMrWf2Z5FprQrSo9qRbfZfak4WvfjRiv/U56u5Hm9dACpt4wCVtHN55j29Eo
/MSXe6r78/qfXj5JwCgre8PNyBa3Ce1DUCwJxNJqvpm+l3hguHr4ZTYCJSmWCjpIkTuHeNhuEPua
S7k7bFjtlnGClgiVHXAXPhwILc38efiIT4VYCvtWwuX+5yphGdibeJpaAImXhH0zFBmwqx4/4wfJ
T7YIEqzD8gSfAX96asHKQ4ywCNpf3McDPBz1BYlhkygwWd2JS0T473AJZvUVLGE/vKpiwfWbPawr
azP5sdMiWsE1lkRA+OcXZS4jKsXcKeHAFz2RI57ct3aqRu5nGPj+6Ix+dtNrpEGkuZopy6fJrBhS
cCF08WpH7tytLs1oxkueC7ZJd/Y/hakE68BL9/Nwn8L2g3ueJAHzY/4NI48LZ3xe/J5ANWgfRbZD
3Uk4uNvaDr0qc29qkPgiUviA0Ov2v9zI2kZKrCjWS0oB1h3IP302MbXdwYudJIEtr6Y+VT6tt/ll
i5V6A1bE0jaxQeUffrmiYY0mGi3I2bXfcjIXjMSc31e+o02d9aZEswBz9otAZiKdeg5yI/qmuF5b
OwVEmn3D6W3OmhfEBkjZIEIYnSoDCCkZjtIpft2t9SjmDKbgBj19S9n27afyL1tINRnw0OdL9gpP
MGVq8u7pw4OKHEuYllrnENxfb21M8Y4EaXW1KVNq6fOGJNfKrbCd/t+bn7GjqyYdm/xRjeaXA6am
NzZFHTuyGZJQ4/0yizjjcVcEbrAuQreyt/TXcY/p8bbocULPoyld2Sc4vT2UYAMLWxcx0dSFtcYS
MPNpr5wVEEW3SHLbob5vo1vYS7pWdVuV4xXuyO2oqbvaeTRkHwj3SuuWRyDYSRMH088r2YXeE5Qx
SYTSzWUyJelulL1/tDxJW6gLR39LaEsP8AsrteRMb/VZ5rl710oiZ55hnaj5RbAa66Itpg+uuPM3
ZewjjFdK0uyVdSEda/GZs08oezflaYMMauQPboasOWZ3a/YQrqlhCpNfPtuxSxXWV59dgchuZlXd
OLp/ulJ/8n+bWl+5R6gAgiOao4tZkKU07blkMqZNdwSkhy5fHgNF/0/Wyvays0HbIkpvZesrT4VJ
WAHL/5lXbEUQNUwOw7tdv1bXLroc3Jr8H7PWLEz2TNzz5SmwDR3x4MHICmX/KwMV1VvSjn16t2hj
JBpBWdHscj4tWS4NO+pEi0BzuxgDaVQEcxBtfQjGAF057AbjyFSrq6eRNU2hnUSdakFTUvRyHi0V
L2aAQsKDF8WB1rzLVmVUROpSNmmianmJer9L/2JH7O8p9VqkZ4g/yAVDGgcB8gVDsLicoRz/ayHg
x2dHQdaMm7DY3TPEYIRPOxr8hTuuco+dQpX0moYY4qxlvRmfKWpICBpW14VwDIRmZaUa4y4HaXZo
GW0wlq5EP/QuLX0xBL6BNbETLvhq49wWLN4NXvozB/ICtLJO0/friRwlFBPwNxyhylmmTIxFhVxk
pss5Zb1ihMOTaUrI8HywagT9yZjFcALsqdlz/AvSZSoXa5Xr3KRwbvaXL7kdhCNvy6PtoD3NiDUz
NFTP1sHy8Wcvuo3KcqVZIh6rgxaXpdnds2CnVWVYo9WzcQHz3idNWpDMy+w9UyanK2hMQUK/0cF1
VGwSDFy36titKPhSpcSPpDAcpeDF2xdrh/I2mFJTc0pJKF85mVWPv/KRDD2V+OatF6K+IT7cbZ4S
Vwq3b4+a0b21AvrdMqSx4UBcPJgeW8dCdERI+t3de8LKn4uiuo8bdnsbi2f0AcwXKLnaMP6ZRUuN
yxf8JdKwSvdFyh/kxFKUNRgq2SwxgOvKrmNlbBsTqks96w/nMZwfPbtwDRLjs8xL58UfXcZ1qRrJ
2uzpe/Dc16uWLemE9gx2UitwVwA8g90WoBcz44pPnpPuqc1sXW6Yd7Q9b5lEkOxWEyxicUNSBO6c
m4ZDU4IupK/FpOi5OFDklpF2zxVbuvIXDWKUQ0yJ1H3glbO4Sd+H6GMa+n0chiEpWb1zIGn1zSKG
7wsV7DXC7ifDu+Cv6V1vMi7poFDRT/dD0MyN0rTPLk82JWjklC9ypFw4yNAODduOytoB4mSR7zOR
DDLva5QQOk1wVmLpz+uk9igH7DH1hsW+JZrVTbc27WkFmcRdu9wRp02aYNC/YxDI12OoVIvcoN4z
hp9hQX5X+iOah0gMQHjoJyUnKef+CLhp073k++ahxJwhYxzoc0UScnLFIWm7mCplky+0jOhpXLTs
TOtiQUfVEJLNL6RPkDVax7SI19l9OVINB+7Nt2DDXXr8G2zDWTOBm4Veo3/daJyjPbmzlSRGmQKZ
+s5hVlevelUzS/bAPAZXi3oJqKGwrzYJMQr/1ydY1Ws4cQS3NY2NneynDxw+XeH1xwCJIAIQ2Tdl
/QvFo0QF3STPlDRjgy17Ero/CfP5cCThflkQek5uDK3CpwFx0iUhvU7PzxJN55FsECzHJS65XRD4
spFkOggXDq29Yn/cgnkgxh3pSTnBddmGEOxqxmBEiy58ldGbjMN5JRs8+2nIk8nADFZQEWpArJ7e
eFwWpK3qDZPkhND4ZUE9l5yGAyOCcCGYRV9G4fN0/CLggmIKvc/K5sReAnQoTbli9oW3niga2i2m
a7eBZIB5An5MLgHOiiSRJThKsHxLJ8uLY9a3VdxlS+XVjj1UHcj+QyqxoeVNhtktl8jMdherV2p5
x1DzCjAnoGgulmvV0/BUwF8cm36ao5PnH2QfbMLcVhtvjW0krCDZOhqyYD7go0JB0SwFBQZnVYty
sQiKx29gYRodidmnkKQ5wcEydf8Ili0OQFZB+hqIe9mLlwOxvcFujS/yHfum82KXT33fxANix1Bb
6q3YU46IZaSoMAr7ik1W1nxnAtH4Bk+94QOZuvL+y1SDyZfk6nS63cA49IqiDNvJXbZLgVBJwFwk
ZvjsKxhDCSz50XVeft25nBX6DOzB+N3Jn+CDl9ekYVmQu6eSmYLHXkIGf4vjBiXDM6VvtYnC/l2H
e0cKZOYfyuJE9NGZEo6+24KDzclFUWZe5PrR7paP9OegT7lpfMiVwrNMTpLgh0hnoyW/1imZ4KdO
ZYuH/fJzeONjvnj6LBITDcgdbGKtKUlS2TyIXt6cSrr24u1sMFswyeFmrKNX1dhWYVNruzEVy/cJ
TZ6m4JCdDTbHY8/A1GpNeTnJLwmVxOyBEfywbMDMVo6uEZ1GLOIrpC2XmPgO/d8kh27tX0vfJPgQ
Go6B3cWhp9CjUXp0yThN85YZ1TvJIiy0QJOAX8U8m1WFrZZhgpo1N8s86Xjk/niCUGZtbU9hzlKm
PWh5bHvT3UKGiVcKCY9a2EGBPa5WZQvRBAFkrJ45guDIi5pei7QCwBGK2hb0m7WIUeg1CWfulKPx
/xcfwfR9QihbOfv7rNNB2uZKMxidWa7bAbGV9LvkrjHByNpw3EBqmTFokMm3WWecVPYjXOU9pscF
bjgJeudCx/vO+I/6B17tUG/fB9TkGIu2w0OkNatvlNQJDjYlURBpX3VaYgLYizxJFhqyaWJBaYcL
W115zJWmkdunSOwiRPdxibeTYIiaHyiSmPHR6Qb2Mr2k13FtYPXLN4Dy+qv6tm6WZOpB69clIn+W
4zmp2rol4oq9PCWOmudvpuiPrw6Aw7vUcxmseFwmPxUXdoiQlLmCXZkZeJqYBl8xUWg/AcQg/AQQ
pnauWaTNtkR8FJElsqwmn7hlQPu/6ALizlSysourWuygVck/Hi30lZP8wExtAEfFknDw+e/aJhl3
YuSpl52LuR0WPNfXzOCKxGF4dFksi8mppqaNM9H6HO98+6gQnxKmi/HPHckc94NK7Bcduh/yI8Dr
E0Jg5zmuH+H73EImYChMzA62FAgoh62kXA9TRQNFohVw9I0muicERQHCrXJGLYZOpOM8NlpR5sLP
4vb/s5dhI2WlVyI565Jiyc3oKc+kvb35n/PcRIrjn/zITRbVzSQwP1HcB+MKtngF9uLg6Ia6GMiL
YAZy/Quy/cp7wSguI4FtBsENFpmp+ymgRQZp1UY7HI4c6ei7QlYJdcBvocfsmhq2WmvCQPmSBTco
JebRb6PA4gofXdFT1AEZA0vKmANyhVdlWe8GI/ObJySvJv7qcnHyrQcxa1w7NaM0ztqL2FO1qqrq
z8noc2cjH6lfDfLsJUJLjjeIYICuc2xZAgGnfeD1+chINJiWXrFINKKS1OzbJYhRR5Z6QXMc1Adg
FM+k3DJoNa2K0vJubVDus5ypQ2gly+NghuMykHkF27y7y5tFKo5nvUeVfSWH/cC5rJET8whqjoTz
qxK6w1yt3Qt+TKB1EPkwcKsbHiWSGsC9M1xXhNq2J9fxKilQPVqupRPFIXTWdaIndOFdfXit24r+
SQfgHUvz4NSlqrnmGu8v2VhTIlfMZgHrTd5GwE7bbSh6azNNDBWsOb0ZPRUekUJQsUayx9SXsbxk
hqojXNB8FiyqFpzZ2k1qfc7tp7elSY4v0YFBBIURCtXJGN74HsyGDngzN8Ca5IdKYE2kx1Vc3cLA
10aiJOianszYGNyk2//j69nf0eFt1umZ+7UPB9+v1HpHKNRs9LZm0AfrnqgUa+JE6uVaSHEbHLoC
Cu2qcnIilRnv9tE3szoWt9K/AOpjYhXwNGmr9NmxeRwypH7MHvJ/9xz+3EMqyOPFo0L4MGatrcJQ
vFuAmcKcQ7zes6JkDdE0s/Epez1B1bbKBj2ULR8C825u2LW1n9UhhsUZ94VVGcfrhHG/pYc+RwEu
LqDJ3TqtR4/3W46oo1UUveYvn5rvznH0BJLtMHF0fNJG7cHpeZlldP9iMzr6L/BaWqdGICVBlr0p
KStL/H0BwZUm2Xw0Hloni0MpSlzBdHtaAp1ffhMMRNryflV0Olp1o0GYYiqR+b7/p07RlcwB1zJK
aNAzltvCASdvpJTnCEfam6rxJvyH7HSrnMxQpw09b6xWXyNvcSymcF+u62U/vInoCtdxtIYCs2l2
nCSSuIIc0SsO0eP47rCd3oaELFumVj6dxfy5XjE1BYSPWcnJyAU7Hpaes9i8ap22CDkii1eTHBA5
JzCYI4waDgO5NFcvFkuM/d4Q2VGfMuW51hIcL21/V/sJ5IFC4+H9pGE/NHI957J+ky3bkPpR+DNn
5N5Rx7idqS539oFXwvzYWvq0kePAdHtW+hIXtILhOda9svAOxhyt/9ZvHlb9FBzlauA3gt7XcNJ8
Gak+S1vRfYqbqChHTHxe9d+9oPhFiJFiCMZcHXBEV44MeOviQsJogiSRtyEvcOH0HT9tcpLL5B7u
w0ks/waLo5Ow/KzoMXySh7xR/V7lgyeubiHRbkVqJ+avanh3CZF56jwjlsev6COkcRPN7dhiirzG
tr3j+maZa+rLRxB/lrY7Dk+OMODTeY+nEjUPrXcOg/0541T7XsfBeDGWZA7kjFZKNbKqwmkVv9Gg
hGK28V6321AlxDJexwXd4NZQQirJQe8Fq3F86SgkvUe61F+feViDAZvcwZo1sCmDusl8FXnatspJ
v0LU85/DKVbyJ/9mTWGIxWiW3QzRDoYx4gpcM2lZ+XWuabFCPc4XLzJNJ0FpZgA15ga28Tq8A2Dg
qqSr5rLbtrpFhURPVL388A4om/EX2YsNLHITKVtFf4M8VEYI1DQhDoi9JWZGOCjS/A558M/6GNOb
qrUH7ePu8QYUPdbD07jvHQsrJrihcN+ghZ5LMf+GwIkiOgETPnuvDqpHeUEnixyWRpmeQMXleGLr
JS/5uVZQlC+zpoAiDOiemPfhWyESwKFGVnewm3DKpTt33YEVYfscHKr0Ss7rGNDTgdancnD72Gst
pzE7rJUrECnHxK3vHkww4CX+3wGbTfn8ib0eYz1fApi9PQbvZw0uFpl38Wl/j5V2gAiOargwRwnz
aC2EF9W4ccIaoWNaFrFlTHR0BaYPfskmwHiO6AGwjR6H4hx9eZe/i6xSoCAvEgGDovT5URPyybZf
8lo51txB8KyPbG+vCcMAT1o3eIZ4oJlP14rinxfd8bgF0nVXX+7iK9GlxnxHlzTSd6RG0I/YEVdj
XaxhDKoTkjq/24a5votbaQAVuquKeZmI5pQWEKybJ1lezKtMg17DIch1ikSH0GoOxIFfzbzTbyo3
SiOpwilQ0d8zFPBO59UoKX4SJ5c06/r5i0Zm16r3IZ8oQes8XO1Fisxoyg2CBEUeVg1Z3TerMUno
L0lqReiG9H0kWCDMewJDPtUtrcf617TCOWOZuWTlUOvg+4Y9+iH9S14ZlSM2ZGVu4EFpDS4wlgn6
IH7ZR8AUSwRyFU+zOkODlc43/2yzUWhNQBm8NqKo4I4P1i548B08dprlm1iI7n2NpbkWlcqGPNMk
J2JEloJs+4cpSnsiOZsGVAL7zaaunq1GPzE/4FdoObBx51DdjAh10LBQ4SxCNdtpYXPpqvJMpMXi
u7aPh+Xw5uO5cNm74lZ7NiPzlmBboh6w979OsSV2SGvmILc9x3KzvEilClqdgPMxPVqzZjD1zUaZ
tBHim4cYJEWQP+hq3IDwekO6p6xqL3Y4ogxNBk4eeloCT7uz4rHjyoYTNjoCAJqYl21fMwSb/gmd
Iis5pni+rUVm1fd7aiOsTK/l3Nboe2pwg+lESaEpVhi2AfX9w9vzyGS4CFimVXr9jzBNN6Hrklyg
1Jwx97w5vtA08oHS00neC9fomUHOPr+djcFw5s5czmkPDmG7VHKCkIkQlXdaSujqV2dQV7G68Ma8
TlFKASfYH6e3m9aQCdibYtMFtiuCqzNux63sbHvYvQ4119dY8jJEIDqDiKYM8OJ2beGuo1upPS4z
678mpkn53t+VImXLJCz0FtMclpAIoxS01SzEzKE6KODOtWfOq0J/SgknA66aV7GnTtlTxNknKeJu
dTHxWs51/YEjEF7sKEnrvUEVSK6CCibRdeK8dp+cp7Je03JC3HCNG+FTO2fQo6PnRMt7+Jm93eav
sqxtJm418L7ijoiyN0kOqmzNO3Y0kw6BniIDmXGTjgviWdhoYavYEXrkptCZNt7x0ivpULjOPkIv
aDieIHgUbFW3IVJX+6LbIwqdMWSoJrp+wxTiFjYLW7WF/lANiZzW50OwIrnb5pgyYxdG/0LLRfz3
XWJ+DzL2Dodxx5SrCpPfTiH02kzsPZQl4yk5/dWxG7I9WeH6SMYiMtRVSAxfw3QyZ1IALEjumyYT
YUao0L9Zy3lZahxrXeYNFd8oFUU/WTJ9h/0liaZsTisssHgjGfPdPmaZ02B0iAxrbT+OtckCmQOH
QV4j4RwvvO5QERdapKtNTA1r0I61l5rY5sOYuIK4oy914AVGc5RO2LGtFCs6UuOWjHmtNvT1WUBL
g3llBeoRd04jCa7uNtMYHaf9L+WAoe73FaZXc8YYUvYPOLGkmYNkNyTwHZSRxHJ82NDBA6rgXPnC
7aG2Kup+KG7LJPgYX00CY5NUqxiT4VqW9DDdSDGcXB1UP7HYAm4F/2m6/pSJk7qfGsHboPFPNlKR
U1rGqaxV5y4JeWo/MWxMQ5knyKXOy0sL3avxdzN3kzKfRAGtn1JNAxJ43bGvT1lmBdY/aEjSSHT3
ODC0IDmXqinemhhkR0BgkDiQU+P3s3DXDvSf5uYJwM6+WsuRFTz+LjGzQ6ueC76yo4AJKeSGYCD5
ZZG8XjlStATgfhw6dtR010pmkka9hvZJEbAMaoveZDrOhNMO6w7Grq4C9Ri0s9R0whY8ZEFUv+wJ
6T8JSgLGeoWdF2zTz54a5UkhDzrLet3a9MRyEaO1k0xuuAIvDkRZKvZMWAFK/Jx9epFO11DURhiw
y9QlVn+XwAqF8yWVFZeesXY1xl7LFw4PeTcZ2t5ekWnJ1iZs3X5RPubkJY2JO3VJkKVFv9W1nDrO
A2LGjX7SuQimDO1o3WQwykojpsZpxw4QFxV4yhTOagiW6kB28xuLSU76Az9q2Se4y4rD6ZxXfwLf
Pf+uRpHTXB6OZaZMBwIiz1KT+giuN0Ie8ca3NvdLp+mPxXfxZ8wFwlLg4NkOZIhXm/ZuCHytOULB
q7DOVcIbuNvBqMgbAT3Ed1XaesG+Uc2xA2ga6NZ17P9L6w4RMMUIVpFPykiHbfeqPHfSbFfTJNwG
P6Hxyuu6jyanaGjMQKYKeMx00m//lzZrlNDvSyluuEYfo1+7EzUV/rDFvG+sLEq4VLp8PJo1qIuq
WfL+VCP7XFl6fru9QZvLhMdpzXtRkCVfq21eMqiFVIrMxSuyfcOV2GTcETsXQHwKDQ+c7JjTgbJ2
KZAnsyveievUp09veGTsCxGPIwC7wicLH/7l8oAyRbk9YuW1OPPRCb35Ba7KV7laCKs/HiejMeWI
fPGknHeY3ENn/UVk5MgyizKCR2cbFYAow9lE7VS4T8wTQEEtYAoE8wrWA3J8mBZNL9m794jxig/9
3gFf+7ngU/rsvLC/fwwtCD8m9bUQXfueWelHPLZv+kNwtgfHIIJBC305hqEwRCEmLh9eV7E6EXmT
QnM13becu929ySdZ3a9Pz9iclwKGOOsiIY4EWMXcmLxRDHkR2ZrkrQ2iy+KU2UHLrlf+zQwgo7SD
mhto1l9+JRMYSP2/IzXf8B+9g9E/mAQRkbRu6Auq5H66VFb0+O87QDm4+erMKAmFMJ+fArqvvPay
hVxIhN7gAILwRSErZ5hhoYbDCWLZAlSiCuK2SO4dBeiTYfF66tSQcGjaDP89bDdqHr8J4w4HPzpm
qP8Cc/nKo2e9clxxQGZNJPVc6Z9ceLqJv8gJ7i7jtbw4opkP+DzYlJQtW0Ie2oDhoLsJHkN0s6Xf
kIyZ91ayqVVL3UMHWAvEpQ/Zq4ovTuZkrh/lCKAP2WLnBduE+HcbL1FssldK+thJrtXbbrAoby6F
d/MtijoyhT73rUnwLSAxS3Y5jzLTl2kga9SEH8ArUCTKtW4D7qWPBg+i7q/Uw9CazU6DVrAsuse5
CKJB7NSca21tN8HPsvz2JDoqLwbx1RXTlWD2SSq9Lf1nsdykT5jpwa446MJiwa0FxARybdmi6GWO
GIioNJaDYm0kyXHQDPPjMIh2N8qw3Zfw16ANtbGr5VwW8Hmnf+RDYgMIp7iISY3uInUItUC6sihH
7E0k0ei0+6XQPrSORolHQA8VHSvqXBoNHZVHVFg44Sqec3qxdhs5i+tkjsKV1gMs43HIVUK8Vbg2
uGkfjo7rt5z7T7zzD9FarO5zkN6T8PXYPvm/WYTWgGjO4I5eHUrS427a4XkKQdQEToh927Uxz9P9
wiBMk6tQ2+DM8mjWIw7/RWrifT1MOYLJinsijm5TZjXNxxIL36/BWBUs6zedfREJIeU624XGjTYP
OSndwouO0JfjlVJjF3Op0BR6KdaDIakyQ63lZb77XEWzhYh5tUJ9gOMypPeWPVY/UD188C4t8TaJ
OvpeEzL90Gsh9FfzImF+hciCTgRuR4LfoyQtm9C/CB94wxroabru8R/H9NqEy3/j2fxko1whyI0J
IhF3LmWjscx4t4f47eNxwmL2im12dsqXkPwHeENE8sutJYWIX/0d8rwlsx8q39Z7+ZcrNOf2kZjz
lOTLdPxiI5vYcXSk0Zp+Lku9IGeR5c8MREiURJpggu/G2PLasolkueyxZqtaGw9+fyXqfbXRokr8
p0PNGKi7bdFEbLSrEw5+3tlI4z8Dn5LHXmZYXuXmpTi6rtnmRBoPGb6K1mbhlS9z5GPmudb5MRe0
kyAaWv9JFfyNBtbgpSMXaYzkKovFtdJ4yPPVioq7f68WNfix78iTOPOKc96Km0tWIZZqexHaBg8b
4KrpeXMlge/9JOtkBchItkX5R0aH7K0PfTStwl6bWahd1xlJsSnOeV6C3eRAXgXKXqO6Mocspbl8
5ldg9oeqIiJ2zodA542qM8H1U8JbWWAGnoQRQ7Z4U0If1DgSKy9SO/aBoC8OxCeUWr2gac8dCFui
v2VuAy+3HCmGTGOOX/xdHWBZlsZukyekbt/rYj2HjpJGcsbQQ+wRXOuyXfaGvPOIdil8KWTwPaJZ
fDdipNAP3aTAOEUm8QFkLKM8qOcF1m+Clmgm8lAJBMXjmZf6KNuJJpUxc1WnvMHPCMUnG2Ptja6Y
o6/ZRglEyYX+fDuxwCN5GemwNu5NEi6J72QKxhFBXG1iQeCRbwggMAUXHv/VhUvtsEQXBAI8jJMO
xCoHmxzyqtD1Ijp6FJwjYkFac03gtRzpOE+6pxjRBNFPtpOwBuVHitshTYXtKjykCfFSy/V3poc3
bV1tEio3POXA/PCwEI0Mxoq622O6eGKAkLeU2EjvwTn6JchxQcSWECyN+fGfEDbXn3MZxUjLHI3O
tlPuc/xnn0ozTnIjWiMG3ujh8Sicte8pR3Tr+fD4MoptgBc8toTbkfUyPP8O6FXyamdRATcHwUmx
cGZByRBzJLR5D8Q3T8Z8t8b7hw/9muKpi4dDDZDZnu7raTNKjP9q+MdKbH5pQvAO6aDpwNTSq2s1
Vii97j5fximNegMsdCNyi1EGnwLLbjJwGBZK7WXBYhp5Y3UwdDyvcw1IP3AiPl/HunrHM0Ybewc3
VtlDPqVDlkqIDfh68RK4D3Womyu9puZxo6m+RW/Kfeqt9fac7T+bcNwVsyDm2frj0epQuezecbE4
44y44kuIqWUnQoge1DTpNX80Xi0mdyAiOFTraIC2UMBuY5lMKdqejXBLYU89DFWy/LQpGUlK0J2Y
q9S/9T1QSif5L7Sm7xq8oLSpF90k1QOtlGvDh0AzS6x6OLdiTu4speD84q21E93iCtG8Ulm8wlgF
ZQ8uuCYY0GorkWm0FqlS7siPqm/H8XxJAxOclW1MqEPleRSVIJ0uOT3ebGJ5pDHY5+eTrOti+FAf
4P0Q++p8sOtJprPCfoQmYAxHyiiTVsksiq1bs/Xqrrv3tWx/ySFtUdr6+mGn3988j6J8QqZLAF1d
nagamJBhqyijQklYXKTZPZ1JeHZWaYjrnSI6UiUb1pmew1ozNxj8kawgCEXvOE9koGB/3YcKcfll
GiaNfIWLPWDh7YGohQVNPMZVNJA49kMG9zYWVDU6Idz1P9J7YJcmLF3nDX4vFqat0p3ttX6Ld8QF
xd+i4LmWwly6QIp14VL9bJb2o5vY1Pssh3xprj86+fanm11cSKnWkgTpLI8EKQDIok8zv7OFOcxa
1NosesRR62dU3Vf+psu0uow3Bhw3c9MHlegPZ16ex8W6ayRINy7fMoVcqrhxVZd93w3bFIufOvrN
V4yZJGwSryuhCY6Yg2kOQEeuQQYthUeRz9TIkSjSuzNx+nNNGNDb6SCKRqU5IuZPfPAZvbpWYpzn
EMrlshVAg67631K9gCzJtta/Y0fx58dlzI2rSUmKkqGrNwbG/ceA0bx97gor0yplH725/VFMBox+
r91UPe3l/5pgQvpjMfs0Es6E7K0GnVKc7suA2Cun8wF8qjZ1cxLKQaLxGpsFLXfeu99+SXwax+tU
Le7hmLcv3l5N9jU9d38O6nH4s5xFs2nEzecWrkUg0UMNdGvAfIE8anmYD8G642xQtUau2RV0VTgt
ht07x08teJzg6lMFXAV+7ktKP/S9RiqGrBkW+9WqDGvpU1VFP+9FEGeuBYUrsVQ+4iCgAanBdLK8
YnEZ/7VxmZcIMqBkESl4XN6MFeX41Lsnkb/GNGz8cNVq+m1eV2nOPqeMmF05glUgqyTnI9GBjGrk
Yu9igtISHEeorj3BOkJ9Z3a4tq+u1XtaFZL9Zwa5se27xzIGVxJANkdX07aCeuPP0YxumKdOSNdK
RWOtsiyRtUKTZqU1baKln8yhHbXRkijkIeYTPcByOmF+5kVpkH5OMPPKEn8k7M/k1PGI5QSPW+GY
PyVingmdpjSD/h3Jn/hWeiT3dlvrQ7kGBd5XV/QI7qGHyh8JT36OzF9CJzQhJV+pD0iIOTPikn+D
kMCYOHFG2+Hy0grU5eiWFEtFlGJQq5V3aPJJosSn3Jpm1o0qka04xj6LM8TFGgWq9dqbobOy73HK
s7mDY4UFlpdR4QlkSMLxhizrhJ3jAQcEXkBrpw7HnTtEEBX4Ajj9oRwLowGs5OFVZ9lgQir31dYx
jZYf+AmU/XlMaz+cFUbRVhHf+Z2ApqSRpbmoFZcMTu8LuXdV9ZrK1XXeOpKAJi1BKz0T958WKtEj
lsjtmnKR3vjxCcpslJvG+l0ajBLHWLbTZy9KnetYx5wV9EaPKwYmSFc/Ddb6SEUCnw9C1uex5oHH
qf499BiR006HSWw71jD5py7wsJ7oGDzlLunhEAl/vW1Rc5BitipNtE+iVTM3XXepwtHKHgNcrq0n
RhYxV2ZYJNbS/C6ooRp7oxDWt+wGluVrDwtoyItEIrf0EMoQsXjgevxxD6M8uUx6Re9m8Kh7Hfih
4bKxsuIRec3ZJTNhl/e04/qNr/b8X0T3D9V0qFjDNKm7MOIjc+uiah5ch1UGNl/m/it14kxSP6an
llzhhqbUEssLJO9NYOkRXWkwGwdVFzMigHXhlOrqdjWWscEYYnFjUl+z60AKp2+y+bSnB6ZGH0RP
dc439v86hpHwIvDzm3myZOP9N39A1UZCVMNWkZQjvseZnnUp7MtkRyG/EWVIpJTzhpvWURra0p6J
H3epnxYKXGocWoJ6c8kdKJpSLt6iVlhQhgVd5Uqx6vJx1ohqpj2Cf2x+DTGSrK4BjlJyKn0kvy3R
j7uddfoVbvXX0NjV150mSBiJFxv7G5LzHYwOoafKRRXJSFkKl7PCN6+n6/zI4jooQuizvLF0TiOw
KnkB+Pt2I383lkqyMWrZ8aYGMbOE6rV0dllxgOeNDqgDrOeA3OIdPupAVx45WyMfEBxy1dmCtszQ
oWNwJ57GFtQTtFTzzFT3ERJ8pEpoOsF9Fi7cvn/Ia4pccL0luG+zFREp+HNCgAlzMl+GAe2+4jde
9C+KA9gwAItWjVTFqBxGo4ps6b2qjFtTolh2BrkLlZ25IgPkGHTGwjqL4fXP1N9sqaqn2li0Q1lX
xTvih69RXNNEouqHvftYCtJWvkfXwGkngFmHxBCaKoClcRL3rrzTMrrs73zvqnNpvuDo1nKe2cOF
soEsf0WfOIK2QQI5ng8GDlUHFm6Ow2qBGD0Y69sJIA+7lnwOr4nIMlUuNWxrK3f+KKfjy5dQGTP8
VawlTZSA8xOjqJdaqpoQq+P+Ahc+CIH2ayFA7f65Bjsaja1jp/TkQBt9XtBMKgS1WW8RqBpGIoiw
zBT5JvxoWgJbpDSjYgwQrPfj6HhwKKZGmjLgQeWcaYLXd2AcVsxvxes3lfAr/nKQQfwfxdzpbsfN
Lh8vrBF5JMjUI3CfR0VDaFzjBJv3kk3t8eHzDYHQEmbdE8DHFsPQy3dL0mcV06akXi/FhFfjHec5
nB0XGJXAjuwLdss7lVzvD4ZKvHNNVroAuCp+xz2tahQxH0NN8kZmsJhQXGnDwvR9NqXn0EYC8oss
M25mrlT94NRishKvwaNBOwrqhChtC2LwqcHO29/S03GuicWnbnnG+KzF548p8028V9+8Zace6X6F
pKpjdSNpfFRBGYnLxbcp84Ai6JEF8HRJk+zMm13oqlNWnELVsykA/I7NpjH5HhB7quezOMA/U8OU
fgzZTTECEz6sUPPP+/OKw8A8qqQk4Gre0E85pwwNwd1WpjamKck/GZRi4hcHXt+K92LoJpZIJzVM
rC2zbxVBTqXrMvKVHOHijioenavrZkR5ZyT54NXLgqYrEKUC7QhV8YAghh7b8BsIXPjYzGynhgDH
z9yjJzWMuw56SISfcT4uzEMpH0b4rmlXj6QoAFQpH+MP2JCWtSltIbtUEIo2snDCaAaY8S/rjDmB
dNKWeXHCy2j2CHAaC/PdUV6vkoUiLvWH0bR675eV80UjmTSzio1lou174VeIsWelgwStZqbcopF0
klNjAdzR4q5Zt1xPiUp05/OSk2xMNA8Kn6ps+LKawSficx/yxjZTNUlBd0L+WvhspDFINu6OaHxm
JD91qzK12AAx5+ulyC7Iiy6zIugz2cANdxdpXlDOcguFxlxAuibo09w2yXYZLG5yAfenRJ/Zz3Si
FK7fDprR5K/31CzyUmSjIVK6n8AqH2yUwvJz55eTgD3cxXAs1LKFTsDKEmvvfwlGOBEsvh5AAs0h
/Zy0abMfeq4/9I1KM71fzBdLOpJaKDfquS2S3ilk6MmAMyXb7Qtr2PsAiMYnDM2GWTr7sR8MPiT+
LcM40TKN6q7r4pYvqauU9c2d5hPNmMbO4X2kyqC60CkClZJ0I4q6wBDRmwbZqiUTLxeB3hR7M6zu
O1spV0Bjzk/dv2mU6ZQqHvAuAd1pUt/rSNKTMw0ltifpDFR5Vf98AI2UGjDx7KBl5Q3ONrh5nQm5
zUinskxfNkWzBa6AoNIfDFGNF1qVam1zDwdbb+0QKbeO6seaxb0FR4P8EXFwsPY8PWv96zD1RH0t
TCz701P3cBvmAOuv5ghfRAghZiJjIyTC+Tnafq0mgpC23w/QEUukaPVUPLDhp7puaX0AoEMGqOPQ
MRAxgSuMe9hZSwvJQ6WCnmCsvzLHos6gtjJj8tMZgyCLu+Y2ZnFd9Oi7QmeTDuKK6yTxHhK+U36d
rJkQF3thx4g+87GP3rirrp6hCHzaZTeIuzItMaALI6j3qg2YpP1HD9hk39rvLRS/+Ev83aUKUPOm
05mMOiGECsGGXe5h4TNSlFxLVfCRWrHpLqXlV0T/cZ0ujSkRq02CqeEAmy60vie/WuPk+pUgHkJj
XM0xkhQDxoX7Kq24CTex44ozPnUt0+uPsjklv9WKkB6x3TGRX6V0b4bo9Aff71AiBCMp6cAkqleC
CLrEboLksywz2vGtwect64S78Q7yBk/uQPNuQpzHILHGQSJ0IRvDgSzibmTMVdl8JkBKs2cAVJz3
vDXd0S92N7TeliV0/74P+korap5SkSrXvQ5nwmiRI0evdNHr2zaO6UtmZevKvTGFsA/KOdBdln5I
JZ58XT9lKA7Dn8AYJj/ZTabfT2FXb4VquS+14BDcZQ544DBFxIguZK/gEvcmmPqYujPe5gmEdn6O
T2Twp1qg7MojMsJSOYKqRiQgfCqqObKbw1mga3mD330rVmbClOZPUI2o/XKCr8nORAwZQo1HYpYL
rGOR/2wrwqF75OoHAR7a++ujnYUsBrCihlWkm2GlploTrE+euofOfGtu8YGXyw0yt81Isy68Dj42
fs3Gjjd2fVlKt/miF+yRmd89DYkYd2doSMONKgX1p01igR90GpKe57uyLtUgBnWiBz/VW9iHZP5Y
vk5Q+4CjbY3KNkImagW066vESXQIMvEkyRlHAJud8pPwxaYB9ZYR3b3yi3hHGs6Ps1VEAD+0M9gt
EGYzqbgLk4pNWhxw2Po9zrjWHOEtLfLQmgg9eAqpmns0NyfWhxZjU59x+jv+81x7J9xmq7Byre69
1wvgv44h7/yYo5VkAg1LUYHwOl2oZmgkqjZ2hfZDIm1P9Me8ChWgzhxtraYuyW72aqJ64ybpXK3k
wv6K6/8bWPI4pkup+I055fHF8N1pN1fpWagL1+oR6/eBFZ0xXG3otmY0kH/5bQfkWIVM6Z3bCYcK
L8mp3p4SAlBnWoh7QbM8zwhqTjH7KhHzPM+nOB8fW8L6dqjW0m2ccUlBNUL2d8ptumT2GiE+rw1C
LDnnJZl9oYxu3Uyou64XsjUmHTGRewJPmY5v9TvaOMGY32cJKENc2KLFAfWD/7m4LGMcY2G+g7pI
yVedkglB0kUPPmBiEHO+liiJAYFPDstXqtYQaEaVRvbo2Y7NiaH46tmP45Wd+ZamayMv4vdcwK0I
98xpbft/tWaI8LKthfaULFGTk2lSQgVuh5lQyZ8frT+SQ2P4OwJeFKTfYBQ0vLqJA1sr3ndgV0Lo
xAlh569jzgsPh52WqAB6X5vXlb8VkabRGjLvcJwY4eMzHgIqHMROhJoio24M4yPHr5y0mLas6uWT
Oe1omH6xaUi21xxOBSwTr0g3KhFT+ywMlJMPEByP59psVjAt0frmbAvslSX7y7MVeKR7Sp5cei9Y
8VaBCT9+MWSliFmOGmX27T+VqA5UfSamV7sT0vgVTZ6DNS6XJTe6nhDGz1n5LeINxvr9+XIpFN+M
6GVQiFZRVHn9BBrzMH/33on5apzIiBXgRe/ywV26RZhhdHNknmEXUZusTJmAA4i5IfLvWO+vRECB
QAZk9wGPzCOzIUD7mOY47/9iGgfU5ffdUHnWXuQHl29XAVLrMRc8N9qArb1p4++TZF1mAAAACqRX
kumPIM+PVSGKO0opbF0ulkxKQOgq9UzlrOq/nR1h/51M8mWjdQtbsaoxby+to75cE+4jAlOrylhi
RY8g+yatBnCWmQiYo4VmfORDaz7YQSTmpBjqTucvQCzSITZmwqOboMN+/i3v30yBPSi/WBh3S2bq
t76pHsuWrf88Hg0rc7Phcz53wVTqpdQRTjLt0Qua3NQ8JNaR+uvk2EmDHZCE9foJUOUgPHnAQOHI
hVB03thCYFwO2UlRFFi2Qawhvo00X/PnYwFzemadx4clfkkSvuIVPTGV/QH5+4TYUeIm9W20FP5L
mlSOXKeYo3DAokwix6zFBQp2yDYAQ13cGUZeq4Q87w1BEcfBFnfjHCQNpBQiygZTP8edT2NOoRrw
wyxBx6cTkD+CfnpwyNuJWR0NzbfvRsOY6CQtTTikzEwhmkfvhceFd+b0m/0bxyIFGnckSXBIdKEs
klV/WWSO7FN8F6OGGXMS/JQF9cOlTsJSR4R1Fp6kOkImBFbMkVZjUNQomEBIC/1v0gyR/r+PZglI
kIfVwO+Y0v55RRExEOGPva8N8gl8EHYo01EgR4rYWHixA+hoJ/X0WyMjQVY7QQLCX6JM7xpNSGLT
erlOQRV++z+8y+f+1jhqF5HMbCbLhNbcjR+LFBWYhiwnZUEdhbiCz8Wc3TypQhAze8+aK/OsVMKu
wWANLAc4cPu379njE+XBxE8Iu6kQhq5Ziczz8L3JbHjyqBJ6yAhZ0dfQ3Eu7U9iJ90F1Me9q5tzz
Wf/CTNLfzh7q/Szaf3Pd7bdPuECIygN4xID3P0likjdoh6S5Ju7+662zgJ0t5qAsYc+8qQbGYjU2
Npp0m9H1JnmYjF/yYBmvQtcT2OJMrW9m0VjZ4+j0svNPAdQ3J4i94Cbzslz0NZhqVZRSEnwM1P87
defMhQTGFHXyLztaW/ukTmOgTpd9QPPc0LjiImdQy9txge38Ix+hSB2bGpKDhK4EnjKRT8y5f2jd
wfRlLFaTwzZ1g4BAs6taQPbItdvf6chBVPzhWEXmROrmuHVyJ5tIN8zYf12IfDztoOTiOYiEPGUI
WuqpneQRFAHHixlXDIVWC/dTn/kl8sidPsUN2OCtnoAfw/yIUcJi3dy+m9YSr4j9zzijiCMxVnng
kAFINhxtfRpp3RR3/aPHC/F/HbCpmS69iziXAnbguYMHlJOaluG8XNVtStpRHzx1W72iw0luROyt
5+3yQBpK3kROY/6KI5IkxGB7Rl4IIxPAkv0tu/j67GaBYaI6zJWy/Wq5ZTpDeHPgPn/CwItdKMkh
6kCCpNJuldZGjNojVpWnq8xrs0ehazALEwr0sNN5gjGItoHNaRjgZCvNHTw2/bEiial56MIuZNIs
rTBv/Dcc6b9S+d1TYFNc90Xs6UR3Gk1Q3yPikfh79z58ZnN8BR2L07nJeyl863oTHWjh4koHBrzN
rqEXpUoCRsFNxILaReoXTKaJzCKxJJi/NBkiuAoY6HHNeKGEux7+IBNEEsTEVrJP3f87DyK3kxqa
Sh8BWajbt+UA2sqYm3HpDeRbo5ZAZm8cVB+3uY+35/ogN8nlD+7kU9VqwF/DHQWj4Tikg2GAPajI
1m3AQoZCu8PEu7MTwdxCYz5w68UV4dfevSuo71PgCu6w1RwRT5rLZD1JQ6wb0EgEh6UZerymmG+M
M8DJXs3JG9hhrNUHg4cWdmK9scG9QYOpkTsiCHl0Cmtvx518S/zYaMqA0pDGpRcMTy2uK4jp2gbK
oAf3+scNEAC1QS1QOME5BrNli7Vc8skQACyGT1D2d12PpU6KFvKhBp8Ben19ehOmVE6+9IcG+XRB
sQt9LwqC+HivvINiwva1QOh4mcgo/H+v5xhq72BYOjdHT70BoBJCynzgen0fIRacP7OwhCF3dJg7
RPjXsjIKEveSGqhUvDSozN59k+UVPt2YTBq1GPQAiw5YeNj11kCuJ3cNCZ6JQszFpxxF0E4oJMCO
LpF06NSQsNAMNG124+v8o6ztnxZAjVtDx4XUwc2vUWQ8A9QF39N0l81bULvRefJDQ1GeqLLhxpBB
SzJ4Bt6H987TbnsbW5mPXa+/AeUhlDB3wM+vsEvbx8XFOAs9IbF253XQofsOyo1efHnoCYAkvz4o
e6rfCsuqb2guN3BizpxoEsSKD0im8E44uRUYTuzDODN4dItc3JYEW0JeZGEtg9dzERfgE9plNb/o
p0K3iLYwukUKc6NvH3qF1+KuhUyIFEPFmC/nQa+nmBupObM7Ecy3ETpe65y+qQp0IwIm6EVPNwew
BCqaIhsn+zNqYH32mnB46wc3HDUh7VSTHmbGsLs4AUQ6DFkWRFJqo1j739uPhdEDgaO0cR14lVNw
Fg/yr5iXWvAscU3lti2aZpAhthPQkhB+RT5+YOl75Tyh6KZuEN+JsMduphBC2GHolTD2jzvm9NPI
ZWg1wlVZnjiUmSsdnetzqQDXwhn1/U2yO5f8dYJKloIQEhZU7ADI5EgEeypLsXFuwPG5DxJI39h+
2CpvehmMN52w3KPLwdnbsPLvKQMgn0M/zMgoqdbrvuyQlQvS9EZm3QLf0OS5xlLjxiLT7n78mcbX
hFBT9L3GdhSWyPP1M5BTAqBSpoAXpoFG4HWLfUa+ngfjPXkgDqbYIqlGsSWpjO6XMHDBxw/9MCp+
6Q8JY9/zoC6rdV8vlJ++xJ9ABCaSXs3+g3BqJ5KFHBgey937KjWPaQ7Pfm+p3/PNt5wzjCN2surk
KTEAWxPTe6jZ2FP/n/DNlrn79++L5BUGdYVde9LyIZ9VXEmizVrcCpd51lBV3ziD4T+GA/+sOQrZ
gDItHkyiX5XE8j90O0WmiD776kXmOz74s77Enk4YmKwR4udcWGPEJdjQ97NPkIci3mVfR4iIgSU+
dU4/JmVL4aMzGSmqBxPiNBzhhk+dHCCpqJ/huy2YCeopz3yRErv/fJ61C8BF2hSiVAgu/PtP7b2J
cFTf6784pd4mEetEeCY/wi5qCYGlT9NQorvtSwhexhB3Kxp2H9LiIl1yH1bBvM+yKq2atcMLtfr2
MtYCoZocIhtchuVj9cDfe08rkfCUyQdHhjDAVTvq2Nbotk6Isfvd/CIWV05kn+L0TR+hc3uMXP+w
v6DpFrHbaNe5YH0+M/t4DgUiMXPzeUV1yLZWE8yvS089bfsg825egHDUit8UAtXehwkAmCP7JrQ0
W99/fn1rq4OmnDOIQMYfvnST9md4s5xI1z7t/WCtme8x2rYtxuMZZGv/enIVk1wkMZHHZ6PFSeLP
mmyfzjFfSLJFJSb+Ea7PpyEL6FCMAuC/ihqn9bxpWCYsSEp18IKZBB91vhHUfV75MJZ9Mb4/x6Ln
uUj5VYYHnisoqMYhAZFzfgl4t8Bx/LsmVAiQR7ItwzBiziPECy+A79t1X3dU4k1HkKpjOh3qcF91
KEtQ+UA2gartxNTXuleZPtxFFoPj0yAnvXxhLYLuNPtzKZUOrkILzvYd5mTBBPOL+CceqXOog1Yc
VAtyZfHKee8l/OOzoXXw45UkheRaxO3tMqBaylzi7drxKJq3TeBRxfYcXAfaFq1ffXuxPx0HRhvk
HO8imu3sGqEaGP5/i5FgYb5r9ke1Nz+v2gmdTscrp/nWND7SuBxgAuuV58XAZdjlr0lsdATXZdQ7
8BQQ8z/TkQxHNhelOhU0KLk3nBf6BfqbkpQa3GTFCJmlDDG/+LCdHLyRnvBIjfYrmDuRuWHy2u8W
7qi8T/TEUZ3YbAYg8pntujstVN312HQ8WhnWgKngeRgAAGxe72XDR1H3Zyb5J36aauaZA5FyeCEp
5ucVMRkt8Sckd/UUlJv4SUXcvOoeERe0W9szQDjMWR8bubvyTAExtNViymtm0AGi+eNpEErWgaE3
caIPILnVOHw4q+zluAwWBn7kMsoYg5Lt5VwqhgtlYvW4X3vUloAuRNPz/YuSIoRn3YT6ALCYQEi2
RSzIzk2H4uiuxI4QzKDTGYMd23iCb7xGBceVv/r4X1/kY9oKLrDMINUbIXSjyNWLSatWWN8d5IfX
LllMBlGZIdGgp58DRhHV2KJ8r1irkL/lJasY2OLvAd2r6OC8Bg5JKzq9UMqW5mWTIPDn1mdPOYw2
wVgmQ0uI6nkhICGrWsMJfVyefYEBrfjokXZbK0aZpaTghBiASia/L340GuE0Ku4YJf6FKleAQXHH
toDDsJ0H/YahX84xlZdngE9eFkCIzX4AxACiAKz+czTK5fcK38iJLWFxUthZ4B1BDbqbncmSYci2
YvHVe9UQi8C1JDXN9zCAQ1KaNmQ3jwKEMShOWEoo3t9Y38dHxCbwjcjcCH5E/RJdVa8nIAaLDtoW
1hxR/vpvqLp+YyD7u6qLM5u9vNDGa1aVMIBWlvpwulLViNvkQhhiFE6j1sdSB/qVAdkcxsXx9BTb
FvGSUN8JpAP/6pSdFeL7sBwV6V/ETa4dsD6leT6nHtIRVCXYMBgQV89LuDditBQ0uiRKTb0VPaRV
nBc4TSSST705aQWxGR2tGTaMWoje0CQMXJSYGzMIoH1XSVthQ9BfK3AiIi0hq2brTcKJ43WCVFOE
/kBwHOMDNv7LTJxdHOfV52UvZRhiTRmTBdnpePwPyvY/CV2ccpxwTmkaWIBJOp9EFVvkC8Qwd090
j1NXF8Cud8y5yF/EAK9v9PT7e5+zronXhlxJM8VqG3asGRIaZWSOvOK2rLPChHY5N0biBjI+vzBh
YFHQc1BHmTuQjcML8LuobQZT8SmSFdLsr0S1KAlHRcAwI91VmtmeohcKcgyUJvH/ooi04rECzkTy
LkLsToZWnCmidVFmrN3lCax4jZmkz1UQp0SpVzZ5y9afNMLP0RIwDvyiX8U68ZbOW2mvzspnYUqM
oG87DaooIQQJoOb1Ryk9jQdHlKVmxMVjb7cGJCLhz8jK+r5/GlhCnd3NBPLPOdX87UF/fQnJD8c2
UmabQ/mqfOb3KoZakVcQZR1P/skiA9AFc8vh16H0RUm+UPAE7Vj9XhqK4MoyH0KMDd1D8k151Z4t
1t1eI2knW4ljLnEEOcIctwR/X0Ppoo+vw9fHWL+q7Ex1+QrrOn55wvGsQLOC3ZW19E3ZabatMGQt
8ZIGXtSsAUh1LgGS1N/CsK6rhi0RNUX5i3G1gi2mXgqeBwH5om9w56aPCDvU6qjItZs1jgG11iDq
taMUl9zq2QFvhwuCE4RFKBM49Iy58nQDsb3st+MigYncMo4ceUJL9bYiZ8d9AkJwR/iyvCqVJjhK
+Qs+EpgORUFsCHBhzTetkNGJZ9Bi+520anUvWaWb2psZ6M9ZvJLbO3jY9fsnl9fBmrDipO6ymOIH
1FTQkEWOVwOIotQX01/r2Gr8Jpu0DpI7fwFHFoBaAguRa8i4aqkQQzsXirfpF5vESWWUTfm8AEVq
3LIrGCbLXodCmIux6gVn4j2C4/nPEgOpR8qKs0PlAAAQA6n4swyz4uRQZzvpvuGk8HbvkSiyCoVX
khHtTGszkqfK8YeA+1kA8i1DQCbG9vKQCxzPX1bmcUYmf+H3yWHZlx4+Vmtn9FtHnx11fzCtpeBo
TV2FLB9H9VXvpf66bw2gZOFE0Q1QplcbyMQTsYUZ0n8x056BH8KzlhaLTnYeA0iUKvlGpp28hQQ+
oGOgSmi8E1BAFtQ2/l6mEKIIgrVPLRAJ6iDdrC1wiPM6Q3UMPTMwwCVl86p9uG8KfmmXy44BIHC+
sEqq4ZZUCJuMaCax/2TmvXwzmb+6cTGvpwa0sBw7EoEm68iWfGa9uYpkEBWaXVyTlf0bKtfmL1k0
UCtd7EdEQnGOIoXrE8FZ3Etc0tN2tba782LtZ0U9SjAIPM/8YnVf5S/IFZjBXBPTJ6gsqawmxsW6
L/0zLMIc0kPN9LWsdzKQaeqllC5oeadfw/B85SwpD0vPAEIA775/5HxTO8UI1+dOBs+7lqYDGlRQ
qbmb94dw3orOzE/svv0kx3yrxVHlwOQCTt0v+iUGeWPENt3VRwxdrcOJ2ButABVEWJzKau9bldCL
nS9cjfo4WWRi/nglb9ms8cxQMhz8HccOY/bHln8AWalxbpPnNWF0nzz6RbHB1Zz21ua+aK077bTk
X9S9LofT+wITmr8NnE3I3RpEW7PUtSoPP+hC2QN9zsoyHSTtce9D2e+8o+BZ3rnu4wMAyFSXvQ5u
jXWKWa8I1Q5GeaNo8WXQQL3CIGjPUpvh1om3jS1Vbjh09a8nAYW0JsoJ6UHa4yaeUvNHPsIT7NFd
URhHxtQ53EiN6iprtFTjHF/Y2ymtY+uwSx4hK1kOeqqsuzh75cBiMAoTbnItZVSBozD90pj5Mjze
vbClhXNqWcEqtwzlKpuQYtHDwMtmDQVqSeEc6tAeMM++TWGPDb7p1EEa7pPOQ2pwZ3ErK7zCOqSJ
G7xuO5WGXfAsn9k1ZYaEhb6FW0Ru1ndpufXEIo5KP1O3BFlyGHAiToz10HzxaQsC45xzesANcYeh
NrUUb92iKfPsNBd8TSJkGAKqJ5/wJ2Rc1hxJzozAeeZKShYNvUdmmZcb07uEFfwc90I9s4XxjHNo
wwJZytnNO6bIvAVIAjAvn6teFDDZK85Wkgjiujr1Q9PdUCtIW+u1nC8N3V9kQk2+8uXuzxdE3rRL
OcVf1TAurguJddk8harLmeotyT6Ks5senTx/VLKtAJUw64AVPQX80MmvhYtYvVU/iRi26E8bUF2B
Ga7NddAxDU7j6whI3nMqx0LmpdjGKMtnRl/8v8BsiWOdLH6DnBIJodkvoG1j5o6GU9Y9DFMPEo3D
hirDaQoEJir05I9PnzFdhAuSxkfVyhYWV7ImpdIj5dPCC/p4gUwh8Wjb4h5PRZGFK6Fpb01qBCvX
1VWXHWfOQTYWH0r3fNMFyqAILcmXBEvmQ28VrroFGsx1eP5nIfEIn40n59skkzXhB6txN5tQQ7Au
VNKmTHFJ5IpDCOpB8CdKJkpxOq5tscWicZpFhrBWdDKqYuQS2YpGTHDvmnfd1614A+Be8Dn+rZ+L
/toEaHKZ+zDwadabvaX+R7brBmIWg3OMNCDeyu0pMXeNHGBceOBHWbAgAKijReaCw5eRHNPGEwTG
XttdKF2L78otMnam4MhBAjYohH++y46WLusZsxmkBaHxuru3P2XQbzX4KFDrT56ndpGN5smzGreI
bsC+IoYAIZQD4krcJTrB4vsU6qd8ZYsnqxr3nef6MbElAIf5A9xnNCQakpB+IBEh1WLDsoCOIc+M
5UUISjkT0LA6AqnaPekF62ohJH1FUc5QlTk0eWjq7xG2P9jf6ihLTuHqykVsEi9vsfKcGl+NZ+ao
UwjSgrCmEVTJAPmrMoi/xlQRYvF/5Kc5cPjKU88JCmD2cKH9HIMGspzKAvgNOQZre0kloO1tqcRr
rxulSP4FHFJEH5dd1tTRtRb0ncwb1WIzpueL4u26IS7NjEBU72OuxQjvEM4n9P9Ywrf7WqXHu0GF
tKics1pc87blR/K6AXyWZTkOOvQ1kBMNy9MwRMdQb1E+3E3B2rd4H+9/9W17hFvtUYwhrq/CjDOI
dFSwbVHJeLIFx+qyEZ08MMPpl1nd+BKGNSVBMWFkPYtvb4MKa039S1qgoDVWtuHv3YIdnPvK8ACt
K2y4I+8+vnYtgoB+zZj9FacEgLLnSEXMxvCHfi4wHiAg7Z9K5vs1mm7ssK0je0GeXOzdTjfqsMpW
ddUqgoyflDbCY5GLzhnntD4tXV4YXljm64Y8ClqPf0o3TJ15zCO/XbtMDGSFa8fWS8G635P0JPlV
wSGhlt5cvNRl01mDMFdGSMi4GFG4f016qks+iRhjaRZXAgCJ3p6BOX8Q9/Ijk7aU9w6T/PzvPfN9
bujXZ82FYUpUczCu3A9XFcMoknsQz3oqYsgeuzgfw2yxEs5DoQvuMtrPgz98nJfPEESayjjRrpmy
hyNU3cUtqEx9ROAX1JqF3wutQirXVLW7EMlcT07oISM339tyBy7ptmCmB+gAZ4cBYX146+0wcq1T
yHNu7gordsqXwoqAgCDNbr/Ft0Ztrmn77NXsxHRoAruhxUPm8B+IpfH2/Zx0XEqprCra1S9UXeW0
nQs3NXEGO94SUn+4O5UVdsq+ux1VFBAFuPuvvCtdkdvysdOJb3d5/x2gtO2kwYZjauP0LJnAqiGP
dAm5V5pKb38vm3z8IvCt3hUSUuqaOjODcejZaLy38IDiAPlcSu+YA0RJ2x8kejQpC4btR0E2Skno
kSCbGbRT6X3otHyU2mb5x9E7gseOdbxdgO7jvvmFmSZ0COARJuc6WNuHWwz6nM7TFOnpep7ZXXFB
V/tDYzrBZ5u62DAtKjEpzW6JFLfhI+pTb+C3zoPi1x32ElpryjaAIuDbV+TjY6ZX3309bN+cNHIf
ow0j7iGjIJEahNwBtwcp3GnWa+1XMRuE0+d+340/hLX3oHjZMGKupV0BzhH5GIjUwnxWvZvmaMzD
TEjtXSXk6XMfz79gOU76oBnRzgxqYbOlOarTQRIeNbQQenNgrhvYZwKI1WNveL73j+EFKTMRvoAI
pBC15oCeEDFDmSL3LqfzVe2xFYnNCgJaIVP5GdNisQqBcZhecXKQYGGeQfMPpP/66UCMQj2ytdj1
/h/1u+TbSv6BkGXAMcgv8PHyCMoQVnzvAkplZFr8tkOXgMpzpuQzTVweryVKMOi24mQwqU+KuRsW
1LDpeQzv1uoJWCrkW1/DAigQp2kjKIIHuXGhs4mEwjQGAEK4zJKMQcIgp51iuIsx1Mgq2b8u3iTU
RiI+QuROcV4/D+jLbpuF+Rx4RLCWHpR0njLK6MD/PJRPIHh20+ZoVWDfMu66AMXFnoDmFxic76kk
ePmU78oPE9TkzBLAHgIlOZY3n6RPnN1HvBk2i57oV6jdZQ5aLFmOfguhE7cj0qSdVn63IBIKT3ks
nhK0q2qp3PJsFbVSVmLz9OKA4Kx53TJ6YQxh7wPIf3W7HHhoCFizEyn6b8n+I0Afq0oZD1FYIy/Y
hMNAMlmw1AE7AKrTVgYYze/ks2OI09d1bCPwMuGMDve4U09l8dpeAZIsvzH6oZjATTa0DPQ9ZHKj
+pjfvmvImyAjpJ61X0rtSYr2jsfr5vZ6wmRADM44UgElhNfAUgHeZ7blY9w5eok1iTsdDgbPIHMo
EMQty/UXcQ3EK/SeOMrKYiyanD7zVL7z38y2f0sWFEZiBfyUEZxLrE6rHAgDdUqJTkM+BdlhOZyy
5do1AuM/6pvKi8uSTvd9fD6ozkfJTR0u3uoZ+jE+Bx9SQArL7CKKKpb1WlUXPv7vBZe8rKnm5cO2
Lwh2Ia6ITa/SIdlxkCi/qzdMhfAXLCW6QEHaTt8MR1NjVJ+pFWDwEfVnufNiwJMXtcLOjgamTcXj
esmvEryPA1JxsL9dOZDOZK/682Ut0WrxfzXOdFWzGcLY6zNRhUfRyXZpomop+HYxvSq9pqHcDc8K
hS1R+tCM3giapNqIM/0CXAqjvZdjO4OStxVdUROEzCe1dEjLYtdLRXIqSrR2SNRUn/RRduajyIpE
2s3ZVp7ZSNvNV2H2T9PBj6n5Gl4drT1zuDRZZj+dXFU9padVQLGCddKuyzTOHfaK2BGgYXr8t6bE
/L+snVheb0Rm/ODzWfrtzLlQPTzDm/zlqEyRZhsDRAgDrmMZJZdw+AmasZ2UF1ERZ2oaQK4CeH2H
Cp6K7illTDvWMkPmQ6ZBn6Vp5elAzgWBX7DyyBaXDVzp2w7OYmLujaUTe6Y8a9BsTHlMrC73O5S/
Kfnw1rjkgN4bSKSSHSPdFqoVR7YnHrqJjIQzXqGiU/7Nkh7Zy+vIkX726sKIEpol2MEAQjr2UuK9
gKtyumCdD3TjXJCuUyrdNdyEM0XdcbcnUjkcIReeAfhvjHT0pobyElfWVcez5BPEsIKU9o6hvwiT
pofaddigL1ZEGzaOMdcnL1oDHoipRpzFbqW2kdyvQajbazCrTgF6jD5C9FNVI359S/f3B7Z+fKzQ
TmBAcBjwrkrNGxHJTAUY5H+Ymhet3P1XyrxlQE6L6d2Lf9JTHYA7wp69Fl3TAgRTZYZiB9a6ijPu
VV7SWwD2zvxWWHGZEDHw/7w/kSzUcRqWKquGzijY/L44JQ8SSasRr7u2rfCidUJ3TrKAF8UJADr9
C4jtQuK60bzzLi2OCc7jLzGVC+elo3FKV2TyXiiqgNtMWN9dz+fHH4lgenODW+6w167CSlZ8Qm+R
TKexZ8JCSlSIVnp8H0LglEQpVN7NMu81ZQoGO0JZvH+gVkkHvX3BzTCjGO5KlFRQqp4QU5B38gtN
ip9s1SThu1R6jvnl1J2jufml2b5YVn1CshEH5OBTp/Tuu7FOR0d/SfNiSIPPrsLkNVePkZLbH4Bt
INbRUQ+1Ip07AKsqMR/xwwzwSRY7JBMdoX95nrAm7FHXS2iuhM+Fp3hUMY7j89K0c2pm7fLylDwv
H7xGaglq8tcC6NtI9FH4UX5stqILHNUJzMqdHTetRbl5Qxkp5MtqKyLrRIkPy7GluasyrHeSQujR
GofxqO5U8r+K462imG1BaUC5j4FrZBQfAKb+/OSgDT3OxMBQspWaUPojAFEPi8rT6mpc332WyG5C
My5NM0sgu0/MYerV0qS+tQ9unNBL0VLY7qYjaB4T3xNEsjz9PbG/3v2V/geU08wS8xg6piInp+tq
RU/xRB5bd5ZKKbYq/n4L37UV+ru/1zLBi4St64miX6YxEPAAL92kwaMOk4lROshnk33U3D8RDsIu
Gar22revmT5mWA9SgjZYxF20chU5pV8ltU9rizTGyoUIRFWjOqkfoYS7vyTGOxzbzHCNnga8Vse0
wqp+qwyIEcyVvyEbQWld8V9uGcBmfg3FV8gK9Yw0p6mjGwPOCzLUhbUu90Yb3JVCj9AQuWYp8zhb
zssvhNTww10SkX9RkU0zSBHfmgHnEF7mlgVq/z0fubRlBq/J5KzEaI2EmFhDsU5yCw5yu+ZONb3m
Xfym7mFP/pMsdDw8V5S4555Otw5ZpsT1/j4KIfA8OORogetvBkcPKg4oKCwHx62CcpjmS/MDCMTe
w5ihwv+3YeC6vz9eoTROjw1B//iXCqGYlGvqvC/t3CLHIZN85T9SZzYFX/o2Bydr80q5FahblpRQ
3YvhgECWp+syTNP80e+M08R6//nvFFYoDw+uP/YtlMtGyy4JHA0h5ySvzz+Edu3xorvnRak6FnvF
+I6HMVnULyY0mn88wKYGXA56uJzxvdcojzppfOk/XXq66FxezRtvq8Wysg31F1b2xNXJnd+aoIQE
1sDYci5lt7tsmBkU9enh4KQglnKPj8xKXnYv0osx0i31LHTO9lt/ZGsZe+AHQ14L/UWq0r+loX9D
vMecqB/jYnLNv1OGT3lr7E1ANclXgkHaHqYzEekp77H+0l6TdfE9aEs+FljsBIF4aStbchopzF5P
T9w0gRwy4BPssNBnih3niSMx+Y9zm5WSB0AelJhxPgA3/i4tVNy9cjmhKIuVldgmwqnw7xA2cz5/
Ji099kNtTWiRElSv363h9d1h7RcBoPf5tvvHIxVVgrQ74ygu+SV5EjU5/USP2TPBhk6NgeF95pYQ
1AZD+QXJbBV2otbKgtOwcune8l0xppZYYLQEBH/FIiHUoo8FRPTDDyuvQyZKsWbEugPJlh2eo4BP
BDtzD1FHQZFOZdT5NUT2v1FosU0aY4XT8ici/iyHrlgceapQs+1Vj1jw1lrooUcVf49JqpJwi9os
KR25oY/qqwV+B6RWqeL66ojfWmpcDmAvm8UKlaVXK2RD/hSHjODfE7DKICB5IMXJFP37ojTFymL8
FH/UTU1BIZLXHEohcxYzdqEncIGvN6h0YQo2GQk+Ukey+LsYHC/GFSC703wUAIWEA16KXZ3T6w/T
aR83UqnrJlVNtbqa+pBNUu8ffQWmEzqKmtW6wP2JDQhpO0RktVlIwzG/QCBhV+li8omjJm+A8aq5
CsVY7qx4CCgogVkksTnDzK1/SgD2QnrJ20Iu40Q1vg1uZU+tKXBYQnXJKRYPfj102IjbXDC1INQR
YLaOOPB73amMPn6PhG0rsilCMu6tZwtDDUSSNbfqJXsf8axw3xz8khhqYol4C9uW9F2zGX8NcXyK
SLhhAT+0qgb4f6242sNIr2LeRdYlPG7OUxeKqB2853syOy6gw7wqFuRmNYUZEPHyMNB0opJK7ub9
Z25EfcmQEp2bSle0OjiMbqAJv0iHi5Er4iobbJlQQo3cXHNz6p3vh65QcLVxsLvYIWSRnGJchOWL
eRsNW0/1BGXwBsc/kKTdJ1T4+jwvhTVN70MNFK32Xsq82sVP/GWEY4V5EVjqYdPd3lWiynANaf4g
gvLTfl9TlY4RGlMQtrA1chs7daOrf3KkRBcj4JuKA9CmFhSGQZJrpXOL/0/af76SlukkS1fA6MEF
9yGoK2MoVz+mOyyv+81E9JrqSSyqc0fJLeO7ufkOAaC4xtyYc9GYu9sNSXIbjXS9BEHFFuMak+eg
RbcI4p/7R6pqrBlHrG+au2lNckFyAzuTstSQqwhHBhRteNXkSB4Ko/u2uCbuZ6ab/obASxPU3FVV
oohU1Z5tbIL2Dol04bN9OvuU6nLTd8SD4WMehizDbpVs7/OWQ/LG5sFxKN15Vvrn4+1n7WWi/2hr
Rfe4g8RBBJ+gEJY78GN5MprcmKjJiP2LrJlooSOvkfar9bUCTDhqnJRY6XizJWg3Xj9SNfCoKYl5
eK2R7HQgOwwZ9kfneBu1SW0NhpaegpAGjh6jSYF+QJHDh0jomgQqmd7v/wKKXsqDLZ0iJd6rw01b
9Kv+50MP7urGQN9EXSxO1QK1PITxp+1Z8/m4965Rhbin2w8h4fKErf5AmQ3bJJTVSOr/iJempsjR
CDHzQoE3oapH1MuK1FUJWdHC6vReZguN2eupZ15KiwMfOeyXLgmXXvQs6ZEdFOrSrslhUtwonHsB
VqM9AmOqPNtCEc2g7TjJbmCXjZ89F+iUpPWwob0AUKVqRVz9g7DJGjLPfICGf4T42+QHoSuOkqMH
vLA14pGAyxv4lTTL2kHGjJWTAcfP/6dZ8ODcQBSi8xslf3NWpz8DIHPrU5a70XPkt2FE9pRXD4ck
wkZjFljrNfVi9qTEKURDJDVTE0KLma8xWSvHAsTzG2QJTel4vKQaYZDL5aRpVPHCE0JgRXuM8fHh
H8z7C1/HD1eQU6lHZbql8B2h0pufJN4sjqtvFejIvi/fJiwwA9rCvmxxmogr0LFLNvIIeV2AzXCs
jn1mac96ZwW0EPR8g12bg3EfHL3mZNaLvLHT+ryiiOwyE2a9ONS2UxhtNoVUnQ3sSFF6OQyL2OIG
7B45RgzJkg1YkcTOr4SEMsbT8dqvI2R2H1W97NMIIg678D3JseDqTiYbuuIUw3W5owvyJTVSzBCh
HH4LlMFIE+DQrQrF50ns2dr4mSfrQNefeDOXxkDSOmtDcDPZZ+uhtpbToc8jlycje+yyU0spddce
FSzj6JdHNpdf9iELh7z5UU5B/B59aRu90wvjy37CuHSu14k297yKQolykXSqTsmdG3xHtCSTakm2
4YJQ+bKtMU0MiTh60Wt4jwMO0DzIDFdlDoeu0Skd2b4cIPzRoLKWk1zJg3opTUWvMXJ4On3SbqWz
5rHiE1LWe74iAONPdIjg9HGire5IOggtAyFkNSNrKPLBNWFiW2Mr25SovSvPhLAbbB3gJNhowxqQ
gAMGO3BVYmost3zsEP8oU0NL2XrcavXbGov6dKUa+rXYe/xA0U3agTdNk3n0XQ1mCxHciYwg+wFW
zw8v5OJRIvnrH2TgJ6bpP2LUpcYz8aQMGV/27bbHkRp5G2b52McxNhz/K8dUtJ30TxsWHcM0k4kx
De1Hs7xmJPRKYPK46LqEb15kmHAvW1EJ4tYTXqPoCruU0rMtvr1UOjB//q31d35DfFjqlYLnM/Pc
9132bbRGUXbJJiaQXrsEtq1QpHMbLxwXrnnWOgwzbWhe14cX1zTvL1ma74boIiW9i08odZm/SPeV
Gemdd2u9EuqMsIq0Z7I3ZK/d+aNMLiPNMkwreVW6+6tSy5AuJXMK+o+5bs9i8Hlzvq3TOOIrnoWm
5vnWpYROHEGnXBh13csFaFz9TTV7pZclYz243pzhjVXEANRRUBYdFQXQ4U5wQED23ZLtKWe/gsXd
i/ErFV/9qVkj04xclKSI5GUGNyA2b6LIEw/Zyh6OcKSG/LwyFK1Ds5b8CjMeh+4GCC95HokEU6GR
EJ02Xw1xRgc7oTbis7xHkDT7jaenJVytYFg5EFRaYKN15mATKxor+zXx4w0ilu+AdWy9k2QQuUcm
PQWGZbCbkH/Y5iWqLNCvqrutWKTXPJLxuMDco0aIwyfLkAegabhDAsOikFkgptMKnPcBEXhjDl2e
abiSKQ2DkI6361BNYlXA+Di23vwSVq9Fa+4xn/xmH7DV6nuU271XTehlrHfTrctamYMHPONg2cGN
e1KGkHNWToSsi2p2lzoP63kKZ4aAVZzEGFru2kzCwfoLHfW9JdNw2s879D9d8tBoB2GAvCAZT4yy
mmAOsaUTyFLijxi8OEd5vKPOf3/k/b1R+LNcxEon+TwAQdk13a/taPCPITWaYPIX4ZfTp6eXirkT
N++rMjgffN0+yL8dLHJMIhV57xjkTK4dyV400d2F3Hya4SlYsEFSi/1QNYTRFCUQHmU/R9WoyP96
b/K5SG49R8RsxCAHTZZg4QBk4ePz0CoKMFyyOhWYT3b1lcE+naxa0wP4vqpclbUSGgrFMFwJfpOl
9qmU3Vnmkbap9NzzOBgyzb97V574Irz/fJ3fn4IDzyjhDA6REmJUM6mghhS/Pn4D2f07ok4CAuoA
NZ6KTi2UhTUbiJN3+EN0NYESJcZZG43G9eZjjnBJYgBH9Aqw+jSdn0MWwX/U3BWM3sJrMBNaOpIY
ZbKZAn6fSP97AhYqSTaGFCg+/Ksi+65BZ6yPJX2IahBRrE0qNfCli9Bpx/03brXe7m1n3H+FEXta
1MrGtwN277d1i73pgV2/1amvtY4/ruYYSJ4BoUw46QTpkMVztfzRBrdvO3G/SQc2McwyYt7EbI0+
y7k16ncGK1FSLzykuGDFPgEumb31sWsmJqqoj6ieSft9W4AQpluGg1zX/us7Vj/TpagN9xhXQbF4
sVj/+FoLJyL5cVbw1WjczA5ifmeSQ72kI8ux03emE1vjD3VjLDRT14swgrnoXaP3MVOTAy+9+M8q
OO1VyMn+1pagnup5iXJoPiBoYic6MfqvgCfwSmSV44g7P6bqFsI+tHGpZolOtPNBpNQwJ5I2wyBH
06wNiWhVQX3vORxmnSIb3mSEyt5jsvrbKMXeHY95fsprVs6yJiFRwyIkJKu0Yoog0jiu7d/49qLo
ZbP38GNtC4yxY5oNeeAP1WGC0ms3/ORrlR0QbIPFIBOTzt9MAspDfMpQ8Drp5htK0FJ85mfTHQoW
GrYB5cTQOmngBgT3tkOla5tc4VFi8cX6Zx9ulOmg4iWd51GqewHsYqTKikYhngnp9DVgJZK7SjIQ
/3Aqmek6vLJL2nce8uvVpDXqogOkjzjwkC+oNSFjbsJqFxfDvSRvpgDvI9Jx2VUaE13HgxL9EPGg
LyFPU+O6yYp9uwiOia7+DZvwhZSvN91n78GzHc420sRNdD5/FDA2WEZRSvhxhC+jBOKeB4Z6d3Fp
PuZIsG/H/8J/cV0lYuMOqb3Iz76t0j6qoSG1LfjNOEyaWR3DEdCdVsYhmQa1uPTWcd4MzlQiXlOl
WnwslFvi7yqiqsgzawmr0mQlgRyIZB3a8QRYtAp0Nh+TEHamhrXEMuImiQRDvYk+fWJRYDvEu4A9
2VT3LjMUvChdJfqZbDLB2s7vd1Y0UTie8f7Jk/UdTKjPjjmFk+D3UlU/sVTQonNzQ20bjYkMjgGe
CH1TNdSlLhPzXBxhvEN2hWK95OobjOcRcofwsl/7pXmQQFwNaTmS03ujBW7wiZurN9R+fpo/hkl0
84A0wNb8CVtwj8IGxSH3uvojBqv4TN6SMEjLpDf1sxFHlgvfLiIEFE90Iq9+2D+Kz1BkIIXtJCgm
TuF9qcl4D/0FF/wjC/qO73RyrsRi5yFZR6LXZp3v6kFeQRJIjAc5rSCfHs0i4bp2hCfGNU8rUnan
wLIDsN7RwexakFlTxRIP4Dkq4EgzCQkjqmPr3CyHwKzBDboTnPmbTyhlnS0/z/qdSMhiDHWIuaKn
wNiL6bIw/Hwl2PN1qnilI6EW0eNAcuSO7LJCv/zEYmvKdgJOZnXZeKB9Ei7CSkPzsou/6p8stvyl
WWLwbtrkVsBgiBdoILJnpEaHnbdg/Khr2m2oKevDQxTh6EAFq/OyXmESZuC4TkD5QYMUIXSXNZzw
R5b1X1afD0PyFWj8QOu7jGvDVxZ7NeVSQxBqWVibAOS77TG9gR0CxvuHGs3HIr2k7RHWtP5psLcI
Tz3wF0WBiZiw2DkaQVO8VTCSkLcVYg6CZiRnttcJtcBdQ19lTBA+QWtTsg7pTq2bg/6vHxt6ZjGC
Ged0wWO2U09bPylyI8N/cml6qvLOoTUPn8HMZtXYkWN4PmcVaK/7bYqTX6AsFTKHJlBpWSBCax78
+Ei0aMNURFNZuptHt9HYYj3HBL4MOnU+aRK0CXX1gbNNn3EFgqEZaW5tTEhYpiwT+kgEnE6sRC+c
0gZAe8Tk0UdpngcyTPrraY6gulXA+zv4u0gdsO6GLPhe46RdouKY6q4f9SKQwkNvdX66cP6qY98u
gbDA5behQDHsZRYFnKh6PpkwfhNzJQUGb40+TDkkT1nlf81qYQp3JkPN8C6Lg8XzKMKCNotFuxCE
g2o/xtCeIRNreMVoBMkLYSUWgwfiUnieWFZXZJb6fFF0uCMITpziG6HtSHnH/q7F6QpN3B6/ZiFw
d3GhO/fqoe7c8PD3O+ype48Hs/Id0ARm4BuSsOMK5Ek+/e6NmPlhLgQkEssEsf8aXNVwEqQeiSbI
MIbN5Y0mWdI6Mkm5XlBA02vLnVpf0DChzeGlJWMvWZOJ49yWN8VJ8olqIF/45HhBTz6JALi8TwJN
sXJw7AZCCCHgxuDHLyRaM42NhvcujDGHeZi+MAojx7NL+ovNNklUv/BaCnLGHAQFhG1Rw0in7HUU
2vtZ6rXcQjUhwJOq8DZhQMWCK8MyiCBlZoZSS+aF5yw4JFxH95TrHP2QzXmU8X7unXzSiksMjFoX
uzoRu+Z+wPVMEs/B9vHfeFnZqCZaEmDbHLXllo2KqvwjUdOsyAUUMo+sp4LN3vtdObt7grSQAn5T
zMsJWVmooqErikFT77PRxwiFYgbINhbMxqbLir2R7QXFEnIPsVEIlv/oGQnl4wRAvwcVkDVjZl2G
tUhaW5YJyzrwFZ6SyyM0Y3UHCtfCgfHFJHIiCLkSzmfqoHgxi+FQiQKbI+OiI/LBYrGAB3usCtSW
Fmzs74s/T3/CLp40LXZUr+MCCer6XvMqWikisGGZ1+YAVdWD/xFxSYoO6G4Eu8rUyRnEiUb5KhpZ
9MO1Br331l7oivVVkvjtqi49GdeLivR0lrocTPOs8LGzDykUNHfy3AczuMepv8252GBL1lhAz/ic
RhDHbRiSRdLGmiasoi0FfGt3YL+3WUk9mvoDIQs+/sEXp06lyB5fnypGoxWYQuaSllm8134LuE1f
PfgUbsVuFGrHuu9jocgKGsOXhYMz0/If0y1Mx8e0aA5F4B+An+mYEKxHOE7t72wdJu6qxYFrgB2c
f/NVwr7raxmae9jVc/gza5879nIY0EVH/vxfRANML/E5H2UKbOYEhPfIJMm4I+l1sW/cQZiGhghz
3peZNzIILsKRhDhg3uGbAWQTDZY5XUbpmmnmfuR88JXTQ9OahxPFcr65Yj7D03xanSEAKHbh7yEG
xkQ8Y/ZLdZYIBUDFKS7rCwsXeyK/ZyhcPUYiPTzsFYGAouTz84vJQ3U0wsWfrWiJ9CrJXV6wlDO2
1zCOg7rCwdGb9VHbVtX1cBWi/9FKjlGJF9PnNN3GxkSREduM1v+6SsFSjHhmN0noM3/2E2Q00idD
TiAr+04fs11QFoGLMntx+ufFFVexLDrnWxYPRCdPFOEhoC0GcovqxYli1yz7Wtc9n1GQFtPF3X6h
9GcOQtMWhv+9ZJSwE24kcmIzhW/O+0efJA1QSIX7qc2mjzvDeMOKh/4glwABelTwcbhXgJ+XmBEt
Eko8TVd+DmBjeAQrWYveDzwfN8Rbz9LHoGsxBCHR8sH5dOxNwNfRZ2SmryJjeVlYjJD9EBD8Hpgo
tjFYZKTFhdigBnXho0RHrjzDJGwAIky7zfOOe6jHBc3QgFxHSU1etZEDFTOGun3HfsWJpckXgLKi
/yzId119i7j8F2P0AmnbSXesDbS2kkHYtm7JsyRyOhRMV7JpoFiPoFB3VaDblwJq4MprcH8HzUxV
4yh0Iu8YSTyjR/uCDPIPOkQWVZw8rO2ZgfB3SUjsDcaK6YfYMmgxZSZkF+bU4gq4jhE/8vsDu7GL
pKzdBLek15kCOgb9601ynG/uLDkduZP7PXSn+CABKQvR/vtzvzIRH0A54CINaGDLnM0+uj6I05UG
AclN+p4komLi/mw5m+WYRoTnrc97GFSsLFIKewc2+BTC6CJl/vMZ/ExvZMCV1THBRcYmgTHWekE2
ep/GQbbYBq+Q3UgwzchbTtFUiD1HB8l3G58EyGuXkFFHvHxPleg+YW3j+gCany1eoKNpHWvz+tuu
Kr4qfJM+fFE8UK3ppL6moin+/SwH/eoaQshNWVo1IAFbviqMDMCkpmrodl32OdmU16C3MlTfyM7M
LwIB5sHBSMDd9wjdyIoLt0/9X1DWlp8DsZ+Srnw8Rbnp1RyBqo+KFb8aKmqvB5vElBEC8QEwmFhf
7/8RmN31pRPiW3/yAUUuS82Uj71Sr4/FnKJU5NDYGL9tisT3yR6bLNrNIp1HdMOPQNYULEYiwv4Z
wbmlEmTfjp0T9ucvAgY1RGS9VI1BzOEaV04abzy+oi6Nb4FPb/ma8VVLhiDzlEXi7ga7WIt8X1/x
/HVQD49InrhQM+qRv9jIxS0dxX5XgOtVrs01VNFgpFyqLriZl+4C0FE7t+naTB2buLayA0cZVYt3
JgVZBgYVf6AkYUpKylOfqmmyLN5CeNV+/nxjm2Mf5NIrwMJa82Hi17k7aSoowaUhKiTnokYg0+88
0CgRFwgiFW2rMcCk4QckU72F9u+PkqpL4GP4tSF9z6cs3TNu0MRs3NzBzhUOUjQEMU0LDlEk6qG4
I8BGUniIu8B7KExmfhTgryMGG8t+MW3+oIi1BoOSNz/wgevIs/IR8zwDQ4elpUHkBht0/0nkkGpU
n4XlAyMAdp40hZpcIghLAWOE0Q6mKJjsxU4l4U3z9qNzzJEg0bB2xyWefb1RTYyubgUjgzfONKxd
wQk7TLyRzpRCJolXfPvvD7t2wtMa4yABtEnTtWuia2nWImaos8DiwlTsm/ysDVhGMFE5wIdnA7xE
Gt397V+wf0T8GrE55ibCt9MiDE1ah8KO92jDHA1+lU6aMiOkpIe0u4LDcpEVwhRcYlONbKnCme1t
yroFAyGrARtg/J6XvxrURlx3BCLNYGrq4k+SSIGLhyjYo8aTYH59nM+YF0vt3eCZvRvbN0cg0V/s
RQYXe+hZTPtYUehrq3NX28ersjyYB7dSQhAGohEpAYtP7di9OzkDrCbuKOaFo4jf4Q8doPiymyyN
NfYswD7C43FcmFfJUlJ47JR07EG+oY32wNNGwC/tSEszxi26KdoDK2+JXGzoff42KehdAffka+fR
CAzFZ18LItzBfFFCx9+MfJLseJ60Bg2q3I6jMjAA/1fzAkvJzOsYhAQuF7vFmiANEplaoZnvR9bL
08aBGERGmDImIMAeK9kc4NKF9O8J3JIPQZucFkhq2COKPKwwll7OodrLbaB6syq//XjR/OwA5Hvr
wPplqS0z4UaJIZln/MuMrByMyIhSL25r5s4VTFvhtkq7NgRjZDygomgu+Ke+Wj9hZfo5UTX5X1FY
eMdXDmDDCBuZS6htN/hPm2WiDrJfEVvgrrSoIQYEslvYXLrUvbiHlgrrCvVL2Xz8RFloyiWCq8SJ
8XOHgAh2s8fhvBYyGEv6ozqsWImFDCP7/0zLsG2ArilFEajurVCLeY7TlMFXm9D9aouZW6haj7zy
lSC/7Cvhk7ZZvnmldn9kSlsYhXy3aggJrln9d09jRSJ6XYPk6ajLv5KzjhtSCDLsUixWMeI1Gxvu
UaHmj+W46ysBQOfysSnmOYqbNzHX6WvXgYFBJCzuxq5a2bmPA5s2nzZghPbX4uIzid+2YrH5Jd8G
jjiQaDQM5xXwY4cwA0drbNDgGyV3/FKW5562gz9bsUyaH6nU68cDv4nk8t7ZmACtSnH0+jJFfKSP
FII52VVThJHJFL4FsS5PcWlxUl2eaEwl4qjoLph3V0cXfISuDPoo+ubKl4I/qScVyrxLcu/4zFal
2xmXkgZmZaJCYM7jFNDOtOBaKbK+6E42EsKWht4Xerpv3RlvC9N/4XskPIHYjMWB3gaWUfJ0Tst3
uuoxL5gl8EH0Ow3vwzdcPHjQxOP9mELFJhEda7hBhb8YC92GXeVAd4XvZOkFUEm+69dwHzj1coaZ
ckqRYUXDMkysM0Rg6Xrv0L28jHPVG3aP6LZ2wEV177SV4uTTYfrmoCjpsz2Dk3aeabT1mb8cGKrv
crIGdktwkeSwtfsBsFWkPMuLL5zDm9rC7W8qEu8MfXF6yTnIR4DAuzRc+JxioIam16clS8sKkJJU
aGpTmXdOOrMC4vu/3xRwDXRhEU5w/PMFdvQmak/byPZCKDlGmeaUaIsn8QsYZmbzmqkDUM0tlg+p
CY+lGKo5XDQuM7rmsmyPKcVQJnk4RvIaOySrGBNKVON5dCJEmubzzMAGLFXcjTPSlE8CVIS7bic4
W46iqF/vbOP5Ti1YgWN3/QAGO94GqFd4icmagR4fHI+x0JBMVthsnNXS0JWIIY4Gq94sgK3BR8J9
2pk4fJPypdZ6xD2U30sCT1iTIHNgKHJtxSVd9QeuvfUnBsCB251wiUA3OLgDchrKN86TQk7Cpuw0
JLdhbCBIt3XCTSdKu3blQ2I3AKyLzgzqtIvZMW37d7IA7tx81I1T3XEoEvQagIQMnD/62kbKnt/g
glIgk+1sHjx2wYqXo6y/NH4CD4RobY9LkHUZyasFaGUrBY5aQdbzY4aJDAl9pQzNHunpFA98KkWM
pdla43u/oQ1hdJrtaaowdMK6HhBEtaGDpy9EPbwKG26sJJCMY+pRDsJ3CS55Ku+ooVDjmkpxDs7J
ff/UuyC/OxXk0xvrxvH69n2vsZhSn2F3Zd68nVJqfmTViaPL5FG4aB/+Yhhuqiz9Brjc7+5xX6Q8
wOWu54FptZTXmGuu7V9My++GaArtf+1wT1VrjJYPf4YpP/BC91VsB27HmMu/vjxHFjcpDWAvEF2n
MQXCHnuE4csUhqkYi3KliPnPzJP1Q1p2DEPbOdX1Rt2Ev8S7mNDBj5XdSRuZZe1cw2r2ucMi1GsC
6iJIs445ajpCXzmQQJdldHOvUuo3JN1u51mXPRCgkpWHUfG32hZGMCnLiY8HL4O/nXF+aKcpESJ0
rLvjPcPxevFG2BPeB6xVu/5EdWk0oDJC1+nUvhNd9LsHPbdg5YhL39ySx4p2iS/PgiLbnkTbwd/w
Eoe5sl2O6ZLwyeP8YhAFDlY+zfi2NaTFU2eXKAU77qaNhKxwsIdxsW3b18M3vY0UtpkD8v5T9jhP
2gCtxhXid3g+OQIu1xlFgW3p8JMB4NBmRGJ06H8reBjMUfVYae5Pt1sFNld3ATxRv20MdJV2dV8n
Eb2B95Dnp38n+gDiZnJVQJVu0kOES35WeJ9lA/KQuA8OKlOdDFwZv7UGMN+H3ZJnnXOqejUCo2XJ
Of1CGauCe6WE8bOvNzrhljiuFhpOzjIQBDHxt5KRxyVsK28ZR4LIap7qG0V2DXAklOZZ/8D6MDA9
gXy24ypim4XaGxN82CBc/6E3Bg2EaueDCBrEfp3Sk/wUVdZH6pbaiD7bE5I4lTnBetN2iiJ1Hf8+
CiEkFTIWvEC9sSvAwE5IuINyLTLPiFE3sTdDLdP19pDmGZjYTQdEns9B67y8tmKRj5W5drcP+vTs
7BmumMKEMiKcntqoeocWRn0K+qWT5HHPOvtZ2mmPpaO0LLyFzdDAIWiDG6c8JFpTt/HfBca8tBpN
xw1pzCovK9+H23Gp2uDtAGj5jp9UwYmxvki0fEErwf2QlfKKZVi1cUCLnmUM+K365g3sAConcUAz
VGoPxjcgE5G5AMrOTtLX5WdUrZcWzvsRfzh2Unjv+koJMaUaTj7uGMFKiRAx+B2jHKmC/xFOOiN8
nhgM9bYdR/6x5ZRWZOdYn8r1BhY7NXrySQcDFsjBEolJbF4Mja8JLFZOCzkinNaQf2wC5vAeJy9o
ta8YorfQ3IdEQVeao1xhPtk9eZkWDrfPdvWRzoYwe55wvoby0GVvDBcKFuTyEo8v2q4Rmm2QLuLc
rLBDR1QUJ2ZKmw6rLuK+YqrNiBk7QdBt2ygD3l/Jjh1/ALI2gaKj/hES5vCh/izGc6/7yP0HqaXx
6CnJQnqjOY7Py4Osm3bMzm2uEzCCcaroRUXzqKQ9Qs6NTbHCB1xkR+TP0PAOIK+QYhXD+nb8EuiC
6GXfLLAPqt513a55EHdY9sO6IZg5MUYQUSr1LIt7O7I3LXwTMrgV+IWtQmbIltxREW8Q0QfMQNxs
BpZ4zQAeyD1bzWNr0cvu5Gefv6NK8hk0bsXXCn4b58bw7/pvvnsWd/qUjUCmwd18SwKEDJfRG5XA
MBX7K1DgO9ysyml+X6IGyjut4vYIN8Di/IOY3STN8+7DboqLKgURjqKMWWu7IBE1H49c8sw/l9OU
yILu/u/q1L2/Ejp2rn9djepWyGdauYFzxB53KWj+OuCSvyOMbq8zSqNterv3OnlaFyRQQax5Nbkk
8YOfyAmKJTD6Rm5reKmW9oI3NG3jJEq7zrDa0eoR5AVEbMVfM/Q3P2ilX8EZB1NhLHC+NhzYd5WO
wOCRRtbHDDFQ4fMMuATzBdpEyMm+urfCA928Rd4Zp80KajOd0T5gBEZ77kXg0KBcrBpZ4W1iWZY5
tGsOVt8AUde8D8mb7uYFY46TMn2ALNTxjQa6HpQ4u8Jk2pG0bHYaYzZxfOJv8BzCk0ocWGiyvIHy
19nNn8TGaDIzMEbWiYff7Tsa/kHXgKHdOfHtRq+NWNL0uHzhWrrJK8Mk39QSe9I1AfcI+MH/7ssh
dS/XDtpq2O7nl8l6nkD58ZQ/yw6CpiPFO7nFhruKBSiAKGaMjY5L17/vqxapNtTM8fXEoqtThTUR
ef/1feMwdKa7neWoysSxi3yjVlHgFYnhgeypAlk6dwkz2s9AW/v+90zkxN8DCN9TLU1iM16qgavv
u6KIwmJ+no+3aXxjLfmutiZ/jdQzPOOA97JrM49TX5rdiTdqNg8MmD2ysGnP5TkWr3UlAByRkUiF
dqzctOyKWuUFUzTxIP/F4D+yJOG1m0b1Sv7FmgokvMpMpgj3fgpgUYwE/Rt7ttMmRhrhx8kZ6lqu
OIuaIDTQLGeirwVL6n9aq4XaZzpYAWLqaCwajYhZ+X6tXxtKLPyUYZLmKUDM6zltiiAibwj3Nm0U
7MwhREOpbIIaSQ9P7wfLwH2znrU09YmDoa74uBd+fsd08gTfdi4eNjfpzrYcwi8WA1WiDZD0/xiF
u0jTa9TjpuBn/ggGmE70YWXC9Ao6Is6a75ULHwkHppC1Ew4bbXIl1Sl2N2MGCOfAIYUGkv+tWbjb
qPtTMaHcC3hoEqQCQqspbkwbcu+1xsVrbP6L3IXUSa+7DZCXEV5m3IVhezb5/jt7lXcTL0ltSIpv
9S3Cmu6yvQaWlrhzJ+x3yWTBEpZ6YAkph8oqQ1WDVsJc/oW0I62rPZ/3PT5xU2f229dn1RiRfZMU
eXAGQa84/WPfqxvzA8Vu6qkbXhSRdqtKlPM+atmXEb331ac2r0qrLKp+rpxDfnx6J5I0tBwkcCv4
+KwY7M9Dsrj4+Y0SpGDgW8MmwO2Ww6ofl4NvU9VLEDJ7x3XxY1YV4ULc5azOroQEHkyIJZdlMkk4
SgGFbhuQdpm9kqGNyZFHxcu0rTs8BTPnF6d9ebkA36YDKHwQ61fZuy6sEWrYgLq3vWW8mIm3Fz/R
1Hn9ia/uMQDLzVWJFpr8mqjELuzz2wGdbubOxprkJpY9PBczzDiUJksc4HwqfSLmMb5wFPs/MXhl
OEZ5xFm79/8m5qHA17O+7y0ponYvdsgoMPoDEHtmUDtxmpePnwre1VCFK5MdTx5QOpuW3FnwFqKy
o7YklpkpLNXZ1Ma3JcVlkwaWgv8p0KDL/96/gcG4TgBc5pkdF6eO1V0HHg82Y+c8QLDRa2gOopLc
WTeVCaKB6063//wjX0eW13lmL2WAnnDl5hgTt1ZnXtjwPqu0Qp3YIXTH671YAZ+mzBTcmLZe0GVA
syYwdG6+HUPcGNorcD3FD+hf2YJEfkRGL3NRNObyDDIYwoER36r6eh+837qTl6ejY29JNshx/KuR
PlHlo7NPWropTVHbVQktp7B75XiV5BS0V5t91lWIWde273+2yzM6f7nIswKGsY3ULI2qGTSEs0fS
BbF2Uwh8Lvb6iLyZJK/IHyl/H2VUHh+MHg2+HOQFLoPfzGzgnY8+cCfejT+nH/XO3T2LFBbf87IY
P1N6VLkOaiyvjQbLxqJjLhrZprHfO4CYARWfTYHqNFBJtXHYcvzWVOeEJTSY/DiHgtf75lN2JiiW
cZPYnS0VYUlyb+B1a5oXXTSYtzcPP5oudxs5UbBD0rFlltomB6kAp0VYCR5eytAbnT2yzoE8KAaw
2WoXXboBjbRBPfmxBy694jS4e6urMh57P0412B6+zOn307NClmGGY8A7c4mobSdBsY+4ZVsV7vPG
pTdoC6Ry/u3zv6fU7T5lNGnnwp/ared2Q6IjJyfL+UYWo/uHrogPpAQ5YxoYpvT99XtyA7TbVLYJ
BqH6NHIXxPobXUlCClavTgZX7nBtQ6eFVrGucfc0CD8gNvxotT8g3ZhxK3z1BE3udOLgsDHhOjfs
ySIKYsd6rSazvGodNTTby+WpdznZYP39uoCIdqLrXHCGnPH7e7Kk7yQU0GvCn9+vvhC2iTp5nL1b
tMGGgxrmsuYIxqKgI3YKdt/IScShnPdutnRlnVgaDS0TrrwlVLbZ7S5SBpMVFYgl1Un/0ojjSAai
fTJ/W6A+0Vx6bfZVm3PfqEdXLNcp7qP2eeWIXlwInF0UGPP0FwyXPv8obechV6r/zbGxMn7Ua/9r
bE1xax8hc6HUg+L2q8dN9qb7SrgMeRcfWYjG22OU+WDjTADXhJ1WqFyINy9hId1jQ+j4c+Z5DPor
mzTWhU+miBofpvZQDB+l0x4CKW9rAva5lIIBaXPIiitda+ROCLwMkWiLCKgO1NaBOLJacO7tgXKE
OcCQOJfEAhCO8PopqCV98hCCTtNNl9HLAo8VHIQwrx4XTfBoahFqqvNG91FaK0TbjuvNxWjJUCgF
MdlQnuTD+qUWjmOLzUB+Y1qfb+Takzb42UKShcAMZBffEgxYfcUFg6vQpaS+6/yQ2cuYK2miU9Mx
oGyg46/9qHlWPw7I6ULoMQG/StqrD2SGDgqPU8GfPZ4TZAB4dtfqy6wVxCghFZWoS0a7SJgCkXqG
cYyr0Sd+jn1qTFfxbKshSeSERm9RaEpxk/cRCGpLJr0KZmvJeVCpdG1mBwWHNnpcNKfL9aBqepQk
yVnV/C4FMBEWGaCKIh5oxYEqWu5mZ4RDWisyxbb1XO8Ydr68QJO/v/7Uu4e/ykGtI16EA56p7gXR
ipnLml+A0sAzt1kpBF74S96S+ADOFBRfGS/+1RDNPJCpcnna6bl5FLsJMUQUmp+yYkbVCQjeMfRj
66rWdG+XZQuj6+eJS7SQUkGI1uiPEXNYXGH0QMLbgglgXYFCkQZSyAauvozHbh0yzj4p3N0K7Neb
U9Na9ZRWc9nwieF/eaSVVVIrPGzSkfY8xriLA/RMzOlbhhTmDxhzlFwmvDim95momMzjI2oYQIM0
6ITUX63+Pe/BkcjML2pXpO0Ogq+ilN1RfyDkEBmLZy3ZP6lu/DF95Q19zJvoiS2ne0jJ29XpP+dI
HFGo3eL8Kaa8gwiacJFvusCyHWvHIkQc09FkkNnaIWMpJDKwhzjE91BdRBIu8ripOrdFGFMMZKBY
hyjSHMdmOjHUUl3wb5SV4M+2bvlvvAhXYB3yV6H3mdq9IC/DT2aHuhR7ucz14sAYKQN4Kp80IoFz
6x/zqLAI0ZR9fHtc65nneAgmyMIECnxgDWpNNz41EEvXxCG7NKFDHiuGfXpALfttvX3ut+47uuGl
oo4152cPrMc92XBTdQQFyw2Q7XddWOyeCrqwHqifQlKoc0I7mcMije9HiwaOEcQj39bwImCFOlfu
cEM6yH7J8ylLtj6xnGanXnXpUHBqNtDkDIeD+p6DRKzxcwf3fFu3POJOBtpKGBIHxkjKKrsEO3Cp
nOirSjv/t3iD3+RSU3pRv3rZNc5HXPkj6En+NjygOex9IbkszxaA3fRZtQhWeobPJd5kYe5qaH+f
ZDz3m6dZO8wzn8B9+yzPKoFoonysbvO0mitZKuQSyrRrpIxD0i7ZZskEYP/yR2eprx7mEorqdPpV
BbCW++lP/fCX8ex0pXblezDTMYwmfD+IN/52UQpnlLbGf0GyQ4pXSIyjCO2sN930d/WSCkAYB775
IS0g1uaa48VJiAllWg8YQ3VF2PgqpzKoo0OiMpW5cyalDXALgdnWHcj/q8UekF/fGK9oaLP8myZz
07O3n9OKJQxeqwS1MWBegCD93qEMMA2XXBqC3Ibr7+9KL9G9YIcIwj7rf1vg9e6hO2LgxfXCXtoB
FSUQBaE0gZ8rurbHBLNUL3ovBZh2ERoQjeZB9RTgOXuI4YkiJSekPMSONI0LaciC0RwAR6c0Pof9
X9bhq145AfJTV47OM+igs0iMVqbp+A0+jyHUeGe7p/fH9tztMcVIVNuKS5E7vHMonE7TZRrfRPxt
SZiQJmdI6DtkdzHb4xBlSbZ2wZWFlyMgHx79RxHEFl394oyjKz3otZ78MUnjmp28i3vlkJ1WYJne
1uEzoBuwtWpfnD7hfbaEl55GXW5wHSo4XgbtHSdWYS2xTLolO4ZkSphHe21DjWltbKKzYja+kw0C
AdSFqPXRtm6nWwmrjaC6lV6edVq/5b9Iksjb8Mj405wqj243B9jiP5oYnrSPjfThPPwnGDmx+mzf
8diHwk+/rRhIMKcCJ55/fmpvxkuTO2RjMn7LWXGBoIiAe9Ut5w4G5oRKVpzdN/qoUUV+jJiZ4WAo
sxxojzQjDJB0eJ1Ki3CJndX6Y8DwfvM/5HQCem2Al2gr5sJXdP4NWur7LqEGzk+NNnAj+C/OGiiw
MH3m5T5Gxw+vfKN12SqS5JIFCEwJ6K3C839MbAmW9WM3Y7mvMY6j9+1ifoDvE3BpquIIWynXH8S8
B6qX4GFoDfTwBq5t8v/xItmcAAvBXIaSdMACyb+248UfGEBV/s0V4YWYknjizgQNLrtxu0es9HJU
SZeinscTsJE5SfvtzhuTOh96mXmZsl9eN6xZASAO6P+Atsx9DZxVZLcyCuEuksVWsy4Pd3F4lQSc
dCT27KnvkXQFjKpWwLq3aFzlEDF1dqdoSNExDElU3ezxBFuMN8kX8cq6iKlJpqGsuf0F9all6Zou
6FVm7bkQjJDL9KFrnxftWnTtlYfbRcn/83KHiyzcMJbfcGsgf+HN8b9RbiNSdaQ+/pDy3BpxKMxB
dTl+rdZKHb9RVOcd7vRcLvdsiPpB4PYDQTG4GCR7+bjHcMLJQuqe9RnbRnaKIOrWDzauJMvXGaH0
MHWvGAc7dDUgLgxavyK9X8G0nnyqFQ4dyOsbih2M7BDekGo+LX4TCdUGfdJ/ZOfXpPzuVgQvxJV8
uaplvu8k8Cz2bG95+FEQP42c6JCVe2d4/YWromtQneNvAFAdHhPU9vwGs5VET0IHv+TzHDJGshQv
nLhpVLYYCEIrkhoyB7BZ5v6pC542W9QhPSmGG7g/y0zGwMnI69IhOsR9CUJaW1jeInJEXYaDKFx8
WDZG21gt1JF0831mom8ozBxOHYALywLj1Nq8Xuqh7cOalzzXQsJMphqxbuVpPd14vmR7ieqY4/4n
6MmBT2yT3sbrVFGAz51r14K2IFH+HL7mKshFwEuiDn3KVCB/te3ZDgbNPcr4hLD8xDCNmsJznTmR
Y396TybneWBLjc8lWIxm1PAaJDYDi64GapvQrGfoa2mYhK8+SWNBXyMnv2tLBiTXN4+eBWxoRwHu
CIJcRmVomZCsWWYAlGxhVIsm1j/afTloHwDijvVKMBxazYfQi+1a/1T1lDfREp3b6zml9Ta3nBF1
vH3TIp0DgZdGeV9bqmuxsBRMs58mUtai7C6fVUoGfX6QFWbgSHub99ddSgzgTRrXPa0Cwj2oHSuy
ehw5Xnbg+bnEdBBrKGCs4d9+VgjetbClHFd7nd46S1HKDt4OetKdJ70anb3z/1r2ZOtR9BtC6T/U
+V7QuPeRGd0qF32OYZuvB3fuEcVhwl6WBzgPYsueWdOxG0asv8wUZN4styXUiqCZuR2QklOwFwS1
Mo3GPNIEi45MN3KMhCfuO6W9QBsIQvOdklkVM1/PRodfu24RP/kUxFiswLQBjO6pfbCgWrUSXNSd
We1a9KxA9iYNoIFnM7QcC/RH/SnN3/rVK3fb6Q3otNMfRR6hZYvstMNvEDFBqQWBNs2vtwybxM2U
7xz6mQamXF3n54zbKCHMdrk9z9fEKFygZIRIaiShyjbZITrRdt5LZbYbhNs5i0xe1gpbA3E2c7Nl
m1zNRVbrQ+cr/2x/He+Rpaoc7538w3xw+rlS0OCfCowe1my3F4dk0dgAOO4fA3ROnYI1qN16gEYh
OKnxcjDGJ+5fWbVFhdpdkiPd9r1m1mI2pvUvsYoVyC5SSR968EiQYesjo9tfTjJGkwbTcl+WgPsm
9hfz7CIrx5LceEDs9NjGVLDGZS9aUchez0s/XI4+h2uDyOa0N0MJy2RVHYHROqlE+tox6L7QBlB1
1EYyYrKeGbVI9Pw9Rebmt11wLFRqESS/jCbpvm0mXpb0yWk14qCGJj+zJikp7hMNOSsvvXV9H1GH
iN4XCjzGnBtAWu8E42nafLBEKkgbkuH/5ltLsoSmvktIBO/9HmYgFPrXTXILa5Ls6wrs/KmkOgxK
/tTfLvkPWGyExlkuNdV1bkRuzJdzkAWPXDGPQFgP+ApYdBUFcwQkYcC+t8VPnj+sWybGUhMD5p/o
yy/HL/3mP6ul2RYD2//ERj+oSmiOmHbPSBno6H+BtTWAxxcojUlAJpEbtuIZ4ukeW/URgWyDMUW5
fZX62AOKzRkTRuqYHR6f94cY0SkPd5QOA0x7adbbn7n120eMpPcTUbeooyhsyXjrgV5CoP52NzNY
uV2J7JkUM/M0SqymRUFJE2GXjO8mRnGI95VqsbzIW+SS2Gq8jpuVjLUfayCV3DulwdfeWZGeKAfT
ghJhMsMr1y/hqbuOgEk/fyB0WyKzfbjkzOPwzdOFIKooOGduyWo3tj3HCxnoOZCJ3+OTXzVrNYwo
SyqaiZqm1US48XSatHxqwM3Sy1bdp1LRxfxERAbFSy8GCoryOAc9au9Le+X5bX/bnDl/vqQaPENW
KsLVCUtkEYAKYITben3dtEjRvkPlrOlceioSh8yEIIoNtxUCDE68gIZjpbE3wEsPGqV9e2kO07H+
AbgVIv8Cdd9XyTWbrIkxz+1NI/uA/SmShMUb1WbVAeGgAvIAWakjXCCJbTyquQYDS4NV+HtCjAgD
RRwVfsGuVHlGcsuiQYAZ7uJqlJZGAgG1n2RkmXlGZ7HP63j8MXyBTIiH9AFJ5AbH8JVM7Y2bo7WD
idaYG9/HQ8MQ2nDBbnc0sPCexdO9ZbOJOoW8my+AMjbUq1Erq64b3AqD657tLXUckDmCwaxV4cfr
qcuqpAdHl/ECaDdVrBRgXgRLMXVLrEWEqz4tzG6SP04RcjwioyPGKqTLvxamalFjaxltCK0MzkNM
r/z1xYFkUbJ6IYwtN3BqIg7sqjRyqWHAue1yubBVLAFU5DvnUoPp565xs0jAhL40C/0vJbtn1UL/
4e9pGdy+aPZnCBSubNaJr8A85kTJipJ/0qpUqHZr4ynZm7uLCmOaW1cl8T8skcY5nV6Of5ceYuAv
wcGm6xyfSpumh6SzK+fOFaM5Ff7Tg1qhV+2capNWctQmCH/a5s8zKMD+AOl1W7cAhjj9Bks5WRN2
DDk1PnKnqllr/WOvzaS6xXAO+XvO+r5goP/W9QicM7LXiKEPM+DENb8jBIcZLHpvWVxjeYPVVcwK
xhRj3Dshon3Xvcbej5dkeXgdoPAxohDAfsbKcR+iHi16X5DIwn7hQND6qnumNHpVs1kaB453a3If
kgGdOlaCzEQqpZLaHWsKXPpVUHZrn1/DHFmdf5dh4vsfMpa95IbVl33cJ12rN1I5AYpW7M0dw0WV
brmVRjCfI3DWQifNqNAwMJPZ/nEWjPInDcEwwZZ8wNnnw/ACMzHqU0SxjxjvlrsHK84czGC6QQ9C
ZXBC43dlc0HNQV4OzmRRyDB2xdPp57ycKUAEA1tPPWqZkyKEzf2o1ly9qHfiQiChHuxu1kVlS2RB
EUt/fzT659DEOXCHbZmct/LDFgCozSOuLCoTzsXb7z6L1AebFOiAI9PIchB9bp83dlnhIANApzvW
aOLN1yLUCIhrd5UApuvJxiQnF7eB1ahnb3OryIv9TrA4bof1T/aPReOP+u/IktJlEaLPSwC7q143
pFht228mfdCrkSCvOd5wV3Oxl7IHBuTKnVvMH5UY1i+WJrORxKy8u6smWxw22i+22X4yfE49p42o
J9tOslxHRPX+e8vQZGuU50BQ6DkUFj1O4lfpr/8tBaiRJeY+sMY4gHqeWQuQuEa7dDV6ivYekv6o
KbtWv59mBYhsQRkBfu8nP8jiLmYltoxISHCLOk7FSh8nwps9qS5dLuv6J1LlIHiepbdtdEszD9RY
keZ2jtiDlU92aeAm4nqUobgntNmgH6WjvgxtS80Nz3bAInkEW9sZ4Uq7qAyxgsWrPoKFIGoFu8Z/
D4x/clmSKxCgHmBeTMFgUaCDr1+AnpqauaIrDSV7/k9bd5vEHTdkVGzRXU7ozfQ460k/XEFc9fWZ
WX+aOVCRdhK0iIrXBVD7O5EdJ3Vg+UBKDs4WIstErR6BgcaGE3wGoQtT9ob7f9EJYsL1Ek/6z2kl
WhBrDKOZvGooIDcDdWvg6V2GIIW7IawVltvF5enBXILi8i0CsoWGtkNN4hE+AygLkz0XUsNM8Rm1
M98aMDqujisVq41HsJiGy1IMeAHFVaj2GnL01BFNtOfrtg3PMqXkzhyXNd47+SK5lVxZExdBZe7b
lGI3nBIWnW1v1aEiHetkDaryuA/uw4upqg06Som9qjvcsrHtufINCKTXnO8j8di8eh3TCpt4yjkf
Z7geRTPlo1qNe8bfx9mgXjHLRvCEGEmcfx3ShufHrr6QGZ2FTWeLKVzZ3bU0Cww6C+dJRGxJNQxW
Zy/j5bBiVqV16aHI/V4behhLc0L2sb4diQVlPPJSadfVcjjUSX7/QcOM8JisAsUdArD6dKBMszms
M8kzQl4V5Lypfp23N/x/PzZ6zXVclalhIX0xYKFBjrqCKx+TOQ5cG9cxy7Cqt62IPBDZqXqWVNj/
BQ6Is7FNYFNJaAmrZFBwzGK7kn7LqQ3HwbOhefVFMy3V/TQnyynhR45yxizmABhooBEh6tAGJ02C
KRH0slywHXnLJy1ETbRWMPV/X5AcMSWzBmJ0CTQwbEfpzhhVrmOv5xYOPDs3sdylDcbR/14/YMWF
XFP78x7DwAEo7RlWdST0ZF3Uqc9hMr1KDAOJkpf9ZRLDw69PVCn/lwXyCQ3khJ/GcQ/iKmrpIY6W
QnmZuZ1iIo7nfUxwehPEVbJlWiDuliSV0xO4dYoHlUHmIWD2ywak409S/jJJPeD0A4udnslT/iu/
BO14EfSMyUZsSe6tBBk8hBZeKLHnMt2SuLZAJbODiaSzGoGv5TBxVJIgPxe7XiG1jcTLBYpm2LRg
Uns1wo4knKfLkkXJCesjAOuV52fD7LwMuZsQE9e1AQ9j7cRj1aTC5onr65aAbUgmBYzwN3xpWkVx
EmLXuVX3vEg1wiwrp/T4bqtOv0xB/3tszq+EQxu6SbWqgaLJBi6NdFzkNxSXi+PK0ADheBFdplLJ
ZTnWkHLTdI9rDorMQu5njK456OuhXXiGzNNzi2lpu1EwxW8cFgkexmlypgZ87bJ7buvJvbV1aMP8
B4SdqzyrL/122oz9ol/55hIC1G3MN5fUnWv67SKDYstbOAY4GKa8ltlkagbWEQ8H3nj+nGGatRiG
YVi/usHjJuWDU0zlXUilCIz18UuxTwtlJ4cBeI4XdgcGzDClxRUYl9RcixT32kfj4NCmY5l2QiaW
U+8g2g8DJZnaTtvj95NVhsXJX3MY98gzzpkPtfOmRl88oAn6v8lpz+/QofgzFhE4e9NVDGOFl54r
Z7QXoLj4WlyJiar0boK4y8e3KVk/4G8FIpq2YWTcoOEyLvalkYb8swg9HNYOayCWr+6vRwEpqFyu
YllqcdWO+xFFDwMUsqAsmYhfP8jBdJ54s7OYEDdshTZ5CNqUs70Ha2Nxxc03/ApmKggwjmjd7Yoo
/uIZsEhjcUuH0Am+nD+fVFzQOqpnHcJaByQNKoRhhfvJtCPwXwOpDUmX8iIZ7X+9dLpwgDWiQs/k
xc4w2f3/dGepjyohRriimRacWdjmlGHHGgO4KZvH7NozE2JJV0lg5Kvfj2CUcW+T29w61O1Dbsx7
e/UZEque5TfgP7uTNlrpiTKLFoW4jRqV3ygqxwxNe00wae7i9I21bd/HtYQbSWKAAXQj9iz+496a
bE3yjs1SUbdLC29a0XMG8a3U3p18Idu4PS63fWzvqm4VqyOZ6YCnJO0Bq0T8LaI/LWnXz3ezhqV6
nMDw+PRJ7+I557LvqUVlUZqGiMi4kmjkvN0xc8om2fwt8ANCKUGTB4MgzWhRZi4MKfcyhp1ezsxk
NmqE3vBKNYYmohlzY5ZtDRNzfnzfovEOlDRPXTgHQEUQH+xmXd53iITOWIliXAqZ9ljM219bDPbG
4pIDN7UOIHTiaUspIot6rxNI9NVcdGdVL4+HI39KYzGOT2IpOFMAaWs7XN2Y1UeiVkNfPTKqZrZn
nQ3Y6uhD6I7C++l68Itnevfw6nKVhUAWyVYaguSV88drnmEgLN404Cj2lhT1fSeXkw+RDuBb9WqK
JzvpQYxXfZVbklv4RohJ9fFddz7426/28H0dd2itklLSx0W2VvqZJu/nH6CZlFkli4ltBB7mp8s7
wPBRh7wP5aeduR8dRLZzPjQGleipX8VE6EKq/6m+G6OZt9DKZvL97GKlYK6UXRSlHePzJ/WHLHd/
iURdWV9ZqSjgr6bDdgv5hMVmDz0hCOijvaUEKI4cqLYWMcwXauudLQ99lRkOWjwpQL3rWWJh99uY
3Ww3csZ2774R+Z3odabNbhm/ZvKfETOpH6G2BaPSmQbE3tQrlctnxMgxGmsrHPS3TVzSnLuTTTn6
esGr19UvBa6k10JHvv4E77t4sr4pJyz2akNax8jBnHXvDIFt6XG9kzoSKdNgRHLQ+b641rm1Gveb
wSYiB3fwFf8xuXG8hOYTTvUwZPQj5p4lYQIYmXn7+qY+E8g3x/SRh0st0js4Bc8xk1q3wZB3hVii
9ShkgOCXYCIhYsQZNrQKrTYRA0hIAyiHZzYa77YM0g7pTtsNEFxm61DH6ea+4alQF43hyUWV133d
WCBb69cJG0saU3m+WTmnlrgx+85RJoCfOFWf++Sp1vrA2trT03+ygxQgUS0urhyyRKYHYFYGOimZ
O3iUDcL1jJKB0gOh7unTwm1wzgqaLXt2gw2Cf/VDCgppuRMYx20cmcJUCw+1rIniGEe99345571m
tSWwYILj+O4A285WJUX/IkqTHxIm7SlGeioVnGAMIB2NQwtmTZbm3/GpE6cEE085u8GZFI6Y3phv
iEAMj29ilTusUO6qi6NFx40xIRYJT2/XlR9CZOoFFHGaX5GShoH3qRZic/Yq0r1+ONcJz/meni0A
ZfSB5p0uLe8nGh2aPlvoTkc/4aNzsagcezeKHgj0R8pE3enkSPxsKIXhEY/7HhhzH837R3vVKb/m
DqI1Y758q8ElRJyW+dhxT3vLUNWSvVVSgAeA6u2qd8aFDJNuMS1RouE7n7o/y3lN1qEnFODPYDBC
dgkeK+z+O9gIqjMM+zJ0DZOq52jYBUfnTfeB44EKjv4OJ4dyGwdBZzb5fC06igAVDsnB7YTwQB1l
jzOuVwVmAsdH0hhpDnZqX5gFCk+JMbpsNDcnaivERywESR/Cr1jyUeEGCh3O93S5WhzBjnbwvnzc
UShoTHjSjYvJB2R1JjJUHv5U+IdFkEHLHYzBu1WVLMU1QBvQr83viU/rLeYc3vtV+zxa7R8cotII
jMOCNXLEZDnD2ae37Bow7YFdr/8dC1i9LgqQLGPsDX42eo7UIOL3P2KJkwVsDfOOL84vHUSw6iAo
l8/9kFxnn/aH/j+2XsIhfCa70wcOuQIfFsS0L9lcjcWL5oabzlfT11FOEE7Qkz+0cwAZA/uUs7kk
AuA09ZA8vo8OafaPYDPcOIamVHnLJKPAdbzsAO2Rkz7Rg69OJQgINVbSmOJmydiwrW0udsHoN514
P3VRm3ybV+PjhyjApLw8lwoLCxjTz9qA7ypL0XSplgfPA9ldOOkGYNyHc4ztPy+UjaSNqDBFZ9sJ
5FD0dvLnpZ4ZUIX8CtVuL9Lbn364C5q4kq3UeNz+FQCUb0Fpv/C+QDSDFYp3fa30eVzFqoQmRFgz
FeZYh4e8Kk26Lbxjm/5h+k+3QnHMr5YoPdWV4sTIFLIFmjsOCpz839xRA6jOHKv5WKlwPomGtSHf
9tlTNibHaZxhhi+pZstOlx6DCCgy82fuwP6hcGfd8VU+49vLFAebpbmHzacv/4SCRLFQ+0amkH7q
0EgXNT2Q2kjttfG4TQGpA9dvh8+8vHLC0Z7V8jTxE8Ce5uYnFdD8TgHB+Zu97N2CreKUIhkoUxnl
Ds8aY1n0UVugwNY1ItbzGlogYdpGw8RPVjyU0IbFhXVyE3KCn+p9UEGahBLpv2TqTJRzhEDOx3NL
4nDCIeUd5AQ2swFYB+Isk45mulgUZcqRZ+iv6JnmXdndARkAjjq9TfLYUk+l/jcYQgwo4aDE2TZj
2o9vB4DCqibrJjTrzeDJiTJrYATriBeugBLYglhhZ7tbE4Iz+lshTq82WaoOcJMXDKfktK3oGWcL
iqh2ytMS5EQfsBwNHhE8akIYk6qfq5ye6tuWFrmLRR/TSGNLlfPb6pHXNoTZX3K4Sx8jndSnp+nz
a+aJyp4gPns6Hc3S/2vpQ5sSlbtH5NZTkcMYFcigi4sFg8dpbwFNDEFxg3MOUsWylVUy9oJY4r6x
jkGAPdQAtqsNTwWI56w67E1UqfQrrKRuoqoX9FEOqA2fGozcpK0Y4tJwh9WteoGyTSTSGR+CSRVW
O7aYTUJh0ugUx1K2/8aNlfsoGZWapIaJ8uFLQ3mXEQ4NLdld0E/mcIk1uibTY8Gt6gwN2UouAoty
3LjpRupyZGw0YzuSAIRtgKPtcTiIKcV6I6/O9zgmNmcBTZ8OTEQb8sDqcxHpeXq8DsTl70Qfz+bZ
1ZKTPp659IU0Q+SF9+4rAMNlPecCGcPhb5gZqTkEoR9qQRPZXR5P0aBhYYskJvaR7juKc7FRrMGV
QYLBIPrLFqBG9JmRBcsVumxG/Kcaj0He0iR/C/QSueLuFjdoFSi2Vq5pLnGEyl/BVUJjvQqRdkpb
Ls56Th981bebdwY0wAsiuWWJp1rcUi7WwD1ho6Udn+g69tn9PSglVHK8A2ksP1lOiEWesYjb4bWM
gXkCjrUAte9zGnrzDnkDsS0XGxk1r3Egw/euCX8h/9Ait6djGdRYgax0mfRCpi2TZyoJBnJdgN7m
tdiEggNl7hNpQ/h0dUE7dXHra6TjqqkA7witNlXI1H+oa3JYcGNLXgoX9sO6n5HVx9CpJd29c4mS
phqGEiHmx6ErammzN06YdZew/ysqhxoXAjJhSLtG5NzBSRQJO2XN5waAuBP9cA5eLiPRu/yiDmmu
qheJlIsXlbi0rj7pIHjybqRGlgJaK24W665U/J4nZ7kfIpDfwpJ/YNliXu3GKdvIA3X+Mq4bPqn2
U6rp2zn7T27ktxqNvyONj1P3v8Um8ahcF2ZxRQBYdDOoHWAxAfhF75Bos4aci6VKhJ5+ak4FRxkC
Hz6IQreYYAEDPCqmkGxvVCELAILFnwqzvQ99Pu41svC8tWYwO8TtwXSp9nUWEPwcV4+WknZ87Wed
QwnASp9aL8OgnQk6gAjju9lR+Jv/ixDblX+NY03oY074j2LrCJ+klki1w1RL1AkKobMAVtakibGp
y6wvgCnX9hCcq4WB636fY96j/YrLunTRyaBm55UxAC/Te25Yt9aVTCv/g8odLEnz0tOPETZHKr9Q
yh8svJio4/cY5AGXxt/DI6jeub3ZKYtuqErQGUZH0q6a61bnDcPdILxtjoSel/jiBMMV7rtoGtKv
NnCM4k38LdCdM+YL5MiDecugmmInZltaw3quwOR7/xnDWxMupZrvUVQsiWwhj+V5n7PbI2ZAKTXs
gZ75FPF2V2QR6qXT7GWbHLk1hhLC9e8eMM91BYh3cjrfRXuCM/4oDQL/86ZP9n7HJoSBfpQ4amat
WSVuOmttePkDPt3jGNvUVVErJGHALND+xHOwv6MpWrKnJxfp5ZQy2wlXTbcnJZ9E+ojJnw5eDdOU
U0HQHoMg3GcQs/iGHKgy8A4jzfVbm8He68V/EqMmTDTXqZVA+h36Av3kYfSy8kVotbnZY+rLx4zD
Z6+H0WfSjMKjHq/w9WIIASlW9/zJVpMozn8CMJX41J57yU10xJJQMnQ/d86Cxzg59ZakqWobGR03
DqkJ1l/tHabhTOFRtmT58561GL+bz3hIaQFST5BPItl/11y0h5xg4KrXZuV2Lo/npFwqG5Kfrfz7
F+ErQp/uGGSXcF/bf63m05ldFCpWHHhclYBT9E9oNHuc3N1lpjfCrVwqmUyrzHF6CHrdRqv+/p8A
ZSMSVBjq6JUU1p/RPeD3FW/ZEnmWmQUr0rpBcr3Q566CPqmlPuHdtC3k2IffWg5HTRd09aa9SDnb
tkfoau30/GjfDM2WpJz0PJ2BRPtuEaHmATjdqZnu2LXAsr5+0kedOQEZqMSqaozI38iB4ZqICb39
l5qD24vmFd1Xvy5UgRnHo7NY3/Riit3zvII6Htx1huX8OCfGe5i88fEHa8RUDiEejGl6vhhb67Hc
tkYDb7ST1BnYD878JfcXZs6ymnU1cBXemP0DLrT8y27FiBZvJqVEurWGunCJqqg5DVzcuFvh037J
YDCVoJ48PGEYMZ0TV4z1gjQVrv7Ln3/HNa47oe2lcgySonFn2ewoR2j0/sUZOnkmgYgXvuvlIBcP
rD4vGdC4R68MNpzbHmnwn2KfrnuxJ3890LC+EkNTvd2ciGuj8NFfJEn0ibE8Xcb6im6dKJJFgwDH
9l70+pB2917JnGA7IrstIYk8CwerJnCHXeAn0Rdv76ADwyOnolcoMClY9PcqZN6TG/uMsPvireTl
zXR9o2KkuZccMvLW2/E7mYtdj4Hj6XXoax8R8qaCM39IcWK9GYyX1KDNh4RxJGTLtx5MueCnaTi9
J1xJKKl/peUs1C1DEBz6GCcrYw52YE6ah8IIV3YtB8LfzUC1yeewvgRFFcJSx2c0nJa57joElBCA
Hg8S2dXRY4CkC/tUNO2k6zid06xrBt8NVeJpJAE+dtGFujhUQe1QdC+KTPVCpYW9LfGEePjOi9j8
QZF+caQlaJc0WCem4W1JjW1u56GWWaB9Iv3YRpYbLthiUBFGD1ZEnlUt2RDfuB6L7BhsxFbSEY0S
NdPYx6RsDixxn288kekqHq910YVvFuqDQDm7zsgwGFd2zjHSSwUQvcw2zeE6Y4sLucBxvG3rXhCm
/S7Xw6CTvztMRDksqu/2ScUYYz4PJ1lrn+59K2MpJp6cA2lEEWkWZBa4aa9Cg5c6Jm5HUcnSHtgj
zMEmDPgV0q4+yaqhpg7uupm1noj2j9yJ8MWxALWEGf+pwrjGbc4VZvXekkKMwu7BssSG363wPtoJ
6tzyIvXxH/qH5UR8/OVL1NV74dSwfEs+2YgERh3ZP/VMHhQkyPx9733n6iQf+v+98aCioyli7O9I
uPbbjdIBC0M/8uyyL2C/FLyxQPlXJHq5zJ1DVrdWWUamWlgmwgzckoNBIMZNncFq863PVe4dmrmW
Eyc03uPNf+vKxkgHQTJsahIr+VKuMCioLETeVbzULVOPC/Thq3ycoCj9i1oo3ix6icYd/HTHahZ4
azJicZbLHoxyF9KtzrJo0024KPCKcdLdSDUA3f3orNg5l8UAy+xlsLoq6MH+Me2UHxX8yunB1YpO
4DOXUrFwChzn2Gpck+/OEU23JMTjHgZ1Cy73jb4VrEURmnI775tTc1UvXtYtlsdGHFo1tuPuTFsj
uvtWFlhd7GObzbwi9mZ2bgGT7pHdib8ZjuMasSt01odO4IExr2Dzk6crkaHJbHu/6LK1xCH0YxZ9
Foxjjha8+C1vAJZl1ObgkEEDpdC8l+hQ+6zcdfuiJcNDwsfgL+U4PZTq6Ilgat3oV4X9t7lJIrE/
Zy5WWW0D5hIYJIxaBs8zFbzTwL2CKe95jS20fbFrgRBSsUAAtOF9XLyUFQSPQmEb1om8+yniQBcd
o22fUAVIBppH6TnDZMBmxrvpOH+q0HbxYhjLcMedksr6Y3K12OA5+YRRXms45JtvmdWha4xUh9zC
NIT6SKw51OcrXb7nWiTVXUg23cgMyZYFe2d79Vw1hw/lCO/ZK2yb7eZuurXj9eqqH+vGOI7x547q
LtVpRBobUxnzu95Brqpf1U80BOZb5s7aJ+NTAQnraV9o+qLgcU7PLphzyRnkjimxwraN6r4zjxFc
rzpXBcPvGdv4bxKpYrcXD6B7cjRUrpzOGgtXnNxuRCo5Sn3BkgVM08haA9D++TQzikCe0E2eCrU4
+CZVRQZDkOHbfqzuMzPKb4cwbZFoI9+eeIpiEckKQzpfbxgSDBiZAdjqiu2UTdN5i8ji7G3uJHph
0QcGbZCkqpDgokDu1wymW+vlwVdRuJakbx2Gdo0fGMqn6Rw/zL8I+5FXuASrFZoy+Uwpcq/SeYJ1
9ybDEKjQu1e8HiyOv5IK0zfg7+29ZENyyt1LbcC6yWpA+xqF2/Ej1HLkSxHUOSpAReEmLaoXewzm
zQlWMVLMfM0lpxy190Cr4q4ScrCkpfVyX8EEtTSrJ6AXcr4dA7IhFpiuMLrjYQc72SIitKSuaQcH
cbm7naESen/IrU4SyfiKsooQURYB1w2bVGF6sq7aQA5yoV6Irk+BZfvaNGK70p5E6481pYHW9Isr
sOocbp7pfTzUCYBDZnPdla4Oc2zq0N2RR2hOmYIXyBtM1FqT3ZebuzmDM2cxpe0DhLLKIqBXnaK9
G+y1TM7/i+RQ2lBICZd2A1fOaP28kHjhnVwyH2Scu6veGw9LKNFTD2h9Tv7AR13FlKymWFTq3GZg
xDh3/kvkO2Lhs0Ox4LSsO2Q9nGOL4kZftKokHK7QCi8PQna0mGxac0NM/V2rsvsfKSY+NedAsfe5
Cpwb69MN3yvJxNukUBBx9JY8My/2XaFHWCDKZbEUYV2euf6IE5CDL87EIdTMLBsCasz1ZiMmWTWI
3+4oYtzitGjmdixjyq5gR+B++AjEdniNbEvbbyNMw12nmBJ6fWiVaig8cvXN7bhaHWqYflrIPtN7
A5a3VIDsSMjgfEy9e0OS6CX/4pB1c4Pz0pWLkU0GrlpTxrd285X7gbFxcS7oQ2cU7HPzQ9HXSbZ9
SiNaf29Oik6twaCk9NQRPrAyUB259RpYtjGwFN7+9wh/TzZAFoMbIotuYlVfzsltD7OapXIJ/Yf4
UNY8QWK/cnnuPHeoLdUDjGQKUdgmK+r/VmfO7qLtC/s53XyThVe23DNFsuL/pWbv/opksMgfjNdW
Uf/TKg0Pxpl3XcyH5H68iGqfazYgbHqfF5fwj+euND3cpnH0GxYgdiVjEW239MPiqRtA2jNF+CL1
k5i3+rG5KPlBW9QZbsg3rudY19OAPCXmFB1sd6/00YCBQwOre2lxuWi52NMh+zdYF2Qod+KjXRdw
yoX6IAxvBKkiwUsc70imD7TE9qJe2P8AKR7nDjuek8Ls3hIZjRYyVXMVJw94WOMtovZ4e7Ij7W+9
g5dS9QVZd5Nrca/djcQywLSj1X2kqFyLAnB3k84i1Zj1Ci2JsTkt+oqm3LUGDXWq4NojhblNRaoa
M5LAPMhIxB5ZdIEOwNRUGGDlSJ0S77iVSIouawMJNerDSKIvB8tt/6TP/7jv+iC87JsyA9ovE3CN
EDSMQZjCKYVzF5IaOptptlfCKywHPXTVAtvpGzU2hmgm/NPpDXllArmJwgAksGXQaG5LTplcDS4L
iyULRFnNBLHC9iZsRNQEcDHqkHpejXRXSPsK7KVI3stppTgTTymB+WL5zanavnc7jzdbNdGfIdqk
3w5c9MczHcVxgrJRGSE2QcgdAPDovztmBby24+ezwV77nYJZCUAGx4hwtIwMo2TWZicd+hIyNm8R
BlAcUEAmTx32QwzaCGUJ72QxEj5Z2Z77XqDPe+jG6jfgeEHmLGrgALNFLjqjjAdFUPimKTBNUs2W
dlREcUbX2y9lNvlVXTy4Cle6QqcCHqQHEAuGIjouUqrFVE3T2NZbvR6LXNMkZfbsweoooywNl5ge
lVN7tfQyA2CKNnUIIO83YtBbgz2NgDWOL12IqxHRhIiJX5EhkbwaV0mwba48yGsEPJFNxtM293dM
fZ7OvpBBQpc1kH5yt1u+VqaFoCA1LWNlMTYnAD2HdkvCD+pP/AHm5IwJssMpzpI9Z5GZ9Di/QKNA
fZfqNKMT6RN68Z8IVK/BfmMZdpaa6wJAhiMrLr7xoZFgg/O22qPQk9N7Wbh+emDJRO3lf21DwKYb
7WQmw6PQj8V+dDF0A6iEj2dChAfFwzf5QZyiCTYwDAATq4187vMeohPYlT4LUrZVBc2Cm9CcYgjg
RglMxpyDTDmmutGGzm6ZIxqLnGcSpeCwYL2DdI0JutxtE9nuiulOmCbMnX6hkJee87Q6VdW74TIF
/4zHjsKQgHnfNmDmTWVI+b+ZG5/bQEY3MTxeGmMR1Ky3hL6KOpW1OTMX0pNlFv+llJYyF4YEzp6c
dUM6nQXjESzFVTlnQYtkx0/SRY5HNheOlRysxv+G/S1eshG1IZINBwKTJXIpDdkc5EadIV9kfeH6
CHJvkg5hULQUWohUBHUVhzs3PRa/9hMM/A0MKxf2vUGsV15/G+gzpzvMbM5AQEuum5+Z02PIWeYO
yKPSQ1xTu8gx9fxQ0nTuPIdIgOOlezfSMqgZ5KYoEzPJjS7Tyomq66IcnFp4IwBsA4UcnfrMFvEN
eqD3npyaMk8l0OyGqLh+qt5uWI7bogFAQZ9idChQ+8OO4NsJY1XSHkC6x0eW6X5LAiSsSNPwkPK4
CuZOGVkSkjiw4QlgoMt3HvrO4BTAuPXOb5Ch6PF4w8RyYoMeEQjck2ufSakWeNCnKQdiyt4ELJOj
FdR/6UHsmAkqnfTeu/J+xkwSb7m0i1crTrAOWfmU66tx8C0Y2GMWiUo2oxbCA5w5rETXy8zVbicW
ee2uqkAILkTlLOFb1SyPLMIlRMo0/9hgxCp+Prh9dWOPmbaJlhTJ36qoWgWhW6h9hiSSKDicY+yD
XpLhxov6cZKcdTnGGSV4cphwaZ6O3WcBWIDuZBmghicW7WbvlpJ8r+f6/M+lZfVd7VsfbbPy0pjB
Tl6kKpcrkfWZFfAsslHc87Ero7Dt6XZh551Ss4ynJrrrFZFjVNyU03bwqs4CeVdvm/cMAMaM5XDd
RJlECZHPwSkMXOJovY7LW/vubr6BAP8cuIxSngz9ZFuTpelDPDNn2kYkTpZ4CX7l7Crx0EKCX2tu
V/kpRueucTkqiGDALN9y/2Gf77jQDZqT44C4/aR+dEX3hz9A3uk7MXVhtha7ZSiQhxv6Ckr+vawZ
4T9pWliCgPeXvtABgh93jLom759cCTjTgWWDZq9z7iGFEs94S2Cb4Mp5K5r6TBeoO2BUH3xYPydU
ju5Su/6TnIoMZT4Kl+IUbq1VlHutvEX2Yx+Fx5LFq6xImeiFsNl8cAU0bs9lSIpliGSBBIYP6Bx7
8RNLm1qloWWVwvohG1r5xNggPkagv4NPKtsYTOSqMC028TddawxilwOGTkgf/pw560VQZDexm6JV
9mr2VTd6LXLx+ZL6YFN4WTwbvjPkr1tWz2UtJlN74ClDNZBHu6COHOGhneE+jxfbdQfUTi8+DB6O
N2ilenrPRkcACeAn9dAkXzcnqEQwYRzd6NlzSKVrLglNWroJ6I7sSDY3xvVYALRuFKPH4dte12NP
sOFrR6fRiHqLAAZFxqnz+s0ZPg7z1oxHtPcthEw1mECbMOZzEyvSwM30lu0YgZkvOTd2HGSOtupo
QrKxG56Sn4mtwlgZEXRPk7J5R+azXhX4Fi/t6t8HEPQe+KzB+RJ01tZgj++Izf8AK6illwEkyd5Z
+cDDXDFr8/baonRsWLVV1h+0yFvksbx4cLIyZCpQITmcn2/UsD2haqWvlYSj1H/Pe7KHDQXIuJl9
BiQHGVW4/5QClG+uU8hapVVry1N7zEc7sFLrV33yx7Xwu+nLqYPSPh0Vnl44VNZ8QBbuiUhcapYT
2x4bFurhdpwil4On3wLpfF2XhgnF3+9v+5+EuDSkUNcAfzmCqpWeYhnftz5EveZVF1+KDwVp8z0v
PVgetgVIE7m/NHiul5be2WIw5NPrWm6QGl6RFbW0TDrx418ghtao6tm66VJf1Iw1KkHHD0PDMJGs
qlgm9Qct0l5zLDgiVbkmfN4wZMwEPUmJvVoe8nbexNO/t5Z4pXDV+A7bNRAhiV8bPi+3IDJLmXDe
ieSSLIiDuktfxzj6HiLevsA8FFS4H5O/sF0yfvDiJ/KW72LDKU12IHD+w7FKyQPd0S5yxBsVk+36
LzkVT3VkMl/ob4aYjsIAKtwTLIN6nmXFnkWwXzijRG/nUyCbWztaJQn0yunFk+uj2iZnCc4rXJjC
hW87ZeJo73bZi1tLDbS71atXNdAHQm/qaXr6NQM/R/okDgHmlnVnAppkWLXwepcQaEuMjHoc9tfn
3UGzRAZN5aurIbHQVJWR7qYXCeFtmP/rxLu10Ym/jvvC27TxDxnsd6ZWTWSEV1qYkPBC7khJNygD
7JzAUlADJlSJvCpKiHeW+oAviy5760HQSx3r6I+mx1hrxRpsbgjlcB5Bhz3w/pErrkG5jhZb7TSV
mSIfnLoXBRpzJ7L9X653tirEKZgakB7CLxpMRpBcgTzf1jR2e0xIIOwEx9pc2KTr+1/66KFwHAfF
wVigyyteTQxz9J91XOyMvhz3NvpTA+RZqeCAtqX3637ek8UbMSH1hT9EvemuRSA7G+hoppzEhFbg
fWEymgXNmeq3YvAHQgCzfsJXcF19+tLA4Vk+UQnQzFbBjKprS37cJNFrck34zIy9ZaIqwShB3rFl
Ng/IHvtP5I++ei8a+ksLxSBsB2HB1tWpzyNPRq3XYCsq8gkmgxns3Aup27mOZob/Blut0mx5aVB0
/IX0LAoLWN4/rpMNWWvzftRW8bEL7/iEZLgxl8OpnLH36MiMK71KXLdmC0qZ391dF3IhDF5zhGvh
EWaxaFVAcZE+FyyKTzWFaHx1Z0CVlAo+A/ppftAS2dpByNzHWlsNXTpCBMof0SzWaaUElISjDIhV
e/B1ssZeJZhnuYsbbnp/QSDFhwSY3ruP09Tkg6v8T8kjdEN97/6/gc2zECvckLnYfm8ibx5XRLZ2
3uXJkxw6Ct6lLJ5ZrBZTgJq4WApbBOeOiXrkkyp3PwjlDWhF9YnrV+SpeeTLsmADmRDb+h90AFQR
a07Mouf2vvy743YesV1bXTArRtkQe1EIt5tsk6UoTOG0tSewKJhZ5FxfVrQwdCEQGYb2YKALGW/A
9tIQKFhWpO/6ZZyRFX628vnleLJXlaeBy89VaPr0tvU68Z2ocVzCmFCGeLzcKMkaAbQfGne3KSDS
XS6iIrnpd+91vOkC8e4EoLtM21+yI9a/tXDS6K0YUk9iRSntPNyon9pplS0dinQrFqnQYkH6VacF
kcbF6SkwqHjNgau5rtS5Y25cOFOBatzqyx4ZzF513513+lK6VxPd5jd7d2SUoTotAVKNj5F6LjSj
/O/z3VJQIoJxAm5++cYczYaExbsH+xD8ji7m9fBGq3Tlt2BzbpIvuCsMqr6cg2/yr3TRqK23AR08
V/yxaciQy+2g37EL7tuc/Lw9Dvv5nC7nxTvqjBo6VXmmmkqn6KRSDyjPx6WjQDCsn5nVZBPuy2Oh
uQS4oXhHsseY9KIS0/td9AScGnRk9fo8Hmb4cNa4WZ5EE4femwF+ebMU98pXXtB2mvqLuOzc//gN
XsYAb00AIaM55UJ+qZBpv3tV3seU86xdEsqVerhsmlnM8UKLpSduNLemKMv8LhOmU1T0YUeXbfuv
SMkm030NF2MQVMh/p06+B3DBiRZBsdlYfRs3DKD8+nnHUNRMSQVx7NpDcaOl8FbecbZr8k4F0GYK
ops+bR6M3kJLaLfYMhfQt0RntOGpE01GmdpeW4drzg8aKaYQVN2vlrMB8Jw/mFBnQYQs9Dm+9I4i
+Z6NnQ2nZMAz81w2Li+x4y+VEMRZ9J0yB/iDtUBg4Y1gmfBqWu7yOV6Gb2y5TVHQzTXWHZ1cWTWA
MnTIKZHVn5Jf6z47sRrjIM7wyX1VFoKlINsKgZSBwNzygL3lZyU4LFsp78RYAwHN3uQ6XDna5jtl
4XrmuYPR3mPsBdM9hpLLVLaTygZbvdDlnAJpcOFGDv2GT+p6igSrisPmPx6uP0AJ7Oe+WyhtIip6
OwHe65aPAExon8QU2TdstvJGYaBqBQ5Jb+GxYEMuOs7zsV6yRY6pc45gAbZ7s668YfKroDWqwbUK
oOhm506XHEbZIwbSTr0kU+0u/xNtopgrbUsJGDgVSwXDTHUW8VBO+B7Q6NaBPAGc/u7ELbQiYfG8
RrhrZsBDdBtLYxt1jHyLFF5UI0IEiSvQ+UTSZBRTa/3XFP71ZYkR1zLtBkNIHpijq0je1DPEXIL9
E+vGEg0zL5lz6vXVB7fL790/wg/xT0JxNWGZPlhvAA5bxVrTmibo8Moemasci5S5SbTPe2nm6c24
ePP3sOoVFMBwwx/bF1vsSXNQaKGl27anMojiW/ocJIZsbSqbVhgPSfvMm5eiWuO7WDqpbTDgUHdw
ki5OK63vtJo5qKJVtU4FibUJvdXOYbrYW2tu8lt/7s7HVv1OhnlC71HAXI6fmsiTH/ZZGuHbnaVk
qXRTk3iwRFp956ShMvpNxAjpKh31oeRf1Oma2aLm5zO0tLw0tspUGtjVlEOzZ1MwFrM3MFgzN4bS
liMVl95O5XZ4s3gVJvX+FaB2bvAX1s3TjRKpK05T3S4NcK3BeD9XbEE9F7Kn1gs4XuN/ILEqV1jI
5gls1Tm0uvKmFIxtcUhiD2CB9A4nRyUpEmoZsG4Jx/bJvcDUXhjZ0vNz/MGZ0hSGzQZWyUDHayIm
tMV7DAZFvu6tjQXqoiPtdlI5TqRTAVe3s6xB1W4/aFOECxWSS8bKwQvxV0Bp5fKSRrCqUUP0UIOj
OMaX9uVzYQbu6RBvXWE0VUzpQgHoJSAN7ymuBDbUvYAeVdG1hAfO07S3ehOwEycdmBQ1NzNrMMPl
lyBxg4ksZXUNyMAL5b2c6VOIPJooZ93Fji42OfxqDU+QMDr4+BRm3791cm1NFHzs9ypHyDwqsKIR
W2nVvwsqA8mCX2M6uo5dOdWtPbRFxAD0S8x+pLJhN7pdMkyVZOuNdOaExxhXTsPeYFE4Pbblv3Xk
fp0pK0QBsdoNomi18b14RqFoZuLTvYnur8himqW0NvvHJu9QNLBQVEQHguB4ee2Sat/OJIQWfySt
Oe6zQaQnn1hwVA5pMmEnrkolSntt322+RSmfZD1FT726HHrDgP2+0hsaBhA+elD4rtUPRGlGW43Y
Fnetr0MUCN2lP5Vt4M8ENVzcmpdKVufinPL6dFugxdhQoOrR8UXUOQCphA2+0l5pI/yGeVDmh4OS
016H0cUlUpozVSSl3+QqBesY6z4GgQRclDWAb/un1s0X10/O2gl5aUqW8A45ggEJKl581Q3YRs2f
qKajC2yf2eYeJdzUTn4FLiuzc4dMW4zdpEvHFFlnL46G+6NojewAXEwiMirE1cRc1hO0ADfwPA4S
weA1FuT5h3x5t2uicIa4Ea0pFB4SJACAXQKLcS735RCEAZ+5WW3pHBNmVWwHauMjfrrPyliapQrq
qYG7iss4Zokz/zydBsKG+QDFM5IK9aJn/Et5Bfa4rZRBIlXj3Ir3UnqZ2RD0HtTbkEEw1SZpR8P1
8CDGX0iUK7Vm9PQhuiOqUgwurgdBJu/eyXLkgukwioCCiW6pzZQz8zUJaB9lYsSdzorkkBiQyAm3
hzdZ9lewtTvoSnB4BfFh85bgi41Ng2A3v1ulTtu8FEEYLPdQbPeQS5PIELJWQritEacuL/ib3iTc
8PjmMif9HhTmqSjXd6ms5HafMQfhvU/FIwv8hh8jbToUSJpo/GFFJdqjgElRmA4YQBdd0tM6kHxZ
3JnP7tBSphXdCaVDidIouXEYrZEh3RPIACdXt55w21B6kTeJqsVR/6K7TuUG5arAkfV9ORYK3pLn
fdViIsIAIeNea/1Ib9Uv38BmqvO2Cf5/F6WI1v+kKUTDwtexz8hF5miAf1Do/HGOKxsKeu6G07AF
BwP1N/eEmlslxtX3wLdUobbH/NeMx93i+hbsySS/RXbk/NEwX06NZVGGdRFlNhTna2iLrJOL2qW9
5dW8syrKCuFe/0jnV4SoXbuDgqa96TonuwpAji5b5+VWPdyFcyfbV1J7MG7FWEL7raJOKLwlv1od
4bvSjATKnipLOoV31cMJ1wcVyZZp0kQDzpBAlbzkbknCRYZ46GVpQsLWjFukr7Eh8vGwsVCsaVyN
4Sh988tcTU+q9/WspH9TsGlzBsgPuztat/xvZf8fVhUZhXSDoqUpKxXeO9Iwyne5bkpeorEQQBd6
CiWZe0faJwrSJE3+TBRadRcNRIpG93GbRLxhuLgKB8QgR8CExu2zOUohxD4wz3athfs3W4/USPVA
mH0Z7e4K3dAWd7SOzoKY3rcSQzAxAMRsfrOEFgkK45isCZMr5PKPtDEnYzEo82y2VxCoCu/j8XfY
LDOdz4OL5qKOivb/HRoBBfLEhiHn73dl8+P2dKWYVjRuWRWhjh9hxURxiGaZOxE5tRDBqHgNzPPt
ovvzTVFpVw301WURfjHaEJm342QUiwu2v8+MgPfCC1HPC0xaifPBSL2kweb2FO6DzH5fAtBjfQ+O
1RHqL5fbZAI9miY+v8DoTD8q2lDlTi82DTifG87WVp9IlnJFCgAgk2SqFpNmvoJWAj0Zl9e/GnW3
1UXhHS36ir9BjBzodvhNV0lhAUvk5xYVgzPsGfNjPTiIa1cCr/T6QrSFNJetFPLnTszvkTxBtU7e
bovSHsgGJag7/c/nZvd5LjA2n9rp4zijfGlCL2HesMHjMKdHEbiFT4UAA1f1BWRfbTn+HDsdi1XD
xWUWwToJkkM7HGgPtzN+DfR11oRajf1wclB9iqpV2VCJf5twcENqKz+Vhrx9KRBtpFK6lNB3uxjo
PXya1I8KCrwNhH0bgBEB12Ai+vGykdnSZoa9b4bKwvzgfLYmCTL2DHcG6XMO3rVUKPb7pn7SV4va
RhROHs9YyU6Hk6oIfK7oGqFUEYsnt7CBxOb60d6julB1qxEoUKURhEsCkQ8McZaPVa04DrlDDDNX
qdpFqe9qtXa5WvJ7JCg91JfnW+1HY3KDVoFbfa7sdF2sdJOYyHyy2aAtQHfBU1BTGyFtnd45knMP
lfJQ4/ibpg/PR9+8s6rHn+V9Fy0d0DzFGpNglS3fhHhjV7y5crPw16NfFG8qyxgd0NCjG7mm3fRq
lERQGue9wvPsMqWZjWdUnqA2dlehKDJ5Xgtvdo7qQcAgTF2E74xsh9g7/jEvcf0IafzQBDKIQFrd
qN/Fn4TyNzaQLIo84fxzBjHOWQRvisjAIoDRKIkK5p4Q2veHbe11It2Kd5TeFGfsaMQvLYUR7cCk
C6vUXS4DmiAcHzLQkSq6OTHvwGpafmOMHcxomddiwE789ja9D95ZrD7csLqg9Qb3EZKmQ+aMWORA
wmDzA9Ed1nq7sai8msaZ/iZz3leCemZB6pywWjsWSsjYO1DmZw3SEaB3nNdsYC4TotCPzGyvwcY4
yMyZbCE2M/yO8CgY9TZnQY0ZkKTt+MIt9x5IvelkiwspNokVDlZaGhhXYZWglsTngnM0WEuIYeuq
bAH0mFivGSVoqkAj6mDbOQxBKxJB9K1yzJJ209tdot8X/tyXEX/sX2Wko2UrIpatY8AFqI89gqmu
WsYuxJKbSvjSDfO4kZI9dmxW15doK2oAr6fyW+LIq1FLVSBjYtQxrDenfxX+s/AdfYNW0MuUDQAB
nNZYGLLBZ49rQcakPJz6JiuD1w60p0XGok8GMe73a0mChL0wn46jrSboGsOtlASGN7WtAne4lwmx
sUIYj5n59x5Iz7XtZDTVaDLx2PwFwlVBf0Anrr8IGF831sjnq3NnEhSFI2M3oryfqaF5htZGiAkl
tKZy1tsnZ3PrsSMnVkZsyVTR9r63psaTIARWhyhEKhw99Xsq67Ll7mBipUvE8mTYvQovDVwEGHMR
V8RtBaao0HJIO11sErLmga+7pUco5ByuW6ZtkmGoH5beU57VDwfX2jB7CqUGqtFMWCaZ7kbXkZdw
OG0vmFfH/R6RXL8QyTQijm/+iigxyTOlR8LFAtSdpiPmGUamgQsIw/fAFwVItugdvI7WknPii+Tg
XfS655oAiVXA39/0gysCPeLOOBdy1DMPZ8kmvhAPCv1E/xWKFSou7KR7RO1eqsHgdAqU8lsp3YPx
853rb7oCscdszxIIxaZbxorBNKwIs6iajBmAUJsoJNqqK9vBCcNYLkxN4hbjdzSxNNRFm8/7hvXE
wrqrxXEKXpyFAO/YgZgEncs3zJ1GjfPX/CzXWgUewlZ8Y79JbjWz9C5zH/6tBJE6R3b0JcHZNHDx
7gJf3AZMFlfvp+McMvwoP7WgCttZKiJokBwRpYEjku6s5GeE/YruWq+Qjgla1BtfbKGymA+S9Ss4
PNLXaczcRC7MkdcVsx48RQ/mzie3ebsnUjk+vv03whbJYkzY0dqEObAtH9bVi+MuzJG5ZYcxoWef
4E4EYWJ1WorOnp37hfq7TObK1NNSsMe7hm911m69IO6vqGLh5BsKgOAt2CGyWCcRjtp+2DPYlHEP
LW2xeU9nqjJTo02OZuIQIO/1YFxTaxfoP0tZ3UnqcRU3T09jE7b9uxj1TOB6UNHYa4OoG0JJT+BP
48/ysWBS9x2LWeCw3lWvjgqX9cyrbOxX+SCNJKoc5URxsdZarn3JhxoX4r59M4PAMpAnZKyj1/7U
yhjcCgaq28LK9d2WcKC3QOI6H79lgDKWhtCxDmEPtSHB5uUhpP2DNaU/7oycso0/bu367wO/knUS
WcDQMAb8mAcN7hc97yEolcwp1yFVsDYAvrZz7Ex7xNCEanKEXPe9owrs+GwuH5NlbUjPjeIV28rw
l12t8xSDyowbC6WSQ3B2rIj9pV2ja9QI1FUQ6hUENboqEa5Qw5AXizX8FV1Ixb80KAOLzh1uGLs3
mF2J5VlMJZ2nds5C+/rzeCv9PwK9T+YqkkWmWrFh06Zl5IgeYr0uE/G2gf/Sy+Su4UetttBue9v9
OV6FcyBFmoz1DQzpxK/GDSAgHmP+NBJmMXYms4JSaLeDYW0Q3WE6zCbWK5Y8kMNs3naWPoDl09cP
cZv2rE2pWFicQhUNsfae99CAf7sMnCzmYcrxprcjxvkEgRFr+xkqc2Z/F66NutScHMmQAhNgGv5e
fuSue+J6P2Kei74QYDX+GhLcOU2H+ZCvdfHS1NqRqYdpKMAqR+nVLZvjYT2jBIUQdMKMcFMHdM74
6OL7DaKg4AJFLhJuwqHuksTDyzYAPPimHJlx0Iq6ktm7G/RdVmy9HL/uvgR9fdF9epyNQiOK6qvc
Op29mm/8z87d4pIxeZtdQd7EUeLU80Bv0jFjkpUOF7twaNv5QwDgpWFDI3edpKXg9WUBpo/KjcET
fcvve84B49oOzjQl+vGK5Afm3LQrreVncLEDhNTq1UFU9aW68oEHAhbDgq2ctq3NRklX2j1a3GEC
Y1tjJhy/jQVp225SCfZ6Bnve8PJAm+6FiIv7eg8vYj3/3R9gvq+nw5QOq7wGETlez9l9scWvb/SW
F7DOXIO4WbWO01gL8RAFJ935y98TeNZME4nW1fyxI5hldarvnFSsvd1LVWPyZsZxAZUQGbZi1bVa
Q5FMmnEYpXKn+Pz7qBie906cJFiLxZWOGpOE3JWk6i1hxc1OHWwWLuhYXDKWdWqEUSwt2f5Ad+ru
MI+EOCGkjOIKtvnkmuWsl7LcJOGrRPvMa6NH/Ag3rJZa4FcHng27ibsZ3rmeGzZ21vtcU8t2horN
o+i21vSYMEP+3HUjl2LE1afgKbO9AtnAZnkaoSljbEeGcJLmRoAlT6c/x6Jo5ixlLNRptdRt703F
OzZGOJvwa8F4J8LucDnG59wX67U75+G1hnFZyifSm7xTEWY/A8uj2bqtC5HEzXM0iJqfwwxzFhR5
1v+NWn+wu4Tk6kH7xLXoYyj8zNDMaoFPXuiR7PjObXKtYzhmvOajEHYc5a1wmdHa4BcE2IoRWlNV
ax7oXuKeDJW3SE1WuSZ3sTl9PVJfuMJcy0Lcbj5m7DN6bTOeWDGozNOQlbCFFLzjsZz4z13RM2y4
ONFalc6XOdVd4N858DNaeP1x2qKvKRiCoXOtFTrTdPn1fQuzcgu1ztku9ytLrm4amMBqI8skHaoL
8YzomafZDkS//ia7Exze2v6TOjIpBCwdCC3ep8ojHnoarv7ypd3AsB0JRUWtp0YTsvKGAwdd1FY6
sBwkiwS9U4Ct2+J/VT2nsVFnYZkrn15E/JvL4ze0lQk6ZY4JNPXN6iNXYTs56FUTlPH/W6e/NtZB
VKPGnkIRsjFmmicAjsW5wX4Wn7E4SLnqLrrZlrMOQ4dwmLzU76DmRHNlu9keeWwgTIyksy4jHm9Y
h47dr9tauKtlWtHwtayjJDlrK+YsolUygzfIhOXaYmUcepj0L96+zpUGDZjHNo+EYGnw4PA5oT2x
FwkrkbCYm098I44O4Oex9GnLMPvXzNGakfcug5s7EZcshbcL/HmqJkfZ2mH2w0PRJkiZkXVbpsjU
VO1pzdEm56XfIh/ZY9Z6qVA/84U8vtFThyqmrepyWuBvqbPS1fFM4RTV8DuH5QN7tbl6xA77vJIy
i+5ixf4w+4NayRnBi69hexSiX/PTClGp3xmr0t/Ewx+z0xI7rfL/z1xI0ZZwqEKUDIJLDMqHN0SW
WxLYb5Ho/zg26tJ+V36il2P9eyAnBQaxRRtI4i3a7SQHP1uh9OIL7i0Bxk7O8fwX+dgNS20m2bgQ
fLrd5DkSDtOm6CREP0bI+7s0CiE47KkcA+aoHZon7zLmLVfS9Z3UqNwM0WpGcM1xD/Q8m+8AlDwJ
vhhyVHRiNeqB8+Otu2Os8d1infBPDmNgE34hPrUgP9/xQNzXOnSAyw9PJZaFtID+SFgtLy6qOJxg
5hcUn+NBFqT93sJI6coTFhmrGs1z3obvjWTSr1sJ6ZutsUIXXcAKy786HASa2C4N1RdGvMw6ZXtZ
SmN+mzqknVSNpe/FEUpq4q+ebCveD7J7lOh7KDI4ARQ5yVm3QkoLLHoXMIVHevYyLjoHIJq4+NG/
7jWxNmV5q053cL9QM9UVzsfFCCvU+hH5ftDKA07r3GOLOdjjsX8mA03l0dmZZXOPQ/BX39difWpM
Bdu4MlOI+/5ww3nv/wl2MJaE+e8MEwGtiZ3VExfgYCYoDsVDJshOZlLMYQ2veOnwWEpudW+aORqp
WO/k2Vbq4zu6vMenBilvan3LIzS5I9rs9Pm++UT5OLfEpNFqEIzS0Rfb4QpUK3Jk18BRgC9id2nV
dZxPxlSEYct2xVn98tIAxE4fAMwZViWkS6BEn6oZfReYcMy1gUNBDeo8gs67F7IfGWGIPYhjW3d9
FhM29y6VnKNo14f3bcGCrdHxiIId4Vo4sjlNEB0FYT76HIBEzlkZExvtADn8zZV5fX5oedtOp/BW
KH0y5q+Aw3Rs8Q44TyVLY/spPePZx0gIvyemtRe4OldwvzgbHvl5RJYoJakUbkvXnso3ANnOYtUt
2ZB0bmgnWZbVSCCaK1H6/PTR2bgNsbTilpQAJz3MsNB4AjPoXbcnwwBHm4PaoIScOFAJmrSpIhSf
a3Z/hvG4ycRJr8HFewwYplMoAdkOjZMCGsad07rKygJUgo9+4+0JyCG0JqcVDV9oLEHgztqRntux
ERWgLmjBt4cstiutQC0RDqhEUSL5lm0F9mSimvlql9RUj63wGki0pF65Zlwn4W9dSE00Aq0eS0Bj
5Xui5bw/EyocC5zQRr8O6gQFi+JjEWFpSGBdQNFW7tPFiKsDt5jQVJIpQ17xUe3ZALtCFxXM1X5x
m440oJVwNhMjBU68fpXIwGaKAihM9gDVLnJymnxrv67F0SxQ9Wnw6t24eMgGTOB+PBRX3ycHVrG/
O50/bqFcEdJo+VpPuIN7u6F3Qq6Dr4YtZFfwsFNzBhQR9aeTwS0/8zJCcPm2OuOoSrs9ngw8MKUq
9dRuPAThC+TvBhNsGSPv2A9FtEigYbvftBtT3K8jqcJqWWilwVkbZEgAJ6yrDKgHkoDHupQGcaXT
7sErwcsFbPaNeoC+ItyRCS9ymIo6nYPooU4LA0JOy74vrGcGZ1OnfVKvAwztGad6FEA7416jb+n3
TsVzev1soAUndfAHDgykGFT+XzDJB2EJirKZTFw/jzsHwOzfIQkuzvT1GGUtkbB2uFtWKOLcEL6i
edN25fbSfCn0UEPi8Mexm/5am5BVZ290xUJ9pS8ELXicZyjjpWZCrbRbDGz8+gUv5fEc+eeFv4IX
6I/ZF4B7UWS7/YIOYoRllx/3zXP4ivdXW/TjVXMKjlNCJP0+7D73jplGGMFLrouERXBDbTY/TfUg
uXZiO7WPDCwpbUK2calZyYspcMQ9pwyrEI1xgZBHb5Kwgz6HVQ9SRNkrUEJommZwSabr9Lgj1zoh
iR9aeEnHsks72zZcU/Xp4Xxd42pO3sDhkQIbB5fDZMnHtyUf5LVRweKV+BN4rWUbEc9VLC//I7dz
lz4N7oqTo2ugptp71Cs/Yvok/vgESjpSsTNsejMkBQ5aMug0262A9l0rq5Yd35uP1OEu8HJ85AEy
cCxJ6JoSRGZEbziGbz3u4mVpw9JYFi/L2yRTZtMTwTlpY5TWESIwxGH4t55AMXi7/b88+EGKBB5n
+Jrumgf+AksEiUp+1ZTo61WBtO0vvUb5foAe88T/FIHiBrd1CFN8OmczyeRAJAGGCdaIcot5yQLr
teH/PoNDh3x3fGbxMCc/4ZnbI8b+EhEea4YE/dlafslEnHkPFr9O1OP+L6QxajA8YjapcoMB62oi
BSD3D7bEw+zAOh+/g6t1WQQRz4sKkx1ecX9VAQYzJoPrlrv9clKETeHajpBNhilcRZ02TKDpJhph
+DfZCTJc+WUaMq9b7zkIPHakFOOcbFsn+YlZRwLKswGSPX/pzDEsOSgl1PuhhSWB9WFtsmrM2Q60
LrJKTcSoZDmcfujAeNXQb8XUAnj/MmNOLVs2sKCpjyITcrzUn3IFgVkN4kkivGWB6+VOe9rmc1dL
iVtLuo8BtogNCDnxDvn16N2IpnOYTQSRiXLXkofHOVe2Sw4UTkz6kFIPwcR5jqBvcXYKfVaj4iNk
wgwGcCx4So+rsnMK+UC/n7xSjkJgzKpyucKAaJWyWjkYA+Kvh5CxopBsmUcgfEIXDy+TcEO5wWGr
saqI8b+u4PL9WyJ5qHIN7UpgZ0sGjteu8jec+K4r6saopSS35BZBNBdJHDVJehfv87OtzSgAzwtj
3UncCb7AcwbFKeDDZ8HXvbi4ZXR9b0S72d35xqR7Qx/MqqxLGz7+lKTiKMJ0zBi6ExD1NjOa9Zyo
6rhYB7hNuDvvZVRPFM3oRDtiNi/wFc2YiQHBsdjnuTUTYReF5M+1Rq9mL135kRNC3feDD6Dx0shJ
um88j+a/aMGhUa275y+smTCK0qjPyxSgR4jh8e9GpFX9fpjbR1TaHkEqU4llqAQf5P2YMurtQtok
EmTiZmCOxTWW4wPpKIA7BCidQwha4ovoAHi3jH4uJYEbj3X8mrQfCaSfycGJv6JNArRMn1p95fXO
wsWdMp8jXwzjO5mQO8wP3eKdtzf6hvSiIBYr3qf9IoRxIDegcfeoFJwAMSmSz/Po20zEWVXMl/LH
30c8P6hHFceZKlt2BZN18OSmKmvZUB7fpBr0LjFIeyWuun1YmwVN7ZXeVNlLbSRnIGJLt9/XZX5H
vPT+qq46EQCE51YCI6CrhVgEhok6aD6vXY/ExoQxjbEqxZdzGdlUso59W1OnuYUkZfUWqcBvCREI
wG5RHsCHActzmS4sdXujn59K0ahipLYAzIJ1a4JXEUshy2OSZXaWh6YLY6/ejKejtkwaEUZLAvkS
gZD2/YKIUf6hCLg6flDA9cHqhlEOj3bzDx6uVVqlIZH1s5BdcMkwaqt/C0SS1lJ7mVcjoifA6RyQ
l/JdPSks2WcxKU6xv6OK0ab8MR71RZfmlo1JN1QessWGwQvVH8GO5goiFMCfkbmAV+ukuxzPOj9p
v7+3qTQwwdQIw4UxlMc5ZOGCHZp1/QmGw3P3THu56xOFFK63pgsnrHHyIr8ucYvTGxxDsVlMPe14
0N7Rxmy8NRCtJ8lic8R6BaDG+KOOVQgaSDv2sdzAR++J1JwUZU6/I2kpfOWqDsU/VBDtt4dy8v7G
Id9wG3kk5SGg1Zn0H/qI2zB/1/k+1Ni8OO5Zy0VTTNTJybbGdamaIvuYMtCeEjPm5rumu5+UG1fn
YQD/ERP1tjmWtxBTwPPlpAOBP7T36/oBrowTaJZLr63z3fkiK47YDCWNf2ETdHRg1c2M/2bzJjHV
bSHot9UUUq4urtXXgyEqA6pkRudiIUHIhfo492IuuBKSHlzaZe1q/o1nxDkyty8p1KUv6677Ml3R
5oy2gbwNShItw7qsBWtYgpE0ZgChQwRZCBnUAaajTg+Nfh/wj15MDJDWnaaeDiLOpfRnlsOfMCVw
uxqMwdHUcxeK0zzLZQuEDtko1I7aueWyFFa67mufWtyjqG82FL/8rd1KXBxit4sL0Qk6ngldaleu
W0h7jOGxOOpYSLd88CmLruRHnbmJ4ynYLbNO2wovPJMKr6qWU4eyz4q2IlDpsYz/HsDGZUDRAmtb
YMnPUqbBB96fV5U5wrhVtPvMOwihwjIkwvKsho1IJDMAHswhSam3yM6DjlyZxMl2ZKUcy+l/PkkE
qtBg/fGXTKAh58L8ra0Orq18bA5qY+gd9NYz3OJTYXbzOoSaLnrBd9a4y31rZ6W2MsLy5wZdh0f1
XL6NNtfhV35XBQ+/UoiM7+kgVvT+pmLU4MLZRv/+uneOSuo7biZJJotAmla7k0bBkEyUv/mY70Rz
DrnIr0OO/ktjoxuX7FcaxORCVrs94LzI5x8k3xtThK+fki0e2tJ+O25SygUfmA3xLfxHH1dGTguE
a9osTw6FLVQ+eDkfrpcIABmfdvRLehagUUoxobybPa0JsRQSt9uGiGb4YsU7yVW0DgnHs62yja4B
YIr2hMeRJJQJ/PC/d5FrScFliT1fp8pdbo0TBo+QEOU9ItIuG00Viwk7yDBau8vQEBZdcuEjig/D
VeBuo4f/558RIYzZiCVK+pnwGNVI2AOLEwAG4goaWa2/TFJ2N9eE2arS51fW88J/peB6Kwojs1Qf
uxoetP9IOStpM+slpRxAPq+06cN2BVyWgDOjbtQCKtOHOQih31eMdymUOfHRxrtrro9u/XpPGGfI
x9uO8QL23ju8PZklUh81tbJSzg3GNz0YeOsSsCKoePqNx3ei0zFVe5KNbe+hCXgus8i/P46grABo
KLawVUDVElTD+kuoI+cOjtYw78rmrfk93Rs8xshkdMCiOLHZaYxBke2i7JmpJIj/ac2vyX4TuY9q
OBmtq0v6sydMlI3T9t009PUQSqMHsrnjb6rDgHdmKaYxfl9xwKMIGOyWcFeQ3b2IiBHL88sfOmOe
fpNwzeCxzwGT/5he5+dHgdNo+KXwEPKrOTCgaQSI0TBq3XtcUYwLy7WIhR0t9tdO260xi7F0Drps
w7BObjNCL8XTh72vNqraG7/0n38Ixl434xObWopRTP+OGdmRE6dVCPdzyEYI9SvvqFi1tctDm/JG
EeMVFHfErFmuRRXsI6o6cJYGe8k8eC0/xo1jH3LN7D5Rf4aZM2rpAc33s7IeXYgb1Dpv4luOv3zO
i3kjacjVc6rIMgrzaalyuCTsPzgx2/Y6QqpCqee6xA+kRjeB7CasfKJiE2deobLVPi8FHYfd9rEJ
9sW2tHTFF9rzCwLDTkTmTMpKXQfMaBGwTy08p3YOI401yQWqWmMC8y3/KO7xwTzGGDMWC2OgGg7E
nS048nJz9DI3QiNhvN1xwp+sGrAeCQA9s++1KRPnsRNKTQkmy/CgrZR69n7PnVXg2AG5JOQIzLDi
iuADB832j2w/TBhmZAr+MAdg4r8+wB4nQxugd40BuGFcs8wWxcDLHogr9mhHK0TykjH1TTmt4kg5
59B6G1gzVyNQaiUQVkHjMWu4we+wqPl8EGFYtVcVxjcVJa/NrImXy5SgwsXUmhlZkjmwq1qeBLuQ
8pIFM/eXMYO+jrZGCoKFNPHNWi071216QGoupXGSbiNl62MGknhDt5B5Msd8hTvWp3c8+E7xyfFt
e9kX/CnMUjvLhONCskwxFNZSsSKZ7FjFxx/cRDDaC2JxTuz9MQqSwk4g5ivKLNZm5Xg5YbqzgKbL
Of8VulBgZUCmK/CHwP0HrCJeiSX3SqZePZC+0/nGLAq8elB87MigAxmavvo5VXZpVQEomKtym+by
gvSHoiidCwOb0fgtI5Vb6csRSLCx2a3pyJXUkTfKnomTfogIIp4yq33fGK3h6R/ydLTaE/X3p4zs
xWhHnNUpbNxCyJYHKjlUgXfzYY3HRMZUnf81q4a/sQs1sD7Zsi0iocbEXQLzYB5KQIwFTsZ4tMn+
8d46klpBWkJd7iliYnKBaEDcuiWjR/IgaNrHq5dE0SEWehaqiiQqCmS8nFcbWyZ1XgS4V9HxBLcG
qq0AYGDE0VUDJx13SQGy1jcdr8ZBXhLaTaXHYQqQRIeSa+S+HeQlyw9T6OoQ5W2K07I9eq2PXkBR
+P7M9YVIAQsleEfI3x38gdPO9KRfir2wfdDnI3SnU9+hOC9luEz8/ZYPMbyv6kNM1XnrtUmOHsDZ
kglGi01qCzaMZo4f27+c77mCdBogqI2mlJG2wddqTk09Nl/AwV16p4FEZ0tn0sH/y2qw8q1XQFxs
rcEHLhyyezaQUY/4Dq4LexkNzEi5ODuQ2hcNIgrbdvtUQNSpNMk1wD3pa78JJsa+QntNGMc8Rc0a
fK/pcA9BTG2ql3AWRYzJwe1wLXYa2FGfxeDdAWSOPmIIsp3aKJ4lGSt92+zR0TU9b4wqxRe0ENhZ
uiFHB4AN2gpcdKOq8IqZYB9k0/whV+7xy89VgSRxv+BQBvJsbZfkhluE1yDVX4/3Yyu43pGADZcS
2XWSBK5zXztsUckXhHAN0T6VnDyuulsKjdqO8sWsdZrQagJbDzIoEbD4WsE8DZpRnx4I/NUbB+f4
/OqAVTEsA56IxN7A1zE1G7S9XP5e9SIbUx2Io7R3Go7JzIstjTgR/s7g39whsiFmpf/G4okNC18y
teVBh22Uglz+eDT0DpzgeGV3moP+sPOB+Ha0Vh3SoKWLoqskT7ssuvQ/0BTaAV7pgmUo/z5lB7+G
pSFIZH5Cm3dOZvScZVrQ36qlHuu6BvyoVndYGoDMjfquTzYHarPR30Ea3Za07DKJCELkMXlMv4Im
i5buKHRrL2RLeBTzsuWsFdCxguSZLjdrN+xi4KZBBsHYy4UrRrCsStwdmTTspoiZXoa+x6TCIzz3
dEoc59JrszZZuXPVaRdUa1Ti65mcJdZDVujXvN/yWIOYxAoRd+rm37aUWQOhiRmP3UOZML3LQsxZ
kWf/ZhVApMUkLJQAar2IYsdiHj15HsJcgKLF/YprC8t4ymEwHzepQPRrVi7inGohPG5exhWsr4Ul
/7e395uNvD9cWCMlDqWK8dhs1Lyn2Hq7tZ/K574CQPip/YjEMoal3gJY0YjStWmtnAVdQ5xn9lpw
mQDrR/6oqgyoKgqc53Ti1nxhuIQvoq3SrdAR+b2rEf0x6jp0FvttiRJO0SqJe5Rh5OuGBvbrvl6z
yV7eVma9PSRY4zKnWL/NShwHAj9nld2mPI6j2Mzb/wT76uCm0HFAhWSVVErgTnVbS+oJ4WiBoFB4
yQkrd7OZcqZxMy/Ad9twByZmdWIInRYyA9n7Ni8DR05+XmqwbimR2LjXy2cM4lUlbcjm2S1xMCbd
xsL3M01ykYLlO2+iLQt2j0xyRvjyMsrYiXpHapvIuv5nv+ZBmRrNCddK4Yg7QZEIHtlMTGcLl0eh
l4JuikCPSK68FDKuVEW3R90aV30R9FzOthQrjGb6medeasosjyy5IVTY8wVxcRXoh/+jxZVk4VkG
F7eZXA1RhLJhJZ1TfAlHROaxjxwrx+Kh9M/Iokih/51qCs607OHjzF79EztRZI8YeMY7AhLVl43Y
psx/yYOjCGrYEUMHvWFOsEuR2oL+6otaVFRZRm7F0mEzuNIlJRBrV2NYx+KBjb+U80eGap5JK52x
1tp+5H7iLIJ4Lr5ACJppWe9URXoSIvKPwjuIIgXUJQ/kRsmVuMQ4ngQ8MRBe6p0jOuOBYmoO93F3
oFfkiGTsEy3wOl96hNqISseWJQzMPi9A3i+GlgDm4rjmWkVsMUXFKFtnv4oLK3vyhKIbWanLPWZO
SkB6VbbhUp9o5H1Ka63KNAUV+3YDqoxY5sRYGflNxxRAdlySxl+7sAtMvMSq4E+1oR9TxQqN6H1G
WmeIGNWxqoRuB1igIznqUSk40tmD8AjrTlABnFhCmPLp6/leXp95tvwfPmp6OntM93Ac1TYSEHHF
oXnLAxp1KhCnXejewgCuD5EA3+01RKDS5t5p1NCZ/JoaV3WMc203IBFFb0Rj2eh+j2tJOCZA6AY8
AzrjFsuJGaZVYl6/qHC5k3QogWpgUBodtgyMQIB+wlHiUBNvd1Ot24cnWuJJb2J5juJC35542/6n
faxYimQHK5pT7mCko/qZKX//ghsKg7GDyutRDHRV2UFdeXdwPuktvQB+Zn1uZlCWy4ZcavVj2VyJ
dVn3143gXXXsej2OkiNsZTyySm1d1ozw3KaDvgCq1TN9wYno+QwnQqf8RT4v3SJugYg2Nta7UUH7
bJ9qcyfDCw0XerA0R+c4d4FTJ4R16/304SVoAxyxeik1tIe/UcrQFYYaFOWv/z8QLiW+Brp2AU3j
iE3GhYa0lAr+g54aoQITglrK5yFlOEbmNLKAkxnuV2HJoW/dgB+LuRhHfU105QiHR+iZwNmYv8uu
csal3VIoxxkBbu5yK7Chd3/P69AxTpX36OfWJUDvBMOogq7VueVebr3knoViSGa4bhjndOdU4Dmd
NjPsIWjAHAB74Qim5caULdcW+GDI4HaDN/AA1G8xy0SMlHHh4w00XtjR7Su5TGcwjOFNz1TgLuF3
ld2U0qo1Hvfi7GqSYzZO76BS5hfsEsOnTMvnhC9sZ3K+o1DLYj4k5M/VI7bxl+h/TamLpeTL0wNk
9KKVJclE2u49PLBrq/b47qvRejI7DTKWiYdgT1cJJ0FkuGG3uX6NamIhQ5KahE17XIwv/P/QdOAk
w2G7SIh1IjB7TtCeyEa74c0Fb0+RLrZ7miULiMOt7Xd/nOWIyq82r607aqsjhd+lL9aO0c0hNL5M
/QgusndmWEXLPF8+tTHOsi8O/crSv2SbdM1p5N4y0S30H1T6Ns0DIBM1EXO2MkSlW4nYyJeIh5ee
sNBdxIMda3jGFPARdzQfNvmYZwjLEo74IdjdoPizK5XDDUbnkOy1TDh0S75HkJKIRX8DpKzPKBLB
O2udWRFAGPTEnGTBE9IPpfrA7B6VJSVo2Uhy4EYWksQphcwbOzUqop1AJH14hW/SGtkh4Da9FWio
WXsbjAMhjnEEkjzt31W6wa3Hd9bmXc9ffxKVsrcOz1qVRE/M60gs/J8xiBIn387eRzP7ekqHX83R
kJxcjsJlF0N6O64so1ySnLdq2CB3eVCc9os3KYzC98A4CqMv5xu6LOJWr8zcSBz/gh2IPeB2fKK4
Q7LJjqRnAxv+W9vdJTDcEWWAfWnKHdh2qXb+nyXE9oOZr6PpwpDLPONcCLXKiRrjtQ//TMXws0N+
nnNZK/ABDNSaWLSG12c1xtTJg3uECNAINStWFfXfWKXiis/Jy3BAU2ajAuVRGecpBwSr0+cKzWod
WoQBP56Gu0b3SwUH/K9trvo+l1st3XWwiLRqCoXDk+rJpodvpic/wCOsbNdVEqmNZY/axAAVhXNP
TVmY6O5cAFB153Es/CdLjQrJsG6CbzLKSud8mAhDnsYVefFP9msq0YGP4zCz6ejr4PYKBnk1uY4I
udmvXZJKS14w2qTwVVZcAUldHpoFIw9M6Jxk28ZH67n6LztQlDoEPl2vyTTP5Yig3vYbR/1dNzxP
2cyQ6JtpB4+0W6/+XAalP7hspzI+N6smPYllaUViz6rgFHLaJQKhWIWCMVHVXf6i/hxclq2HePrT
qI0bsG5F0dnH+STqXsGNOWyg8YzdjAS/3r2NzGE6LuoKHfCZPGmhey2GP/52Zfj/7mwjRbAWxxkb
dbxI1Ad13mFNEp6BX/zOUfZyY/pfHFMA+bK/q/dEsIyrjY64rKvL6he1eQpudRyJJvfd/CTZiQVJ
fhgv7ctwA6NbuUfuzKQztChJ7DsCtpN6FhcFg6x2qsl0rH+65r3v/uwgfHYIH7j5bqlPyIjtAtBO
nbkotfK0vNmDmksXS7q9NVrQkiB4ktimTBZoddkl455O9lKpFvuzCaxGLBgLDPysD6XwTrFXUQM9
ui1xC5eoJKulGp/l4e9LIyFHWGvk8HCZMncH/qVlFTMbOKFPUgfJB7kWbPqzmq9IUuNRPkKFGfaI
tOBgw3ZJpNITxwSr8XCNCjqbC39mTwDJV+92RXrUbkEaZj2virPhg/DOXsB+tkDp6ai0iOCe/DLW
Bgqxxp29sqHUeVXi4x3y0Llg5Pn12Td7XxzZrV26V/zt8QGF3UCBEtiksPF3BPjiHuDSM/UQJPnF
cRBI9I6Z0UArr25CW/ATNlSuQv7vQIWE1ZffCsZWGlxQOgI1lnpJK41kYNVew/DSQ7bXUikyUG5S
3ToLWD83WgDuCkE1THRoEz3boEjX07gAcIW6vE2cFXrs65P2uUo358WEJQa+gAwSUGeHZW4ZA/ez
0RTRTtUquwX8y5dCS1Pn5Wi6nflyloRhIKhYf6PhyqwKUQYUJetM7JgQr8yry7eGiVM5prpexTsH
W6oRMMsAeSE8fMBI0zXR2QQuiOJvnI4ShIsFBdLnlT19Fszks9pH5dT6k3GHmD6x3RRDe52LH0ln
dxkLTdsJwFr6f5ZI6p/oJ8VPZJwpZD1KZTEVhkNMwaedTbXGmaYPrYdl+KASc8lcVun4+X9s5gXR
g6uSN4CGANKlQk1bjKBkj+8eFergPyz1GwdHXLEsZczg9WUUScALZCdKJtdd7VNtmHpQR172qqvK
PtutlL78PP07VRs+S/a6avtVW9DzdiNHElVrO2FN8kpIdhBiLB0fBDXF9h6KUVq0Zvkdkx7QjKfY
4H8j0kQzHDr+6sShjsdONSiJRQ7TxtAmxV+Zs0SMNC0YhXtXdM28iAfBR1gDL9IqIi8ZZjxwU1tw
U0w7byv0o5E8Kfl5cq+cTZN2OO2ao3l3dqab0c3nQ7HALs0NVA9lVKOhbL23eaUU/nFgXouVxshM
ppHjvpwBUN+aHqXN/KIR2gGEhDzbnt6KMcc/yrQ7DFnXJnZx0rLsbNEIfLfhz3mHbS1rTzROK5QD
WChXRqFzsXFQz+mu24a0/PhUHSyDqEUbU+4opL7NcWk6Ypn+eg35i3YznxrCyQX2C+gIqkBIVyW/
qeEPfHBlupDK0uaVQhXXrtE59oTmQsibgruRqP/5AK5kgLboLsZWC/tiCasnbRxM0HoV0TxXdhg2
j3qY5rG61q/SQOvOvzHka1hLcPtT/kKp2b0SejhFIYZ4hojEN1rtkmXmaWD+FD+KWyDcsmWbctVD
MB2e6Z9SKcYKK9uAtpBE6kcYWfXd2xqW6/otTy7cM8QV2o0rcWahgWdkM3Y2+nwluSHvDhU25+Ao
oIF1/7TwsY0aRDVPVHDdf5Jcku2d+NqzT6Yw8WRD/U5LY95nJaftqEGMLhUcaZP177fZaPwvk+G3
fhhLowHdlDzt8FPmBwt9mMLb3vHfAPVODggDR4KZkIVwl2rWOTIK9OUADkwvRnMOWBGfNttQM1cR
RUrTV883nNDka9lknJd6JoewZBIYZxm2/uikyuAFBG2+hm4hFQcwlOgBl6zsa3A3AfoMU2ZNlRjs
RQQuwiGgJ/CqxCNN75Nej6Q/N/1aS13eFqaDRAKSsMpGzD66ATI63btusWItdg9XI3TwmDTag6Uh
cEKXk/u+kV3E2QNGMjB/dcLTG/erotiyelg+DOnsCt7b2tw61ZflCs0Hw1uhiL9chXB/Jw8ThmKu
97MJuASnuVsvmI1hWYozWkVlHfr3z6dPWB6Qyqe3nrYFmvY9vfyvy+PX8og/t5RL843WI4OUwsOE
gL2QLygOFlIwaZm8kuuvuhf/8Uud398tu1GNtqZj21cgqPE2tEjaEhqVEYAot7J+VlEnIolwOHi/
+DxLreSdGiQotSK32pihk+AFakomEn+hHXlaSbs3rf+alab3o5QRKIu3Uqhzd5CCOMKWlJMBFUry
m16oEuhRkJNjQLLeZz0cTeGzHko+0H9AUDDB8CkFLrfLtv4jUhFM3rkyBXg0qlumePSABhkw5ccJ
eFFBqA6NotHp4QqBzsHVMuRkG31lc4wBpYh3CFeW4Sx3p2RmIcor3v63xWP3tDs7p27DNp01zyYk
YrVqJC1goda0Pj0MkV0hSXkRaM3G3RHwA15ocPXE+reCcfi8vhieTrNvG+AdlujHi3z+aAkwvb0w
0Z8OXTMEi/zdb52j5smbpVfztMdk/+qtB+SiIwSIWK8KPnGhIloCbENKOnxYC/qfntDGNn/411As
lhgQuZ6qu8HBX7Q0wb5DSA5kuvxMthluIuSCs1Yot27xbjEPlvJCrLrn0BRb0IwG5UqqBvDSEG3q
ehPu4REfW62qxlhozeviS8l1XZaOpEl6CJ2Kb8UcxblRzWJZt/pB1m8BCRgovub0WuPNTuxd8wYt
mwaR5zZtruCHngUAwQeiI5WIf3xMBBDKc3Nkslzo7nCjEkBm0MecOJNhijKGYV93m5U8QS2/y8PX
Co/Y1NkfqMPcDluSNeeEKOqYRz00wtpU9Jexf4+j4Xw5QRHzoaK6F9lt21qCFbWqbYhT/iTVR594
Y//P1cAltW9lu677vYBFCGuK9K3zbjzQI5vpM/NG4pc4XeMLXBIDb/B9iN5yS5/Ax0ZlM0WPW6pq
9ZCH5bTMIwXMuDSdxXIiveYBk0bg5NGfS3NCK0fsHs72MkX9/hVac4iWGECeVZvy2DjjPpN3UlFd
Kmuy5T357Drv1bXt5VdMBS4PHw+yaLAhfB/Hr4m2pABeJAG2F/FVeAioLBYRtGt4BtRKS1Vuwa9y
tkHXMNB7VFHa+fooVF99RQ7pPZ2NOmVV52kmeTaBP1oPxjHex1hNC86HBpNpy4BbSu8KfN1kvKxl
6UrDRFxifJPd3/7v+yh+aEzOR4lnA1m89BndJ4VjncHKDmxz2+xv0Lubf2HhFKhk9+8kkgDvAM9b
2ZukpyvSGXSF2sFyYCEt4/rzfX20DkEk4ND5JTcF8nLdgm6+UGb3qdnaLBYaLw5Qx2diOcwMdXwM
lO2xr+AmW6RAn7Wg6waK2C8h7LJ4wAqFujUxhLN4E0WwJJiKBZgQJ/sbPoCfUyc+eLDkQji7DkVA
1NcvzmAzebqGD6/VUxKGLdiAva0+a2qwjXexZx9jvwTWbx9lL+2SZe4+7fOA+0e0/dol2ixkQGl1
QlLMFQ82qrzsXaRkxZEmaA8Vnf/9AXC1xQ4js0kJL8dc5WCaM+LMFjQH0YBq0D3rLbkh88fXYUrt
Q1zbBncQJZLdQeOBJZ768KhENJ6N3CHJ9/PZzfJpFBoSCNAseZzX7Si9sqXJuBqDD/C72RCPGcU9
KITSd7HruiMAGR7dgXJzcCfWZA0RfhgP4xZp1zxZQbVs6V9dIQQOzfEbFCiSvi4eroO2njcjBW9P
NzvmFJhdc7uMhM+Yyjd8vtNkjE3BxWnhD7+W09tLrlTlk2Wc5gLCvHLzDUkV1ZJuAGv+a6SGe3H+
iUTIK+BXBw4YNEBoWiLY6RJzAfEsMteFri6uuIpFeihgkP3rGPXNbJgW7aBcJ9wbV0Jz9kEbQXhA
lhkoGwh8H65BMcUCQjRxq6W9EpJ/RxEvCvjEuODr51Slkk5AjHKXbhBbkOevR1AkLBMkmdVCCsdO
0x00RNt4k46TKyhokFzozUkU4PU2g5F23OfPyWKcBgUIC+7K1V3WTy2uB2C+BhW/tKLbmaORV194
S+VqWtJmEcZkowhVJyXXTIzSmzKD+SjTMgw3SqKsoIxAYeM9toLIj6CjT4MsTVmJInGJRjqhfG+M
NR0O7iAYIgFLC5IrnUvff7H5am4AOjuVdMkWfsvtR1qmOy7aXVnxlUrbtMUrN/yj7po8hGBd4eU7
U97EdQwtDZedm2TDpJ4reApXZwxOpNeXaqZ5/U12juTOU1LBpAwRq6+OlZH6JsyowaVQq1lcG8dz
skbhSi6LaUFHqtMutHKrtLDYgVL55qiGY4h9YeqJg4BhaZtUNyHYbqBn7yfVUOpBypkpyISq9rsX
mBnF4390homSyZVnwpImfGdLhyXyIHlQonxFDWlkFAduTXiq3IrXDVDLcBr60/rE9T85ECB9EUJE
nQGRh4+s3u3qc5Nkjhkt9XljvYvJVLiGLok38t6Ogyf88Og4f7foVp/4kNQ01c1W1ITlnPspT5DD
BqMVZSyBBKxMEf3vwYtAY506E3AYgrb8hEdwz+28LyJuNe+21LlzgiZ/KjYtbxSFa0kalT706SeV
KLB/TXz2k31qYSd0HHxToSNEtkcexRDfSfZ1JBDji3u2U4n0is2ltyql3ifxFUtUCr3XdMbbNssA
WH3r5bXl3DPrhRfpmu6WrOeGLXVz5oVascUC3VD9W0o89PP3U55BXWZwrSLn5gFLRqHhovuLs+o8
XYKMoiWogfwKGGBoyG2CQziX/Cih4YsTYkGYU7JCLNIRslpueqJy1HNNqO7uaiRiroeoNfFcQCGT
MQ9j6DV/giZPh9lqGvicKqHF6y4VktJao64k40WPGM7flOvqvyEo9fiFi+hSguZxyxSQai77em/9
HG8fgV3lVkhpbF5aSSdaD9RojFvVAwQjSZGrtvmPbq8koIPNrUbdn+hIXcSe1h2KloA1+f9BN5ol
hzN8KoijZ3IdoxGuUTw2Vsi2Bu1ekXWB1ZPbZnZlFGnCJZRUFntmQkwQgWZtmcFQGwHNIH3gbZiE
vv3PcOkNUzbMYm7DUgNJhV29PY/eY0vnCMQeQvLTvMqQwxIyquCIDyM3mMJk1LLF4pS2XDaLSOVQ
yawJoWSEHPgoZG+x+QZg4ss/dgMCmvKweff5amc3tzLDgccNlV4Wpk4/M0X/8vQ6Yri5Z8pDsGPb
hEekTondSwGvNxzLTqsdq32Fc35HkxvEwtg1GVVa9YflKUvqfBV6ARu+JjHBgEOCOYwly2s+BOV3
yFJIVDV12F8ngy8wXHnCZc+XnvBQuqysJjbyBhSm3QoCHbuuYa0rlTjwtc4js/JyKckXPpIoCQ/V
WwpPkwfBEv6ixy5tioUMN11DplAkVzqC0f7ITKC5w9L9jrHzyMkI+KO80fXGyHddElVV5X2eaGyR
S028o5J3RhF480Gp4/k1HQrQ+rX+54ZDNOSu2iae2W4bJ18AX5KYCGTVDrFdIlxfw/FxZaH3kNAh
oHHJFJfqP569L5NyvxhtqqoOq5klgH5wwUjAUI9PWQrvMSWnep28AW3nJLO+VO/Ly1xoeo8fbHj8
cI4STbzI+AZyEnwQj/Aw3mfXxF9K/Rp1XflUixh7VEfpa9M83otbHKYD57IxrrB7/moUl31QCaFg
0yNqAXZBjfZ9SXERbBdSvyfJTFgb5MxNMvrfkwc53SfJuHi2rw2ucPv6M5hASabT8nGERAAYDrkO
0GqBHYx4wI/XOWDDE5I9pbe4RhGh/hMRNUKO/xZxYB0v6x7A5vrr5MH28lPDfq9yjso9nHlDTA2f
EECzyIXoyCPB6T02B+Y1QFfeTQX407RBR1CjQ652vNqLDG9/eltrOhGFsUochTSHbM8sGPwGNOUq
7vewTL4zlZsEblq7Bs4vyLru1mjx9GYHiqnYAq8BLiuph5KA0u3ZQShoNSt2HmXToItNxUdo4unK
ZOmO90mhYgdy+Zh0+DTKSSQAeArzrCNUmg2bSrhape9YqQtC5IgyP5kqP2cfNMoXu3TaYxrPkfIJ
WUtlKyBqzV8XqLbpZdyo7C8dGvK8BUMgHBdDMmgJDQXb/4gbBHY5v8cLuFauQfG24WgkVF9cH3EO
l3Slbo4UvdEs7SVyMuwNnunjhxkng1VKJZDo8aIOFSHooGpaULRGRXoMU7eFuhmpSW7KNC5eENtv
5dp2/3pfI54tCZfPxCCrdB2tqPU3KBplAD7jeYDmCbLYjBk9Q4fcSYcGuEXWneJHdu2SJX61i+Ez
5vGip1lI+6RFl83h1CpRNDb9DkoPZQ68ZmP+eKRkjc4Jg/VLM/zAiZEr7QvamgZv2irkX0z+nM+q
YlrbrznzZWVXAOMAJSiOgZtbK2csDSkhnazUgLafHLl6Ixcaxu+vuLEkoiROmGlHCFyLYy/hpm0n
K/7sX/CqEtLfky3Q5Witke+rSFH04uiOl7bGF2xENWZ7hGSS4cDINg+3rFAo78EYqyRKe24BioKR
0IVSXTWjZsVwqsoi9MGFEvR65x+hNk4we0PcF5ToQOdOshrvxKJ8XyxNncJqbShzRH5sTBnbh9WB
o7w/xOJybAi/3Uhc2GcVMVUj2D+ToyQ2NmYRh4S8BWlK0a91ME4bj+SR18LH3rfnO7mxjZuF9M/5
oyhADVLySxsJna1Cb7Mr1p6PpKXTyJq+L3S5SCAHz309ND3xn9rJlKZ8W9CpLa8AsW0Z6OYPEy5n
rSqVuzPDxIB91MaR09YJnWt/aqAWLCkvICVGH9eOaVVyJ7ysEdKq0QsmpJmdww5u9qz/U4OHd8Gr
CdKg48r4wiKleysyq4LfqlgymxCaevOiZjq3l1Ep0UrXhfGlzF6ULiNEwZVjiGXLqT4p4nenySzu
jU4pS8VmfTgWqe0+WBW1YuoU2RMvXKkYun22+qz16CyDd9YEdlKNn9twJ3xMdp0FanD4/n5NK1Lx
hI1fRepmk0mpuzt2ufm+qPI7P/sY6SralFyZv8pkKxA5ZbNVM/dShdLr5NRH2tuGdBs3qrJaMMBr
d3CL82m8riPEroMdN6K5yBqhNFu28FB3Rb+KbcMWfwwgLbuyPy0qErNE/1pA+i/xaKDzn46STI+f
vW+GAbW9yAAspOvZFO+8MxqTgcOjWMxI+ZpXIt4X/tozvVLkhrlecoIp0zU3nn5doJ+Va6m7oYAU
zi5mD4+a/s9Q1L6ZbmX8eSQDOi1dz3rDitHFf03ES3sUcBo5NwDPm+0F06MltjndMuj1jPpY+d4L
gwUSZOazYaucuOqUORz2kFYKj8WV120G1MuhZBzTpDgSWKS+TsH0Jw3VqEqYCkX2emXKWszpnv4i
1OfOOXy3IepePah3rLLMQO0GZpQzrqaeJKfWHWPhsWDc0KjqkGwFiPv/EA7q8vFlquzb2aYYzRmn
X6mapKRjgI2KE5cPi5auKzwQ0/hdAnWZ6end7Cblr7pnWqGipIMEHNDl7VEK8UtQF/k6kZVhLjjt
x3sHs+Ddb03Nef9RduJPsoIV3LKCNRiTBbys0KxNCjBcknu3yGbKlNUSJvAOTp8kK+LyQkhPZlpJ
iYXi68wLG2HvAQADa66kFTVSdnAmjTOgt1lnUSVzS5RSKVXu1HO9FsnCh8Z0odyAr+U1F+9JbbkF
1hb142nKl9ZHSdBt876S04QIo0lbEPAKhSwikX6Y1EFCHylzUW+fSpp1WIdFyZMvD9rLk61O+rwW
/1x1fgK1FFD60jgGEJ+q+Geim6RhjV6w6ELk7P3fIjZo0IZ24JvuRgYAAkiS5mJl88oxY2z0al/I
antUdZLoTLk75fIsy5B5HI1ZLokrP3hwlZwwoZQY+srBfv7ktYDoo8qle1XrsBH8yDPudlZQ0t5U
buiZ8P2SV6yyDns7ZO99RuwgLWD0ZcrOe1+DCGT+fWPkITIwN7qG+2Aym+f+1EOYcjEfes09NcGh
qjU1SzXOQbhBklyh89xoZc+8u7a1xVHZcknikzAUazU7q3F3KuPk9pN7jZkGK6P3WpHAXY4EWjQ6
/CGcbcQumwae9uPJgXYykfm44qK/I+8o1qE5aqX7Gdxnjrmga9cZjyJrigTeqLRbfimgl9LJX4nq
+lMhk9KQjGP/8jc0+DAVz5WSFRns3TUBSo+Ts8NqUeCrryQvBcOQBoLHhK+GrpWRP+UPMByJj1VW
4IPObMBPaq3nFrXDeH/XzqcjPfFWoYabvv/w8ttRZMXnZNrwfjK6wPC2d8NatWLANeMEWWykAWXt
8BdkSSQ1S7TqTSH8IcHm4eKH/Myk1XtTcHAjEhoziNq6hd1ayxUbhvQWuDtWVIwsvWkShyhF6bKT
2h+MWsFBl7lXATlmNnIBWl5sOF126ZMFROofmmy9tmo3MTiQbJfjD5xrggFthSNYt4b76lDGrGFu
cKcvoAuRjq+x3xG4mvR9VkD2bcYbavXqk5KhotLhSwb2Cup1eLTT5DBOmFN4g7HEZHsc8yHcKJqx
kGcFrXZ8C59PXw6L59sTiLJqzst600Xi7WWdLPbwiNjOKPI9h3Vl5pi/zLlIKDsEiZ4GBOJyq7Mf
TdM3QNST56MJLoI/M+k1hz1Ht6Sim/rathSyTo+ZLHengoUZOpPmaNZu4xZndLfmzVg8fv8db/0M
7tQeWlZhdHia5d0fyEGB/Nb3Rv/Ji2gWHvcCbrslRCe5bhhPdLuiqKDJq/2KGhEtKHwdWqtEwEDJ
vhXNwLLI2PVd+ziskJUPTdguc51v2BE6N0lBAytxO4zsQi9h+ypovV5/VHgShecdfmiuq9ESakMF
CGED5fJPIwKl+tezGhBNjuuk7TZCxbA+N2nHLMEW3ed0RB77ONjsTF4PHPjkI26gDTp/doLKdE9C
/jhS7yDB5dm9QLNXHgsFFN6mMfw59dMcBi87q+M+evYH3U1aBmDTXXcRng8c3jMgbKvn354gk+0N
KtKNhtaLyqpXUr+w09P0ccw9Ef9kwAuW7Ltq4304/mzg9kM1OXjxhG7lTRUsUmJOtKqwq8D03TxN
w3x47T962d8Vcn6pkl6EA3uQsCppMjGhGRxtX47qdRsq4rYr9lme9pDBnjTSu+NtmiHtrA+jlIbT
hM7jF51wkjvrD1Qi7Y9dw7tB9SQqqkY3g6iRsTJHPYuvJ5lrZ/Lw6LFEG14GJVgFnI8t81LbdBso
lXWPw5LUV/U8lZ58EKO6CBojIkL3XBTm6kGH4Wn3psLaIOFIVmnmauQB0HKuKZEshJCLz/cWi8Bb
gOXC3gHO7vrZhVaP5K5a8IJckyTfR1v6RDkmCR7VQuXMKuiZtku7DA/yYzP0SKdxUWQbOGr44xJA
8jqvdwbHLlK3WW0yLBn3X/zwVorgcRJgjqjoe3ED4Mwtmj3LNCeMylCDQmNrTFb4Msanm+ELloIm
sDqcqoxDQGxw/b3BlS3cnJeuOy97kNwW3eyvSk25ZeZbMF44ze4rASmn4h9Cs9uBmq9qY8rgM0v7
cSbkWWL+fjpnf06N9jr+FQr3/18DiMVOyQD+SdEf3LdAGxGjmTJT+Ecr7Ykvl32Kz9MlKX4pMEnS
1ETX35BnvK/3PRYnZVeOHXZcMvsupJSC+7dLN2wJWCCl5+O2nHRICUQu12kgjlkfZpnCg9Kadg/S
mGNIuEkmHXrHDHGeRekn6N2LBNNCmh9c/1Hmz2W6vKMK1B6I3BTWC0NZ/zEwU2z5Z0uydS73GopW
+byHuBVsW94cBnViIb9RYCAaWb7ywFloMPKUmxNWv8ChY3QnPnfPnB/MBkAIkK/A18j5WDPpKize
JsDlwR/AkFWew0Y972HjHBwwHViiAtjgM3+LobbbyTgqlDbwvtfotaWmUW0w5D6+ZpwpIEZM1hq+
cfwlNJNv37VJT940qUA4bxz/hJ39chnUv4uJl4rldC1Q+kiaGXkodprdQTrBpowxFzDGxDQTKGaC
GTMqDpd/ltO7C/N7KXt3oUqNnqiWVBDytTFO6oBKcojQlH4sCm03Avrya1AOq/SnDjeSadTuZ6gl
MggyuW01713NF8RTIllxw+ENH3K31bAqq/SSaBZQL5zQq96oRjuKsyLSk5f1YPqIvnTVtamVIcu5
hEA+uy1BoS8VIAtC5tJrlazVAH+BSC4IIDzXcycnvyWdRYTv8R4MgClJkS+h5jALvgGqfsi+1mCy
YjxcGB1II2MYS8X1HkjW1EXlmdGtRTUHo/Wyh+MHMgDMwEK4GqS+A7iZJPnzjwfj9M1kBr/CRsEn
s3FvmDieI9D7mOHE4Q5hFrjkLMDGeCsz6h1FFvBFzchLjxJiLSUJY0IXK33ICtZatpr+g2FCFcqD
QdJPLbXDRjEAfbK8eCfSJ/nK4vRQvDDMD7Y1+x4zSeDXmXnlAjkUMbuX+Cjfv8mn/gxBjm1mwjT0
bgMBKnFMmbfMpDrRPtalIe0R1gSZnwxWj3peo8Sp3QTQO+SWve59jyNe8+oJWCsQBDVv/l18D5SH
9msFUoskBfgKEyXiSMiRyiL6zyoSki6v6CpQIewMC1xqLba0gD2is83oU/E9YnLM6pxVz9ESWsCD
LMdpAyLq18ZqPp4vbbLZa03hhvOuCUi9YsS0lIPwPrRgf+6kgOm7rwqbbTTp2bipFYL4/MbdqZ7l
iA3UMVt27Tomv6iyTqzx2iTMj30UANym61BVEnyC2OtjKzwtiC8NETKmrFlImK0/0Duga+VUfKbv
YyttbdYIpHE4JkgBlTAB+3PbX0a1ruksH+tph/skRiBU1oKtMzdXffTrdCGq/eJ3+/omgT3Ln8Im
/OOYoDA1wxeD6R2qfSB2x/EGlUUUEY9t9w+eYJDAPgwJ9TQQbmTvOCeMu6GWsHBYn0C10BsJTnHC
7cPJ73Zi+apiSAciRrDQapMiZZDZoBh763H63PpI209nFjgH7dJLuAQqv2psV1Nb3wFyQLkKhB75
o4VoY4DYeoThiG2NWXyg/GqJHpdHAwoNVli5s2CPT1grSrjMUPEkF/Rko52opwFV95Ofi6jzg854
8U2rK7FVeNErNgAGMDBwILzwIOdi+Og7mpYnCOUPMl1wDsu20iJme3nCAgVl7Czmpp6zZN3rGcgF
5oEr5RRk8FqlBCRGUmiol/3dVPHE/+HdGxWXXIRCsh+jp1I8RusDvCadkrIWk+2nNWKMB6M5uljT
CAtnNyxgYAtyLQJ6wqw7tAmhw/Jat1C6DjLc9OZrO3wLvN8dL1uhJcOKa3ku1A51rkHkfFgn5Bmj
Qnheut59oRk6pDuQe4+wJj6fnjYLPA198Nf7VOV9K0FxGWoZNOMBXcAKknSprC+1EnZBlSfGahfC
CPjI8yC0LrNG4XemyuQgv0ADc1RU/ZIRe0zDyZR3rgLu6xtbar5nd79ppuJaRYjRDw/ORpnGxrOn
R4NoJJkDkcXSpdDqbBquXu3Ii2S1dj0FLii+lF25eMxzd/yJjsLv/qK0dVsFPoPiSt657pXedKA5
b3nWNqhpWy8ToSBbiO1LZqYWLJMJHW4MDdAO6TyTdZj341wg89okVMA1Ia3egJRowwkUrZofnYCP
t9MCvXiSa+Zu/UU4oCDmjHpY1aYuFtALaQsSH+IJrg/jSayxOEQHBSgX7VESAE24bGFsJOLUwSGF
dENOh74U+vnmpLrCeN4feHGFvFi7p+pr6SKMnJU0jDlKP9pFl3uaVmTwwgiuk95+Kee+Cgm86+sQ
Irt1P85dL1P0qz6c57cPQXnmFwyslfkWtsnpl/+h3KeNdMDSuzwKqtXkGOEytSBWZ1/tZueEui1A
/jo9b2VyA8gqRoK5whaqZnjj+3ryb61P9DcemXWHhPH8yfxEKru52PgqgROTMWtR8ifMVESP+PFS
Yj2rVn1TJGx4L60wBIV74/pL+VlFaTekP2hAhVCx+EvEmL7HDc6dvzq+VS40Ht8TW26cdC472fkG
nkfccJ08aOHJ1Bm3TN/JF+6gKca1wrz/ov3iudU0rTcspid5jsE1X7iOtzyBQO/Ck5sLg4pgtxAi
8Iz0Gb31tU4/OPQseaQeE3jEg1c0wEP23jXhCQsP5bxbEZdfottT3IuwcT5W5RWm70TOw93xaLQR
npj7bLUVlTVsiG9BW6xkifMENNgbTG2iefu3+2kHuUimJr6j2pnzQb86lricsdv3RFNnruzQl2l9
rQdlHKOcsc3gNNt3prjSGps4l+nauDwRH8bv7eUgm8zrZuNQwxfUFHMZVgQW2EPIeKVU4XEw1XFf
Q/0YXSxakp9O0jFCJ7vAK3XhB8v5Np/doxbgGmoNfTnd6aXH4z10WslaBhb9zSgGE/+oCTOKgyGQ
Scr43c2T/8rjUfqkAQ1/skX2/ptAnP9GAxNFuqZ3oLllBJ65eTSIGinhal1YgawaHTdwYL2a920w
Qz07nPYFlOuX+npo6V6Bf6jTPTe+ckIqqy3BZwcF5h3jyLs+ohRwrEA6XoIr0tY013u8L0dGkRhx
3lNHdtGfvgNtVg6sG6tGm3V+V9rgktje4eoEhNwhBDInW8eOV9QdZmh5PTwT6qDUYWQKPieQz8VW
BkNWSQE+HilSLyNWheERutSDkMxxVld5+1njToj6Qu9StOC/csnjKEjTNMeLCi+gvffPCaf5MZaX
lHQW6f+/gMLssP1Lc+Cpk+NsDBiXVBDnoucWWuaRWOm5F7J/mhWywfHih5cJAV4hCksugEHrKIqM
h5y7wpn1W1zFWYSiNCConkJENo9mrW19qjpHL03F9P+R/QpESjE13g3lFTOzl5ey8n++lya/gT2W
i0xwcaAOKCg51HUNKpAoUY3nCNBVtNCQg52ieuejzqceBimS9UUQOTuos27Gc6PyYytsOXejnYWC
4GWgIXLerLVhSoBHh2+BJ8kD6djvt/MtzvqDw0nsdD/L5R8qSsFQKGsLt0f1MWoc7B6D8l2T2Izl
vz/NEh/OJGDelqTEDR0ShTgMOwSTeGhgQGp3L+cNVUHMbGsYgchFaFh9Fy2C71UgiG7PXamnMyJI
MqBU1ba+1kMAqacAFxnM+gVLvC4ICaYTrTGIEdzkyJsZ+imquskP1x/96DXZVhWDxm25z8hITG4t
eI1RoBVKShM3CTc0udSH35RnDGHpuHY1b2O44ySYP/Cr/85p+Fj/1qTUW11/5J0KhEmU2vN/58bh
BS+7fnF6zRuEJV8rkhJMDL9Ob1A/CfRCngcKogdyBOur7sN8HED7jyGxTK/t1WQ5Cd+gbrZY83e9
VbNhdi222ZY9ACpmtHF1DK+p4YCWdHo2DENcvbGt7hH8/ToHpBc4VdRdFkWM+IknFi4NYOxZtjZK
JJf60P4l6YtkX5m2SB3sU2JN1egjaryCbkL8R8Qkz6DicGW0insv/r+cZ7wZQPnyjT7fqw/Kolwm
583ogCk+eHatN2Efe04Utz7PVW8+IX3+2FVvBTE1c+9EozFQViGxTBRlPEhDdMn731/D8zCfl3RD
w8KoXyHEH6QPibxp1iqcUIxzdMPkeme0AzBd6gmbfHtNAMG8evVE3nZOzOj37wmQAauDLtAHOq4w
0QFOvarOA0v8hG80PVDxNeh6RI/6vksMZZqTGiHkBA0mZc8qNhJiEo2RCzHAF+4zbxx6i1JS/e1/
HiECCfJCHKWaYRzAZs2kIGgVec/YkZKhFtbd/9YcqsBqTtgprtatcB7gpyamNb/8AL+MKdaK0+/N
N2j9M+ZTGoFiKbCBDh9w25afay8fVemutDOcmIa9UKwoB4ygwWCjMhOxsO7Io1jbD/oqYVZuqDAx
D7zQNKUeeKdkLHvCqyvZ9ktq3L1vMQR0UYCQQzEvBH7/aZWQlo8aNBJHj+62MtnA4laA1y3vozCf
sfpdI189gmQqeUZqIDglToXEN5+ynL9l+eY2vJEfIlg8CtBWDXupmw9u09e/TYB/ADBZXV52qUZz
Me4SRAwtfR5CxF+PbbpnhS+/AGer0vocojvt5Ct8bhp/BKYixUeKHFA6TlpMzexLP/iKZ8Vw1itz
ZQ2VoTH0RuuGiKJMJgSyk5dwB0mKU9brM0P5XAimAKCFIUrBkzYdq54PTsBhoI1qPmkG8ZA2CWgK
gobv/+WU9Aku5TVNj85fH1haRg9w0LFl5uqIyWTrAcEE0aZQNacwlZjE18nnuET79N4eVmR0rqw/
+t/YjqNSN3H95QYbofI4+mNPQ7HGBbc0jBS1CbxXXSJkm2Hd1o/tilWwcNbjbLQ+k+zkQwx2XLlF
Kv9g7zKrNnuEGhlZUldyCS6r0ifCV0zZeFoBRfIpTcTyCluX961cnLLuHt/vzvtSf2vOf3SBDndH
4+VJbxkybICBbiCXoBqFqegt5h/I8kmHBXpQm3W9GRvN035KFJ+NY41QmwIJm4Y+jUz3Q9zol+4l
AQ3wr92FgTQVqMHnzAa55UDdOQhU62Ga7KNcqfMMGUrpNFqJ2ZyR3VuudvvOiLlWzquH5j660L9e
Hkh8CsR/V3Kf+CFzCPasZGF7ANIf0dpES2bWJyBQlhk9dLc3BnLbt9rNB9rY/iKTeZwR5WCugUIP
99t64UnYaw6ZCiQijSbhqZo9bM9UoNECvJdTAU9KsLI+aWwFxNo8/W7SdfpjoiZZz2S0xy1yIBm5
nvBO1v5Oe10t8WFdyGgln0UFfJKFgdOBrpUScWDQ1S1tyv3IE/LPvwngyLJVBRUs1bJpgu9NBfXI
mE7c3koUtL0bsRDLhDF6lhCcTnPv7OuAQffLblaXbtVOKvBIV90ZNqr3ZcZZQ7jtsFeyAOwYwYhK
RI2lQ1fZbo067Fz2BtwlkXm9A5y+hwDc0YgcBO1zca1b0T+kxY3R9WRWdbT2nydQeuu3haFYeO96
taE/V2cngtBIbOLD5D05mhXzp4jYuDXsOPXYdW93XTSe2PMef9edDvGAG0zX9J+5vyZes2+51+z8
vhp7s4zAGgDPZQT7XxtjABIsRNGZJz7WoXAKJz2H9UvyqjrKucpUfydNIBLTCdrH0L6cZ/tqVtcq
1rSQVEKRrgUbN0mlqpjOkC43N4KICMdj8/2hV65+Sc9mvJy/McOZAm8jvPTUR4ZrmmbIPcb0mK70
zFnb+wsXw+EuTtAOmqWEXmo4Q2Q1Cv4zrIsVADGgVk1Gg3ecysm+cT/Ara3JHUYztKR8NFJr+2f/
X3pQJgvbmwTEWOr96x0JUZrylwvcqLhvbU/FqJlTwcQfB1tqwVn0r0V1blptniaNvN45XQ0VSxib
kVF3XJ4dGGWKDFrNCNqUWIWkk6Fu0rxterNocYE5pDCkJ1YwqWCQ/lVVplV6+wCScDpsaVMDzyVM
yd5T3GykWyX7uKAU7FRHET7rk7gXcDBX5EuaZ4SaAAwjAOFOrANwa+KyeCdEoGsazQuZmzAYGrOf
15ynaXdaOx5uD+R3GaM3g4sadsRzzdGo2IwjNdD/119dRuou9cddYUbsCYxHwh8kIirdBT3NfCls
wp/UKSHULnfmy+dQA5ZZX/je3qUt9RT59nJYxTI7spSA0OGgrreRjj81JtPqOibevAwwGDZr0PyO
w5wVR2BNA7mjF6GNQ/xR3ts1Y+ktmNKD4QZQ1BPyZu2lj1zzVqrhCU/uErxV/m69iGt5YXbqplfv
n/LNf1kD14EKwWN7M8kcWajbQX3jsq9Hk0mB/K9InWQckasJIB0fMXlt2FrIMDF5/FSiZ+Yj/92a
DrCaO4+zL87cwO+0W5raAuDHAxHKRS/hX4SWtKpAgsAq/FZJv0f1tkvibvvNn2i40fHvaQpR6EDX
URjP3lFYv/BUHSfbKl268oEf5cDJnTv9zNB2XODNCKW6sUNdisiM/w0sn7nysYsAHmWS7ytTvz3n
a4bzGSOG9vlMCRqGf8RHkg0DRA/QdpqeA46ZhzBOywTQmLXa/5NCCfSzQ5mpIBIeiR4fEdYtMhnw
wYV4tBeQqPbaz7PrC3o2qjosfinAdFK/CS6VnTztYGZmJoos5vc2l65PUXaL8lvhTk1eKwIDBOyM
qTAKUWPbpkfZa/r0AYsnZ5R2L+hY5WzQxxKkU/gS9BGKZgx5m/LJLYiYoQ5E/ycyqJwQW3ZEqJSi
zTpcCeM84jXm5BZPHy21FdHx7RwJprdAdKMctkibDhXIKTuHvL8Lra74IXFsdPtdIYKbuFlxH7gM
8rS2HGuss4N2T3oXAgA2t5vKG6nTI2fIzJSspnylWmr/f9mjMxRg6shybbOQEuo9wiMC6yn4dbFh
Iv/S0qSdc9vyWW7Y1wPqgXaqH4gDdxCaFLNhvWr4GqeEJJVnmQpPw0XUAJvDoAN/awQ6X76oQlEH
Qd7h3ab3cf2dw28rk82dhZBppae1wKeC1EYzfzEeou2BJGpP03oo+WFxQK646A/udi6T5jf4kPFr
DQNWz4IJixVBT1dSFxpZMnF+bWHWlbMYUtethiHfyP6PxeVpMI42mRz3aL2WbgfiPjmQGWQIfW3P
ZKcI4SHRXWp9lGb5IuuC5F2Zv6oFOuvx9/E40VUXsEUolPSoG5/bMZFq8jyfnugRwCB16PXO4nPt
aGXcTEtrx9+Ys1a+KiHy6kb1H3yNrJ20fSNXu3ZwrZw8Ztpfu46GpXGvaGLB/fNKmUnr2IXZM9Fd
u4v973qfKXNDS3OW4/IKCLkvwnXWxRfV4j+dYptbHCJjq8lddazVb3u97bClWefpZVGozf6mdiT1
9YoLQxBQDWyNZo+qEIwAxBZqtQPMaU+tRxveS48JDQZEQEOUxn8p6C0i9fFggyaJXsIUOgLbbUtw
k88XG/YmYjXN0kuK/UgS/ciV/cTcjevk2eiOUuZKwj/et8vDlsj0r+6QUk1KGT7O/yjB7aUa2A9d
T4Z4TRIoJim4v3aO+b5rHQSB/psZRgKp7xLJgxEKVDYxM83WgMEs0bDhltG9EXbTzKb+VrAwFSfP
uZDsp/7NGfPYtmrX+Tt95IbaxrzoR+0WrmGSLVucCxa1fzHsr3+o3eO26Nop0Nkd4dIOYXCfjK1j
6Lqm7xMRNGBEQGp3OSSOdF4m1VXFD/Qi8gGcRImLZB+9ZIJL8oS1pNdwKMrhaYEUxKTkqGCrFjMl
o+aLnSpRLx+tJlWCJARk4obMsD2CQKtw8I/XMQ2fYysSa/BcX9IFiQyVNWaWQCAntiTJEqBuuRMv
fKQvmrj3B4kFC6cqyU25hGnPuGJm6li9WcwJR404YzxY6ceoQMfvwYkbqVLzdD3IKOSK3bgyKWAA
zy4rkQJ27RWskK4Ljl12A4kcodPklkRCCTAFZfRm2F4IeRnQ8yQYU41liCI0SmQB7binWQyoofCs
rA400Pxb5cH3qc1aSpZsK2n6KUr31yzXv0njC6B6Ks7Bw3o1N6AwhZ//W7JFkBVOMDqrWNYGuo7c
qq9O3Mjx/JRF319EivwSAeIT0NMiw9vbDl9rXBe2svEcBKZNxhK7mVJdKtUqw6Wh8QA8kGfmVkCW
x1cBWW23/zMt7YDhU4vbhAHtZHkUWk7DBS0vNYalU2xAwqhU0bF3/eYI7qGlN6AEo0CoOtWNgWNR
XZ5N4xzlqm1N753kpwuf0K/GQiCc/5CHKpTRhcDnspBPnfB9sbds98HVCydQt51IICYuIW75S3/T
TQicUu5Yx/VznwLCDrvOXwnKDRBO+LctyZUYlKFIglF3+FWAicE9UBWGNVUaLf0T7LIPysHbX/rQ
rg4BDFSytOLFizEqW+/ZLMTAAF7gRyI42XMk1OFYoLoL5V/iTXIDvb4HOOoPMnlHW6HO2+aG6i1Z
xU+yPSTb+6DmRjsG8Slb60smgOUF9YSIV9zCaIybPDkJWQLyYf6wGJ8gcjCaLj4nTgRXrRHgqzc3
eLdcZS34LdjLJuxVJmwtuxm9yMIL3sR2fnhbfXXI4daxPg0bbpLZuxUFz1if/jx3cVqE4+IKMcvB
e876ewm2eVQyXZAxHGJKRMU0JIxhjFQVUsd8+IfTnD36eBr5Z+zbRLz6BazVQnHMSHb9IrUA0QR5
IY3w7UhJdTykFzgu1ZJtwWtx6hzJuYJq+WYW980cdgL7uIyyBtVbUYbm7Xb3u2tQUEOrGJaQL4+I
avoABlv32PCUQLLbxtkJ6attWgkwxMtX9Dih+LBJB9fGF04kOXVCwdFvgmVoXKHkXDIQubUuuM3/
UDzSXhFVPqpK6aW2hFWH6KOHSMDPKnGI8Pp8H1qYTZ1djME+SdbPC/cbvfov7EtvPo+F2TpjAsDi
C5Ql7xG5BjWdhb1Tkk27fCpYwmh6g/xf49RHkUfNgVyo/Pc4DM6zFUCay3nm/CM7P6x8qa7A77UT
QvuFW3zrUmW+PfAfiYwNLrZkRdTYvqoFsST64AB4fYdoDU89eumMXpE4B2wA2rXdFiR+DxMH5VQO
mKVgUyrqQoO1x0/7D7g7UStEDHHG4wsVArb1Gm6X2VBVx23UGDIajLvGjhjG33+qqMGHesZDqh3u
HvSX6BG+LyRVS9G8lh5+EuBaaoxgVyn16KW41c7CwcUy7gKQKwcbI3xGEY39TQ9R7NRDJBERObL+
XrhZ7Z5ndFZKAQN7o4hC1caHdcNccEGC2G12XzNxlEY6mClSe8wn59JoL1uUKcV8aICeo1iORMq5
QJg2joA21vvuPUoIs5bMGp8N1R/I1ggRFsA12BBMei3M0zovUgRrrkbWXRI9iLLAyW9ueUoPw3PK
gGrN1unPLTWLAnT9VYfVQRqpAsh5s53TK1gpupPS2Zh+eNTe8BzL6xRtfxaiw8RHhQtmwIO99QQy
hgt/9rLSQTiWtb8GThioPzljYCPZ5iEF6UtmudoLi50d5z+59FYzEyL0Lwskh29CoZQimPPEizVj
amiVOPFuqigFdEyoVkrRAVFm7Ph6WcIr8sa2hv8vmTZ3JOoECiIHAeXLivgkuJ0EBPsgbssC3VX/
8/lfn5GwTCUpY3CnNdfM5DhV7Hx1/2WLWbbeMyIShjaRN1sXKjpoD9QdtkJjJEJI7nkb+D0tdcS8
/omtnUARw+ojWYdjkV6kXt6/JtHyr9uN7RcPwIZKg/tcRI19t8cQehm1McCGbWIxmOInl0eHZ42A
Yxa5u5HBLnczlURZJaxjsauQ+nMvz+jlC9avakcJtLGoKRmiuw/OdttQKct3FsmkqmSOUHaWHxoU
WaTHGMnzQcGcNQZXH+rqoXMfWzTAWLLYyjJa0G+tEWBLrEC+y1CAWUdANyeNK30d8vBtOtFNYz7V
UPMBQJ/Nx5VE7hNTJEu7CrKEMweSm9QCsTjy1uLzgFl11L/LjpgflGQoFn4GGGzUzts3L5B1hVbR
6I8wqKwQYmyFoswrDbUNwkZTN5XA/8SGhJLgbOTMPKI5DF6o8qMS1eP7bDKMojV50ryKdqoMyCpb
A6nHuDFEJS9e7lp3y5X3OG3PdEoem7bCEso7LrBWGFy7fvDdsjmFrwvPKXOfMjvYYC+cZUPZxXJp
n5DmuN3z5PAzQNb6NSAh9UgXUmJyynA/KZv4FnPfrSBlEpFAjHqZqvLSKc2JPhTI1HFtf+l3yQh9
ke/aJcMXsEgapc3nGzo8XgvODe9t6wSU7lsB+N1hny2TJdmdm7LBigWpCoTykqPmobBAIiopPD31
vaOyphl1XxZspx344ygefeVBqCQunJxytXdKoDTVgkAIfo1+VUeiiW7EYoxwOzGN6yiAmSwiHkqV
AQds1uIjyVcf/XU21fRnT/g6Q7Ioai0EzTzYwfKinhf8z3Ymxzi7U5uB5y4w4d3eU9c96Ap4ptrL
ZR3zJ7nf4SIezYFKTtnogrPRtvg27rwBqWrRSeJFDkBvMxyeV9VqezHT5KBC7Ij6GHiKukm7civd
wMYjhM/Eq8d2LWFQYdxsSwIKeQRg1zifn8Ffx4IsK+11rXS3GM4h61YPAE4JTcSQBBpG+E7xNakO
+j5B3D07OlN/bxfkX9FQPY4zkoIheD5e3fLaXzm1Pw3chpx1Tl00F59rH1FzSVA4LkCZnyZLBICB
Oz+fRRuqdzvMzPkZRIc1x95Std2fHQZqhPesC85MVwQFO66vHr+/XU5+LTCtiwsM+9o1sUW/IArT
OOLqU0b1IFqalUvy4pjGXpVouHTLn4MmcUwZVVAXd8jvQJ1RUd+R4vEj7PG3hQgny6WWu3r4J0gD
8NstSo/aayDXm2ya7qWMiUYJTofQl0lT9/aAcZsQ+xlG9POQv48Kzdn8P/xu4O5S1J8HfDZH2ok1
mGed5qC7+TPP3rRFo0h6GXUxJPWD17x/68qZqDVhevv0Tr7tR3rZbWSS2FgV3BJracMobE45/BHj
yvQUf/UC/YYz3vAaZHMgbYwFZCqmtHX9Yr2mOn+cWiSwDIBnqAdFVjilh0Yh2yPkZrYzDeZgdHVc
Oq9K1Aj1bTZcy3wexaw6/O1jc3o2cTuSfAo6a9LJ8xWCaj6Rr+ImY9+gXdRWQboLakDRLjW/dKPv
zSf17clf17str7USQTmE+zi8TmfVr59cdXA3C+7RYEncMSfRA2KquAmSJjdpYFDK13KCRjgyb1tw
IPbQ791KQSDI9HZDQ39Tx0NzG/m9kLLrEm/RZniihxIOaeXkqO6aVUfFqaBHZLGCyMy89ex5D2DX
v2mrxJvh6JOmTDnfWLQfuIivbbDs5x4+e1rp1dtYPWRqZ2DBIvA9exzDKaKClVnxgHtP8vhP3emo
XS/vTD2aUtDfbtwuJKzhFX543Xc9n9wApf2eDOVHuC7rB4gQENyhvEIJ9QBo76GyprhYnZPuNSi7
F8y1iUG0yJW6ZPqiL5USWt1mLFJ0eeTFLB2lEkz8L3R2wTBAlGaEdNGuJ2fMoI+p62yF8eO3jCxE
sShSKaiG00AVMhCnMCczIDjs0uFHLsGRBb0+s2yyvMNWBG2i/RFZ5uwFttmcOGpFVIM36lT/Yalq
SBKQOr+5pH3QSn5B2kOwwCaNq9G8EtMQ3DiUbmRXLtPtagWOI7SkfX6NhuT8vVpW0K5ZHKwQY6jb
C7Jj3IYnDq02bxQFJ8Hkbb9kthjFCtKJRDaJOESjfNrYKY23tT4VEYBjfwj/TjuRpl24Ru2bVarg
4mrBd3R7NJzrlzMPGoLPTI5HZJOG/zitAmOp1bynVizbBTqudaOGYXa5/WjdzobAD2Bx9mCiGYP9
6V6Afh3C7ZQNjWpjEZ3k3nagwAEGC7GCdMlTcHh43CTrBmn76b+50u/489XfPDt2u2VorX0qLtp0
8gnP/L5PGAim02r8dmCniWA6dAqWLt4QCEoT/8J+rvwMLD724k+nCUS5XUi+S7EJivW1IL30RqUm
g/NOMWagRHE2ww47e8k9I9fx4KO3z4p4md6TgB7eDHdc5aUgmMiIX3KaadymiJgkTdzzF5BeZlgF
NNZk04dQ8/G4r/3HWEcXcxbeQgug3v9u1xpSE84pk1N+hgyICg2MdEw9xjIzEhA5/D1jZvSCNklY
sgZSJMSUYA8Zkjpfy2VlbeQU/xC/lJPY0h+ewsj/h1aI5pS+zytK0ZHBisPOcZVtzgYmBwInmKNU
JT4I4+oupkoHZAh+Cx6LNh2suTBHW6gJisr0JadY3OM0uNj6lqDegOg+mIV/J84/eSzo7X5py5sf
WEn4Oa4uWN4KTd8bHGzZchTWjpMtTgD/IGmZDVwBi4CkEdrx7On75QAt6qM41JvdjM4+Ocs6OMdW
gs/ad/BcOyhmR4OyVsOEOblulVLDLb9MeWf1RElQxwVydpsofe6/GtLHSRgEZAeS+sp5Y104M+A8
utKePGIrSyGAfr1srOUZ07HykmaHId7c4OOm/2pur63zTJaf2bc2Dvf15qF4y8Rh9+u/mZG9M4sO
qHYlZ+nNvwgtkIf5iIpGAhYjkNhJ+054EHPGGS+nrXatB4+S4Ry/heabDd8gUcIaQRBuJbbbq9+x
g+MsZIIunWCnqCkrgWNpmVhBN7QIAcJcgARlklkWqOrcGtPCkBsuWCroTPo1S3DmLtLeNOtdl940
FCLbXxOTFAhJT6wP1GhhU5+00Gv4UHh/MEC8IPxZvspyZxDEb/fFqFDlpnKmYEVr4n8drU9/xBhU
lnLEWWosjM88k4WbP1lm0X5PFsSmLPD6dlUeUukAEFMd9XNh00pIHR66urZVj29MwNNTWekmnYhw
v6GaxM81DJVFy1WnxVmmYRSNOXL4wW7MyIrheUYHPom6NFeL18uqz2R0c2g6lVGMTytnGGTzD6tn
5Khsfg4MRAx1Fl/h1VAjYfBTFnjrSHFwShst4DvEzorb2ZuPnZOcfHmglC9yKWjER2qECPt1Fplv
ePraq9IsLBxkFpEgCSg4mcFk7nLzI5DFNveInGOc1yxFcYBZcQifgJgaBIY1exn1wsb6t+LVpYR2
Fs9xqOQ65P5GXF5REge4FhmprPGQJ3yqCbfXevWST8Dhq+Kg/FOKsenJmC+iL8O83QOUhZzX7d8p
+YNEi8UUtr3IQxN3nOwPguqotuBD++whTRQVPNJPD46HKu/RgY3dT96XfDYOj2OwGE157FKFyBz1
9ADv4R6LA9IlzIs5uIW6wtg/o89Dlb2qCECd3yVLST4Xz0wmLI64v+7feLMFOUFk95wf/TA7PYOE
Js1it4tabgeEcwieCycbyvWfaGfMQhIaeS5aG2pSjTkNg+aLhJJOfHO00bYhIYDV35yqgEKJpf3a
cYRfIb+Nb4fVPg96rViJUBhXYoSHGNs3ouZ+TMVkgOXrzRpvSJkEQjGAGSlWVjh/z2HgFJq+bMR1
F64bkAQK2I9ot8bGwBnTaPpzRYyWWa50zIdajWDcloe9kWybHh7AOb6GHolXIzkxcew6FM+YHsyh
otgFhrWYZUnHEpjSRGLtbsYmUnZ4PadvarYEvS3qFXlGQcqBVDjWzpIVn7NGc6CLbHF2GHCSjjwL
nfcfiWhw4SOG5M+/OJy0TBIsvwRYQfquG2Yy4BHE1VaE/HCBHx1ppcrX+m6HhatyyC9el2EcAjnO
6Gf3293LWzVzbuDHlooOWY6z0eEZ7lShja7FM4w+mfH0cezg96W7ikBWI0QkOzTaE0EVA8DpnZ4O
bUdQxHKKZLUaNHoB6AXCSWGZGA2zmmbqWtICndtY3dBUPzQ1jz3Qa8JRaQYlYTMBwZ8lltkKo16T
uGq/cemIhCfDHn/02jBXpJ0LwIl88Jvwcdkg5x8V7qTW30wcadCfuzO5yAb8/o2bh/XwpN9XsKQI
Qcw9Nf3C5PVwtBLHvD0uAqhJ+T5g5eXtvZ2fiOOS/RNS3NvUK2NKqv+GBntrhe8G/NcK12diMhQW
CTR0hgz7HPl2dfHE5Oq7gdRcrsuomLCdcI8MmCDMMmE2x5NAgvoKUtAYqC9eTSYilMef/7UhXPLv
zNRHL/nEdCFHpl8hrd0Gg49owsEUVmJxoHcnTKruSFujoNDdRbt1nHZxU1nmVXRTyPxO+o6pfnk9
YXE2ZyjDdjdfDYejcvZmp1TazR+rSbYUy14q3eOcMsPvANG1PHOoD89ii2pWsnwupiNJhRxrsqK4
ISqltQ8InFxYl5elnNtjMuO1AQCyK0vWXHCybWG+n5j85jzVfbA1ViKhYcU+6P0OxfN2bT+A4UY/
WJTblXsXbFiWvA89GvLzvXRtGm4a8Vt3nyiVTbdx6Ck2M2Yd2yETAKZ0wSA7mOdr7N7m787Fllej
0DcWAyfMSetoPLlLpuKcgFDzhh6jaAuNvlBAbmUu4JeD6FDbNv5FpjkyVw4+o2PpeJouXpmO9aBj
6S5EiUhAdw90b4UjdBdkBgobip0MZJURBqoSA0Et4p4kLzYXCRokjDtQwS9LoA6qMvVbBhMIUiuQ
6G5V31o9oEULATT9EVasM3jfp205diVFxI1oT9dfr1YhHgaV/vNGNYe5UP8T0705hhXrKmEGQaOX
i5yJDVuuu3FJbejRzTo/gTcXEyzLTVn0evdVYG7857ed3YVkMyWGNaO2+tMe2YspMN0Bt5gpSrl4
CQshL0qBOxDJsSGKtNcOxNzsqiK1YT+HVXZwj7w7RtA1nib/cVVDrW55vFU6HwpBKyBKDnv8tgaZ
9tmFVv4tuS1d9vdgtyzaCD2M7/j+HxhIRIF74GmWsKZQ2rI4KAfYjLM1fHSOsfJIEcFcEtjXhg38
5j1ips6GXhpeN58FSL9Tht0KVg5CmtXGc/2eY2UCI61qv/rtTCHcrNF09iiW2Eq4rmfeqDgxaHhU
fOHGGt/UyXi9qePg0dDGxHt44qHeUiFPpT+MZ9e1nN0nmeR+PQm2MtPAU54LLDIiQrDyjiIcydkb
+i/JsVFlbkD5Fb1sp1STyVf8MqjrrldaQctlEo9Js2FvXLL09T2vnOOctGdHybTyoeSxy8J0h1Wu
wczZczbonzgZcV0NQ18Y9c2TOKXjJDaxoC7fh5d4ScTzqbNysqOZbQdOOwMDax1ddoVK7MZEMJ0W
PUcZ2njXcabSsbw3T2RQ/rGZOV/tl+DA00B3hJwSTHTkDl3kYbptW2+rpJFoKZntgyx8JUGW1p/5
WyBXbMEwoM72UfUlFzlhl7JMTLFRUePv1P0N/nD8/bbjq82DxtKXIcSwELQSOqLbCmc1xWlv8aXO
xiE8Pf2OD6joWH8dkJvFTrzR+soHGuhKWvM4Us6U/mQ0d5/7tx3ZqmSbkKRFgTVgSHLxwWjYkcpP
sKbHfWUP1bovJllzNn4Ly4fboBpb8ly80737KfCQpZEK6DSYYbo6H6VrYLO2sfaCnZzXybMzGtJr
kwbAaQbsabcerrSO1+MKVM6vQjSrj8bHzsnWDZo3INfVhzOvV9Hq1I3Opd4RwoiDp8ZLbmZ9TQM6
ib597cRvN/UVaV8yWC1fxrJsKrPoCua7iZJ+Mm/astK/dvEnZ08skbaufqaqUSkXEqKebfvN+yEk
Hy+99im8t7UcoM5XzmFGks9gpsZRtLNoGQcr9sp+Te7t3EeqkEwQhvwiWW0SRzo8EP2S/U1ot+24
G8GGis8Rgm6n+8dz6BE4nEp2SBYq9RoeEGcMUla/jcQyp1XwyvY6EIUgd3zHuHSRAMYgcAAR7dMr
qMwmg8B7e4sTRWPRQhNKSJhzpfk7fyQ7dBVyDs2OUbqUipkiztdvBq9QAO8iUWNk4KAscrEtXhzx
zqASWjozy00PjOcsc5Hz2DbUlu2+51tMm1weE9pXHOgxbLsvGgNoxqPWWVFlid/GgCigM4HvLlO+
d4ieyjz3E2t4U3nkgyv5bnFvZBVziKxI1XfgoX7VrZMAffBsa4llqRIPEYvXCEtqbG4LnL4eyXNF
5e/Cbmb1h+mEY9R2A4FqUhOxRIkEKRJ02UX+Cp+C4myeW23Fn77m5CK0E2T4zCu71i3MMveeHOg5
j4K5AB6aUlu7P1HV46Y6cjfk5Vkc3hUdUQwu41LfWsNkEx20+MwwpX3e6F0D4FIgiqo6XUURN+pC
YTZgDzPllYtrlO9IBVq5d+gha7XfA3RAxPean60cicjSJv+vGxpFVMYc9RknOi0IOSw+ZUTpin14
Y7aaa+aA+EVp5gPsKbwKg5vqCSjmJQw11CWb1VIWzCMrw/EkfVrR1KGu1ExYozrBKy6Vsgx0THgc
0L/KoeIR/vtsb1FQn0Jdv6smx1wJKVXoatkDLJnjprUUS5BQ5It/BHT8RdeHbVvSGBuaBJzlnIEw
6bfYFpyX9PobLpbFaM5b1m+YxEowlgWvzdzrZX2paWaJgF0ywI+Fxisbd7VwGJOIr6Mhgbrwq3D+
k+L1JFPVLupHYCJ0g9KTFhvvDE9EVURBm11g49Gl9r9A4iAYoW1Cj7KhGtzSE3yThOri8ZnUXefp
wSeligE035pWjf7O1A2MLeVy6Y4c9nZJKpUZ96O9iJBD+65TWwfiPhnCyRULhUXaR8yhS5f0iVTd
fIlD8KO3qdxi6nVDm9tHeqsq58TTsjOmTc/CSlLp5w3TsRi1vZ0UyDgjj7M+fNylqQBHFP+gno8U
Aq9eJxRWyAmyY3QHpwPH09b2/SeyNVeZ/v9roKMu+Nt7OL8DGBA3HsiirbRhZLam+xs7ExPZqpCi
6Imu1+WSMN9kuPow6wRhrdbAxZrcDEwuwTHiS3B3imEXMacM15h+QgCDNCQ6/trtInfy0vmFBQco
7hbRYF9XuXM+b800FqFlQN/knQSVgPaANoJEPuoWQHPKSZa6jZgvK/c6XJMCC85Ku0XWJnmCFr/l
pO0YOiMYC3SoRAfrSIv5og7nWy8/JFo4Qt7AXlbm/Ri6dEchS7v2F8mHoKNNMyVACoBrABNcHhLe
I3wNx1SGekcLKxV27zYyri0Y8aH//VURnyBmCYHsImnXCONGOI2PgWJIBFo06s3YeBUt3Tqy+8Vl
bAKFSPhwOT8Y5JmdjRNLxFOYOGJ+nSL+oD6alfQJ5mwLAA/Nd3nQUOhKM5WM/sWnpzr6X2aJchmp
NhArDfRPBtUMlFoyWcZO5KxYh7Gn7uYxK1FYfAMDNWJiVcnRyI85mHy+y0P1QL/No41DNPZxAP2Y
sJmEAJkUQ2lhiV07cqOducrQUiTPlp0cjMuj4xQeImkWscHYtfdP+SpcSt8S7dv4Myb0kSSqVK41
V+0EIZxpYQbVM3kDW4iOWlo9bIWpo+aUfEuODXg0ZsNh1eXcn2bl1SCb448pziU4lyOFgoHdT2u/
hYwHvNj6kicDFEs6Ei0emfu5tlL3mz1BydRex5D5ZNgx5krtcrDEhUJ8WjMoWjyFKux9pY55uMla
HFaFtSVEbOZDujBX6PZ6AcKla9wPJBfcVodjecyzae52rZMb7FbFFP4sg1XSkTa66ou76olXehtS
JlbRKTJGwt7i1SagirGeLvla6zwECh/URpX3fQ13be4UTCGPxekugEhjCP1/AfwgLSjjekNTSu+g
5qYEdRWxAvoygcV+/XKJtG1YzDJGy3VCwl1LNyk56EPXyAHZd8XbAL72yuHwSWbtsOlQo8TPn3K+
RvFYGFT9b8lSw0ZwmzN69oByjHMeBDN5tgCmk7SV0xLTNpdImsauDe8NoCoIhApK4RSOYtqSdRvs
pIXZF6PpUy9AF1E6MWKh3ZNT1Ic0HTcMV2DLzC326ZjyvF02k7u1pw1OjLy+FyvvdDjrt+Jw8az1
6QaDebQ5ZRsYa0XW+KlL1/ZG2de9PLpp5y1F/di3zuDa7a8cbxP7zbphHywgophtKjIg/YBsS5yP
hGDGadCE/mfZzvALDCmk0bggOckPjc5Xm8qPEDNn03TGez/BDJXuKuvtFVhXhpMGSAQyTsS8Wb7/
P50mizGpaiXKGJrNH3IthOAB7x602/SbVML3bdB5hr2hVhC7rnqD1CrXpDTwDKHypJfqVWph+HCG
lPH/fg2sUdPLM+agN7Ouadh/ElQ9ZkB6u8i2zRb1fOvHvtFtwhUo2CgtyJd/Bs+A1qj4zLbdZzUe
TOHS6jSkv+0ta6J9uWFYIg/WhTlvgvVa8BCUbnYd0KnAKu3ZyItGeNsluz7msE8ztKhQNqYSc8WP
JKS0fcoGvfwGgfwRJzL7Bn1QPwpZ0qNlVXk/CidTMc3iob6C8UTe7nR5lW+Kvk2wz3TmY8JaBik+
Jh7Kml5hKZjg+6MLExudCLVwTMjVpiH1ZCd0A+RdlR1kFVCN0PAxctd03rR9bB3MjKldoB7q7G0b
by7o68cU1JtEdb1xng8pacrQLRTTrp6Gm90covcQfPFWxXVwTbb1IHNCG2mlN2aep4fSUsiRiMR8
Jnk2ahXPQLfnsvtViAGZLD4uiPxkmX8kCBm7tRjmmWvaegKrJNJjlZdSeuXR2uBUurapc2OCHaq8
NQE93HDZiQCx3mxI1zYJDztBio4WkWlfApgLwPfIuNfiyKQrIGrH0G4adMB9zvjvBYCnQV4Cxttt
8BzLiOwMeEHTsgby6XuBn6eKdlqWyUw77GV5pKhyRjjApUF5d7/CwxOGUzAFIbmTHo1Jgwm6YMr2
cb0kpYNlebeMTNCLT0uloK7e+vJuAMOGWt8kTUyl4aFnKIm/N2WrWTUBrAHDoYope4yD3doNdNT3
4J1/su7He4ZEkPbpmJgh/ak/CqJIFppir/JPGrZ+5KOWKovkPVFykZpIhUGlI8Ti3pTSlRctMTt9
0RRwWUR13el6BVk8jIZ3rMpoelxDO8yKoEyT497lJ6/h1ZtIli1IrrcKgQMLI2/Gowq7jbeoVl2U
MVJhrsv1ImhoNHft1RZBI5ff0fKrKkKfVI0uZ0TDLSw4+SUy69P875YNZw06VUAwD3omFOS1f5jq
o5uCbLEorkjovvyOk8QbjfBdyffyUDc3PzJszpitgRm3w8P2TWwv4zM7h86cmVL1OLlp8d72/3H5
D1Nwpdg98vYtRsPwn+XNhNdO+JhWWyV04SrrCsXl4+Yq3cgrkMx3zu0QqUVlU2m6MpldDB9OVWe4
raRkvxspJC+kYe4Yi5wQ/FzEVu72X+SSdKIgp1NZmoViAbJnu3oGGAqPO3KJ5vt1Wgxn1W94FTcj
/mWRaXhRFdViFYYaHkcHkASdqBE/i1V9hyuHyWowo66ygX9yzX1t121tHLLgqAXN0OEkuAGYz3aW
vk3LklmOwI1Tx7lYtd1tqFBaT5CRHEtcdZnyKpbmSpPJAI1OAKczA/FKDr2HhvTlKK/ea8A7QZd6
F+rUCNH8YTL1/V5bCvj32JjQPXSsWGHBp4cYDgzOT5IYRNPGTt4IAIQ2iCMb23Psnk8UFasXT15W
+w/xKSqg+ab4QecneqRGHc8NQEdEfuF6fkJAxTzpJN61KeB4oX1bSyfjygvsBxkKzvq69M8vgMQe
oPKsfNi4g6/41BKIwYGTu9PoN2nFdw+dKvs/ubK32YfO0PFDv+lI/yYkkfXhAvqqck/pKGFHh40E
UK5wZbcBVYYL+eXZOfVV20tdApzDiBN7+2NxrobVG4gg1fWXVi43K2gDP7rh80eONlK/LmGnC+jD
2MOx/ktRxDPmoBRrwCSlXqdDivdWjL+9QtpbBisRLJm2bblARcCnNcJlP6EvSArcw/3Ga/BVDpyE
lgNjeOQpuYZQuoM/kvnEOUtXDRnBKzDYv/Uz4QcYjAoFbWDpBAkSgd7akSJfw8I2b1acb4gNwD+C
Zup1DSLv/MGy4/EHc/NNWBxrEe8Wd18vxvNCePeZ7k7kicyY4vuTN4SerSb5fE/J35lKEtoRhTts
QoCpxHBDfWxxrDOFC2++GvXk38y+pq2s0TLqzXdVIyDUfwlyPHdpRR1z6rVIe6WYfbf4rYxo0ivg
4QMb+aFkGSFRw5OpuK6rel8tdTnBTodJEoZ5kinJL52Nd0V5PtzBa1UHpOfbDDwPbWuGc3f97iW4
4nT+Frx5LVYMYOsQkMqRuV/IIfkuni8fKrx0cIXu2Dzr1VevidX7tVF4iu2YOzxIzRcdeZgKj7tu
8vO8G4UCEV0DXJOdK4GQGiqco2q9xsbYf9iakX7eCeYth8Hm+/La8iD3y7648x5AOeR8P720bFh2
0lTRbRAfCQBzzBkbCdsJ1uHHgrUxZXTHIlaET88QV2Ed/BSTS0yJxaGr5QrcQLJk7pJx5/Uadhlm
ggILWlwF3g1hYRozn+MqcKiPx//YhHaxhfOBkQ7oJRs9y08U1yp4NyNAaZ0iMbfQTlf2Glx1WpES
PJR+z8Hc/7tq4GGN4tk1TWSq+nflJTCv7YadqrDybqm+3xBGP1qOxUQuHXHVVnmLDj9fVk4YX7V0
jQq5vffZYz6pHQh0ZdoFhHF+N1NTVZ8c/3Ao2bR34RO67O01HuGJxUuQupl8ToC8UpU7TvYTro1K
FbPJgoV1sXpah7tHJeTAdMdWueitnIEC4BUCc2Ms2HxOdjzeqoaEmLO1sN+aO4ZHpCw+DrUEamSa
IKmclnldctAISrqAVxAJ/4qJeqY0Ma08FBc9VPgyQ767IMwL7PI0tHzV6+5h0WnNPs9zOzzpEjHX
0xrEg49RzmeBLypfqCV9VYnhjMpWWIqHWQD85A+02jCVAwSChhcdrCH/3wn9PaDvjU01IqayPljg
hgz0gUW/0kf2GcCEBr3V3Zb+b29IAhBlMIO3laanofFyYnx6lb4NYEV8Vc1esrrD4+eMnstUI8OT
CqN70tguDFgecTrgMI5db477s8JRuzx90Rt0mP656v+CzDjMp3oCRvXP5focDMdNSo85I2/xqGEs
kAd84l41UNbAXj0TF/5INnZU4c6H+Jx+T1HUJtvWVVMqScVREQbs5IOo8JCaoetrmtR13fnl0YGc
Jxx6YRC8Y0GFJCNCsgsVvK87T4rxn2hbu0uXR9smMbGydzBX0H/sN7yUmgfLkm6sNyUTDshxMq+p
QRCmqNR8AcenMHqUSIhW4kfH2yy3ZgBIzywKCKMcR4QxxYsnsgk1LSZvCuB5/RvHSUpzfbkKkaUO
TQPdjPYQLrPCv5j/+QjeTc9ERqAMc+VIK2WQjf2/hO3CEU7QOvGwUoHaQgmgPOjynREQIERKvZmM
2G1XS10Li9ykfFq1HCAqhG3cr83JtmAPAlRhHO9EGUcmGrMviwy+VRPVPmvTANQ7U5j/Eg/m5J0x
sSG7q1L3hPsCbkpc5Ns3FzCTuGUnsI6nzI7xwN0ZUpIhAI945O5wuKCNXa4F+pnMSx1UG+XmOyPi
QXtTwZM1pdd+Rd9T0jl6RE0HHMR42gVE0+RB4LfGhpCkdxMS6N6PbC3G7NjA414qfcxN3YumkK0r
uE44daDo25kMebzufeiV60JU7nBscB04UKLu1TqytyvjbvASsKfLCHnPUUGLltAehZCYi2Vm8Fir
pzW6KEGPWilCB422Sh9go2NIS9qe2vkN+CttTbypOm0vlgnZrwhd91Vu5bVH46/q9fYKdV3RrpPT
7AgxT+reggZuz3qaARfQRj1fesOypRjuGw8NnHPmWF4achamwkjK7SGxHnpMVpMHIBf1OtkJjh5g
Jh4NoaWSpYoKErKfyjkTArfBvoI5EL9ikLUL4T/fb/xHRnIDh6AxWzNk5gdfYeKf2uXsrf3CoHA1
HShnc7IqgHCGSD0/PKhEX2Zwn+VMw65buPnlONFhdD6VhKV3+DGj3IxP6Gx3OASXFSB8oFO9jJai
HxJGCsVIn34+It5Fxvp/aIM3sD24MHc48kI6MsL8xA6viP1X8KZQDwBiquZK/3T4OYsWXlunv6sD
KSUQx7F5l/vcomKXRZWcSxDSPuDlz2MsHeS7wZ0bDmaspHowgvy5jNgnaqW5BqJP3onl1kGCVr0d
bhSU29AWdF255HFEpMvk9/5FUEU/qLeYsL2M/Gsg5IDFxdywmjD8Tf/fRZzPjnmnfe8mmm2Nfnb2
8fBiOxLRZBKPMjxxtTLv4pMMKwtsIzLlckLaKWzsB28PAOtOyZMYS14pDf4vPT1a+694jd3dobrU
NIEvXgnR6bNs7oBvNq8IFDhQh9spREL7jhHrd/TAHa67nt8Qp9RRtRxa/Pqmv8wa3+rHY2xfQUUn
1ZequgzxIvKa2cSMqSfFbMQT9l1EqZ0RNpv+Ebv7+sNyhhoKpdR/q9IZp6Mklsc+yavxTXSbL4u3
nfVMfkCE4YbBh4tkF3DS/ZY95xjR4BzTHPUYFC/VQWuAI/GLoGpfEPXBn73iX6GAL0Fz/9R+GFOc
4b6Pt7W5KCLQtBeU1ZjeDy65ikuc8/nfg6hUBWy1gqRAmwnZceauNUhE//klK+K/1dzEKQ2qUfo1
4y5dosuRbBDSGmVKOpqFPdiJ0eL7PH4uZJoxewOV7LyXkLAq7JBa1qvcz1/zj7jPGAluuFgyvRmW
KloApLdRXkNCK2hjUc2ZeF5JFCu1Ad38cDlvHv9Cj04ccuhNJLMMCttt6GLZrQLCqCR1/3KFQsnQ
aIbgAeApYvdQb1gsluyVDoFyqVNVFxg53uSxzOM/Ru5tZ4KvHaFLKuyALcnNNQsyhDvL6yjZRPas
Zd3QHJVSvW5vK2uzc04qHmeRfobZ08yXqYeJKf82LKl38Mz+Rqi0iI14+vbuWy4eKbtZAWgi4IrT
lGUFDz2qdjK8zhwX+dhhp3cvjvT5SXdQCwwei/dzOm/ak09w8gmSEO/+Q0KMEhOKcd61ILs4lWqO
Y58qj/Mv3dCneG7Qqr9EZXnTtGvY0dj/0xr1U8MHsNMtYjHHcOf1+Avm346NVCAS6IjFHm+67bXD
+l+9FbQjAZWhKg2NhHUnZ0b3U7Z1ZElU1v2IqBZV0d6YwQB8F2+moNuDtLpM3HNpA06kmBkNVS7y
iwZ0/QjF/PlRAaNPD8gP8KjdZnXlOjeiRXEf/42aXELEOWWJXE6AtQjotsd5AS7jlz16WninO90x
y2rSXNxP6ZdFvGqLIAUgntK6si4Q8+TiRuI1BK4Yl3iSIODQgDugxsxkHRRFy92DyuPg1Oc1kljS
tjn6Fy2V5t0/PGq3fxraPzrQqbCdU5KuDFqTelEJgfflJy1pRgD4P0EPa5OWsRIwimSysJ6JlE9s
K+UVqJ0McQnGTZk7eoIqiooFAMjmiSwkGZuQT02OfZAdOGEG4zpc5fQllAzrbLGzDdIvLdT6Hkrr
xv/SM9iDt7jrgDwRS6zJUNI5+nkjtFVFKVMJsRTNi6FUzp5UELszTrs6fy1Q06VPZEj9JsehokxI
3AgoeEWGNh3zq5DnAXEQX2aWh7fRAXvlsGr1SssKelbXTxB0UMsKuG4p3/bHae/7nlGxWrNfayeB
IWh7IVeR2npOsSPcmaJjL1y2PAJroW+8WxIBbWEThmKv/HOrdkcYYpz+TyBjj9wN41qK+yZ5pWy9
xXl1l/GelA/XDvyoPlNzbow3x8tkKyArLUpTjXKbSWryyhEsXwv/IkkEKwlS6sq58dMe3izYKHCC
MLW3zELdT4qPHFjduQuTgc5F5OQ8Oo6xDMv/ey4Gc7S8+122heXsXjHpfZwoRn1znJbI7+g7egnI
yCzbFY8C9pSkbU64K6pdXFUBxbus75JNRd+HN9oqFHMfI+VsrEHZIV9aHRY5uCjbXSD0SLjeUREO
fl+PbGuPEJgbHPy5o5C96AY9wDuxp8Il4NKR0+yY4HBI/LsdKENY77oXfRjDXMJ0kKItAY7uIV0I
wsn/gsgegkLfiMK4e7nVoYWQyt+zoxhniUkHfhmfeSayxUUIrWuaWhO4qrcx2rBExFPVizgYtnYj
Hkr1ZDRmiK3euEPH3SrFyqyzE+92olE7Nd1pyV8vFelZaAftzYN8Hm3mBSbg1evhXkT6B1Xnndz8
lLopyadqIIeH+z32mC41RPUT8U/jL0Yxa5h+TPuk47YTX4kNTlZH7ukWBGh5Ylv6i2wZgI6P7dwE
hErXEurQCPEJ2qSbIHrTtrFDVgGcwkEOyffjQYNhqrpbGzQey+kDhK7DOA9Sl/3eUAELcmIyv5cy
rhnsHEqd5ymFSsXWhdbQHbVrpt00hmuAMhkjsrrSfTOAcvShlaTuzTbOoShzcY8oA1mSc0gny/w7
m3KoTktBAWt60Jz0b+caO8AUoEERsLtb7BBwSCxq8vffMLa5g2p+b7gry04MG1Di2AtEFh8RBz3/
phptJhhMQY44nG/5RtWDGDXFzROgEgR4mjtQ7kNK8nqP7SbPTjxgvUzdSwj54GDvX9HSNJHb64L2
1DxdwnsuTheuzvuOqN43D1yQt9nm80ggkDQPMXmNffX9GSQaaCrhZDdaBO9+ogzz+1uggUt9th42
BdKnI8yBAowc0LxB92s0JbuicDtRO3u4XgRuRV1n3SxpJ06Z2Chb49v/795cK2tM33SFlUltx94q
m5PoE5G/1xLL3tNXccylcxt54tHR2o4zAuYu+/YCCnHNqUMRdxv8ubrIhrjcvUywTvNlAGjLgsTf
L8ZHDOURxvfSdgTNZsyrgrEldGW4+9N5ZW1XphQn37StRJDIp7vOxQZNrEwgNHDT3brSev1xPdKY
0++G4D72Z1N/2oMfEnoiC0BQeuN1CSMjHPB7kJ+1dfJYL/1+lgmDkvjbR3UL2ChpUP2SyDgJvOSR
obrgScS1AVQ5HjL2aSEeqzSl0fvQ/IVASrjg3veD+ykg2Cy3w8a9W7cWC+G0yXPGiDqQLTxnRACI
/o3O6FDCpgYO98ly90TmHktZK7a5OHeIIqhwx5a8VRfBKbnv1Wp5SL+yC7rT1b/Ws+1iRNLwElzh
Eff6tPtpHaBXGWS/S8X4exs9iTQytRYY4Vquv+sw9DjPW5PXZdTZMLLgqlH8FziA46H72vwWVk42
1/XiFA6Evfd816BuCAavPcF+pXfFs/v4qtqj2++IvN+TfnY/9chYw1euHpaSrVeMn/LLOPzD7RaF
thw6ltcSVJWgnCBhXO66195vw4fWuzQzUF3BgNpj/jBj46BfPacJ5o1k1EslqZwA1dxCf7eA/lpO
69arkj99HV8lnHiEy3LPdBqzBtbtnkby0x+0WpLs47jS8YYZOaN9BEDgbFp6F+ohBn1c4c05XZLq
+yz/XJ+0wXrkZ0okdz/YoPtwQu9rGwHyL5EbZlvy72TAbomnIh7JpY2OlXYJTssqmwf86WqLntty
jXdbpNV/9X2GWdPL784aA5uEPibq8jBSx/6dFufIJGQpy6dH9JJsIO1agbLQlZ9pFm8fF3QWd1Ed
yJU3jvKAeeK1qm2q4pIP5KC6NkPfGoRWamw2bM/gP0utdt4ROCJnO6WnSP3s85CD0HeL4hvbqrIz
L7kj+e1kEm14zCaJlwKB13t8vo7JGMqO3nLtjNivD7h9QgK+SERGPmAZkIxBQHMp+SGR2HlCUYSs
+bMbCKl8nnfPKBy0Q4t8JQZ/BYkLll+tIT4AOOTvXfYt5Lizg7H4ck0ePWdYntixg9rVNZVM+3vX
WZCkVtqOHffXl+5ruajkZ2pidZPlaagZyD50MCwqUsnHV60ZwLD7zqyQauLyKyf4NMbs3JiwQJPB
vSpsgFKYtL2wehu2r14VcpxgaHKt1mGqHpCzGmBp7j522fsH5d4pT46FLbzWCu8OVqgh1h0QAb74
bwILpb0PTLGRMJaCRwMbx+2GsFG6EmaWf7q5pg7HdXgejPTy1aLwpAgKxt6Es8awYvSV+Rnf2Wta
Lg2s04FKndIIM9nEyKXtCyWOWL3C3jjUf18BFsGfwHlkNDSW1HErsDA76czDX6U3KNcHfVNmPrLf
/W58elHpOX+OszagXh9c1OSlxLl/gZiaMDxn72MfiI6Bv6nFgY9tZm/XVb3Eqsykwoiv3lV69TdM
8bHm3gU9UJQTZQtcWSb0Tz8pybXFOQmC2byVNkKTVXDSnZfxwywu86TW5EajkY7P15PZH4NDbkGi
ljYALKSoFuyeTGx8DLDOgO9vrFWv7Ea0ln92CjoEytA7DtauyINC4nDBpvge39Ar1Sc2A19eP1Ed
qgT+0sO6aDzQkOQQBIKPZA2kbOo5wD7Xd9jNglZodDxkLVd2OpBizMyaIJxo/nJv/BVEAo66ljp9
zU6LpYqSkfgDkn4Bg1ombPyOSQtSFRj/WK5Iy3dj8/+3zbgONxI9/QYjFAjE7dxBg9sjCwW59rKW
k+Qsp//ccZk9EEAVLJGgKWsgaKCEg9nvHldbj+JEAEDPuDhr2grXzfRbQqWkJa/Tq3F8TC+7rLv3
S2WBlK8pO73VfYjpWsclXGj4zE2wnj5EyJuVneXMqysUmI6xYRFUQ7/F4VWyXuxBuTEIK9W3JbHa
Gzg/NEjgtxOr0QamwpvLGv2fuHFER99d3b0SksZOdbYFaa4LVeeDJ6fl0XdRS46HJFVwPShBlzbb
KVcj9r2cnlx88kGVtWf64PBg2RAl1ATyLtuvR15HG+tUDORf7JNMwVFaEBf7uxTx0empvT0ouYOH
t2vXxIukVw7ov05yv3+6xaEeqqjS3BPZcCQpMoBsaQBCa6VSzQ7MLU6Js4tbbVIsREaLBFL8n1ck
4jQRPNi+X5Vd10nmwW5+6e0Szg+v6ckLgqmVBJMtJ6lSDZuxTvdQuPLQsvQ0wxj9FchbjugMIgW+
JLu9qmR75LtXaBIhVWJalUCh8NwLqwKNg3l7ROg4/Ru84tKQ3N7MHDHJ5Bsi6QmjyfZV1ncx+Ucj
V0n/jRUMhMd1j4NWkov+ASzct5eXWgISL7oCXsexBHJAWO7hZsSqezYf3NNSl0EoxDuwSwVEvMYV
wKnOsMn8GA8w/5dJKw0Lr8S+Ru7+UJmyfJMhMex+TfHwrbdwO9Qg9MImczy4ECA83KDcFncdmlpT
ndkxJFyPHzxONJraLCs8o4gsS5wfiNrQGBXHlpWRUhLMcj2V98xw/E9NE8cKJdjZWk8hB/1p4/5a
F6/GV1Idily2C4MxedNCHpa6ECrdjS98VUniZYb8GrXpHT24202c7s0aHy5Hie//fh9e/BlNFLFM
psQju7k5Y2VJPi7JekA9LMN7Poe5lRgp2uaVg7uFH0HKp0NdMfRH6IILCUGJYN3QcwPjiQ6x2OMC
q8R3hbBcS6pXbLJe+wdBBRggNghYIbaeA/eyo1Jybnutu3Fu9DmOoqBt0JymlyBVLbFLb9rnYqna
2PF9BgXddRrg69PnRttTkS1jZjYqoOuHkNsz+UYOFKLq7CgqHqI2mb6qy1Aw99sA/max09nAZuNJ
O3IY7k7Ql6bRhZZNqnAd97qtvKCOYsbTzKoMXz2GbIpBVYTJyihvo4QZ/y8c2jI1MxlmmV3EJZcf
z2lUGV6shRv8AzGzGiVWbG2At2X4S0USJ8R+SARLeqHVk3a0YFnBqkB+rjvwxRYfp5I0ypJ+bFgG
jCOuvhvrJX5kdGwt/XNyWZY09Pdd/mcbe93BeTzPBHRj1PFdl3IQSOgti30rTSKGonHRot+LIjrs
6uecKkdrlWqZlhClEgRo1qr7vjxUSp8OthM3iaHS9S7uj9RO+GB/tGUyHifXLI1FMu8pFm2unJch
TS2LGmRbv8//tVx5LQ/G+SCsgvzKwbvw2EEvLHIropHJKBrG20DAmgkcy+A3V5DXux3ZLDuFbBYm
xX9QlAgvw0EHCSc6Sx7/fwCh43VNmvCvnTVn+A5E8TVVOOj/mFpwUHBFSzwsXAPxS28U7nC8fk5r
qIz8iqBBm4f3R+REVAsDyhQXWOhqLPfk+m0J/M0inXfj4BR7TYopbFvZvRM3nxYdCGkWU54ruio7
1/vzPotpYPKYVV0RyBx2yycGbFabk8pHLqtMFGePuxzF7fs7WvFbNYHd4acEYonMGv/vLxQgU7zH
djiR1XbhADNReBNfT4on5wlZUifmPyw0QarQL3jxsn8KsQOqdoKxLqaDjNpZFKuz4z1vQPGGrNBG
v/oUvf1rP5Ke/TfLPyeX522xjE+Akwyf/eEmaKvU1MqJqNJKCRCKwd9Ti1ArB8jZAa0VlHhefbU4
S9dtAchd9BhiuDB+zM0VKwNDkL74cFjhk0XRtJ/sL2Wvm3J2tfRV3/CD2KWapGfUuQggUGxQNXFb
2jRnOOK0k1BNZZ8XTDMRC94X6y3HlXYDZFU+BLsRyKLswAnXLlxRoKr64yVaClWMlzaVArRW7HLn
4dmVyAemnLy+0psX1J9VfZBadSRhy0dzoca/tXZmCefeUAy7pgiCk3OiplsaL8Iu6CCzL29GxZ0Y
q9Aj0u6BE7aKiFxs0IVcriTUwuQobTb6RPGwQD064MkuSIZ0rGjKr1MeAoy/boH+d9cafqdlaFT/
ub7/k7Ko0hR9dnxNJlQRT/q0ecp4VLiL4msmmvcBHkkDlTLGbY8ZypB2Kp7AvG+FdWLbVuRJpIZy
ZOnbE6nf69LgpnL85i5mJRXleDYNKC0Zg1jkeAp3lxZcJxfD3uGURamko3oKzMzvHM1W2/ZhGNox
fp+UXNCGt4+zhexe234TWpurDu4y1/iq5mTAL2S6aInTtmEnfDmmCkP6Ya8wjOXexHunDIZMo/gj
8HpguPmTVazir8m77UvWMJuFIyluTG+P/kvqOshI4i8IVFxJMvsalBRa9fSrj5i9yfwAhPBtfVQk
ssybJr7x+J6Fc4XiSFjqiJW18t0gwA/VZP0lubyUyDENVxDY+zajYqcpaVwq9b5veOE0ROl/5bsw
kcc+PKxg3czMgdHzz9/fKyf9DlTiyz/mcrQlncHLMP4oyGop8HpALJ2sZod4rgn8yw/ccLs9lfIj
UMUmBH9fls82WcvOwClazoEvXGxBYxhusopuxUZme6cwWMBNcQ1J/7hcLaP1evY1kt7Xm5I5NbmU
PFfeYHne4WwNGsOa/e6Eijni+dd3y60+lwJKCTA9DfiJ+DQ3MVUwe/q0N0FZXJ+ZOw8T/UPlmh1w
YreG+cEB2wQq1y8HNbZ0L1hH/VzTyGkvcgFLdC60VT+b7aAEXDsf7BKt7uBtq4WygLn/zrXzotig
AxCb0EeMYg7p8tuKz/6OcMYeSy7ApPQzzLvHHPrJMZOi9wepksf462OethXaAJ+CcGm1jUhdMDlt
yiP4+o4sQdr2/pP4IYJFsqT3JxLhBXQVjfzq6bXMOcynLMxjeGO7JRBXPh7mGSt8V9WiJNF9uhGq
8SkqTUfo56SFnUDaElQgSyhxKibc5KefYPlQeTFurmxgCymPjfJW1APTBP4Z5+Bf5q5bty7PhFo5
bXzDEPjem2jDt/9r3S7amabkWlkPvXQpb1BVjI9ngsNmjqDN/iq6DMRATLKbmSjmaBVWxd3IpHwu
tTRFYptTLi2WYQbnKzu5V0RSkl1huhyizLs+HqxNHmxishSLZ3yLXiD1Bq+6PGUGSiKxNwtHqWpx
Et7y8dWEAVvwkxUz3p1yvqwKyDqvc0bew3RCSDV7k4rrfMH35FP4nHoe5xUUdBqv4s4WrXUt0fOg
ptO7kuC63/6LndRuwZnnnBPFe18NAYLt9OscBGcyvcOoRQonm7/ItIo2HmURjLYDx9pie1f2ZsfM
XfETvsNbKlfENo4/Csr1VXEhaO6SAvGYM1Z1pFDHiES31IjBz9HKxGSBNjGiqoACDbsHy/Xbkeig
bUrmXov+D+LSE2a9XdnZhWJ2d4pbZF/FPqM6aC69iRnEav1hH0Xr1nbQKTohRPCDy/nwAyL4SqGf
43t4vIYgVc9LdOk28XHPtgd+7Gsh7+MSrhsCykHihmtK5uPNUo3Tcyh4QXkuN+7uhuHooyAspKUW
5P4SaiuyH3lc3QKrwgy292l/F/KJwcUdr3E8t5zKLG4k8UCUZSkZQpKqnwfy8Fh9Zi0Bw1HmJZVj
dP9Kljo5K9hM8CvxNqygR5fUE7Y0IaWOlmypp+U0UYa4xEvt8iogBJSebAUJAjj4uDqZKyBjaogG
pdmMVC5pHIEXlw8pT2BjNiWIVNV/l0OznIqQa/y5CFBWc1lU/aE1QAc1fItXhNXXV0Rt54xLT0Oi
PsXIvllaKwwsM/A45tLLYZYhLOYcXITEkDv2SMXCQcYp3lopXiFm0NYFjrIEFICiQPOSZgIl1vSm
e1kPTXfjohv2MX9Mq3A3dcvdxuOfTe+lKLE4J7OKnHg1m8QxSJgZgtnOQatPCZxHMXCjhpCwrrId
MMONOJVG8EboqOPsCqs47MDhnTHMGJsIqpl/+jyLx3vqlgHMti4fIiCF3DRCpG0BWh+fhVM5olFC
plU1NoEw3UDly21drob1wzh1OxcTWMa6pbP4kjKvfAMDSatVCJ5j9FVoclZVbj5P1kK7gTs/DPoA
7oNTjXI7zoJMWY+NC59BHxSLxioairiTcWdZD3ba61irZxYYLqiQsqVV93iRPCFdxSoamA4TCNaA
LxFnt8jM6Gn31a45521gneHhPz47EShkmPTBMPueb1vDAfnit6Gg4ZmL0VQx5ODqe1oGBORqZfhM
JGaQ11c6DX0rKHcXt3ys0guaVb9ilf9hCylkNIuIXDu9HJEfiFo4P+h/OfPN7B260/my6yjBZy8H
xMsmmNFTVuVm4AcIo+bUo2d+cNyXHVVlo55WLqIJd9wPlPmrdeg9sxlQMMF9Pew9wupiDXV1gE/g
4h65k4BGSWLGFnHmzKBPwLyAODB/9JuC+YUFBkw1nA4ctIOPc1KVPIsfdNVwMcn3VUDO/nYZGHDk
Tw+ji5MBdnHHORtGAZ8J3L1HhmBFy68PZpAwt8WkiIo1Fq/UL0BX1+i1pyTKTE3ZQ68w3V0sX9Gh
nxsBTbrxcn1Cc19SBetrWr0Dqt6myIeb66JLxWvf3wpMM60Rz/gusExyWpyvgsUTlaVgu/THfqvf
ayE9PslaydgiI+1/1vgnmNGclk11DF0Mz9L1BAg9myqwdIepDhCdkcwplgjxGkQLqW3vJ5TUaX94
dSP8G7B2naFjzx3tm9vWBrCr4wxe6G68tQOPsi7WmDpLJxbq/PZbrzSUFOHwrL6rzhAbwlUnpPu8
uYTjnoPhYxVYIwmhaPAtIJe7JX07p+oDRNc8tq+RlgMy2v+RsI058oYlhbTyX5sYb34DkSs6fChh
MRbsKZyKZnrgw66g8A9rCqUv22k3YmST2UcPwsKyZrm9vWQPxTioDHv3dRDSxnG2UMdvMeUy9zSQ
3byuquGM4Mci6ik+LVthdjoj6a6FDWhA86JA/MQJRcF/xvbvaytULFb5h8XlaK6KwVaPgLlshxDF
Fgi4jSgxjRV4oAxF6+P2Nxa6G8C7KCpnvnLR1BmCzBBQH/BjLQKSniUwa5pM6BA1To0tItSbP3le
I4cEXM6imBQhnUBkr6N/u+xlBlj1rGFFg/8vwFGpMWLBCp/q3pBvGWpWCUnQCn4xdOr3FtT6n3l5
Zfyr/ixrN7QUc14FcZIJYKcuk/3OQNk/24vGVulzKIvdjITZ7+QoztksPsVL2cfJnNv4zo5I8sr0
JnKH6fmaOEIxGpASnkesPxiHBIbY1s0ICgFTVMOt+87B9DNhCDj0YygT0s+HvswUbCwoQEYWdI7T
lhmctp3Lh541ufCaV8wDCr1QdtVBxdBVdq+/7LeDH3dCbTC3v8g9UmQd+Q+a3xtyfQThYdsR0xqm
hMFsuVTXMQhmi+Naa005Tx+PLTFD6tCd0DcR81TLC58QdrYyBv09FLKvkr4YCgW6WB+BdBHPRywK
HzqHF6xqZ8v3Q2rLq/4621AXuPiN6iZlPh/sgu/UmJR+FSU8qwxQ/vzq1bA/MAyvqUY5aivUOh9I
Lo4aAb+2suZYCS3e81NzFaoRwOA5M09/1DELyffmXfxM9+1mgUXsoxCZlT8kQJGsgiIjOc8F/9LX
hfZ83Uyo3oU175hAa9GlxlwzY8t6FRnP+Asswme3sLLUV4lRGrjrRiMnJlO6M5HLMWi0M+7cSJ7v
CoOKHRg419xmocWpwLYvFpqeceKKvBJNtY8mq0OZWQUGFVg8WAhMY/3c4eKud82ZZrA1+Bxh01bA
/U9caPuJ3sSQavaxwjtOtnaBhpgxCH+JmeWt60X6hLA1xswe4UEsmT64UEjqu0Iq/8jpxUQ+Z2LR
b7+z0M5qhfm0FC6zRxr8bbQwS1doyvpsMLNsILUW6RwxIlRb3axFckBJiykeiJ9BRHEhVNXAy/l6
JGSgBPv4kqx4eQcZSZIBtHQ/6TbL5BMMWC+RoKpjaffAaHQmZi/SYjwcT+hHG85scYtO5DYyT+wA
Nqqmh8UUM+dYL5rIkVafs4+KDafGahhd2D4vRIz/sTrGHSFOOmEh635iBdmaXS1lNrNWEbIs9QYs
u6IA7SQLouXOSVoOPydPf30b1MZEWbwqJeYphI/G08LNR034BxDLH2+IEQ1kHkFKkR3dpQNT2ugK
Axp33SR2Y5+V8pgJZg45Uj9STuJEILKwnBFLWDJ9akkueyZVuZnLh77kK0VqKjBjStnZnpvsmH7K
DJ4l3HiEQjD72NyIwvUnaMo4bi3Bjvf9E6w7RQsSF38dTt3gVz8mADii3WKMPhW4iqxyMxxdIV8U
8CRRm3uzxPgpfwHyD+hnaLQoClU2XFawXA3rlzPGWjMSQ4MCjg6pKCrZBcNYDucWKzzcPTSfc9H5
s1WHHt2VzVBViYH5KCnmhH3VE+BGfI7pVfEdQEolVlf29z1mXB1+MbgDln1qHcScNRrzwOyD+813
UFP1mbxk/qW9oZxV5CNNJ1+WUE+8G0CnfzBAYPYo0XuxRy/igwWQ2XfEIhgyiustBZHXiXj3Azbl
/yXC+E4YkEzwvZROyJN8mZ70oQRhhB8J68YyxJiVgZs/1dY8QngN1NRCtUI33RHfx9/wdZ5me0wB
1jWbXEf/hNgdsqYD5MjMuV6TKXIzXdmc6+I9szRpuBjBAhRM41Eq9LYucgyXirUUnIua9YH88yPi
wJLZcaVfjzHOjgeB6WsEWW74xC3pKqvrJDo6hkxJZ8lkAtasoRP2G4dB/icDMKDuHpPFpMbtPdt3
tP0rROIdxTV268iGB0Ke2ivwdOPTLzo/oDsDPsQwqSTVzaoUNCaaskbHl4P9mZIRV/L1e9N9eIbN
wPXQTja/h4T5FJHX0Ty5JlqE9xzNmOHpVY+8s8LonRFw7zg91ChBpq+Bsbt3Mae3vaCM0VSARXl9
EhoVrdtoGpMooWN7Anod9vldQ+8iba9OrOY/QcJlFC5db71Ii5cPwSSP7y3Xh36ZksNuEML6zfZK
IYhuqvIeLprpfkTx4204biafpmgGtimaGOpzxt4BWxJKQH3Mym/KBXgIud6Sa3dHjXjB+003dEAn
2b5R8vi9F7YLVhEdtD8QJWAb8vFTFaRYBWMSOKYVhnpUs/aQ5M3thZnakbVk7cmR/lzSZhPZEDpl
ukU2Kv4wC5YOFX+RUtbFin/YuIxTo9M3SPHsFgpFXvo6TdgWdLbUw6Y1eJc+zzUR7Nq5pzXHw0/l
sSLkgR/045ZYN/L02E4nzrDJHbqqXtUI+Kd+MArdvc28eg4qDVvuIzlTuYCjF0f3xhkxeZlLH/d1
wPEnH/beEmnVt/+bFTLOUNMI6PjO1Eu4CZMsPdnmbfMSGMu1EJ8AZZPYTvc4qlCGdnNNJszhepJt
sszWr8Qrwt2l8vhX/IJwSOxoFs9bFI79u+HAH8VEm7ALvKkwJ/+9EXCPidPHkOSxrcQ7h/nbJlZ4
aQjlPKv91tMaaelCpVsbt9NKuRQJLwR5/ivE9f5G1kLfou8Kyr1oBG4w8MLc/LlFaYiBxCqptOAi
RXDNy4UQthkKcsNj/zCIDy8E87bmPr5bUHbPZqonUXg6ITNBK/J9up5JYyjfW3DRtKlCwSyEn3hU
uVm42iFVgppNEuk6t+Wfu7+4GhIsU67sSkAGPv9g4UXZ4HjA+09CXB0ZN7DQddiowiLEh/hRebzP
zFlpUR7rl+huM+iu/zyq+q+glmhxUIxId5z4wPlmzuxgzv0Ml4VKAwSFBgSqtH2c5y0y4k2YN1HS
nBTAf4I1EZodFmt38C6jtibzNVofwmIxEDcD/magcTK73TOV0c+NiScM1SvUXhYvc+L7E0EuKGRs
ZIrx+4FXADIHvrdeQG46ez/BiMuMwE2ajjg6i5FLM2lepLOpN/drRiFbH31ebMZrCQcgZyWSihSJ
lQDqaDqq2I2LyCce0Df9G4uwZBarZwkww+PgWWzPBB6Rxep1j0YV/Z246fabQKzMXVJMETUqRLOz
vt8OB3ARqn/BW6WYI62Ckf1e4Z8uk7dtFEf18Sk6JPDw7qHxYpqu4MpnBKJ7XMbrj5CNTNB4uEIj
iu8FX0AZbQh6lpD7/h2Udt/ApYJcopMnAxjCTybqXrZ2BWOzLjVhw7r/JVbToo/Dvvw+T/HE1TiW
RPk+pghUohNMdLR778KEZLdH36QqzqsTfl0caXGe5hjE7+9Jrs2BKtfwKhTFeT84kdg0OI9oVcgQ
xRaZR/dtiLjGqujkKLDrHS5SUFOiTxiSvXspLdlzAh9zzpAjjW/9XWMe9jwI9e34Y0Ak+eJipC40
EOVueu9nWvUNoJazYVPceguVDET78whdD4UIl8qNYay3qIW/2p+K110OMCecAKwG0pw6z36szkzo
pTjhnjWH2NTbYnttTL/j1d/H3aSUN5NsgFR/lzSDBm2iT7db2FwewuvmtMmWLXtxitYb8uxSPigG
U6PFHAe7O1lND/cVFefyW8HPCtIwx032gzVF4kCo6m3K4u9sG5CiOCQyfoyu6h/cjgRR9yg2DrqQ
7J3TMON3956baT7xh8kIdbiY+YDrIxFVUdtEhTtwo4iHRt5zaXcOe/CdCWqk07KLbdJIghegavNj
b60QIfR2aLZ1IDEvKuXJc393xf8la4J4303F3xOMAbOdtXjtusecL4pkQJGzYCeOy1uF8ASmKqnJ
d9DJ+aGx6tRb9IrCezXEMwy+TxqKVgQFvK8Hi//67WesuCptC6rBMP48QxVPt9RB8ZK8E6NuJgis
l3xD+qUYjJU4LrqL3lw3NHp0b4ZzXPx5mdAqtFVpy3y09E+6Y9HK1Q8Zm1uMBLZQk2mtw+58kJ6x
gqUp9n34GrfxhhEclwidJUbulsvY7SDKkYe2eUvusCZh55Hth3054hAuGK0CW0Rs3ccFZdPb29m9
hnBbLt9r5na7GwJ7Pb0gKu9Eol4Xkweirm7J3TZREDWq144MoMYl4V8n1Vd8fQiDH8QRM2hAABgK
yzJBoY992a6J8J13Sg0mQOOlYW4uKj26LCJ3TMRm4rdUlB/vsbdkVFH0Oy9yxbesVYoO7UtW0aBO
d/3LskkltMocWZUyE7N0SE2DZrjsm24OHpxvLk33vtLkIcq2nXLIBFMk0mA32BmHeSl2tmzYnJ4t
kB674dybg7SkTk4tJc7UX/SEHj7bei6D73aqPr/M9GSeQ1XU26X9UW0VL4RGgJND8vCi/o2wXlq5
wC+UixiyoSetOElNuCORxL64agSsjAl2D9ylLimlwvyRitJVf2tUAuAjrz7rf33ECfht1kORcq28
i3KXuUFARFS75viFgz1l08CyCepUv/cayyEcCc4kTdeLUmNmAFP8dxUmvPrrYLXU2LfBXTWrzPGc
yigEQR6wJmP3lwJATHwU334ESRmEu+S7B+ZaSgsk+Tc8hPLOfR8PJo6dPnQucpTKa7+6AkeDPcIE
LPbDosrlk474G6Y8VMtUarxCBMia4ZIOtG6iBBkbNAIvLdaZ2xiMC3eLpM1wZTk8hMDi1qSOT2KN
eZjXxFhfAmf5mYLz2aOcuMc38ShrWLPnHMWdqy8aqU2Kvh8vWmXODtzi7goJrA4VM9jZpdvlFlCr
Lfw7gNcKZi175eBw8ZEKO11x5SpjzdCyaHCGJeZ8ZKKCnGl6nLRXsiD2dj4gtDaSXnMp5kUsF36C
UFNdPKBWPsjGt83FRcrCKX8tuySpfF65FYlz8pdfaUXum+eHldBmmT1dFLIEnj1xRqzYevJGQMGx
c1oGr7MWfAiYaZBzLp2dwitw3Y7ZC5QagnXxXxzpjtqMEX5TViSrC2DEmSKXylXsQLuwNeY0b1UA
SAQAFxp2e7StLpYjhLCpEAWzI7J2RQb4RaR5W7+w3MCUpSfbF0E4Av63B9L0crHoS+I09hSq7Cdp
eQnk8iZ6HcsLplgHslCHThsgnGcwiRTOSJsEvEonQP6wVpt3HJuxlYqJSH3kwkjAKVYSHH0BYIbB
kLwFX4muP27b74/+rH98QSHIwX2Lr5D6Z6dkRcgVL0zYclU2oCoxx4/gQ6xfwMk9kaIvu/Xl+ivH
//sbleT9BIcBNQ8eTuotHleEOM/P8L/2BdmBCk0395I0qWuL39y4EkGiIyJdRJ+IzbaF3qIWvIHA
MFArW7Y/n8nDaoVTrcdKQ9/kot/cMvm4qE5MUbaw8ueKn0bDl80xEKMGF7iMKXGqjBHnAMtLe48c
uh8XM/TQGJm5dxUTEmLF/SZ17nHRXXBN3feWEx/Q7DBjupZ591MfFVQ6/zWgeJRnxbTTql1mSqkJ
TpdR3t9Scg4HbCOBD7F5AJa4EXgOEpMyYBptS0UFczCJu10wyXouVYNZgyrMPQzUJ7bDgeTTmu60
KBhIJdS6dH8ywklqKMb9O8TxuYEfsJlXVkWqB4sUaKyUznmpVAuJoOlT+dqfd/De4qnBM6auZYVp
ZNOPPxrgyAwP7CvTPP9BZfXPl1dz3fFclGgJz/qSw7ytCCcRmFEC9HUpSioe592HbQAHFjUdTHKW
WESN4Yo9zZmIqURtqtPP3ftbg0akBtSJ2Cks8luXmk6Eg64nPB22Qh5X56X+J8ka1KnKJvQsqH6H
msZBgYyTJrVfNuiGS+Vk2YfeLgnD+mJUeJY2j3oIigS7LVMgfipoCbjF+0wxpjL0yZq6B8G4BwB5
HOSZX955ws3OI0wz4uQCM8eWFezuhP6a3hYPGdwVa6BfjAjPd6fkfrVEEr7q6wlCbyrayBVNveDh
LXUKhdQoawBU9WSAuS7o20dKKbqYun7tDgL1cD5EfvnvwPujSBCJzhNd78tHFtD7hzrymZn+gSFy
z8EY0PN5wJJw6ap2G6r4J3dPIrb7gTaGks2izgIwEg5y68rCASSJkAbC0FTMw8yDJYg7mzS4lRZr
O7oq0Mu1cHfppLd9na0p3rdGOPPvwxy+xdnzInF0QyOfhhB0KMzxdW7Gw40lXTczjwG0WdGcUP8Q
kDpRF4LfKnPzJeYSCESlBIsP0nveUGl5TBnGUwrn3Pf/48Z4Ea86FAVshYFR8TrNOQ8lTGVRM2xD
34jpJR/Me61S64Hy6LhYP+Wcvt184hipshTENNav0a/3qYC5DZJ5fH8w150WeSgxJkgr+0gJWRlW
yAgVsdW6gUPCfLUbCVyOa1AkC1hdrsVe+Wy584G/thiMKKi93vwYOgIDX0G73AEzCuUT6uFiGRR4
xTeUx0JealuGKl7E5YjZ8Saxvg0Hl01s/90ixRUXn4Q5hhxNNi7ZCFd3Hwuuuze3IatEKmJcreqC
rPWFhMPkp93qcH6+xhGL/CXFLhSOa3tD9vQSEUQ8OLF33XUYw1mZsPD2u1EMfRyZDwcUie4vXv/4
e+x9RAIIccJTzk40vImwixS5RoXe7qqiCP382LwXS0nc2ScdHQuCaDje7LWV7OqfaFkY+Fp0rCqj
97qbGcunYDj0wnY9yfE2GJNLaCW/0aIVPvNZws/P6DqR/Aco24Ut7lt0HffbG8CoE3xgnXcdM4hw
B6maz+44f5beVFaDSwQ5iOkNTn1GnUKMX9n4JlHOA+szczvVpvuYkLpKyE3O9t5QmQYOGUn7OcF1
o47mPS0KkMdyzlTJxIHQ0qfMtaNBNKZ9BwByMJYop5RWSkHyyGCPXEkOn1JOBYqPB0aSXnUGjRuQ
iTi2p1hC/KOEjawQv/HcdNUtw8laIzhqD9R3c98njT9x/REf6QOh91dmrZTzdmZF5PKV7FC+a+wA
LulYatLgq/NA5dEKpwBEvGNFW72iGQTG1M/hAeJZWjRmNdHG99Pfpm3EyDU06BaIshqTiDtqt347
kVvr8zEzGi2W0JcTd8n71QVXTCNr0hM6QABStU+teEkrWWqSEGujch0OmktupIv77Nsu/2f0LI4I
9dOcq1vd/X5wvg77+ddjiimFJrtN++j1rYbwiW3u0rQ1AjvRC7NZmKI5SiCfsqxXDzTTsreiWDpw
KYxvwvdqaHnKZgB1L/JFDCjtAqZrVpN0M82p0zt/dUCPlFyoWWUcxnVfnmoynGvbvrM0CVoMe2Tm
qEEo4dp0e+xtvlRZvVE4DqE1HG5n2oD2ygVf2Zv1reRjkSZU0gsZ2peiTQa1OYEU0BVCGFydGReb
lx8Y08R4Y92hBYU3JggzAiST6h1334j+QKzeZMthpXZoMv1IJ5pymLxjtsBNihglXy+8yU5tRybg
XAaFHu3H4NU00Y+RBPFDLBcHQSfO25gE73oi8nTcH1JAJSSXvedW1JzOuY/KkUXu2N08rQvVWFD5
ZongbJe3Yi8e18XAC6Pxu6QHj9WBUcepeXRSYe1/yiFhUeArT/NQbfXTUE5jMo8Owqrl8njpt0h5
v88snpWmxT/KQFZeDrooNt+uLyWP/Mf43JqcuzfJu/VGHt5TEF7csTct3Oe1POqVYUf0c+CJj6LV
UW9GkfSTFzwePv9H5PHNVjljqHidyN87zqWc8KC08y+zhiELjJwSzeq+cvfgR3iNHecNoPPgtbAI
C0TgWp3AR7/GEWCLbXVhj4C3TdFBc7Jm13qVp6jyH+jXRthUgF6KnFfkAqBrzOHFr4QD3vI3GCbc
kbvRvyVaZV8+Gn6qAEga+ajx4IebXZAx07xTMhrmL+6BzngLZiLcXIgz8XA39ghDxsDeTBvYUtN0
nGSlVkuz4i9j2Dobvi//HcaEQ8bgO4524X+LmlkJgteZSSWVd0eY5dZOmayxppQgy/aM1P5betQl
2RADu7DkKVZPi0iC77SGy2cH1Iuem2jtPYQk8HCTg/J4IkE4/Q+961C3/R6fywzyO03okpb+nRSN
+4H/ekbjSKDW/7j5tV1N6e4bJxDSgt3HN/DnZ2LcLV1Ud5mS+v6Vzkr2LcFuvmg670Lge18bifrt
1DzDi3pXSMm0LnqeyIjccENUd9OaMrItJ4KR+pqyCXefnwLsmiG8S1/kSmpkLXbZcltK7+6jdFDy
1urOXyjY3Cx9REUXeLkKpZ53cX0P4hcSw3J5cSJWNT5PZGQ55eCnRaC2qTr07QFbJP9EttpZ9jZx
5/8sYI0EindimdRbNTF/IEyYb1cEN0Zh6+0TD9NJkW/43DF+w6BGSc8qAOdBnGGWLOde0ONGAqOg
ic9dS3BNOm1Urmq6ZqrzxlUBEsBHtW4rFOxy8v2ZReDKwQ1dCbsgbmAOP4gqf8ss0F+/Pp9BqA5c
IJY85GZthKNya7Jya6AarpVjfcBr1UE3XQG5+zuXEYe1+uVFytbr6f7P29a01Z1CRnIfUHwaley6
PPdUXDSKUCbTyTJx8PoryxmIB+EI9Kch/6YOjIJhpIKoVkVgrhTcgfT91xhfdQI4wN+B+/I9bBXO
tPOXG+8dc9EnWMjPTAT3bqjbUUM0feWqtgSImF5v1ys3mEIQSgVlPfD4aiv3nLfp34Ab10KOUnHW
zYQStSTC5tw8RaBQx824Gpvf9JuVneyXVc3KIrsxPnxcZbFusUfT3iPy7daJ3fNCbwK/MB0CJNWg
eTTTdwWhljT/QW1wV3Crw0QChXA0vFPnncs6alUz+JCGiQlLVFGNoKF6LUMI4fI1qMTJD/O0Aayn
MSeddw5v0sgiudxdF3osU6TChCVhI6zsoKEvSIMOZ7U3eoP142H+YhO+z4xaabv/DjJT1TwVtqXX
xJoRWO2MV7/R3Upu1Xq0XZkzPG+7X4xXvuh8BnHqCra32q3KFEbEEZoeQ8jKBcXZUtibwWjdJX1y
ODykxOcu5+yzbSHvWVhTjuHrBfoV15Zw4gMoCgd8OY/gfgXnUHKSPea/NvPQnxYMzYoDRdvKamQo
HvOWAqf7VWsm8JhuSLFYG0YE4UOd3nI1wxpm+vqiWO7XZIe/rXd61J+ARbUmQxG1QeXaqcvQjQbu
F/aMk36kwoeIjpD+Uploc8XUWJM3YsYkstHZEmN/YLDTt7g8kTJkwNdz9TTgpPt55lcurU7I5Ddn
a8eOBgivPt9MkPGxOdtJztK8yCgvYvRXFd8K/nP+5pRkU2g3jIMffjKSQIb8uv8narTCeFBV6CVC
ykDTKYdw0gXpLOZmXCl9he8p+vlI5nmTwmbdF4Vup0+kVI/J4EQXy86+ijK7ePfLd4GFxHvwAVUQ
dO4r3/x2joBCk4O69JeddJeGF+pboHpzX7DGuvQ9iDsyORBjuXuDyLMyqm12pRC9QS3ZKGnlrsn0
/3h5BWl9OvysRyXKXPiF0LiGwy93WxUdkQMjOjkOLUHqOND+WOHX80SqKl8tPFVxFYLnAEymv0py
7SfrjVAoaUz0VUNIap6GBFkWaHyXAyyPBAOWfibNfk3lzrY2qtiCR8+PJFq4FAPnB3z/4kZBNJdg
TkNegZ9Ntshs1ETHKhT0njN0ppiHKmAr/v4qA1SWQoxVjFEawhcKMx0VZ5zRvufWsBKuZHE3do5U
BJLX5PjnL6dP8RoPGfEc36W/1i2c9RprGgEm4CngQJNU8Hk8YvxrBNgG2hf114fv7tcf7UsWAZ60
gWo6phCGnB4oNNnQI6d4IVldXTHJAL5ltgde0tXb6ryeLFfaRHKaxmFxM2EL+YxBN1C9/crZxe4G
iY9e/TjGiJL/B7q42WUaqzAkGksCywhkIfC5VH98w5DBmeVAWUsMyeCBaVzx0GQiH9L7q3I+8ZGn
brY4vUIAQeks9H442R7QBhYLJkk3zTqcBYw9QGF0mTzcmtenGXy9ErgenD2VSecIhdQUX+yC91oi
c7THqkfHIGyHxFN9o+OPhaioWKziQXLuEiq/WoxFP4I1c1UHZmlpvUJAvZ6fmmevIKsT5K9amgb/
845gOg6477eRP7N8zqYwWOohlxvzaJcoSU5N69fPwFMAh1CyVVQBuaLZFrK/k1o0+de20eXM1ZiM
MSvyH4aLYmX4BARrV0fxluLUqzTYIbghkV8LGATEShWD6U1xHy9HNF/svr75m4k8IZM9LYNWtFaP
e8Zir9XS7Rrz+4vQLkuUKt7D863O+vvwmoBw8s9GedeRCO1jUhik2NEB1dnrbfp41ZwVRJE7s61C
9QXg0LkDpUMyWo0dkMGB28+declNKk4urIMzULeBwyC+L2P7NtzmiCmmbEZ5EHsFAcn38XVvYQg4
H2K1HqI2Yxt4rUdbX/SAyaiBijRKVy7fPdzfpGd2Urk3LRoxxKlBK9IB4gW3I02D4DF/YfCyzNKE
QYkkYAAQjLa2VfyEF4WkbjVormKLSo80gmhJaB9BeVWJ3KzPQfP9nvapXRXTbO8bQGcLhzYHEo+/
mpOYx39r/QwVUbA/+Xhvc80JAump3i9hLelDDW3GEXTew1gZg0sMrEqpFrnhaFhE+Pm1vGgE6sDA
6pL46oyKae/HSfitRD6zcu/UnxDgeT3uWFNjDsWurZx2PkYgj64hWrwkQoUErn8vMtKo7SvLLFCJ
2iBwXYEIh+mzL7P0HbWttdNKIp1ZUH4BogYlOi9o7jOeOeeqG9hcgfN+l0a0lVAG6k9Is8rflms4
dizBMdF2jk4GvH7jLqFSAkigrKhW1RNB6woeQpExwizxhaYD0P1bZl16eNZxqKIsO9ma5ySQV/jN
MN3M2oN9p4ybFg216VrHo0cyjty/BJSrN+DuOye+th5Z9FhSMhbkEqULT06db91a5VByR/7gRKgQ
W4Ff14pO+Uc6gFbkpSkO8N4CyvOpveY2xaWmTrNLhteeQTfobJq7vtWO6v2cRkOzueTpA4Yq7wlT
lzT+Sq8OozS0JCza0c4uC1CKNzDXYkWwU0CDhr1HgmMwAkiNJ1dBAeSTjkU+1MqToxKWRAZflod4
MfNj7WSPDzmI6+wpqkkywg+sM62z1q6gfhLXbLO9GhotcfMwClTEQDyvXVHgjM7Gm7nHMhUv0i1j
cHX9K+jTMKU4kZYcoi2aCiHxsYEkRSM/3SlD0Sq0C8Gd3WXjfbNDC/E+V7yR0ADq7tOdaKgsBm46
SZtuBQtgffkPhV+4nlpA9YRzwgwgt5hl4v6qAMqZraJ42kEOr+x3kbg3YWiGTCiGUVmeSmIsCd//
Hegxib0YwlHLwkekdD7hrU8ouQ58dKPFzMOsHto+kjv+IAG1Cd/507yPMidLMGRLsjeVslrNxYvI
ZUyo4XNv/lglwGixA4HV7F8NindGoznZw5EekgDeSOak/uBOxycHlMq8/9OBLlNYppmRQM5OSRBo
IY51IHv8PRqAEbfmCZZH3ghGFOapRGxCrqbDcUthc6vZTgphsyX/fLcfKaMAUAj/eGT5EL+4BiwP
SuostLGtAWv6WJVdycW4DktIBr22+xlFWMXJ3fVBjmgibmvHcS89fCWqjWGVxjMLmh7UoJJP9K9G
Ak4ze/GPamZP8GtPhqlIrfBGhfMZAsEiwKzqsFKbqrzhpyK6xoyQubU/YVrbE9u5MgYWVZyGOuwE
Y1WWDEMhNsai/UrVsKImbSjwdgBAt6G2WRQb44BxwrtR/0lFp5Y1U8z4F29NJAgi1OAtuP8vCAS/
dOVJvPcC/Gp/Atd7Gcaa91oa0HpHNbTzdngse8C7Fa+9mLNZMkEAR2udPS3woKb4pqEHOcW5hNco
CgWXkCRhpckRA0EOiOGov1hZTj1BenVOnc3wPKGMtnFzF/loQhQQqP4RrGye1YjhKeQUVyI4PG94
qU+2nKpvnTLXeU43IzkAUkjezW9jbexuLZnDoPZQCwzqaF/VG8ZVhzpFGaRRT7/gGaBjmeGEW/GW
lKjBjrpFQ6PFNnD5LpfaWwjPyLJ3V/4mg0vfyNtynOPZKFqaoDDH0kKLa70o/vEZ21ADfzQa3yqi
F1c1nDgiDaWkQhJfuhVH3jAQDuWbv1WsZ4bObUKW4BldFPWn199ftfOv+MyTCx67q/Fpq86OFlu3
5n43iKGdwd0DVekI+7mmS8fpNSVWhER6u9LrnramqjFfObpHZ7tUj5e55f/H/TMvvDwHjw/gQD7f
r991JHFpkPpnsj4vT+Kr6H6vedKL4/qbLxrTM2J0SABkdDdiSEuq5cVXVsrlJR5tBkNmTHb94oqh
nAMj9ZtyJE4B+/HbwclFUbHomUM0DQnHPkv0aKVbsnQX40EAJyZTInW8KMi9c1/mqkqA3SN1TlkQ
P1iGrtf7JizkRPCIRGiv22Zws6DfButJRyufu0sCjkGfvPltqV+jNk5/ZilI63UaPoXNjRsvrsmK
BbvRgZ5YMDWXwF0jvogi56wC+fhagCHG1sYwn4uSupaNxMo4nPINbEhEOd7eIzqNzn04qmJP4G5M
el9Xi6QbZYLjylbES9sfBt5MqFmv8snfHgB0t7AHXIIFjJJcJZOi9wu6LSyt6Xbiznx05OVZBhHy
7ZaMheT1lwz36gToYr6+hQqq4jOoZcRLvHOilndZ5eVeTsJ9/cKLuvUUCz4PqSxEr2af34l+/O1w
nxhiIlJT2sddGXmx4c+vSczBgkGV2ghPyGrONkVjzvrbo7INEL270y69Ubm/vbVjnvR2+oJ8uMIw
EeVngaEUh41NH/U0cPyMqDkW6r7O0gqVU80viaS02NlatrQH0u+gIyilDHHDovo3IlxgoPZnP751
FhxL7GLrBh4qgNE5NPwEo4KAR3ETUCBPveCAkBUkYtDeJjQ8sIDSIkP3fKTbl44+4x0/ofkfZLKp
mZZs1LngJ4iHuBBNofU9ApzblcQlbtpQ6KJIV98A9Q5yasg3s459lBAkB40z/J5Zz43MRr/jKx+C
wmAE/X1ZyrKJotdcuLxosRCD1oxPt5V71G4uTfXo9rMgcwlp9NPYksRu9W8meOl5M+KGaXOSJOf5
T8IIKaFa7HeJ9zUk/Aqhlod4QFy+nlau12nqIxDOqpsCtoNncQ62kOG6+J7MyQE4LM0yvBcDcL6Y
x0CSQSrMzqc9kxHNggNTu7i9hl6HiHzdTidB1ZtY4/Vuz/eetlqTSKhP1MppnX7ryVU4/mDTkL9L
7W8Z3563oere2jDBf9lKApxfssRXr7kJz8SpmPv/r6TT2URH1ZaYz8K9AE4/H2CWzqToUMCesTj4
r+ZNK3FgKPYJWPjuFwTlcyvuUGx3bQwRh5lXRXi5/GiXHGTFC90jKzNSAtYp4DAnS4OsYEXk9nLo
ERO3LYr6+FXK7h6rwXtVjSHSOrImI4rAPhFmFVlXMirJOM7yMCGmj7PryL8cTYlR8DSsZBRxBd25
eJ8sMYlqgt5dAJSveOYX/ADVv0ScdbfjoBnP+Dm126h9Wg0K82C+JzBZI9iUx42wvpYvaaZTcuOi
40xPnO37zQgZ9pMoiQflHb25z3OOZgVv6mC4ESsK+aj9bs9LQQjwHCBel1T4ZfuglS5SYFQLTe2i
2BXpNsYC5NdNS9B1MAb4mewiD3sIvc8ZSu5Uw/Z+3JRb1cleYsnP39n3tdKyocHmrqCHQ7SdjUoC
O2I9HFJlZtoocE+aNi0YP0Jaksj1q7uVDziapcVNwTSmmymSKFwEHk7uzruhTDWW7N6FNhZtWDTr
npdBk3IVdYMOzHL1dcd8lYqoD9Mhwmee2igy0P9SZ4Pkz0qdmqiykyIfA93K/0maeo87lCuVyyar
/hCjuH3wETSxW8QS9wrjaU0asDnqys9dGgq8b7/D6qTBtg87h+LIjnEHXNo/SsjKjTC7KWXaTBue
FFTiqiqVaLhIX4IvLEGiE0Fu6JpGM99N5Jpk6wBt9CchOcS7ZW6h2bunJlE/M550M2NY9OhsgWwO
YH3SeGg2pfK6HrHKRR4JrKQFQZ9D4v3D/BkbrFcCx2yhRLSyO4+wxdp5Hra3zW9g2PxOLgpCDB+H
Fd49hmgScAMqSy7v59ahBHwWr9Sg8QuKqzEZvwCGXw07N/pYiqHUIKviEz+NuHFE4b0cNquC5J5I
JoL4Rfm97xQiGTwt6o+RXW5r9QHZ0vjBvFwZlUAlkNfZg2ZJ4dj5uNL61N23y2UKKjHIMm5L6Iu0
qWfYllmn5rggnT7W0+mVSJXuTjeXWcak4TBft7fG1X5aAGtWQ+aT21EruAzxlfEfWFObrw0Kk2Sa
W2vqIHPfbt8PRuUR0pTJMZzCGVqaT1ka7aJeVuQfkAf18tUQT6kbYY6LhC/vMLLz6i8XeUO2vOxD
V3TjplzWgUxWypv405pHw1uOAJ6Yzwqx4SilKG5EfyVI/V7KgOMrZNuAIrmUEY5giF7rVNQB5b4O
2hpS0YJqeCV/btb1w7Pm38CFVlGUv0Ou/ttth1AMBucJbMthLt6so52t0uGf5MiDquaELpBYhvkX
cT0SGX7smzQPo7xKbwZ7rSQ6c6xKmXFkJ+w6lLUk3JwTezaufxd4k44rTqIFjeV73tRjWUr2QSt9
jsOKfIJaaHDPpQ/es9azPIktAm/rjZPEGeongihVZJKMmMCP4Y8uTzW9Hf8bhnBMuhaMxBlWgZHq
kcQrB8Lpvm5/GkDdjFeazuDXI2R4ORoX+SVfJ6mYGUFgUsBDAvHlPBIq0c1GhOmmhr9luOnhZ/H0
cvMZiiIqxzlsxJLempDUqGD6OZO7AcERpEU6xQ4myxyUgUApzYM+ZLzVPgS3LMaZ1a/4ZjyBH3uj
oRxsyZsBJ78tAL4YrV7kx8ljIQxj+/k59noN/qDFLHKOykqyA+ds1vaedF40d9sbTNQyUYhMCawe
K0IPNPHlizP52aq4Zx9Sg7rT2Fn+0rVbDQKlZ7CH/Q2woViEZ4EZxtUmEl+q2u6dQg79IwM0smYb
IDCxMkhE3/kL4G//j33IOLsT+xd8jx0w5h8gogjdpE3NaXP/eIClhw3BXgCS509Xh3MHMFassgql
mDKyvuFkJJVkUlbgXewcyIt3DUL3KnHtLZvLBCTcA1ikj6amA/ItPCgQdi6az9Zx/XtMNNhIyQJP
5o+0xd7DkOOcrwk7JrJ0t5dL/+/7PDCr1hAV1PWF3hOaS2yLqyX53RUz+Fd3OIi2ZJOOHtHdXYDk
Q5ed/cKLXvAfI1oUWMyqE+5JSMYX08rkMo8RacSCSwvfuupgVlc9mka9MOCdTYW9mh8E+ypcuEsO
Lfc6jgoZzqAIMzGprqBSwBteFWSRHoavpzZXE9hMMb156ovR1ekSlYMztmz6L2AEVoZi/dJUwDCl
Ap9Gm6jj7lPlf3apuAr8nCQPAPMZjqdfghPCq/lZdCGRANX5nDnEWOy8Bb1Lm4xDMzzIN6sUenyT
FKi9YvegCh9JbJRRockjZ4fv2CFdGLAo5i7vwiUztFGAU0VMxZkDs37QmacEEWfRtHjIMZqX+LSM
Nl7RFwDA+HY4X89zoxvpczFVyP+gYsrXfWD7u6uygup4p16z3+tUOm+wSXtOD/6WAE6YZJD4k188
wu7JU8R5FOK+KQZbf5w+aIBU8NTis1HHRj3tyJvVnHxuj70cYYyOUSyzqEn6urO8Jom7lko7Trt6
8nsXgxVii1Dx+Gzk9Rlc3KHMDIWRxCQ9Rv2Er97vy3LHCGu8AoyuC73KDyI28u1N1QBRFJMKwz3A
E3Bnb/G/Pg82rdIkb/v0Xq8pvivaUXbFPxZDwUDQP1mbzCadPbsLTaeawxzBDlznyEAxLxqkdqif
QFTHEb266Q7Vz40o++opbDUaeG8KmNbPZCh1j9cHrcMkMZQ1fmrDrYRounNamKDupTFk4F+LuOYJ
km6NhlroAv9BhE7PDjaaJUa2gT9OaZ6ZI0PrXTXmheKjkubYtr7E5wzYkua5zxXweEj3SqTzXLex
a5N6UcYbQ4Rb2/nrrccnNFvByran+U5lq8mnmIEAZ9RH6KfWGLvRPo5HetXMKsZeJ7fuqBWJqjG6
HoUx6LWOI/QaRMcOGtQ1nLGl56hsdfKXcEeRAZizvMfpT4O2g7eqZyGaojgFSDm7BL5WlJ0yRk0g
XIOaq5JLhoJXGKjF/kahgzb1jonQBo2D9OwfuzDNk15ShhpHQM6M5XR4XewF5AHOl0n+b3iFdKIw
mulgdLpTT95WmPbJZj4yDkh9hovnNS0zSmc8lcl/rxnVHAInhHFJZowO5SdJjV7Q8B4VigP/GyC1
ew5jf02c7sUIWIxgAKoHq9BMOJbQY1qqg9H2uLCk21+1KK25Woz97zSD1BYEiQRkxC9Olh0es+3V
6gqMcu05yQQYi4q24cBBEQOor9jR552VshXEOLlvzl4Cm9mfo+LjPPikBoQgx/w1niXX/9U3nIZE
THZM6I2iz4Ef8Z+ln0JkUruzAP0wpNBMeS57Fo8vJLRj6iZmvbgU4TyghtaUdHYdtyyb1aOmS/F6
sDrBwURbBgW5DSduUIfQ92NBVB6A2R29vSnE5wv6bPbBG8grAInnozB3rpX8VEgx3p3ewmfddg/0
yDINJ77fX7yeeZpyF2JCXHa4CEmiretvAZcbLkfO/sgUA8wCGbQoQp1mn9efh2EdkWUwj4y9sFPD
qWU/l6MVzr6C6r/SSLnCN4pU0hvMIIUsKRc1DFPtBPjlTmDhF1blkESfhqKJ9Rz0BtWoTK/Bg5ls
qKCHWMSG39bvtzkQqeKl2PGc5YVEatVMVvQ2Fn+11FbffHmuez9jkMYUZpt1Bd26re9CrYpBAY5w
fdvhaDYXVof5rbEenKDZFRD/OIE47G7b6cwqQnFHGO9yw5xNzFwRYkN/GrcpFZpB4wzSHDOaxQdT
Y5Uj9CpxZ1BDE7hmMcr7KM0FKfHspYV/srUkVwRtwjr9uEyig0jqvzOcCluYbQZc3rqwTmLjOu5p
eDcCd4rVqRh+Dql8lsiQWIHQPLkOp9n4+SnNSGXocIMYZKVohy9gueB4ThOtlnERBkjBazxiqIkM
fr6gbD30U2z37VdRFVmk3mm9+fJmpBvRIxRt3x+nQfFIBs4t4YqjxhhO0l3ucreYA9lBhPO/Qcls
15+AolhG4REOp7aEPwOD8R8GuCsXuNYUijzqBxarkbyLjQIm3OarkCBVJd84yboQQf2FJfz8wstR
B5CbGXL3MMgurfIo3f3NrEes4vO4rcVdzFjsDhdbknK5YUaMj/lD3yJ0LmcRU59GRFXBjHWWcXCu
Fd1GxQc4EpLWl4aq2uetovZwZ3kb5PC3gIC7TJ5u/fl6MYLvTaQ7Ki7IDdHoSQ0kpry8qGSOuz8j
kKT1h4PGqWwqWFZcqbi5b+h7IT7T/qq/XcF05ehSJeDc+54dG/pSzFcE/J3KVZzssGuCfeuO+Nnz
cvuD8I/cYGGfVo0oR73Oj2xC3zu7HWWCXOR0XV/sbymNP7kC32KMCGgI16sKMwn+MktECdGftyPc
PrwdMSoS5TqI565nn5oTLNl6Hi1DomXc/2J2/pNXlVvwayF/rV4bysiPBbWyks2njDn8Y3DBXeBg
QjvH/6fT7vt0vtDdsZZMy0QT1tQqV/Vbq4l0xZz12EbrSAGMueRh19Ojg9ivX+FnTEZdSRSvcfit
xBkShw5cojfqC6d4B9zUp2oU+wQP6Vfd5Zf/IxjYSQLyBekS5WdudvAnYuOc6P5d68VjGE/KkAkE
el8N1BRNIMoHh+16zUndH0mwwMTmgljUsrbxdsvkb1EY/lopQWLggSPurTpkV79Z2sm4vmuYBcAb
pN65PKwlh2vSLF/hXuAqtSg5XRUUzNbs3CNtob/XtRa0qYtl0KbkSz9fjpVhSW20iW1FeFs4idqX
O4toyxszLJwqdw7GVqNs6PaTJ/h5Dxl+kauTmlAJggqR2wH9bTy+h0+k9xIq8HGHErdY01lIfq7x
VJujnuvR3jaMXfrbj5Up58FM71dDCCyNZUat4Wh6KlwLvKZHbJYfm4A9b29JYb2rQ9mBahOE+Y5v
AqZUqdsTBaFC3UtOp5D/B6bI1Fmo3IpjNveJpNBj8QFPKmmoSsRvp0C8RSHX4oRGOU3UD2yluM6E
frfedvYADusvrOrMR07GUjfelZftGnJLEoc9hBBuEDG79SYZO9L0Rr6bfOPuiPJNAdJPmiyuh33J
GJGfUhg0nRrzpanFYmLJp5kxesNMyHzoYKe860Dz81RbFpwkditqud4D2QfKzxJ3lR4tqON5IqCf
1jIZ0kpn4ajB+aq0xvL72iOU0h592vYl63nYkROTzlc8OPVIiXJqgpBXb7t7CxfrC6NNyMNdCe4U
VRINhbGjM7YlpcukKBfeKZZOHzHX00NeVs61nD5zUYC9VVEO2CgoIfOXMMtVc+mM0yi02e9BQNOz
pLLoufdy4Zb4gjuncnfjZrmIsNUSuk0dp7NE/YfbyheUCVse4yMQoQMeun05dLb9JIY0xTIV+rFG
GAYNfH+0y3Nw/nHLe6j3kN9xC3dwoM8Yvp2dQ5Hw23nzFNtcuInZvJX9v+aSmG1K+mtvR1tH79mI
2dkwxS5nIJQBqTDbrRHRqwghtDu2liKit6apcs/SA2OcUdghoR3Qr6ySJfPEsb4Hfwjde3nH7S61
IoHjGCQQ/MKYObf7TxV0gBATQuw+/vBkY9wrz8vhQz1QyIqV/y61tOf2mZC36rwMfgoBe0ri13sf
t+m+bS+zLKg1kCiscBPfqFYiESDVU2JZo8iXB0/2zZ2YsRlkQAUYBqPvXbOR9HtuJN02kp8uysvn
LDqvb6YtF7Fg9u/U3ZsW3r4Y0cetv5QLk/XBy2rpaueGeygmxEeZU4Vo5OYrMLjyj6BIjhnYZp0d
Qy8OfVMOb6ZPeC1w+w3/lHs9sdNiksXNbDmcR/rZl7VTTN5lkgTWJlfsJ5XjPksnNJe1yzc5Z+GP
l0btQZu7gg/bLi3XbKAT1McgNWP0an2qj13VCSVD7unO6XmeWNkWZRy0klzziBkEN3M+Mdkm2q88
s+2GCp0TffSVIbQNxbd5AK/CV2wfC/7GLzI8hKqzPjmuLMIv9dtzJL09/Kpbnn2x+ZkgjJqcPIet
Tijyn9MjgJN0DrSl3lPonltapiXnqpcCbOApY4u1UTnlRkd0Rqkh3qU8b3KIlqfjiLgGGJDwW8/p
trewL+Cc9WCL6aZvFbcOpE0j87mYmUW7mGQqJ78NFtNULQzWOMUAzLzm/9JlZhTzWAVK81+PoCz2
2saF1s+2EXXCXw1hOQtdWmJ9mql5czJSlsMLZ0drsMGtPD1Qm4fFEb0WzaU28hNuFc5Jhz/1UM6T
t2G6ppIfp0Clw7E03dkAhMA++Lj5KBLm4J4OkuVvx7FsovNHpyarYZ7ZxpkCX39BhR7e3sKGRbwr
Yqm3/Lx93uJWrguu94AmfBv4DOyIX5Jkt2Co7rxIMYIx5ZRSVe7qk9hNDeWGSRJVPJZV/zYg9NGq
OAAOKYve5HbjSz6wrNASyr7gxTW9SLNb955yN24iLvfM4+0Oguh8ToPjEFF24QoNliO8laJKNmyg
3dwDLPImcEkbCy/iNKe/wf8YdGufOxBf7fus8wVLJL3Da41Qb1MMksVZINSCTYHiVxesPt5YP2ii
o5/tVPy3aO03cfUACkshZfs5+ImcWGsENE/xJujWlfVogXgKzNOSBcq+tI2YUdqShYgUsbPTAjLV
psS0Zf6jZxuupKEDJi2HUc2iP1CdmbKg6GRJPc2ztU3ef1tx8tXjf8tzSbQUDzNPNbSu8a8UItRw
xfcXlIc5WDP8BY3Gf3sShtTpoFTtShLFfgQN47yPX/dvu2ZBWQZC2qNIk+3Darna0lpT7dFoN2uR
MoCQ5C60Kvf/+17y49/uDiVcTylDHlz98WXi4qMDYWix+gXCYBEr41KtST0Qj1xGH3hheI6XDzEd
jbCK2jF+eKXO+sGpWpT6EeGPAFuyDnYbiYEqXmNH20zrA5FAGhxe+ESSkUhUFM7Hj2MzOkT1mqe9
pW1x7RkhZUy/wjUy43rIlQicf0SBhhSV0Tx46DAhbJY/7OAz2IukdG8XvwuWb3QmsMOoL8AR0kTk
olKtemDwZkyjWS8Oy/ra3rEfLMvh92Q7L5PmPQOzQqTw/WpjkV28Bdd+1qyIrm76c/F5dD9wzyLj
3AoTbCOa+xVYj9xjwE56CSFxtCOatc+7Q1Q8YuaQf4D8qQDFQ1eP6WWIahqpYvfr8BlwVhh5xNqD
OUGG0TLFv9YXl6R8J0H/1X4AOkgr/4orZPRTwwI7sZLGXO7wBLdEr/8FP4aFcCJ6h0hOYdzutdlL
n30UvuJA0eXFNq+E8gE8UxLFY7OYJs7bGTG4Al7a0PMcrIe+FZOVDQJKJkoHiQRhXA3WXBjLhtVB
vYzfZ/sUm4K74wLTQhXBy5c/eZoJWSf57Zf9bRoVPsFFOEtxt2FhzKs65dVHGG8Gll/HiUBQS2Hj
4I8mYw86hYvFoXWZdUULVKAElU7VfX2e4roctcI6KpkLSeNZgoLrGLLBqTrE9cqELpQOJwMRb3uC
hxFmBNzl9FF4qg8J/y3Zx+aoE/5dE0fNhinY9Tio2MS5a6sjmeoFxKvGkk6k3qIdQLAsJZaP5svx
iYLGQ5doxm4VHEEqZd0+jcLvYwbfChNeWZb2vRCmNrtUqfSQqXlvgg57+SVkjYI9vJn0OFGXPChm
iHF7lqe+Xo93WCfFxl+49m3MEA4SDVDMAyKh4OCIYZxTZCoua7b49Dx2sYaAtgkFbfvKz9t34iYg
eKkGfqAf3QA2BZ2dGzzs5hGJnfKZa/+fZv37YZZczNxJfewLQz8aBuhRmjLO5ToWI5mbtmcydQQk
bkPPQVivcNhUl3NDEuWCOfjU4qNyaybp+1n+jNaVzE2xfQipr+ZQgLZxl+mpPF2h9r2TsGpIrngw
Q4sgMsKfXmCtO+bo3GKsbEtEPRXdxOzH76oSGoL0u8pPdIkBG4ih2fBO0vDvGAqsHwsAKBvIc2aT
oghYdMIuESwz08ewuWYD01lQ/celv/Wfjpyb2J8y+MCooHMfLbXfklb0tAeIhy2R/OosQbevNbCA
IfNICDktO2JPARJnSImndZtFjSjNk8wvEkK8dMlY4HsxL+AHtJvoY/wZHTbBAGjaupqjtRJRSDBv
M4nTLPpdBQAaibacpm1cOFnQwMXRwzrMS10SlIOc0EU3iz58eBNjcMohxsf9FxFq5vCdEkKgUeeS
+ft2BiV2RdxOSOmg1jKLHg5AdrjWQj5Xsn7B3galLV3zahQXfc0ocJVhNYeLAxqJi1AOFDqXz5W4
5zwhwO6xbhQ1BmZAwe4VoWMXFQDkku/tJK3LnrbcuwhXyQfERFomsBsPQBiF8l7FFghwj+CHbbsc
B6EwmKxA4x1I9qe/BBPh7MP9KHpZkR5RBY3ASSeJ+XNbBu5p5b+mSHPh5m4ghzw/e5AReH8Pp9Ih
ZXRE9ayN10CZkgyMX2L9tn5FAu+sQS+47Dj3U33JO4SeEsQq6yv9EZE1PTXPaVIQWhUULdQirC77
hORR9wgjfq0t89KdwlqErxA/alyi4WAhDU2bzBVlufbNQQF192TxN+USIgiyQ8mhjCnVC07Onm8H
F3wyQ0bivkYEvKG0akxEXtwSFj90NDYmhMZX040M4z9f2TotqDP9G0e43U9lCVmaH0Dj3DldwXY+
9JASahGsx2qfuL2JFAA5nw+qTWZrSXa/8YL8xM/9uiiFL2c24MaTPbABDPyEm5vTahkpXbPveVzA
6j6Su+fG1G564G+HVjZ4XQj8ok0VizAgfsikW2tJWJanWmFx68kQTZVVPELiW3o0XPHhLcxagnjq
ZHHf7KUYqZwbomx2/Tv0zwzndn+90C//zf1Ct+ifausdA0kxwti8Vj9acWRLk6y+J/rPpGXAvm/e
obmPSIaFnvvYfszpMC+oB5fArUWHDIltga0yiGPBLkIDtTS0YsZd9zHXc1/XFpcldT6NM4Gu3+eM
QvyTpBcLmTEMk/FVVnm55iJ8W4ICE+37SPyircKmVzT37Yai0Qm8VmmCSIHehwDlAxdU0rptUj6g
oPw6i5Qb/WFV+UdyfcwDs2lYEO4McS0YHsHwNlzttvkt7uGHh0eW6Vu6EKaQO7KF0MoeaaiWlwOS
Wy+lnK3tJXvrsa1XUk/z51jSY0QtnB/1oRZEgzFRRr1H3j7NvuCXuyKjuJg/GjWWjNFKtCygJsqR
kcADgn+SfZq1HAuqgaS+8yhBvZvWVlD60ZoHd7bxAux8yJhs+8/fpYnI5QL1jIisHUOx0nsN474o
tAu1nMnIDFUtkfMq+xpqXMwCoS/6vrHqZ44YmIDG28O2co19am9NizaL7Hd3yzUW3O6EyweKtPXj
M69T6saSNkfa4EzkBc25nmohl4JfTmOFxSQ/FwFwcFUxwvsg5lo3q1jme4xIrvax8I1u23RSGnoW
3Y6OWgnD3zW1Jq55Y3YnmGBlXHACt9xjQ+kZb3gkUrbrtaZq4IT94++xwYF380pzPdqQzZl/I3WL
s8gQjItboI8gGc93H9Z+9y1tYaE8g4JwPV6wPWdeP6oVeWRYTv/spCqnWZ2WupsI5tUU0s3Vb9wv
nHy7j5GHbNZ1Tvk1A0OiSm/jAFAWD7IHd/NoAjsDcwWYvbg4P2Gz3r2WlygIEJLV2ruwz178G0N6
MoSuk/d5OOCWoF5m++gxtSnfb/eFzMB0Ft6mpE+6NjhbCbFX9AvxpWhuYlRpJcjYxJxemhTMRm1y
RkKLZkEIMZ89A1dV0Jv6wQlteYlrINPsWkZRnV64KptLa1i8EO9Q04ywG/0g2R75unZH7P8gBPyc
rjmyHF9fQbXf9YUTUMjQYJjFX1Atfv9chDz5m+aLidzorX/LWc8K3NyLUiRRL5l5KZwihxKfnBqE
NzKyRPtAnR1JLpecwJ1kZiMr11GIJOoBaRvw3TNZT7Ep5FCAzrx8LFpJ6e1ZQ1NEGvCSotHmjr0J
vArXwxi4Q6GPwfifiw9cMU7kfeodvPZQEdUcROQ5FWv6pYkjAaQBBX9h5uXSVhRgWKu5ZUu4Mq44
p9QrF8M3RlrK+xRznUlB3prMJrWyj5REcspCX5zr5cFOPmfh7gvEgDb1fhPw3UjymH2uPE284lPM
bPfF1PK+pAajsAwHDjQQ8PwdbY4rFVnzjOmIiFKkz9KMPprGtoPyswq0pPMWybW5vH0h2/qPH/bN
zz2bDuiYMQEgJK05zjO1uLzQ/OjDqZLdGoBOrnCGm+lAKAFxRM/njRu6qaa7DAGRHbMc/C5lC5r6
HATg+0VGvhVY3kCRxZNQy4psA7wHc7z1WVn176K8MceQXgKvj/FVMhKwTypIkQkJmfbRZc3sgvbY
hre1w6l3WY9XIaamaSl/PQgH0PgymqE4V+V1Ib1EdhmVdAw1SEomWZ3X1qH5S21z/ic6UkuDtv80
5F+RIKWLjqvws46jHVvRTetU8pDF9OgOM9CSJsSN71YXpRfQonpA1Wnx2tTunnQF1iKqhYVZdKTf
9HYXZ/+fgFxC5cSjKnrZu81+d6XNwWTUC6fvW4OptZNRb0TW7xxTrYvePfxuXl32ZEqQECeHOQ84
KYOS3wY4LO97k7MRtiLS6LxF5taSSRKi0gtLVZF6sTnrqz70pBe/J94nuRR2ak68Pappruo92Zta
IFdf233uwf8y7OkTkyNmi5xTf+RXlqoavReh6lY5+FXMXS7YEIuRde4gR4IhPQeFJNmQcPLkVHqN
V7xLCqVdY7izgIVpfbym1HA/+y3tgJ3badNnreEVYTEGzHgI0x7k1Bu5DJkFt1D7E7YQUPOS6YsA
sOI5K6MeVePe1aXR4H05+EB7TN7cHNEWbw8e4dWJulAAViMTcqRc4G0ezHiVzwW0ctn0078zax0c
mmh7eBYI3eUZ7Siq84zR9gPBBeYDYkQS89GdTQIoUlba06Mjv60BkHMgKoUfdTeBgyRILAFaGf1m
dgf2H9HRfJyVAB4/dK99ejlL8+Egzq7U3vfURus4NdZ6Ky8CzRhcAOZGr30nHMCNGSTIa2+Ho/X6
4jAKdoryzQO2iQuAiIjmWxXii1vdKr1jJzM6lrn8coimGWcjM3eA4lLK7kYOZ4kKZnsBnqYN0XPo
ukrSuLJNogOazskyqvgtfNvR5v1tSM0DmILoF/BteYZk3vf2Om/1t1+hj2DlOu3yEZNt+aCIMlDU
RLPqR/mSbMsLQdtxtEazX4EUBFSqGXIO3KjQ5GnfdZQdll5BHD0uiQKe2D1XnN7NCzlQReVYW7jF
HdkUDGbTh0YlPLsNtvIaFd8xAM3FwXNRhtI4sAqySuP0Gf8+lMQGWPKmC8WUwJf6IDdXUCgLlU9z
MftDAgqgEqzzlk7lT60L3aYll5W8DQzYayqR1QJ+sHJqC400wPH2a3BLocFbIKxK7J4Hroy5FmfX
R+QqLhXSBfcM63k/T2BTylf4mE30HXhilp1u8b/vg72srlkJ6+S0/mUBfl6VVbsZp+ErgCgpMkVO
9dp+Bi0nh1zEIBohMMZ2PcZBdkrp+u3T3mKhbjJUSGoI9Xgoe+2jvMaxtp+CzVLF8/TTQFluQYvZ
yFqsTGf59MAu2m1nHd3kZAQyt0eXopreRvqcDIaTqpt/UUFH1boUcVoohQ8mRlgzTBDvCoTCH1Mk
pDW9n/S4NRF97SZqE8Gj6W8ZGx+O/IjxzATwWsHgNIuQXEHpapIDiGBcF4HxIpfGuiEG5QmroT1s
ux/BI87LfAd0/9y74F/3Ia0cToo071w/WwIuvu5D4/DH5nhvKX6tisu6RPUplQwMg47Hc0ts8Zj4
en5LrxeH5fs3uNTZ5ewvsANm4sYKB71+J2CClMpkKI2j5+DLYdbpr2t7mtJwDPprTJGGJdXA825z
hNCN3txYrdr/b0pTG+WCHyaraQXDMc6QhEThOFkbTgHfJdJwCwRnJzG6f1rvmdNEhH+GbMxeQAh3
eOlFDiuwrd7fV93QpMB8LDJy6P5lZ6WidPU9iRC0WtWRfGEHbYvx5jTrJ5leqG1vs1JpvsRiSJce
PSOgY9NK2d19HqsxYG2Ht4SxcUakRV+NjjeCM1nhstklSWWz7QKBdCLxxXqfexBBGNBGb3DnwHAW
RRBkNCdWapv9VOfwRors3JjqkibemrmPavl0w5JgW8oTP2dHW1uB1rAYsAZyP2iHi0IMDHVVfpwS
bdXjER71feKO3C2MNxOsmN6wMXvuBXKPsvfMDdZJ29J702G4lQ7U3eApMCtWNY2L565bqkXVPqgx
WvOZaGztshj/cXdMDb6//m8o60TDsHyp/bRPSaZsA77+9rECxBDN7IbxOM7QrP3XOhgbQNAW2bEy
OWzpR+7+hVsr3hHewxI71NjE3XbKsBSC5HjqMqUy1y6mjc9VZ/CR6pcYffGRaUez+StksAl/d1+k
fhXH4G2yh5ASvjrImYn5UX8EZFnmK0W5LVCf9IlFJjTV6EAGet8LgcRwDLkJRfpCY8KGawneo8om
RP931ZmRIqIlU3nDYDSgfZ988cumTc10/K/cmDr+4RrEvL9Zpb3I/UI90C+pmdV8WRXtz6SpdMAE
hm9mKf7VhSQaFWseE5ACaQF2lFqIBKQuf1YzYhjZz/0TL3n1kuEompNd3wPlK6jJHJPN4AgiJn+l
Za0Jz1FAbKEm+lZAv3AcgHHoeODyyBi3n9Znrtawulk/tqTBoYy64j7//ccBvmmYoqWBa/lHOkio
j7pdCSA1opXsZ9h/Tbk3CLI9f5N7RpBDpa9yam15aM8D+j2TlNdA8tq0bPYvuSd8x9eagLgGWqp1
Eg0+jBS9Ku62vrZnyZNz0GQE2Iecqy6a52+wlnGXQ3jwPv6JLMquxQ74xw5z2q7GUGUnGL9Kwju9
DMQL0aE6BdDacXhQN02KAV2jqS5m63iky4FmkGw6tPPXMkHPdAR6TwnSIw9xOPUauyXJK0BjviXg
k5qnOCrgmeP4xak8ZNX1cq4o1yMgLO+ebJPInMbtlWEYH73zU+dLBIX1X6tWqwHdQpNghPoOphwf
bYzinl5LKzLTs61GBvYQbsmSAB7NQ0FZvB/iDq1oCQtrKQK/jRKIXmuv2axxSVs+XjsCHE0znSv6
ThKebn/JUqq45UO1TA2Po99LTt6soSvyhV3Se6qxOVBB1ceq1+sX+Fxyma3YjAhZrtVHXWy1HiWk
Tx/S0bkvEhGJYVMdSkLNQBxvbRi4TDte02Qg6ZR+Ozzz76rvxsVE62KkZrp4/afxYPLqOZd07lzE
jBbg1Lxk4lKhWjR3I0Ipz5L1Az4FmUB/N+zGok0ZPqJ7d63GHw4UZIfiSXm2iKYeFx8g5yxgn0T1
asJsCQzn6lBN3nMpnRwqC6Q3zxBHgMmL5slr+Rv9fEzJUum/hQ17q5ay0CM4NyrdVj7N6gngfEKO
3LlyUXZ10ZrgdItR0VDfwNTJElkn+ADF/2f894afI9OOBwEK4lZgf7M6OsUDI1VqaPuENJXYKwHj
g8d3nWhFxhpJ4cv9USG5U8TgBDmOX1JoP3od3V1yQDYzRRoLSv/eKuBeI3gDQzleIxNqu0nE8QVQ
+sGTgYiKMUW+X9WNqYg2HxUu5Bd0iZNX4OWgIua80YDWXeX0xX9c57L0TeMpXx9ksXfRaw8U92a0
PMY0k3IluKbUOp4FmYcuyf3dQ3YZh26fwBlFtr9Ifk7SdJEC0XlztgfPuK4Z7GAssjlpi+ynZDPj
cP/duI7ezNF7VtKEATiaIO4QcM6CLXL8Ke7H7Eu1RYOFy9ottRcC69x3hvj951r6mN7Lka2N200z
hpRqSQtl7/Q6tnF5sT+w7nWZ5iAT8BSR0EhEgXv4qQs2InBHPuJK47Nsx0QyWdL8QWQer2kka7EW
zLmHezgv2SXaCOH/CNVFQvgZQGbrGWWAAnjjZSdblqhrZFbAW/uTkP9hinBI0pFHTdTQdRSCBT3b
jwRVdgOBWOV0JRw4p1wtyByo+gQ4NqqF84IZJMWFxe/2n4UoJKCiCK+xjpHHza5CKg+tiNIkBUNd
zFKTRa4aYG0sJsDZSvBr5zzsTVoI81YFSiTV4uPzGoUOHWjGX7LFnYDlAMcWI/uahZ14UWwn9J96
EPl3RqB5fOt5HjzPQHW2YUu5adSgw6NHR4B2Cp7MZ4zHx5ixokz4SZ80M2yYZwm4ue39bC6Qxqr1
ACoVcjwdB5EHxNJaLVwy1U/oLWZSt4yhdl330ybQMXx4lklFy+A9J/iMvlbXRhvN2AYc9qaNpLNo
CwGL0/qXP/RMPv0U2rNwD10sWsmjyDxvxxTbREE36p6oZ5Cl9DaepCuzEQM+uAwW/afCWEx70Q1K
U+wmHYN9SEKCnOqd/L+WD/DLMbwBMDf44h4Epu3xB3ZsfxVmAIBLdKY9DSa9mTgPmDQ/nNK8JdYG
/jH+7XtRQ+Tsg4OV1WWDree+l8BnxcAinleDJMhlf2N0uyRzk/6cAriH/P3KI7QyJJy6gMx9iibu
aKBblPE3M3/dHICYIFRfAiQxydD2TJH4l7MTFkmREj6RnTM9rl/9whxn40DIwBhtdFRjRsTZFF/Y
lKZOLgdsGf2WOFT78muk4OmQKYyZQPPgXYsLkzBtFaSNQ43RM4gE5siwvJ58fsygMkzpV297roRT
Cizu8QPV939Cl7hJ8ivj+2Kb4c2mFtyfUu3AexyU3wOLYWlOpAIufzxqUJ0WgIx69FDlY247csre
6L2M69Qsp08NBj5CiCnly0DyKQau4myN8T7Zq4xIa2JRCNa+JvVMDJHeEClhfkLKCauHEVby+ENs
up+4DMMOP4uDyFto2vTP+PSfxg/OZvpJAfR2yxO1kHWlUV1Rh2b3r57Sgt6dKTH1qGDtDFAdGtVp
YgVHheOBHD8Cm0/ao2fzv1RSoNGUVftTL5OF4xIk+nwENxbodnBYPgjTKVIPFfsFKq9xAiEfd0yY
jV3e5gikXhGEWZ6xBa8wtM8R++cXAXC/sOiP0L69qDcQTgt4kbOVdKS/1EEs0ItS8pdX2CHnUV2I
PBwNvbEIvXjfURN4WwvUq5sCXU2RupDrvECcR5echSfaMivdBwVpZqea9NtQoGQA8+Auf27wGw+f
eyy/KjN7z0Mgy96VAorse52iVv6/WqQzPeGaVpE9ybFwkWGkzruofFEKbBm6Yk2X65VmUXxoIhhU
8lmL0ZU47D1gznxaintCQK/p+Fb9puMtH/EsiSpiFaCz395zlBu2yOrMPOltM+C/ykIj/cPaFQ+d
HT/aTf7nHjSnr7bYyv8y8RWrhXmzQomqFtaP5GGZCLIiVXZeDj2y7fwvLJxQeaA/c7Cx3cxUFv6g
Ij2wQlzx3J1h7mD+a6NEQJVYY6h6PaH+S1hXQMHWTc/EpnPrQF4jvAkFagg/HjYc6IUnBqkheMIP
ydiP5WGaCAcD0JMU4Su5s67hjOUJWjlz4ZUV4S2l7QdcJ/V7IeMfraAMhshDJmX0Nm8f8VLJGmhD
hUSCa8I94o1rx0wxh4y0kRbF4/77D6natC2mBnnaDMLVKOpNMkrLVSfXN2l+J3veGC+Zqrv3Vm+R
UFfQ49l/hrvLAQF4JQ78mGDe9hDxUcs2yw+0+Y6KXcyqeL9WaPUSoloQcfWTgT3VyBC1nYOO6+E9
VCT1wWcrxHmBpZ76auFHv3IWuoBhegZrF0rp4vJZZ5208PM9kdrfCjnOEablp88xDTZtHHzMv88h
wUewulU+PbyY27OtB0Hn8KaNp0fbXdqrFn+DbT75Z2fdSQYs5j2YUTFWPZNc0w0XzP+RuJlGcy3Q
d2VQzWGwzQprLbSgDbGMkwrnBVWxpH8Anz8gIk12n/hsuZO9LnwCvPHmDxCFKCKjNSQgR6+wt4p6
Z9WMkxrafyvme4gjq/JSthV3Wcvh2MvqPtnt4MA1V/WsJZcmRQ45D67Frd5D1ZylllI5XQ3DM1tG
JYMTmvMPPL53FjdYgwirwNgV+zheMBbGcb8SV8BDhu4j581Y5NseJV2ajjzrsQEDRZEVbrffTAS4
SpR60VZ2PRatc4CIFDQBOFUIAdpJg3yydfq4m727qzGFkploNvE+uuTMeAEfHpOcvtsaeq2wxu8S
Cf4sOXalzXi6rMKwfsGA/G1h52LXTZxaPwTG/O0BCh1gy6GMYi8Lh3YkHqihiZh2oEAHqxGrTMh4
jKXzO3eKAFAn3vbX8V9PZJvXM41w2l2SOcr6b3c16hHZd6OwtBw8ux8eWdSYJACzyRqFP+j5EaCh
oJHwlsLch5oRsyZd3qA5cOryvfspLv4RY3dwUdWPsiolm4c5oKs0hEKMKBzpxVJEhAbYARYCOLne
HgdguCiCw9NiPWZbKNiYpdN04h/9TRqntp4lBnvXLqu4Vci5mCWHfPcDUXO9GkpZgVhn8ZPQKxxC
huiWw6+7vlp5irzDqHkkIZkl417q8vuFCP+cQqpbRw0Ylj5TeBULo9yA+T4Bh/MLzO5ivgKABkVU
Td56q7o4xkR/S8Gg674KXY152pfPnjK/sjDFhPWvLbexWGFi3sQOW27lsQUQKoeJ+MNpAUDyzSdw
X69NMYI4iNrl/IpEN1Ctsw7igCOpvKjXPnkI+CBslsdAINZUkSxXxNbLcIzHhtQRiqMhcH0P7/bO
5cgClL4twz/7L33d/YZChyem86kOA19Kj5pyZm/6J4LS+5TfJU5eKCZwJTM7D1UZMjLEkS7ZIL38
ar2GD7O0KcEM7tyBn4b1O5LbA6KLsn5AAPM5ReRTXndHX4XQxC02f0RIegzsuBIrUId8d5hZ20BV
dOJt5XCB2umx2KatejnznJsm5O7taYa/1IY50uViH1O8ZewZoIkhXnzlRAN2XqEhhAlM91v1k78z
7B76e4OqmZGpAcqdqpu7+juPe1p/kqzJq28bZKKLp3m1OVAnf/CK962AuaxOMTr21SgeZtHtQBFH
rC0TjpMLv8BpjURvbgWBJ6+MNu7dVTtPBFTSteAfMqpKEPMzLd11LYraSNHOofPrCJCoKMi+7EyE
bkhPMubiaCURQ81NFLMfOyodS++HnkdIU4JZh0bdG6FiDs3Xs0mZWS97qx/+kEK7wZeHDf89Cb2K
EjtoxPRwC97v8jJMqclroxWPekxH4BVND2n/VntsNBD36hxohdnXxffZsMiAQ33QCNxRVkuLe7US
RIul2OzRV9xmuABLrB+TvVEUXY4SN50xRZcRSI6GEOQx24guCVSezkdhuE5Sxo5D1E2WsIKYXMNm
/pz46bYFvdf6W2DnJp3+mw8H1nocvVT+qd2UeBZjOV3qBXU8iOXnkzjME3iW3agtZKOMFawQ8gsd
4VjZVixA49rYZqur4rphstP1LILjMLqFr0ecGtIRaT7bHiYtmXQFNzevqPtuNn+P90o3cHhei7sA
gdwez7IcPIagG+/k+MVPoJcsmOm8X7Lteu5b0/1z+YMAg4t1LoTLSJe7ZvoN7A1dwYfmNq4zGUBG
ZTt0Z0yjVNwdMAcc5WcsVSBzaHiKbUMeLdAjvT5XNrrjoQkNXskdqb5DSZiErLBe83hN1cNDPvm2
LBPmUOyUyJfj5CPMTAOT9gGBH2bg+4sBonPOAjQs6NXJjCflzPHD9vaVIGKeDwa1/980Vu6IkKDJ
84dqMcMyyA4lmlPwJLfalUxUweFb4oXzBndO2jD13nYBPYL10Z/tHu/HHfKBiRFa1nNUOqgp80UD
r2XiHcr7W0KUKtTl9KXi7aUO+aTJ51LbCjlcuxUI2EZjGwuxYd08gWO/Wx/1aVW33YWy9rT2xyPQ
yERkvLmW8iOnkP7QY3MCUDY/n2RmsmWSpDczOZIpim1CJt06H2SMccHLFzc4kuuXLQe91/fMUjG1
fd2ptjvFMdIgNgIVn3V0JjCbjir0FKhOmjnpsk9Nhb3QDjjJ/rcstvhB1uevlMxqB4T0oUzOkLGY
xIoUQxeDqmR4cA7NuLzbWpPMpn+3rMrNDwV39oxd/LYpbb1ItapA/6umUf3FgTTBkp4MRctoCs0v
HFVnvb5ffeVXDXJiyy1EdurH9Im3E9cc4q0+XENhWvjCtrk+3j0p2+4HTlBfmEFKOK74aYNbsztH
sA+zgmP10Nt1frvIqQsZOFLZ4D+uFbJ+WOllx42b7S8YiSs5xgBwwBYeBqqPBGjNE7+uhrLUo1Uy
b4fhvYh6rVMBUVE/EvPiztQmOPhkyU3/0vHCrbX/NLfAU1DWR3q9zDRD2ryFvKRTDdpvPZpiscHZ
2wkj+dBrL8Vdnr+9HR4XrrDczHtO/rUSrN/mWW2CG6oUkk0V3k3eTsCAZnM9Hy2Sxxo3jZDTaGCi
qdXLiT49R6E9HI+Z15hH2Knch6M/ROaB4z8IkhnFIsk4Zk0HU7mL2ZXds3GDvdrBrpBGSLP0lES3
BVSZEbyzOysWGFks2A02zWx4fXcevKyzGolbN4kiqHKqboUL4chx3jpVht9fzj2nAwNoe7AI0Qv0
xP0GRMzzrfJTERmze0kgGCQO/eX4Ub/2o2FdGsWNk8oOpDOsSjZ6I3kAZNlR+BViFC6ReWoSxH8X
JJBkhU1MMFCukTzL7Vu7O2EXhinDofR+fOll9Fcz8zzHDvMNQsw1/bkE9goC7unTCbXHbX2hcWx8
FNOp3wjsyXCnIZ8yFN/pHlWoiB9wfW2NXYgQPdhdulOUSJ2yULaArXtBfoBLu3P3IwJ3jBNEKtuu
QVR79c9oj6k9cJ2E6BUOyGnikHRjP6P/fijiQux6hDch/KAxZrI/byRmGfbFdc3HFFmst2UDw9PD
K/Q8Qiz8JaC8N2YaLBBaHvXj8kVuz+p7r170weOdyoEUshiIznNS/FdYbaRMwvNQTF/VdBxRSOv4
JAjt5FEWpDT5JGPq8B+C7onshCeR15ZjlsOT65ImLV4qilmkVAJevZ/aH30PYEdA2yoIhoA1GwT8
Qd99q6CE238/7Ar3Cv1WdDKJEX1mKQa7kxEHXWbOpn4bhIs4YQtc6hAMuocZo54XVMribGPs2sfz
k4q72zAVlMQvKJOZd/7z6/JzxgFbhjtl/OTrESaZpUQ1PNTGaaq6F6HoKog0kG1PfZhpoKiuB8V+
96jHlRVdL52Gy9ReB21L0qYbXMlYrzxuu+Z7zeVkUsCkllNum2Gj15RJiKioGXHcIWvooD+WpT0r
trWVe0IOg1vjrJ+SZwPlJUVu9wI+eLiYVMONgqDf/Ho2FOBJTUsFGnQd80nMkQ1S8Ehftv9dHM4e
4MzlxqthKZQbxCGFRCqVWcfVMgIDraXUBvoA8cyIOSrN1UjSHKeJS0eYsdt0sh5rT2ynXZnxz5Nx
J4aCSOmKIsg6XzqaLeCaP8PJUjbsArh0nrRpWDcdFZVDukYhOBc85jHV8Zlk/toTxSPgA2QhG3QN
Vy1qL22RU+7Pox0aEqttdk92pRvhJAR+46OZTaskaToHatTCd0bCBt/Qq5VLRZgWf+y3HZXy0EFG
+0EYWlBpp8uXTUhV0/ef4XsQJ4JprCuea2xcpr3ebCMx2CJUeYtNZiK9d4WvDXwwl2Gp0okSIrGP
WTm3WOs2dffl+0J/Qi8dw54G+N+5cMOipLNr9SXVDus2F2XJM/R5LS7ue5FV+GwNL1irUPz8gX8Y
xjOZwC39VnwJnyS3/yUHMlBFmW5CdTXsNTtMw33xEB/9BdTDx2dyMzQyf7RVIGo+i10ktlZbb40A
LIhZUsjurP1cwvL0wGZ6OpY1A9bE24FlT0BHEDTR5pQYFJeVpjAY2WGQ3qqrmgl1MAyZwCEn7JIZ
dMwx/yK4sz6YOsTxT572cpt8Zzy3ZHmk3cM/jedD5Jl5bLBIw1opmG4e3bdBz19mSqM9dPoTYyVL
GeTwm9BLn9rKvHzGhLyStFV5tGJGCHjj/LgIxnh4HDz2yQHsfFkETQyHphDMv4Gr2QAUtfhSdT5/
2QiU2oalq08/It2ImMVIGGKvfPIelFxH291V87iHjX+/yWp6v1MnvRk5gGygGAA/SL8TYZf703Wi
zzwdnC8b6ujkIL7TvHf6Gx0Cp7dvHpL27fkaQOo/2hj4y7DmPH44OEiB3xW9E5PUUI0HtUlHL7iZ
dH3R70HpB2wLdqG48DgAq2sUF5wiDYqIaawUz4rGJJMH1koLnbo8LzpoHQ7VvQjw9rh07heQcbIw
uNIa498GwmVpDjnVSLMyo5fWZtytZfasnGATS6Y7vQ47rsgnI/yb3j3H56/Gnw0nmiOa1Q0i0MLW
kU3IKMeaFTtGBcbqJk/axBTT7tp4SG5P7fY6CWNOIHG7kjMHhgtbUfKy0HQAdm78+fnN8CKIYGXB
8tAYqlMhcYnzMVkwJjjppR/DsnAc5AgQoL/HWT67A4y/xeQbxNdMkPsEudoIUGDO/obmuPE6rrV7
Wz3IGbq8m8r5J8Pmqjk6nVrvf9V9PmoTiv9GeHlvRcWt4r/LE/cOjFLhm52y0I6NX51A+v4eGa7M
cpaBUNBnKjGfipEz5mvvdmpuJ6H7EPRsOaZYibZ6aBuvEOLRPcA3y7oGaTaIOrmzKfVXN0/kovHA
dl7egwkZKbEB498CbllqyRxD3RVhancxzOqIGgfLBvlewDAuiGvZ0frdAvXOg+VNa0BoTDKhRPPx
usohN1VNI/ZPnE/5cf3wnJvmZELhRyifsXARMrTBffJ3pYEc+7+f2rF8lnrekACJJ8wLmEXBzGqm
w6bUIaPrwpnZI5GFgzxvmMqt99jDp2TLu/ZKCf588QySd4FKMdxTWRtVI45MZY9Hnrw325rsQlHp
lO2zJ3Hhq3EeyJJ954gVAzCJXAJSllTz8Z7pwK8X+xX7hEdAbx44K6/buW7B8O2M3kram7md7xXF
J78dGWPjXJagoX82J3q2kT8TSCSOphLiUIQV544rvbMiVsR2wALfhL47tv5XU1YLb+ZQWIa4Ybo/
sVkQL+IVwiM/0kRmXaA/9/b1A++SiRGpVhdn7YOEDjgiXn9uEKSitEUcRjO3vTJH1FJuQSedRMzI
0DcwLV9Z0+RkJQA5M01BSdLQ0Ur047dQrEoe+9wv3IsOM8P7hPs+I9ed9RHVqeXtQdo67HVy7YUI
sAKNvtEJxWzUd99PMu5CFDME4rPOdMr/sD+odzsBsgdgK1Lk/z+LYHOIFg6aVMBIeI/ls7SxVcRp
JhOyX8njClIRjit9XduIz9Giu+njgYRDQXiMliTnjRqIjjIBnXTbrACUewVxVQmiPaqhCgU8KdUJ
zKoKzPBZR4/NJ9BCZrOWXIYrqVTulTNbEaRxk38tO3NMppwVfs4Dp38q2F8IcXK8JUm0GhE3L/GW
HJVJPef1vWVF6vLeS3TnXMJFgQZmx87T/XmBZRBRmdgC6fr+G3gvVcipv2def+75XNaw9B2kVneB
sIY4pLFxc5YSabBRBEEbAkuW9toGArrDAP0j+ESe+ZRpkq/XPFhFO16xX6PTzqga1+JlVrORE3qe
iHYdKJZeREfJ2UN2A2l2PjR9anv4zjt5AFvhOPtqII7Us6qRUTKN9It2sNuAvjlnveIgoamI5nU7
9y9zKhpkbx2fbEm9sDwFttIa6qUPEmnalbc+2NIU+eF5gvXQVve+l77wtTh+ydmvfMG4gMtZdt8W
ubnng+JGnXlTKo9/BuOQg8GZ3Q5KuFS51UF3BcDSUkAqWnLP3JrVvrUDj1fYIc9vJIfqKHRGEwsw
q/PBOzL0gV7NIqF2R5/tntvvkJ0PvM78OVhO0hyAQeWAQBe0UtSlAFg+xdeBhtAeI6ipkiBVaMx8
OrywFF/3OKodzq7P4mVq0Y4ZG8XEh1HVYQcbu/2w6ifkBB2IwuThGSBjWlLuaD++flwQH5If63Ch
iUlxirLitnZwBDDsaGAa4snfgN+xZBtzfcZl7I7SINeIVyNdTyzf0MyBBQwmk5+2cvNsfiia/bkh
eMLKMqjI836ouWVmMHm/J3bD08AN6ZB3vur50hSRPQJERo62Df+B03iQuVHpean8leGQJQIJV0Bi
hCh7H+y62hfaJ/a7weUT+D/UK5W83EXwaCdqe+OLroV9PSSdxyrP1SpALowL0wTityAU0CJsQIug
kQ4tXg9s6cUDO8WtKw8WSqjXLqzpEuz1BttIVabO+n93mS+LJPKZGOp+r5N+6OL+Wav7auK/Ulco
FgCGUHX4fmK6ezSO4t6dU73ifjmKN8VzS2oHrTNnti+qHpvAJSu3vecGh/FgX4zf2CPQMm8vSxF4
ZnwNqEZGGzc4LI4AzfzQ1Mp58HLi+CtvT2tizzzm/1v74ZcQx+lcPE7J0ZpHgKQLfhPWC81d1UUi
ggXXsJW3lTYg6e0um+seIIbUwi5AdsXZSBUlOccYrOHbKGu4vIa5WXj5neYGx57aUCFBCM320Y3L
NrO62K2pVsnSSZTzfcS76+s5pYtUnezUJk++mpz5HHMqA1SWRF91JvmMFUTU+Yui5t9Vlx4sH0LR
cfkf+kp02zBqK+tUemrDfd8c5hZlphTZwwYMHjiA6e3OpQlK6+YECl2xhkIi/NhOFG1/9PrRmJrS
nyMHd5Wgr2RsUmbJ7SW/rXMpLRbNG2HUqxTswuD/APSfx+q7Jg45Gd1+A2TfbTd9V1kLQYGGb1pO
e2II3MiVz6B0TBHURWh93Bo8S83iAut64Ma9pyG8ZlrbS822uYor/OsRnt2Ik7wgRcqX3I/nS8/V
nkATYrYvSgR1yozqetU7mSXDfgrpjEb2vc4Pn1BOjiZ2HHOVmkcJaYr/PLAl+7rvXXdjGGBGV6qh
sUY1YEgrNXxtyGyPdKng7qf8m4/6QykvuR/tQcJKVDEL6lkm+xjnzytchnmw+nrAiTa2y/ihfu0g
aOkX2nM4FzLCxgEzO4O97dpZCZ/tmEmspxXDSNexzpWytQ1BGHnJJRwPTc4xpSyMi2T7UzK9CSxy
m/kxYN2VjO8DRlvne6FcO/OhKDZsB1jFCabnldPNkQqFWSgAuQhq+XTcNB2DDNjZznFCKQfrTYQi
toZm/4t0ALPlgzdumvf0yeLQcvFrUrDg0zPCVZkZirA2a63ZoluMTWbzOe4kyG8HbUMrDaUEYNlW
KWHsloIt6/jqPPbCn+TvbovR2u0dr1V9aduUmQ4bPKTOR54WR+Y6QNcOYjlLqoOWRgIAMPReB0Ak
WTEAa9HT/8e+PORbxz9lK3PeNftuKiX91cWGS/geC3i/tft4eDt27rGBN6obs08fnZ4MN2ccaEBh
+mMVUlBJ/0NHsQzVGxuMUQxgVRcpEUWC4OjTJW8a5odA3F4+in/w22/3DngRcG89TpOlcBTe06zU
o1tQDCZSb6UPzgpwWIb1N9R3H9/Y0DJCTDRiRDUW/wIsCWvEpjlpOxg9JAGGVAtDws0je+SAr8di
1irio+vffd5NdG0BSzPd75WLWWWxikJ4wp9ijtGjl1mPHy+8rNi3qh8sU2TPGb7KvYJhx8ZlKYMB
wflJFATRHSBxX8E2U1tKxSlb5zOa/j9PZmd7Vj6cXpYelIglJijAHUPEpArcTtLlPMsh+NKsiwH2
s/k5R0/D//lo531lK038aLrQDrrrRgm4+486g2GS53AyxQnl6CgE83YHu9rQncYMSWuqclmDcj5Q
1zmbU8BdeKBl7VT5xzwYGK7aFtfEy7TDfvXs9puRrlTB+trreikYxJ0dGsBJXKg48uGPcxk9Waz3
PkCVh1eMsPtdL/ueLT4sxG+4NO2o5BqjMXGAzI/4atkrhRDE522DN/7B1uW8xBigbeFHhUQqT3l/
rNUzjSjiA5+L3ihPgpW4zIDAizCpLQB+RqaUI7FWrSxOSkamSujFzkItAXjpLe2Xns8A7OJm2nWc
tSiWqxVQkmaXU9VTxyKLuB/7aUI4FfRegBNFL+/fWR8/zRgSzBj9VUmoPh5yZUF0ZSPqCtU6UTcK
RlUWsEQAMBSoQ+XThwv7aDNv1hDIZHCY14awL/WyCfKv3AB2Yi739p5Fwm/aAGhmM5NqrQIytFrx
f0/Cx5l/yKMkVLiG/tx2tgXYDcrZdyW5uCHWyf8X+mhVpuld4MA6ooDUpg1ZVVA2yi8bDjJu+mc0
Py6ZpWJyLHuajWegp+QtXXJG6JwKkyyEhGiadjhOaS79iMGlvxSX8ICC7xoXk+uhaYR3QjayqdOP
m5KoKIM0RMGTGed3JYd1DTJUpAxCsgCD+Q4dPgei9235WIV3MOI3dxM6jE/1S7XY5/wpamtPsMyN
Mws1H/Blsr/g6MEsN98TV9AcgLhAbAv2yUtXrh1CmeyJqrZJZ0GgEKO+Rw8KH3CLpN+ag3AiJntv
jDXmRmTkpMsbKao4Tt8B3rd172XgXoNkpT8hURvebRlv7EX6MvX5FjbxbPTWBfv/QpOg3J4fHT6p
wQvilM34NywaSLd2ExLy03aKK64p1f3uXLXzmDQiwd5FfKicMtY3nbzXCeljS5XQRKK4XtJfy0l/
n+P5Z2lylTPsT41VNkc1br8BpDJyamY85ExrKlcj83+hfAVpgPZWVlh6FRwpefdnpvzDUyRtbF7g
OrCKRQLkxtxgYgSSGKMQgg9qoLrAarpeIf5YotOiXuvROzUov4LelZY1jgiWdcF43XxKIsssCdG0
8ow3nJ4BhRIRoW9jaImx6t0LEBbx46fepJqQXKJ+72FLk5Sr+Cqd25nKwonZWib3go8Td42Gnvul
yTsuhTFT9/m650S3wXpMOsN5Og3K+MjCDWO+LTgJGUjV5SV94SKTPbUB049thwG2BhuzJNVOhS8E
G63mT8XkSTU3cD31pBeptfJc9OWyrSXNBuOOSGmsfCnPSYat9Cbvd2ErP3VyPvgt4wK3FdcOgE+V
Tv5usPG5DvoLOZuxYXPMU53W36EkJH86qky3XFSgytUVtJsklNi54ILw5ibwmdA1lkormrj55lJC
0GUF35M/4Yv3tDuAgaj2mDUXjCkz7aBEr1U6DU/okUUZP/bUwpfl1dTNl/k2ImKLeqmhOcjh9UKo
4lI2MZCGMm+IBO4RK6hawQHl9M+NTb0KU9U6u99eWwYmhgb9q/o73txXPO8yU26FBO2R5jUMOExZ
JwZe4+ulYktRL7RsAxFq1nx/IPJrS1iSa//LS8TCOGQ5wE+u5JRfeQQoMKVjkXSEg19sU8EE3dEC
3rY07SpsjY/dyyXWLJTKriazykB1uIMu3FTTzTSuIowQGn5kN7fTccJiFWxjd8TxDf3JWHEk6Pre
+7U3S5u/PhAFneXsQ5oGg473953WXHO+OuaJAyhV/VB54IY0ynnRrDAiH3q7uPMHIqnsoQkFjSAO
6XB5xKXe75E8e0DspS5Wu6pVmRlOPbfGdslBp7SA5NLUCNr1mED+3BHcQ0ac0mBXJTyMHWWv5Nks
xJjIQizM4xE86Nzr9x7XiQsp7IOQRCleXq3argO2hM2FJ2UVSf++rIcMyA69ZaQCOfMSPB/B4Hy2
ma00DnEPu/NqWduJ3QHNADMlMJcib93EqvKte4ZM+A7r4iCPjHWT88bv1L9XJQ+IbRjbwIU8BpLL
Wbo6tAZNFe14EMgLRa7K32BFarRZQ9Flq3WoKM+XH+7/rSIalTfi72liGmNOgOsS9hqbrAEK1f2p
z1YdaTOBJnQbjU5p4EqR0/3RdJU7ZKcVhZSAS7MzI1pKIw3WkRMa2EQGxgu06TJFEwpIqpQUmrgL
30I8PE/8Lqs5vFZ+FcLdL0CBDeTH8o7GuTH+uuxColYRs6oZSjgKfUEaCiqaboGb42f3+FSksT0n
thydyrZKR6i4Sr34Y4t6ht5Q34jSQO3/wZzAiN7vCm0frNxD5r/3nF6ovlkz27t/Utsq2GSqym+h
gdyTP6Qnbu3lyYKxzNC92kiSFvsDqN5FxZsPsbyYxRJb8jDdR0NEdHVF73JF5E8VjFgCpEm+JfHI
DN/Snx3+CePmmZcFKN/BYC/pu2nDsipZKgXW/t2qpFzjeeacmYMx/jcFDPjcozNBwkLiFr0mSXYi
+/5LtS/fmpq7h7RfzRPXBC8m6S/Fox9VBRYxE1nghwOg0xWNT71w4HHXbCAarXRQh+mU4Uk/jQ64
tJaIQqJchsmAaD3GLVoj0qOZhqbuZW1Tn7oAJdNUeqNGLp6UIKqSCP0BxEPg23Vymtb/6EkO8bUS
MLIz+b3yt0f50nTAlys8W8dxFTiOWkRAWWFMMBPzc+jSTU2BERD1rcYVWLoYgYlr8NxvNuwSSVbl
uOUQ2hM8E9Ga8eK/XSZeO0xynt6yLFOud/NPr3yqNjnULWrdBeXaa2x7L08Bb6H4wgUaosbahHnB
yAI/fjUyDZ3PWcx/SOZ9t7/aUvbOckwQUHdZXGPNjtnA3+O0vgNJU+CxFYEJ6jgTLAeiXXVLAfNR
jRdg/OrXnLwmANwirfOPDYNoVDoq4x85ojDDrMNbbu0jbLPiovv0duApMgBOXmLAHKjUWaIhKsBl
lD1Dp6aAL/onzOJo1mRA0bNxN1wuJH2ExnOHSJZG9zIcmkAEd9xzrNvuTQ5CuT5ba6Jfvr8Oaw0+
bBzOvsCmHsQPBiYGMdV0QWqsAp9by57utm9ChgNA4ULUsiY2Fuzgn5uSFxMhqezZVGbtSMYWiBGz
F/lQCxhTD1xGdFKbhE7KcVrrfv7q2tVM5EMIt+NkKuNSJLf7ScRqEVof2XgiUB77GBapY4Pt3FZ4
VPXV8K/K/HpZ1EX3xH831E5+R3s90SGzg7/xsRorFeVBoUXQLs8TxGYDsJB7a+43qfQkKUUTgx4q
otK/5EbxBFNZ+CVAuoRAne755WJcf+BdhQurVmkILL+luxvqJRF7uHdSrelGCIiZh3eSv3Ala72s
T7MlyLUyiMPXMt8hQxerpEJIFmOiM/VsAivdJ352A2olRCxhPZSll2FZ0AGRqvqcYFQK4KePZBAk
gwCBZzJfzKgqCn/R4kY40dyIul4LBpppIwgT16shFOGc/PipqjP+2XMd9s+fhRLmo61fElFuk1P+
6K5f/k5Qr5zY/Fs+sKsLLtMOwn7Jyf/HhQYHzDlTWFqXP9D+Bfwkq2EbIgwNwzVwDmumgVB8OO0Q
gM90PC9+5bDrJaZpeHT2Ao6d+lG03DyXZjIi66DM6xKeKV+kk+D5CtXU49vs2H6yEoogfqvvX0y+
2t2ABRk5dx/1xlwmOg7Livn4RG+0+Xqyx2S7zyqqSl8g1aP/Gc9Gf6MurTefT6aYL3IVRc74lK8k
JxnrVm235L4/JmAsGfmnmTDVndv/krP0SdhwtRrYtiU0Jiq3aei0lAtab6XkrptA3v0PYSAv9cZn
Lam1iaoOo2HmYn4gP6dWSYlfpB4o5Tiuw4feMvYWsCSrn+XWVBu8exupPA8dyu7hdmt/zw3DBd60
nG1vSWNUh4xU3+d94bbgmJgFk0i/J60aSXmdahBKys9PTc/9uj0JwiqdZDtH/Rcz/aZOeP8QpEXh
QDVZHg6Gs62tsQI5PCDcm8RCOHLgFwK2TqkREhqcY6NEn8JvJtPoBHsyrU1kygPKKm3NL/fzbmPg
VKQj2WqE58+EPX+3Y568X469lVZng5cLsdDmwIiO25tyAGXQQVxOpMl1bSrJJgnVoswovH0/9FIl
VGWu1n6Bpa7e54iafm0tlB3xQzT7EN0iPkJP8gSz+VzwNNQO/1qK2L/IyK1J1XpWHv6+D5K7886p
4uJyhDgJdAalukd+Qr/pdvpjCiwchkJx3dBKGREFxgLI83fG34FNnY5KiIKvybXzrmLm8xV3Sa+s
0z36E7n+RTHBlWwYna2Iz1672FGZfuZNellz77P2N0SaRmgO/GCjJM6bbgD/MOxrGxun0LryBRGd
SP9o76kVcNkcd2em7QY3ihop3UH8tKySj3e0QDjKp4hQFZOBjGCS+KvxBRWoRoPlw/S9hkZSBv9U
u+7UrUOSnQKEz9aJw3gQgbyOp9PpfRyGCjkmcCJO0MGZdBXK9qy+wj+CEWhH00naMAPO8uTgQGjc
0IE4oQA2zGwO3gq+QQq+3Yhq3yuKUbPf2m62EVdSVyR2y+xgiT/2J3v8Ji/E6ACr6C+uo+hdWrUb
pYNRzmwWFVHObbtYz6PVjF87NMXqEZXIfv1nL7RI/sg6Els5zrX7GHOgproq13Xe65/HW5XQvNYY
r+pVRoib8hSe1brIfIZRSb+urwPo8MzxqLd+W5w96ecqLQpCdsTEtnqRAtIMtb06TQMrizSoEjNF
waufLpOBBHmctHlq0fK9sRchjNj5H40zg5FHxF7VeD/ec8XhyRQNZCPNOOIpaWCcmLU3/S/LyCs2
+cv4oMiOfMejPISXW+fr8U8no29PfHnKrnqWO9LwzXOrvwoTZL5Bori318lUCWdEyfqtK3Q7oti4
/SyXPOjU1PsqM60cf7WXsXDLQJL6Y4eLAcxyEBLdhryDbr9BMnp5hkbff8V4AfkLwwJUEiOKE6LD
V4U/a8Vn+AQZjlZtqiMeiPwT01bi3os5M6BAhvCaP3sPRMKvXMGWlhZJ/HLKh3ruzPGxQthqjtEz
BFOy1lnshVMPncEy9a5OFTAboEC+/TujK+DMXGsVBDJ/frpeQiBDCpttbeFrVzCZ/vTQbI5gtZfk
5h0ctrfBHocgKKGHUPOKx/YC8tlZvwCiWRTylfQbOWS59SUYD/vZLUclO9x9D+L8dYe+5GXVE+w6
dCT6K7b5Rr2gB0L1TbxvYtizUeyZURLQOX9TxbXcDSaUchZ4/q7lwn5QnnNFn6dPXnlFhrywSco1
F8UaAdqEZJ1cbl9f2t5RJpUVYs+wml5pW7KyBY5ok9MLlYEiCyoko2uE5x2bDVMZ4Wsis6VOtrpQ
Aupum2NOAUMOPPJy9lvHd8TfIy7XwidaV0nZ9u8Sp6kbLPhRAYBpi6Dn5F6O8S49qBS8aad8d2sT
IlFmpgGgdbNWBQmJs6euEWGNKGSBVaTG7h1WGqI1Xqlzj0Yp+Ra98qA9oZ44PKWLCYWmemnfQyN4
7FenZxRCQg+5UUCvSRKtI6PMZgNzEYRPlZ/SMUVuiqBST6jc1r01qOiDmcD78ooutZqRLPZ4q31/
f6002jefXJ21bZ5gqIgN7Bh4CbsVNwJUxUVbfnxPjzd4aMKe7JBBzT0uTbnbe6Fvxf1lyfngYrv2
kJCsGxdsB6/6mAdtWVZRL7qmgdUU/9WxDQ5kPD2S32elV854sioyaQiwkHq+dRCpar2hRAZW0dsm
DO9WjMfeoF4iTKSo57Ko4STZzBRDKeys5FXt1OyGMgzqs4aTR8gijMS0Gw9jfW9OJ2Qkj5hO20Ck
KiefX9rM328Y2pk1vRZk2MgwPU2JXhAMU3xWWINh/0fxwweO+ujt96RH6rIjoly5eNVsImyZtZEu
SlefgETJwQcjJSa/xBZZUNdWgB2sa4V6cr+Mmk5ZiWwMO+FXlzxW670ZYOOSv7MCzMtQXmFfxXje
zuCg8anDx2cSfJ1M7F3lqpOORlKd3sIUULObCrGT/ruckcD7/RZfT0ipKn9QM8G4ansEEBNcvuMO
xJPhZ1wHE6utnZHIC0xJSvcC1xHFPDkNjw4K1vtjwDDMOGONGxxBZEqUs2s1V3gobtVAsNpRJnxP
+yma0F8+h+aGvZcm3k/mj94LUJUMWUBPIEqr1Wn1DB6alojWtsf8MFRpOOpDLasOMvTPOHj6MYG5
IFUT2dsMO5fYWTOIQRTDsVG8LBjGL4aMsDuexAu879v31Nyv1Y2l6OeOSFp0leuyHECvV/qK9ueB
YV71M24ayutAEh8Kbii0MSdwvgfyHYW4DlvPcxjjnvxh0Ih8m7k7YSz9wWffNlXhqC/Kz+Wm6xxS
Ifsl/ZDCiMyVbJ6on7h6OC9sdx+FSGzV6E0d3Qp2oHYJwH/HV66j73+/O5f+7D2GeD5+vrXkf02M
5y0GGbhEj2vfe7f7Wesv4+o6TVZEbj84RgKjKtc7+bu5P/lswXg+G0x7jM5BNNyX8AkIO4JB4iIo
WrqSeXOOsDuIAkOdfReH5yDphD9FGjXqcTYMH/gVLI9YF/0dCapnNs6APm8uKV+dwmLIpLyAj/qG
hQdgigwZsUSK8ioWGoFcNRz0MYkL92VYG9zM1TL/bi2o+HzykqAKU0FOo62NkGF5NINXVXslfdao
kzccGpmYnu+HbvFu13liRMkYEQh127lzQS7VbKFetpYCNROB7ZTLAyVgzUW8lRKaKWzEZneiiXS1
McPebI+iXSjijUTaPAAmJsaZ82n8Sp73FuQiTU+5HcHV3VG1fAU8PNIm2gAuXgCg5ADbW7inLmJ9
eIfVu0eo9mhunCBxiMfqOBzcg7U3dt3k792GA36bngAFSESV5+oc6YNpE9lXyNrnnpLwt5Te21Nm
WcqXojssq8/DZDlxCZZXV08v0nj/woFKEbuEM7mPieNq69QtOnJaBW/B9e1OndfYhT86RLpdnMlA
6ed1MmydldmbHfwR25G0UNrF8oiIS0jkDwIHhs800JgR5WTURk909+BFD0YZiBNyacSTOOsybj49
D9RHmpSOOtsJ8yzieme1fWYRBQ31p+undqtBor4PM0PYn0AfVxrh9uJqqqRyQ1rfBgASstscs+Ye
19QQNwO0V+ag76/V1P7Hbu0GEK8qTMTPMXFJ/EpZp78dE9uf8KBRUzR5MocOBnN3zTu2WgdblCyD
hNpDmCFbx8FrYu63Li0362bHFX4AaOR8CauLIbtwfPcARjILfwOrwWoQ/lf0UrxWSqU+mRWSiapQ
zxyJ1+zWDFiVAzhm7kPNY9OE2RSEmVnu33y83g3zL7zpllwoZTJEred4ZuEi4hBVIWKA1EJVcqZK
yB61qcNVFPsfUhgPzdf+GjF+x9/BWmC7iaDG1aJpV8V/ezYmht9uMxnYG0sWrUWngitn4J7RQlPP
tzqKdZ5fQVE6PpiSffb3CvzQN7Mav5mr95grcCd1Qz8NaDqkwl3uXpjpsP0d14Hszjwv7G5+tgPb
Qa3wZRtbBqWPOPWZ4ooRxgrMn0NS0ccwj0I0tDHaWzqjAe2jl1IsFcv30rM6Nr2T21doTxY69qay
l/tGAAKDLfkJcfgX1hOZtPwdRpN5+I/+snNg5WojPx4e/ZbN5Ji7HDunukkVIftXWDJp5Jhi6rs4
rUcsX6m1P99iW/rtYqdBRBSKYI+Vt3quGyVn2xpVIr2LGvxs+vwOy3VFSUm6TORhz/gs8rSnaeIV
1Vjk4mX339vLwgC39WKy9IUCM1KJNfh+b6i/VhaLhxVb/p1IBBa+m4filmjwTidYLFqfPG36hBtP
OuDTSu8vgF3BK9Heg2pF0KAgWuHb8ypLkhNoF6cWaQudDbKD/S96YbiWBtmtZG+f+Idia80DdSEt
a8iqJ2drFFOgiH2k2S4pw3hFM/us9suLf+5jbfN874IRPzaQbWwVea2AikIRaN+T4H6sVXAUjuHt
IAwrhH+RjqCZlIp7c0hayA4gVVaHqlrdySQWwHDqEygFo2YPYgkNhhtMO45ZvaLTmlc8viBM4QdP
yYaK07xizpJhSlHnwnuerRUs3C3LfqMXq+Pf3ERlQFxT9tEp/BnXI9V4V1jQz7JOGJxBPS4FgRR3
thvKzPOrm23bQmG4PbULli3iXJvFQ+eBRbl17A5OST96hGEUOHUG7w8qY+QGEfU9MhqGNZDlsJ8M
forTSnpfanoGyTFF2YNb+39s5gPkYR6JBCzjspQaQqJYpSImRevxVsqVv+e8MYzagH1vA2M1JCux
U3jMn+Hfz+kSLgKiLu1UIS+iWp4Vz5kXxPdmXrcFMPQXYH0aLXaMPAw2aIeagc0KUmSGs731WkYn
MTnO7jNc9PpyiZD4ZKGWq4qv6+gckbyiZY61RIRr/lT39XJBAjNJ6xkoPeORKeLwVe11hGNf/i5N
jxkUW1PYoKf96+CwySUQDALogAnVQ3B9FNgwP2maoUMc5B4mfi5b6nnnJ2zyfSoOXpr8Qc2PC6bv
TnKLLcQPr1OG9VULfIuitPgoHbRI1AUiKCQnw9G71QAPxKn683kG+Sb1KwgtdfKken4rnsEo3sX7
5MLvAKQWn+0AYXc09fblshanVIkRRdQ5xTT2cwqQUgb1ewgbY74JO+ofVe9vawRjM+/jvUMGFGoi
HYD+0TDPyMsY5fb5BytkHHVCv3jh8uJwLmJknFeL5ioQoEIcemcebcqb1yRPxPj/+Dg9tn68J5l4
IO0vPNj1BqPsOwPfqtw9j6EWBBOAs6PpAmeWw5JkO1V/pM62fnBYTHJ8QnGuqYsnnWb0bWjWlZM/
vHeIvTH6SKq2APH9hCvQ6jpPLoUHqVsSxeEb4A85Uc5lEb9N1q0EH7S3jwp7SF1HDFPHuheQWTIt
6fw5K5fxkcNmydvazGPa0qBnzD/H7sKt4gwMzSIu6qAjOZuNe4xwGmzBmdYVT6ZM9N2AJCiJNoof
sT7qgZZxveN+DTAPGoA1nz2asmm6kPXguXWLDjHQHEdySipjpe4w2cOM/4jKKIUWPgWosIl2uZJY
NtjSTsE2hTOOmw+NiVqvcPDZoQOViwiU/FaB0mGRS+WhUYZw87F0yCoBbq75JfYgH4BHh87Se7Dk
NzLUJwDL08YGC/AhnBrfuzbAwRQd4s6TJBnD1tge75WqktYXtqnbDwVbm8mmhZ22w/FpLhxxwpWU
RzYaOHKxTWsL2tpP+5AwgNDJZ2nq6pFr85GNaSrE/RjPtC1tqiPXsh0EQvQ/pslqO02Awp+WoFO9
HkremA8ZXez7ay9mj2bnwx8JSGMgtxQkutH9OfOmIXNCWdNooTz/B/nDXnITVq6tc6yVnvpI0PHy
J9V4uEiGeHk3wk087Xsh1ZSOZfJa5Q4nVh+U6jAPdarjXppl+v8dfreO1v4EfWjG7mKEkh66/Onw
CDTYlTdFc409beWSeS0btoVSuX49g6yCAh53ig8yBFGqxjlIrybBeyqcC9WGK1+NH7fb0zcwbGzC
/ykhVOmOpW/PZlu9oovyBHoIT+ryKlqeyAn8QkbanRthhmR3F2VpQCAHFemgdewG5k/nES7bzyuP
Vxzeg0l/dGk7JELMiC3F5R6lLD0RP2jSvbF51V7rWVLyQfdPp+4yRgP7W07nZ9x3CcqAj8I6Rp47
fmYzxZePkeSI/2a++wcg7NLEwdG77O16CJszhbO9rRM6YpAu0dt5c5sknpSCfO6jqdohKbqT4T+/
LEgGqgcTBHO/8VmZnvwa3eSGFAk3hPDzpjYWNMXyKoQ9YqwjOhFazAJiu1lsGbELSpRL12FgyzDJ
HhOs4WfRv903iAjprHmGpSXjkpgqYrjgA321lBgECp+m+t7e/HWk5i2XefsItnK4bvOSj+SXTkZP
Q16+YpAcvrLPSH+f+yhZJNHFETLTc1I6lFKiAS09OHZKkJj4HaJm0qRaxxSjhBPAlRH+NiL09jw0
7K2iz6ERd1Z3vcsBEJnFbMntKUW2sVLzGCTZtJlE4lOpMmEUhYKsYicv/8LrYw+KUkqxEmYyl3/L
CzQzQBv2ICgQFLeWGEGrQvkAR6qJBGBY4t5AeySi9kdQkTnMBk+q+b7vrGAx6/RdVJITnaf/ozTs
yDvScbkB9qaRAMkViMqA5a6d2lI+sn5pJ0ZByh2i/SYMU1fOmcNeCgEFEjRxCALbWM4fk8QrGRsr
hDgoDSXKzhkhEMspiiRRdbFUDfB+T0ZWSQlWCnSDAsCySb11+jG3AlNRnHSLIaBa6lC96GUFFu0l
R4qxKbAhQeDUejwyHhrhsImxDnC96LjsJuKmGifJ7jOTrwqyIAM8CA0FqXHSmCZBDJqyj1kCdB36
D5u0xYcI6MSdMKLwHetReyB7ayHNcflWAJaHLayEIuupYOoqVHlxndVrXIwb6gZyl95Jemq+UoY4
90n1XA/dAFVfZ+slemq2AA1VtziiMWchMz2YeZkarHhGeUnXZ0HuLiLD2/iAaIeV4p/KtE9g3ZbR
BF9rfEiOfufiUmnL4LD5Alf1sR0mngK3SnmzFphOMihGL3KyFC7K09NSyRO8k05Rb/CmJz1ezd/+
tHol+T7LKE2g2weKCElm/ErZy9uCYxYUpfde7JznppKgqkV55W1VAIJBOgvNYOMbAn7YWuH+06yn
hA5QKku++rE2vXo84+6Hina4yXsroGc2IeT92xXMVC8f9m+UfibhyvKIYCzcDyzj5GlY6O9IaR08
Bb40ppQHXvZZMavFm1oj3CeNVpYB2C0tbmpnQ6RuoaApL1s4Sfv+g8DBCiFbCN0AZ2iMhJTxT0Wj
AixemJrKor5wOhtATM/fgzilrRXdoHv/wRQgvQz0djkpeZeabDTiEGdZMibL8YJG1Xr9fg6Jw8TE
grpAo8yMWdTtQT8Nrcd67MJTeh+7mj2yFBq9xzgx3L1qrrUigY0bs3yVhE0qXNlO2YRLczjGVPl1
eXWOsv1QFpepVhF/Po7AkO7JGVKU6Z6ZlwsfMdH+4iQVzxlC0FFCe9W4+hcvQ7XzdLYESRFqVq15
Y6HZ1GUttGRo1x9ALGLM+f5MKQwknes82aDZF69XTMQiNvRvk8DWka7Y02IUd8USn27bWu8vcyfS
9Y6ejKvtKl+x8iqkq+tYDp3Ao76AAvGXQfmhl/tDvYH75DzyBR0SMM79FPZOkumnqZl34+c1kkYr
XoxJjfst7/w/r1nW4y9CJpBcihTFkz/H4Io9rObsMl9RrGTLGUOa6ECRn0Lpjo5kJHR3Gfy1+3CE
e7q2qtwR46Z2sISx87L3xhq78SEbm2PVq4ig8gjQxAah2jd7WUaYE4zHKY9dyT4kgRdZyyESWkQ8
7MzEhBiR//+HWPxMBOVxM34m6D9kQpDceHyUOcWw8m2nQ6Lf8yPZ54f0/LFC6NUT17iThSJ4z7Wv
bbLb0GSlus27uj/8mecAzpgNroen17vbbHF8O1l17q1PaZJGxZ9xHs5Wxwn3cvpA+mlRmCoTcIQ/
H1QZR7y5D2wO6wOXqZDVebKfGn0aUXsHaomSX8zBE6krtFNFbkz4f8ER1buVGs436MlipjBHSn8K
2scM+jwCWYWK+54vW1dCnWIFwnPrNh+RnUJCoGvBkpDz4X1TL2pyBgvIqJj86eQLAI1dnCzw17Rg
kCA7/DJDMCSo6jAnDcPwM6rELrJd4wPha5i2bgyW818Caon/vhCNRmXP/d6G9SYzFiFgvTcSbHAD
XjbADjehTwZRQHTdutiWibkye+BHGUt2Q+fDFSbrMZolhTkb3WN5UGzrhHFl3qkY9bY2m8csHcTh
V74ntmK5uWwnZzeM+uvcwiLlDgP0BA2nTek5/OjHi6T0ijUQIFKH4P+O33OPBDgA5OdKRMdaz+Sv
+5N8KNtzJbRHm0M+PZgWq3nZ3LtZQualDFNVMn/Rz8w7VfXY/IRPXQDLJoDLAKGBg+Ey4LHb+RGy
f9PECIX/B56GQfbmWOX/egC18YKF68xa1IMfbvh7CqodhZwljBegwphzJtKUU3iCzEXfFuYxWoo9
ZVhQpJQXzcauPD7EqEdNMibB+EVp23ihlHPPn0X1bi9SY7p9MNbnS6IVNoGd6oqAgWRYm9SvWbmX
RR2ZQrsyWDqQ0p7Vb+P8ahpdWWShk9ywD8TppBkl7DsULjiB9fPbCimnRyU3OiCtqv4Qbr7lG4Zq
OFihcNa+g8jqVosofjB1z1N0Uu2lp82VTaJ8lPI4Iu3KMArU3gCNeVOqXCknacIornQ6kV8H2t7O
YNB3exS0c/SEnLfFf1SnfcPWtt3RQMrMCTeZ9bON1VhLxtTEhaQ+yH401oInaE/NUYqhT9azqdUU
GlRVcu8ZeFHsiJn/OPAWkW9bHu0qlUJdFdqOybYJ3qlY/m8BzfhVeCw/6D4SuEIyhhXxz/ddtcdI
ntAO+XTGbYTmqIeo14ie0HgDzDMUu9sCHllIiNiD3+YMT2OMf32k24YIrIXTqSbNqKIrx1fnurXc
1xRNs7QeFaVuuLfQc+zxX4dVxtrZmxTDTyfyAsXKO316hHjscVh1odgziosH0e6XAIOqi99rYYGd
x6NFb59AMnMH+QvxNwIbwDort76xwdHfv4lGzLRXy2DR5tw9aTeCBgMe5Sy55Dd78h2LEhcNXhiC
KydWBF9pqkYQxovk1lJnOthQVz7MXx42Qn6CEixqKih/ipyThu7KMROgy+dsF4Z/jS7A/9DI5hDa
HBgWuNEESOwP+Uwl7mFk4h1Tcm8p+uxcXPF3O6QZ6FJYfP9bMIgIqhLKDjBhcV3kKLDMCC2RASZ3
L6jwwabIxKFrNzQS+/gwuK0t2WPahHw6ebiKupDfGxlsfj+1yrY5jYSaRwmlGa2w283cBP3F7Vsm
T98boojrpTyjJl2v/zQP6NVGpWAueJCiHnF9cVwMyGxrCcDwvLAJ6PZHAZLzPqPOHjeOnwtTd/nz
PDNCjcYJ1UPupCJdDWfawiezzbGJ2lAqLZ5WpzWEGKc3jhNzHNv4j9dWVKeBCcLy2ADMp1lkrgwY
SwK2eNsuikPv4Gf7p1l3v0TthyzRw8I89zQpWOlICvcSXch0lXCk9/D8t8ZOEU/8IZCqiHMJrRzh
Q3cE3ikfu+JONtUw/87xtMb2pL30sFFW6avW4Pp44hToT/5feqU70O+1NnlmiuzA6odz8VAQtg47
EP22AFD9JGAZSW5W6papRNewUfciF5hPojfsDwZiP0cDjecr5Wp+Ughda8gYH/zA7ZWHZi13c+lc
XY/L5XGvudhpem9NHMu0dQb25GXl8gp8cp34wF2qeLyowb3CVfA4fhaaIHOUiqvgpmW4U9L3yfTk
Q+LDynnIxBE+RqImU5E2kOsrCEhvs59x8f9xhsDxXewZ++8e+5O01KxLl6AbmaT1+fNVIMcQBlxm
Lv6g43kGyjvWo8Zb3ChUxQIwHwo5+tX+LR2Jkbja9n2rSLAF0TQEflZ7el0OnW+9Z2t2UsfXOYwP
8XJ5oQ4GcGaMM5mUpu1xX1l2e6Zh1l08hMn23iFYsL2n2XWZyd2rzo/LIO1YH+PuvEYeNB+J5hQs
y7e2/MO4n/M6ACPtIt8+XuxYIDQx7JrOuKFRdpjuUQ7321XE9IzGjGdQdowlONrQ4LCDudbnOJ54
wu+c0rhaMxGl0sBFq5JA5D0umognLXLzUuEhiLoeLRT2bpul/M4tsrP2Kc45PD0gdxAsf5IlcPe7
Q/R+tfZU0w3CyWErCaU6zSdRC+K1PBXYkdq/MXFk9U1SclrKbcNV74FhQ+CeuOpgZuucUPJXS+Zm
AbT3oZFv1ZLDfgGTIMUQRYFadoa7HfXVBi3JU7SP93N4DNkcf+2PkbtMTb4YnIS/JBtUGLzTEKip
FecJRrUd3/cP0daVDMOIDintV09MrInb1Pdq07M8j35kUFazRjSNvHrNtANIDKAz8ThdZl7urECr
qLW9epABHj6kGooGqc3JT1PqiY0+02RqsAEPIJWbB4ZOO3U7/igLJkidb95zYlDI9lKHzAbD3Onl
Au7QDHtFIQdQjFSg31B3LQLwDkO+pFqt9H/8m1MhCmM1kV6GUtj7fHVrz47kxSBtH5iJh+UFaL02
oGgo+92JKSZYczX2M1Cuew/i48WPPmyQQAgDZ9OBC76L1V5kUD8q3TRlB3V/Ee6NCPPnPlT5wf1Q
GfoMbRT1kIcZ1pkxJfmYm3dsHQe8NRClyZlHyNQNsKDqyz+hccrVq6Mw2Rev4qtaXUPjioXq/iBQ
OHi9F8Zqgpmzzzq4afh1fluWm9PCo26Gf6AlVnG5eb0rqRuJdE59iVOw7FQHaYlKAvkb1rieKHMl
svqs72OWATe93Tb8VMJ5sa9x3fx79FcQgIBcHrYwJ/zvwtyjnkRPCsJ4DAkrvn0/uC1ZsdbUAtyw
UaMC/umKpPJ7j+F/r2rJIzROkNpGoQNt7ko4CzygMS1ncdVBBKo7BlXw0wbfRmhEfMjsxd54bDna
qezw1F1xSOvJdqh5h5Hx4ADV1fQgEK/W939EXcxZV4Pd3ARh7JqPbiiIPZ4eeuDF+DG51gD0p6cL
pC6y30fwV5R8n5NGvySEaoJY1mKk50ThLuv2Kj4CVzpk+CWGUkTE/ePemOwiRWxhbm+HdzYvRPdN
4ctqcSG9gQuhvv8YbXIc1AUb6Jo3FuCtTAx3RvxUbQ28ORiMEkJKBmwt+ej3FhrwB//a6qwO1kZl
1CKoILwb86hJUh6RjJ9obM1yA3UDelOfF+d00axuECv1XGfnvVhVGftHLYZCm2Tv4ChY0ugmN8gR
vOkfs/a54xBbrUQhhjqUc8AdonMGFuv8FYMU7coV9ugLKl7kqLv/lXVAwO5LRImH66BdNT+oJkKz
jq8GAJr660oeu6cnkFqUl+DpBNOKtjOaUHjKrS5SDWPWokRCk9lQECN71xI51HQdcpVm0S7vwZ9Q
1kD4lUlszpSs/9c8b2XImkRMSNvbwjnP3nAY2YKb6GcmaK+YppTlfwbJou4NlDtWixZmCM/bNDLl
n1S93B9ihxkEEyDhxOlwgwhIn4TvK9+BPnXfVCPnPlvGc5d3TAgRLYQVyO7FGmWfeCHcPD3SaK0n
KBecX4U+H+RKiEuiKlGBTFEqkI1Ls7vE4RfQBlUnYgVmVtyWGaryKMl0BrQOb0aaqrFzYfcz1VDt
S6TfKpF3aCfc/CJMSp+IJMcQgqfcHA5dimzYU5225F0KSA2hy0m5m6DJO2ohfaqH+ngpKOo8IPKJ
NS7V54tjOS9FHf6P/1XwH8dPQA/iWTnV2MWjVdu5ZF6X4hnKpy6pdF1mlnLRz6Z2csW8HFJucTrQ
dQCCWzMDli0M2QiRaQdkLawLgtt1zPCKHG2N/IsPBNEJfR772pZWhWRsQkN3SJk+LXGG43e3OWu0
frboixmln4r3sLl/G2CalyaOafHsDatVldQLZ24Vhm47kKvVYIOumrkyLQORJl6AV96WI22D3hvM
AezcqFylfEDqAUPBGxHGRQlemaGVzqcyU08e098Y28WHt9luLeJAWaCUFN1WV9caVd61m0kigzZ4
qoCLxEHn3lo5ANLK4wwL6nPprcktrprXFCCPGxu201elJJpuBCGiKmZrwowj2GK+t8CzYU0TkyuL
pVq50+kKVr0oAhPxpIxbVmho0U5jUvgTx5fP/1YnDczBkUJ7zW5HtIkDBjBLYavV/xDT36lue75y
Q1SE2PsvJU5yA/L0Mp2gzMib2BhM9f7H6xJ7N+dJSYploKw9aSQVxSijSXFvxN31oPApa3F9182K
sa7f0GW5NDc3X4FadwYsQPIV3NUAv2LV+Jq8WzzFFx+GhoWayajMSbtIaPSThhASyDqmdPrJgADa
bCW6N7hCevmxKXZHv6dMIPmATth3R+0x0WEb1mt6eX72cPBs42bh2YbOouDJUc0b0f+e+QkBoDKb
B23LrOGXKxET0LC0hx6bhaUCsamQI2ROBtGQCtwoAyXu99O5d3lXCgsVp9iZi+uNqcprgA3uTnpB
/ERSyej76Ye7+WZmh9Wm75cdGbLB2oHnHrPtHQtt8EIwaFZRV/+8zWY0HbYDtr4YE9cE6IG4I3wp
c/9z+86JnZbsjMI2/1fYwpYL3qGcdA33TS4pj+EV8OjckJ4szzb+i0S1lN9oI9+IeWFr1FsAiOnP
KAen/BFXZ/dTVu9qIGZMyLG13nU0nJGT5RP10lFQdxxPYYguiNAttJEoa9KkJ3BCr1BDYYVh+FWZ
puhitv1yrUutlJNaY5nQo2zkmN394lXfbMxeuOA1Twc3IXBi0UlrGrBgAgSF/F/QhlwZ2gCN2wlM
tgXpB5bcBSxIrKcBQRPgdIviM9eJBFZXWPiDb6ok54duGDvnLsXgXz1YfYCtEV5i5br8w773pJvG
lZrglFJEDC2aKE4SHWp2ZcqymoAGzr7DyqOi2y8ZQhJftI97GZLqemNOX55+d7e+joSjW2FIXqTJ
l/t/WT5gNM4ZQ3rFzFOlWXxMLLT5NZTB+1svtQavZkM+c7LvSBOpARq9UJWSVOqKutYKoCRRI8r3
zcjbavnh3euHp9iDHuMo5IjFY2oIBRRELznhhIDv8E+jY4pIlrBRc+i+OVg9KLwNb7M0YBeFoSux
8O388gqDnfGNjpOqdqLXry2B6QgPb2f/Z7fGYX7do3g15MGTdsf4GWzXONB42MexxrR9TZUBLTZJ
mRZq9Al9dzhccGyjK/Z4n3E3sOPDa18fEWQZDnp0DqMAGVvz3lvJYiKhQptffzO6vcE0aoPwXn3p
XYIanT1ioD205xV3/jYjQIBtbHINPPLcEp163ftGT5E2Js1fOeoGhla/kz3Z4+WvqLADVUq5aUGp
owNyGAk5at2uyMLjJPFe7YN3urmXr8WpS+HnUPSKK56TVd7suIkhwLOaHdg335sB1+dRm6lhMGLB
r6ozCEjSA0sZrn0FYXQasHQbZCH7CYSYfv9iUx5Di5e56aU1F3D0RhJOfge+ICusUdt9zAn0lHKk
VMiegn0gXMQGSt95iqZJats4i60vth4QIyhMGtloQHqBSxf2o0LnJGujHbugcnRmdZPIBePD3PuR
DgMBzyqD1HBpgLXbteLhlVt4wBkS7f7wXaqzrDVYu0tQ+RaHvpIgqEY4T2+8/GcGZJgnywHDyeaT
3lTUpbCFZqvKBvEtGPIjZxIThu/XXP4KZVIzFa72j8w0pQw/uMn/wPLkgu8qY4mZycN6PXFrIIEi
iDUKdb1bROJQ9TDh+wtMwwWtdhoy5Z0Wt9phXcPqxees3qw68h/vFwc52MnRG31y/5hrk+BRT5vC
8kqwFSSzfDeHP5Bpahj3duh9FZNNiG8uhZ4OxmNlLmaaACvZZ1jawlmVLeQfsuhdKfEqTo+LNHSJ
A810K3YsaE6q13x8gE2w07W5VUhZRBNnUEDukyvLABDWCmnsCVn9BRnh1EdSVSLWadUqVA84wv1e
E8uTroMsJCr1220BhvywGLj16mWmrW3/HaDBeXCkbGjPYES+wVTuF6X2iRUPhy0oJBt8/+cCm7Mo
G6yvkTHlV0D1rQg/3tZmG86PPjq5po16E9DmvX4sIFq5A2MnSwkEUNAO2LuO3T9oIx55kLrtlURZ
wzDPmFs1a7Lr9fzN6390yPJqLH1xGxcDIIHMIWawjp3/CftKZGU0rSP00aiIbj2wDTc1hOgbmupy
LCaxYy7H/TmUAQTQ2FYmCxCgT0rUGMZjH/lJVfpBbWSCBGbPNUIDKUIMS98irZMtOkS9HQe5Zyj0
tk6bQcOSmBgTO2kqx16fN1nAdpTPTyrIshDlxPOkSPd628wH0fKLQAGGwjeyhokJiwBn0eBsDPFF
BvHBxu3z6422mVfUZnZ2J0cMvDLVD1P6vh7rpBHXkhHh9rZimcsri6BkdUb8CUw9B1/mpUnRg7LN
BB369qHx0eR1S4yGRePBMJSTH5ngIAfA0kgf6M4d2xVpEXqRwu4iw8nu6bAmOcL/nxlxwuQ+ZuiO
3Q/EubL1OnkRrdztX31PJ09Nl7Ywt58ZNcAI+l4i/buzzAI5ZJpPc/RhIqP3WFMs8D/0A51OEjQB
woT9bqySUiUHGS22ymwE9EWrgLfgR/E08oR/Qwu1x6ct1/6oERtwq3QGMLgU5s1ysjtWiECue4wx
bOLJynb5udvApBEcSNmWdv9Ghbo0Dy8bBWwbuDMwCwLnHi6XkeVVLS2qsJLGChn+j3HVkWplAwDS
Dr3TY5p9aoNMZ3HJeEHIEAmpUKRPSFdvLluE82cIFJkIWzIxVcdKKt/WAmQJKbqYyTMmZmPKqQez
i7I3DJSjNIfsWvFz8lr4t6NCyj9cKrhtH3/tfoaU3DWzXtTamCMcVZGZdl0VbKHucmivGX0sy0WG
v3t68FYq7/0TwfwDkazZMwF8YCLOhJgw+jfGWHG2wWiaK/4K1OeU/qPEufd9F/lvDpO5yfCLK3xz
lqgIn5DgchPfnvHPjwsRyKn9Bsi/0hgfgJmReamuarNqYQMCghcINbjJBFqusfgLNSjfJpA+1nM/
HyXUxryER+PKNurtYG8DP1vbJugYr2jWEs2//36SKVtQ0K+iuro4yaKw3dTaE3rFbrFlHzo+ocCc
fa7tRbxtuqa4IMzvdG7JDzCMsbJybEjnw6Yh43pt87M71LP3m+Q3sG9hGd9VDRwOeRIsYQ7ZEKtw
E4EngVvIfsNUhBiIHGp53XN/EALwSJUow9suR2p/ZlnO9uivYORWGZlg21uFkAUt6fo7sk/7DKHt
ObUe3yP7ALZQgdRpiPUjely/i8vmybKU4/s9VNvIyWlHLzgR8HJQPZvzYx21bh+wnMGspzyAy+fl
dQVp28EImabGWH+2roU7AwodnqQjYg0OIhjWamV5IdochyIoruBU4DnPanbglZGgAcwtlrqVds3c
MNRukaiZqlCB4PrUoZXs/3aD7hYtrapAgyRM3S8+Eyb0Ttf5XhB9ZiW9xqo8/wkDKMzlUBXdsSoD
lIdvOY58XrMZelGawQfX9dS13+zuIpPA6WFmcgpE5Jmerm1K3gdWLdKT1YLmQ/poom5+Q7TE13eU
XKZX7kNmDL3vaXp483eijUwTw8eKs8V1KrKd57aBDJjkh6seWhQIwj+za4dXsiMALjiYt3w4YyYC
PcpSaXCl0hljA1YNnRe4rwMIEL9M8o5tBtQkOOikOdjxWekp0iPHTSqNoHKKRxqJ7WRnF7BS2Tk8
1qe3nHsDAsUm+udTYRiin1ve9E5DKWinubG231PDQ8X2Z7J4Lx+4ePdkF8wS1El4NteYks4Ofwig
7+lcLsBL3Ni+5cly+Ku6V5yQLHwXN+TrQdvHMTknf+D+J4bH1zfjS7g/mfa7ClBoUOeTRxoMyIR7
GJqQW8w+C+6LEw19INDHF8rL828irt64P4xVMEkADOOP7xw954DDfBWfB7NUGV73KglAuY9vbTAa
LI/NgyBfzyS0l6TjshDVjx6HpgGnsMB6VzcqpZwbLW1INmIGaHJQH3C+H3wa2DRrhD3sYwHlpzK2
XZn/WQPiIP5L2RXSqyTmwAC3oHzgIZ30go0Ic/r68IpsxygP9M5kQM7Y9pAlaHFfzbmTJszPrfRr
eeSq4D+lmZA8tqWaH2LePwAWiY1HsqEx9oiR3rIJ1aIimf8oXifJ+cdLfy/jFC8eyYCgq/A5fGVQ
8Yyk3pdu8sll+QAAUwglxh1q6TeaoEatPqEp6SbTGPTQffPT1e/VDB7IevGcBgySqtn7x9MFAe36
Vf+lcxJqTgug9qgHGcS7bm06RR3Ufi0c+Ze+NCk/Dw+mJ42QbYpIgJkOC21bPcwBEwbiJvvx+BiY
1p7ZDbaf0Jlu4ybqbBlv6fwj5VTY8Xzt7RXnK7vRNDkF2V+MTdooRMErfl91T3jBwWfkgcf5i256
8ff5yQdNCERROQpUCKZnFfwUg4AI0ksDoWDJbBc1sfraci0cHv3aBibGTMlyIkQYFKM6Pkq8o2BP
A8wf8RdjSR10sS6GRJTxq2d8XPjfsPnMtxXjfdIs5+7gdYJgV2UgoKDgv1M6j6nwEVeIeFkIK3Dq
JTAMTaXiIFGM1s0DD37C7a6E+frA8H+R8K28SRugT18WwOmo8vNAw2Os1bVs50P+QNZ2FExtIRMc
jh6VQ4h280IidZQ9VVhNj5Nqlf7RJArQ4xvgHcpAMh/G4DO1hQwpZ+wm9EcMW4p82+jsBWzKQMbF
hChIsS4lu+6uFHgJkYkRjfFBU+Cnq61MS8qN/JObghotZ4W1fmmMRSo8PX89wffF9mmBKVv1eJfc
+Bqdkf17EBMA2Er6/q9dnytiqnCFy7gl60iUpkzzoFL/vEPaz1XxmPYFe7eSdeF5WA4HyAkPlNik
UDM3fr++HA2a7pCOh9BEAzYEOFCA7yT4PI0aJ5gxHihjnTq8H3RU4H3IrNmcm3jzyYot4XDGffyG
QIh1mrnO27KOSwYb5NFyIGs0CO9A8f4i52eIL5jw9UkHwJoZMFq+DD5bag4fK9wGjsKJw8HvrZbR
3WBCOceO6Ci5Ys3GllKa0DOBBQAYn1/pcY9Mi9g53uctjr6KD2CsVH+RbvL22MY0q3wYCfMc5b9E
K8b0NaO+LfaMYHozqwUy0zL7Bqss380t3MD5HiarUntM1SOd36RVGvG6HkgTUQSd7D5nL7zGCRqv
LXyp+45HDFN02yCHHOC402ImRNGCRrDBO7A7Q+7gJmyNHo3SDTgi5wdL3m5++pU6k8LAUH1dMnIj
FF4H74cd4RqwyJJ+0Om2wVR1swmJ5DKMnTIJd5juaLgPYhziofjPNyF6qZBBd1Mmjl5Md3V3Bvog
PBI+DjiBvJajNR+mN8C3NIW4lMcAmofxm9hzmcK8H+BDAKDsvqEC+cZ52ld9100vCYW7u0H9qCgS
ykVHTlxRikN4j0gYxH59e/LyBCDWerh8ohFg6RQkoHhuxhPzfiyk682wYnbvhR+m4Cn4N8TtZgVE
L7iCRqFtWVTa4zNZDW62UooaFnSxyiOoTdbGMjZMriadPrsXbR8pyqBoIISkuGBQrPVI61BLZEFf
4TInE1rYwNeGeIz3TWH7XTuI1w7HtlaF+Exd7qDw7JO8C1RDw1Zaonue5YcBzvEuRNu7K+4mudn3
SJmAMtzYnDArtCSD/fzYT9+3YLK1Nm3+sqf+8gp3qM+0gKTwn9ZobFgDDGfplgT2TgldZIpXu9ld
U/BVC2t7aXAS8qoLi80mGR7gt1+AbWC1lwUpVD+nvTbom9Pt+jpWyRQQDdjZw+bl7zB+9bSSVFvv
r9tvNEPsXV+TKyYFRz8piwGgYcJ+/jmFsKhhkRObJUnmIYrC4W8If3d7MOmEEXRNKz915Rz10bzN
kaP4PB0RNpTbRUsgABt3/CPQzQ8tYD6np7uFaWa80f0L3fLEekXPLR/AeS8wdXyOL1KlZ5dOrUBj
VdmJ947qGDFPC+twZbmtWyKsh84eY3F50z4zCLYofol/wQ4lzpCe8ZEkVKrg3UjFtYO+f17rR+un
OoTHhKur7ICwiqgJru0VgFqtjlhGheDUrsndjJNm5TR53epicm4IXCI7G86qqoSjNtEjlkpruda2
QpVGeOiY2gUhLWBa0k/24oG8C5GQZw2zXn+cNNyNogDhLXss+znmZan7gm1FGw4UlDDWngB8LaM9
ZSWwtnX09DGRLWiGrgv+4CWi6j5T6qkdWQgDQDbT2jdvIIFpqFSPayVopbv328TKmCpW7Iz6HKRY
7Tfb/u72jj9gJ0Lr0LITj06JywxUKND5ywYyLSFE+nuBGfEdzT2dYTkhjQ2ElGkUCmeFNRx7mekf
L7RvQ941AknCTQfAnz77asQQJ+2aS5Vre8CeQMKUIG2Z2gkASLXlWmVhp29ujjBhHbxnXH8byAMI
4+W+jeKG2eRNHf4MLq3CZbEVotafHIaeyjF0xlrKK+h3XQxsfqLW7AjF7oAKtPnhKCPcK+cVO/aQ
fURAioGrzUVnEqyVtz44+lKFyYBpg73JOvz/M2gNsnoaPmtVhBv3NzUqaBsoTUWyU6qsSpII0JAa
with4LWRd0rnAzik3h9aoJE6hNwalva7lD/RMj1Gl3flQga1jqRGqbHiNMQLTvRUqY5s1tFiO2iy
dUURk0+zbk1aqORgLMOw0sfEqaWSEvEhu46tlpHIwz4grm543JuRK3+yRL2mwpHW5tkqdSHJn6Yf
tAZD/gMh4ukFB/jG34eIQB8dCEd3TpnguTMMYSKE8CvTEJH87roM9DE+o2zLewznEr1uS3pRMmZ6
vhRxPEcWNXhFALO8xZeF9wUGt2hxRPxfDg0OVg982dsDpyS2YuC3bbvBxrdRat0MS5XP1MctHZeZ
mVA4aROR0KXWGEtG2DzYNpFLThZO20N2qu7Q2AGPkN89uC8AUzjrrXzEfmkCZwIGIr5YF5vsPmWZ
lXva9fF9nhvdwGmBxEshdiRU7nx0hQ/HxrHdhjF8/af0ApywP7dfbYCpp52/3uPatE/tFrlxzU8H
b87g7Fhsiq4p6cx+0VtOfgLtyvBRFtAIFeaOmCnSXXfj5qhTMVw5vGTlv0Ij+LMou5XXnz960MQm
VpFfCyCGpRm2YWoIPq76ZOCav+n5GtYZ5afleeyKrXcOe91qzN6J99tOGX4QwvK3s7e5ZxORDHrJ
Cx/m2bWWppacEA8xJWZwn6uQNhe6LBXJRSx3V8Eq4rAk4Go3gIzNxNH++Fhv3CEm0M8O64nenyp+
4noqyrBdn5BGT2yLYlTK1K9jRjETdvJTytZGpH8GrnIe/+5n3IEnVgWxI/EQXZhg5U9nip97N5Ks
yJfGf3PgW8JJwxan5hod1CPVbI3kuMyjhykUHiORxAPG2TbMCzwGaz7gCj9QhPistyud6VeVp9ur
jkuL+Q038Y01blgnKEUikBeRWHAIgcmXUsZq8oUat3SKYiMudiImHuDGFW+tuGIAJjgzX+pCCdwX
Klnm77IpS4iK0tbqqgTJeI8gWzUMioe+MjJlyyHkGiZ3k+3GofB7Ou8C3y0jcQm+raM/qc67B48H
V2V5OhRdJ1ELKibXzKC9OioKxSkJOylRl3b7CAeehi0MuQFmEhvqco3JJ1iX/HVkm4Qd6mtifgZn
VWtXx1vpN3kYkjfMT5UFQ4122KqZ5BSmCuy8Z76VDBhbTVShRn3IYNm2FeDfVOwleAtHsWqJBB2P
lWGJ2LotrYP2WT7Q2ZGCpDKX7eLeZijBel7gBCsM4HeyYor0FIXcWzbXf8aquTjQcCw1QymFbh0/
pX5jne99mH1K9gc8HuGfNOLIMzAn4R4lJXvS+cWrcpOLV0pRTLCWpbGrAZkJOoA2H9JJy3p39BBB
9dELOlckoJURIoqBo/jHcfUVbQyVJlbvO95VaX+tH85mzyBXXfEvVzCNv41Bl4K+Xwe2ssTTZqOF
SATSwYXx/FaTOG/PtYLEckgn5lwCsnvHvQyx+Owz+nX8ew1tl6ul7h1rGz5is+8HKtibpBuauBCP
zNb5ehVbE+M4i+qJWHqEetkBiKXFTJw/JNaXAN9xi/mv92iFt6daHOEcaXtEVvPLJChPdA5z+Pbh
833Ke06hyUTfWDQ4EtmpEGEtZH0vKJ5waWPjUCByzEORHlXKuJnOAs02CWHhd8CPY2gnPEe5JuDP
RaBW4zGj5Tc/kWhuX3jpDXkBAZFvLLFM5fQk6hfsNINqXRD7sfK4ZJPR8TSXl47GFn63oJRoJ5+e
v3W9N6FeUiIBe0tGpS76eI/PkKPKUwC7I7G6aN7nIQzU3yL+RaYXvuJVVqmaH8f0gaoRDgfj5kQK
KFMO0MMnGdowGqyuuWM5EVfSVYBrRv2D6NGoQixhaGZ7hPE4cPb6L1BFvGGD+rfjirRUscU4m46R
ux2kjj37XmmRXf44BJ45Cayd3xuErX9JT9HLadbRGRQcfOXHBOX5lCjgw8bOImniAOZCUyKe7Ayn
NrNXDScRg6ZC1zpfPJHGYiJx54MuYsKwlyP6Kiy3gQTuF7CH+MfSbz2U/lNwT9MoFeQpzVh3ahfW
w6ppA1IKqR12zP0rm6bFJq/gCcvip3wkkjiDmT8DcolEsu6N+vkO8IvyV+PR7vx5RXNsN9k8vJx9
lbZ+C3IfbWYcO1Rp2/Ddl7v0B/e3y3oPqUStZlPWeeuvc2k4RCgYufgvyQ98Av1bAzHR+XoRXLXo
sa/An2sOXhTHo7kgTwYJ1LbuZpfQIVVgc1R/AiDbmCHIVSXKB9NDsSZHFJTTkwC4JmsLUp7p8hCp
RRJLFddIKZJ8wwyGttXfYLLtI5b4dTcfzWj21qpgZGuw2wkaP28OZq66eUrVd7jFDrqXQk5pKK3O
923R+1mSht44YktcOMBub6B+/u4UNDG+mwg7Bd5qLHJZtFxnLJkvv5E6nHXksYGqIuy65u2YJfw5
Zu4j/n6pKYlU16grooN24hDMQrymDIXOS6HZDb8M6CanZCwdhBVGdoH1SKCb63G8Qi7Yw3MI8Wxl
pAohZigteHeVUn6qx8oerm++bexIi+CpOIHqIcRlvMA8mm46Wj5vUcSiU+vZ/hk5IWD20d45IyS1
UaakEymQd6Kb4fRB/wpmsDg5fC46T8P5gKLDqzcuZx6NV4S+hCvc/ttHZ89UkMD2f0aBMRr70/pK
ajcI+SIFmzpxenKFT30Y2JkUvSZHtn5jcdCaRkI4HEes5+ysI1aKKP0J1jvZk7Jk+SUEEr1wFUAF
YA7ZFFKwBM7MTwAUdE0dBB0REFbDMzCHqB/ORquA9ANLQMS6qnYl5+QXb2zT6AekXWMMWa8DWLxs
4UbcrB/DaQyIVzHzzSTx05qM6TMBH234waRBp/jSgDG2v5fjYc44jY1DppyCO/o/g1FrX3qjkzcL
Sul3uoqamtLs5vH8IndBr8bh1uNK7yTIY+63x0ww2qDTG3r8qTAJzpwXBWWKQXkCUFX80kafxIe5
EnXXvZljlx7lC2mYgEVzRUaKBckOtfBQSbf28y8tOiQXNoR/ZGD4jownNaOT824Kl6XEjMb5rIK7
U/3PtPqLP8ixSJyU1l+/pKsFqYxRvpnFGj06Zun5fbH3Zd/LlaEbiAplvEn9lZyG/XjVYR9s9yS7
58Vc+Qwj+LzLB3M2lTIs84QrZLqUNQyuEX5+/u7lYVjgIgvwYPFNrYybCXGAnUWidjgRkhWTBQSc
qTcFUMjEj1A+BQQmZuVeBuYBnx7RmcpVoryqX8IYSYjwtk1UThKPK/nielvw9TNKU8ujFZVsfwO7
kpfIvh3TxsWGZulhoPaLteXs9fbSXjPg9CaOT5jD9tK3C4+VaPwAjKKh1D1ZVJ1kKpPhdEtxL4J6
0puFnyKZB0nW7b6P7WRdkdJUmD38ZoDq8bpLLE4HOdsKg7y/pberZ763JORPeBHEWkAJyuWaxke+
iH8FJTAOyPCaFqwT2CiKs63xDh7c2MrMQ6Ohlc+ioTBjVaLKlKLD8RfgoPLf6uVhjdbhN12kS2o9
2eM+KvMtNrB0w2MT0WvlxDFn2FmfqEcnTJC/rwlTf7TVsTJy6mO6QHPeOYkj9Hy8GZM34yKyOWoF
T0QCIUNQ4qlLDRrtQI0LmDD2KTU1+O7vevcYkjF6+Lp7g/N1WUqqN9nGtB/ndR84bT9bMI/vZOsJ
+kAxnstmJ3+N7tnHrOFz/PiaGjiO/Sd3ooehumd57n0JeqfM9fusxOVh41+P6e0b9aGb1WzfuxXC
pEN1mPsnpOpiTeH5xhaIF+yr+ADCBbSiUCRoMf0DvCMySWRq3mpi3pkvl6ZwJBUc++ms/ROfoDEc
+a1wDsP/vwWOcEzciy3CRq6oPrbJ0Rda43kaK+HRr5/MlwqugzImafmw2b9oNdmwDXbC0UZC93Cd
rcxLzzanFQvdLAnZBfuByzjK+Jv5N44DVG8VXZ2MRu87ExrWvYMU9453aJO3WT1BeZcuUMo22rZb
nTNQ8Mes0yK40kzxYVFukTLNAi8XdAV+n4Q6z7LPNcKdsnhc53zx7+U6wLMG6xBgle7UfeKtKTz/
rq3OEU4B0BjCX2lNPYy6XBELj0o/NabXbp1RcCmBaQIW9I5QQRIWgXyt4/dyo06lBZbAYtMrEPpH
0olNPRByBzjSsA8EenydkSf0Ju5FfouGtNAedquiOEf8ekLFQgCra+fsP/h84M7fE3th1vZVHPDi
Vmi5lw3+3UKY4rCClHTuo25GZul7lLAy/4DkaY8vyxmlGwaFjMDnvd4oWrNn9Z5HPty+bwqNkp3a
ajjabFUXnDO93mlBNQWspBgITGIcE/tqF9oaYk/BxX1qrxt+EAVXAznXCCdfhQk+FoijLyu524L3
vRIyaE5hYw1CKkPWnUgMd1F7q76tZdfMYwMZfBLqBKTyrANhxmEbgCVMa3KW+Lp/rgjI8K8Xm9VY
zhVyb/FIl8nkt/KE6Sqz9msKVVmA7Lr2TKrgBqoaAeg53GbzoomVOQjyKScPiLBMmDc/RY63mvhZ
TkaDwG/kVa7FPEq7q55JQalV0HHbS50CbQL2Edz5a/owGTCHk9AImlMJsx0m1/5i+mP/ObahWXT3
rjWSoh9PHmMPlbL7P+0VCW7CWqFEkdHOeuW9wUT4B7TZJEQT59ACE/lXWd/hiDz8JlL6eNQ0jI0W
5J7dYlaPSxtRj7I1vNSBPT8IvJmBP3NrrFendwwCkClc2GOXd/aLlb3+3L8S2Wu1WUpOmlqrq4MA
j6LXHJS9tTh723rdUrCokd5lFTXq+KlnKb0Bnb6mgjeZuz7rDqebT13jTgPzAnXf/6TOLiCXUTn4
z3OMQuzjX+lsGKDo3VhkZuLOKBl7DeKb7QMm2ByTSzXHSDTvopKfrUg9TRZV7g504Zl0R9RozCQA
mQVD4UEQmYmR89xlkoS+4CjkcyJMl6ln8px5xtvE57IXSyNQeTBuwiOvXDik3jjFJ1S8tWWzIVqu
7vgO661090JByeJJ3tVfQUFOUZn8QxuSBF0Fcol9BJnyjYqvvlJhGlOsbZmrdEnR8hv0pzuloUaB
0nysFoh5AIwbAb6/MvYg5mUEWy5jfTXTNxQVv5zB0j2wwbpKgfLiUTGQ7m0vuUKerJ7jdNt37nZJ
n8AHcZaBtId8SKXTRXwYtoGwGH+cxtqryTDpFhbRCgsyYhADZJ42QK3NxzBULh6Z2vnnNSONP3X4
GsjbcdECa31kcE/88BcEOXQIGcwGRgdDP6X8Y5x06j2b+2Nqsx/Cn4jEXpNwxPsKxL3OmPTRjnS8
FXGTAdtGP4aNTCi4rrp9XFMELKCvYPUVsJwTEep6L1kAU8ZXtw/o7QOqX2ooLARYXCTk++/Dzc5B
W8M5BoarE7PaW6SGNoUWpNC8FZnKP+bddSog4dRZh+aoVIrR9G/6ii3CD3vOGZM0U2mm0k2oOisc
nxvGI84YRxUvN8XWh3zUpC5CKXn8DxLqDs2vMoL71W1ZVJVu7rbpx/j8A5mr+wGJcDZlKW1JWRsm
LieIeHGb/bxHOZeYwTBgont0Vn2Jm7kz3i7js35bFYbz+9wfUJjnn/YN3qbmNVouFfrf7PjEpQ3B
0PLjTwC7zhCnPXNrsrj8auOvHRdWCvRXSR0/+T9cxBqxrI3jQIVNfGUS78bGKhgrz3qUDZRbYzkF
bWgFHOYTn0vTiKu+wuMEkEur20eOMmcKm6YSkIdqVldGH3030VqAK5I3QxdTkKyquz9PzdmnVn3/
5osRfetsKa6MKdfa7YMZI2q2AAgKNmW9xDccQjQCdtqeAjBtWcT8Fm+glUgtw5dskqZizauKvOrr
pMSXCvMsZePXEKsws4LqcrRNYO1v3gcRJoSuZ6rhM86WMbwZTHch2vcqszfhQCcRzjRdhqRzybXl
s6Fpbk/Wnwf/10WsMe8W++OxLFVCIdO3ZALcQ201GYCfvIILZcRgX2Jvar4RR7/9wR+J9HMrysfY
4hCt/tFgZS69eHEVfKDjCGKUEoTFbNGLwB34rmtr1WrLHB02cWeMDrq9Yy5khHESBA1vPpthDsNq
4mDdT2zrKzcbw3VCgm8u4SjrxokNQsFZTVUJvhaC0GIxapTIgQq71zQ0958zDkcDmQJ3yTp7yMil
hC3ElQdgflmdRPkeSgNb1hhD4VPBK2O55PE65cVmW0uLV4LojXlHPRzvrDH1QwE6rA7t0BVawE7n
4TaxdrrE5w51sX32u5YA/4WWQliJezydKUbXnQwiv348wI189oIQXtyiUycUG2yfq9vbIwiwLdZU
bMOsQadg3E572CkddeYURf5t7h145BqK27PGcubRnE46srS5w2kdRL7XW1vh2qL2/0mi02NWKJ1R
B83vOCReVd8pvMgC8++DbnXz4eKsjcW1Ygm+R25CYIWoy7ebSmSnNP4rGJ52515zNbsZjWNMOW4+
dtqQpdc4s5v3wyOtt1JVpspoCZwgiXGeFQCRziAaia6Dg3k9kwa4wP0u9NY6tsN22AKv+MV/9bG3
neZi51cjmCvuvXU9+GIRcp5aDR1yL0W4zgkjoOEKCBRdNceG8v+cFKE6NAV5QqIq8O4Yh/n3lbkT
4PpCnWttXyce63ic19mACgcebfCZZi828etnh84CnhemCKIbOm9VD8UiCY8qpHRvL542VxLoFHg2
QicAaLgb7LDUjgz7RP8lgzqxGLvzzb+413yl41o5efXNJ++ETZND3F8dzVScnrletvLX7EoTt1Vl
S47MxWpL5eQf93oLNuG/ntkWX2jnzZFoo3hX421ce4XKWKx1Namo8K4+QzDFrTGXzJ+ssPZFjw0V
S2FZpjxZDeXOJtCa1Gay8ASJUkEnyKCh2a9oyKtYBiOrqwZ1+QtlPzzXwQdOY6gHZagNGUdNuRKT
gugJ+JIZRa0gXwjPhuf9vPMaLWHMXwh8K9euzLnxwFGtbEcBM1I+SKs8gR8krPfgc2dd7UTYJCIu
S1ozifsS0aDfqQeqvQ/N6QmOguBv/qCAdxYyUQ1JG0Nj2LU/ZbnhuJMaQn+d9Cp7kzc5jtbZkBAo
knzLRZvtsVJVS1YhuKfYUWNhi9NqtBxVW+FE2OPZNEmakxDcD4/vivgwRpVQPJPUxQlhT0R1SP5x
sEbmQG9ptK70vOF32o1B5eTEqCP0cre7JLVc50+lFvRWfE7ZyBmVrgz1xtZltmYp4EIIpXfNYHPv
8XHZl666QlSvZKhocxDTMhBByBSPlFKu9o4haEMo8DTPjw9QPgEkHLWYxgck9YFUM+e7Pv+hsy0S
5JN/0D5Wkpy+QWG1Uc2H+z8Jw9tHkdPGdxf3yh+tDGtflVYdBMVzHoZs7TPTOmkhAA7XvrB4kpz0
cxhHz6YQYCDAzWSCkN+X3PMoem9+JqLu2p/4b/wTcDxI/J9Ww02Ypd/AXH0bcxzNEIvzzIiY7Wub
hB978CMBYgAncNF8bePPQUY4dHyKjWoZ1szyJLbv2KDWetifmYroVZL5+HURdeDwAmEj315bZ+t8
l4cKFuDNXdynDewAQ4jCraOa8jBP5/WzDZ9bXzZnLuI81vv2FwEmfkMpEj/Tbp0QPlbDWuljxvR/
U9mBcynPFYddHCcyTCC2VIqmcSJ4rNWNqeDB21OedlA22IImzKtOCCZQ1sIk3tbHv+3bZ23nVNYO
nyaSzqHBw35WeGVFh95xZ6flXlz+mXMmoKmFQHpgDiVXTvZpXE487LhHhA3FPbX+w60oXH39ilas
HIJmQ3zheF2CKxGLYQ2fjNmZO0rjrPovY427jI3Y9Xj2js0e0YrJ7OOB7AxfJl1b+WC+a+dMA4k1
zmZ+L8E0cUJYlJubC+rv2Fa9p5x86jWyoplVktiOB9dm8J0LVjfUP9UfS28IaznM2eSrEd2GGQ6N
DUEEQJlEdy00R9Q0+vdph70WzjOhWVnL/3+ECtoZA40ZOAyKeLaRdmX+gE40FDadm2PwFGozZXWE
PgY8O31clL9mHjV17FhGSw5sVdPUJGXbxJjnPMYILgQErBK868+iBl1N/s/bHlQz99puavFONU4I
mRR3elrx4Mo5wKUEZyJc4znBq2UDFOu7QjvSFSEtxvMPaQBsH65hapIaE4pmTFqNPfMfdX8D/uO8
Wu/sKcDjDU0tdQL4IQT+3eSI0WVz6432bs7K3zBcG8C+k3Vl6qJD6Htxnxj69J2WrxmDuOmIhzBm
tARQskg0SZWGa4RPwvYQclZeYRqhGSQmb+hoP25Wbs8FLQgt+DZ296TQr9I/X+uLG/wFFK8x25In
tUvF3n1fTSa3wFIY0haT0JgQD6xCzwX1hpLI9LwKuz4ft/rPnECY0syxsp2P5dfAkciD3s4KZzHS
TDWTpjVtU8xdqriWZjO9MfwEZKcvmEhI478x4TvkqoItsG2bigg6RLVFAnDEbRJvX9/42sIG/U24
0XFwMrtZ+kK/v3cyFDSOQRhDFnrwN32DmebIf2HtTXNifYG1EIwC9H6hHadsE6lLmSyYYVTCk5N7
1Xnoe8bbfoZM2In2/Zw4/we348CBMRW0ZaKZi+SyIJ6OJk8BrA2N80GfCiRaM181TGxMuxV9dlsh
zJVDZCbeCsKkm3QR6OGTXdiVeUsIzBzHNkqf3FzdwAvck0DLYmFLi04zbebPvDdNU1MD97V2Csig
GW5sVGqJ3j9+RVjnuWLu9TJhjYUaccu4uzbzoeirCzzMqukCVfRGtl8RR009b/ABFJRHHOrORTNh
CId/ZcvAAmx3aaYI/ejdVPemzMjktxVQvLtZUzpgeTYQBRGHtZ5c0evOq1E4duT5Yj48ZDV/0y7C
oUfe2nHI4zDaB09S8lgPnqg4ZHtvGoiABDvIvSlJpNuKGUG/2ZmwhSnfNWhTzeRu+mxCFXpJMjr+
P91kOXXep35e21nU8bfXm6nFILuhhfmuHBH0sjL6wveyc7pxPJ7B4To03eezylouYHkqc/a/wQLQ
xt2Fx61JTUZ+nU56NrMSoVXpuwMwihv1RgplXd5p5dxNn9f26eZjdJNnTeDP8AFgYiI3cPCMAGKm
Xr/nj1t+m/T/w8c1+JbK2b2Dgek2uopA8qHoaTrJHMhaULPO/T3PFRH0zzAkhvEyfn9gE6cq99hx
esqAkuVuf1xktt3NNilTujaUcSZZlC35FIgJsgK/0aG0mAkWm7PHSb6HKxBNApX1HkLiEXQLBRLh
bC59tYNekzLaWAOCUTAYQ5hRHhVmTYoWuC1c+PFcIb2vD0gLx/THI+uk24XHxcezdZ049PWoeTHg
AN8+CPROlVOadcDH3LkIzjbSi1lzP9altoqpiw8xux3p2nBMz4gb/dA+GDofKg4h39AUEfOD8i/Z
fSseyUSMqdEOxsCm+thFOLp1QTI8Po/oCojJ3PZJbto74c+icy/Z80qj+I9x75YgT65MnavN2jRG
XbeDsrhPXhFyVv1/s0/ZzjGpbzF8q8HfsQYhW2i+XWRBf6F/W+CzO4pdIgEQyu8Y1zIYX7IBaIsl
ltRv+x9mGQA0bwNheUGz0nADAVscBVDU7W8zwJB1QfVH+yEEoX+yUYoG4hn5rbMw5lDWZcQFAu5+
a5HqAGzdowfbEZ5/W/zxYxKL05VVlGWYvhzCYs8M7Cj/m3EQIErLxUb/9DM+rPAHYdA00y8ZbPOJ
wdMBjmWKXEfGnLIS0UiAFnDIZBfyCvBWGL8juEziwo4/Ml0Rrfwo1Lyh5ZRUuUWMcwgx8lnrDONP
g4UGZsABHAsuIDsLuBjt9uLhBWI8JexHSROhFJ9zz8Xd+bDdADA7fGY3Z7gM0hLa4agO9usmareJ
HKNALx7uxaiMI1CbfYggDRrsAHhWDJ1JSIn2PeQmfUcrFEjr/vIkxTwH5K+ETLdnuujPSDAe7+ka
U3SUWwYawsR33wmUzuXvHthI99n9Rtve/Xf6niLt3MpqEBxhEGyp/5ZIikIS/IPwJk4TMU4hdRIn
HJg2Zmc07jmWhzoRvII5NIpkHhUEu73LGgmi924xCGmmNppJOcx/onTHewGQooNYpAwhhmSVuJda
NfB3dRGYJN1lElyvdvTOPMDASMYVI7RPrXzqtqKYoHEdNwx7D2twS/koVSzktJCTfAvqoZihMUd4
EGjcVSHidCYZiv32lSEZpWhJD5DT48fpIZtCbRCGrLIEWNKtG6a/0wccwJdgzEGGPDhpr45LQt7B
BHMdLE4iPiIUGiHXDFIU/y14JgDHyhnUh7Oxyj1T5zwe3h2AcpK27yAsZt/oSmxKQjXSecHWjZ+v
UgnsRleUNOr1K5t/vvQChPOBseSEhppw5fxzZ0LHlBRrh8406XrcYu3zNBjYH6mF4kjRaQUN7Ovo
Vf+JGafU5vA4osaHpwz87hHDKciy+t5waaCFHvPXmXn3xCCQg6qCcJ9WhmWWoNatwDh+sT6O0Q+Y
7SqAL7ESeVWXoFbt7ACRvPObR0eZAYKDPBXski4GUViyW9mZvlNtVYm7vzYziJZK9otdmV2mjF9a
/VHOF3tqFtsZvZhOU50uqNyjvCRpKOyra2CAnzUsmVoTcjRNTPTm4OHZnayAn5Z4E7mZFzKZjM3M
tyM6Rr8mXF2D322vkDBFMYRGIZ7m1KmRFvpYLXAz7l7m6Qeu0T+1ResmIw5xv4+vBuEhoHzsqbY1
uezK+Gr/ngddp7SPu/Mb+Rg+n/gHwjI7MAYxLKjZUgjmAFnSF7e5IwI0YAvqvGSLUp2dMtCLJes4
6TA/TzhY24Z8A7Vhvr9wLvZrb4T7ILvaZt6AmVm08Ue6zfkrs1WBgoUZqI8SlM3F/GP7jwBvxg5b
IsjwN3KPOcBPBvljWoVdCJiaoa4+qjFHuEK8PVrV6SfVczAvezNelqQ0VbMsytL8ZsYF4eVxJR78
3l7YEdPfbI+s9JqmEXtkl7bJod+LXfkKt8yVYGKodJZ6pK4jmySXXIA9zrAbmMVwiqcEKng1Inp9
HIxQSLZlZN/caX6BWZ9b8w1UdW1sa3glSGdBfIaquO2OsDrVoo7234A85Oq9b2YWgRma1qANNTkn
g9AgJnndnYXZTW0jjU4mAu4RA6w5nxbtOUrUXJkXuv7fTs8hCkJbKWKv8Y0O5nMfJyILr+4Ujquk
xey6ptDQ2ffqAqxM/lV+mbjKVA3WCs4MS1FJH1HU73u9vMnqO1XddNiJA1uWX21gsLdUOT3TMUYW
ugdayAfHtQk3g1h7bZ4YVnnWzXi90xQK/f63778Jlq51GcoxIl8ne6XPjeUkx64Ikglrn2wFd+6O
xGJ+TOCDQqIX6b78PS7H6eoKRhWEfk4rcm6RL+G+EhbQ02gRIl2hMPzPsRUDYqvfxx2ZPFiwoe6A
UnNEyfqKr32lTYCy44ZQWJYcwz9SNqXdnK1gbfjzX4H5QneqzG7YqnyDXrbDNKDe7DN6Lq7Nojob
MHw4DUcSFX88xni5yVQ3PMmd7lWnJbneO3VGXrKz6sVI2a4DZF6QLtI8NgXhyZcmsDw+mTgsiUW2
ZA3jRnXdbyd4bz1Q1iKYCuJ1SbgZJ92G6sg8Uo2CqBRgeX3ehNHw8DmbRaK+vRhLVZu8Dsh3ORip
gnw0DX/sO81PeNCgoEe31sGmsBiwgDfjaNAsrXEnCc4Oxc/AdvH4G32Fpe9p7AC8JQwRFof39Cnj
zX52i0yykD2aY2kZyMwbKo6r/NYm5u+cxCF13CHur/6YkXW+S6RIZry72/VA5A8DLhQ4xBGBWVkc
COGhEGACGStUBTg0U1rxmfcUrOBkPi8NdRoUTPkkGQV5zxPc1qP89W3W3wOTb1C4jQWPbytzIz7I
0gAMdtB/bdmrbVurPZzkIPZ0lXS5gVrQQtYRg/SiJTvk4AvB4pcqG7oEahJQT3LTXIgk0wTp1xQf
LIGuIgo/+KCs9sck/ODspbePd+Voio9Wj52qGdWHb7Dj1fz6NEI+lrrNBMug1W3HQaBzwvlNmIEI
gt5/ekPHDfMACl0xqLvpy5xc3RMH3JvbbqZvtOVUjt9Ec4D+UwRS2AxMh3jYgqujH9KbTuw512nF
AcyMDFdM/e5S6o8Bnfgo3cZTGMiCeR8bQAkgFDJi2RsYkNXc6eRyegqAZR82XyOKo1gh4KGP9oc6
bEAUKckKZFygmxGy8DYu5HUfY+d9lEtZnSXPGLM5f2a3ZCE+qBqxad1KQBxUNM6YY+4TEHLK2DOd
K1N0U0HEaHeZ7PqH8Gkegw2OXJZSeS8I1lNvEF9zxAK2RCJqJ5NlsWfKqgEK3Be8fS4UiNOwIKnn
uSk2F3C7S6+5WrEZACkM7nABTcXNvJBIaHJ5ky8gb+2mU69SRKsk9ScERtVVyUsZj0vIUa6CrMq4
/24qyMPglvWCeGqJktjoJ86U+S+2nlxdmxs9iYnvuNLF0PFtZNvjd/XhrSAUPD3kw5pyg0TnRxom
DJIM+72fAcbUvlixu4T35u9VPnHHlX97ulpR+5zGP/j4v2+LECiYdVaBtYqFqDMWytmI8/RBPfiF
8F3eYbgLG2hSpKf9XOk6t2OeYMMgj0zkOZfaXBnsVOcRQtoySQdOTRCLPQAY+AsdDHRDLQOgoRho
k0Ma7QBmkksCc4+6vEHERx1XE9yWQaQv3ItSR3fiPRgyKAqLCFoJhTo/X5zPGfxakt4XnG1lIHx1
GBdv8YcX1RgYtDgGnTb1TKqx/JFnsX4MPZoewTHkmdF+fGgowIvngkkcmggUJnHg9+pELD9w8j+d
Wvv7Fkjb3B7BgGFYC1w3i36KUO483tUsixOARJSPyCAqoFhIIpca0g5uq8+LbOiEV6eVts6lYU10
BwsrxFz2llQYHpgvxNv9xzsALzQjiXL6L5V2LxF2zCil9KEZ2pSdq7iVwWjencBUhzcCLEZDIWNa
y6nKj6WJAW8O12xtrVDt16YnpeEN9hlv7me4Ps3KEZuKUa69Hh56rAuCpV+kQwtTTGpGHSM583tC
sSHCfKAEa1zGBO2qgm675kX6DOINrXlZP/cV8GNj3BreIx9Q4Iv1fiGRIUMzy2YkZKgaCojVXi/B
wAhc4DjgspEMH9AtWmt2T8sioKc2LKcMohsbEkdz1h0mFckJtMVJaP57pzP2by+aunX1N6Mdi0l1
dun2yajeMjop7i+m/pLXvW66h6C9c5Ju5iWUcedd0Lqj1VuppZC+QKTE7mGRbgfCnRjXkUdbZK1Q
e1oQOXBeWIGCYU313rTQgYF2g49MkGGZIFAU0xwbg02ygrhUEE9fJlbVlFSu2O8+jYIsegQ3/u1O
JtfZiQKYUjwqG7ZcCEf7tQVS+dc5dag1mg7CxtbRew9OtpFrtvECh3g7Rnn26tJt09nipsfc+Ue7
GMBNI1ZULUjNghpYxoOlZ3UCdN6hJNwezmxp9bFqNwjIW7cs6bbYkmLC8nXxLVdxhU7rVVN83QFC
6dfGy6RJTugVrfZ/vcqAO/C6zxMWj8G26ZsoT8jpW2SP/VXV/jY6r1Xl/zWYk2idzB/hl7xZkJRZ
qmelNj1E/Y3wRoSiVZ+zLCaDVa6jLuA0VpLgeoR5M3rp8LwTykqwixRZZGbkfovQEKNyVqV5z+2J
8sEs4eVDHw3GLWZLGAEGFs5t3lbQNOfEt58AeAHvrlDEJU1xutqSGDqwIENS4bsqnxA3WmdYIWec
zONC6EUR+HMYaIQvoN3KWcMaSJDuwvo/TiyekscTLdU7xK48VJWgaOM6+ICyN3h+EMR9WmmpTn75
d/CTEp77psPzrQVmo3Z2DlzTaL7JfLnQZhMQd6P07aWmmzmdtehbMA8bwVF6wHvHz3g8im6FL4Ym
RAolbiHzlw1XbWIkRiUwouL1CYQqw4dT0sqeAnoyNNjkO3CZvr/38hFSgBzju9ogF7aoQR08/E6r
xMoODZ7bt2N19bCb71Q9YcHBtUNgoXZdiQpc9h8A9C7buCQ0JIuor8pYcgczb/J2W06RSswW5rXN
nAMdIZBQFezrvHe5jvp6w3Bp4vCNkGW2teV20fj+/nmYsZIbFuIGyh+MnA2pqdC2c5suz+o2l8LO
x21x7jWo4MDVSJyvgCdWbbsZT9v9/3t5i/lHdTGqC4kXt37J+coCjkhYoVUj/sjpRfLmif5ZLJQm
GRX4ia811MX3jZcjonovh6ozUuqIgC4iyVu0B0e4/t+Rpf4m5P1eNpA0ZK1eaprCuLlDuCdqIBzX
P26KFb+l/snuNz7tOfwSUiNpLvjScg7RCIkxSVs7wLG6ljefhaAKvPhC7hExqel0rLEUUl6LaIuV
4INTBda13qE36m6sDJthM+iMUy6yc7OPU96yE7l21QLo5Y+u6oYbOBfi0qfNuHR1M9cT1NiTroAK
33pg6AsPRKjcjr/ULJ6R/X+iNB5+5AJYHFZOmyVTBYgLvz0Mdn/fjd+sqXFdvnkF5CqsBiOdMFpb
FyrvJArCdiKWA5HIeUhRh0an5iMPKrVNsBXfETPHlrOALSzmAVdcyUBL5shUXKH+dsBUBE0SbNuE
ik0VoNOWDxWJJeifUKiwjQMG7ljgapJdzdNxYl2mlWx8RoPX4ZVed7Md420MaG8+1FUIX3B6SwFn
xaB3INP/clYQBSKPPYAe7rI3QDiZXuZGO94M31GBjauTaPEL4ZL+j9UPRUmuX+TwfKYsc+M7qjMr
yJv5hLEQNu6SSIa/zs0y0ebfMcmnSf9/e9Ea2JlDk1RTEvFQ+a+6sK9DJJyMUls65wqT88hq5bl+
3pD/JL1zcnDk/McL8Q+8vHojbDnAg0KQCGA7fpY9O7lEvYs72Sgs8P5ESofGESDZHWvAIuvDGFAS
c1Vlg6NgS3L8uMHxXMfQWQXnhdBrUhivsZA6ajvzGYRUTyQelvGZyvaSP3vl7pY4mp1rsx/3D73/
EoT82EiVLBlOyLPwJODqjf+Bb7QxAR1PITHkkLbSxXyLEGrvxpIe3BXOOqcDZFSph5o0bAp4swZ3
ht5FAdt5mEv0T2hscKYc3UUje5Q09lMqu9ohEAmPUdEBe/wrBmNwTqDncVyPMx081e5JuSwHFDfK
GVoq1lkQggAd8KPFHUV883S1/Ywcatpq9zR+VMLB4XbHzNrLpCbwq+SrrmHjFDmzquxs6ecrvsVK
HF8hy/QSRX14KTL4lg7UaOt3ZBHZW+jINtPGHfuIHfuMlj8Lzw2vURK8WcypBTgJgSWY1QeRzVHp
lfCZtZ7rb7Wo7X0ia2QzBQDpAxlgv3+RWu6U4dbzRCuQ25aizMiUHP7r1124td/rAanYaPpJy5Hm
cPpvRejjNNfhk4o0oS+pIRlxoVE2no147zRyjtXHziJH/QVlAmJgJPpuCqzoV8GM4uWdr2FYid0v
LRGFdqjuoIgD64VAOwlTpxWHwL/MdWruBYEk6nX2wdk5UhDW60+zF1aaVssgaablBhP2yQu2jhBp
P7b8FzGdqi2oG4VTu44T3i/VJeiXheEHGbxNqJ19sZlaLiw+yWyLLjOqL/v4UHg0pDlJdG0+u+Xx
pz+AuoUbruSkDU3yGeV8UfvH1P8DcvFAsrFxQ0BM0EofNp3nKB+/DvfVbG/6GbPId3e1YNppE2Lt
94l9wCHm0uH6nqn80XYutMcTJsOnlrJ3OawiikmR78feAYL6zC7PhNXajbBQgBx1f5kRG94X60x3
YQsTk88ZvCZoH/8rEcmVQTxpsqCP9sVAKCwFcGbfoQLN3WDqhHXSH+q1MJovBsO+ZVF7LE4KZUZw
x0CR2gCzB1iLjxXnxb11VVEBjXoWsAqclwlV9ckFJK9EGB5G9vo222ZGFqszOoEt5MJnc8ZouQx8
hdIQAdV7M0A3jjHIZGIzXxz2oJr1+oP4RbLamDQ8ghIRot8C9ii8g5kMYnaVbt++gkMXb5GI8r9b
PaGbsVxhqv8bLES9PFIHjRZDuIbFqBLaQopE66ZJylUU0/LJSwnaSv9JhZcmruUKGWNL+gHOv4wr
XfhwD7JZvmM3wHbmLX6Xxj3y0bNUTvqGiAHJjlXSpcp6QEGjuYNJlLIy9UuVoQuKa6VgAu4aI9ie
QeIjbj+6jE9KltAu2oCYfIOUsyK0YWbGPmWCCUi3e7tEbJpHxfI9q8uIdOpDNfTyE3tCdeNsQ+Ze
BZJ8j9gfdTOUFBPPeABaEpTw3Ue20Sxe6KGGGGoZHaPzAhYwwee9iFkT9o8LCuW4z5S0FoeG6q2M
dQovFBuNbwIrSrnQjCzC/HYqrGADoWJa+fAsxxk7+qg3P/U2qU0av9FDoCQdWh0LUt9hvxEANGWK
0QDQFgTdmWUjqflBGCp2UKQZ7OP3qNNlhoPJ5ZY9F4/Fi4ryoNNbte7TJEzqiOdGZTQmr3z6gSX/
xnTsu4VCKMyv3hEHVVbx3HoJdXDC9Kl95GBr6wGSv63kG5Z8G47JCO+tK9zHbKqbN0FkjN/OzfHD
BVr666ZpxSB3Cu6QYprEU5ZzD0938y/IPBBjN8uSBs4DVBEZTwtV79/a73KE3CmqFl7QZdUHIOsY
WSGN/C/zik2votf9QE9WtEGBRralPlZLIsdKbx7uN69loEqKl1B0wCfcl0KurVD8qxnH3VR5iOk7
B5tqmlAjQOQZiHCqymUQv5nnxfR9fR7kl6zOb2nXCFyR6AVeEGlx4nMgEEXZffpWf+g1kJWHc9sE
bIRxN8m6jto5qAGehovkE3TBb5h9sqAZdbbYt/T/Grn33VLRMEq2visJJjWm6ikglLeN0oS2j+f1
QctnXKQK8pQtFJH3uwvVq7PkLNeHIUmquvMutOggjCYH7VryAwTrRu/RJ41W41HQRbzZlGlvG2l+
F1D/UM1rIQW/x2RxiVzqc/225fZ4IdC6q38280dDSHuoI2CpU4tapwObTULzX07cjPEntd1FPfXP
j0QpILsB6PY0tI2kcUgY7RjUldzW3WI/Ucx7K4rsiTxrG2sWgu5SQhzERhX0bY+OHLCWJsvdp2WL
6As85gmnyBGLaim7vm9QGO9KxpM9LGSA8J0K77MvclxD+99KYCq0+h/T3IyXEwqqcU2s+YBrTp4n
RETMHvsHvWc2mItxSqQuFM+j6aR4RM8eMvz8eTvWgVbKw4Dr38sxDSlN8JWNZMFIVMwCjfq0/ech
PG9bmcmxiAQcnNS/TJlLxqK93OqAamIaaaoScHn28X8ts9NZksZ0G3jpqfdxr4J+I/zNDXgZkkHr
6z38KaoxU39NkIXL6EUmVmnkHAlcpwmfCHn+iKewhKH0dxL/6DyNMqcKDCpoWMtNfS81Qs7h0Ton
rdpDiSdKhaTypczVibLIXESOfGeBhsvbZUX4C5OGIpEPVKr9Sc4Bkhy/XXtbX5BiZYwAX++mKWWS
Dlv6BTQbII1NkXV1pXhUH4fHw/GDEvBt1fn77B4go02rLgt40JMESoCtVWTr/kJeY3iOPPocybfO
i8YZFbOmQAevPTTTg0i7XYsTxpJANm5P1Tgucv7S9zmm6C+NlD+Oyy5ZXiD0etxLF7Q/TAl3WCMp
7MoPRS1eURjO8fM4RN+2MTuSNiQqyEemWVPjPw2vbYZkzrzfcCd0JKsJtDvs5U4VVF2JaENvq5xU
ClcJgbn1QqWbelfuOEHNSnyybuFcknO16i4hNZxlq771PgB2sewgRLOh8Pbw00Pp7iRaU1F4eGtL
Sbt4I1nuJ4MEqmlZKvdlA/CQ1C+WHyxcP1b8CYR2twHDAGvlITFKJRS/r17lo6UGwMGZBDavjb69
6ZEGlpdoaLTJ9SuceV2n6Rz6/Y9tRHaUyOQkv5ROuBnOXpByftbXjaIQiCdj5Euv0bf2gfhWMRk0
h+/Pq9bJHqircdlT+ye8GBn0Z9OBQtl/W7EdKHMMCxybUed/NJsaJcEZXYiNXdrboI6vt3hP5rZE
P3jQD43f/6EZuOkJOeMX8AE1jQQD6qaYNuD5yAv01lIx92dpBsdGAjONJpVA1ewevcHsZQanGvYY
HedAhpNzIkGp4ptOhonqP4E5aaRh5Hl+/7sCvvDc516GFENZbrMvnSM6VjmDU/QtQSoyyR0D0vyt
AUFB+VXRnDPfQUzVeU5HtvExvOsESRBMo4iuesS+JLV6ubqsVjNS247xxtexeG/bDl4+bpoyjRii
Y96W2/pRVd1t9whjVedP3ad7ofK1VWRoHS51HtaiEEksrKp6wHEwY8e0hoQgHIQJ4grsG6pHD9pc
Wxkx7irZZIpqIu5u2YJLRWwCwXulz6ryY3GQXCdArvyDAGKJMBLpBQML/D7w6NxVZ7sdB+fRmxnq
yHIddNEQxqEPX1HZ2eX3Kotgsmx3fhjDEQw/W4BiSSqKCWhTubRVJcE6kzJpWRrh2JPawOliLXTt
T26cIV98GrLzVk9YShpiIgccQSyQPIZ5YtWj6a4GHdWDQyCjT0UpBlAwUeUPAMM/veGFMRN8ySrY
jOnniaGKt89YkrgrstK72CSCdnz4kxkF1z1hmi4YWI8unFi79D+yO4DgAcnleY26GsSZkPC+MwDB
nniLwkkszRAMb9Qs0qkXQuA6NBnX2IuvXMAEP6/4Z+muU6fZEuxT7LYh1TsawvaETCk12dIXkAHH
Gu4TbFnzkpLlXeb9HID3Z0TM9r9PzbuZIDKcCbjUChD/1LYyTXNB881dkcWa4OD3hE+vDpYL4/mF
sEahW31L32eFMt725aIrfFGbJ2LsSMKfOIX0x3Isy45ZTlURRlMS12CS1j9S6XPynJLb6yLE1hAj
sOofp7AYCl3rQmeYi4ESxmIyT1JP2ocN+s8qz4V5zXmibllmG14rdJgPw90ydBy57ePgoz88vZHU
ZD865kOeLI2YBrzg3JV3y8FnaUJ9RzE9QpIH/8Q8jA1yyYs+Y1UwE0OcDgYNwKWv59ve6zY/5vcr
yUandVZm+gREo9lur0Z5DW7fqwc69Ktxj5oJXfa2l49zADA5KiJpk+4BeSSLn0pLyjuvpUd69J++
W7kFheLGC8yGHHGQHhvCa38E5RkPi0pwZlqBm4bO+0x+EhcFll3FQsN9CwkAZT3KjvPPqK/i1x2i
CzL8y921X//aBVvAeha+ZODwXfn2InozFBjZwWViM+2goViWy4pEozJxtfJoAU9v8gu2ZjiFjqfo
9nzuyBGzMKvsPJguf0XR2H0YeLi8qcG6ArCeyVs6cB7Ak5VxvwOpTPwiHKBl1tmntxDCXmybe/4s
vuVudOOMbW1dDa5Ke5dAF+MA4xCmzvMP7GwvxMl14NOYLgA2t49PPxaYVAy68D3H0zkIPK0p9xhu
Wg5IAGV+0D+zeUr+PgHEHLXDNhKQAp/RIeb/AxTivGcFNUvWYgkTC6tlNY/xj56+YfMGUzj6CRi7
gdMEq0owtcnwVkBJvCJaPg3zo8MuLdTvHgJ2lp3txYfBSvFRkndCloAe1ge8H+Z9x7ui9GdTs7VU
GWvojsn9Irr/hLBCE1TycfVnBdVSNVJobT7q1mEXiq5xI8/36FpsakGd1TaUeV9bTiQbUA5NyniW
SxqmYtxDXplIqtRIJH2z8SNHV+b14MJxrbeweYw4moBU7TdGPOaZS5Mo50GRcRvTMZYj5RufStH6
r3F5KPdaTIBZ1onIacobe8rbRyww3epGg10srJm/KtTTNyY7wPHrJCafQkmWrCeugxxFVACtKDsz
nmbKxpnRyIlJ1T34vBn/SrWGWnZkgXw3K6UqkF+2ogJFK9W53alw8xNb02sXRtySZrk820O676qP
qJ2IUVUqnDbmhT1hn3eq0lZb74z1OZf6m4cTQ8cpzhomspSz6VQnGdaAG3BNvl9LyvIQA+HRVsgl
yh1Qz447tUlNixRvtxXMOmLKYUYvMRfEA9BtBy3pZqE2yHS3ekWUiQvVVFzw6j7S0qI5YgycuQ8Q
kF3++nvjipYhZGpdpG4hUTkUOm1E5MYEdGdKTDGdldZFFtFu9mJQp8F1Mr4pg7V+9Cx0mRebyNNP
uSMiK8DtwvOsWX/I40rubMlMzbMzD9bGmxS88yBg9n1XYgnTHEZOM9u+MEzaqcye9vJmikk9WPpQ
4npb1NQjC6VyPIsvwK6oG9txGW8fc94DrueJgcJQbgMjB2I/vLTyfHcEaTayV+wuO804HxpK5Glu
ETKESHrJv1OK+XpxFeTPkT6HIDC5PPjjBGAjmKCJiCFHMmv18BPQaMAaF+h8gKGYRDlN0xl+Wpse
TKlksxfAujAig4+SaeAB+/uw60t1+R9FdrEQCRiKFCo0S1lg5lFBTEc5PaVjMZ1kuODqJ+Dvw1MM
AuDlN6yv2jVUlicJiwsLnSvLlp0Vz//sjgIcbplUmpjfIrAIOFugbvKFna25Fp/3d9GT+5O6zmVA
YN991htEFL9ebLamxhzxdTprRKasTYEiwT5GBrsU5/ZG7AGMAn+UHDIn66sOzoA/Ll5Rj1pZayY1
h9wKv/wcuyUALTJ9NXsRBSooe8B2f9ngZPqHKI14mX5RHda784mVwwDhYWOvwlRHkTkegfNBAt62
MTDmil4ybrkLMWFUGgvOL9N9dndXtT82Im/YVZdP7USsc5fdCOFr1PDvQTIE2xj6bv/VSzufI+Wj
z0Www/Q+j5rbqht1M7OuCpSJgm4fNZ/4Zdg9V5Dce9BDtUQ7Sfbxl7FRDz2FE6HHNfS/3aImLKa6
D4pe4L6RJ54d1o/5aY2gP/HxZE4LNelq9dVF8C2jR/tK2ZoLxPnLOTKUtiJrDvherUhqvDJa8SR7
pIG4XBnha4hGRY8MnDhcvy1jGjbbCHX+nplzxyFxqBHVtYaKoROtfJ5V3SFU6E0lqbu8MRXKTC0Z
JciDMgILgIKdHwI6K0yhdgxuByNmnO7/N8yt2DzouCRr7VMX9Z5YB3Og8FJbV6lqq6vZ6LvaVSQr
QXdqQmeJkzpGer6YgIHQ7EikhkP15DTflrXZUeQKZauZ0AqwjJsHNUWvtCg54ZSC3x9Jlcjh5kHj
mzhGWjmPJKw7/vDuzyt7Im215XCrI+HrvrTvE4XcwSD718crYmUgMNiAClTw9KhkZLCYFEM34o1U
j2FI0FHYvVLml0conjQ/cHZRWOSxpUkFzDB3ZCPG7zSBzRpV1182qPwfYo+qLXwww0YOGOr1ebYn
KTHGCvV+R4U8fzzUrQtQ/qlgisWBzuET02pMDqNCr6FwB5J71iwNvVFUDugU5EwYO1oMJBwssYxt
Y0wrhTfuHBTEzPtz1Gcm/c6KBc1JobSl+dV6YeAl9OnX6iUd4oM78obFAQci3XwGYa728Ro6dTsK
xmZvoD915TxNwk7ZGfVU8B5jfFIybvI9ZNa1Ws4TOtxEPIzZz6XvdUg67clq8wj50oDJjC4GB0jT
77MWlc5VCb6uq/6enGHLR400jtsEUiAxZTd4j+tt1bXmnnVlrFgSrAdViypvcXo4AUOMh3rF6s7E
Eca0prsBjqbXwe0ox6qCTViG/KlSUN9aG2Srw5tmSPVmdgEh73zgVNFRYMS6/DvOjR8HYsK65tcR
ZRJF/LLWNdjKtAbtnELvZmPtNXATCgjAxRgIWamXLZX0aE72+axiPuxIRZWa7TfoLQWff8oFlTVB
xByOlUz8ny+kug5+c4kGO9P/aUpdWVdzRd0D6Q6GppYoXKgGp/oa2wlj9r3yhEC6EXiYEqGuX0Aq
wB95f/IfpQ54Ja2ta+K8BMG1YhymJd2hTEyR/sjzbGF7C8OmhQRKgizsJtIzIOgt0jfWyDzgs05I
kFrXbG6UTgqEYEWH3sXWncMEzQRvqQQxiCmLbP0s7g7eCQa0CDEat/dL5sKMWzg21d4VfnPO6t16
MWtenpk9PilIVqt5aUsqw9a9YCwhMHMvEF6/Q7qb+WREF7NOQbXfFI5iEZKu+hkpp773/vL1FXrE
GJDcpZ2P1ToIZ/MdCoMfh1/tw5tvgV563XTBFCjyo9vXnAnthYBirDT4kSCxApn38YY/XmSVLLJA
F7thOX7ngCXl/Id1DAxHuVwb966//khF3LUsHZR42WAqDIXwpjVtuaw8XyTBxttLHS4OpRJXVcZd
0ZdF7t9l0qTvcw7DhFaf4SRU9bOx1fr6JAPfcjt5wbkf4UKovVZE5UxTNmihnUF8ALK3wY1lSgGf
CSQq/UG/BlmRZGrCtG2cvAIZFlYmtnt+As+6PSRZDOTbDfqxmN7jj2JjRcpDSu0k+klEB4Dc1xZh
jJ639ruFDZiNxaoj2YLqi6RebDQaZ/tnFGTSM0l12TogZIW+DvHbM76POXMzj1mNApkzwibTKFG2
LXHnQ1/OGZ5raoqkDcWp0OtD5KwaACHjBOup57mNwuMCVyt7CyDLarnNIG8XRjeDnjUX0vbT20en
pjZqOnl1U4F3JBqovppPy9kvzYKUx+O4xxmKHR/jVmvZcepDy75uojvyQgTrEFFse6gjB8N156gQ
AX+LAvtZWRZbr6a8zOwRlbVG3E81XjqoAMYgc2tuSkI6hZ8kmZ3C8jIn5om8EBXL1AS6DompSKx2
m6dFhbbYiaob41NsjFd38dyf1BzURkqWGqFSUaczTYpfYFCQDF52MERh1kFqBrT7C2w4fjezcnNg
B+rMOCjoUk26QHtuR9CFuXj+Nkpzxn0Gqq4HUC/oJMbYIaz2TgPT2pfalXV5GHOImtECEw0ihLxp
wxAJOkWxQ6ivoFDMKJvBdcCIgo9rDvTsFPUs6Ef2nvMD2oM4qJTkgGylzISq1MyK1N+FErr7/k+k
hjJmFO70inJb8DPPG3VHR6dJM/9teIxuWb7/0ijh+s8YuKYSZH4Vc3J7TMDrGmd3pXhfwy+nV4Z7
al31exK/yUVCf5239eperGbT/1tcRC0XDz3Eyih0wO7B7CJPKL7Ek4ERjigr6T/naEVUtd0Hl1hD
6/+JKxmjnfsuwHiXu7G7v7saZgpixwLdWuE1bJmLH+/4X15/XJGpemrvgktOorXCXBbA4/AWte4i
Pnk8mToceH5fL8bVXxk7iXMcP49qS3o6pO/+DaQrYIpHjPyKU597N1yD18Rwb0wpT3+l8AmAP1uR
3coFxplkni0ynl4BRYLTLyp64MBaOxneUjZq7gKh6qK14a9TU6UiJJOsADEZ2Z7+p1zNI7l8gbxK
gCJW2PYd6iUNNJFpcUyksW1RhTge1nMWOlVeIe3NBEDDLHcpbeSdMChDNhrxi911X4L46+Jx7rQ1
sxRVj/DsCRl1vqJFFg6VPwzkW+f97qNk1u8sbA/879nC6z/q/PJ89f0D/VjYFzdBVoA38wJ0nIiM
05Hu00zHmzGtSWBnn4NsZsT5n23OlaSN1NjqrJ+pOiY/MITEYEKU1yShfXs7jbCt7Uj92Q1TmcXG
Ay+M9QSWfkgF5Dfc5befEBn4z3voXEaDVmR2fVGvkw1kblSv6otKfbwqFMpETR8G9zIBxXFeXdHi
R4jCBYBW9cTHd/BzSiQRTiN5xzE+w5XwaJNWlpY2oPfgnTxDLu4ZrkDX0gUQewOmlxMNonOrTQVi
XViZHW3R7K17/COWOLSo+MhOMcohU57nBYsmnKDslQu/ZWKf0FzkC4uDTz0uS+qVu4VtgTmsHGFO
KiFxu+ba6IhwtQ8Dq/Kzczoe+uHAlVLesK8PIzDr/TVVGZw76LJbP4WmexsBVht7O7izZ+u0zSAs
Lu4ObToMaXiaZUaoETYzEbSgtaGRiDa+gbjQtIfYwuFACo/61CwW6cww1TIOpdcvgS6j32cJsprG
qcerA4jzsFmjYKi5uHF+1HkhjrF0v6cfc6xc5Q7xGkkIzj/2b7Rjn+pUmM1hiXRJ6+vm0Imb9SBc
qRyCp8FR39bhMhXXCQ2j9yiAyOdF4yru3Vl/RtcPzOkIdSt3ipDMEoofhpSo07y/aqwklI2KVifO
824Zw9HW7i8Lq6+kDzKd2cKL51bcPKZCWb+5A8fCq/Hkbgsl6JmohRXl5RqnZ2/nLgGEgboMoDgg
gb+/7zy7tAMqPnoFKOr/+Nn7zeicWsUfIa12JkGHdWcW/ZacVDmtWJMINCBp8SQnhQUDM60knrJX
loqhyZRIJxpo6uM7RfxH+L5X8HAQWZYuATo7dF0qFOA1yUxuCAyQ0YKFIZPmAHSV6frYqFaVC6hE
fvRaWVzB3hgz4auHo2J4B56CqBffF1VwOJ5Ljeu2VWO6xoXjM80e1wVB3vSQLU+xgANrXAinMyBn
s+b64Z/Tn5ZPUNCHCN4s5m08pLHd5zm54zyHBs9mXP2TgGGVcMaww8v+fgLYis1Z5A7pIHJhedFK
aqzYdq1Rq2uRo+D8ma1Q6TeYrONhbtVFhu52Ur5MG5q0V10rtsMkTZ3+Iqitt2g/bq8g7HVQt8t6
x44nX/kwaEHe06+jpVvzkFvAgf/vWlkeZ1OTo0MpKvF4IxXhh89olFujMuahPKU5HqWvDt1CLBHc
U+iNLgkwHvQPhbzAiiXg/hs7UYV2XxMJXM2RvtByOthpR+tg9rIiLzkAkFUGP7Q5GY3WzDVv/i+B
kWZkqspwOYaIAolliswz/HsBNuTJX3xrGjJdrFRcnV+ltTsoG+bC/yO1cxojYYzw03/R8RuLk+Zo
mnViJRpNvxke8uFz1dd/RPpIbTXelaf0eGmkwZph+z2ZpPKnWQZQzoaEE8yZGqHbS1+GvsQ1xIcT
7o04nwju/N7fvAUr0XuK83q2WecOJijYdzWxnZ1FapVhCLB7iOZuhu+w+j4WNZ9+xBLa/OvjdQst
ed5nn9sbgRZQCceMF1P8l8Y5mESo1nhUFHdd3EzAIT5Yse9/8d6HbvKMF9dYnhB688krlTxT5VQE
V/X5BeXibKJzfxI+Wa7b6LsYIv4lttxjgPqUXmQYlaxlXFwacuMALa6MYvbomIxTAYHLBNc9t4I5
HZBiHNKDPHxlD7zFsrAY5lIvwuwRePRmXXAcdZpnpCQCQqKlTdvjikN5EdPKGlIby/iDUVN7wi5X
Et7cGxGQLZ6z5fbcw95d+sa4vbdWoPa26BS/tuUsGSS1La1w56rwjQDg1Z98tMKlIhJSoNEM01yL
RTVtVlDRDhfYDA5V9rozqIir5XMOKUF+q3S0A90I3l4gWOeEZ4XKADc/Y5HY63+i984PqVT80DAN
DObfBGn63U6BcjoJm83Pcv80vqoEpYQQGTRZkD8w5JYWkMQRyRT39DxoYpwBxE5EAMbsPMK9sypP
s7B1VL8O5IWV7cWyN/P7mEA76QItrxHG/d3EQuOXyQkngDHl8SoTH/RfA4PLGc3QdKd3CldGTUCl
A32KPrmDMkwwdofbCJMa4AtpALfvjhob5+rgneSpRjfIp8mGZrB0XxssCfE92yJ0vZqrAqLjQ2NS
tnWQ38/yOz2PioU8zBHy3+wsiX2B31l2rrSBdcXvv+KX0s+fvh8euyHoIZX56unSq60cfOnjukj4
1cLA4M7pLrlkkSNw3LGD/15d7k3aj+4o/WAgUNh1Anu2HQbt8zzNu8/sSqw919mf8y9KiuhsJJWZ
vhWavtSWr/BOhIxmOsQ9e3r9ICXNCvp80b1+VHGvF6nqVHf2i92nUhp8VcIJ2Onvw+oIFhp5XtBU
AaLc8bHMAm+xK0pfxV+2PBelEVvQkwhWuKZHkFsLQl4ig9qnmSSUP/BCUnQ+/a4a+Q3ph0XE/lrD
SUBWffhrgLJRHKEiXAmQ+Sdm54gh24UeZryD8EELXldmmkDMUv0GDF8TnaJbSfNOhkdZftywgPY0
J8nE275Lrk09jjC685uj+YHwpOwrrtR3VY4IJE5L3LvjBVu+pq26m1CnE4MegvFIKzsUFImgtnTn
SjTcilKtwXJuUtmTfLD5MEaRJpz1ZR88vOBnFSyqxIekH/ZDbTu+4IgnA+jgSIkfbCBBYX24J0OE
a0yl7metIx+IglowsqaSEKc3YC3TMa5eITbvnFhBJMwREjd771FftfF6vki26oR4gBW0FvAvYS1t
leyBhAkjtLJ6RATt7cdDn6jm/POTUC3ZIyoQStbaPDss8bH1fkb1LbfvZv/QTELtyeuBgp5m86U4
CHxZ6MmESFvhbOAO2JA7Goiy+v39ttkXkM4rogvJztl22hsH0AsZROk1E3oMGjrzH2yqrNShwSYs
Eg1oHF8QPwA0ZrEn+q1PPiVg4tvyaC8/FQ+LowxmZVfGHp0EOIB9K6Xq+MHRCK9MIte230FyG2hA
nhvcEAB2jcvPkCf3NnlQMAT1qlfZlQ68B+IchmYU+Eq/F5H8K3/jR/yLPEpmm914H3MtLAngxxvB
8FndXmXv3SQq1hEH9HO7UBfggcj0wuv6QgFg5Hw8RZpvwDbUKJAVoVe9UgPDFBeFnYUet1Ovncl1
upixvCl/2UAWsRhGHt9Hp4edYs6vHA3SzLTy4bAo8iCCj00c3DpBbfNzmZJQ4H6QfJmr20/XbNjE
FsDFGccPWzDCRr+2rUo5ArCFOVlmrSqFnY7MTIZXZxXI0htxEJhXajjEPzbxiyszajX/Ay7+zPUw
lt2lqg6P67lvJy5QoztoV3mBb/9OhHh4VqeGyutB4RMxDcPQ0sDYKVnks4M406N+rsCgpFJ0X3WB
/7CXC8wE3uJ9npWDlYEIaYs0K+XBV40AySM64jMmAFZ1VUEQX/8Egp2MLN562CiPv0JM3kzYIZp+
KG/yhLAWtN1uqf13ZKHqF+TkMJw/7To1X81YDDY6Vvw+F7metHdh0wNfSQrJUlzt73MyEak+cTfq
p37pm/aDXMkaL/2ytfD9sDnh0gLaJlI7C1MW0L9ZXNFtgCYiJGCm6JxT55UCmPycio6yhy7FND80
KQqx3xRhwwuemsyPiyecsrGD1Zt9F8ccwcJrft+dJFxe93fSN5i07+FksKLf52lY3Qk3Tp9/LIDD
HoKyMSRQ/nY3zNg7cbG1Y6Vqnp3nduNuKkTLp5Gyx7wGG6oxX+HQYt8c2AhTF/T7MfcNviBKJbNv
QMRE36yFGHiVRvkOxuFsFcmQiWhJUlAZBBuKNQgo0g2McVTh0aQQ6xCXNuziUamVPDbWjRhkMm9x
B0++nd2esG4NFSmWr3wAQvID2eCQ74Grys5DF9k6uWmxR18244eeVP0R8pV1pYXnM8PbOpna3rBH
qjvJXLN63UYIk6OIjCbqfr02HzFlXrmanTFLw32Csk9FNL5d9BBn0vaIbvONnISRqIn5G5IE9mWn
QmwMM8MxQV3oYc+JWf8PJaIFcoNpIi0ua8M6DRerYVTMrwhQc7vlRnsdmrDFSkkGkDlTfDo93AAq
/2+6AZalX3P8xglP70G9qcFS6pw+TjwJ8ABLDqvVn/yQlZkNt1S/be2VQ3GLCQ+lQ+EBWcaBL43s
ByLLsrk5sFdCZZNpDrXPWvtHWAALjTxeOTy0RCfGIEaWFQHG+tShCGJXaDtk+k8vLZDEBmIwsrbu
8SoN2oXaOBYEEAxU2nRxaf0R9ttr+v6T3jiUDyR6JjyQ7tHis1G1q6uUIA31F70APVLvdVxGaMLE
C/5jjOlKXJMXfg/9JmLaL+LSkN8IkiJ29CWb7f5ObPjpIu488GlHsXSA/TeTZDDLqiut14VLVI/g
g49UGcm5rxW4Z7FEOxqz7arj+YX0EO8PGyNaBLnaltAXa8sDkzCBg6FKTeELwngUKweMvqDN0udi
ADMLx/zIaIwPBQmA04LvWkYXhXK0hXIBopuD1z4f+tUL8OUUR9LlwX4mn9QDJkYbTWkcSLi0eo56
xs5LaEBGbmi7tMCscn9mLe4XaRd7+sB7F9CNLspnvobz+WpBPUh8NMsQQPlzULCzKGxpi2+IDiHw
bfTj8CEHuynPL+5Rkwey+vCZeePGpMbz/Lo/ZSYMDzs9IId/sKN7obEZERr2rISSGjrQHP2fqOTj
9dQs2AeoQan+zGN1//mgj3YLOgbVHzr/9p+CkWr+Aa7JHWenodCEeuD8hA1pozFIf+qs2Wq9uEVS
cJjS3olVV79N9jsks+Xj0yKp/vBpGAY2/rrcnZXfIEI+hoCG1uDgrM0LM5bOBRj4LQ+lTRM8Chzg
640Fr8969V7UtBeuNrGPYtyT/VdUBseWruWkwEsx3HjXoVuLOeJBUzfpIkgJ5b8woo+Zjs4tONsz
OfcODdnacSd7h5dKC706Ga4iOcabWg9ZiRqQB1aNSNaPj/8535DHRS8FKdNp0mscgR2pz7HoaUAr
nmIRfXt3IghsY8+qZs9eK2oPkE5NqR62G3H/yWO8Rb9Sx9NprjxdoLXUs9Rt+8XwgPqbHBO9tYUP
Me0SP5A5iO3JU2RLVp0CBDr6+L9u/lC3hbT0f9TepQ9cIzmu4EF+MufHePWVOhFrOjjO24/lwRjZ
sLUUBmSLqymxMcJYWv8VMScH63jTuEE0uOLYq2fYu6U02X90pTe4Dvu/lEdly7WMtjyCVJ/ounmf
KP/M6JWhfCwqVd7pY3lpPyl/awkeAjcqSMhLakLdspdW/UGqZXSW95PhbHt8Ta2Mm6dO848esCCA
FpxfTUEQkHLJBHNTiYpHQtMXsWlOSPVlhD7sc9PuCnT313LgWW8cZIvZGpp5hFoNqmpollElmkFz
BhlC3YsUznNeEgkOTWrwczv4ExY6G11RNn+vpo6NC8pDQzx1LGeQ0Jk2kPItyPCgodhuzdK20x/S
xhymh+nrMdhE7JmyHKo07PawsZnK/L7o82HOhtZuOyjKQc0DYi1HgTVY8JSI+kMH2CRpjXA4mLMW
4IsbwZzy3feT+MPgMf1ny6+MIcUDB6uREfo0f07yEE+6grLqhm4kYnc/tdesRy2K2YgJ4caWmePL
i4rYpBTHWgmdG6wGhQESVjB5urB0LnWHsC2D0XpFT8NroWvVbF4YWGbK05WNhANqyl924C19rap9
XbYCDqlQ6d8mWsNQ2haUN5eVP6oczHUCiZEJN6zSSPWPvT2swy8KpOsz4xgfChkzeF7FCGEwLQ7e
U99TA38LcrQx63eVBI8zKoZke3y8KKfOeMX4DoX5zJWfNBbhy9KGhhG8S0QYA1Mz3lChBWAGBBev
xjPxwfzdDfJfo4iLHfpmEbncd7MCkrd0zW5ojv5mzYDEbd9RhvDkJkHLDSq8Q2hJhjTFouqME/VP
ed0ne5O4fn3pfc6Yy0Q1x2k1sj156MhoQ1qIc5KaDsaLDrZzKqbFxuj9pLnQ05x8amZsnzAbt63X
E9jR/kAGeaURwOp7PKvpeAFj/2fDVIuKZ0Drk4UIDWgvrx6iRZa6zLMLPP/jw6rusaUU26zuRw/4
VH3j7hzJJRfO3UmM3G71DpnPB/bcpKQyRBv0INAg9VJiDph3O567C7UXVS1C4uif3Di/aJNqobRB
ehtCF/hJLElHA+7TowQM4IeH2RPg7YnLmVYeBQCpZpPbqOuVXLjubrP4wG/Ff6xBuiK84wMEyAul
/AO6pmJ+rH3WzO5P5MrbvQfCugan+7DugNp2oXqY59W9n6zc4ydK3WLm8les/o2c+p9e9bIkt+Ni
MvZNUNMzRI2ZPbxqlEG8n+e02xHp+u+/BakJ70KgifEs2hqZtv/XrK9FIQ7npsZ0tMcFe31ploCS
sdfjkdx1LK4n5dmWSeDMzc7jELCpRolhaKEIqCtwCb9uxoHlWg01WlF5kq5mF5E8DdwOYWbuoXlM
pF03/PNWvIf3BFXgFiXr2dTg8OcQHdsz9i/TMStWDgmIsw6BTK/WY+11NDmWH9Nm8Yoq59OCIP6c
uG6b1us9GEktuODS8dZ6q2SmOzA+zMHLgmslObfJ+gBshkF0vc8wWxzt1EXr9VPTT0ojmfNkt+zr
Tv2Oco7e1bHcGN0eTiTZfPi6/XdaCrjp3QI1rVTfW3GvLZVFQeIn9C5x13CsvwgVehHdpyB8S81U
BdfssvFY4dqQ14RDp3maU72QSOMvh0bHLHteyQvCBIytdf6aR9ujycyWNpTNqWffblMTqUOjJUlX
k0RwZUWP6NQq83JLl4W/pxA6/xBcKJAMnoPaGhjS4GHFtIh2ns4ZNx3b8x/U5OzgGwTwZunJJom5
YL+w3CVeAbwwOFBDrhZflHcmbITpGhCfCBs89tWg9pByXKWuGrhBhIHV1XCCSzo0jThOc9ZpUH1e
qNSPdjT9pd+zdNxmfOLiewFZ5X15LCDUMggNsaId/+gNCcvos0pYMRsAXYoYSqAd0eSyD1ijdlEu
mHObDfxminjlLe7nDpBewC0D0BpSvzjqvPYFH4blkUn9xS8naEBAgHXrRVDZd2aukNiCszyrCOhb
ukGSsigeRivpSZKlX2qbWD6kGotkFHx0dV+E9rYEEaVDtvSPAn7qkDmylXD2AtK8/dkz7AOpPBSy
gHohc85HAv+FtQ6RfXZlaEW3yjZsg5pevIN2t/vkK02kAwT0Vhsx52Zakj/ApEM6I1NUNUIFr/uv
pehWHyFB2VLLLU+WX5V9uX5sS0a+wdGVAvAi8XCTsqDe6UHFPLRVy0Euyce1Drw9f9KFkW5jetmC
LnkxB7OyQ7orzWE9o1m/Gl4fYRCTkYOCQipq3QyP7ZfCRMF6uxlhEhS9zWKU/m/OUjN0XlBiL3QB
UsGDgCBVCRtiNksx7y5heM/KfKphrFJVp6/ezhZJ1+Rg2y5fyhvdRpdonss78tP3uVdu1eRI/72Z
+I/ki/aAG/doTbhwg3fP3GuKPFBActKLAimjqd3yV+L0CxZwHYyvgbHEroPEdWd35jgzQyeDxn4s
bK3TbL8sLvEZkAKjn9vasadT8hIJ9/zKo2Ui8RYGoS0uR8G8/mYFK1dErfG0RGzWjDVeqW1XpKGm
iY3BF3OzAOqNDHVt0qgawBvzTrCoCqBERILOcG//QtbN6g66I6JBy26Q+qeAktAn2jjk8yZSyeMm
mmgbbGoTecRFZnRxj7AfiRs9n6Loy0+lHjuQL/4YVtB2Uxc3fShEw7/dQXpRD2aOjWFka71H/I3p
F9ytPFg+TAYSvFbg7pGt7vg+aFyvpc4zG69tTPAI0ZTdf1XQ6d1GyBBBxzI4ebDDJuQLE6IJOGvJ
1taPD8rT6UwygnZeg2Yv4mdM54KyWINkjv2UveIrEfJZXtEFD+oV+cmBi2UjdqGZXTsoercqF739
pb0rqpsoWlFaHQy4SoxnvDQt6VYYCPdO8uCU/6YKLPfkUjNxnnSL6IQxu0heaPn5hVGSWAL2gMG2
vpGbYZBArnDpiL5To141mqEYUSNbVUW9ibKXqH8wlTRd8zoe1uV31HiVqbVl6yjxHMyE5j/wJhiq
K2CPVidcQqNipU44TFrpKQGiMLHKyo9d7LwgtFCV3/tv8fz/ND6GtfK71DRSI15vBHDQWwL/iX5Z
Eyxl3GSbRql7PAe9nRauoxEtWi/jVHIwW5MV6E3XaaXtfqMfDJGbv1E5fzsiGVRgFKVH1ubaKBxm
r37UQLepnNAU7p8v6+ucFn+lREsoua6iWmU0VoEis/zPHdb46d70XOpm+39q5xKNtcOzPVPAim2z
CcMBA+qd9mHanm89pjkFmgJeSmjMmov/FplQRIujUTPcPvHdjoPad9jcOb7AElY5lHQfK+s3GEVT
hjDrKSNlQ4+IfBaDwW1H+YwmtPVdyJzlwCSCG6axcX30ZmRDIlcS7Nt/m0BBcOtGvn3/Zdmdni4X
31vh1kXwQEeeCjUQ/f97+dbauZHyqnQAidzAxn10AuusI0cExFgh93vUHSSn/Hdu9jqSnH7BaHtm
NJd7CMv4ooGBPy5X3Ce96Zi74zqP7oOi+O0eHvXbsb9/Em2ogqRPrRtox/d1GLjDQXIiU99f9sKG
SVlxqodg4JalTyZiD7/KxwTwe8LCV6Hn9JfixjRedUAe7s97+hIrSfuqAqQfExrM1CGTEBX2fvZj
cjwPyF8NAhg1kgm1I2aeQrIGl1u0Kf3gGOyvM2mrVPNc5Ta4a+D+jbg5WkPIQgk3OW+RmPV+uKco
6j3ZsoYAbwnfRthSV333TwwBglnXSpt7VCcj6K/dKXAdxuDMpehNUhEuIexP0EeJ/odHHMOfeMOD
XGKWj7tcO7Ca1oViaA5MFs5WWlJOaYAB9w7Hf4l9jHOnOmJtoc0hjywcPzpEeU/myGm06kk+8eyj
gz7binE2uim9Iv5B9HC8mBKnC65S/ITkf4Naf2ylADWW9S4Vv2CgPSfTx+Fhcme4BtMEhbss1rIx
chzzkjpvcHBQRVEhQ3xD5wGFQdaP7ur44gQxmjWVk8WFfQneuaAbrH04jHjIK60tPhZRXY83qqI0
Wxe7FPh/5eFgTFloBe1HR7cbyG5XX3wjxJNSsHs4Fv06G/cUIb8pWBJ9YPPoD0dXMvnoGWA42mtg
I4ihudP0OBOhPDg044rfcX5HTmdCWIoS3uMYJDmWOgPjdwhb2PMWWPv9jfJ/fg+xxJR3YqDQW1ed
M6Uk/wA8hWbQCzeIhDxXJ+IHB2WXS+cxeyjjoTKoP1g5yDLTHi1IRc/g804VVXZm4SeMzP5VVzKQ
/eYCYajiXv+6hOQWfdXR4mgbt0u0/oTQrgqluFU7bNfv8+4eM0Q4npDqoZ/TImiRTx6j+ZkXZmA6
+eblzOuAFZ+Z71sbsmaS2EGY2JQnotpNZAL3sHz3Mlv9HjUsQPjXkShGNkEovYvbwD5rr6YKAVh6
zVlwh9MU7qAuz4Lb0+QKdE672396tp/sKMgZgXg5KXx40JlHYEkloH7FNAQYiL2cQ4bRPBR8P2/+
cNbnq3i/vwvD01V4UOAjNUPpV16hqPlYo66gXHZivWDoOiUXYqup2BogMQJxu+gPuz2wuDFAGpFR
V61l7aCqpTI+WKCbIHJmQdRdWgDAgSJtTateVLQAXERUpahU5b2UkyZxvFz8D5HrheiAUoN9nJVV
5S/woFTyBB3+JWRwuqr7TxaalffjW7C6aITzLBF0OSfUN6rgMewW/nTsCZZbgwKEm9E4C2TyRuhS
43UqBsT286Gw/BObj1/siF/zo754CHRGtLJvIIhOOHWqMysa631Y4WYM8UjbEpJkykD6iMVk1eVZ
PeZjB9WQhI9xxywXnLG5mHBrz9UpFfQf8m07OX2IVxCJnzsQ/bcbKtSLfC/UHqE7Mc1pLnGFvZRD
FIe0b8pOgzKNgiD+wNG6tmR15LjHSS6/N3FMzoW5OX2JZm392q2jAf3++/xq+qOi8KAY1tTy0+JC
S3PBMEv9f+XiInwIF5mpyYOVUG9RcAae4RNrxl/X7BGvNWyLi8xQsfYrmUEnr9JNHi7KB1cdFEtO
vjHdQzwOwZN27azLY+fBEO6Mm0wv6QKIm3gvDP6eawm2JzkcI82Wy7m2pCBV5Y2d/o2BTJYNyjUv
Yu715go86FXWO9U+w/4pgFyAD1BYf+E6M3EwiFUkMvr/2jLuWIJWvZDQ9kVz9RjZ0DiTbWbz2xni
JH/l8mFpYF4yzqz7xJATcbBrXoFfF7j8AraLapmVAhy1SmveAQuKA0vAa7MMY9C/YEgHgPYUCJ8w
2zqgta7ztwwLuf77oHHfxMg8r4cyILPNaoH6DlShH1Kd1zI41jVkgXlz/2O5C0kykq6TNRYuqjMP
vSuCMh5Zfgjy6k8DdV+9dHe3xmQi78eBjrdDmG7O5ORDeep3HSOYTIohcQ4vx+jwBFjRhJMCVT1h
OgENb545pyqWHtFa5QXHVxnClzdxazg0dXHcMXQE6JIeXyJzWUudBJg1/mS85aA7lHeowGeIfbmO
B2UCt40LFKdaicijYWhy1KVG1i91MMlMeQA0lSY1/a3Ztjr5MsLR2aUdoEmMTOPRgHFzcjhpjUB/
KREJp4jfIBH1kJvjU2rwjkAvM8sNBza6AWAk0I33TzqUV3qUWZ4txYlYm0ccUWbNQiQrbq4xzIt/
6tdxHmXqEjmQlsRS7b/Wq6rE+hzUn/JIq40THN7El/btaNsMJ4R0vG5irXMFpf7fd0tArKi+snjv
nZsdDH79N2KIcQ7HP2K2vxcF19+4mIUSsgfuBo1m8vjzPcIx2cWGS9G6x4rdpg8JTZuxtcNuzsy4
Z4JY7Hyoa3FxqpETfg5BWMnqMGMuMLgpPXAOsbVJQjCqr6lil/Z8munwr+JAFq4np4Lrqrj9me+R
CVuterdBAv440pLVdG1/E/6UXehVR7byiTYCZTAgC7DcWlrKvh3eCitP113zae7NwvAvYuwRYp11
vVLwYW9v+vuZTPdfF9AGeUZFXKdbDAVBcteb2rKj2FMwz4adQ4JbcAPytt3lWXR5Kk6cE0ECTqZj
w3QJ7mKE8T0mCNr+uTx5kQnjXqGrGX+mTKJCLL5khU7T29iAuys04zCpG36ysAJF8seqhH7Kk4f0
hgBuc9LHaclnFzn7GXiR1y9WBPNA/ZvyAEgHSxRRQMaiuCoiCgYYX5Aj4X3j+KFAbHr1izDfbQ9c
AakgY/Eo5tRzCYsaEVJ0aFc3KIVSVrE7iJinuIPybd33g7xGAeWkNaT65ZPiYoyT5UD9y3W0s1KM
tkih1a6AzDt204WD318Bgc8KkcjISmCthP/mJjpDiogJ+9pR1lMmt0pPneu44U+8va7eGCvrZH1Z
zFcvolyaq+XF0rliRb995nm/J9yZqJ418XHXoUMrSvR2ULjLibX7rE+oGgmfmfNXQxgZQvxWJtE2
p7/t6uLN6B6OjMtOyft/ZZG3DIhzf4Q2RWZT+OpnEULkvHhxEpUYm0N+5oMXlW3ERtq7CIsY0Sfx
QGrkWuxmDEN9he1K/O2RFnl1pNqTNGSNoMIMkJQBoTKDDEvRSgTv74SgNOqmfzb0Qksj4Yf+A7Gl
fYXDtZUpbkp5liPTOaCYY9mGlWDUyutiLnz4fIHVUdOVWyF5o9FuN+rMSJJ6wrah3ip9NALiJQkT
s1ygCJe3h/FPm5uvEdnm0Db1RtO9hSvx7YL/0Bf9Mti8qqDiG+TdMA1x3QGnZBaFtLII+x1Qmvdq
6oJiVH5BTTKhRhrwSoIJnj8i+x8N/NUX/F/0icD6UroEp6U8Cgzyscn7JaEboEuN+oFXedN1E42j
KqttOzItc5J7b+f1svhA/KXzAIX47BYrqS27JJdsfs1v1qtQYgU/9N/01eGJM5bBueqt9DO+fis4
yshpRNPSXLjI04II4Uy+VvrSYZggZArqqSj8RT1Wcy9CiDxjHsouNJ6HNx7P8mTvtO1an8INMIwd
EBQzSXmeLxjm0de8aBMnxKYUoVwdlu3KEWW9YqABWZ7PAPllDQHb9SRGBg/xdhMtvboXrrHjP0rS
x0vWE4zXVtuDXLf6NISoulrepoK+nDt3W89FOdCzTor8GGbyz8nKp/gzwFD1d08i4wRpKReGUtMX
fw2FfVJY2oOfUzIfUpN3IwkXFrwisJycKdlp6U7ROOXHA7zzhh7S62RsTLoV9yTUTRTWaDDnkiZg
gjEN3tQ1ublEsCzfzG/ZUu/j1J8/CdWBkuvoah12Qk/mE4cNUn6HR/vjU5j98YmRGP7Vg/+7RR5z
xlXtPKqJajlaF9OHRHp6Lr7tSuXOXDi0WcFfSz7uyaDGg8dullb2rdN1Re+1fwvnud7IHBocHZEM
LfUarMiSs+xnjIDuEcV+FCwM3CTlVQcgqTGIakywQTwaTxO4ldfHcmgEucaVFJ/B99uJFmPzum5j
kQkZ9ZEguOuJFkc50MoWjM3D9Y7yBOhR5YFliJXwaIV760gzBJlAu0V6l670MHdyeyLB7yut439Q
jZXjXX7RzoKbu/QXkaOBtMXYl44+UeDWTTL5vcmXD2pHPe+rmhg/OxqxXzvar04YHPO9Vww2MGKB
MQlP91Gyz+T6hD7cednqXe59RfOD5xyY/jMtPmNwxdT1wwE/a5GFZSFZSuxkHnSZcB0fzyAee8RW
54mpGwazPkpjrB/7RN0x+jWXL+Inx+oQy2Olxy3ML54bPXcRobaJ1FjGpiXWwMsUZR25LXKMOHke
c1vrL9AcE0PuADb70HLf2ryjn3/kcLpBUqQ1jMaPQNdvKwxBmASqP2Bva0RrO1Dt2RvTfwEf//Hp
JeAaXdTks2zGgeAyvZz7fSSqkFmFB7+ax83fkuKZsHfy9+U2xRl/XtCKJyOjkfj9lDX2B9bp/jIX
whncKOpmJTrkILeGSpDNzOKqNQbQrwqVFlzdYodb9CQBrDkua/NaNjeLQlyh1Rx+9I70fGE9uO/u
PyoAN5cxDxYqfxa8e/Nf8GyhHkrJAiV06KeJvZzqIc3fzU5I7k4+f0eyy0Avp0R4ljXh3Ci9sd05
KZ30S1TeMg1Z7RtqB1wiUuMrwCr1rcou3B3v1XTMP3bTqfERFEId/J59czdQzmhxkR8kHyuwm/Wq
kaBxQIwUthnAt9xZJRj4A509YHi4gcqfLxWSKpjE9AtN3Tex2b2qfaCzWxQG3eKGy1Cp50os2Ecc
PKStFHbyLSvEaFx7+06S+l39f+U555iJXjDjTfowf0WnCPeJcyIGcjf9uSZeUaaHolF7Qo0b3svv
/53n3OFaSqbHB2GyMuDQaW2wmSNbHU4dKd/b7xPWMkcwquJg5l6U24fau1FprBMKcLpfCIrklfMW
hvIJc8C/4tXNXWml4YEaK73WJB/tGU9iHR9zfZDzwrJRI7ViviGvicJYa7x4ug64aG3bMQ9AD9Xi
FdeaU24mveu7KGm7wu9ytJSABoci63ycb1i68B+2lCf28xxwfDZmOeb5wdyZd3DzdIhgml3cFfgb
Py2j+xF260g8Ap+TzVwUHEpETOMaYr7itMKycHewZEa7TdXcLEfEBFYkqpEmrYIuCVPxBvhduOZl
mhWdXOyNgxwScuZ8hLiBb+wDEcvHsuXDUkSv9rhNSSfvU6KZR4wo/ef/6J3ptELgzopVOGT/ri6I
dFPPfpsIuiLgfGeAhTU8QF6BlFS0WoFFviDDxp40SwNhU8dwKPl9FpihDx2t6rmmCtfruv7CxtkH
Tk8Ye7H2e4frWkGPigJlCweBMIHkrK5xLLvZ3Z7krvsKQgeUlqzjrhOYqIZZO2hWFyVoCPZ96kjJ
JhEsrPpo0MQtndo/pq6pB8PLYOfTWJRMAGoMpEfodvPLu6IiKIqfJefyeqo7gkQZEzKsurDjAnVm
X/TYWmhqEFqXPa32eFhC70HtkuDpagMXnic30m0eEL2nuBHz+yyQMntWOyWFHEMaStps33l4hayx
1zoup5QWXG5mHYLE1kkK5bq2MYanEoSkHg8LLwoPkjg2PDYbxar2pF6nsJwwkmh80+ffHHHBQ5DG
PhMHr7ilfK3reEBxwSLhcALCNpKrCtyLFX2w7ouHHTBUTzZ0ywCQEIGoh/d15vNIXKGwDUYGj7LF
A16zCH4Cv8SqJojF/Q6Gtd0rEg7ccRccSvgF8SeudunJSL+xOlwS+SR5TLjQBQ30fATwm3ASRxP4
+iggxfXNH0n+ckvlo9kWserBkiEVv9DYWDlRY1ioC4TRTPW14ciFu7Y8LFbJ2OYtZX/6F3GD5HmE
FLUeweyZ+bub2I3H0PerfpeE6Gp5WH1UshyVpCsNk+HDUSFihGm6PejUG0G2LeWPU5O8UhYrrPHs
AdFt0RVrHuWh/TAtc12FzRDmfS+FQL5bNwSryWLP9l1/qLOxtGwdGvZMjxdtbJqbZwJHU5VaYIuN
fosPcgncmrVxocs8RTGI9UZUHrdCpivse4er7L6IffHfGnhaI0hFz/RCsl7f7g5oMd+PZR0gYJQH
yvDRAXpZRrl89FljHAdLXYHH+JOfzmDrvLheyYU5jnEbpzFXT5tp81xHbsE7WkCVu8/SODZtzoy1
pCUv4II6gBt8xMRq2f2mVYUdBBBd836Izgif/lVBceQNmSWUMh3pPG4W3LnkBvOvDcM7HGjfGDQn
rq7SFJ1QE6WmNsgSN1FtwwYLbEqOHWI8jp3U/ZjjU729+xhk7eF+fFSGQbNckHLVkkpHUUg1G6ao
yCVDBYCEQlt69HrlCsWsbEcs5TCSyMmiZClpXLrV/83DMmjIRkFj4A7V/0eNupCrSSklWGmdHv1E
Y3PLHKfhyBoPfl8wyoqVZV4m25CLIcr08HXrfLRe69TIDed6tARKIO6B6YeezAEEvnNxIDNxp/Wo
mFiCO/1X7H1/XAz8P74uEuYBD5ClW4h9t++D6KliGrWmVMo/TQHHqgrE88zF8WSn7DJOAFlR0jmf
Miq5uk+Yhu5fSBK1ORs4xfvmPMkOy/6ExJ3DLv1b2B7MpIVdlOdbrgjUGlK1YfTN73HbbAiZUQRG
ucisHxyA0aTCJ4BzqQdtltE53b9y56m4UPzr5IfenF2COzkt5iMn7xCiwglDS04KpHGe4g7sFKs8
x091bCCzECMGjZNfY1n53HjTNPPhChHn4QA2HEYkDUgTaHYjgvMCgLOGM/GjfaoF584aGQp3c+Vy
ByurXRoYTB2TWZOa67ahhaEscweDl0RcI+kVuKdXeEYoaNcUvr3FSMysfrddt4fHY1GE9R9Vw6v/
YPz1iMzGzKduyxSt+w/Yhpl7Ax4uvzB3yx5aiqKO9F9OB4J5TncVk8urhrHz4FGiJod8ZpmiMll6
RcKPPBnRRWgNNP2fzfYXrwfyCEbd2oEMC2XRllS0zIDRdAG9iak1JgqeoehXpTUhL1WtZQpxNnjg
+vVehETCjxAYEdcTymoj+76NRbX7HWPOAA5ZI2S226zXvk5TVwsXZXl4aXGCngyIh4fXD6huCHD9
taI47tMpG0iyK9cb1QRt9Ew3ZR9Pjn+0IfsbPGkJecmhSrcHvThg7DRIMoLa410GAO+7SVdHLXcF
gn4sgHGv0+PRNHiKATNMSQ2Z6hBD1vs2LRWoPpb4/VLgq9fFh7PITrevVIuKCrro8evmnHsudNU+
4pRy0Wyx+SQ0rNiCmzBt1uNRjm8yHu+GWY66GhrpI1Jm8O8QxOZtHJP/Lal9A0gTlwv+Iw8Siaf7
VlHGPUMZl0Tyja1tS7xf9TcTi7koGC5nfzjAbEBmYcHH9JqDpMYCdUgsjAyhdoDCFa075pGjHJ0U
nDzGLecPPKKdkWljaecACfpxTVCuPkVjW7FUXaSCyAOTFf/PIsNNZGNsfChJzHSBHRSwJxXeMCgg
BAE8M0tJJMW2vQGnWYAd+GBfG3qP68pOY8mPkgG2AAiC5CnjrYBELRLhMn4Y578lqJEIAzAfWsVr
PHAvrXbFRVz8S9uz49RYiHQYNdaYxaDE/BO8/+srJpO7Tj4O5pr1CYViWPup23Jo2Q52kOREYtgF
JjRkMembBhLGrxy5rktt/TCQcXRs84ygCI54oG47xDm4ZgdloNWTDZDeAp4QxMAkXrl2g5mEvPHB
JTzoIoKavfL4U05XYvv+yI9qQ1R+9Fwk99gpHQTJqeifnOevNjmucTi1QN7fb+l1L0Ck2BJj5LZN
Ut7djN1Kw9XA4enum0WDBwdIHGBstN8h+wTUXSUcZFCIUGH/rmCBkzJWF/Q2di2ytCxT7L5Mp9fO
j8UHCNflBeyG9zR4fUx/FJJSjUuYDFyBwAmwcPffnkDLSKgyk8BRppP2AeN6MjsrLQu41HfV0wq4
mHbiRIkiG7HNVgDttTBQzjGAba50IYD/Sygh45EJL0v5WJYap4w1J9oNkb6L1gT+ob1OXLWT7uLu
5oYmE58eErHKEjjO8dOHAaVp5z7q53ayitXjET5rBRAzIA48ZdUPe+fGLdWFRadxsd4jR95xXkgi
LKruK4tDaOsQ8zPnc/G7/AeoOyGzlCE2mjPccoef2B7raW1o5LZzNnH3jK3ZYRvFWDZ7vM3YY0fk
yU2rIp0SQpr6+uK6as1sPfa5UNXAbDXJcjLi3zjD0t400XpNnzuDv5IxEJ1a3hlZp35/SraM8Dvh
iWMAn5o6bF5rbK/R/2TogimBAL78fzgTwk4nh8D9zKOBRDhWXhJgOFlDntagUZ/EKEcky135nC0W
+c5HEgRXCr4YBy9+n5zh72R2039Xm/tER87w7o9bhPUJwNcaOCf2YXrwvVDMeVyFhowmpIJfuDQP
k9ycnkwD0dIsIUYk6h4aMYg0+vuUp8GZOEzxOlOf/nQcfd+I4fQp0A8LedocOK4/TYp60Wnxi06+
mubV5cLgkMK2zuRrAUqgpaV9Ac9LTmSV+5L2ShIU4hgY2CJUjqLV5AcqmmKMonLoC3HjmrKS9YYM
Y6p8bnFUymqaYSjWzgNLoAg6z4TmAPhT1osSitK+4HGFhuCzsXJVsi7/+aCOgouxCeuEYsFuSHmO
z33WcfRKZAmDY986Qf+riRj0DV+9QHUorgrJhLX8cvdZnC1w+6Ktl7hchlFIxYnD2XIP6+CYwAKY
Dc8bOnevVU8WaUm3quzsLWzlwKn50DeMbWNfRM+aBRK3ctxALkr5fDqsUjXaV736Z7svYq+6N9W4
pUZn3g+FR3lcVpxv6PaC0qkA+L/83vxb2gB5gq4iKuRibi6J+vecd6948XRJczeP8alvr4OIgigO
wzPhlOcveUGlpZryBh+F1GLJ3IVEo4gjcoii6JSjbRHVqycWQtBVI6APnG7YZfuEFVfJVtkThrA0
QHi0m/jEV3HG8T9tY3ho425FnFiJixxJbySt9+cx+73sRQBBCIMEulkvPdDcV5b6U81C5WBefIVd
5mE/C9B07gemEjGVXFywiG2JZQ0SsAwZpIPnebclJ8jPugbxkzQIhnME0/X2HYe7Z81OLXMjE4V5
TIpOvvWI52l6kWrEDzk0VPJn02Ibrec1eiuNPXl6PP1nSYzd922zF4hcPYgZ7jb6sQdkkSUKHepm
Vx7FqF5kGImyR//gRlmgG1DP1/jiAAXtmToNkuWDJ3EjdDtJ8T0Y7z0FFXTiWvbAzAPV5dpMZeZz
QMi+qsTM9QQFkaY7J9VUq9PhIP9kDCl+yqk7erSCwoCekjA6WpXJ4552k/9I5MOfKI2/+59X6pTT
WBAIUDowhO6SicRwNuJ/L9lXN6hvsMRKcmytxWeBqWJ/xCgzesbjxgS/sDgVBXZ78ibIkxjSYmjF
aBOFqJYOLjRZcAJxDXCeNBAdUTDtoovQQucBcCaqLF/kMjCrzjhRK3eEkZdVIxhcYxAUH7VKGSej
WfubDLPHinY8x852ZAnIpL11UevsrFl6V9b4+m8Zs0M/LOPeQxHUX4SiCU/UgMpxQ1CjSwMm1t1M
IY9i0mmrdW1H8oP0DQVBbG7qWf4kU9I4Zu/E0a5iX4Gfn7en5vDmepUrnbpnbyBVLTzrJuadsTc8
Wqi1csjVicOUpPkMMUzq82jjG1GrR5b134daqJQTgf2KqaWZvwyQ98vCPbcQ+ra2Id98c9HnwLgc
35EeHRmzBCglEifM2vfiVXruMmAyQZ+YOnew27gKrDjZ46gpaTtYp55pwG4IthZDcnqk4CBdYqM8
jO4/wdcoTMr85em0WWiom94qPByzk5i5ga+O6pFrmDfwl3qhbPQ8oAu+Oww58VQi2/h2FDyhYWBX
llXem+80ddrMQThGZUK2mzuTQDGOEMzR8Vt3xLMWWbyXQvr5/wlJlmKJhgYDQXWYCk3U2Wfww11b
0iXzOU0Iu5DMedLPqffOcCxN+DM+JYM5u8vZtEYlct0/jCW6Gt/T1DhobuAStg9oSTfwtA56itG5
FSMz5xDvxthiZxCv71QSy5LZ7lfW5xJdliFbr5yQi5Bq+A+P7L4YHVpFWgaewFHEW2FN+O8HCg9n
6Xqd12VtLf5nY15q7Cqh7H2PT+RtSfZxPPvC4+GT+Ib79eMrSBkNTvOjbDz6co4pjvj2iT4R9gHn
w03zHJppVTRB09/q+eIojhaPqauempJStxNh56gDGMBl7Fh7SzaeiEuWppIs+07VykPIv83pmBV0
qBdrXuEXMh5MmVWz92cz6PtWb9i/eAj/U1un67e3YJrd+dF3c8pbzEXBqD6319BbmM1ng/dkBNRR
7o0UWwL4JGtmz5eyeGJAkt0w+GGcZhN0eCwEJ4jzmtD7q725ashfQ8DCQSilYSWvvzWGv1cIr20B
XsEt6kmth9trTdy3FXWXM3azT8st6Xo5p87ikZGL2XPRZcTLkPuV9qqFUTeQ8P7iTeL20cM6va9H
tZjFHegiADVAtbjJOdy3kNNeDMlTVwySzzpLOd7Q1hZg9ArWlOFkLzEH93g/MysqyE3FpWnlZJ5Y
xW2tNrBtPO2npRCG8HFvpR76zKUYa0ievi7UJQojWQAsmjxsU87Log3FSQKgr64LSL7KnAj5vyRq
4/SuOm4N6VpW+mFBn4C8HUgfo7C9wVPud0QfFjgtFX3PH2IH9lC430S6ck1QTtBtoZgtP98yzBFG
rj/euTiP072P6v6NN9d9WRgC8IFYdqm0GrvObKY3oe1mAyWA6tg1hEUFeEdbl5uf4jkmOaM0Z54z
gUp8jIuEhxHUPcEaZx7q0Gdrg2YnCIZVsWV3foXC5i3PNKkGacuH8IUgZazydt8kaS1N+bACwifZ
FJGfXgGUwKW0ftCcC/8/SzXxZTSHOHNGGaKsTv8F/RSrYVnNfec0tvC8cjT9PfbayLwdg84rqMvA
i4VudIWbq7NDKSkin/IdxCcLhro/rZQy4HBpfr4Onf8VfoEiOTAiJB5yxiO/1LAVJM3N+HXB3o8R
Pn3QwEeMz7Y1b/nwRVlyKT+A3SNK92+4SEg3RV1JREL1GYohHoIG5QMhAiqiNabwc+nW7+yaL+4r
9xsyR0AYqlamT3j9sIoUSdrv5opoOB0ynjtek25TyEaHWo64riejfaGZY4jYrBwuQ3qCCIitwJmB
+I2AkeF83aJF/az/Erp/et94PqJFoc7cWQZvMncFo/8WU1XY8FNzO5hzH0L3b2Mb8U3RBiVFJEpa
//Y729HGnIbdD8HcuElwZOw5y/8llDDEyPlXjPXZvCoWooOozI1yedVakolHnebvN1zWWJIDHlrM
0jABIj9jdCYUZkKEfCkSFp4sjCsiRNplh7TATeoJGN2pnUkXgwIxzjkySGaKpJmhbKyd6GLN06Qw
VFOK459tnsjzctGsbYRx0ywVJ1w1yt7Wz7tj8BkIkGFcpt1i6K0UGMU1dts+/pXwfGwswM2kKNqm
xk9j97DgMZMgjTaLo7Uej/uJWftpQmWCh7meScgdTqJqvRhnLE2U47qxZL7skvAB0huJQKY5rcd5
GF0j8HO1ZGTMfnOcA+ICvJ4gY2QfZZWpAldNyBgH1k1xqqgZfVOd3pdWu1RM+Sm9j+9CdwStBTux
0jNCCYVzcn9gLx1CTX7jXiiH0iqFLHX1Ui4jncT3FU3j+hMkc8knLUtkhzDLM11xZAk9lxUGtoL2
6dyUkGQkDKQDKdVq1ipOH/nA3bMpwlSPjt5igAjnJiXMbBN3vr+pY+UiVUpPmKdcuqQgyWxfImQH
47KANB9MI6RQgIh2B/fBbR53nbotpVbRgkA3pIkn35My+XM3nSX/OY5MZrQWwML4IitTjR2Xlk/H
wTwenYXNwMUMaNjtvr+Aj5VI32eA++l+QRLdrCvqoxStv5OwcL3M0QBMV0dNOJVwhWdgVoYkrGMn
THhZBirzJoTJxP3WTJXOrJi+WXPul0LV895B3l35qtPSBpzeZ4mPVcsGFijTecCrsZsHF6lfaNX1
A5+uftVKCmD1Mao3yGpHgnChK3S/yGNpAKVQTqAkXpYHTUNaifgyDGYb2Xpgy8CPfXutPSR76iEu
BmRjfD5lEFd8DMjIdlx+YfF/3RX7SVVM8eDWXQWIsgJLTJGEH3OmYIb5+LH7ZfEkDyqOwdAlyvJN
b3lbqljR6zneciEql9fjmidKEdE8b+nNegYZDU+rXtur7SBdFyE6jFgIV3tgXak0dBoJhZZRSeWE
8iGGtY/krdM1vOcGPIcK2v5k1VLkBxOLGuDHxaewfzlcjoHgrmHCRpKLUuhlW382j3FlZndDIoJ3
qf164oFB1piB2c5PLADZx4mimkKmCL26JkIn/xprWGLpTOOOFuryUg+Fa/9QbhKgVdH/IA0gPaoC
s/FMcAGpsKyMCgoLhZR/P6Bf1ToKsi3LFwD/KRwN33vS4rKs0wZT4Bt8IA7MsZdKXxBiUccBMBHK
MQaA9xpZJLJq+9UUFYUZxYDjYV9/YIJmBbIU4T4YslFKM9ePE9cnyV5rkfjA51GTJ2sn+oAghWBg
ibBH1ED5bU4sbwdVdiBe/MyGLOr4rcsmy/ACjpFfAkkG/1yJi7rf2OEIcR6dwu2peJ5ShqLvaPvW
lGUVPi61px9ztWwwkFFT/sYj88TEqssGC60sSZhgT5NQ+GIUSzz0z9dO1Khejd7ZVUpx1YiugclQ
jChLeRwyfAGbHiURF42MY7unwJzJl1ekyclsTAMCcnpiGysygWviDUt7yY6sLndv4NBJJ1QTACst
9MFa/j2skKFIuZyKCkM6IxpLtN6CaYz6rIhv7FlF2uJl6csXpnFsJZe9mtPKq+LthXLYiHVlEfr7
eRFgZ2loUiCaYTGtQ4zpecdWceO91S6/VTlDrz7edJXSpnVDX/iAW6vQo5VkPCC9IcNySoOqs3iQ
Qdc4svv+lImurxd0BTP53wn+33MPfayowzJmwgUBjWlsWmfUKhmKfqUc/JoX1u26x60I4okkDzdP
XswPi9TWHBogWKO0mJIRl2sT8EqS2rGwrdIX9q6BqCMeExBSOHtG5XC9PNac0pDOYnUEgg8ENQOS
Zjak/AYGqLLjnKyGoQ3kzK+DNZfEVqbalLIRe9bFLrZvC51dMdsK1f3fzY0OM9N8CpE/2MEEhrX5
oWGKgBt71IytcsH4pWMisPgl5vyePzsnFprtjCgf4hvjC7RiPaNpUsKSJXCzekxUTGKyIbHjqv/2
EqN31BIgFOOwAzo/Wtk6rqUWj7s8m86aAx5DuQDiJKD1MnyS0T1J98k+GkUNoRtejx56DS8Cf8Tw
ywXp5noPAD0B37bNEa2X0QkWuTvveI2AG3ZDhmInK0/hfMzeSJRRnhSUbbOw+OC3duEjzg8akwgO
8lNiX3tSyI7WL1oLPqFpb63v46ROaQNOwPEHaNgRedkZqxC5jxEWHEwkZVY+KRVFujutqI2Pf9ES
TDasWEnN2KxItwK5LiP+RkxWPZOxB9X3crX+7cNE0OZew9tfG8QuZ7ZHqW/kF2YRelUkCtHGxBVQ
Ai5GL34aLNdvcj5tUtml4i/UxzYf7EU22PXt8kr5+59B+tfNh5L1pWP267EgQfvS8HYU/y97Op9t
cOjxtRT3LSDhDLNZfOb4D2WFxgwSGE5jmiknJ4dSiJKTSMfZhq/6hXZ/tAagzUGSIlXWGYx0cucJ
blxoYqQX1TDDpeTGxOXAZ3bhiJUXwPAUW2OKl0oK1ch6CswUXeNbSdBaA1QLsVUvd255vm6dgtEn
yu2AWuUwfL8Zn+0/tfRWDWH4SVbPpcLcq4PNz1fUOl8tqyk3wTU2wSFBIxIkTdK761sqJ9jiCFj2
DF0SE08a8EE7mrZblt5IgxBmvSU5+UWNqhMvOYVaP09s8zBNvFdDL6wgU5HH733diuTqA7U7ZCN6
4bR+HuoIISuudk8EXGREA8SyTrtaRHQIsQ2LTniHm3qXlikMsUohaHOBQycmREUNIfmEHNs1Bhlq
kbyuc2Gd1u1gX+l2DLcZukPkLKfQx2mILvt7Z8MErw6d8xqQUnlVBZpA99wUPG0Wv/KRjz+0spcR
nx9rECZAMZfXfcsKWDrQ7h/xqQQdQOvX8g5SPdfTZtV3hun6Ud2yblgAevACmO53aVUeovAKmY0v
Mm8t0dHPGA0if+PMq48Anfayl0Uz7fEwmyttn6KAyZ9/xOV3jE1tgT9zukAvQlvIXTUN+vSVYWh7
J0wZzUs4zwGGc06NPndgvjMhEcCvAjne+6QodV6CSP7uoaOuNvAi6QsGUveO1gVc9aR8eQXvuq6J
cv2iOPqN4luNytgmVm5A5AksrHA+Q5g8M+9/Sx3UM/kSK9T0TOPEs09UgnxyGcaXrn//KJaw4OdQ
sruziaszR/vDU6ndwWbNYg191DovDBLTBgj42rWRnKZP+xV30jOkgUjOi04Ws8ZO2TeaOvK85Nb6
g9Af7ZG0lB7p7W5FNYBXoryj/DnYcxwG3Q8SOeLWfGq9TdUEbG8Z4OJmzfAxcrqnkzUCbHdt42cL
AziNGFYQr5kRofQoVNO6PgjPZ+/aJBUgbXs+YHjn3Cca0YtIWjE17m+V6DZi90wOzfA8s2KwrsHm
oFus285UMG4HZUCVF6nVnrrsbCMrlElQcBOyLxiixJoAhaH6hfinBZ/o0su1PXYgSYo6dfK5b3bd
9krbjeoDljNq5K1Wz8ymzxQUsIrCwD26OgkqfXvB+8R7L1ks7N7p41So8Stvw4x7lSikgaBkQbtl
TtI+BllYU9fRR3I4Uk6owuv8TwrmMctJqMpE8qla69gtSQtsRfUUSmvgPbk2YODG5Qk3E8n/8SVu
i7XyWqR7irN13lsfltDyQ9/LgsrR9/o8U06BxPrhU92uVQ5V23E2pLDr+BbAqMIw3DMpA0tJrwKc
+BQsCn2U74eBdNrf0zJLOJnrdCUIsdBn9GbVhceWBwBLjMlMZN0xt29PIcC5rJZdsSRYqMB1qBer
+2c5uUOndpATLUKfBaMgmXVrUd1DxswaZlFTl9nWQHaPVL2JuX8G6jcNL60sopilAGfbfUwJ4jAf
FAhsRerZkHgKcC70WUCPtGM4N7AXmhZ71ieGbXT2SywjCq2dXZ0tDG9QyH5M1zsw9u0va6tGIhz8
GJ1Q8sTy+YdLsl791995tjuR/Az51QhQoBxZo21gJYKXsg5Tmy/6J4kwfwFat6frG6wLdocRpb0R
QY29FHeF9JUOZ58ByReIw5IZf7Iz5rVE1ogNVaTTBUMGgNl/Kn0XluEVrIrAg5m4EGtn11DssyKc
1326pO2hOQgQQ0+10FRRgn/duWJsS7r9e3jR7e10hakgIc1NQuAyZljmoPKASen/AGHEnEjJsx9S
sOfWI97ulm61iwcQRK8Vg1mAJ/4h7aZ4C+APnzgadrlOlAIAc946VMw2Ou/dcAbRWU6BYlqrbjAL
sy6NL6ORvdr6ytYIGEwIbpkYWtsI/PjL4QdLUzSICYfFZ818BkiuhN+ns00pt73xrggqaUdb5hif
yCUQlqZk4c8P6ZK5EUxb3rjCOFKhfomUYdraae5nLgjpgA6HBPCtmVUnOyGtHbJPfRBNRSg08DUu
2qiSmLRxQKHDNZMBKZrPinIpy0liuxEMDHmnqOFvLI7JVzdtY/TmvpsXcETJ6wN3Yw5s0Z3PBuGu
4hBmREfKrut0fptzrQZt7dnVj21o3522/3C+/3j1gOy0Wk68OctI2Mq6iJMQVat4AxGAyvSZynw4
JbRds4e9XWsw/7UVcej6dl0He/ZeTX5STKCmjJmiMaRsuQ+MYzbzZh5QpyJn9tddM8AKTaC195Mx
mRWIqh+0QB0YHsDx/g0fEYHhw/7/NKwr2Q05us1l2AS1nDyh3W7Up74DYDLRNJ2ptk+cBQKMo1jk
mqPnsbertEB4OHHcMJNwweoZjc7h4nMIejv+HrQmzL0pHAXCo2lFbaeSK5MVjxO5ETAjfu5M/hdJ
1qN25K8xEGxxO79YUc7sGjOr4S3T+0iQFwVq3K2vBb0Gqlqlj8dd9wahZoRueq2/NgtikhIgEeRa
wEEMSDLFxuJPL+mg634lSwdkGbCntDfWmL2mWI9DJ7arBBpX+inhk/+/54LNK7v6pfxM8HwwG+Oc
t2ffMqEyQDQwbInvBg0pNriZUUlLI/JAFt7OQmcqXLZx2XpYHloLT9y1uXQMZBlwo4NoN3i2DG+o
IlK2Z/YFDNL8HIsoQPsXVMIGRijm7q9aPhiVqunDpyR5kHbsxdvMA8ZF2dyegBLcTDFePu1kLSk/
kvu7DMbT5xZnmoiaJ4s+49W/FwEQPlVIIK3tWQbjd6GzlCEwOzpPyVGKnFwWKXaIj1QoiIAvpLjh
kJDSKR791Qg2477I/q2SrC9Ow0KIc+8/9nYFHsXUA7jPv4Vq36Rogq55BCQA/3CUk46+jHgSNBmn
Sl1nhCrT5FGCEt4+p15cmzMJyL8078qikYl5F53FUijeIDg9QtBhnGfzPnAo0voSh1Y1doheM9vB
Za4ofVM1MvUessSXXpXF7H5WN/V3NdJd3Cl3geN3uLD+Im/M+puOb1pSvkwY9gK9AOAvRBYaH8RI
0q41SCoKM+ChMITIDM7chlD/RxOseJv/HFbe8UbOjzigLzVddq2CvZQ6jKpKV8TfFnHI5ZohYsgL
zUhSkzIw8TnDfcAfOpJwoHIa/GjLhbi02mTIQCoFWaaTBV6f9/UiuQfNbPoN0RMbNHy3chmBq5UL
ciCfi9sO7izNIjgomqJSPBaVswlUWdYyRvWY0VSj6KCi3EWo+Z/OfeMzOO5Vf7CwG+1WTn53pZI9
m7qzqA6RBcql8JSjrhDn3T3o55Dibe/WvtTa06d57iQIQsrv6TzkcT5x0aMANwv+j9ohgcGxmEcw
ntqXCY72kMd4lg5mXRdVg/kzgnSL8m8lD7xkn63KJs5PA+9FJzAjIynVldVrIbejPFeGeATEp6NK
sgxLAP+BSASn1YTfUDKKYs7CGJoPDULBcpOmlgzOy1I+B7HSzmVAe4johBuQYs/gCiuZzEhyJ1/1
XcSUZ2zmeJRhhHDm1maf5ZoSF/2k+PKaYX0lxVy0K2zZKyKFqVO8tL1VNcy9MwmwW5ssxeMoI0DW
EJuhce/r8gfRDQy8mNCfad2H0pCVI05oUJGtCzdFsncC9lGTpiQ9LzZcEmePZzfzmYe2tJvBjxz6
S/j7p4U5zDcW7lXwM5D7J+s3GIp55ZgnRhr6CZs+xXHnLcjRwBKYjCt56PZDrc9NOzzjZSGu4wAP
NYdTH913HuQIOu1wrRxKf7K/yAq7oV3smkvt087sw1kCmzF7wF4lkPahPdIq30QIey84w2L7Qn6k
YZIaFTw3hffTjFBqKIGhpCr4W+Xv7ruIS7JbtyQxSKRi8mMeeXWSNnApGkBbFAArKj+WbIqcIUk4
kjwmTJsAKXuLSO6QFXKPG/LPoi5+4RB4HZ+Eielr/cPAat16hDPOebyGl9nuYjJ2PsMTr5GVAM9s
MwZi+R2VahWg67GfMKKC5lET/JVN3WjZSkzIbnVdLBMGHDe7qQBf38DFQNAuwSsxXzaRwblXq1Tj
8zfON4rGl00X3AybjJElaqrwZlPkI17RItksaVA8BeP9bSAdZ6SGnQCINOKNF1G9ifk+SiFGl4Cp
xZOdvHL4nWiv4LLrv8SNg37GnkIasHWqsdRXpTC4tYxruzOegMPTvDOcR8j3BRM0xEU8AzO5AByP
wiUpwoFNGqbKyo17YCcQVgTBuYlfMpz1iKM8NTKVbrBY639Nju97Rbneiy4pQ1frMdfnodeF/2KV
Jd4IGnXlVE0hSljskPHzyoNl1Op7LJPH1aG/zr2PmLKGG6WeLb/5NYM9e7Mhhj4jzhfy+r5JAb67
hxgpGmSBmec6/mN7N+2orphKg08IHXxYHHCU/gQNzCsXz1sOWMXT+WBGOlHQck752UHnZcRL/H9/
iN6V+ckspk6D9SAHjZFVtj48EdwNP00aHl0Rji2PMKNHgoVWPH296X9vPriJEhd1oWvL11zdDFKA
xvoSB8t6qWHIgEo2t5XqAcSGWDarnfqxebCieIQPxQ6unmReo6DDqwPGRg2U+uJDDZQyZ/3di5m0
q2JeddxPmRzU2PEPLOHDzYEeWYI4BJBelGr9Chir8km/3jLCPBJSv+/Gf54H9cEfevNagLXr/W77
YLLkY8MHz1HFM7fLyIC/QFeynYg4YANrT0/oUwAcpB5HLzW9Sp9mEXFPjKahIiNTtAUN/2XcoUuO
0rSLZoa7dnTgGJzskd372Ywlvt36InR0rln7rao4ddaMOeOhX+vQ+vhW7bzmO4nrFoWlwSS9u1s1
eSDppVzGlAj5qkgxYcCpSIyzPZjfzpRUpyOF6h0RtRXNiGqDfkpps3Nqn/hM21gFyU2PIBZW7/AV
HJmQEFPIoY3vKs3y8QxdF134LihjRejUsMCofgAVb13KXpYIa7nrYAeg11BfDAYgOacZSvbWqVdu
COob/5edqVWOKL4GkJYmrggM5rV55YGzJ2oGvjCOJtt2NJq1p+Gcy0Hy2n/rGoeWYoIAf7kJsHwO
1u4+yVSYv05zSVbzMgQRbK39kaVnkj67vLPe/dNlQtuclU2cm0CWVknvUufNUMxp0e+5wYzes9Y8
GemI+Eqt/ekAP7X8oVACZ7ZTer0i/cL7BDHQNQ0POtxU9vZJtU0CVQTCScNBX05S7LnhKHtkzeFt
GMOE2UDkBGlyvk+9DN6hpALbxIsw39Coi+9L28+aG3giLRIfXCHi9XTZiYJ2nO8ILoX0/DcQg8NZ
EFJzGkBsphcYm/KMK+h7/cbcpSoLPDmGSInPtExh5kj2vebpKbVzwboeXRIYSiFxJ1+4HdHEY8PP
gLeobJ5jBC1l+u8VmLHt0GC6P7y37vHHa1yP0Q0ouxipCqSsLTVYNTuHHJkZ+w+v6XsnDMZhsE/m
5eaTmAsX9QoCyK/On6dE4JTaK8d/8IcRjbZeUpYcBXzsMWgc6r4S/qqfOT2vadHXkQDIF2q59Dt+
fXeYkL/MuHHp5nXcCWPnphKcZ9SpgUiK2CtL9ACMtVjNo6PFKMLnX8rpmhgMIv1Z2zXWShkyzijx
9pgJrEEP/FcIZOiNHrfgnjxna+F38U3mAPO00ztsyP6SIVe+7WawpNVdR6LITnZWGkgVPPkBr1fQ
hBFveuvkvlpr7DPSxhJHHwjgyCrY+GvFiQaspJ5stU3egNwy3GHHfy5zawUSrZxS8X2JLnLGnmgS
Ni1m7uyfMsmIArnURthbXi95QOA3zOLDM4QgAW9VUXv4DGVfbsIEb9CFO+3cOaBQEbDjCpgizakN
glrTpLEK8+I5BTiBDmZFYGo+m+df4YS0cE3p43BjefG5HvLQhoTO3w0l3SHNRGLvZf8MK/VBFDNU
p2tijeQKGfxCLaTCzZVyhXhQnmPeiVT/tDwbGY/jDRnEXONIOZ+arhQjJaF0iVDwRmGAwYt+aNbI
/LnF7BMRKTRx3C3+XkCFoHCBoVp4B46VMjSPogPLNL7PWJHM6R5RVRrE3v6n+as3cYOkDL9seWZl
tZ/nzHYvFRNJv9XwoPW6RvGgHlVDszZFMmz9NwyP6RC28e0/nVdqctvfHlDE4CrIcnHfj6o71Hgv
y7JiNpHqZmmXn72gPk5edYqT/ApKrfYl5hPyayS9hefxSFdpUzW20KRZB/QBSPRkTIjIMwXugwnG
aQllMbR+9+BMSM6syhbhEBk/eogyupw0OWGIY1iz1i7+UNuihD1Rwu3uva/W1X+rTjY7cuBpVUwp
DZrx1BKBuxc1h1iaC9//y9FHP34CV94teKDKdmNC6AXEBVse2R5UXUrhcTpPOPcWhH+16svz5GL2
fs8bAqJMZaXjqM4LyDLpqlwbuPFOLmRINHrh459iIk8H2YPLfTitCodq1+L/CYmLXs567P83HSsr
jgf95b3ulBuh4YYQ3h19Z7SRGQHBaqWLUTdK+BpiXbEA24RXb/oQ400txlKpwg79hZlpBPPBsbFY
QWfqM3X9Je0djVGjFlHjsjVVBe1Fr4u+LHzASSCARijSkPaa/6CfhCn0yWYf2upYdAXnUHdaOecq
clSQuGvZ4YaVJZNVALriU/qZDx8S4byjyISTuK8WJR9f3L+CwdxA/x+pAE17LhCrTD1Y4B3uaqPP
tVlYFnz87uhR0deFN++bcUEnoNL+oM7t5GRDo3uYIXHIhWqSBNs+P2cBFT+t5gvvDnqsemUJ4bUk
Q1yyUPxfqVqnKvGNRUMUOxvM8dys7Ene95cDXrqJoPT7UP+P7vVSM00YMa4Oj+44ObG2U/vkT7yd
GuP/9nD4SPB3uUD4qqTOLtr2mvKITkteoYuu8tARLNqnB3YRLAQI3UecAzEPAiafeolfxbmMM6en
cB5X8DLcKgnCNdIn4DmaE2FQe1ijA1egthiKSJEvl4FCxymxHSE5jiXSYKH419RlmV35BZ7nNSU/
pC/5Q+tjtKkCT0PwN7t/09G9c6Koe1YMJ0kwkdhYhXzJqwDX71HUJxD/KH7WitB+53cGdk0ZVypW
44fw2iCaKI2YWRj0cRLvbCXLFyiIiiYVjWPij1vWXLTYYgtkJJVq4AOFnEQ5EupCzFBQKKipYc9M
aADe99F+izD3Ki5NiBUw8fWhsBQngcHr42+ot4HJJ7/ioZvc6h6Zt16yVtAkoHmK0EyD/G+vqj3V
UZoLzKLyywBJ4AJdIzYwyD/k6VHh4jRtovvqSAdxA08YH3ezMCJKk/W8EMyD01PQt7ifr6JadNXE
4p+cf4o31NqT29O7S8rwsYKMGXYeckS0zzQl/Tspw/Ik2mQgHMWjasb+ta/Eew1H/cCOrZ0VCXhn
K8UKhd3Pu8bTwlHIR5Vwap18TlyD/L97ApTTkLu0upHn4BmfmXDXRFbaSiix1fWvo206xBtW/DT1
q3GjaAFork1wXC/sLn7p8b/Kd91wKdMA8rDaDFTq2TczJ5VPyDXsW60Z813BzuQjxytPbraMl12Y
ZhkNS++vwHynN6HxIyzlPXp71Cmu6wlicQUXNfXjgKJdHddQRJSKKoBWpIzzigaCGT9tOggjZQ3J
/mnnFAJ4JTPkRvy1Ql5SHGMzhJWwX8ujbOaxgZxRPCRtEJrO+F+DQ+7LVN14xu3/7ULww9jh5axm
VrDPTYc9A/qFCOf0EKy+0EgJ/D576ixwH5f5PkZ+J/Txc3Gc9LW9ttPIbmMPrDHd/nF/fOa5ORCX
OTbHEHSRh0vKlhJEpebb3wMYCotsDzd8hYCww3QN/W2MS5XMWZKxAMIAOQ/DSX/zBMo1i4ox6MmK
l3dmIokTN8eQdzu+Tz6q5wVpVpxcOOfCddXXD5mrDe1DORRXe967IYUwR3Dl9FXUj+zsJHk9H5gb
j+CMAuy2F+cNff7TR23lSyivDzuNQHBgNWjVeuy31/5U7gQYb6dLG7lC5YMMQxTOUmMaizn0Smj7
w++LJ+SJEgpEYBT18jIjCgDz26Kio4r3Kf9z3COYb74tsAe/AVlbyaBikOx6PsqX4FJXvN7gWaH6
aBm++dFe0+MEBtpopreiJyxU9T8QpWHtFPpQZWYIbsoYGWpmoprqzHyeK9CMwvQuQ3rygB2n4Mx8
yqzUDykudKTReUPbOPrcG8PosfK0U6WyZom/5AoUa3uJ6sXE4f3FiYyPJ2vo62Xyk2ci2dX6LxWS
MfkschlM5bcIcDCZEMslkRuwt5sfn1yej1vqj1pyfl/EyMprZeLnLHQy29XJlqCUyigqL0VAIQmW
/3LsM0Wgfeh1DPkERkAlcF/px7RiKWPMNublmz+8b44zFqDEPeZ3cLSoNDotivMULj275yj8BgIN
abvmnw4vpw9trkE80Hv+0yxni8k3yFOBlk+IcjYtNko2M+BrHmgffGVYhBBiqLAsYzdr930gBir1
d8owCb9KeZfKrcxa4jz1CMAKqHDXBg4LDctzxAJmMJiafPYqAN8PuQxLHFsBXfmHT7jcRJ3yHtUY
e6f+hpivYP0DHs9iS876K5MUXsQCChZ26kYEnSeu6wz4CmFK2q51Kc5TI+doTC9+NpeUIjIRzH0W
SuIw8KQnBJv6NTAaLJDfUfpL03G2gxRMLuCD8AK3ifmb7b3AdqALsCUbcoSWUcU+G45I4QfMUjDY
jLw4wBMnmCYWIrPJPEo3BSwOQeTKdyYVX365mA+Z+gjPe97MtRvdAi9lOsj7Y7Wdy24K7kJ0d04h
2U8UZ4Qmh1GJ9TFy+ei8d+CFiTpdgZquXGk2hP9ku6B+e3Tlsz3X5Fw04ELW92gdHL2XzNmmcrD3
byL9Gko3X5HjhYN6TBXH3ia8fkvGMknER5gsoG48s6tXso09YDsoZCHH81K+uIJb+wtJ4THvmW3t
wU//U+ynnPeFLzEKhBtKfnC3Du7JwtZ6Ful/vn91cmN7g35KbJO58YaGHZmbKeg0NHJ/59toDA7s
PpqkcemOeOc5EOmlKZiT2gnqLxtkPLOCLAhVhD/u/xu2kR0/Sdq3Rm9z1gfxQeIaZxlCcQCD9sXS
thVX2AeN9YZ6ykqt8r5bNxyup2KTor7vDExR4e0V5zmJ7xu5/+W9m3aNmycCLqJtY9ewFSm/xbIr
a8dVGhoq69hWWf4r6McXNTLTD1g/X9bwE+OXy7Y76pWhNmswaJW044ATG6d5qQOUuS1F11uIUbU4
D29wAPoXBbNRIi+YJNUvfpbobq+UTdTZ6ezqrGApUDKsk7aK1g5+Zp345G5wfRSKhxsmxC6DFbya
08QGFM6VGgOeYJjZ0vfDkLUtMP3/N1/BKlvCFict5UX4byVR7/6Ne5q+fThUpGce3y4bPjKtt6QZ
EZZcm/ZvvQyumOkLFmlyZU4+0ipYRR3AfY9gva0RlkEDWZYd30LFaHt6SQJGQJhVC8GqFaBk48jT
15Um6v7rTyq40S7UX9bJZP3HhTICMo7JxxdZAfvg/KOYx/wlmGsWqKJ8xANyfwf2hV0bLBAbxzX+
QyJHc7W+KNy/0ramacatoQG8FzJ4YXRYVOreIaY2ceKwrUAk+RVMzMSlPyzeWrX5YFhWAh4q1Vy1
dLceyKe73kL1cl0ybia2Ryr+mRj9+PczwWr0Krk+wQZWANCRstUp3RBqaTqnRACrsSaaPt0v/iAA
yol1zYzVmyeZJrEh7ae4iwUoO5cvDTnl9DxKIB5p0z0qunEfPdtq9HQ+lSTAt/tz0CEttd0YjQvJ
IWxQ1ldPdDpVizGVA69oHVMHahrCRwJXpxE3WN8T6RbvnSEJ4lpR/CMtki4s9qKUKmSpCd79axxY
d2ARwf8Td7nJx4A4Ukd88oxvq/E7hzYSQMeVdSC3sGYv672wzgBCzTgVCsMLkebu0+v384g8J3Rt
fztOWxabkIAPJiLxP1xCmJuTwO4OEJbTMDBorbVSagTPkWpTYu+Ojt6+earNmZNtAnDjnDnyp5hD
uAwBiACKce5n1Bd8Xw5JitHVxQNjq0tFxxWc2A+URnIW3DvedN8pkmxV6BB5Iolkx95veBox396D
QsWFLY/N+Ld7HdqaENL6XQPKm0/mVB0vW9gLJUNwLW/cmMQxtnIJzUcxBylIaMPras6H8EVhCF/a
54UqzaSUrTANcyVGor7ztHwUqYsgOgTeMJj2xfQhS+PT1narI6j7J2SAF/qbMai2BZ1ByW/inZcQ
oZuFhf8VeJq67bREw1weWiQwvTSs27B1H9ccxhepPlJHrz8vpHrVvXJx/BdiWFwXYQRu61iN/KCg
HGMTvIY2NH5cAf0k+tiWN5EQWYs2H0jJ3XPJI5dQfd8u6qALYFVQCXtAQNEp119rdLlCCK4N3eGm
b0t078AjHToafNolCLs/48ykYimEQ4zZToeACTk8CNcNFX/1ODFdnbyKRwVKo9rJ+ZjlltcSDe9Z
ir0nurQZGiz8WoueE+A75W6PXrDhFAjuOx7Xjl5KDp1vS+SfjETiSlFnsrLX5ZKgueibJPJKG1g/
H+Iaeiew2EESs/MihCfobgGDIFO30NMPsdTFNuGWKpj+xFNkvYeVzn/Xsya8rNkr/NAB/M5abZtO
KJGHXoVXz5BWoYFY/TtazAzNJWqM42fx8lSWwNicRMzrKgPN/3sz4VnO7RzJuU0atxUqh0aYmtNM
VG/8vxtFrv44pfUnhaC2+aSvHnjet5fpbm4MQIIDW95KGO7nuTpjt29/GH2zuEKVMV7P+hoR97HD
x1AndkALscTm8Psw2cUzYlkEL3LpHvfBD1LyrLX2IX4MIs/5m/RT5foQkNwntCxlWB4015DT/Ucz
iwToLlKdwG7Mh5tFEhFBA9vvB0aP5M8ECZi4TUMX913zn/y3L+vs4oqD6zr7E9YpNOYUFG/XeZ08
Q7ghO5VzADhQYL7mrkHVd0ZkrXW1vQD9in77U7eiX4dDM28mU/G2rNUgBoYsej92LVf2VwgALjMx
rcDhnhqyWlS0hW9AE4PtFwWhTmJBltoPnhOVAoZliUJaN/atAdV+/zTlyeCV5QH169ZrEnW3eS5V
7I7cxvUWCfB03ysyoVJaeBMb9d2AIxeyotBvgjVrYhuNSfR1NkLG/RVA1rWXfcirliYzSerlR/5p
LMdAPeGhYhdjtB4r9B0XTmbvzsLDo9lDd1ShyP7kL9tIqw+b2CrPJk6CDNTM9NSxTIwBVlojmGfn
ko7d7UUSI5x2cxJBeQjqP3Ll9IGWlJtegIMcE238nB9ahuJwCyWXlYXbZNaiu14AXMkWJELprjwv
0SsXxslETJPIaHmo1YaQ+6BQ0CRKdwwPoznVFh7w7kVQ46A1/g3dpT/KmyNHd875M/rjFY/pR6bm
hw3qEcQUmiMCNESeMt/4REi8oaTWodptbtDSH3l7YmoWgNrA98DwcZMb0NMyK6aCIsXoSF0olRLq
PWbTVKJeQoXf/QzCyzlzobTqqqNue9xod5nxQIeNTHEmifC/XWCtH7FeH/mm/9HLn9eS5JBjrMSw
PUH8me74rPz0UGk7comkE1Lc51XyID7XVnXLRYiXDaUjGkyHr+9b6ywyJhUJK+ZDyqnbk4HbxIVp
sr9kRX8LiPPWjolKZKnxx6thkk59qcdJsMaUQviovQet5uDqD2VkYCFk/6gPq0hDlsL5PH5+G4P0
nlWaU4Pg8RxhSniZcMPTu6MTYWwT1PO2pl7YT2RaN9p/8u6sJOBVAyc50Pp+xV4ov1OSDkA6t4RH
8i9TvV6wkNeKOzYosl72bXGoc1zr4ilL91rk5ccE2sl6IE8trbW6Ye+noCcCfv8SYc87CwUc2xFM
dRZvfx69Jru2akDouCAlPoKUiVvv8aq+19VjAQpf0l6tuf1Gx8mOyQLMd2lqMJA1ILpJ5DTsruld
Mv/TLeYOMFlj+bHEUPtN6LmadIbmkP2ym6/Jn9Dcfp9KxwL1BG9t2Uqh/qtGg3UbkwHDQVnsa3p4
kRHlbd+SBk1RkSKCDOc3w5lJKYWyk3kwQvMzseJmVfn40JfufmHx5OlE8GwdBpJFK3ohG+TaTFDM
VWAYK7FfiZIbYu84f2KqbiLjiEZz/zCijV8knkZQYjM8+IGrt20M6IdxUWnZJbr2SPIzawiwvZId
7tYirB05e7TnZja/7ZPxGwbeDXhDKqfVZEPYwHjtwvU5YS1UsZRcJvO2e+Hoi8J8/sHw2/r9qu/e
I2oTmFP9hda37Nhv3KNkpkqVGC1BTzv5MJHEoBJUrZVgeVojVufI7guwqT4yV9OdiaKZFvXemnKR
1OrSCXIpsi6rlWbbiBp1DHelQBJCC1u1bHLvGzIciukywRifbSU4hcZ8vbkF0aBfSJkFk4YpRHod
1en/jQpqX2ArLAcSbUPu6mLPX8mQltET79zYm5cKaFnEm1Q5oYzY5v8MRwZSVYwW07Ggi1djhRp7
jDh1w9raQOiHmv5zqbfiyKr2ez6KGB0mpSScUTUKRtwwL0nWbGtKg1i2w6hEOI5cFK7RR36m+0pv
Ndthk2G8x1jECuqpH057Jzbex+KbHMpEafjbN9jOPL9XCzqiD2Jrjplfxnp8Hwo6CIJ0HDCyWLWY
0+HzUxpyX/Lum2HoUePq3pMciVWzokrSgRqNMAuiLquEOQC9j4mXEo8r9BVUaRSy78ub8LV+csgZ
/f+Hpwf7FPdiEMaDS3t0vGwIIJXSRh8ktBBKiWlfXgMloLzb/9sHmaPi5CJwQoi42MeK+wQhh5xS
IiB3DLZ1mMrBv+tQr7zrkp5EZmI8lMIWyj+4mHqSHCz81MQLCd2bvwdtIrvUZKZaKD6OrWHvPESW
1x2B062wzZpbtTBfcSqhKbGsQFBIi+GMRtsNLg4U5hvPBbm30nYyvh4WEjHUfNJ8QFy0LgbsEpGO
9H5Pt4gXbYxTq3I8JzZqkv44j+ixNP57Lp6SqlEYVeBnNH7Hok1CS+SLihpBHz+coSwNiPXu36//
MnsGsqqp3vReFxn7n2hV8A/IxuIYBuuA8OQkWKViI/92KT2L4QVyXiTfY0D9Naj9PHJySMUhAvtP
h4zava4YWoNEVKxm3D3Rx71nxjzSNBR0/WZ7drilkmNvfk/zSuN009cG4ukC8j9bE+fsrHLncjaB
QWeWAGlC4tfFridsK1PHDfL4B9Reqer/7thyN6aaey+Adk6jMxy58CRp7/xg6SwJdlsP0dYiD27L
lem5tT006ArPuJ38KhdjNO4EPd6HH4LxV6FYIIjoPxc8P0hEXmQYdl1Nbc01qr57VZ70q010SUCX
uPW7eNOIVRO5fo1VBin6BkmDNsMsidPFy6oHMsUg06KAFPc/5nMq2kFA12vV/ynTddKt0R8esrfA
ApyrsowWCfbReaOv5+SIe9S1StT5JzU+v9kAt/pQMgO80ri2UNUy8iNbrM9lNs6jkrSBteAJu5er
mLb2gQTaBBtmnoC66UdmuB5I+u84Yd59tbSzZmwfyEfB0xkxlTOzvrqiuJdVzh4g297OX6Y4vSCI
bMIL6EVi4bnh1uef0Q9A5FPbDH6FavIJBr1DQgeBEWzYfPThK0mWNtEyB8M6zJKlONy3n7KXCGkp
KsdHIO1bodJnh3RnK94W/uYcRpYoGFkSl3NmzHv4xYvH8RdiPCp0fdsZMtp+sA86lKGM8njAmDKQ
PJQ336qXAK1ziKJzGhxdt+DgG+TTRtM+J+7DDs5qp9RR43IqTs8K8ahsVxPRo5YhG/afBKgTsAZl
dI8do8SvgXlNhpnSUtEAQWRJ0LukkuySVTLiG3kqK7anyFPb6Jw1FzAy2zKFw8JrOBPAHXFxx9w+
uCoy8CmRYXZgK+pJtKQfBST/EWzvI25SK1dImAX26bPLVVPA1bXLgWEpGw6brV5CZ3Xg2g8ajiYL
kd0RitXs79Owc/bnOzcAahc7EpkZ7WyOplo1ustRcI5pk7rPBWQrU1GJ9yvzEgnnyqpFKL32ttsk
1OrSKD9LI3Xgfvu9MoAkg/bVPe+sD6XRFw5kkGrroSQVy7jLJxGGKzMf8z6KH0RafZQoCMeBLrTz
xjIHRg3ih9yawRL8NgD1ml7PMJ2+WZ+HXEHMKlFmIp+IY/NVG4uL/Of0abqnSGgYpV53sLqYer9i
DTPa4AfUu4KtWP7fS4cOgQUUmmXmy4b7BAc3DrrO0UMtoYGlySmEtr4sSv1oJCxoXptClj1hC7t5
7Ve2lEZ2ZNZz0z/wNUzwEg/HAtJ7iAjtQzwH+lt/d8ML+3vFo0M7uJfQtU80UqjL3ROPE77ZVLZx
I1YDnRAQ1U/ZaAkkgI0Zmy0QIMW4c/Y7dP9ZDGQzpS0hhYftJWfY2qRvrC52L2b9zKaPC0rS5Mol
eVSXuCVZOqq5Ph07dDalF0BJgk1P125+BDux7BpJnlEa1LqsYAlWfRI1lEv7XuTpoVNdvKvkfIyJ
zTMXJ9NPhZdjji1awdlnoi6uwg4TmL/1MAtgYZpME9Milq+7g3/0u6OsICKICTcJiwsWHqdzLVGV
Yg2N99TRFmBN2NHIAJu61aL6ykUEs6HRM+ycSpMZc4VqInomdnkRLIATQNIDFGtlnCDk3IyjGtwg
AdQsBw6LGcQYrWMcsrDh4OQmY8Yu2ksFQ1lI65xLVLhWhZNURjKoYuMsbWAuJVegEyud7+l4+hPQ
2vBDqq1XKJJTgISqR4CdoGnnrOR6FcyCDNvubtojr4Wt7WLaB5VOPhDUbu1nAkDX/9oW1a9tRmmp
DWsFxxxILERy3h5pkJilhgvSDwrwVEXP8apFvHZhlPfICqbb9RtohusNhh85J3ukDw5DkqGkNnb/
9LJm6m50iY9RfixqU/kqTiTDcYKyNJu1ED9rwpPTaeOD06Bo7yhjK+zlTZcOMudXTuc5a+FGl1I2
aOi+BhFmXQ+kV3UMvA4OZx8+9eFkcXLKHPJDgiW4+G5VXgS8lKE7QiszAOxdM7Sp8NogmW9K6oG9
G2oJk1TSZ8DLmBMuNHkolH2uaqfdIYAwyr/2HlMWS14TUcnpa+8NkhC/pGNOpr33J9sJ/dgkn9ef
yXf014aAqJtQoVLxnlCetf76vMTrMEK3g/xqj4VX4kDz15c1dzMl0703bLBydRtq3jeqmHNnn4PR
FRbk8JDCtwg+3I05ANDE66761xsbmpmoq2k+Owv37jofdZI1xFgHRrxzgf1Nd8p7UiT8+vz+ed4M
jsgMyxJ0o+kEqt+6nkgVnOtdtx47esDJtvsl1mddRH0/HlT3aZG2/LgJcVrTDM2QR498CKDgja2/
7tj2uQWWu5nAJfNMqD7z8b5yfuLlR2V14hOxU2FyS7kkJYy+HHZmfGfrktsUUnMrm3vANp1NYwfu
KDZwJA2BjpGEf2n6Zxf9OfzAgAf0ph7Taw1wpASRkb3lOa91uqKU2mBOIr4Osoc4f9coOxV9QBMl
6fyZOUKAKxJvQA1vBgw8fxPvXW2UyG81cHtxcZ2DfHdbytmFrHQnKy+kEBnup5TV5h7hGOwqu/s3
27YbnfFVmpq5HSvvLtjCxcYwM/EQJx5y0tKq1/iAvXXFX7JA3yNyw55+AFAPFLJuObU1RyNWziyd
gjLxggG+qQrm3Mr3MIAMIzWptbxiiMGQ20XkDwRP58pLVT11tbQRuVs0JhcOrgV3QfF9fgxQLbeA
NnyCI+MFNTRLpDwc9nvLcLcisDDDzofKJQbtKR+60zLhbp/TttUEh1LUk2DpFSPeXLgVuf2o1/id
yheU9URVXb5kxcsgIyFnmsK8cF7uzMGLR5ne29wCggZjRlHzLX8oJzrzoH8U8Bao8GomtH1tSVGB
mpfeTgSOXP9lBYFlWi87o8aQjw9dzlvWEQ6XaNmLXSDnAK3Z634o9OVI+elc6w4JOLvjaYc/xzXh
DSAr6Dz1Vz/YQ4Ns9ZkROsSm5iqJl/AU3dwdNH3+Ttpjiq3IKrRsn9Su7A4EMMpKQWpkFae61hY9
BvfgbILFCFqL/QfL1tKxMfcYPwHBfsT4Rd+ombEoT7lyiSEoAZ0eCrlnSB6+8zrw4kzSGh+zQFvH
56Wwq/QTX14SZTsbdFxbVG83Kn6nEc4ZyIk2vUJerBTBXU625iPzkTW/1svL+MiuRB+9MjOH1KPD
SVO7f/SPkLPBnPmaRj/Ob9s7NuI46hRN2inq0rt1DnPWGPO8vtH7dNgSllqgcZyEXPaxozhpDGCx
mVT0SuPdBktrftKwRvdXUgQihOi8KMFcfigQ9CDVsfjfNjlRpVVNj1BYauYWbafhSX2c+9jSe2A7
O0FvHVVnh85awhI4s40C1/W/f3+qBfy1ztQFlguBJXD8khdcIuE6kMXEzAw+RC1Y47aDRuhpViK3
cgbZ3FnWkHXL8gfuDZ4nM1ImHQsSKnHYTJ9xTwox4wUoPzrQQ3WpY3SV1VHa0tB32YexPMgOU8GY
ga5iSdbrqG2utCiehxPW1ANrWqgviQKqHfXkwqBTpetfvGcmq9GP6z52tecTVhqgUiyXG+AL97Mk
XgjZ8WIRJEuFU5EBDgkH+IEAbRW/ESfLDwf+o0TuPzSEKKda7Ubukw4AV4tLwJGq0szCKADy9omQ
lc1nXrI8ue7lR0KevIEMJSltZq/SDjVmGWGrBJuVMXwv97cukG6JDYK/ZqLIdA1w5r/wercJIZZk
IL64ouwq1CuAKkx1GfE2cSpIW7K9rAA4a0Nx0tiPh76JKXL7XpHyBTTV6ZO/oUBClm+5CIEobGxY
d6X2mlIjlGYFMXdOZPPlB5yPJyGTzOpSTmVNMrdI6XySfxZUBoE05UJA3ZcHuBRQQ3GHX/bfMY6g
+6su8Ne3ASARuJsTNbkbKjtS3l/Gef8yQSGa67Pkzw8H4eqLgizjnjz/SNb6QT4F9rTu6Dn/747b
SMg+842ZhujPXLCyfXqLZMzxSytN45upnHTnbFoKlVwp8nC3U5DBBSy0xM0z345eIZAH4OLFpny0
MVH4rYIlZ6oXvP1W17BrA69JmwmcTrA6QSkPwN/H6PBl/SUOx4rXwnKEubHfG/BcZ0BOwpIsteqh
9DzWP/9a8L61bAxnhxyD+04P0FqmgcKwsjd62yatCZsRAvKJZ644aGQHpVDI0IPOdtB9CDVmtNQZ
QdBTIKR4dHYX4tJQ/DapEJIc3G3YaVkxH1nZDzrNxtB1nwyPDBxAGbA1xPb8n67UIBaaR5+RH7+O
i8Va7HC/cSwEuNcVOTYFYSTW+EdQgY71i0EragT2+TRsMQqHaj6NTGSZi6WH+YBlOFrltocNRDB8
1SR+oij9pt2U8J30odSkWJYqdoihr1VEqrTAeiWqljrR7TqwY09FDXoLgK3N2SZpAeTIFMlAWViN
8ewXAZbFvX4Ix+05xO6a1YGG+MrBYfz64rcLJrsZOX3xGQpC/hXjRJYWLCQ+vAIVeMKy66JiqdSm
gF3d3cvJZGprvCHaB941lFY80qgC5VYY6ABM673z3mdZbpRl15uthkt9yp2nfIVS7HTYs37/3X78
T6NawP6X+mVP3Qku1lOu9L+xFoV6aEvS5RalsIToG2JnJYAMo7M5NLQ6iHPWYSIFtrwEm8H5mCJI
k+fjV9L0yfE3ujVJoEWgWQpkQB443dOtZsA2f7J9tSLVHpbH7zfJEv7d61GAHInbYPAfNSq2TKJf
2PcQ5YhF4u3u5Esx5fLDJjEm2JorZjQDSLnCjglMtiNFA6j1/WbnARBpMRKgYrfrfMPREN+T7/ku
nN9WRGdFjJDUPscSiRhC11EHY/SUMF/qr4Sp459L+LR71XiIkOdgDSG0VTt/Ul0XrElEyCEx3QYj
iFYu7HyGwcKpU7Tf0ACVbA8aSZP384hz4tNvp6z1ekR6CPQa98/6hnrFatJjA3UgRfS/XUMaYy8o
1LuUbEURxS3wXWflonncADmBVgPFSHZyZCGv3zENWBddS6CSPc4Opw95L/phP/nP97K5NlciQLMC
SE4gi5tXeXoL4Z4/GjsDEExQMBbgUy+r7kc34LWsB6do7VCnNE+L7nvM/erpKyGpwM52RdFEHBkY
wDtQl1Khjx7S2XBnI1TJXqSCqrerXs74zHsdJkbd9kVQHfevtAwegHOMVnvok4pGJwdQKvJBQon6
ScqZRovavnQ6lYReINuaY6qZlQdiT7tbu7FFJdp+UnQkfeHI6oZhZvzJs/3uJwSG6kfLO23H0BC2
qzTJp8UFsKXEy2lgaKMVrz9G0sIeM1bZbvGwx32P+9lb6ciYK7Yp3XkFd7rb1T6QDNn9H+TNcXaM
waB+78xGlYc5oJ46MENZ5wg3fTUXWZBk2Byo/4ZChrOZD6+w8qWHVGluTPrsFpJa+QyBPs6uoFky
NCpjN2AnLxwUlT5BVHrP2wtZlQdmKUqvSdR0AOBSCx1OuGCbZHcHNOthgqjo7apawY9EBD1U7FRx
oIPXl18M3mGHcsxPTzdMPV5R2Kqaa6vFwyaMt9591omWcSrdSanBHGe/pnXnv4WOQYANnraHwxSj
a8NIuiS5eW3ic06Kumw7KL9p5SSLpadRRM2pqv80GZspdQ56jstsJU6MqQjltmKQb8NB4bz8R5K2
XccVqu5MD4//TpfgHGhX9tvgXOFYkSt7zEoxi7jy37OevontFHpzAdncCq85CxQ/8Ofcw7j7nuc9
t3BbVvWndywCQlMg8U0Kr3kZxBk+hKBeq6bdG9QJ9q5K5m6/Jtt1ZPgw4zUaMOu4/mrqs5vmnTEL
K1ZTdoziGtIMEWaM24fVty4grP1pfmOPmawXVHTyF24FH2M1cD8oBX7a8rf97cqt6WLRv71G1FxU
TlInyRcwJWAyFmJX56nGMlJG8hStaLVYcG0RD8IpFXi1GqT/D9NqlM4EkuOEWv+OgXzmUIWNQPFV
g4cQwuDUzb2cFFJJH2nEit4kbX2SnHeedU6tDj3ldDJDo2T4JuHeQzv8uBvuO4gNX9nXys74ZDYL
dwvjryiLFW+TMECNHwnyV+RSrKgK2o5+Rl8yI3/HCKTwEZR+pDoccSo1l/d3y+P76TptLJ0l8GZG
UJ3Xqts/+CrimjrLTfPsBVUQMt82ShjTCRgJNVtfdanCX+LkiXZzgaTU6Qcvt15WluLkea/btAjx
IULwTe+tkBhMcyzQui28NdRd9o9YPIUD5VYqgc0hNJMZTlpa8lLFdXHLCFKQ4loEuUofoVwUjqT5
xQcOfXXY9EWwPSKyIoJ2RyvS+lxuhrpnOwo1T38QH1lCzKJyERHN3UbgfxD+OrwKLsjh1LOmCjMx
1IeESHFwBs3YxeICSdllLMnmTX6iN6ajl0kcieR0ykYeNg8zMfdtGcTx1pbQwLKjc5ZUUVX4XlY3
ZsawEXtVPSrkLmK3GaW232woAxXNDxVEVzbMaXREMWxIW1dLYefpkKKBEBLlqvEJEhvO2kdWdDtC
sZOlVyMj19PULDPV8XYrIfaPfgoL965UTppR8tF0gCh6Be4sccTh3W7Y0uibnOeb9KBL6l2LJqah
gE4FOnxz+2xhgfjjf9kjWZCb20Q0do9Rbv3KKURqv4BFQRC5DU2/uuEUY9k4WI5SC0lxs0IZRFj4
sVCsuprZ9Q9rATfOsdAFC3BU7S786/n9EHiHYw8sX4DLiPVq80FObyfs0HfPs/bVSu/+b4/XJpjc
Nwv/mnwFyHdS0NQScPpVtPovhULPpyODXHpY8+l6d2liLmiY8Wj3RtJv2LPcoixiDYcmr02kjbB8
tOqY/5KosjBZ7vwhlnmND4b59OZiE8uaLtx5eVPday3ieW4uZMzWTQdVSbPdCL8RFOjDCWzZaN21
gSdIfu9G9QkY8+tLikNTjyQg2rQUKIncw9CYbSEC4o8F+7T3xk1Ke5mhmgJSaMyFM1xLAWb5IbSc
LPVlDNW99r7UC+Lt4d/LlTHmjS37Z5EEyLUkHSiQVrCPo72Ihc/xCsYk5jOIm09igolfP/nETE5D
G4dwOKAtWRn+7D4TsICYe8OMJiO3d1V/kYYx/3IYYNT5r14C1mC0N4aH4tC6q5IFibxkcgIsHj13
WDFYN+SETt83Why4jnJSQHgFsLHtofVz03nuUAfyTZ42jvQb8XnlpX+y1lnt/ZKwnsgchRNNDsJK
W0wHGJ9tlJ06jJ/3BIAbDushRSCk/Fk8yXZSCTk97sS4+o1SkhDntaHiK1AxboO1EOI12lE3CM9r
speJMi1yjy94vWlVc4eT8dDCAg4DGhCa9hZMxl+daqTyWoACvBOxQj2zMypBlpp5tHRjkHnpkgDm
2HGlSfXEBaP/L4/WartIF1V4Tm0gWuHMmIC4FK90885YM19U5AcJY+XxNw3EyBRnOnK1lJjuPJMJ
pURABoMXI3no/8clB/jr61vMCL6ePc61LydVykTUF1E7YGkfsej+FuUwigQynWjmEI6Uk2rUBRFu
QBaUHHpUWtTd972L9GOxX+TJ2xOhg3T9OQX8ldZAv7aLOtfKEDyOMnEt5SK5qhQVteUpSHK7RsaY
m4eLJOP4SvMImG2Q5fs5M8ooKS1C5xLSb63zmGbUQRC5MsEoHWPsLoBc+aMlen+0TPmwuFwPUA3O
4GXsHReHk3BvyDPKhAkmGQdymn9TuZC86lsoJRpdggp4WbvWH67FgplLVRlcqSku+C7CVWe/tG/x
1a/q38su6IQ9ZpirQqdbsSoO4+miKwh7VFtLWE4huIVTujnlRwDDOP/91fXWrud81FQfKOKg4FsB
+O9ew4iRUTd78xl5DU0ZLf62yM0MGZtohAod+vomYVho+bjsz2l7g6PsNxpE7cZPm+XRbkNRz2tp
AWgWSr7JqVd0xFcD2tEswuwio3UdTgt0EwcbLG3WMbq2eh8TZ0oKJAi1X5RoEkaK1wvM9FMWmvJD
ul1aBy7Y/mv/XQqVaf/CPMM8U4N81hKPY9mM8kyWfWnycAJPjlycW/lZXxLEsyftnJ/DhTyhX3t7
1FcbK/vV76MTs1yvFBh7ptA6uC1ZyU4qrwISeRR8AwNrMCCUOLqvUFURtmGNqdq3MdQA+DwReqpb
ca3RHOVV4+RB0TIEAf0RpqAzDMduWJDRaupuPQPghm2A3S17+gv7HaLtLO9UDsqQvi+jNoEzdl1J
Ab261KtZLkrIjhNZGE7Ao9HYvOgE0VYPmL1ItQ/nlvtwcWnNeGf6TQYIUZv9+Zg26CliAYhlVARD
VZ+9fNfx/+LRU9InPE2qr9NtO2jXOfRwHh+vJK7XRV3GIjmsXWAud7MA/1bghnC20+85e54bCHJH
18lHy58CF5/Zan961hhrcnLcFkPL3Jt0uWJNMC+vAk0H75NsJ7IH9ZRKef6ckSeYHU3szENSkLU2
HUaf0SVaTME4ROU1dLaUrMAl+Iwr7vjspdMspF5soi6bg0mAM+TunA6QgUgZKh9Hk6ZVIERcaiM7
1tqbc6mnzYEiIJiFAuF8K+MVSvNr92B6sB1p+Fku/79cnYWNAx+vzuLb8FjEovGg4p9WIcofK9hE
VlpJdVjp2AYW/bh5V8rqfElA/i3sDf1Wjl9UWG7GLl+z/WNNg720wt0v361ilETK/weTck17DR/Q
dQp0kQSXFilStMPFVjM8X+atT//YnULPIKl7JLqtf0mBVoC2D6uRA9zYayBMHUYAgHCF+oVFl2vL
EQMfaTQ5oCEL/uK6mKyP4Cajr43WmKgDobolEYD8k7gaf5dNeWsPNJ0f5glwvpCqkxbhBOowJE5+
54xpF+ZvpFR8ihysKbq0Klug4uRccMMHvAvziUD7ZMPVBPVzjeMf5OTuSIlHOmvVRsQW3QzEly3P
7RJKAVwp5huSmdsri/cFinn1BsOMULSIkjjZ+cw3VTLa4Bg4DNpg0OXmtJPIK1aGK2iUq4R2ymUO
N7If2pIuooV+bNdKKbODtHIPxcr2whGj2yyKbFs1PPdfjLZ/RdaflmuyKjjm6jGPuXIw4YWw4C/q
hLxKiY3PDnEaFy8x4KqeIFsYlllMGFmJcNXASVN+is21fgOpZYpGcHHYLL5WPA3gW1inloi2+VFt
FWrcplb35dZYIdBSQrYlTibhLi7FNYPSxjkdT+8L4V7ouO93Huxwk0RmErtHWKLan8EqmvZGJ/wr
lHOJrbUnsZPyIsG/zbYF1G1DO/E5qWGPOOD9RZv0Qv4bjB1msu37ctZ6aYALDraFSJvJi/7slf0D
Aq1qYyjHU577a9urA8/dFOAI2d9VxH0/Oex0t33MAG67pfqpXsnSOBFo9aQuPe5PR88nPOsXlepQ
y6FqEYWZCcLpz5Qwo6CP3Q5gVv0ToHJAP0T0Zs/p8+irINa427B+mxm+uv6Zj7ERW5rVEjxIbUqM
ztNqLk5iqk6d6kFXw+m+3h+kKI5mUt2J76jYRP/vzHRWVigDKF/G9bwyRqBaFoUzi1OJN4qWS201
uiVbOHYS6Ziv++A2RK4u0Xy007jYTfIie1m9SU1K6DnHfE+n6j/h0Oi6vABsVwHsawXMLHsMckCN
6xYINjmYP1N5Vd/D6iYHINU/ZJ3/Ha5yJLQZQr+7iJFkXdbUArmqj7d8cHQ3YS8KoRSGLpBBjQds
cnUY2NzPC2/GoIoWE1wNs7Ln8SVQ81a+k3ungNCmMRstNzmxzAdP381QkdCTIFhaSYJwP2614PGE
Ll4HEGWCJZxOQj4IFxduTJjaS+dVg/C8iyyj5E8UpaBKA5qwHoiuqO0rLDjq9tKrye4OQzqh3m7k
EF3OZnwKXYExqsw+gaxWqvGRvnMLVHpdz2vF9Ea+rQKePYwQwmrfS5GaRR8QljSBNKiQktIVhXgs
ngY71LXOFNWLew7n0SCThujSAhVpQRXZraawaeWtawImZBqUDVrTaZ+QDGiO/lyorR89LqRZGkFF
fHsgarSNpICD5TASIZD87bCo2fahdCJ/1EBy6REsOlxTYv9wa595UuKgoSH51G8C/5v+jhGNNbrW
P8wgVb/sIwvjSvAwGfnDHZK1g0F3q5GRKMOGgM16gmFG7nF5TSUEqHBXwbOOFzAIkMXt3xA258Nx
LG5cbG8MLFxAwDoqbQu3xo2qzZJxX3YUDe4WjFY5Bfu3BfAngELKNaa8wUjSKAfkWDvtESAsML+t
438bwgUfYg42BlhWWhyi+iDmWBX+nkHT5QIpP+61zCIr7o3BR8jbu9K73xKJ5cgkNXZSZaeIjxT1
SiyVam0P2Ml7kZczKcEmMWcEFKUnjx+vYGGZufpzeIFLl627GTOc5Y/wHOvB4mm897EOnOZeZ3br
sG5zN3bA4uTq/ieKdTxUX0LL1ITkD9H5eiHJWeXbYDwXizOri8OpIq4cdw1PHEzMiTKaYLN8TCq3
9BIziFOioLV4TDxhOIudtCoflBDLQMsF0Oac4oIr2jXHBKaVN9W9VprOL1ZjpZiY9FYBVpguosZ+
UYuBW675gcOb93bhPAHVigv/gKmSVZrT1rNRSZQRslEy6d4E9PHxD7mKPM0CXfUzPkmgfffmzCRL
zBNzO52JYks8qMr2dwD0tRM93/3GEGFT56oyYg9IU+/Yte0y4XVZsn28UjQHOTlKsByOqzq59w8J
CZ4N+XUa9WL9z29ZfM9U4OTzd+7aBV7KNeMqtnN0wFI9Rq2me+JpTzLPVgq25DpLOZxv/sFFhmyU
hJehyyzFKbIfgFwPvWQs86r6QLTgJrOrRH6jNwKDkLG4KZ3CVyc+ejmZ9m18H/EhAdZZqoesb6E6
mryCzKxiL38KGX1tZbCHSfpo9jS6hC7+feYje0POA30XJKUQzWu4Mt5T9Lh7+oSdXbRyIJD0pqpi
5bm6DLHqKhzgIpq0MPAsQdTykJJdXLCXaGOxQAM6QcSYgZJk99+1pw8o2an3VVIqRjDyAjmK3YWe
hr5Dwu9J4ttyuSVREWhXWcrgGypfEC1e7f6z6sEEK8gA65TqQR5Ih03GXdluoFugv4VfHwcRkw2B
r63FINPO2rkY7he7GgkFNmFEa3grod+s6eo6SnTH5zQSbqh6OKGbrYzx50pl+dw247NarESlFn5K
1Sk4JaCMoEfxInqKHjuiV16GlqqX67m7lh+ZhsqKknASoMAQlc31M7/jQdWLnCXScqLyYaZDSALf
cjIkIpXEgePXduJ1/T80qgiG8PlGTx10BUkWlgPlZMlgqPydDVPmDIOwX3LMeF6kDXjSSKrVTy0+
YU7IEHcCMNiDwkB5DdrrJ4zJPQTEcgVlofGgl1GZZaNOonFoG67t4JRQtCQCh2p6fQX1Bjuh6UTq
gigJRZy4QlFnTUVJ7Lz2Asr8Y2HS730Ihprpok6+i23PA2wRSEW6i4WH4z+SLzb+uxXLtLnoorxY
yHYwyr7DvbH1JNIx3vv+AG1N2DidDMkosp9mRVMdCZYz66t6nYjSjnrtUS1zLb91WPOinFhOHWdD
d2J4retZfMbHMGAsU0W6BoFJowkmXqF70LIVL31qGDnU2okgDTnGXNgeLw6NFsQRzsQ0tLyuMJQj
va8OZs0fv75WZ7L+UzfEUQii1aQRbEJ2GpK0cuBr74mHqVfCb4ML8EoWWPwJGG9NtUcD3izBsWq7
aPa9LdU9p8+N9U3E95akt1Q9rZTZOj1fNCJx3r/hnA2GR40PpoV84qDJCEvXSXrUvZHBGT4NalRA
XE4kq/kXB13J5FClFHye70EU9P+v5OfxTHhcsxx57+TubKz/00zMqXwBizmcBJtMNNX4SCE0m/eE
Ick5mc6Nw2hkLz4/6eGDyagEvLTbqpgdEIun+SXVfZaq3LZcnE6qPCX5WnVoXKWCaC2uOef+0yaz
1TgjCiJsMXYyEqjhJLfOL3JTgzcVkHLUe8+/oym/KGVfT6VPQqvtYuLgDuerM+420EHIEiDuFnaP
2uJ1KEr/kKXsYypfV1oyjqe9dGoUoUKXGWWD+ihcjMT7zusZI/y8+DjhIgpFmkvFiicw89AuYbCZ
5oH0jRnHTF6Q1Q07fWFhiWoidwpznIfn2Qsm7Hj997BsHR9hlYr02LH5kNJh51yChR/QU0P+886r
OJ1hfTq3QV3Lz1aV1wKSrhvoBoFyo6hr31QaViR1rkXo/l/r+N95LWZNFV9VajfdXGq/HhoqEUHL
lZ2Agt2PLMCnFLI9e8YpXzQ/QJ0O56NXZ52gwR/MzSFZ0X6bitWwGpJx3bBGzMkBHSX4dI9mOHhO
dtxvH+w1jWf2WF/XaL3Dh9F3LN7VJUgRRvNmvSlWCbpwJHColVwUenxY3Yqt1IZpJuUdVgSyarxx
0AE0Knc170xvYkkATp/x+2S5kPchFkTvhszE4zBZtz+egj/0yWY3qeKkSgDkM/S3B2IryTLQWrvR
FEo5Ner7B5EVhz/I1xstUErgOv8foGTaJ5rJiCDKjy9WJ7SLJQ/gv7F31e6xXyJj1bk/1x/gQ/J+
OS5alL/lMl5hY6e/KP5YCDDfQTCBYe7ZHCltxTHpXqTj4GDR4NK2zax6rJy8P+Dgr3t5nsf3w22M
W4zC7B28zY4Z8Ank9tdxHNEQTA7pNIA/A2lk5plF7eESgkxvnB5Je3j1UKwLLBM1+/fGYH+XFiyi
T1Ndr0i5ltSu3DcdB6GOi/2F9FSWv9soNWNL2E3AaHJGM+C7cRbM/ZvCJf+2bozgQn4cyttZ0B0B
0ktlW2n/r33++Z+Oq6DzwRA/D7VGLIXxZUsh0u4Zv/vVR4qXiokHuS0xXJZ7/moyydy385IaEYbr
dozzb3D9O08CqPBneZQF5hVKcuEa4XjgA8WzxC1+BmPcEyO38P1epwSnVjc4OjAc9iUUiwyeiUkn
09j5KboyAfE8gwoJBWC4Six3roWznvYKAVNTj//rbk9Q4AntEXJbS7ZQVNAX/b4bkyvf6I215XN/
b8bqOu1JtljQVMssNVWAO3wKPNCjEOMSaPPe+AxkEY3rUTE3J73Z8HCBHiJwgWNLbrX/DL5QvmiN
+olklVJGOtEX8OYbgwY7Nbq0H59rFE5synv3a9sapGsEBSAMNqLuQlJw3t7xkoVYzdAdh3Knxwqo
4hDGEEczMqqVZNFef/1HsigBTLUP1NG+q7HflQdlDJmQFYpbxz7UEWMyQSzY9S1E67s93t907G+J
mjuSLqI3qCD+wC8SO6ZGfV3c4iEzWx3SFQBla5QFRgpGul6d7RyvZKNIm/Uzb9RCAsOfxYMeOCoX
tzJX+QC657H/iWj4/Pwq/NG9d4zQWU1AcwlN1jfQ9oWzCbi9GIPI6+VCagg5wsKdtWuS1UuEy/bQ
IbOE4AAGYIZ+5trZeQc8y84iW+Jl+JqiLDlZpnsBOc1AeShpxVsYZWZhsI4YCAYmq0l1uk6Yqshl
mgmVyMj83kSzQ6B+fGG3tZqQL9Z2znYmQdDLd6Rbn4wGW59UZ6OhyowIjqqdVISJnYgH6U9WKiVy
XEDKiRHi3WVOONiZ5CYSrMQmv1TLcFRG3+zNStBkoAcxknYA0oRjRtokN89Z1g5UZcUhjs/Og8uu
vpyaz5CcGe62tu+FtuwM2fW0yJAD3ieI4GaC8bxkmVT9rAivBr9c/4gsCr3qx8zwDGQxOGEOEhDZ
rWQGHk73wof+C+VdgxElCQN/RWyFUbe0HCdstyScpcg38w2QnjLCYIbSiVJWW2xsty4LCuMAJxyb
dw49o4KCTPcN9Q0sBzdq9C6nhfULGuYgpWR4KINo3S1QR/leC0lVAxvgDtDYNdoXvx391RhjYEov
wtrnzIQYZujWw6XWOVWDAAwveKWXOR+wPj7tohLxrTysyg+HyrpmI7ofCX3IC8NHJFns0X3J3brq
8aZTKitoFwLQr+GDXO0DgnsiZLazve69r3iBd1qLlpoqpR+kOK7z6QU0KEhDXotuvC8SEuQ52Dcr
cKYeNM7tjxk5jpTJPyWE67ssMerrTPWB84kH49ZuwfjOsK1AJIjc+EgNTVeKpqMx0+cU9MEfYUrs
lFNLkJBpFgDkJ7FJsgDRcbGTFhKEeB+o/E8DCsDzifiJxjt5cSPU5aYbiLxS0K+g4MBUvOZEihVX
d3g1DD4MmFKbgCIKZw0xrgD8exZX3RDCAUPLs8FxoOggErLvHq7wj4armLCYAsOky+daBxiOOLnD
1fLML+M7Ltvp4oUmUuJvFLOC6usQZdU7Vf0dloJzYjxHh6CtopIulh9lDdLG02/PK+cAuiRwEw0A
+gEaudB1t1/zSu7sKMX4bC2EH+y2e3LQMPgx3oCWDhytEzepqYSr/+49yT6qShCBA2Hmf3U5+4v/
hRUi+I8oISVILHkesaFjdZFdaVRaDNOWHCLR0TyshL4dqjlKtKwPLu52VE2Z3AKPXNxaaGCk4x8M
eGYDsfyFMOBBzDgG2UJY+ltB7sj23wII2pISft7D6JXyOevvTXT0VEVnx8YMn4eb20MNdJVOlYXp
7i2hf5ucg4lb0ThTPpcY0AvHq+9u+5HRx0X6d7gMCzuL90AtQ/yrJlHwORnbOp5yJF4ui2RuQACR
0UUijnyYev3TtDMG+O6tlz4RUeqwoyCnZ3WHRKZGMj9dVBtXW3kg8hmnpfW3dUCWnvPfVFq6jQJY
wzolEaEMAE2cy8pmAkK8m1ZpjhlDvp2z6j3mDChKXmQIuEmY1bn1AOC+A4jxw+JtYhCULkQpsBHi
oq6PSnc/Ci0tzMOCA09y0IkyL6y+j62g0bVixp6ih7L853pI3KrzplElTkgPIfIy9wP7MvtO3T+s
AR1sflZW4vEJakmoUrWy/jS2wk0tcsaosojSms9ZFnEuJdUwIS6pHT5U3CsHjyCPvIEhDFoGay4+
7z+1jl91YvfWnMGPX+bardcJM8QXqTmwq1g8n7H6fHrwQ7j1pROaLrQnd+Cqn05xa9KLhS1QcQEp
IMiAcEiWewJySqtUuHgMla8I8N+gtn1/dtTRefqaauEe8c9UhW0hYfX36/d3BTKzgjy5dNYUfjZ4
lMRR0041yIxJWV/lqBt8HRPTQapYs6L7z+J/HFhWYFTcRR+mOWT1sh5C6IvGdrrkhrf6E0pWGZcI
KbWXiGtaTDzOC3KWPW8hzjR32g2T4xbSoyeMSGSF3hlW9gZhUbhbE//PcaHbvWXMfjOPaJDjoqA9
mjG6x55dMPzQc0O/+A/XJ3T/kucc79qcBirT3ZZBv+IWKYOyoMelaUt0OFLaF0a9lQKla4IkFwgg
S0xW7AveRwSlfZCahaDb67xubrOYdE74cBDoa7gKH8NUUsQqNKSz394SbR94mYdXGhCkcxB3HQ2V
RP0mRKEPBKGyDF2yIVU6HZPaVSlcYvU6738UAAVlMJ1R1mgE6cpBSSAR7QWD5X96w4UjpHixzsMP
bselYU2aWnFygOi45B8mU0dNHmV3NdXUlfzxCBeTfXwjZJMYjih4hiVRac1x9/p8GDTAvXD7eMTm
+mAftT+dAiSf6X4ajGiZPxFP3wY8mDdpxkCmGoGhzMvu9b7DmDjIpgyX4tHjcibAMf1CZJk03N+5
kZO/xApt8fOFACibQ/WdsAFolYPiboMLJX0ayqGMiFjh1NT9JGoRFXRuUUN0nLwd7CjiZ6mVZ83j
3cBirj6bnucZIxN9uRU/LrtL40LFWllb6FxXW/dTtCvzT6U51qfUYA3lE6qiWP3zWVTNVoVk+tc4
cxOCXpfLDPgrDhBWyVZlTdjoFayY+aliOCq7AyuDxkFDHjCNV3joFe0Zgyzdgz5WEE6EViTTx4cP
iR7B9KA5KTS5kzEc1NHBOBdIrEeZBKHUIuARN+LxdyjU3kKhqEXUDhd1ez8xqJBzzzMoxO8o10Fi
MWuwKcb4Zl0Ei8nbe2PPJsGFvO5qdqRRii1sd6ErB/joUUv8D8AqIwMkDGOvKrtsrladk4Nz4T9h
/W1lVlKuH/ImKeVEO0nZsLyVgYfP5ECYVnYcSoah/SmvQhe/WUpPv6z2Wjl4X4Mgs36g9mFKNqIv
XB61u7NNq5dOSDO+4T4P/0JsFrmSznBeBCjWTwaJtp1zdB2slZJCPU34+m0s6qwC/lN9Fq3LssI8
o/dQ99xeZTd+zw6Ppqyr3tCYkFdaglYzy+cc0NMt5XRAzqIbn66RLqV0dlhUd0ZUj8t924QmK+tE
LVuyUbk0TXwXWk5WXs7Uvsh4rzKN2gpI+PGFT3JuNLCJatxDKIvMO9BdSIDEON0W/yb7WquqoS4f
oAg/Rffb9SVlCdgEKG+XmDaoek+xamV7inL4A+jSVzbx7Y4Tnj9LNMV5B2Ere1pIW7KQDOGJZURP
lY7Kxo6P6wJM4PqrnCwxt4+e5rtfcuMS5uHw6CSYqO5UpraCTQsrO3MjYEgEeECw56xU6GC8+dOB
ASSE3qmG6zAWAIRvuqoCZj9a/m6WOhm4e24JbX1FG430s4Zz/9GpvW2GhGp9Zym1fhSMv+GhX5vu
bpG/tTx7R4gUGgTgz1MRWdQdH/ssJhfF+COCfHV/TBm93+Q8yk1ocEnOfmkpaZkKqlt6pIcUTiFr
1MEYNkOitd2P4hBJrrfdpFRAqwYIH/Kke/Wf871YLL+hrVmP6E8C+wEPx1HZw5GnZPFQ7c8TkfFu
TYUbQ4H8Ymyku9p96P35TQ34V3iG4k44Zq1dOMXZt2BGeestxjWnDmgZP6hnyH92EKDP+2+4XIqI
9fR5Fq/iDc1Dt2VHHYealrq39HbKJM+YK0xoxXH1UKwzI0mx+VMNgRXM3dEdkL/qsqlCR/59LIXm
TiAxB5FGXuOdCk2YNBM4vwkUoc89muNjC5/8ctk9iKhoGjVIqd6+ljO8a4MvN7NRqgPCb8zR5156
LZs09ZdRg9AoQzZgbulE4RQk6SLxw51zI/th8+kQ1lFkqHLBr39vFEiimATQx6yejZpu8Hd7txtP
ZotlW5R9QKY8YntIrUa1fz4QgX34xK9DNkCb1KVLxRySCrcMNUcVoXZ59f0oXyhNDCTZCyfybTJQ
ZtuxgLgdIwrdIkH2R2ddr8VBVXoCoWJuvOHznP1c9U64I1cMNofIbo9I3k3jiJohjnbWTOb3eNdz
pR8GcqIqERwHxh8ZOWwMMwUXP5d4f//PAzTmqbsVojDg82Xu+dzz3BSI3Fx0D2PBy45SmVbeusrG
Cfq3p5bxvW6AMPIqpYJanfNa38FYRn952jBXCawC2V078P2w9q+AowxIwj2aoabcM/5pZHQUWyuF
sPiBClhVijsZf87vl1hYPeXBzQJFyA1Ur3INZL5B0mfUXN5b758KDmT/WFOjIJHsf9cpcQBct68s
RZ7TblQP7TSduR4TWJY1XW6fIyDRsImgk4b21+rgDunT0x5Gaz5ZFCQ/Ok7UJBJmVqRdiw1oMuZp
sDVXq9Auckg+uK+kh3+OJM+ChxysL9260Py3sHlrjp/h/JLBnPIqAUvW84madO/B9gcIoBrltune
BQ7b29ORtI9c4MHsPi5szqOZK+CO8Ixtd5Z6TktKDuxqE85ISiw8BDcP7gIlX7h8q10QGDvsZsUO
pb55Qq7IFzS/gS4sapQbI3RsOt8BB/uGNv362aZDzuz2wlmaVu6jdrO48QyeOyI9/+0I1pJr/Cc6
4fjvKBEpPK13FM9wGY8BOOJhf4mMTB7XCPEbirPj0M2DGvaiquDeKMhCfVNZVb0GUuT/Avwb6fz+
fn4SJqJWHLWsm6gOwMhLpcxUDzq8B9ak75g/gNrB+ZrRO9NH1aDd9xGJiFx/JVHz37+jI6SeX9da
DeF+KDl88DMaVvd3qPJhvPq+nSjzudBdG+RWkON2e4NOZ1IiulOIjOZN8+QVF+p0sJizQT+WGLud
9BPW9nI7gfStgmpwGgd/FPT7f4ovf91hvqVDJ+72aqKrDAvhR8P1A6ujr9w1AycDmFtE0K66MibT
byyUVfwV9fC9k5foPfN/7sMogHNo2ZY9rlEvbQtQK0hAVWRWRoFivUTBY+5EY+xB3Fiu0n0L+YDm
hWLjNXTBFZbqswRL3hiC+vPY5wegzyZbgF9pfxz0xhIccK8jRI2nd8n9o/j6QtVjTgsXDyvshblk
TwGGUEOZsv2AZ70VeVIF7eJUk/ycjAif3EX33KM7HRvo4ptmeC1K4Rp6Ay7hiIupErsaLO+M4/33
GBp5tRTIdmAq0qUZEpqqYafz37cXA+wI7iRI9Hj1EDss1G0Zrou6pPRKJs5SxDbluamv48qI1CjJ
LyVrUrLVxTCjNZru48kn9RXewis+tlWxZgzCAb/vTXFHP+NsY4O5ReSRX2wryuAiKM4GBnkR3VW4
QSUSIBXESbwsfkG2eDTjKQXnoUdS8nE3AsfSi7PGZL7A8ksxGm5xm2qPnWfkm3yuSTN3JCpgPZm4
lqUaO987mvg0PT+oDPIJE3rsDT3XGWTVU4Kw1FnzsRJZwuyInftBNoQ2qrwCDaBDU5CaZkXWYMj1
lQQtYnJVchZbQfX35lqKRKqSzzOtUFW7yw5K/ZonVUVlD8AJFwONiSq9hwdZgN1bl98kRKfia3K6
kAwrI0rV19AOW/y9iumnVbiWJ0d0tN9gCMu3By4302y4zmnTEfviDFAV4eWiZNmco0Ci5BU492tw
yZABZ9M6XZiX5FC3dAw113PdDOh2doQj2NCMrGxFxb9d6sfy/LJzNbzilmBmmXCHZVKAwjg3mmvt
hc3f/FPlPli0duKVl+SD9PUbLJ9YYyUUR/igjq/is6///B5ImJ1hp2c46qgj3DKXjxj5dn0w0Fe8
uj19Hyd6/C4C9t6UICQUEVTsbjpmWQV4Wvq1aQ1ttobWoSTTtK/RAIOd6rpiBCMAhVfSHWXTfk3s
VRAwa+13rbtiSOgz6TRZNbIuBr5lnDjgqNH6uC99adtBI6qx1nn3VaOFkrheAIuEnB3xJvE53VH+
ZkQVaJ6T5vpnsbTvGD34BxWAVLdAdJsBzKIFmNCGZSEHZpIQ0WoyX0x7d6ZZk4/mTqn5fKaH0qs0
TNnpHMBKWucYqP2HH2wACi8E6H3t+5B0KqaToSsQkdAgd3+M4Ev07VGKvCGL9id+lStOdsMQlUgI
NCg02qJP/86RSgqypn168J+UhH+pkgN6duJrF3gZF5NS09bzJO72r9QS7yFo/5QgsydMmnAZQmre
X2hJQO0k4z/O0m6Srt9rH+kYj7YuVY5C5KRn/OMvMwXIFn5SogHF2oh5vIRMaM1x+zoLtz1wmw6f
gp70NU63DP9zWHd2JEpYwseFOa/oAXKc8tBaYhhmb6Y8LRKWj5nxI3tYwfyWFUVWyeyEkmzWL3Py
6+t9cD3Y8OR+5FfTxEXilUKO2f1urN1IIfgeiT+ZzNke/oqgaeq3d+T5hCJ2cJWA8zH4TUJdFpqP
awn4Y7S9+xCI+ydH6Od6VFzlkX1n1ShRpBXOg3BU9Jw1pzljVJrfsrp41hd4/gQXeP/wgTY0DxxC
R/bglORz341lc7eHaKF3kaSXFRssluGVh6oMSRss6nmr9eUdmNal7Ta39+hnRzl3L+rAk3LRzPoW
XoEVJcLU/394qWVcXRYZbJ7rykQZuxxOBFwu7xPV/Q/6JGKxyuOSfYB8TOkEAbbGYQG37mJEN4FJ
i9un9jJfStLV7hmr2eGP1rj4aanYS/zWSsRy8pLP+0PrJ4LhSRPR/JjNZ8xxIJdWLu4UyhEpEy1u
kAI9JHUr8LDNPPXTVPz3F2cRaNGqduCbO7gwlMAzvDvvc1p0lB2OZ8zT+StuSmY2ON3AnYqRjKX3
2sasQBPFdfS0gudGhUXfhN7VutvruF+GWp1Ni2HVQk4p9rmQTuqL3oqecwTyQC8qjZVyIPyENW8g
IXsIc1zj0atOOghrh+QrsqkJ++qm92jXA4FLXybj35u4f9Xgeumsly+fQrGantRKjjhTDzIFc7a0
GD+C8mOcFLrr3nZRGPu62q+zCDWwDohdrNxUgOybU9bkBQAUvtzb1kVP8LsXrVYtzyNirhbD/WB5
khbmxXqwq7fqpiclt900ZWOELLSRLVErTzn2wEvJoXJTQ2sIfcJ6zQIH9v9xPtwmbmoX84SFEYMz
02gfC531nempdEUHs71hOgN2zq1vF299mW22LoydFK9vdSphLzOy9PlaonGF4zRJtNN5EUfe9JSJ
RZ38kfXbGZWN8lCdw470nJCKrlncLo+gFDgklCrpvJLuC+K6EkRUBh4tVLNuNlZkmuZdr8f3v5fC
6PMHn+vjhwtrjNfGap4bfjcIdhSvbn4Epszq1ecYJQkHNaZ747wLbSpmCKPtY/UHYRqHhnIPu1bW
EyHk6DqlgkP2jmNjhVD2THlFWo7xfJzkw6kfBziXASZ/z2lWwzgz/hzJrIUFb2+QOJ+IqKTR9TTl
woEILsYU+vRnfdcOM3UPXB/TGfVfzZmzlQhxnkD3ZaZ2vf01YVLXcwDNodIsToGeMVHdWe4aialv
rLRqGj4V+BXUU0gZXkbdG8Ods8u9p9aE8BKAyqWBzEil7R9FTVavTNl7Npx9yhWKO90L8XDVGCA6
hSzcIdk60AVWhhpS7rO7JbrKTfPW+OagMUHD4luBjDfZ8UEZRffuoM5TFMXlb3FUoqkhO121UqR/
Em5fg9fbn9IfEA3OSOJN4JB1ncvhoXCjMCkAVH/vR9YAxHv0FMiXacS5J+pzDi1A9uIyxTYcOzAk
2SvGUMKltQCECItSwa6md1iT5MZlZ1IAxi+G1VkS2Ter9ZtzTYcEq2wSGDaqT9VTri1bhQJNKnMP
o0aU8GgYlATdTOQxw3Timxn3gE2x3B+s2PY+u544gAXYkrUPh73YS+ScpZgLp/Imf2LyEIBKLmm+
DFMPc8k1mgyseXmw0Eox+mJvGSjEH1VotyrCc/+uQGW0vqg14tgMjrjoYX3KNLqBjOgBoPDDB7IV
zh2jPXnLU78fSdy/PjI3PxIR3DBHdq6v3Co0jrJBxdX8q/W/YHNUwK3Dh6FK1DFQgk0pK4Bqzrg7
4RdWURH8rAA0eruom81I9yRvSJYvGE7x4GpJCSa2xVcAO4HWu+uO3muc5mD9LSh+xKNqednR5JUR
JcxrSKK/OsdnyrnCL9HiFmdAfXHeDM0KFodOgODAMGs6VHJ6fchTyVL2rC03l5CU35AyXYh3fAz3
bUkwemDJvJcKqJVcdNrJOZhANzykSZL/poVtf3rPBQvQ45lCI7Ju/nSQH27g7tjHjpXlcgVCkKHZ
7lnG4E0lhmQ6zBh4BjxiJJVU5RhO1GiaDq8n3Vb+DaF7mEx47bZY6QRJwnEmzd5FpCHxk/kiCROd
hoIw+6J81GIh2pkXvnoNZ2nFQLq+BukqAh+snhuVH6wQK1N2nEQW/sPRySjD0u+6xxFIb5oKz790
YcgC8jDMEYlhq4vOviTd14YF8/20S8Qnm/iQFCGFunV21+JoFvRrVjbU3pMvCYxxubSn/D1ff7nr
wocG+/SWkF7bNOrdSg36KCkph+in3/wgcz0ufR9vyKHhb8Z/+4w8Yenby+LDucHLcbhx79gdR+8s
bI+QNt6tgrOZauT+AstCGoWNtMw0sV1hExM6KU+ZoXOm0g8BMBbs/LhgvNJVwrMai4YXCyXtCLWv
QwyOLM+eeNLJ309zrOWTtUWEuJUbALDj6Fl6TW7OG7hBM2uWYClDJwDqR8Pzy150KVKPFDk0IvWf
bwieJ4IMYxO6GwRwVjJBx/B39VOXHYpohtoCBEPXYF342eeEuHPwf6xZqMmmVTV/PqIoZ+LV64rV
Ze93GmcexP5cdNvF2fZsByl1aDoN5tAGAHkSGBbShvlzP8kQUW/KylvdonCvooh1oFuySNUvdMMT
/+YsHVqEOfeZ1BhN+FvSWeLEcJ42ap9YkODtaaw9jyM1YTerpG3r1fg4fVaatT3x79GVBHHAf+ip
KohK5ngcYkuqkZigQT9QHHpxaXInJSE5SrsMC6FrlVbeRm6Bz3OncHFATwPny5qzcpUwGT2+oytP
63U8CSBkjYPOA/kVcopE1Nm9XvWaN+hog1sUS+vmAcN+Pf2vkwf3WIxRxUTe3EWIVy8SCNRmitWz
zsy/EQuvcso4aySrk2CSgeuIZObwTeKCcM7b+qNQLZzirZg3abyu5cTNAg75Um/PGlw4MiWnZA/k
mkWdhtjonp/Mq+VQreMYXZ/DLiDwBpKAFoxEPYLMfaxNURrLInCzvvddBz/19N7bzOs4n5nsuKwj
JOKEOQYqfe/xFfxc8aAqwjSxINEyV8YqSnrFtBDRW/wpTWUCUGgwEu1kDZVIasZif8j6bu617Owi
hGZk5OBwzx1ipHCOdFG0uyw/y5Un54b6qjrlfYvdKsEjuzwrjJaB/JcwawHTw4/CSi9UoAzPYJo0
aRQGoBdsVpKyT61678FuuLrYulX5fnilbZ2tFnY2K2655Vu268tENwacLStZs+5p3r3i7Ait2xha
alJpe1ftJ6oJTNFyya3/pBGCvJUM9EGNJqrtRy4ijXJZAC6CICrLCugcwx3i1DTD/VpAk9ssrVIi
DQJy87Ilbn1tW8vHSEvbth7DqbEasHBLBCBPE69s+Bf4vM3QRfhmmKBJrfeN5Xrsl0lVPfaye9Z+
yqV7mti0vRqGquPu86TBVaS2y63cfUeu8w9PdJhvoa4XuDLLLjnuklEoH3ED1zOPoBj3IfaVKseX
jMopF1fD/er66SbBIvmeqGqWsq8Gqf/v7vb6wz1xLb7hERoleqx5/xGH4+AxHY/6EViWKvAacHDF
i2xP79DLhVnY4wB8XyxK/hyV3oeXulgm1REA6V0x/xI8UFSiRUATIiz+p5oLJHZc79e1+noJ5zfe
0sWBmccuytk/HcARYMAY4OokQg5s0JarBKfa2DwTpajx/6ElRh/vDKNseEJkH0wefq5wx1ajN/fZ
A8HgDk2wtTD6ezPGq94vgnIzigMlvQrvWpOAyMMnW4VKqiiEveFwuHX3RIWPyNlyUJ18JGHDYrmx
ToIoQIH8RSYRd66LXt5CpxzT8UFWROem6paqxfG42tMtHq98XmIsmndYQC3x1bQISBxxl9pQhxCj
ol8dE/Lb5qAOB3MRiZSzAJqn4RJm1HP0Q7te1VoZ75+4Phg9uOlVCfusP8itSren57AIJ5kkZ3x/
3OccYuxQbztUResgk7g0YOq6I7qcOkS6bR81RHNa2vpkzCO/3SKDnPnCgO3RJBeQENMANu4Cw2g0
Dv5pZVUXxjbw4wrh8sBk5/JLdKWOebwiPt3FRM4ycIWBt4p3t5sbgTAyMR5lBlTC5gmKvg1VfBwl
1cZYzVdWhV0SuFI5Hg6WTiKbjWesVZsp5nfU0R2kZaJwl00bsD+8JlXVjl4GHj3WeSepzk0dXWfZ
ce+z52balC16PIoI0As6pPAPgbjkyna9141zL5nvRLRe+jn01rGmKiHP8N4I/renAgpAfuPw+16+
MwcBFvAt0CaZeJRhT6orIFCaCuUCNq3dmO+qoufvdiYl6RiHKIiU3ljXCoYP5o46zbnxlCSDRzHF
tGHYHhocPXKZvieVvywxS7VsHX7foWzUCFmph89jcBjim985ykmiF+WIhM0DZhUIICiREDw4nDLl
RYDyPu5UgUIAvLlzx2RR0qMQbrfeICV0EsAGnK0oETe4r+3YeRg0W6RzG+bGKKThGFioeOVcejMt
5r346QfG44qDkC30toG/J/2Ue6N6CsgabnBwrNcOet8btdRSZML+NhgK4PizmvSFkoNF/U0aQXIj
aEzK80kxEhNBLa4P1HlcxjvD9BxcPaB2cleCfm4adrtbl52W9Wgq/Y/3dXWEHt0QBz3iF+FN+ygI
2dfvcKICSDiyshW7dkDxkchqhowb0nBd/+O+bPd1x76fZ5PxQiaR0BafjLTyvpFjpasBMyw2NOAv
yyz8mesNV0dOmV0OyMqP7gKqCIhmXeOYEAtiJCd0d1rdcDoq+SwzuNrAsPVfbSV9a2mSANiMaDGe
rioKeNtcFVCecwiSHmnqy3yid7FbD+/gen6baQ5yAUhKqtQmu7BLAvClphG/EOhH2XogaP48kEDt
uaojU28dt4ScY0wpxSVpEu+plc3MDu7XtOLkO7HmQadzfXxQ+6XG7EHEwBhxB+Z+Z6C1dwVxxfY3
GbKyyRClvCDyEv4fvNssx/UH5UP3Plogrg10NWc9WyQeb5LZkFqQgnP7zTwV/vubQGXEBNz1lL7w
LZw+Ix+pFH45tDqqJ9xcA4X9tjFMN6YAqNGmK7jSTZfvSQE9MHSXp9hHL8Hu9HrWovUpDM4W1dYq
PTd8fBrXTTbnSKWBHoCXlcA9+733ZMm8irxMyF8emduh2c+BHPSBV/vzIhWRN1ChbTRoj8mUkqIs
c0jhBB7PT3i/twF/uL9uzSh9nyLJRjBErB+Vv6Wu0ZNAUFDlGbPX+5BgAidFFTkPlV1r8+OuDfmo
QTchDV/Hvga44zJvXUyHh6g1mFEymyfm16w6cl3VQzEze4eHFfp44yUCdl8lrJ0WS75Fix7MwBde
luQsYDLYcupyNn90vQ/PzapHsyc9Yt/GCRiG+TOjQwwyPoUONpyfya6iJQZvxyH+JFjAkOHHeuKR
TGAQMLGTWopI5bG1KC/i/hixIf/JBhaiqh9R6xQ/cKZWih+hFBWoMykO7pJlP+8tb6hv5zR6dT5o
iBFvIOlNmridOjTmgdsn3SvBnrp0u+BtwlvOLgCPNMBJIOF7zZ+MBccWqGpQ0sYd/bOGn0mUUyuY
qm28WwMZBKVs5qnvS+Iou9DyOfxoGfhY+5BH/eNyNMNwu4EDaNYOclfP28DK797B3SRemNfO2L4f
izAd5nETDAjn64//VJvRo8lC+aJ80kaGza8A8hqnQbD23XIWODFHyyk+lCWhFg0vzk7sWj4W+qlL
6LFS9+ODTbuzylvMEAq5gRvxwfuxjB95rbwNOy3xabclfVCovi9kUsGe5vzhMtLWglcBJWQtcdVK
7ZlwqZS7rASCL2kNr2w3JpN3FYbb4XohC2YtWAmo2BVcBwLG8Kt0YO42bXPAKoER/YsAnLWJwLkM
AZgWXS6EYSOy7g06Twje7RCQN4SVwX4YQA9J8g2ooelOIL54XLM7mL7c5UJU0AQe17hu4B1HFN+m
Sy0N1Uc4OhLjYAc/HlCerT1kPsCH+o6MrC9kGRqsgCurgcVWauf9CLKOVUzGPxlD65xf3er4EP4T
gKAb4W8AyaP1mrxpeiWqt9eCOlU0m5veCmp1c8jiRXKgaltJdCrVBKE0vLo58YjZg5DAvoTcodV8
A6fk9RSgd8YDrJQGRBl8MJettUJGIEtHENoyodenznBe5RA7fzaRmQDGyhqodQ5aGgAKb72bXors
3nO/35PJQFKkbFAAFfkAAjroHz4oepglVSdd3D5zj/Ms3BSwPv5xMWwQuPbGJ2aUEUdBiGZIeMgL
MEtDU8nYiHu9kUg+jk8ztHXKXmwRAMhI8xyOc9oBLH0Sgg38NTYp6pOHhbgQ9tOw7yRiOTBCcrnc
hfFyjpBaVD7gC0LSmXel+Ly9Exd1hVSwLDB631cvA1L8mgXSx8JXqy2f/lan3xc3oVc0lZSk/saH
ELOI/mQpxpDgTBsLIkO3TQ4ahtNxvdno+0A5PXuF6btGuXk+l6aiFLITvxHwaS0GVZCR8pzuWb1j
pFhG/IuamTb8sCZZGxIPFanQkY4KEtDuSBcE6YjafowiQ7BbEfgz0Yup6Rk+Fr1J/Hz18bHAZIGi
IAfY1VqzNeoGBySh4hguHS0vdMb3/ZnoZ+OqX6YbJY3th6hUmCmWu6mMM2IcaecxFiX+nqHy1TDo
5jP5KyvwxXD1UxWHp4WmWC8wKHm9QrR8sT7gzW8Yr25O8WnbjUA0sLZaakf8cMT2SsKaBoXazjWk
6/e9Opq/0W774KCFWebXKcSE8C6qOISJljWq+x5mOSxXJRhX5B6/YbEu3SYG067S5rtvY0SgrEur
Dtvsk7/XwQTWMnRzWeayCSFDbKztQlnIlaiAvTk2h9RngiavNPzUaFHZYfvz8FaRHk7eISYASgfo
MM1QY3LxHV93y8d2duE0WE0v3mQ3/pK+tJpcSzH43NczscpfPzLhesdXNEIaY09KCf/tSJWuiV+n
PPC4mrfBdFBJqCvOkULVoWc4S2BdtRrHO/3wUXFHlWPhZd2MiSBgAvfmFtHnRiI2IMxunxEPXQwX
u9iwNSSFEk24J6B4QzhCnaUYIXeCnVqfRfgpSbMYY7G1PvzDr5CFga7vWNB5PbkIUdMSHoF144fn
IzYt9+BuS2hDhnN+Mec3SJ9lAqyL6ZeOfUNmY71m/44b5GmJfRi8Nl+75oLJ+UKLEjsOaivnR/hi
f5RZBtdsQU3dd+jC00Mhq04LMBBcoV3CZQADzEDMoo4eIi5knS0Jshb3yHtZHReUfD5Gn+if3f7p
ShKrL9ynEBnuIGre4BzHLlUNJIT4qYdqY2/Lik4ssL5rrk4Tk8lxKElFEfprgw3m+oIyOyM3jKbi
0hpen/E4dvGft5RyPOCpm+PPv9eV86a3mSn54spDI57CdbHSRk7KMjRVS7FGWWyHCjNryPOv0Gev
T5BGS3mgze8FXQIhE2uTa8o/5v6gJZoDoJ2IyID6cnXNwxYCM58t082XMYvcXOnxJxfPqhg3GCDB
P0KIqUENBLWPTGLUGcZgGWrJgXEcgIQsPHJFRHPJ7bhot5QIDXSTtgYyjspTTzM0belVuVswshtG
exmhSsASn8CSXvtFe5ebf1gKf3M/IU63CPvnhqT0et+P9JcZudBMmD8ERkxDYEFNCXdNEcNCYiO9
eHeEtVn19nO5AR6c/kuo6N0GVPfPUEy/xaLP7Ya6Zhb1UiWCegv5zgkPcfBmJ76+VgB1eUTefbe8
2003Rm9lIQZHhVYPJbWa1TX/4gQU1FuHNCbPzqZQcu2QtdbegFG8/ipNer5XnZoAnPLRyp+lBLMk
6a8KYf2DGcM3zKUpn2oWF/iJV+tUcl6LRFf1ICd/dPA/15RkYNvL82kNw1+NNqMQU6QaRzRy1U2/
30kjRvbdyY1/hdRWbg17gU04lbH7Jgfwv6YOoo/Up2fOlDPz+wiJsF0sa/vdu8pjS0J7NiJYnAJ4
aRh2Epsh99IY6BtKTeKWJN7DIucyZBHykgQ+uRSbUtOYRR3OaV7CyZTkhjU8T2OXX7fAsZ9e/lPa
tYU/3/gyXLpGs/Q2USia8pFG7ehM4Do8v7aAfoPL+rj9nXxwgzmCydwhdAny3gGHZJ3pdBN9Asx3
/IqOgMyAqtf9t05Q4ik1XSP27FyLBMIhwLPUkxNnk8NACkW0nfdIgU5i9SsZG1iMFj6leSfka8uE
LEjhZ939ld5QMvchHmrMFkYUedjRcrh5XE8K/l1KFbAFvekDCK1xVUZnAz9ChErymUaDa26H82he
H+SFCFXw4Y0JuDuwsvYqkODCg1LsbWrBCyHIE9cz8I6FdH7lqBNhfPnBCvGk8Qqr8BzZnRE1pdQd
Q/2stCXY3LIPlrGytOTsccLCHl688W5QYD0sag6fGRobtg+g3WHLdSnEIj4nZQwvVytDcA+mUzLb
9VkzZ8/JUH0pfDyHY9kMzB+ApPYZGSvEEuRrySpCcBVj84aCISxgRGfreU8EcFQfp9nxL+Xd8cB/
YbKnN0Cn5bJpC/gcVsNb/fjeGjk5fmCMv0RuD0PMFDf703T+Jeu0TWotdkmoziZuh3ydHqNuyz3P
klpwkQo6mVyFZzwrVexuZXfhIqbVy2mZ8kh8hyqrroQCj7AUrITCXei3df25nH1/bjyRI6rNmbPX
oMSGpX3Ko3335tjh0Ez1jvnF9MWNGLrn+BOlz+EGi6vI+TL5jO+275kNBReZHzLtKDoieXUqbGHN
K8cx7tdAHDZFwWqAXgR5xj33bfzYE2EjOpLkMlhhtM7VAlYf8UWqMd1RI0oLjXo/bEnkOA3M+B4h
pLsUGmQlv+V29hRHdhdPIOX1ia4kBirS2m/TjoGvQpnROdjIW606KEPn8rcgB1nTu9zANa9abw3w
n25e2vxY3deJPYOjxd3P6yn1Mn0CPsDFTWEFMnjh23fDGsTJ+WQnvM5qJEvvH2ZI0RkIVCqzAgBY
IbyEYS2mWiHwTcCSU5vrI2EPSBfFvZyaRdJnv2TWpjvsiHfT3xbwinPSwFW9fG0oaTz3Nd83/kM8
36x/1mvZmm8tWevt6XCBB05o8w3TvAU56q31HNbuOPnYxR7dZJ7Hf39IqgYaP0un7YCtzl7EsOfM
Coyhtc82lIZ+IIUA1sSC83M+1ohBxGtjCZEAwbK8Kc3NKkoptxurhwx5KoSP0puQaZl+m67+42aw
6YaKfH+b+qdNk6m8lMsvwKNeox8Z00nx7I/1l36JmRCdFE4lHYSo8JYP3jQv6Y8FanqEGhTExR3K
2YGNhCVz8ldKcQcOm9Qz0JADU8pnIBZElAu+TaTUubdU+2IBnjQ/it752yMew4BzOcaW7zi4omxu
3Ye2eGh7WXRC7iox0wM1fnol8Nz3DYtU9WBax6XXFKufbf3qux9TcdboI30A4+cG8KA1J9BJlECG
B3ZBo1DJiPas+aEQjiYecpR9/WrnjqFZcTldVHQWZSsIOHpxEFpthGhLUDLvJnDmHvOtiLtvOU8C
VyVmB1lRztRjdt2C628Rc2O4Ua3/sn3EjcKulbgFPr73fcm8cWgW9Q9TWiRBh0JS7dT4djQlf+l9
EXsvZz3l+Kfn7SazOtH0iamWZzEWdUPtX7xputP5+TSiZu4q9klSW84d0olUdPYunSM1c2z5uBHl
/qbPNNmPCcpzKYbP1qe+S7pDIxT4WH4i3Xq3niF6LDHh6N9++s15jdoDNCNAh6NCbBw2YRABRZuU
SDl911hjGRx+i9esU3u2Fel4xWwSg4XVqOl0xWOgCS4YC4Jh0HFBRj5vMv7k4IXgKXT145ag6cdm
/Mnf8nnAxt7vkbrHJw79gyGKbdoS8LHn13+H60foLo/7u1zahE3QWM8PlimcAexEhM+uZsdHLYTC
a3Sw4SGyzORGhyYn9O4lxPWymgKCmpGhEb/VmF6VhFfvjuKruEJlDgSIA5us4rZHuv1uwlrYPCxK
SEXGihYJwnDieHUbQKqfUzioeaysbKPZ+9TdlnTBLeIaclF7qNySbg1G7edzsagziq1anlZz8vsf
wveeO8awIrX3pgxptImtqdR5msEm7Mye/THI78L1umO+85QdCatmfkN1+W4tPRtKPCbaMhT3PSut
ZLRCtSLkQAhV1oJqNp5D9GNueOlkfQ0/bdX0Wh2QziROQDAW6uerDPrMcEV2S8gOf6hSTc2DfAyI
Y7RTXDUv8LUn7NBTv7R1LLsu5RI17tCBji6hwTUwpVAwrz1LCHSbui11dj0w3RXNR3Q9ruM6NKMe
gR+qN1gQlqvkwifiuHGq98lo19M506kVWZx5PGoE6fYq/8ECuyxD5EAnQ20g3ku0XJCwRb5ZjlhR
AIfxis1/9mS+1Sc0ZyF+GeDrywtB5Zdt5GN545dpi8aQhQHdBRNglibI3/vxV9G6tOr1d47wNg5v
YN+niwgCoH6Zvso5ysQ7IENQoiUFmQ8c8+BG/CZl/OM0vICgebpe6ajCb4qFbg4pmxYKkIEVizxb
WQqTJ/6pqTR7PuhXlFtoFjXHkLW8fvQDMFA3SsevgRpp2/iXC19UkcxaB/ZnPsYZeg7P8mDneKgF
gTTSlnILUCETm4UmCkBa57IlLC81tvUU2YBpI/rUCxDHyjhclRIKJWybhtID9axlmsxr1L1hMFdU
kgH0Kss4bms5OWKrLIWI/78iNKg7DlK3K1fldBAg/pOfwJbKlA3eoCKIdo+3d6WoLvhy1u8RtxMQ
fGT9I/C4ADisV5oF8ansxIZw/feqKyCqaus2dNFUF6asblJrVS8jmPEg1keupIdPmgJnTO/F2DKX
m+9iF1k7gF6X2h/mENCTIaMgH0GWSmyhD5iVGHJCUQKKCJJb8ZqlVXlLFa+CIvtNHRx+ovq4XAU3
bKqOpD6Anx4jMh0LbfUfvqU/B3/hSIGSFZpHBsCOAnsW/QbN/u7LtIiMimPvciTSjIwDe0pmo6uO
yqGvT5fgB6+qUXYT05AJYGYq9X5/zHt5oz/AECow6sZ3j6g8KwUcY1n6sC1jM9zrkfNdUaCcnVxv
vQ/tQ78X+BwA1IDoDlEGaOqmOiPNkkIGMlz7tDgZA6L5B8hjbi1X0ZWdTUcWclIBUID/rLvUGJEs
GbiFSs0LFRsTk2SWj/RQ8KWHNZYi2guVhbDwxnxcTxCPtd2GPVsN6VjQnyYIaIeThFodaeV7uf4N
j2/SPI9NdikZAvgaCM9wghasF7fWexOwrA41QBNk9MhA3AWGb+1y6fPVkzbORYsvf9H/wDmwAsGJ
RB/1ubITWbJIqayPZoxrkQrILOjuqlMKuV+Q28eRpjOUZCeGpC/spchMH9ZNnNegShSzNsZhEfxO
2iMmjXxB6FnPZ0Lz86V4QsNQ05mQ1aRh6mBepkMHXJj2U9+Uoj3FWhXRfN30eh5GQVwNr96WzUIn
vPULQ8DTGCdMmEAeZ0FDXs/BSqgjbBe2d1GQqHZs5oxR/o0GMlddlTpyw8nNMDSh4W5bUyf3rgJG
gzlwPFhsvYMWZhTyFBTjN8DmKjiok83zaGQ0t1ZxZLj4KDcEuQuE6zO3+W4BaELGBTIZGO7/7W6L
9o+fL6ZHjd+qDafwIeyoJkTiJNV4bXySQWc67h4DsxIdXip0nZF4k69FjaywMOW+hwFICI7G4Ot3
eEoKNUbCWCgxbLL/OGvVmI5rrGvrr5zfwS4YfGJrjjRUTLgAsMHMU6id5elYaN6PRS1iq5D5eSOr
aht8fi1YImYEuvpfziJz8tomdMMJibty1RDIc7QFHPYXzQ24fi0QgcZA8fjPAMcb9E+tmVQ4GPDP
tQDq8NU/v0XrlbNijjvk+PgPkh5VS4SDGG/KgvS6zcy0wdrr6EfEKnHuwfCpWvqoUbwFOBbQaiLq
CvZjcRcbmPNZIcGpjk7PYuJcWaKIOh6rSWIsYUT1+egrssoaIRDlxoLFcir3Gm87BcbclJ0pPljY
UISt4WI9SFnKwFZjOi8SCelNm1Qv+3IZldgrCxRrwx/XpxR/8ItcH7/xQH2zf1aPNNvEjIK0M+sg
MhHqLaccNi6SsL+OHadikxapZySKWnh3coHVMoVyAeQ33NVbMBXT/fXD5nZec8TZ+PNOizx7U1W1
yDSeZjm4UYOkX7NUccCjbE7kx7pCezXLCgSYLYyiS4AZSKv5s7BDgcawToRCPZf6lAKQfyD4Oni7
qJq6IPP/D3fwOdoExi/yGwv5sNvZmoFqsLuWifcMH5PqGMpOjM7lFON/vqyUqLbxWDfU+2NTbwaf
QWwu6iNcm5+OvFjaat1PG16Nbjfk2f+jCzsg6sJ7Hj1BwlFytYOcSu0CDQQfY2T2s5vwascoAhve
9NYvVrTlW2Fwvh5jyYDi/90HzXoDVz0jFBpwc59pQOvDoYBvNoh7zUegrT8a11msYnL3wrjyHsTT
gIwKa8T8AwP2EtGhLEcJKQoOJW/WVO6+xXMrMiOfTLp1wTyRVRsPbQ8fvOFkrsPHCAXPj08j3YjR
lgZCnZzkp6gtWfodgBvTRXUQrW2MZfMCqq5mNMbYFzyyA1yKmykMOp/ek9AS5sCe3BvsMvGUzHut
Gyd28rwfd4+9lAFwCxRLCtPUqUw6SMCvva0D1BXSh3Mmm12oSNwtXjCsltY7wLWI8+TYXRad0P8k
PuK3u2nnDHedJ9E46V91Fx+iKRVBUBdIi+OebMHd5S7BR/txrn2YuaAEdu9oQHHNAnp/43SR5vaU
NgKB33WV4ePt91esFtYK2c9/79V/n8Afh2HIrTL0OmtA52F+ujWBqM7Hb0M001hZMjoQ0HH843Ts
q9z4lgIKUrcDp0qlWpJsmJw64gj7h8rDcYV/VWZXV7LE7Omag0XlxH8p6/qSeIYSIGwaB5E0/uFY
mwU0lZCatlx8jMtLxmaR37AzXqiU+CYcHADbyFI5d1Q59NzKPVXnFzhuI77tb8MgiIASfGkox512
Z75gKUcOm7RKnl9Z7viby6Zv5kfKSfbwXhL2/8j4RySTykFUBWok392YXm/hEPADV4psunOwFKcy
FGz9yhbOjTL0sd0iB/Yv9z7FlcVAtKaVpOtFm/F3Vo9FhnmwvbzewxGUKAGGpk8bGUSJoCtHUtCN
sUut7ZhThpUQarJsOicAbZfwW28W+7pcKW2O0ZNtWa3yFLzq5QhWu/qheAAUxRf734Lxj4WxjnCN
UwuJSe90dcq7TyR2vYLVjTVQ4S//iTW0JCb7y7AwdwkrH8LeVe40xlvQ4cs6j8AkoU3uxTtsHa88
xeOyRrtX77vylTpQHtzpvK5aX41ZRHCUnOHmy7AowHiREEIMP82MdZCmSnyUa4Omk8jST9IOFPA2
WrEgOjTSaPo7EGXCHnY4GtrP+8yq/+kDWFsjyPbu8ZtNCiZ19+UF3DhcRB8tpMzOov3UCbt57FcB
uN3Yu9RVc9ArmZeAgl41pQeF7Wb06YU2Rb0qhqPmHpyAUXRxXvi3G3IQkFvSadJsEaixR/9CqR1z
Fjft8HSxqzJZbjae0t/3UguZ1Qubr3uOYvGaLG9389AECK4uF4gomfOaJXpUKtJ71YAYG7c/m+99
eaLnmyBiNN8/OCrG2270yPqmx1a8yuxcWmHMfzzeCBIOkFloS71V2F4Wk6Vaf35smk6hzWXc6Py5
Jw5KZ+jd3bHzKSV00n56vDzArGuMZOkPdlEwOqTAfZsLV3pa7Ekztz6koaUjSpMECrmZ0gQWGJ7j
qn52cSKNWgVPLshRTXfja/FbLu/vL3qc8TshKjEHsnrlaHEutPvSulla/ow6Y0V/oECT+fc2wJhq
iMoSpS5VG8unc/Zm0erY37teC+NImbzUx2DxV2+Ud4VOkONaaGY25puAlc5TIrJ5D+0gUDXXvAJz
TFEE+Xy1cNythxWEZpkwpF39yJKloQB/bp7poZkmCB+C2OfVrCgGlLaL5JD4qW6W4KofBWYvkrdk
r/nYvxToWM1ac6aUTAqlcqqUJyV1mVTYMaprrTZ9ffLHNBk7rwa9rsL3vLnQlvOzlRRL8E88TxRL
aRSOdFtPYv2+opmGGQ4KONDTPl/TEeyIzyYPIAHjmVe3B+pSizRHJRTD9F+stjqfSyIs+amDaFrx
BL4ojfQD8sSCeahkmLgyL9xsAanvhYP/XbRAkBe1+yeUf9JPazXhAFW5dUM0QF10iKs4HeIXVki5
+Gsts4HhmJDiP7yEpUzu39BqIq9IG/bEKQpScIYGp1oOXAHK6u/k10FIOKYbWz/SnLxybHbdnxlu
GaCex0yUViYlkgUnrHmkFIHh4KAaoDExHWdeCXFUOUAqz5bBRbEsmRSPBFN12r7QfikDLv0aG1NW
yseQOF8u6g7mMFty//2x1eBqwfuHKNgnpSfOEzpOIL3GFAaOjIT2Z8lFp5byJ9mDGXaHD02TWe2Z
wa0GesBVPtrUx1rNoR1/VTAWnAxR23sIw4eu4xCX6k3gKMZ4Mk//Bq2K910oRPFj62M7bB7gq6KS
Ka1U+Xead7ed1wnqkwUPDD1uv0QdkEDwv7vwb+v5aXqDGF9iZUNK9K8JgugHl6FiIw/JeHy98To/
ZP6Xbmi5fdExgDXFhUKsbga/0g7cRGKN9/APuou7AUQ3C8Y/DGou+3i5lIktwfaneJQz6Dicuf4f
Lxzaw6REy2CYO5ru8s3LM+Z74170+9ZsR7ZAsUqWFCm+ws8WItaLUOw8jFgg+O399nirRJdR197e
k7XEpR4NbedZqYMrIjOVskd/aZ1h80bTgrWqbXWWzAQcONBin7noEIGaxhAW+DdLygzjNZHMx9ry
+nj9lF/oXu0vsrfP6tPeTq6ooc83wEqVeH8y+QwkAojsLPh4x//hiupO3zUrbnzOhQNyXrSjDI44
XWp81/iUx7mdTKNwm33bat92rsV/iRBPfNIw3RwT7tdwsq4GIIKuf6RUY/8Rvyb7COr6AdFOi4pS
zzYTvCbbss7Bg9C9DWxoPNfIe9K2fAyeLZPnPK+csh+jM99HbTvj9CiYIpL3CecwnPAKoHXlYUo5
fUFACVBrDY8PBpLhcZcUDLqGPq6E8zK6J+yqTsngs/rRX8tAAi0q9lj7nztE8I5XRmk6wbXXz5N3
M3amwBEW9n1u4sbkM0ByF4q/rJT4CqCR8N+a3GYej1o9GBZFxpvOH+vcQ8mlIyhlMB+Gc8Kup+0a
M2Y01P2YDJ6pSjKTwY3vlKVryU8cENZrGUFZ+VlEU6sfhMyK3CbsjlqtD/64eFAoy0qDnBDVbGe6
t5/0nthV21w9DRvCpdo00WLZ9+hrjc3TmdNioyLtUwRiOdDald8lXdQhANRK+rNU8Ug1xM3YDZY5
dIJIL17esVVDvtiEWm7o+nqh5Sl7FV0zFyOKaOP5tz9gtrEzID/1vuyaBiRI2pq280+UjQVA8kaB
jD9YnbEmkVGmlQBfAKHV+pAXgJLqgUFbjBCR9PHUPUsqiwqUVGGLR1oAj45LiZOl0vqMzIRLSJLK
aoUZvAT+uAXR7AKGOSWdv99/Rdq4Mq5+nL90Z8sFwnl+YNCKuuvTAualv/l/D8SvT/qZ14Ir/tAC
9IQlV6cev+nnSmnc/nHq99jXhpExsEovhtJLqOsnrIex7oIZP4faGIMiBhefklLWX4WnqkNMSurt
SdY2poyidj5AimQLtYoMI/B3cD7MME8laN2rxmGd/EvWZZ/VXntWfYkUzbapgONitE4N5dnUr+2E
S+CjBWbBJy8w9XuYuy26Rl4z6Db1sdV/qF++jcy2xmH3MqBYw3/UUiJWaWND2aXK1vJIkZ4w2rXP
OjlKoNfEmV4iT4eQlhZtxrYhOYht5YtDSA8lKR1RjYysvLHQknNLfOJrox+TuqiZzCQxUKIiNAOR
yWz1fcCDSyhHG8b92jIJdqCgq7rZB5yba5Mp9XODtCeDK1l6S1WbEsS4d4OJucbAs68DAFuDhaix
n2HosTWeLS9tMsAmZVoLmnv4x+o3POYF0agbUBYBOFIJW2tv7BDioH1p+TmPkphBzy8v0mPXtEzF
ydcDV/qhB0Q555XqkJPWfvnctU+sI5Itqw5bPoKHAibak6zIO5bDJ3whwcO2vpq4t+SHE/MHjcMV
mDKMM/w0L+dMOKdKuDiPlf6pis8F8CZERo+i9DuxvBjZg35mhZCJkgGd2Aku2CXU9yI6mmyzogj6
mVaV4eG3f1Ie4ZsjQ5yxLeOjowhoVx+P4NW0jHgyuWDmjzrH3B4Eg9Bd5ivNbfOFFFdu/CploVOx
RazgoVPDF7g0bhHaWyOSZ/b8n935bfmfCN13EndCgJyz4fl2yW9hDYdbx+QyG/Wm4ycR5QUPB4YJ
JU09bm+45yzdfUATIprcJMCxnujfGh5s3j2IxDwXL3YUny9FyHvITib7gpXG/Xqqm1vRet2NbR+p
DRnssncQ4Az8XPDYU0ktkgXM1CoBhMdtoeIFbj1aFCsXE97gS52ArW3/YR/wZ0sBwhpTKiTbFOyM
TgOwqHmDsgTsEZhmRNWEV4lzFjHMS88BMK+hzehX+VFMRTpSwQwzH8vhFy2REFaPT5gpukibQp6N
z8kl3h4p20/thZGMRzsJjKFg5TL//05du1DdpH7rJojq5oEjjDC4yq1x+zZWgOqhTz8ZloVA/V2l
1HU2jpiL47D/nBsYdvWwvPEwmociQPECXbrsknpjVtCboDqVnmG8Hp+W4nviLfxzXD3XU/bCj1vx
CUYOznSKo+UrE5GKeQOMh3LtCzGj2yTbOBid54ueJ+MuJNdJRZ7bBInRt9IB2uzjoLmuFGioCGBc
eN56Wpxw5xm7HZMpWFNOwIyTsvriChR3VKoJZBH5FjVeL/U0zTeIZsBkLSLXbIvVy/T2LUBB9G6v
H5S3HkzNBY0VdR8SQfD6wbYVUrGS3GZsnutJhJfCMip8hv0D3VaPTlgjwG4ujyBgXz6ca+7CKHo5
2Cx/sUYAAoFV/1I7rZcviuY8PiPdo01EdAOxJTvpsfr7SGT8VS1Rzr1sXtQ6jo4YVybYnyaX8x/i
84pnOv5kdQzxpH5TKFtSt2VkzbfH20N6KKSkOLekCvmwQUI/5bQyaL6ypD8qZdNmljrtZ0g0wer5
VtdxUARgnjbL00QEr983yymqWKHoQU0uDVn6ooNI61pQ+EHPGBxTr74d5Deg28pZVUUrfvuNSlDW
xpxC7gwIaFG9O4Mx676gp9WJiUKkWRChAPr2JdUmJxzgHdqIyjx9mCuDtk5Vvo0+nLH0cfWrTX/A
pdagCRoVMAKsy8VEC2DDiUoxujQSYD8vqMmrBurUofRR9A2wI/g1U/QsQP5qnWiqeRWx/e1S6zF0
T3xJ93dAWxQ1g/6JFBHmf/Aj2y5zxqe85IsAq2BPKIoQiTjGrV46CxM1QYTOUDAvZm0wiH08tGyA
BQ4Xr9Od8GX7I0EGA2dg/8GT2qmKld47jwGIj2GKbf+o4F/iaY/WWnP6YVavuLdvPG/oJ5xQAYFw
5gQXRCH6dkTEqUjToQW0VxZutffjLs8qsqq28Dg0N+sB1O0+pgS3VBHaw2uWIK0c2HcqNleL/aty
tozhRRxmRwAi04v2vUpw7UKIlV7G5UYJMq5MZ2Yvp5VW6Xo9Uyl4WdZCkcui3ya+g0ofBx36k9fS
TmTtFQghiPB+ExyObwsh255s/ml6TGkrAJz4jod2FfufiShSqrEbwA9fp6+g07ltpyjplA1Z9umT
ujsrG1rCk7QdqlDzcZL94bMtYeYzO+GHiX1VhVlvVwHorakuqnUfN4IA5SxaLD6Tu8UusXrkvNqj
qUlqjiD5GYRFCyP5HSBJy4QMHdJa7BtLRF4vaGfzOPhUHRsyp3ABcr+OOiwDNqgL9mY54chlc+lt
Zv7S/tx+scJB1ESi7zStHoPqarZjALJfhbNy6WF9zFNreIQ1HhyvvZDta669QgLNTLZ5U/cH2djq
nIMw/1BEbdW68KzhD3UcfTk1ldOZ8QU7Tt1p/0X6VSEWWzE0SCQiF6TNBj+VVMYOzTM5dVZZZWHN
SsAO96gHzTya8DBpg8whhHbp3QfCW8aTRU9qL65+SBF156GOj0uOnkZLJN0LHD1/s8J3Ofnh7jfa
fF/8pKglubyLrUbvTvi1vQxkziMXXU6xBC3TmLujKbwTte+IeDLdk13VVgI6P8fbYf1HBKk3lVAX
PVEJcq90VQTeEjxRNvdTFq70/dW3euODgYskmZZ/7xwJ5H7xG5e+E0YDabFu9S7VuUB/0X7Ucn6J
imcKvbsWFDth6rtFu9oZlulKXuUg49cAmWadpzYNaBKo0Nb38oISg8p5ZiWKQHTgPNONnAukWF8j
peylIiGTTdILsjYIA7mdi8fzMSBjhq73p/+xJOzXX7MBdMAKr3O8WKeG1LWc5EoEr6uhi+7leRsH
KH9+ksfAcoP4OiyW2SMQhWvr0D+UJiqfwzNzPQ8Ax0R9CqQeAJLC99t34yDAYBzXIR5cyeyMQViU
ya5M268MCaFHlIOuQJG6kLvnpOUaZrFrFAje5+zEa6UnFLGGSPYI1gs0IZKFZeqxgOSZtyIq/ywN
xJwQcSoKSI5DX+mQ7wpn0KkX+cJH501qn3+c0jmJWKgTFri+tsi2rO05/hF88epuWlHqONoP6WyJ
zDTkcwKHCSIYETjTyXI0NUU32Fc0XD9AC3o5cnkx8H6RTTNTW514zPBG7jId54HWdyP85KPdFsYK
7/jj3wZiZixSPxSAZN196kqfIF5MFoI7eOBvbJoJywZHTk9A2OZzCbuxUq7ARn8ijb0LW4wl0epV
empxeXwTWJo3cY0CcUp/wsjJWbmTr1H8zf6JOHyLCKrmD4Zlacfw32KcYlu/nH9Out9VNEDTlPMb
MIuKRuf6nnS9/q7MPf+hGMg7dSRVvZI6IvtqVNSX2lpDo1N5uCJlecKW2HEgHbswhQRL4+zwx1tE
hd4Xr6wWtIdep3E2D++cHLYE5BM9VF2Mkva7f33lNRWNQvF3G0May1nBXeqtePn7oHfYDPgeZLr/
QQsg1DvZtDYwum6Svd+yiOz7lm+cx3o6NX63w19XaCUjEzCgpl3fEjRhPctloVJowOVxLjKUnO+q
Akr3grvvwvhaPHjek8gvhgN9pLXn1BE2GvxWr002uogrDxo/HhPYuVe5e5QV1pVg5nUQYeFXyWwe
j47nb+gyzdGrN4NuB2LBQ8N0O4CAnokH42xpX2B146REk/bjUINdarI5wV8FEsnV49EehDZLzvw4
q3Pq+JIFSpFLePKp9SdcD2N3RNpNYJynVyL21Czt7YpwPgPa634U6YfErJ09UbxoMeC5QFNntVVa
v1XEyRWAxG5HVvQcGtN7TZQiHejpRMxiclEd8QcGZENueoVlSxbuh6CiuFTBpcwlVwIdjC9PF2iS
Zrm0vLWUP3dkUlBKDEE3Jd36WOIi+c7H3yEMSFjvI8YqO3HNeNZyFNqifO0Iv5XtQnCGOxxBFXuM
ZFpB7t+xJux/8e8i8g3mSO7m2wCp2xkG8/B8LRpmQnTOo50JeB00atdHw1fq5DDunGNykvTJBWg8
QdajmZk8VJvhhggw9cHkXezlQsmZJ9YsoVGjN1YX6+H60iURppMS2W1j/OY3XlSP6/7YuYRXwGbB
lKiAyLeunJF29Wk5+TbS2bDw0tP6AEa3y6LkzvO2NvaJYGBhfbNp0BztPp659zRS7KuDoiL3oUEZ
SUGjYvONSYmO6eJHAjcZb2mS+bW9+4cKAuNOE6o5zVIpCOSrH7xWFEcMj/ZPjB0fjmnAtxteOwYx
9pUQXINQtL3qwL7G/m3l7lDIEMQuijS7fWuEpwbhEbhIyzJ1gBij372RrY/YJ5rN/tdZCCvcV1OT
PZSmDX8rCXqZkuOXFejBnLRDq6I9fjLpl9SvIpfTs0O8ZfoyUoNOAybqn07KW+ZKfY/DqpVhgmcb
uhz4IAFDHbt/iA6FJom3WD07knf/0ezEtLSL4SSGLFhGSyHTkikpJ6ZfyxF08p+Og25JU6M4Vocu
q43VzxoHUSlrozTcwWcoq04fXsgiZ3HVw8FMTOmnYVy7C+h+SP4b2rUq+q4NE6m1UzKJcubj/q7o
z2v8yCAfA5XZtHDPu4dWD9k5qS+qyUA94OQBhPGvwULXtSzRr3yy8ZYVi/Kx9sAjuKdiik27Xf+7
3HOZh5YC0ypN2JosVHi/jSg+q3SnXsSZ8TCbsvI0VhCOaeG9/xh2ly8sKKpRNiMPq+TDidRHAgzf
y9F+d1pG6+UNcieSZMrkw13o8I56FhL65V68UmclRKiFwGLRfPkP4L2/oMn1tZ/3GxlHWg3Jnt8o
DIYRSMX7/+VcUShhHAs9JmCM4lI2Jjb8QSqYQ7ip3BFhAQWTRp6G1hFezEFpDvs0m2Em5EzqhOvt
DMp5n3UI8GGf2q85AhRLH11m/bZk3DPQ3BvVZjXpNdLLYwCUGzmctmUNeWydChNlBlvU8RZRiyM+
6EIBzB8JDR+qmKfRBhIZEDD6mgkhmPBXUeWLxDFd4JEc/Ljigyx+o4nhknPUg2nQr22v4UFtjeVF
3oCOi+h7NmywTwh7HEEMNqn6EatI8DbHvaosDknoFR9DSNB4MR4+bvH4nX50+S1LhcVQV4tE+2bZ
Zqjk30RvG4MSvomyCrCKErYvu689ZVjLlMDNctUoCfau9D/nSQ6QSwzOZW08uGpRx1KM+WeANvEV
Peq4CBJ6KQFc7QCfZddXVcAMaZ1GWpheeLQoSR9on38BhEF89kxMBHwJDJDlBJcZZChB6zt+bAt+
tkuPiw5t7NoTLi5sXUXl7Ln+yLJVHmgA1sDVwPMRu5tYN3vpLqkrYxuuuF2LLpc4YAYNn1IpPojG
7Fitx8a7NPeuCG4Bra33aEdZPB7APgJV0lLQTM48FvGD48umnGpZHFeXKZBAttKAi5x+J3v/qMO6
nE4QKerMLCNcSlWG4TZm0Jv7zsoAyDRd8KrKyCOQDfDzJsdItDbFg8Hxr2sXD9iORrb9LPKcqDjI
pIa+zKVpcQa+JkM0qoNosfu+c2rtPqZdVhkXYTC6CqgWqkh1wPlC/x4utCnw76gu94huS9WQnkYR
5neS1vDtxKOwFPvAx5s6eA2ql2QeoFsUpplUC9MWqLNzRr5ANMUO3jzA4xpf9Zmc8eEpssTNCgel
BQ4kmDwRFwLsFidylJLMYfWrySpxwKfR8QytRDAgjDxK7T41G6R68tyP4/JP7z6Z5LN4sCHa+99H
xgGBjA2XtlJR26uUav3hfUFYU7FHtIjpr/7fN8pA6b4HcB/hYjMUzpiIy/gQLBvcvH0ZU5/sSTK8
RTawmU6duaEISgLJz8IFOoJoW+C735UQxKOFYKilhglunKLJpqTm9BLbXVCX46eXSKyYE+z3pgfH
gIWH1yR4hSLIs/svFy66hgmAJk7V+Bq5HbchGUQ2tFH2woSI/zfLS+wgwUJzVtxp98cTOGZ09oQr
R6M/Y/gakfXUCQQ31hWTsU7+Gba6R1Bk4wHLuBYd+cg9UMuyiBrMQs/g4sEFNbxburJGWorjmorc
P29+5kTiLUScMnesBMCw6lh9+m74BEsgGa06VUhNOXfRTcHsdzPn2zJsi+fYfaMdh8rYSVpk4yin
eId1mWZ6fgKVFAJIMm3hxUCcUmCjP1So/LGS1lvKHc5pc6g93ifJ9znjvS+0DbDzF2XH/ySrUkbO
avAoCv+F3HcNUEFjEhVDHPEpKESRK75bxaRMtYmPYnaiyhPn4cO5cwB5+bLx0CwwPvEXjgyp1sO2
TNw9ptpqfYLETU1lsypH0FQ2Z3ixvRQO0yAKZyb/YhO6097BL+7xukha+8uhjHZwB9vCUyAz0m/E
0sL9bm0Fla5PNdH2NLn9ErqozaurdpRmef0rFI3168tK9tcNi3FronfMs76FOlFuRzIJMhevtGZJ
1uY2/c3tCYBuXYEiHbBGp1mk1T6/C2lS8XDnInsbxF9d+eOoyXeZhHEsVDtj2Tcba2aWeDp81nTg
lyVqFf7Jw6KwhMq7HNB3Kfn4vvljHCZLZk3HZT3Pg0rYfBvWzuSmKyoYc1ujLJ8AfRMAdtnhUfa5
zgi1pSaY2f4k8JFlkep1RncCmqxT7KYbfUYJrZe9XDWFuKUOkZ0+CP4vC5UpWSZRsEKrHvSPXfui
T0aEBN+5bGvWYlpF4kkgwVTsNUTGLI32iuzTmz/wdU4vrPB0gVCthEFboxIuaA3SriVbxobBmnOv
2XSpHG5sIfQkVPi2Tt+UhN5ePDUSQLvYK74An7E5Z8oGm1cyo7+tb4X3LmZILvPlG1nmFU7bVrEC
xzoL6UgGW2kSRVspXyjNib/hqF20KZMVSUZYbD5QYsU/ZFRN0evNKnBZuo5HgTPYbsklerUNL/CE
n9+Dc8RhgDAPBgxSw5R//9UjGAYddVrpHaMYENKhWNcZYbCu2SuslT4cl8Sbl5XRxNd+hATcpeFj
IZkBrQX3RzVHDIvfKTuYblq2Fiy3i/0UQx/OUGhvX+LOL0Y8Ay8AjucCYlUG6hQ+wKfXw8ckYDFS
uWJzx0a6cYnfxS+Hgs/y+34Lx6eQ14BYkbVgjH44eN/qBlsotqwkjfdBpPV0bMJFQbqupCaXbepE
mAWnnGBm9qeUGJcf4J0ztpXz3caagIHZGuhYDpR+LKgcTOfRRAop3Sh42Dddi1/7fiv/UGTgtM1q
ZAcFgXJUBXyStW9OkxRwfW0H0LbnmgArB0FKLVfSMrJnlpU/EE5+SLeK3iL8pBiCvYhyeMjImymm
dSJpf+l9cjjmNCaX4/ZdR6wFijHBJioRLBg4KMNmhg3+4ssv9d7nf1J92x52L+slycPW0CWO5/C6
axGxWlw2LPkAP5B+AR4e4WqkVtkKu6jey/t4IBPndMpRhw/wQZnsKETSvOqajlQlk3GkTix85Tby
SqFXeyDphAEbx6i6xXZFp3WyoOTgIWJo89OX7DVkJnEHzVITIlL2NEqwPoWYPP/3roxzn7BwqcgB
febuJEcUdcEBx2u1DzHTK4CFi6qAi45/FEhBVP/ox+5jtNYm6SIqZJJrjkkBbJ9+ccnhsCOJ/cng
cGxnFYiYAE4Ab7JjiSm98DlL/5XpCSqsKCXYoPiYryreA+01aK67uotmIOU/reaZwp1u6wIPWVHj
R0E7FVyTvMg1MaxM0xA8Lf7cM4Q2u99QwPEhvGcf2nX5VceUNuqCEG5q91SCLoP/oKHkiA1POMCh
tlIRT/IxfDG8UUw8I95apL5fkiVQbkshlii8bMrqpnSPefJzxcQW0/l9MivpcUKvTGfk+ozTgl5L
BJDBYDOnywUG/BOScdipdexWEivAf8YC/BngCkpYjApJ2jujyXp0tJ7RZ9X9GO8PXv/zVvMLUdX8
neD+U2F+2yMXgeaok9wD5aijEgrbmdWEOh2rFptZajJPBI8fMM4SrWF8r3ST7nvO1/yWxZfYyhyC
mN8ZGx9IL6913iIIbs3C22PWW02VTPXWfoOixr40R+71k6UdD9N2TlLCpxe18uJ9EtH78hF+W1iw
6FA7plIYn3XnbRjOGfzxWKlnR4Ws/MeTTAapLJD4qZ/pyHY/OOmDPU3to8He2Y+UAdlb89FR9GJL
wiQ+wASi6ccaUl20GJJl7FliWmmR2HDa6hlLq2C8iPl2Qp9DFO44WN7npVSxU2F6jKoAofdiV6S+
rgLTUOyFxrwPepDgRxS0XrsYKchmxKPBfgqqNYsnRnk0s/HTO/2YVvmj0oPPKKZ/bguOebZeQRfG
Df+2CZ2roIlJw6vbd0rABtJVYJetOgg7QiMkJBK2dWqA1TCtSPuk6/Gv1KtJ3sI3gLmfBbuYtl8w
5F+eFmKrgxBRJfYBm0U2VM+d4np2S8qwpmefvsYt4Ww48xfYBE/AfZvIfkz8iyVTdMDlSwhIuQx1
nhvpRrty9YaaHttMEWj7ULHZpjkDE2u82+UHgLBy99l/NJTSAaiirBStkwQ+d4hVXZhw3COVps8S
i3DI0yKgHfUXUMXPvHrUXgnmA5j1qWYMJlisWJy1J7EitaN4lWCGaUFD6L2OokDU11gNKwk3nSgJ
k8DF0C3wNiNedgz2Hp8d8AbGZx/d5rDCSJV1UMPoFkCqdEw4WEv7FjWDxQ60Ox9qtngULhTyXaIB
Pqh0pC0+qmkJfNEs42i0Sdmrp5ZekBQbXbvzWvf7lJ505RpMsoLeAO3Nfv0qilEkMoepHPUfAB0C
QfjXdw2cL1MnfLPESRFVgfL91rIMg8Ad5Nhoe94XFIC3Qz2Z28qvp0iooMxQ0ozKsJMbYRIPKrF6
CFRwep/X++zhmcWzZBeCz+QD+zQxeKwTyfmJPh/SypuojDVNIlcBE3SHn0A6/lB5e7vp5UKz1cWj
lLQol5HbNnjdNULTJZS8UT9U30/erxVNo+j2h7XlH9Ie9Nv4As5NcjBs0EP1LjpN7+M4/UAjrtLr
aNwen8aDYmIl4qJvk9xSoZGdWtLWKsOWxi4D/0tWZdHVgSv6VS81DacLyNXOTGouaM64MDCBMwKF
+v+2OqmBiLk0RV3bsbssXGVG/nNkBa421jj6EW1GwbxHsOIslVenRNNiDKRIGafUIxLcsOSg5c+A
rZEKfCMdq1BE82XrxnXl1SodPzpiuF0c7P1Hx5z9L4nQ8Akt3OLz3xuzCpx50Cboie5d1a3Lugis
x2jQbLnvmNYM8nnf7nZzvXhyAZFAc7t6T4KKRoL2RY9chqnEC2SMiqDCedD57n4s2yQvYjyeQVtS
AfWNAfZC1O2Ah4vOq0T5TDKCHIkUY+0Zg2qQzM7mt0GGauu0FKk8nMjCcFn1MmAXQehmKzhiDJTU
rdUDH6HXxbtDxDc6FI3lSqzftfiOn1TuKLaEvKGyyLGirXJzW4HWMRfD3MeDcNVLlffvtPZD+/ur
BLtgPBoz0pLONgcsswZwwB2klQQDt29rvrJIs6OWgcM5U7Mnpn/AtVIE5WwQ6JKxfUzeMpWMgEJI
k+QvpgEvpkmlSHgAUM1fc55s5jO5743vCvyWlPFfhuiYfPB6P011ZhxgryA64zTMPf/a1IgFKnkI
BvGZdZ1GeaucUYBYe54YERDZhwpF8gQTuFyFtCQUqzZSNZK4E32K/k6oQInkTeHRBu8/UoLUiM0W
YZRxMonjbOfjq+zFAPDpGOu+UrkQe9pMp1aYFrIOtIiX3Wycq5zw6R8a6zoy9cR8BkN5HTIm7390
8ImFT3JR++yokjf22X9kf5bCy3JVGi37NBp5cj4if+v5/EbK1mA97wyRyFJYIE7nzO9Zr4bjFg9Y
GLQrTqHQS5mrfMtTX7hHgs6sG4/PR22aVjkYLXIzb9iDnaRzq1S5msoDiB+njdnRRrWmZQCK29As
3UzB8fdbrZx9y77EiVMP6NP7mTe4ArSzh4C31Qnu8klhGmBEn78tKvpHruZDM1TvDMwIa2E554rh
s0UIS6yVAk1w8TOcFz4AiKnVqx+fPIOUaeDWbmMC4SuupFIcU8zqwB//4PGGYNu9JzmyCzzA2aw1
8SGWVVFPmCqLmCH49Hc6zuMaIaUR8HoyJa6WgrIpOQJpODeOqNC6ALwaS1gYDmGq4Hf9NR1EX5AP
lisrO163lbeHnNO21ts+WNTr9Flv7ogCxdLWJt0NZQ/Rhih2XfQqAeykZnNwP7CoarOUBpembJMh
kwqsfh6LxSSjafGCiJGRL1DIIlHw7tzIN9MIxVjF1R85RI0kEbqtm101Vz+mzpMt2xrpPuwdrdtH
0B3RR7nW5VFG6xVFmvw1I6fauF1XZNTjBJES5FdXYJmudomIyRCIhGLsH5o2nfNYOFlS8XItd0mt
b50A3wIb4OgpIsGaOG6xV1QOGsHE3qANyk9kIztnsuCbCePLp/0P/9g1/qN0/uAOKNdj8P4OGuQz
P7R6QOqllOWsV7m8JGD9EhAqmoivRZPumKFF0YalVLS4kVuhDNIBtTIM4eGTUcx5h28hxmDOE3Q1
oFsGhzyngypHLJzH1z2NH0NRd4uU5fIZHNpL4uH+mDo1kHAyuQmPa3xbpc8z/gKtnvGhzDjpkn3A
BgHXxYA2KEEY5FvEkl+dmxKd43zEWi8f2Mngi6g6eyuapkJXCaddVbZuJiSz6GcR2NqoE0+qaR3/
FM8wZAMXSaQCieQxPY9GfocV/laVojSw5l/MJaQaYT3VLqY+EXN27KYKSWVZbuMWJ1uPjPZiOPnm
HX4Gw3P48q/s5wsKCIXOYZRd3I4M2fci106tRaAt55Uh6LIZopz+jP1kJHfkV+870/LQvAZFA6jw
lDEeIYMugvrlj3pASs+Nb3L+PytE0fwwze5N9fkVyKJ/WhsoYW7agEW1MMxE5JUAic2P1lEFRpis
FIEEXQUUtA6sZ7kwjj5y84uGKIkj8EXLGtUiuOMtsDLs+vPvZaHMeEP6Rprser8j11qdqgTQ06p0
MzMwj4s66wkhQfjP6xM6NUMSlZGwdP0JzSjknH3kPZRTu46v3GQFervrMX7QW+HCyM7B9D3aym3X
tGdkpps+Tr5+Ahl2lkwokYhsqZT2xIIP6CAkHk+PCSohhKh1sziy3FfbUQibRUJgTLWsMUnCO6f+
Gdzg5IDg2i7R2F5jl6CX+PS8bdTpdX5Xwb79DTw3TBDx18SQ3V9vOAff75x+V9I4OTLtl+xp6uoa
VueMELSn66JWNoHYIasXJvFszMqibkafNiAnafyKfhtnd2R91hVRS9jsodTJwwQZ5nyFdp1NhMcU
chlvz2gpicWbScvhEh9HU6gtcYs8LYozCA5GzUZdKJWWEc9lnMoNBAp4B3b0gmnJ77A2O+KFrZEn
2BOeAfiUEEVZutd+FQLYNzrswmZdek0U46DxwVM2slgVn5s6DVdW4TdxZweM4YBeI/rgJsvxxcl9
MvK1AttlPGrH2TDpK/ocL+jjlDenv7XFwaFLtFl14AiFbrkHb/qF42IMyxL5uhRgn3/u75YFqfDX
4Mt1EU60gPKDrAf+2Zpv/NwiG2NwMpQWwUPyAA2z8vjs/WLUWHviDDQV/YLAMjvMhWJnsoGpcWvN
vSktrRuzHNYonwwBA2OrU/MeZ2TEquBL5LdJUK+DwEghwLeXiwzRCFD9THI1Pv9tjgDFjCUqAVsH
/bywUfZOyHHVCpDAcxvyANKFYYjM5IIXmLkliuxpn79SkciOz8yFIN0gnuseKeSRuVnH015BA78Q
VYBWvkQHPV5m1gQXRr/c3QPPGvSeMxSu2tmgeND5dpvZBXuGhHODfj7Au82hwRdl4/z4zuS5Eulk
yhl5dnRz53e4iEyGvFVKTP4GMWOfPexiV6u7130r5kLD9WazFVrzuNd2bVvs97YcbmyjGUy2qfSB
UVaO8Iq0Ven7+c+BRJkSprtuVfqCu8GoYAwJvwKjUe3yZ7U3OFu0lYEpO3lqlQxq7w9RNvyeqZKa
N/am8Ovt2E9jnCY22M19Y3LURNsjyaxi4EDbpqRVTaVTgkqQtWQM/mrv8ZER8QqWpxFuOXjEkxzV
3EHLCFyZRQEcPIQQsuK93iRgTwefnb/v0TC6/poT5ggo8tPnteRjaFXDD5MvKKhGHEhKMehsrJne
Wkn2RBqF0iqtrtfwEx19p1dtKcsc4HY6LF+QX6U7gf/0wSWftNm5U9kuNDjc2wnenwiKetRdSi+1
LvD2bLaATIPCzjian/x2YowY7reYbNMOWkb+qm7F+hFW45Kw/W9QppfFTYn+Pc+IZBvMwzpI+dR8
oLdRlqwY5WI6+91ZVAzQ+hCFHi3s+4R76cGzbsvW4NQQAqaufr+0stS2Q1ayEeVbB0urjfcg+WWt
vRaW4O1Pd9OplyHR+tCfmzD5P850kA93YJKvG76PFPzgNH0OciUFkCUL9kVOLc9XIv0UmQH2nHxl
bUXrMgueRxVZPvwjeCsJE0ZqR3xP3ljWxhH3jWaanzT99vWymI/XD+wIxyDUKNs/h+KGSpN0Fm7D
qyn2c6NWnMAZxLmVIDCfWgPMjWBNF3r/Wvh/Tq8rsOvj6EPgVDh/fR+pI6/C5Rj15gGTX6FydbQA
b6VyZ2qesYEXzO5/DSzwIdor8Rvxt9/RiNuZOwAvc9TfVzAwo271li7brVgW5qdMZejIvUOW859p
0RTaiajVkFfmjMTlqdi+yYTheeycp4js+Psri07+y4PntlaUfx2rq/+eBrpATHA1DgdvC/n97G3c
rVRxByLi4bt00i7H4r1THLJbMx8NIt0NPd3CifOr19WL8eXD+C5BtDkGQKfzlFkAS+T/O+wKAL/c
0CUE91OuBYLFHv+TMJZPJUCU8YYPyItdr9vYfZ46KE6HlORTfrn7+3VwflN4LlAueb0mb3YvGV8S
DGaIeIF6spMBXKQ/1VZrPf+BVR3hC9zmahVWfYpDRptNpviugx/paoORWww1lD43eVHonmarGwa8
lb4+MJTZW05Vi48JkYJm91sG8V1+fwyr1fLitza75vo1WOGFJborCWSe09ow7adzfM93txoPR2AW
vNfAB/2FO3KshfGB8JRHvnkkw2O5JSU0ffQw/BoNjExOWsLCnfOw/2qABxjnSiyfaba5aCZ7LXi3
n4Pg5kTbqjdCNc7U9w+/6a4sCzYUgnxxOcmJvmppn48ax4cIyZqhM/f3AhioRo+kRJWSyisHwtBd
xliD4pwq+7eADebL3qvplNotZHdJXxDAMLkYadlsjrNgJi0qhFLELmThxS04T52GFbZ84eDMDR9b
7ovzYsZ+8c61CfJOyCxO0eHfASAe9IHY35U+LaS/QOpvxtFeb0tcTxj+tN4zuHXvJi5WkNPMtHac
l1crrgDmCK3+t7W3l+/RY4y+nI/kuoNqFQUmdA7qL9L9nPll1qYxVFlODnnuRYPvId3vs55JvtS/
tDY2csWm6J6S/73crI8FTP6cXneZt2RZkvMmhEWnr4FsVQw4mhdx/5xMK0yo1w8DqqdXAOEL6sUQ
4+oZz+rdg8PfZpv0VEGMhnFCZbl4T8arb4s86CDBhoy2FcsDRBK95Owo/JqfTJ7cuIFK2Qcb0XCf
KZh2zTQkq1pDxOWVmZYUu57/0EipDO5roKexCInLUwdcQxgb6+AFcDaethTIRpSxQZkmRCNMsD4Y
MWROMWUOFbcp7AFAn4cE4iGQgVyEEKZPgFfdeCgaPHvXtkzYEYlnt8V02qo5bUMxSFZIzaDAWwe9
ZBN8lexLJMIWmYzwe9/k60/9uu7B0S8rJrZjo4CO4fdUD93gNxT10Gvizq0NFOYDaX99amS3ZlB+
Vv/Cv4SJ29ngWuJUjb980HbOA5/HWOjQW0nfAiGso8/Ix5/Rxvto6bA3bMow/ru8uH+UmU0i2vjB
dThMOj0dz+BatoC84ZwI4X0weiaaHadPRAXQ8VSlS1kj5risDviYIGIl5cfyg0TJ/XkfF9zf8pdq
bNy7mN1QkSLcbBOnpJMpx+2+dBtWFVxvdrIcephQyWJ34IMIVCgXpXP+z9ePaGiZi0Na7xaZ9lxM
zCw0Vc1j/hoRmdiynYnvXmTZN94WnU/Sy1a4JXZcASo54sxem0xp2fhQezUJmgGLKiEEoTstMTp4
uh93/h3rl63p+udHb6if5NfFCEICVjRMrdJQ9K6nhrWFZEXA8AASXaStP3mP+vEBRl9V+bEyt9Vr
Z/PSswENOsarXiMOM8R0braVEpOgHWV3t1skoBrFPBxuKCZt4xvEJp7ssXkNyo7shyjGsG6D0UcL
dd1ottrLSuMEbI8T6Tc4sJuwN+cPMTp9J1YMkjaa/Nrb2b+mYfLM2ztbKVgKl/SHYMswP/9G01RF
5zfOqO6BqdrDbVsJ4Md+2+C4RQ67w4k4L2NfLULA/KUIuU3G3wPvpIqs6nqtSMNOiLVyaVB5jy0h
FGujZvgnLJ53ibUX3m/jjHGKeAEGYdAKMjO1K5hztzOjiDPJlUa8jCiZs+5M2PnQwCBZO+s0dvFB
RbqdcYG8D8YJ9+Qd8G7RPKmmESBbM6jFcfj2btnaXVhX0xUOzokFMeRWvlcKR4qsI64UdNodnNKF
MNYc6t/chuLx1pAN1Zk/8KR5NOePq0ufW8zMAvJp74JEAtCbW6wDZ8p8VMOPkQ81ERLoYLqGhQIG
HORJz5A3Oqx+uJbqQRo/nYOep4pahVMLm1RrLRCi3Wt2B2kbdv0wZUJBqy4cnjKEXyWYoZourv+g
BtRT1TvXgcKC/7HlxTRJSo9xp2f/hE7sQvcpzwww1MUruOFwLDsmOzLmnn1WXJ/8Dozg34LIvDrM
Mj8xT+Teim1Sz0NBE5/CYgBJ5kkVUMOZ4xguGxFtL4rwwfeE3JkwyP2YliRdtO3TK/SNLfsC1liD
HE6zmycQgFDoVcKR+GVNRV3W/RZSojRZbLNFN9P4REZklE/kbQUaI4gcMxsiaD/x2l3MK1GcKEz3
HKdZb+abCGhL96pT362etGqlCpjBiU5P92vtkPjbUJOFpihw3mKlNiKhUpQu8enNVjHbMvJy2VPh
fvCswMx+ADah3yRGzLZf+h+zZerrVm9rMJ0Mw1I/RJoh3+4C5FN2SIfNL7hyf/SlLHcJIK2JrcG7
/7GOOMFqLwErE13Mn/VOuueE+6i3nIsfqq25+hv846bqzI6rsXKVfSRzLnA8utgzGZv1P5yxWTEX
dOh/Q2rlS/eBEXJygcwwHBoA2jqXRhGKASNulvX0bTIj47zvJsAkM98k3cmNxcia+9u5NGhlfvbU
0bVPkSsaRY161XZNHRLOws26h30YvMyzsMAkJB1bRl3jhGtFBEFT1oCeESAS5wD7qeUS/3Px/9r+
zlU9a+ZjjeYcwXc0K+/G9WORucvxQjai5mKriR9mArlrVXJVU32S5XgNisFufgUkybcWGMIz7Y5J
NX6lpGheB13vwYwmYwLG9Ar2fXKJ1kHtks7A3qgMZKU7MEjK8SRURtJ0Moqp+AT4y+QvBlEt2Tn7
gViHBIgW0B6i2Ju9M1GzLZnBqYN5ONX/ty3zZC5Pw4pdEj+G8kYPYTudWaGGfg/DFP8M00Ob4ziy
qx+y/mfPabZhx3Kl6zkzWYHgggK/eJp4FKIlci9CPC2Sgtw+8FfFNsmb1090V3U8MtSYaDh2FYgI
IPszgBEDRMPr5kcNeL8nGeFqtwqmEWOJdMxZZ3d1uOAXcnwGImA+rWyWj3NFDH7IUbk99TTMhnTo
aEeZpUdTFgYILU4pcMvLoYTIHFvyLSSx0pNfOs/k3S49LVZ9sIrRZ1LHLK3pr/RIZ66X/1ZHBfvf
Hwqkg8yj6QpGpu5V8ncFop+QJHOvpKUniEX5Y5jWMGZ+SZq2cq5VclpmY0UbVS7M5SRiLoNd5MGc
Uiqy3+bLok1jgwLf97X/y9+mu9VVjxmqIXv5XdzX7622AcFYFzId6rb1+cRQuK9EB9QHd0SPSD9h
mCwXuzj60w3h6wbGea0MYbVC3VOR9rDw9cdSMQeiy1CunNdasihMZCpAGfKKyJ2LOggEQQaZnXlA
psyXAV77STNFPxKF2JuJ38bTu9OJgCtD8vHoFE5kpbHNc0sXMaPv7juHU+26Idyma3LJKWZyUj4G
8pC1l3kEqAI7IZz1LtdCEsN/t3BYkErPp7zzFC+UrpbV5OWOZpB8GRIM2KxHxS2bq+Gm1+CrzW5t
9AJuzE5uZ3viux1O11JZaVjHceFFeJ4DujQA+Gz4y/x7q2QHDEqHRNiZrWddFTmM3YgNi9O2E5Nc
ETVqdTMHgT1V1uOwoboeIdIGS4In5Q5Zg9YqVinhfWm4dE3vAH5lhf8bB4rEp8LyGgdzBGVxhlIH
Yt+cM9pazRc7qyOM+kJwh4IfAoG/7NeyjGGWB1jDh5zZi03wR33ncgjCyDY0/W7pSsyqnh8cOQd0
+0qBH/8/dB1wMOozQOVgMB6nGrWl6YhQP4K6yk96oQPjJ9/Gg5knKTRN6ZYV7KY220OouGd+OQyB
arzflvQNICRlOvPkcOmYKdTC7iliptskB9ORKW/vDKiF1tdZL89f6ebth01Ew4N7iKxk69SaqRUO
krTfq/szUBGwiSw0BeacRoTAhISP8ytoMu57W5lXKWZNrmkkQy7M0Iprwy3xQT/qnDAgpF/BF2uz
4AR1btr1MUak3AIdAc5nDOlqUJCiuR70fTDCADVZAf8Q50pUCrPMV/kCdTjYNmoQBEWzvuVM5h2K
z+mHGBgHMJmXvNmN/dbyHE3a0PkZnhVszK/cR12plLKOuwifuU8IzMGwUV/G0Zdg4Q5Ssg+azxt8
q9xi7gQmPAEUoBjV9cmkfsmNKTWM88O1RbIPE8UYAyGLROC4ZKTStr+0HXRPcnuZkMfHqasQQKIv
h+xCLVefjbM1JVbODu4vGiMX4a88O7+DdtzJ+UrWOhf6Z8SjhJaHtaSwJQF158D+Cd1PzgLbCCcA
yXm27uG5Pm+CcqMcCK8/CLw3nwfVi/cds6sMN6eVbsJXD0oYsTmCfwexOjCmbB+ifDLR/i27zGun
+1KtOdhHHF8deeBoG2STmmYmCEhFwIxu9rV6h0IBky89n3+CMTY6i8v/ByI1Yv52KEuUPZqeULmP
W2B+PEEHx6QIs6EKoJijeyq3pIecPW2GfgQ9cCZKGNguwqZd125L62W6CnjcWx9DeUVelSPrPi3H
3spTuZ7DNiebkiuEUgvH3EaWQJKgTcslLMTDhPVyUMVNQyMHrw1mCbLpalRFHzEzjcna3LPvqfhW
IKAVWRx8yFBH28dcCC21Z6K+1aCGXgv12iDxi+H+NMPYn/ntvdK23LhbKYAiTV1LIwJPcVwMZkw5
byVOuaCtxifEeeTTpigrVjqYwoAQiBL+ZensrOn0KXaoozxtMm8tFHmYr608cnPT2qHOYDCBwteM
WTrzrPUAkWFloPPoE/I4xLtURRu2P9i1nPYM2kDA23Yn9XGvhJmuY6G68wgUutUI4+pFL9QtcjWx
I1+/rjKkfgX4oF4U8qQo69xeCSg/oge1a+gMur1LfmBpnjImmYrurgl0zGdj0ZRnBmnEW2WptZoF
nn0Ve8QrQS2xFG97cNSz7AlxboCYnv1e+/l8vsvWGpywyh93+nb3vZEJu7Frl6B0P+JMFqzg6UgW
doPm40qGM/GUM+YSxwQ6gaYdtlOlDCMGOdCd9Gbfz+I7J14JE2s2hxIdivbT8KTpqJ4sAPiqdnoG
QQUuqAG9OxcSVwpUa1eNlDJuW/xz88zjH8eN47ohpQgH/fce/Fcudg4YrXNtZO6YNOs80zHVKixL
FRHGYo8HUKQjjJ2kbrfjlj6WxHN0jUtn9kl6O0xrcniEjf1LhhZ7yfofn4yUGYZ7XsJFq8R8spQm
sVlrwm2ZybydHh/yRcBbMX4udULsbYD0u5uFiVFImR/9IUwKG3Bn9ORaq18Kkzyb7Rnrt+jcJFRh
YQ4H75Yni7Q1SqxhsfxFMwSox9UHzeWjx0/CTetZLeFro1PAu2A7Wjry/v+cAXtU9q9aoWF0BwI2
Jw+5+M6diiMOA+Y+XkHxZlN8KbQAl4w8Hdpw+KxgqeJRJCS33haLou5D/aVRgv6PR3M7QSs9Cdfo
g7UWbyvtgtB94ZeUcrCKC7RTOn/6RDlqVvGzJ4BuAovJlv1eHxLFNUvb7loaN1E0icWbh8PP7tXY
+kKi/v9DTviMnZ2s8nNQHoLHWg/ZDkQEf9nNSjukSSVhNUa/uyZ5piCypyDdSbhZhjD29fNFEEAu
ctzLIo718HW4x9SX5eBZxX0VKdUQC/ZdMtMe9/lMN/EQOXEcqVPScnY3EQg4DSVQc8tzHZKRBh1c
gwPRaS5pIVqT2iab1jPLbaO53/L18+GJjQFt0XP3q4x5N9POi5bGTDuAfWrWV6kna+x6DMuo1nl7
RRF3cK3CSgNwo6E8n/c+r9+qweDnDPRo8ZwWyy6lPLV9C61V7unNUxIYSBIluGvqqxaYMc5GEy+d
8KoCT2bdXoC/3cYnzn7RfK7S1J4abSB53uXU58G2y+tV52v89P4BkG1bTEq/gs0F7pQg7n2q0X2v
JIn3zDuAO/k60uCSUCNYye+XYQysaKuuRPEOntBc8ZfUPSvXM4bHJBUkWiwODMnYEBu/+umRx4KG
hbzY/HRWbnxcq5Dqq4bmd1ZKPqK00sXq+ISbhfeBSoH0C0RT+exKyaibLAySwhHn3MF2P9mVX/q0
KnZOFIZvdEiliuJrQ2rc/UdTnmx/e3U5+omJ1Ucd/WtcdPxcRwrlBNRPefuwi27/Miew0Kp+wukp
K7tOUpiUicQ++R29kZoRXRWDd25L08AO/KyJoM3Ty1HUnlh8/He6CVRu+l5Cab4B+Z08avU8Su86
Gy47VEXyU/AmJ6XJVWZOIpwfr9Gmg80fiQZhohyQYbBKTiaNka8ZWoxPsZ6+7XBgLS7HahU9x1AL
nFrpcOM9G7rzPXenxOfQNML9QLwdweQ4CFQXtjRL41d5/Pv5+yQTQOofvdvryKu8/i7Us5MZPplM
/cS6cCm6/iH/JpybG1sqCnVaCoxHpUALI0YFi55UYaui8FZiwig+zNdhgLdUw1I8ZE61VTFGZ08y
P81afwNXqd00mwClmXS623UB3H4ZNfmbdl9OhdkhtWbIRWLNLBNZ2YaH/o6PV06diT5K62g9o1pR
DXDDUBqn2UlmD71kc6w5eBdWHBou2wHx/zOFkrhNDN80u13QbgDVK+A3iPnzjMc/5N9fkWpM+lm1
d2QSj9krr9Skklr8XU4Jxp8lzWSi0V9GTJwV3mRyFx8NjH3EF3t4LCSb11BsZhevkkeXIE0RPG5W
3gWqnVaQfUGy+WgdZYjnp8+AOiXOHN8G+K9WkeWPQ1V/kZ3SyigeE4vaxgviUHwmZdBrZvQqzoO0
MFPC1+3Epc24HjNA+G9G1LvzFrIJhFsseFV4US/I9kz2eTMKJ0hFzDA1KiWc/nygARfbwU4moyrb
+1GLlkjFS5zQwWFVyoSFMppjiKA4g+T7fZ/jELaJgb83ZOJGFyNuEBW9h5wnrRiQgWYRa8Vj0HXB
fzdzkxPbnxAoe9PSvBz+hMdUSD7sCnJlBEToXwNhvWgIxHxtTGpkS2HmQq6CCPUVAJxidKTXerqy
mYazI4imywgV9LIaliK726RlvArHjxDcIWhk6H3yfqd2Dr9dD7Jtf4ae0LJAQimx75G3moRNth0G
uBGTJvsaEWuqGIoGOG0H4YOz89soCWQKTfLSrl1loRK08tZFZJra6amvkGGUL/AwnlEFiwaRd11s
nSBvjEhULXqdoeX6EI6SnGUmnEWp5Him9xcUHyGE0P6/vfExazipR0aYIlTXuqepx4QkOOYYuSAm
ksjT5Jke+qWWCHSpsJCXMpQGRo037HMcCCOFEhXiJvXqBtsRH5g2myusWxt1tPRe+fUNL+JhmWQu
Hf0B4VxzJX6QIgX7dco3FLjrPb7D2QmJSziaVv5dcCFsEjpqz95YBIDBEIlSD9SFn7yVwEB40+k6
F3qqZ04KO7OGvVg3sUYDrDDAMQ9Xjn2KMi3OZxSgamfCPgiJCzNzi2nwGKbNuFU2f4c6S3sjEyqo
/f1CBK+lrImOXQDVmSdwMD0nbrCkcR5CjfvMfz7ozt1QYr0N7owaXJBD+kNAmb1dk/mV3frr0dT9
TL3gZys2GOA+r88ZTW6/5sCtqah50I0wIZj5Mb2qxiS8t6h9apKR1KDZrp5ZUwMqh9DcklBaHuDZ
epmF4WzHqj6dwqq2n328D6ZXKHn8d+RNJEB1fEMBuw/E2Llq00lfhlBIf1s8vdfFiof+ej1E7c6m
O5wlevJoiBhQsjr29ZtRx+P8LuAqtlhsNiCmE6ujL7febIG6jYEzUhZRc29VkiK03IzPo/UGZpym
Mz0pmMAEazxqj31aohUXTtvPWf8ftTc2/5ncbotuiCFWG84mjhasC6S7nyLoMIll7lhk5mBEsSDJ
5p7nylR7C6kp4bOvloo1GwaLEI0tpLj4+7AcdVuO2wP7DhIQzGqBpYHNgkPrWsP87ax1qQm7019D
WgNVztXJtw2SfeLPaPX6zioXv3zkqkLgT0sWvex2u84C9e97Chv6H5PSjiEg/OZX2whIQ8s+e+yR
/Dju8eg75geSaS6AEGSvL5SqVT2v6tbqp9oTHyE6EpnKpUX9W8EBiaYhrQ9wtl8LF3JAHeJnZi9p
jJIX+leJ+CcSfKTPON69OmfMUkTwdR+wsmQfjQNsWL4N9C8wA/9VJ4Er4Bh1i31hjcS5fu+/zj11
bh10dK72JFrGzV1yBwlz0EipM+y5KBZK/rqjGrkzcaFZMQzCuzXNUsO3WhJWnZqE1lHVKt/GgwQP
IRukXkwvxtGhtvJq6xCAfyiHuBULbJ7JlHeWed93A0VoFZ1eTW0juek9mR4W6qbLeNLiVBiHKAAR
mtrZQ+MiJu5btErp/jVwdTwu3MhfToWzWaJXd1gSzCOZN1LcktihaKVPsV8hXuG3lxY3adeLi6qq
qWOx8zOuc2JI6SKQX1m4YpFI7KYX642cRbF3hdgP6rZwUmf1iwBBBzn+cGES2gBnYloGRNoZvyc6
ONWUuWrkDQAM6wZ1BnUbkiDZmBohxNjHe2h+tPWCrUhjsaNjIx1dBxTu0TMop0l1DNY4pZX6zoZx
UI2hZfcNO4eJh8AyNtwjuKjzdx6YXVuK7cvrQmoxonyVsbHVGZ5WREynLbxAzIp8ZgBlK1PJ3pu2
a37s+jblkLmYK4UygaaWcF4tXEAKx47crQtIBTpQULQ2OH+yzbhqNvZxdZT6JH3xgRC8ctGyQLUR
Y34NGiwxIGm3ldruIF7ZOyLbzAn+IZP8ocitvYy3WTpNnyOEFOc4Hy35MjhfsvLn0gQzyYXj3Fh7
PCV3nf9/5f0ZSpve1B6oKUbRdtO+TnCizirkcx2DUTgJOwlM4ckdTMXHLGfHAKZRyxRT50SNiCdI
TtZRC6X02lRnbG+CtXNl9fEznGZLt8HEnSncxCQR22NIW3/nbLWlQEHKylmLfk6PE3zg2dfkdYxR
NYlXbcWrq2kD+ybSg2GsFm9p4b46CUXS9gRj+enmlBttOEgSOV1sEneG0tvj0cI9lWxS3CFv/PLp
nmatZsM/Dz8ARFABqHVq1ovJAp1ox04XM6TOJxpXRKbgkaaIVw3imn5qni9giTv2DLIme1mW8Aid
Uo9BdEkEkdgG5Rg2aOABERGxpOJ1Z00SQI51lzJEUMfbEEQuE3McVbsm88W1CJxsuq5408q2XAmb
iJ6O9amHCBSGCyZu/3kND7c1lUsxdmy4nbqd5s6snGFEgccvhRa0v17hI+zURE1odL4vp3fbYNZP
AmH1BTa/dAiPRt5vTl4Rz0LGX5ymjkNrcjPhVx41cTjAN/qUkgZIQpPTWGlfsZiwbZTq+akSlhq9
xS0e1dlzn/JaiA3zY0jmh4KI7V1xKIrqwkLkJ1XHuf6LY+PAvixDh/4h8VN8xHWMcEG6kdi3mMJo
NI4xN9GIElSqc1N390piVn93oUE9lTFIwWMBhrjrTRMqNLS6HK5xZ/mnbLMCK5vvvCM8kba3baQN
U/2P0cRdr0a54XPgmxGClZlaczpVPolEFDtCDBbQUEvMiKXdbT+trzAtdeZzVy6t5nfY7x51Iasy
R9AfALvnxHP0q2OOWyvC8XQXztyIW7tgWatX7J3/utLYdwdGisidS6cgp589kjqWs52YZJDhRPbN
MSYneJ53NZZM94vUide1OI0TOWTeKPZhbIaMeVE1xKcRUV6kyggF5l4eDxGKG46tIzN+u6X8H8h3
pRlLCPq2zAc6wfACr9gtsFyimmzQ4PvTAzSCm/LmFmSua52w0Uk9j+82q30MPYz3GIRCzsItBDD0
xO49J7FAPEOOd5iqhY5mRuX5t4FGmksBKYSsYBtjhN5dyNbJv6zSlDBQQuURFx7tpoblGjwdsLUk
FeUIN6/ONkRZg5UmVfTf3r/tA+hd1luLOOw14oELj9GqiD5K81Mz3QW3InPjj2kuS4/whE9/BtXJ
ykC3LmmIGKjCSr/MFHfLnrQQl/e8DrT9WmqH88Va32uK2t6tuyeCZeVBoqX+PXflX81OIJBxvVC9
xQXruz/rMNf6ZHiYALQIEzbq1EebURqlTCVr/OOIsicRbSTQ2OAswC5LkWJZtM1I0fbfOaOPad+C
n+2aqfKPRIcKoRamATlo21QEGU35BEwKqoNAtfQgvHTUwCpE7EM+yJD4EQPKX6xUQDzmfa3CMFzO
79lK7sOxbNJIqyKL5lA124URvoKncNDdArjkgM6IANvI3/DC8Nhgq7g77yHdrtJ8l9aCcJl20faz
GBl9VHsOyw4LBTf5YZdynC8wHiZgn6WCHO/Xl1MftMRfh4pKdpFW1bdUs1JzxJbF/KiL+uZJakyi
Vpzjnq6iKm/Pza6149+1GchUqI1BK3L2eD7631K02apWPwa1WM9s5j6uEXCUyzq+vul9ShXTAYG/
IOvTAIvd06d/vYaZc/ndfl/SNNaRY8iaap0julmiemoftP7wCLTH6wGcKyi2TKiYpiJ/MUS5dyXv
5UoOWib+rR7UUzspcBDejloghC6+0rMG/xV3WT+NA8RVIHpeb8JK9HZXcq8RrL8fJ6++1FeuWngj
PpsCozmJW2ViTHQi3vMEOVamSnledl5s2GEMMWq3BJiOzYnY5gb0MCKm1HLWn2A9ClY3jBAdZltl
q6ci6K06aUrKb3T96maaLuXVX0n9rR+xYkP79MKZwo9NhmjKCREMYnaWX66eXXMHPPsBIUeivnG3
N7QYEXOSm/VjV/Ra1eDXGsr3KWAn02qPDRWq8XiuejGAM7pByj+odqIJKLRaC0Szm565WigfjdaB
NHkKzbo1U+ReNJtGwHR0vlJivkKnyPSDw95Etql40X2ACEsG/Uu9zFfML3ayHgC+6ve4KVNP2dRX
0EV6TADw4wPw0Bw+l24FWic12QMh+O5pqgIVfDHZFFw+JbYtMug0IluDaeGv9Hj+KfBJu1CQbSdh
y+LzIKQea0OunV/imh5Z6exelE1pfUgUOGbE4X7hHOz7UyLPD3nJqkYJohBrrP8V0t2pZjCoSaYf
3GaAWrqxxQMh0x8mTZCrHOTa3Nxnxz6ZPybt+F5ciQHbTqFaW4YvVcAk0lFf89XURVI4b2lKe5b/
b/6CR0/UadEeDJaPeXei5Kh1bkU4v/KpQzb9WWgKmP8JIupYIyBIZbSJqHVzO5H9VBrNLyaKmnK4
uUORAZnxNBC0tM9vdmoS38wA4oyBtt+GJP53nBjX1DqA6eEd+trcUiOq+DKJPsvw3t3vVQ8wQktZ
dBpDAMwcqzKcbBHnLtdOnsAAN8p7t3wRBFoVsMhHCCVomZ7+XNzHx4Qdv9JUl3iXr4/OQTCgCfLc
9Idi00AAI2w6HWItReEVuIJcoV9WCaPWD2qBsCfHIbtCmyY0W+qayz3/61gb5tqsh3K52yf2sNFH
TXc4u/7RbWsnx3GsYuaKKgevTvUniRIweTkVOE3at8Iz6dpTysBxtEYtAA8L52xrHzj0Z/ksgPwP
oVTUKzDzVESTKJhkZL9WjuYfiWP060fs973DWgfV9W3tS3oa8MpXUyOVpgU0WRubUZNN1rHEP3Po
eIQljGx32eRgpr2iDNB6y3cLse2quMOsjubUKOsoYlqJQBJ7c+PLlz78UIYG4SB84PulR8TI0idb
6jMCfQVT6aKvMuTFHQU6DVdP4IBJzu9FS9WZTn8h7hbRwZf0i+/wDfS8dGV/+bQFvaM4vR+PRiWf
MhkNbjfGiIpC0+F4Ldyd4DrnmMfejQu3w8eUpOUOjb54IiswHQ19UMMdjHtVZroSGjyPwPYHiXli
g4zJ1bigfbplpl99/IoXXKs8fO39OcQDg+eCw8knxbtDcGUUE9EZqS15tdUV8l7p8xcgy32v73QD
LVL0qqao2B8XCQJGzZRK+xsbLLvyk0vLXBd0b+H8yLKyjHNNmUcnZosM35WRwjCg4fxt4o5+0E/j
Ak9yFX0f4Nd/FoKqMRyW6MdbMMpHx0LH/EUYePks0yPqNnNjuRu24eJRu4I8QBqaYHuCosgWL2IB
JjfYCg24W2sBnVoFe6h3ha2uooSNaBIuEcChU6JMhVFJ5DypEZxCTmBS5Ixydayd1ZO8BVoaXdXz
Z/gRuBbivUH+I+GtGJKJpU/TV7AmFWF942O31BsehQ2bi6BF90AkIT3SRwbiYyv+nikwgDqesk+M
aOxvpGd52UVal0s5wlRA5k3r8qQmze6ZGgVX3LzyD7O3O13H7Yze/aUrFdJqZcJ9zIq2rxowCK5/
1Esru4WUMqSZF+KB7hzBwL/GMfOy1L8tyRcwlG285iILbPZdi45oY0L2c8/nbUtOLusra8mmTAF4
P4nZfvXRVs97va/ND5o8CHuzroR6VIZ9fEHxqgt4KYxpqRipdo4vp2V1S/hDzICMYG9KzvarlRdR
D/NJTr+ICgnfnjN6Nh1vB4a/K51g76FIeSxsI7+iGmQkzIctnZTnThlR+QTHT0/i6XL2EOPvw2hE
4oaECjl92V6dHmo5CuARxJaisZQ47ChiVUUd65/jIcAY0yExQF2lfRVjYtbgg8OnoQokugMoL+TK
Ff0wz1kmJiIPToYrQ0z4fwMVouquAim1eVKJI69dbvs8o+yltNYGDIHSvP+TW5ndOfrgOHEECxAm
fGbgH0zdA5AatrykOsaeSAhaTz9VgCSM2t2obKLFcNae1eE6reh+uSl9jqGgcq/bOfZ38ClVzA1H
Zhkj2Rrwc2kWxuKWgFlR6CsyXQLs0xRDv1ctBxJjqEOyRdKsZBJMZB5ESoEewMH0fQC0JSajeReZ
2BChmxnq5qoaigfxW2jt3WZPQd7QtQIhaTEDdZSsffPS3wQ9PnysRnz+C0w0zhQuhCGlmcZqYchh
Mb9CQvKc74UfFFTbIu1h/+hbfvX/AJQXixQJZMB8hEn0zpzi4stGOnQ3G6jCsUru4EgOXu2PEH9s
WAW3B/egrVWhJCXPJ6cT/LigadZaP/+9HqS8rsqwE+/jl+DiFY2SilKj8V650hqTM9vY3Yz1lX+e
fJebpP8qgXCmd7jXeEog4A57wyO5WQIdP4Tte7jsw6qvUF+Xqs2H68ftTN/S2lgJw3TS710bLKzq
gSa9uDoX6GD7GprGLCIS2aL72Efe1xnFhnbDMPhAoauo8LqLmhr7fm9qCRR/JBdqSONgk1uXer0x
jtD/BmAIGZ/uq8Gho5YJ2lTGH1stTbQtyllpZQnoo+Me3fEypAnrh9qrnuLg5TzYcm9JKD+v7bUu
2c6gAsZLg6xuB8rmBFMB6lStfUQMaakHvCfIMzKNABRTqYtrLQS87rhQx1oMk7zQoDCpdKjfc6Qs
dxOhTcYCoPklJf0g5IWl5o8Q1dXFCyPM2MFCcLPJ7l9ttu+TZDNyoh07vca8FMpmCvBTwbi2rWd0
8bjoTu9UThJJuZEwiuOLY5j1sufAapieUIaf7MGvFLNvzkjARDDbRUqQgF/KUekQYFTqehRJE0jV
F2x91NRVd9oqmfBZK+e5RCa/ICnc7QFGnLBvognt7ysx6Aif0aobkelv9EiiKQOLdSw5e7cXaIzi
N3SbNHnvTF5qPIMPLHz2i6HHlRe5z9WFl3u+x9MgI7fyKk0ZORteOQ69GjKKYIz0g/FRkWBfjylu
PKgkbc51b0D8uZU36teTRYWEN/INFfnwLKK3cTMlBvOZbT3akazOQxO+DQbPWvDBEdZ9hUnJkvyj
9FB0X4YlYOlKKh1i2N7QSJAHS3ayeJze1VKkDt+jTi0Cl3eu5F25AL041Q8Kh30GffAHFdKw/3CQ
kuAnFRFkdDlGF+Q6sKIk5rV83FHdfrnB2mS67xYx/fwjmcgw8c6WNc9soT08LIZNxz0hRPuY4V8t
IXUMegyHyu8gxT2Rdv6MNamM3TCXK4i6usGApAauKXVtUAK8swpOg+o8UwUl8Y6c0sxhi+U9mhQY
wcLglchL4bg7JCmYtNNEQQ/QZ2FxuPkK3ch2WpK6vY2p2ew+X1vz0J+8v5cZ936JWB7FcF3QBrjs
8FZSnzOhJCKRbXJv5y9S+5+XC1mlLv7AAJEmfWpaWG+X+wMJPuTxIlqP/nRmFx9l22J2xBxVW/+e
Y2VylYhtSooLpPrS+ULVCgE18iyRdyooHruiXUNGm3rG6SAWpqLlYK84Prj9Gk9sOx0OO5wrVeJ1
PP48EhXvDNZmpl1rYVyKnJ8DplXcg6AMuWfCdQdQOY5QaO1M2l3p2RTea26nzi2/fFHoX0DhIFJU
9/N19f8ma/YbvBOmIoUcpy6EgwGLnauErh0U36dz5Lkst+gN7SOrKDIbH6PIgW61GZf2lbsDNB4+
OrfQBSq8EfCM8ZcVIioenAbvhvWTmbApb2nSD7ZmGNzveYJRkvs8TRpUC+RxZYt7A5W5sRBuoXuz
fQ34PBK8PoGDUevr0HLKc9DCuA+HqAOppaT/O9anMbgwAgmtx2RUCwILBvDAmjBoeAvrE3AWcor6
PiB74Z8l8ZLLPahJD4rqjaHGIYJ5b1NPTXvVyw06b66Ohg34bIe4l/GrytkTspWC9R8QL3W7wwuV
KVVFvzFRBV10oXhf8Gc4S1aiK+7D49HsXyQuhdS6WfnGBR2pG8lq6yzs7KJGUrUWxrBtPhUg3U8n
ieubVLWfmohZZcHEun7F0a7bQF/GHLq7AieSCKBpLnymBaH+F8NNyTxPuSwSJHPjsi3hdLr58kDa
yssFcorlo593ACzMYgqDd0C9HVnykxnOLpLp25SDwPmCQ4y2Rc6I9ejXEFKxEhAclCPSP65qTy8B
7mBwfroaXLHUnlsPjNdOGVYzzw3VnhHYL6VnmEV0Qw/E5BHemM/8jhj8Qs+PITrCtswLu+AjtGjT
mw67/QV3b+jcVzheu28CzndBxSGpNes/V5XO4PlbmgoNx0rM5OnlXGEim7sfwuVNFYxCWviAkVys
iAljFu/PWgN+/zfRoPmcdXEbRDY9U0iiP8+6BsweqgsB2+0A0YJyy/HXtZXme86Mf7h5YfaT2FqQ
VzjZIXGc2bnRvjPR6EsM1ap6DKcIg8IICfbqvHortDkxQojFU7y+f/TruNmH4Xl7xQ65t+GbNOy/
8Y3WOsUPr/79VYTeFVSrjTjj+sD/QCPxVnG661hu+d/2F/PeM95HtXDqPnlHYS9jQYckBEyt9zsD
YR8oPfQkYuXfVSN4R9eH1tvxyKqI1d+tvskLIUAVpuIl67q8Zbytm0lgXnAS1FQM+2oK/oEhq/+O
3xKWPSur5UX9wtgnhORvbGlVSWXZ2MPYY1W89VeBWPfOA7H9mw7Y15+sfukGdLtR9QXS49TnqyDi
m+rANsniXyJ6YNYuPPNQeHCOb0FlLAgHlosEeOmortpWygdFkuIoiOS23PlkeN8ClSTA/3eSLckV
6sk4vgsqxpuspvn9GMKp1v0pFJaFuZC1ZRjXTcUqes3bMgXVkrgFiDeJQQF09KCULUQvWnbyQfqc
SCJ4qrUdpouKvETtNvoMkxkFTSRz16LFxzisdGLcugon+iEs9Nk0MMs0i2vpWL/Xx2TPfZ1fM73O
IPSA7iwDYF8jdh7LfUmNbmty11s3fR1r+NKuK+Q35RUMiScEvn2C7B0kNN8SsJX+rE0rc0zV0Etn
b6RMcOjFXV6qObuPQRcTp3fZUPfqtiLIAJ8Irx61scCDbFjxdppyeu00378kjjKSJ2iCaz6VnwTV
Y9OjABP/DPq3Dkn82XIP4QH91d/bMqESB2d01IhpkF+7uyqcJa4//kNSfmzEk1sO8R45hk4Cycbj
S1Afw3PFtjZQKM8iu5OqW2hKih6sYTRiFNbPwWMBK73B5Yx4BRVjrUzbWTbJ9YdtuhoHy8d9i6P9
rWzpgO02PCXW/tcu5qS+qjDAbQt2hSuMpRGgMW5ql9qvlKE1KY3D5n0FYSTMbg89ZxUOAoN9Lo9f
pOz3JpR2lqYSVmwqjLgfoIyLLHOsHUqQQ34pg7A6eqJYqQREt/h8cOvxe1WcgGhPq75Zs3nXVndP
8QccjrdsoMG4z61nnCbb23UZF512XHp3aQ0jUPaM9ZdtccEKQKItcrniJtaCvjH+t4gvynEjT/Is
2d3ZIrBDuDkhflkWA4aRKUkAAdciNlEBn5X7PQzL1WpMiD7R6P8e2z1CZdi9C+lS/KQq+oJCr1FJ
b8JFNRy4mcSWJG5ux9u7nfmQWarll0RXJ0joubXulrNrVLruq/FsgXA0C1mUxlMGqZ5pU5p8bYEt
aIECDg9WMfNi3gKM5Hc45rqZZ30XtIRnH54hsootTJOYFGPhGRlA5KLoZjea+jS5ho0mXOKbGLk4
9S4hLSofYBJyYTPJ9iTmG4Y2o0C7IlTMri+gVZF/AMo9GCjQ0jww20/YyW6nMrU+yC/cGxZGRphL
bvbGoDhXKnbUL+85pKrvKmq6YL3IREDC3Ez/sQ94xtRHtDTuK9C1Qwghqxsu6iYXa0weEUIbb7kj
7L2j6g/jiEvZqt5ds8o6I/O8h/4Kg4+VeDSTbgsAgTjftUxw3hy23pCxR/BQo7mnpbekMilui0cH
a0108CFVohc2TVDluMrG4DVjcVXCFATPG5hXUBmUQs3A5MqDCtNEOcDKG4nhM4lOmxyJQKezE7+6
Biy7dvsRbGWdobZRmt63RTiWcGOH99DOcLbPVSkSAZ7Gd+/+KOyfzcc6OkYbSsjBpWcob+i38txn
pPqR01XDC5qdcveEBoSKb6XLYJPiy5S39Evh9sVsI3FP82fThM9Kt4uoyfUkF8ZI8De7hLWs4/mA
+j2Lso9BV44tNz//BIm1UY4R9mf4mSD4WfzbN+fCjWvZki3VMmQ+UxSvpt9hAMMz9uy028w7dv6V
u0Sixe0Q2M1dYOcK1D5JppRgPQmqtmLMXvzsxwcptLQn1OQXFgJ3d/66QbO0fsQfyGGg1uAGxSO+
v0jAyMRBBi3sI8eeZXl5Xu9FoTYrgf5CMlJ3QRCgBcpWw0uMplhbw1qjsFtzABtCj15dYh3bTt0Z
BuTagyekY4IsO35bwCC5H1ogpKzDfrDGNXMGAuLbpVnsJGcZZkQ0qLjV+pOCjLXPvx4D2Zo8ABxo
48L9PGhivU6rUCIgEy6IMl7SzYPghLIPGKhJ5y6IbDq02dq96oXHctBGisVPVdAD4ifeixE6ZqcW
RS5Gl4jeEvuH/fMjvM7/l8lfiLa+o7DyGNySoNOi2Wy5kfW8nCPQ99moTNd2QtVrew7rpziEdR6u
u4dS5ykC19p1ZUDaZ5+g/fFtvv2ttfBLlCoywhOFTgC4sNL7mPGVnFv788/H5mVY63o5DPbPyfL7
9/dvVOj4TvYDmA4IPH6FYQmYBU7Ry7tFJNgD36QsuCjZ6tfkNQBtiLmBTRiwcdvxP2Ox701PXvVv
31ikqMp8xgHDMZ2yacTTXDLbba2dhqkGAFrpaXViTIkM3I2EOrb7OvzWuydfiZlJ4q7IVN7jMNKh
aZd4GiQxn+RSyWYmlzJEajiZ3+sN/csVDoG4FIh4HEfEmFwe7ZJDjfoJ+6iQiWBYa0xAdet4rOI/
aJKBT0iKNJwj+yUbaId8XgpQoEGpXrdF1NW7GqABxsqO50yRN5uTJfuw8m1mT98lLRQzk6Q0199B
XHOmg+gcVifdVMZwujdCXikVdXLi/3QPtcfETzMw4Kn+2RDQuevbdKsjsMQS8lrHff0qTKMrmTq2
PuTpQ+VJ3VZJgkHWFGCjftbz6XgfUK8kn1lJaadSUxUQQ9jey/d/CfSZTLOaQQjRMhZo2HE653Ho
IXqy7Ic5zgxF9gjJ8QEfoi7DEgMcPL6wWAU025zRgRYhVBghltqXCZxKXygmSGHxPYWj3/3vtfCK
dpUZ+gdcvRoBIH1Ph1s/jHKUfkOgtVdlY9ao6LQxQHIb0VWeVCWkLjSAgzxineZLot1F+WdqaGIA
bJbG4JFgmjRbqCjAxSOUttJpQgcQiXdvBFOqGq+g68znQGS7RcBiRuPxHGz/pBMcKP6zHsGul5j2
BOSenxMQCme6jgKFZHP8Jls26V+fY1VdgX1mUPYNYs9h/vuG1QA4wPWRgxCwbJRSfaFMngH5yEYO
wehX5QHheKqaMdoE0YbOoNTGWwze6C5vMrETz35XckLC5aTDYAp0GdA9YadZkRBPtdmxK2DEWhvI
I8c4QzJX/Y1y+FQN4OPpedDiULEMPJWUP9iFTLUUcRxWOucGKIAY4Re4mD48ayW/VZRh9EVMVu5q
ZeMEi6WMw9K/sFwEXi+8WMcaTrUTipWJd7bHBco3cHQUzHg3MrRKUFnDX7kOogbtKiJ2Ywwr5ChM
iiiarTxbXPMxF95EYUwgOLhV/cFVsUconf/eZjTU20EboL/SARLa98UvAFnWxfBgJqLTSTytQma8
Gybtyzs/Srk5m8meUK6WReTZagZiVuDuxIe5YfvkVSrDY3VoEI4cvCacShW1GufdL0aPUOGNLSSk
+2+6TBTn3SVAzG/tTBE4wJdsjNNKGNO1ZAMDldvPqZgckoUfqCitDnXDqmLsDOzOLDkUo1008WgV
6HFYwqX4kEBEjHP6ALUjvx6c0pYa48ArcX6cxziFxeAZJCWd/R2i9PVtg4fTJJjyKEFoxwxS/pKs
iG/08lo5yr7oMAfx3MLVQnWpcn+uwjf+sQ5nrygHHm2GT3ORnPOEniph94xpx6v3AmrtCpiBYDcY
OTLN2f721uvEeLwqRlh1KvpmlohwF7LQ+gdLuRyg84mTwsduimIYTOdPvi8E5rcwdg+lLgMVg5dC
fu+4ZS3mZEQAo7Mq3buaFC0v352bwy8h7SEr3VjyHamgNQWOl9pzFw+42tEP7afoH+3uzIbT/6IC
Wimw6XBQNzyv1COICEvD2u25HRPEVCZU2oxUP1aAwhAPgBgouju6KCPn4LE1jILRQeKznuaq2JaD
ATldWMmveEnUYgEj8eySOhMEj3t4u0QPjJqJl5Ei7ckZB/t5NVZMCX15u+n9deWEQFayVDeA1PJu
2Tt0pMHPLA/7U+NaN99x1I2lE49kzv8lSBg3EGBImtfugFl0/RXin8sAd1daim4FX9l7fGOiB1+n
JDuqeotQJsomVkF4i86hFmjihbDyJyEGVkRCv7Hl3UADEfT6XMPUHCukNuiYxvtkG1eRqX/l915d
+XWJuuDa3EnvwpeGyg6LF5jZQDlOZ+uYUg4qJkI6UP4ntibKq33bJWR8KhYZlRiIkb3lJYT/Wxur
KTRZOQ3pwJ8Gi1vDZd5NexaDOslf5/O9D156qmlE+Y4gOT4UPFD0jFPTglw7IhO/vpDQ9JrczBN3
j8SiSNLVJiC5ymUCNOVJapj3KSqZJ3wj4IGWoPtMS3dYjXwneYF5fhddCmI7JI5pMY5+RV3ezF7R
22lxmjcTvqWgD16hV2bOWYp0OhLb4NlxWpJx58xb4A5IOHc2T4+dRWUC9neN1Bc+WJ2AX24YDKf3
SyUXHA7tleDdrNLFuKFyLeD4fBkSSXQSnVsGuyy3KKyRwDdZzuTBvIOJet9UPAkGh93+uCKEzfwX
KolJGznuHGc3SZoD3yAvIgewMqhwjYbnZYW7EMyS+zI0M8ixgnW3cIHkOXvIh27Kw8bPAv9VQSkN
UifsTEAttjf2p/TqAP/ADVns8ibqcD57ZsDi32SjIlKO9zRNfMS+Cr6I5Hypq9VOueE4kVDQ0yKm
3IrCeKIWTu46QGyNMA+59x6E/5cdNB1SvBmypL3x4tWuXg0fEAe6YUnpYel9eSpyTh+C0zFi/WD9
Dfa5I61L8SSJj2keemVUJuVXTf24B+BmbApUhV33BiRbmzOAG9xQvRMeRvJ7A6vTsVMmOYsyWTYS
1/4Tda7Vvlu/24RGRIRrfIDWQ4ts751y6qtTHIxS16cd8gQM9rvZ/4ppJoXAc/7e6cBRMuiXrsc/
CHlifMXBszLa5tDaUEeudS34UwaafrhtsZGNOl+0lY4G6+/bpEZ9h6Pfxhk0DeGI/wHJ4ySiG1+5
eHkpkbMZUbd19Yr/aNruw/P0s+xGZPZAfG7VLYwRRBv6jsqDbHqMob5ysheg+iqGIqzH2GrHc68h
QiBO/dAEaQGvPoIbPKiQW8bHK2dcZ3qLNzc30F3AFKEH77asZzbv0ZMVQoJIOV+qrK99PFJ6CZCs
cGa3d2doLgd8ziYMJBQ60gRXWD/Ev5ELWkK+hCOfoenUJDdNuy98c2TX+wxsIzxibyycUngYEUZh
2YDMZCUPvxgOJp4gzV1VajJl06kMTh1qfpasgGzo2us/8P4Cv//FTRIIUCnG0xD+Ixae+hlJBAeD
XDZaJodLeYP8FcmvrxfV7D7E2qO+x3nqtG+QzQWq+XKKmrzNxuabFsYyjR6rufPuLAQ84dLi7MjV
y+ogKw6DoNDJbnc01Ki7RJanPSfMDwH+5JqYHONebW7qAURbDHYTjYlexkvDTLvn+JBtmMH9bL6c
VT5VA51sECch4VFp6w5iKEFfM+MtzU9voBUQ59XK5jAfGwAwvq0IxtPxB8MYtOjdI3WHbRJOgFFM
RCu2CzNm5BthrINNk6FiAGEJycDkWXmURDlIXxlIAnvwrmSQN+4OZK/FRWhqi3wMPc3U2w7SNluL
DWmsuLuWmJip+cklea9G+TCzpuppYiFPsWNCRybBs7qIXKySf8Rxq/0Pc1LwcvtDhS9s+pYwh071
Aku6dtdDUAPEWOcJdRIyfVODLv/XyTN0c73UhvGU+hG3Rgvq84xWndv9uk7RZ1i6fS1kVYMFrsQD
c9E4u5K3/qeCVeYciK67xPl3i+k2GooSmhgBnt2ru+jem4xIO8d7FT89eIS3X/vekRwqtucIVQwK
MHbtWPoAIJonSjlbk4nGuZcjRUg1GSrWZSf4XqeTvF1vDPng8FaRdx2BOde5OeOEsHp3Lc1GIUr3
74TIzVUn7+oLnylk6plyNZjweJmhqmxBBv/zFhPkczHSEMckajM7gKHA948jiA15oPENKFscuKYG
+jx3ugnSDMW9Ag57EzIXCrLLTNYyWsSzs8XVtn6q80a/FI4ME6bmwHgZHyE/gz7DtGY/JQsB71Yc
oA/VcxhVNmJTj/3ViAqeVHtTKo87fYWzQtIb0VKId9jvEFgN5uXbAsBTbxKwn1mZaj0MOjM9g1pU
Y8WlG0CRcW+yZBQ+3NGr4AZs6uvgNt8o/1YPNHhO3YWAnQB5FU+ErB3JFg33f91aNIYKgjtZHDu/
nImHyu1Y1tdVBgl/4E4cRZpO+HRZSk1EtfueoJvMPJFnpdgvKJs4AfCOC/iPynkQsUlvk4RafLDI
HN4khRwrSJhBBcd+gIe+we/vIhXfHnCikUKwQuegS6AfRy3LS6HbgCEcq3CFYmi3pGm93++hKpiK
e8RQgmqKQPhtOoBwk28jbyTUEaR13GTF4IPeIqclPbYHciKNYoZeN7Bxt/th6W6agKsnXvpKB7pC
vxDi56Jv7dUynSrX+6S+Ok3ovqmyptBPjntr0lHuXwsXMdh95XQkweIm7zL4Zxokg57UVgoQbBOm
nMbeM0Dic37WDLoBnNk3REhZWWcuvyWB9A7X5TE7FsfQpejVDwzYptguslSuWNnMZtXFusS7KwXg
a7e7q+HPMBTTVESAqYoXrt+2MzQV9KCIVWQI3ZlVpyP4Zv+icy2jk9QpG1PZAnKgxb4slsbpzzBh
h7aU8Ul/H6+kXFmzK3eNlE7WEUkQuvLNWIbWx07xrTqBZaQlJ+uUpGNwmKM5bxZeX17eW2hU0CXA
XUePoIfvQG95p5/n0dZAUTrMaEYDpU224Q8dM23CiFJVjhQTd0sPF+CmNp1iwuVkfxAb6Rcfhj08
coiuXb4QjLE1JTUgbBNRJ1aYhnN5L9s9ABI+Xob+wejciuEQpYM72HbG6I5lsVQtJODfUNDTDdeC
NngQFiRJLXrPO4gq+Y8QEetWsSClJBkZ8vSmoYsoH1aOLTDiCuUjoKq/TFaMNna8QamWY2hFORDn
Kv//RaFVU/M3vc5HqkRB+ZUW8g31fFb4ckM6PV25KjLXXTT1jmNIZFGmca7y/kVxmTvZcCS2MwIe
kuMfaG3bDmibDAfsrXufQrRW0LPHsTyHS/E79XRivK6izNYzWfgV9BqflnGpW1WZ35AaV8YH38ke
TkP43v2gBnaU/tP8FzudbA2uYslRxFM7u0uvaHSAjCReEnV18JlEjH5bnB0CyMf4gcvdL7U6Zpd9
5iot02C5YO1jZCIGzOFowWEh/Mzfh/VFlj3sbqpz0LNSrpVGLeKVYkwQh4Adj8ydlWNFbemOPKJV
5ftfpp7M2elITQaLSJB6BNijhK9rdDkGZvCnZzQzluFvwPtAvTBW92vwiwt5DB4jYlK/JVkKWsAW
I+Jr3lzjKsw+5LIAlm2b1PMmU5prxLoVte7+7BArYFDtuFKSB1R2wxkpIEs3AOtMkvufGZdvMXi7
G/+vU5O5Kqidbhs/Q/67j0oZvKajpWV/rDhuhKssNzgdbhMQW/wS1zS5jwod603VOLD8EPCwj15B
RkwsObOOefzDO4BrzRsUYUTojJeUFO+eZT+Eli81Op67jFyhPLk2QAEo74baYtiX37XRE2TJ4JJ3
RNi6RZ+cYFXTiuSG/GA/0TC0irVpXjMFgHHX0l9jMfZg5zoDY8m1gbhFj8c9zpNlM2kGpx7DCsFx
mSY4x/UR0nZdPynceQ7rUjq4FJrWjLtIJVtQJo4RU4UWJY0hSx7vqW09zwjo4YZZYVPdp/0yKVgV
eHKnWcAk7kjuz9qAnGEwHZ16wDNd4ymjpwfAECNesMZreDG+EI6DHnVHfKapP2A+VY0tUTGtKTBm
CJtNP6AFqnwPiN9fwPBoyCBfNDYNgBT3njTLCca1BQIlNvKKaf594J+W8nWika6MTw9mfx/VbJk8
qBpCTzYrx9WFTyqK+rBjA94VzP6fnV1TY+6PmCdpQVg7a4cgsjmGJ6a6dVjG7uG3fH9p7Qz0R3Pn
n5INIbnLs6WTH3lNAsv7M8Lq91E4Mg0lNDDaKJQN6v/Dfs8DnNUhEBNUA1HVmy4KQLA416HyFUfn
nzInFpTMYiywbbbJiiYTzT7BZ/IxMAPgid+vBaCp7NsO/OGSQeyZdk1xVmznBby0gtUjbCL0uxTq
HCoktu1B71fbFMCPr1iwFNOlvY6yCZmTAmDL9atOloWRjsoeB4RQd2w8Dx37j/LFe3q/DAdw56MX
MJx0kPWECcpagSK0DOBntsPx4c4LCKzeEjABfuE/GJs73naDRoHmJDg72sR026+GVTBqw3kvmSHC
TLvOAL4jL8JOBENZEnO/lL5IK6VNo7znNNALlyjEQ624nG8YZfWSvgJt9JzRi1bYdeutxfUwOtI+
qhzXz6YURDeaady718gq6SvkktrowAqv0PdVeVqY6eadILpKSqKqBmgTYjDqzkWL0SNzzAaoV3Fk
FeDntjxx7FH+66F2K48pt/nvUUbokTU/vPmY4/ExIpzSYTy4wpKl5L1/Kt96kMhIoJJZZTChRVlK
kjXakufTZ9jBOvbn+MBxFbTFsaac7ug3stws3VqWHvMGaFWSNahtDQY9cm+TwWEkD9uwnbimZljW
+i36t3WNjVJ64nyN1XzSbBz6liaapbtw95M4wdq4xRrdUUaGwLQ44bF5Z5ezaj/E5YZloglA9ErQ
fJ0xxBUxj8qkkfr4a9dTJIdIvEpADIAOmgHj++2HISdLtPVTT9j4iRPGozzBQ/O5PiEG5EDzSVb2
CxQjg9QKi2BPcEKurHWhqjCSowVcKhw/z5HCaSLBXPM6KTeOr/c3EXQ78LwihNSPVQawo82hvMWb
zYUWcP7gQNRYW9YX4QlSfgWbfeSPIBdzSiQCOFAF/RTWzqvLqpEfvgM4ox/7+g3muGL+DtBEROGO
+MejdXiWAzSLtdXTB8TRdNd6M9VQrrIceAj4bSdkegaNbJ+BY/b2Twir2KQttOVKQxgxe2bk1JHx
c5ZFrQO6rseT/qA4xbxG880VWK821qEQhHpklydM887AaV16bfkaBml5f+Q7OO+grNGk4qQfOeCn
b0h+y90clmJNtk6YWV1LIogRZyz76sEpvq+F2PJlQSYVpHpnAY4l+phxm6ir9Ll/lGZXgM+9WNNb
eSSLtWZ3E7v8KxisHJXGbw/3sDmqzpqfxnnJPDhre8LSAtvCMoGOrB9YnC6wis39oTrF92Klpfce
cCdoPd2Gxuc/WYJmeqf28WEtQ0vUvKv7QKeaRtHgf4v7j+3UkFtoLaEfxSnv2GFQHXIeEYVa2pbj
3rNaGJfe8pFdYNCwPEvkp28exkT2YxcmGvpcX/a3GjxM5L9ug/XGN3nh2yptIfpq4DJkSoKzi3QR
17mD7uQQjkYBqXmph2vncGAR8rVMbn7OFWxWq3Xpw2akUQBcs/gpik9KRt9//bIOAt3xxelwW96K
4BV7ajg02V6ArDSchE9ujZiDneHh0GYElD9YQ5rtBVVmmqMAdgvknZNk0jxtxNa2VvX3dyo2hGPK
EHCfqXCDJSn/lflJtPBmfw/7IcnTTRe33LEJZQVhyXJRL+SxCeg1pQgZLoKKSROQPEiSoDf1WjJl
NGsAGZEt96O6eoBhw8YOKdxQWdPe3Xxnhw950FEt3gShiavKkqWN5AvgCg8A8mcLTx+HqmqFuKRu
fChpkf1fT9ibv6zWSySU7g5KV+7JaNo2NooXir/4osEzT0cq5/OMsi73wAohvcPDFu0gHDTVCUUQ
h+qRaXjDN7w/+G7jdV/ysRyrXy2IFxUgc0fVEfUJ3IrAGgVpPGDU7CHSsPHCUsImcEE88T2BnY6D
vOBzyREkYJacZdCVx8r/uIbdYox5qzDHf2a7PD90vEo13dph0JaHOG37BtK0jMDrkO0lxg5ZUOeM
FeBMygQqN7R4s3u789+bCH6Ey0P6wnqX4BqB2wnlbNZFzU0MwAndwdiuGqcqegVC7m2DnsZe4qCL
IO9d4FaNnEky59f8k+GzovOF+xCVo/mlQ0rkAPipvROEbMCan/JJHlTXeYpu0zfRkkCLB855JPmk
FcbRTI+/YyXeXoduQYwZcQPaE0kqq8MPhh2VeDm+BvRoeb+4B1mydn3Hc6EeS2oyaik+SvMEXx7e
dvFInRBwa2VAyq2bLNl+E4gPux0KGyxoyTNiwUjbasGviq6CYev7kObkw06vEIphYNCrpzxiOD94
3q7u/H5jctENjOe5yvB1rFfJnJAHRa6MgUiHsNQ3iaw61j0iBeQ7hsJd2RzHGWtq5GpGlBg7/scW
Ias4uGBoKMfYiina9B3cOJQy0f96PzLMsBhAYo+F8aq8ZN8pD71KhYrclqWHihUgQcDFGO/tpFkN
6hdmg7ac10WwXToIGDqoQaDi3vmwvzJPQKQNiCr4Uype6n6/yAB50JtuBcGea+psr6lKthfUnDUu
UsdrJP1APHFBMSqKSJ+v0zEuhYULAoqEFZz5DwKINhcBY7tp0MvxMbAcwZb3tKYtC+JQbjjkz3K7
tFxu23LTIy+kyTgu5e7dduBa7bHBDweSVXgCxfDRgjctsr+Cp51672W5T0hfbGzYumz7zDAjDIHl
11xH1aSQTAEb1FDmY+gysv1BB35YPaSLtq+jgu5FjKoLzjUtSuTouJwegQRx8ZAisX+Y0Rv44Fsv
PMTjVwlHTjDhVzINr4iEPz6hllFvTRZ8VqZuRoSfzmBCR/y+K9NqFCBn3xIlyLox03lWw4aQ+hyf
vwoutY3sktbfswXZn4H/LodpV8n5fmvc5iG29fUA6lQGgKXSMJ2z2hIevlmepxB6xXvWczdorBt9
CzyG29kocw4phIYja434l9df8Eoy0AEfb4gDiVwS1TDyKz5R07isrcZb5WxETc4Jt7rjqkY9NzlB
uQ0keuMI3OVstTfYXjg3seRIFluO8bPeTOaSCSUo3iKbSj7X9+RLYOIr7HLt7LHmMhmWpIwcuujm
nS7A5RTaO/xGzLJ0Ac5KBrLSTCNCWIF9DS/EJ0jr5I+w8RWBlezB/TjPRP0ON93CzmCBhkQxuCBo
3zBbA67ahLIGZNlVutT8S8hbmflQspDUWiPRaMT6AKS6MmpwEZSXkjIgbM3YBefxpW3v+DQWWks8
qAS/ejlTiMkgOZN8joWPGBcfaXP8NWvOmCHZiW+UdSO2mrRWRJ2VkXRiYbrAafEWhjJHniPg0fzZ
X3HG54MxGxs5CKOHNFHaU49BobOIzaG3hofuWV4kFjzwQsWEAngGZZMaHCIC8kghh7PjGvf7Pl5U
5aPx4ZGePkPrXtOZ8cif1tQAjak5c0X3pydROYape+YsZp4MzDsW90WwAyx1SHTSuKiUSSteWSSf
vby2Qp8tLsIwSKxL7WEpIAdo9+3RHww04fMubazExXwCBMPTRarWaSEWNKB8KbHjMKNjjv/64oXO
HJ6IYRk4axQ6LTgvp5OhQAbG8TIp4gU510UD9OPZ51dCFR9r/CRLZBPzuheHdmep9ZlnvTRnm/DQ
czRRmZVxzhjM7ASBS0fkAWvAqT2x4DNY6ct54eP1GbALCfq8alPeXWwSP4vmK+lhB8yVxguHKvsf
jAu9Ato/kI8b54Jrk3xwxwWx6zQdcGAE/ntzSm937psGFhj+JB5EaCV7sqCFUAjN1ufK0zl3URq3
4VlbDf0LWwaa8tb2Rgl3GCD86yp5nY0iaAWr8G2jatK+DDbjuNk+tk9BkSuyw2ibCJJP3tdLp+6I
jJqdoyoBqJ4f2iUQLhnkeD9XFK++nSLgGmuzUWzFxWXco9W55IX44j2O1aQD4U6F6gRQ2x9kJb6r
t3agNoD/17AntRTgJw6u0dzNQqlJ7Ic3GrY/iVSazIrnrCagZU0V0REwduEVbmalA+nKTXWLBPQp
8ojcRjdiYoZeduLbbClVvjAky+1233tsMdvl1n0VJauxG3JteXNGA6FDULkr33bLS9UU7S2fwkIV
Weox03QweQUwB+pnfT/8++9GoLgWgoPSmL9wm+zsv/Kmv3IZXX2Z7pgK93bUl+OXLNYQ5qxgoY9J
jUcKenw5FHSQ64cpMaBCsvHZOg0O+XXgRfkzxRAlvSVxjt8zxX68HQfRsIkzazib5dSF+uzKCzKp
eIj+Oaookx5tCGeneJdk8xhaPJuJj/bibmscxJs5h2mII4t1MfWGcjd6V64RD7rO12/GgtN57Lth
n7tekjZVVIGJ5MGDXPAm6Fa0y62rUadNTZmc/u56DeVOCUw/nFUyRpSm780OTxaVOkLRJrvehqq2
AYsvbrQovl8HuCtHKsjmmGFcJdUGwRkoVTn6FGXk6kuXEFdaUsz5ezXSWqrFlShasP9RbRUo5u36
MjUZ+v9QgAbseo/BUI7hj7B5iTAweRhA3g5kq0Nuq9SlscvbHF5TKX95ZYO+/yxY4XfJl5n3fBYj
j2G5fnLG+VnuNluMNtcPi6SDk4JMaDHPO2+kIqWqIH1MVMMj4qKzH6Jw8izOXLJaAQjVNvQVPGvz
HvHDvp8/kiqG3BPsq1mPMIxbVJu2OKJ3PBbdzb/3Elk5eW1An5Dwyvv39EqrrePvTvch4PTEBktj
mUJFZkYnWPbu70hZFNAb4eH74ppaL6eHFNdYABj/JRYUV4SlaFU702sTc5QHe8Tx8XNfmbc+ASlZ
VnWEk6ieu6TWy/grQ1MouOg9q73cS34CRBIPzaFRUGIF0d9Yp6q15dOCbvH+gc46Q6wSAS3uejxT
97OzYognBp3wiedj/ujBotsj/RjbYt2HB5keKjls3+8N8cZWQ8s3cfbNmn/ti2E/vAb3yOUjSZI5
ISNGpsZ0HiS4bViYcbSS+JxU9LTC+v6yI5KnoGcJnHcyjtK+qtdRRtTJDZMSs9nA1L7aGYlc4nzv
Nd2uu5qXLaZLs+U5MXeGG95qeAEDkjqZ3X166GWT49rKXQvCrWqH0CO33xjjHRMPwYNJ0Uvd2qFE
+M6jYar+SIcIWG1aj4vGiuBMvSKaIq4sx+SnLhxmdK65umRGOeBphH254R8an9FaHZuMl03BVkXN
5b6F5qXwXBz+3DJld51d0Kghm16UF3fS7sR2lyVcKSfUZ1l+Ps5Hd+Sw/GJjiEPt6y1tUOu/b1NC
3dcRTMQqac+EKZgZlF+GXwnCWVqNar2jLGjgRp53oADv7Z/MS005VUeoWtnts5DSl56eR/rXUU7g
OVpsV4BfJ4BESlFn9gEeUs45rhSfKmbB5nYqRgnfxbeOm29WbEe5wulGLDzpahvWlA8e1Fxh9SyP
ErUCB233Sv6ZaVgiQOv9Aiu5Xqfzdw/jkKJvXn7SKaLeR+asMgtSJNUDwK+nuFFyYQY6F7PR8bPI
I0AkGOmdrPiOwt4N1jgm/69qQC8z21JjKyJYuKsLhNVdSgsb6Lvsqlw22NlePOe/8NnVvLBB/K2/
+7/IUKNVets6wHKtOc5fByRIQRnxuuJujE4r50kOTRIzsL+NDScwui2HgW8r4S59mtkrekt4NNPK
jE0ZSweFp55OG+S15Q9F8Ft71M8DLPINC2g9xxFu/f4cS2hf3E6vgruQHbkfSLSJ5b07YI0wWrLJ
Xrw5P8k4frOY1tYir85R30nRGejh7EYsm1wAwgUrUJsSfX7VjstVBwUIYbz7+sPRjnpXrnZD63GT
7ACIBWMPQ6GjDtcoM7cPvEdupd7jeSHm53/HnHuVEiJWPX+r8iOQUgNhl8vY+8O2hYPukz/xTVrm
n8mt31MOzUfk+6+cK3e3RwsXyqXFjSvitUI82Hl9Jkcl+mGbnmdnZdu8zXW5FB2RMM5MbJgvL9mH
ZeWj/AbFwPBqmAAHFF0mUcdFo5oIxcsLGDgVkD2HwCzPdCHjP0QeIAOVGuhk48OtVCS5AumDMHdv
6JxrrAKUITMejJbBKj6fhl/is81OIuqQabOu9QuwwPOevRsp+w/EJYIaKrOd3CMtY5YsdDCCWXsX
Voli4ULPmHVUIS9Cak98PuzW3wiXzBvnv15H8CalTvhjkxiGNPBQrvU0YiMAMm5ZjGSmw5JRKI+A
IUDThRzWFdMxpB90wJUcPZf4fDd+WW1a0x8jjhYr1KRKlamFzX2Y2JYSjKpbPEu8AjkVLXW2/QGY
LfCqji0yCrHmc2wOLCnlP5TtqU5D62GELqRQKkpf2SyPirsgvDPnT1K3ldNCVE0PpPeZuE7XqAhq
s2jKOzoGI+oR42jVdjQXMb7ySV5RziEP6Bj0HEGFowklNLqRixE8fXMhV5QM2sZ8QMz4gMJp16ui
axfiosfvZwpcaTex7DDXL7fO0z/zzGGPRxZ2L+o1TTgzlfJSaJDNhFTKSdwyhx3x05jcgyO8qe6R
GD8BNUYUBim3O3W7dOW8ZC9LZdBXQTyJrt8bGGnysgglflWdpJlf+eEzICpnSAwVv22k+L/51dkD
0Ah+Nz3hCzkziEfUMS6plj6NI1n3o34zCidqbZ/40Dx2jslSuO8cBf2LCNbNTpyDrfkHcy+XBi4D
t9/S1naqJgqyzJoHiY0QfAgGiIV5aZYruUPo6F2ASfb2MVgTMxfuVtB0YLS41Z3sx2f58PF4CDZ9
tfhYV26QUMk8d7SCXWXXjh9cO8cfiY14OQ+beDN6ybuuz0M0fy8PIxWupNZgv4Oj/5Ga0TnDCeuy
YpVHxWOO90SF4pkNQrxAURl/eUss8hCZF0LRWPorVKmRrF6PhYCBDFv8dZQNY9WtxUbTZJaC+e2I
yLrlUfukLJE74XCF2KNdxHkkfxhmfz6sp9IQ+UF4P6nzfyb0sdOugEIBdUx9JhVqTSvDn9sWtiCK
0BAdystsu1SwwMr/bujrUvPKcl8Ish4VuCKMdrPyPsxkqqp0JNWUaTLkMypulmEiAJRWiTTpoaU+
OgFoYQGTs0EZnz4ESbtN0giQUy+P77ELzyWNiw/nLKfoen36Nhq0BasRFaTm0L+kSBomQuRv4Uo4
lkxsazCfMhLcl8CsnllHtJmwav+bJA8/dfySQjDueir5uN7tKKX4tOIvRhm0B1ewItzA4eSwEHHn
6HJMkJ2BexN8uf6uvJSfR1IbCL+xeqxtGSR1mHwIT3/jVOS6xjkm/kqAgWTKeO6iJFHbft5Q35sb
n11a/VOj1kDJYwDdQJPoMmtNsk44hiqbfE11K9qCZyLGsbTrPQQUC2EY2pmVvvGBwQzm3qEQHi9D
LGACRW+6hJQjFrljBzlLM2yUbO0jhwNyGp3eRAKjIUzEeo6F6+9M0ts9wuPIVHbYsckZP3BUyAOr
k6PDsZiZKavfPADcS6Y1eP+KP/ReeqUIlQU73zml56rs2mKktIsN99q7RgdX4gijbEJRWzB4NrD3
fiHk90Zhnon/QgiYpyWasZCP/nOPuTc/+pv2Lj/azVwMrjppA0Zjk4IJYiKb5TdhHQuCjZG2aja7
Z4i5UUPr2wrz1QMp8zUAehQWRHPxKPDHuqguysCrjME8gkwbsGAkSA6MAt7h8dAqjNI+3Lz8Zj8O
VgzxPUamrLVd0dDoJrQT15gT4iwrxO4jM3aLRfHId7CaBx8D1hk0CSZ97jMERmTyk1/dzZ5dv+JB
1YR6lRgwI8P9rTAo7h27Ye7zBsO9ndwSwOs9717nU8+oEoHIvmDHdbFExrYqhBmRFw6XIcgM59j6
jQbJ2OzH+yjqeBIiK15lLSK2WJ48lJo/2fqy3Xzkjen83Qdgxc27612TKRBm0Mr9bR2rujME8bT3
N/ckT65pjP3p2cb5mjSyWWHIwxn0O0YcY9scyS6tkhycbrCQBXS4nQWEhZRTPLA90crOZMaUQGUc
DFsgFFTWPpteUI7VUKBSwHfjslwxdXowqQk0JJKuRvdk2Ejts++0TDNZpdOETzDuX39LroNwpUug
P9thdLkpelbiqDP3lgGMJze2d+X6esyRnZzCCwZ8jOrYgENJF/j4laYHKD9zHwZAAv22rjois1XX
kPzA6AzjMeB4CQrSsjBMoVpj6ZGx2VVkTsjn6MdWZaKDAK6//fq+PkMbnulSFixiCUhL9SbciWHT
57Lwklr8/J8OzHRDXPSsuZe0A30EZte4sD3Jr5LKx3sowWLMxxIJ6KhaBbtXkONEs15M4MN0KSob
QVMmX09eEoAn3DO4tp96h+ajIspFIyXgJo+Jl9dy+pfNCiKkMzwwex8lukMbBPzy9SNd5NzqB3rC
DEZq/0KZlqCTBiHdHaZ2UbtHsLcNybswyVVPfpfVWhYrClWREl94+oXOBfv+7gROuiNeoJ8bnN9F
i7RpDAptJW2n2LrK927pQKFZFdqv64MRmQvgx4rOle3fhC/1/ALcPaY67HDb9WC5rBcoYAYblL+E
EEmflq73oL/T9F3cKFgkyMvcmms7fhMcRAdcNio09vYdrNaCy/FP0ZByutCSuFZLY6JieRBmaXPM
lXRCgSaGbQ9hO4Y2u07BlbbihZ3W5BlZdHnD7PJjonqZ+Q21PJB5wfQLj3/HtaT+GJBslEnqO3CB
4urnSxdJUiQNWsF5LKeXHY4hUg78os/hJrSRg+yLfOvj04LK5I4MSh+vFnlxDdZGMNOu9zWoJ2cs
yKE92OGfP9lqJnkAWtna7AXHwOBkz21baM0FMu2SPFVjMpkmeLWT266RJHNqmJ4ZjrF7C01/w0cL
b/RftLsU2l/tWkS0sRY+dKdF4zEKB68yrZ0xu0PB3y9d3C4kNLVz+hxu9HvO0wP02DDNWsUFwU61
k6t2gDw3xaa8NPm29w/MnKz6CnN+DanS8sKQNgqniGiKYkR9meiKxS2U3oYMOCg8ueYXmSyGnNzA
gBdM6uKmfRZ0aQb/yh7XyC/rMpWgFOu7+jzpQ0WynB2SMyO+fWDirgTEenI5aiDG9M4J4Wgrrufz
vw+OZFeapWcMuLfniuYg7Ifjb4rLz0Hao8S+Dl3uBoTXy0Q9f2IniZJdSU32TAFmCA5HRSMNRqaj
/5++GwtevtSsS+R1U1Lp1/6mM+luuTwp2uXhtA+lswyYV6Pqx0fDvTTlI/XBHHPgzrfS+kkaHpJ0
rnnqmJBqCW92L8RkDao5oEqbqqZ4VQ65xrnkFCF/QrfP577k+eekCWVHzFUr7KeQiHV1HZc9PMr9
LGnScTJD3HFJ0YCKMDIluiEbbJbxvmk+oqpOCoXKKyDogJGQQLoZET19CWbmk5+X+baIBPwVgVce
c4wjESpGGW7C9TFpUqUiiXq112Vfm3Emanfcx3WXREvdsL7JkvnuAz2Rp6DZFTMbMOTqSMbh0uSr
QWbO9LERny3SPGEP1HEs/klRQ5E/x3EBTMISTOYmmZbflaXPAHGQo8/Qx6vaxbXHosaeMPbEZ5/+
EE0PmLMSfKSNK9hfSp5exkwnsGCEcj3hC/qK+JbheXwlrn79fxirc+gBSh1+9TQstDujF1J3LJSg
5rPoU6gIe9aWRsY9n2CPoviKAGnrC6n/bQPNnRPI6N1GQ6qXDSrqBtqiODfoR7hKCTS/bQtn5oJk
bb6OxgTEuj1P/r3mYztSEh15kC3T2mONTAM/otC19HvxNymgPpIDAarLo9WFksBBnE8ivEERuWSH
T+r3XFhkgiK6hVvioSftVwEIyLsTUVMF8WCppUjgRgPd2FuUB9nqyS3G+YduhxgwB3WOHX1yLOUF
5oO5e/K9IXiKwENe2aRTiRszPKUqVfmeRfjsUWOwr96enQH9VsGU9boYjRsaymXrZUeQwnYGZ1VT
meQvfqZR2lIDT9SK6r0dbX/EdKQDjTjG9bbjzvJZG+nDgGoPzXTbQV6ORBB6XwMTQjWrZi9vxl3l
I89FKYv38sqpMnML3FNAEUv61wsJoPvE5Zx12+pdIGF4SFteGJHvcls0rumWtfbS0/P/bNFIvsn9
TW1QJ4KD+ZEE8LbSXt+fen3Ndfd6gxeMsVuLVKJZOLgnN/ndE+j6O2cISXJXh3tCZMMrH0wI8UxR
ZTr+HX4OWv+dq+x5HiotVKD74JiIoeuL1yi/3daZqD/5r8oecQQIJJAG9jUo9PAh0HUWn+eHIPJ8
4ktVadMvb/RV2VZHM2jL2OE8Pz2hbe3NR5RgGFlK0jt5R6TATCWVOd61uQ6WjJKOJpmQIkjii3b9
nNa2CNA+3/oHmvBhFFJ5slmlVx4Kwop8o8h+wNVzHztf0iFE4t/JtZ6i2VmgiYX3b3OHq3QnmQTU
O4CHy3Js+5THZm8gIzEkG1+PRhNUnGDCNeiPvdrVAwTydafN3EgH0umfm6pLj97rtjGChH0e16wc
Szx6uuID7SpXdNKCOhoCmnzK0O7tqtRSe1ZWkNToO6KJ46qQisYaWcJRU8mZaLVh16+gk7IS+BDP
rsOPzEEyEf70qj16zIMYV+YtTT05e/Wp813/EjU25Eu0J/elcDf/yP/0fgJov8oWXaNGHiHXbYfW
m6Ih/xbHZy0k3TzefgGmyCiSYpg8af6vcCVS2BNkoCaYvrkVs9rRfhobOM+JJj/x8h2vxcevM3oD
VKNCgQioq9EefGNpg4awieMqQ78A2F5jTEml2AVcOtMeqwkoqmYOUK/m2bx29579gQ+B8bBjDcBx
82qRywv0Bv5p5qxpvJdXzARd6sI+Vcbgma8Q6n1M3ilrQxY1gVMxdPoFpqDmWzZR7g1L7p0ZglVx
I5a27WlEPvS6OSgGuoDlZmWaYGa9qdCHk5Igh1e5gMmghTl9bx1Jhclf79LLbVJ5RLAb4qmdZNKM
mSyBuNLrMOLVXcxYwnJE/SbL1rros0i1s2z8oqHUMD5t3H+sFgAy33T/C3RjTlHQ04OKZq32qcf4
VeuEEkfX5fCcVMVLrsDV3r5HJegn0KcCGOGfzv0TTXNDjBiisXlrXruMZXf5e6GUYJXLD+hb1i0p
ZcxUaYDgyXAcLpfFtAElZ2RvkEr7yjOnx3MbnyTq1QIgnb/+u3uQQKqeFf80xCCuGItm3ZK1Tggo
LdgeI14hnEUUlK22ATwpVk3CqJgoFLIVgdjpVy7KYPy/Q9v1mrBHnODFchk8bXwxJtrdjHNc4fNr
E77iTekydkxrMPFC7j4wn/xWaM0tOtOerbLh2rzaRP6fkLy5zdLy3r91AcxFCs9icMtV76SKwSW4
9fDMrKHZYYQsSFpm9i1y7u1m6C7JqkC2p0d2seEC8JfKCujvb6Td1V0yHpvtZF3Wjy8njoiOPkQh
WCakBOWLw6AS6zg7ieUK0GoDcfFBookeQ/PEOjijYS3tHnJYmu7RxITtGTyIeGwdfXlZPxA3SXWa
nUOQ7flhIl4lg3fvS2uWCwaEaayadZ/mv5lDisIwD8l3w3LtVlcbAqYtY12HGbR9NL6/GBaFDeC/
c++vXP+vjZJebZjZCL0KAqiy1F0FmPIlELVQ0XVXthuL7OANTCvQrzRYp3xGGa3jTB8+t8guH6pq
fBFoj2t8z/Cbmvw95GlOVMUoaog+XuJIvlPN+B9ZTRXf5w7j60uZby4SuXe8HxK9qhFJ5eGL1X3z
4vtLkksWrdAOd8kMe301SJKrzVut4IzkW713n2U5leUuIKAJ84JyXjZrPkml7LZVB1MKKG2Z/Cqy
yi6t2M9HcUJ589ISOqMFiisn04o7/yMxa3j4wxA0P4wnJPF7hnqO/CjRPmej0ShlPCsNYp7D9Q4m
AUafxlNNuzpVA2F/n7rXYJI7Aqb+g5CY7c/dLGfSzuJRE1vHbY+iaq3ELDXRkLNe5uDLDYQsupd3
PgJRqyGlZk1IsA0BqFuyUsU8WHBYUzTXr60lOtgOLxrVvvLbNp5oJTTsGVCnM+X8zKkEdM/CiZNi
qlomDtzxwgICgsulDBfMcxHCawx19vfoW+ujA9KHeNfIRlDDfv3T2OGBVFTUeHCPOXgFjJN0T1oP
sIOCChaRh0v+UMOY4v7i+0aonNUZu2C+mNR5j227rE2N9wKcydXWZ0QoKGnspEY5/3pns+eKTabQ
uec57d5scDDg77IK8VZolhMdN/Y9wKI3cV4Nhm7DODEWGSEC5wwXd/YsNuV/k6Y1u1HROy3WRoDk
7tOKkWAnpskJZKyJsvAu0uGvZsoCRqMQOPyNcszTWd3GWV0YI9gzH2W1mzI6suL+mfmyLzrWiOJt
rr57dvezXiXwiH6P4u+yZ7NYnyxtAZGvz2qIMGh9pS/ghn5xNqrNrp4lWiOCWcYQJ+efRlvW2phS
WdXnQavltPdpCrpemOZgGkndia5wQJE3iAZ601YBpDqlgjntb4kqgmm4usutp3RvoIm7VXgQStwo
qtf1+ZdTC1RlEC8jqNVcNcw+HIRe6rsjk9OCZT3D69CowSceYFSo3Q7BSVf37V0B7YrbTs7DsXbz
7qn8AtyY7rylcvBgAiEFlphBKFV42nX+c0tENnV8/9wLoMnQ1yzgIpKRG+RQoQ117ynb9RfWCyIF
hkwbp9ykIj5cEvF3s+vHb4m2Jn4ws27ejlEppiaVOpycWodHqfAd3EYZtr6Rg3z2GP+ZVevWqdy+
ycdW2t4tLd3/WnxANGY7wpXJMW6ki7seDR7kmhP7sfZR/DkvoceTV0gd39Wm/5fkXgCIblUkTWLM
7PPdBIbinskXr5gCbJmd7lEU4ZrLvT/PLMRU5mbt+aLqpIbf6Skq8/nbsqoTTVPnbNuMAqfmL3Hv
s64gL66GY9iUIzy7m8/Z2C3MpA/EyA2sdrh/5HBo+PNz5KhqKezTPfbOv/KUNBeob/Pyh+I3wx2T
xhMcIEStJe6qkKsSPPMh3pVanAlX+TDtPNRhkFqYFDOi5M4M3qrd11AZlTOkBLslnYeWQReHvcnS
klK4gygbQ5ir+U2CEFKndTWyRuJQfF8L0JIJ7VzZlcbJ9JMh4JlqWHZ3afj2jyg9x9HqNpH/9CAF
7oyQHdC5Pdn9FhGJxAg5rSKnwkftyQnV0RCc1MjhH/qusrR7JOHgkl4z0ZrEjNPKSjOXbhJxLHAO
GdI34rzyoKpeUTrujdmbw20iewLMx59gX9Ak63HQoXDeqVeT+o3HpbAc98BJo+tSwS88BaoEb1+M
+XvJbPu4egBO/qUOe65CwStJmxyyn8wCfhKGwhBk/eaZ1+gqKUda4TcShaiLxEDD2J8iUcVWFY1F
7/4LpKYvBsCMCRt3IHH5fNBY57qZzYR0aDqLdwxsq0pYitj0HczR1JhorwJz0P89uvaNCr7f2XMu
fLdNrMLOnE/LoRTx05ThV+m+/bxohMZH6mI3H4tJ54LRhSrixaf14hkM1JJEE7icB28d3lKcx97M
LwE96lSH6cGpRSqXiUV8FFP7BiK0rxIEH5lqJx1UvqaB76yiG92xoCf4A/aDRFrt1/HdRg+blM+6
HAq4q+3J/ZtsaCVfN1es98Nlc9eW6gE/2SaMizBGGdwBKPRCQlgUA8LlY6BELeNX0An9A1Gmhsgw
NJ5ZG0liof9leQl9bphE7J0kqLeWVu5le+EC/7++05YxERlE/q4ndTvNBqGlirk3gBIzdp0fI4xF
HM+W5Zx6vGKFBSKzcEA/JC/BDAXm7ZX8wE35IIQ0nMme4HzlZ5DyH7H/KOcI2DCSHIwAJ0BDHOmB
QVtl3Bo98fnXIPam7hpG+q5hXbkZ3zRVkM8gXRZkaHeBOOdcQwjiCBnXoUO9C/VglaFcLOQWizKB
gBzPYnseOm68m8hh0qSHBdCctBxLAD7g8L8X4xyw9ZCl+r42ZTBPSaJ7cJMyMMTJAF+uzHT81B1g
zNFp6hjwf+vbVWouxmo3Rs/Ml4YAL1GjXakh0EQaY6hbCxWSEoKVGPR1O1K0us2oZEX1bQ6bzryz
mQ3vkVqqxY7Be/N6oFj57N8AxitynoQVCeNG0ETgcYO9Fc+H2FLRnAixL6dxMXE/RRLRBnxclJ8z
OdNqNfHfHmXfXfVW0ys4NT94w995ODF1fR9vNoBT4dzfclkujOTUoL6AA3xvCPEHFk4Esi/A+qN/
GcHBylEY9UA4HQrRjaCFB2siQeDFUdnmYvT08Os2W/6iT7Vp+Z944occ15zKY+DtFOToU4B9XveV
eS76q+R3VR/xYDEwB5UwtuzJW9P5a1sPVRjZofLf0f+vwJepoV97NMjapTcAOp+3gZLjFTKuKOoP
nMBNoW2S8sW4q60UptCxlpj/PSzt1UBdxEHUCQND900iFv8rz91MPlAMvPn2/MfPt7p4W+MTmvzG
ahIs5a88Qi4l8dDMT1ix6wK66oKuUrW8hSAlMWhaH/2BC5h9MSak8r6y7hTsdg1/Bxx6Y2Pqfqjf
va4xGyb99VOkaCar7TbKRGd6FbUPZ3U3csOz5RhWEvGWcSX7rB7HiCai0LzUKrecFERqiKe3QM8g
LiBbWxXB9AovfBw9EkJIWP0lruWfx6JfGXMPfd8gZle6AJQrpLBPjKnT/ofj8rkYbYcvvKOfxrpl
W9dozPgMaMYm6HeudZNW9/wFQNN5ZetRNDO3j3pZsA7v6tYgaajUZ7+gPWvNedV7XIDaise6Jhym
6Oa1aTTvVeB8FUu5VZBLN4PK4Gi00lqEyaQ6ROzRwph/BagLGxPlIDeD24d5KdqgwWdZjAkUSdat
kCR64dAymVVddda0EcD83U8yVJqovBbB7kmYuv8rgN8tvtDTdh2jRCCdLcTRCzt0S12+M3rnLBdF
y6/wVT/erfmdeirXhmi4oquvrZbnpivZ7cqfVWYOOXF7VN8H4XAss3KfP0FYqUaEvisBtr3EeunN
Ej/yBCI4CU+gPWKLSEvm/2D3DgMHDV5jhF+ODJiytrFMnpWcGcuRDE7Yg1oWwy2mrxEWPBGo16Yl
dq88zt21IZ53FEF/3p53GBbN/i/+tquMQ3qrzV5GubehQqgqmP2i3xw6hqEJ/Qbw+9pm7kDEfOk4
N/J+JpAAfM075sDC8KqaiwR8A8/CHxfnmfVCqGM4XwSlsyi0Fwj92uVdLXMZNazFarhr2yOwMxKS
nH3TgJjnzv5SoDmpSt6p+bC3wp6nJ3end/6ZR/Um0dgyPSilpoptOuAx3fG8of3ejfiGzAintlsK
YuqwKsnVYY+sewL+oARcLk1kH1eJFhergYksou2rBkAY02q2+ex6Kebwj0QjL+LQg5K16Buv5Ami
LqIoj5e4j/v2jMFNMdr2kI5HD6a08NjaN1z5gZsUXgbOOkMgZvmF4j4W9DgAsYjSniCR6VVESDOp
I9poadfys0scPXQ0GqFF1Q0Z0nt+4l3d/SOrk3j/o5YH6Mmr12X9vdR7gSKBLcaMOucZDtPqRp8K
KU1lZFWMXK54LNLqsIum+AnmJ0g7XNT6qggluiua4MmD58XDMujQHzPAeW0Kf389M34lFmpAS36x
6Jh40FTrI5BehP57LeOSSTqHLqiKFBwL4latk1GbAV/YQex/xGUayqqzhN5/IMZoG/wSSeQK2eGv
hl32A3DojxMLuf/ru1JPyAPr++k0QYc16YOjreTrbQjQXOSNFdxWBId51MVG8QKVmznWpYA8ieK0
ian1cKR1lRGFpz0kjxnPFzJXckI2CPBfds5D2K/rykPchQ7+cwuMrqIP5gAB/DPIBh1Mn2PglVZs
hKeBUo5aKdn6wN8kgialStP1DN+smonh/oW4HqrdmqSZFc1kyREuteZcxeYB48MOxHLfKnmv1Z/O
jdKCqIqvxvXtih7ms3rKOc2KpRNf3hAZcBT2wZ1zhCe1gpQVfaz9OYxp06TgR0c3FxZJ0WjwNtjD
rsPkMi4IjcJlt228x6ybm5YC4HETUGxpjVsBfbpb1QSyoSkvz303r2PPKnnmvFVi2h2q/6nVTEIC
tUpv8G+Xd41NxuW2VCV6DIqZZVj2cjvtZKCxAbq2ZkzbJJO4gCGzpVuTd9l6qBaeCmZA648T+EB0
KHEE3qFIqCsms6XCh9+izUj3XBijImFq2fpCufB95f+Va+Ljr+h+kD7iSCPEPnFL5uMXac3ra1rj
/3HPbYJRch+xfke79v0wpaS5ysJRlr/sXZKJexNplMMC7Y0eCnE3Xg9pzs4GAVX2zxq3u16qUDlI
FEt0jOmuH2XUCLXx0x8pzuefeWcb85tOMRT0u9B7G5MiDMWxWsL9OCVaZW9eert04L2G9beMYZ/9
igLYgdBEqNEalheLw9WgCvFh0VxAvr9/sU876VJEa0ZomQXslg/zuzNH3+bt1pqLRvY2TpxOR87s
+bnGzGH1s/zQ+OkgdfV9lRmQLwM3jPoiYCScjZuR+aOawlK1p2IVIjDvXSGNLZ+nyLEWb6dJ9ibO
xorXeVevwgdWWeTwSIBoGel/++R2WlISlBmVzMOGbKRDlQpuojqdGLIlG+Mw0lQUtwvb/+6htz/V
m2wrmHQyftLxErZuVNf3jym4qdUAGj/g7dMI3xiz4sL5uTjTOHZ9sjDRMk9yIAUVLy7/mbu8bkYB
h0EYbJLdxr0u/QjRBXLUPYO+Dh9MzfqTzEdNyXeVuWfWZvB31HG0xz3k8D6aWFJT2tfRqc1ok3q0
nUgDmqF4Oq3BJ5lyEQotDW5hViTScX1PH9xR2xGD2bCAbNsEiyMT+Sv4G3ah0QU9nn4UulssbyxB
svSRMbBTh6ZJPoHKm4vRgCy7uci+V3MlIxVCzLjjz1Sb84J7qJ4ssVsEbLzwYsPOXCsTLBVGjb9t
1GF4NserKD7/8w+jWTG0+La8yyUFPIgZnjrAAnWHwx1gEPtXEC9T+tsVsCgedNjSkbfs47IstliR
S4T4OsBxK8MiL6PlmSZHB7jJwnwmYXRU598j6ABiLhd2aTxFEFSL6OtJGfgyzFLf93PT/zvm8XEA
4guj8a+Sfsbjs39CTeH8rOslwydYjP5HkxTGyLP2UgVsyFiQpnPSYqSQG3tKwrwiu6W5V2sTaXo/
xZ76WuGkxUNtctZFL5LowW+40re4sNUM4kY3TkA2oz3FV3SQO2nXzUQeAIPnOoLJoagkhpu0Fo+9
5L0bIOxOWxNTPMfYoUEkyWWZDeSwe2HUgoYMNf7LMCb9+FRHNlH1VEMYDeVgW8Ouj+1IAGei93tK
Fxtjh1h7nC43ARX85u+6UkZnwaJw25thmyD/gyT9XEAFZbs3tNpU69ICkpCL/N1fMmSeiLYzZm+T
6522O3HO/5QGkh5ORcUGc5h2OcdbhAaYzYx9aFLQNx2IqqWarwGb/LJQobD++2HQzv1NMLAhf5uJ
X31P6PA2gMJ/a0R1GpJdrovWfNQus7QDqMzskSa0Zo1u4XH4LpHroBfdXcw0lxKNZ4z7rEIPTM4C
UoA/bR5b17hUETd/MzHx9pWsDQLH/y7f68nhTUAwYjboGhBeS800w0PgVjFDOwDk4De46xnDdGyc
/2n8+NfTROE+fLSBdlYTvNEuHtZ+U1ghb27DtXQbBCQ6Z+IJ86wibz2PJWcZiM8pOv2BMBMZIbJ8
Yy/UJRNms12IsPFACR3ZaxdTu+t+I7aXptHqPF8wFxYFwO7iM/QKVyHYzlS8QFVnlQcIFzY9jmCu
QYraypGewBNgLZk7IYPchtvLTghLCUW4+uD5wQmCozKg+Pi84aN4d6Ljxw5zOuggZN0RBS0knkBE
amcX9DWByIUADukUNtH9z/UCMZplHNJjtApWrOuAb/EjgKVMLiAdsqlHjYREcsSj9Ouglk182FY6
oVEN9fuuc7NhTK6XeH0F3DPTPDsOVOSFOjrgYaSNoC/ANwSVqKo5AUvjjuUCWHXNjC7i1kmjxLRH
803H7ONfwPHDGAP03PM49o+wi2GVKKynodk2rZPhwhXuRHXHISJPwbdQVwKY4rXD90lTUmYPBau3
XGTVSFVEQDj4kb0WiCK3Odo0zGI1IrDpOdaRbg4awDfl/nDjQqhNqVUJZSAcMjhyWpFoeM1k709a
jwJnLdikkHRxiwoOvSsbqEY8NaAw2XVCvPfRDy/DFo56LL7Jx0d7+P59DSt8y5FWMXndeAR2o6EL
sw235iQa4dYXS3ZPWnrT9UlipDfOSLvWsqgetM5SVITCF4qYt0aVIJ4xkyVE/bcxgiMd8Jzsc0fZ
qiyPeP5OOx/au/f+hu1MYUjSbZq36xNQihCCVZ7YdQg5qVEM5RuVd2xpynT8CMm6P10DKuB8hY9u
lxXOIjuzpAZzsfhRdEjA/f35nhV676Hq7QQB+Jh9BXpi7BAydHGND1uWvciTud5bLIxgMRTAq2+6
F9sUUnyTh9qP6lLLL/mHVRw0tfuDVrsYoyLk3z/BVkDk12igFtrJHXYw1AHksz+w22Dc+gyfXFwm
D8bE1EejtIMFkCCKCRmN2hqv1HCmqpfhmOl0mop9t3mSW4q7jWZS+RwJlMzqUZGHb4FqQp7/4K7L
1K6AL+YqqFQ8nrQYiHcDXuH0lIMdBk0WaPObNNvHni9Xyz3k5w72l41CneuXarO5O1ZJsuxUwzdW
gqzDb/amSs+VFEyYsafkrWmbV4UUGwzt28fsfZFXTe0c07EeUCnkmkrtFDl1aVgtow4PHKRYCRyv
DXqMypmPP3yDCkuPtf9ewVl4h6shEa9ahKOCnt3cc0F4KyrlS1cPpWVXhI9i48mMhFFXumnw8PSd
ssPGGpROZKybctdfIQ7hVis8QIwA7VE1S8iGqi0awnRk2YQmI2tsS8YsTO4y2nxvwOROIOfHvyXv
NV8c3uDsXXslT1WzPMpYXvlJGW3Gs+bonjEK28xSjsD+0ENUlrHa3Rig0IDnWEZMMO6Ic/W38SF4
fGL+ApVoybS2CdVM3mi4wzFIAIA3pKBk30BiHQtfgmNGREnJziw1/qWeOzZGeQtbKgZhS4AbOFBB
UEaBu5PtdWUG86YoIf7l58/FXp0B3Y1Hkl5ovd1saxxEac84ELwF4manrMwfKyeSi+RLbb7kHjpV
aAFE5Kq98bB5VVp2Iwq0nh5vzaYgcC0LsLYnT4UUXKB852cNBZ/C5sEQUMJl/X/FCvwWphB6Ezy/
9G5Q6l5px9q65QNvLoZSeNcdhoyU8t5mKXipRtKJaLdd2cq3B1O3igzE/Z9cDDcJHPUo2XBVELEx
E28LLVlG3nLPmIBGjKM9XKzHRWbBASdhb8AhLD1BoR66waZ7nDDhgutbK23dLnSqtYRcC6KwziIQ
J9CLCAShTEdZJIW+PtEW0KBkb3yyBxz2wI/Gvru4jRqbAhUVsWrGLVwqcJuSKdGn1c1lNI2EFcEE
N9C41EePGZ/BwQALv4ZoYJo9+TDwxZiuzWmKuFEyzcXmqYist3iCUic6lfNg3aEZOLePO1MD6XJF
+gpaU87Ulg5fWv0W3/TD++HqdtVQOLU1QVXGxuCpRtSx7gYp+aoUgIj6h8qLbJJV07KUVU3Tjd4I
GMbRB2Zjg+oqRYuZrX1mrG/TqVsneS8WsLCMUxfQA7C6jekgeDdEJ+FzQk+jrW6kZREFAvvAfzzs
x+I763oh1Z/zC/rgEFGkxAilXKB6jFccmftHIPMTYHC/IBWizp031OLfkchjupSPmo/b57IVv7/0
L5cWppbHGCRfO+Kdikl5riXt+6j/naHx1KuQcop2vV3TSg2iwQcomtZwv9cb/FOIAItDjE84y01f
2ZMzuD9Mm4P/0fVwom2RYctKH8HyaecpH2gSGFGav2YlCOfDbL0KGlBPCi0hWtgLXpCRq/KoCYOR
EBJ2JKfxtBuclvojfhJjnQKwqw3gynoMzDDWywXRzD6SwTyXuXfMli9l6QaCiX5CsL/f41YkDgm1
Omk9N7t2BCm8Byp0cQs461f8O4Y7PONcMdCv68hwAiZcs3iN+CPAOyTvKfyJbt2FJ5JrkDuYMyc3
ZVT+0+x6ptBxOVWQ7cqaK+g2vArGO69szTfkfRHQhTyuoQbj8rwH7z9rL/HNRie1xhOLUAgT8DgR
ST/zQtgTuH73fgCTP7J1M5IgVjzxbqxVoW+DcM8HmHi/48zComOmzikNCWCPAD8V71fo6XakWAU7
RBG5Oq/j58iCvxVVSqkYSkQDEWWBJrXdBtD60wK200jYychgX9zlqKIyABqoAwwSpYopboRZUqfs
0P3sL6akLNK9gXc0wjDz9HUSocYIjc/QGQlgMMoGKsBRX3d5QO+Qg1hqC+xuLpanoUczkNhXJi2W
zT/4Yb0M/NetXI03PYJFsQ3zlrlNeBdf7ZmFr8kcjdhFzm2b2Rdo+irZRNzPEG8JZnK1vBLPFiE5
pavj2lCC9vI8ddrxuzVT7KjsLkoVEzggBHd5fcGFUxJb3wCuRvmN2smtP1xwCMumsT4cYsroRJgw
9sRIBSZ8Pxf7gjF/Bduue+Ost4P2doRTAH1w7tb4RLUncs70HjFJjsRVHtYzQtL5nszhsWBqF/h2
PkueZgcleLWUJdf6EP5rOOrJdEO6WdOg7SlOZPX0nFmZKCDJJiHckNdykJDL3VJKAtY/X5SIJuRc
Xoie/foWfS9g2InVfai/eeyZt7FRtk1jnU6D/PceqQDzdhptsoGC7loteCekjpFURJVwy5/dVY/n
Cw7ohNO9/dc5pDij0D8mtyMV/zmfGV7ytascCEBxYR4ImWvvUn28comXRxtHdoXlYAhKtA6CgGfA
0HhBYJoMIXpm5XKSUV+rHKsGf8UXHgr9xKtvuuHcyOgFGDK/EhxNmoPaJQzjfcgWdPWxzv+rASdc
ESSa055/iiCorJNUWFUWOUIBD9l/bZHGWbpZHOornq0hZYZSCmM7hInhB2ljZ0QGECOtGiM5Xi7a
bPW3UslslXgJsHYVHbdicvayJUSxwiyC73ai3jH3Nf4a3mmDP7Gl6svlv/OrVCzrAueAR2xfF82i
kBJWtS62oi2YGcCzN8bizNicbsOD8rwtKa5/1Bkjlie3HdH0iaXFMxIC1zPFYlccicY2/xUECBE9
8FqcCFOJpoTtoBElVlk9a+VqRlGFRFo/BxfuCjqquOJievS9FWKefGixO9VYxRFCjRP1C3Mzn6Hr
/x0t3tELOmwS7CmvCE2OEPY61TWQUfef77RxJ2uKaOebOZ9Q82k+sYx3qL2j9z6RJrFk/6FNvFKN
sFFiKeUhqTz3yh/LP8GPFDALCOMt9JbNpzDLcJlGB12CzNzXnUoY3ug6TUfyJ1VbShW2xsEy1osD
3fuX7noO+Zhxo03Q+9y4sxBLfqMyc6RQmZiO/hf9ACT9FrfIBC8li3kYBzqjmSnhTCX/lNLAdUhX
vGivqmQS+DfTe0CaVXl9eE7CxHMHpxlxWBf8MTewjhTrTdK85AHgi3ssZqHLA/7JWF9GDsPQeWUM
sxE9VWFepI3w5y3HOmAGLCLqbHFcoO9tuCGS/5oYXQEjRQ9or94mAHcDqFm8FSKoxkYj+udPxfGW
lt9HkeRpWKedjbN5ZdI6ufWhUZao8sDxsn8iWa4styaILlopQd6wsFwizT1bplVSnOlNyM3CD89i
o1zA05fiatJet3F3R8vgdk4KLhLLEQ5xYCc8BFQD04VreZk8ETKR/jfeLQMTPLFIQZkA9z1Z9h5y
34NZ3eazslVRM4n7ewNhI9gMdf5ldmjVZDYup1/2qLx5tMZ2ngfUIcQ/S1QrXNtb/YbTfe7Ve7vU
w+xKaW92sStwkq1DrgR0QtfIWKprmr4+9DPSxcQmuEgpqKYWAkAqRFZ7XyJ+/w7TOYGP5/DIPGaV
3D03+3KXR+UapBE3KFImMSaSdQC3TpdrsMDnLRy2Zb9jG84gaXbbUhBVSNJ51JVClwC4tpXVp69L
cmoOxpDI3OHAeu5fDl1//+NHsdUmc7hcCWcO++g459loEriV0tKiUH4Ebymw0CMmiYBCztCPw0tt
xXucJ64qFrWWEzMs+WzkloZT4R4NxZTB/1L+yVtQ+rudtDwquE2E1ZPuwgP9F+vS0040D6qOOrXD
yZbNJ9mluidEvrZH4aKlAiYgYnUU9kj4v5oZupa7BJdYxa4f1GeJAz7+Hvj+d3mSsheMUV2o0Sgn
WRSBvUokWwbMCC9qdt/M8sc6cuQx+LpPDhre2nEgKP66XyqjmNfzJZIdQODQfaqO7japW+HRbZ3t
jM5j72wJ+MHi2hwdNwlRg9gWBr2trBtmikd4q4KGnTLB2trvxl8K5zTuHXcLZ7dVAxg8GJrt4NQB
rmiQFcqnvRK5hM/LPzGk0hKrNFHziRITf37mRWphMQ4tN4Pte4WnSHNd0NE7Ued/IOGDBp67Mrq0
6duuQ6iMX8rAVo1qrdZGqaAWIiwKOFx6rTmgHNNhccI4SXu39a1hKvMkbWmrOekx8Jw/pao2R5L5
01EcGY0FGJpsEfNzbg3xf5kt72JiQ0gWvJJpHgWlOKympyodfW7l4iLmA8U+mvInjq0xowDv6A2w
FHEOSIZOf101hWT5cF0zh1XrpvXLAMHCwpCaqO5wROgMjAFsraJwfht3L01xnDpPltiHIdCgGLBA
aqrHBeEoMoG1xdnrRmxzXHHZ6tq21vv0Suoxmbqkpqb02vVuAOwKm4Ek23u/TIIOVdfAKZaEZlLp
sLxcnNbXdqvnUwaTGY509NwZXDXAmlQluTYRvirHFh0fBM353zNNVIclXgg/ZZvPJael3KHAESZG
CbhDNwwJ3GBK4kvlelEJhkT8fLN+mby3d48cBcaoHS4Tsa7BiLZgr7gYT0zkaJT35osGqNo3+1EE
fw2NCId0EtyP5OEZToHuF4+DX24jP1gSrjwRvYPc2S2H3sTh09U6bb2sySeKzII+1H+f1+jIpqz6
NSZGPUZks4THXuzWkheSNN7Wei+uxomAlp36fiZa61odCcLLMR2i6elxU8JoT2lDHcaDx5qwUDD3
u6Q55UcszRCv7H02xodHQHTvTMB5P0nroT2xv7kyunrDjfblw9V2Hs33vXy/kb6SoSped2MKEx36
KMfbA9aohZ4gRyb86+x06SwRzwk0lhZGezXEs4DgbOAjR1U5l9oMrM5ei+aoc1S0w9jrXYTqItke
zMnam9q6kDn3Q3RgDUJP1gT7Q5Zn5G35jb3Q47+Yqz1x6GKJDHSIpmwzDcoEg7nIxh27bemGpKFF
eDhM46+j8mEjcznvLwQnvbroTpoHpsC7RmT1o5u5Tx98Ugv0/oZve0aza5UPNDNW0gNnF9ZKqSBU
n0f4QyBgbwzVusM/7HKINGwoF9qhi7CFNTtu+Jg54eP2xpSTDkIH6zQMs+Jull5FlaKTBpzjCpAe
1HZCZC5VnE8blrhZSxIzl3Nio0UthEyo34pTBWD3qGhTeK5olppUZJ1+3hhnMs90WpAJmalYrtY2
1Gyhfala/XpUEvHWEC5JnCAwIK6o77Mmrue9+yf2oEA+zGUyNQ2kDKgYYDEBfLBcHjGWR7UnEOuE
k1yRCYhuZYy+EJ92wcA/jkRERjTjGTGkxdhddGltnhQ2/x8b0zEWohO3LwZ1hRTnVBeZraLMsLDs
rGbFRQmYpegpuST+6di5cCmDMmr2QjMX3guPH+8t5w3LyXkg/TgeHwMVVA/noReKWa/gXwOYVaDG
wZoT4iy+jD7FdWVLhxfLpQuRzSkG3dncySXUYrinjv8KAe/UcJ5mq1jymnqkgNfhjG4bxs7byynS
zZc18xb7EdGPNCnhOWYDW/K5rInldzAqhp2DHkxBJpcVKPAz+LTx8VkrDSjtsC96UFrcKCqL1M68
GHnUnQOCJf0n2eIawSlWePhg+g8fphCTF2hFkmclwCEAL55OqX3XagWpKVhspj8+VuRwPnTqMIH/
aGeyfIVlatMd07u3ojiYePPu65x9dCJRubAFgFmgRymHPYXPGOYjGNJJUc11uZEybcN968c/opLc
xZH+8m3IXukcg4YvK4nx4Pbaa9MXLBOw01ZJxBLtpXWv0WJLglU2e7bunRzNqxE272AG+5oO6hX3
qmHrDtAuXuSsMTyon9HhoN/bFNHYzFOTeuTZ7Bf5rBpmRct8w4ePqR9zeXYGHBlIRFkDoDCHpWkg
kW1PzQSU71LUrV+R6bFo/uKieHdDlwXK6OdbhyBEtj5PUpVbU5XJgeaKeOl15U5fo7bUPDCx0jOC
05rdpyBhgfW7wgxZJgqfy9fN08//FG4yZJbN5XFikY3nxmd60h64SLToFiTXCXGjJKIGNVXSigFf
guii+M/hIw7wxo/a25zR/Ch/pEViJySi8ZLnCd2QbWSk577V9RcnHllkT+c6AzPwrGb6VDYYc6Io
QkKpQHJ2ApLxdk5yQ5KCI6Cs3ZixGhQQpC2xjPYtARz4rDiHLvuOv/0wFHghkrYeSwkQtLb8n4Al
V+IRSWi8vkkL21zkCF394yBa1hmcl5X0MZJYpsmHQSvFpFy8N1hQXISp7/jDF1crY9+xH25hEG0M
Oz/kJ25V89d8fRxAxEtW3Stx/F5WS2jP9udPDNQWKJ8zR6FCuIra8mhgVodiMgab9VDaItxaw6cP
a3ahmKkcDKVrGz7j63aOLkY4rF24isMD/eeubH5QQovbkX8yYYAmILDPmMhDh/Qd2+pdWBKd379R
7IvwSWj6//uKgNlDN72jF2foOvFikADKicexomw75ZIztVy36ofzv9La4LEeRhP0faEVTqSQc+tU
MD1ijEePkACqhTBCnRQISEfmc5A+9M4+UJdWU1mXbT3C7xURYRbHcJRAw9hWvOneuPCWxJBpMfbK
efH/01WtuOF4ZrcykuEW8hWeD15jQcGtc7kOCi5T1zQzvRYVRzRzr9hwycyn5SUs9ZJzQv8au7Yn
ms6Ij2mgjNIHGqvJTPclrztim/BADrmiA0T6hEMA1K0bX3eAxNqDKw78pWCmgcsTnA5xPa0IudZ/
TWTVU5NpJFk0VYVUD/ToPgr+17lj3Gb7g59GHuKJsex7UQXvzRO070OeVD/zoIWkbWkG3xm1HK6N
x95+DiMmZ7PplafkKREpjHxur1a46N6GP4l8WEyy1Hz5pSAfkcOjPt8gdcvCkGNQAWKfZmJSGIdZ
szbSngyx+NPNmsvoFk0CJov/iqnb3024O7znKvzLvf+LCILo+sTQFwP8YJ8XbqL5XbR73X4dfl3h
PofGQ0bQpgf7tHb3alp1IEuj5CCTQ1AyPzG4qxxkThaVpwxh9TewQEk+uSd1tdru829RCB1+DMFp
mpfDk9pCLf1FzR30tC6x4NG3ADVsQLQrQdsvHE4wuKZfO+SQGck002vsadRrckXnT6ZcgzJYIO/d
xqO8ZrhR8hQr9GvipPfTae9WFDxmHkIGyeF4818fyyrElCYq5WvAohB9xYPGtXDRFFyDqn7YHssu
53mok+PMqJyX+7s3hy0Rc2w/h9MxiW21TSbTvbWEZM/PNZjSG9a0RrtG2oxBCPEgr06xd5fxsh0f
KqcsiXK3hdFEeN0z6pkM2XY6Kq6W+yuvyPaIcpwFtHnrg1mxohh5gz3SAFbO+wxTHPQC+Wvq4m2C
ZRj/QOa8wmSZXBM8OMaoWaAKb84zZ8l+Yy/y9gF+VEEfzoJpqHlel2K1iJLfnWlFIXubMIvwCJMK
+Vs3Z6xeu0zTa0gpn74j3lcfxFbDh3led5SdQg3XIQm/dRwRLt0XDRkvHhD1fcn9I2olzzAGbfRz
kGiMB52um0EjbS6f4LPqIH7AAFB4w7rOOvJI8Agp+xmt4mnMjuLWQRVO+sx/c5EUILFK7R9p/j66
xvvxrINW2clKLCs74JGIC5bwBTVl78K8IFz3vSvQ8kQg7EFDssxt11tqwtzNnMavNY5PGTUG/ob9
QhJuy6PLwHJVZ0axsPnOm6x5M+3iamv5AYD/WGNsKS+jOW3UpSvpXcF76SUmWzxs08ESCHc2Z65Y
6XBBmFhw3kB7kgwKSF9fcpsopghqTcFpwdy0fiNvUUtVQqF9GyJTSDJyvVYcWKmWQjbnax+Cw6aw
iKFKmZyLdBK7awNgBBvKQgJX/JER9T/GM/M7Quu/nCidfIvncfj24uNcWQvgvOyfzDasyxHDcrTI
A7AyXRNpz72+FEup0rr+nB30aDO0MJlgG+gxn8C+bUpEypFxHeBDBBKlCMMAvbSUGqgpgn1U+qmW
zteT2ThTh1UDjDMBJ4QOCrVwfKRxSlvJ08/VGf25Llud/X2dUQyG7lQTUYdreNugoBvKm6rmVK1J
uEzwNrithhcaaHgZoccMek8W5uYxFjmeN3lXcDLD2Y1tCpyjJ6ATdeqtIbVsGD/g1YUyA+tbV35s
lTeISyUzhAYS4cogVI8vbq0Q8qvERmGkNYT+j1O9ZSWggfbEGduCK6CtVM+l7bKZxTDeprWAN8S6
5iH5yIk6DXhqqdFoelJRuPD7E2AHh+EJWMUg+JmVfuHccnEWMujunH5msnRpqfOLS1dYe9t1UMiO
FDaghvZFdc9Ei+QEv4CyL24q0r/9Kza1mAiA+owNwMRpePHEy/9BjT2475ToQ0M8geVtBI0AIUwk
2Fy/AR9ottM0Sm4TbOwsloOXWzqBesuhUaBuAwZZ3ApCP++U3OCTPLeaMEUWSRRwwKfKsrJgBRZr
jR9zEp3FwTaUCC0SEyUyW66s28kft7zugltZ7Tm4VZT7L9Cqlsp7Mm2AQC9UvTvUg/wlSN+R5Di3
QdmEDIH7NDqmGhlOF1kHiGQgxsVH5e0ffBhJGdNk8APD1iDmCFbe1W4gQqgy21sttV/IpZuWtAs2
4H3x3A6a3rMGEuyq22zmXfV7UDz4LnxlV5GUrIDR4qMSdyTCxIk5mUL12P98CwoZZ5qZtbnddbpM
Lp3a5eLbzlyqxdTjzzOEWAs/rpPE4zD/kclzyp2RMG+TafcgA86rRQQxA7ppIuj5ckA/uOHVG9no
bylgo7VIoKaOM3zwHG/f91LZPB6xf3DPMZkRs3mI9jtNSH8YJ3AwZVeYze6mErL5MRFwIluM5Nmj
L47tw6ErlmX6kggIisb0ZNBfZCLNdFcvfkKxcYLElaAuLYjA8kwhbp7uy2kIp1mDfGUkA1iltGcC
W6DMWZ+d4iSRzA8bacBDa9bmSYviuQxHGtBhABpAJ/xULDS3rSJVYTrKhVZ5r+bvEYHgGSDINv2y
sxvU+fp6Nshm6YQO0TvvudEseuAxhvuPtt4jfQJQW2Kdw85IZR5DFpMj6wbGaT0qx/67BNUMUDVw
4QgRc4fzx1yF8zA3N+BuCy40cJQvC1CTg8kIKXfyJbxI2RmK5jew5b+jTwnBDNScc1/5R4deepeM
xhknAxHVbJJIpFPzCIgOiUDkoAxX8FUgyLVb15O3O1x0IdNwJATnskFcytYiX68+z55oxG14ij8x
Xz1J9D0/IIJJHOfl71OnLERVEEIdLlaj4VuS7s2m/Xbq7NfLqTf3XY0nFYl9YFQkWStTT+/fAAsn
5pPqqTo0fjY9XM9ACUWUl55aReqbHnYfT/9OyAM7J0vTwgHJh4RTuA9Nyp13pKOwa429C228Ydm9
+D2IF/Ygd2dqK6rn2o0K3+f+j4cFYIiep1RIH3YBtCfecOKmWvQ5YPK86tvOS9c2HMoopDW9xVqT
g1p0JpXQtd7malTbwJIBm0CH0/r7jmRxv1Mn95XsFKKkKL71npVu03fhwrVnxN6nLQqxKGfFsZiD
n0G8mLZHcd3c+MPsCxO77jqm1i38RrMn/dINlVJlysoKpjc75HukMvoRuG7Q+kxF1ZjIH8xAr6bs
7jn2DH5g22QWehugFe38oxizX060RW0isqSAFJhUJF6GnADX2O2Yak6yVDTM+IfABT5dUfBQAyEh
5N7irOxyZW5cz7ogP7/iYHGzV6HK3+2F8ZohYXgCGarCc5ABRnR2WE6yVvHJ/qN4P4Z5/OWcUSqH
VTLZnkpFkZEdjL22nx7tGhI5L0RweYGqCtnmNsUFWQUgIuizHfgUK4nM6SHz2IL8g+unuhcHzFB0
YI6MzEoYd8dr4v1JGWgqaYUpQ/hlbH//vznxR6xMIzXNlrxzjV1t+FJ9dcwOdvup3tUvv2PRLjbm
MuWMashUKN+D9zPYaOPgyklYqfoY/0TIf2rsaH2EJ3Ou0/pYtozjGPz3/HS3/lOHzW+1TW48R70v
4UCjFEGnqdk2zjAtu08glvypB/QA3jRvWsPwH5M4QXR7W6t8lTZO6g4AXtiVRtO97R2JlvlJFFml
E346flNCw9nTkhhi/vQI+DKrqAE9247Jk4tjziix+PU8AiyGdUFza/xMXV/OEoXpOpf99QipEA9s
SOI/rXwTveD15pJEqt6PexWP1lACWR1fS/x1Tf5fN+ZLBMkiNovpTSqEoV9Dsm63uPR0z4QBXjVQ
nY28S1Wz3BmJ6Oux5JBSG+APOeQRJHdVRZJVXf9GWSWIDeCaJkD43u5Gal8iObjBVMTTlL8cCpqI
/wljOSt3c0HqDnGCrbsgpyFSzcDJ3s6jpjrItDv9qWUf3IOfxEkz27lGxO2PFU3RYAlRI8XnwHDH
YkoJMfGsOxN2lo4HAcpVUPqkAm7jRsN7iCY1/5fgJwrebNh6UUFbQL+YcAJZ3aRpRxwMIn0jiZvb
3zlN8/VUSjwZCmhaeqXQ9TZp4MW9sIfGDfMoIUz2Q/UdJlW8hEJfMRtgDzqyMmPFZy4CUmA5kIvL
MKIhEKWp07GAmcq6Nvrz34Xy2vHeq/Aai2z+qbUWHgfFyYaz8CEUmD8ak0xSPDIKikaDJ0S6Pem4
Cf8tc+muDKm27+2KwSvdV+ajx3T9fi6i3pNuVQxa9T/wAyfzMro+bhI/XMcrLa+EafCTRWy39cZK
XvofKnJus3i7+SjtOLFt2M14WiMuVSufdtfaguuuAsP8C4ulKaiJIwuWFx7nE17wge045nWCGT83
Uz7q3dT9qLwbXakCzfn+jB8Dj+6/7X+DZA7oUyBy0ZlCvoqUaKVToHKQNd7Q3u+Lg7uTpO8BzWN/
o63/sweW8+2GFh7sZIddd0k2hYN2gOuZZEnVh/k1RX2Puv6xHCPK9MRrapFiujV41BfiAmMWjRSD
YKk7FXZumN4M4u1G2gL2RO/EaMvrVLVW+8KLGtvMlqCgUMPX2ewcagxY+CAX8Ok8BFxD7YLLT1x6
SipmPN6QDy6i0K3gLzuEyTzx36sDxuBLh40GxVrjIcgF7i5it1BI7jMcfZ3+aBt8+8PqOhGncKZ3
Qr4FQr6CfYm7ZgFnbyyukGOcN+dyJqcg9G+LzNMRphrx7bIQkjFnbMwTaNVQrErgvm8JUQmnKauh
jTsK8sT0Z1C6YijGR+Rpzdk93Mg5T03ws40tYGIgQvdF41S537FZZWhN0YvPdlVGqBFW7Lh14Mdf
WCsS3mSIlEbbSuv+gN4OO1xdweWIVz67qaSigE1D2l7EP2h6nzRtgbhe7Qvs6R57u1w6CO0+KI3k
ruZP5VJFno3fqqy3E4Aai+f+dxffl4OuD7jaZXDSD584hu9gf8e7HUnn4YJJIrTjw4B/tD4aWgGi
gOVOPasTl8y6wuNJ8v+ixjtrUTMT0Bvn+FvwejJnOHxc+NJ3ban6q2CVTqZNIEpyexuN0zvg7fCk
mVplWKSLTvpiIE0nkz0OJBY8H59JUaAyqyEikbpP5bVFRkhOVnFaYjVtP9BJSQYNiPpdI10LMT6S
qf6N35v09AKoUqHOCklfxPQ2LwIYx+dkkVGV2J6xlUVq7jGXYuIhK0NTKQfFAQ4so0xkSTLolRyX
+3Qjq3l9fn/pXxuRpV1BzOVDGHGberEHkp8RXJH4s2FjKDSQgYJ8JVGrNbpkwqGLelck0qGOryg1
EYnf2A29+GKpbiizOjZmnPz7sCK8w5iNSMnoQYAreBNlvFbil40RilP+ae7Ts21fJ+fcqJq84peL
tPJZSVM2MwkbvNNgn5WxwbbvC9YrZ8bjYUj0Pcckcd/nDNapu/HTWq9S+comLsH385BP57avWgOQ
kh4SM8XJJHjg6lqNxJ2ZoDEfPQyUaO7u2TbMU+xjBD94bCIqmKqq+YuEyY85Sw2rFir1BQWZ/bac
MpR0M2AUHLyswearEwNMCWzB0KLiXBUGdhWUMqOfnoYbeESSNf1lfJWSu1CexY6R/aBYVByayCvD
E0sioAfT7ZXXWVY7508VwAJSGWa6qXNUgIyknOXm2RjvwuFifHPlb2/K+WHUl3+lNw0Ii06RZNbi
y85l5PGkzpxaaeJcERIXW1jqAD0Uzh0TyFvS1B4IHtBterynRaGqJiMYaIaEvM+kcOWOGC657G12
sVhZiBXoKp2NT5HtD2wakHfM1k7++LDq/BGXmuXSySt9FxsjKVhJSZtCQVXVt4DD5YRgx82bRfrf
1M9uwiace+FDOjpTj4EqfvmQoxhyLF/7KqgwSfHb5591MudS06a44Ns0OW2kBLyQWcqHEV4dMUPG
KqzxBJYKURy8r/c7DO8cBpGkQI5ZKQNxKJvZBKD+eUDU1XlKpnyjJBgfN9d2PYToqunSFVPFbx6M
jc0yowKPTgsUM4/M3QwVN61I3JZyADxttO4TqUq0gREzDX7nNEwEDJD6O96wrwV5CjeWsG925bCl
UKjxz4qu7Fu1tGoYpk6WSv0F+VTm+7yBX+/NHsJwSzB146kuVet82oDHaO6LO6dc03eSAQD7VTby
W9df7rCGJX5cZ3aOuY+TibgPGoGlFuvoCNSKJVqSz5kF1r1vy2MtyBFo0u4Jgq1VVyPzZwD4d7K0
wWzl4lU/J31ZiAJ9VCmJfvCwJRqEZwrIE6lsqWHNayx6jHEMLBS9k/fxsbSHotx6KxXLn30cw2ga
C5Euh0m1ME5T69J0NmQYqWd0g0EJbaboyh9hEfZR4CLCxkb8HNC8x0l9dimBj8XRsJFVNSnM3L4t
yyumwdLGXFO8wtvzE13U7psz38Jh6FL/6A+fJzTEWrXvlW/Lt/586BtXteTlIZPUa5GZuajnIRXB
BmiWp6SSMEq05+HyhOOoV0vloh+nd5fKrISJ5V51K379eOjpZQK4fpv+CoLdI3UOeqPH0fQJQWtJ
GvhqM6EVYqf7SfE9haX9oemQ1aUtGSx/IcRO6MSbM8md1lKg8ldtLxcSkOo/iE0kMdhCvB3hAGrb
mJx1o34jXCEvFBFtR/cKxA0xXhnDU+HE7PM8WmbS6jTvIFXuoiC7i7ZFcspntx06rzitoFPs7TcN
IKHxNHs3kQhO5+51f58BF7/EWlj6Ct2JjPpN42p5YUtWtYm9iyhO+gwkwqXP4+EhTXHNwgmgROoD
cthCAGlCS4jLJz21hwht0eNLKUGKdXmHZdzFMIzdTUKD5vdNZ/GJ38i97Oz90fUyfxR8ZN+i6bDs
mzkkn5cCVz6LqCeaVOVKXJJkdEDgnSxtsvDHzi3eVbU2Y7HMvD2mHZZ3gP4PVOp+KoHVKjJ58WE8
jwaxbsiL4w7+pgPBcb4XZ2ChEde8rSl9fWj+0PIIsTaIzoJLEhCGaO5NqUL6Zvtz/QpMyC5yDLBs
dZoBYV+NZZe3PcXTQKtDAuZsRNo/LFzoAKKkNquqUgDV53PPMgEqubj+ZiYv+0MvwLNxdS/bXoIe
PhzbyCW7f6kvBVG4D9u6BVn+AZkBWMbvVOjIx5fZMx9uhUzUQPEU9ihAFlFBCE7EtWwH8bwHFu7p
pSVbPCJQGEmGR+/AL3C1vYLufXufEZe45+q7yXkHSxM7PjeM9AUiDlX+PZCECyIbaHSsK3DZwOhi
vIc3JWV0k8wfGrwHfuVpBqy2oL9XAcPZJ3ILBC/GqTz8sxhHiABUw4WJTRtsTBylvMU6jtZrGiDe
+RTWFTHOfJ60DaHFzc73nIqnN/pTJR0SPSTSq4zg7/IvYPVzmd8Oi0mibiXhG/KMfRhjEZDjVjRD
x6OK+FR5o8E1A1/mEBZxhSkPBFleIFp46ifqdta4qFcTBqWDNxLLHfbz3ZiqiVudLNZ2U4jb0+ic
SIFcDdHMRApEBytNErQbB54aTMUsPev8BZcgZ9zjOEKxJwd56Xg0eFLzJNDUs+acLpv/jISo5tvs
BX4aD4oodK84eYfwUJ4edDzxaQpqKur9AHl6zwYmjt0VzpVkkQR1pI4MF5W5aXfYpnxpzEHLKKkD
jGhEnxCSu7eW9nZJlgPGst2gsBiuUn8FfL4QLFvWGN40qScWiupE1sj/0POGhzHAonEQ38yVozmy
Jb6J6eHxF6m3Whc6shoz8DydEgndFJHW2/Xitk7wsnRulK+ZLz/FDzCw62850M+n50oRW3TuiCQH
usCqn7w8KPdfOze17HEaUikoEaGblz69XMY75jI0G0ea2nTxNx7p9v1VQqUATGnXkjKo3AqrB2At
fmAI+7hAZuNPv5o+7xutzsbt+aaYBeqEKLt7Wo/ChNrdkRPgAOsxyxCdnXm5GNHJYyam7mFrkykN
GhpvkTcVDsUAteS2+XBcVZ40WnvPFGuW/h5jB3fjdl07ZShZBhNrpV1wWeozn+nO2tsk74Q5MFpF
ZR/2uTs/GYrTt5aGpVCdQDdKwfRB0VvBKmZF1uPmWYiIxdjUUBdWep0W8KH1M7/mH89+7qx+KmYt
zkeAaMdxb5N0s1j+L3A5tJBp9sNFxt4PMUdQ3khD69KmefrYPbWdzzl4HWSESEmqiPCsg/bfyY78
TYOtGV5x0LPxJrAHQIv0x9QEf39Y+x75dHEHauAIQk8E10FR4OlD9VtO5JW00rs14qez7P1gdleZ
XHfJlOqE5ErlsJ1e7DCf8cW+Tu5ouiPc/rEexLVNaU1kMHAUGDQPEiwx6PnJht8kyn4RsVisOMN8
UwGYMoYQfqpcpneCbEfbpO/vDcNBo0qWWBXSQ6xKnTC4D8z7dbhEMBGucb85wtHparBM2BBtuwCq
O8KRg8EMP+HlX1zFMhHowDxGh55HeTBLefA7ItzojMCjhs2ThbdfnGx52/Oulmm+fBjBvluKNnkD
zV9MI6l8rRiTq0TI2/eB8Dj+FGNowvPDdyJYCe4QARChFgJ6T0fwBnKTyJs2TG8302r1Gdn95zjn
D3esi1toGLjoohYbhHW30pNAIV9tQuEVdQ52C0tBWeE8Vf5zbT8VZ3DYn8aqxEQ0b7kF67rVmB4g
PLNkUH9LcJJk2fX88Ro6XGmNd80WRk6eo2h8Y7HbA4hwAcxK8nLrpyNmbC6k8AbDmkafPgr0hQNO
q9PHSZNnRlRtnaf2vvBlSr4PrNuB1Nxpu0zTc8QWTgDXnepuC0tvzoaztsqjUn2MBwmNOuG97N5E
g5bCt1d0f+IFI+Fy8538//rtCD15KWzNmuFzYEDxEpOVw0kjAyWfop/3psafxvZ4h/yWTQb6rjrE
MVkBsGRREjYugzs/yxkTHpkmy75/g/ln2iBRRegnh0fjPdDy4zUbrLIV9RqEr2yArqB2loN0+rHu
0qIgTVTlGuhWQX4UeC/8Q3j10Vq0xHZ4wwfosbBb2v74rEP3atDZmfGpVJF0NSMFqfzX1QTmNgxM
cxYHvPDywiJqAAdy3TqvuHYYvw7m5OURzpA04zGe9yi5KRjHHAfBEVqRqZbtsrMJPWoiaFYXP3WY
uVdZFAyOWd9/6x8YPmrBoPPAT15ZIqMFF3plar/rhufj+EUITmEBIaZvBCj+dR8VilRa7WJsU3jT
nmjw2exB0CjjAhbwHs1DFtTTPUPjGzaBrhoXWZVAeaJEo8b6QimWO6Cof9Z3gE3jvoyHGZX/x31M
eo/YtPltJOf2pxfCxEzMjR8s8zqailcVbvU+UUXwI6g0KPIv2/509krxY1Jdow6GXIl0NR4zUUWE
MED2rcVUBzIhAyeanGs4lUBLntE8P9NcdHRS9Nge8aotkzvZKelfeNDbjqOrK0/Cc83Af5l/i98o
r7ICIxRl6+fxU3C3s6RUq+BLgtF7rDEY+IjiV0LL4p3Y64HorJ1uDYR1VYsBwNF9jWFOo+jQ94VL
rJr/5cYPJWLrvc7sWaLAatCCghjgS3zIRPrqc27uDOJ+TdaKetL2u9kJZ/zWg4Hwr+z4DQPsbj4z
19Lh0423Jwp6ihDbuNXwWCyVq89J7LFbGAngKp7tRJdHpGP/UGCZD2iq17ZC84V7lA6oQs0/Bs0W
UUs0Tg0wli+qZd0Y9oOzq9eN12YttUUnWqfw23NmmGBGxqzPRKTRCbhXmMYfgKK0OaFeR5dBtm1W
qSgqTXIYzSk3l54C9fsCQRVYg3cnLI/8qwJPubrqfKtXxdGByoMxg0szqMN15XHbAyvxh9uIi7Mc
mprpZcLYfh0LYDyo6B2DnilxdxmzKZ/65Sj4WroyOal/L8E3HKldcJeG33erQp4TlRTOj09os5La
VKmtveL3Jlz7dDqt1z4Y2mTpd59rV7BivVUmPRVnTnCQiZoY984cTF/3dmXHm/C254nQAhJyQRzB
f6w15xeXszBlXkGX+X8h3XSrviQwLl3SjSKByPqmmAnOhGm4PhJSQr63IoqywI5iujj6anxE8Fu1
h0snWBXSgXmzsTqJpt66vm4AvCbuaz4u+xLsRupcbSqr7GVuO30IhCmhIewi9vs1GNxWZ/gH6wGP
SRUlsDgI7S7sSBdUcnrGKDC/JNM1YbEcPMAiQsDMLYKCScW+5iGE2HEYRUmrdQWMTExtb3g9tohg
tFbUE1WVPc/F8MvB9hejM6nbIeGPIekTo1RkpOZTPQtoinPSbTAArNLhPoTZUVSp/uBeP8/DKBve
t7crB8v6LjNJwTlM1DIO/JmKlQcdV+V9n3zjQucHUX2otVleeRd8+kVpucCJXECFEKnpDBM/CE7g
M112/Va9j/52Q4ylRe7VqwwLer4ktyl8WYAjS2O+ftGt58t6m0EoyRQN3sRZvLHYzXGacIGcoEIv
e+OAajOjJJUTt7EVm6B7RbOe/OYaNFurpcavOBm0+9cFWMZex2L+TP+3NqkGb3Nnhit4BoGnoghe
OkyUhc2MjZheO8Niv0X4kih3VRqCFkaKgHvkJ7gN2v/dQ8wQOaTEYEwSr9r5qmQ8C2zB/sxb0hV3
PqE8I50bERNCdIkQS2FilymgSdHpv6dNs725QPv0aqCvMal/MlGoemOz5ZnpGk4EbadX8+Am8TSc
ZS1a+kpofp0oWJGchbgEefLX0aWBtOQ/YpZXAauPJOMTYOWgUVZC97Pxz/pkQwKrni9gNlIESN4/
LH0zQy5OmykZGRdJESKbY4ne9iTqrfdmlnsIGhYq4QIAEvDI9h63JaQE54lkm1uDNBPsB5ybMA06
w3egVoL8jaqn8cmAzLBSxigfqF6T/FbGpTDlhNJn5uooxZ9n4ShbrrlWWOfkE8U/non8fKbfBArq
PxYCg8Y4/E1paYXn/cCJAPRY7BCxFmvmTD0WDnzlz+8xkdB/8fUSiiuLVpXfO/slhGv6O0nBjSKh
wJ9oX/l7fsudL7frNeBWdwVcIkHVPeQ/bwmjcctyzUzmQSV0nyhpH2iup+gH5MG3I/xPVq/buTdj
7YeSGj5QVY6N0UnOD6Ls9jw/bZ1DS0gqsiMC095Biy7j8fQkPeZFpyiMNRUhfrLKn8uJZjmR7VFL
GjdN9MA1wi3XVUo9H3QrVRYGLH7++W0B9kNOk4ZxDZsI60levzH62VmaeZUhrx3haubivPFMjpO4
dCZ+MZV5UGzV0NaIv1sTa/y36mr5XJn994DLiU3stFalrljJQJajKM3P6n2+qhDbfloSatBtF6Mu
uwLu0C9LlQk/f6vxTo2kJ20OefiPmlm9V6AwnPzcd8KCEKwoWm1blmPCnc899N6V4O/TcU8Jow4L
+tTsK9bt3XmwrP/ZoSbqHYFqlLyb/yqtznAYXbnyMyhC3jyEUJ0Y1i4czb0xiLVee38z4VCyqLCv
GZjgEcfAqBb743Ro7TY57HcQpCQxitzYpplnktjijnsuoeo4Or4IRMnygqqVFEpmrAFnih80mJQ4
PdkOOYOm5EwB45qDljGxTOBXIjrbsh7salj0d2eVOxE6n7F0VbarT7IU2Hyjkbwe/pPYxEsWwRWR
wYAcdVU6t739bbhBjH/uye/CDeoaEiuDYPDNqwEmYqm4oORFUy6LOeqvOhSNVy2L0kR+8MQQRruV
587ex4GcqME5akDiBJ9c0lRPlMxAD4SIjzwU1sYxS3/uNkZWsJe3OtQJq8E9Bg7v9LflbJBXRYDI
9BYLPrNniCMUP6HNSiLRRdguRpC2nEnQXlpx9FhIkYElnIBq2gftmoqUG3VkWwmBBjAC1RNUWWd+
hbtZX73Flq9mM8jR8Wk+eD+D4aqoMiijI8CrGDww3s3rHyIxsRBiblz1aKVuvkLmWZQHcXp6PC9q
OY5diuToyfBDmmS28scbBWp3x+RhkeokVXtFLI/lOcM7+WY0XfT8oZ9MDF8AVR0kWv1Z95jtKdct
VsAVAZZljMr3BaqnP5CIzrCSyU8ffSXLeEhljm7NKtTGeUcNTnQbW8zl00ZxY4fHKuYD9fy5enR6
5Tb1i2QpMaHl+a8aYk52+PXe7khskdH0wTURwWxNLWNAOlvMAq/lFsXqFmwtmGHdhvpcum2m9ej2
8ggaervqiVLoOU92Ex7E35yvSVPxuAY8934mOEbKA+S+6KZKoVAwhBEKop0ELus+FIXPLYJW62wX
W80gAXj+bf1aApS1rRRqvQ8JWllDHQJYac3veeHdcNU8vzK3LUEyE4z+tDFDInuvtjN3gYgsjhzr
m7gqKzVf0/7B+ut9duHIOJ2GINruKy7J8k3hjmGIWW8DkX9MHwPWBxEhB7lQ1SkJI3ZxSIBDsRPN
nLE0moZw/trXEZKmmCJvVYpinf/mEo8TQAUot0pSLM1Aux6sjvCcK+J2Sde/QPp4Xn2v6Po1Hzsw
YnEzmlawRTc0HltCo47258HCXrCDnyybwlX5Ku97o45gUlyWJ+K+pf266b7dweCHqWQwYvNsOyKc
DyI6eG3EcSWJSH6INOiaP4vZve+zgMwZGtmRGieXrhVO6zg9UBf8W6PBtly4YwZENMG93jltjAO/
073iAzEpxHQx2WNKuHdg/PlKsBi5vN6cQK5SUGdIM30D1Vb75WugVBP6QuLyM5CyIs9iHaN5pXfJ
fPQkp/EKY6WSSrPkwGLN0Vk0ZsNVMAbMHGhOHMniT7VSRDcFbyTe6pRMOqTKVMk3okaALTtwtMSh
+M+irvvobGl+UFB33QtOHlfhqZC69DsYtGNU00V4oe54/LRgoa82+/UtOTVeWTeTPWCga97Wj1ov
wyxx/GIdzL+0WwHMoFciOlmTyYD27fxmZ155l7bz2DMoqTTZDS8zr7ZDvnF6pKimqUhpabgIaCU8
d3ZR1GNKP32OyNWg5x2NcSI6w38PRwfQ6urP4Sd0l4Va5E7TxL7fXhDWWl/wI3SCLPercrP4duPr
IGRyx+lWhqh7bT6egcZFsQoLiy2zuoutFJkXtnfkUjlylCA3itrPf93GOjhc0yY0qZkyaZBRCkAL
p6Fvg4oo02XhaWgKnD2bmb92xc08XaxNl5tbwSpi8halLtEJalyTA+BVTy48cUcu4EaXldpHzNsY
rv06pgEqvq++e+t1Y9q3AbOBuN0qVtcMB2Fgdoe1uuDCJWl4MdaGkzj1z84tOCeCNB4KLYyhV6Rh
DYUh6F2fRugMzMN2YSSSsIipus8aOGjtg1332lFzxxtmuC+iQ1bOr/CDY3rc1anSyNOmt06kUdSF
SfA54Vg9bxkEpQUVZUhmfTObGveoSNJraDVvK5v11BY3n2abGLVFBldUeWFRW09STxm/3snjpkeV
0bSZh1QFDgFmJElto99lCMIeEbh2W0pkx7HG3AL9ISXbGjDfFPRSUo/XokM1d5aeao4S6o8Ts/2r
FGJvx+xTTBy8oYLs/e71+JLQH1op8XljXKuQYa+3fRF6pe7+spAauL+jiqkwZQ01g6K/qE5Czx15
qLggUWcRcMqwU7dliPIZj7hw+oB+KyTwROu3g4u8Igr3G1jhFLSAZFjUZw1oQ6J7Xe+2Db2Owwuh
H73VnY0uHEooVAbtoBNGq1ueVQV24AASYI8VE0bwsVj4tZEXeDuGGjljYXJyQO0PoV1Nl8PEAxH+
HkJHrvGMgW/bTSeI9UTx7brKp/Jr/OsZ8NQAAf2FYrI5lZ38UjOkbnPF+ArHtrjCSv/FOgaDg9HD
BlmXN+sFk0l7cCK6C8xY5lcES8tELODKQzY3ivyuP1aq+UFGjpXDvp+R6AE5KytpHpt56x2mVnPR
GCjbe74yKBD0/h7bQVaagOTEjPDU4xT/eFOzR5kiTCDQH6XrEIsEw8KJxqPtLNSYeSAQcsYCfIw6
Uw+7YQ18sJx7MG8C/GeiYTOcRt3J0gd9o0ij9L59LPGV6apWnnrVvv5SjgdwOdsd5e3StKc/ToiE
DXkfy0PYDgP41xgWnzTZnruMk/iEZzHUKQhK01sCrF136Aj0N1foYIlIewUpF21uYMoaPe96Sa+c
Cypmmxb8GJ4Tb3hbD6H6Txbl7vohNnmqsA+7mIUYyGAYTy2iDBVtWysrn8tIEa0s2SUxBsCRtvdJ
5gzXzCiRINOJnipNBtC60O1aDwG5U8LjcYXTDXnq8DJoe3JYffwvSNrv2Gl85Tu5Q3BBBs6ldMFx
xNyezPZVWEcWaQ/oHhefq9iIeCBgV2q4f/HqffE9c0N6DsGqHMXskkbLaVwGgpVzXcm+PjhjSNg8
7mWYEgrKOcQOK/9nP+ZMLrLiGjwVKTTBqBH+2NCE1u4CasFxFYQleyH9z2iIDrBWBCriVnAke0tM
qA5RUziFwWIlwnqqNqAwGMJ0gKdeBkI8LH2tbljX9xmcMaGWwMpUnwR6k7L58DDL0d46m3PZWnjM
xkkVoss0kwEBgZiOhma3wXbXVl/YgSJhanxZdmPH75oKDvL0CnlxyQbX1cp4IED4srMtzaUgVtPe
iSNWHIzA3w37v5p/tThRSAkUbBIsLzkms2WijHUelp2ik966vi7xd/Ae0p7p7spr/CDTbZuizlEh
Jiv5P0xymrkZp8U80D3EXVnzw4NxKJoQgTjTIHHK7DcRVWg6smieOrKumyoMl8o1dsWdU36eRZMi
lCzfejaUWw8uKI++cgsTtCRldpm9tgTmTL5ZzDZz0tP2j7GmV3bwzecf10t/uLj9Mu1/l6F4ZEsb
x0JDn+V12OlFDh1wqu+WoRxQvih4YVccTe1Y0V8hDxmOEhqF3ESaJncrUI0P68QQeNNuIvIs8SUu
pmL/3arFwI1Byp6g15rL1xDKp+vDqsJymcQqDTzlvtuul1CcD4T+UEwISeYB7DXh9h3ARE1J1Aka
hCVcCpgKi6owO/yo2Ym2ic0co1amCLeB44kax0BWGnFGnBgRErOjSV1swprUSeR1AHWYukLVTtuN
sTFn10PVvuqpur8YDOOsjPtwJr03bKdW9v4haK/ej28HoLQPMcHRXX3D92ZBv3DLdRlJRHDkUX1j
pcr9mYS6HIm3f1tjrBMQeg42X0DtDEF/vhawNp4SNzPa4AQgn6A+kdnZwRzGGn07/2VM6Ke5wEqF
aHYHRCgH+TWp1yGR2ubuUavtjR6CCriPDlpTH72yScOHZkEINiFpzs2Ddh+TcywcO1i6FWAeRYg2
LA0Br/HiehWPe251yW72ZcL2bBDt6Wc1WdMGSe6OmVgcuKsuvVY/yEiTJjQF/YCd9sVos36mpBcv
9weHd7Z8tHPpZggg8uNa/tBpV6wI6uYwzp1OGlDz/HUXc29s5g0HqvX7RA3ycf5iYvjJd/ijnVqy
Xm9yI1UJfeCeTHRxltsY/9eeBaDwogklqpWHXPwRE5+QW96SEDho3OyBXqv3SbLCXAgrnLhp4+bq
2ja0uzZEDKdliC9JzgDQKMCkGmVemj8AMIfkrZn1xpTPERGY15dl4BFOG/A/7YwrJDes/QEyTDcq
ZfvA0qwUbYCWtOtQMGLQ+ZN0WxHzDJw4O24mKCzYmB2U87VQ16IJ42Ys+7T2cKAWCRr2ksfBmqOx
S6Ny4FE2S9q4sbibV3ueEx9ApOl4AKDPPBwlJ/0GobRkRuXrg4PfYhiwtNQ3knG/8cqHg6HU/wqo
0g27QUXgEloMQ6ju5KS8/lR4SzzVcR+cFMlfOLmO0Y+Ik5qG9cZv6RGBYp26mETiyQmM+KFTKRqf
OvtGTzNoso5d/Yn3vpKcLnj6shm72ewLLQ6TFtyj0JX6u6stABr/BUer/FSeQT338e6tfZ48Sr4u
QuHje6xFAd4IIFYaHd3Jt5xoSLsnHYFgfplOtVCj83N97YTtIx2jlNNjJyu4IysDLJSQersNtYTm
VzYwlv36aWl5Jv2YmLYdoAbIUGPlo94l67bBIwvwlYXIo8nDyjx6Fld3TEelNknIjZDeV5kTzpjf
T3KeK1h/Md4olD79I/I0/voXEG338y6IaqF60DYfmys4aG+QNc5jlPg4nAok94f1JlvbqONbtiP+
rP1LdMe+ZL2JDVaHIo8LRe2jn8pOI9q+8hqlz/wjwdXSx3meI7bKRTNYUcxmB1mDmwKT+coW5/9Y
naGg86IXZrh2SgjaXTKrqOR3qqNG/N3vnvP9FLJVm0fvk6zxHEYdeKo++cTtJT8ijmhy3ntF9lth
Dc3r/vea0xqHY0TyuVkxJgIkYn0uUshCSf41ghAKxmuxEmwJNupgB2Uoh30tpfDXyx32FGSYoSdx
mhhiRRBwIfv/NJbp3QXIuc1g2h5xRJu6x5rOonHk0rEyI74ee631zLDSKZrztHG4MtdUTA5bxZxo
Fd441fkEpgq1rA5pDi8QT2Vkingh8IgBkGd+mFLv9fHwj/AfWxNxCUHCSvsPBf8tfEbTDw/oq1JW
zpfDGKEDogPv7YONH2ZQOC0XFkr4J/mf3fMyw+5kFhmj+vFBNcLNvK/NBZLRAyDHEXjN7qZ9XmC5
Phz4nhXRwbwPTzXb2tkuCC/CevpU6JfCKS5ooPrjMsvgsQQjEIMA+r9EIPwzoCYnieNut6TDlhpy
Co9UW47tDDSS1rjA+oL3NQkEIeX/gUiXwemK1EDVW38pGUhqtAk/XDI2ivmS/THRi6n5e8HN8bVL
tZinCoA/TtZ60TqyL7dKQJlEXZ7lFO39mn06YDEyF049Jb3T/WBlR7UI8w/HOSysQJAEU18DRYhZ
nWPQ3sxn1UYiyfrr2bO81ggxMP03MAPXAIOcZAZW16pqUKUdFDwENIN0NpNYtaEZhfe/Luwygv0K
iQv2n5jvDpmH4OvsoymAFe6+pDxb6Fhd4E2oqq8pk4lhlYUlj2I/F2SHx4aeYTiaq6yf8e4hr6kJ
JXRTU4o5ImU3eiASmvMuEvB1l1+WofHw4gVZG4XdaJITUWhDJ8Nt+rJST1jExjanq1pATxHrhn11
mGBM2tIliNGoeiK+g6tZ0woa8+hLC8KFYJzJczI49zafx2yXKaATEWlOeQWuF+ynVb0K5H1SHUrQ
Sd+kQSuQIVlL038mjlk1T0+2qi8H/KCRP0U/MPygq5XiAwoXWIw9YQXStlCHbkDai/em1vfp7hA5
LxQ4EGvjYNFIhoCGZVG2xDdzZDhiznASZd+t/OfiBrlAM46Yschq06mzIAZVW1uT7pnS3y3NvFDE
Bz0iP3vNL977kEt+Ud3O0CNdzR+X3GHe6pfeRLfqcJS/xmKEZx/Rvw2t0sI8bYzPLuRZMPYFrNOr
FUM5fspTLcyHBAl5Ky0TgdKiCCNHK5DnyF3qA0m1eeCkCWVb/ZhDAyd6m3WmmKw0lYAHSI81YRai
CwY+b29aYncQYJ7y57BliLZaB+kUkml6SNwZ95N1c9mE/fOgYA8/ufaOnhdCxp/GTufZ7iotZA2I
rzkrLZLi09AL6cHx8vEhK58I6C7vur7lzHF25EQYxfQMje7PTRS+6X9gpyMJU+i6GcsYNErPWtdE
Q13dabSimF905gDu1Xz4hL1QxIfujiipZAu8LC31E0gRd1bEmpmt3yxoF3ggUS+1sgRmg+X7fcfI
nVlQkKmiEgWFilVYUvMd7/Chf+VmmPVmixZgovTEeecaDZojw0593uDNeTJxWBJ+BzpgAE5nebA/
XLpc0xTnfu95Gm20BFvPdK7a9Axj6qv9kP6YTZWgoyY0/z3k7OXDNuj4j5jxvThTz2WSwyrkm/qI
bPE/PAHYlhRHv+ibJum4+/CY/5wSLuyniZctX2phYA03X26OTfQPYkUHt6BQxqG+dRYxFWObBeMW
Dzzl3eopDVVzYKAYAU+o1e+YFI4WpiMU2wN7oeB+0hvXUJvUvU7zHmXW6pWE03kbqK82A+gb5fW8
SIPzlMzu0hkqb+Z8IE0NSRgGsHhoDiVntTe+kEWs7hf4/oyZdZ7aDZ1jaHMCHBJSllcUT+dUU5OV
aWKNwchNAXPK/VsdmtBTfEhboJMduVGsjpmwI4Ad8Rf1OTIjXxlSwwfZS/LeL0icSQVrDx5qCaOD
Dvslhis8Ky5S3LDU5knKKc5V0FfAVQHR1vdr5XBXVYBWna8tg6dccyJa0mn0FfCwQ9ttg2Qg50Zw
yPLsOVJjv8DyEHh0Ds7T9TZ4ZTJrmQIQVB4kq11qr8+9dd1ksObwt7lp7rhA5u2TNqaWgqrtm+po
0qRnyDD8ma0U8RVDV8vO7T0zjiliISGqcrszktioUNRDLUwgk4cajyfIoNka1VHEmwDrcILIqL76
zRi4PT0IUfDVKkXRKhN9PoeAA8Zg46J9C0wfGNY7NFy+T0YGhELA9rkS77xqeFimBKvQT8sQP2d/
GW9j73ClDnohQoQR74r2M8cKh/9Vg3l6B6eO/noJzRafeI+FLdpn2KQw5Ua7FDEmc4exrIIiEZuK
wHtjO9CEVFOWL3LyPWtY7GRAkdfZFVcS166Pd4b2U3XuUa2O9dyA45RhTpb6ZNJihzZDHQmef5gl
YBnvG21iWDHAlQAbvdFYFZ5Mvy8ddcmvgiCrm4WEznRQ2pfZiYGZEdyQiiuQf2WD3Apy9nwZ/WQm
AXci/2N6q6JMWh2iL73gEqNDhm6XMgj67HGw1yb5GZPZhm0HS4mg7mFhErxKWow5QYbHPJye16xd
Vzh636oKSGLh5RJjCYkyi7DSNdJ8Si6nkwqBY9W/r+wbBh7QQvXB6xJT32zGDhv9IWRqsoXEGwmR
VIWxbJGcPTUW4FY7V4x7K+UmZE9NADNQTh0K03c8gOV+gy2OfkiENF0GGI9ThA49uqRLdHHbirwn
NJU5VKHkb2YHxxf3Fz9127S2wzQUJb9hopiEE+MbXx2kA3h22JGhqcGRb2yf8GFOvTCyVEwAy4ji
gNFrquDc3nbz2WprO6wOn68Ry9JNphwX+cNAxB9Ck+iNn43iIbP/RZ7RIgOXTOH4/Sda+N9oW1Om
53hoKo5VPZ6nPMzWooDvBUdeyVwQN4Eo3Y3+m0IfbYnhr6FFcXzJX5kkpsrWgEPe2DtgEoW4r0Ah
R6ab2n1wV/imrgArA0iQH4ngVDGZR6hea9RGo1orVN3U/fSHKITeDsgSeWkwwLu2zIyVfde5mj6i
Z6YxouKv41sXWUbC1v6x4lxpCJQV9UblIXoPoPhW5L1XWX6IsikrsVnN1sVJvibxOVZSUyEdz+jf
xFy34b7obaLOD1it5D+kJfuyq/g2US0tSaBCUODC0AALZpPhDHi3cCBua9K7Tv3qz9D1jugWoUdM
BpmDOsdfWz8Y615oiBzpcHSeXMt0XDJisuYJCF0l1HDxSGLgn85GgacIeLmgZmhkOx4afeTo0xYL
DEsr3h90NYo+IpaBH95vZntsngh4+CZ6Ic7f6NI56i6ZIdWwbjLC1S3VsfRHFSHNTKXDincdsKFp
BpCm50Qc2cGySTeNHwLkqV6Gha8Mi02dZhagNPGS0ef+qpYykiKyQ0+aH5GlDOkNefe0tbYPhs+p
n68WZpRbrHHEC4L7IidAz4mR6N+WwmrilvrFvTCsaClvcp5LbE3BomQo56en0cAW1fRWNV96fOCK
cdmX5Ck6vGNlwIC17AT6D2QZ1tcKoUnD7wwP2VC3sKm5mtzFZROUEtHjYTT4810+wKc1CEr7INwc
iUg2BB6zUDWg5V+SrntyjPqdviMExL0gOnQPGQr3WOJQgYD4cmEmz13oILfw3EmEAvuczryVtBB6
YZrk7Gru8qy0n7C/P5vXRaBd5b/NuslPRhlbH0JXbEu6LvdMhvpH1ioZS0JJm3dYIPY5n0SPepmk
wsUk6liRI6m73lRaAV2UcrrJ29KDhAYo8NIgvVbfL8l1rHfegVtiOeOTnCBo/WAQ/qwlw80UrnMN
NkawA5wDwITBOUiWp5DbjCIHnQbHPKLN4NzGiRcUtZio+ep4qcxuzAmQGXhAnmyrm6F9pyUwuJfK
G4Gv0SISxxxPtRZQR4Xgwp40ETXP9rk3AQvHqazzWftvGSBVDK1qZdRcsnd+MfWdjZfxVCVNhE6C
TV0W1dL35mDLEBP4J4t9UAqZm1LcHzs28HQCZ/aftdkS0jgJ7+KZwaJLCHlcyBXLWyAqgGdaKgf7
Y+RMJBgFI8f3b5XCSK03jnukiywSCsVbUXmR3Gt0QSvamzSwC+NwdOiTtkwZd6xNScsktd/5noJR
GVFQxjQRvvBS6OAiN//TkON3xWylUnEcVblA+mIOIC56gehUmm0WhVP9Sen5z5Yp0wewZpYUww2P
9JF96sS0s5rnIlQPXihcFOW99Q7HtLwv+YMgk3QOzzK23J3x7+j2h98YhT+B1SCGtfQHbcZsoEaj
oTzlgV2/6t+1k/ReBAHbmPfTHFXsnIqXkEehy3FVDIdlxDe1CCGzX0iX3D7HS61Ca+UsZ0ep4Hq/
jGX8BcJ97QQKLXWE9koj7M17XlYN7DcJlsH3pSMSFuO4AC3Efv82gKPwA0TZC2VuN3N/JlqQNlmX
7qAfRP79hg+FfuV+QxqeDoNPbClPyabcZOwJTWKZkIeIOQlBT2kTAWY05c5k5LsH0KhwROgr9iY2
Vp8pc4Gzgk+cl/FJvCYmEW9ydxtGfAPvOmwjMAC62FAmLUjAYixo7oxWH9IBmhCYE+VnQRmiYBpt
2rO434nv4QQS2pU9yFOGHE9rvrdAD5tge+dkUYCD50iLUduFlW+vstVJTlYhvAoOX5zYULnN+LXn
jNPoGXOW/bnw967N0jJWVoBY3W89KiDjPkPlYC86nMgLvHWu+4LVUmVzdLfvAGSQSQ/EZUB+CAaW
z7P4yxTNipNyOP6p8rA9ttPWJY25czDMPe6Cxy/FVztmoOHHJwmx0u3t1y6XzNeLdKaG3H3v9YOv
n1o2LUlPLrUd0Ct6Be2HN1hepRYtIK5/Vum2hVFcn/jOt9p3v30u18N0u5rG82P8xME5hZl7x8Vi
5AZn1HWWBd0qdFPMhSCOFdNf4sHa3tEFmu8/jIPD7smrGio2eSmNHPBo86svi2KXLeoQaAEF4k6n
of5lWcRvKBPCG1gHapEBjwRKKlKRq5tT7Icvo2uVl2gQGGuZl/zxxGX1Gzfx3I+4MyPqeXJx6PMo
lsmnEyq1XomR7SPsAik8eTuI/hgVKG3goHaW7owM3PAC0tU6gHmpqUg6Pa/6mkSRKuWr8tTLwgJ+
1tIblnozRg98/T73le2HTtordu1wGtN9BJWFx6tTNYNaYKkvb85r6Ac/EI/9c4822XlRH9lBOLhk
DN7LkSf+McBU8MFem+N8elJKmZTjvNG8HzG2jw4QcgoA5kzN2TcPKSqM8SYQaw3GOhD/mq9qNi7v
3KlEf845DyxL/zBWb62ZtMBjfPmxCCr363acQPd4Ee+Z4ThHTcGkjP2bffWxZYXkEeAxkVDRecV3
SZaLUJkg9nS2FH+FIMZ2f2966Ea4Qz+qEXzgpBAZrGASyUA7uujajlXVeUifqlJ52mEaU3RKlwCD
mLxi9ePL/kG49xMQzrc0r0RGzl0tv22sAJoOc8e48pJVn6kktaBBikHp1Nc4UtDsPxFHraPaMB5C
Ir2a0Mt2JEnjzhPln/VRwu7cIHfnETDnIcrIRp8OMfzDRV+/0Hw4JYbfcLoT0pP8chHLvmwcKJUZ
p6lJA+YTDTjdnVwhr1K3WhbEQgczIw6pM1LsUU/IWjUcZfkXwUVmVeMjxNgW4Og9FBAkQEV1w+4I
lzZCmXWF7vjusnP8RsYIJ4aWvftRoFI/+lGNpNHCRyeteKMYFFSRFfSr+8youdcK6WpXJtZqOYxr
jhuuPiEwFF0jw1+4DWkA6WMvflslrAE+9E6wuULXZUm6AO6AapfA8DpRtA84werxirAczTXDWTTq
fOXTi1su16wlPZIGAZGZ285AUtGFnVr0afM490taWlKqcXQrys4ApJ9Xgt4bwxp3mSi2y2JTsl4t
dWLfpzkFKhAOx5QNvk2jxCyteMuUy5ggYzs10WA1ci4VQpQU8zJSSr769bFgPPAbII87Hp9WJc1g
w9rBGp3B6ukuC2BSsRpN5GxVHe+sgZwdYKFK+luNw3Kqf1ICmQtoApvBsKN/d8CsiOM3xXSA48HH
S+C+0GpfQN3PiPWnANqvDwFYvmYoTzvVpOEsLWsU5BIijQgfZj5UkYmkBGKDPbcB4OQ6uT67V6Oz
GeCXDrddm+hjOvmvc1H/3plGCw+4/5EV/1VrouYGxZpmSINVeH783qkJMdAGwX1nK7bxIuIMEQYB
0ELa0POzM6JU+EIDZFcZoSrV9sGO5ZxiGkeT1LFIgL7Rhdmeom+2V/yJ/x2kwYarJs5A2akEoQ0R
/eARV6oTVs3hxpk28y4lkVNdpDLcgGUQi9xWGzSw/8Dw7pX2RRkAH2LN2UjjJjF24DmjsG+lbFgz
3ab5g6YjxnJxeAqoM7x3t/PFnxInGZEFizo0ih9mbDzZr93W+AferxdOW/fiX5omr5bFCDZiCCYD
CewTdfw7zagibLH3ZRyMeABhYGbBkPKl6J+SAhsrQ5Ee/UDuIk4cyGUtkWZ8lswGoYjPTzvjSWYT
DdfhQZ7nnBwJXdz5tdW3tCTEvqDqO6lD42MwEP2R3K+5V08dH6HQQORtdtu6Mpqq+0RJslYJ95om
LdflfJKy3xWkB5qqpNwKwrS25OhNOOx+gtt8LjwfqAjf00k+MReuXO3cIRP9n3rtv9Z2BThvM29p
LLrKOfgoEKPdew0QShAqltXYL5yFpzwi4bkuwU8PmTDWYyTTqF+oO/mBpLhpwokrnCfWwJsLgPLK
+7AW/eDZ4l4I9TrffTZjditOHzzbsUsSq3VBKK+TelSJy8uxb6CubALqBFk4AS2usftt6ZpG0O/g
vgjKIEij3wzQpWdpSuaCJK+o+BbUr8udxLs4VrP6cOl8QX9xyfiW0gVCBjFlF7/IVwN3TSyQtpMA
lvziAQO/SFLkpdsLaVDPr0sk4rtXf+kdbSYHstF9dBCOcne862MKpXL17C97iMdMMrmm4dtmMH2Q
UHZOMU8zQBBvTXW+rskd7VTJHTqm3H71OAa5i+hvIfdpSu0wOHH4DLdrV9WQ4WfICmLyO7PZ6mFe
KrqtQCvBMfkapi8Kgtne+OwzgOjU1dJE2OrbV0EeV3h7AIxikx5w1CM3kw+zKGnDp1q0r3Nb+Wak
NVxaoU9AbnwNOONIY6EF+9MuzWz1Ymv0+QuYxsH8ESWIXe2hov+maW9VQLEZW2MVjRwll8k6ZVgg
1+1cCzFrM9ldO6MOkLhSGbCybDeLuJUlplmFTIT6aJs6cElvaVAWh/eO/LS7Jg6qi5cyg4CdpVGh
WxEpgyPlQsu7EDkVsttpzx/vFPXfgFFfBT4IDnMa48pNLdLDY+CPEK7lc4qt69gGd+VGH16PBFLD
nE7xia03QD+mM4iURr4DmNuOuibbqAb8yozg1aHb6+lQNeQg0jBwlQMrkxYgADEpqUv0vDo8OaUk
HphUkN1zCdABloqy05dFt5LnJKHjpgL1D1LEdM5HAi+n0dTMOPJVK/uLorB7RkeuU5QoO8KOH29L
vmlogWKeTaALCNXKyPTyx+ZgGKli0C0OUiwLIR6p3M5CI66Ju7uZk07uikGwCraNGahWtwZn1ZRx
Uu+5VjTdenP/cAzSuWFjmVzIrBe4iN8DkE3cd30WkWDHqIqjbc0c4pkZe6/pwaUJXhPXTxyUsQju
0lEvdwD+ph9S8SUEr8W7w7yUXyQbSSvdPgiEGga4waiInYN91ZkVVYRG+8N/yjZXRG8ZEjHZUIsO
qtPDwgflM3vsJVsEbQlGSENBVOv3aEDYDRlYHpayxChgfyBP1ysKjRHWXpcymXoN8J2GTCYvNhc4
9EuCOZ+oL8P68FZf7QFg/CbtkR+4R40BCEap3Kin4QsyULNHlnEC+VzPZWrG7YyjtVFXc3xo8/TJ
60h2GmOqfa8O+HuT8s35b6P8zZkTQDwBfxMf7eAmQkz5f7x6zQ1IgdwWYznCvd+WXs7huNtBPeI1
+nvLPKFS7fxPwONRk+lzL4eQ8MPn/Lz8+lgWHGALpwUhYDC0sF8rxuRMwkAPDwrP3gpaT5Y52zMA
GUCxE87sQEt+obSh4kr3FZYuAUg1GpO/KIm34J1Y78w/eU16/ufUkW6ogkFgTHdd3tFvi7XO42fP
AFp+NiFmppZMDyrFq82gbpmWLAaBQ1ENlrY88n5sPg9nkG87WalL7p3qyhARNDp94s89e5M30R/P
f5Yrv2UEOfC+NHc9dBbQnCgBOFozb64WquGrRSH+fff+kx3D44l8qQN9hYZXCaZu9a1+rK0fWl+H
iz2rfVhdmiq/Q5/z2KzriboKUn5kYAQydliS6628ojTi+54YnEJfpzYasCp8jm//DdGO+579zl/d
l9sQHVRXREoFL4pGDOUJWaXsvhzEeQn9NEbxhAdEE9i8hPf0d5hfYoaI8D4PKE8NwCuyX1kov5w6
1DISDr6zSGYwhhs/ZLbLzN5zk+L3jnpfsMfwXiIciWP+I7Gnr3fSWfssvY8jobsOeJvVi17/iXSM
C40tOjrAVdRzBDrNqSs/UtJ1fg3+0CSHDPcnDSBE0KsrVDQCC9pkkPdm3/NqJE8reuK16EOUnoJE
45SuSbdgZsHvftH7ZMUAKblhtOD6BN2im5OaigjK3o039Z4VplqRhYBVK+qGnK7xME+wtJxRCzgI
/evZ65DtAZ9DuXe4QYRGjEoOA0mwDrUbNp82brMvmzH3w8t0uqXDK+O7ghw4RrlALvf1gBO3G4zT
PPP391BtHcC0RMaOwiGD/iVcAlP1fL7bZgFKZ+QkbEwvBwisensvEFhmldCj8rKBTMZYW29F3ZKc
7ccj/NUDUDSWNW3/B4ZIU0jXzUJzwcSARIHCwsqksR2U9mwxoaJeaI0y32qGnklPGfIEJ3z8X1Jz
8PnRANp4NoMC62eTgrQzDYtqfhTnN+QKRUyDP3Kz2smfwK3OXgOXSy+/odsmO7KucEpwhEUG4c5w
xEvIAo1/1eUfTpPXK0xonbtpBRVtvgAfsc0WYiBdyO34X9XcqZqXFJ2VRCyEDb8YtLWSp5jzH3mB
XHGOkvpwdvfgDRhXWe/YUOhEJbqKM6PTorSliYQ2PR5xlvUIuzhlALsMKBkBnBOJaPtzdpGjGQuC
jA/xjcZa6/lj1KGXh+sD2RqQ3qNOpjm7t1y4mbHSq9n77rQ+Q6NkYENUoTBqWnLJHk8733SfHtfg
kW3zXYorWWMvrQX48/czlcQ4X57ulCjLmiZbjsYmFSEQ9yAsnUtpL7SCS+pjZQHV7VyHgrPRLqtQ
UdRWt9L/XUvxnWOXM9dCQD25re1M4S9DQoWRfVBLxuD7BmKUFcNdsbTfsgzSW+TL3xL0z+daaKX+
4KdIJFc1bjIFD7i+0ApOW2QBSWpsbM3fc6mclQQtyv5C3LAwT2TtzKVdraZAmPlu707LrlWY0Vn9
TZg80mWNkz0mwr4LqG05PqPxWxSrZi/VZl/ydKmzyIhq/xP43bLLksQp6jtAU6QpWnuK7ZxYRUq9
3SZTYmrbiQ56OHuWGZN9h1IEiNuRifwb6i+qNv+Su/PkleUaqHpyrLgXyYdhjlXlU7ZF1T15kgGe
gO5ODCF/h32RPVKiP5jpOsz9DPky3kul04julexpFCBC8fV6XlJFfnpUrkZei4wpnFnL/YNH4taX
pBqNqVcDFH4NtYeb1SZI1jOpxk7n8wpduTh8im9td0J8V3f3dJkKIBqcNr+jG+iQsa4er7vYum0T
E3KuXMnHev7bS+/MtA6XK0x6Tih9ecbE6Px3/yPZpd9+GvgKN7KQh6M2aPxTn3gNmjUlemfx6C6z
XFmCYXztjaohHpDKmePLKs9agNEsX2wJZBZG728IQCAT7io18bdY6KJgcfcle9Ws2/UuCWCZCqRF
xDhM31db5z5f7OTb9yBB8Tfvr8Njw2nJPY9ipn7VVcFn+H5PfnCYpjDV/LzeIeOsEzLhypH/V6MM
B3gd97uneiqfH+aSuaLS9eK94fNXJm/ZsCS5RV8r9cAy0OFQryeLmYP5lIVcYisAfCsvFIg0oSBZ
zYAXxPqq3NGW7OANuG/0R98w5ZtngbAyOz4ictM5+4oFctqj1CsD9CyFnmJfnRN3/xcVVt1ZDHAA
cBah0OnjhLSfLXSxEBimEatXxA57W/Qy9AFqCrpk0Uk1dKTqJXgNIIGN5mGrKAIZXZ6K0NhoBUCX
iUwKU9hIwe4GEzgGXm4kic+I/bFxfAqa4BJlSGrBkOQZtaZZ0tQbPOJtInMZaKIg8zIpzgh8CxuQ
rMkJnTRCwuDH1mR7zLexjleL4gZxPQwCaei9QyXJaJH+LpM69aGhc4n+vKinkXdsAvHhEGG3a6V8
1xSTHoU+yEV1J/NycQEZ/YXC2GFEDwZcV9Z0TUbNnpBHOzSFBSkiKQYYdPrDhiNceqVg4/XfFrRt
BTXwrYV4nMN9wvlwAFrcxc9WLYQm99GcqrqbsaZ7ugQCsOW0GQVjCS0ag4d4bobI61JqhZ4JFUvc
6+ndFvkLskJpcQpKeI/eG5zm5zHxGcdYbqmbbKb3LtyYzPjQ0CBJmIFhnbu7D/Gn+zIZtQ1Yujfy
AVudCxOXLaahQHNxuYLF2i33RW0HQjAuCRwdDrjnb6ZnCC6mvcrVP8yq6/YJM6pYqUdEotEfIyjo
3PmUmDIfHxMbe4cTUQfQsPODh9j1OVa1DbAGtLL+JmAEPGRx9HmjPbldqfmA7trk7U2xhU0cReA9
A2tyW5RXFRFk6uGF0suiIXA9CJRnl52WQ1QIhKhxSn7QziHINHVQMdWZho9c1VRO7LME64aRGqlL
ZTCOyXDQzSG1eSz6STYxNIhity4peH0NlySWUuqa66zfSyjHsQdXm21SITVXdJpH1azVFz5cEIbv
L34POG1R1Jr3hrxfrCPhhsNtVVxEbTmJ7D1y3zQgnGjB7XTLeKehYx4c2TJSaxZn34dU5/4yyaLy
B+q+tgwYDRz/1pSvjpobdSbEJM8rcUUxwhT5VIw7o2vvmJoBVPa4vvglV46y0Spmfu+vm6upfmz+
Id0zH1P9R4zMZNdzMgE7pzd3YnM8zgmy2aLe5LQJQFGIO0rSHjiSiPFfGzGV2BOScjuciJoj+y7S
xhdvYg64GYTU89B+LFEm9T22/nXlYaOPd5xyZziZcqX4NWo6S6XXv6GOL9xgeuDLlcfz0gV68wRW
LTnQd+HMDofUM9guOSFE3uYae//+f7S4EY1oKxhs+6QUhBhGVsR3olNIhSFoQUTEibEq7IiworK5
CmlFnuTZT+m/mAzLMAZXjI9cbqVG67huQP/8aeSoBGTy7m5WI9zTmTFK8O4+YCLzaBWVbv0Bw5G4
oART13p1kPvxD41hKnYr1Xa1k6vEQ+RBRO+Z4mXmGAI4KKjp3zGP4WXd5+eGgb1Iv3hdWfftnwkM
Tm0HEjwfWQwPmAVPnkiSG9dc2IsCQu+f6+kHyFZNcOFVps65oBDJMtyJkqypKaBvfy1SdT9jRV9j
1f3PGlI//zcsA/xd/Ee15udCjTGwBKMw3NIFoXitGYWrB3Il6cP2txpL8iGKZ8aiMfP8/h22KMhv
SoK6mjHEypMH44JpAYt5EivPI4uXMElBe+CHLeRak7UtjjMvX002acBpMy2A5kFS7b77hfiFfwFm
UotDq3WKm+VC9QkxNxmZwlkDOxQeEiOMtnu2EscgSSYJfCiTvm7tOJ9s7Ss7g/Bwwr+BJYtlgDBK
JhAa/WdEKRAnsve8l9/jtnAyi/tYIwbgE0L/KytJBhKznHVNr0BcFk6lC0Q9QQC7XTteR3FA12Zo
9Jtu4oRhMPW/KpTGTKDKSFehpbwcwKKg9Hlaj8pS4QUaF+k/1zFbtNcx+11UPXEz/AkSm1gEZynN
g+p/tQC7VO0nLCfcGZ+OO/QNzX1jr7yfZoqadmRNmlnLeRAEjxcxDL/C4L+JqcsCR/C9GAb9ULyD
OgMJDZiI7XWoClKrQXGoWOh2loDwa7/ozbda1FzO4jRlPr6FqWZX9q+FXW4KqZHWDR4TggT5bmJm
O8lkAfw6PFS9+VgHCzQvOVYf2cYWnQ7FkdSbVdMGbt+nGa8OstqFRppLZk3737XIi0fxDmThlhWq
rNYA5y/SX+qA1lOSOyQDeM/nK1FVA7ZvtXruOLlCrNiKUv25rzuGUSw9drNPRR/+tA6gzooWObd6
FAyy+sD37sODI5m6CHO4OTC173ME6ztI+24jlyUYJ9tLtfZFe2vXIMYMJxhvLflpCqzEOoD/nfyF
e8wwSo/VTMxyoFpO1ZweJKnfZly1KHGEW3N9aokgpjuYDmHhvf47GJcXfOQwIPII/4wnyxxDS+IV
BvJoVoSVMdAHPq8PPifxSa207/nzxVgtdRoZ585f1ZDO7PiiajBs9F1YH/Hq+SW7Oao36TOye8Pg
vXq0hFzTKRwEcpvIryg3x/XxRPafmgP8glttOu19PE4x8t82c0PYY9mv56B+elQnyFqf0yuATcNT
/UI+9pmSoqufcpk4zqi/ZiCv++PybjVPuvisrhjo8vQwwdBN0fv3Bjrc9K7BURmkaMupWOMz+46M
DqPkoT8Qpu7QyDn+AkllOOxP80wT4h6YJKIBHXb+qDsRoLCEwCCw5/JgRB8YGsbbwI/t9rrfxZ8a
8BNWs3z+H3vW6noYW1QEmg2Vd8O9SDeMFv3AWjt6dbpLctzBoc3fkw8YbB+QZv5V22f9fli07ltl
apdpjCmPdycfHBaBzl3fkiE2rm8MPJJv0GFALaVxkHEpcDIGS44g6PwgOueSuduPWWumPKru+a6B
PEDvSbZ0vdbSKtzLdjHOQohSZDU90w5yVt1z8oFsFhCgJA7uWuu6wSzbRgBXfBcreQNtKEqOIMPV
HquZpZ542bShchOt1qfj3V7Cs0Izs1FhjursqAt38Zvw1aFmtOWvzge5S/nx5SkgQnXZR3tYOsSB
CgaY+90ZskM1gAhx7AuKI+6Cffjx51fnEW8QmWqGVD2J4ZZQXHm52HYmAHPPdghapf3uWOLLbt2T
j19gZb9bBm4OYo4kNFRZ8QV+lBF1kFFP6rAie2m4chQslT+WPsxICxkpWXReS49mTzGfgtsUA4bg
mhDvZ6R3Ua2mjg2P7OgRC0inBF2FwAcvKK4hgS8GL1KOO2mlbyKqHLZs0qeT96Skh42bhbxQKTbW
gipkA3HatPz8WxNHYqG9YK3XlNi9KXLRyh2pUg3h1r8esx8nJpgrSSp5monQDk/YB43T6CtIbPsV
YZO1GQSjRC7iAczMjQ7OdXUDEnLPXiQOoek9M670hDf4vZYt7PJFCIcKm7zvhHS2ZKwz3Lku9y4k
5EZ/jyLEJZlSUeGM2PPfEGPDAZB1LK+psmUhA6h2oHcVL9rZh0jVZECfJBe5cUwMpxR7Ya74ytFQ
W5g1nZaa2yM3FL77WQijt6vzdiVXLy6oMUyPuymPkd/Phk+30EGlhpllR5E6fkY+JBGjvjeh1QCs
j8KjJe5wyfVoQX1CGeNME3PlQiYwpkmf5jx/Sw3WZBTutdaRMh/nfAohO2790MaLPHxaFPmyhE/x
JKTZ+3ZBOPYsFFSXepPsVcEOMo3NLhGcql7adcZGrBLHdYtNJFTeifZtJbN/VGOC4Fr41wZH/VUA
ds1ZRugW6Z0kdv9ViRsTrCXv6UaiJo3Zm9XZD6Mzk1cpOtXX861NJqe6YiM+qvnd+jy2u5mPrNSK
dXyoxZwqljM4XAVPH0cNsp80urtDvHAMx4pHw+T73035ax8IBsIj/dX/H4v5bJSdVZhj5wy+x8df
pvqEmWuIaWhzxi68Q9sIgJRI4b+KXKq471N33PH7cDs4mjGOUtEHPcssJp0T1wjBoanODhzWlAhc
/jTg7Lcsdzu3uaeb1hsPBkue8d+Wm9UtgELj/h+6KnRg9WIPi4icsQlgKicw3C97xqBGeh4JoeVp
caE+iEZeESMph3C6hSQDUiwNYcgSokvIlaElt8cBURYVan3ddfpR3+frJLZq8RD47ByRip8nImv0
lRcNy6Khgo1uEMpFNgzQ7y+btkiiJYWzYVgCS4FEAuusl2hW6pi5L+i226zd4iePIKnB6QPmX+ML
nhzEzKhR57X5bJXU2JxITsB/gcOLiGWKf4t9oaOP8IbcjX2DojHB6APNOJ58efzogKkfR1G65bDn
9I1mOlXZMzj+fO1aRn8/3o1JcuzDUD55fTtthW1T47TcswCw6/DX4m+mbgMYxndHg4mz52lDVg/F
w0RnyS3SOfis7bcUvt9WIrS1KeDJiyKRlEA1mNXpexTniDmjMen3eo+FP17UmepeEQ/TMVKyrRsj
dU0jAFNljtT3Du2jGuvcR2UeO/l5KiSYsqG9k6y2ei8aLIPiQsEpfwGgfCT65nKRPlpTsYEPMiHL
k5tNjCKAIJKhllM5VWGahs6ILsSJyD/OeOCQd8w2puwGJcycP5lVucdxUz7kFIpo17YX1RxJgJz/
Dzgnzz98UIpQmHcQXy7Tjj5xr9T5V7lRL7mgl49UjZ6vX29ou4JGJbCl6Y2GaUkjeAuY4n32Kcr+
LOKl3PExJ+vPId01stIjMd9wHuXQIG5/OshVl0LdukOtFggytueGAMc1AMXM1jtFB4sk2HlHDoJ1
Q4T5AL2lUxofSX1QNcyq/OWtWALOvEXz+ZxnmewdCELwmThrp0EMaytFwAzQl/qmx/cmaNByy78y
R2j2zy14YIL7Y8anQbcMRwWN+C7PdnHAACQQCCW3OSQiNkHlrzP1vK5nP4zEqKE3LNW/aI+XK5+F
SfJcjJ024NrHwXpkyY2eMmMghL5ClDh3tawJjuYKPfOepFEpnRGqXMT4YFLITV11NAFGrQYfbMu9
mClVfxnHwfobGOkjcmg6yRv4TLnlvyXfG8rWfQheHkV2kcNU2lzFqOxG8VdyAvlKItk/iae/+lYp
fcnGRZ6OYrE3COjPpTwVOWpbHPBJc+ObJi1Yyfo9qrDj9bzPAIDP9M3K+Mb+N3kna9+eyXDanVKt
6N4xT5XFrmyMuhOHS3psk8fwhU8Lpc8dc4YsqiFK4Z2X+bhC8PkgUR/OUQd6aQICUOvRcVRoV+cK
wPdC7nxZbdJS3UZPcr/U7YzRcHgyZVSojzbSsrPcwPme/y1xWJ9qEhlPA4Gidyj6O8ygEv1NCSWZ
8QtOSDk5s02lnC92mWZJwfuQtN0D6yLYhelG73TXm2ebsUZA1Y0/GVXh5nfcDYyIv0lJTZk1XmkD
gajufwMiguju2lAfqUQZjts/8747f6pdbLbK7gZPzi8X6olGienYcnzRUmHRzO7K23X2hNI6GSiL
JyRGtgAm96rwUydoaRSrD2bSL8CJiR585zm5F/may5ETAnvamJyzqS16bieVypCEVfa4zqpk8UDJ
ByHoFv3xkbgixgOELeEEm9Lag9tv3zDQi2WwL0kVYGHD5E14uWDEQABLu0OY5mXUptXwWlvmnO4x
mkWMPAml+0IK0obQuz39hbhGgkAxMaDYoLsOGXDJrlhAC9KcCEzQXcJMwGOyLRNYreoIlfMiNhtf
9ax/GV2EqXr8o0+fjgvygwEwvqhRO4NB3j9MRS4rmAuGSVqgPt3iKBnqt2MpBlXroKsKO7UdLLA5
sPRkmF9OmYOgjnlxgsrVhkCXEZOYFX+OA7VWeEUVKvXz+XwXfvaGF4qvWGXNaZt7ncT8gjF5K1xg
Zy1e7RNwkLuuj5XiaTc0u8a7C3ZTZr43cIbI/zo07Kks4bpKOeSQXNmmCi556AkSFkJpbGthkWAO
Io6v2SidQh3zeTQ7U7q2NoXuqbPhaJldo6ecB7fBNyocFDpP+bTK2l7Ir4ZFElMk+Ju2b69z4RI1
8fjjE9hOZ8viFLDjLKp6LRlRPuSVlE7L985i721m7wCr4bkPScIjN37KYv2PZ6qtNrYqpTCPhU0q
oWmpaSHx9IVbsXcWJUgmo9pcGeeJqeRXmZWVM19uQWrUh+lgRtKB8h4sEtljC0RYTYK0UXTbsMlX
QhFQ6Y2QHWFcwgO9hgeGmqARfRGAKuIP+wMNwuXOSW9JzFyvieer1ygjrW0HWFKwf8m3Qc6M+ynL
EELx+tRPEf7aIFuAcoiBUJQ4HlhjBZTdY7F3Wu5SMRuksVxHfGjO0hXtrfsHLpr0ke0tdbcSm9/R
1uOzMAKLGainsKdOmE7U5vHG91geu1r2nu8PRAUvf+ZW4unDoJkzXQJ0kpYf+EJNAZrLWRnRLnQe
LQvn2y0NAyPOZ8SXtE5+KWdLHlmDur6IwCkkQ1ZcDSjyy4LX+l7ahGAQGUhU+MAj8vhF2TsUygDW
0U5jLAm98AuZtekgyrlFHw8jJ+oBFKCS73bjlwMUY7KJ380aoHvsinQshuyksdIJrjIGKdpigCs1
+/+mUM2NAeV78KjfjF63rI3uUEve/eRhXGHDIiHAeCVAWkAs/KPPe483mNIgkTtGVN07H6HxQekx
X6wcRsVxP9tHnxWbvcctptN5Fffnei/qq1foOGB661TsduKZiR8ElO3sQTdTmwPwY+S0SOI/CBfA
Ea6wa4718UBQE0jpoh7jkE0lv8E/Zk2G0NrmP8iOZ/QwblMIPK68ZclKcL0E+YyGP996dj+2SvHF
JopLIfm4W4uITLe+TZBdlAqCZXbwGfhu/ghbIlshnkVT+MdI+owsuYbsMhAK2wf4YRHJLZ1+YjxI
+aJ2RFsWKHyF74vOmV78a/O7hywMSe+lCqWMo6VO4cJYQw0zSb7qxpfjTd6y0onuBVtvVlEo2BPA
lKh87TnYtY/xb+nvU4wx7UaZIfhgBmmD2CSAq0S+db+dBzyJTZ+UTj9Cojy2hC+YmlOPcqvzqwFw
f1zhCgyKY8PVm90DRJWUQsNIFBO6HhI2sO0/vuZ3duFSoR7PV76DGRN9o7R5hWn9slwae3s7XSu6
QyJ+gc0+nxEfYGqpz4UwrfCsJaSWQoVOv8zNOyGQgL/ThqMd6kdCr5lVLbB4Ok74xJ7eCrV6XQwN
gYsOrpu4rJU0onhk1Mwt754v2SCUHZaFn7PnwD8UrYkw3UFTBLdH60dbsT/aKkVUCoBQggiioBYH
xukPM30+aWAPe9qv+Jv9eoTKJuE3R8dY6qcXv7PXKQIMbCGiqlY4Onaj4SlXE9ds2cpaEKQzeaRn
UOdxxvvy5VtEPDdkkCDGhoM94U0U/+05slMCRPxjMb2L3/KvmwZLZmHmTc5ppUBs7J8h2VgNswPO
oSr+Oe9YR2mRL8PXXaPsmgR1gZP2erbTleVun7rwn8g/VeMWUBs4WzgtvxmbzfICTXiZnNQ+CgV4
5nWWcoU7OqSannmIk7xtXArkp2asqz9nBrKzbc8OG4O1iBHOf/cTUsgTafHo/T3FmVq8Y0BHzUjC
mVCQ54UhkNUaOfVFnB/hDbQxEm4t7kvW6mZz8ohKMhoCaBalhO4bqajtNwrpJAbnLKdM4Ie776Es
MSQBgz1y6jNXzQ7kNmZGJHmMmEGnCVt9ZPva0vhHMYJK+TYZPd3WVtV380XnpurHb3nMKw2d0KeB
pCtfnmabB4SYXKQj/NyPLO7TOAezxDH8k1RJDuHj/QkHYGzH8azCKdB5ULfUlJn3WleROOo1A5jr
L/SeHGf/DrbE+3cEPqknlPD+8scEq3jDJlWnepJRGRRzR7kT0VG6JFuQaQutiNldtJzXeFhB7/aE
S4GgfNLxMKFSIjF5LYy64g1MdbW2/PjAvq+Y/IufTjBGPTz/+KtqcVYHKyfS7V0Ogjk0XBHjXF3d
exegV+NcArhgB1nKT7z2x1nXDWzkTElq4cFyVecusGdUJo8kyQpmBF2FZp4j94RNPhqjXswetrni
TmHdPO71Er2kyKtiniNWjj55AAHN48l3U9fRb1Mi/DJ+LdrEBABXjRF66rjro9WEBwuElUhbpuwk
cAaTovlh/MiMKoG5BQcFy48H4J8TQoOOWD+ieexio8U0plmcg0CzdD5/orkgcSbJba2i6HvPunyL
fkneKxL9s5YZSRJcrC4n3xgya6mnq6mh9YgOxXXvAsanBkwSBudHupRduSzc8M+f4sk/VfefgqDj
ysBCWl0kH+aSmXu/YzWyg56ssMuksyZq9h2KJPhsphi2cRPFN16APIandAtKjh8swBrBEjvlr9ki
CeJg2TlVrANheHjCCoD2eMx68TjQSKUv8gygKFILwipSj1//dfBWkuvBngiqMGmrjO0m9oYsEDDo
E0CidmkrEQe0RtmNRJhvqUw8s1DkJWzqh4XgUSDpVpf4zcRIAeklmLSa5buyDf1ORxXQRGNeendc
exl9VaJuEjF6hqZ2+kcOTAoLQTH3pMN3Pyw/qDorq+iwcNEtjF1SOr+On+6yW0izOYAJLpMVZW8E
D58YM2b3PmS+HpxYMhA2F+UrYysKvz/CBy01CYiwG9CLlmMBhUlPXiEYx2qXrZ0FZiCmoet/0O4q
VrnnsfgiDltWQis6Z7Gnzk7nl6Cyv78VGPz6L9ffYkXeygN5mBf0HUXrJmmirnI16zBRWKy1D13X
N2eW40nVllJPrXQfFkdlvUQpDTVsvkveKLPDFHbUAm5nI209WYLD0tQRKuI6B4SJitdDtUrzkK0B
5zNbqHKZ+LsAxpOUMH77e5HNGz6PrL1dHlf4rXXuQbiecxr8uklQb+v+gQWzx0dRUAx/I5ssmuEQ
QVelpqB7ybe3rfH4Hsm2oO0mdMt6CYk4KmAkm1SHAhSaAzvAn+2zCFf/zr+SbLK7WNtV+PkLNoIM
IYqDKKN3qVkGLn+8Ti2RN/IG6VzgvbkCWibvgp25npdm2Wo4a6VlW15ePF/yY/KLP6wxmrpawZ+9
CmX7Y7hKFkRqV7tnEKnZEG0Y44a5XLs4j2+jaSVIPqxW6huVsQ15OxRL2vu+67R6G3XFc477K+Jy
SrIJnmbzgOFRJOE27SFmy4vTdbVNu+bpxz31X8zpQ+SAOKGv24OJgpC5uTm+oXmBXJXz3ZOT5pix
4runesW5VwDUkAYQvWn3RpQcnMLaBtyEjrG1VzMnOzyvEkQ0FcRDk2LlrSZ54zbOgkS/dpNvCf5S
qM04zfHmfUyMQWCskUAggpyUrObS8tvIC/mTuXADYGwBAgYZhQxYv4LATCxMz8BfN0FJLHoEu5Ht
RNwqEIqS4743r9K8vs4whOF+Frq1e9JgFCyvPmrFSKaBHG5S5wCr2MYv0ga6VMBiG76wQuPP3DUo
Cd0ex8I9xjpl0uXjmuRtTVQXYG4mharmEPre+YPqc89tmj36CvrGg2YDdBKhT1BWxnqV9PZqNpmi
FergIihedeFOafRIwPgS4oo0o6fQpHIuQnv1oTyF/amsVTXeeuHVP4hcK3a2BkYdxuY/j+KKehiF
WOVJcPY4bmPc4iwo6MdiweYpIp+3BWIWghCcWYJa9Q7Dy/kI+cow8x1rMzJeIlplYOJDyPxJ2YGD
EHqlfJUKCdxfCPuSSJmPr3+ip4IUrPlyvktxGg4TONqbURm6WrMNMKLJp+oA852cJ/jrnz6dywNz
ucqCWYhCHzKWTe76UOB0qSceNFgxcFa15wsYKObZjvQCCZrlr3lWtVp56O/lVJV55bu7PlEJdZ5F
4rvcR+tnUU/WE7fmYnSUf2bo58oW5MaYm8lxmEJC1VXVtDfFJkbBS9uT9wg9BO8qwbJrw2wbJuRf
B5cTyT2CaznZuSRsZeT9xnMHkSfMc63Fg7QI8vTMI83fNB7gP2v5VYyy7NS5VLRvci1xLbJj7n0b
hDOL6HhZ+ndDE+Yclw3zzaqJyKmlo06MNoEAq8TAQQSVyo2ShEQTJTrB0sTTGEd6llmGwwnuZIJO
pLtrF3GW/g55VJ/P3B+Ev3q1Qpf0QpQW1L7KAy7dxQpEjWwAS3/sMTmS90mN5w1u3cTiXT7TiTgF
ZlDxJo3lW3HEkBD6MQTCzVBzmBJBjnUUwLpiBV2nR9yChXuelZrCOXsYUYY4zUKVKF+GR4xZ51lp
pB/jsF8+YTK3aeA7EKrYRVPipPCl217aFcKbLhBAemX+MI/wZ2lIMelM1wxxRDr2K/l1PMhHLay2
zypzYpL/KRIZiyU1u/pN74clIPEqmNOg7HnIBFkysUS27gOB4RqLKo3tRImVTn4dmt3DiGn/9PjY
ArtAAbEBpLz2SZA1jyY7F9caYcAymm25ksMZ09ELCaHiOfnCxlV2nb83mSqPQAkdDMXNq5Q+18Vp
Yp2NIriN7MFJxbbdH1KZXzAssb9xCDnXUp8+jcv5OTFpt3fqs8BRa2V/fwU2IliYcR2X3iKiAib4
Nssl7ol1KlM96Y+u0C3vozqK7n2+0Aoj5nEsbGdTKG/8Jr8oY7eursmCYm4vc3FpP0dRKVELyo1Z
fVJB9RwErLlqCEsWHnhFOJcQzPkksFKdwUtHJSPbnjkFe3Jb0B0JSLOTpezYe1ZehY1zsjCNjuMw
Q/2GvBdL2rJdZaJajKUAm8tOAR/iFVLcDleCkZndvEY7vFKSRm+2ydvgTChfwjtUHt0x1zhGW0uk
p4vBWdly3twQPmTxBoMa661up4/AgLHl+EVEH5ZPfvB/PIIkGssAL5fkPaYFvFmkTPz5rIyi8G90
YyzJTtzTvmO2r1+8ClIdg1AeECan/MgbmN6G52iiBhFdtUe/w4UrRlPMWX/6kly2sB1kqFMy4MaQ
PYNDGTjP+tj038bM6Ca968vA9ONGR2nIc413iXit8yioT92KQ3hQDscdIve/jtzkAeeA4Bmlb//s
eZopCis7eOZALODXVqKFmxT3CMHnF409R+bA1BhPGE1j4eBB6BJIvPmpZkxGmQHU+kn2DkSMM+Mq
K7Ky7D1tT9k7US7IP31TQ5mmEkGOsp1P5WnOZ5ePbVqINejAjWu/nKrymc+qwQSRTscCgaZgEgBZ
YoqiK1zyJxJmfmsbNSR+rR9QmLhRb1bcDM2S6IzHgpByhCNc+9bR1k+p0exFGkTVkAEgQ2z/hU3c
6RjXXoJRjGA8DQWtWPfH+1DxYf2FJZWOUxGDVAK6k40OrsG4sMath1wDKdyVgsvIwJNCGqh0dQmO
FR4GYf6LjPc7y3ZA333kWA8MPzXuvXHZsBtJcqs+3UHG9QE8dWkbeGC4iGQFFPpKqVEbnJglfJSb
BeMHFfSXd1d+ZBS8bHHeTgEnco6vw1d752QB4bezAwRZFatiGI9bZpsp1jBM88+fcX7IBro++xTV
gCz8VNK7QOumCEdrZIMyoXh5SStLO4PiB9FAc2ggn0KGhu2VO7o5cIcY3xsOVbxjpx6ai07wlLQd
GJRz7hxw8lbj+fxrtvkBSSX+QpDTVGuO5bhuJkn+WuGycBlZJQ3XnIQmCaDGCXvUHXe5Kx5hqcam
nr1eL6EAX64/Jtq2kQojovYLCwkccuyIdDBjMhqqJ9eLip5K0utPS54fnGYMjPsCTWAocqCme5rl
VgWuKvmQBMCn4b8gYBT9ty4VwLG+d16Jjjwys0o7rClvE0kN4yjaeDwIBe/TywYtCS8/2g8L1dIL
gUgtgvPsVsOsfv52lFpPBlPGWd+KnI8aF2KHu4gD4d6UQrSS1e+/KDtg8Pf/htwRr8yq8Y4fludL
HCbZ7hRzmgH7e2vrrssPpEbN3lQaSUK76+6ykQNWymF/o8m0ADIqOlPrcF0ZwGtLAOJJVLmiPrVG
v9irdJ8si+ITvyNUsYyNHVxpTIgB/2XuDz9ODlWR1tUO+yKPlyfD2FoPObuyJBgZ6rd5Ob3m/TDe
XW8YlXPX1XSzfxxFPC/vrKw+7tWGH89DJ63q93fqa4N6X8bQKnBQg1z26s9CNcCPM7z6+uqQN9qi
VCtkF2WSEri4Ko0tWH8qg1mFsFYPsSxUG71YXOosZsdffE3l2N6/qzKD9jJRtHgoGTmsQl9Qosx+
4zE9xC84u8z+rXFUW9CwdqdINOR26z94wOb90fj0RZiiYZ7itnSWEyFa5vYcaDCFKiQeQi7x7k7I
u87S/CZ4p26Lxbfrilvn4er7qDrBnT6ykcNdViM9AF8S6AOBvXpDlxu7QxVjHgbLBjvGe0T87DKs
fWZeB3REO5vvSez3wRHAP0KZA6f2K1uZlTD4iWxcQvIAIwbJ5kfAAvWeQTtpaNT/neGcg3zc5d/+
DqAHAQrQTwcZBDsTry5fBTgrB0g/eJ1Oo6Cn18NQb9XBT/DON8gzRxp/vBlfvu5RigKQgXEVzGMW
pIUtbNk+wjZd7p1F7EmmSZdl1FoUjg9uDOTKWCm3iiub44mDXu8e3vOcSbN+lgmBoPGfxMrfUdXW
YZZrL5d2mjusCYFNRYn49IhW+bSipa3DZ5HpojCbmLhvLKzC6T+nD87mMAojUIHHEUN6ZK8jcv+7
R4zeeJ0Q5Lml5Fmh+RwoL189ZL8YTIhuiKEXVf8i3KavusuJi9cvsqUVsADNtkYdIoSJKhHFhNEs
aq6Cjq8jrrhwVuBJSdefNeIh0+8ozy2na+IQ7+VllpieY1Egc6WmZqomoTjrcs8Bjs4DYofjLwGA
DPb0HT0l5FI/rQkLHfepuHcd1VF16VD60CdPMVhXzLGIxr8X6E3Qd7W4+V7MVu4eKZILryU7qbnr
vE8Wt4YZHSoIdqOGo8qu0ZvQkzdv3DzlMv4vatOnDDfJHK23HR/ikqE6nEsYIDZLm8t9l9cP0VfO
FNp+DvxVD4vHx+tOPeXYJL/n4YtjNNb0/Js2juln/ZwtIzb9Jc+kZzfV0oDKNc6P5I6PtNtmKApQ
ZPMIPmrcCvErR90RJxosCB/osPL50IxxfJdBxJPrT1MmfoMsm62/LEqoIGgdRLVfx8byv21ZQCht
DxloRbjCHzjxqB3IesWLdLyAqhK2+MTuKjWxvuwT/+x55GPehyioRWKTFpwz2hL9+O/dAqVjZWWQ
0jViDL6o+sgUqOcehJh+MGnUWrmi+S20Od0sk6XGSW1lLaXrs436cnY3ELNEGZd7MHBcpcFTvheE
fHhFQ2HSsdeDYRFmmOWhIfyuPgcn3jjzm+oCYumI5Li3xSFagMo5Gbq+LqVRMXO2Mqxo0RiezBNF
ajnKN6s7k/L4wkMVz3rXCDVPJ/8V1zJOjhlFFPYdeTy8Bkvz04x8gg2hRd0pbd4ACx+BlD4bSpYe
9xYWdagXgwk2f5jQlX2OsGKbv+cqyKyVSUr/5goDFuGU2mnJckWfl5uECf/PY88DvbRUKSTKak8k
81cIMmJrgrDitGFhrYKyafi6oYgHWBNG1bsYjgGSHEekplUKCV1GSDKN6y2cDlXNF78AaOm4fIzz
n7o1ZAvDNeOGdjUhwV91fzfEGviGM1KDrWLKcNZZodlvKPuBDpolWkEssYWDx5Bwx11Dj5n7eZAJ
WvsCvhIw6X+b6RmnixH3JRiNNMHADRw48eAQdnpyuiHFM2v7Sz722SeVlxErMcol2HidATt1S8M4
TExWHOn9r+eJoc7xloSIL8xHcu8vnNxO03KehQI8kNhYmZvxsv0+ri64TRnq9O3lPj7r3NaGWkAl
AvAwsn3MgvIe9tAcPJivMcR3nXpa9KKrcFZBlbPYJ5jg2hdeDgXH2RUPdcEWHDDirPBsmos1RJnf
NeTRVZ+lRnI8FJ94BmE8lKeyhraVdW7FhP/dJA0vV/hQGHkHHjz8YiWbAcKAzLvU7iMF8F3vRisg
lBaPn/cTUaa3EbjPyF14Ok8mVLIpHtYUaYucGMIDclPb17IKAK7Bt2KC/gto/UdTwMpzXGcxiwlC
RgqLGfVyiah7DEg3gTQ0/doyUV2rbHUmtmzHzqI8euN0QY2lSCvnxuW+11Dq9NURArmQHhDaZaqA
w5XKTwnrCF+fwA/2fHpSHKzIRQnYukqhhabHTgLJSmeGa3/LZ9Zfk9bqJa09gGgAWEUmbo+jeaMy
1pvGRTHbkFQYi6WLPgESANyjCZi27E12FfamsATU/h+FvrIJPJEfSqSdIB+YMmsieK+HrJib9wgc
yeVVeLZVhB5acjdxKwMJEWieVMUhGiM6vVicuufgHNY0NdwSJthf3rf/loKR2vgAf0KvV1RDxaWT
ajVdW0kj85ZsiSy1PgiINgfkgS5H84Ze5g0r05KQwjl6gnxT4nMYLhSXPEy/JuPGU4bQ5j1A5mrI
gj+PtxwqDHgrPoN6tYE4Q5DbU6UWNr/0y1WuNcdusNu21Z/QTl4ETzJZVTXmTJu3ViFe2ENNB8IO
GIXBpU+q/v02hbk4KdlVYgUzA45ZLRvnH3ofunwuXVyH16JZosHhD8uXDkCo+/RuNujZrO74jX+H
hqOD3KiK08FJOrytUF8mo5NXUuJdQags42Yu9YNtN+ni0VNuokKofpjDkWixgwzPtJrzBevjWedG
PHXoghl4XAK7o0WY+xH/RSJ6OYnutDO9XN8c901lBsLlzbYmEqPVpeuigOKe29zFRUSWr6roIN8A
YE42ijeV4hrfHY6r1IskAhcOBKra1cmsB++Fd0QFvsF2AiNnCccN1qgDxzBgIJiDOiVqDGP4kp2s
kmm+zVOWCwbO/rbQMUJZtAznsmK3o31+EB68HjA22vzBiCR0X7TJtCh5EBP2iAz9EXLS2tA5ji38
xCzSIHqm+xuYdavR8MzQtN4kTpstQ8DtaORPHWMG++VqNcQTTwbU6C7dHSaHMUtQqf3Dj2cZoGrZ
a746NdZ8ZZ2MhhIuY8CAPuvpghzuez2/wj9f73ydJsVXuQ7BRRx4i2eFor2zDq1AMaf8xTz9a3kT
5xCqQoBNfeVZCRydnE3Wn++eCzxHfLOQNPFtAPNk7UOSDwR0Zcp5h2eUqvkqwnXApFKPvSFafUyq
4NJAyCWC7QuzLcO+PcOzjUoHdgSzqFcDtZW/85iZNneXrL3xqPGqQ/vL5qXSnFrfV0YlJh+fPCfz
SbYR9jtO8KV14YnrBx+ZfxjeLETjMymVQpaHL4WPWagZ2jLTh2JavISNPu9PhOEZ/yN5QM5PbraB
30Yx6B1r2JZlhVsIzfX/GlhzdNaXqHXUY9Px3nW++ROnXzEwixToZl1nxvTAw8xjWb4erw2OS4AK
LWJt+jZ1nQRqvv6jf4wWjIr+BTbsjMVDCYdMAH6iIn0iaxdXgDsCuUdvxziJ8qzOtx7xnq+ivFnv
f0yeSFhrDLNffXts8JRWjQGUCbCOuidl1KmTqQ/kMJBazvnmjAK7M2vNK1pJpLK9iFm47WZgDpQX
WgCAhY7m8fRLZ3De0mvHKvQmqZspkQvxx9VW3mLoUc5ZnO5XRvB58yLrlAP2gP7bCgCIopo1P7jK
5WD/56VwkqsVl7OYzt7MtZ/0iXlU8Gmg9IyJbHzgJte+i8I7laOGgfxtokGrT374Y0UExM1vO8n2
jiD4YItQ3HXzOj2jYANpsLtVIkI/FYnD5MGUMJu/ulzoSERCLSozMz2C8ZIr5zVff6CzUH879i87
Dl6/SUgJH5Nwj6yGSlGBWjZ7vRim/LFstwfZtaqq2J6weDSewjU2O3zyHZEF0ETofCwM3YA9Xuag
jCTtZ4jAcpowOXzJkastb85dC3g+HuW8xbd9P2MhaKtbGo+MxTtTNlZdedmYrEeAeAqJKEbazV+a
Z5jpFUomG2snl8MxVrVUj89e/ik3BqOkHLmHNHwTE9dTNiqndTI6Q5eI4krGqENBD5XlOI8ddCJh
zh4QZcJoUdegslFmHR4INbK9hnMngNouVO1AHYIVVrftYlERTCIsCQIk1TfSh7B73QhGCfTaf+o8
qYIy+619k3/mLqi/ODTzEQ1Yf7cPTWNPlK7y3sotXPslBcXfa6PG9Q6PS+LhqWXZjOrgZXaKN2r8
QodeT9mFD0RmBWkGNh9mL1s81WMqJp9VO89jtktALH5AtBovHM0QYTPhP3CRbdMwfeMdtJlcd4En
3vcvU+O++UdCWr7MvxI8qFwFV+GM6bBhX2ccMTihhX/7fcQJVSj5fZgksiGcPoTh2kL5G22mgkyi
GUgxtDC4Tk0iWyKx7og7uf/6cSfjAZGtEEmYXEvLIjEQHM4OLxbXnUtp5K2uxkoKlqkv1KlSGgZJ
bPYxxBsHDuepPZ+ig+gfUa6zPdCl9w4xCWtkrgWou/fNtV//XLThTnB0MH2IEcQRuapx+H8NrUEG
5ohzpZr0OfPrw7UwppntVWbWN2IeVJS/2kJKPzFPHgvrGTfxS5weQyniolIDreYi9LD1pKQLNxPW
Me4wyv/iMIN3OXSLxm07bkfEENdhMIDknLNFzI/IcJ7Q4AVbIhcAWgeBad0JGCtm2HO2ArPDw07W
5w+bC7Q/rVwOobokZoLNoT063U/XvdzrF7RguiXNo4RsicN507i13wrURliunlgVCWsBYYSAYzd2
Td3uCIyiedMNUXcEUD+PCNZJzmgRlebxr8ZgCT9NjiO1db0bLNAYkswNVxkjW5IFMGCC5VULSCsR
+g+cz+uCA0nFkS/0VsCh5XKbQXwCVrAUtUKqn2Sux6k1lQj3T0z44xlLIY26tzG6VuJrwIpK8Z+s
/rgqs7M4/wV9gx6anekNZm7HBWlTG+aAZ+rA5p59JB09X4pjamxEWSlQFmkOVSTo4Fx9YuXgJ1Po
uybCrxL4Nz29M4QdRTkMLOFob7wSW7edB4PtBLbtR36M6/tujnQe3YZCHqO4WutFw4DUGxJB8RmC
uazAGSg0OXtLLuyFAY4JqCihv2uBHf7/tB9VeA/voG+Nk5b8Jnm8iwD3qpHeLZW5VUhEIdEbvzlB
1iNvjKQw1yeqTT6zg2QkbICxJj1jHsV3YO+SSq6OXq+L1ASyzEfSNmbT50ZZXmVqnD7a9BwZ9YsD
ZK1KfbCqKWW3+l5XxiZliOMIw8czLqlyHRyBh013z7rfuASiuvPhBeA5iMA3ingHo4wmafqPBp4b
4lYuTlMjhsmpNBC2mk5nWLfTfka9XZdYaKgU6iMP5Vs42Ks/5GYbdJ2GJh4fhHbDRYY/6x80kyLl
kGtEA8t8nZheDtokuOpk79wAlGUfeQYXJhwyuHINn/Qfj7DjwUa4UwQOBnovvR/NCj5R+hBRd1JW
lAGv9vHXArFbDifETnQGTui5f2xc7vxE/jBnYXjs8pijK38xcUiDn772ZFCAmOLw9cxejdK3oDA2
Po8yh60dhBsP1gd1c+sq3rmbtfoGisqd32tSegHVymXNWkct9ku5ntHY8vaX5QFpiiP4l0tostpr
tZZWReJDJ9mPz5NCSH84dxmpPTGicayRaYXpMGXZzLOc6tvi0HhSNhAr3M5Z68f6WBaAYtUX9svT
kBXH0Y4CZZXdOcxHZiTJm0eU7FO//FgV2NNTNMteGkBSDUVkxnS4FoX3MKSOizMtZ9B1XNC2yt/X
252Hbqkepo5afMjUU7izE77AV1YPuO43S8KOeMKQFMuCbgYCaqENXlD4hn8/PicqkPgrQQhxxIff
uU2UuVIQW99F3mvVu/aHDBbUDgaQgKrPNprF5OdlQXeIB1fivtiMv9UsdewF8ZYR7aTR7fY+A1xL
ddGVN5PlB58TN4cP/qajXP1eDApHRQouQNqWjMKOYy9XXTDsIs4oc+hTqdhXErmsqZnQK2hmQXCH
w0fhYuVUTJyjriGYqaB78dl5nA8SiByO/UN8vGY5M5kVT5mp6QBdDJwEWRPfTKAzBnfy840onFuu
Cji/YpWAulA69PAjypbEP4zimB09gHJfHMt4Hjb1zE6G+J/AuOzXUAkPDV2i5JfmZ+h0ZUwn73Z8
PM+BXRn1v427oAZJ729bW/dNfeT0ZaoY11U3HCDteLMK4LOk4RPzI0z1PLZIG4sY/e3Q3RMB7dF2
eI80xegCtbtzm27uV5lchNsyRfPZOp09WfeCqDNvCfACrgovFnHEQyFHNrIScPCzsOUbo8yjldre
Chvnw/8cUAEYI03pZvSFXCG+QJcwpjIgaj8cuadWa4xODpKeK6zCfRJNnPH2lganZ0w49sD4zuVD
rZcOD5226DWUW2nW8Jxovs359ixChsaVF/JogsHGD2ziWNqOzEItujM14ZIk/DYNkV3plzIeydfq
IXYbRJkVoca8JC5Qgpn35PW+kh4VJ+o52jl0erh6BF+Z9Df7BVXWrkj4VGFmhozxjQK+wFRcFjsi
1pC5A5Xif6wz6ujY/zq1spI/I0kuugceYMpFEvIVt3Re2GF/92ay1ZrDQmmx2gZNvafqRtsTl/Js
2FYsi4k48yKfQskpQPjhkHLOPccxa9NSPTLjlIzeXBXFLpOyK0Yjwqz/eE08GASa4ZhT7eQR24YG
qmqxoLnTuB79kHeW/MZvswhDjMyN50mXsvb3b8aG49vfZomkPd5WiABMfrGswtxaHlrmXe+ZGZ7K
8lbL/XwYr7YmrvzZzmkaRYvjjt/+gLAZb34/xfR4ux6XKdjdam+vPHbkAelo1SSGECFv4PLmC3Nu
ecM7izGUYqb5KIYbGXWqP+aeZKJiImtBgT2pSa653L+13WIPlX1bskKYhQku0yDwBnxAOtP3pUrH
Jyft9NVt7xAsUbTodhmLtKQgHM7VOHyAt/iq9h/7d4S/LHoQtRKYn677Dc1YAsQNw299opbJe2jY
y5vQW6zqhDp7Cc5lYaqouIGSknNicSDhZlJMO0yaPgvp6seOenLw9bmUYCEc/puFuR8Kx9WDqSbg
ETWqeHDcjRyUA+4w+pLX9Em1nOEAoF0W6Lz2CR4n9UX8uo2+SLWi8KF3UxH0GS5ROgy3yb/hmoBR
W4nombDmzxKS6xILwGO6IeGoIUHju/u144ON3LZvexWyLSWMUnlRSeByo2i0y2vTffFBNgFFXM8k
nwYZQwbGkq6spnps24wPPz9sGw9EfSONdQwXtfxxVFYoUDHvyIQUWFCcLM/CKC4Cbb0OI81+i0Eg
Qw+dsG3BVIgypRQ+nAOl+sxbfLm94yrnv2ilMMSozM9tDPhPLT5oF+MxqHyMozpT8fGZ+ed+5L2g
5S2P74RDdYzBgNlfIfN3HDvSAt8kF/a2GRjYeKR3sodRVN9AzUma5lk3z1jNu+yIHj4/iUT4po1t
smUnR+lbJDL+Id7C0da1xdapG5WdOOcLvOn10Prqpf2WpYeFR+Zkc19yCCeuGY4IsvdUiZUBtOv+
YK8IAUSP/3F9KAx3a+HQhJEWSg+9bi2g7tqBa6TpcB8TU6mLTfQKCu96Lb2u/ZG8zrLyy/tMjq4u
TyOOyWKl02KVMSnprEBip9eff0f4gZ4P/Ilm7jkYUiRnryNiWOdWHgY/1cx6dae679B7oKubsTFn
NQnZr1OIQuYUdgKE01O9MCtyPZGqc3zLbRPSF3rjnJd6e03HO5f/bM+4b2oR9jzVXC0FmgucPO0l
tfaNa09wUdPBdDfiK//nJCLmH5mZj5KFiAkpbKhmzaOifjwVWVhWf6J3PjM1TNW/LyTb13uMpz3S
fRL9TMTpbDdLmyKgw0mgOZPuUZIUSQdjPl2HyM8GGSa1F4EExvWRvPKtiaN1aPmmX8drUrrN7eI6
0rEvyuCMiVPk8d09Sg/uA0RHKfnTOkzu3gH7KdG4zoZF2CTtAspP+10C+IgiNsvQaxgJBzN47rsn
dRsQltolJbGlwJoTyeUuoJlj9yHRTndDGRCyAFpcuiyQh5PPvzKfrWwkO/vqkKsY3Pn02U8L1rED
id70iFfUhkyy6PWIlX7VhqkcL3koEuXubDNOzINtLT645OvOFzXG0TRoUAZYUVqKYA6o2uDOAJjp
gLa6RzxdrcYLn4Kn3ZGvr95J1wkLwEgg5x2+RVXFR2ZiOVBWTqDEGmMEpRjgX9OF3mfRqXtc++0v
I9p9D16Gv74g51gnIgcISfHHHKTJ645hZUbyiuFl/kbaKKN7cCJlnOlAzrLpIkkTA168oFTSlQDI
BrS994KxUeqmBuVime/GagHgo5LgeU1SNCeTjXmE2t+oMOuKqArgjt6RJi/ndJoP49wbcGB2oSlm
e8LMCVnGWUx/rcOOhq6wnVuyNUxO8wLqBFzjiNKP0zurZ2EC+41Q/kk1/5D1GkgOcBpY3ops7hdq
LwrkYwiMtmyIDjIPKlGdvvi2o6T/a1POlWWhfzeB0P1vW6YHy0X74EA3GUMEVlh3LIRtFcRt6159
6i3KV5+hsI3psxImYqmdvoxOOc8FKOPPMkhzDZQg6xrZHSjy9ovnOfS218dLOEyj5XNox//CZYd7
KFZjvnYsQsIX2Nh3qRtZ5C9C6l+7mrQ1KbbkP9Mzkj7gGxW6F/uupzorp5JXRWs+a9lu2kqvGLQ/
kJU+DQEf6FC6k/LTDSSGN+NlMsEq8e160huzhwnOBlXeL9oyrIYxmneUVXTDj5up1wPl+rE/2xYz
MkzgbLSfyiMqIV7ZjOCe5rR9f+n0aJUTYa1AD23P5emsufh8QaxEIaRKrxhwSSL/cL4tdvP18nsz
0WKDQG3V1+2S9dxJelQ9+kXtro7N8sxl0h+GIoEdrmhvCEVbucHffGe+ZciPVb7gnAfdhfffPu9s
kaRe6LL84qrUxRmWk6YR8fcdWk5kYYyT0Nb3UT0cQ0+6fOIgcv+0h0K8iuCheBZgT8IdZfrSfPMZ
a+92lXBowk5gmnj0kCRmw9uGYR7bRbwrjtECkHTqjvEGcpUUw2FRLP2BPzD/ywuyOaF70ssvhRMt
Xmzw9s6mWePLJz6kLrhpWvBT7OuQCpXDwpXYPpXyWemRMBlz4h0qYuXp0bb5FDvYUnO1+gHSrlTW
ARK66DZNaHk3wfqwz68omKHoDhVbCTf7ZvSWVI4y/Bua8977tmMtS4iQuc2Yww4VfeFksbXBImTx
DK4vIAqPaKYKEAS2F7kmGXGW8jCnKN7EhnkrBMDooJT1eCi/IlkOmucksBZzRh+s0gbXtQzS/sdu
tQ0SHL4LBc+BoWWduhtG+D0HCj5eSHBXBXE9vkgvbcPfDUQd28eAO5FOsbAE6mh3Up2zLV246NvT
YNInfp0cBz1FxQXzn5e5o2nDEdcuSOrPh1miM5g8A7DooE5i8vyaddOc10JnoTILrxV8Ts8/93vP
YmhPtjwmaBypVJQMMU5yjmMh5lZNDZuKNy934hIxXXd1V5/f/BeladMDLKB/+mjhkmINpQgoRTzV
qTCQb/0C8dy2yFCGicBf1HLB90j/A+J6tJV1twm26XnZrDT5jSCNKrB1l2EPaFjrdgVWXXAwEESv
bRCIvRVOnfvSF2inqv/cJpVXaRbjbBeTGyI8Z+yHj1kA1itIvtkoaibbNok8IJnN2Ry8RawiLQrb
MkqnTqGZHjaQdtEeAYU+HPKoYgRk3KAJHdhsjvL/ogT4r6CbpzLhoh7W8tOjVGOVMTTHRAm75MZV
yS5XEc9X5n9TWYaV/tWemTo5Q7p6p2fv2ez4tATWVRNME+appQXfiNIzNpTiuytWN1qvl1I1AgbN
LfMpAXFiAOgKG+JJZbLL5wOX1o1h8hOLCt+z+mnXxe0uJmxU0dO8Sp+wll4IEDEGdBBrocMiXzOT
lnWQwFfN0RT4czjNo94WxKK8CgkdCL++2bMEOdJfh/iwf2XVfM9maruhbESjligHZ0Z8AhijDh7V
fat57q/xQRgt71sThjGbYjSky/3gkdM3zf2z3574/qGcGFuMPZegWnWtVm8RI1RVyzhKkSEVS7pB
2ANSVnJeCQ/2pyghku/unn/w2rEDJhafrJLw3YddbGS9uoTh4HoIuwZhtTT6G/+rSS7XwsFBZVQC
9upP4bLw1NxUgSIPKripduZuEIkBmpN9GijJL+HuUU5HFxXUsF2O2hGBzO+IGykqs4QijhDmXW98
HFGEdXoUnZAN30thn90hoS5H02HvoS4Dbt/8d9DPyh7QN/wnKMBKxpatDfdxf9ydJM7LNnYyW2kO
AF+3AdknPO5ZgQX00oWlmpgDH0kWHqVu8P9DIsXEYdcRbzQNcnjayCmL3MX8u8QmYtLv7te0KKkw
I+vFH/NouzQ94r95fz1w91+JiPeKze3WBEsIBpdQxdGYPEOcym3O+xiYsunsyIolqtBVsn6mo9pr
tiX/6CL1db8cSjugwlTl18ofeBM1mcvm6kqDXOruJJ6o+vga4jDtKADG5JaR1+5RXGOHcIXhNGTe
zf4T+BZSqjdf6ajKBfcGb8cq/fei9FDKBJTtv0S46uWTdEsVKqSOCDwjyq9oIaZoYGhKnzdW/z7k
4JKFroDgvIMkgZLTulcAhI9KMAhy/hMD5jPftHXFIzZFB4daE4hw7T+ShoPKq98UZCkjW+vIpaHU
zjw49uJdXIZE+D+6t7BtCBDseCp7bs0UOOXHkFzE8j+DmMXPT04myLuPoV0tPAMi2BXxHv3qOV+d
KfUeYUAG4PifKI+165jq2r7LfXpBJBucNw3b3TF6CActAEoTuSEyRmv8p6SK+ju/xU89p/aE2Mli
ERZbGga4ahxYlaREPARIhL9PbIr4jpmmuwWLoxkkgbqLGvh/LabfaF3TTr6iS791U7uHXETHuOe/
6PNdldQOp+Ph5TBcI2evdhJIWH2jc+KT1OrbqFyAmgGzv83+QGsYEzYk6UD1PLwQYJ5M8KdMom9K
Cz63+kCoBf2b0Xi9e77n3z9OU2DAZuAm0sZ4k0XQhP969PyFct70OngD4ve/PaNVHZb75czexfxx
Rn7MrDKSZ9b7Gxg5A+ba7X6ib0+xtoN1pnLffKWD0MEf/2rZWyE8dKStAr0jNFtXrcEbiI5iRyMc
H9ycxuTNeaafMo0GiTN9bctz+AjL1TEMnVwaXGfKd0qRCqfRk0RZmkOTKMxg1ewdfe97mqbK/zzz
0aPheFeAA3X9Kz4d90GoxlbJwbP8xUGtLn3YofrogCFd42Xfz7wimEKTGVQZPvlSfgaAyvp+bAoF
XBgtJYU+diSnBG7NjnPayKiDGVFysTz+ZpR7+u1Oq8Gj2VJ1eir5Ophi0WAbOE/5w+PKRCOLKXgv
dh04lXPXkcoEMR85VATGDVF/Kp/D0GoEJcOfgYecV8COOP8rDO/qQJCfUOmt3WBaxfEhzffdSeVR
qmxX+bAg14Z0fFMmE24IFxCx6iE5gQVjGkEVgo9xz4C1Xdb2K85ulz9GkOIDeqvP0RxGuBa10URl
JVvAersut7qmNfEXxWEwZO3sK/xePwyKCzO2oKqrZguyo4X1MzXDcHHVBJKNSlOZhXQ6hvwDTw0A
AkxEqSh/zOuTSXY2S0FrNoP2M7RtTpkOUbwXJ9C8UsU4gjudJpJuZZr20OS8xDYaxrSW6Xxn1Hps
tnuRzB33emGoxkh4ZYvp63Keq/YUirjPzXJ46Zhz5/P4VQqy2pv7aco1CLwUcYyJYSUuTniLEQqh
U5TJjey9kxaXbJVH7plkbXDNffLMvU/s2tJRc3DSMfPovdsaqytD68l95V+N4NzgF08I6tf16UZE
4EC8MQQSbXJcgTISjs3FH9IsPRq79PJ8yquBzc4cmikIonJYfI58qtUtf32D521F9U1Pe/T+uvbe
nacg+hrmbSVEOL60z9c0EbK0RXClh2luIv0lN4S4rpiibdGiWhRV3ooJ0ireVinADMGIB3ryh9bo
5QhNP6tIre+0nW3Li9k4xwCfabpPK+9TDZKOBOIrCtV0DAHGRWuhbtw8HbwJ8MJKlBL+loNYJ7lN
zantsIV0YReWrHdo5h0gx/fZWc68xfaw5teQ7nHo0GgxKVAGjy4F+hLrWdywg0GMNw2ZxX/M33u2
71ilW6X2UKlHlalelSEgwVn4oufcv8u5TGlIxb6qeD6um17fQu8AIqY2FcrvkjgBAtsspQtAnZ6R
9qbs/kak1xogDPND/Ow4Pymxyzl4El/jYYji8t4wE9mB+fejQXpKGoMKcRxPHNwjz5grAZpxpjD2
E9FtEH1fBS3asQ0RUT9vZHBc9Xz6CBLaoJsGkA80jpythWDoXHUH6fLAQ84UaOal7MWVMqQMIhY6
FHHclntciOnK1P51FrTiypnT5wd3PBvJCCLadQEgjPv2/jELWRlPJ3kYwrnt55F0+X16pXaxCCfs
CL3h2BnxhcGzQxgIx8qtivftJhyz0SDWGc/cLTmVHuJQHfzoraBGU/7rRGRXOLZBP0E6GhJWr0zp
oZbVltJUdN2FFdU2A7AuydesF0ZY0IpH5m1MOrs5A4C2ZlISHlrjYbzCHp15V4yzog7n0PU5ct1S
e4k4r3yTlrd6ONh5ZiO+d1VV60JYC9c8PEUDFnDCi/Sdyyu8w7lrVgLAaecSeqRdsMxPTC9Q2JS7
hpKas+f4Ays9riKrQFZn6AtU6NGnwv1YemKWwpKQy9UV+dxICLISLGFqygi4adybJSvnHEqKuGTr
MzAytt5QFGaDpsI3KTPjO77GoMGDVIEurLByA/q8qtIgKDW00W/gIJVN78Ec5jLpAZdgHcZ1xH+9
HxVXDAVipm5xaGCFDgJePmZVmCpKzlsmPxtJgXAxkDFgI7zRew73pzj21UTfzrfYFSFZD6+E2qY7
wzwbzafNDy1k2yxxHe1AWsOE1xCYEHzGn4im/dSqpe2Gpbjf04qY+4Ax39vyCK/OhV9amr8Y6ISt
NZpsMIf5wSZDqcKzLxbfjJjzeRlm4TiTA2qRuQuFbbwN9Embu6BwI9WMg4cAodXLp8v/0uAaVRdP
av2JlStsWSugCO1znWraGFD+CYo5+iml7WCyhouq6AeRAf25ZB79Tm7dYJppZRPNJd8Zb7UQpoIa
i+HK1PI2TZogyxATuGB1O1c8Jyy22qgnNhMLW1JBkabYGIoTcoND6Vf7mjGsvJ2U6H7GEQvDrZET
wuCR51AhaaJndrteWDYrBao9cOhZyfpTll4olr30+bFrrVbeNkiMG/iMSNU/r0SoEYPE9yk1Bn7A
CO4VGtA1RKIV4k/ARaDBXRtFybFwbsyhYkOdni4V8VjdA9l+85FU+rMLHa4+3W+Y3CdlGRK48/Vo
NNELCS8QCXHp7/l5gEMfK8oWcUA8YNVUMe4bI6L039I7bBidXEAm486i/pX5LhUWv8dfgJLkRnqQ
X5/Dv/XRvanYEXUJRhXUDzaxkd15nDlsFn4pWeDACNxYvGF08ZABoDeP3ugOfHV2X4ACHh7+pGBf
50jlgW75gK6C6vTcUJpSPUSCVyQA2BUgMyrFJ/njF115TEgQspmp4SHFZBAYFxVUxHlZFvOrk62i
9RM5WXm9W2GQrRH5/evAD7ar5BF85/Urz2BQfeeKyLOXxg/D44sQr46bWeS4zKD6r3Y8MAanwrwG
U+WYjlKFezeWbs7j2bU8Rf6q/wiudAAP4lxaCtIjRKMOZ8ioD00F7fZmpDVUkA8AR11DzKUNGXMh
D4L4D0swZ2GemzZ7k4Nr4BY5XOA7p2hqCVzRlIOMogIo9XFbxNrk1p1y55xH747g5xgLnBUo1qUB
5rwHk6eJAQ7QmZfgsXEXh00yPLab/CqfYak47vLUWgW/G5hYLWZ5zFKhvduDgoLZXBofUr7/bHN/
P1Iz9kpSarUqcYLttyOuTgNuJHV8X0DDqHPO4LrQh0whv5vs1orfVJ0MWnR6Gnk4i/Lj5Ebd4Wm3
30zX77H5AXtbhQi53CJ6KIPFonxjcIz7Nl3IWjl2tsJb9+l9MmtaODTO97TFUZA09Bhlex5XRtCv
TodDi5Bduwy6TaVl1f38y1sWVeIIoTigPyeRHCw7WrgFEq112ANEg6AEevOHAgaNcGftXi63VHrp
RdJjJoETiDXdrAQSY8J1JNgUp2XjqBQvNguv4Q35UdDhZ2i084MUzfXunbMZDpmHIzKPt34qoiLS
6DrQegzjeLRnlKfLasgbyDMP6qsms6J7r3MVEw73WEWumPLQdpGKfLAK41iTSDoRNhSe84GNy9FH
lySKPqYqHTfpXjBuM0+EkjNe/VoL4iMIfvf0vzkZ12HUJEKFUODsQm/GOksyyjhyA/bjz5ccfnwc
KaUr2jrapL1bMLa0G/XMqveDdM4dIWUsIVC2eDKV/r0WZyGCUb6WkRVlsCQCZtBzdK57/te2stNO
5AjhScKPlP8r1B4RQaapOI1TSQAxbifW6xS9iax6JsQ6+9ta1Dc03lhwOu4UB+SMI+LV70WnIfgH
dy5X7cleS+VmK09UhcHQF91FmAdkU7GlkJ8zLSOeBtVV5f6xtlcupH2zq+1lraHIl9+8IFq1q17W
8IGmTcUY7APzJ99dDbTnXF4XzzvEzoW3ydUDY9f6Jd2iifOtDyQKrxE1LI+8Yt+luP6cWTmQnqmL
jqQl3nS7+uQ/XyaCnx53axkkB5uhUkyDjOf6u7cPe+yPq7rfrrJOK6lPFvymxOrfiMBxIrho0VP4
VgeoSc913Ot6h5iiQ0iz5r1DtRQAZish0Yq9DfWk4PGEy5zvIreee7OHqQTbK5mOyY6wjhRDnhST
l1HYC6tKgPqLZga0pgCXdfhQApKjDr7D+YFj6j+s41ZCmnxMmseU85Ff9Znh8ai4JVidUq7d+hOb
RRAUs/jvgPXe/21h5eDuJRU0zJ+Xtpa+vnrzDSbLTjjapxkkZFarQjRkM7sRvGU/KkXYyM465NXi
vXBKde0cPWstK3b7cpr8mXjBWGa4xxJr6vKTQAKDPIyWf6EszYdGxBfY7x2o8Q8+Xb1C+4b5UcJ6
kQkk25XrMAJEIqcXWpqWroWefUPswucS5EnhzTZYhg9ZHpq5FzhiTHlX11adGobJWc80cAx0H2UA
+d3LGFCtLr4P9dfNkiQc/lJ/VZue3IIx5k3RnCNLqqLFR4fdCo7xhqgAX7nxRzaof88MNYn3ewD5
CJ3YZpExoOx9KR6UrmkktbTklokc9jm/4jo1Oj+gRJWX4bwLE3zRpY0bkM+66Llh6i5VSnHrvtpU
KxZRWDpk8Blwr+B75li2g0TcrKnlivihZsdDv1aD6s/mQV0EkRIFkw/HG6oeh4OZ6Q/RpUeyNR2j
1RoTjZwOxgosV9KbS86bpWKdFbSaMDouozkCV3tV153M6SEbjrWEEmPeWMLQKzdy5xfd3NzGcLpC
Qxhr7Y4I5MUYJcB18CV2Gi3zRpx9xBVcTsRkKzPsKT0zRZx64CiKbUbhTSMqg5gnrWpgfE4yadB0
ZTQxqQKgIfaTw2N3MVe47wGeTiDy7JFA9jbbV72nZUBhy6DXMu1ATr4FErab5lMWqiQrOiCHF8MO
1aIAJ1sMNeug0GowiXhUf90ujORiZWGna4HFXtWNltt0eVyNtP3I/+R77ehR9V+14RAixBD7cXjb
SVHvg98C+/6ZFtS88ArT4klx/54ztvWdSC95OZfCxFawpMNvB1bXzL/kDkF5QL5wSwKwdxO2ZTzw
U/gBMivNwnM6ESyblOfomhF6kVzacxDZsKX9aDmGOWxTvGoz+1DpCg7F7nIDe3sHjI7aj3HOWcIt
t0xZO6FwJnLTB1bJFvu85vsV3eiBst/jExLGM/IaDdAiBpTd5G/ySwWA7fw1lQKgWlnP2bvxQEsE
8ClCOBVcp+KKaibrmJ0Jua1MWu6lFlVenEx8VBnKfjsU6tdPSscrU6Ub9MVj5NNQJLfYGQFXQvWM
/WKSHsZXLUTZIsFPuHFS4XXZ7SlnjG/kesunWQBLCy/QJwPBHOOaYm4ItFRDslIdCAaJOw6cYGGh
zDOm2tuC12ddFYZ3c6dX0eroLC0ydRIPPJpPxyrOA5HsIKVmRW2Xm8NI0wlAJcIsl2PsjAUVAB7l
Bph5ub5A0dRDmH8IhlfhJrWwHgQW07TNejJI4hG4DheUk9RY0fJmRSVsvNx/LSnBtrWK0phsz+kS
QSkWMXYoHgHC2BBbPmGRhRd2ogHEJ3OL6a3KR7UACAp4TKcWve4LNYpDehasnv1tblEtsEe+qEzk
Yqfngmuo/DRTWcYzJdrTuXKiZA7K15VuQ0VZtF2NiSUS7b8FVdTdOFc0B+OnhgcoJ7exIpBiG0yP
BAt9PEjFQvoXOoyYhPzjBqWPtiupjhzYNmeDqbL0xk4+w0QtcoE64gnTb1A9ZQYIYxPFSYND2vZ5
8tMmX6snVvHbFK2xaO7WNc5bWnQdcvAvfumUlQtSh6Ikx8bc0OPhPHmCydWjWSbfMKogQcsud/gZ
nim/biLUZwdQyJ0kSXj842ZNaXiPbeSNiDXauJXcNG358vTmTDApURpPHS+vcWiQZwAzrP1IlC5C
DjJxfddkWcPXCZvjGWTvWGQSkwRgWeJDgSE3Pth6wyYlQ1GnkEr7H/q2BqOCYRhwZ6WzFNpAaB/f
bkjEoA1JUOfIAOV8tQSuRLtkoI4NFVSRut+Lv4XAgFCrhT+/kC4w+Qfi5EuQZupqFkoCeuEgvEnX
zRr2L7TIUShuKvr0Jlgs6uLcVVC46Mkh+gdd8dKeToVt3O2mB5TpNoIvaQX1MeN4zx9CeU3q7mfM
MTYCkWb6NP/yUYjVXr0Zz/yyN/dqV07psIauaNWSanotEjF9xWCVN+dWu6HC2QBg6A1UyhmmvNkd
+3ZeudmjJRNzJl6pkvfDD/28IVo7a7UgRQPtn7EnAtd3/UlKx/NjVOfoylg9SQkXeQjcgDEb5Ha+
55ZvlT/pl7Mxv0ADmkO39dWyBS/7og0oPecaukxJLDkhDrJYcFpCkEjkCMuu/nBqdyDpBsF1rDze
RYvjSd99WH1LL2mJ0Q9iU6LPemdPgybvs0VQB33bb2IVU+S78JrKXa6dYPgvFumxb03rMU/ba+1C
PYmUhUDhzL2P63ziDJuHcBPz9PK+MJB7xBkYcRfdjtv9REFu5KrztqDX6N/KDoXfeDEAaF5yjs81
4kqpdbBQ3YUDb67QunryGWyTpP4+p8EFBN0Lpo4FgJf8OHehvt4fosz3tsCRlIceg6phTGDbHv02
nGQ4lQ+ZlGn4cpOlrQdwNyGSszWtt9Rcc8nffJYoy76oJj7ORe03w5lnNyCciIUgESX8JZ9I1mS/
SvG148YGxMBw2o+Y70Yy48zFX67lZJovBdz9PrG3yBGAv9LG9ZExjmLhSLuzBRNsFiJEm/KU4R9t
ieSC3xrqWw0wp+bZm3omRHaRO5ryZmcE+YPxa68K7Wypdx1nCjj2dxtE+Cr3USrGOtKc1mW4M6e0
oKwUwDwF5Nacl0kbGYBAQX4CVnXOUfhI1gnNvoWXFmQ8Hh05Ehj6nZ+a7mzMLQIgo1sgMeHZeETj
NRTUaxUM0MIbbt9c2xFgWhjPqxAQpR0QHcXGF1joSBUi8+3N3ZpR2CbpgW6YlhxhhsJYxJP/Iy5A
YQ6I6R980ApqJN0OPkHnNL0lcxOqYMwbgpXidEC5qU/VeWxTsXMic7Dqn64E42/Wyf2Hef3GgrAq
/olyFcIsxzMLRxb3aNg9loNAv8JsGyarq4DPLkttUEbsqkTKpd2HjFEEsrrUk0FmOrvsKGZvUbLc
A3b0X+11Wu59f6K8G01UrHbgEQto722Lni3L5tDJGL0I1cN2EPI7BkH2BgBffJeCa70OJ+3BSD51
Nrqgq0HkjxATtgkYI5IEuKMui2tmMOH6H5YodiF39T3ueb0WRpIRabaEwuUu2h04Hw8XA8xUGKLI
BDAX88UX+gXkN7hhltWNXXwi0SKrdqkQjA3mht4fqtWevtVRSwUUTsBEzuuTa1adNnK5x0K2kJ+O
3zRkq7St3PDGUIgG2zrGtTnU0VKio5BnHG9bzZke8RdKuy8KLU17Cpz5zjUJmSJDGCYwjf+h0HW2
ohdSef18XndAtGEgnJg9PHehkuRZeyeTMeIXQXfn7rdAOGAXB4VPWEX0ZdB7WRN+bxY14ISyCZrW
gC6b35+9sOjAGLAX5V6k3zgt8I6v5Y56w2CjlEVU/+fmljMa2dy31KcOZde4pkiTECYZX2Pb/axd
RpH6Wn/rnSLA8vL3AJkeiEfC4gEa4UYz2xaj3mk+axCJhkvKXI2FfJrGeR6BHYiybSZwJS0QmxeH
Czq3mvTmLzvdndWFoxIoXdApGiNcDRjL3vrSJbopnmwxjSCir1C4PLDp0CM/aSZTVvYxihIjPjlc
Va3ryMzg8av3i8pBKXK7qRHOhuHwTzD89iPpVGNdUp400q/vJOtvIyn9z1Z3WTknrmLatxcQxVqh
Q2xrsCNUK0eyFvVvFqKwLEnGW6HdnDkXERmTN0IXcfhMHeh8KrRbRmMYV7fhrAEHM+YqDRIW+fC3
BzgrV/rSOr2CED6H9H0BgnYPGOgceTp/3Z4ds8ZMwma66B4p9lPcx1ICuwXaXPYTHaqZYLdy+Q08
LXTt3N77nl0CWF2NjZFa7jmPBp08OCYJlHjNZHAC/GE0q5PtxzfY0rAoU2Kk4oLINY2F2naMVgbl
8OKkq/ZTujhzye91bEZLvymrMdMvDQUeAdDr20nAFusF9Y+yAKd6cNISycm0mqVCQGb84GA+1b52
+QTIaFFARTSXLztIjxkLmOuaPzenTCVxRW05eiM1JEAdOsqzwHarivsHFa/yrugtZF836APeYSiS
4j+Fxw7f1Zzc9I3+xr8vx2JvZfhbQkN0jd6y3brOo+oO8oxr9VODyKYzfoFSU8+M9ygPeV00+IfQ
Ta25HvcveqJNofwBa6IS1gaU6XMt1jaXxiz6R7Ht/LKJZdzl+biIUR2eYDrR3jZOp0GIaPIL4S9M
6SqWeV+Qc9M7t7w/l6IYnEMLp+935rCbI2INJ+lIyd8miRKG2ujMWFGhgLHIj8sFABugpVS94iOl
y0PqsUXZsgdSp+y89NhQ3Lpmc4XjJ4IXnEXwXJDN1ZN1UIqcDhsi8ekmAlc/tOPLdxygJe9yEksO
Y9d8dO8Zn4eL0Rkld1TKJXvSVUERgzxOguLwhrGPJpz5qmHQtUZnP82txQYY+HSfDdDx7h3b3igE
vJESKvQWlrAWvxnSD5cdGT7uclt6PbJhihrOUylZRCYxiibgOM+QbNZk0WP2fQWKd7CzhbGU/sYD
PdtChmKz5RTSPb1456X2ZjoqHUTbNgU66I0J6uz1Zx0HM1YUuVoFMKBRYgImYFucDoJi3bJa9YXE
NRJttu7KsNQZbs5hs8hhuorI/B2L+ooVNj9ayOfmlubc9FLi3EcTns3caSs78YP3e2AJNOAuTa5A
4/dbAE5kzu/rgxd1RfOFcR7Fvmhv34AWr+U1qQA+QZDRmbUGwX4WDLlbbElqQe1oT/D6AXow1qZD
YzAsGBfJ0q/4zsb2KMuZ4oKEVQqQfmW1wbhMyi13F1oxjrc0mGw2CbSyrewzYdvpJod+b1vk8MJS
8Uv5Y92K+dRnYmtmuuPwbxJDyuI3VJLE/wFlzYPK5gfsSH7KhAjhjkN+HylTeT7dfCnmwDrEdQSO
nExssMxn20WaFWwDjBPUJd3lK03I45BwMPTLt5dZvdEE+foGeVS/2KTwAmsFMeH4OiVyao1Z/0k0
vmUMe8iydCe2s4pEO8cE+GsY7fBedlF/Q4BcLrD8tL6ecO0ZhjlQWX6AiuhtHlPSs4f9tRHQr8nZ
DSsuecVvQJjDoDJ75kGqdB4s/ZQWRRki5CpDQvhDhdYufzsSmwhNljCZzZvEVj4fmO0ljduFUHdv
Zz9iQznmdaVrnqc5+1KBiDlan8matitOzcAt1kuMnQtuHd3EHXz+gDnDKCJqv7VtZGshLl1d5UA8
NXBTNtYC/xSVeES4PD7WE9mJW/54baCYv+g6fCtQlmtfILbSfl/eCCH0v2wBph/WU2LSro5Lw12c
9hzcEZ0o1YD5Ts5ZWIK1Pm49LSP2fZPZnOmQS3gZMrPC211/erIm7l9OIncRDh87R9eY7JFU94Yq
q4IOAviypMJJcr/KqhGekavAbAPoqI0dLg9ntOzgSwa4L9xxyUZlaDSDY+44rAvcQg1AM2mLmM7X
nZgh/PA6r1Sb8gJu6g6HIkDuSxgROMkNaEid6ysqBkyoIM8ec430l0+gG6sj1wGbKldu4IvgZUtg
tO0LhZMvPntEc++eknlFHaJt5MQ3HsLVbc+h5q28zgTwiqX0hIRcId9l2ubiGsnErZCZFWaGerdo
eS0T6sgRIbD56D2RFIiDzNkywTbzwK81v+lqf2Gnu6Uq20yXAk4Uf8GqBm2UDyNS4zKLC2NbPUFe
WCTYeFGd97lz001VDvtdk9xplpX7bcmYf7/6KnVTid/syFnsDWpZr2Z9+B2iWYNPpjH19Jx4ct47
6BQz5rRe9AaOnD8Nz/4QG1pq/ZkRM//CiHMCv0kVjPgQJnFsVNljri+UflOU1dMPbRtWW50lZyDi
LIrglXMij6a0BLYkFd2+61bGJ/QIqSuWbu0Eb6BJy/94limCiN5E9zCziyxhca2ei9Fw8y0ougGV
Phs7yCGpqUlxNrH+HlMrXG1PSTjypnlnhxGnOh1wei7Ph2xpUkT/IuIa933mZac2f/6x9CUdxMVk
PdiYkn6jFZhx8i0U6LS1C9V3wJriMdsoy2X2iyYoWRX5LNF1HkJ8ld2Z9/V5w2rlmR7wMdnwpshg
EWhLLCqZP8K0++TybiDAlVpIuRp+due0uK6Z6dTU2ALbC6+mrr3XEicyv1IkceFwQJjn17EhnjiF
OZCT9OA5t0BnK+9Rqst1BhK/6Zmys1W4az9OlJXl6QqawWm8gdcbdvgC25C/QSgxXG8WDS8hPDaP
/0MyzbgDgzGgu6ot1NaQqVIA4WW9M7l/SyKTUlXGzw23LpeyOxGLm49IT+AsyRK1mMc96sUewIMV
r0kQvcWb+/Vx7cHGlygkMlFvhWPlJ12lsTFycJE3n7+tpqj9hZng8XJVUagvTAO1kRhHLIQ+Zb/5
nbtQqsVE/qwoLnAWmg5FTrcaciesr9NEICRSTBNDhVMmCqVd5wNdD2C+nbT5yqgoeIFTWm2dQjX1
zH1wthNzmEDRga8YyTDcx3ogvrrm3B10uhCslM6nI3/73pL6aoLtCfK6LYYmiZSuH9QIiIftAWPK
mq4uH1vn4bldiZUwWsZNsvSyx1hPn6PrMqYf1Vndwx9gGEwLv2OF8xxEs8wB/AeMtmCAlLmBC+kz
JmDZTR4nfXSPBaN+M1Q59eRoJrF7SNv+rZUbA/0C/TXh2UpqTGrcDi25oQ/AOi6tPAEcgrk3lMdd
hqBm9YpF+1uWh5qhOIfaH546nabS2IQm4RGlkb5aY//W+hEdMpsjiAdRiYU4FzAB2BAFD5Ttps0B
TrLJq6hwq0ZgE9Y32pvOkbOSQxP/PmE+mN7PKi3yLM6rsPyvzsKnCpqfJyDM1D7GAol216fvd3/m
fYdvm5nECq4Jd+0mWSf05aSIknDvOohNBJudyaJS8ZH750ZBH/fmERF+IyOxMbREAhV2p9H/HrIT
SL//XuFwSK/Choze4lVUOcBlsSNdBWrJp8prAfQOADy2E6b2y5E4nU/PQjUwpC1MM4qEJQyuckkI
fS1WCmllLo/mktrs1mjdvwLRy6/NM8b0vjrUtzFabxE+u2Se9H9BBOAUQZG0ezs90p1kNAGPKa5t
Y326Ggr3qHUvwkukYC8MxV6KBwzw+NDkZ3a69za/uS+rrgLksQOzL2xjgGycpCn76Cgh3W9kNPNP
x0dKrsQwECf+vUCowOeR35LpGjFpMtLC/pATIEp9XkVCDNrETZJmwGslyIoBlxjx2sjYvybdwW4s
Pn0l7lBXdrPTd6iNIPB1DE714fU0s0ShUb1cOxBG0+lmxoNhE94lBeTuCfk0IrbCz5HEUYrIlpMK
7wURvO1e9MTlPdpg1Ll2nHx501eKR02TCuyaUSIjAGHgaT78+5ajin45oVx/fMlP47WAe8EYJ3bi
vzgfgJOCTyigLyjw8be/7xIT2RBXKVcY5DHq3KujCnkQeYbX4udgcQr+uWZ4ChRB6eb3jUSDvbyJ
5oPAqzMDNoYg/93lps1fNhluh3iogwt5iwW+P1PRHMZsu3/its6W6tJWjMTbA+89/6GS3X6r+49U
HsNZXvrf3y1pSe6MesA/ggO9CZSPBwkbdxFvuOXFA8K5CX/vnmX8WpbCKDBL6pOy+rY75KS6w09y
EFLmOK6IMiZYTpm/ANk21imgMLXE7ShgAA7PIVGgcxODBibTIYhg8geJSj/GqxvkLSyycuDB9Bqf
uQ/nWvRdR1RhZ1Ugn84ZiuN70k5gMQxNDyLIhORVU1qSKm7DubfeyFBTulpx8aNN0ELMDRnKPJPQ
HSGs2RN/BLpVcDlq+R8Kvz8WZIBYBMtUqdyMYUbmEHJZxH2I+9oyBYYpI8HgQksI4onjLmEyY4lC
3t8YExtBevqW1BUvoecv8WU6UKcmDfQRsII1GhWfjVrfdRxxbMUbjHLwJQLfYzm4GjkTLkHJbWq8
jV7+mJCSkuG8xJhGuQWhYr2+8qREbxjZRX2TcKtnPF8ClB9uFYfIdD6XbKS4qfBKdueAyKVN5X81
abs7i2x7eO/qDGlj9/8sFBvtwJgws8dQ+OLn0RgBs6AAK6Dn5F2HzKa4BbUN6LVHb0hcYrCxm4WE
NUndagX1rNG8GUWOGW44BxVaO+l/no4+1/6VMFBg73XBoI2CJ23f79RT1WhFBWpDPu1oAgAQX6ST
l1DBBA+JE2u9MHEwO1vX44y3qXH75+qZpBNommsP6/ULmNSm6zTOZgY3zM/+lr5rikEmUTOBc9zY
cVOXB4EuRD7bYhHLqpr8dECRwVx4ykJsnpLP/LUd9YleyH30tdIN5i+E4z7dYHsrwWrhqdfRZxnM
bqgc+go7tOPjY34aZqcm5AG8Zxqn4PhgcIbtxgY1hKU1z4yznLzXMYDK/j+MRwLPFHdXEp2fm4qM
VytB9+YqdQLzKGTDVXpnkVsI6dNQtDsisU/W1OzOt7ySdgZul2/QPZ/xF+TscGo5J8D9mbpjlY+b
z/n7jmHhh2neIcFn7FWwMa251BORvbTHOMMjp/cZSVD8A5gB3gvkM6Sq0OYbICYx9IQeuIjHCUtw
bT9iPHnKA1SBIK0AfZnGFVhlTK8CHQyt8nZVigMY7Ojl0GDMxlLrO8nJbWVVQCxwcHSgWAznh/mQ
IdP7r2iKlEaTVisow0bI+rtG90XeK1NlvUFEhRF6ILXvfoVjarusRb7y8UpNgYKf5PCNl14rmU+U
cTX7QZlIZBv0tnrDkfoFrSmNmmG73pZSIrrlhf436vCY6jJILNaAAtJQtj3XLnVIqFXICOymN0ek
rEdObnDDZrefTGI8GClFYJEKQeb53BLZehl7aDlGYLfFM6E5QUeFmn+DkibSlHppF5gTgvWMuOAh
9do8BfpkV6c0WlQaX4MkvHtKK3yUAiil09QFdceZe8H00Z4PfDrG5ECYgrgSIWBcWO/gWmhLCP4+
h43zHVrhCyObhOyEV+1CrD8f/ilN5zdmCruc5iBkoruhZlzFqZYabRCi3XxsKcbpPND0RZ34aUzw
oOsSid/RI4Jy/ZoAywiheif8aXSAzxhut2sVV7UZZEyg7t+mkowKM3BNq/vgkfXkBSO9e6f581V+
H4pdmHbmrNNBcHDI0pMqb7+JSVy/2QQ+yQxv/G1R/H8HgTZ84qFHfZuoWl+nPjVhRAccYwr4Z1s/
OtQ6fqPqcRJaIs8nNsEqCwCicouLw4NMzepOv5axtQF5I4CftRn8azHnO+Jpo2cnWNWQQ0CRhycs
Zdow8tE/eM/0A8kopzsDf+Zx20/4o22IPrRtPmDiV2jQgwRaYAqTgDXIqJM5fZgUbATzfzysZHHq
yy8McdJOolI9Qyg7DJNsmBYY3Ue9OhJw46AjREzX0scHpr4b9sFMYZmbdO697hxvxn3A3iwUDkc0
DEFaE+9Y9Tz/HWQ+89Iz15Hlyq3tgOe89QNmlQhXj9OMhBrfcdQa+kKzDooEgQ0rJdlnwVXXxLW+
jaGIR1Y8E2V9Y3SUGcLlRvRdUVs4Sg/rudSrbkkQvOVvwV53kdWYkJVi1qdk5d3n2AEFzNo0efLH
VKNpLyFpiSz+h0EypS30lSFmRoVCZqaf5woog4PpAbuKm2g67CIUcFQLZZ+QfwtTf5wmc/sCB1Lr
OOpbHLpiOsWJQ/pVfKG9n86nwXfwQEizTGIEu4OX8He0gMG6lcuVpmxgvi3KpuhquXD+4rPiJGYi
zPY6YUcEff5tjAVyc7JtSOUPfjGeKWwz74YP62v/5WFitsQ7HiZFYtfTeRM5KrMDjz0pwra3Hz4U
hxFTPAJ87XbJCgkFq/FlDyIoxwd7ViqS6Csz6p3eKdcPLyIV05P7vCxaFsCe1cH7DCBKXV3DQ5ZI
TfLopTCoZIi9+9ajMWfwMLuxPKIUHozA10O8cb8/wE8/Y8OqDWVOS3zcFIl8x++PmTvvDLkg0X0C
Hmm7vYBGqkdcptxl4OP9+hbl/lH1DOee8HXcaU24K5QdCbHTOHXHqWsEBhH21vyfNnEz+JK+pEdn
Ryr00I/z3L9+JQjN/MciICVisjoAoUImyFDWGbLSjiUdBeZfvsZMF984fvACGlwAxZYrAY/100VO
tjh1WPIpNqTE2UlxKjgdn9knbS2WjUpdxtvavCzfElu1bdbaLxLr7vjZkCVHTsPxdUfIFnQJ3cg9
HNxS97Qegh23eSmnD9s1igIfkg/B7+XGJ5OkWnpR4ZBmMH3Kiao0tYCvmbWaEfnvcDluQQFdvqyb
vCN56GiqRmkWp2WlM+odutXpdS17+vmiRurCNukGXzkr/gr92oqBjP+6fBp6zTCyNKAda2mwQxOR
WAbHI7QxzhN3KQJqMnMFGHonJz/upHbcZH7NgkJGO+BQtxOrdHZX0LGaTYNvF6yL59op4XJhGN4Z
GdVpV6QhysgExolv3mrbQ5KHhC7SEJdmHQ27NqlbOUD9WnsvrWNYHScWnNJXweSPYwwjEQJv48wO
kimbv+LoySzHR9l80ROs7TsfioYFXyrI8bQ3tGjbVJ1Q1X0KC5PzRhh9CoaFym3D3phiYDYtSeI+
yloWQxUlmvwki6Zin32gN12Y5ujwhQGbhp9P7acznG6+OKK16XMCnSFnEEJlDiqWNz1XcvVJf4rl
z0h0JY+vZjFZkJDDgH9Z7FXujlwGsl2GGsTeCKksi8Yy+kZcgdVX9Be7tD45tHrMpR4HOHb06J4V
LvSpNmMMaQ6PVl4yg5JI6mCtyKG/+EwBm5XtdpEabDYgy2ajch/JYa4NwPh7J+/coFAoWrLrjiqJ
6imkelVqCPwr4vc+HC5ekY/u0Rf8ymXtrsLHkQnvayUHkomMU7ZUMouDtCMu2QW7hoqlrCRe+v/a
JDS6ApRDBngk1mZOSGmyb3/KoSig8GrvuchKvRZ5EPKFivK5a/6ju6fL79hb0WwW/+gPQRXzU/Ha
ZKpxUEhexvknrLhNUR0FsodnfrBPu3Gm3Rh28LBXJn7vYx6C1rKXecTi1gcvt0cwxzNWE3xHUsyr
hE+rzo1HyLdT+v7d5hMM1V5B2w5wJtK9/3LyvYDZyGR7Ful3XULYx4VhxWhFuiicGVZTMGLc3lm0
yub3AJyThIQ3Rc/+0D+7ZKLdM8c1uuI2D7ZMn5PIQjHzNa8EKOUKqJvbgU+utxhwjD7zWnJeKGSP
u9nlPfSSwbQRK0/f6R995KEf5lrOHwlAqlm14zS1aOcrR3p13KNcSzxp48HdUHjonHxd+nExM3SO
vFJbxvI9lHwpe0ehRFFl/1r34P5Fv6irqcdG/X1ycEXCFBloDhkgDDHfS5GjMPt0bE5Xq7ncR8yB
nhM4pAuPZ1NA6bxbIzC97dFJZ6eE+Ll8aLOXW+IsTJYAYRCYD3fNHivtK5wioOMWEKvjtE6sO8qb
aYuAaDKjmsV5xSZXjNamA5OSFmQHal5e0OlQyQp4dVvnr2YcVspYPP1BFQMegE6v1I1SVZkUPZh3
6q7JNJB/X1ryXRPYclpd9T79LLRdk8My7jHUTBVjRG43HPqLNO3gYYnnlqML81UTifq48Wm1AZPV
+OCutlAabCcYfPGDoWyzrv3e3jhlKJFKH26UlTUMpJ2Xp92RfXSKhrCUi4QzfiVdWc700tBg/XNm
LBEW2uPTrY8cuzR0fXAmtQZIJwgv+45cevHctcXZooCjlH6a5W3K7Gw9He1UD3evt/XBCi2hSFfD
wk0NRKUo+lZJQ3S16IiVTJdxS6tjWwJXsqRNUq7Ov58Y4Tgi92sghfv3zYvuQ3qro+3oHU5jXNQ+
UCghNp9wY5tJUEShR/GG54+OdKuW4FGLX3qXqz1cNVIx7MUCBdxz1GdTquXDQHdmcDfmDxQnsHSu
TaOEw45FbuxLme7kr85WZugcV8gfJOZfUFz13FzRSo+mWrwSCbU5dJ3AbADQJJ7WZyz6+/6mpGoT
6b1mvRq+QoRt6++1RPddGOVD3nIbfk7blZaLHzhQvIHMlyRgPHCDBIgXXeaw2JtVAeBFPIx9px66
YZ0PjSPrPN4wfyqqAERlx3BGWuH/97v/1S5Abc0Nm9pRO3PbCYts1l4o7Tai4e2gNAacgbN5d6XS
X1Y1nTTFnE+cGmWOMlrjKYArVy+8GnRBDcO45g2L2HJMCNktqMQUBo5m2UMkBXMYv60dCMbZOslz
UxWZbrxBMA4QSlWNtBT2V3f+wMNbhPYJW2npkHNjVrHJnInecOfLin03oqMGgGgS7QC8PQ85zEIf
sDedW7VXO0ytvIA7zIEpGVuq/xeR4J5A3fhpO/mCbQDNFLGq2o/TR5u1KoHIDvt382smVwN7f1pr
DhMkjk0R1fBI6DsILPi8F8B5sc3H8GyvZ8YIhjRTuDHIp44rMAUAZSDLGGOhxS3pCnqs0yqpJPQp
QJ7AfxxEiJpDSpp870c2mF9y7W8qoih4EeNjGNyzTRVVfbuhPL0BpQHzOSiFGpHAcNnM9jIH24uw
mkOIVCzs1T7MrYWl2ocJnrvo9x0jgpLW7DJoL1MimFzpz+/IN6oQMXvtpJrDwSeSCCfMcHYFuOAE
7pqOymmZRE8YMvAMl8h0TdtbQWRgUPulJCnO47mLtyCvnojbgD6RL77OIU6rms/F8YTSNZK0z1b6
e1g6ybnK5SOqQxGdPJCNY/mBZ23elYQhlzz6BusuOoVgZPMI4fU2w2+YlcUeK2pJ5smB+6hndC+Q
XElZy5Fao/mYQ/P8qCCnpdptjddbMJBEnNKPjC+bXAAlzOF+6e8THvd+LXdu2S4tjlrMb7QP3kaG
qZ0jxHWe4Nn5w8vYblpRIk1MTM9F17qj7T4SeUuIlabnKut1NyM4Xe5coLsczvoSN8JnvHiDOhxS
Y/n24QzyBvKQHdIHTJ2Qw5cQ8YdbmX1dJ3kYDNo9xdYL8Z2B3o847C+WDpc8rWX8v+4vCNC5roWy
nBmktLhvx+qVeF2Kk3RWuZbGCh/8m19gpgLhdmmDP2lAgtgVu2Bfr3ASV+15TNnTy8xAA2ZScFty
gI+X4Mua8mIEP0bBCQC1WbCacePqePi3Qdr8jevXrGLudhxEm5dCRzWTPqg/pGmbLMENUKF9RuuP
XSqmMHl5nwny4PqWBROLOyyDF3ebLIqPxQ9ML2hjuk2qzOzG5udG2i95rcVzZ1GwNjNqw1vTqxhs
BrSJQyUrmnluftKXlAHWJdDn2sH7ufWb8YoQBdHGizPOhyq4sCxBOWLOAq5CyZJH9FBaJU5PDuM5
ZszttLgXqbpG0BiNE5ccEK6voiTIRh9T5GFZahNf20MoAhitctyTXDzeT9S0eURyskuLeog0vSUa
Fv5ponsSzShq2U3yrT7OQ6IulhMVAEq6/EQR0LKKJSiRhCWx85Htni6OBHYCN90qtejuY3Ks4Job
3Og92ylPiqwvfdpVIYy976hqeVOyf39bBHdAA/NONbzh7skdwhiJDwqMlYhG0r11J0pqYYZUucDR
TxEUumNgVxifYNgbp2Ed/6x29yEJPXCL1ANt307XuM96g6zRdavrI1A1CxxF50lPeW821od5m/nQ
hBNWmjnwWAKJvFWvLxtLVWoM/J37ZYw+JO6Mwc7vbF0Zv0FCQYdI0T7gu3gNKXlwFF/L96eF0Kap
H/NUIpXQuoblX02RrRNHz/RyyN5UlOkcVVVTLT+5MsKVqOWEnMCWFb70QC/7RpEm2BTDX2iTj2wX
FL9LWtXWU+92VlaiS7mG8IS9NW3lYDSUlbOuMgNzHls0Ph1jEh/Evii+8OmWFXupojk9/N0LMzWr
ReSYcXv38rTr4JeppBYYn+yqDTsZHrun/ZuCHJ7r8RCcQIjumRtWogrycEJ4vLNPKixX7Z/JJHQi
pEIEp1JGY5HJ96ISFvlWFgbxk9/oUZiGBWsDDHTG3c160FHQUuGfNGnsNoqASaJzwcFuh3Wbs099
uic0hyoC4S57yD7hAsNJ9iUg+/AaapSaPVPM3A24ojUSuwNvHGjbJ4SL1VXcIKOre9a9I/z2C7/I
lJtQOWGMFdpBtnCRMnrEerXohMHZckzns1dRZU8z4WTx/6KXmLkyMX5QnLZJaQrbZhiLqoDwg1cQ
tkMwNgIFzJSMOew/Vmexzzf1Wy1h4+prc39lGZdYjq7581oUF90BoDzBNLzTA17uytqjg9DhyL3y
qoICAe/zMGtzMvpGVOyiqOuh9BU8ZvpQZIczLlqIXoAZZodLsd3ext8cDADDK9hUcaNmzE/5cHda
cYIaygFvCN7sF2xwV/UzmthkhaGPzI7MEi5a3mDmcTABSgWkUz+RTwhE8TXtXpectz0IaOS9Stkk
iFkBrIfwRQTR7wdmcEvwhpiLQliPME3apsn9MTQRfZK+1qXC4QqByNvuF5LN2n6nEoA7vwt7YtHh
ZFY3XQtzaY8F1qR26SLQZMl8qs0cpIKI1Fe7iDXtMYJtUIY6nPvCcRc6tTQhqbMirOarNEisVwn6
0UZ9YkkT8frlVlf1jSoBvYzp2U839YGMVydRU96Gk4XPNYwimPoiUYyHFlrXooPNPa/XEXjSdIkM
5aHMOeGD+mr09Me/Zc5A7GWrhx1okbRBLHO/WmKQjSUmr6SsVx4gZ06Uv8DxV3FrIyOe7cEeX31D
uS44wLSh7AJxkNnLWSgfVEjgOLqSoVolQ558/BdBUz+HbOInjV+atEQ7tZRbEkFWRZglv2DBoGfA
vGxgWAHcyd1jG3cObV4ReWcwg5tfL5n1ptspGF5EdX8Fs1S0pItYf9UNiFRMvpIzDzMtPddy77TQ
YStYrCHe6bz38j92KrnusF4Cms6fL6tgArQpT1+X+yv6tvQIpdW16mImZSHEh32aSiFIhbTjxGlp
LV6qscuCk7K789ZEl2zVFdhFDUBTPhLTC1flM7YXs4nHr3eh7Gd9lAd04Okgpba8e0yeUPIu35Xg
+F+AdZzHbjSVA6Bif1G0FOtRExZBmCCNyPp25MvdgTziqV4ZnHovZnVnmYqQDSqT8Z60sIeC3KN8
3NqcinB25du4zCDXXKI8DujpMAIowjEDNg2FRIml9+JATj/dWmAksDrcvVpkyxWsCiWgllVF856z
hLWMVKwHJYcMuCW1h8G73Au6Wyo089SfbNJtlwLetP9vQWbUEyZ44VMn/5QVguuGpyTv+7yaohEG
46RkHLLdZ96q0kKra4U6v/Cnkevt0m+8/JNt6NbRhTInhkTi933MuqrGVVKzOpCHUpr36KtLuqFr
lfAdz7+d5uuiN33rDAGcmqyrsOqi6F2BykM30vf+e7BsHO27t3GrOpiNWMhdfGvdlKB95/QjlFlp
gmdFEDAhdM02vomIs2qZzWhvWfI5dl9FeX4/zwaV4hjRfEJfPChk9w2rbpWl0EH0q0fFVWT7XNHD
9EY+31CletOP93emulYse13xeyRdd4I738bK+9TbhhoYSXJWRVO6ALH1RVPx2nQGDB1wTIpjig8n
6SAmX+r+jZccQAvfC7Wnw7onid1IYFi4/0iQqC5XxcE/Jlbb33YQBks6Tn0RpeF8+2usAI6ZV5dB
ZB8QOTTWDmcoGXOUs3Yhhkviq7182d8+ZSmkDRncfIj/hH6oC1WPUbrvo6Cmmt8M7TlGgfBtzIWy
CfTQDUPxsw59ZSk39ZU4h29oa2bIsrwtg5xUX+o7avZt3VMvNRpi0pvGZdV+CIPgtByDjWcLVF8c
bJI5KCy7idzKxZmisR8I9BSptQmZ9/YIVX4mLvzEvz1S3zkT545jIxBcXQ+lyYqJeG7B2I2ixclq
v2OiRvZWAfNGdl8vk8MLmTlwevhCQbtnzaUm6nFrBNQWZ/1RcQn2ez+eK4qP5eeyJ521Rwn35D2U
+2YjV3PfKS0Rci59nWqkJCUDJTR5KqK7rZAwbTKVtUjCfWkgRHv/iyxGexJYB5DQ/xjxydEiJIyz
vPtLh1tdNqdJI4pld2RMZSD6oLwGyT80+ek9AoW5Kr4ZsmY8Fm5Wso0bvCfumEiaec2tGS0tFbi1
c6rYsBMJKLEJWRUueIsmBAzL9NMnFYWiJqanUXYo8B/8tZLz75AzHIm8U1dZtcYrrOD9kRCXvksD
A17/pusOR6WddQ7sRCMLyJJ3UPoOkbUoTuBnN/RSmVlk4JpCJJzVuiFw/RNXvBhhbsOYW2tIhV08
jsixo3rKDI1VpPotnSd+v5F+jj2mvAGkd9apRdOyniW5sDuA54rrRzrYdcYo+qoYuDFgjipXbMCn
NlfopQU+4v4S5ZcZJoEbASAo/gBTHVSbNflAEcpnQqkIC60s5mcCDC2vaQmUqRe9yKQAsN3/I7J1
3eluCi0PUvPDsn6D0v9I6PWjhjENlyf/QJnNGkqgRajQaAjFSeIsKvbdKRoT4hOqXHhnHYRKX7n2
WsC9B5IZYXxp6NEW8pSSFzTUqye6fFJzkQ79NPk/A6o55yvSEKUbHHtY/P1MnP7+g6pdZIMR9Kx3
uuXPaBoDIZXmBAPQYL9i7wJXlcR3nUFpY4ZxjldfJ06VbuEW/G01JItO6VdGpxkwoiY+zHM1PkyQ
S+pSuw7IJnyz2BgfXR4d57Oepy6Ey/xTBmT3YtneBPgdgsa8rEAmMeMwG/1FZklhCXZVQWLzsGRH
ohUPvBPh590N/m4HbJIIxdUYVoeVJtFxbPnZV5si1caRDqPuytjR2XmotED4BJVE0xgJsdBO2pv8
SwFxyYhSLScaO+oLxi+QbDPyllfgLl9vmqdAYA+a0M5ZRHF6klAbMJA2ezf7Z9Qyy+4tgBZPAIOS
wle3Xb8EMx1AZ0SyOZkKzSvCULAI1FRkUL/S5HU1Mpqhcc09NBv+gnq7YR3fFboNR7mHW7+TI0JQ
/iiieK7T+5Ol0cMG2oMXGkySpexdqs3vKIii9VEfR2QcnqLzOBf5JB9w77jPnN6lbWjttPkuU+PI
0ABT46qDv/ZroqcVNhsdWRNN4qPtJeVzZ/ffv4GA6tfPcvHcR6Y3GmnGGg9YA5XSLlCaLjSvT143
ZjyCb5N/D1bOSZ6jFz+ZY5vWOJJN3q26rm+a2QXKCLe9JVLLpK1lP+ebRLHBV3oudrr97YikFIJa
cPLy4vW6t6JdnBin6CMcB02tcHviPUeeOLJWFzrjcx/b5/bQariQJpyPwF7871pxJwjOXo9GWz0v
Gf6/bd3rVkvWeDBCG0RTEqU2DbkHJ4xjSqmBhBCikBMW6d1q0B9NuHL3x46/xgl6WFwrSY9+sj3M
YZ4qqTkNbvMtM1RGKMfzsLsSJAQn2XJkQUK75xvAIMwePzikRzYF8uOkhVeRF0W7crnyQdAMbvpH
V8tTMcQDHApv3l3i9q2ipX0MDUYZKx8P5qZtTBKQjq1+pd2AB1EgWVtUXe+J/iFFtV1RvyjvXCmx
tOvnhzKvdV8JdMjSI2NoarKDV2m1/QADmeTnqGhSSqlkzFNTwk9J1+I7ivM473NDtpmSieA7yLKq
CyrADglP8dz1amZG7yZPg1AwgvWhoNNccrPvsDSa4GF601+afX5dWRGlVyZtZvLtTsc3O/1TMN9R
JS4bosJqI88aMgmJHZOUGzyXjvZU/O+Ym9WlSZBrbkiBVd7Lqe9L7Dln6wAADH7CzGCmMvllQuh/
iNDT5dXFhP+bujhu51rt+mySVCC+Xb168K7au0uwRa/MDkyEb8rmopkROvlPJtss/Hltn3Yf3u2v
pF/XukWjKQS/BgyM4QoDKVQIEQTNMWRxWmtyFWdJwLdt1LL6TdFZfV3+2jHjurfhVDQ4Z/PHqQG6
wFwWnqes9LwIHwLXYvXo4gWqMeUfLsfmjS6vL1vDnGwNWxOhhyDIaRUOcXlsUoBs/yrSSf5llzUd
8Cl535VLV8jB/2zeEl4OXWGTKrCDiX3iyZ/x6HRPDWWbAu9iDNIWaaKmzvuaMfvVRFX14eeMkl7v
InjRItYgO/OtnKcD3pmPNgun3QqHJRHer/kyO6XVySkZm7tcddYZjtM3eTi7S7bDXyE1EEb9Ql0w
GxH6Nt8Fb4U/1aGyTvEwgOD+ZKpJdpre4ba2XAKWdlKAPlzFdK4GxBUxNNlp5phqS86b0pATpEh4
oFd/MOtWJzhvvsiWfAonMehY+2dECI9yxzu0+dLLTqj9GkR/4jSmJko1BglIMVrQ5KQizzuCXKX+
/MeeGIkHgbW0uYZzU/qUkG+gA+p70zZRTIThl0nokV9UCRRZ97mo8gxDdHAf1FkPWEuSlx5PN5gJ
HwpwsPMACkzkfVlE3Ary/iPcz3kUK2R+C2xJq4Qzi+gfqEfFJEnLTgpkUWV4ZaC/0sYuaceeIQ6w
Z+d4Y0aZZ8UhsUUlHC3N+Sp0A5xWS/ubKTY0pG7jVFbgMYD1RjMZ60SsRH0o+bLyaXwli3mcC/MH
/S6a27jhkAyUG0h1FbM9Y0vgpzJShswP3DowUak59zfb2z1MtWu8xeGRAVg0j8TG8u+3BkPb1CqJ
XZL8Ml508zRdYItRJ2PHrhi49UgZaD3Uqei2U/hCS1yGBWVXy1d9n4XtjzjFtC4oFalmgpEeDJJu
sUYBttj59G0F5chvnEOZ0owKGN1dRL103KeVzRs5xkTFnIP3JOjByQynMHhEQosML0PkfH4bf4M9
LLRcd3KFCRRtteOs5du3CSBRRSE8xz9dNADfmigYgR0XHvIydaz/Oaslue6Q6Kqxas4mdtkZxV7f
O+vpN2pDh+XmlEBNz/jKdz+DTtQ06aBOfeCkfEvj04hR4ZP68MTUfkZESm6QadzQMOpW6Hcsyl9V
xPBvfOjPxSSuZZje3ZOWzSIVqGRPi54747O6ufDXW/bwRuMbncjaYVJLNGg/vMELiyIcxT+gsGo/
DKti0xJoxSr6GaDD6AmHXmh0y166l9KzL5MK+J6LeXEgXmADIuOE+IAUNtLg61V/y+sGKI+cXHvZ
9X8J9RKjXEu5X0f7an+BDL9vMS4Ai360ICMSrrEhlFHxJz0MkEt7rjaDvzVbj8yK1uCEqp3U9yCy
ru4xHjSoL390rm7Vr12kpBtCX+nXQvkn4tDTZJuxRYHs0rHRE09Xwb/YNcWPqOA0aXb9uLXLYemf
Vunl4Ejt4KnaF28LCnbmTIPqnjw8V3xldkNF0G0gWju6XXY8ToPAZNpk/P8LqPLeF615Amu1SQVP
aCNURLVIQPb01hEXFfD4wI9+SHfDXc4dHnQE0oM6zUnPb1vIHmfolE/7YjOTXHJDJ/NCTDYN4AVE
1db1s8Pzg+jzlncvCfs5i5uEyyKWQOMM6NX0LyF/gA/rn/VvzcrWjIXRhmz3A8d8kcIK5JXscH0j
tvsV0UNs62nZXxpIgYBT6uoJxJ8dhIsM33ABAwlKUuCWild3F4cS/rQ1SEKrKxMPBWiBZFBQ3S8H
Y+9Z/r37RGAhd4S6WPn87CHC07XC1wFV2aQLmdMPwZCyr8bmnZlhwrnPqGzhRGC6pli2V8PD6icM
aM2pDQDKdPxqhwsN8uqw4nJFv2tmPcwn6X5L0eeQIt6ZhoyxVOZmRmFGQ+YBlOWt7xTDfKo0LKEI
i2BkDAHYBky20dT81pqvQQVRpEY0unv6v6N1+rgMdAuKSRe73d+Rg3/sLGQVnxOgzi57BA2UeySy
QPrtEsl2ncQaA6QaMdrpwhSZeizfVk+PzAAn7J5GszDeJAPrPR4TAwGT93DqwEQRzS5vflJ74xcY
WmVjEy7m0H8sJuA9hdr6TF6fbD2hW+crnZhwXUKvV3hjZM0M8wevU7VZ2AaH1W2YLRNehfTL1nUA
th57F8qorTzieCRq/odKisfigE7pCPaWDE/Y20Ct/DjLvU7h976XqNnwsQmNFW+gyxjdSBIboIEu
ESWPVit3CwP6JRTclZshp5NWcQmeWKyYSx+1QPBUNlGn9C9BbwIdk52zowsEoG3Zy/64AQh2tV17
MrJjM4Ig/fqdu0K39G7dttmlgSLLqSKEOchIRzNbrvYRiLVIdPFFDWc5PTd1Tzb9IlIsnBHF6hGq
HgpE+NUBPRBSAsu9T6vyKxl0WLAJ9XWkZ6th7hXmrKXVAFydWhcrRrFRO+ibYcM+mk8iKzvHarHD
UmfUB1+Nsugj1hM9SElk6LDTXCiO9k8hlokVjdOlGYyv6a7RrVoVtExUTN5yXT8umqPzzjTGzit+
XARlsbzsx2xIOoFtLpd7LKunbgFhK9N1KPsa+tZOXjbjwwlNGt/oWjQ5bKck95Ku7wS8gtL2rXZi
rvyJLBo/3wV9HmewFQqGIkp9sMU7f26Rw5ypqfq4mxBvv/rPXbcu5nw/MagkO5A2iwieSgBZTu9T
UvS9mjtrroyjpK4Z3CrPa7qilnBrFA1UaJllBX8lmDroN5tCoX7WEauGuO9W633v1FJhxTF16BXW
RNV0SrMDIn5quc5WaphajhJl+CHp3men5IRqvJBt0zcKjJ/jDWo+uio8SGTn1Z/NftqXuAWPLJiq
08KDNxY4sa97BYPAsE/tlZzp8T7q3Y1tOOcuXRakRHP/o/3wM6Sg/mK15WRTXsgYy+hYilH/0HV7
jyafvd9j7KOtmoBPd/5+wp7om8v2SRU/YTsEYLIwHMtg1FCyHXqN9Oj0+pILdJLIE/Knn5VZze9Q
w8xjBBhFlAHpkJC9PtJxk8A8lg0v9J8q0zt55bnXCpkoUxnlCJsTsADoBHUSx79911BMmMs2MX6p
0owpurVptmOhDqtYTjn7+mlnW1wVyNH2LA+gNnflpwRufQugG97L2qZwMoVD41bOUcivA8Z1SkZe
sTXe2P9PyVvSzw3XTp4OLpvDPRemH8rVGTHabpBcjQ4dE0jtUi6snjVVGnE6Fi95dCig7QyyGCHB
QvL2xigoRSF6nzYLJEHAV4BVUtf+NsmyDzpTTYNrGl+xFimwqaX7ZRi2R6rSmOLHndkOACJ8fp6m
GfczAX3U2/zR0GaXQ3Yiiuk7Fb3wgAIW23AhGqB8YI8j67+wlBD/ao2gu2RXjhyaArnnEHleXxrK
I0WQnLTjdcoyH4pO6OZdMBAwJLCU1r1sd70zgBn6sr+cFyXs3kCXZze3l9PMuNGndBDWwwkkgELl
vQ+0DCgpe8G5YNMwSm1fO6TA/lUmFtzVrkyTyDEXC4Piwyvjx+VwlLuJkOKTHmxL04cwzsubeg8m
O944z24xqbyS16JYBT+2SUFxtYi6z6GZFNoa2x1bf5fam7SIOkJoiYGUQVlf1NoY4xaI7eGNV6z0
86RMQmz+JZyckECicO6nubQxq1kmKYgf6EK/jrfkfELomxeV7Isx0+Cj7RTVmCGVznGWgBJ7GFMR
gpmdN7eUhKPfHlQZcBVnwuXGcSWO8sMkglCoc881IPtC6OCjqVI/Je2Zx/wss1j6MegZsRL7QNYC
7iU05bG94XNL/AucLbwyHHp3Sn33TgvVXajpKt8rjhUg3a8cYOi44MXBSs2FeJY7JzCsCgEGIHXp
bbiIkihtw5reEc0IJbSu2AwPsS1FOhIK8nvYShv8ke8AUMnc9uwkgP/5L6casSdGiD8RtV9/z6fW
rThBoQk18zwucmbbpQBz3Nb9BiDc7TuWthvYHzEg5NUG4+Kcw17RSOhCXxP5Sgi4y24r9iA+pJAC
jaEuT3eP8qARySQAVDrOPLIh8kd+I6vL/CuOdCA4fZKHA6f8yw5JsumVQRMTQtIKcL5DUC+K+2FL
3uLT3E5zp4kHFk8UJKCWSWmAUyyt9EJ/vxub5/ZXF9CuhA4lkkD8UQY+11Wr4c1ArRq5hYqU80CZ
Fs8Nrtiy3YqYFHUN+qIq5aonOgVesS5lv/RnoKt78kCsAD2l6pEmP3sestZoi4sVsuJm8YuRK5WY
mCu0IVIdpC0ZsNNOyDxNosmBU/s002CBUktWjzjYOYi8Cb4Z6esO6P13JeGa3GTphahf/Y6aDDdC
9QmN7TpOyb/Nsnpu2vk6lAXUUGBKtLPwqgtyPH0xLWAfu99TXDedCU6nAd4w8WTNNR3wdg1y8JkT
VPnhTcGsnbnmLcsqgnm6Al9lgFOwtecd/cKSKfn48QPMhUfd+FIxJfYM0nLsBC+0mkwHnLjdd42y
gkryH/GSjIZMYBmNCnNtxBbu2Kqlx273TfMhOBlGl+tKxTH4dH3zrObZ5MUVfRFadiYrgShbh0wN
gEO9hgrjEnlab1OA39zoNYXLB5dAelJWIaEQBG6e2Knpp2VRpP6iOPzOjUuMBOl6r0xwQtg9rSz0
BNh2BlPkzPl+yRSs0HPjBtSmc/wnCOIt8zHj24P0NEA6If9+u8jO0FiewY4vfAfiBavfAnFWDyEr
MpDXI8mUtQLMIwWB7C0ACHLXQBMHt+QxJ+ztWgkaVooXFzuojfdnwrGeEeMdKjNb4WMjOer7Tw1S
NVTo87Hnjtl02u4S24RRUWKPs7JMGBn8JeC3HYjcc1s8auJWbYxcSjfbXfaq2aq9/im+0AeUb04F
MQrpKoFN/TicL19pJRx84ExYk+eXt3WCTByfig/2ZKJu37So0ybNggDfxJybkLZhVLWYdoHk7RB3
EksJW2v+qmz5DNV2aPNSHFYMfClOav6ZEurdQvHbrax4HdJZG22DC4yh5KBGg6aU3OnPjdn1jP1i
CvlQeMCMiw1lYh4J/6yF0Ey30fcqQmZF1e7iVAERdVeX6fKxVrL/KhfJtOZFcoVyeUd0t2TeB4Up
LBP95gstK5SnLHBq5eWygntZKTlCNoM8mZSMhxcSqIQS/y0G+Gd/5t7nhJW34//g48vkigDdB/O5
6lcs9YLcH9SXA5iW63DneUsIVN/H0CW1Y9DWfYUssfg/I24xDkW2mbJWyaB3lhwqDT4mlLSGZ4gB
asgnAkJS5UwWROkRxV1YwJTEuvZ+32S/29ZQJg6OY3WSXiN5/7O04wi2uB10HnweSRAM8PfgazcE
ZSRPMuYQmmzIdEhwqsCZEP3ODyQ5EKBWJsl2U1S/6SEqc2xdfUEM2nFDXtOf/UY8ibwM1w2/qGGS
sViAEVM51yW5nZMwisA4UIk2JxG3QTTED+zpBaFBOBoGc/bygyGzaoVZJIi7ow2U+70PBAFRerGX
jh7lzVWqED2r0rWOlywFEl0tDX56BzdavyDAmHYo4bHK/QmimBxB4vmiZONGvqDOFetl5BMQfakB
2fGC/pGwLcEcV8Wiat09trQgIteqXVpMLkcriCDTKx+DeJslbgajf3dPaRSqNFW4vpm+CUIFUnmC
H8EuIks47aQYgF8TZDVQiwrbP5mK78urvIV37k7oFShodeO4vu5FyGrubvakgscCZb77oefwOP+H
N653V/xFZf9R/5tk51Ofg3aDZkhaWsFEdd48j7eTEs7iNWUBxutzjyNexcn1VPlhWAECj/dKrK68
71RLIWo4pO6CpEhBlL0hYdMeWyq/8+w1/uy+gP+tciMMB0rhWpzQR7XG4LUk4AEuAB+qsofNEsWA
eEOnqF5BgonlGFChP+pAyIyHhNbnpIttSuZtJZTrjp7dW+965yGsd+hImdzmrJKipFe1qqluP76F
6C1TyNzh3cisa88+2DAHn2+DGUj//lThKO5wUmCZ6FwPskcM3IQXOtJMPuiy3ljytoNqYPYuKqAc
iyvtsfgqc485nYC/4TZsH4dNmvzJd47yBmGE4GdD6dk4ABDr74XrV9UVqFdSyFPn3zpORmORyp1R
ZZL522t/Wa877rWwnOFMMXUhdVwr9sgJk7WEDmV8FhLxlnaFxaEr0X7IbCnQ/1u+w+mnoEWYIJLW
uECJt2Wd1JfbGieP+L0z+0W5HcGnwHJMVKwxwBDzt74rXjxQHU7768V8XfXbdMlgK6Sr0I3Idg4J
P268NmLXtN4ghtwx13s1ZxSlvApmWW6o4ZBtjJNy2+dOlFEZCx9+IUfthcgCrLt9gBCwnrhOFGRx
mS6JZiyH92QQpVIfdurG70q+67NDEKRPCJW9NhTz2a8s/VxmgV9OK75za76Xxo9BxKGNbr9gJgFH
xWR+ZLz5GnZjk0aWKMKcFphiaLvuj5C5LR8t7xxPpco1+9Te15WfFuFVk6oE4oIq6HDbCI5bfTVg
Hp6Cn+IdywazvHevJJwOjOYUGlMBNzVe2ziIR+6cApKiq/xdNB6/weu8M0bdUUDHWBRQcTjt7JGm
heFyCM7FrrAC/ssBA2O4bRQ0GAvB4T/ySG2to5cyJ8yTWZ1IqQV+6ufHPzvb7ZCQf0zreyQKvoiI
Mww/I+fNCgEK+gbgrFLjiE+PGH0+gcNBq+nmJMVnmhJBhYCQrh9m2pcieVr9cxOy+L7nzpuG/L6V
iwT12xi2Le908aWR2hfIWbvKj4lG5J+ylcJYIVSikOZ3lKeh2JYR6dgjPt1PrScx+UFR7Mz+9JlU
qNd0T0EoYSf4SJqzZpQfDj3XNfyp6YOO6de3eMW+201oPOEIy9maN9UZm2C+njxEYlLG3QLOKtw/
h7/sjbdhI0S9WIeGauACJ0EGdCl1RtCNElxlo4EVulfcEQQFS/D7cWBXTgtAK97HCzxcomPtdz9z
aH1/MPuOifkNT26gHtMZ9cgY2yvlejFHtePz7zdQO5HwMim7OAS4PqEVFnE7hEp+XwfJ2NxdhBWP
5Kn4AWePBuPy5ELtHvg5slc4+g7kHyhl5hE7CB47MH4ArpCI/OZXAa1vX21UNOxeNivzYqvGAw0k
A7B0gEk3o+2m4sO/zl4BeFDLQ16GfWPgyzTFwnmW+GOBF2Q7UDATZrG5fuzNK9W1sxJCW0/0PKUH
bm4hu0WxNZ2m/uQwws4gBowdl4pBuZNjxgBN0G1PpMzxxeeos7wRAyqqJ79qGtxEJRPteEBqllad
gJIWVQL5kSmMayydjTWsFtsHZI5h0W9EWHCpoBbu8eFoFJCYeekq8NSGuTSR8kIXjlrduNwk+mT6
OfNZg8X+7z1qwwQvxNg7oxl3AI67rV9iQFPhdYtT/oGNkjSSiI5/kvPEOSU1V2mX/LjiE33TJd1p
Harvz4sG/YDrA7knzSKhSSFzp0nlzyShj/RnPcw4cmoNaXs6BhRJ5ryEXjRPh8G36c2Lzb+a73Ts
kHxDVSDN0dgLV7ghruiBqkj0LC2Iebv2NBSo0vVmHkdTySfd6DNPOS4VnczAcdk8cjZCV/cH41OQ
tF+b8W+Wrbd1UQjBOrfTKu3AYBEt/0p6B2/F6H42QbuhqCelRTqpyfsA5FKgVo+ItkHobMISLdqP
XiIBql7svtxuxqLG9ponvF9HeHh3llpoPgrBATNfB+dyxp5vQhdE3IaX3byH1JAyHRd9RNkrviDO
2TGr4D2YoJMJ5EL/hsRxW7Ed+V8XVnQXpyyd0tTbX/i9E8cAKGs2c28k1rIG0wAL8ixZABGz4faN
Pm8rfc5VrhzP6dGjCDXgBbn6BpXD1nr2PchtbhiIN99xIy3LtLxjtvTVB3OgzCfhwQy78rw7srPd
R7cHm1uqctK9UeBfnY8cj2dY1j5ND1g1Rm4Mz1icU66Y9pQYLbrdc8xMKRYRb02+N4dVpYPomXZQ
XlYcftqWd+fsDL/UsaTvntcWrDvguuzkivU+wttfx7pt3xkx1G8+jVjaRBW1m0/0XCPd7rYnKhvq
vRexPiPYwvRWYER5CZESmxw8IJejv/STrSP/0h+/sPG4RhXWqRFDoufuRQI3WYBXJIQNTA3h99Fj
LSf/bDsuAv2IuAzxQuJtm6kppU1aGGU7wh4mmf9s9hDjZPISYywBgRum1gLzqvK+m7FacHdW9sBc
WDKLW8oovf03GbD0asTd5clYE03UQNY9HvNLw9xwmpTykT5S92niROU6GD+MXsTA/tlefQh4RWza
nN8JOemDvYYj9MSJlKnhRGmN9aBSXcJ1KNbJHgvsEw3V84OmtcDv8bpOASGSyb9jQOlFRNMNbZk2
Cb93T/MFSC0qCT+VFODLJHpzoAsrR5jHMpu4k7o39JqihEuVgY13NwfS0fCBuSP8DdMPdimM8N/a
xaW4YCU3yynIc0DP4twSq11PY1lo7t6dhtCPjajcUDbFCyuW6izEa4SYgcyiZRkOQf38Dzmh3RxO
CDLSRokaIMYD0BGBzpZ4TFZpl1wKmHbxAQ7D6Fr5wQTS8EVs1qvJHYDWw0DzztB3uPX2ot6/znEX
ttITUIRBeIpDa2FVyDqQalMNkHYwaKcZn78DJ9ku+0DbfpHub99cwf4WF2J6owjCz7Qw2JhVvr6O
zdoW8Tdl3o/yQ2U1kArGb++BUooFLyordawJ+/8moyIGPr5tn46JDmuRrZgPpYOmK4uakXM/t0af
6iG5lGOcN9W7rrxxbWPWDJ4jXpHCXJqyAjVLh3pymZqaeAKsoXHLBk60Bd5K/9puPzBXugpp0oec
EQ8S2VZ21ssDTAW9klhTG4ZawHK+aA8PezyMCyFyhA2cYYl3FDfwWjdBV30mfYKVRHx1E9SYHGcz
JEksBvbm7SrmwkvGT6FADD2EtxmpPvE+f4zzL3c1uYopN1h4JZPJFUk/9rrQTLp7kA+9cpAg1dZF
QXnSDt8gW9QvPowkjBt6oeoNCfkY8Gv+9Ty2yfrndYAdrarKHzn3IaOF+9gIuJ5jL7CZnqgIwwPt
IpGwjGJgJancl1txUNZdk42VcGyrx3ZbeG+uCe0p9ylDs+80VJFX5iF8hXMaECh2bwS3qzac2CeE
o3DNd811imFws+GXW4tcaPgs/wNnNuKebndi3wlfZfSbneVserTGVeW+iPX83nEI+gvmTvUeX5dA
JPWCKe2g9tsYmcpFF3kFoR26pi+lD3tUySjZC75fsJRngaC7BBbuNj2RcrXv/MTnufuPH3urRTLY
Y8DCF+kthNCuFQBf35BDH2ZV7W9jRKW84YtfhR9Vlh7joNNxSt2vHlTTsq4mSekw43RK9E8AkXaG
71tSOd9ezHRDkFOX1dPCNdqpy1vt8tQO6Q4hVb1veoDXjmJXwELcIqR+JLvDtXRB17GUdJPnkUa2
YHx0n1OaIuKG84uihWt3Ayj/a1XA1KgJCOfxfdS3uFfr4Sxe3qGQl/2BoexCNUvlQFOmOrWjeH/7
VY8KZfZcTw4E8rp0hG8xLXN7z0flDKZJzt2JXHhaZ4S9yEp+L/TpiAFnRih7lF/TM/r3uqqcUnPx
KLlGDsWb3yjcKlkm6/nBngQn13QXJ8Qy3GFhUqauAkHxZnCZynlz6E3eTlLSM7GjueZFoZArGGeu
OZxIahXG665RdR1RP6dQZB+t8cYSBjmj8r17M8aQqXQjZ/F154Z5rj49OG3dGL97H1KhPKvTbbia
F6Q1LSj0dBhsQn5mOP2yahjqgIN9r9t6/yGkoaESVpdUrpayty9Lj4ZtiyCZnnq1nwfU4cUA4Juf
yVvtzpMEB8LIyzH5UXNcOmZHh/iZpiwC7GcSaVxLHUqW41Tz1FFO2QdJf7BHSwE9zNwVmHHfZH/+
vcbNed1sCm/r5pzxJsiV55MtsNzWlnrsPn4KUtWtkfXnRU7pzFcwG1dt/Y/4adwj5QlZBTjivtzJ
inEiG2NRB+cUk1P5z728HwoJ8sJNF1otedi0aeogjMGUqCNLVwVIj5FLSgJyVQa4urjM2XdsvFEF
X5lWr4sD0AKNxYbpLJxhFTVey76mQ4ljtV6482QDUA+EXwb+erEGXq28vBIx8kVIdTVA070fMqp0
NCwXh3B72ZFs59YFvoyum7RU4aFzclzwydU5mjkaV4ZnC7/Db6TOFOlo8NkbC6qlhGyofdIjzbaI
/T/QFnqvgqBVKMRlALAvtMceJcrV09Ea7JwFucIW2wk7csCtLRMl2WChyrxyN+jYQnKM+iP597PJ
LRLb2qMdikVekgrexcySewUoyPPDW+wTSnid1BjUCOk3ioZFGUIOggNFgdtXn0wiUwOKLheTVJF5
tdF5K/mN7/Aj1n24vlzfTz4/4EqYaXpKzVrK08mUdOYUiL+8G72Y6LKQtg7WlIWaFbzCWb70AVkD
hvbS9fKqpI4L6dSizRTWkgzXYBGrxGIMsYlTFuGuUoz/RF19j5Mn8aC2nI28qahgjzHtwuZELuDf
hkngLSutmZLOP7lPFHFUPjpltVstJ9zJNbQqBoKmrOuagek/sjaA5uPXJdAccIUJ1CyxJn/Ny3+q
RCKh69m9NxwOxPbXUiVnvF9RI2X6SS+RC7I16X1hDQBTUZs8pHZ/lJiplHi2/6ZI/RSOpkkFeuho
PSwe4BShK5xeVi/JI2tnBUX1ZCdTqttjraBiIM0wp2wXuWzWU+e4N86ChIUhrmR71S/sKqPkfEB7
f5zput6hhuZx9orwIBJFy03cE0Oix/DaVc95UQipELJlEud/fu2zlRspU4uwMLR4o4ZMoIDid8Gi
Vp9N3VCvmNT189hEWqgWPUBV1b50VWFa/EiOC2Y5fUgqvEZLQBXE4z8kp3uR3+ToaOoTvQkW43Rh
pzz/PjceWgtTDW9LYYBXS3cAc4QPmT+WLF4ChPdx/cbJVLuu/p3paPdOLaC3hUMFS4zYFqCTed8o
2nQ4sCmKpRaz0FtcyWD1TNip2ujpfZeY6Mfz+YEVNdLwTavXs0y/NFgQXGCqQr4JuWGcHA95E5eJ
LGmQRelqvBebzPy+XHutmEBclW9lPc3razS1idVvf1Ap+lms0zqZhs6PZbinDFuVRPo/udBISpvV
uInRlppGbxDd5z+CikbJ9/2MIOktax7sLa4LEnAdMJAHMyjHcJjdhKTWQ48EpDrtVjcsyE8K/ecH
jPvXO98xnROX39bJ4tMM+IgZTeuOAG4GfJWq3ZPI+XvLCk1OX8DD5ipgoWK7krf2LEt0JuuOn5rZ
61uqk1M2J+QrY0QzKlUfixVN5xrW6hMMP5AMYJr6eEwhBZsOxd/bL7U1rlBhss1RyKaenGjcvLqq
zKEnm1gOmlAt+dSwm/PiqT9RUmHkCPHoqSHXBZzDnZf64QDCgtMaO9eBXxXPWBtqxK10+mWfZnOQ
CxrH8DJhE/J2lrE8/uCppVDphPG+dZGqzArhr5q2W/kSVvu/+z1LzEzv7AyN7fSw5GVQpoGoWTzq
tqSnmsysS6bqgKNkXNRDJ7tb4S+asrkkWvFKj2e9E3TNQf7DOV8mPrZbWGiOggFjKaqXXsmANwGD
EHa4luUKKmAuSq3VQYwWtYPfSm2ARladUgf1coWaycuho/topsE7oB4FEphrW/iH5j4vMfj66fE7
A2kr5QlGcui/7GYnJn/uRf3xkluDkYtkW6e5npze6/XTkZL+xHzmGhR1X4HZpSL/jAqKJEbVdPIZ
XEM48V1PhZ5TmoXr638Vhd6lnaj5mcTt/UeG9DY5zeAh8mzY0qswvksJSQEnRbM+Z0H/tTWzogiY
uCLFoASTXqshnPbeVWOcJgFoKMBAEGjgb83yAtHDM5FKL1KK5aJ1gs5dGeLGHpOoSlXe6uKEsT98
Ovm/eSW/CtiFB6Y6pL1rhcgGtw2ISYlotnvrdlnojfAfCAc5MymufVe25MEiyBx1Ezps//U+1eiU
jNnHFhQC8Uym+mJw0LHCo3oCe/266S+0rC8HtryIcDImPDpGUHHiaCe89gWt/rC1TlR0a9R5Y+RU
TlLCylqx6K4fvUWMXnZKtkPQFoSq4qbw7ZOe9izAT3+d5k6fwZprvJiJSolOGL2D1nSrHAI7QSYK
SKMholt/bXzfuAXJP1jOTo0zMGdlbfoXFGkPllqApiPLTZyY2ip2cLX3UE6hmCxZdxcts5LMNFa9
8Y+xFfCYyotRNnU1yoZs+BgK9hute9PmGES04bNFz/xsSgeGxNBXFIPI/pcVHk7OwZIOIlKYF7ea
UwPK9iIgembA/yXygCKOFNTUv+91jpb7zd/D0JUPqE0Ha3tMSKjOljPkzmYtnUC0+0337+414JHD
UTwBSgk8mvnd/mkpP0vM/iLmbT+hfz/fVC0mu+ZTcg2bryWIZ+bWu7FC4COjJViMaFs65rdu5qac
4BE2+53r22vAPSKL5XLnBKID4XbxHSZEJ74QYJE6z+vyuajawM0RpQYUinjbOwORdxWspGXYuMz9
qKruWjYyoJzjrO4VOJsyaPx6dn0J487MmBRvEOBA8OuJx7oA0joMJIp/M2sd093VADUUH0AtsWGu
WZZMk05gm1LEFh6P668nbH/xLcUhLjXnrld1ZeVQiTROQHQtz5wrLk25At9CmlbgsZO45yMpifJp
iy654sYPWYfCO3ZjrsEQGGKW+i7z96DbQxw5cxHdoBQGNXR/LSOdPHCl3lsOqofbPSoxFxm3SV/W
e80bQK53CUUN+OAWn7GeegPJaTtq8e2lXeypQGIaZxW41yLOxqZj/vPCKXKQR/rMSzLB2QJQ//JT
6yIjiMkKOKPAiZ2pGaUFoD8wfflEoW4zaxRT9u0adlFQ6oc9v//cVCi7RC4En9ABnY0Pg0PiIjPA
QGjqTvHIbN9R7n5F73UWIy6ehHtO9+9dEK5Yfq61wIiTd7d5LawseSito+WTgscA5h8ekOtPBEMb
CoFv5h/zqc+yNpU+AA149MWi45MZLjxjuu07C3x9qwjTgm445Dd3kj12jXE8hcckXs5PBHaMlEVx
QpJ3wtU2DIKDAWBKzfsWf4NEwnEmpZtErwD7Fck5DqmrZsdWj1AaWEah9P7dx5L044hgNrk/YXRI
Nn+z8VsFgI/TVsbSNO0CFZlqjIQ/nnrhXymAZk/qUxBVQwq+bFhcNGqQZhGwx8p4clRFgw7zEYlf
/+vBABfAC3w4HbMJN50j+YV7WxcjF3RFqcOvuTZBGm3nXGw3wVAuwp1/NCfSiqm02YTDsU4ydLm/
Hern2T/skpyamrCZx6VocphcyblaSgMM0NDb9Kz1PyoRMNQpKc4b1FT07gbmWJWL0/LehnQ5HTfv
0snYDPKyQ0UPU1vQoVxVgTJK1+1a4+hGFfTaCg5RWQFUwiUsgR/lenNIAvO/+yIVVRAExLuGAOML
9UwmMMzhZ08krdkXASPgK3mMO6bF86aYSn6bORpG9g24tsCF97qh3L2TGk5bZN5o3zHt84DZmuC4
Xl5r6oG9qpn35KbP+j0WnbTk6brRJmTM2o65Ho47ZaACB1vSfhyDU/Z2cY15+7UvRY6lVeIr4Zb0
N97PlHp/PGL00sNm8w0NpBhaqGFwu8W7v5ppzVd3YRjBOKl2+TCYKWM0eUiGZIYYEyf9/BIdG7yF
5QNs+YjBlwsGnGfABex6sGAyH6DNHLXrXuU+IfjcTDGoWv3g1tFIGU0qmqXJ6PBjXm6A3RFRzqo+
KTedoF30g3ihqkmKoAisv8wivwk5+RSkv9I7WIZJ4T5oHd20u2COqI9mrWmb+8NW68QFpEhuDfud
Cq8kpVf7exR+txR4Sy+KY1RnK0/G4G3ciZ47o0nVSbFyD2FwL9XG6jlSRC3TiM4HBPPLzIl9tLp1
/wt4pU0qd+NeWfijF0+CbhbjQ1iaclJhecqZLP9I7/krrWx8paF4nKWYAES8mgifvmp4pMggEOON
yNB5kquv0EjtKXQRL475hOsezS0RkHWyh6qRTTCy4WuLMgwy6C/CqyONbCjLjLbXSxgVOKxHy2la
CN/YoRYBBCxGoKcqsheF707zvcG8J50AV3OiegnfsCZGjoXtXMzvfxqxODODH51TYI24Lp6E4Ree
F6JJr4svxomKDejMElCtI2EO5tZrAZu1g//0pZ88pC5q35uLiVXNOti/fg40nmmGc3rqa6nXoBB/
AGFL809dPLAkR4n7p6U1WfNuCvGgkWBW4ZgtIpmGrE9kyMBt2XmO1CE6u7VctdxVv+AFTb21LSXh
G7onVWrPZhfYNddhg6NMmxDxxfzRjzCDHNngkPqGXcvGjZdppAoOKpYEkmby4O6nzuhxtdjJk7Sf
UrzT2BY7gBIBw4e0PYIGdNHjKJapxZ/vLmynROefWizME7Dw7+PJOwYkWeEvB75NVJZxljjlipha
4UIUKCWQfAwK0xydD0M00YPSQPgYf5zuJuW0s0Oq3T4Ka1CIP4a235WM9XJeov1qS6/oDYcYDYtm
744dDG2Ilv4muJ66gzGi7YyGH51vqrRMm8z8GvMmHDXZRtMbO7h1ESfZkDJ0LIivXQ3DdcxdRxBd
xhELFq+0H9EIcj6xC+Z97gD7Vb6EKhAlii6oTLaI98nesMNiabeybMUVWj6PsHiNRwW9Kv+rwDJe
9kvfapkMNsBLR2rtWAyAB/PN9+Lk+DXREmGG+U5vs0iWMHauvGZsr19vUXH/0ZuuK1GXtrfJ9Ppe
LWN8VEkAB3YGccIY4oaWdTEfUP4AaoxUDxMlQAMX0mUP7VCHzy7ptPQgzf1wrwHaQEgjZWo1Rc/z
dQdeiAjNT5D2vNhyxwV+poMfJrb/KLP6ezFmY3pjgfLnnKqTEKE+Zt8i6PtnxEw3ec/N06Vrb3ft
Oid9YJnQK0wt62CJsQS1IGuQrVeUneBt6i+eOHoMHfr7tuPDSUfPD0titcUiveyawFtf67j3cvo2
mj/hgz4Lfm6qyjEdjIxoMrW0YvYJ3G1nhDNO0b6XlQujWzHQEOfI0/eC2LPKN9aiGkSKp3P6/1hA
qqns5mqt2Ytfx31EH0zxsew0BcJIKxTPqWWzZFStB+qgRNB6PtrG7rEWMrOqxiAYVgk9EcWyo8GT
wQVN3W674zAgTjyyYFlEIsmWZFcu+btgjG7nZF6gLXYkf/bCoooEsppgvf4Q3VTIqHtOhK9lvKnj
MSDFk843/sKqargH9zfMYTsI2BHvzzIq+hCu2nLWrgqsamHNybX+9HKvCxf7zaJ1874wc9A7DOXN
r+tUHV3dUWSAXS/ItlXr+7jzFn5+qMM6XUAv1Xtq+Eleos6hz4COt/TjqfAnk+Xlr/SthsdSMVc4
HZ+o8D9Iy955ijzp5+bFtUwyCdiUsE/HNC6TyHeXG6g0/qXK4pCk8mHkrSE2tg+22qsc7jswIjDS
YDi03uOFFlS3QmzpSG6JpuePIihNdYwcHqUBYNIznVtlWpzYqiOXnMHJ4QSRAtj3vtIWNQk9Tqgw
VmCN6j8qHvuVk7a/oLpafIN5IIUr9CGAgc7ZfTgBXAr6VoISGFazw/owQgSFBSbLKjhXzfSD9trU
ATW0yZ0YwlrWJfOsOoOGu/i5Ed/QZQlQ5rXpIppwfMPIdJmh/CVI/eUruKPJ6enEmxAGykNRmxBY
y8c/mbyh9RGfZSSr3j7Cygjcgb283K4NqRjveWft5pQip1MUdTUn3LMLMU8QFkEvYaAVzsery6Wg
OrczKHpT1mETTUDqNhZdAzminx8vDRXSivIKF47Ais9sGyMUxYkYNauMqKnW6Oxv4o+lT833B2WN
ByjPMTBXyvzmO0czmAJY8brkUE3UHf1RQ0ibR/cBngjxcuv51RquLGL045L/DbyzoKu8D4CIL0Ly
azLTDduSQlb2nyEIdiCnMKwzzc5QE4bUJDXzVRWKdnIcLWqcI0qEMy+wMFrV7IQmJx8YOnzObwBa
q0L7hqMK9tw2Igi/JH5MiSVucdVUYR0DEugw77b8noONC1HeSo76jXnpsbXVax8c5IvpgpEBly7r
3O2DMk+n6gToXiiP67cpK2RJgjGLBCtBT71CW9/ln2u2E3PYe4Jd9Cv+JR6cgn5u8yMi7XnfeyUX
OWRgzBSSjS3lF4xUO+sHFJaJRqXkkpCOj/WbOwbz9Aoy5IbEbjKmsQkY/wzMsvQxR7arV9JhtAc4
w6ml8iSkA2NjeG3k6xTrY+uHx1TClrTkW773NNPFDt8yLBCkhKU6sR5huRtfBScU8YUwytI3yfjc
z4csS22aRYUdqBT6NoQdR8lVJ+1L61Q+ocoxKlvYiVs4mb5EVWLQaHyuTqG7flU38BVFOntVJgOu
aS6Zm++GlBChMY7gSAZ84xFwstjLoTl8sCfDLDObGt+s3rCZdcG8dZsSe0A93eBcrwH8ZkGr7pIf
RlNKzr677KRolAghKXmKlmXtmcxCjiVMyMmCsDci4+LOIqGL2Fd0RtKYSeLXTNtr3SrlrE07BIiU
yVfQv9nkCN2eBt14Lks5kFxrfiwtzOw4wcdL3c1Sm1bgZhqek782cL+/EGnmZqD0UXvQP+F1LoB6
DsJTCUNF0OvgwvKRbIVSvwuoS3FvGVcOcctn6mpVnzz+IvG9AEDdJblRtmqDehJEfwrgQ/wvrKbQ
5+Nb6zuh56/8NQK4LPsvINRQuawpzoncPeu0+3AYjm+lERAyGFFh+pByCWvFhIFdDcBa6dkg9STh
OtmIlmMRfC1TShcWa6lhtzGOTiCr1Vl43VCQN5LJhVkBYaCQAhCbw8Kp4I0KHKcS+xYzLW/HylkZ
BZuYNetsrUTeFCQG+/VOuEhu2cfMoCA+gN/Sltum/09uS/WGDd3QpR+Em9cbLE89TPLDWT2angEN
dIh/443JgNyp34mwe8rdFeWRX0YusMpOBzFbj0nbgAx9Y0mpPZy/f61igFDmfJ1WPVMmQ7320VTH
bRL5E4xkkmHRnpN93Q75RXxHjCNVEriqXQGUZM/ZS4cT95eS42OQNzXyqiEG5x8y7RZcKWGmC5rr
HRHN6jpOwzUgtwAg35nWpZ43Bvfg4SexDKApPgLxLFBOM0Fd1YtATgNpoXW50UaHyhsBBRs8XRxk
BDV4Zfd5g5kdrTwQxsJxiPrEeQnmLWKQe7RHfDfFEoSWbs9BD/Yg0ReIjODavZ64Ij8YBVHwNola
5M0NcWEDQUEXrCgPT5wkOn950n5wLqQC+L4PjlH4SrtM2trOfJI67EfzOnDDNA+krUpmfreRkCgH
PsZ9CZ+XBg4/xHXetWn8QDgS4rTpLl6RnQhTzoZikd8eSeTXnhBnpVNUyBUyLIzoYpVb6QJVUAER
vydnkCaiPYYDkRII28DodynNpQfitmdznQ/YVj8/b51mVMSDMWxMyy8JK+dGhbiehdGjFaOJRh13
fDMaDpFvpGB4zROp+FKf16XlvqMF+xT46wDvx7DKF41ZaFCcpaizJi7tu0xew5Xp6G5inag/VpdV
H7xyPpS7UptOzZRsbgeXOXToPYl+OB3XTeAE3QeRt+aaGgz4KT9w9Go5OGsTF4+3v2V2No3G76B5
SLf1HlA4qBwwn+034l8KpKoXJpLuK573mXd7dN3K8/MPK4fzrCu9elq5hK4yRnxAUsJUFuEMcFFR
89LrBNcWDnOqEfkdrCU3kDTWcwbS0bQY2e9Ec6UZkWrksLxjzS5hGV7Sa6qsGtRQh5Mdeye6bt0N
dAnVkzjFDXjwvimwIwKeh7JWUS3GqZiIWhKTV53Bc/S63kw126KxtbYysaqzH0R0f8I5yMT4qsin
lwAeSqo/BM3dtauJSSPNPUROf+f2+zYs2r/01vnrfDQnm9+8cLWyJWznafg/NfcswTk4VZ/gzZrE
ulNSHAiz8ZK7oG2pOdodE+oSsUiOj/kU86c3OvTx0jmgx+uf9zBY7A+faVT+jhp98iP5QM8Jsf2f
r+BkDMuQ+m+HrTeOZHNYTStWT+cpO0GksxG7+dEc7l2lGlgHV9MT41kNXgSPssjU/mJ6JamOmYm8
paxNa6TjsIoao6Jl0yzfOg1fKX7Y7NoeZ9rfnStHFQmWa6/J00kJ3Xt2OznoQQAn8wSCOYaaiM/e
picAqn5qgATC3VTwmdV9Gh4eCC6EpATCHT6zj3fPVnKGUUePZhLZSjX8STAIgQlKDPfuMjt79o0p
TbqKWVzMzzhoZkreW7ls7a5n1gSyf8ntkCfXv++1/gNJwIiPwFP9241cLu15U9+Yvrcs7AQFYw39
Anhd2SNeJ+Nh/lCJuylnXWRFdIHCaHIm1jpYvdrHiwmR6F/ReFVj3g+FdLEt/d+lMYwnr0ORHXi0
8WwWc5goK6Z+Z/IUSkPGwBIipMVev1lf6/sm1PR3lcjdXv53TtXwVOvoRrz4eIKZsjPL0Sk+nXVi
iZc0LP0fSD7BYymmE6+JIxkGf9li7zBXXeWpe9dajOlPV4FrZM0k9fWO4cnz7ypLf7x2yc7uLAeR
Hxm/xWKU3njLGFRqKq4ofrJcTJm4uriSTd1BIj/yo3nqGK7T5Lq+rlWiioz4qoPR1SdFfCj4aCf9
SwDVdiqR5G6sRcz3nAi2nRnsNBQSancRcBeslaZC3oN3bBLzJwyZ3di20qmwzbtsTM0dqo4mfXKM
/nNODFl1wD+cxmJ8n37o/Skg7/GxzHPEVjbjcQoWhO2XRhUUIXJAJl2oN2JoRacikmM2lENNTdQm
Zeq56uWLCk6uV7x0jrQWHtbAtpgTqlg1I40sfZnHoXCfJJTcxps9Ze/6kMX80nQ13l5C85X6QHm6
PqJkPBfr4KnhwLNBoaWMskj683hYj4CJr/ZW2a4DifkeN6TATpU3MTMsgAQd7+4vFUY0Iopg2hcK
1IH+Ilif2Rbb+yzqcMGbm/yh873T15xQqzwroqUFrsFHzjuKgFTM4GZxU9HIptsjQIhFZMtmoA31
o3WdMvyxb6+QlpC+iGCyUs6UTO3RwxXbWT9VaCfRc8In1Fq5wtkeK7T7lZ14nBrwCb1P+wMdDa7P
FfClITOgXTGEJGZT/n7rYU8O90yDnCGypkckWZgrRsYipgevfbIA6FkQmiZwwb3I9hMe+yABaey4
/qkfR6129yGBnDaW9ni6LxFXpCXlol2cfLPGSsVWcAoX1GlAunEW2x2e1m/qHibHeWLVOV+0nqQ+
VwWong1tJloXEulDNHkoxy9e7Fcq7LZx9Ot6PMjmsXIWz8W6NXiQQBxEDNAO7EuSo3Btpcb8s1BH
Rjs8vbYma6gYpV4t4qyZrj/fM7cyncP8XUE2HihQOuPuNM0LK+NB2LMjfRCJXIz4D2an3WC4pEUM
yBEydMUN8YDzzqUTnTRerEcFyTekYWTK4Ax7+xyTN2vbNvWokE+tBenV+gBfNyYqhdOcaGEwMqUQ
8MSy9XMOwon6NYYEPEaJPNJ7mxFpvxt4OexlgwhT2hUrbOLGXhbxrqDJjhJPAJN0zuNwXYH2jDSR
51sTWO2BDmk0+yAth5bXdjo8ZXFSK2R4m5Fj9Q7wl7l7IHA5jTjI55Fk0zU2/v5ZJX1W/TGNKB6b
DB5ufYsQPfAb60NPzCt00+t832CkTHISqUULZ1fNkiMLoIRXdvRNu2TmfxVAs6za6ImobzpAoW9A
zpM9zoITwkFdLi3AP+rM0NAca13dS5l2nSuWAofWomfVoukoWowYALs+CpT2zmSwrXTKgnrJBtJk
NZZ5myCcTgcdNYR0mX+FjSUtOQIGBFurfu+048Xq+M+5NOVZE7fq+KZIJR95ABArRnFlJg/LQszv
1pYViKzCWSwlogkc20eMEOi1v6+iJzv2rY2Q9fqe3i62HbQTFEvVCBzRAsIK/GJqtwq2QDzlj6o1
ZEhHcBHVWTS6bQMtSZ3W+yewx73f7KkVBU0KmRKNfN4+5SU+K5UI9IagGTXqhEf4liy1Pjhhv/SY
C6xrR4yaHTjH4PnZJnrklPsEoVLS2lilKeIz2g0sUS17+BWRgOqGg45L+hhUzrYdKMkmDEyxTR4z
LSZNUcQdlWlgljLIL5oAyJx+YliYjaxoQ46KbAmaUVQFDWl5YrcaZ+vcLHgsGExitC831SPvefuV
NUAvjD9nYNpa7bUcW5LRd6oE/6UO13lfRiv6dpfRs1lhzUA1GXIktBA1vXWgYevX5N8H14DEf8dt
0leUxuaJpuppZYDL23EdxopQFCx0wNJWgkVQgQ4zQSkP7pL8HyoGqQu7OtOPsiN3LbmYBmXKIAQ1
ChjGByGq0p+X9tLfAny7J3z3LsiQFyUiEuJCOiKqHkQWX9hDkbrxjQZmFmhBm3cNxDhpF27e4KBi
/mbn6hHOGHxpWcMaNuBdS6OVLNqZlKnbuBnYzNQ5ruRdARLkBywu2H+wJbOJeuLsf28sL+y702F4
Lf9jbDDzkHkPhLP3cAzE7QY8eXxpYuiyXgZE1NFXGr/MYND+nzWsY5Z9lHeCAzHlR8n+SyMpVeep
QssByBvhp1jmXM03173yCScDMWml6quZ1D25Q10LE8n0VUadlHQ0MNDUmjy54viX67fYGEDQll/d
34XEysmwx55xLefTUUfymETM+FyAVcuSEBTC5a4qKHtGyxCTIttE1ACduEtq0wp+/ZkSK1HJCLB3
REmpEvswtEQeiNGXvtuIYujOfNAvWpN3QX5Px+8u3Axfhnzp3qwpSAozbwtrAznDHJ4S6Esq3a+6
rfN7zWlB6RrFcoj3e4KahHKRJl60p2qSb3WiMlfz9IEpIXye1BrlKDNFOSgpoejGS2Xgga+WMhM0
QDZLFJ8SefGyf1JwXVTBlxub5tyK0E/8PDBTR0zVPjATWjIMHhj+Q1G/mJwkgf7x04LC30k6phn1
csZrRp3Uc8bqANTjOFtZJfK5WQrNqbfx3SBcoCfhYy48LJZTDsovIMVKyjFJ27pqEtbAdvaUHbAe
mmsPlg7OJzq5J3J58ex7fPerd6HXf7QE0/2HR3ujw7kKdIFfGYDfq0mDlJLe/DKx5WMsjoYPqcNX
sDPAW3pHcqigXEnJEgM6v/YGDfEJO/0oRjBMzxLNPowe9IOM6ETZZH+yGGyzMEVc444tja+dj2Sl
DUJWdcDuq/Fu34ViXsRoQuFs7h0Zg0duJrkOZRvDaX661IojrhRXzUjG/TIYs4MfmfsZ3+QsTiM1
x0ykb50yPdY6PqSzxm6hEtxYDUoO6byReCUHm5bIMNpt1UpEg5RgSNvnIz6YsS3xK+q6jPOw5DWn
eCGlZ5s6CVkJezGCa2Q/9pbaxL/V2JoCmvJaVuZLnQosA+LIye7p7MYpyc0BIoyX5DgEHN7ydJtT
CTLa/F+fR2llamJn+CbECFjHTmHvoelnVwfHMlw/piLwGyHaWtlg0BEt7idbHB0cVxyNuPzH7H32
/GbY50GorNE/Pg4pebBwirHIuUuIWyntqaYFAseTt+mOWf5IFvlpVHcbUSITTGHB4slhB0TCWKQU
mayOJuMxGIECCSVbHN6I1ohQRlpiIMBKNOfsDs/W61uSd3mFZJLSto7xjQjCJ/VHoPVcPE7e2iQ1
oGbB3QwqSyWlCn0euI1xkG5HoAQHGntrMdV+a4ix4vnXrBZy4LrSwd4N12/EoosfiknLGjCOvqYn
zEsJtrzynadLX2Ji2NTMjFMZjgQ1I0Jd3vaDpICSgg+4h99OeIL46/xNDXZKgenHm0uWKpEvfMak
hKK4ByKHAclgM/Kzig3ijhsEtgTXCiEBTG3y4HeYtud/dRUdJ29nw3yC3TA/c1YCYqahiNPPWYE+
6URDOSJnTYRmknUEyW97QaQuGKOrvn4MmZ1amm1o+g4E48Ss7+GV/sAH/Dc52XK3vNK0VkngkE8p
lRkIxtZrMxqyGqgo4WSmClhSjYX68M+RUdXDk0oJ8M4DtTTNtMShN+WEQOecFOzNTQBKMQzxRjI1
UVWDsb8Yg8L1mP0ZHGdi9UeTGgsYN2IHiInreSNhTVB5xE2ie8RtvuzXfWPB/B/GnvtJvh0cqP2Q
vNqB1f4IcdLippeWfTNyh2byI88OgV87SHOhL9MtcgnaJn2tNTXZezfgiwtpKWI+Z5yY4uQTT+Oc
887/GRgeZwS4/54ucSEuSvNyEYfxfkP2GEhsUOmdT9iC+cMSQGhvsyjaWD/bdc7WCMYzxspeDM2S
VGaSJ90VX7N3l/X22mZ/v7WW3xgmqzcQY3p+pG8BR33R7cW7i+S+UENezPKtvA9NMjEu5IoMRgOx
gxFMGFM4+pxKleNT2veeeE52Nh1GO3GisG02W6CMlgytLdehj3CtFIaIUf6VEcLinHkxjzHag0L3
om4VEcERlHDPai/o9jPAREm8Jku8vPEVlyAziIfP5kt3nezMKEkEcF0KJdJp1K28wx+6j72jbb8l
RV1lTVCv1XlXxsYuFKZGzHFDuQJ3UTv/QpIY/OL47840TviHJJDQlyxkOGAmeRhB2rA5K+SuzaPP
Bf6mN4xp1SOJ8XixWTAtSoVM0wj9mJ6IHjjGZre0ymBDtIXyg/iobrcCrMqGYGnhpjfiPSleSTXx
DZvtWL0KJZzN4uKlSMZAZP69zG3rMI0k78l61JdDbWYc/R5S1kW5cxK7HxbboXHhTNp++ak7btf6
yh/MSlV2YM0+peLluCi3JoDkEvNkVulU2ALNvepgSvSDApr3owP+wmTePg0d8q+GfQw7dHn3ZoVS
riQhD2L4d+++hujC+iwD+mCA57otAeydeS95HhMnUUu7j2R87T7rpK/leiUvzndToz7Fl2eKubjB
cYQvpHXJ+IdOHp96lY1o0GsPRsUVUK79wjQs4vKKN1etY8i30gaIBPeB/QfJiafEgs0HUrlw6ZiT
5eb4F1EshqWC5EXxx/ioFMoNvsnrB32U7WoXRHJSpbOq2n335bvHc1f6E4rP2R2XLCagKqzVkI9Y
7Mn6EQgY887+t2FbAthdA1lAyNOVKMvLD/AKDhKzIpNyhcQSCcWdEJv0NsdafNKvNdQ6fTlMXPvg
+zequpbp6kC3BONmYuceM7FE2h4TLIcJooO4o4eXwkD59yTf3/e/3a9a83BahMrp8soGYlT+ke4b
T2/kje+Fgqsaw7kBNjWNhAYry/PSjoBj8ASFXM8x3VR/bixdJ/bRL+/ZRetegKI6cs6zlbhtxyZ4
gSwf43PoWpiDUWPz0wBZs+xnDJ6iQ0G+T0mdDiHKkBrsFD7336c+gApAfOruF0+OMwhtcY2dphtD
sUe1JG5cEnwQgUAVEGSedL/WcX5YbZ2b/fgPfM+k6+mdhMBRpxEtLog3hWieaIGyZcoeJZHzNm9S
wABlaL3Ma3gHi005IBCIvRTDEsQDLi7iJCdNAEsbSi6WfKrMAEShM5TIGY+VnYkNcQDB4n1BKSsy
JM8saSx4oB0MnUlB4Z6lZRqPrGP8rQfxJveRQFwg6DmEoLv5R3QzGwIxh1FTDKoU+QG98//rvPac
nil8VnvDZw3EGgaeqlHTxhwW43PlQki0rtvyHOsA4pnJFl7OL2E/oFKslXZO91eStYx4Q4E7kmOJ
SOpzGZquYkzSJawd4YoEjwWA7MwLkxzJlNMsLbCMc++r5dT7U7GHBjDp0QQCoROS6ExqbKWtjthf
VxZvGFmwhNgQt1FhxgD1yk10P6oBiuuUTTRTNfvfJziH+DqSDZnS52SszUGRC0VKEfa3wcDbJuJc
Lz4pOLT8BjEFdB6vXVlFp1QLJnLzU4d+eI7yvMEC7Em86XPV28YkJzL7HCyC4hmP48K84QB2Aks+
q1VX8lRhOAviDeNAH/jeWz3NvnfPNS6CFWJOkgsM5xCXOt+N47fSzit945GT6NRxnqKFIvbK5lFj
hmbQoALO/tsEB1oB3d8+5Q5LjsmYuk1h1sCuTtZLyfmgvUgmMMrd12anlUCFhmdp+jB+V3b09uz0
hqkzJyCMHXbFQEFiGpTZZTtplZbLZWBgFaNtNblXHNtYGAZD4sBW0HMjQRlMOoA72E9OAXIRb0Qb
mOWcSLsEyGR2FUyEnwO24Ybz5utvPW4qs3v8rcN2Fo4+DLrd4cQ4JEfLucESkgkBMdFPa7gR+LXf
Hm3ETPs34t/Syj9bX7FCHnReUduMnAXltJOtVZCmfncgOP0AAVB1HhsQEGKBK14jEW/ySViTExjS
3StMC7wfe3JfEVVE4fD79pxWBXWcTJ1/TLYsqqjCyEu2pv9rfEurcxoI0wfNYW2RMqdCdQmY/4GT
8CVuuLceSvlMj7YB85/D2oJ4vSBU6KcAVOEmCQ6z+LZXuzV7Q1Z35Qbcx+6y2nY2PLQzgmGltuvz
fWh64Q6fuplTHl7frbcKM4/+nYYIGAeiW285ry4dRkdizGfkrYm15NFvithJd/Eewbszgc7IOBxr
mQVux17+WUAE6tp0NLkm60Llz+Jz2YTnPaQlAthTx42gcIwAyD8k10NyaQUrqsK6jI7RStumaF7+
sB8BTCr5u0iNF2su0PpjN68/xc5vs/rEtEQL9RO0c1CQzFtpPEIqVGcOel19hhjh/58SmWRWZo7/
A18USTMxJu9sIoMS1I0tnuj0RNaDl5/X3PPg8Q08KBSwfw2rZxZmh1JTSUKrGEAw65TytzGwv9P4
jtOnVcnIDyKLjytNv3yNYZDr2BACVZcv+pKW96DIUEdnjPnoO4A045d0jBOJTRQIvccdTaEUheZO
Q+pwkHeJDDrUxzHnAQD2evNfBER/WQaRacuSU/6YscT2yIoezlmxJM5I2an7fJF/eOeJYmHijnot
qrdAeps40WyIChAs/c/blDk9P27jirdf3Wx7uK3X+axfHX8M3zf6OysLuun9jqT+NzzAb/f5UsbI
1q8ha9ntGXrZ3uCHgKvEFXgYGfiOvdgWUA19nxibA7R9efur4oqADYlyw59qQtE6UWUGDyNuOAEK
PJllJGw6wbhWjo3GpRg5Wpltfm4KpTuSIbIFlRz4E2obY9SEiFjamltzU+bXg07sfF5wuyCmwcvT
6yPsn3Ho0HxU6v360xghRJZJfDyouuTga9Qi8oU34/pPwnopMwxc16JpixmuRTrAUB7azMgFFVev
JuWC2NpUzgtUjii1xR6+VUT1FL0c0OjcPL7lOMKy59CgWWbJtYlQGmmR7BfbSIsR+sXtccCJjaZy
S256BH9D78lMB67goEytOC3NTlkhscgvw2v0XxZrHMgVMizPTnylsG+RdRI6+SlvjGu0DuZKRScX
5bC+c8srrggDXcFmTBOvU5lXuytpE9DRzH0ySmOXeRNk8NcxzDnbmhhpmzJ97hinRfWqOWGP1i0j
yY5Xb+vUXT9OHF09er5s1TLcbh+qqhaRaerdqmLnnf3ZTe4UosZ1j47ssj/WrjkGOxUNCld/CDeT
gwwy4RgkuMz7/Z3ZC5ubfsupwb5iUFiJjC/VrjRd1CYYoK3m0Lr3+E3IOENKP4cBUI5/ZVqdIKsl
gdJW0QeozO9pi3Ow41Q2CXnlNrtufpxRyVsKFU+KkeLrL/jiqGQROFGi4YhXCFKhpFXDX+zXEqyH
J/zEb17I69mylTrPp3u0g2/F2bJM6lJlRNp0GaUNM0fiaBNC0tnY3Nth3lA+i1DzG3iNrghkXBbW
ypJGrYHMWh4L5oLVP/31iz8q1WUTZ3BTGxD0FMCqFNUz+X1xujzVh92r/TizedP24kdF6Er+F/z7
UFyUmu1oirgVMu8LfcM//LDfKq0aaTh/J61aGEvm34Zqqwy6wTcKXB11xN64iotTJosbvS3YXVvH
Ef4gYFLuZQx9WyyN7AdBfpVymuoo/EdJBrLwbMMpP9zz423OqOWo3AxCkOsHIugs6wmV4R4WOlHs
yj9VwoOPY9CfZ0m2mhYiumnj3Wb/IXRY0YsBewx0iiFxC4Mwe2X38D6OcxOFr25cQM0Tb0gzZBSJ
xva1AlNwQM0NvKF0h1RG1yFoMTC2ZGY+TWt2lYzZQMO8Ch6RZG77b1KCypnxKOjo/fi0R54bQvME
07fgmhmMYw75PTXnlrYOuJmhN8zFuSWzxK/KrbiE9e5l0cGwXiaEWJYVHhQc5W03Y87Wc05vFsnG
RVr3xgOKSPBZNVH+WA01O/Z2uGWqcv4nOG5BZ8bI1Ps+AmV77AIvDhLVGb4CzfCR+HuE6+DUpp+W
KkhQnEF8/bxONA7g/QiA+Pjs0Zvl965lxE8jelmiTrXcrPV/1smxYIDVA7a9yBk0DmVrcGJerRkb
yKA6stbvbW1Opap2vQBoj3pcR986j8kET8VMU2joaKUGX3Qulfb/q4IW5Li3QL4DXopYrxv+zP2A
oxATM5deDhy6VCmVreO1ic5iBd7XD2lOiv+21xqMRkwDKnk1QU0wAODFFabXCN/aPhY5bFExT6p7
UGXxqzDiDAjxCB70NcqcVRv+HzVYimzXJJ6eddKDI/7C4CvXaFVFRS8lZJi6my7HbI6j6KArbzO9
1yqTQYU3XJaS/kaNqQC7sQ3Q/BpHUcunvhtbwH+MMFROTK03gh23fBPmxmYCkisEG6BJs4NJDTZE
WG8GdtH3ZaISaaioeN5vf5IPLZVuo8D1XyEQUmEsdKxf+CAudly5i1MEUZVCCJ4AbQM4UuIK3G+5
3j3vrtIHfn4Pvm5fuUCvCgZTLXkMs2Blgi3VKmI3bB7tNexVzue9XAWzxPK4ZK04qYPaGZianz10
w5bVqRc2EALtg1aNu26pm42nljelEkkZ4YLYRXh4sR6E36+PlSifgFh2jKqe7wtwzJpaRpLGxL2A
7RXFvD4g2bcE8oa9A1hwn1eluf7nICBYbRlyUHl/+xOKBx7clE+ckrzkavWT2PcidBCteN3apgoo
YLWZJBJunfwq1lQaUoZBTO6Be4z5mBtUrmo7uF1xpnD0j6a2ujVjmajAELziJTUxhVGurcRVoqeK
BTMX59zU+akRpWBijqhgJ36C8UtMuWhD4yWzjSE03T3Df274fcsW78YcH4F2hwPFLtckEyRzbUBk
lvPx9Z87/wJ56tHaNJTbzbeggYhBfpcsvKOy8sgkhtXrW8djfDhVDfN7RozmBocihn8b4u26rmqf
wjnakUv22lis7LOnpdyo8v6Rdacu2K8Q5GKTCA4pxDOPjJXjNGGXPnlLbW/FRPthF201Z2knGFAr
jShOkOqvhG/7CKsXEPoo+nDdZNJt4Jo0YZhg8uVxfP1fYp5ecv4IQtascRmiT1eRByY6j30XeSW2
eqaZZOaiuR4ttSM8O0ULTEwUm/UcRl6TKbw3KkNhuRAGVJ3+BKuatOG55oiaBaOOJF7767hVsxiQ
MuM/a0E4wU7pjp1mupwFhFhXOWdQZBvvzVN/aEWAW08mEMOlojOfVajm/V+LIAw5LVcT7kHhR09s
W1aTP/9qJ8de0LdidLNgur4DN7Z264x5XnQ+rB9sPa91tEytEyaxJbKUWQJVsU7LOsqJXswblv/L
cSDY4UGSixg34uFb6DcIeOvll07wtAmiNHtWKaIimRN9lHqaevfKf/++GQvpGp5YJZfxb2OpEP/+
KEMsXCD4IrPvRBXwUE2rZzxtMEELb6NwCCHg6eFac6UYnFw+7SBc3bhii6dLkyf5L5LZQ4KUR8zH
nATvOZSO/3jra1PxDxklFifpWaqbrkkmY83XnijM9lT8+lCvnsuPiMsBQakvFTnpIyevZHOulK6t
6eiHztTPBpHJb5IGjI2orHqv8y6xBFfJ1ZCSIgLUV+zxBidvKUynfgvkecSHnnpAbETS/jjRqp1f
VEePpwKJVGV2mITkrqZxQ6V8tGv0txv9bzMGauvGXueGCWveyC3vdR6gmrb7Hop4A55m/7tZH5Pt
hCqsRMCEcwqlZXLw8dK/9gKhUE+/UyRwZs9XF845Z93awgRPKag1sntZnem5oswOFD44er6UOJ7s
05DKGzvttP/CKt240RjQ2l4r5r3UMaVgRTQapaBSslC452p+7m2eW+NgyGcnWvjhbmvdaTTXGjCJ
q4FpoVj237i+kr1V+L5/ivJySigi5VlHKlmZ9SUcR6mnR9p/9KLggwb0vCnCKpxrQDjhFlp/+YLS
pYC2PZABhg3VI45BP6zmnJoXYtrcjXY0Wm2weRVrU8pIi8jyBAUv58UWh6RWtVd56Bqzozm/QrWb
GguoBoQQBpKsHrevnC5Dvci9Cla2OBJFMMl9AOfoOrYuT76VHoI+VZhT6Q/Ipf2akshXW+TSbFuL
8oKBxfQxOlLmpUYoYXF3530uGg2obyN4erzLB34SqJYOsYycyv4P/H8nVwkMrm8wVTaoIN4YNR6X
Gp2EaF7k2wmTqiOVRrPDqIRBuvMYIjz9oMnXNqlc06yVqnU8IGYXqs3xZ1eJrkXS5ZXljinWSv1a
CnYDH9DQ733MW7Ae6MLD+EqlgVBr87KNcrp9Z3A5t/vB83H9Q4F8HHQqjqZ76U1MFk0EyeyJANam
gHmE9WfMoRMawrdBflGKFE6lO3uPO/CKF5wIdI9JYJd0xJFiTpnG+IK24yMKU4YHN5fEVx7sIG1F
XGikP1gGIOduTxtbxd6UwAlb/cwslKXvgW3smhhoqB/OTmYvQeWLTPCcYix21xMoEghT+FG2vNXq
7MhFXhgPjaJraajcm5dwYRI0tlUCCw7hhvIuVijmYZNuUZk2sK9VamlckGBPd/NDrzxvphFH2goY
+nlewor16fmOAF2BO7kKM8YwtjuTjojduOOn0hyD+ca/Bf1zMznV8HSYvu7Kcc9680Vhcf1CUxR2
hZq3m9IAACOQj8IQT+yS+bsgYvpX9bjbsc+1FQuAEHUbu0hAPMCgWfxdO24esQe27DesGh4cbdZ1
TP8ZNkgN8Ea+VlLitL6gnu4EryYpx+ctHwGzwBDuSj+YtlTZNccKZxTwipZTCJXInfwEZzLXh3XI
WWYrrX2n0FRR23pSyJGvGOzkvuasG/Dy+i5TFqhWgrzyeIAmVQ6Idc6XVc7tZhr94jkuCtmcllpF
EetqE8CyJBBauXXZBHWKd/bGrl/yBtwHjR2lPadkxnSoP+JAN8srHLCui6DdJWwDEuXostlN2tUh
iMosYrPSDxlgyhz11vY6kbDaCMjZqRbyDAujGryfjv75Aem0bwDzNnjThZWOSUQhJp0KT3uUcpYX
ID2s0ZQcMxPDo/u+c2MMXj8sosfZhMeu7+qhU00ixLJhy6HAqY6bbBinQQWxhR8OsnS/CDjTTheF
QDr8Ram3HritMg5NYWkadmFH0yGmd/ocIX8k4ZI0Zk44ddBn4g47dP2kDTAtrGe0BVqCUltD703p
/YcCOQV62uWEwJAPp0k7xkgdjvi1yIRter6Ohf7UmOHXj1Ab1gg2ucwncGrwSHEnx9NYZP6uqek/
HDKIch9SyHNX0N1QP9NVBIuE+ZtgEMCoFbLMMgJhRCS3WhlnKcVKGrTe/JLWn+IcWVbZtWBzkTrR
vxGUFdRLJZYzrWt7SqZ0QLjB1e+6jPrEMLzy7Hl1yx2fsjH5JHg8POb4qNEmn47FZLwNLGGuLDIC
3ex/gpfGFDrN+Y7lxizrSHJzdp75GIL5ZLuCO0Owo4i7yp0sJci4aSoX9D2dhoa/Jm6F7rUlC9Rn
At5g3CIieDJZuBzaIR96fkW6nfle4KIPXmrIC4PJBGVqWwi4tvou7ZZA9oJ8GcoWQ2R0uoCN3Dx7
lKViGQM3KRxYb8ZVbfCy8kUhdSYOSqYBpUjwS7/QTfZUjNfV3n0iZgoNmlQel2vQAwLraI94nkSz
Ivulgxynmdv48HiiD1K3U9Bgd1V3YCsu+UTAm9XoFsy2Oda0pxCNrPAwuaDIZx5iFV0Yp8oIfuSi
jmztdKBJKlryayWPWCtcfK1+YOvb1bsvk2s3MILC0GpHvB7QguAO3cJf05jDXan9NuZjqS6HDklk
q3psJgbEG7XyDub+Ja42SRUsH+FPMhThIVJZVW7saBehQAfUos/L8xQZMpG9lDet1mBRlkW1x85P
iZnu0Uqpic4UsY7Hx9EXEMt1MdN4q3bnrq+mSZl1rmOKWx68W41NwNKV/KEH2dA/KW/mHJieCTNl
olNNY75lea4EUihc+V4Ri1pr9vd2Y+Ic8npH822l+6w02ZHJe5k+mYZWS3Ekp247JHjukE+SIiE8
JbN+DkVlap/zGvsDVGaBFpXip7tauJ61QVS8lFsWy0nRrrDdwYn5cR0lLWIOU/lnr3TvuPnq/0rd
7fvfE+Kd5o2Q8e8CXgtN3nzArJoQEpNWvOVLzfgMRbtkHPvZJLp9Q88dYFQY5FfBNlcmNMAlgGcR
gJC/k7BK6FwtBfO33zc/Ch8DW4k0qSHo1Css54yF+3PJtLHySIrxYgqTfyB6Go/DVHq9jUOPS300
QLxsffaY41pIQJawt+LfdbwGbApTQg9jRCQLJrfURQCcXxoehLgaMiHDBoeeExpGlCk4u+v9lYrX
R6tkbQxvlvcy3YW7WOE1l13EUZUxFnJKCmrfzbmEQwTRDhEFXxctg8IKtwuhU6Pr4HzqkmQYG3I/
dKnmdIMVzyYjdFUcG9IMCDpvKRSPqs0KbxO6UO9sNEsoq0rlR/uOba868wZvtk5QPDB54Bu2GSZh
sIQfO3vIwW9FMrc8GFH12urk43pycSb1N1NDATlwtWUuy0amW/DKT0MNfcLDvaAuXaFloQpgJgYU
m50xkXYPJRditjP6NUeMrMGgHGYYRwtnqveu2P3mBgAl3ROUmS0K3Tz3qQwjwZwfNP61gnUzDTyC
RGe7puOM5XGpBuBSq+CMzAxN5VG4sswwFdyW8xoopxEWVraFLk3LlCTyU0bmw30fa/zXYdqyLfnh
JlKcj61JYQyXcOW/jaWF+/KvfLNwL8LEcU1yREVQF6F7dm3LwWP+P64ZclAdKC3eJOMzddTCS3Qm
rpNi6zJBn7WpYLkXrfbsvFdkAo5hiBdOfsue0jX3ZnEgqR6khA4Mi2PlqlKdhGmToZsn3J5dspFy
tqBB3N/zdeo99seHmc3LKV4aVyUGXZqVpeRPisJwSaa5VF+BBGx7za4XlVmPG5Ro6IGDvUkAQYrS
ft24k4X65geRQ88QvTs4icdbQCTQxzBmK3nbkYoQUwYkcjc7nKKR2VXj4SM2BfALQ4egFG0CrjTY
w1seYzWqlnkPDo3NmMjkWJ8c52nGWDJASxUgt5UzLdC+BoWrIi9t6ymxyEESusI7l/bVyeysB6cE
a5nzfNQ6ubx3x0P/jr4wuoqgJ7bzTBwCkkExsYnhcGpjHU0K2gBBHtDnSM41pHYBzolmW2c87TR4
IZKyq7YP37+eB3lkIWtpiRhYBG+q4+16I3VjJKb8oUfpDsFmCjlvCyXqfSZL66A7FkOnUs2sJRhu
fErj1+J96U2iVF/RRmxVnohVyNvQ7zjoOVQssobvJldjvajltNlrePhzIO8R6maRopi+gH7Z+Hca
TTcKIFcEf2EauYitE/vL1tZ1bKFp8kvCWpI5/p6/0vEKpHhlqgAYWM+e/Pbgr27Z3TRMkgKYanIy
VLtul2qXkXJvk0j8SKgjh624Hk1huY1bgPZqS7VHC0rkKk8ScQaqW5Cz+fcjQcwRWPZT3ktRNlT5
O8CTVtak+ycS6LOlL4xU4wiStKWZ0e8Un4ed5OA7zfJWzDTDLVkP/O/x5H/Twdu2ZkOCvpfgXE3M
dvD5d6VBNKpQ+gsNuMr4CdfyjdakVKSaJTleMI92NXOJCUB0K+EWsw7C40/uEhkww7QSCDqMJP1N
ZB8Un/wz1yM2cJH0+49Z3+VFDulNFro0+GDxoEHFf1kw3pIwkK2B7+cA2imTVD2aVG7NhcVC6KrV
qT6yDrUBiFx+u2UOq24gcvPCb9gbusYLII14RQLoDgA8Qah42+baoU0TX1GqcNtzUexmshEAquBy
ugNBbY5H/GjnOInJ6Ry0WYocIR32al1jzLA9By/j/Y8RbE+RLMch0YO+OqXllSBdLgCZALzEO3sL
2w+DiwtZQ1yPW2WdQWd67qquEUKHlSOtSnGftyhLGKesiN/e8Qmn44Z+1OMLkJ788PteiDaeU868
V+EteGAYFmtGwgVXwbHKTBbnuEcUC4//EjnYCcol2w3HZWnz+Dj9WYsRpscC+bg8E/XkYwyLnnS9
5hrh/F8XU+6oWpCQ59xVvaGhy5evxhTfeC2k+Tk5CMeEGobxV9wx3frccrCKiWBS2JVntzhxlQ+T
FIJZl/kjRIOywbCwm4RqotwadgFr+rcTAdsZ8ChBmAzi2w34hmG2OaiatwZjRvUI8LaNtSSKv/82
/fUmeMnUx9PI3HgQ7gfTVmUsEOLMH9Khtm+XZQ382vDuHFEZYROYGHdkBJm4+6KCSNyJ8pWt4mB3
iG8fRhK+7/TWc+w8vbRNWO+UxTgD0KKkdDIc2isSkAlCwXZnX1zH26gTsrWKIrJ3wXqa4ppTfIXh
KzKR3UZkpH4y/CdzU87XfGMW9WZ9bfRAD+RY6n06GLwOeK8SPxSSftMhAyFm1U243rXh4JLVGBAW
pqPegM+/5tN70LAsb8rDCOOgieigukICZeUwkHl79+J43NdqW8jTDRQZLaB/uoqLIY3GV2VLLI+8
FgL/1ZrWxMl95nqqbui4hWg6i89ARWmo/tM1pkxn7Ytp5lkwPcI7sIrnjVbHH22KnBcw07o0T4NB
4nUiFYFYjyurF9r28pQgVsHxjGOvzv0U3siSRv110lxa/XtTla2x4jtOgx0WtoHd+RVOxDx543lH
88/sU/cQpTjaC2ijHxcdQYMviBqB6Z/Ozunbwqta4qGUpOEhJKbLNttDD5vB860b5+/M+C7vOlUz
WKn6Nbh1f9+WUvqouIPrPlIGmaCPV1vBarNP1Ylmc2i0G03HjT9OJ05WET+S798rDNyHqrToTvY+
lUQMSILuUTpjBAME7ytGdq/LVoytyjjgo+2SWbF8iXBplLKrkbQus6zFhrCNTphye+s3L/fAMSYJ
GzdQgJLuKStY64Q7K4ZYFP1gEviTnuxXpqJEjuLQCiph6jz7mesPR2zG8dz5f37CojUorVEdjTmA
P1XbZzAP/0STS10URTs/CjfXqfDLswM8AMzgz+4G1ll2/h0CQC8VK2CLJtf3wkbRcwsdpZTlf0TT
mZge4zums0s037Oju6gdMQe3QbeqYjbYlgH9LBP+tt/JlQ0MQLohp7g7FDo1ZP7UH561Tdae009A
wQCqjU99slQ5yIEsIK8CtV56RkOdWerHddov47JWv+HVD2Ekq1B4rqcHnI8Mfo5fNofjMtCqLRql
wD46cy1Y2PimTwDBjTuuUdu5R9qsO9qCmmZ683jmr1uPWkv0VUly78ix+C0sDhiUwfNd4OmpIN3J
55oHXzJsAZTskYNDC39s9t+irqIZGn8267irc7k+yrDRdY2r8HdFl2gIaPONhmZHtz2j/Fkilsho
eRIv0rO5egsJ1N/9MELzFr2WOyOfHJxL2LB2kSqZnY3m2KesAbvNZLfWX5VSwFC5SzlmYqW3UBp1
Gdj+h+ZTajlGX717q1/kgKt5o4KAFUzt2GBA8Ov4o+KTEvUH4VZVxTMXfPKFyAEDRZ1hkXzbekKV
I+NI7qYonYzMH7+rY5Fy2hHeqmvm2497vunQ0riSk4ILIiHvQmlfoFYeAqkGIBcLUj0BCeK8S5s/
bFn+L6tg3mqFpHe6vWHVDAnkR8LLvkGH4BIGhXhoDt0RRgOduETOewQw/JZBHUBnf6VYN3tDNSmE
e/S0aBJO7bKvl23ojPw28IOUWAxjTP1hld+qHeyNYSLLpIPpYZf/NcUAVrd/6b++h92N2GhpE+38
G3C0VeuIh6KHegbSaKCoWE6392jxN9Q2AfFAMSlbwwIFWHZzBZ+NdlwRx8WZHnd1YtK6xNpGwdLH
UKx+iWvlsxrnSvf9VHIxUhrCf7NLwYbpDpTLCXVXhSvt3S95OWstkJo8wbCzdNtbihe0eZgDAdQu
vCCnoVIx5vyYU+A5swu9nB0jRqTQ8kHNICMEhX/wM6JErejEG0gA2ytlZDVbxylYQFUI7X0pk+Ce
vErJLsH/TKiZszTKdDs9vVNM+Bq7/NDdfYstb3cGh2Ka9K1y3atJmEJbYtNBhhigqctuVl5iuky8
euMDc5Cn8LSJVn7vcnEBO/tOr62+x/KY4/dDKjc47+uHZwTxMYTP7wA0p2pFCKZKxuhOeiQ7jlq0
uSnNFzTpNM8wUCXK052x+fZ6Tg4boR1DIQgb6mO6un/rXDip+VXA+9JWVvyJo57xUoiY23i8y727
JDnwYsbqOS2U+uImCLPDusMRn5AY90aX6qbj1AJq2ehX4Zf0s+6TRiJ7ZD/PxP4ZtWiSqzFqJW8H
1uji2l6ykhNtN9dtfHOq/WBYFCVfL7TIe/QzrUwdKcoP2wg67HY5PuND+J0W0Yavzh9Q2BownUPq
uIwvg0P9MAvvDw7CvB1v2jHkg8zjKZmPS68sPbnJCga2l6iNUzsGFd7ZsWSQb5Mld6uoscBdDX5j
kEZWKoWYvefzTAlDZ37G7fAEbfsLpIphMUwx/9a3gIDnB0Jxcc7jA0WZQkdJIkwbEfWJYfONCEuu
fpOBJef3e5ru83FCZck+1/KoBQ2J5jl3y3y5XBN/uNdkpIKE6xLNYjF9Oyi9woO07N07Fa8MzEjq
jLRjkobUQ/w84ohQ81gzk8j9c2CrzfT5Cc/hM2N6xK1YAze4Ia7wXmMbIp2o7iTKqhDJuyi4q82s
bHuCJBIvqxlGo28qA4DqZdVJd0lZfqsH6GbipOnPFbd9GXhbNYRfuuyqv6IeXSoe3VcRGKzs1GjN
IDXtHHx6xaxNQA3rjV3icosAW5vbpA7njPUk4vH6z+ai0FhP3qcyKbVICsOWpLJEE/6t43VO4T5z
a1R9FT5aetDMwQeTucx+Rpk7f7pJTBG+eduftDQEDNeiWf0ig9PAUuCWD6jN8QTlvzb0A68VB/Tl
zKZ6xEuh6Gsp2dYE+h/HHGtC2pzHIUoP3g2oBINlftuIaHhnq3wnDxaFYmTvvWFgEL8PbyNJ1Xn2
55LHlpHOHPI0zgZ/QzP/MR+/sOFwuY1zJm3FkZyFjRO5hnx9qNyea0T8OqNQgmr84qBqNLuXayPL
gJCdJEnWdKrLH+h6Fj+To3yGMEufDA52Dm32K1MSuTEnXa+6jupyhSX0aBeHGf0HFolQACS5mijI
fQq2a9YH0uVoxA5b5ty5aDpTmWMU8r1RcLsh1C6UwnM7yzJxe+eHyllBjKYzVzaG7C8D4BZPj5/c
I88mdMzb8ispAG6o2n3BzLJgjX1Lt3rmrVEFL+rbN3Uuwqt1kgQW4WOj9yqnaWaGsn8R1kjylUY5
VHbCQwI+zkWma9ySUy5vsp4oNQJpJmL/XpB4TjL4qoQomcC+JbEvRciWSnmKObVPH5MZC4D0stBJ
cZ6YXEePnovMYUz8PaDdi+dL7tZrIMImEBXjmTbeNlvzGAAeekxn3/ZLeMitiWJ632JDs9LegFzV
Vwr9NkheH/3LEEXfFIozXVrbeKap/q5WZ7P5oCkko5cCWnIciLQzvYfB1J8u2/wgi3R/glhqkRcZ
TIMv9j5jQJvagk2uR2GE2JYast2HB2MxflirY/KijryxRcSUCmJqi1woE8i77ylP1FQ24TyLjctO
nn3cxk7MCxvF88NTBuAasP85dmov7DbtdZdl9NW3igxXj7qNgUFQg46IgW3QVIHml5LAX95lALHm
iFtUqRnWdfnGEZrwLHpPDAiJwXon0T60n65PWQ8tQagZaFBGa8U2BDVrvssbuzfLxP8p/nRJR0mt
BlcftD4N2jd/Mg727uWbD+2v3a84D05d/8Or4BaKoV7t9gLm2rXFI4533R4Bl3bKJ3FmO+880sO3
qHTOlJ5MZTWi/t5FU4N+s3ejz1G9E3Pjre82q65u8XPJkHth68PdkZDH8ZWIYbgbh5G0W9v84GQV
XlyMnfGaQMeckU3rDkrQ1RqRHSk2wvOz351Bb905Xflt+YdzeH/9jRtNMvpHYn+DG44AFc/fhBQa
tY4Lr/MYFJVJZc3zNf71vQ2hLwCsfkb8/EQ5yh8IhD0Br5x1nO+2RSO+MhTRS+4+VrtqKqBqRSUL
gSBnRaPh6PAMAlpsKFNV2ql5hEwpxZTBJQPE1QQA0qmOMOXf58x0r/7D0FTbv7KWbnQ7p/lmoamH
tyyRCOpPmsrDLbAgNYI2msi+VrLqAKU4zonL6HHRcpY7g3yAyTQQvnkzmBnq6RjVzpDM8Y/RkVNm
wNqlWq259MXv/53t043ufMXnrIfQ3hGSRMZWldU44sCdRUf57up0xcrquJivCE8+/DMo3c9Z5fXg
nw70BYAlZowbBRt3ly1z/7+mOVmsuJ22iLgWpfw3zNw88iSrPrAgS4YBvzMMJdVSGN7qxBXnN4qX
Mo7yKZodbZV3q3nWxISIZbOQqNeVYgvW+/3lF27PZpq9cItQsBY29PZQ0N2PdOli6dqLKMDyDnYF
5VDlKQkoIX4KMflHLsQJrxERzdQpLfg1OiF5o0A34XSM3FbunYeOh3y2OMkmylJW+kGtT2yECs2Y
Sg+dkJ3/R2JU54O9bZBhBYo7Et+YlbC5Dakklb9Int/stV/L2237Vba/NwNRUf31ELgBgXv7el2X
9IbH2+0DIjrvj6gFzGo4aNJXc3/VlcESXhydGxNvepqEJ+32/LS+g9N3CS2vKvUB2F+X3mbkvts9
pdg6iCBXErdTB24qU29BbpTJMgC3mGsKRqyJJN5cIhazdBWJgt11r1KeF7NXHkBm7fr+lSVFDPSG
nAilN6hzET1AjBSdhpMBpn1imGN8E+3xDJMJOKTpIFCpvXg4ImFJ1Bm69qMPaj0OZDXg462I/a0l
9ePdk16HX9z+OV2Ym/V8Lb+Ez5nZQDUocWlpIBVky3nHJK3Y8yIFujFVzHioOVxvdE2NwDlgVJzs
uXH/Qt/A7dAFHeuctLBDku3Ez3lKh2uerpIdRqtMaKmWHBVXh/gjDnrxF0VOiE5Ao15C/p93tSM+
WilG118OUzzIYZrtdH5MZvbYJBiNLk7dfcazmBNj7T/ez2C4ScHe3nAF7fP5jpFAnL1/+cmE6kRs
pdsir3rDBZfOPKkQBjxgIGoViqF2DaYLw/UPWFo5uJdqDAaxMfYzm2NH3+RPYgl5U4BirhlEzsoz
Yxp4oAEbe4vqu6exdN1UqYboieTRAtKV80aYaHfiMFisFaQutkcGeUZTG4wfcWu/ro8WwuvzBjmk
gGs5UA6o5k5Z4XqwGwpzHt4t+lHUzaemeuwLdMSoHuqrs4clVnhd4fOdPty1E3yevOWlmdN+4hC/
WbXZm5IXxVjGThUohkk/ww8pWz6F9Dv34JUv3wmcAnAt8WqCy7A06qoCMI4eU32B1zX1ftL8h2cT
W7sj9zw7rZksZw8Bw6WVS7BAwLqbXDK96/n/cuvf+makEg9xJHwO/okBTj2gilVRQaX/bgBBgccS
MQ/Tgu8pAbz3yK4neDp/EjmSxWyY3OWOW+xL4Eqs/mWKk9JmzHvGLhI7N+ev2Ssxd2nwyq50Xaf6
rKp2G3pLRFWVAx7yUwNeUQOkCDC3ECf2NjJd8MhzOmYhyXW3PDJLrm3190DQwrA33ZlmgBubqt7o
pOH3NtE41Ku07q+WhC4CWxYyoySL0z58vjeqf8jN6EQllBV3b9xsOMae52CXpdt/6OiJUSS6LD7c
PA8kcAsoPDDyEz7lGYXLpP660QI1VW2T142Wb+3qNJ00HGPkQBm6NJc1xpoPd11icEf84/5bAYaW
W8nEPHX615V73qg+dJQ8uJKMOajBPhTs/286bBPWXRVeQBijB8rVsEf6VE5egsP1lOru9NsXovOa
RfsrPEV/hZbRybvafjZ1908JhbBg9YM9KsxygHjAX07rtPNWI1plH167zO0+z6hxtnKCfQytnmCL
LB3jXSY8P7Pltcamy1LiI3yfBPnaYSLZDEhKnVNRiCjRc6BCgingMXjUgFPsuoLnIBgjMSzIu3mG
3IUR18qtQ+MkEUdaJ1udST5aStg0HliqH74n/c8QZJl++tCaJ3PqF4w+8UngCvpLBO8NoiIdu9ev
nVbJ1Iggzm9Y3SG/XpEUZ5xRmEUFi+HHI5bKpaU+GjZ/ktwo9VSq5JK+ZV+/bxjuISvgZAb81YAN
+8T4AT908mTqWrPVZYHwjnLN8sYvsup83/MMQEzrQXYyZf40kGoZRkhYOY4Vw1pz8gUoMJnbvpDR
XNyjeKa6XzfQn744O8D7bejHEnMAtE5oA+Jw248Xcqm3tK+pAe45VNXiTKVdpdSq0TqdBD5u9fPx
Q7Abw08UqhlJOZMPvdYxLwliFOcNxqnQ6faJasnUIcSPjbnA8dpVRXjMh5+PKiFVLYzW/fDvdglC
D6QHt14W+jfavSE2ttcMtGsj+vF8ybQ4zBh3uboi9BfivdNXCpwmf0hFtD/j7RNmT+AxhM5ITSO9
hlKxi49OH8FInvbIO+uY3127QQe309JuyAfiN+fKWLVxTSu3JmvgpuId6V8QZBmcSqb7sWc/AJKC
S5PVCXXUdl06whA5tDjdHpibxOxOY2taW9zflWSg9e6UfbUV6+PLtKsgsppw4sdc1Y/f7aUl/2WI
xNxFE5NGpAVALxyc75UgW4oinC+22TwI0PleO3T/DxdqYeef/MC38xpMPHUyG99J0CApCl0gtgMZ
y994aQSF6ZvE8Al7iOpBRmZnhOnzK/bsjtBXkG2dfzmwoPUOAvesrluBApdHn2zLRduSAhHP/2RX
fjP2fLkUhpiOUseRcuUwLmfhxb6OwG35D5YWcugCT3oGeVltlOmeTkqx7LNSGETSZviKf6ZagU2B
XT6oH42M6iFOju8CD/MDx3PZefQhUiiGk7/At0OpGtmcYs5AXgODb17Az3ubsFtqb7wOM66OmyWl
lTukakMK3yTNRn9tFbL/L/8OiDYSl7NRdNDajJ5XqfpRaytEPhdr7NTfILt5Vl75ybTAZbtWtKF+
dCbZ3fuYw9VaryyttZoSLBMofufeuCrJBXzkXWIUhXeNDmMSd5a4aQb4jin7R4Do88BkGbyiXphV
59lrk5Uplvb26GtOjDUmaF6nUoQZ/BmnV5Tjd5DH+erykLRhF5Xzb49ZluvCZmvMIF3uTXV8V7wf
10a/YQt7ZQLnUksZz2U8iVNnHipqNenP4szi9Mb1t5vv9HfhOFmmjCGHf0D4NbJqUct2suntcGfR
VHGPrPt+y0Q/hU5uN0u2fguAVib4tveUuzfl+I+FtpWCUKaE2h2CBPDSBJU/+KB3aj0HQCWOtuHZ
DqfM9kEC7+SWNVtdcQcujBDpsHn6wJzU3rfgRBeXRd/CTP+E74cHFyVYz/uulorzLmwzYl+NeRnI
PXoUn0OIf7+4BHzoD9XeMT+/MZZApgE+Db8jHJsLWCtv54bqLJYKu8nWnZugSMgU/Llvn92ytgTE
zW9Kk8sQBF7+AHLrahFPIuOKoRj5K+Uciw1oKKW+9fgHIc4Olmbn3LkKDhQffgO5GxTiM5Vn4QuI
Zzqugim3q4V9DnGls9NO6keEeShoRUKsAQ1/QMCkJZArTpof1/HzqXKc+NY4nvf2Q6Ig/P7AnODT
N03lEbZWDyYSghg1XI8YlRrKIoC3PWNBcHmac31zTZPo+VsWyz38ILvoH+3ic4EysEw7AeR7is8t
N6qco02uCIxhPE5lAwdoo7kmsGr9wt/L/w97GTy+stOZ8tWf9w3L90Jz416Qb8navvlPWVXFA509
xXam4faGC5nCdKhN+E81st44NqIizNobuxlFBQxbdAsmnl2muqsRmEGqGt7s0WTYe1OVnzAFW+Um
/jTUdSvlSZsOkEWPKDc1qWqsPaVz73faReB1tzYKqZBucOBbn42zz4pLN5SGvdf9+kM7CD0+xXoR
mjqmFe7z7NfsH4w0Xj4tp/mH+U56MpKItlXZ+U9vNqlEqbT6WmRcLcUA5ecjz3KMqDdktidkZT39
NRRLbpdGIHVDf+SUZ4DgdZ+oECU1mAIHZF54qyamupXlnKIfCNknhEpjRCQXUkmJOjJqAdsYdoPb
NnkFHNn6OgjtrR0VF0dSkxQBtIWmbVl5U2pCndNY1Jr/T4BPi61YAQh3pS0upQuY1WIluzRVmatv
MDYGbKBLwkjoVqLY8lkHLTX0UvDGBlSnyDjmkNPO2rjew9T3z2RNNFwRjIqvjFz59aGVnyOVOmMh
dVdG3zWFHAKvNIH6W/ei5/trjXXhqzkbUWDa3UVG3oma/bBjsys/u3IhDpthcJDqowVPOfOQfcdq
EqLhYRIO1z78w1/Qfn4fMzBQogCbPlZ5uA3wfwH28sWWN22WVrZWVkLCctegi2yaSA5m0kVFY2iq
jpgkf/diSQHEb44UxUmghQp04YD7b7/p0Rc5fvwSrZG3Pk0LMKYOtIP7x3tgt1CoiEb6Ep5u8hES
lpUWk6bmaAZL+I6xkZhSDqqsvnyH8lFUF/3C2rFTp2pXwSRleGtR+GwaxECSFQjTSlNJd4dnMhes
d29eGDYS2/62bwO7Wsa2pq7l74MyfeGBD0q0ESmMgFU91xK6KCpNHmhrzfREZPcxzHn8vSiJVDlS
52SWeOTOHjx/8le9T/LiTWSObV9MPMlbvxQkNYjlt2Hiz2rkfw1KeR5FMtL/CdLTfSQxbCHCWcQp
eaS29gcogjsHK2JP0GEXk4QbZ+bSij8OffClyToLWBpT0WlDeimbUgDeECtcXO5OCedtjeuzqneD
oyoPt0qx9cwlG9E2Ef/lTKlGSs4bZItBVsX1YucMfx0EpsnGA3WMyVmf6kBw2a7R29utX/h4xcBD
cV2oU6SfPXHklCUoS3nT7B9G/itzUitRTZ4Sze8tOe5gAt+2qOu3iXV+hPK/ny9GlH9HQWLUcSU2
KdiOAdIE6C2grDgJORGliP0j/Q9FU/BCX0ou3wl2uORYckX8QHP2fKUGNdhkTNYb6C0Pi2pdFZNO
USqdfn7eH8r/kZbBW/1YQ58GQDvqsx49wbsvLktA9WrmwNUNwmOR7e0agosBmcx9rYhwjIl//gDT
CrhSu4GHhZiw/pDU+M4y88Z1ZDjvknsWsUeD9+VL1qPt5fzLteNiBQsNf/kF/bqWjV1Rwxw1Xozp
WMOybWNKg0W4ksWzCgf19mjp35a8/QfDNaSuU7c1HURHEvwlZFoAN3tEcV1YTEUNwmqdubhlyrkh
MM2yg6VBKKvC3YtUxnkTSLkxlfPhqXOhZM1NzmAIlQLQJiYpGUaPoANfSJou9yzkVmQID0YugD0M
/mpaOunQiGtT/K1l4PfwaOeaknNAo3HQGf4IYbw+NLPPqVrnHlI6j3fHS2JOWL66kiIoz2GI5Jq3
8U7jZ1eb7Y2PluT59LzcVtNUVsA76f2sI5GDBhsvhXa2jhAIWUypMun4KKyeiocXceuj3Mw2isSR
U56XjRPAoq3nYt6QLEIlx/EvolRbd93Ut/gfYG9Qm0UIEJutSgg+7AjwgQnStJOaILFVVLnLM3xu
RLXcNnKG7Rw10RYjBms9QjW6DgacIK2H3VTfsLQ8J3zOjF+psH/HhRx7yGMNHM733D8yidxoGw5K
8PrvOgr48CGSJXztCNoI4x2rr0tj23rSEse9xVOq58f0sbIriHp5+WoKfN04ooYjKg9tVBGmtmql
bsvxO0bqGBJIfpeiKDcv+Z9ScNgO2IBehtp7FgWfpFyJJ0NBDQ/XepNp9OIkGIaNJ8TOGJnF+TgV
tbDe8THXyO+2jnO9eaBgwjtcjoJ6zY1oyp5aK08cNIJiiUx92k/Z47+1z5jK5M2p/Y0WoWyBo5Qv
Ocqy/xYoAtIr57skcCY7WE2Qaym+BbTWdhtpPQvNaIFPAm7uipg+HixBHfQLKGSWsw09FfUSJqEs
xsc/Ij4pC9n4fuzTb/27zewxtHZ7jtHq26GaWa4ksNzZM60/knkNWS8JVRFYnPjTTQWEu/snnFgW
dp97sc54XRnsVS/LcwMHfUmoN8fx6gBPCSmPCqro7SNoJLW8Z6nHIcrv/1uw9nTM2RLqWRSuYAht
4S3MNixT0TaK/agg+0iUlw7U72162Sq0vGz8llF+NoGHcPhk2B9/4C0BlMKgpsPOpxWSOMirMBEe
3Umcc5Vwd+ASZU7BKJ4BCJZMvVTH1EUfLGTnhgrYsTREa5FhrQpJU4QB0Ma7mtbeNXjeODQGP0zR
0V3n39jRu9sUz4jKyrjcDkzaYi85IAINqI1Tuu+Dm+sEylQ02t8KW/VAAXtjqfr0F49BIFV2PLzc
+jncfOSaxFq21M7qr2SvX7oYuLzZv+vFqNaUgs6WKu/iFCqsbkHec6Jsg1E2lghAHpF4sD+MkmFT
7ZPMtWwbx6158bq9gw0cLJ38VM5NHADjT7pIUiXgy8etftLcKD5NLhz4tHtOGsROozZJ89Np2aVE
+oka9A0jdlspQ3CJJhusm3F4pSalw+wCw/Zkr2GQzLPbNYKWycTLB6LYr523QGPDaBDjScekmpR7
yT6p+4rxPSHjYDclActoK7zjpmMJjKn1PXTCnygNZ19mayfTHnNCfcu3Y2RJan7nN4iqfQt/0v0W
vybBJ/mkBJkgjEnQIMTGG+elmslXbLcVEuStDXpdGQHky9VsoZvU104zKR5L7MwsxHgnoE06unrH
anMhU6Qi16wbd45bMtejyWT9ng4dD60bjwN6ckMj08BXHD2I8NZPNZTVVJUpSxcTWz7Ngk/gTo/D
Ys8x/cpXB+SHYP8ThVlBhdpoV5IfqpC2RVR+NAvYmiopWawL/H9ZoUX0/PHNL1ToYyLEomaTHFD6
8uhfffPxROs9QKrqGYylLQ5CgJmdUerxlc9OHxQgJsH3dxOvDiS/f/ZzgzRI1PAk9vQpjsk60x2o
ZbL6LOcEPueJ/zk78RdPsx9YOXZ6OTEjOd1ReQ8hR58aS869AQQXqLt6vu0VOeYOLUTWc+oOsuWo
uvcMtzpZxKDOUvdSuiuxcHQfOm4G6LWf6HbOFeCUncoVVfndA5qvaR4WF0HvtxcwTVZe+ng2lDRy
vHn+7WQ6XTT6mOBQHCSKYMMhutrBwSgUioqKpuEDGqr60xHjtYM5TmjXwwpMeUq3bKgpieQCRVRX
jxKJ1LDo+EwWWkXfMmBiYlnm/z+kpWlQtVArXxW4NhpZ3Iq5zoGQd2Fknh8SNJ+rbNLGbAsHDuVR
vzCQ8wafAAM1RfnlKOxLSRoZslPUKogs/zJ7ze+vfx2ns30N1G5cZO05dibtMxNlytOA+LJBz7e4
2u+CqYNLo8ovarp3Wn2IDHpCGyeHfX6BJ1K4EUk0rT0wnJzpkKsiUHWu4MwOwhIG54iWDJ04qU5X
RoI2eWhwYZVGKjFm+9MGOb94rozUxn1fATWU2PofRjdxNqZkNfe98ES9h1sWnq6E1XFFT1Rix1Rf
PjuHYnWwfx6hFMa86lwdocng+loQPp+kxXy2qvjLElRVjimGbzDlu4XflIS0Tjsoub6iEuXhyECp
F4lH8R/pl65aspMlO8ccJIIy9hDn6dEwkNd4yaAafyu3luMysh7gTMIXu+3X9bHFu8AtRB30JLny
B5MHMCm5Sj8Uu+9CJNlpKzUal5DSX4wvTbBqEZD5mNM65O/z+QcBZzsnBVirbNK+hMA2sC3BZnUm
hOmSvzDwW5P1siX5KFq0ATY+jjAFnHZC1hbXfcCX9+xZ5vkCeCeAr7DUs+O517REDYmFB9tMlXIr
HPDf96AEBq1EZO2rEzE4BQOZGuldMLFEFtWxhf6xZOn/zDFZYZGpsBr+o1wvQ47SoVkYjBHIVQWS
tFGxh9llqGbbniEaEwvyrV4yeIwQI/wMdxkfaeZFZDn6x2bS+to7oeQ0bBwn/pXs2kCG0RcQIVyG
8et0PddN4sHjf6j/GtDEsD6fyFDBotI+OlDNitLP+vBUYsG/1tf+fyj5d6HH4ZhM+5kLeZnuqkkI
Eov1ZNBa2i0tVRPpnmdrz77Z5IeVMiryewa8gVqm3xyDzKEF716e/N3XlnJMrZFj7JsJ/74D8l2C
oBUjh3hu1xToXN0B6CXnXoS94KjVgt6P2stU4/LgLX3KXte+6/l3IJI5DTrgRo2FjeDlo2M677z2
FwC1du4lKDCiiE9RR6XIWgy2poQt11v3cj3yNPevT0wiJX0pwQIjd+sxtcyeUYDOObp2XUAlDMMu
gi/QPZdsNUeHtFJJAs3jrLZtiq+WrNOZsU2lBhxBE9vaCrQZy7iOrX5MttZ4XvBxcV0MczGl+WIS
cTIX0d+5l5YWstgaohYuD/71Jvuy3z3dRKMbeHBLGaHXBg0DQX+Jo+2Iouh7D7/ylDPt7ZG6hTcx
QrFX4bW0+mZS+RgcpGmiZ4dTsTlRCB7A0OmKG6WjZahjmKFOtPWjJWdz7LYTm9S0SySl3dIbOLtn
hx5bHdsotHIltmSUudiy7wjQpoNUnNBs8uYEQVECMf9myapDM+PR0HCM9753BQtFgPEfOn9Nkm2a
gt7R173DabIdcOFEELS9hp7B7aYDstHppIWFewN8vBeUOZGz3X5ek7sJWZuAJqGGc5lf3vWHMXto
n80nMtYbC8mK60KgYaOD02JM2dhQE3ssjdYnEFu0eEg7BiWP07L93J2H4JI0FOsaI56YVSwCHGg+
KyknsfR4WEFl/SBR7+HPtm/kb6UoBaksda75iDftY3xtw+wkNAXODQT2Fsc2fe/iu8rEOkYo7Mp4
BMgSWVvfZwIrdq1qsMwgMwtZsyzDflgMYzF7CG6Zk8OFTIJrJlqHo83eKfzXOh5rATnsKqLyEbrb
bMBoCZzoYJPaXTx4tLzUNXl5fYOCi0REaAOHLkPOXXSzH5vYbqRbzKNRTcW9JGL/UaXxDMVADgUx
G39Sek6jLKjEDSPgG9aRetgb3inVC4gxzUN+LnXazAkQLXDSq8Yz0Ar8ZJMzpe1SCgNzLkWXwMLe
twcXTiifuAfBnrFklC86pZGCdb1wa//WNXydqCjHMHxbUpVuZyB5UxDqx0zvvH2SIwFpnO3Oe3g4
PqM9oM9KnymTshSSn1UKAeV2qbj/sksWzTa17rsuegjmR4GO0tAHv5UWvIIeFAt77lWOiFicfFI0
uakdzpvL1vh2fO0WsOyepLMMXN6LNs5I0pSD4pbCVI5A9e2tyJ4LJ8EuL43HPU92e3ED4kp8P3IX
1Mnq5YDPNS9pDqS4E9VESvpy4ar1ftEg5g+jRoi4xZXTTYLYkoZl2aq38bo+T1XiH5ruS6ZXbUaR
Vj8zx0OBVzFgaPyoc+LsM59fGeTXiRcr8Kmnr13ZKmHroq/FuAnkq5gHlnWCpf8lhM983lVR/GB8
rzflZ79+szTFIS0Z3Mw7Kt33qJdpxpBdy8jUrGNFLbWoKW/JKgsxnNdbRmrHzc6ACrTyahcK1eXB
mjXemY90Prwjbo2V7Ki9AX2BTa5pYPGgNHryVzgkPScld+zYVGMPlmkkWM56wNKkOngvH2/Q1X8z
YJrfeE4tFstGK0/il3EFDVYnHEjE4NEpaZDyK2DsPx8mBbi+P8A7hhVyKkCcZmNO6lk8yAnDczAI
GX//sG+oUt7T80C25mER1f59eXm3vjyXhqS0DngK2fLwctLBtLANsFpwJw8GaNtU2ia3ys/ZI3XO
loHkxIag2aWBO8SvwA3p1Ai3huELc4VLq+zNZ1H1bmyHgrmbfdZItQekDB06PEB75knmvk5/AHje
/WTcZA2boRhUhf0NNVfnIPxoor7eQQ/pRtF7I7v4GeJuBg4ir4QG/CXxPi8U1zAxIdUmoR1iE8mP
tXKoruIjPec8fNmC/C5MQhuyOi73OgMGq3sD+8/R3mGW8IynIOZwGTlTgDfKWgE3RLyxHEawzcnh
vHURn7uOs0zM/AsIB/OjuV4yzbRtsNFi/VkvFzWldEU8b8C5D4Qllftkmkz0tZfGD7uaOB5XN3C/
6FvJdmb8caQCKIvWfSPb2GCC6wWzWWfTWtBn81te4tAgZD0ef9lybAhmv51ZOJqLqAfjey1lwFgH
JyCBoGogBW4pF+VBk0xj9Xp5XRYRmFpZYkg5QIOEiSnUbn3O+u/sFwSp1AGYag8lu3pCkyTFLs0Z
lAlQRyQHdP1cbly2ozZ5bZw82An1Wkh7+Qe0LShZH3YQW66DuaHsyt4QDU8KKrG6iXJNpY0Cse9X
j4tBvZAsxQS7mGo++oSYm6NlkYWviKXS1LuHe/DVot0UI1O2h8rbIQINZMDme9D82VhbhQHeSzqe
Ln1XS/01N+t16+RjXJ/XPg4ZveV/g29Yl2exjFBoXRdATaJkFtOV4nph3oDNMlo0s0GopYYhaZg7
VQTtg5orB5d9ceBjLMuQhr86Mvu+L/5C6oDsH/eHbQKerlhH+j3a4Iyf3bige8df6XR2UTlyjHdf
PrqwL5tnWXJsGRkDhRvSLexlYZdj51GzEJ8As2nlSHQ6g8Tu+rixYmGVofuPV0ijzFprMVgh8E/S
1sDFr7nILWFJA3Tcxrk3FuSKA1/ZCT0aBKv/vUPzV6k0CJPRSCiP5wQnPpvVnFPB+Evyuq2wQ/44
oSfXecXmanyCubNR+CjEb9Jrd56rDFuK3rOPUUAOZKLR5S+vHgngXsGpkmrBTaEIozap7eChtfga
Qxfi4x/8DrM5MqelYR8lUKI18l5X08m+e5j+yugaKf471H3L5ICLORyEFndoig4VEiNmqOlLJRz7
uAJvfd/UV0jte8MCITwnCNi7HCPK8pmBGWtngMPlSOPsE4YpmkOzvPnIjOQBknvFjZkqrLSmVnXG
LjiZltnvHgrCJVoweMKYyDQVBw5L9b0CGN+YRsdFTqICXIKGC6adjCJKmIJZTwkoxjuIiIRXXk2n
qUTOtXsaeg1w5vwcJKjA/H/j1n//0aUmIC/y5d1Fr/1xIvaXTJs3wnJf0slpUEo+CcItis22d2ZG
HtYMtUUkMCZCvv/70vWE8CZrWrDic0+6WZCEQdDkjdunBRCaRXt/4VXOv9Z6EQDfiFb0qI9xhSEr
iXgam75nCloJAosVEh7QJspjauXJoNpCsKzj2ZWWbpqjQ8WrGSv+AwSBeaeJGdL2n5JuOHtEpP9S
wGAy5nwzqhZj4dBrMhAG19ExzG6Sc/jY6ERu6IawsvGVPN78CLboGmzoBRWHBNfT9Hi0syHmSS0K
faF4t47b8LAVcJj9MIhcvMfIO6kGIWrlhrpJGoFptLIh30CJgw+DB1CtE9jRGwdezCfuqpa3X+p0
Q87bUgIgaI4KA6ay9THv+e4LZ7AQHudadgZ7MPQq2Id3xoJOPPn8RdgY1+L0j59jNFirvaDVdsG1
L859cwzuIUigkPwcesJqi/D3v1RInURSEl8bF5FnMTXDy3Bcr39Oct1vPFNpAub5zNGtl0WP/Yd6
UbEk3cRWYdpp6k4vIHgZQaZJxnIHTVm5ctxenlLeiXWYCijglQLU/s1TC5DJ3/zd/jEEGY4fqsKe
ep0E5q3xVkSzJabT7qMObOgz7cxWXX6vvqD/ZyRQk5lqEqxSDuS60Nc3GrCOxDJOM2ckv3xreYjR
TFFYL/by+9fSUzwyF4DpF9VCEpG2JnkbXBIRrkoMg/Y48P0QPinLFXuC4ePnxaVf/kDfG5A6v4vw
YeVaDlO5XMUxdG9QwbzK9i9v280v6efOMnlb4YisfWIna+Fm7eNSaQ0osb01ZP88cZE9gC19OOg3
d7yLODi+05XGP2B5h1biR6YaclEvZB+7LgDKwUv+T8fNUdlMTKz4wF9hgXtJCCDrwOT43ktGXzWI
PSwyF9tJSE1wSBthhLTk00vICYsoedhsE/IgwDuzBgEsGaxrGPpZXmCC312HRWd9KuFFaeZ9f3jy
12W7v+4HVsi61vXEaeemc5cPctIWdVr3333oqS4s1GlraUp/tSgHLg0ZADBAQJmFSmlFByfXLOeM
BJWUijsIhEQq+qH7IuJATKLIzhRZ0HMw/8c3e6Wk+7NTZF1NZ4l8CZnI/jFI8V8QcMJ23WBuTTV4
dEuQhjfZjOF23xDjn8pVehrL58a2uBSIC5/e+Ry1GYmoMqU6r+pANNucOOZ6ZhVHeH8Xh1ScsFVk
lQivp9yjvyZjxJV6hgqnRIxIPObrHl2Qu77BlP7ISFcwgFCaNuNUpkzxETgcSfmNmQAHVb1+dcOS
xsJaHIXOUXRExoQaakWdw1z/MJ3EwzuQpLD6jbguts4VeFt9R67mRaHDYmw+sG6y5rzwfi97epuk
R1/ICnd3BsAaP0NRE2ELs96NroHSI4R3sfeRvjuj70TQtBbwee2H2iwMM83pV8/hyN4u0V9cPq8v
7GHpy80wKEE1bpuDMkWl39FYJyL3z0ftu2aRQ4ftQoTZ5G293pZMTz94PmzofIGn1+cuH5dS/sVh
9Q9VmGa4N2uGKgdWCPHUFgP4+MP/Fkq6RS+vG5LsD2+H7AbFp5emOK9akxXBKVAk/KF2mh0t6cfQ
ov7CP8WGvghMXbnRDAPcGrDtIxzUo0BSwBMHTxcoO4hW1I41wPR4oBOA6zCyYwTen5fmG30DeZO0
FDq3EDSU89v/oRl65wO74YtidfYQ+DcPbyQDzaqDnxkmYUMXpchiX4G2ktvefkM72FfRCdAdGsge
bGnLthteFGA37AXXyR22Lhsjz+jj1LtNq21K1NOPEq1hwiE4mf9pp4kyAo2G/Ija5jj2eEtcJvHc
4hiTWA1aYrDthXXe9WbJdaPjF4KF6bdHq3WkLJhwwI/Pw4B5InvEHfQ0Ihh9wDKec+bQWEcz5G2a
zIZQuYeyh3CK6u4VgJVGCK48kNpGORnvDpqHDsfTaBbcNJSEklSVlH8zJonXx/mUM+JOljBOlLuD
9kKfWNeokM934bBDmooTWzchu3ili6Ww3BFlXq/Ryl/OmEfiCHdtn4YgxvDHfuX1lSn/ym90jlyc
X4LQRIr6/TNmhmk5vpCupKJxCVjud+OSGR1eT7NfEK4/RhZx4c2g9mIC1bSbvHF4rzNbqnDBe1VO
9UqUcDfbl7I0TMQLuTWjejXY6URc8rGCXEgrRSlDoyjqgQFU2N8qF9gXhe1UB+IjHk6TbL9rQIwg
SccvGq+a7PW9KGx7PJaPx5f3+6MOfe9VjzeTfj70vqKQk012fE/Y0UGWlWc82pR8TcAsTAiw9UCV
hIIrKrdnNoakCWXZ34aKw3sHRwS3bQZl4ajvqxAZ2SDunUCjvaHS/XWIu9W3cMgVXoqjBRTMfFdW
aN4s9zsw/Ff04EzTZhzbJN48qOLrpqBjoCOmKE8QBlcJtjl5imLYF4uMr44tyGpetw+/1ImJMq3e
wgXZ96ZF06kBlho0DVld+7g8/rglfaL2PS+UE21yZVcGSRLnEs7SeuJx9Kkf3Wbws8mFvwXRoSzF
1cqf6lnmExG67MDxKvU0Z+TX3gXAHchSjpKLNLENSaxfrQgaaVIShIlvJYrAbpxNamVkCKbVPePm
lgXB3WZu2zJGZ/GR10h4CpXBpancySKFrmWrndkKWdkNIyzvfGEcT2NbY3tXNHzOMcixnUTxZLe/
FnZlxaZynmTzMWj8Jf1+t6EqLHJb2ZIfjo81ieedNMXulGU1jcDXzV2iwChOkb+8209567X+/ebf
YZZxTk73Am3k6+Gbihpj+qsClVEbasg2uOYTH6rXuu5dwz5ogBnLhoHkUGd48IzSUn5qT5m7GvpP
d5DbSr/h1D4d6gxsxzHwvf/vWD2V35J4qQjLnAUej58wLp5bsQbTqkqYnLLtlpz6V1jDUn7N18cS
regfAFuNh9BkWkXuTVQ9FaoOBeh+6cwg/3Ua2UnhytcAUZzCIdvLv6DZPMtr31qkteETuEjqF0bY
Xh/fBI1/Z6lbmMAwaoaoxzO8SqpK0FqzjrlAbeAtMqvtoUmwenBnCL0G1x4mEOKcoCP815s6etir
mbGe39xdgq3YKCbeaz2R10ASVtXJ2AgfzMSG/o0zj8uot6zzGxpJEMxYHgiIelgy1kuBhU8cDJRC
fd8I5vKD/rcekf6OliI7ITfUvq9dCMQCVWFbFzgYQZ993Qz3lT0yO41aQ52pRRfSNaF9k6BOXil4
0CImqy6LJ48JZJpQ8eEqAAAoT8XZehikDYfF+2n0yUf5HWOuqM7ijyVqyoLZqH0Vg3xlrzvhaQpq
J5YGzF7+lE27HTxG5AwTJYsLebM6T/dXTjr0mFE4Je6sXj2L6GXJrxwra6b2srz9qq351driiovy
8mAoMb92ozvG8zylhbexnuFx5MXmtf7CjIC4x8IAE43o7yVriTKg+0R+6r/XXIE6hy4gfUHbjo0s
qvZRF88LKholOCf4ttvMHXycTmFqOMpDPqDomqFPEkVHq41VwKqlgo+g1Vr/3p8yJ4uKQlCS8QL2
ldTApnVHy2purAKcTxA0hqWJfaCkdlQOXu2+KtERapJe+YM0ah3WD1e8MTBMnxkeF6xKbZ/LbQFn
6A/wxpuMzyH/k+aqX9BFhDH4hw1ruTdIwvxYDOtceOS4OhUpyuj5SSn2uDsV0/RNZjbomNDkSiX5
OpyCChQmcd6+LxxqOz+JlLRBdgrY6DKjswOs2W2084KBtYr9j7/E/PrYqAYyGk9sfDrhDEd6+jrI
OokzYV0bO/34BFCMdr+v7rCHplJeaujyRAkYQ9Nqb/Fa1zKDanHzx71RTP+nIO2wfxu5DDG6F8w/
Vi/S/RCsQ1vsupC8O6FdsoiUvDbI9jZkAN54K+zzUKBC1opFmFx4x65XD7W2xbvebApUjGyTZNXI
4dsk9N6OEm22BE/9R11mXkD+C2MRYSWfTLLlJav0hG6GVKUtc+GQCTA6exQg4jzIulJ/Py9LSQ6w
gWl04naXGNrxteu168spKfuC24W8bsmx+VPl+kQqhZN/0kOEU8atBVogJVisidJMni2+Gx14hUW8
iGNCJ3Ovt8ays0Ops4x708VnRR7bX0vWYOuhM5Q6HnGpYEKYePpSP2BG9P9fclOt9kimmjLAK3Vu
YND5Y9YTOGoNnwo3WLFbGv5VuEufgXiqnJLDaxtm2uYIvtBjelAVtPiWOlgSIZWGlDh+w5L+bLV3
eVe/bCaYgeWoC1CfT4L4QaUQMNOANzFVztkBJoNzOBHS46VFLdjsLIuYCT9gyXpghO8iAxqG8Wl1
vLw0TGvQpY9y5ZHQxAFgnuMDfK3mkd/pJQog62/6nsObxg+WQpKDCFEbkfgjiT9xMmLA5o1P7dHv
KbTu9qtQwreyIOUR0Su/nNh6Wx4oaZiQ46xTzS6knlphzG3MQhP/2LF5tPaqYq0kLVvkboB9ZRT8
GPMfzRXXtZOio07nDKJ3lW/9GidRwXAw/kRavzJYF/fPiuwhs1waYUNX9NHhCDUD5nHy5h/SITqy
0Z2+iOnqYHkuxWTOvMV/NJCm91z5o/f+MCAuMk4ujHUkB+IDsl98z0zaPP6zag8zUy//Or+09KtW
YrCWVx4NRN685D9CNeYzNW1M1HAUfs11tcdlYc3r2fIhyVJ9N31G+5sH8Og3IRfuyPeQv60t91YQ
WR24xTbzsnA77ScMEheP4Db2RnkGyK9Gz5SS+1Q8T2h6C/gLOFcneoaZTXEReF0yKjaadbrZMy2w
k0wOeiJyKpM1Yn/jBuXJqecRhcJZq3gJRVBf8CyMDYmemu9WSDrJYwgMlv7cK9TThgPu0eu5MNDY
C2omT5IxvLt2qDmXlnHBfc4ts1z0JRzK5qRKCvMBbBpD+N9DnkJR6aYg06+XkYYEarSl8aEx+FQb
PsIzVDwo3pWsTTjKKT705sCxBx9KzMiQ9Ol/HaSoQJm1k6JPRS/PFTeBBO+GPBKykjmIsb4fGmY6
1USve//qk5DvP8zUxQfwlJPvh28sC0zYsakQnNPDm8Qpaep35mABSY1GyUmzqiifxfrdfpjagUyY
YZ/7M9JRP5p4VWxe6wW5A4rGHYyhD9NDEvvxz7nnHWPj/uGtMsHowhf9QI5hqlog7/H5+GdsAqPa
SD+Y57P+o3hsX/866eIuqmBd+SsgEHHBYOymuHQQZMY43gwZWkfXUgVzVvoJHgxdl6gJuZFl0LJx
d8axNp+2AO8qIw6EzJSZn7Be11WWKLfWI+LSZNzlO94N5PGmkxsLfHGYA44DffcfqeSBZmxa/0oG
le49lytHY2hCBGDO00Cu/mrGVRHNKHKYhywRnervPVC/f6tTCk5UgyNpZf2nF9TzaQ5ftxpa93y+
8NdYMzau/p+c6c88AiwIwK/zLo8XzwV80QVXeHHbQHtqHaLAyu0X/9v9e/8OQimCUGwWoJv6RAjV
M9AxIW/s5DTB+mX56MsFYbXFiHZ6jgz58dVp2EGz0cBtts8freyR6NRHlwd1+vTKEhGQ/oVZDQZJ
I9S/4AOBOI+AausG9pEBAXeUVANLq5eU3qaebgHTHnm/adD0C8gAfMxxL+dnUftr05N8UZ0qorFb
vzU/nW40By04HrGJPt+8QRiKkPMLaN80CGnUc5h5m+iZMBcPZ7YoJkC4zi7d1S0OHm0Qk1msx5xQ
iiW+YcVLMserfLI/LPIeB2vuJe32tk5CBUsinm9P9YLmfb0XiMuNcsAlONX8+uofaTcqspAb5CBJ
gjhgvl64jmfD3+mguF/NMyHXuUs/8iiug6rFo/Aq1n/DrvfYD2XvD2KsBcJlj5/euyQzo+lh9uKB
qpr02s9cRHoorSqXtg9V1EUVAK5QKM4ChneWUf3efm3beRLWcBy5djQANuSCTyPEjaLwpy6oCCHA
vl6w12jehsrwkHm6+FFQ0TUZdvMF35yX2UckpMFfE5F1ak2mXQR8ye+4lgArHtRDNwCFclRIGG4C
OHBYywDiJzUNa9yon2Umbgf980/bNRMuAykeh5MptyzsoJJvAWrHMV3pEVsb8bqELyZZE8FUiCDu
Jj2Co17gTyXrN+HRV1NldG8sQbF5gD+B0xaG01cLleeTLBe1igOYKtvHDAqy9kLQo3fUyBh3N1YG
0GVZNLmrhCrFsufB8RgCRhh0FwiWg/+wSUG577+diTEh0XY+qucF4dEXhXtUser/c9eCHG77vq9q
o8Gc8Z1ji+R/4eAkB84K0mdEKUHO+3d4GzZ2ZqakFMGYr8Hkz+GPWOlWuLKhHXeK7hSmakx89DCG
uZXlzn9mk6fc1R/Gu5O3RnCl4NHMZwOsqAzO/FwHg7RFq4GgsZ6s3Uro8dpvpI5T2+B02MREnSql
8Rqef3FtpiV7Nm1fNggvynt6Jghdruy2Upfn/aRT8eXou0rm1MCUztC3jhomXQ4aRO6xS4+RnJyg
1oN+L7xzvGGEp+Ok0bmLa6fdzHoPYqbaoSSdv1lL60SiiXCRHczZ+UTLWYniGtN1PcFAx+3nbPUW
JTcro4pwytFSfrqyOfFiqtxJU41pfOi/gLTpPl+K+FazEPp8KnrSgG+Xl2oV67rv+g5fn0Wyp7qh
vWLZ+Y6K2fjiHMZp4DgTvCD0IfZmZuwHp5ISRnk3xS9YUcU7qO5QhBahA+7tmIKsOMLTW36S8KJm
2YLAHFQb6T8bNc9vc88IodUyF3Xi5fujFuKchY9l+pQnlb64r/R9C6hRiKRvdim1McRkX/r08UmT
1qk4Bjw+yuWvHw/vZO94LSOn6vTWwAQ/HaVyNFXkjWimpCcXqTkcdScUGQ+XzAcHMUaC+jEZ3UFl
P4S8v/opug1mgJv2scaBVsLEmho5nY/tNwalUjfalaiwYziqzk4SItnCWiHWU5v8Dm2ZpY8wJryK
5qP1WTsA+7YYWty2UEuAgD2CmfxSbWxpQ+elG/QJ7HTDGZ7W0ygPIBbpvJNUnLsHF2pC6g+1K9E4
SH/vVcMN8GdB+IRikAxmsTPpGcZsleb8UIfe09HjqcoRV6Xl+PjbONGPSEqDXkNWQIp1XDGqKgkX
iQvRvqAB1rpQQXTrQY031U5DnemwfAH+XJX/8dBbeCamBhQbFUvYSwz/H+I6WgfSjbGV85Z+1U+L
tcw3DnIEn6KmWshEp91qbxdeDW3LmUWG1NBYfs/phN5ZXxUYZIHVWkPoKOs5ZXy4RNDyAInXn9tz
ZCgD/tAv7YFXd409/b9qJ3Ooh6v+40L68yTnmTsdnj/QhzVimBIXL3tnoXZ6YR1ySjqkkHPm1N9j
VOBfh0PA1Y/5J/KR4lq9rZNplmsBzkZ8wjDIx6bB6WLDlJePNzWrxma7EyaatUie9B0hsvIqmcPE
j1+Fnc82yTTuJaaTdDbs1PkzzyADMV2xS2Qn21xx5JJsVC+ADwQ462v5oyKh8n4NRdZRZyt+kkZ0
Ff22UZ6g96fSOrtU+vK91Ofwiv3altYvTCkTEq/EQInLCrH+8dVA9BjZzih97PBbGi/4tiVWQv2C
w+/j2TWVcHpdRVUFYZIofRMDZ7TuFn065g3mpNBLNhCLZA1PlEtvT5qL+QyA3YxqazXj1fJpwAnj
/j/i7Z8ZPPPFy0FNUFyAzHRcrZUOhplxHt8J3Lvsr13IE5klikLJuUSSRXVcP1eeSbZUgzZVR0Lp
nqJVGL0AMDBacZ7OXPo0Uxff1+0pklE3lH3NsfrfYDhV+Sq0igANGbcSJEPAsILo78wEqFbaBZ5i
HMNOw2uVIpR8MrID6dpV4Y+BpHGonebOpj8nfubpZU3qAlVOwJKghby2KIaq4+hJvpBaFoYhuRpQ
/H5R50AzQuwO3TE8LiR29RuisoJ2U9YCFx2ZkzOfbvLo9szwMqXE02vXx2SqY/zxCWa+dNO+a6eW
7oH2os3+ti8vmrRSwSQXws1Bre7mG/mzbQ6MKVBU3Pdy8qDvd51uhgoEVCp9GDjvBJ0l3l9TlnwY
6BnorOAbTAAf5oLeM9CxZRPSMaJXYkvbGuZJTHp+vjcXy3QjznT2XfK29MBfGSrch3ZjdtxYDqE+
DlGXgmad5h+jr33WiUUFzhol+c6eMXR9fV1CL172hj8YqpgUO1RsLUXASDyZqT5trEjtaG9ATYU+
s6JWNLqhQ9Ni6StVcrIiMqlq4S+oC9Hbf3VO7sZ49G3kwg/6ditlAsZZF6q2znJjMKhJDCcGM09i
CoMleCOipoB7rSGDnqmaecfa1uxLuEclbYr3Ogc54V2KbgVLmG2i2Eub958g6L6sBE3xm3HJgQ5m
ZgpPgpymQatGkLnVL13shKhSlu18Thw8XjEvhXVIm4Mh3LGwlKEiOGvL2+PLa/MzGhEMbkbIu6nm
3Pc+5cJK22L3KWWhXOs0yTf9LMBJEMGAu6ZPxfJDDruuWpvBsDWCyhtgnf+wApnn2vTd/aGLbd/1
6ovYel0dMUz8+nf155IpVNAqH5ABsdsfh8SgprT1+FxqE+eii4QvcMIs3/P7BGfi4t6IOIe4jUg/
sAd5xvwS6cFaIll1aVUqoiZC2M4QjdMxuycWGQmZVMQVvP1MIjoz/Y/hwaDkZFPvqD1TBWuNv244
deJPLWIm3wkN0uW3N0Hc99A0RCqVjTatkNHQJG9uSzzzEYNc9TNF/bQL4N6TTficmcBomQhYh8qv
jIGDfcVV+wxJRJs4Wl9aTDRYLajVWSJYF5PQEG35HybBNaLnQlozezS+DjS85+CuAybA8k0jBb4I
3l4A6jvP4Fqr6jxmXZDU4EhVvvP37yAIYJnaq/tQIJ3OWlTbgnaYTWrJy9ujJ4/smmR1+wr9Kfeu
bl9m2eS4B8hGy2fCRWKW6mSJqoXWyK5M3cudQDLtqu7BfrTDORqxtrASMU5RRUUbn48vjfPzwGY/
vEEZtGpG9qdtbf/GTWml7jCH7+WXqR1oX2x7xCGuyVSkpeGlxM6MSQQhffh2pGK974Mj0qZG4hYD
Y3FHl5zJq5G6Lq943bZODLFOnOubNGC6iEG4/YvES+sCzV/1UJ1aG2KOdSJkLLl50NsOHUQkixHn
aPchJD0Anf3+coT0qN8HzQdeAHrNgoH78FFhomltf5bVicWZqZWOz90/eMPwKDmcdMEiSn1CQn3T
bN7c+yU4+6NS8Zn+OK6AyGPXtZ9n8uCsduJIWQPLyPEqxVUJMKHu3iqJA4A0/9gahrU/7y2Hmq43
+KzGT97Rcp3z8dnVn3rtDr3EnX830GRIy4AUCoBeVGq6jALA7e+rQ4uUiv9SReCxL6s1pzczBJQf
x9dxGRwrDmkra6xuqEBT3wBKuJVencPct7Bvo8aDoOJOXXpO47MCGHdSmavTnpxFwNU5AjnphkC1
Qr9IsdqJrjlZMDkay9F6gJdfDF7jpYTWBetCygDZPhij7gi5GvrHwgN4areV2s9BEvZXn2U2MNlD
HWnInhbJoW+3rszLy/0c8evH6pz5IoDgRzNaAZNx79HgmW+d1s3JmLWDE7WzYedGN5XUjiHIGvRh
5+0bhwrdtA3AgWxpKnKJ4Z62q+5rqydGg6l9G5RkvG8aEJGRl8paDioQKeOOlcs9SGmzJyw9b7mR
OjBWtixxtpJtj/NVGJGx9bslTJayr/JA3OUERGrlZ7SwvbxWN+qh3wlr1aXN0JE8MU19Uky3AWKv
x4jw6IVkRng9RGbLpcHp5qUNfQh8KPRd2oQNMjz9341NNP2zufth7RTFigjeRLQCA3KcAEEb+3o4
bda1O9JiudGJQfaQmfmQbDdUMeA2lH6DBGQXcTUgnYE+A+vy8t1tHHp1ukBYcY6NMBqVjz1U4GMu
MsORg7JmWoje17LyMDnQjn1Ug9hIDnU5deonU/CGAhKzuWe07tAkPQpKId5tlSoxGHYGMSEf9R+r
xv0FqMG1WVBrAJQNH5VCKSvQfaEPpxNYbP1luRStxExusNb+m3ZLzKCsuVeqmLLTVe6Dda+1hvUp
8eIIsviPVKWQr9SVGppqEXccNc5AqjpZ9mpQEjrV6wkaffc+2R65wwZTkHyHsaoMXqd+TJt/cTNz
4EYRyDQWPl7fNTCgGWyK7Tyc+iGZXrm2BFQSeKWmbx+Wjtz5cazUGQXyLRPQjwHVyh3mcUOuihBX
FhSco/L23M2dDjcgNTGdt8djk0TQKFtH9tf23ZPi0C2iBs9zVsvtYlJNiLuGBVOEfjiO0LFEtVpy
seJgMn6fCQYB2odTT/Jq2WNwXHwAh5lb5lrUeBu38zo2t+99UJ3PzYy2dZx9+ag57j8/gAsSkJBm
ZNShLvRZIF9wm7T66V4FnPZ72pzRnOd9S5Oy5qDhQycZNPVCQHiilXGeHbkwxXJOOtEPMdIrcJj+
5GqayBqRIbDqIGZXcVrvOmxOIQJ8dFzjAe2QoIyBF2/+1N8M54EPByz3VqInfKyUaHe/D6aJ/Md3
aJdOnHhYhDPO+cImYmIQl7JAWQ/mCC1lhcZsHu7Ija1IYStlMcxLruKgwgBXvE5J8rovyR82ZYt5
QMiykzOlbGZ1RFBnqLIh2cSJ/8MY4NkKlI5VhAB3OGp4c7FNc8BO+VuLbIOa9nrK2QPL2m0w2mp9
qtkF+b3HubIjscg7VSXfxSrD6oieZNrxHSbcuNDx2MsnvFQ9GMuQYmuTK2DCL9IT72uGRrgepVlE
UUXkvZLcFNq70/tU2AeNrDiFH0/8Q2mbbfy3M40kWSQdMMe+XLaO+sNJ4gtjTM6edKaewpBjgeIn
jI1YgvsWm2HgsDQE8xT2LVELxFEJ3fz1WME0HW2oUhaO4cC2C6sNqM74FWZVz9Ie1406X5HjglQO
wiC2t+g1DxmfoJvXiHkTn7z8Zbg1g7efrGMCKhPeiCKbYdSe2/DYXC4wf/esE+pS9T6/bPd8+Zk5
/p7lw5HKgE2UcMbDFJgAZbe2yZlBlG0QCGafL3o0SNoYw2+KH4VvA5XEnhvWewS0MZ5/TeTOk2RS
Zg7kqCibr/P1dsN3j4CW/gyqr3OUeYvk01iKSucvUqacIKEKOYZdA6l8DMnDYFguq2qU2tO08rgD
hKAgaDCIPZqbWGPp3AgLduQ1k6G0AHHPlgQMP9zW2gLuBzwZDGOeu+h+imfyUi6uxhksYrpGmgKu
3PFeBgrtLKL4t+8r9aaJQziOgbivw7PWCpN1HLm1fJSS7f2Fds/vTjtYbglLwmGuHyzQAOe1p8Hw
wE74UZUtv0vx7S2nJ/ArWp6YgDtYapxQgvokn/GC8yRj67zbC/krdT0nFxEIKLPc3QskjPqiZEqh
gNPoYHYOprKA4U0wLycf4zhAXQWSKVwnr1wPWcYP8B/S2iJSEVbhBQizSttnHmQUAdwDPIZ0HxKF
jlQ13JrHhumYI3hlLy2niPjIzknaDPkqqKnHXRtjgWDJk01Hn0BKzk9pkf0YJpJnnRXG43dwkpf9
9dBe0lO17+hnhjWPhclSuFgXGIiCRSPO07KsiBMuY0wa/dvQAx21u0il2fFeGfHubclagHNoRiFQ
UOTHFXZY73GecauQGBVshhVwioggqNwpxv+hn4G2Mo/uTZVoCao9yb4seCi8zAzODELjo+nsA/oM
ivVsjOv1imb0evVIa4wu2Qgv4gCSziXvxCRqxfOdrRCbEOYOG9/zGTnP8glPzmic0+BOM1HfW2bd
ECsniF2leXymHT39y+KJbFRkxUXA+Ml154GO5+9SB4QbDHevEH8Rs6J8CrQf+o35CbOg2pKk6CrD
RJxAY8+arFBdvF08YhTb/ntqu3HPuEhmencDvtambEQ/YylToe8zCUUE03ogZEKV94zmOjfyKsve
QUWUilSs+kZ8/gFWbeVNZuzuL4Bn6x7OXbphGirPgOtR2R8uf2c93CmuRPocJNfQEinCgyFPaVX7
mNoHNt+fn4z9m+NPsOiQFCIEgqxIzyFpR+HV91r2P/gVWqXkkOZiPgLKgXZWJGDHAL73mQechvAr
C8xzknajeKgE+zmK7xth50YkCgpFGjWivZWrq3CfeE9ZtYyqPVkm10rZmuCpLiHMOGQouSkan9aK
t+2wzH5zd5oWSqFZMR4MLjEcqtKM7WVwM2/Si5nBOFwNQJVBcXGdmd21IrhWR9Qa8w/lJpTXDqWz
XwljRumZfDHnG0F2tXrDkTjYlBp3BJXfnmBLG7TIja0RuIobDG4Xs+I7aZRWRXhiVDpvckJdMZ/V
SVQ0xbPPyUkQNVkkTUbGNxp9DW4SvEHqQE774IYpULbcH0Bp2+uJ+lWWMSScpDRSlx9SZ6HoYthl
I3a3hkddD6QUloHDEItUA7jBnBC5+V7k5cNT85cDjzRiFqQ84GDlABJBz6/SGuz+5+dK732EWfza
8R6fhuySWIcHTiPq7s1bRG85YzTuJhFka1kgr5OrHaAjI4lhXLsfSsHN45u09ka1eUiCZp7uww4M
1jXKoBpUbmXkl8O9skJvFhJRvSAEQlf5G+y49AE9/4QCglr+h4sM74usV2r33aEmaL3C2uHfCeeu
Nb4vRUsN2uuAYEQiQkaYxGQYixusJazbKMZ/vQtqfKJK5E9yIJfK8NvjUxnxIILBRxfm6xG7NFu0
En8ee1HZd93kY35i4FrZajT5jvilzj55FEaAiLI0Cnxaypc9ujEVYqwD26SA7PX69VbZx/9t0jKM
FkKJDmsSdf47KYxXdSucW30NJC/IXYL6+b+7eXUTCS5THRKPnark4/aSObVoA2XNGAq+VvNpJmEv
1UqngThnF21i9TRRWeMcWQgoHm6tqgWHOzif3CII+UKLGQSoCXy8R/lJnCd40x/iQbLwmyPUAcUo
NiWd7dhFYhdmjEju5ZnEweJnR28Wzzx6dV05I5DddPUXM+Qo7vG9lrfpNCELLOHHvXOwcnd1X+01
uWy/vobqrduhrZoR2x8oiOqLq7BrSW2gDk3L8mjooyNEF3wGiiytcVgcKGexvPKzdN6+okFkArEC
2h3fPNQ9XfaehiXAZulZ2u6EZaEx7GUDrmraPcfYyr0rMbaSWu2e3pj/5pH1ahJOv9gl0YLwOo7a
bczpg73do8VtxASI8krOgGe1pKNEPW3ZnTDtVpr30xG60vXqd1FbjakEEfFEBud10KQQHZej5+FE
xYEYJOJIJPfB31nO5OIv7elInfR8+PMDaIy0xCxZB7tdTzDaGPbWO81o2IwX+UdGAgNEW/yHh0JF
8METt4hOQ212Jdv0tDzLRLHH7hJcgh4pEEYP3xGlxfW6PHoS/ML8ua3YnoXNdlzwf+amnlcsEllC
C5d3Pg/ngnFK2lSeDsIF+OoDrpMZZJFtT9jyCeoEG2FYM/9sQ+UNsL9VGQMys3+fAuvL8GNzptVO
WDjb7UlkXESoj0dnO7JkGjYjb7aQnXWaLk4x5MvgVmYrwjFk8iR1pKNfR69aOGP/W4LSZpDSwjvH
fSQqN4iwv74btaHvFclRGOoMlSEx0VkMbZh0coYNWwd4G5LPhEMS/IXmS3TRsIMk/S1Lepd7mhw0
ECAT0afj3sr3oLl4aZZMOE1ooB39SoB87zsWrqtrxZVQQOvTbkGq/YVCbZzTEaKQwJTQmP3KQ5Mi
rEmIw83Gz72bakm++d7vLZXfTZYxm/5VG7ryio2IrMNYLanYe+I1fPoxzCJlPPQjK7PChnZy9Zx/
PD+m2Rly9lCUyTD2E27kliXDGo8h+a9n27O/1TOIragXn9pmrNsxTk0vYPFMA3/zAUh1JfEMCfWk
Hl2oqQOD2LXS2K5yDBx4brkdf5IfJPsC4ihvmES444A1ij7f9zXP6mX6RWQKrH/QZv31pESt/SMH
McTpww/ek911TUpoUKiH61ASY11/k46zf+hDcj+1LNDifff9GXQ0QkhH6wETBPnpeAV5F33Vxmd4
kOyWBBgGTDlb2qopsIVmqWHIhNV8xjG/1FznebMN+n2nFmFp2OlmC6JQNxYvBnECdgCgFYiunzu2
urLv+iYjnoVRO+myxTVL5ZN6Q9zFEGvCWdAfvtKv8saXeNTDGD2xH2cs56DufNnXANG1uQu+tx51
34ZMP79MbXtEF1OsQJo5uEX1XOFnHePg6Aa0xwgkqdFFixI/9QzPtpemzgM6MEn32inl4V/eb7GQ
wXTCmHt2QnAGqsrvdPgagzMJARWxtj6Ju3hFOvfGY4m+XOsQObmpMK9CQaAMaHjiUHNK+Tkl8YbF
s30LIMA6P07+/fZQtT59b+KQVAwXUMjhpm/PVcMJhqL5naTLJQqbgK2FbmcFcQP1CCvzjedlfDet
8dRbo3K4brGdy9FjVK4P7l2pckTJXJe1WicKQqge2++X706mZh8KBdDHVZdcXoNESC90gd+KolHP
IzXDH5AN3vru+sn1jD/UYJq1PeovChhX8EnW+xSDLjq1jok8JH3Ba3gzztQK5uhOVQ+64KNbygD/
zsabPRKd/bEdOce9pMKc9p7VG8RJqAoRbaftsz2SwMaRZvKkgCKEsV6V90DudyWOvDAIMBorczmq
QrTAd2hhTo2lCU1rqoA5AG8y6k0eO4nUrEKxYgzc2GPUWaJ56EAZA1s+tU+V24lx242QQ7dQy5Sb
RWsi3AP4r9LpA+gL5Bll3FilbHNFgIX5MPDkX4bGXNBnWRpr3gqS+lAb28vFD0oljlJgIPWA7WZ4
r2MtvcoKTblHLQ8kbL8o4Yw3yjewrwLUHtYKiSN9eQ2MZuP13jKtce3uqugndfQUf+LCMm1BNQC4
mbaTtAOsxRF3GVluy4EwDjbjDJcqgtH5kUw/9hVNnAYX/+X8UyrL86Rq7nN1uJJ+o25w1n8xaXKG
TOZ4z2e3PDkg2KrUbJnQWKRY5xP5XGv8cwDWDQjCr+zhEoEXXZUvjlT62lkcro0MSzyYBhaKWtJx
YqpNcQWZspUjvK60mzdko46wbPeHZSLvqoFfqiZj9w4SFAINxRO+Gh2Y4V2UbKFhwhm7WILOefrc
MKxiFN7+SFCcBp31dwf4jJXciIiFfDhyBqftQYjdD/S7pUMBg7H7NFU+siEMPo+kVTfQER496a6t
ZszYprdIjTc7/+K91JN5XyU2Q/L5BJeL/nk+NKWSU1R7Y0awYnOrip9aVFypAL4fxCA4UPLND0te
raddu0O/y+Ima0lJHqRm7QzE7LUVQtuO7Pp9cYvA6EqHlbp8e4ZW+KfYnUoVJE3HQEU/CMvQ6Oho
5wkbyq/7KrSldKKsCNIQfIq8f6FpWl8PaTyk5HWKOeDqJq2blfK9EuYKusFm0WVWz+L798UN0Y2S
fHr7yTY1Bl37LDcK6EzsdslTh/xF4+yFTeVq3D//lP2JTl7qFdRmtsgX3OdpExADmNgIl8ca6NCa
A4ksTRTLIncgg8EtRFq5/OolfKrkaVXLAUjMaXPmGClYj1yMWQp0GGGrZPsmNbm62nU/8WXN0Wa5
0CebJDJqsuFqsP2Oq2fUB81Husgm9RpQ9gK3IKnlcqKyp+7SFp29r/dncHX4daBNDWHILA/IOhMP
A5EF5XVjj84Qx9TAVGBkhbRbtLMt0YkPsAS4RBgefqNj1yMqZNCaJNUFm4fJq8lnRfpDfDRGa7HJ
8aRou0OnNTHhmymLSvW8Yy5QbePKl+zlsczi+ox1UsL/8gevKHSuN5QbrbzP1XdxFgW9bwcRfvp9
LZeY4gZGNAlyzRtaJnFJ/jAtEWTtwslirzgKpewCnIkcVWj6fZYBraRryFgKrSQKyMxQVzKbUykL
Tv8Uyt3Qpb77LWV1BkFs3qHgJ8sV7SKJxkT4HJ8UHkRJx/zWqxNHKaLy9hdoD42YONA4bmM4knvW
2WfRDAbgtapj2SS4PsxhxivzFdxYQ5IhWAn3HIovosgVnDBL7NLS34Yf2EDEfkpx93ZU+B3+RigS
fOQ4xAuHtUmEZPh55Oc+SWNSZrliCPI88r428yNRxu/wmh9A686CfKwg6/Zi1mKcHVyhRm/PuJO3
93zsWIn3dx2w63eiWcedNsrWVMZoRXSOcwxztLHt/6goNpUH/2Ig2JwdmMZF7embRIbxsQnu7KKD
+LhOxMUOlFgdaVX8epAniRaBS4UzyykVg4UTmz8oi1/A8rHf4uSwezgvg7klLTbSgKQIsCt3J7hS
kuWUZ6zXlMJPuG6Shrj0jYDPPN1wQvwJSOP66uK0w5NPSedFgwPyUewefMtPjCqX0aPACs2oxNwB
8T5/eg/rsG7GOw/rDB5Ocx8huDf4H/T+0y3n71QcwB3RmnX6rsLtjwoUda5TKswV4QOEquYODzu/
v3NvusarpXfno/zB5YL1FoGcwOC0SIWBD9ShPbN7LQDigYNUOsVNuFzDvbTQYJlMglth6huIl+eo
FsDrueXMGHxE3JrsYDRqFteK6mKj9uu0gOsvyyBNJzRmgsfAThnU74VbctYIdW7KK0BgfEOdynUq
hmwrUyVmpGQ+bo7/YADb7TF9rtkOzkkAUbR/hDFGDDOzCv/M+/GZcneTWJclENkyLVgVRo/hLigV
M+fCR/4JLFRapdAR4gcFVdvIPWu0QEfrFqK+bQxICOOoMYgX023+uWke0Iz2ZNBOeh2DC2gl1Rer
poxzmRlHhN+/y5+JM1GSfLnadzhh01R9+0ZRgAGIlDcm4wq/2f/nNo/Ee3SPRvry2lmiFAq7lOiz
li+ryVMPYaZ0aJb4oZql71El1PZ5gbwuNFIxvcnrGF2xy3pI6DZjziPvQFZ6UfIdbs1GeMNGnNJD
BrU6USfDOzZMMYJmABOiBeDfaq5R65ljFLpoFDVNzhEh8g/njOHaOV8BRuWYMuq4ilKmNb6zfuEu
YGb/Ssn3GYK6jZzny0G6WfcQ33MMZDLV1kUsuwZwfynP33Lt5AV+f0+H0MHp/9rUKNsUuyXJ5z6n
4okenkxjEc3mWt0rOgCxEWk3dmqOxtYsNUAEs3u/vI3rADzjhpchvH3zVuLs7aaSgmHUU8wv5jr+
woTm4216/+4IQnkW4g2CLJsY6m1wwTiRCsNi+BhEBT/x3imSe7Jhxa4T3xabEIHh1jBIkMaJ5pWm
ghOVcMsX/3HRJzfxIs2cJ5N8UFY7Wfvji0xZLZMGnE+vH4Gw1He0/WJPf9dXHAM9MeWqt9jz3QmW
VURnZGP7Vom6zhXLfNVhpgjlu2OmU/5kXnBhywIGyibpXElzrxhGpsQkDnDlamrfZFUI0bcPUCay
dhCkoaG+L7/jd+4fkNwsPgj3oD/AVY589vtIX34D+w9jv+wvEcdL5QU42aIvqTQfaJkzCIVEkNjf
YljV9LNQOU3tVPE50kP6Sj4aIbCDx3maLcNhC4Hp1YGKg1VQR0dWmAdFp95NeIBko7ksR7uQnlVp
rHztWp3tHJxGtx6/9itLWqFSZM6vg1hd43owliTT+Y/N1ctGPTT+ONK2XWVMbny/Qo3eUV37ZJDw
rJtuORkzD0OiHzCGwTpjbvNeNTak9PXpjodYvwogq+GvtyW1VMkEVtdVpSoAB1bzkA811UP5F1dp
uED6UmdGrC4l/1NdLAo2/g6l0/Za2lEQd8DVnt54hsXsu0iUGc52/ZP8FpsnQLi5nqcHG9lMn++j
V6NOGw9OIog9Bjg+OlGLSCbDyZN0I+KSeVP3d/QRJIPQsePvFdX9uuxgRF8kTmPF7HoX9n9NCX8H
jClggfCppkSv/tnHTF1Y42UX3zEg772+UKlzD4Yvn8YYPngiX5gagRMehy0hJ+u39gpRqo0Dq1UE
iTzhvh+lTci4VvoLxeGtdQEs9BORtsXc6VD7hQxgj0RtoSQkNorGP62pmEYxSRM2SPPOocsYXRoe
ZgCN5IP4h966yGNeDHP7hssiad4DB0eidMK6Yn42j1uJmMAv0OsuHyskzFJVcd7q3GdxRU4+T9sI
L/9pY0Y/ll4NJK5Wy7WBFJlLisKv8AjPqdRg610kqj3DPrxwWDd5SKeYyK6z9oQ5DNq0xCX6fA7/
YgFWgJzCKgc6STiIMXXOb8MxISiHNY7wcUNwy+Qr+RRclQ0rI4rYRvNynkhH/hbsH3bKajAx0Y/R
Hjlwqzq2hT4cY7WkDUXF9OH85cPbMUJHIBxPpQQe3/oUASJ3a+2UioZyN4UO1xpCatrEpNB+LIKL
C2lzJIICMOFKQV1K2CVkhN4K1C+rCv6FPG20Ym+3fJatkBhxew4eRK3t8g1lGtgvlTbm2FV23LqX
Of4a1EcEKOIY/4/d+yVfqwXLYq38eZaKEq3Em/zATvXBoEoAp1iu1xYHqP53gAULnq5jZSFCtbl+
je5vO8SCh2u738Q0VaiGsu3q+7YWrvBYqxzLVfCWw8wDO5EeCnl//U1nV/XAEjqBJorVs4BeLhTV
iJA0GNW5ls892KYhyjdLwuga44PkLeCRipvDzNhdz9fPbeTVWrvqtsYjEy0AcSaujfYKBYHZpmPx
D3HxS3J52+UIv7mWBFzgk0axVhPGlwokp7yuJdxkFMIpUWRuG28fr1EnBHr2rnJbcamLeewg8pTc
yGUNiJCwGOyM/WsKpfklnBnZQLyLaq5gyQLPqXci55BwGBC3bgqEPULxZv+VzDXJV0Dx38W8CQPe
FhaamBxhPu3bfI2woVJGqHClH+po57PIz0RRL6Sb5TTlfnI4hFNtvR6skZDNeev6ajoMNZ/1Ho5d
EsfidcCAgOxl0VQTOmX8hUfrMtTAJs562fsr78blBpByoc5pv5mY+5h/kiHgrLqWHHBjKIeyUNaI
WvK6fbPHGnfTg6gYfjSjbzaTj6POyMpCT2KFIlfPkN/zrVZyJXjybtJknz5vQb9K2AM8bMnybCgA
Grhzy4APclYevFggjn6PsjB6xJU5NCW8e9Y2YOE5SPWwpuO6uwwGBCd9T7C32bKUaQXhsdlzGJdD
JjyUOXuTr19d77QPgVgUJTWRTG1bPOw6JQVA7eh/2nCepWjJde09bSJZtGWVBzO5alM4INzl0dNu
0tYd0oUtWlhT2hqsrZCzhqQP6GXUa6X5ZxecgIaMzecb+e+UiCbpMxqu31erWgsvnAVN/RF8NxOG
8V9KzZ7SmQx6zNl9Ab4eIbCvyCMikIzv/3dQ9RnvtckFTIoKdIVayrwkDkLzFIrsDohMNqQLhWGd
abL0HzDtOPfh1m4rszxeciZuDM0IEdxwkUxb59rZ+mmS0wj0wVo3IIBJZ0Z46sgt+Nf8tZdjDXEn
iVIt19E4hzPohA1ZaanMcLNQo9qDHvTMq3HkyQRNUPkisN4sLPobQqILEF3CuXuHCHwhK5vEqlbZ
/je/LGcVvWsKmK+98N6I8do/yZvj87oYrzjiyml1BsIeypVGcNG2thtpVGJ4vn5jmacBVQcPPLSr
iqwkAEvEal31gecByjoE4bFjlIvd5C84AYa33Grqa2mT2XD8S2oEqUhdlbPa+nwqi7dIopWvphsX
/5kG/U7VOcAzK4v5B2AnR9uiQ1E6o3RJA8ROTWgZ/iRRSZ7nvxxM0+F38YbVDZwL4FmO88mh9kDD
0D2XcERrKUGIg/4cEftbnsTIJjT2U3hh2sFX0MtaiCavtSdm2rt5k59TQHCjdrEqvaCSz7uE9WjB
S/moW6LMXVtuw6OR3lS0CCVvn8pPPGqkDBwnNFxb0bPIzTbUbh7gTIhtMolkB28P0Wyv1KIqe9NV
bdz8eUjUocuUuifZkeKmFbhdG8o628vY8LDJcyxC12dPD8F2OU7cGSmWi6oDa4ri/ihxsA2HDBQp
o8yhYN1j1CMvjYnu808mV/Ucm5Uld6feBBLVXrdZD9xVKAhLfhDWalxcWIXCMs27FFgb1yf6Zp6n
SVI85ouZvb4+7ns8/ev6EzjoXuLxVqljkSCmjC1mkesSJeFW8nSwr4kxFCwRRgcr69nrFzVJZwu5
em/Fn4WfGi4b0zeWSiRq7H+BCM0WOJ4AzMguleNNpWC304YDOKbvQiW7kgvFRTb9YQmpcG0pq1Pi
NdTZF13xkX1TEYsFyFcnjVaNtHrYaCZSCm/z37SDSfXWSx1J9Jpeumr0jaIOrgTkPNi2YF9RAfdH
tK1VCAitytZVaPYlMwYHM0bxwTlcNtTmjU6wi3Lbf/uhO17cmqKlt1WnTtaWFl/T0PwBMjXdbq3e
r1WAoVfJyTmELpuOaELozbpmqPnhxjAUYH1VMpFJePwi+cTdJ1U5SNXM8sIdXJ6LhU8gBkYQtNhk
6D9ErpFpnlI7O30YUo+tGsaRzT2vESh4Q/auIQMBvZdxkXuWV2iewPVlEARScKT6Y0TknFOdMm83
8nTSQ075toGeC6yAxv/uTqRAcueDVUDchryNpTX9obdqfW84ieM3pCWkY8w2KQh25ajw5d0Y6hZj
J7XQJp48KSaL4ZpDeFLYoaSxF2uyBeC3Za9d3zW3WOHaehO/h7XeXcCACNrPvpdS0wtlwshfoUm7
YhUv2ExmbnrydyUKXC+sxEHo/S+vEyWZTVIoehsopO1RVH4d3yj9qQqfEJij4sF/26IGv/Wt12vY
+7gEVix1068Zqg+QsfKFTe3Hr72My6js69agNTkWppI44jzKfS5N01q4fiTNDk+xT2xN7EjvZFSr
oxWKv6H5merMdZ13KSi6h6Abgb7XhspkSv6yoznp8b7okEzE8SrmiKLKNP5kEwuaDqJxgr3ACipm
WcweyfaWkPlA2y6r86r4rE2TM3Gx8O2ulR8mFTLeIPNrfp9a6BcllpTwIztTMmCjPm8BzL43tVxB
rsckOVDMJ3X3jR+soLp2sRwS2qqw4rV9xAHwqnW9adkkvfAeKW1f0H2A1NXL3NPOlwMBQiGtX7KZ
ds66Kcr3YOcLnGGAeY7233pZrvaYwbgCLihzE8om6G/dDp20GKObwLK0LF5K9WNICo7prPet5xVG
zyo95O5nEiYi2R7YMQQ12rapQxRoC5fbl2C/Yn6OPkjahPXT1O+swQbJusBRsClqXy+4hs9hBtYN
uv/SgVEbeQT54Jh6SRAzSoMEhXsLd0U7bNqOJxIzbhjUqtWsS/E5oYEU/YxkG+LuAMy5zEUgpMRb
1JjkqoTELyATBCWIiVhyPh9vlVb5/57hlAUGQjsmm6lnlbyqd7hQ36BXkDAGqatbdqH9Zm9bgzAb
X09CSp/BFww0/BDP7UV2lNGmFscQhe/YW06wt5g/0VSODIkAX4/HUqzGX9rONYSd8U5SSk6YrBdz
BzT3I+mowuGNNerEAAfSqm10VzN+Vw/OYCvTW9BbNCR4+Dd2ITdhXnXkSBt3ZDl0qC1o3TBaENgc
o3vupBTmU30u548rm3m/qVcyfFrwFe2zHeYAlVG3MSiOUuFqeBUYVLRBB6m2z5fzPJXXTOJNdehn
vhtMXHEnpoymzsYQhzZFCQwrzHTVwuuFd3MSXCYreqeVYIEs6QSp9+cJ+ZJ8L2USnG0SUsnbGLIB
Si4Tarz8/HfYFjUssID7GEy/faGydNXNl5GwFLcpvRNjosew35FIiOBv20NGPLEhMdJVrut9+qYj
Z/wacwvDc+JbMxas5IA/Ul4gpFjts/Jv3yywF4Aub1F12KnxXDQp1McUcZ9y08Jl+mGJS6+m8oKS
svMeHzQuIpSlg38vgE8GtyDmb8G6J93rMsIfD8NkHeqFLPRems5MLtvisLP3X3gBRK4DsrEhKrcB
L7dY50wtObNGuGVO0qMFA5YRKDCeDcfoG4VWaRKdhOKZeY738Zq9TqAHESjoxgmHWmQhcr+cw7MV
7w+nvk8PDXIIwvn3VcDJzXTEA37T/Cekg/9zLqDT20/z9PzXjb2ufxzEMH6K8Y5DIS/XSy+FGqnj
lt3vGS4/+NA3KHJ8u9Gmax8MROIXJZMQkW3nsahA3p/LR/89/jdTfaQ8oBxu4vGON1vobZCjVMt2
P5ZWNso6gE6hYAQO0EpJOxQ7pZ/zSNKktxJz25Z0vofe1YeEBg7BNrIIHX7iROuXmH6l0A2p1W40
HpSWSJtt6Bf5ziy8RWX6fGMm1QRN9471l5xAOBzPiZ+Fc6ZsEXQH7VIpWJk14Yciew3aqT+2NJSo
nVZpmh84i0Ibl8+FQF4x4dvssn3XhT8J47NGRdVokllcDJZvQzU/ARP9v9mjOXRhdFv4AVAqaOgO
pacMrsZTCwkKYIU4+zINbxPkQBJssXh4k9+HbYYWKnggND6NWTrSphGiYEm08FfA6F+S1esZk0hI
afZA2dZWBnz7bkPrdgd0r/J/7CZ5dQhSDCbKmj7ssdRhfATDEZ+pMZp/XUY0ARac8tKzD93nzAwS
cApQW7FBY/8N4eae1detM0O1tK32w/5Ew/26NJq68TQig1dgsHWZtiMMkrFL6Ifr/kOKZb1NIXt+
vdkw5iyCUkIftA9p9M1ctqlwkV4n7fjganL/lyKD9VKQOl03dp+dzDmMCkaqNWQsPuq/t2pWiV5D
6YuwYtsKSVUz4aaHfmMaxXGBj7zdPSUSGc6ATC4hJmdqFHqAQTcpxXYRNXajxomGUg7xcNxK8636
ad78U0FA65agRDyyIsIl4vhSZWyQt8rEfGssWEjuk8MxuBAdOKvdxw7gnwVys5NskhKpvohbvu3G
/jvHARmQF0YeHv1SZJwguDwSh10w0pve7nhgBVPuLOfYCu9a2WyQwPAbkdojnoPIXaOHB2mObV+g
2l+/cHc2xdvhia69V+TWN0yYG6m95RQpIMhY+ysk3F+TpVwBDz54NxfRXpAi0+h1Evf7PmiFrd2a
IJacYLqSKVfyHOIA4EhCU0ES2kT39G4TiH62L8M/s6jReNy7ReJ9qzdwP1AaV12QVvHeMoizxP5W
/jkpNP2M4E5uV3Hn0LvqjNUTfOhPQxniVETnpYd3mjgkqUPl3e2HIRF/ZeIn5tC+uxsp+5pfJ6e9
iFPPSI2BBXYzAGKGCl9Wem5E4OIdgbCO/CcABo2HX7zONIA5KpgtBVEZCecD2BPqT5DQXkOaMc+2
DGiPOB//BVOqNTH0XBoPt/aG4zVvZzHHUNnXvx8EGSsD9/BD6g1E90wG/Q1V3W13ZiG+qj760XBR
DQhzPV/829ayBGqc4teoyLNAgMFEfpPsDKKSVqqmjDy+QtBOLCM1ilVcE6AJCZMoHrX/cOGXkDq+
bZbl4ki7WxN08TUruPvWaAAtdPW6zhTEAUy/S8G86IewZCzHx7TQSxWhYuXRWR7pOcw2Zve4TDpT
TkSL/1jNsVCQZYhZqcP29ZtmrcxVRrIzTHm4/Fi6E72iv4N/PWYOn5mYM4jZj/x3beEVBd11qEpW
2agbTqQfqDoryH18wMVceKkDlSpejcZSkzx99FnIM68sElq77g6wD1jbiAAP48s8UHoZp2W1NykU
1ay48UuKlaE3Jy4lBdvv+P2rSjnOO2pKVxPhpbiitzP0LZdGTGY6E/65OYxCBJ7q+44EywyS97Yy
jXpDPkCISTmoYz7Wt/t4MxgDPQiJ43aEl2ey1hRZdwmL4IXDR8uRqpeH617cF4jGMgcYUd+92+WG
3LaiA1Z5fL35c2cpXYS9CMULX6Tyw09vr8Oo8vDS2Hozfi8jEOZdczLb5W0qxpLtVJLqKOfvaE2j
JSzlUCW2QV2z3M4VeZNKcLasEdUfKI04uePr8j/pvnFbZUoPa3vW2f8ZlM6GB+mOowK72aFl65Dh
s60yYqaU0ufqOhto1GVfx4AUW6TXZLN17fODb5bmWFox5IJdSRe6BY0GoFlkxZX9nmeMFXcXDgRm
vzmPr9d2L6ygm+e7SpNUifu8L5snO2A7k+yPlvjNGPTF0FruQDAf9t425fmf6QQa+PuOsRbtiRg8
6wspajG1DC20C0kI3yLbqXV7ZQZbQgELHdiDhLPw9pg4EMqHcIx6rcZs1iumarg6BoKDD93bgpza
/8sDa7IIBVuaxQ042P3wOAYMjbDsa8J+/CnCplrH8Wutm/fyIs+7lpkDVZlW4Duicun9cSpZOrg/
GYivSxy9mxDmEEUGoRE/b19wuazuXFp/p3M+l4EHKahI+LFXW4zuZZlFHPmKuTznlfzEdI4Et5wo
O62MJiy+zi+s2JDL2db38iG6JC/Pu5WEmWRWY8y7YaRtLxQGyL6oOa7XYrxQ3iv34+cIaAtMxxOn
gD8C0EeyUS4VdPK3tqIrniHDI8WIxTuEwErocq+KOH56tmRtPBKgGVYEOjuY/R9N6e7aSrtYYzK5
8/P6L/T5fKCRS1t75gDZpFYd7p26ioEA48EuQaJazzC5FPhnjIeJljPSD0eLfIdyfB6OsrY5pPno
2lPdaeOychbAdQK1eIzH+qcHa7i7/C2XlHafQUzvpHQ9DlVLw8viAmJrD7u5PIS0zMXMhHBKxBaX
lQYdbr83qXAyGMihlQm9+OCdqcIlcYgR9KuC1wN/PQGzIyRnH5sqJRUhpUbRI5ElSUL2gpGDt4EM
p3Zfmtc35jQR89V/rVXAxl9GYIJhCJcobRYRVPPolV196p11s8mQ7oQgJwF/fRQdpUF62h+uMGy6
S7XrCo77PMoGMghHZhr5QX2GDiZ7htqTCmZWuzmJzq1ehmLJVTqiKjjEuC9L2z3r/Re4hipi2yoh
XFPesb0TmPVpyq7I3bGDwUZWYFD/arJA20deUR18zXcO+6j4wAE4nZWcR8+SaFRmwn3PyUkZ8ScC
6k9cVo0ZpBIBMB9QXzRIYdg6nFTUyZbXVAz/xzlvS6itMQ0EB1AyzfwSs+rQzWniFpK67k+mdX5c
PasAoCXh1Ijy390YU2O4zjK1EUQcZTVi+sHCwxK2sNScQbwsOBTVm7AL/Tf8PLXGUiKp/iEdHQvw
JSU8jdScaRdj0caeGCEXOEA4fLs7ybdKVhOEyX7GKtTP+JfXYOUOKVnSfws5IXI5n2pju7FMtnIL
kWc8OP2AmWapHBQE4g8X4VkaxxoM7h+z7Rj2vqW/WrRTqV+sjVd/s3cefUi5eSWst4CjyjqpP9H+
yLX1Y6vjAEOPd2NO2W6g4qceZIPepXE3J5uuJJj93V6T4m+NoCuFp920euLklqQP0L5GVeL4wVDM
UFwd9l/rrgc1kjMS841hCCLu3DldXD9WTMjZvm6nQnkt6IfgtMe6t3Do3iA485nkK9pW+sNApww1
6xW9a1JCgf6ZuqteWaoGsCw0113GJbjZzxWVfw8uHl0rDoFwKlKiigeJjYj4Ur87l+gnprWj98HP
zAzmcKjr+noWv8x9M7+H94da8kpJHZqqURj4DNEHeWQnvMJ4z8bob/xZSfXYNaTOFDJcHcsI6E2y
DndFiA3Y6Gs94RQFOG3mUz0/0bN3otWsEoBX3kFodkHxN0pCU6ao/Gyq0tEDp1lsozCcB02va0eW
SNK2borFYxxLU8R+MVNB4kV3yMLydPvkSfzp8F7adI6eVpfkg9wDDxw+EvnOx1URNZrAoVRXNVn1
BXiIWEhUaY7n8uWUnWXvefAMC/WLh9QkRxI07GkYthshB0D4X7Y/8JLyZzqBV74g+b0cdZzo0CWu
KI7/oilAY4y4c1+FPTkuGmyFRk8QNIskeU+LlZH5IQpDwPTJmxeJJu8PrrOjgFBFYwRu6Cz0Wf6B
Mev+foDsoomdnPbvZ44xSl7iPqIKHdJTbVhmSJyXMN8Iv3tCDW4h+G1DIfmcczGKArL/9rZykle9
ukkXtHmqg/NRbHRBz8hamIux5BSpN2/AVhVHWbHZcY7N9bHUeyxSZXcatBG+AXuczT3jcZcxY8oY
1D4KRm/8GUriBzdeUvuQUpRS9zst/U9kiXBaRxO4MpRfZ/mmSEuL//Qe082InH7FEJf/FJUA7Vf0
0LkygdzbMCxDvTrc1v9WxXRIozPwhCyBkzwaOXoFu/LQgxrqLI1Tqu2moO5LEa6ALBzj5gDaJZ5O
pjkpFefWnidxUZKU8UXMmYB5Nlw2678Z1jexG/D6ZCcURmEM2eFsiUu+5DpHA93c3W91PyebHb+n
6NoLjktWwJs8OMc+/pWWmcUcjl+ngSQJXXZxeDBPUoNNS0HVRjsBOsMqt+K7wu4v3wvNZjWaVfmU
W6yEcwcvo05ZoOquuHXST0Uak7CrWsMZ8jI3ggCBttGIMMmhc7RYYQfl1iVXGK6XeqwTlbMLn+ZG
seJBD6k8m7GNo6Y6vEarRPeaIbXGf7Ec3WV0QbkW8kRyxW2fT4pgi8ikqlGAW39fEVx2xzMtWT7f
O5bpGYP6C86EblSkrLAg+bH1zaw+rLuhnjQo/E6Be5KfGQMN7jJ4aH8NnQjjan1bYWgMKC4p0F49
eGWzn2LL0S9VTraq9C6veZKcg2oN61S544O8xo7P2MftG3GT0GTjV66bJxqEZbG+IzQXAgeqJ/Kx
ygTdHbEb+1XIftO+gznVi+sMmCZb76BVCbjCs1RajpIjZyS71MRPg5RubvuudY0O6Eq+teOzEcYy
ar8f7jxkiOAhW4hLAnxaY9l5YWXvlhXsYluAh5xBn2DF0a2FOlh+D3vm7qAslIRuQHq+Zl9Det6B
G9N0AS8qrPJB16uxq8tB3aCfGZj+E4eMOR1kkoLY4CrhcbL0At/UQOH2dY5dXKt61gT6r0kVxMHg
8rlwISGEKTmLH02b7gIxBkXFrThMDzRojefG8rSKuuuzReCKsY5z+Unun621GVohnizmM1BZrJwB
6dCM48DcU255bS2kWwFt1xOxEZs3F1q0sOEndbRE//n8z21Xh6Yo0YevjnNVPLHGUKqUnHFjYLr+
+iqHHMxFrUDo+ZkMMIIkXgNpVp2hfvpOfomIbCgZKKwdAuhXM/MieL1LvgTr1FDLaZuiTM4R8qjn
HPBYRGv1ycvwGdVb1ZeA/2eCNw/zRVmDe4Pn9zKMjDe/4887BVX90+bYTkl7xp5o8byMBbDzjnM+
hpC26XCljT7K2A+cdTlTnMr3FlifKqy3dUnSmMlJWimxMOndNYbVThqV8hYFvwhwmyGmQ17S2zX6
/0lvje78c8T8tLrO7BbEHUc7gYLp5CZ+GVG3mqLRnA12lvCZPE12kDZvhESaNDhd+7aMMNJuXY0z
jKBQ6mXItOkJfsfOec4Fg4QwqCgy3ZnmFg4JhBzhQVSbuNMkjGgTuYvMxruzaFRc25ZlnBESmF8j
tPFu8eryfX14bMKt+sgLLaKqtJHmJprQ5u4x5VJMRmf/eCJhVpVcn0RjJCjgenOqtoQv9HsKWsST
ySLb7UVDS0ldTmc3dVhiioMbn2a/fWCeP6KX19SO4iPdILsF5fjmmx2+NnM+65zUnJ3/+1flxVZp
4NuiKbnLq5NAwOJdhQHzHTmOuHAo/A+0KOs8Fa+JFIYsiU+wCpPPezLwf3ZXMp0Mn2w0XEWTFk9P
JBiPQkGDNYNZRjBkpESzrL/OWzls6rvGdpJCTkz5P6Y5QdpDpGi7p/3NfEPJoaMJ2Q9NacU2NOD4
wKx+jlMiT0jZlEemhUzQTx3HsMvkv9dn26kVoraM0D8sjMxxlp7eikWLpIWBn8A7YHj65nq7LySV
g6KD5c9FgDzd5MnoBnX+m5PhKOqNuPwSd96pr7D6tpPm6lvChO59OAq5+e0Cv/q09cmu456nWtcx
Ff1hz2qBfd/dVOq+F4QpqzIKF6d2i5Rf6KcqL2v4zji7DV0NXEyVEkmNACcCK+FjYN7JsR4evJRc
v0so75fFoDmtN11QiVs8TXi6zyHOPlszLpQC5xa8tUrV4S6t7O4xSIKpqkH5fTnMUF92qp8eQGae
xdK38xgQsRzZWGeit2LAjhIGthsjlPKuABXk6maD0K0UHr4QPLdW1s3VMpaO3klBs65pqryAoQFe
Va8/TxpmL9e+eKPWBT1drHt7/Fgd3jNChmZLNrSmu3UCL3E+ABfcfgj5n1uSk4uA6eSlHzdL35YN
CJnuNk0JOrafbJWochZQPgYf+q6NMURDXc1jwC+Ybuvr9rWxKIIzxeNYtdUmTazAX7H7byXMBYnq
uTDCy2a2QK3GBEcBMm/MI6iSaaepUtgQ9BY/iWE0em65dbybV0AHTWmDw0SkVoGaDa+0Pb4j3gNv
wvg5MjuXaqxitlLbCT+vgV8yXkynQ1TeJbfUvJgNBJ+NMAqVBh4AHOe80a+1nQswGwAh/PoZTG0K
VKq32pgKtHO55F2Vh3Eu+ocgKfZY2uDtdINN+tcFAeLAU7Au3sqG9Qj2VITDmwei0NfoI5meBz2w
0p2kdBSb1dKcf2xn53To0btslM//pVOcPWvDTBTahl5mEa5SbR8joW1YoMBRD4PUSLZqxKNWyBFC
KAcoF6hAFCCrsm6jsUQkL04HVOnU5yIgk1nDfvs7a7IScKqTBxuwTfMXdQHJoBcsvh15IHnequat
Yf0cu63O8ataey4VRmXo4v1o/a7hLmMF07NMXG6gUHp9BVsi4+SsalO+r7HD6Cogsm10sMYoQ+sb
UkE8+7XYZzqx1pylJuRwZXjS6GNqudpGKijwnRycPzZio215QhLbqM1OaULwiORjkwxTIJdH6teo
58ltudXpUH4tGU8uP5l+674kpUH2eolTeKaYCiLFallfQXdQ/2zw7Ba/tXIlZXJZllOkqMbG1BE4
bWLXS86BVWt9xj1mfTZooBtkAPrMQBYXyS+dkRwWWctn8hj15L5rQkr/COgqjC6d6h1KHwIbzlP1
iEZqrUA4f/aPIPKZd/YKic7iKpx8h//GtgVnouBMTZtvC9ILSin2/GN0D7g7DhhbmPVuvW93EAR7
mDrWVcm/YLHtGwazQq3iTw31aPtfEEBsCdu4aycOS5NHt0H1zxzetP5t0vlfjVbiTuN/KGwghQSx
OOmNgHqGx/vOJynLYN+/cUYLXs9b8K0hlJfCh7O2je7A6rGC/mCyg3znQFKIdDjBpq+gj0ixY9ID
WCdChBBO6N/SqoZ4pXhJ3F9gLcM6PeJYcbNwuWEm7e8W4nfW3tNG2UtEVsKrq47pf1hJ/gTNigju
3IyuYdAz7GFeZGLnAvw9UGmuKgAHn9btAAb2YOyYw8EdawZDdT1DqCNnDQLFsV5qbFJl6rvtH3Zp
mPvVOaMLo0KhvloyAkxyeIkY+iH9Nipkv4NxxGAvJxiSajECktY5ZJ4Eh5hE9fBlOILegehjKHKi
gTPHNnOR4guIWIS177cllsVCNfwmJHG0oWshzPkbRn1+42kxftqwtgqwP+ufZNC2Zr8Qc9tEvvJ5
QbVax/pK+BhAhB914h435Rj7cinRi5SU7WX1FXlbQvpttbVUTKnr3hrqhqf66ywangt2IZqAuD5I
GILynxwChBXcjSEtT++jRia6ByTussTw8BftTBMhAehdqIfLzHPqM/EyC6sSZ3AAmKdw4T+aYmH5
sq4EKVD3mpPtjfJySZwZTOFmieiwghJQz9qbteWbAzlCk6p/rgupyUx0mpHlJSBGojBbLvZlZKaY
Fd3NlwH5wRiaJVKLV+PZLr//6BRn6jqJAWP31e3QlTbDoQXItq8UUfXje6pG7ISRRhJX9kB340zB
UPSwzI8uIlDJbtL8cmJEjL+63D7EBOI3D1qMDzN8xpAi/KVxSVvjcy7Xek/uToj5ahIia4TBX7fe
8/DUWMRtca+wZsUu4CIfGx2rqkOgWq8ra90getgXAun5XNugSomfNDgnbTuh1dL6Ud5uom9kbq3+
t2AA7PcPjRPizFHZGXjuY6RFI3w6TCYplQMAFY+b9ZKryBVtbn1rs8n7SgzyYoKpO5q5j0Czvwvw
q5cNdJmhH/sZGzzUZoAnFF+TaDLTKg1etJUWSmgGrNPDTudw06NgZkzzUdbHmmltaSLJvKe1om88
x3nm/zr3zANHn4nXy+0lzVQJccMtaFMvKFksyWWxDATx6kgfP0nspwbksDSJM9VHR4j2evyyFg9p
d0yFi/1M54VaI+YHRKod4f7yWBHUmchxEpQIju1ulLAJFxbJscG9LFoV8Zm120CPQ3lxCn/QmZPk
WKerYYBGWKQYUz0IrRhHlSTHhVrvof+L3odRWWwFKH7dxZEWjkB7lEgjZrHn3Fr2r7yxfQpHjmy2
luX1yrKpQJhTXTcDYHdpdMM99plYmTPzxQO2BzomjbtWdh6L3sOd888ir09cfelF2KsAM+4TIOno
veGkuY6CuN5w+sth1dVywy+Zp7pfzTtetIN7GPoLvsCaCoQTJwZLqXJ/tJNNyMvkroYR7t4n0Env
Bvkpnh9X71WDhk72gPnqLOVMvaL0zuSeMlKd4ScCDTfqSr3O860pEeLqlqANIFX7ZtkLcSNeJaMg
PzYrXvEhs+kN3HUl+uodLvZc/YH2M/ONV/XzPY6T2XFTCl1YceUCU0gMLqOIxZjttJrL/EteaB/L
fy2pekly8V26NZ3syAvU2VPhm7hwaIFmnc7c1juVSkSkhAIl7WKH40+caMxs0l7MWRIDQV1Cvenr
HgBoEu71gGQEOzaUgMHbrhvGM+XRGRdKiLGU+m3wnG2qBi2Pf2y3TJEw42ays+qPZ+R4o9kAl3vt
hhcEIapOh2aJ13z4W4Nc7rmrjcE5n85SfeoqCPnkuPH+SWKHL8u9Thbe8yM7j7E4R7pNP0pR8jl9
yS5eo3zihdbhzmkNj6ringPbwuutdv4bZiXH2u1xfF3rOptnAc+kWsuhTlOHk5PBiBJc8RE7wGoG
oJiHBXEMuX8zcSEDYlhKoKt1vo/22YxdQS0udst9Q1MAIU4G/WOCGn24zwZ6HWSNfnrcOfaB1ud4
Tefv6TugH5YPGZcIU1btFOzUygs8G31NWaHdsHedlB3sFyJxuR39tAFS7JaKL3ffF1qMCay4quPQ
DRk5HbW2RHW3LCWwUYbd9gQlrMS+nXZb+uiRHZDA0fUh97Ur3esxRHG97ZRlx22hwaRT+Fb/fzp5
X/KlRcyxFJBGalq7+MI30bWoyQOSOgt4AAG6ogMqtdusCT8dlQRs5swSNMOMTLsAD8MSP7YlH9rR
nJ+2bVBKtgqdVIlJaDAhkRN+alYGEzYrn9yntGqLIVi07j3D0Ax5CsPHzDa3yQBWJSAuzBwKvcuq
Fz52EQbVPyqroO9ywdx6/pJZc63v6t3AladNLJcMB4N7mdc4dH7oZVb1uxqJb0nLEbxmoz0MDsmN
M0PbYP+CKvdJmHrcaljDYdtW0adHJ6Yoty8Tax+5aTErI1srh/pxQOdqE+gxWBGdcH/of6a//s5O
TCezpDP6+6hFZ++rMiCO3MZDe7iKLKdUKHFf6YxbcWWctPGwcAjrUqe7VAXRImfhcVRwdnGYHKmc
5DiHkl1l/6NVQfHt3IrBqQWgjZm+8J0qpHtrFECtnXkzoCyC6IjZdoVXqsCccFgCH2Lk6uvaUjwH
FX6DtmvtRM9QhUL7xps3KJSijWD6ORxzjJcP6DNivugEKUnW2HL+UkR8IEdHpLLChQAbzowxr5Gy
rqG2C0qpruRUXva9BQYZ0WA+4L94fFq2Y5CcWZg9Iv7qY0jl/IMEQfhP+kUaxbf/M0x5I2s2hFtW
w1a5GcKohWhZDPb81ZZKULFvD+juJN6s6Ut4Pk8dDAtvyt9eaJIcHo7uBNFgKLW/pvyI/d7/E+BR
XW1hNrWlPnUZcOkQi2CBVrmaF6e1brPpaxbUysXasAUhR9ehL+HuEKSdfV0HuyafqZ/aYokDD9EL
nDYAXDSviTQiXDJsfOB/R6Vv1Oz5msGrdeRQaDmJz8KaMKLmmAxl89UpozUgHRoFDEPD7fpNS8Fy
DsJzkv6ccDg77RQoISMW3tFUolCV6yEU1Wo0PDvwiDHRD3Jz9HzR4+iN/SLM58xt1iE8cofRqZSZ
dH6/XShc51lRvYdLtKX4qp1W6lnwsDY10FWoJgt1PLJ8poZ1vjBBQxofnEBXQqreyhwMrvLd53AP
tMz7tmrBbyzaq/tdSlP++HAy84SIMbrxXLqvPTn+DwKFigyXOAb7bAVGaYsVNMMuobTEJDi2YIH5
0GlTtnaF1v6hNBBhJppDtsqO9G0h0NWkV42/SCTXZVXhlMTsZ9AYGPj+UzQLc6PrLAuS5rweWsoj
DTG2YmFxFC+K5Nsmkazx0nVJEiDgswJgeGiQ+isXg3jJdoQdJdYRUwEANlcq5vS0VAwOqgB3eTq2
5vAFozjDwnxFwgt1B+kL5QR6GT+iWRHSEBRwqo7f9pflk5y4KBxJiPAP16G7Q5JUm3CNL/iOtyY/
GNFmMhexc8leAgZzkeQrFC2x1HeKyEM4bbhoGw7UBpHmLWESMdyCrLXRP8pnESluYsE0dt4IhiA1
fBX7uCxyq0UumkymWUtSx5sbzUrt/AA0ErECCKg8IW73VX5YODKM6I9tyb34wEypOPdmFdu2Hfgh
8Wk43amHCwA8aU7wuzLbcg4hog5cnew8QXlJVB7GM0RTnyekMXn+spAPkn1x7CJA3emx7ubw2xlq
YV1EXXWAsVgRidMVsNFeLhp0OdshnZGdC6xzag4fHteAnQXsZbQdEBXN8xmK0VyW9XeaiunpRQUC
jXC2l2TzptBVSP0vprLmKZuMNtk50SZ8Z/pvKSit9o4e4M7+szt+SzHbepdSrYNBcswl/MlaglbB
IYwpkhh2vyi3zV8YNZ0I1EveUStfMiP79yebbdU0vxzikqn+kjDbifsbfXiOvfttj0x1r3WrT72h
uQ8HAQagwO7jUiBiDAI0lyXVXIkT4+etlpWbGwE82tZ7M/yAQI6hIfkKlHVjlr++0ZpSOOAiF4gg
khtwWKEjkTRAnYhSzh175hi+aDPC8PfrnU4rRS3ZBAxUwFyx4qwZHHVBiRoyHRfSfAIDdk+nt/C7
uuZuePCw+srZ0nxeU1b9ojH95CTe6xMDW8P8HjVGs31atE0vru676TxFAE+3cNkGJ0HPpi7K1Ddg
QwyAyHg6ZUsjglChpRM/yQbed+m3/mN2hwD2Io7a+GoOHB9z9F+DN+oTuX5HRDsTb6LMyYqRFKpM
RaXTFNN78b4gECPOuvzpGAyM2YAOaSnw8mVvG3ye/h2JXL7DdtkYqJEKvNqS/Yy+1liRkwN3rGD5
Y3YNCNXvTrFWK588OJ7hBBqC/Xd8HmWMcvTEyHsuPd9YngthVAMKhx8O88rcuXjfy95758BeUWGg
vShoZvu/RkLdBFhu6FgJvoCJHR3Q5VuqyqFMyELn9lmcC43gBHq9jiEfaiu9IN4sqtPnvB2vyX0R
VE23TGBx8ihuWM6cdKZ9obRDx1/1buJbFETInsw3BXjS3CFxvyA2837xix/pasSuQ/MKt+RV4YRg
5uwwy9BVWS/MKntgtnh0lMBCmecvIjP/nITafkd57+2xu/R3HDgp3pG2AjqtCxbXNWt/jcU6F9Xg
Q8h35lLurHpJ+vlLJERDmPPgAKXJkEn6sIbZUoNjmAETKgfcL28W5h2CIATzLUBFBzMYRSSfGDdE
fOCC9DZthKlvCe0Ey3WTjntk718cxoLLzcnb5n6ZxYyhUpjppfF9/tRUgqgzEdkyrhLuOVOy7oHH
dWz0FJcXsZpBnCwZk+GzJxEp/dKHsODbZvEiiDiMYOyW50lDSGMdRG/+G3t8tT6NhpH3vLRdMNHW
6Zfi6PZ//cg+7TYtbg5bCqGRU4UQ6gDxmATPoi0LZrnzcq/HwQ0OY/X0O8ahqpbD2p0mMxi7gQrv
+o6PKP9Uz7Mh5QlJwCkXGPcvvDWE6qnnIdJo61MbmpbOU8YtUQXpTw99/xFsRUVwZHybu2FcTRQH
h6E3XUJ8Eo7ra778/lQVE9mf4lJ3B3eUu98DvprWeaP0O7YGBAAfQ4G0O/QP2fYAG5b1I4HI+Pd2
m3Fm90X3OFDGPpW5UXvRj6Ho8xocIwv0wKBeBbcSGPJr2f9lQXWBx43gI+zka6YF9AO6PZxrkHZu
b2I4vJ6mb4eXzjgjDYlChP0fxv/U7Gg5DwAODUGU0DeJIV5Q56+yxNOq86w4e6geB7y0HBSiGtt6
E7OMA9pw7PzZ1cGy95fELmlQsx7ywXKom7P4MtTQmLfq/g44m2cQwRw8GFs+Fvw0SipEHWeiTfiI
ckZYpBkjrmWCUyWWlhANzNUu9ld4uE3R2tLoaERJVMdoi6GNnWJdyz/MBU6BqHCbUhK+tiq2dO6s
Hhvw41n9/7DyyTWmVJyBWTE/SweKvAUuWsL2+uqBIdibYVbUJDtCRXCXLgvTgPivoRUwKJ3dmeLc
vJZ0FWhvWqRrvypXRe1KzCQQcGK0qm5RcLaWjdUDjDVH8zjTocVbM37Dd8qdlg9sphEvQ/CRuqBm
6O5fKxcPp3Yc+VlGOW6vwLGCR7A3iLVrM0Pq2tCcoS1FGsWBBsVgb7Wh4XhAxD6w/tuU86yFigJ/
vnQ6M8WCdhdmV7luS3+7HyPSHGb3zrTEqu837kASh6d5MR8sxvykyFujfyyWqIWX7YXUa1N5KtDo
fSeT/TeISQU7LKpqiKuV9Wy/JgmZcxtwNJ/NqrmBgCoGYlEB3kGM77dU95CafWAEDsMjZud2Y9h/
AQp2h876BixPMLpf66CYtUisVSvsXszzNg06TyzAOSdKg8psokfn9YSpkxl5jo58lCL3jATlTuf9
5VHkYRdqQ9dcdi50DfxcADlX7uKsjnqhjrjlRtTeGITRyCn63ycIbVbWiTxP/O2FPNAp4lR8yXcB
bhKig/GHSQnTVXSsxIo8RPG30nHH1G9K5UoGPgMUFXbAWfEu7GFMJw2a5r0ZMut9oElfDdJ3//av
jQbA3xjU3/yNkH0/63v5z+M4vVHaAGbujHyVboRlBG5NRoB1q35Gospw3NbS41voo9c8gnFtPUbN
5hvBOz7quW4xWvYVHwQq1bsohQ68vUgHmywgjKwjFLJ4lgWsddwlaKPIg1LA9iibrDBSRMVqQ2MZ
EGaye6+OYI2/RVFdD8WOpjjuhy3WPGOLhwsh7CcJiqgjcEFT2cAg3JgGlvE0Kpbj9NMwHQUHgu9L
SPSKEXVOTMtIi4oudR6ah1I0Ue6Y6YWr8JTlWGFyi19CdWdFIh7oDrLJZiNAaygQriiVA/uR6kPo
v1zl4gxb0DZIcQ/hxelQr5EwXYtNTyF/KdjIm8LtB+fjRjlubVNMq6eSj+oZx1hLsqdpsGcaBmGj
gYR2lfUg5bClYtFhc99s/H1eTsPj9v9G44rvltUoiIqPlU0qqKQPT+goyOh41T0B5IoTETRdN9Dy
E82AFoTUbTOjrQHtR2R8nxupRDRIMYcqTUGQzLmDrEuaeZykffFsZHJMZREc2FnXGtirQq1Ojf3b
nIlYeAJkCe5eUEgf0Povk/RCzMsByULQMlSW8JGrdHPPWR6YdZu0lujCfi2UBIOZ0HH9Dthxb0B6
Golh8gqf5Ppgvbz2eEc3djvJpY5fTSfoDx4N5m2F+WuX7YesbDZOjMgsmCagmwbEHE/L164VMETY
LVMO+GXNgP2U+tbtwj0k+6dYu2qhTb17Fayq8ey4WmKVgHFMNdVTd+Z7hXiXEX+qLDledHe6fY+5
Jz4WRGtxhrLzvQS4DCwCgYTEGb4kllNk6v65+RdC2wH3WbBtM/la9DqpvBdFU5Vm/ltiDl3lOfTi
rtesHdF/TdnOPoPFpMQokIYZFw+ktfCGg7lG06LIi8iyCS5nkL1tOrrSiYu7a5PVAscOxYbCkSYK
T13C46rqigvxstPbzvLuu4bCxZO5HTXKmIhsINnjYqwxs3/uzuFW1Dy1Hb8mGHmOrW9C8QdvQ2cs
fcrJ3Uih23qgEpNl5y+3JE39TXrMT3HkSepoTWlWtL3SBD0uat293krNLlREP/AMGenBNVRwF+fZ
WSYZVGi8udbp65V56RMt7i9gTnWH+a76/uGODgMTrKYxG/6rFsohr2lS8kHJvZjLTLyY8dtN1n8v
l4HHh3qEYkhCdtGC5XwwsCn6rhJ2WKg/6RbUcPdKRnfTqVjQeTPKC61rB75tH32ZfOO7YyzzqrVN
qmudSvDZBuzOBn8X75lAPMHbcH5O6Exw8HI4rUjAgXAMxaAHI1VvgLMniaPnNgcgNqX1/VtuTlqv
XAZasSKKfc2GGyJ95zvrJa92vUlTgKwkIH7EDrq/er/Txkdi/p52jmZsfAtrh7fMFUT6/fQCH8oj
6S9nlhesJVeRc96dWYwYxel9ID9v+IUvwb33aPgHpfPs2WE0rfUkrtUYiqFs5v/EQYjtvyM5CY0K
RnC0JqJ8Pmpve+7teKH9yXQFj5RFDX4S66roo2KlIKnoKKqRBawF32Nx48PV2BqlrUACtuDgRCcl
9F6+UpooDV4hn24vnIT+5GVkWruzkCj8HYYNUbiYGMFm46MKu37THlXQkkHpFzFfTY5k5uMnoWZ9
m025bcbLlPmmpeh9VhP+AZrNXm+qfdACFsbjeKLq+R5lAyqHjFRR+HEKUppPrBeriN4S/UODk5zQ
rS/UDPg+7tJnZ53cwkjKF9IAXMV3UtUgk8X1I6W5Gv3qTu5mUQ8lbTNUNx1g0m8k71AjW8JH8Ugt
5GRcUEIlS8oGS7RYgxn6noGyxlZEtaX8EcJ7AN6ryAo7gOw8AUOdk2A9HHM7p8LYUK4gErRjEtnO
NQEV+xoD9JZo03P3FUVdUYjQDaJryRf9GEogcJOS6WBEkodLVU3yeMmQhNbVHeETWJNqo/TFCycN
cCrdAts/vUFJA779szW3CnFyBwWhhsYBpcWL7zYinptMzzRgGlR/vlx6A2/stwmcWk3lNlheKdJl
1RWGlvXwkhBBmq/CkHBL3HmOOdvEWDDmltQQjeMRFlzTs3jaVwP2SEcWFTZe7H+q2Ks5Y5A9Nbg/
VWRBXIMwieuNX822hvITPcPtSSMrJc2LMkNts8H8TrHDOknBvTx4sNERbpc2bADq1jadkSnR9biD
RR8rofKkdcUOueBRa2Du5djUYxJSV1xQC2ZVY1cWt+I9xObQsw/hxvvMaU18k2vmZxIb8Mqf+564
p/vb4xyAIzyBhZKw4W4Qf9J2Do2RX8StGLGr/Xarm61UauNENe9EPFO0HhunhdZiNkzYkdgWfIO2
52NOXtbSFuwLJtZHhZR1js6y2qm4oHfh2ld4LrU1UAOkN/eBb4PhdrB0z+W5zQRmO0SOBcmRKahy
ZmkfUDrJui1KoHQTm7WVVcb8LT6MTWoCbbGIqtn6asu3JUneeAm3OOEyT9pO11p6jm7+TX6TjDH5
rWt5+k0z2nCeLtB+nXmZxtVMyUWOSiPew4jTg8c49FU7+7oxRDnFkUh3D39eT9HZxJciL8lEAaF6
Tpu/mAnWJpJZLMI+hnuYT8SExOpSMN7/RI7XXo+yKQcilAFiY8y6JkUHSs3rWR6NkGgJ/Avrh3G1
XbLHlI6dMQamA++q/JORWr93nuQ4IAL42PchVKk2I+MJdrGUuceiBKSQuHb1xX8HI8z1HAO59rbz
kOHx6nUh3+wVcOUUx/GDqvH6IAks9mfUTVvA+fN/lwuVv7IdyW5SQlKpEuuqJ6BkmvHoR1KunzQ/
AiuSaJMLNknUkYYXzXTISPnjKHOrF4vfIrv/U1ys1sRob8wv5nTLOHPHekXhtxvPKaX/gShkKLY5
Hjbm7NUzx59bd/5PQ77/Y9elsJAqFk7OVkfJJR99E29l0vtbNwxPxOdGKI8axA5sd9OEdCp4hMN9
o6onchkdPy/J6uuXc93udJgcwFpPWTf+FJw3rMGEuCzFl+9XlZRISeoSeSYJHCUow7VXus70z+v8
i9aYdzwbVS1NdTDKg1f4kJ+xmQOMQjQj95RSx2osUX6XaLRBbhWyx4WcbRrDkkaQIa2NnO7lBagX
tzlg8sncMkcpTen2vq45CFfKwqZlyqOXiYt76gK0BnLbR4Pt+UuViRYKtaLcPphHsNkH7WyjaWP1
F++jMC4DpThe6amBv60y4tQc617K9RdLQi3vUFNfCkUuFa/B4YIcLSG99PwRO84GkjIuBtYYyBQ5
xXaoI+MDhKWT5cKktRSl2ufw1yYcqdb4iXvKvP5LNf39MWRx+PhBUQ3rMCPLbipItldvKIHYDQv7
nLak0Nz2fQMRdTqwnIhtkdNkDc4RG8K2LDHRLJp5v3yTxvBv0586mnry+2CNmSLEE0ma0S3Sh7eE
37I4VMqCbX3P+X3d2FFarx202e0NyuKIBcog5z5aXeATaEDeJnY8O6i6/l+BJ5wY3JqVCPNfCm7T
VznZ+xSjyyR0/a7vDs2fP5PRL41JBIpjXC40q4ChV4wGCLpNxU9DNr//HpLAfGJ6DSKcLCEI8PV3
V62XBD1a84UwPQA5eC6x3DzGfDS6v7A4BmGHmWLSsqpMa7QtRclpzzdHVRJpabu7UeldZAlBvQbx
hlGaqvR4GNRO07WxLwj8+ZGQkSjRSuQR4j1Ar0EkYx3SNKwUmKBoYVp0bB/5tNzVPzptN7TD4VFG
byxmP1HPaAVt8Hw/vC8v/4424H+NmvUCn7dpfrY+9+02fgP0N0wW2D9XpvtVYQtL67Yfk1f8j9KQ
RXJYT1s38h3ivVxWeh3y/Se0oY1Lv+2NjVqfVCcpYGiS05juH495OVFMqXcfogm/jAQ4BFGP63b1
y1lW39QbMs2fS1/XfOXF07JegEXuqrOCUHyiJoIXCJvEFdibzRxv3gjlAInSXH4+8ECWRWkEZzSQ
w+WEs1sVurYA7f78rtstXSXFOwjULHpirK3q9P66fvFAqump5ffWJyuXEBMSYFzo1xqytO5jEx2c
4eEKK1L7snJ52ZjRI+ehCEGbs5zi9Yp1be2ucdf1TQBajd0kMPUpCB/Eh791QkMv3MLHG2wdfkLt
fktu7pQlaAYCup0AGWWyxUxUlT98ZXQwx2+9kQ5ffkjDB9fhj8yXyS7La1ysSbTQxTcKGt7QouN2
NCe/alp5tcNfenOANtiynpRLaNCLMR7KLgmQdpPGwLqy1ISGG9qLzkyZ3ojtnVefkebkyCu7lmXX
A2mmVYGhl7WBgnB1fs6yD4QWOENsfbkd3Gkbqqtk4QyGJ7CuWV7DwLeVvVY97JrG7Kynsrqpf1kD
uYZ4XpzoheyBW9XB3zq6tOE6temWeWrAoLEDf81y4c92i6AGB6TSFcTQf8s/j4ZRK25g72YJOoeF
SU18vezzd4UTaVIHjz+XpPS4hmFeO9uXXXfHZNhwPW6C1eLu7TetaCvVYdongnC7MX9weuZBvoWQ
QrTTIsXQ0XWQIQi7BBo2UQi524U5NVS97bQDgig3VMYhS0nSj1J/3mGfRo0Itld1d9dch9PwIzo9
dElgA59VGFlIb4JOAvFG6TNipFA/UTtvemOEBggjryLb1L76OvJ3apl/helPWo7aF3epXajXl8+2
II47ut2dMOL3cbWvTXPYyArUN3ZojeyWlD+UVwiSNI2c6tAnq+hhpwTZ5CHP3SqvqDhAgiPq4VFd
c3FAqCEPBYpoKJ0DXSnTzhex88nShvcUybjo99iMPRQb06GpS01Hp7gj4xJAd4VSgxj/h9Y1+f7c
2xUmjHs5y1RV/x1//hVvkJCtMYoT8dTzP/yV4KvnM4uIDtL5rfcDPkQu6oMmlJQAHRLQvKzN/cYX
kMuRo2kQfzYWLiffIqJJE/vQE9M4vLIhN3HIz1B/uLnQfrAQbbJj6Lvh5v6uTndh/SE7LKabjGTx
+M8E7DKmJ5pFAWgIL1s42KsBE8YuYx6snTl1hwinOcHGNwC7ODJDW/xMw93pXUgvH+0VJeXjxDlx
Ut31IUHxx4dqQ+fbkCLZHrMChgyOyfUzhAQIfRssYeRF8viq4fLV8x7jcaV8OvnXEqOBUlnO5trn
3Y8cxsg6FXufcEfLFj+X+AShzZTi0+tKeZX5hPut7Ee8HuA5UEyWmVUjFFV97mrvMROOalZgVUXZ
wp4a+utXjq8xrxoW5xtKH1VFCju86HvY78lcZUolx1Wkt/MoPyX89lhSbK7O4BbBuJSIpU2ghlR3
6YbP1gT8b+gaAt5cKGeTW71oKORUQeUtlyEH08IuK+1xIJ3fWyMh29l6WUz0nbt+j3iiXv3iMYJa
qQsgeshFejQ1vc4PfvbRjNaF0QpMJ+oecAa4F7q/qK7L2qPXvLtD2PnIQcGmqvrP5zTguaROhwkr
fDwhTnT8hV+nfY1NYuCCk1RFtg4FtOh7Oq1SdwsVYxzm9DzyYEOlQciV8TfraMJC4jCl1rk9VP8y
4Io9swHbLyW3+v4xREkLJwsGXnHTBoArU5b3/zfiCX4Zg49uuOLPbURALoZxfyk2xzLENc8J7jmM
B/Jz+bU2G3kDa6UF9FCi4jweUPHFWRj3UU/TALTZbHfh95mBf5Fptv3y1/IN93oe/NJu2rCIrcUq
Cq0TveVLyHpgk5jaqmvWuadLL6caV6PVbiX58NHby8pLvOnpx7B+4ACOIV0C/xCKYlo36dznNHGY
MRbBJQ+wKumjaquCQ0K9Y79pkBOUhqa9eYM/x4lzDHGkWMw/VxMIhowcOQG6Q200rBdfDiXXqCMk
U/LXMGczayHH5u7/vGdVvo59oGaGI30U/2FKkerMbGFxTzKDWRNwslBNkYFOB8RpAkikHn5hv6Mi
ZovLfsq7MNV7gZwn1SyAmru4uBUo09irDzjfRENgVee4ynvUE1tZ2RhyWEXk39U59uF3KTmMiMnd
9C+ZQApOo766JNomfhsi3Us4hAQ1jZrCDUpB3p+Kp3NfqdYKpLOaUIno5bsKt6DsR71x6w81HDWh
VcPFLU4HP5SGUnnVjGQXpcqbwuD1/x9ae2GI4NpWnFKQFeT+s/0k5PEQ8ewfIqcK5BTqN0qaiN+5
IbFoxIKhATjYbnPqz50daxZ0rF6r0TPm646L/UIDedqKYslA9f9yPi11lRuHpj4/8n4mOPe//XqB
3n3qAYIMoQRzoa5vwbCjNymoGjXX6C39800BTcmcc9iQr1AiU+x9Ot1f2RJUyiENbaMnA+c4VkkY
jo1hhTOtsolns5BFlJM83Cc8scNSGmBu/Q5A5w+25yjnPTjyxUVqTsfj0WwCT4BIlGXjnS8iCp1v
KB78PFH0pbylOd1KZC113zJb8uE3rAUYIOSK7GLYNK4nwuo+LA7c3gTI4v/jbumDzTyh0G2PO8PL
62bYK1K5pz8NHSlivc/SNMdJZCOq0X4/nKWYPwVBLhhgpoAFYOn1zgXn8F5vjDUy9JIdN7l68Mt7
jwT2EOrA3pZ9uX8F9bG0t3u9o3TWUE/bm8N+l4/IReHv2gC02WFTF79PtFi5KFt6c+sr07FrlNAO
JCC/GZ6BeMnI7i3CGuExyWW+p6vgOSvmd9ztotsAtF97x3Ts5rggxHklLlxeML5/Yh2iBaDAx8d0
k9jg5KZjlUIpVFHT2caknA0hvTZ/VqRIyfIIUgxES7VdnC2g24o0T603leIUNUk7hQVWXzqWTJOU
G2L2tuuDcuuQvPLuX6zYrYD95sP7d3u7T9c6z3/JPl526geA0IFmbLrtG2Pe5xTOVy8sLrpZrv1O
Q9pW2NF52B7CrH9n1eHBTIxm+QQxNym8YPLhCRKru1vI4PJISTAn4Ph7gW8qfz9+yN/VPHlJi+Yk
zmETGA7MBKj4NKEmFQgZzxL7g91xZAFW54pbFsJdUE+j/hVzaF5J+bFolnVbhABhvsPDyIbJ0ICS
1gWmt8wCs5a51fzmZN4yFi+BCy+jtfEMWM88wf9XA7uKfFo6TwlZSri94Z1szd+Z0GogZPgJf6pM
06LT5o14VotkZ8gOiWtNzTS1jOa9pOcVFKbZpGQ0JOGPguUM0ZJ60bPlHVkxCf/jvF2ZjPJHDokz
+5HD9Z1XiuF0nx3IYxonQam9DiJGtvu88i2Dpw0JT1uQVq5qBDoB+mfPKispCaLVblbDMFyPOyUo
fVYVd2wDv+KGeWhd5GdQr4BzsWBos6ZN7bOR2BmB1nCvQPEPA0rqlk9geCB0GHjA7GY80F2dT9aa
dqf5osV9I3HhFDdtFwA0QKcanmyjVejOpRONMhWF2Ekldvvzx5V419/saZg9nTXfvqzb/69zk/hU
5HGd1DmE50o5FrJXYlCMaexvBGT8WjJ7PQXp8Qi/U8zy0NdajQZNUs30E+yDo3f46/Hh7n56hq/I
pulzn7uIKyEowaN9PlB17Gy7WCCJG2EkuynuZtMQtd3xnQ3BcXJrASXUg2onl0C6Hxo0XVM0ooO2
DQ9imWNWnPlbjVcbGdMe8o27g7oHi3+hlx7Wwt+4dHCB5/rTnbH7jjm+wGaBLglgNwysiBIqgWyk
4g6ZSQvj8JzA6nJ8HFfY8KADKev2A8gztm6iYS9vnSuP8HaxT3c8RLp6BZB2dP7p8H86PPVO9/VT
RoDpFY5+F1cXh+8ytEw4QIJWytAczQAO9pPSGQjMsSjRF7GHfjT/LDbuZ7M5XTAERuJ45IPE+XNm
TWX24pfu9W3YxNdpMRIFDdvmayOpHwT4o10Uw36eMOzFhn3XeB5YJkPBfi3dVjlT6cw6hirO16rP
VSOAa+l0SXT+sgeJhrB3pch5lREhOPerdOSNXI48QM0OknObGdwf2ttDugQcNOYFutjGYRlRBXr9
F0bq1nbmXLDKVzmZGRDJMEOLyBDdq8C/9VnWApIHS9EFy3tSXQlaaf7abupYbbkcoPKZvW0UBIo9
3uFiBGrNhzY6u5nydmbaF2//uUks3R2KPNLb5BXSnGy0lafS/xX/rRWteTZ+g38T7h9kZOohFyLp
DxMho4ZOIF/0+OHNPwEhG4yrycokZG/qWuhmyH6Qn3dDnQNTA0cmi8DHSBWeCARGdttNO6lGKVNi
Qog/MgAAQYx5xNz7IyosLdQTpO1ohSALQxg4xGDcPWj94R5X7GVB91ng1D/1cvyRWI036k9Y33St
FHIa7u1ptBDG33wBKHsCFTScO+EQb+OBcpjpZkf4gT5PT56WD3pk1Z4BCGdeYrF75xLzXXcAWtck
nXFB1LtHBMsTdfqfkhipUfvHo2l5WcUwXJO5JtukDgjLejt4CXl5ckAnLw477efKmbAWwI6zy1rz
DbZ8is3s1eKjSq1MTxU5PgvEezOOsZLyPgqiQgpwcEXAFeWc3+Ev20ej0dBTMIvfwokL+nK4Ypee
cQClOJqKPe2UMqTQb7XYLp/WyjA9JC9R6hpnPOyOQdnX0vb/lcJ1pDQlrcvYOhAAijcZxQBls1J5
CBwiL1Gt3gDtjsGVvPEn67jecgKQV7SqngJBkm98HWP+ePGeDFDl69X8O25AsH73TRSkqyaXh+Aq
UXy+7sReu2LNrIYskLbUlsK8Gld3O2bLokXKQAL0wFughaKOrX7TQmKKcIvQadE83taBS3cSHkDd
hnuX/gCBdiczaAiamGxSRJ9smqYf+nClk1LtUjjOBrLl+oxGliiV5cf3MJTpPBpvB9qswX5yHV9r
+EV6oiGUWXuUFczF7OudU//dGhSENe3f9dKKohTHhxabyr+aYXN75t4gIteW2xZ+Y0OQSBzmL91P
7PTg4rLhha7nVxiZ+1urwezhq0qO0aLsvYUuUvL6e6FYbA28krcMKieqD9nQcJq6ehtG4dQSim0E
Xe16KOHGpJbKrw7h+RpSR+MlOejF4g4wAl9/jOC7qx2ejiSYilAhOw1qF+toaQxb4TmwIv6p6cXf
G6U4SD2aAlPuaZE7Lq5dmS6z+2gRRpkEjOhzUxjgb5ctluAA4/nesW6RDW1gDSVqdyPDL6vqKdrW
dQtEQmPK7v3vGtjZo5+CaJrgMeD4klw4S2ISPIhoD5Y6CwKHCQAGHtV0LZ56Ec4SYNmyALuhjhxA
UwVBJo8O0TeioYNuxIivS2Hfrh4N3q8bTe5hME18gambX4h+1FMEhNXKCqytMdIbbz4CZMaNzcXd
UfIPn/vTLOmKvYnIyMfvGDj3SgWnmtd3h3s1vzJkpfVJ4qKy0I678z7TWwu6kg2AwswVQLuH5zU7
09FFUyhuGCTBkB+GLladdHnHdQqgxnXrhJTY4w+4icgmFkSB0Fb+KTFqvdM89m/aO5+bMimE8G8d
vuL5qiWTgjDPt08eyM244w5ZOE17iwkvrjTahB+Sy2CrfWQA9Uh8JmNJmeuIRjkMctepfjMyZOQS
NNeQ4+14csRNOK7VRgwqhZXDz0s4cVIPPN/UQl/9aXRXZMgjYod/TOPnAi/WAKgThmbah/gr0Z/4
I4S8eQAytZ694HzMshAMaDYkP3aYG0jsdP1et8H/oMKC81GXQ+FT14YssYjPbfIINhqG7+lyQ7GG
J78rRIcRH6t8kfbO3ye7reVQR8c67h4PaWSfy5/jvWydPirOtNq0u4cu+3ouYzaj4JPvkVCY1Bvj
CxLzAkIdG9kV+ElijtglqnIUPUqnaDorU1ajLl7csZ1f5O30VI6BA9ZEDl++obOkS50tcAXi7Xoh
OpHLsa7vvZa3c2jzM4BKvtIpzlc40kRgkGjnF60NZQ9WYnZkUslG399GsS1wKLM4p119eVApUNRf
XnPtLvbKqIrsYFFufqSU9Fcv3Sgq9LIr1tADZI52Dos7YMmCHRsPB35Bm7UkALKvrOt/aONhi3Lk
wF+wpgQ8q7u5h3toVbn55ohsiW/ilPU2ZSHTelXXV7722mHRO1liAXOoGE1RO7qKp6zb+q45dM0m
HipCSg6vtZ8zN87wHsm/P9LxTdkrqNL8682khgv8g+bIO2Lvm0zrJd4HAWyyudovoZoetJVYMccA
VoxwPQa82TnD5Oy6LPgpcyd9VXeA0NwH06277BnW8hHqwifNXV1A0wM5jM272SqRVBiqMEQo9KfF
mhwG3XrkskKhG+xoCBjzOaRYcVJfpPRyEkWDi51dIwrBp2yR5RxKkH0jzz+2cH4GzevqiyNeBXJc
bm8JN/VzbfiNSDPEQjwHMRiFRrjpUE7XQHqkHQSPdfQ0WlxPWS/veF3s3eGgAhY9uRZjTBiiLWll
ae38aMyuHMCaZTaZtmF0Ybks6oKTcDHQi0WDm5F+ySmJ3VBbZrjfxZBfwy1DWwByIyoUaP4oU0yP
yqY+7Fw+ovg7NmjUiYY70gU01lEQ02TJ3NeT9B3pd3DqKSF45bWKfRTRmPmkdYWMivV8aqCRnXAx
N/LLie/RJod2kZRvvOz2GuzU6O7aYiqFG/LzSjVR0+sRVO0o92hqh9+rSpy2MgNlTGoeVQW+ofie
7JvWinObs1e6mn2SREN1qqM0Dsv8xM3b6SD8TYckX3plZ1FxsTH7FjERVNDiJ/94jktP89FrGDOL
nmWRg3H+RHb5zo1Mt4QFKf8A0jpniJA8w7tKyO1L63dS/YZLeFIbziKdLSRbsGpKmCOWW00FKc5U
UKVxGZq9hmzJ1Om3I7/26wpXB1riEhK1u4p2EF1QektZHIKaYvDIxynnYs8FhDHYp1zvNYgsd/9S
Js05BfFsl6sq/9cippmyUhdTKr3BX0HINFz5uhxhIfG9W6I1q/6mXIeu0DRGnJo/2xMOphrrCc0B
oI/OonVT1oVh63Eee8/+di3doOwUjf1o3ssuSBcCMwYjvufGKbuOo0silj0BzoK5KdOLp+1zMnKk
SjswXMKjVoVUUQ1SSVS2zFnoudU71iPN+zbLyMSIeT0Fxgu0HkxNi3nkcOBGsBMqHNW6O9tNVN4l
mbogLNLsqWfP7YnBbvJdXPLFaixSxOgW1vCNBCLMicbhQGHvcWaS0tmCA4BCmmsuYcNJlTi739lL
y6uvmOQF/DF9U4CbRFGV7xlft5uBquUoo6s3DE8iuoPwOzRQquxJ2QAUfgwZ9+BwfGQ34IRMZ1i/
kBnYz5z7mZgigSnEUOdYdB6P2KjLJtKTG5yRo08fzvzLRpWjxtTKbF3erBs/vGbhiLSUMrETTSgu
Xvx00vHwsc6PuyMnrSugpFvE8gb4JLZheArVBN/fzWubo3jOhew7r28NLqBCWrR4xnROTbwItmFe
/wbEcn/eHRIZtUjhDiMwtUVNERanjOajagUewtVFNMHQnmtdYfjqcj3Y2+6wLyR8zRNEUA0WHxZp
Dumij+ZcCXjwYftV63seXRUkFmtepsPRZwgfa/0zx0003sV3X8d1pAOQIb/0RVEKW0joYxQUhL9y
x1hkkpJ6LevbiRa6sK3b3VP5RBrRzTpGPbbMjr9p8YdMaD6srXNxqIg8H++kKtabZnZEQHksj+u2
/LbvNM+fvPRShpcbfonx/Z5ufO3pi/ZwHrLF+o7Uj05fWZkJuJbK2fpIMiTecbcfknrgBAjqSsqI
xopJE0yn2axV1K76oDe5II/AKyhYz9dqjBDfyloI2XbiFy2rOa6tJs6htpNY/9N46XJcZZR+DQv5
SbQjv2YGDvxu4p7cJUycCOxzmXYi1bS6kBFE7NFBV7sG3if3uch8JE1H0dORKsKR5xqdLQQpdrgA
8sfBLQNUx5A7edmDF/X1BwBzsluUIvr3aiW1xvMGY9KDX0pDNkfWX8QsIpqreQi9XpyMSYn6fUmO
kwcx5PJdFm1ul2mC60oJGseim0ervqFtUSESdVsIqsv7PLkwd0aHFfq4praOS5a6HN4W13q2AjTn
d9iljdwimnGdflyLz1eCJQgI66yeZprDJfgDD+n8edTTC33RHlZ4JedUqLdWj3/Dd/9VvIprPmPd
sNi3JrSonTVqr20gg4LVu55gf7Ys90rmtAgEgQ/mf6nxE3IwaBav1F+9YMM0xVfi57OcfvVU3jF5
iMniQ+EeIqOPM8sAukgtAbwZ8jEWAdcioh/01VneIiRucYCV39dSQSt2FYqEkoZv6DBb6bHT2L9t
H/CB2HSfFKHl/Vj/ABHPMaU9STR7Ssp+H/Zm5bD7d3mOJmFBzdCA7E1Y94Om7gEe3n/MxDMGPFmC
GH1oknA+yUxt/wT9g8RLTInS/OoN4ur8lzVwld+JMuzjs7/QNO43eEUr5/m855ERDzIY4CfN55du
HI1A940h9tgWtPaitK1OhxJqG/f/A0UCa1/fHm2SoYrlZ3lDKv74q6KZ2RaGh1xh2w8fDL2fC4MU
ZMnB5aUg00POyZQdhkCaQigssnrRx5UccdbmrL1uDK+ghRqvbwqojFO14JH7HCy/FnRQaAIxq1Z1
z7v3DoB8Xl2ErNXSz0zb7l/Y80PI7/kfrIYRsHd/SmL1OL4fkuMlekb/xxQixtKcnvjrpA1ZfLaq
KYE+3WWDscrNAEGIkyuJHSy2x1dkAoqJu+enQNtmkiLxZ3+c+o7QwLdFPg4B8yPBDrm7tRbiigAv
UvnWFu8Vk60FpKLvIZaGQsDOvryjWb+nPZnbMpq5UQ7T4Rnr/n3Tsv9ZFSFr9KaOGihslU6fIrek
jF4CAV6h372f8gyzDy5YHdmQnbxNkOkVAVi6zEPeDjFTXdQ+tyC+6dDu72+o5AVrgnjnlmWdCr0s
mLiQxMvcE6xWQFN9iWu1RiyYS0ryxnoC///SKCgJ5yckA2tjai+nESge6Ev5BxQUV7y4ASI4c4bV
MJ/7OuY0y3f0Z45GwYFLz8an9Af789RAbJqYDTmQE5QvHoBTn2SxfAA7LclMd4E7WWscl3auJuCP
NNkP3IK/CjGzicJ+MEDqQV5eX0Uz8L+WVJ1ma9BoB4YYSoQDtvpoZ/E5GRJF3MIcXLCJnL1K4kj7
WVue1ia73PiWnpEv43u0BTYPiJ5bCHF7tQs9knVYzAbQ69LDSdscQhlx9gMLB88rjWrQe9aqGnm8
4XjLULKwb117Vbi9HNAnbBO0vDbalOkgQnbbh6o2Fer80JCMdeRvLxw9aBe3u/3/FbvvHrR0/Cld
XRI1kpFLd1kbb9QiNH4GBGIxkxtslL2hj44a/hhWaGDsyLuyffz4EyIY+wKSBcgQAT0EqRnhIGs8
OoHJ/Q5XpK20ytpq3OqypSnj1e1sK9/CSNLX4/fy/+qs0sh6tEy6MjXMu3bxOdoaQsKQ8aHubA/f
jlXnOoIVDa3cE7OdRyAwQ+ADvsT1h9HjmLI6VkoF5sVQN3pUnhpiAOhSIRKJlaEQTZLgYETfjdUp
lX3BA/OPvL1WQ3MqFtaxxzPMPokhxQAuG51xg0fnRHNXYX4Z4++57NyVHKV2iqgObTs0aLNq0C+B
MfPxq6IC0dyTZ3KpXlyoUSoeaaq7sfutvoEZaz2tLRfWJm66QFsSLerZppbr7TXLYxw7FHnZVxmX
5D0TggYuimP/WYNo8AzXhd8ElM2EzC2/nKte0LEMGnkzZMmflwgfkL6oPZsnOaU7LC/kQLvXOis4
TZ/vIzfPfHbV9aHGHAlxtSnGHfFFvp55sk7QtvJ38Wk7ube4pZVv5CKy2dBcKJk1sY8HIbsK+Xm3
VQ93bgdgDPIgcokQUSAB/941MU79MBkb37Y1YoG+dn5uDEKQ4QkYcKXJk/qXe8gDJxqHBADzUoNe
pv9ukU0LszDo9MAd4ttStvY5Wt74uN6nn03xNlek8jlN9UW8iDQYYhc+nBtMMNBxc9MPVxpIC196
7nuVoc+YPY1I9Hr2IT94iwV1NRbkZYuLfxbddwBof3HpF65Do7xpm+CK5Ry78iZrzZbU4l4L5D7n
HCD0iILi84kN9n8uw3zPLHPNloIk5ZNyPdwOwEdVz/PNk1QXE5FtzI7N1dSDK/ROhA4LSA8UUHki
tLHUIf5bmKgGlNHMQVjtOGVDBNUtQZIQm/Jl7H5Vf0SJpqJGBmiDBf1UseV1CSsVpG8jC1RWDLN4
dz4UBRAzvbX/XxBPnlzgUzJO/emibTd6hGvISh5dZRdILeYPryEPagGLE04JGN0BYd9x5S96vw7N
ZDF0aUaexaWa21/l5gcwxkiunJFEl+f9llOIZH3Nswpqb3Dh3XrUqE8gX0mNyCFNg0fhSfL3ZvTn
2aG2g26vxioe4pmVJYK2WHDKE1TCKHh3hozohVvcCak/enkOJjul8FEdE+OWLdapgS3JrBVGCJ2i
cgspLm2Su6HYXx4zMaQG1Vsbx31oW7E1BV4AJa/CS5ds2jbWTSnKIl8Qx+qUPF5opJdZkb/QkiEO
62u10tbF5i+vVaXhRR+vIh4zeCnRxPAPNUAOOvP69LKyp+WMY9AZZywQLc3QI1NPuEhyn40vr3aO
8R9GYzN/EmYvCMab66jFFA/S5SsVhS1Izo69zd2jWYxNXIGvuHFDh4eg66D/0xwlbIrUKLYo9Rrv
Ql4MufJ41uRKYxUBpb1wjUiQvUOYHc53/gckiC13WSxO+yQisIz2kOWaqZbSkYeTYbADAihEIzYJ
qwhSm7DjEwYk8VLYgo8/g4fnNT3D/TtqDGTnRnn+IZI8ur9Ce/ulZZgzD1VDGsZE7zTzxCp6l6XR
RIgGxp+tsCXI6ldPeFawWL5tx8EQdENt+x9RxWN41FNus1ymbTyRmhTXzIH+kpqK3FjoIgbY5aBm
2H38F1/tuRLgVNxfB7KYlCQhjU2q9/+DEhc6ueCdQeOCA814++VJqN27isevVf9wxzw36GDkcFWk
nUnLuTHrLmRFP8FMWyj9v6w8YdoHLIGv301Tg2ka2gd1Mu1pj/J/InNLPc5ymTzftwBuOqzDoh9o
A2SjALz/ZBzGKJnJ6m+cIfB9GPXGsVdeECNdmLBd3nlB54s9L3CHUJbzS/NceoDkUDbZW7PaytsL
MGcjb4J8WJvZmRnjAkZt3aaCTmZ0TXoECfYa0qiv6SfPYxVQz89a/xHxq3I7CDBl//AZSR/w/FKj
d1aif2I8gN7aWmERLl9qrw+kITXrtzwV/l+W6ZfJCWOhQtVQOBCVz4j5GNrgvYge74fAhQwSc4+l
ikUc3H+o8zGo2vSCD+ZdL6ySFUluoQtrSkRN2vkvmusWWdAPyk/s9VS6Hr+U0Lljpu3KnQlTD/0a
0fG72oVQ7nbwnhuW6TKVLyEzwt9sJ+IhwhXjks5XvQkRsaFogj5DNbgHdLq1OtfGHLfzUPNIrFgQ
6EORSQJWcBd2pxjGLe0J6NTwOLPktLycJjmTZ+uzC1XgafHMLlNi8rd9TWzIvBZvvANmB/yge73y
ahUSb9ztrJUaG0eZifJpcEpopcCzdT/kKq7ypJyaH2cKjBOJdpcogdiWrgIQ5rfTyany+rGv3MwU
EVZfwNUZhdlgSgRH1i53ODCbH2GrEdYyEoOXgWsDIXvKfj5YUUYfS0zClR4N2eOLLEvj+mcVPvaL
abkWxa5sG1pj/aWXU/FAC5cZyq9yPcddTsLLh9QsqCnQK+Y3H21ugErDcZbXs/IKNe7NfSbIYLxn
nIFP49SprBq+dfyCbeLNzx92wYlCgzaeS7HhvbR0fIZKHUR24VsGq6hRn0+bXbPkCwWhwtElv/uG
xSRvAfA8YXdyeeA2oMM/P07R9YEhxNQqBZmfGSeJimcrvCHtJMkR4x9EuNtQiBIutvtE70Q4uTSn
kFVK9RI2dd6CQGIU5fS2KEWDfW0/PFaA1DDtB3oypxWiIqX/gjcCWX1NsEjyCol1ZFdHoqUSkwzK
F7xAjyO7xnKSZS/MzhKMsstMX6amuhWV8ah90h46UDC7pyXXBBQbBVwBi8rhsM9lpqimbNVy2yTQ
aI+ZrAJze/C73SMv9YUzOikIk8tBE7YpYGru2YdY+TLg00UraYQJafqXPhIQfA9AmIzFw428bv4W
MzvZ8xSJ7m0QYO3RqGZKIQqeATfPLo3+95pnIbaH4s396nUQN8IF177uSa1WJwlaNkJUJXRmB6XM
esK7MJqZ8ZLnMweKyQrZWAD2bMwKTr2CiuZTIJd+oYV31CmNL3btDIHnD2dCjQm81MXROCDnabbY
tJjm1mvVmYrbfIeccCurjrRuVKgU7CAVV9lUz6lVCJG4YVtZ17wcYwB0ItOzxKKv77GgjVfP7L21
KJsFEXDSt7ZoPNxXOdCsqN3inJHzIJuxEej+8K0wQbeL/2YtsJJjLh8oSk3kRyPLxwK4HggYZHHE
CkSvhS9oYbVV7XZMBuk0CwjLZhuns/fhI60qAh1pRsRSp7BxEUnHHTGuP+1kMplAJc/v0XpvW51X
XBOVjW4h3QGATSHyYL14YGEjJdh7CtUyt1/fenz+SBxrPu5Jb3qAApGmyqeszPnVFk7AZMP2rYO9
oDIZhstcCYjB96AhzbkFrdKzXWGPN/9Ha5CUO9d0OKwRwKEpOLpBpTTIMdEKDOoHsd+KNK39ACkw
vPJR5Ita3aqSmn3AgOrEVr7YRlU6LWhV0PyPhzDXIKIe82F8Skwn1SaNMAIUAZ11OaSPrW3pLIQ+
wXjwjXN1ivGg/SO0t6LY4fu2XjhOPGF1zyStNum+Hx7elCpZDMnmrKj2+ENwnRAEHq1SMOZjI6pS
mWafIdtaTcHGc/07iEWMLJruBahBdR57JgggrtP5SDMa54to4RiX7q5OTjOJlunjtHtjpys4YPDT
mxC68ECQiFmwGQv9H+oiLRTjbbBAEnHMfnEM23CtUxTY4cdznMXrWfX1Iwk2AaBK9ZWthFG0QeT/
ENWV+XJVK9uvxIOkI3F8G5r4uz8GQ111Eu2B0RjWAt1BUgRh/G6QMJZ9/yOAHkqnBP1q/GomNNR8
xoikLg3LtZltTh7Dzbl3KcNqssgdyIxbBiywVuzZMjvgmdpHjHv8dJeneS/OIgXctxKuH2etMKHl
qUXYxMKML/hbbusBAnqTZghz6vIf3USRjQU2Imzm1ptLR228mcxtc8lyPsBpekeL/fDOLnEXFK18
gQG3AiI6jeOFOOZLK/x8IH08OzB/kbckuwyrhZM8E3oGKaA7jOsnL1MXfcLTEcKlEdegD8hCNf8I
ZX+PqIFjgk0BtSnmPkKbP6Q/4egADBTcXS/kzJKZuIOQ/1eK8jxkONP9ZF3W2OHOCa4ZbBbnJJ49
qN0ySyAjsuOcRxufU3jPpI06GlAOVI5UEcKPu6ne7h10LkI6MNAVA5XGy6cpRZXTjpkUYLtaZmGq
xuji4HaB+N9TeZ81crauhi2qoqNlhr/oIv5aYbayskpZmDmiSbB2HB0gUJMzmQ0bS2pBn3URKxyb
Zf7f7VQfkeJwt9WxGI/PnBT+N1wAW35nILl8eMBmnJvo7ky578+oPl/PoTAPRE3rlNTxCJulMBDf
w1uGsTa/QlqhfWVbKnpKFIktgAQ+YksZM5GH6ImA1HBeeB9ESYYE/Upvp8J6hv9vHCSTzGmLVAAd
+YIVuSvNBagDBsqAGW8U/cnhScYY4BoZi04kYPm+flOC+YNaaJBzE3aPL9YZQLOVm9gUR31O2w6T
VoIRpKBl72K75cgKJ2+Gtkf5sk+/bhnELm+c+M40MYP6gVP8lL5S/90Eua0Fr2HiOvxwrMBgD1NB
iZ+A7EbrPRxd4ooxGK3UgxlRB5xNL82Wy5c7F6k0LY8Xni0GaMENv1JvfqX0y4DKLC203KfaX7Uu
XSvzIsQd4NlA96uH7OCOAagMvJsSLDQXOOALbPGmjiGRnYeNqzAc9A2BE1u8seGfDOX5E7Gx9KFd
03SOoCGh6ZZWvr1Ipl2AR+4VjPJBJBI3AF/CuoSaJBO9nR1WtHttjCtxDiN8rKMGEog3tmDrwqTl
SzyKk27VGJcKoWpDY3f51d5XmKmVgUFhq9OQcUmkE+AxJdQu6Xmu1GC8aE+gOmHupj0H4bjjvvK2
dGN54DndRHLI+WtSUKV2FxImob5H+ns2C91ymJP8VCOS+ldOzy0rQrBEAqLbrQGc1dsnfXtUvkFT
ZAvhNEg4UYHTNH4LUbfzoEQ4XH4Y8uRmTyAC4t2yNVzEIwC0nb5No9RNfABEycSGDO3oy+WVfjdl
AcJYNgh7VYeaO7CfkSaxRCvCFe/lB45ttUTkQm5eDXJ1s4DFaviT22oKL4VpgzyM9cNX/w9aJ+RZ
a6L/9iTcuQK6Qno39PlXNH51fQFL2dBPG6id6ClabpF6Y21Jko+x/d2XBrQ1mEo5bCtPpgMO0iSX
7ss+MukisNiyIuMeoYoQCbXpPrmnQyBvfQH6pniXvsjOlsBEZ/iXiHJygpJhLTY7+s3vjSOjXY/V
d27WiJUUcWqdv/W8QDfZROXg5++DvnlSKoQo+jRacC5GhSNKiW/PGyxGD88NvFsmXZBr/btkjsHk
vFxVVUjN9PhEvPKvKueX4njYIhDVpiW8KMHpVBiJPXXqKLwH/vrUVm/P/H2Z3UfkXRkvW8jMhgN/
nMz6WI+NbEAq0wuR2oUi+APftdmSQtZ/pAAHY9IqyGatLtLX+5uMKK00sD2OIi9QYzpt14HOnqeh
jKOhvvY1H3kGNpB/KcMEZORpAu5DQsJLxLkEFDQousbH7S4fswf05UTM+Ef/aaUV8GZ3RKO5Sjfj
2WwnG6nOPneCrVUFi/dGdoPsZLHAV8PXv1NsxUSg7fPhSrSggaRyqDRrQgpTwwVq5JpXDETWNWDL
ehg8GPrPxlStDkutQKOvvEBmuTmFCb9ZxPgqlf6O0PrH9BNWdAQ+ZvBVpHsDNltSnQb3B2BqEjET
M1oLDeISizxSHXMJnGDIR51LiQoRB3ibGodzD5USRWOOfRtx0qKYIfezPvVSUtrABonLJeJfoWuG
14Sb+I50TKnLeePUkY9kbwx3lmp4U2JWT7SNwYvrEZt7KytFdVOlhUNi/v6dGb3Bvh5sIb6HXkZ6
EoEYfs2M+hfZs4Ao85nzKFyx7tSeikhBweOCjbdzUKdmy/7TKwhssKVxUBT0B3urHf0MAFRglbNo
kOlUMRKiF7lORCjQCPfJtaCSEhvI0YClpjdC4YKuqEwt3GLrnNoKy23oRymxNtpLrgwUkZXUkl+S
Z0bKZCn94UYDIjsKBEyphhe9hdYOAaS9YA442aQ/WuRECgIaIX6x/d513Iv7YQlcdJvM5/IAgPt1
rFX5TU3pZ+7Pyy2xxReD4aEeikdyqpYkDuX5XHyCrUmiuXRBdHbUe5azhwqZ1JIHTn/nhgIPKRPm
4SNOKll8tSGC0P/C2MhEdGmYsquTtSHLLd8UP9XpP1yIxevub9QOjJ7Wt+/3Lg+Un0+EffYBY4tR
i32jmQ+G4jnZIward2b8UJuBuiZ37jOydEWQMOxTitLXUCXN7YP4hRG8Cc8UxuDvWB2r0zivY00L
t9Pp8BCZpA233+jrkZb9fvAKQxQYlfEZPT8tS//ncBWcEJHnNM0zcFmtTKBNz13RO3ytfn3U903P
7Hbu/rXLIIecsLrI7ohFD2dg5jpLMj0VDcZtEJqzbFtzVZhm9p4E0U8KVF+Squ2foOk0JIpKMzh5
Kgb7t39tcIGcyoeptHgy8/Jtm0Soe7MDW6PS5ZLOYDULy7j/QvbMGwzlQDp475R0t/ZtSuv4HiZX
pCVd/kUCe408Tm7WCQqqoHMBddJwozSMYDRZr8puH9tUS6G+LM7sGZotjNJqcSuwSjUcdMT+GEQ/
T0zcmUuYv/vL2IcEGbVV0n+IzW0HNin7lEKar+UtlmzR4AM0W9ZFjZ6SCikzYJB4UDKA+Rto1swh
F+bArnsQtptpaf2tqRCHZKn9YXnreBN0LN/20ioNcJ88enOX5V+HeUwb1CVYvQZVq/3pU3maoe+R
yumPbCbRtGjRU4z6lRbzstUL0xlP7TNjMCQA/HtBt/hZuxSgB7ZN3nkkBYUwm4ST7iVbXnl+Pr6U
iKFUpKdH2rpTx9BgEMqzSSv4EXVYFMDzaZ6Q4JYx1vl0TlUt6g5xUH6VQtxq5MPfLWtY4ESQ07jt
HD5QeIWC+WhhM5n3Gez1AEIXkmOyJsSyFaTCJlPgFs56BEf1qJmFuLMiaaHdtlcKsJsRcAa/Nuim
5Fj3TbmZtcO3hqyCm0+Cs+c38KSk33jsYBj5BqU1ozXiJzYb7Fo0PprRJ9E6D6AxFdywS4cld+6J
SToq90wBVjOG3+MSxRB3eHY/sdDVyXfHAnbb2tTgqgWF6AhnfV+XnFAJt4Lm35x9i3765rdcJiVZ
Bei1E8NIZ5Lx31M9EnqMLhmlxcFqjfmdx3GvGvCBaFPWTorDYj5F8/WEYMpNK2GHPACOhUWTpxZ4
mNOG358BgMuqXz5x4R+/EkeMd/RO58nDMWz0qElua1USXw1FKbu5dpVA3QTyfRRMA+7POxbG2Bkm
4lAfp04quxi/sr2Fmvch8VNwb6+m0Z3pq5AWTMvL8N1so27jErkZuXp8bug6KzqR7lU/IIlYUbl2
f5qrwEr+nNb+jx7nxh4I3Y6Un1CZS68/PhtiimC/aZB9YTLq3AVXgXjUd0HPKxHOOv5ufND7C7lA
1QsUHTrz/CZFkrEGpFydpiRA35yj6kwgqSaSiiQ89oT4WB6RgCcGhn4B1Ukc370j3OWJR+YfXVP7
bCyBN1MLM8muk5a86fGNOC3S6Sl0xnyVXBKdGi2cyzClgsx2xcYpkA55u6TZyo80pvk1ZCOSKBYx
N1Do/CKeKk5odmkTp+EM63AXtlNNVBnCAWHBbrc2JKJPG04f2I07kCedUN3OnjZEhdMm7KurXmVm
uRvrlULHPNjSxG8GeWRv12ENRwrI34l/birkzHD+cKHWoJvcbQuHVVreiKMoeej+x6wOCKG2jkEb
yzWxU1ZMdJY8R1/pYAXwVjGHLRKmhJoZSKtf9bCnHkulp+UMRCFxqHuPKV7G03GmGiJM1jImHul1
v1+hN5xVS17/g0iXpd4NFMmew5R+SL5yqjj1CQiTBxlUd3llL3VFePDDHRwMPavJr9zWUcD4GShC
qYDxsDFg0HYpu7QanLwrcZSalg0KEifwSo5YP31whVoKEVePLmXkWd1oYphzlZgyhUv7eaSwqdoi
XAH1Dswa/fecbeGJkDqohtVf/qLNoRI6LIX6JWHMAaqgT/ZnI4wVU2OZ/n3/v9WYjqAcGrGmIyKe
KqKdjxR+ImVU3zXiPp/J+k4PFj2yrIFWG9r+A2LrAU9ggqaoK8XqKWiC1Tli1QI/McE8pOjaB1Cr
1aHlM4fXjQ4GIq7cSzgZMs1Map01kUOi0bs1d3CnLnGP4twc47zIGhCAna36syP/9t0jnYhEWRTd
JDXQEKk6cmJ9h8++GB/X1vLf2mHhYOuU+ckGqdZ89Y6nDueAYo+RIYLPDNF5HxKaSDdaC1iNwbiT
PnHBpRpPA0SNom+0EWAjlm1I0qvpps514XHuGN+MCYxmlNKieRnpjp6WKYEEhi4TUlfzDu6z4C4t
R6CbSKbSoNH4dfuiGk6Av5foteFIhaUIjKH+39nxbIsw4yeLHGpK+UczmtX0fb8V3FRjGfHes6tk
jBvwKJxPIPTZhstK+06DCs2hKLcAzopprRgLsTs6L4TI61L8rY6o975qs1BmNz274x4M5ktI62H/
bHglvFO0b9pLY9xaufXzJsCLy4KAzcYOdX7gYpfQJOi5vb9U9/HILluakQ/Dw0tLGQ8ytlH1WVT5
IO1nTVoQsu1uqDQF5g/CAvS4UqOrpTdjwj0TXco4DAf4DmzJaulHQEZUbI2znZ3szbt7T81H5E/j
PmiMKjL3/BXqqvRIAxhSVkJTtnLzxlqOTOuDM/s99VrABNMa01KxBiuaQp8lw0GNgclc9Au3nFqR
2i5LW3wgO7qHiLf1NBQ4CszIz9MxwHRpisYA6yH1e8r+UATwQ8laNkbAVeQkiedCDOSSkAmDPZVX
FP7VreRdkz3U8cUhFl7bMUSJCx83oNbg7RfsSKEYS1TshMZJ6vAb8IDJGl+ZA8bRh4q19SG9IVCy
U7/17mpysZ3EepYfuRpfa5SH56cQpEdGz4MhL7BmhaROldu/2ghIeIJjleVkh/oMx+cb/pTQ6o1N
ZWNDm/3LK2yZuYD9VMXvQmLc+cb+LErVHY30qFkJtqMQ2op+fYh5ON8ivxUj9ScicKs1J8uMCYbh
/sWGOelEPh503xZgi7fbGjas+RL+TFqOvbtzjLgQCcKiltQxZ2vtfjiEwZBqPhQo36zK2Md5NH+0
jBqDrzmQlMKGJreCcGO7/G13qs6IiQzpU8dcG7LL63iJyVLofsh/cpypqPjXh358+LrtLh4VMRaG
GWOHaMdxYkslNGsORElm2UeYLZdfVmcj0Xppb1KltBfF9jHfpDOpwoQrj566+TApjEylkGzfBfAw
pJsRKOSoZRik0napUdf+TtfM5F9pE3EIyDrEvOiR6cTuowFGGOXMp8FXcMU+rJhMpHhTSCK4ssk2
Fm1zea3d0qmmJ0oF/oaJ0NH5oCBd8w1xSH8diq0gHDYgl/KbpOapOIfSB/QJZs1pqvwt1C5hQ/hP
dIV08kivxm0UOHEc2S5f1zFaulR5NOR8kzyk69kOB5LKWpnK9F91rpl7OZIsaLdHUT2ACI+n6MQ1
EKvXfywJ77SIZ21Y+O1PxaLoqiVEUa3kySOURQSUGxrsedZi6qrEfKqFZukuIKBxJAqhNHY2ujY2
M9rprLAasTKsjSNxwyyzD0OQGs0UEbv7LRd3AnYb9+Lwrp5CaZbIoNLcx0uMz5qOjXnilnsYhzty
/zOd/Qdh/34OfZcre9qzuKWzHSC0KKCrfS5v0hUn3eeQ0lcXLxFe4ZmVPTDM2EBPZc0tt0XsCtn3
ulDcxxlNlnTWx4GnIkHKI7IvfIVuIJhSnfTofBXFy1jgPjzuFgVqB6mbRe43Lq46+U13OtaUg8z6
I/Hk3kJaAxiFi1l2vCmVjNk6T5I3P+Y7bAoJF79AAaCKfdQNMkR8TAn9A8gqpDN1ZMahsxt+F+gZ
XuH5Jnc7L4IBi9TQN2FnzKt8fgrBXq9Bi7mnBKLZZ/oym/+LT918sz5hGNKghCpFPKdrtHp8sWwb
e3vG7GcFSgs4QB/zx8hiUEww2CXEcaTukWsPqDz4iLxsJViRv6znoeyBisgJk6m9q3ArMW/LKR4L
onGP5NADfZzaINz49kYl6jnx84tf+BJ2U3p8Xj3FnA5P2HlCGyCUmFNxGAURKI3p6VGX2mDeadOX
fLHkCRIXgxqtfbVxPZ55WTlqJacdQT/ZM/RP+3W9mFO05FJH/R6gmNWMhWsNdd/bmRr45g5yNEnV
We6r3YI86fmRHervP0hkBwMGQf/Y3TZJ8bC/MT3hzdtAAWhCLOHK/qojjuWWuLD8GRCsVCpexABO
7XRae40la6CfujNqFUvk6ZT7CloQNo59/szfAslVxzZ+i8JCFKl7LkuxlQ15GckCezJNVLm8R5Da
lzyITn0gQ5v65WPMgPwiru2HA5rATV8fzhTwj2KDISli6eKEoOSjF5ZD6hMJ0TxNYAmhmWHQcCTz
YpwQJL8G9a+aE2k0DNc7BZ6zEdcSxPyULR/wrdR0sBPXiV28ELCa0KEQBF3iDcnxOvKyi1ztTFBM
dr3Zvz63H4SHCYQPtqtoQWmHAkgnDeKATTT6WYn+KGXS3T5RxvKZFY5Vh92I2L1gyuAZgxo6G+Nh
bagHwHiZRF+Zbw1zH+l05oBGsdIAsfNWExOGFkCnjvWJU6N116EzNgy9iP4FkNQZljGbN/Swee6U
Igrtr8NRsE7SX+J0i78l9oqLV5mi4iJqvc7ms50n/v+5sQKD7t7OcugANwDrlvmQIByhPNpmBwIG
axb/O1ETjuJeH0YsZh4KeISFZgUl5E/wUawSvHFA4WI2HCHsSjGt6rApAl45inO/z6luVAxeq+uD
BSdgRTJ+g64VcGAFOD51vof74cgFFhPVCioj9vMgjaFnbuvakl2nFtUebKhkJ4hFZDm37L1l30By
YcLW9+kKw9gSqsxaqc6av05ALRsdQ+/kT1xC1D576eCt+6SL/1870xKKD6vO072cFRsBgCFHLehk
wKzQc6dM0c9m+d24bRNhzdlP9Rlwps/RhSMvp0kxYYDw+STjdq30qf7MHhkU6VI+5CeJHruUY//2
WNC9RQ7RuvmQHnaU4gZHMPz6NsrGwioHeqI4RL6CBVDXlCeeGw9JxCcXC0CQ72gJjG8xXB7P56qd
G/IQVjFEF07EE6BipyFxhQEBMTh50vrqwEH55at6K+eqxJwQ/3TY014p689RYZQ8eZz1QCMdAqxp
TK59veQoNNxhhyub18lb7xT0HD4+WN5WLrL0qciR58ogo+UDsO52408hNObnoHfyih7u9eku9kiB
zV0Uq66r655hEuRPWglftGF6pu0tQQr6K59tEibZ2BUhTpkoV2U8CdC9kdpb6n7OwFzgcnSRNm6A
wnKdBzlbYQiNfPqd/CdMP6/18YjEGEge/VHMs7SyEIR+eg3zuA/0HpOFv7POSQEoBJCRn5uYzCjv
5ZL132PrJWCeggBEPhlvaYD6h47F+f3x2YwddnLRI7zlK13WjfnxpBU4CYvq6sv5LuJnS2uQWZzT
Qle1wxE6+0cAOHfPyB9hYMYPaeICnP5DjV9+VlG5Bpt7zS8ERxlnu8s3wVmcV1G0fkcAJKAUp898
yXSyKSABWIK0hNdz36LTFtUMGure3FlWfFJ9QQwXYQ+3pSOmKEn1vNDorjRwV4juCmIwuv5+/Y96
wDBspr5V7/yQMORxm3WKEWFDpuvvKlWsYTXpN9vzuKGK4zbaHhlrb9hsVXOFnYglPNPCt0yIxnuN
e0lx1rNSwPWt5sRTr89DPjP2fmszPG5WdwTrTDdxnRysgLdzhN0pgn5AVESFrrFBTfrTBNbCsAHQ
dguH7ZA9fWoQqn5PEtEhAnDdqV+/DH8QLqgtdN9X6pQK3HsOYdL1gpQTyB3p2zsVsihR2tmZElYk
85cXFqEn8AovI/JbiJtga2mFuGmm0/RcyjgAnVPkKA3N+PGumZ9UJ2pGc04vEAkW3Xc7QXPrkjn+
82+D7waITyLAaLGBZjU6KxC8vEeVX4XjdVozIkIrEjwmUUkw9bs8T5KjABZuvjMZVLo+YuIxr2br
ZI4T4bI33uCNeUD+LrjK+VzFusLHjSY6Z/zj4NwXlN6Iyb7o/CzhGMBGgU35Mi1lM4MDpOOZ7i9N
C774sbdvL7G3WMAvI06jHR4N38t+dxoBt9Oiob/7v0lZCLE2FpwpuKHp55gHPgoc7fDRimEtkA0I
sSUFs9b/HYpZUKVKHbQ1DEM846P60gcLETwNtKTR5njuVktr6FKF7hXkcU+KoUAshNtwdjyFy7oc
pnI2aUQrZ7jShBLyF+NmW29C8a89Q0M6JekAG75h9AIoHCg4c/NN/NkBd95iTSmLPeQQYV09W5oo
ff+vUbptYYh9wEWspWFJei3TVTOC3ubB43vOxI2mjgSHjUWxMc7a/aKAYl601nO0Pwj1xHWv0Rj3
WwaD5flhSTMgqQtCwmrDLMFoWwmVG3Obsmcwn946WDGQutgUSX+qAMjUyXqJlwKTFv2y7HIekkk1
gg4cXJ8o6waac/k+hnUNzAYx4sM+t6d8qTO7Og6HMopJ/eSHyvtq59lVo/ww93Rbewcgtp8X8TCi
SvY3onIdAmFJ/GLoSUiimNINDR10MklJtUkl9VB7oji7OxIjJXsXV6xqHCScPzkg5+tDq0j2zG83
g8kJa4S4tjj3Dtuj1BTsuYKMT9Lp1E8js9RZ37NYT06USzd0dp0ufsU4Nmhze9XsjPv8IvTcM4kX
+ukfBy3lF/YwHobM+yKbnvMhlQEl2WoEckg49P6NNt+sHkAi1eRo31h3mOsSUAHB0hhAFVfBV2Yp
uJz4jawoFGqZT3ZYazRYnYfgRfPUsTXVJRgPczj8BFr46T8QBbXLzhos9EFjbbH1TvDdGVsZa/Ro
zn1JP6rkBWeBYXqP0pQ4BtyQgH2Yc+JpUe0x/NDeNAGOUhxJUCAI7k1PrAN/6wn5uQ8V3aqEf4Eo
2JeRToafdzTv64xJ/htiUv9tNfU59e2lkfm/vJAWeYZ9g7fnbkfHuge8zifR5TYGOdPCtPTif32y
dkt3yFt/7p10O9oJ8V26fvgn4c/lF+hNnwYI4Bw+miR0fZxuPxrZaHp3VFFa8Ro8xPqbHd6bPDlc
OUpenFOoYMdXMHBSLG1mBuKYsoyGgltTCjpCK+VF70uwCeDHFSjAdytkFYoX7x9BgBwlKqBGwvZt
/ZoOaMFmq2Gv84S3Yg9ZtFDWut42RhNfk+E2XE/zrIiugZTHvkybsEkGXJX99mgsz5jl7BEW+0NZ
YAoIj4tWDRs54DMCZ6mtFA1ilaU+asadIKoZPKx7UkCiBlDPCnoMFiqn6ZsY0ShdE3ku9z8AQ558
x21QMzRJs0Q6+G4GnkcptZs+TcBo3/JgSdkp20jxmLxkdraY9HZ8HKh5/qpPkRCpxPYn/Dxry1dh
zOnzXQnPgT2IszBYd5IN1FeUBSAoDnqzv+ZPUYeYyJCCtutBaqJXlPnn6gcCDEaOKZw/uCBZ6nho
ZTfi5YQ1jNq+F4vP5KhloSnXBh8yceHaNfk3LaLaL1i65VRxNEW5ovSvPQq5VM/NCglSfDx9foqs
RSdhLWKfej5dz9Rrvj+Z0FlSzV/n+8JDhIB4NLzyWC5ojOtOqlV2PN30HaD4UrwLq1y3mhHkmkZa
hEfGEBcQ/jY+GCiSpnPCBLJig17tPR4h2LcW+tRTcRtPqRVzIgJnfQzX/NC9CSfiyKcev/VdNDIe
FLby7L0hoJFS/u35sedXxeSi7KRz6FGEJe/7fjxnqH7hKitZqYHfnAB5JoGa/X5XINPfOlXUNJAy
24388PnA8r1GnpKqg7kiAmu349qVk7ZuztpKD2fhBWbCNG+6mIyD8w4Rfan5T53qnCVTBfGoXP4j
S4KF91so+wCIadFeDaYEAgLQB/7nGZv1Q/ChxC6mPMLtJqx3IJAvV2LaFbJ5xW1lgrozMT9JwQHv
PIs+XgFsYCq8Xmv69822C6El1UjFG9eS5ceSfMiIoMPnTOWTDzoxvn6o/ho5OwrQypGX7N7fxOlQ
6jz0yQ0MNTw43o+5zsXQQIIRHVuRxDUheoKLnrlCoiasLYqEUW8e0MDCQrXmjiOWs1KdmKLP7Tdm
BMX2KNnx7XUFWzitE13cVyXEa8DrDVVLR6ez2P8RZ+vWF3ULK/V8N0blKHjKmerYBa06FPaBjflD
D9eZVfSk9hVxa3w9dntHLhd2cIgp4pYAekuErsGb3pTg3d9/tUHELrAeVGPb7KLGkXIh034GuOTx
sMXAVhzRNt/o0kvxid9XcDUCFwj1ogdcUbtTuekMc2HFHpvjQbayE2vf/mBtRXEZ79k55uvSJf5m
cgVtR7VC02rwXX8aO2En3iaCFpJPLoKOGZusif69eqo2k/ljodvexCv0CqmhR2BNZN+JWb1ZULha
3EEZqAkgMbGIUxNdcuTTR63EZ4CJ/JpknSbTnhkIdxYhq1Oo325rO7SUbVzGYOju+qH1UeI1yPUb
1soqVS643X9flgCXB7Ryk2zWk1GmQ0p4fmjZVZkFdFk9WKkhJMuZcvNOJh/lP4OtjrwOkRLQa769
3t2d5I+4BIl9YVGrHEI3mcSjP+APPwX4UPTDYAhLhcLvfsUjKrSEQLIJ01Y1u0NirPaL5TY2QCCx
JaUxhq7zFcpvvI9Tc8JRxrkZ97L5sOdcx0ICWBzQpX40ehIXyCn6YWptQvaBIYCv9RHPIW0SKaVi
xWbgFlggXZ7G7C4hFauItcGFyqq7Y/GDYuhMR3OccA4o/9L4GH6A81fsrO3RQtAwg+qqewIrTttb
LThaNNJIcpupszfPO4YjKeotVZFK6ZxQ/UnNSmzCDkoFfeAPB6wGHabac4JHuEY1N35nDo2e0LQC
r7qQWfbXTwz1Pp72A4XFpA+/oIhT18BUJQha+vm0oju46/EJY/GjtkqrrFFg19i86xmj1TvOuepM
eiTU5XGE5mg4tqavAeaihh0/fYnD3nxi4Zi8zg09KScKDynI7MNCbXkavjQQcO3hqP8AsDDiYRKn
CuQEYamvzgdkwfbXeim01jkTvEb+Fwk303WPPHyZLwHnkYJJt1sC65H5CfZr6h2gL8k/sVkpKLLd
5cVvIQh2T2AmDwt867zXuFGxrttVMDPBfQT8LQ1JnYurJleKLdVuCFMMPEH0aNLa41H5P+BdfV2S
2lpKqXVXPFe5BSsWzd6NM+35+wx0nnGJRFWawKN3GxKo/fHXYjPbhyI3hAdRTXTsRqg+0f4DptGs
gfSe1Cuc/HM+qdomRXyoaODZFMb/U3xkgxYtukwlsU3Q/6NM4O4cohtWtiD6Ldxphpd3rR0FPW+B
IhgS8b5tN3rRR06Y++hhhjhL9pWoREik4QcReEnbzJMckO1ktf/5zW2v1JaX77q1qYsZb/ScJZbf
pHwI35dBr9GYAFCfQosxLZ2VM/QU7A1kDMXsmQxJNUvs/1IBsnAw7oYCDgsH4MlF28nN3pEYW8H6
dB9Y/H7z/OYWH43ISSapMkVAL4FPrAP+7Nx5BDnFlS9U+6ypts/x3G3DGlun9CyWXP4wen3RHtOa
UuVdK+iEuaNJP0uwqXbqwVPiowSpo9mfqmDDMXQxrRjqiYtftRG8cKk7RBmUyhf+nD97L8/PIIG8
btMnzC4/BXCg+KDAld2UvdgBH3C9qm5n0MdT80ITBc1rth8tumtOwAlh235iGlsFeRYKPJc1onw3
DVxOTEmNjaS83NL52HZlkdkspVtr8Bw+JINjAk0tl/iBSO/4pO7VeH7RAJVPX5j1/xccvAXlVinp
QUQHGRLOCnP8FnEbpYhj6j85FQEk7Vh8gSJVUO9YAmkf/c50Uf6k3+spnWmGGdV6suzvBAGrwiTf
A7Rv/p+0nvaZGMKtBEEx2ZjLepoZdqhC2Gl+V2q5uzhOKqKpPiZ3kgrn21syBkwnLGhVzqJifzja
VohfKXgrtyZKBFoo4gALLR0oAanaWKBHkbMO+4Pp+0K6u2U4v3NmE+FZUgC11QUolTgS4XFkDQyI
bN1fGmhU89TYw5RoeNnpUKoQRpPJ+MPrF5MQ6VvWkOlEH/Ni2BInGfhRgWnv84ySRwVbjHrxq6ux
+pzI6AxmgljDNWOGwEdGaNWhM+ocqQ8nPb0Sv533wI2QhS2X1bn6C4JJmWgTBLn9jShlssYDvFE0
iOEq0EXh8gUBWcnUPnyA3A11MvXViclg+HsanE1cHT5r/JzH88c8ANT3IiLGfcb1J6GjGi0mHM4d
IsY3JTyJNt498KvpYv9qX2B/K7OEx7EeQWkpZNz+RVMLddTrY2Z181G/MoLBUwJOtLjsCDtI+VhT
riqSYmVnnqWprP4yEEK0wTSk5NZ9bW5I+Yc8mB/GFgs22oflKhfyVX1/GLsBXTr5AJ79Gwt2Wky9
+Oqb2+k6SsT3HRQ6NYm5gSo787acTt23uyxEXaGWoj7XJsiPLqAFsfHg4MUuoMDB/EXr3xzxdMNn
ekn10LI8fisnIPA0NUcC2WI+dcMN0kD6M3P2AjMhQL5my+Thl8mF6Iwg+NhIoPZsyL6UJM+pgeOG
uQ/0lX5pIbHJtYumUIbXyA/5Eg7AQ/nxWBCWgd4dTNWw0fKzSnLsMy8d5w2Q52lo17YiQrQHKi3i
YNBaSnBlIWzJx9jyabOpe8287UehxlGc7Wg/6glUNHfVv+RN0FV+YezfBX8C8MIv6IBSOBi1aoCR
YHlYqZIksCWgNe8GQn5qqnMOQkYUb+w6prTkSOLdp8DyFMSbxtKHohfiDAHNW+4KO4WAgubM8WHj
QYe5hSCE97iNIWP+9oOfyknFHrKpmvyHhKYLNQ+2UQoI50s7Bn7bxO7lIRpl5jF+HGDWNjNb9XjN
eW51FoR3K5xXwgbcSvS2epqqC8OJe1PC9uDIvToeS0oq8Am8/DAsCiry6451koe9m90rmgYn2laB
fZvQrJVyWU+Z9ElztCcwYCTiFMJm24Xe9gYBLbdrn8E4t73GWfiT1S8chorSQg/o7fjjCvM3mw0o
5lmRSA7MEIL58SzrCj3ovDMpeltDIAWJSf0jLW8wWoqeoaNV5YAh02I11qj3790kbPq7mTO9yg7w
qJIFiL7XOUBkqpvjKPH9IxDeebrKoX0e2ZEswZAeD3ZO8dBpvQddA3NfnFPdB4D/Pk474VACdId6
BHNMC7yqJ0lVxp0szMkzGuAhms2l87/BJ8Ylqbe4NTPZFMsrYSXZ9xFpj5elG/MpVDejCpk2Rneq
34SLiu/F3MDCi3Ty9NMW71wQaiyTOf2qTJ+SkuQOSYkNokTf0LSMdi/QWoWjC12ipouAbPZlPVJp
PA+0sBMKLcP2iYeLfUqW5zk8Fy0Rhjc5YVXKhrOOcMd/6gUVyEm9zgI953sNikOVs+iKflFfdjkU
lc8zlZND7ya7pf/PO62iHh/phT/sgkHbCRqg+y4fPY9yIXmK3ZfuG+tV9OoaekuK8CHo2srERIoL
/Yof74QbPPjOOGPWNB8pMwkqpj7juuQeSrTDW/XlVFkgqatzch1NoXNve9jNTLxSGGLhCvBqirkc
lYALcKqBWPJGyZBNw6kf4nnOalAmF7Z3ir1SREvPdvvdH9fl3uBe2kCuhCAj4KN6a6dGSyb2NVJF
ZWzaEWKIiwIKnK95Clq4dumdje04MdACo3OAIgz3m3DV71m6410sh0/XpZ/Nl2jxXqtj/AFvWXTd
fHbqANdCeET/CdhoF4QmGISDRexap4RxLotR59bzERQypSqTM19or7x6uEqWfAyhZPF3ickILDmU
4M2Y5UxdBx07q25gGU5tcb5VVhFi051OP3O/ZtJ90cqTmOCOk8msWnksHjruvtc4A03mybtCj0By
3cPFhZZSMYsme4nteHje+KBSNhrQoH1FmyhTNlYvYoNP1mRvZHYtGjTZ1MASSR44AJdf+DRWdCz5
0wmxf7B64oJg9wTTr8j2//jj1cYHyPKYzEdopIj7ipYjFXDRQlRgf9qM/nbqSv5KA7/e6xeShgVs
bMpOaFFeTfQRFM5QdQKqlOcF7Yl2DoedcI9jXxfnCo5aunL4VqJf/fEmGb4TSfXrXNjeTJTiFIvD
JiBvJrduFUmVjgSptfG9ztdf+1+zoN0KyEkwtrxGhz1hshQTRwEukIj8yfzzu6TxSLjz55cGlf8q
/Z3gnN9GB0YMGM86kNdUOKFHnotUe1iqt1yd7cL4dMbiLohvvPmhk+uDOdFDmiDnR8wNy+Avbk6R
aqEOCOK5rs8HSrguvLqqLjyBOQeyIgCrfmNwdkqVEg06OcN8LaSQO+t+sjFIA0TPafF9yLwCV9bb
42eRui7ozMmcb6V3etfyeUlIojwPbHXr7j/KGNVCJf4KQDLNe2FwgSEWOPDyuUY448DyQoIooUzI
ZHI5IiD/pJmePNGPk1+e/SKsah12A93IfNW0cXOUg2U3deh7fXNwJChyd7qLvUI34cXsNHZYc2rQ
ZG+DI6yFhnLguQpsxhcMUPVenq0HdxbmIcKylIZN/CaoFq+U0wntwQ1dOv+K6GrfaMutWp5CCZK8
DwRALwmdKFoiji1iPhS7SqePXUacHMCl5Ip+VJnJt5mY60YojMzvnOfNrENcaDjnNGSjq8hYig3C
/1mJOyFuYCzAlnMU+hGqs8T5fElYFagSZRtN2lik55Uksh4yrFDQvJ+isEnXgCRznFl0rZkOIu7g
MPE6rv7aNUKu1zhfsOeil2pG0CHFVkWRnkCIiGL0jw9wq3tDEG87cXbx8lfECDWBYaueY1XHr+FE
SsbE0Z0r+3eQ3b4Bx+5h0ZWdVSpCcRooXu7WKWw47nvpNeRta/oV6ASfLHcO7aFyZIFGX63dMsUQ
ff7M1jJwXVFlNfZA1gbkdLCOj5FhZmY7McQQ+nPzj2enQ/kdjfXO8Lx/UyIZmttX9JFOsfAieyLl
9lVzf1dEeGfE97xcyQV1Hy67GBob0PCoMZhg9yBTf+g3x21cvrOU+rSUlkAux3qJXCwGEN4OK66p
Zg5DiG3h1V4cErVxHWQPCK/BJjEd+ZM9I7eSwJbceLC9XJ7pnBAyw2hzwkRVIjPKL1Nt339t5nfj
7Yy1nbZW6MXNVE+cX6XEAL2xlbgimQ7OSSTAJ2PHkZKKzDxVFNCWxrZn6NP82r0E/ImwS7+KRH8K
2LJt1iv+Hpvl2+Z/V1DBfAyj/KHjXXlqWYl67Ui18gcZuNzGrE3sAkk0BddeIu9CikUxVrDkZcaX
a1wj6GduONmx1NlbZh5zob/zmz2sK+c8lRAlxHzX3LIQabTUMvEbTjbCFdjyTNxVQ1vFB3+3Hva6
tHszfjRaWE7O7Z+ZIfp+YCIE+4cBmvKOBKeXZzwNCWWRs/VnKc7Cybj+TsHKgYFhsUdjl8t+eFpe
6pIe9QlRfKd3eIGlJzSCM0gowX6kwi3t6ihe2kNqHr2xcvVFtHh2dvZpGBdcULv3PCducs8MuSt/
QT+BZ7U50kRXPaIuZsY22v8Rgu1rVG1rU1qYy1amERBIjlOT5l+G8TzFU9Q9UcnjVxYLeh3VjIzf
ZaktEOtNGpCvjS1X3RFJ/jF3s5rRyjfyvc3bCYHP4ds/6FgqyqAT/A346RQTfFP2fxt4pafxXFRP
zrECRb98YlsBIOVQbC7KUIoOYhTyQ+s67cAT7m3AlQTd8FH72aKygPdgYCfEdMFlQr6iHbYXSEVZ
QCtxaExsSGQ7ha7lPmTYlSU7Cp4uOBBrObhkuZir4FzyLVIQBtTiwA8q/fcKCft1k2gnWaDjwFeq
iWVOdmdhViG9iibLTlT/3bAhYlwcJF5PhKvGVILhgjWSdmpjGjU4Q9s0PTydF/Xe7cUnI2G3AoYw
46KDjtq6BCbynIqPSESjtlGnAPN/Cq+2F0WMWXXiZhzyZ01oJ7AeiNzkOu4yp548L9+bPCumfpT0
YR7iOWqJ47L8BN/65ei/te95iXMha0+nGuElr9hY6J4yr5AjQTn960Wsg0/0qBtByYpJzcj/7+cL
5xJ+XdJJCvzKNgqn4Tm0qPUO/ZSet2YvyWTN2pO4r5qCS75UiYrU6lNanPFdJYSz2zymNQy7gIHn
HkSGYsOhOzvlwHzdxp62A0aRs6MfC1xYDvPoymsHx95o+hcIyJrJpKGrbb8xSdPH3fy5XfgzsCkQ
h4/X8uNHOD5vZbpfNTnn1mBsAyTJZJQlnaVVDngL21qFd2FYLfsfv4b/QveFI/nIx3Jtctkmf886
SKL7fFrev/6P6lYh1P1O+FbS+ECL+5nMid0SG6Hc+lVs/FJ0cjwhiOSnPp3kCeiaCgcYcOXaNO0D
yXfdXYFcuGQ1rWaEtpYRqZMcjQW1s9k5PL8fBF+1nGyvguo85DP+mMxj8Wc1aJ3sT1y5tXZ5J9RS
NRlXCL++FlzK8HMKmkpIOoqHrci6WlLtmJox6Q8lVWhDG6h2mju+shpuO/sE4dJEHV0p0tsr9n6c
DCUY4DDXd4/niZ7GBahZYQHz9E2VL7xLp/o4SHaIUctYZHidYGeRci6B4vGoiFXcJu10CPUav2eE
en8h3Y1drxsP+5HFWuEQRReMDzB1+8I6P9vuh3YNh/0/7TRjao7U4md3LorhS74Wt6vg1JAFx4EE
yxZF5JhPtJkk1541OVLodGfuYk7k3Yp1wvPxJDaaRbP22vcyrsTietT6EM0ZG+h8XMPrxXB38UW2
O+Pu/2cB+pN3X8gww+rpIBJzeN05triWdtCsu/vmlsqngiHfq5/atcyH+zOz6TLQm8uUVvxoA6LZ
caVIdu71AOOPS8scxHDxmFBjH+/LBHLlxzPjjANWspHtA5f914C31MpDCL0kENT3JvTQ3M+GvDSg
wUbI2JuWB/edufqVkD1ucsHHMJu1Wv9yyDqjfCqUYsKz/NB+vYPQ6Ti2BJy//2N+25etLymwC5f2
MA9QpM62U34Q+VLhrnuaMdFofMebmd/bwmz/mj94VR9q+zgjOmz7a2tPMJrppba9JM/FQU5WG/6Q
gfrLpdD6de2zm7o4+lFWS18KqzdqH4LTOGJzbR9VpJ21cFlVulb2NaaB/x6XIk2q+KR3swplUJSX
L/Bw8x9MVfVxsdBhDrZm3Iaae27oG3SmY1Bo1eG+kXxM6ppf/O2p6TbUN42IlSpUdFg5UH2qCpvR
J5gJUkS2aYD34hMDnjUix6iqUzv1/jDtsXTOrfgkONPEO84KscvHRL1x+Qz/DN5kLxOhsAAJM6E0
KN8aS6ZWRjNQQ1N4FuHd01SMBwsITtaSTQKH8NcNmpR2dNdMKvYC735x/B+MO7FmRmUWZ+LkpGEu
d5utDd5PzMhNOvqQwOx7iTZmrqRNkSuZSUSWaw4GKgyeu3TR3pz7LaKpnRMiS7TaBWr06NO1//IT
kw1crDHCoSOrt8LME8+9ZbBtZ/Ssaesj3YVr/D/7QaF75Z0Y/3eTpe5SaR5WgPpHXhdWBeImGmvg
vTKxPML7IVELushAH+ymO+DhidG3fDzlsMcswjKU/jmsMFJMQsJOcHnYQ3xc056ugRr/tlZbDAiv
rjmn3jwjntcgVFTmeFyfHH5PDR5iNvYjt0o13Ga9rld1TdYoHMU3n11CQxD1XPqcc8E/27i72PkB
esiqizlH8hz/TG3hO8fJPC1DJn4u20m2mXUUK3jzx8bC4IRA7KdnRkJd4werRqIRB4PxfGtk5wND
t6J4Bp91Fh8z47lVfJDqJVcEFUJ/1lZlCJ/8CMuf0jlqTQ02IcDcj+vkU08+nGgPTMh93OTGSGF/
9KxNEkYtyMK3SLV6Fz7ijQTHt/dnH0LKp/pPiXKa0PBcQtShAOZZMxstH/6pIacLcyyGJVV1I8Ff
CLrQwWPkhz5ePhRiHqSMxX/N/xBN0ioyBSCaH5HIMIofhlx7kkiZGJk3acjQGi40sVGFxyAzCVAb
CNAcB4tHK1SnuekL8eCzQeJrfBZ2pIe8XrKyqbRWRBRnwKH/zJ6dU5a0RKwTtO9PCCHAgXMlV1oh
xYdT/u0J7+b4II0By5l75oKbBvEMyDAvphg3cObGvsGw3bozQFsLHT0rHxI91D4IuC4S0WQYhYUX
niGj/PuuXnbSS8nmnltyk6zbguSg4kPnaltb2qTbd3yzjY1L4ZHEIOZRnjhBzo4fmeNp7eT1rLU/
3HJpjez0uLuXTmpq2kLMkRk5a90PSs8j38lEoDsgojQoo+5YTIreQ6KT2LzVZXILzsxliHLul7+G
oo2RlUmj0zlGFw2mOMYKMJzuxIu+Jym2tC6FGG52r5Yfwj5fWe1A/xOfRBQW25+pyxakZXQLsxV8
WbbfIv1uvL+WYtnhsmm9nbS/LsAp9d2h2hIOE6oIA6zvtSk32rvSzpmXou6/PBaauxvIgcbyHmZb
s7IUsoIP6SSnIeqTxjhQryrl+R1WuWnEBnggeeG8s5iT3jZ/upfKhf0QxewLVLdOkQsLlsWSk6pB
6ts0NgZwRuXj7FaL3coJJOwkkDVUiYriiynHA4ahh4ZY5ghixs6rxnPXMPXesOHbphpjok66Kz+4
B89Q4HV8qjuxavoyVdWqczjDOBhjtNlG47MOMb/YBwtyzyA9yxa/YvRsUkELbncQekXA7i8dZeIJ
A8Z81kqlMctBBrh4gdt8doH+nlOYCcLPAwpK/00bRn1X1qmwYTq+yhohSSoG1Uo/09j7gAKu15o4
E0YNrXs4CC/n4neP0x8k20jXXjCf3itRSwR4GfUpW1/gOCovo7TyOA3XxCkx9Db9ymJ5kbSgakg+
EVNmgbDi5N2gdNsiC3Yx6w00HswYS7a0nOFWuECF68umUOeeNjIOBEzWtQK8snmUz/MekiX5Pp+/
1TPrtNp3ePzZLDQ+1q+Bh+ZeoVamy2Hnd/J8GkxCw0sDDWV/dUnfJQ++ATW2CtnqxjSnJlqAzfPC
UejIz/x3f8TG5uxbf9dYea1mr5fuX720f6yS5jAwKY1hdF+E9BWP6NQYlI0VGo/3+Urdg8hAb0Eg
2Lxrj27tee5ddtikZguf6ruY2P6xqSGjdfCtZYKXaJ/UmLlCxoIi9DVHHd+y0w1FKVkR8IvgJqHY
UQms19sekawtQ1VqtugcdQtxlXyWLCKi8x3HstmprFTaCajNKVJLI58zSchuGbENcGxNVNCiKfyr
A73diFxeTuo+D0RNQCA2ZpapTuLKMK85YcQrif2aDSIy7FKsuiss3FABQM1lKMdmMKqWhsMn+2+C
KjTGvISm/g+9PR2AqtmmItzHVucTcDCTbxce+GtWfp9gnIvhvggQF5roAfjiplkvqT3U1n3a+loX
FGTNYdwpchshO47d35MQtc68jMV2ikkZAAfAGLa6kBWSLi76kfDrzDnHcw8dV3c7ku0j5Z0aIlIJ
5+IXw6KncZeCiez07GxDQDOqNOvrE3lnFnWnY+KI17ULfAXIXQJikfGMMfft2Jj3y4g21XtS4B/G
Ep+6ivNPCsuVsT+g5+IjQpC401IF2oZvmcsMmATUPr9ws7fgO91myVkwZieY35tfenemU20JPC9x
ViCSd6ZEONazdWnCLXZ3W3TeyZttEzYrQ/bT48VPHmltYK/1/dMlwv2aeiE9pYpLj0HVdnncX9RN
p2wErF+lcirj3p8VpIF2fvnQxskpHwQDpxweJLO65h5/mnHKQhf2tlJk8FuVeQ0AUBnvheAQ7aqO
f1Fo1yIirv6ORYXMAccW6UZ361HO/aTe0rdvzkyCEKYwroafUuLpcSU/MqtG7EgkJm8jx71aFzJi
QpK60Rx7woWw/8IU2gnEjTWIcSK/Tcw025iLN78LK0U1BTFYviIhq7cb2BiHwYGH1Or05EBcSn5T
aO+oLnF27d2tqWBy87/rpFa9nFwNgjcZaOwlirlfHrH1kRwUG6jvxFmCEEXvz/5oM/Kcgfho8yWl
o1+JLVpWRGMFhDbiWOSZJDuv0jI0t+lR8fRUBs1K9pMo1rg0K4sga6IqX8CaxBACEU9pfGzmbi7u
9ptmiUPYFVOpxrfr7VbIJWxePmKGqWg0l4g1Htm8l8UUxBLQvfi1jQgn6SXcwgZ9AtHaunt1K/A8
Ys/WFo56of1qQ1gYBCeKdu0Fc/XobyffkLrAr2WjcO5WPDbB2YW7Z+FR5BUSr4GykbkRi6csQdws
GAe/ekISACOrnUwqdc43Yu4bld0TVTDCV/iVwgwXV/9RYNOKz2vzSsSAsogQYEvCYv22TmaVjufU
fxT+LZDoTnBTxut0tixhT+zIFgibG0uHcLIVMdtgrGpAn/A2SUX25sn+rNDGmUUPXBoLytDro+/j
C6lI9al+fnzrOOOoQE7F9XEFvo5XDSMVv/TKd2dRikuRQpEvQCXkEFYfEQz3BhQ1/k3+9RfpClzu
mA1IJoARN3zBhOJdQh/szUzTghZt1t6HaZEyKEY9HiQZ5RCmHYVHRlDnV8APn48fHgqUcCew8tBv
cxRIuuZkCzFvLxpX85hXi+Tx5cMaMYAXhUmLSLak5Cm9PtntJx2TCE+lu4F6GmI20HY/Kdow4g0Y
winchOZXzYnGkKI7xkhMVzqphDjjY+Czfv3Jvcagfrz8IacaIH3DHPX9BFoSye6dP4X+p+voZkw/
ee7FDWbH3ehnm837Xj7aydoSrfJzgz1P1NSOSheqWZzJpMBIWBqccf6gBbtESGSJv+o5L7FCejC6
1YaMivm4iaUDx63MIwiWnLfrk3ineIu76ANXw2tXYPJxLobGaooPPK9oXhjacxHpBbeXOQVPekAt
WgIz8LfeIBdyhmSrUmfHzvHXg0eCkjnETd+KHLWAN/PSZfmV7pfA0+uRQWY+BS74scdM2h6YwAfO
OOGviks1FMrcz/dtpuJ+oXbLFvOrP7++FiCcRPNYzkTeJBlGxSCa7Kml5pwLSlZdORW/lHqtYvZg
AodG2pQjG1fpwLUVrllTfsTrzPS32sudgnqzoX7khFgzUQQFKR3ktcYMbf+UgLt/ZG8HIgvmTRqK
+9kd5EqyljAEyqD0oO1xRUT34yWeg/5w/iJPgbNATFU4eoUO/E1h0f/CgcinbkAf6vmnuofdJkNv
mk3SMV4fOB5prttMOj8xIUB+mVdumpfJzpRR7aH9WpU4HtGhse1ENOV29KANYVe1pXhZeIH2xOgN
j+OCeXHhxIKyLeJjDhrCIb3tqU2EM1QGCT6aW2MLCeeNseSPQmKXVTjO2uMgU64jnjLXmAI/X8TV
OYhD6bnm5SQsDS3SI3h827JRyjAVqWwr+ovAq3N8Wt4tMZeEohVQO3TCgVK3OobmxG+9n5naWRC5
OAtScIf1esl3CRpSo/Ac8lqleDjm5qjljE0gmWVtFItqmhgA9aiiZMZrH5fTTVoPULcPVgdkWkLD
wt3Zf8pcW5l9id84Rjl5cO39I/XsYTvk4Htye8Hi2/NPBvklJJHYUpjCnez91W/mEf2cUx5uxm7p
MY2h5KrCK5Zf/LjkVNXDYvw8aUTwymdapmFnYjmUqTfS/ZoimNmyVt+6rk9LNd8sJW9v8j7h0XZH
pGiasAW1FEwxPlf16yJf8rU0QcrkcqUh5RMw6sOXyXfHc7rDNNqywJKFVYYwrIh+wbBb7izdr/aL
1T3Ct3Z219CLTWUDFaprkTxYDsJ6q1U+7K4g5nRgF7RWhxrWtByLtK85mCqVpYiLFWILsSdtq+pf
IQiVPD4EbN7k4XUiqjQnsOXyBOTYE28noaBuKT6KDQpA2kCljIDd/i09AzR5Bcu1LZcNPcZxGTOo
ICjgg2Ea1LUS5mODlQvvODz/BnWpSf31lBcMnTwnP6oFSACGGZN+KjoRejr7jDQFa2IAOMYO31Ov
z9NbuCAar6Vkt0eJELXoKFXuxpsn+Q4sTyT8YluJ4nUefKJhGnj9FkdWDcCQDTO0oOl17sRvQs/k
dX8lOCJiupwXnaR4in7dtBG5CEsVVdPaDm+bWoi/MdLF1ViVh1u8kz6gvbm77MeJN1LWRMPj5WBc
1SNpT5dtTROKFbWoOlQ9FQIViSH7ZeEGRxu4B9NRbsX6rvhkqe9ZfCZqLqvBzBBFx63WM9TdO4ik
hjQwmU/UGBKdwFMreFJMCaePlBZIWPBRJzJL1fklJNf2DceLLRneimFdXf4tKMQ3cwUC4jkT383V
lPAeNYlKRMDYJEkHq2uE4JyLoNwoGpRxmzsbZO99EO2q5Dr/rxAUbWQQOZVMKvwBILrSr6Y263k9
gHjgZ3JwmOkvKRs4VPwjPwSknj7MtOGg391rfZjZQFoYzEC6lp7aRl1Ms8w3lZmGsKOpsZA5EGfP
Vjx6wE6p0AHdK9kmfDnUAs4iOB9dCKze+vjBF1X9mCw+rYdUIbQ/MH2qQkEUiq3QXttBBYGQhPev
x8nBz9AJmzZdqt5bdaV64ppQ6XF57Xk8STigebCRjMeSb0NaXWDA6kaRYZZgcZoWo7UKZVgEeQHA
a7nwveP6e3Rslh1PcuFw+TU8eOz9EEBRoy1I0N8n/mJEvwUSLzK4YpaNLqYM8OKPSbeW74q8Llwi
C78tUIqiGYO1BxXUe5MGjAV15j1wJt1Y7Eykx3dmvW4FFClej93UeLw5Zs71XTluToISmHiyxZ2p
ngayFHt0+/po5rapc1gDbFM3SVa4edYO4ox5YK19aDPry87sZskDoLUtUU7TUXCqeJLYs89jA25f
8o1hRT2w9etnaGj9j+/T2sJUbd0K6X9PLQNP9s9OwnAaW/8OfPZ3oITFFv2C8keLQ0t5xvQEybr8
kDXRsZVzCqjcstllree1XBMJOutmYXqo0/4sh3kWnNs3gr7KNzzHFEneibjkym9//POITE7P/JqQ
F50kgyCvKxsOcS3wAWM1F/NMQiO27joakLSaqIqfzK1rl3kssB6ETbByrKsJkImNrtLXumR+yA6b
O6QacbNkrrgXaG9Pllx8pZ7vMydB4JvUMw72PXhNHOsgsWuyFAWEzdfvP7PdOCs+ft22sTwkFF80
1D+E5qYxrD18Eq+AEzDnIVLid2knY4Ty79swGsSKRuFMUJAFvH21brQALGeldymgoSM+B38Dddr6
2lIOEImQpeMjeo/Q6IRPjXbJxZWLjlPlJKW22q/rN9jRVmuSIH5I9+l8VTy+4efcTIJytvb4tAD7
6qnwTW/NqGYoHzszwEwTtNKfPzOf/pH4FxGsvoOeD0fXS7xyrz4NgS732WeAjkMo5uZmeg0F0QTs
PObNARsPRNrWZug2Hq5eFsHn+Jw8xxNx0j01V5IKqH5VTjzI8nvEt5ozpKvkkbHA3m8pv3jsGt29
ktz76hKnKrPqAf7VrlqDELEabunGhmupZLQ21zSMg7uEUYaYsARxWOUlAdmPNoFKpy0jRGz4IZaM
gFlikHYZOHwjo5DIpa+rF7Jq0GFppLvWhpLmg9mnbDojw+yPgrEX7QQSxQsKuZfiKRagzarkWEzT
4JtWRZll3UDMTiMDOeNKVxrwBek5xZtML9HwWTRIjguhxpUXQK4b1X6E56eXI09SqwLatHZWrrx1
86Mskv4J0yOThL/7PBkB+25minVJDHF7LHkJklEYfQl7KU0CkUAWjzkwD5ucbDTVyrV19GlXjJPi
jyKSrgX/V45g19b5rzj15sMaWtZz9a1J14BW7SsW1pu/ti7optf0HKyj96UP5a+tvTIMJslR5C4w
umS/u3B2uoZVobA9y+toLil8bOyVEgM1KQZSNXT60ggz+z5ws35+Qq+i3Ru6C+ccQ0niKce9WsNN
cZHoNdcw88ZIoEbdFh9UzoQVjpc5At+2dUkoaiRf6ZJoNK/zzDfJxOi3G1BEKAIwvovb2xg5wZSy
A3WtcnWCw8Enp+eJ3uZMehIhJtlFuP+kbMGHKBdU84ki3gdLM2Lvrq6vsXt1Wm12XWsDjShnboLq
UWO86he4B2KGzIvy0+Kgdmf+Je//zzzpuhtwFtrZ3qrBbZWri4WnoTsnHBlh8cKHN9EPys93raEH
KTz5PMoAhm2mbqKb9Z+iou0DJbMDsCc2SWmM4J/3z+C0bIAVwSIWGQU29HHHHn1KLdK/AK4NdBHk
/z1q/rFutHl/UJotp9bxIu1LjaAlDWlqzFIb+kxJqzE1NeqsCpCtCU67C7KSmhD+OdvPFuNqeI7c
fISe7GjDCgon/K1yQzjAeOdG+S0a3mM2ilpEJcp6ecPAVwWeHYfClH3DrVZZxxKOMYNfW0B9SM/A
hg5ByVhpIvH0Fm1r3tHP/vWWNFgLR7Pd/JfEXnxiPQ5up7X1GdgKcQL9Z6Pq5J8szCS6vQDVoxA9
S8qSCVx1o5aVDV464uSOTeKXQG3pELM4jHNITimgOYG233/3e//H03U5ATb6/f/hUvkxb4UkMupj
Lznxl+28YZUGg29KCqQzANV8azXtbvonEVq1DCpO1z+dlhm7udObeWl5vH9pd7D79JiPDC4I5f0W
G6ws+y1FDhAQA88uDdnLA/3lBRCj2fLf5NAZmM14RELMDx9GaTnZ3WJIrAUbcb2zx4ImQvJ7bRth
+apP+uidlOEG47yrC29htXfW5VRekqcVbenO5aKeybdEZg5vb0YTpDTsL7PJMq+PEBzIAgGLR00v
hIrsh18/N31VSF1LqqnfMoTo2afCAaau4S6CMHg8fp2y7KHZ4U+ECWyDj6ntkpnk3LkgK22bpWwt
aLfPPzWFbgDg0JIK7hDF0Exmwhk8mzFx2Zs9mTERUexgMDflrYGnwVSZYI7yB2ComOR4Qor8nNaf
OVCvPHSPicgIB6GMVryQYgmhmOjdemI20vYUSMH1+ugON+gXTz2ASxTlh+13VgQLw1ADmHFESaLd
+6tZgb7dH5PqrQQE+jqfDS4j8laa+zjaaqnPZZFFYuQKz6dcU3AsAHud3in7bvvaqhdRDNXvWMrQ
eRq0+nMbiv4hWzLWJOge+Vq4NBXU9ghaVJcIZ/+wrZM6UC/FV7fJn5Rm47sNT8nWkLBkp2x4nE+j
roRo4Wqyn9kZaUgxwFpqJBeFNOd3vWqi0I7XAAg9avncRC90irrEbTeqEfD8hpslpFVHH8INM/pO
sIS9snwW/Q7kdqYbff5aUKalwRzkXip97JR8oXIpXHNUHQ+MCsqjx4NQWaI7QzNzPYxv1fGLRa/T
4HI/91I0Xh2qpwlDIBSec23wgtE14pdirxhyBrENzsv2LLfKEXddtS0xsdIQ571S22bCKeMdK+rV
22PM4F1zovidX7cjfEwhrY3nni/QIPfy/1hivmY8vz3ZASK0DRAid3yxTaxN9JzhlIPYX9hh1mDH
sHWZSfyoAZIXbbwkTmhjE3EN4Krz/YIv1+PEmwIZCJfkYqlHZZrgYQJ1yzCBrbMucG3yk66xr8NY
mCMcnY2VNYKoJlxr2SwZFUEL0gKBAeeip60NLN6v4R/ygqgv9JFrHq+4V5JIyz/RpNWXsbFahcyd
Wm3ZBiMSyj4qm+603SC+MBeh8RVdHaZtf/yi+SuKxeYfdxkqdizyGHo8MvFwMo52I2wYJH/VbNqY
obSBwiTfcZi9AU2MI0cfQg10xIxaWEo7GxypXJODfipKTWCw63K7mpS14ArUp32rrHjfGWDDQjtS
z4DqRlS7Bh4HD9DdMIIN1PO/CgX2j93k26VqfIALZWFntv0SZAjIlAZcQLCTZKhnNNiLFkllX4A2
p/+WPo9C0K5eKWR7/tkSwJ5E/Fqvj74aa5Ek/3YwSlPuP/cBLk274JAKib71ssaf6Unfs8i8Kr6M
q4VGG1WJPlaQGrT4glb/taYGBkToYtwrcGCHa2sWtI5qDiL5qAShZp1uTbtTr8Hzpn4uFQ6WsaES
nhn4kfJCwxe+p7FSmUqjQk/62AYeQN3LNOiIWAh2s5quIWVGyyyAZZPoorvhSmnhyLn722S+DDAx
YCtcHxTlWtRynYvQa8IQ1gNkJA6Ai+yY/3emS3ZQNl8IGLwy3WGwKbDqdvg1oyfy2lzAfu8y0kJr
B4Ogch+FC1Nn01zEZZanAkzsVza8rDu+prdMi9wywqOJ79aztxY5qjFKhGrK5Id9kXnGPnKSEKTx
TMoEtq3NVtO9FXCbKoaJdM9w2GGTXQAos64MsM+1WhPKT+un8jJqyBxGlltn+8NWveB2hFlmnD2V
PUZ46faTrApD5btr3Qp60Pqt9DYXuEPT/qF4idvJMidclnfJqXzpgj/deVRcbWDueSkRTzlzIOEh
j+ncffu5V0t4QQI9NqQcUEk6s7amuD31jKILxVh+RV1U2WV0SI8eoe/mL/MYmll+IPKKqmZvRTQn
dIf+WdLf0rMRpOEv1QP3Qai8wXtRiBzOWaPWy3j+cY3zyKjQ/Jtd/mkVl95Q0YYK3ZbGU9zAFgdd
6SsrRzQJzsWFdu4O3/61TPWjr72KvS3iByKpko2d7qg63e1/VZthK6MuyN2SBFbqKAsjZSrloaVx
Dt9ems/OpdZSj93gWqk6QqCdCpxeLkdePpgVZqKaQbMyz45yfHFRvBqk4DwLU91DGKp6slsweEEo
By5H12gXmqru6foFfCclMsg38aOgy6vT8RmbjBOvKFJ1pMazxFpa8qOJf0S928BOn1xFyyjRJi5z
YC7P+/hpHV/51ztt20M5Fv2y+meuhqk+e3t6XOSlxajUpk0d1cexOACKZ4qoFTlstT02YK4HQhwn
MpVHuKG2z7Rnp4oocMvjlv88ZoAdBRdS8gvmhKzushQJH5xDoVBFIMPa5x0eK6w7N0gdwarUI0h4
TsBGMWgTkIzTyUWk3M4m3pP7KUq08cRtfHJK4UEZmJA2F1M7lIS+cRXqPPNnM/7piLFPQWkZ/fiG
yremr0zSu2Gm3GmuFUUQ4rUrcq/NZacFVbUBVNRR0YcTF0dli/63JoAN1ecpQYbGgUjTCAqExi6E
3LFdY/vymy6d3lgEPho4BM7ozOeuVxBYKZkUNWfM1eVHb3ur1DHerV/URfWyxpIW3ZuuVzM0hujC
ySBNeVh9grnkcTx1pE6jopvMPRZVnqpLyKDZ4Yx5S4y6APeQlB6FJ4eFp9MCR1I+QymSt1ICONyQ
t8w6C9uHdcqlXDVsJWmwyEB7JnQTkGOX0NSZ6EwoZBNQ20jIs+5MLTHprYAdnLewdfkZwPSDba0D
7UHrJXO0yRLUxW4GZTYbshUmpxUJH5eBEhbd4llatnDzaX7FDEmQk/8dcleX/FKzqgFAcRWMFdIR
1wgFYLH2XYvLLzaYkVOZm8OrD0z5DQA2SOPAf80N4jQIW6+i/NDxc9B+beCyl3k+3b5brFIDPAQP
naROVbZHy4HM+syWdngSFBJK9IPsSW3hxvKpP04heHeF3XnX1XXCT+cqPZC3onAcBr4psJZFWxP7
KcSCE1s43YX99bnsRE1s9K5n8iBk5EOQipnRU7WmYS81ep1ulSCHvGmhqNJnOfmFcYimiZs1X1eK
NOrhD+B7NNcVLGgq2bd6km+LYmkwN7ZShemazMGjt8DVbR6rj7kdAQHjU7WcR/WsvaBQjm0mIXZu
iyUrnRYM655p2/nV5+S6wfRk27bid/oUMxiHBSj/DcCoEzckfAn01aysfFGERERkdzaZAb1MGYOP
TcxMqvtkJVlfTy0B/YoAdPsx7TNSh0ijLGUExpgFN7JxF3lP4CU2Oi2ENzXSKcasUgoPKG2v1bWP
ReawcvA6mZGsD9Yq7I0VyRpS5o1sF+5Vjvzt0SSF9Ek4iWtmec79puC6/cL0EWb0Sbl6ha2KXxn4
MzRNyYYQfRgx00KPOsU0BWINXnB79R1ei422KCtfIeOHdbFF+Kz9kMtRsED+sxrgahXW4+znQpTw
tNuBko8izEn+ObDe5XzJ16ltpxYZbpUXXd7clb98i4gvBGQ5dYN6KOE58stamH0ybxOhVQXHe4s9
lju2w5HJtnxj1pLlurtkxzki1MzlinUvAFnn92PA9+DFefDlB2wh/XY0mwEs8TjKykmeaNLGv5p+
u9LyuYmCP8NjUARKEriLnlK0LxlpMGiNe/W6cfyDBQGI95TClxFTpxMpUBgv+Zw851dc2EidMZZD
5XplMADp84higLErE+KoE7oU0BsUhda511tF5iI6wCcNnE+n4OVlyKgdHH+zodP5vBCHU2n248OP
A+FrkTlIKDIJf7FY3cI7dJ4QddcIN3QrBbEsU+ry9exDrSZNqYDULF2SEVlsZLCsAvXoLiArjDZi
Vi1gO2Df1mqm4P9Xq7yylyYdex0YXo7Btc8wk5A8ZMPRJ+3DEHbB0ezwdVbvVoOKJQt0IUr5tfrU
yeBn/9nNNh/KIQ113B4nweMWzIXeYi9BGNucUZ2zylGAXKPcia8E84ulqlQidqy5S7p4rK+LZwd9
VaJrcj3iwLr337RxV9JKx+pNKfMhZzmqs8rBZjPzHP4o+J+WvKKRVvoBHO8D0WoFtJgrYSCyCH6l
HVcw3aMUTQ9YZtdypm9oDrogKOFimn054AfwnHpUyA6JWN7AuL61htMSBdj9iRVRNB9IwgsjOY8B
tkLtTz83FO+Y52g0riyhfTzvRZNjyie/kqaYMzdnMUrX9oe2/9QkSIfac26GrUFb23/8xzs5eqo1
0JisYjQy0RLcFDQ7UNS5Wv1xWcLIkPmQJQUHIss4WYmsPyUuXr4PR8BUmFpmAdhPSqsFL0p4Kjoz
PHx6ZftgDMRXd1tcvw7efRz32PWfCzma+qx7Sl2gWn66S5HyeRwS8PUBHddR9HTLHNF09ZBlhTB2
Hi57I7pA2I25vo4kaV18dpbk6GPhHPh9lfM46Sxtp8UR92eqQD5AWW4AjBTkUkAXPlJM4N2f/Xnl
eHn13lGXkETB+XBc3NcZzLJ/ycVicmAto+KzIUIFHitxCUqoFC0aRtNminuCwFlFsu8G2EQbPpge
BYdeCGtFPkyB3OY/ZLbILbrGFJxBasSJboBILk0HevmLm0JahjN6pahHSWJmnFBC6WeNhOWdQw2t
rXBQa0cRitTWnuZ0xYtGOEfZKrGu18L6Mz7C1WSkxHDqh0tIRp02UqB6k31Ft5Nhp/KmUqcRKa6k
vQ0MGG18MnkHco+o8mnvHCNbtTYb5eFKBEmBGHvhcnYGN5MYUdO0nr5flbjjrfYfLF0AC1t5aXqV
twNRrkTBN+dIpRORnz+7QNcxjJMJiYSF4cFpiT+kaIcz5UiGHJtpnwEkiT9Xr/PMFrIaHNk0rO8S
HGbpPliUTXbMEm+yZpf+e7JnUJiksaTJAsdj2gzPVpOT7WwV+ZwI9Lixzpy1Ua4CHVh4i41hTexb
j3ylkZ1IgUFk4N4X2VD/QtcRN02lq4INo/WMlINSA//ZVG71SuRZ7uhp2igASxlPy/AKKpMJeQhu
9QG4shMy8vIF99Pouk5EqbNjsFmt6xZ4eTy9v9F49Q1A1r6+BTkqqsK9dsJFs0DNnn/RqpiOz0ku
qHLolly6ogLxtM/DeM53Gfjo75gejOGdOHEx7OntN7IdI3+1nzaLGYL8U2bvzzp0pjldg46U8Lfn
k6G2xRCqJV+1Kp0FpRaCOHGflRucrsrfzqv3K7FidT5e3HnacwwIYhCbWzGbyG3NyZt4HGYKXia2
LuisoFqAwIp0ha/9ik+ou4QVx3xUWfxis19hXz11h/uGZAy1hgoTy7nvaFL3OYHOT4x051n26s+v
Kg58DzqY4li5ZYc9yfaVWXRT5IcsUM6fNo7+7/yym/TDrRKZOaKAIcpoASc/ni3oL7kw+KK5UtdN
2GEmO8ZeMjDe1/IoXjjdLQbFU56N/6bwMtzg56w+4ZezJGsSjLbV2YoIHg5eO7RGBoBgjRkgKbdT
A/iktC0slB7dG5xtPJwpP/WsuAMm+dLrOPSGN7CHHfUPGB3qynbCvpWktLP+w/ERgWvH9JazdpPn
r0FLqqHhLE2bhXTXWd4O5Ra/buKQiTJrp7UmT3uqa+OwiZqqHqD4qd0gw83NHYJzGmkaMAiCKDga
5QhPU10on6wQl5hzhYKezU+8QjF8+eJ73w2aB4XAwoO61DEzKUF7LR2fDHMFeXPX/bvXlnHvw+jH
grWrm+tDDBTGxH9A7PxGTWw4MUxSbyypawe5r7zTFv/LCd0E0RiR7aeZuYAE5EPe4VHPaRcNt4Ma
2OQw7JkhlAkSC1RmlqZr7SlQfgudYupDYoQQVCNQCY4KxEKTWyk8DZCZi92qJ2FloYHg8CFFqon4
6azkXK4BzlbhTx6HhbX44G8NkTySkUnmZVAqwyupcnTRZZQCLY+ydITyu6WHEuOiZe/gPJ8i+NUZ
SFdD4LMoj9EWuEMQnVymkoNgUJ+wbfDct9QvsIU9FjpTRzDzDkiS7P8Wir0tc9+houMWQR03XzEo
DshchXywB9wX1jO8Wwaww39wJTewZaDROkv5kmXOfJ/JpmCibyM0rzr0u62ghr3n/BO+Z4TZxo0b
xXN1D05gfWLf9xjsEwEBblb0VK/tnyHw70gNmYgnGkummOYbeWjUOWKbjlZpDs7tXDfQlzMdK5cA
G0bydBm6MxgnuVVwJGlSvTS83nyMUblvISb/8KDW+sZCtT3a2W+AgbPEzcQJX9xHXwOsjm7cV+aG
vwonSOfyUKwmIBHv99sThawJ7njnLA+TtaUEjZBTiiOB5AgEQ1TXttuBMXdw5zpG90QkXYsBOhpJ
ILbsT9rJTcoxjSt/TYE8RwSnA1bzS2xAj5Dt4psOU/J8EBknfz4PnEgw1fpy9SK2yv+Kw+HwuI8e
u431PRtT6GYp34GYNwGw7Dmvzhsx5Xdn0HNG6S8fjgJyafre4w5iaeFi0WwiqiijQITTcrUG8l3V
9uU/r6W0jq+fNGnuXrV1pRTzTgcufOwPKAw4/VNc/JQMoaLcKGJcU/YvJidHUg2euVyIdSA7o6jP
EyaZnbSJMcHgA/DGeojvlb93Hs4+vNbYHgDjrSqYpQbhKJ1oQQA8FIJ9MeyKZrElvjCXtAeyBbtX
fveIbAVap5djgx9CqU44CZS2r+m5mtQGML4+o5Qtai72+NTP+K1QpVxxZAg8qetWZZOOM1mMUqqa
Ts4ytfP6Fc/U4AXKv3ovL8gqQMfq5ih2kGw1jJ8Fs0Tl0IvMLSuzaXFatnWM/AbTyCRP5mBDeLpV
urn3RTcC6HfQLClY+zvR3HueNzntB759OUcRkEf72q4ZCifDB4avRklDu9t1sxJdnPrZWl14nUsJ
gylO79oqqS7yqFBpOElNkUxjHMnjuFHbFx84MlocG7FdKfMTyl7goXwTfE4CfGc9j5fMzRraogcj
9QrRMwSt6L6liTnkOWfuSpqYmPBiv8I8XZg9/hQcYqnsG9rwqXLPo6FUV6OYRgPern12/0yQouJN
Qumu8BK+0cwQzYxwfc6d7UtDEkdDbJ7c04oE2MibWG9A18liisRZhmCwuFj6VQYPwHP57vMf/af+
IPQl6ZKUBu2qbFBbuW1DHHkfrCrbVA68fweICYPiNL+qrEAZIVUsW88WE35hS+kFFQK7x3tgTr4s
P38OlLAAmhB7v1UinndCXNnPvLiH7Ih4dTGdyMXLv6hDcmyC+GsUyZjiAqqSiTMjM3vmKj1je2gU
UITQuuY97WaYvVfgrtUwauAJVFXT111a3sLWkDlAS3y7yTaYK40jw9gI6qpAxD2lFBtzNze0glNs
7q+sN5g8LsadveYmd20as9BlbOXY8QKaPQh9PpQM3hz6AYIsBJGLgqY3phI6Pm/eWpVhzSg6BZLs
9NLxf4d3sOoEgGFSC3ZTcxNTvt0XifG35H7IcOMz3CRsMRn1gFNf6Ln2xLbLl5kOIKcEfipfQuXt
Zj5EAQ2Jd7JJjXbs5iYu7VPQPoQAwkX0/M4leuIGqzdStEQ398xFOGfiCPulKYhX5iq55Ly2LqDG
A59IJmT2axnqfelCYV7pONNSRTfQXC0eSJetTsdOT9uwmk/UeujiqO/fOFE4hPC1u8rUlgLm8xlR
m8leBcqWCYe8QtwftZhYksUipFKirARJisPBcVVEvIqdgibrLbhfZCoL5ImX4VFFERUkJtHo7fjZ
W3cuATxrbut2vl4tjBNPP7htqPOrwnMPx4mQuiNUeewbWy3G0IZycjzhO6TtTm1YpIqi5yNtFqRG
nP1VcHo76r4yXRQXq3NbDIdcDr0vhuv/BlL7bL4PZHD4nNoSJ90yCf3F0TO3PLVJr2uL/Ux2QMO8
rPJlRosSYSXQ3DR0wKVqBhzh7gtFOJIpajv3RXON3L9cgp4a70Ig8Eh86RWdJUMhP+HgX6swupSt
HNrGbhR7rsIxLeuMQP5hQNkXCC0k6Ypnf843Wxy7cuvDu+85lgWZRJcBsjCkSuFE5Rk0I09/+Elz
GujCEQ6wfziQ3eNKIST+c/UIS5gfGPGZRCnHv717AXsWrk1EMYhfVpvk4kiZcEYbL6uc5IvjtLjJ
bQ8Rjdc/WNGqkHDdfUC6MnSKCcEdXL7aysTmpCxmRhEUpGRTflVt6dyrqifSDUeCo+ryJ1uDVxZA
WZhGL9wxooD9xqmRGcsb8tqgqZhwhI1JImV6SDAvJPIAyjPZayUAT/b2K/UK1Jt4a2O+8BMlN/D/
1bznbLDGKnu5uPa1IF74pZSAmHBXNv5TdBIyOZM1Qd02mAxnCrxwrT/N+/PBzG0sk59kirG1Ykud
9K6CdF187C7QeuaF0NFdSCKVBCoI6MaOcHKqpTssxxqBvCGgCzZ+SscMMT5Rmx3bBusTDGdUw0ZN
oM+gwqYYUhIlRL0MFM/SE1VdzGCUSrNZVR3mR6fb7EzpG6MJJ/4oLUJVsT/Zh4Z3wMO2JnWDpfDB
ho2Is4j5O9Q4r2J7gaOaZYxKmBkNintufFccsWNeTDWA6ViJGCfs7+6NlqGVjnY6vNIww1HfNqoJ
4plN8g6eEDK2cHL+lPxZjnlJT/9ni4phe7Yk83Ehjz7lhDYrvs6j/8Di0cxsbPuc0F8KT/TUsh2/
94Z2Xu4f0Uwkso2IF7j7oV0sYefuk6MolzgbAJxsSMtTNJrfY0SfAi94060+ca196VTXTh4k0cPb
kMxKm7ANbf7ii0Qrw92LOuqmhu5i8FAds9CG8Uk7mGklgRKDK9h6KmLCNpXI9nUqChTjvQ2eaiue
BrUyzy8Atw0cts7iEh8pNodLpoaRFEHcJmpsHZlfj8nwkIzGuyFBnHWgHkZFNY6UadX/67QhvW6t
SI+Fk+vYl++aCK/igIATlo0yEzWDg7He8Lw4SpzouQWYC+/wawJwVnKOBdNxCIUX/zIqtMd3ztHq
RVNFlBH4LB6UnzipD3dC0MNV+wj5veARMEiXRDepyF7UM4Nnx1zXaaCCPKEr48GlwAu+API4QErd
DUufHZ0/B+XlkhziYIYD2GQKIqLGVwOep0UfX6vp5XRTCz1LnUzlMaYvzhe1QPv0V+rwPz9XASzM
E5+JBuOn7MTqorWvwiMe5LQrXDxh3vrgFKBqy+IF7UYGsMUVjuxo3OLUS9/tXApHDPjmFxDDjram
9K9cka9E7CNKICJYNAMTTu+yI1aysDWgPuL6EsUKzvpK80uhzAg6Am/InGcV0bhQ+8YPFT5gZOmB
B6qHtVbNUr8Mwv+jjDWBtmCH3xPIOHBVgaIa0XPZUW2CwfDHXlDw0J4N1Wt+oxG5DZ5NTFBTYiO9
mX2zboIgtXu+C7Y/jTCXnEObYziUyxtFadVs/8K42ZCSb3JLgL7M8rSfw7wPIOXpW5yb8O8fXrBw
0vhfEEU/AjSZixYbUvlSwlFRy8AKpXZ4uQwUQNcB7YoCQqCCgHV5woTwGZNhvqxKJSnY/KWw5hKU
xHHZcFTS/FDi3Nt+rTDlmkshEWqJmgVCmV8QL04V6YTL2aTGeVP317EEFHt8mQ4k1mfPQSToZJAv
huXnXSKM/OVk3fsUYEWLSeRvgKA4ma/oI9ldAZQmrloRUex0+ezrRCt61FInk3HbVnt0UOSA+NPX
bAkiC1MyKSmiZaaQJOpf8rKQC4BuvIk0cMw4ZObmyKVj7GAhiSXUp//9MZkGW9DrEs935qQFewfn
/5uP6mE5Wz6IUcR9ZJp4pbPpuoXRecYtDb6g9AwEaVBvJ2Z4NH0KzsnT99gKOfq3+Q9ni+NOfmyd
Bipgv2PXb+gppSji9z4Lv5FnCPyq8BVBFK4Oh3+flbc1HgnRxUzsoCdFvOBYcG6neLorwGoVweq+
UHN3mPbc6FACbS624yb9hYZ0sRwhwxnL/qm3BNgNE7jCX1Ru2wJU6XhMMbsS/8PSPXkKk5wvjWgN
zC/DJBPrOdwFlLWbZGRlbcvLvdPTJtsgl9BDBNjOGWOtu/3q3f4XEzDQwl5BEMOLe6ojzGpQOoYD
ccQs1/DgfhnIvPLxLjSHRyc5Ru2XejnBMAu1eeipAcV/dtJ7IcZkfJqqGpg1zKf0SfxRP10h9bid
gj1nrdsxGiXZ0BVyTLnJfXA8nsNcsX1J90OYPcJt/DcJSm0FcSspB20f1W3gjMsszv+L0fS/9TYr
/XkWjlnY9gaI5wx6akZrxNDHsAh7+ITupIHiR5uSXnx4X2ntfmvQntMp4MfxiKQVUtgX9PACm5oC
6RF/tn8ba8LckhmNGgfQ+iyS4GB5UdTnuSOJyHSUgxLz4n/md7gPISavAXZixFZ0A3wMhnrceB7k
y3Woss7N7ydeNf9NRKMF0lGo9RmNeSLn7oRBRLbuZCV//pFBRsqAI04lk8f98ZNqYmFpvgo+nhxH
tl8ZaSDy1EpC1AaiHpuxiTjSHmJBmuTI7rYS0FVaY5F71bNqwVxdvjv86sIZqiH8MCH5wnTvgfNf
q8Yl6x0ndErLRMvh6QC3CKe4L1x0drd99dhq7fCMFl3qLEHsygMqsweMOaJcOB2RbE56P/yCGqOM
kIV34G40+o9ALPzggwr/gbv+X5SSXGp+CXDywKvzZRovpyGT6ULoW0Iqm0HQRY8/nf+kkTQMMY3b
L7wE6y5OFIfzXbBaRi7gqGHOKjbkJsFF6E+xj8d9WqOPiA3S6EC7Ou/floJRsCiT6h2hpY3ChcfA
Oa/rnT+FrSGmVy8cnU72xPlZya9gP6+UhbwNZs2mgtwUMaPFz3ddw7qDQTT93Eda9+/8Ymeei9tx
UH+043sZKe+4T3iaPaUReoI+7G3dNC57ZDZVq9xXjk7nHST9WQZV8P5BKXs9u/meZRFxco74BhpO
uXkVKjScSEN0ycJC58GsK5p9HEbCSM7ciNnQgi+SzjcaIrQqP8y9LQUHWWcyhzl1Qo+x9mC/Fqle
g18JTk0KO4lIxKpVXLQ4DaCfFHSjcVJ54x+DcYIfkMQ+eJeYHpQRpJdtf+OP8DObnPze1517xTq3
Xj7JRBkLKGES5zubNh7AQibXqMdtKBPcden1t5vnX/31FOxJPSZPL9iXpUtlXZs508zz+J0Gt2n4
poLGcU7+VaEvqSfo9jLYb6mDozkHWhtYzK/p7e8CoV3w9JCsCsM2zda3WSZz5ilj0UhHfqUR06mm
gECoUr5L8B4fcrS9E1vYW7i4jR+4iElpF95DxoS8d3l2u6+eTsQkMIBD6+MkGtTAVDsLCtlO3rBa
jYCZTymeksZ/ibWeCVsy31Hmnc6pBUJxtX9jM8Xx7Grer6QtmdpdJOTqWTxob6f/nQSHZZtT9bQe
fMWAoOjbkEZN7oCmpBdiX0ObUig/ORV+mSk0maxv5l99FhYTb+EZcN9jpo+lmjSLngA7ruSiJ0x1
ngWDU1H86/rj3/0Slxsh3uYzDkwLTuRJJIRANPG8BV15OwfJ9tZzB0DisEXtSabR41LR3jK+qNEz
AwFMmbqQkI1cjEOxrp9IaUhF45ww+gfKKSfBgwWZmn/OP8sNRM/Q0Batx06fRK89lrv2Z/S8++U5
YqNFTKp+yEN6tmJr5PH0YGBeXIeVSiw7Z0k/q6zZFXZOeJ1CGECMcImkGWOy7/08Y9UAM47O+kc/
Sxvt1WgClCUJ/8DBZBZLPBKUs5luKeBBYQbuhHePcHB35SqUIR9c3SG2j/oSUiKF6mES8CAa/MXK
7EUaq3DlAzk9Se9+OQbrWJt8QFzS0LaFRJPhn46BpPxi09KOh4DDBBwATMmOtWXKmkWepNQO0vVu
wuAP59jLhVnZm6q3XDFADthjuX76w92YVQovrgU+KGfwTuQ/fS2zvqEnIoiG2jNbtNdoMTruCKeQ
B/EUFPGCo4255ZRfA6e58rfuRUyRZOt6WPIszEZ+CIotYv2OICjB0OwOaEmjwTqqHIyWWzsS+Y+K
Ieow5JQYLPJ/VmrsZ83Ea6i87VP4IlAlhqz65R7nmBRtmgXgOz5SLTr3MK6WuR5sRTzeCMvRzIgg
mDpyDEmjk86H9uk9k24+bA5/jqsxUeFNTUcSfs2VLeIrBWKn0R/hf8NDmvN06apk1igDgXh4GWG5
PYXmNZggtwn05JRyZshU5n7fMXKM7qtxmtw2TXGDn3AWe7NVzWImqNFTpydi980+titMCEdcRCR7
c8UOkWpPbqCWfVJ2GysRDutoxG5dFPHphnNiE+j+L6J/7e3bqD8ouFjL7HTStqWPgG/oWruA6XlN
QxJKGeZeQzZ8+sPwjkqNFsWOwlybnlMd2sh6h8Ai/TT+a2oqo2Q12sOK1WvC3lpIdVCUGvTx5njk
dll2pKvhkScV7VfscyLyreKMzlwcUovB2vQpS/M8DUtaNY3U05lWJxmMpwxDnxs6sl4o06YpRJr7
IHLUicAk2OkQjnRQRRDTF4jge/vCT23Mu05Vt3IbIi9oLLhWBqCo5itR528AAHvXyzrYJeU8v3/O
UhvmWXXRRmUxFhlTWpj4NKza7D6cAPjNR6Gafof0EGJKsd21z0nIlxh2zx+VyLyKLhcuQU41FFTh
AzLoh1CWk0tjv/qabNLf9QLxEJmrcR0EOINBRfN3WlxtdMtpTuoLqTR/01Kajo0wIpgqQqjxjtx7
uMIPZ933AoFigFYcZ3TeEF0kUeBBJvfljgf8zK+fOxhGom8ZAFCeWi+aaOk3A5dDJ91jFAIAaPlc
yCJM8mhc1bEGgH1UXQVEU1smf90YHitl/aXLdBG1Lq+76A/d6Z4tLR8faURa+uiryiY3XAHZAPv/
yzp0a/YLrj6SzqPAtC2llufs3y5Rn5J7uSVx7Api1OuEFLMESJRY2m+3LwAU7SWSfX9gAh7FAXYo
lKpWQIX2BrgBC+ecCTey58DejLvyLzsV2875MYOX62X9sx5rmmN5vH2zbmGILhWfE3TVDUIYKA8T
WvV7E6jkC9sbWWQPlMkp9lwZdP+vwzOgjX+3KraiJuvZpZ8iMd3SdltkdI3Z04/vY3hsWMfcfo/X
izDmnqFskNIOjSXsDSDcbaVmArNnGob9qfzZn9o3NO/IdAvk9DLSOwlkQDaeurtNS6YF5G6lvOdR
pNVfCpjneyNUuntMWqmdCzNRnSuTWduxQnJD1opaPv/2xGUez7IAJatdzZF6OB6sG/sZyk2Rv0jC
yvhesohAS4WCt4lxOLmpxmxJzxIc5LdMQ1l3S/QIwEwMpnLV1w+JOQBpCibEsah9dcX13rbRZSpS
JkYyUDTs0z3QCRTvOyNI+Wit9X/qlsYvoBjCje84QDSdrJP2xnKrz7QD2uByRb9scn1uND6ApxDb
Ot5Xm3EAnjG/CnkeviCfhk9SSmL9yMyP7ZIyl/2MfAaYgO5A7JWDaMLI7zEK4zToYRaSBCF5pSMf
8Zw5N+3IeHdzqexyITu2duKkesk1HZ034mVAlqhQaRXX6wAQvEpo1I/08keH7f9XhtLVnZQUL+m4
6/CRQlyB+sC/SxvyHKCRQ6uPU5R1uBCPRmE6KNOfmY6abIO3c5v4dIITzVYcSmbQ4EHlfwtDTHhK
i4cVBpp5iXj1rZu6Lneh7S7hHKJGavBJQZA9WldOTZSvhce9G6JnBSKPi/eYqDnIOXAXfrIGmd65
q4nrxoO1bLlUKdYXTlOl5Hsgc+JGzUL2pWUQCsrh6UvgRtJxjmclLPrYOQzfAU5usDpEW4THKcsI
FAhdisux/ohOpNAxU4FYpU+dlWS2+M10xLaIW8rEN039v2MJWDpH8aRDEuDCMgPsgshZmOgj99kw
N4LhfcMo75lYhe4jgDFFiDMD3+vtgT7KXUXDizp1iM1A8GurEOLWZSqTDC5h0IaeSwu9tu5EsRjK
XBFexnIRd4/8aW485qiZDAYy3PP+4GupX1AwMPJXnxIqnqJ+BhPxImcJH/kifRPFlzlMNYtWEWzx
O7T5woKbzM+PyG5HLjLsAA6qGExmEQ8I2R+l/7pcbMvuEVdukX13MtrvCENO9V1LoB1rM/FI+2ru
PEDbywdvef+1pR5OKrKwGbRVltbkBtcsJ8uMgvuFB/Ye5awxTHT4fveoA7hs36FN0yZCS245Ara9
V+L1JVyMmMb9QKwvh1liQYxYmL8VXvn+ZBYgVEIkn5Df5QroVo9Pz6qFQvFVvTxa45LQvonKYHI+
21b0x5sOrkwa7apg+88BpgyUVmlAbpcktIYmtXCb599HDluWVgIaTmfQ18hz1r78CvW487htlAx1
VMrEOhD/pzx6yoThHUWCjQdRKXURYIcNOq9M0P5WDNCLqWXeEpjSbe1f5qnFrUSmjGbM8aaVOGMI
ujM6B7AaVQ77izineaHHOPtV2Rt+nAZejh0KrEimnYY95qm8zDKU170sVk7r2o/D6hYeRnTzSeee
Y+f+LIFPbMo/vLJnawHTH7rqZmKnmbnF3RPg1udZ6SMaTl7QL7G09TJ10rvQc6Ct7S27grtU3vGg
jy3y7jJFjvy/6ATLbRvElsI+lE4W8mzskSv0zNMHxZO45Ccg9RennLp8C6lX2qjI7IHwVE/+370E
CdmAZJCjrgHzFyW7328qrx+evbBwuNk0xoukrUrOrJg61QYssCM9S8TvhNCkGKa7flVOsPkjXShu
MlCiz9ea3pbayUiBiFrLlimp4WiIYcbHK+ykzcjB100XlUtCg9jW4kaMMN/G3zorb/rbk7VguYyD
Xcoz99MWl8LMKblrxONSw2kZpX+0Tz+MnkgFE9ikZ7kUVRcEwkEooQMEOs2WQygt+0VwRQRbjULX
aA74Ruu5OFiV2RV1ZeClmsxR3sF/9nXaZKTk5fmenITH9ied2aNDrhkfyGMwmtTIylwrt44gDl6W
jQkmfEeAygNlY3ORy4N63i6kBG18fuFP9v0yHuO2uEhXAuJIEjPCtJsrpVJtbxsuO9gtenla+9UB
JnBchbAftp7mtOd+9O4ct+iVXx4u2U4zin6zTCK1OFZ5lgCwnjSt6B+e/aMZiSzUH6NPOOeg+E0u
MhDd5oTlWn/mAc/XOaZJFkC3QQl8OZrp2v73n+zeqT+vPr9gwesw72hBX1ZO4hvKUSkcqbCOQMzn
Nd+MA1fU0AkY+/9nFPYEXS+OhMGtIrTS7IgpUrmOt0fCXownAErUL5BtR+EBYgPW9fqshmR4C4O0
em5u7Q90q/X3LmQObBgFXRm8kKcEKbcVT/S85w1dcZE3MiNHUN/JLvVBDPJ/YUv2r6kDxn/Y0Ooq
bC5zsn2TptfZFOpw8Yi8+tq85mlPvv22WE25lPJt5vyFJoLTd500kxuSFeE91pKk8hLczcc8JqcZ
3CbUI0f9ZLRc1xi+7gXfe+M4oaIWMoIj03t0hQ3kjZug1v/7eIMv+1LLIFZNrhe3B+vaRnjL0/Jo
7YxM5a9IvepXU4GuYnD3x0JfBAk/jO9Owk5pw7DS3CsjSWXWdJhEhyJZcMTh7iPZ69AAlAdg/fJa
+oBrGuyxcJamMWpaAKN5qQLJxj9uuuQCoh7b65uXPuq74dijVPVYP6FCVqPlgQhO+ORkhALWIEOp
9aZcrY7oIjT0RqDwzavs2luidoIpRvPWAZPy8qCt5MOgatOuFI8m+0vTOUXa2rXAKpFAG203s40+
m+x7WRGfde6fVa8j6GwQh8nLpqkPQkssjKDsaqvMRBWbThPApWzY5lpZ9p8xcwu4An/eQdi4kF09
RSAOZPlK6k20Ui1LMZuDd6NkFpvXkC0LmzizbgifRWathGMy04j2aRao0rOXqiygUFBJ9eBt1CtH
z3DbgjmcknNGBHhhkqY7Povz37wn4KLLiyopJCn8DxMsR2xAUvRiknDv/pXTBUSj/u3uNLAM2Sdt
BJSl+pMomQIg6dgcqZ90uWajS8H9VHgbdX532UFEFmPTYq7GN2WyQES6WffM6HabgmhqUTiK08PV
Fnhv2nU0q3CkYIvTUQRdwdKkHf7W/ydGWnYkh/qAFplFkdTxw1bKfFUmuz+S0+PuyQwlgQ33hKYr
cPqWf8SOLwZUJ0UlQgDUjEqawgCre3ReawSZsGd+lAWQ9mSu0HYChlMWlkiWsO4xjCxTue+1mM40
qwHLiAbbUwCORGfZG55dZOa5etKrR+B51tdIZq1eAWHE3pabQ0NelfogjSH6oJfdxR4eI7JbDbB2
jUAF6ByckvksyBivx+aEpfjPhgfp/hjlpU0sL80G6YhHBMRQ7HCgajf473Bs9vp1vyBe8p6+JLiT
OOVpmqIi8fxrWewsJPXu9jBsQottwJnkn4LaeOuJq3JDTMpO2+GO8Rujk9b22ch6z7O44sofUYDx
dGheSl1O7QyxnlEQRA7ijL012QYuog9OlHV2noquJMl9ihXLLLJUNhy5+R71/e3YI8Pd7YfKwU13
QGegKGkREDwMLzNcNXFALs/TAoosKSTsHWSVp6A7ZfrRML1MzfooC6ItjjVM6S4rB2RKuM63UypR
ZDQueZEyCoK27wvNSzCcPmSsiIR6OXo6rXieQ19nBxcrXeKXzUzpzBAMW/SOx/4Iod5jndnqHH1x
pppibImVvOhI+Out427bG9BcBr2QQ7jr+DB9sNtYOkbabxBhPRUkl5ZQdlKhzNicFLtpRPjiGD1H
BtDQPOr+CLLAv7wWI50+4MLSqPsgQWBkJOPBNbzXJKt0uV3KHERDLdGdmrg/h2jOIZVqRD/jz4Mn
i7e21dZFGlAfdPTrkIh+qbm8eBbsqIx9r3v6DDEZ1sblKljU//+6ZHNDhGd/VRF2uNyVWxK3YiC8
oSknMtd4ZFu7MVB1UXg4ASnT+xMa+3DSufWPKd0vAwvCJe/vtNhPx4g0IvDcZwWjkuCcuB4GqUu9
KiokOelquWakKmCEnR6DgIXOcsqDbq5LpnIemb7Bc4DZ+ybtykYgNjbazpW62tApy6PtHwB3qTEh
3c002vOUcSBPJr/HDyzlkIFXdzKEtR0ZFemVvv1qerMDmByazCjTPEDbnysIffBM/oF4mSs8gK6h
snHkk0tWHv7OaCyf0zwwINTmsqn2LdDy4id26aF5PpGGSAWH2T7bf/yerelwm9yZiedT5g90Gnyv
Ia1htThOglVDWjM8lqPCfsYXfcKpTfBtBHTeVgaBSPa9Cdr90tkH7Nrz8Mn9rpiA0bMN98x6M9ju
o6lyCoft67K74Uw2jcKzP3CNvTdbI6oUkoPzwI/G69pavUMgB8TVzwvo/HKCQcYHrgkP1UXqQxqY
1aB18VBRHqUl4Biw3cIzqxgqCIAnT9yq5lSqofOvwF/IP2IYDU34Qt8i4n0iVUH3+D0p68H1btiz
kBJ0B9dlnGjNZADKA6n+utq3uppajJaRIPUKe0TV5VkggY+52J5+EV/4JyC00NEBUFm9aiC00JhU
4ppYw1GwQYqYLjFnKaWCg+TVtuB8wWQsqJ49TpZ5XAnAP5TnSuNf5xHD/gjNMP96uyuquZ0AzNjL
KVz99MJIt5++pDcrdMFz9YvR6nGzVJaI0kPE/Sq4wz/6RkwhzjMB/Dl4kRHTDqp36oDW5ZCVCfxy
jUEG27FzmXwRTzWwgffXPKsLY/W9FAxqR1Rm3/cLxKEmiRdr8P+kqQGBPnEDNmkYWcabYA6YMYNx
Inl3O0KzQdiWcTe+tHMg04D1By4jVp33e6VfIwN5vo8hFsSOF9rgjm0AQE+HCwKvCl4P4EXq7zun
0WIyTlOg/mshn8NZrTuSRoefU7JSUwu6ShpvtlG6epVs0gglocwO2bZT7bj+daXXSPDcmpGMqTjU
4bY+Q0NROxq+BDQsd1mIjFwDYDg5Lc9bvDSRoFl9rwIXC/hlpEdonKG01e8Os/ZeeN2o1XfqECRJ
QDndEHHjU4hIfzssxtxjvnffttZCgE6dRNckFqdngAY5QwKv6OpBto8GD1c6uqS6NFk0gCLI+v/p
djBnjbv7xySo2O8dF/HcFsL/dpcWOkFKRXjwfXgY4eeTxgR0rIWqvurw8k/EIRORBuyP5lgQakpU
a5OUX9YfzWOQf8RS/FQum2W8jSq934cVzqhiYujQumpmwfHc8Z3mEDyc60mV2d+ORcy7MUQgoDsZ
4/GYYXOCiwqRv9fUkq06LCQqrsEC7N/PVfnXCGZ1nndpkWfG6BlK3/TmVbTssp34tK9ewEOelg7K
OtxwJg2AO8f6Im8ThMpwkpSvKxvwiuIctNNAaVaRibjdMpVe1kEN5ASAEI+AKzuGaIquyiDU00mn
w2s4bb0zKC5Hio1N9Gw4yUr9ZVqyr+10CWLT/3PG2dcvj9VDt4JjJ56/zGxZz0XsiBzAfJud6cJC
YG2ueCyVM+baK4O2WpxqR0VAsx8YDT1qcCnr+BrZmM8e+22yhzOrxCESXTXH29Zhr47tMDfPy9WT
dzwlj/vSJmVXn3EBJKeA2uazEMl+kGbPDK5iMeCaOOvtSSs2T08XDzcYgsI9nJz1NzbmHkAxXh8B
stX/89ZxG6H8DOCewSc1VVf+0+FxIJdxNVsacZJIJB7R6VG3Gk0slxn383+abygduHUNl8MHkOpE
pOtYFEK4CI5QjO8LL9PaYR3SarV8EL+LtUb3WBOnPl2SNkw7TpgHOkVIcRmkjW9/ycmob41rq5Dq
3PiSqFak4oanLWOwhmexA3WDG6Hj9d26DfxJtP6kaFF3f1TNCxJVQ+y+PpROFzWVzhgl3aSL6kA7
BBUy32sWNVzNZZBX0pRsyNe10x0QtlY+zAOubDIZ43TtM6L4uwshUfDhai5gehL5o1wbB8GNzprY
3CWFox28LBSC/rXRe70q3E3BwmQcp8rE8D7Fq452o/CgVLlpO7k5y/c+O3Qe6A0fk0eO1f/wDHwv
q5YXrbXNAIne3hscsiLf+v0g/evCFmDO7OrNi1tJ00ZzIEE9gR6wa5yNLx+w3Su2jkKCtJievRi0
iwQypOJOStDu3e1xH/QqcTCIuxK2o7XPpH4Mi1QIS92zBvUljS50PN2+bYIKGItVg26TYlUb6FSX
ut7ETqnmqg8uSOvUBzCtqZQP9n2udG4eluGFrXDIoPHv1I1we7+Eb9EsjNpnBqDowLV/nVFieHW1
nj/4XwvgPdwsAsC+pTyyJfqQ6QoU4152XHSN3Q4H7C8aOOdGl4hiAepqLIboEmlrSZqnhNgbAlah
LNW8X5Og3tbqUf007xiHld1mtsKo+F24on6xJujPK3hD2rGj+5k/lnEp55QYafm9exuo8EIu9IKc
A8CrvXUhEK6FDBlZuJFOiEwxC/hBCeziEMLhfGUlDhY34EgmGXAYF5g1ypNa9xkUAx2C6jVAcvwX
iYARmunNAE/SZWQ/AxVWnBbw+StIwPyHyZ2fDLxDLT+KOLHyGwVU3IAtkI2bet637aJHA8jnm8yH
8SNbsPkmGe3PO3+AAotlsNlZu+wZJbl+OP4UcNLBWjMv4v7g279liSugWbjgTgS+fNiD/IaXRAPy
ABgHnl40/sXWwUBSuvmCCoh5yybBZ53LdKkNmHZcFJvNtdDieLbdYwppmqo5tknUQN3DTixUpQ27
no71Vxf6PR4sB7sPCsTsjioW1J/Sl1Ep4VX9hmubFhpdB5rre687dQqsyj5dCLS3aKIPh5r9E0vg
bNFCCCVecMzlgW80vdnEOXW+snYl0+EFTKQrVBL3tkXIc97FxwaupUEblii+oj5qdyUkSN2Gn53Y
p3zWJ6vX9dThloUwf1k61Pfl+G4GxWVjI94r83GNBxKMAiZSmQliM+buGVEzvmXQDSCdsaC7GLep
exT3CfqK2yzwpEEXAmPaxwCOvjJXyqnRknOqvyjoEh5XM8ylJoQJbactpR749+lLMpLv3h4bcKub
GzaLFlYPO79bXlEyiLLz43n9d+xmG88/K0byj+hXKjUPMRopg7w0sEXvtcWNGczW0TderOjgRgab
fRY6Q6aH6cRhEh/XPx0GrxX1JhsXLctiUZNKDJjA+lX02FxDmNGRG/fXFV4vLXyl9qG//KwVsXPi
zhIF+Os5OWJH5cAZCYfzDWqoYfaBR27OAh2tPecpEiZ5Pkgt/JZyG4gEsZK3uN7jr2mUsIt3JLl2
jaEklLHAUPWYuPb4PqQ9hajVa93iuOExjsgBwMBzGcZKOltHh7CSp7GPYo5zpEIQXWqmeBl6sR01
sbXgO607XRAiZ+GG40GOduffwTBAuqfsHAIxWAatYmwKIyxL/6HP84GBU2jKjUfIHdNPMcI1pCv9
Ca/H3vRDLYDgRDZzSdqWEAvgZwP7azBAeWjBNwJrwZx4KfNYZ6CYodKJ+yj0dz2Ezjd6re/SpJSz
eMG3gDNmTMq/0ysjX+U6Ef+qfvjBvHvSX2gR4KzbCE/c4mPwTEsqkedNEN9+fYwvFfKETr8dHYyk
sjo1M+4Pv0OHpjFACLJazG2DuTTpUUEsgQkQo3IGzT8MZzmpzRqxc8GesHAa9AX7sy6rB0mRUIVG
NnFpG2YKGU6txCdGltviCaM2Qo2DaUTWn5R3R2KmGI/pJY1O0QiUB51tDhzD8QZRwx5OTZRzCiOS
wTX00A1yoK2lWcNggqxaDfA6VY31g1/I5R76T5pIWy9JZUdLoMmBH4IF/MYhPWnilkgkJeKvWg99
RWKGVqDSMMXHqAO9l+l8Qysly8LWAn5mlpFpLOzHKXUXwzooXZ2rXniWUNUnxj4htO/8xJbDrFEP
9l0l06xuES0VvK2v1Nc30mTz0zU0lZyub1miCRhjS3NC/HtowbpxtGKqXo7mwWExsQEZ1G5j1JKD
7fE0pL86bbljI9ZxgoYMFt4rkHlQYNNJ/SeS1hrrOhcM8+Hqz951OoEF4L/gfgK9MGXSUhN2iKf1
UW/mHIUpjmoe7hyrgWGVmV3rN05rs1Xl6dnxC3Vt/oVG9PNljUTOo1bM3+5R2Avp0QJlLP73fKmy
wPN8hRSbGvWRf1M2p4e00veBQSb9T9QGtq5AkEKQlJIPM2Na+dH5W2jKVMUizaudV6DYOZdB+2tD
AOLpZ7z9WZwcQzFQP3r2t0IX8/043W7chireUufvoUQ3MkDN1mpuS2lpei6ibuR8QsImsYcwc1El
3QdInnW2c6zeslh2FRJNk+TlOnjCaOBqSUtPQfntlVEzoRDtaARQsFyP+CMzh2UkStRIS2oinMsb
pMTEjICoFfyYa7o2skL1r9ZidyB0NLTU5hVyLdc5oQdABF0gs6ARCc6DM3X18p/efGz4sN3L5KZc
aQYFFDghYN8Pqpqp0aZim4ATtUQbZ4v9z6fMPZcDWDPUtAGHEMQVuvc34VRjgw8QRd7SuDOo7plI
vZDjTusQ4yffckdgxaFi4utIn3RbJ+Abmfza1UtabFEwnXhfgW893I7qHwFioCsZFvZBZ6v0LJTC
49GzHQ2YbcB2kZuLAFT3Lu7ptDg3y16MTdGxGmgqVJWVkpX5HD6YJpDIgG5TK7jwHsHhUdwri3QB
LLsyCaKOhw5Bd/pRIwLHvQEhuHjydvIuOcAYoykD9pD2qUbJLEdLRuL2weCYvDlEgqRQVw321qtB
AeLq2ba6TzUsecHXl/wlF1BZqzCmWo9EYh5ERlsBokhcU5U3nRQnPq9je7MTEChuQB7f+42kEUOn
O9q+zOUCxMrD33HtJrXs8UGQFCeedPdlihx1ARMBYo7WBQvnDRyyqT5b6Uu5SSfcNws3DOV2+1H6
imEBF4W9afr3rgKrrO4athmqYq0MXLgNiWDApFPw9aDDk+sSr9getan5KshBNTDIP9caFOBnUE0M
nxpZ2SrYXlAHTqOPt914wjeJDL9gLoRc61xv/1iaMey0QcmGagKDvlWB8RTSRy063hrTaJrrEAtE
U8/FeRxovRDTFpQVSLa+PFGWQNAXRfdqNGFK7GyywW2EscUu77AIoBrEYy8hVMx4D/xVcZCuWN/+
w8dER+HmLrw/mxbInrXs9UiPRgK5eEa6C6louFZa+hdZCfcS70ZTSPolZoo44jeI6DP6/gIdDpBu
tpKdIUrN8Dxh7wf7EpQbYfy69CSZ+jj6VRlcaNriI11DZ0TMW1p0H+yS7vhuzd0DPlEoMUM4Jusd
pj9835on0gHrD/Io7LdOAz+eIUSDnDmrLpV98BeaEO37rjzjDynOs7lRzSnZGMj9dJDy1pmBRwMK
rsXd7adNL4i4CtD9wXxdTsmRZZYX4SEJdUj+i0amRvs0mkNWVsGmGQPNV2PsszhpGh72SppdX5lZ
6nWE9Yuxa2aZKEWkX09TurtaqApLux9TbykK/jA43n22QBF7Vry0CVSm4oAC1bMNaSM+l0Y4hmGb
jr0/ytoGJQyw2G/Auz41XQ52sys7rOlvICxcPitkYFkzFJ+SIUYIBFb8LHe+0Vo9zvSgE7GLUeVB
2wC5Ehi4RRugwZP/GjNB065YOWPQhlMLQ3w1T0tNl3fH3t/UzJzccS2TyBPev/gF0M2TFUzON2eJ
nbMpSOS7df4V6c+vNJmcNw8uXxxHL4+kOMlSf6Cn7ZaBGMOKU4fgxAo+oN83/kmgYyNSoj18+0GK
iSQvv0qpQML3YFnwtCOczDMIHm8EJH+1/4yVMWRYEFvmZssysP50+SXnf3LBBJFaZYoFFFdd0Aij
7FTUAkBIS6L+rLibXMMLc9Wzo8LPf1qX21Uz+l+LZd6RgNx/cC4eu0GqglOfLEdtQ6EyjXsm5IsQ
IM2kI8wQSOPFTxKXNdQNR6tJ4vtEA5WvfQiN58J9tAOmeYvd9lHjjMU1uS1o6DYogcsFDMVOa88X
pKsnXuz5qWmhrJWEmxdaFUGyGJje846oLQBlU2NXZo5lT71qy9bpUrFq9br3GNcnRTU2GZ44a+kd
anjKhScDORqqyqFCXwnwKbz4zuhnl3xb/HbMvhUjs6FgrYAXNZ5AbfC3goIbURaqnt2C7xPqc74N
LKSDXmCygGyMlcI6DXbrd9wE3o2VvGod4sMqiprumSHgtQL9qxjHxFyNObCuaVLQ+3N5zWlFcWq8
6+iERIS1GnWhQ8FH8iNFhUVhtk2Qi7rbmrnf1OHY7StGmnmlpnDVr9JQiSiuQsjlV7jJxujkGmGM
67uwJlOE5sujG9JYcTGhEjCU1SZsfe0oP1ONqEa9vPO3h7Cuzbtpb+fF+/AB5ty307FTlSDXTzBS
Su4t0IrTvi92BDTrr1sqRnVmJrebIm3rOcI8MEbzcACkiHOCqPX65K7XzjxIpU3O0FxW3srES47O
PrfbC61s5YYrOBq24wxI6HGAR77To7n96uE+imyhtJgeUVe7rDH4JbHhvjPCEgrSahTlT2FG/XKx
jdHkm9pwSFlQ0IJJq2GozUCWZIXDH4KbfKXAu6Hhr9/t13lQxDd88a7EPl8fLajFtp9UsodqFtSQ
paJH7hjqENAcKkG9nHZhr0HY2inXL/UblxfqAAkC61TMp6yUIES6rS/SpFfeFekiEoQ9BNKC9f54
cacCK/HDG7UPFtZ8Twjc02JZb3KboYSrvhdlFaLHODshuq75oSffUdoHKGrajwbTSWSH8+hs50SJ
cbDeel3lQUH2954P5EajTdMNo1pn4HrQ7wQuODL2iTldiWIGBcnNyNgug7jX0K1eYPcXnjzFxWFo
Z+mk0KB348pCrA/Z6ol06ptCFRrkeDtTwvM2aE4E4+uH81/hAHZ/YK3rRoC6mTMouk0iSymWtmXj
LHAjAPL5UwOedkKctcvqyLn+qG5rlacpix5kq/EHgxarqtCmtp035oZtV6yp7VytKhiLxcB8fQan
XnCoU0v8m4SQBZRj5Bh7Gf8NHAXN7bki8O0BU5YlN7jCtI84lhhBCAf3YGqNtjC/jHlC6epSF7Iy
3UoVYjPcfB2bG3JbW8aGyZylrZ3eYnFuyhuZA+OGyBDCyEm3r1v5pjp9tESsOprRxI4vP7PuOyrP
SrkuSWnueI/Xo7JzRglcwxiBERpnGVj9kZRnfGl7ANf4FBaBHU1fxNSV1jiQj4Or5ZDL72Kftze3
iWiJu3IrxYJUTp051puo7KByYKBKtlv0zTBq07y1kvVSqXgzI1hjJPh2O0+hk+U8l92irVfGMj+J
QTAbFvoclEXIghRJlChb+C0FxFqJHnEJEACNDNjQlaMYuHRcNeCbn9FusZEzPFOJz6m/ReqCFJ/N
OwrDFGUuuMFuWsiYHCCHVbYdvwfzMA5rPuebwSA7egqtPhK9YJuJaGgCAYgy0W2BnOSBqR8QAG/L
AC6gUeUOvHkUNk2cP+gK25IPxdY0RSSaGHYNs1MiW4JZEZGEgCeqmFCUU4QIuaGL03b2ZeGibvhD
K1pU8Vtr5Js3PSyusOmMsjLMr/Rvlh4EPsY6l5RZp+u830c86fjX7fla977+NWeeHjRxxW9lmthb
dEAjWaf3YcKJ+66WK2M/egUw9k8Y7Tmoo94sZsPaPQNsDvF9VGdS6UnvBiL6AmQLTg40hiD099wE
8ARiK9Q6dC4oMOMfpxBLHNTYdF6XdQsld3fq3lPX39rixHQvQw6k+ui849celKqHzmYxtPXQdFtY
2S/1bCQ/0DgeaRcO99EOm+wW/t9qk7YBrOI7vABwHWatWKS4W87Yc7Oquh39EVjgPbdPOHGhFIqS
Zs3U5sIyZeDdFMC7BqZXx3gf5EBpIC32ptQBJEBZERrddZCHXUOlqxcVyMoPresjrdNx5WJD4Hz6
Z5xMFKp3HkZ2k/0gmO/mJAazluhdxewWxQ4+825kprtW9HxGqg42ZYZ+4Zik9tkBhpdlpUX5ROMK
PgBVihF+stc5lNKReYVWb4L/5DHpHePmY7axrzikOZ86JN6zXXyVSfiEx7CsnrNVj84MMvCBkx3S
3cqHtOfiF+sqa36DQCZNwApPpQt538QibijbT4HdFvB5W0rr8GWdbQI/7wVmaSq/0+IbumIK0yv7
JiqfpnCQzysWkAV+2Sm4YJ6TNZFuGOYL15lxIbUZoLUz4Jkswj3a37tvdZE4f0+xsjzPKyPG5Psc
I373O8kk777GBC+o+vIW2pj/tp43FUERGX5SugZpZkQBcAIvmNoZ99Kf1FNi2W/8ZwX7abAgbPLO
Qc6Wa2xZenS1lf9n9A3XC5tX6m9v94IQOSsaUcsqYtWcPZO/SIPlc6eDwbw3W9QyqiYyzWhpdJzV
plPmhSHBlOjpRlaXR2NH8HBdCDLY5dcKCHl4yy/9Wl8iWSG4JqeJmeD6HrW5fNTEtjt8x4vqu4xW
HRKF9BoHHfUXXih9ir/hEhjmdLd7RJn6sf02PiivLxrq7w+TEewbGKo7G5HSvNSV+dhlZEpaTkbJ
PDWoSDT0STYyQAmm2+3nW3tBlzVAk9uG/BmlyO+6PI3Grn1GUfWM91RyXXgsVmGLUS+thTxAUUsq
kFlTd9bh/iJj4Qw54CndCsHJ5DuZH92rjNXi8T+9A+6cD75R32bmCwRZ+Ssn1lZq7wnqfcEdBXh2
3+6sp/LfqBFBwNQn0RInvtw+tBJCIbZoErSL01ltGK8wPRp8sXhe7YCIJcwP8V9qdjlV6JSXfaXE
t0lv6osUR0YZOZ2uqVkC6KLjnL6LNWsASmB7cN9MOZu/8hL7EPbMIgihI8tN2cZQm4rrjcheGXZE
exQM+bWE5Xg3BshFfGXZlFglpVpKKpsFsPuJfDYKcj5cBePqVpYCwKPzCB/bdX54LTvEs8VDXWq/
iDLv8KgaqP9TyUEbvaFercnAzgmNwldwrwcj8/1E2GePllVIlhn/ZMBaOO7GsMCsDdSWXxWuWcfV
exdjIec7u8kWBuc9PGN4pGre3RWeHKJmm2MrsG2P6rabCF2BPVha78zNjKo0f2DdtSMTtnWJoNcz
YOdsKSbCcbDGSVZ9Nf02Pt9qxRdZ+Ua/6dH2dtLRQVVLtZlHg2yntH1lC6z4FYMhB9OyB6ceEVl6
yvbkysJduPI1LJQJz8IbYsdBA3kUCxFWu1Sv1ECN+yDX2Ma0tVStFuwhlWO/lxlZYgVzgysF0Jk+
povQAxpKycko2vJqslccRmbHlw3wk/XmTpfiVtBHaMPI4yc/hHTd4AVeEa6gTJ+93QRNpUklWnXU
P31JTEUBpyK+48qnu3fgkeIeKZJfD9DbFf0I543XY1oyD7Weu6CwUdEngCuFqmASDvPWgx7omiEA
478z97wKkJrq2Nyqy7uZnmVxxjXotpuqwBJAfeEFrLE/RMTY5EMMzcqGtj4dbebNRjqSxHLjlv7m
VvAyZGfXFaJZx6DLw7Q+Nm5wrCoDyy8xfeQmfL3E5vzEnOUAg22B9YresAkrTc9C/4dOdGl6KCW1
xqoPD4QXP1AwwFEtG5u5dHAPy71sDp0i6mC9mT2E2MoDzDJ5b8M2g7nLnj9Y0C7PjlLq5Oz2D3v3
yus2icJf3P63UTCEOH/3H5fz6eWNw7b4ZOaVo/Cijgmdc/XQ9IzJAju0Fmk1qr0QRHeEAyU2KD+L
2+802YHZebWxRvOckmPm1sXyXcygpdbFLPNElgjsZiC8GchFfZzKj7k7rvehSLbEfLfgwrk+2Bvw
xTAqVj1fsEZkOk3dBYclO9s9rnuWNsozHfjq9AyGUBRF4DfqBUpMaOaKXxRinwh1LWhTNMlYSz4C
0v8w5++nLtIo1MYbllrC6UKJYvPkS25Q8hVpjXuHp2cQdZw5s7gmqnTQuPhq+tozJ6HU9emRX4T0
E+ylVX3BXNZWdEP/hYvCDrHB3KLjq2Im162SCRcdxlZMOkKYzDZ0MxQEFWjfMFHv7VKbkusXpd1K
wZtxdZr41m7KufkfLrpQKOmZBeeCGdyET2bvjxqjkMsdTGFuwK7NImCNXmo1QNWBIVuxAko5rVCh
n25vz9OzTv/1FJD5kq0dFZNAsoZY7aNmJljlb4QpWs6/2/c9y4kU1en/f6chSuHZP8pxlban8hfN
PuELWerf12mSfEkp5iOrlYIr3U2PP4VuXf397k+mD/8id0LeQ5OaL3mfSsC+CR6sZ4KfR6NUU2eR
aNOWBptyC4VYknxexvja1zsGKcuhL+hltUXygVcTmmbt3QV8f+eTtSIK4BOp0if+LoJkPy7dep+S
JKEC/nSACgbezEXnCiGzBx9TfqYKhSa2Fg+u/yR+A2Bu12mtAHWtO+vnZvnv1DPmO4A7LGaY9dtH
Dl+lhnix5wc7PR0GyoZFdYUxflyjPmLd/2S8rld2qEP090eRArDg7p6I0dG1DnNNJJ0JONFCxPYq
FrpyosnZIVAm/15JJUsxhzzLu4cDTVqQ/Q7lJvhmc11IVFpDjQCSdLmIFMf9KxXCacFQ6dkpQX6E
LTGoyhl5BPnf4cvTWeru+NQcvQJLaFssYEmmFq4gDXvGHJf61VCmEtw9Ec2eoK/cLCBG9PGQoMpc
oUmyXJGfZYyTZthrUGPDe9NHmSl6LTPHib6KKWq0SHJ9kddDGmcqNKkb3EkjAmG5X22q+IPPd3Na
OyOi9nrDgerrkgFPL+g8QseQRmr54X83hfc+i15zn9knWkEjkvtjlSQc26JQMHlc4WHXrcK1qgis
iMvCRINxf43O0u01kOW5NeQmrwVQ9y45OA5UW6EfyEdTDfKJW2zISYegdiL/C3vhZm9P9EkmJyHL
X7EJzMIDX6HqpS0jEJ7A3WeYRgBvktvyag2MCqFsEipB/Rlsy2n1qD3cpuOQ35P12vty/jz5g3Z2
s9xZ9pKGmxYoCmJyJojZ7SexqoYv7z2zjW5T4MTY5CQfeW9M2SPYApN6Q2LyOSgxS5GPeuqLqGdv
w62jzxw0eHHuAnK4HGeSDz05bPLU/L8xtcouVguw+gy8A8v93of7dQtCVIUPrg28faY0bSJk6EJt
c04LB/RjgMx7etEXGfpf/KyKzztvqYAtA/Sx2EANMtGx8XqiffCg/96okBgqdbZjsJQTIt7Jmkb8
OBuuSI9/4458DZ97ukMUW+OC8fakrKP4x27VBUAUzh483JypuugWtlmOr1RQio+jEHemGad07OZs
s9KyQM8IS1thVV2tSkMCcrZLIdownBca6NsHRcHASnOGQlThEeGswDMTcm3R46v0uRS5P3hfaPQZ
n1imMtF6eFdTf+YzQ0DjBXFwUqH0ajwXsO81s9PV746B4qZIKaDn9FT88HAWvlGI5zSQw/Z6VJPb
U1//p84GwR1ZxuLvMZnRQaCNNeQNG2MOrvLIWcDTXNpopuvhZWKsWES4iXnvPFidUS7/HufkZH/2
o8sM/tuQx9rqqYBe6aTCcPNMW0JMO7dtd3fGUZsFWWUpoowEm7XXgDwCMYoyMNBI4I3l48RbmSMT
hRd4XLp4Thbg8TtdMDua/qLFKkUFFJ/A5hv6vTwh1aEbUgr76HcZiJ14wrgGR2eKKbIAkFv3a4oQ
KdyVOLd6m/ofmq4ZYSf2CXlGPQVA1Sg6Ae0FR/o6Nn8vNX7ihWVp4R+Z5OLIpjQzbtV2otY3QGHP
/yx3S4HsBWdk72sa1XiKuP8nMR1rruMkDFC8NVMDTiRIZ6EQmiChK6w/myxMyfjdPGk0Abdp26I7
acgP5jprRdWnK25HpVXtHA8s2r4qOvmXkSc14QkxEMQIo2a77L2RCruSaU9DFkRnzzcwSEY6VISR
ly+lrsk9EzWi6W7byfMCZvuDw3WtH40LN6VpnehsEu0u3CpEpZkZ1AaD++0MP4xOM92ntCIBqRA4
zBltw6e6jQPl4KGwY4TES4MVEovhg0PfviTm4oBU9T/yQy2UH6H0Ec555Thc7Ec7e7j/Do82s4Sx
nwIkCDPix2fn7cSCi+dHxaeMTthuUCvQVpUCZqzN3zXoYDqoh2X4q9X1TFREAbhbjRkHjmoY8ZMd
FrwlhpGB++yIhfZSk37D7JyIg+JFP2Ga5xnTZ0O1YjrsKtemkUFNRg05cWQiiUtDmBhZgu8sVARt
KHKBBB+AqJ75mB8x6c0lER57H+ymBJ7nHtwsHwKuKnIPTV6tNmzobPynCu3RRwSDVXqn8MJGqdt2
v4II3UVoG0jbAVLdI3c3sluoMy3olSe98WnwIFDulFkTFzPpqTehrTBlcd9VoDQmG2iHvyJITowB
cbEZXtUbQXQl94aA6lXzeftfYGSJhjfnY7TitRlCCSlxsqDpUmlbmDNRT5j09F9sMs2njbukFlGw
2v/tKb2+/wL8wLKrTUcaVmrCzhrUivStV3KVodLVsf3HhxRdXcZJ6mTNCrIEJRdwfZb+YbFhgVJp
kgK5DCTqxMlXxLNruRlPEeO0hF9XwalsuW39IziYtsCDIjFZvbqPDBoacbo+QccS5at3XqXEuN7g
ne9V0f/E/HSiVE8rEXVB+xNbZ7q2Qfgp2ecPATCZaOniec4Qw3xBazifUV6nsFPVs17JlxkKqrwx
nMNicC7USlZbjhv5DXBEfk0w2Gjbkt/hijRSs0FtYBnTGMVc6ylxLCpPH+mAljSm2doDokvwjMpH
/uQj3bDSGDP+1ElJL9qXqPcSVf+uLnpieEDCEt8BdpVPWysg7M9NXcB2cxtIGPS4IZXdJDJKMOJp
iHqYUefZho6Nfrt1o6yo8ZFKZEg7cwbvWwAuQ7TwleRNIvq1G5KMHdtugKxzQRSbrdBlQcTD9O8s
HMIVYGIGxt8leAwc9yUzz4gQya4CAInLXkvNZ4AUg3fuQ4huorIcuQODr0A5aECs5kznHhLj4ptH
Gw71cmdrDp83ggfs7zX7OFt8HS7vluFA57kpoKuj9i1nNXTLRqTKw9/F8FBPxok1l8eXKWyvmKUB
267rVTkUyXlzy4m7Cz2Pb/1BmShkSX2ngtWgCQ9TzBPCSow8PDeYxCUK8pa1PZpyjY73z8IIJsWB
jgTwfIxj1owZz3wwqncJESJn9t1DbcilHlyUeGO6C6zaAd9vLdd9PZpeX236iP/fdSm8Hl3mYnVH
OKyU8JgIJ2omSWv/RQT99t0rGLBQ9kexmBWn9CF/heo5DIzKzfGQTjSkOa088pkpTP6OrnUpVn1k
e9BUn7p9dg0EBksFwXcbOBusjF/TP0+l1hizmXdbTIPC5Q4lxXy8jr5CUmw2HaGY+9GjKUWy53C8
KVZNGMUHOan00DfESguhyBMSNwMZY9yD+dirHdwE9UyJY9D6erkasz6e6K74NvkTqrTB3QQII1CQ
Qz4KQmUhY1EWfKGdNmMkM4CYZzDhLowKtYq5/eoWbiSm6eeqshccfZZoIoI6Pa0h+Yfhrv39O6R8
+odOiV7/4I9+hOa7funwyeDVtT3tyQjqM7mJxCeTpGFcTsh1JJbLbe9EFPao+FvCU8SBpXxVtcG2
y+GGAY05G0PAKEPf8lwqbYqS0U26AbkdqSxe8TU+5SQ2kaZSuq39s6cKTy5SBjGIYkdROL0jiQlg
00AxYvPb7UhCLwsJxmiS2UlhI4erZsYfALE4JB6ZAp+bK2IRQxUi3kHNOiLN6HFjX23Yz5T3M+YC
dUOyNiM6WS5SaMuLVHd9I0+GAeEVXEaVjdfPOYO8CMJqVJ5rCfIZMQ1/rWEM1ta3QbaW/o66ylQu
n3ulwWEofbPTOe21MWRsnsgO/WLqSXDRMiAkT4Tp9QJbo+amWjbOdS6KLOBUwTfe3I+vNOnGKO0F
pAn2z9HoFPKxnPgPYEkuHUl4wB+lcsVHby4ms6E5ja8HX/rQN8q9Pt4KiIqmUIPnP6PCjGU3/Hwp
1k3s+qdk1BDS2j/p1fUVBFDYHDv/0dls4MSu/CV/9adj4+CEOsad4lMrPthrw0jrWbmw9BO8BFBO
p/XTfyJCfS17MvfQVRq09k1KXowlKn6pMLGsoqTHlBTlP/pT5T6ZiIVK5n4xPpyE8+mobG7hYxKu
bXcG0uXsHbfeFe2JfaCe+LS/yVKjZOulnAArCiujPHSO1OKt/2/QH2BFJvd4U+BwdH1NVRQhVJIq
S9QYgA9qQQAxR1wKmKmISQYqKvrBYTi+QMSH3h3lUjFTCoeH3EyzPvAa7mzoAFUX/5jPCyPNPqsB
2E+7ZLhva10lHS3c7qQBrJoXhVmDFHAODWQsIODlU6SVQPtBOV/GvPyk4iUUCYDq0RcygishhJY0
vGfGSQ7Ys+hHxb4q1DsTv+/taZUpgcDl4AbV/hZbeGCCJS1RJdQo9aieQN6VkwH8WclPEk40CoJS
Qws1JHbBLd0BfyuUzC7+EQlT+6TodXpHmizkM+WMAsHk2AAqvbcdcM40jGhL7t4motLf+X4Mbv1/
TPAmMHbvIYehkLaCQLcxOoyQHfaYxrF6cM0N50HRyshVbVZDWKTLpQ+Fhs/HFCdK0Pgz7NSL5kse
1QXQJ7nxV7XTAbxPI4LW1L1p/ypdbf7+mV0Scl/0nhTvzpWE4ggfEz7svpQ6xOkk0wfsIEPhUUit
zwxaRz/HdZA2i14VeZhoLOxANeVKmSGhYslvSpq+ueVy5qyFxJNM1oJ2x2jYUzVIGFYPyMQHeX0w
ohjsZUfBNwZp0Pl1bltN53+TEduhZW2uEo+7ewH3XOEQ3ylDvA6qdFGMjccEiPFc8lubAQz1tYDo
7o3V2o6b6Bm+Q9yOsmeCcE5exCXiAXLdzhBp8POYiabgP8O0i6j0TOIhblrBtawFRiat87KT3jcp
Hgl75j12w1TkdtPiX3mFTvVbe9QG61juMffwNo0NqPB45rLDYisBE9fOfqvFMgwpFMM+NlXwkNdt
XIHegxmkQQRGbUHcwLnfwAPciZHZ4Bmb5EE5Nh6Q5+4eko8UD/y9Io5j830k9kQlTMqMa/rEkx14
tETobS7lA8JWFz8mMze22wZYJu7wH1O8Wl6YwAgCy8v2GPOmji7FS0t835zVPEW/Dpr2NK5zCnv2
mLcmLI84p/nJooIsd15OdxJ2jkS8uUe+fyOBOfSxaaz9rE2WaY/tV4Rcu8/YOaBGiWzf6x6LeA9d
+MSucNdNtBAs8G2hjU77IGxlXLw6XH16Moc7Z/3BEGIV3fS8rUdn7qo5sT+vM8CB1dYX0xv2hUgC
mBoNdklc7xh4RmgEjsAh9N7qDxuXRyHJVRByXTJorBZFt1069DMhY0xlu0UN36/BcQBaLjARVVWG
RX/g1IfqQV9khmoIEe6wzVCmB8UjTLUA110VSF49ri8B4DIdjzsU/wQBmFoZRfU4/5HOXRwqY5Av
4jkALhZSk8XXUhC5r0hi5DI0Ays4lMbrB5743XKCtU+BMI36H8S9Pisnav+hFlfhN74DvM6yJIhS
a4rG5g0pTsY+HFfUfFZdup+jt5uGROUlLeH2V1sPgqGkJ+vj+YvGugjBDtW08Ult0dRXgz39FM67
rLDFOr4D+am045nsU/hw6CPJqZYMvYNWT0YhHoCuKAln0NhQzLFt+OthcPv9CMOzbA9GRc6f+j6w
N1p26JwYMPMLlSG0ixJK7jWzvLIsAcMvQ7pk9sdLvn9wgSuOkYTNboHcKkeQXNvy9lYPadifLY57
hAv5v/w9w7i19yKwFuVcfoBd36IPYdbcChLcDK1f0P4LNXSFRa/Tr33MlEs6bhXSkovTWikUJsI9
2mTO9qvziymrzfXeuELC3wWfFQbpOqXKbKKiCsMjpn/rkjZNUMUD+ikxeMDGOx0uEsBMAfa0dkvI
EzcfcgDp5KNDe4IFGz6ad86aYhIgi0e4nAeY8q7dZG7XDYOIyA0/1mMVlErFqVeNftlMSla9ZAAW
dIsaZjhjXYeXsPXTLncAo4QxBMp9XKur6NQkY5a1DGhtTIJDQNq2YQBayDHWXNR5JAO2lnCRfXr1
YgaWdXQyYLq+IQweQqSkUT787fUehIt3X1By2Fc04r+cLkN7xqZzthiu37GBICyeumtoy+kgNzlL
kEF784yTX5tgoIzkhiPH+WaPQoA82fvnLgvIVCv+6v6Y57kfTitnpXPQDIv9aYRuCkrVRkiDfkGi
6DdC13HlCFv/kiBsxoq+ounlQNf5ou/l2zG5jlGUSrUOzVfQaTY18tkAfhaTO+LnthsUqVkHclCc
j6s1WvmsUYh3SVdD2fG2TwAUfK/uPvshjNEULtxs9tj2S4BFbRmZXDhmRtQjIc959Meh9tr7SKFQ
sxiOYhckD8huAY+ck9PxuZAkuN4E2HVgh7QJF5gz0sGSwiHicif4uXuvpATM7G1feOEPRssMSn8j
+CGx+orZ2IIu7NGUI4t0Bdjj1e855h6QAmcgjRj6s/5jvlWZMiw6bXbtIP/3dU35SkIBPyQuw5vx
cn1mGkW8//c88d7GxK3lnBZPA+bqTSnwrtB1IdcviXraKxlZXNiuP4pQXXQAYNxWnaLFGx+QTzKX
h0tXFZ7dnWSi2LZLmQOPAeRrCa2qlXI4uwbKyiVV4BAWemZKMIXRf6roZnV741eJyGq99/jZYWh1
3LPTI/CK4JnURJABXIiK+dUxtL1EXFC4k0at/Gwx7b+6u+yzSnr69drLvRNpRP08H59swvScrdXF
TG86rdzgVkEE+qemyuYEorro/Yhbel6WXKigzDfljFz5FH5wyNiy/c4srCiQcPglzVX+8/kJmBr+
bAYq1upFI965ZAReJ2bzpuDsgD8yb3Mev9v3WBTL7qDRIRVV/hRB9N+g+JkoyJR/6mufCgDna/e4
6TaYdceqz+m1I6Dt83zj9+FDql21lJfDvT7iomxp+eWt8BkBSepy8dB0HP4l75a6qJEgT+tgWlM6
bSYM6ZPF+SjwTPMbfHqqMRBfgQuBXEgOwQ0Yg40YyQWmOXIQdw4vUuUoBs4qaopCnu4MFl7VvIQt
hI3X6tRgKxl1eg+8TBhcCzv+BXIWj9YkteX2Zvy4aksHsru3BSzvoiDQHqH+RegL3Fh9aJiwR7uV
pyhfgLKLfYXtNrADRF3C0ah2xILndjP0f8DaK79vM1cY9s3dn7JsyNwRXfIYt0v7MJ9e4KE9dI33
SGOf1VOVpsewCNldZPkUYupPXHogqoKvq33vP6HiPWuCNJujVY6k/YNBgL4vwM1tc7MGLbz16pEq
x2jzg0WnD+jgDzB/0kwdL95UASH8bQ4lMlmVs/saX35gB/teGlloeXIRgxkIJvaQW/6oc5G1G6LZ
fix68ChAjuekNETzc1Rvkwo918Y3uofave+lDOPOjMU1HCo9bKNGmONg5njGIGygUaoPI5LN+mbP
ztAmR3+CiNqoMW1XSf8s8ncu4gXBfNFqo0Wvr9ijH6GuKHzkY3dy4kHYAVf4Qg/jLNmY769ptvjo
OOrb5o6fSu4ZDQLoml3o50zcdZtRhXLeFo9vY+0XBa7ahiXMnLDEl6s8uezln2ix6hpKvQ1Gq3r6
aWBSn1nJXR+nwo8DkZj+/OURlsxoESpnV4xStb9wxTFcuAi7HHizNIl+tnbCUkVXSYQ1KjrG7JB4
hGVtbgxLfk38DwwPNMbm8hZbZZEOnCZtvDy4hlb3yAAM+LSLT3YJvLOjmXXscf2rQJF2+T/zCQQk
QmhMlMK5p2tplewLRG8GqlPQeXQKbfO/CCHJ/ks9Y9Rhj6B2OVgzcMHRz3KIpwjkLoHW9XvDnq65
dslbDqGKLFCRtR1X8dXkOgbmF64ZtUARARJ7Ka8ZgKTJKSSJZJ5UrMordWqaUF2pJhdHc+Gg6wFX
E4jeyyCxc2VFWIwWsiFAYZ3tLPPibTQlFw0RT/RA+6AHO56wPMpL2/8StF10XH+Pd9RNiUf7OpQh
ItfsqY/HOAcIcH4e2snzpdofj90AVwdJfe9rSwCgIyUmO79rZlU+wzttX8ijhWsYnzWvKy4mrwtc
4qA0xv7C1ct+PWzYFxy5DDsrypDhW6NoW3LjyZJRFGp4L+6xKmi0wev1watPEp0w+wz2R4tasQlq
qBMqCDLlR+umB/aYcnL7pMQ/txgoi/doqx56CLZmEqPEDHS/lkEsiZUI70NVCpEtsGf9dyq/LGmY
dn4+9m2A66dBp9SxE7jUqFwgs4DYoG8GnsTeLX6okLygC4cgfWs+5cqSro5IntnaA0gDBOfx0Gfb
pmFZ2L64j81Gf1YHXhilxSXHnx6chp6CnafjOOR1DycyP/EqA+iMXVUt/dky9Kx7CbV+V8htfx7I
A9pcAAcQehu7g0wEeC7p1wvLt6aREuFBLfurve4ZwC8yQifwwzXvyylVkTBsHheEWWmXlOXMwgFK
hU6AKITmqXL+iaOP3DGJSsZv7VuL9sQY3loEOdWlrzmcrDtadpzBgsb7yjpNUmqWZ9eXiEuPq2pf
OyXesMmcXyxTRKxEd+vybef8ZCLARzTRBVgWtPaPyW/ePc8/1reOCk6fHox6USNOuopuGQvnw2aw
FSYZos9jDH+SJkgfstTww5lVkgTmEPibDpvuAnLSJrFoqoidhSpyj0WKiyOBNNziZ8HoBf4Q1wjY
P+iRA0R+DL5/Cpw8b9GeWv2TE+rGA3twoLYAph2SUClbFQ/r1JWai/cLW5oDsiyI0QsdenlVMynx
WO/3w2nWdXhvYGpOYTfjSap4Gg8ndZon9qkgiUtkjgNt/fozRqU4QRg6Rqg5FtH11BJlCyqGG6zk
7Ijf7GHkRSvI5UDbko3P6Oy6/L+kTJchI+u6LJS5emgx0d8nDMD7XoM6S9iDO03FWkXOcVqEFCio
mB0qrCAuwHdU7vQlz/yM1xp3Y7s5HDDzAY/PwVcEVasIvmyrGKDhvPtAs904iBUrksEp9B7wOjov
GDBOLfYlMHBUVBf6coMgtQdp1lgCTEdC4ql2ifAXn4TvCSZB9P+qxesU6TgM72rKZDwOnAPIsNFG
RFBt+kcHLXnjMqYyXIQlKB7pJOqG5SvQXTucjdYGSaPCjZa95NKLz9f8PxUMP3Tbuxer5/+LJKuO
1nCE0XQF4/wRqVGSarI3xJP3+KFpVVaLva3G0m7LORTBaf/RgUFtHB7K1ZqP33I8+zvjSGLp/yPG
C8/m68dEydwqY0ZJ43CN/vifbJB3/aHgljodb4V/uL5cljDCUDh6G0yeUq8zQSGEmyURANrENZ2t
W5ISKYKbk6lbPqZRVJ1JmSZxIh7d4OtZ49pjiMBKiJoGCuohMtXDodBdYbRPs0ZeDgqdCP9O0sJ7
fTHtBeR3myqZDHDfy+akGBSce1+MyMpLjIAtQkQVpB3DJLeLF+V1LY8SEnUK0lmaeZ85V1DNjgBI
QjtgsFeBovHgATfK9WnQAIYA4M+5pQ854l2igsqKLlI8IE/Mm+MdVvzxIrKcYMgF2vYL7N/MMS8H
Z4MQQLo6TfmRgW30EACApp55XYhk2kIY0W+t9T7+vZQpUanCbPNwKH8/ekmaMIjh5Wew7IZPqXMR
+x2LiSdt57dOFmtzulnfycfWGdKjgjsDF0+EOGmzxkoOM21ill8GPbN1yMWQO6O+eoANglJNRbwt
sTJxx7o5XHfBmXeIlxmo9EmTUyQAnZRW0MUL53XPjkWgrjU3QYpkCWahMtBS5b26b++E3TDmAjhY
Qfa9o/qmNmkLF769D4Twxht58v6cL2aiNOyKS0/KtAYzXCg5Cku+1ajc1TF1vT2OG5Xp2Vl2/uIU
w5A4O4KKu4QEc0UZXieB2tmgDYoQ5+3qSFVO5aCHrL7twsPKXkp549x0ulErcWsu2kZXEMYICiiI
RrMseYGlTWQC0yJR5+ZjLmX1KhYZOO59HkGdEM9GIs/bBV4hnpgx5SvJo9NtD3cWPl6IYDfAakgi
Hqb4WmeIUlcEoGpGTxdhIGE8oTXhFvyXjmJ8D/WhjDp6izLQ/Xc+EuocnzubzH6sVAq+FMBUFQi6
J9y9zSI3DXsVzEmwbq2KIaLmjKYs6Fj3FNzHUYXU0EiCCR8OzIBT9WZ44FlUhlhEjYdjjX4rayt8
UVSsN4YCbsQel1vOffnR8rIuya/Xpw8G07GhbUfpIqpn8gIFovR62GTn/ORpprrYc6JAqyuslg+3
F7OPWVWxBJ7gedWbH9SVFIgzl4ik9nrLV243Mvd8lzrTQCQUVKfoy53ofvJjWE+SFFOKMG9EMqkw
TrWsY6Y/aIsp8/orNezHQtUWULX4ONXMZu6uTQSt2oiTOU7Ge97tFK1miUB1EX6PUTOBfctGt1Y9
gc4J1xN7y+GLlOsibRAbnuzZ6ZF6ATOQ2OeNjXDK+eNwk1xBn/fOKCQVwo7qN1+jrFAQVl1JnWJ6
lys3M6Zjgulm8ENkVTflJyCTATOESkba9Bo/Nb9E+nVKSdjv0UI3ck34aATwVT3gx0Lq9UnfUc92
9WvAWGlAonQkhvoi+i7kG6HMsiCjThGZ28NcWMY7rHJT2vt/S4+wKneeCh1urf7DiQMtRqUk3FgL
n+RDQZdOHGrJePMNQiNFsktTpnvhQfQYy/yu6/B3Rs0mLrqTsUWhAvorV2C+OAqSrMjmUDsoJSuh
8AW/8D7UsRbP/QRWgINsztShjHDD+IbzkqJPyrPb5M35aIlCOC01DF0FlqvMAnW3hsYaA++4iuy8
TJ9S4SVf+Sm1tM3ZCrKl2k4i6Nvi6+xTq1RJwQjZm5axMKRbkD9Tm+crBKqrQtz1AVLMhdd2Jqzl
73fPXYT+jhmCQ9RBlK7fdQFy6+f65R1q+CjV8oy5+1LYJg3vX/VbGxccIJhGpyl+sm2ysJpQ7O7y
Iu+judx1Q1OUWfKU9Ng5FGtN6ShkfxF7jegRQfmzvwNIGLRvJ8hMgQ3ZrBpTk0wJhl5UfsVRpIbp
PRmaot/Vuz+wzOIp2oQkIO0RR1uOAssHlhRxifsCiN5YyMSJuO5mSaZ1y/92BjUUNTuLpHM8i6ti
w+At1fdDBbyvExa0ZjlUyPCgP8bnwQhESk/9xjOsfirB4K5dxmPFPYVEnOUeL2ietj053gLUk11u
z9Aw1DebyosYYueeibDEuFxeTGJrkBiKtaV9J1bJZzaf6/xt4YCLplO1lhxFYXZscKLCAx92sLtN
jDGJMTZcDeF3hzVlIyTfXMgX33hxLoS9xx7uRartPUe2XXmByYOCUAT0cZEPh85q2YTnJUofYCO7
Hejbe4MLce2Rlchw4U1Kn//Qd+1yOJgXYPbzCHg57BfCool9O/Z4Y5qnRDklhoOCKu5+qb0UasFp
lTocn58pLsG3Op/gSLqZLzE2Xq0o1UlFKQNYEwj9AvKCXXetlbXcQN/nEXp13EbEQZuzbxeMadzH
0Mom/lwceAYDrlAYn5X1I4RPnpqj1xa0AyDAcDRK1MY9Z/CRGdPy/+3M04WkpLywDmprz0QVTN+e
K2v8eC/T3WfFGnqyB6PB6/Ja1vVmnKkpap8EZgvglLUXFDTcKZnQeVbsFHL863Crl0EgaE1nP32m
WK/gBYDC4GCwH/2+a2is61EOAWoDesYe/2cMY2lQnL7bzQXHlNCpWt0RGNmo78d0n5gZkCyB/Ehw
TcXF52Vw9BfWTTo1hiPjgoL1PacOlsPNPzzbOtzC5oJcsRHQ/fGPMYPOJ1dbKBBc0JJI1iyvw8Eo
CGKcCgXCtoPlJLlWVhKwznvfcxWD/FZjL3uXxkhF8dzgrFPAWDHd/dYupzXxSoDn8p1vLu56hOSD
CEdVmyZ+PoZPee/dVWek+rTaVX2wXE6DLWKSmBnEWwpk6z3LIqyAhYE8GiW5Koc8EtXPmJfxf0sQ
SJjKYHC4nFzbJwMlFG9vL+/YECFb3cJlpjycJVzs78a88vwAiOfDC1uI67Ebszk2ht9mYTkE8tbW
Ad83frIF9UkII5NKQQdrDZOojuptnpt3KSx94lqGjY8MckNhtACfyja7eD6hiuSpIwI8DoPUlEGH
+2M6ZUcvHj7u8GkgakGOValIcXWKbkmgXIhKvzs0Agk5Ju6efK1u3+8k4c8E8tlOgypcrCqnlv//
agyh7dOv1y+KMWOsMTD2YvxLzGgvnjFAwT0u2HU3DuYsg3u+kXLTD9NkTyTLt87Vpug1FAuCfjJV
kAhuvylKz6qw9ut8rjaSrbfr+2PmMeefTx9yols71o6rxZJ7z3mg2diN+XgTxzkOXkJkqN3/fiAW
FKap7EuA7a+3MSHxlalBi8Nkd3Ri5qxNQjHAohhAlwO6t7BQZGOBen/wz3RriKbH7CeFYgjg/mU4
jBGYFpFhGVbWkO4qdZqaLMpX2I95E3szlhT3Tbhk94OYLbtcK+98MqGh3f30rYGjOYTH6c0f2hri
9soDUqt+1khOg3ueWB+qWsoP6mHV/TTiKKFNVNABYwhzI+32Bmg0FNjpydWBY47I1lInViipvGqi
Yw68fPje0+BcxKlY3NHzHcPUyW07QTQ7d58y02fP4Vb2ONC/GbN9NfKa05LpV7WmAF9AjFWOGyuD
3Y0TLodPqvf7/2biKPXp7SEMSvqCV6qn4r28FcrpQ39wCg/E4qvGdBBsF0FyRCZebJjuZspUL/Ls
5/wcCoRmIV5U0vz9xTfFsEtxVr65bSZUpTZoq56qdpCvroPHIqxeS+VFXJevEYUQm160m0ky/v5S
bNzK404SESjbhRpDV/kTuCzQJLsfS2NUNYKIHpaMboZkZGMSTVuX58rakJYtx4FFF227A3Wx55ND
WLCpZ7FKDCSDl4bPyOdjmf2z17ZYk5pG9Nim9iWHvcpU1LmY+02Kcu4t7IWYECyF/iP4z8FSewQH
kQDjQMctxzIsMz/h5DBTBZM8s+SVWmWIbFchewkUCAiz4gL3JuTK/M/RwHNuSZbh+yV+WIhDnq7L
j5e7Tl5npY8xkCslRNHLiRFTXlwjDegbuv1sgikZD4m5u4lT/GHU5P14hsTK3UZSc2eYSDhe/bLV
klMp8/h9OEYUyoRxL5A0QjsEzOHCjAsEZPhqeTgptvtSuq5FYbM4turc1eHCArhSCli6uYZskdIv
N75KYMF63+BsQsAAE5rE9chV9mVzOsKWAlnRwefzOM2c7KP1XEYmSt1ak0wQwHsywsUheU896fTD
/ZGOZTiVtDrlEsaUqI15TDX09LPS3EthQ3eO4zWbwH2mLrWw3AUpuSx9gNoP5VblLwBkexWBYflp
zxuGoWjeNdJulRiH1xxiXOueuOO+gxYMPLdrPWnuXmqMv7DQVHxeG4tOpffvnVocx/b2Pz35wu/M
vMfNwgGa2hiQbOYZhO3yn/sAnDywaDdpKhdVAl8RxsgkxqcU7pGn/EZ+gMFSmxN7gxeZVC2nORRi
ay0WbO8rSun0Uw4hOq5rk2PSvMF97swduShzjTkV4YhiPC1QdPc1gITYLRfa/VXH4gzsR5FCl7e0
Up7REdNs2tcI6CQCJOeLJ4BLFD/y4NgcNRS6V6c7y3kEHioNx/FIjZhH/DTpxp7jhi5AKtzGj4Iv
tv7i/tB8aTm6vTCKEuTDWuSODr0JDeDw9jP1sinl4QTbNsuCFP+chV+7xdCvlDNvHvi/Ack68X9U
tN52b6i97JO/lv2FGR8WbIGlysHCjrrljlkbR2Gh/NBOAPJqDGUUCrFEUOaMK4C6TO1jCydaOT7x
4FEYZnSglUU0H0DtMYX1RKEDkz+xcTMrTqnRNbWLhiel81o38OO8zG2PdrMMJGNjpvPMvWQhYiOZ
nkkpxSnfLNJT02k3lVUuWl7Xtlpztx8ZYatApYk4GYqNUw8USKJnEFrfqrs1fgUs+PXUgrYiy0L/
XvIpwTbyQ2BKIyiHJInWhmj1CxClPhNIBR+Q87iFsYlhFLjtbL0ROoPolS3AT6IPFR9sJ7ovALZs
4HqpJlVTUqYV+8hJCe4Ihs+Q4sj43DCxd84Q+PpifrhES2MsXqpUj+/kFUjv7AXgQ9i/FJ03DIuU
uQbA5AondsspoE8PjBYNIDu1qnRk+VTm7oEwxY3yiWDLv5dSmWGBYMUPG5e8FJKz25kLDUVpSPy+
NYPk+AxdjysgqdoJbVH0heblt03ldQ1Sj2yPZ9K5XT1KM7Wc0Yy21UvEeJwoj+mR+zP3ttV+IZv4
DR8eK425ZcYRFeuVAPXzmcHY48oR+JKRL9nf+VCOlQR4Oc+dC8bYpV585oTZLjqKnDs2/hmMaQnX
oLlyycWQC3AHxhwxlhW0CdxgagLkaJfTriFBYUlvRYo36THchngCZiQsk7DUWVLi4R7fL/Bg0SWZ
cUDfqkQhYDJEecoV367L3RHVbf9r+Uj7cWNtX5/DSbzEFXtNvYdKi6fPtU/txg3ciHJGwpVvDPRl
gjMtJW48yXTGk9ET23MJ1K525FjeaGFkY/Q6BUqlvYK1Y0NgTqN9NaF+lIHzjr/s1FrrjyiCuy2L
vJHlphKecUk2vxU8uZ0PJ4z/iwZww6Vx0c2UDsEG8+SmBLAFVN1nlztlhlUaBadgwxfLlinJc2GU
HGp7j4iAX4Hm5zlFEjK56vb2eoqrYzhAyAMLyMkyTywJ+wkfse9vaEngtXRXMBYn0nhH62OPKzQN
FX2Nkq/gcgDXlxxYDv8aWe8dn1RvHi8+H8KxSqpyfMunA0XUee6fxL0cJATzY8/Wi/BZPInvWQJE
dk3Ph+Ir2WtCHLx7nBWk7GGJeqKSm3V25hGGv8spfNbyTgCwlt3R8NNVxjGKvoJkAb63OmzyYVbI
5MBDdYKepGbbAZG2FAThAQ0Cv986c5p7GzIIIc55XCGERRanYHi4SVDZNTVEEG7UBGohA+VpMGam
dQL1SzjhqlC5y8MBaCWCczcQaKNuDdHpTuORcBpgZ/ECGtdeeP5EEveTuhfXfUV1aooCL639wU/O
eg7+oBHWDASU9eja4MKQj9rhUhJFknQsDy398fMAFxtQ6D9Uf3JgNIc5mkC1QCIlrmA6dxnXBw1n
1D9nmxv3eXDCx/hUEvE0q16eUi2GEDudLyVAaDbC9qXiWtS+gKQAwrw79zAZm+e96zY8V0QHGVjO
QZagxga9xwhl9Lh2sVtBDn0HelpWgH7I97rLAjrt8rlVMQii+4s5uP5bovOjkOS289q+fZyyVgqT
e2HFcN48/3b2C/7OuRfdkRbUskAK14IOe9+ki3haI2NVblt1Jjw3l/nJO+5sB918Nyb+Raty+J65
Xt6FVShiQkxbkjwFDFJpHkBuZt6ErRLZivH0wFpzz9IYrXmcmvUx1xSRCIi1Q+OSnCa/X2sdCbsn
hepmUPVxYGXg7TEpDthmToAHJvYRKXJUWRic1Omaxerpc3jxdBbrW+SvW4zwZyr/TjCwXF1PAf1T
ohWPqeBtwL1SLgd2mQDbCfbCUKuTPcquXpsxQAcgNoVjryKdCmFnd1xn4g895Ycle9k57FD7R/kN
gGQJ6rsqqQD5VlyTqAtXTxiUDi81o4NpidkaOPlxuTFtD6g+7UpOMtbnpGqPTYI64tMbqFyydCqi
a6PV/Zg7k85U9Wdl8SzS4VM8UZHOre3tEAr1oZWhngjHU/cNNd4/za9onkCUG26zEnGadKkJ8rEs
fOrT++mGSJ0/v3XB0q/2Tn8I9OLnsA4bs5tq7J6UKkVzYrPsjVec/2clC7EvUGA0ZTJZQwzyA3Xl
gXJMS7ql9HwKKxo9zGrU479msM7jda7dqqfeqivsL0V6oPpzgjqoH61+W3tFGIevhoficzW9AsRo
w49HDGBs35G5UWmKGZP7lZxRBVelD+mZ9eQr2pyXci3TCWGCpFIkJXsBMJceSbKECNbz1g8kndsw
eLOnPZfS56ezQVZvyBjfusgO/5txhCQifm8f7pa2xWYhHMNfoEyN4oyUi3GEbX+ZzISWx+W2bSkE
rloRENGfvaLvCZWiKW5aZRJ+eqtPbkVLwHS1R8XIHLf1T2frb94H3eIInPsJPPVi3whaQ0a3hnRO
kUdszVuX451UgGr1XdMjQIIxs28Wna9rNuJ3UNwS7TH+40gWyuL4V4JoIcRL16UFU+kIkGqxzEsy
qZms091LynzjZqSi+rDYmUR1otm6WnO3yh3E1eL+0QNvlAEG9MQVeAVm99w1ra0kL7lT5S+Q5Je2
UUxbKNktGO7Lbig9g/AXQpHpAFGZXCir4Xdy26RgM1bsD6RT+C+fe7I9JZuq/bKCgutJtIS3KLk2
ggz+3G5LTB3a9MydXRPtNJsbP5Wu4OY0zcwUoJP9j9OVoLGQLWvtxTX4E01yqBCBxVyw3L722dAF
6NRDMBmIKG3WX3ntk4K7Cuv43vXmSIjg6Zg0jIitrPt13KVQpsFqWgTB89Hqxghnvn5dbHHyXO/Q
rUGXM0SDA4/pZ9o4MpoXU3SGkoItIddGOFYApg7PkuEr7cipHtje8BS1+GZiuWzoSO58Tke3sW8v
2WTh9JRaB/mHWJXPJhiKHBTrvVeMMqjzmKBpCF67qlJXe7mOu+FbDZ5eEgE0RjJnZd0B2IMI/lTL
WI4byWxEYLFJf+MTXzCbMBdHbHD+GskYhH/sG/8D4dqoZosfTk27KHGEFFkgbyj3fT/As9Y5lhpd
Xv+B/s5HCt7FOb+FueyMSgTHf9bZtpynmVfxLhlZkfKIYvFHQY64KcbVmCZLGISrOv4+rg1l6c5t
kJupUGQR9Ceu8i3wgTEXH1c77eSFPWwerJKWlum/YcIGNuAv/W/8IfgOW5ltA4MQsNf/8SB9lEYg
1jg1rjGIIxycNFe8DE7Un80QamVt3kssEpMV3BWRgV22hEn0XlSdQoLmWjlmTuwDsI0ByX2EXPip
N9UXHDKhXW6+cVdTKqtHKhfjyTv+f4UzEsURX+EVP7U1Kknh+/PLUMoPBzpVI3JIWXkvaqafab8X
7DtJCcKFo4Y0yrB8ibEKSgq84mksCOV+l0KfEGAwhSTzGsWWAFqrObsx3fGFXSftC+45xLHVL0OG
IzXIzZ6cYoJO6ctaY62I9iYGKvrOAcLivQIHPxbTOMtMkwCMHcXkQ3xYSOASDgKmQo7ciZaXr/O/
qNQIUOZ9Z3eSbTYvPawLFOE9Czb/did8UwntNjMSfVo022rHDyoUDVBTANWLScV6K64AFaYstCb2
LInan7iKL15my2kp3jNVYSTpZJjWURlXcU0kbVAwKdU6weZ19Auz05fzK6kKNyO4a535f9EqMwQo
F3oTGzPdrzC7RSFqanH190mHi+qR+lsxp3R3fY5s/3dZ74P2W9zk3BQlq5od3YWUn+mWH4fcdEGQ
rvl66FW2eIfuhoUxH00Yo4Ybun2kswDU4EIdRg/FXH3FyBksCb9RShIASP3xdIdFWzNLQXXi24+I
PPgFHP11nn12NywqG1Iknjn9/Hu0GBva/nQmgojoMyEags4IacZqp4xvS+cZ9DdnRsYtSTFzZ2pp
94FQJ3hH7uZlfzKmXqci6GD2BBO4okSUu72/p5msyCxR51djv4AHvHLFz4hEDXUKR47NJM6qdB5M
6jXm2eM/G1TQlrBMcoLGjTk5wqbn1uAk8nywL/u34oe4MWHPMUXlc0pqRKeKlF0bPAjkl5mq//2F
nnKF+4WsUBb6uuIAiU+M76s5PgIPObNsVsZbVTyjJfYKltYece0OV5kpL7geMJSaT5B2L6qG2AyC
soBQAPzSDnSQav+tjXmC+R+vieN/pi/16d3Aa9LxKlcm/xhAe/Kp5hnAqBgU8y/ElcM4qKk3nhNL
NKSKYIFP12q7o3lXY+OAuTyagawVbqR5VcH7c5QKKY7RDoGeVtvmY8UzmEel3qSrAMZNoeY4QmSk
zh/YOC9wiayPlx0fh9VbkF5pqkPZVNoWv7yqHRp5R+ZmoBhhLmnYjojhZTJJs5OJxndMouzZKe3K
/Airsk/bHCGyJ9pznovuhaH+m1sYq09eNyHRK3G16BPKwo9/OPQIjfkxyKS5d6D5XAWMwKBQiPdG
3w0BRBMTjZLzqAlbPG1c9SysHlfqzETlWVxXjyhYcLUhxAbIJNGuQzVnD0UHUDt8QQ+iyJZRc1zb
5YOIcZ0ZnbFbr9L+JhZpZv3UvQRSJTFzoR8svqoEkFqD61Mk/kW7+uUbiH+ymJpOStMstWT7iLg2
GeW7Z8T+BnVBa4WI3Td8hqlsB4cYL1sf+fZ9G3WW1RdkQ7n8//BuU+MDx6qT2OEs6sA/FX4iFgBu
eLxzs8OoAHrwRfiISzMoXEWh1s2yn/GPVVt6M+zVVIQW1hzeoHtdggK4Ril+lLFfOgFixQCEXNOI
RQaR/FXGHu4RUhiNIqjXBBug9X2lhMqkn7qGkxvkjUEnCnF58mMQgWaeFXZAJXsCnzyoqJP47sbp
a2ROVlv1Y1H83O/4M2faXpVeFADv07hyt3RnGJ95VAGvkjhhpGSH0Wqn4UFIXBvcbLjOwCFps9QY
b41KaPUaipen/BJIwlhUl3xiuhlbTpahoLwXjxMRYGS7l2Okzr1ZFXnFPbf9mmEb8z6wJfSNIL9c
lC4KszQk97Lol6tpSUc5MRSlydbDn8B1XYDjyuIbQ3xgkW33FKRuYwamRpEQ8oFvycj5FcT6Sy83
xfi4YsqBBtTbmF9W6l5rHqHwIJSvlC7+YSkdKMr3rGxcFOmgYkDC9x0fqUQH19hR/TNgTIM72pBl
6lyeM8MnxVFk4c10Hq2VJqfwOAJw6Xz0uuGY0KNuoiw601XyOrtWVYcrOrP+u2RymTX5CUhHce1M
+3rYcE6va5eAhyYEp93Ea3VpShJ+LCS1Ow7ClsSw6MlaZ7vgfqOY1NQIb2a0nxdokFiBYsW3Pace
764I/RCLjCOr5Ih3+cfdlGjN0gXJEfXtIV7vXFoIlkLm1O8ZLTwhTJf7Y1lwRi+Ljgkys7pZSKJb
NafJvGe0gJ65U3X2/kB1xIctonzFXAGMw3BHpGv3A1tTONFzfCjyJDKA0MarWhEEiofn2+S3sduO
q4YlPTjZEChro6qwvKpS6SukemoM4MezPJ/sLrqfSVO2SbFivHMZR+nuII8NCWG7mCgOQxY6b+oc
ZqkRPlVXu1TFoVEaEUueBq7Wqsx8Ewg7zbALh3UfVeRO9bZcVzPC44FX+yZKbByegt7UZTjJckHt
Fut4muEtxYEZbavBK0mbKYt6pGiLn0j4IpW6aoWxRu2xGs8s/DsSQhQReSJEXbW8KGTc/lfCMgX3
2lUpxlPNkwBAZlhCZAkbjvw9mGdEbJuEXH/BiiNE0vGHFASX78p2+9HAoqPFEPf1FG3Z1vH3HQji
p+IP+cQwgF4BA23yxQOiQiCUbTQqbwGHEI7dVM9zM/fEiXoNpdvJG6kPDTuE2x+RPBsTALxFy060
3BeVjJf86MerEx3WmJmjgYSi8TvzLq+6KcfTve6n2bFGCKrcJdcY6RbJO3LMHR1KopORaoSBQCcE
kvm0dnTjbG2r9bu3AhokEW1NBz2n+Z37FBmqUzWtSYbAdYpQV2m7zrSY2M+3xu4Oe7WvpVFW7Z73
dxhP2lxBbMhBUWUD2x9xDv/rQ9+9B4ZjOysOOhEGRKQ1GQhZnRr5gpdIVpt00Oh3Qb/58EthrtkG
vrYk+yFc4/YAr9mzeP4rZjK8LtDe14wBjrVV43iWZnWjgBUD8whUMHqo27YTGpMNAlEoSQECqZaG
lLDk3JXroAWl+XLOS/Epb65NMFKJRIFWoJEmgFtkjFoauYS5ScxnlMzjKi+sl7O8jvokeu2CO0iu
io514n0RAlKPQNooak5Aw0sxS8tMlILVVYCQJGx+WWhuPUJVpQLJ0Tj96a+OvuDUd78W1UtZI9/l
fw2BgFWQJ0g9LkL/QQ0RR1yr46PzGClwitiv8frIdbkH6vD6L7aiJHaWgztzAqcrtRjLWl39lMSY
sMoVlPZvq7vC5qxQyPY0QgGc7+pY1GLPxe7nVKbI32x+RM7RkM3j0FlUB7LcOMcNKGhzdyUmcgj9
QRLc3JODoLzxv4FuFwZ6m0eRaz8+SYrwSU3NdPFxBw7G3Z/hN+7heAQare38o5GMmSJ+b4ZfXvIa
NnPgjtwLHOAk3+LHvait8BBLDgkbYUASk3PPYkT9lnZhom3rRzUxVKkWnqvOfu/RkOIW1QjZUYFj
cvOSgcxwlUARUrbN/pXYw6tHWn0WAPG7oTPCmuU3f202wORZ4zLwLkYCbnBXJnHfdbhSZm12yDAo
0F5UGRrWeaSczdgAvaPoCInX0qmu2yIlEqG8EyTvdJpQM7FgPwD9C7RSeEwEcZMDIEXDqFscoRbq
KgcmJs1xKrGG9Ig4NCBEnBALJ0xMjqKYg0jF3BxtUXp+INsh3rHkYY9DwoqLj685T/zJouBt7KgL
HhbPk9kCCN9QJXvqWNTaLU+Y+yhgw0hTyxf6l163gAvATlCu2cEz3+OEItCTSg4Mny+9++06cvGy
myeHCh4Qo3TAc8pQlaL1dvCO66A+KUqkbvHNFO4S1aDuEzDVz92ZnZHM4akWQveZ6z84BsTMjv18
G29TQ7LyezqZrihmO1A2iQ1cgWKw+nUtt3aOQOPrJfUTsKdWbcr+Q4yPJ9YjOM0VCvPSpTPfn2m7
vZuc29wn+j1SaitQtr0qo76VtCsF9aFbAKnO10kk7wFDqtISyqdNtdReEAE24lZ5b2jgnHfVbSmG
xR5PKat2nR4+cyFiMwzSBFS11V50wv4Z4Fk3VdidSHi+t+Xzy/+4F0Pq3Z4694DSnmiThJTIhtJ5
6ZopQKhBWwkDKX6uqhxm1Y1ESVTgXPC3m1Y3YGQ3ribFOCZMFh76VepIIXJ/X+usALxwiz+8Dp/I
Qvk43Qqo5biKP1k5eXeS9hRY7NSmUiL2AM7kp+Jlp//oSPaNT1xrU73l3OWOtjcsmcVFakuaJSC2
o21idEt5WjIB4eJ7A+DVVTgb+Icsfv7i5NwLwDs+nfG86BIPLZ0v9xFWYLug1QHpJMvwW/K8lhec
JuG7TO+1Vcr7nUyT3BfOoHovAL+StDoC/ZyMft296iMuCSTrl+FIXYwbBBglDZvimEy2cPFTzDo8
NDfo6U/ZNNBrCUQJa/dU9KOlmwEYZGp8AN8viRu9p46sZZ81inTuQ347HLFbYthbziLPZR2TbF+s
/YrfgRPkzj8xiEFiEiPTc0JJkwyTM7zXLmffepPHQnYAQ5jeXzL5PZ2C6ZpojIVHXDKptpFnIAgs
M3YrDDuFqPLCmXSAl4Tu02f1FZePOlapH+uKfRh1QAhPNive/37x6Qj/vjAFHhzYuj7njQtO/x5H
IOECcPJxHN+tackdd7Yf+rxVO2wCSeDJscK+lSmXh2KYJp48OxhXK+K3BMHO7DuDqIi9MjsrHmYx
FL5imH+iLV6BX4K+rHLjdkZdZXzi/Av9alqN4IiEbsGqmdDQpL/o66ESrYBZaqWVkC8WYuHRvu8T
perfGsY5hAuTanrKaVYcn9iIFxm+/VbVaFbU0CGmyQkG5VuS/rSjx59Jy9PWqmZ5utyD+RlhUyJW
8JRVruObbpTLLNSfJr2B3C8zACpOZC037KGYvj8JhZdJOIjM9sx4VdV4WVBDChRxt3TqLDh+NBWd
KnuikYWmkG7n+VxC2YSD3QU8f0VjkPf3w3C28UfgK8F4Gb4WStORsrFJFE5CjkxgDp4EnrYvSIA9
BtQcRo+IrG4QtWu1gUAuHoRq5P1GiPtQXP11lGLYLTolo9y0v3OM/PT/yB8uJlPtEJa3ywlNIUa4
DZESOWUPOiTfRw8mI6z8xEFaWNgxAk2qKX3X/2huB7IJLbcsU8Uda1FN5cAPhcP3qY02o7T2K5Ow
VtHCipCS/d3EMjFH58fqnLJvikVNcVFiuC580SRrUv4H0W9EnLT5kFeT1je+Af8lwW/s5x6pSJUx
gSQOtoOmYBbcX4NdiJhs46i0f7ONcsOOTAkd6PxLV1BYzKqbTWoQSqW3jXITiJX8wZ51Wx8vV5Xu
OGgFjJ1ZYU6QysStqwzP5ofSNZ0JVm8zBWj/Qo7imiQCktkqQ/DPuHSUq4WWuO7XSTx/Z8cHNbpS
gf49NmisSgq3lM59SfO3y1mg56Jftww4jynqOB3d78D7VksPtGp/1MqTMs2xweYaeIPu7uyI/YV0
82C73jG1wLe8FJQgaYqvKVgbr0HpqU0SA/GylGiFyR3AtIvHhJ5FRZksWwIrBxbdKXTzC0hqAd9D
3I/trJAIKpXUFyhfuOOphQ+pywBTkI6ifpKghv5j2rQwNRgapZLLPqDNj93cfX+WINKs+q0gUuEh
I7w7Hd1Z9bI5mMsHvzw/iyttHdJySedn8a4yKAJgZ+ZS2Q7vuqcstT142dlz8vbeaUu1TLGdXOTv
ciwAtzzyxMkEMaVXHK6hsQppH5RJ2WQqE4pOZXdQtDqx+JVyhqMkEA/TqaZzsyM7w7EX7F0FvG2F
GpWsUZLx99P2nq/NJQUDpH1ZDnnOLsoBJCBbY3k3bCzcWpGyXODJaBXVvIhDVG70HHY4Jjs19riQ
WfkZKwwOzb21jTEywh/YlXsmgKpHLqRnav7YwL1TcWggw/ErN+PXvPiH/gW/hyZ1AndTmL5CeLOi
kPhXmGRe+nzoTV1VmLPlVAPDdyYCgaHOJ6ezJPbFd9/JHFL1695zNAKh5/l7gqT1OROp8G85WZcn
pwmILiggTCvoI40jOHo011ar50UaGkY3PogdQmkK29sIw3UiNPxT61tVYjWaKZVa1gNpDzr3/ggb
OetFVMnbwWPtqKUSB07KUg/IFwmKffyMb5D4UZXlLSl1gqeMWBkB2e4ETWevhjYiNtJ1WhU0sjwP
l7H27IQo76ypWKl+aeToZBwL1nGdU0ZTldLqWLvjYE9uJE6uIc6U1B6zMIFUiZ8V08jDqA2c9JNv
r0YM3Shqae3wFaXJLZRxhdNBG3LuqSIYM7Hoq6RxMHfE+lVvxPHPphs1XfpNVVpfp3+Qrm5ncPOP
6kh4Vk7JbtM9Q5dtBPV29d5V9o3mhKTSM1eRlwgnnEZN7enncCxrgayPerM+Q57HKrBEBxdXQfwG
AsvP9Q2DG/dfCZ5tHYia0qX2XDg4+ONnGwt8KQNBXLjY9tOr0xruxL9pSSSLy6Fn68aMRh9bN8yK
7o1BsljmqxoJvkoZ6e1XnSvGMw62Tx4gLzPPhvJBsest3uJHFBy7smRMrzpjnSxuchDvAun+OAr0
OwThhvq5vcR2pw826ZgN8xtaRoNCI13ah/dj0/sv+jutufmyQuXL4JRXsonY2kM7YU//YwwBAkax
XuAplb/bZXkLUy0hjZSOk+kmCJcRKnWkdeqNH0AREhpw30G+QkLrfR1jQW/rBNYYccAmDP/iwNfC
jSyMkWhBka3MXhYEzca2d0F7t+6lSnt/x3G+EfKXZn4XnzSaAUCFU24To5CUG6dUl3Z1rQ64LdKI
qZHvr/Y+O8XoN4PYXcuJ3h4TCRDNFWvWEMDEY67Tf+pREJmu0bS3N+MALug8TXhrX391TbX4nY9C
svFkjXZ3Ko5e/Y0yUaaNNTsaG1ypPth4hhORYYaF/kDW+wxVFrkAE4HWQjxqg5uhIv6Kzhe1cHiL
BlxRuJL8BLhFf7nA0t8ovtrASm1Un1VZ0lqBUp0Nj09Bz0Sn3haZiePk52S2odd02lfAo+KUq2C7
mvDxnl9xDMzzwWwRmkn8ArMaj3VY761sohR5hBNFIgPLUAloG86rVRIJWXbfud+znx19QDdLDHp/
ADeYNElKb3UNiFFV+4atKt/xLpeqole+K83BhJb+LZB1sCSZG4xWGWrVDEDer78h6eyihDZW5Lva
BcSS3IDicrAqx/K9bCZqXKxWKvRIYIh/8zuaL/5rfCyWmkvekmQN2UuISnhIngLUMAnAr23vaDEX
8lYfV2dWzDrue4PbvoI1eQYkalR1PXByLqW+69wNOgZHt1RXGz4k6pejEIvfjtRLWjpiavPrwZmx
q1KXi9VrpgIOMw8oACnYA1f3P3cDKduxvs6b2RmwFnXJjZzBvJcLYxL16wADARxjnidTTDxzVrnj
Owne7WTAuS7CpI3r9h0Vri+FGH8AM4lGpb5jlB59koQi4RJUtHQadsw3l6LIzXiJ07CLNJrevJXh
nNt9UfnKgRbH+RnWl20d0XOlooc3EBL67H2M3rQa2fOoj26+pjvw0uJUBf3UAhAV+07bIhy8RJHW
aIOqPkCDKKqIcbzCdmuW16VsW4m2RwIEKDMfP6c6DPHge59Fjm9v4iBIP9T/TRh0otLnw2vf9KjA
Bo82ybvDQaune2G6W2csoPfQdMpnlEvN7uaISYsZzGoVwZWAQQTVrkhnjNdDaWxkgBnCcUNamhJ+
25MRUEat34hH0YLlvvN7LCs6gipVd5raV36rhGPL6LGmuxTmFk3Fo0C7YIyfTpzX4C+b8XoViQuD
cTnFaMaiUe4xaserD/AdeYWdXKbIZxzMXsyIhqvXj5Voi76YoGOOlyyvyts8ByBcdgIbZ3U2oTnW
vZ3Xxr2yDAyOHZxPQHeS8+sRC5FF4QmpqwGnN1DOOWSRonBPDMQ4Miw4YdMgFSPABG7IWjOy2MMr
fn68rJITW0eBwF3I69XaceAquWeCatoZUsc1k+iZkXO9F/ZpXVtY5koyqXLkpJTXAGnNuzS2GPNa
A+mDfPebIemCYIh8tr5kiytwHOA/UeWYUQ36UhPMPMnlyaZScQ6+lIaqOvcEwwFFXj98hPpSvIEm
tWxfdbLtkRiNb6SWAuZBRKksUZDfxSVJsuUzJGC85uc4JMcJ8WSsvNImF2lsVgWM+vlrh5cusXr8
WX+JtYcuI0DqMfwQ6kbSG9RBiuSLumnLSgK2/sBitRKQRJWbs36bPBhIkL4dwZlCiC8TGDlaK8M0
h7pZKmiBL8I9wSPjkdaIn0gI7Kbl+UygdbTCSrha7Wo3DmJ39d43E76rCxRgnZuq7rvGyqWyTUUw
HS/cpreaSxiKIUkYv/WR+CtuUFn3eVxjodFrIDNU4jK+vsTXuU7WslGmm0qmB0Zn3E9tR+FpWsOm
FDzUsDK8i84FEh0C1qaSAbn7bhjmbqOvOOlX0sRyUqL84ALBWYZ55fataGsHP3C1X/i38K1OwTZL
sz1slDH3NuTyw0IxwqivmqoB3RMS6Mp9Ka8TA8B+7BWyFoSej7rF+6DYuIAFZjPLxHQrM2rQX9/1
pEQmboKfd2ZTBqYBNmrtsBM6WsxI/sSGdeKyfqdM0usUuBPh6o1PjPQK5czgL+TZdNXVS3H/BiSR
VW0+NX9I2j6ymUw7nlffAM5THrKjloKgV9u1EZLw7+RZ5S+hzrFFP4P9RKaSZgAGkAyB6kGO2JIo
37OcHUdpAPZdtz5L272dVOIBTepFTlDqiEhm00sTP4HKHFDNmUpnfbVZ7302TdyRWLBcxIZKnnND
WdxiP37utLTa56ZjJCqtFLuN1WScQLmWTeWqhOOb3taMS0Fz4o/+/NIkOCRNyjNuslxCyeKxxwQ1
lAAOupRRRrgjMXzBkhUrdj/tPY/xzIQu472szLK22kmosEzTFfiumq7X9Ynhm/MbdpH/uh5ttRTC
m/tA37fZrFdQGyThPvfhOM4JuMRwlnNxAyuUEcfAeff/Fn1BUoFzdhstRbP2sjz867O0AZTe4sR5
Q2ah+ezbER/uI5J+4Im26L9Jd/t0tNarE/jWlSRy3xbc8dJDL+eKt7qNDKgYUwVLVoLsBH3X/OLl
P53XZbfUx27tDEfAOQnAnLaffHL2cB1MgsRdZpe5B2Y2wL5f2tml1DdyRc8jYApvpWvolme4wz/7
qDQMGHWipIrrI8wWQFElphpToNMdUMA1CI3bDie3zK91EB+2t7e4jnutHjZKM4iwU/zRWGQmv9L7
8ifPlQFWQQIPTpKBWTw2BKX/+itn3TJ/r9slCb0HyOpwp9QpQ9lpMC32r4kltWvU6/l3bvrLuYkr
KYnXYVZh7dpD6SeKhxBLQoYAQJM6sF0KlTZB+ty9IVo60fSIc5aNkXffM77wdMoJ2fpmxVxXxtv5
Z7/jkvWkfr/jo5L2cdEL89V8lOruG4KWNP6nefX7qv7lhPlVu27frEjl7e8MmQ/3Zn9DCH/+R2Gs
53Y80tOmbCFouL70nz/y1bt8wOyw19Qq8r7A23syr/IrZKSFjKWlsa3pVVIB9TyDERQUjo/eRzHS
NSw23F5muv5rtRs70UtIVte0iBG+gDY+f7nYI7N1koMJMcgg9fjewFQm3iTeFdGY2vnWnvaxK7wt
Q8IWJsbBuqGtnqAfOHK+tjE3bjQm6w7uB/MssYUPAupVpcaK9muQYZ9RiPqm2GN5wltTZBg8umg7
or0K5mcEr8+wUx4jdZQHfkVNdtEKu4stnwOrFoM+IQbmmsSBUjbSa1+o/GoIcZcbdeE/xwlSZcde
4DNx0XXaBZYn753m3KUtKVA/A7DWJ770qVj5UpJ8ODNZh0RukqB+XsulTGx6U4j1edPSh2TYkStn
ORn3gIppZHWZ79ts8Kb+HQsQfWAJRNhm0OFk03/UJWwHqfZsuPIbU0LPY3kUpB4608mU859QMl3K
iD7f3qHQPq2Rj1rJSvoCTRNA/4yKXga3ig4aGDH8vZJxdw8fSblnaMFC2pcQRkYGg2XnTV3HE40h
TmZYo5jVA30lzJN84N5HeRZoaZiVvRdXpTAoIe91uieQMWao0gRrQQQnZfVT/YCiaxJPkIOKFico
FrmaTNjMsTqpu5Qrs9CtfyrPIQkyO/lBLTTmYNYePlBC+YiczSi/p2Luhcv+ONbJ/nyPw6HrfUOd
vLZNDLWyokdh2o0fHNB1vTGLEy0dJ8nK2IrfoTBlhZDJy5V6gcrPtQmNJ5+DWzQqLqX0GD6JqKf7
ahcdnMi+MHEx6zYvRUhPIYukWzIu+V+alVhNOQDxvKm2Ah1drWQzgIhfV8THhBn9F77PRz4CmgFD
omNgKmI2/MABhsBrfySKojErRL9vP4rHIIhXAj39Sz6f/HCM7QKhZBiihXey2Z1I3EwCf7qMWR29
Sp1dQGMSdLu0WT/tGTP9qupms9bEI0adHdGI/HSKJVCOW8AaUz1PErLB8TyJ5/8nytAPZZHznWLJ
inHBL4SA7l9VdAh9aZVHj5YSq3RUdQ35jPkEZGy2r9wcL2LfdqhjJS2zrAcazlA1i87lBxPr1aLC
ET/gEKXZMAf/6IXo5xAdy7nJ6waVUmqmqGNDneqYs7kCYc10sYrAR8u4GJ1MQ0RWtNcpPTYGDQTY
3KP84yNq7bcfKVE/NMSp374bd04PVRFmxZDjESvqF0i2UBkygc8lmoDLjQO7NehKK/Lr4UUGKdUA
NoQKc1ro7alYYjOTnsEYjHYt4JTWYsanYdTM/1aGbw1I4EoDWcQURmbQK5HG3Ec/AK0Hw9RRblYG
S1yT6cT0PLmLuZ6srQY7hYtOh2/VNoMY5oi+b1sV5zt82E116vkPozW8OVk+ILC5VMeHGgC/Xxuh
zMzxUwQog6+itr9t42N3w3yy43UPYSCUGzo3lpRvXP6TEIRJTUgUciXnHaXUhuzmxbyP+SemiI2K
73gB/3t091kF0jC66khixfDabvUQ3hja302V+RR6P16KqAitQSd20nTV0w73fSFihGDClR7oOfUk
zTltGwRcwV0d89iwqnDTa0pBawlCLs4uWuA1XQQtaA9Q+8pF3sVe3XbCA1LgbEXORrEOjAjjFh2T
HJtTEH8ZAWTMg0hm8Y0K+/zh02zFwMVM22Cy1iz6xMDzyAMVlcAonwuNrqLS6BrNPLu6luQd1Dfl
y3N5E28kKuKi0qlMQDge0VtKNlLSwOBitOaxMdvaBCPecIa/SAWW7jNqvJ9APGi4XehEg4vsg3SX
wmFbHkAzpk7gvq6I7SGrnqU1amL2SillfC4KT0Nt76CKUTU9GcunMbmaMiq1lw+Wt4zPkF04radY
dH8bZPDiENV+GZvR1MlX2Nb+m5rW+Qe0Vhyst4MBiDbcn9Hl3TfnefC6x+vEEuOpiK5SR0YaMieG
75jb7gAAZPYT5UAOhKG7Jmdljarv1SX9L/vKDOCwOEWfbEXdi07uY0M54gNtxeG+Nkcx8klr88DL
LtYihDImfcLLYR+wLvok3LCV2c1nO+HcDrDf/pFvsKRSSJn8vdcwiwzK0RN66Y65M6CI1n9w0sXO
TCl1KnCrp40RrwDx0TIAlpS7wH6zEDce4Zkbaj4ruQ/oO9I6C5Igl7d0Se/4dt9ZC6iKU3pMCh5x
l29lYGY4xIvbAfpAtIOnk738Wb0xc2iyksraAq+yVmKXrw7jbwQZPmHNZkVChxBJu38iWGKQ6iGZ
4YDgOUblX0hdTMNsCQeUN6/9VZorUcCSpg1K6bHfo4PJAOZgiZ1h5wRXZfnaujDpXTE4R6InpL+c
m2VlKT7+Uxbn6N46cLAH6OA5AAmRVriKoBa4GBuD5KrMQPgNrbbRjEu14qOeNUBSdyZVOLMLWIrf
TRPMvwi5VQCxcBxlgK4m9TIKxFCcqtmyBDGQv67+pZBrYp4ylPBOWrB8/YqXYIm9Qkp+vtokmsCk
PDP5qMu8vRSF6rkkiuOFrJy4g2e8EHnc2Re3SalEC33NVvXOBxooZYpLUPWqFouNtDpbne1q+XbV
x55Ry918LOfqpr2uW2sthRPzGE91WtyC/pba8ICz+/hv2U/rExTDcdodctTRtHv4ImcFH+xA7G4C
F9XGcEZELeiXn+8OwbNRmVAXrXCjtJvHLK55c0PvCuQwwd0DiAEZ5027FBqBdw4pOZZr9alSO3fu
lCBCRaP5CqNCzy7YG4R+Gd/KYFK5UNl36Nc7ILMOZeISriaEUyyOGjaoGySgewawQSftni4YrTks
JTpfORI4iS5Yhcy4rZnuZqZ+ZP4U5Epc+h5GUZPoRWkz5aprXSOzVWF1SYtYMN1jsXyiHuc/HOcS
aVhjRBoESeFTlG3ECVih10NFarJt9bXeGBnStxz+kgBM57GpRL/rf2MT091CZW7G0bjVOJkjFU3o
OCqiPB5zh8+3zALdohpkLERJGto17AjReBqQT7S7rDM5mzxG+yALWTmRCyo5ShrDD0SOkdBvocHn
TOgdhzvBl0xxQkSiotmOWQzxN8B2rnmmPwF60pR1N2DzOmsPnTiBMyJcTzPCamX6Zi6L152ZsWhm
hyGTv/3leTwqCaCdOj8B70eDVQR93SZFjCi6qb7NEUEnouyAa4+9Zr/hdd/cr77I5wNOgvo3LFJz
E2i7/7axtHPwbJ2wvkwieWq74lPRH9WEUn+7JWxn5TzofMo3T5iDqnKc9QFcD4PCLTELBzYtfzft
TUVaHxBpV9uvzT09c8VhLSeqf1H18Ld02nHIguuq6v03nW5OjVunAseHpy+mJUZ3fsTqCag6U4Bb
9pGxHF8o2VTWHmTxjMy996kmA6tQvoVSfrmI1FtN3D3bALLnwPt7Zn84vm2VmuvgPKX/dk+mXj0U
GjQKJT5fC9Vix9fN9S4KYb4afWDrvrVUgFRvqKWtYfM1XQIQp+auEersM+grc8zpkqYcmAZiSTlG
qwLpNyeSFZ+/bfF47nCJXWllHHuz70DA+2OqVs9yB8nupODKXRsvCVj3vE06eVM6/upRuz6pLe9J
XUv9AG9W56Zv1GLQvswJSM2HRKo6/+HczJv572E4+TmRqDNQfjRJkZ2BMuc4FUNF0bkppSLTLaMM
hKGjf7URtz0GvhTEZrr4MPjGnrk0N1RQYbxLofVTQmVjAmWgE68FEcORt2P24xpaAI7pPbl45kHu
ayqrWV9D08H0s3GL7xBvgjpxtH40w+o4uHw+JYhZtKj4LrrJlmqw1lz+dDWcfpd3Y/X1RgAQSrzM
XBJAU83UKJfrFg/VbwYkDVSH77rQkmuMHdXEs7PkhMY7PT5RIYrQ/hvscAmnzKg3SCI5+H4iImuJ
BBrO44CAJ2hCdrz0bRyfzumTNVd8cCCftsM4YdAA2uLRHCoCmSG5f9czmrI245zxlk6BCxPdfLjC
sVJXhlImFnve/nrDkt3KSGwWTJkJ1ZWMYID+bv/tCB3cGrdckSEdDQMZXEt7u2e+3fcKodWG1EfX
rTLXL3QiiM/s1CxSRdtVPudrLdNig5WLN9RDlcLNHxTfA4q6h9Fu0GhgM881fSnjmnoDPpkXZSRY
fBQidjJ98VKZRwa/cBlD7tHJ36zg5rBJoGr20O53j8ytRRVKuuoqA+BDVTZ6sTJRbnw+neXnNdld
rpoTfeZljLfu8iPSktBgKMtVU5yZfbfhvcoFgRuSiF+8Ipog2zVfbzhgz9IUeQOV+28ZvRDRlLoY
MhyDJIP9KWMPFM+Fk1mwSk77+Vz9pKNBKN7IsKfHftW/bt3r9D7GpYKfOw1v2K1hqGCOlGDRcWJ0
sb80J44IJJhOHJ93+gLLGd3QJMEFCygownXeBlK11yhoSlxraEMLbwJR9HEL9vA1zCccJwNN1GYS
mlXNZPvniRS0fFNs6YXaZBC6iRIRNF7fWF0N0czUXBNii/z2YEVl6H0k5bwYwxtvm5mvnapn7khv
ANxddeXqszS9sLr59NEO1OfVkY0Obf4m8+LJVfYByzdL8mUKUFH+Rd8bnNTqYD15hPcHOgBX8gUR
hu3fFTfQ47m9XN3mBb6ALPezazDwAKEEkV6ZK8HYrt/kZMEdImBjd4eOYR9R75Ja2hqpkhqdnNI8
WnwCFTb4ZZcSYOHHpvVxMctA2yXrO9CCnwEJfrlN69xUseLxgmXKlfA4Ym4zbDEeWWsAb9KpPxke
iNevPuRlod5xgcEzD3xB2nn+xOUaDO3yqtz3Rln/xkj4mbpcMC5NpWs395IbE91Eo4hP4LJ/lU6s
O3Inh4x4XLBUMLqiVmVMplAqwPdGenAnLOtL1J7dk/kxM6eibR5QT50vnvhasJmvwVvQLVoD3lS0
Yftz2CivdxDdwK7iNhqWTvOsYhUJxWza1UOCWH9xAF8H4MwwoCRA0aqg3Bc8Nb++uFqVLk9Xpv3o
q7Exz7k5moT+96uAbXt3zY3jqMd8asv2EhvGc/zdgJm8hrGwYNYkYZD/QeJdb5EZ6b80x2jIz09/
XMIq49LdrmMIARiY0X9Cj4qD52XJaapu621bx8fYzV6b1pQzfR/STZLDA6qaCA8DWxdOywzCCOCp
5qjBofEMNJgArEEwQ87j0RTik8V5Lnjxt60FhrFbd5dFHlMcb6mT5yeB5ANk7bPuEXk92QDF0mXC
TiicupWCuw/in64soty2YU+BtmOqHO5WgPW5/D7EKmoj89nELfDsSAYHCykZLLS/K+47Vsdkl9oU
1p4kaWbCkf1faiKIt5R2JoYZCkwPpfYAiJJqOrmcEw+rnNS3l1DWWQVnqa9k+Z2hjIcQsOiZSuod
YwEWCV9F4IfMNUdirwhAI276ekQQrerDMQEo85WCXWTqa4oj1CgvcK3RpBmsCZ0zB7O6GGRTif1c
r+prLojDvcUmV7WnD64kdDLXN42q5QVa/vKeCPH2JSWm3Iftumsg2FqhRqGm8+meQ2TxykpS+3HC
bbJJbmMPC352ac6zzLnQzyeQTZolHmXW8S405K9zO/xpWfzTlN2ytXRdw6KircNqHg72j91lH07P
RlN6hAP59dGygktZDs9wuMDSYxZ+lOcFAjljNpsRY8buV06vP2rEAAMdTrFkdp8gNBaWS0DVRsQ4
8heZPfJjJ1Xm58wVjr+J28gJZmUszpRRiEZ01CvGbZHNgqo/pMvKHG+6KDwF81vsXs+2erJfXg/0
HNCFVqvgZ3EyVH8GdW6qyakICZVSfbBlycLKbdVMLn7bJnqGD89qg4vCLpTypQxX65QoJQ084MUr
GDmlZ0wHGNomIr3BwU6W0Iu4a7NmYkmuTq/2C2iOI48L9FyTHrMtfEnqPAjVbxyvs5jz76jXmbZT
tM7a1/fcFSH8YYgT8EWSFEuZQO8+HBfsW3VUNfSc/HZlJMqOUYoP+zCcBbmu3yQ+MeKMtvCPKlWu
HgjUw426M3MAjQo61KPKhWd6WXIdbAv8LY9Q+3Ug7CRLubehUe+tPLiIY5r7UhLdlSoEmpnuFLUQ
FJGyPhPxtqSzHfuctfbt0tHqmFQKWWt9CyW16Oau3+nY3aQUzaE1pPRdlgQqnwiQZ+7FIy5jT4ej
ye5f2oKI3YQAIs/FP6QfyLlLQGSvQj1G559GX/bKTpW44xfSaRxAYtJUg2vRPIallPRiW8rJJtrX
JYPH38g4EI3zTMuWcCiT12/4gfQ4cEiBvD7wsc2c4a4EVZwkRqEdc/JEkVxqG8uobCBucSE44vkE
BCs1M0zzi8DLlCv60KYvemhXNzgDVJVnQmw934etKVpTuU7S5IFOsZ3rn6M2BJYIQbzNtP7otJA/
3nSEwWBk34GL9G9DtrKB9v1SY1ZO6f8ihIYPfSnkJh1r3ibXnjvNDSkDld2xUObl3VabXMCKAV07
rpa9mEFS0Z/kGWrvr/XjjH7Zzontu1tmh2KNDio97gBz07ZuwK6pCWrM0HlGj/euiwkvHLjokv61
x7kovJ1mW7SVwz/DLwLS3OSuIsyQkEhf3wTwfrR/kj2ioI6jp0n+NRXYzOJ9DOVWKw5iwz0nJVzz
ipqLA7JymXRbwWk4GYvfjsltEIOZ8yKmMDJCJ4iYlPoA4HlBb9dbExWc2WK12NXJiR2o8lNIOr5S
q/OAsX0NskYTMI1TCuz6sWPnDBaqsURIkJSVyYyX4Dvr7yaH0F/Rc7RIrcm0yDoxMk269FuAdEau
1QYtg1NiexrQzQdeRR8QxHDzlTyuJd6bHWIW5+5dF6CbzrscOg5vRYgwDFfYHGl31BIYsagu6OEg
bOLR4GQ1diXfkSkdGSILV35/Q6bI2G4zuz9DMbMSlW42hBolN1ybRYxlJiQRoYI0TbCaZ5tgyApM
BLKZ4XN6RtuAmx4clIfsDnAeiRwbupJwl4+CQeVAZR3k1O9KviSkXMVHpi3FZaezTjBEyxL3YGhE
gGeqTYmGGz+lCj009qov0l0htqqbaAUrvpZuPwUg9zbIPUsNZg9HwE69w4VrUxmeAuMuvOpnwk+U
ZdVRO7FK7p56RYC5+FCs0gcxP3kysofni+KZXrNhQn0o73PkAaQ8A4GnBr5+JXFPhnO+s5flhO5U
GngSB+NTsBgh8OtmsxoFCYVSQ30TXs7PBoqPJ3d+LWPiK/nx3s8ArwHWcBN0ictu6vVOADZqw6r8
8YZkAmoNq+rcdryPdVprkTDlz+2QZAysPgZwF1bcsf8STwnEUC2CDvJ3MRG6Q7OWH9f1rS1Wgbzo
DkMQ73RM6KxSCEwL+omjBdppdu3pfDMKKxC2bUEd+L0Hx6n4ojbaPsMO6OrMZl+26PNNcR8k938r
4yyB78jCtLZWnKGv02C95YqTkbCsqUxw54DmuaWFlEDKQ6dkmH+PXBuD/2oI1e83dh+0jb6696ko
CcCsYJIjKFPl1Vb8AdHBSROpaMXIHe4wuSc0phRPg141SoYc864AeSXIqLd6TWP3KpYa6Xls5wjP
AFwa6dbnmez6bGeb+66/Foykf4uvwS2W+CpvyQjQsUMJBASLNZYVWP0KDwWpz5iV6iNT1O8gp8MV
kZbi6AqP5vRGZzza3pICXehdRlC81q+ptTG5rMl7fn3ml9G6LFau3G/454f8UR/kOas0x43OlQ+P
5M3syqt+9fsvITm8qIWEPepm8oFtFBBQP2X+KtSSFcK4O4qbEyvUDOoh366IY1RZR97nUCDwvd0S
nna4U9EgEnP5XDrb+hXfZwl3MMGX1gKcEruP3mN4XaIR1mcjIF/Ik4Ju4x3YKZAC+/2wWh176lul
AICCtfcKJFYDjokCn8Q1pN3dfvXUS9tRJg4RoYnvLaJXaGr3nj0cZmrlGkM/nEbGjMLFIMzcjGO0
2hDXnnO0+4yNdyEgXqc48rS2mnDQGGdetmeVLsl57t9hxSPfAiJmJh5qrmR8f7QdCoV7n+nr/se2
QZdvjQUtCTgSZdZt/EYSLUVFziatlgoL+cZaOI1iFMoTol54gFDhNaprJTfPIjHn/wL+hiUqKR5Q
wsqpRO6f2dGgw52OQqsv59pqCXjRm8v+W5V62/GkXUyC53b3WhQmWkmnB6RHWYVlYn2fC/Hj/bBo
UaIS+DZW7n4ArsKvg+B0oAq8mnaeH94PSDVQENy6sffbTmEszlr6XtaWPGpGRG/0g2+BTuPvOWDE
daCHN8Bg6PWNh3cUXUJ7dQ8Ldmt8UJ7vsX1Ftf2YGp7ft0smnD5QvKTUQ3LzJWJxL954ltBjTstf
uwTzc9CvOPwNcZNpntAUyc8QyqSPTIMasT8H6Ecf/VL4WLq7zuhJKmdngBI2cxJ1ALUpO1krLd1k
YRojNMwdpppdrCUULxcwrVkwkbg1pTV66l2zhSOJEdroff8ffMNp+bu+Ti0xk4jGHrlflfpappr1
L/gP96H9V1b7Pxj3m/xoJU3SkO8Z4qZulRwz6SUHvFf0U94r/75JKfmnNRfnI4u+jWj2Ek/jLOgO
l37qlo9xrNV4njeSm4+8fvV5A8gjcXCLnueZUQy4g3gM57Yi953K5ChFgi0EONaUpRpWxMUo7W5+
Sd3SgtPcklushkc2L1PcyvCMNmfaYuXN2eoinj5avqNM4Bm+43sQlUyrUupIb2nivWGizrFsxwo7
4pji/ZFEN0gE9wjP9R/jDzUSw0EZZjKcTE422OIMLJiFhilvr4PZdkkEAHl9uiiIzspS0RUzl+u7
QKSuXggptrdqS1SaPDzTPFItkpWB8nwkW5EaZC2553if3zbGY/XRVZY7qnEsVJcyLoMdaNyvSVkB
o5LjZFCcLuUZG0TdQq44FNYgYrYBZyQAHp3Pe2wtCOegN9FOammQiB/BwetHk74jDlFqj91rsRkH
QUKEoSz9TNvNRojVyPlCVobJJjqJeu6fbVdwBJdV2h6Io3b17v1GQ4kAvia6Np103aopmx8hDbfD
W0kEO/9Bosbtwu3FPiAN7V+5BnQpV83uBJX85Kp1YIFZPSHWPR6t5hFt13bwh5laQSjqgjvZhXp+
+U8S6905XobqJGQJo3yhQoAQHd+HGFumBYGP47rGdf80jQJw8ksIMsfrqdc5vpnQky6iuzoFnQIO
LDglSMs568y8705sdSve3ZBfg4s7NjMDy3pgs0TvqaAXq9OhP8yJY2QIY38Xpwj+x/WDmJKTL5v8
aCNKPtBOdLyKjnplldWRty2zh/wVTR39emxoV3JXj4NLOTe8JC0Awkb2vDGUr8urRxHNfbRHR2kJ
BZpAQwVEqeKBSFK5JsRGApuHoxM6IPFKL5Z5rzfkJ7C74USxhVkt2pD9pmIUCxJHzmn6cnxeKP2o
zqphElN9LVpS9bFRRy2gKOp1abJx3QbJQIO/cSUaHwfGNOZRxvqGy36+V8wrQuCcCicZisHGVZX7
QwLFHsbPDOEI1Bcuv4Wir3mRtLVDlxuCB5mL4Mbv/umkcUGcSoSQqD84z+bMs2d6A+3Xadx+V2/d
T1sP1s5sRpAdj3MIRAD7dyhlrDwlOH/OC2u0jXphQ/j1KSQs52I3NOT9DmfDWp5bNZ8Rz5xTZtaE
KJawAd/LfJf+JkvpOcNacEWuVNRaKZIY4DfOSJXXLCvv0H2Sh7jfzvWbUXB1hy82viF+QnTJQPG2
hm9hosNTWJZcLU/Gz9FfQt0ML7psPPadhIcTdn2bvdHMPuNSavhbbnbk3bOhqd7JaUP8DRlZczrF
ll1GQdzhTb2l/BQ7SVi0OU2hUH9hKlmaFZ0LWIAk7K/1+OJmF0avd+g8jEAp5qJdPuIhYPUteVa3
+a7v5GAOf4xfC4sR1J/dlCaeib58mvuQC+mjPdvCWMnr2mXurAZH8s8w3ssY0kVNaAaTxIc1585C
98K3YmZyEGi4/BOJTIHQ6GHqpd7+cazCqJ6xqVe+h8789pi+DqolGHxK7ZoIRk3qnaSGr8VQIfur
IXXVukgzdWFdCZrcsD88v3pMQfWglKUUvGGgPYxnaJo9vCD+Ul3ycdnG9Hastv2sUFanLR9+e6Yg
yVxTFX+SrtTruDO24B2vYid6vjhC/lDe6bjyC5J2MwkOIkm7tbF8mvdhCCwJmIHo34wN3ceDipKY
vN7+LSI0waWk14W7upTElASzXQXbwMQonmspKdRSwr8h1/wjR9fOHz3Ffwg5ZGH+qs8W8tRVIb1f
YB5tAGQM1F6clIKO0/LJNJscLcMvNSxBlCEiLlU9FzyN2LHKN1DV1hzM20zNH+ohpNDocy1OoPVU
dTNXMOamxPIT3OT9kGzuDBpYy1Di+78kFmrTDlh7JbAo8yiJcyxTQQsYPd1VWmYaCdceXRHiNEA9
+UPHozazv/kMCwQJ8R4dEFaQMjxRoC+RZkkReY9ddh+egLI2KYaFq8Avzss+hPjAMwTLioJg2yNa
hF6TeoqyWYJh3PiTsrgKRgdG4n1O1juOJnsPBIM33cw4qIX/4DFU+yvA798od83NbpGqyywHrRv5
NmRWF66xvy3qaMUeiutpalKzawFySSRe0eo7ocFF+AX7U4n32boALAbbx3CooTFH/FNzZNZdskWY
c2l3thgpY8eOQDTWe0ZRY+NoqlN/N7tCLnjvv2YGNH/H5C18rtxwTFXQEdxwR+9c0zY+WD459v+K
V4mal4gQZFo7Y8EB5eyGKdPXjH63VKSXvrY3SwPmLab9skmusDPUj+ss22wv8WkQgu/jgQYqmEee
1EjYSOc0sU0OIDnwWo6lP3Y7SE1dAozuju2mae+k8ppoXP7k7BJfA6dg1kv0JFTSH70PSyVuB5El
u40E0NjRB1t02kSLG3xk+EqD+0+Bj84MK/gKDAPG5zC4SWh1+jka98wmWLANhu5pkwAQXcDu52oG
RdyqEwCyhRi6bbKuURYnIZ4klr7b4JoJm2PBUFk6vLLipmiTbOqljxZu0KNYcOy0SO5+m9WRwHj8
BF5nMb9WRUWh6dce8wLHJe5AdNWZ/qNU00Z2as6KhTWuESKIp71GgTnnRzpEklUjeVCh2CEdenYP
fd8B3KIb3fDDc9jtnvsGutwcnCcyjyqt9+RTptXxn/GSqTakhN//EYdjGgvzmcl08LpUf8giaUKL
+0fqQ49v81SjHWtwIYF3dsZFKcz0j/2g1UV4hCd/tdrt5vZqW2l0c5X3o3fkWqIAXIafhH4KIasQ
R0kvUla776GIB8tCLSnDlEpnAixIcZcwJ6Ler1Akf80qwbl5+quyXtX4ZnYL+AB17eXuc5AhAePp
djJqZfZsHQ6BUydEwulCFj25Caw0duf5HbF1wYtsnSU4tdw1WTlzk+XKiwYRK4Vvfn3ePbf3wHk/
YSmqLJ9rcrzx/Wrh10LrkPTVIO/cpXRaPPNHP9s46VbnQYvh0cCnb7Mj++vteJXOTLYJoWIO9hQY
fvBJqNoDzmYVy89IHOUz28QCI51+G7HgnXzo26SnTsTVed1EhAEfYy9duvqoTHqJEveNYXV4jjRy
WeP/uXNrOAgw+SwpWBoLbWstIJqqimaaKZ+nDROcIh4SRLqMA8oRQaTz73g0zMAtvnruSxRao26v
nfwJu0Bj3cy3y/zOvi6HmDGdHThyuABitBhbsdswbTXLqQ+9v+UXJpZxYCUc9mcWHwsTH5Gl05LI
STimOhgARamhbOfcksjGvyGqy1AwYItmbUFAhlz1oGgIV0cSRrMo247QdJIaJ50ZtVbFufie6wa1
a88eQFPws1nrH8LL+7wyscmrDW46j2qiV19bCdR2OrwsRgFLW61T0FttGgZ/2kuGpmkUmfiS27XY
WeFSEMK+Qzkj/Pkk7zh82XyPVqfmkThGb+P5B3dgCKefa4UAM6CJelOcjxpocn/xTZgj2rFr6lF4
7bCDJ+3Pgv7kxHWaAnOXZqGBLHhw9qDenSquszYD2hNOEkdFmibsAQwXAaULpC6tQ1sV3n/xSjId
qiO65l38zqDbWuFLh/Exu/7lBF5nbQUx3ZcI1/0tg9KEBh2AaX0wBBMW58FfWue5I6zVp+jlHbxI
GnWaP7AA7sALKh0m1yEnkdK4Cos6vaSGNIpDk0pu8mn/7/JPv24Wl8OftpB/6snkeCISteqf+nyR
b3RdCqyHLFn9WXwll/ZgtDzvniFeAi5uLInXH77JPKTCK5YYtjawhJ7aF5Sqq+hKzoYMv0ufIdrz
EEnz4xI2ojTAiN3ib6envbA5BGjbnAkKYPc+4tKWLYBc/s27fYhX+Hjb7HYJFQrWm2ZhDixKuSIG
VUAUCaARJOmk+qVGoahPzyKN8x0FCX2AnERkBR06rrGZR6wnf3BDIWXvudZeERKOfYCYs5qVxeEI
3LjIOvuSJgzykU1qmeTym0gBSXdmswqA7yth4Z+wqwZ98LcQABmhVwkRSNlBjpq2q8xDvE4m8ic5
uoPEfShaJ4xnx49whXixeAn+CY8x9DysURSMHmFs8EFMcAjrmdA0Y7bXkX9MWXG4gM4/vLBPzulC
f/MsMBRRkhZJh4Krs2iAB/x6kqulv/mEnV+GMHkaXlghkhw6j2iPhDjxfIA38JFZ2ZbTYGaO2jv0
vUl8iDked4NEz7lW3SQ+w9lXhBaAizv8vsbvCIiBTO453TZU25Xm/nHbgrTrG8RPBkzbTHNt9Ozd
ca0kdI0F+5ZSTPwEBW5N9FvPhXSoH9GSwoH5PdNW3H50W0W8P7NT5y3EyojIIp+Tz+04cutN+wGy
Q7Wfj8wmLpakVnI92WLqn97mmujjCENLdmvdJ9lcRq3JxeD+qK1hbXPs2Hu/EnQCA0ItUaNqjm/C
oJNSq4dEkiCkmYHCH6V8juTWiBI1KCXbyECGIVw4OgM5f6HHrIuyf+/I+8vlfkG8SlMIMzhwEwo+
/l5yE0Nreo/7MeEDvR+32uHzYrVEjmUNCjLNs0dyl094YeFZKbGCY52eRXuwcBSpYkUxTNcACgOm
Gyh8n6a+PPM/Q2YQXcGTZ6zil08LYpajVLoJwGSwJ/y1AC/kV5n8RMwi4dh4Sxroc1pty0zk2lH5
e35ZPf3X4N4eoPS9A21R10ysJmBGNp2kYM7KH/fkEqVQbgqZTKbK375r1dO2o4YOg8BRqw9AAKHm
6dW6yWfyip+XfFM0lDG/KGe9i7UoELdCP6VplT7oxBzadpePsnjaLXWa+/N9KfACMz4Lm7PtIxmt
M7r8QNkWSXUsuq5L5d3j3tm22gv28AgCNe9M2IfctUMvATi5VMkRMURhKpBi1lcEtp3ehvnt5Bwe
kBf6uwf0mNG7w1PHL2VY36aTXoEA3IHfBI7+3G4cqwiqmP/ybsywIemrB/g7OYyEkPCmxuSwywu0
Hz4RTRDAnPCj5R+FFLZ7xiB8Buv/rHs8aWOkSqY30kAwARih1M3QQSutqkiH1J2KwYppatOpbWmH
D7xNiVTYrh+xuJrSBFeRwwyVAVqu/HXvJE+ZD3cCkgnyvyf29+jOZKTtKHqaB9ap6xHTtKwHNNRe
uT5SVed1X7jQHTgYwtebtGcu1VgD/Bt9Xf/SWzsqI2u0XHb7BHjuLybLqku5eCSXRL3Kl3YVtS9f
KXl07zav42+Wue1yq+01OZ9kJCCffWoQgol1khUYm9JpOAuWIZ9A+TkcVcA1gv0PYtTVYc002eUN
iLkbPnpaFq3Dokt9N2oELNr6rsPFwZPxvAdb6YUK/RscK4NH78PrYm+89SkgGAa0DP3urAG3RoZs
kFT5YdNCRsa9H/rAv9hzNfMWfMqSN0T9FqJOXQey7gml4M8Fkz0AWiT931KS8xPb+R72U81UI8yG
QPIhb06MLzOrGjGtfaLc1Om5/NN80yrno5A6gntN34YQC7NpV7XR8cdsBBATQ8w5qTm9PKERjtIb
x/dgDztuPuetzTIajU/+d4+hERUK71CL2GwAatUjTb0cneUpsA/+BtB6Xc2I2afGLKc/woOYxFZK
UdR+UL22jPOcymVVAJAYU2fsM0d7ZOThC1krqkDpaA5jeaf/Oqp0xujEP5WrwbXNWNrGg8JOXafo
wGdSjV40bgzNT0oxhgUPEbjGNLQCDZmblP9cZLPt4NOTPIl76lHH5gTX4Bv/ibGiNqzFbT2iF/D6
m/znSuizzprFLFi+Ui4wEr8EOMJkeBijFW1oS9hjVf6ejam9G6cAJhGNMLQTUPzbPWjOQfL9Qy7X
HYD+h1kTslgTNmgFj/MzwOutfaK8Qk7gXteMU1J/Xe1PGRq4mmAwjKZl40DocPnMHs3vEHKNKt93
iklthWtsbOCCjpqFEwBEIAYKZaDwgA/TXpaP9YhuYJrSZpjR+i1j39yUZm5Hokr4RyQVP17BGa3F
5rVmj4FWYs3q1Yf4QRQQBoJef2KGzmBy9MNZnNn0xtHAOTjzj3TEoRtMPnySis33x7Sgkp4pchGZ
NZkOEzjNurErYnWl3DzmBLpNE8N+w2qrW2eafLg1cZPmjkmjywwegMRk3GEfU8BlTwO1cT3eGFwX
/d2F/C1W7r+eaSrIi1amV9M7LgoLV+Odg6cA+ypKkbkpLTqCfIJjioWfKPHp4pXWolOzLMvbC7Gg
PQWSN53LYwQ1kSEkSwJT54YHM1hR7orICvHMji6I/Cp/i1GltPGb7gWR+2flHok7aNQhY52Is/5x
rZyoBb/as7jU9WlTUjS9ZlH9n4aixT6wfqUnCWqq501KusdhNNsy4Kh5/vsi9m1k75sJ3wrSBeqd
UFLfsEKtPS5ewvgHcZHiDMuuh8i7ydBmhwXgccDW48gyg04zBQnGr0rchw+LBb/0IuvR1Cn0bJp0
u7y1iZGa6etpR8NMzp8eOfd/wJ+F8Y8M1u0xt0+kmkRGeEo1srdhL7V48ocsCd0UjmSj+eZrXfnM
h5bcOlqAiHDI/tML/Fv255mNJ8Zpz2ibSEZRVc3PdkPgyyza51kMBkgkYC6HOjjgn975AVyLjAlK
Hh+o/bJAuSN/2wOTZWOgrOepVrxreOjn260MGghMADt7mxFonaMazny+kvJD6wVHf4W9MlbEgv3Q
EClXrY6QY66V56hlMaTrKhrS1dfhLQYNLKA4ylHh/tYoXSKIt2cC89DchA/HcIz63O4WUPNdDwXD
OsYE09xMhcueMVKvLSTP4/wCtV3wPgCMbYO4wp8455gEpoSvQIzv3j2saOs44XrAW9BeNmE9XI8/
TJhpdaFepG70zW1rTDb3TNXughLW1zmvQv6oacvke/GnW+u781hRWqxevvL63eE/y7lNoIOnJbJo
vXosnpkQNKSmzUZ8sufQpgWuq62FedG1g7YWPfWMx6Z1fmvuxU6M5oare7U7/YSs63QXKqcp4tV5
IEiS5WMJxcmP0jxFT8f+bQawYxrU+Rhee7rYGHrGDJvQ6JnB/3OvNrF2NYze6nO/RjuIhA61uatQ
OvaL2p3eSPFBsKHaz2+NZcgbZH5FsdYfdKYb7Fqmi0PeJImjj3SmiaB//kQM/3nqUhIFmL4nOXpE
Qhvvjgk3ZyYKCfswbCeIxcuhtAT230vdqk8styxP9NuTcaInLskPjW1mRulxSyVPLZBGzZWFHG7L
5eDG8dBdxioGKg2v0vwrpvFp1xNn7ssC5MUGCSPz7mA2teS+N8etWMZfiffeR9Y/OBxk7UmdGtX8
tR9+ekpecGhppUYj7XHnjfsYHJxh//1D7VEU6Qk0uSh2TpM0Gk6EGEcwZg1ExU20YnVulv4OBhN9
KszqKoaFBM0pp37+rHvKRtV0/Z3ZTSZ2masbhQ+Rof7dhaxhlZM21LKEpEQ3ziSQf4lNtOF8zYcT
LSX4O0tCJBh/Rc3ADoXWZkjcrmSAoC/EkSeqPbPT/OaxKSvzbeKu/0UAHtfzR02tIly3KZJdOiVF
t63P67fbVjs6mDToZ6EcuIbzoMwaMaspRo24QGb+kaSbno9O0ZjuwNJyDT0tZ90Kd/8w/Ay9T55Z
tuBdoQIGWIamdEtNFRny3fsMDta0wZtcOayM8k57pfwWoJ89zuy1JTLIEg6599qZ31xXwdx+2dHb
gCKOrzJ4iSdsHrGq2B3VmWwr+vMmLnQYU1593XpfFMfn0ChRcAfIQC7n5JG/54WLh0mJ3NoumMso
jETj5OOB6eqnzRlY2NvSQ7+v9G5U3baA905Hlb/SwyRcU4xSZ4jrRBBUnPthe5KVFGCCEJXl1qEd
bL3zP53AysFWIcdUtnfkhPdt76K9Bd33UTP9XtXAfipZrIKXcBwkz9+daEThhwkBIO36p2dkA+T1
AWg8lb+wEk/GVskUGSUcm4mi5ljEUs627Bw6EFsQyFmx6NWmvCWaOXOsjmQ33nf1uT1zg3QVKufq
vZC2PTPMVcARFlv926MmRz4fRW28NtCP+HaAK3WHV4MSewb6HEjm6LVCLH+qCYILxd+uDG09gIJt
MPGxUJeHf+DZLxM3NGxM5qwWk34bHom/NKKrM5Oa3isGaWbIFuJBPTFzzO44rLxh4TAg4kWhB0nK
W4lXBB5gmQrtIB83ClseCEXMMwg3ORLWnjueDICCFct9jKS75LiAHSx8/XOfQFbh/Z+He8kbcsi3
mlIO0fr4Aeauy1PRs1q4DsrmiXzPvFmBOQ9F01aCQtRPVO7WRklnkceAiiVYCB2H2bS18fI/t+Vi
3r1NgPKsN5YUi1o0eB6einiSEhBDF4Gta2Z0XsmOPb17ZmStTmdLzv5/e1bip/fx2m4aeZzBQt/t
hGc1nNd5OUb9GJQxVh1ub0fTiKBYdbqpK5BHFONB2oi5qZLYc//GNPLvh002gUMsZ9Merzdpk6rP
iWzrQZj8pV+apdRXceq+tIPoTr0zOcBrD2Gxf6q+RGm4pxh8BQQ4lpXd+RLgvA7oEu2IR2OzKO+8
oBWZzDuZlbNPd+0EwlAFP/X9H57fFhvAR/5hgDM+s/SVUFm35/9wFEuej82YR0RXRwpAbKAgBki1
0gkCdUdJJexHEydnL6LH/zOJMohYy62SrYI2iV1Z+NlA6yxFpcSH71HHVmWehRXuaEL88BtMGBa0
HdCq4Fbs8LGU6e95BFx5IbYnpKA9AndZJLhPve8pLJIPPbCwjM3zvBk9fHRbm2M/CS4PjqFaskbv
7LPuKsxnSiKkIucOeupy8/trlLB5FWxIH+SKcsGrvOnoVFY9fOeSvtgUEj+HJhhq2NSuUfcDwuO9
YZ8DRsHxa2HHe0KkS/grTEEOXH7NRrmA1yzDn5GKyi4wSZ0HZXfgxUxFvJGvQKgQD863ecfuz+Ww
B9ewNBXgVSWz9BjKO31Kh9hoASG9QmR+0XYfBBQUfEGb5t2yeLynwBWAX9/e4xoU9fJrZfyUdx75
S5IW261jPd/DSPtBaPEZyk299LGTdiHr4uohxPzLTH6D5k7gvgdTsQMVzMZJIlKOPDa7F6vMw/+h
U4t1EB+s7juzle9uUh98RfWbSGPtz2hG1xw6M3kjZNNyY3SXGEB3pcfn/yRElPEV9TSoJrCnNS1e
c7rXDR0x3mFaZ16hwE/JhPm4CgKl6nj7llyj4Jf/Ao3XfT/PjS+FmIPoXNLsd2Vu9EuM8835w5bs
5xMS8vLHirkvK2Y/pHroKB4FrH3+6WCRYOQ6u+8kJmAc6Szlr0W5WYazzT+AoT6CqOY7fScEQb2a
76f2wA8aWGKsXbYsZ8rgpLN6C/uGm9f4MIpm5Sngtta6wK8Aq872blUtiVI0ZmYq1w2tc9bhi+bw
HNLeblsV93yo/VKj21Zfe4k1O9+2Wq1GXSoanx5exrEn6VWl1KXXCuw8DWGv3Tn4WEdoQz6nz2Wb
3oPs3BAXEltsHKmmhGcn2DV8fUlFcQ/R+lLPcTX3SuqmSlqmRO9Q4PY7wvBHK6gQHCxmqcb5698Q
9d35JevEZ5DDQvHkpZhrJlZp6AJy0exlw6NsJS09IEiKUxFMODuM08x7zVnpMFv9bPRanw6zl9Qx
XSfm+9TZXE7ZxT5gmHzITKCOjNiN8mrDUP/6jajxstTHEQmaEKEAoCABPOHrH99tJTkwvQtPOYfw
UFOMT0V/xQQD9+2j9S6uJmcQ2IlODD1cz/CoSOH8MLjmh7YsD8tFpTqF+/bv8IjMRK5QgeNM+ZvB
dzES9bOgaAd1kG0xCyx3i0/ztUaa/uaoMHFUX2ksO9p50wTuRnScOWeAenVNXyUfENyksL0Nozb2
KfKD2kIsPIPVHLvB4i9cMZwWnD/1jbXAmjLsE6RzE2bYV/2Et+dE61gQ6Ir6okpel9j97XwShQkf
k4rp3SMyHoSgz9AxEAU20sdKwEIO0EQXal1jsLet/Sx+VlrOWvhWGkz/pIY54OrP9olC8VeT1W/Y
81ES5lax8TSG7gn2SudQgFm9Uv7tmvdwMQH8WNw32igJtkWaDUx5QGZp+jD95nEbGC3VG+7rE/FI
f5pII0cu/44Vrtb+3uO81j+HxHtGUr189hVsXwGfnDpusPKsTxSM61pWUyMoYv+4voJI3hYOvsOA
T15ha6nZaanEZSjR4rSohIXocQoLjMcSSQyu6o+Sl/X1KaH8jxY6PyD5l4qhh0Gua5grUCk+xT7b
nKKqaue7WvuL88UsonScMQ4SeqnaLDjDz+CfakaBHftWrkL0+ePsbjnmtDJxmGciBQEid83CsXAU
fh8S5hoGufNiIPOO1BEy9fpGxZznMv+VQyL1pGLZBlmNo0TiakI8U5wwXTGanidG3/qfVB0gbxY3
RgQs+0/toD+fWIxTtw0JXQR8IIgJH40cfseaSOIQ4yv4/SKSnyJR2scf47Jvka94nzhT1dRbZyXg
B5AUowKAXKBKLU2L0GEZUdR5EGglj8l9ekwRRdq/cWPDUG6L+FVhGTpw9aWa5mEio6URYf7abDfw
m0X+B7pSgApkoCL/TjDu61TEeUbBQw06gP9Ba/3v7EkbcDwZ4HrrCTG3oJhFOy/6hL4ZXtJ8355a
fj6BLnakWcRbCDZeFIxIUPdHqVvstPgXMWL3UQ+pYSOpD04TJRhTI9/swBtsdOISX/q8k/94goFy
lRFPI/XDe0Sc95iCqua50xhZscDWWh71+NEiPDwwgy8do3AOo7QIoPejwBOUknYUYdjni2SIPj9R
bDr5+u95BdZmUMJn8HCS8OPyTK7LuflUXsHN8M4/WlwWojpPyAyIoLCilVNKeqH2HilaxCjmIV7S
3WnxBvNUxeKJaxCFdrQbAIIaAFDYmaQIYGgi3iVSt4x9iFikkU6oLbkmTXzPE/YJFDdVg55E7UwL
QHYomCyLuE1Ip3vFbm9CXj61ElfRYJQasFHZgtUBIuTf+nrBMJctxEWHIn5wDUc3WBmmVelIycKI
Gk100kR+mlSG1kqAZTzD+JaClFoUofDpf3fQeDhFmwxFsx/xoVxSEb8W9El6bjmtIyns02zTwrSv
N9poSlipSYJznehR7fwQFObUmggaayzj7EYhKz/qdwgodNaL0g0aeDbDbbWgtgDGbptnuDl5//vG
lG+xvSCAK4hw63GzXUSpXycSZOLZCJ/rzFs5yHNvpthaJakD07vz/RFIyXiteEcEhDtfVLBa1N40
n5nhS3PMagcoEaYCQa01eEtwOpG7B99CEpigpPdrneT25lZsaYoeghLLFFnE1IaUMhqm+z6cn9lK
PBoMMIPie6UmUbjqW9BhkOHEckZnZwfshMZazw1FLKSgRFQ5TfDo00shE6ot65jE7zvB15aCgzLu
9r+WHbRNAP1wSht7ReUeKnSjbRX7nI6Im08NJjyTgjlPXJbHBmUk/CIT3F6sHGK9NlkLwoHg7+4w
gE4kHX0BTRTBQJNUdDcCemuJ2XqU88s4Riqx6CsbS70/MWcmZNwcEm4OLyAbvTgEZmWtvE4lbGq7
mEaPBJ4vIR2/HI5Au49uY8BIGKT5LD3LLWVq9xxTD1jLg8sTGzK8mcJRUduLlP4JAfADAZ+T8LJC
qRkrshTN+g5dRp+k74htm4nCRW0LyPAdvFtdqorK6hEkbDwO2xeeRNhjl1cCYQFrzqN81asqVmuo
HGpHDmg8LfdYBqqrWRPblyhnbzUK37flr9S4O+AbybyOydvTYmfUnbuYkxXT9MMMFu19lqp8Kh17
BbZzk2y9UDWg5zSFNkuVsEhMJuP7HUp5r2ekcR+Tz28bgPaxUSdN5fzfhrmD3n9AvXtBTJIM7f8Q
UxVlS4SpCDCf7PeuHmQo/0rNdmlRtmqs4ioUtaxdclUYcVP8zUhmz1YXkUzS2f4Bit0GoBD5iXo0
kFTQWU7982SeIoQVtN9e7jQhloEjFlSeBNPwQin/LTjXLoPf8ecVfdJ5zVtl9hs8vXlXPlU7HEK0
SpqfeCgF7x2RR4FcTp1bGFZw0pi0SXoNb1VJMQBWPHL930m6EzZxcfL/T30kMZwcrPsBOT/2Dn7Z
/FLp7POgruk+zPvN9JHVNGP4qFgEAt+IWJ6rskzsIvvVgGXo+wFL+kJuriVPMsoyqhVhzCYJH9RI
M4cMcwwHZGgrVRW7Sny/dRRnmXCKZ4/CdobwwOgbIGWTNa+8z+6VjkRBLjrMTJMAxvI9gYxEvt5G
86YLHu1qVFo7BV+I24r0O00eoZ6WjZ/8EeR1We+LLP2tetAzdiZBT54GSoQzSgiD1pWXLISHowo2
3l0I9p0fqSgnOW4aBmE8x+JDjWsScdKtOrqlKUK1wJBgF6CXHiB8M6+ZEslAMRHq329AQjmY7juo
mBwuPrtQdecjI9N7t+A0czyRIEuCOnFXDydbN6aHtqc3nFobQ2Pf1fzAL9d6AFELeBWW4nydRPfO
+ZbapQ2XgxfE3vZFZkSNfgrpaOAYoPJkLwbJ6T+sfajNC8f9aUmYVWAY75pS9S3CQitoRvCSe41f
Emp41KE6oV9mx3TE43ksBCNooIncBX5BUEOKu72ufp2ofrxsGzlMVmMBe0b9N6g9834m3Ov0xTwd
vJjgb5Ls+S6XNiaoWpB7QLF36tP7vUpjeGvZqG3VA+OVsgqUA54rJogMFlizVKaWIRLiVF9Tb46i
z3KkJDbzhVgFNXV1QvRkOjDUs0daWR/1tk+/b/4sKqH8ZF5a/4Rk0CaJFb58qgVQapCqsa0cjasR
Jl5rvQf89PULW6Fpv21ds2gHQdN0Akxk0PM/iQ1v1X5MUvp/XwqTZexF6FGFl4dk29OJcoN5ApMu
T9tBhlyrZxCiolqraKXcfg8xlfONotR+z3ppSU3wzQ4cb0M/ujHxHqp0826/A5YgtCUkYJKFYH87
ysy5QAKXXifQvDoqaT/gB65Zc5y2vehP8Re5MlLna/Y8NP1fOsK6Sg8sxNt2G8vHP4rej8bilxiv
JuMHa1kw5RRrnGzzjZlBo/PTJPs/DltU0q7I96wDIz5qF9PiDVFe/DMCeWvMtoBpjUTQGZy8pYt1
OqXQu5dX4c33GSuemVD/30KAjA9z9SvkteK2Dqzizib8qDbo+h7IhvSOCvbCk26jqkO51EMukjJS
75f2rEY+jP8bK6p9/tY3lVZf7Ko4hSg1U9mBn6U8uDOuwj4yBzbdOqnNiVPl83/lBZKgki6USRZd
K6oxIdFoOKzZlABuQ0g7ivuoNgR77VBZc3RZfNzNMpLkChOseUBnevhR58CXYeyEOAjQuHoX8rtj
IiDUXLYuahGMq5oKl8FjlbJcRxfIDdjIyfikmSW75F/I15qN9uYZ1drTaMuyOvLuXJxHq6ov1eP7
zfyngXaBkIJxmh/MiB3NHlsqi2rK9366s+2bqrzY/bwa08qyGjpJABZgaw379MeU3ydqxS11z4YL
u8GZDIv0Pa70DTeuK+FwmbXJAyltBe3sr/E2K9lG9yCE6qxsa9s+MOddl/JYQDG0+fDQ5dLm9FUk
zhsNlBcfGcJEv3Ifg8SnkZ8GjAW3cFsv2JNYS6+GsFkhMSRHOGocX34PquT6IhPL1+sWcD0vP2jB
oZG6WIT3KyaawffSfJO1JPpE9NqL/4J7b96e4UbGPxTXksR9NMf/CS7auQetH7YkyYglmy6JwUQp
nsChIH6UYIzUoh7EMtxTSl2xHawPqWCvXyzwttOAUZJmuBT5JQHkCaF0xftmwQbDAQVqJDIOCDJ/
TKKqSOeKaCcZMVn1a27ny8tcniWSnsvGkpubB8OsX8pyxoDDm2ChQj1PFEdeBdqpvjFs2K05UKdx
iS9CqMDNA3uLdxuEcccOFmdttDv081lPdEQFLAJQtCeVCEfsYXcXsjTbjxkhFjXeVbN8GuVKh59f
ABNQO1hiH/qQrqyIJhSRLyotXvd7IeAHdyI3eOqjIo3w10n6k/jJEY+SBa46PWrynm1H4y9lyKIP
g7EfzoYOx6vBzBDDggJid74ElzomEAwpqWngH+Em4Z+yhC4WaLRHNP7E1rPY5TjeoC6wY9QqHDQY
RzfgPH8em7jKkw8OxUOJLk4MTqPfbcK7R3WLx90GKgyGsTp7sHhdTf/Erh/6UL23Sy+EjQ5zrmOi
iv4Rhg7s1J9k+Tq3dP7PkYtZ1IR3nfhKViTrDWwp6YqIMa211FNJnStE/nNo7TrvKYZln4Nt3vvN
Xj8MKJJcAZL5YG3SDHN2w9XY1LDhiF0jEl+rqi+lKdyyWW3YQQQyvbufObXOmPS4YyAsPskYB00C
tC4lywJomSvbEpIiodPeCjl2XxX8rabyXljQ3s8L3CibMOBpB401zM3R4L4QiM/oOrgRUuU3irlJ
zoz99Rl5/J5CLp0Mi7GsW8fOOkpXP+zBS1OkQ3FJH4fI4tmn9VyUcnhfRiAIuKr/2Z0qqsGhpyKv
OJswf/gA+Y8Q59woj6HL+cUz7q/AZ6Tap2ImKGIJJD0iLrJeK7ZPzpqx93PuV0zcvT5Dz+wZgU2F
S0WOSc/0jUZluRmVkbsTABP4cRe76kXHrurH9Q4G34x9IBIV4cysLQzcr7ezC4OrcEzY8+1T+BoR
b7e2+/H4OOy4h2ksDC/kT3Y0w7WH7O5P/zkgp4/WF74L1DqbHCYiYsUmLkMyTXT35q+Jy/hamK1u
12OwA7uWAmmbmpVGEVwrKls40iqB9wmiHeb8K6PhFL51ZwKdod20Sf2ytbhmSIV5tV86LoVNbx9o
x0nIEFZSda1Q7wrbM7LS3CmpJUI5mmxSvre2L+ZL/fb0W5bC23jHmuv43a1WBCqTnNJZTdoiGesQ
mZjJPR1Lb6GlHbnyo67n5GI6OCM1qZSsPc1WPTICgENLZYQeSzz/bXLAvA33oKNfJ+BdAtDOgwHK
1frY34dE9NQkkvo8XdwMz6EByeqXaM9dC4EEh+7ehplEOR37+hnHHdRmRYNrQ3P5EUsiIFIyQPbj
kL4jvV52xDgqfpntrycEYf38/3ktJ7uns1Lpj0Sgg/IeD3QVzl4CF8PU8ufDeyIgW/Qd/Bm3TbWs
4QwMQpUp5fLVH4/l43KbCzoVsWzTBUSJCS92ehQYXHGP9SNt3rIHFdcRyeSItAydgovA7/Ln6vPo
tsj26jelMo54Sp2gNg6ZrVW61qnqBeyCC8omeaBi03INWLk7gNzIgBMpCYRYhk860vigekfT6AJ/
nab/VzEopVhG1m4pD6w1ltNpTmlpODBV3GJxNqQxWg47aJW7G6nKg/4Kiv80jPz50/gDYgwrRl3/
50ffHE/eKIu5BUygDyLkSam1gYzzOayt0+GkhF4AU/MIai+G1cqdSqUBaboDcSTmlhQZObcUG8HW
QpDfGkrBxj/2HmZ1L/nJHd2oGZ0qf9Xq69lDxNtcyD0bBAGU3MqvhvfLO2aRGSET42hjwZdUU9LG
sX/dxy9beUrCXuahqRQGuZohUykCXTOo+9d4XWoL+07U2Rwl8GyL6khyrHb4/YOOBP8tErsZRDtM
N1ewWfhWuYLHkGQJltqB+BIR6WC8lT1KQ0JEcUWHNQVl0Y+mC3YFox6sxfwcmXDKytQcejGaoUB3
fqwqlZ/AhDCZv3Bhaie0WGRXkDuw14pjl91r1eEToEFCYrEYfWqqTQ+NqJ4f3uB+AmeKnwADOEWa
mWbgWGKUQonbvJlqOr5aqXFYo3W/eKfEJ7qJQTRRhcStrhAEnPeQUITpBPUsyKAyavyRfPy0rp5L
J/euds0UYHJQ7sykAqZ1Z6WuqZzyM/6zXrPyQE6xdqN0tqR4A4kEn4VbWywlNcYgZ71lZoRt68Hh
r4GKcmi+/MY0pBtL242j3lsZIrceSUeqzwwQh2yEXc4HQVdvx9jw/dYiXVpJcxF1RZKqpOevchC4
xGUh+icVhqluUh3dLjVO64ZX6F3P/HvNicAdfwsm1yXIUsGOZMP0LshwIQ8Vrhro2K4u5z5W0hr7
4nIIVr6RLaadGZ1ZcFII2OENew3o20AUZ6pzFufVzp0q/AktEnCEYWqBb3RqyXblG8UnCRp6ksSm
Gqb9e8dCBNPOIdH0w+wpCr8DSkbshcYAAIM2XGsGplVCd+tbnhBOCFnDLhSuAhRWnCRpcaX8rbWs
rc6Ep4uaaik8VZEdXwl+PX4zlcFidz1LD2/UY7OxHOt4KDgS8mUuQVOZSMX5GLlVN6sWi8jFRSwO
nLSePAZdfNwZOJ1BB9lWPdLpe+ihAhPf4d8MtDabC2FnE+okM7fUb77kUmuiWSBMLpH4ohzIhTF7
D2haeA7Un8jVlslS0ggU+76BUDQhrmb42udZuuqadsDV+TV6Ksm+D0B/uwdMtq02P9vqEzFn11F/
7/mcjNO0SNJDEs8LRnsjhJMFCHOTYh162R9p5SclGRZbG34w689FiqBKpZoLLLrQmqtLjYS2aF1P
lxARpDoB5gKxWX9Ht9Wyv2I2G3uKL1+j2+PdcMc/QJDR2NBpp0wnIKo3U8qqSCkFyZDz69s1nahz
fVebColhtw68J9wzDiciEH/v4ff/SiVuf+C1FSbhl1JOAzeIrdcQ7W3N+RGegT2ZFJGg/plYajk3
I1G5ibWz8iCijR4ZCVH94xx60v4u3iC/ya3CEqSedZ7M+ACMlFE32YyRLnfG3R2poaz9SFR2J1E7
EPhYoRiTvKJqP6zyvL1j8hEqUqrWiXijczCjIdeGk8cLUE47DNowkgpF4CVSSkENduZ0Bf3FqDW6
WtDJfL0EFm2fU3vu6KBeh54pWEyUGD0I3LRYo1SgYHzXDt3qaoVph0qkA1hHuhJiVoh0lJlTQQnr
9OIUYuRLxFWzzDW3xDOaqyQW4iNgL8ach3aZnG4e+6Kv9uw0KzhquIs2EcrOyFdR9aXuxWEnjnod
a3UJTUeUGaAD2TowaS1xXpOySsk+KOIQM7PUMIQt697xg/Q6ElLjTi0mfIRN3yYcQCynqHCq5XrZ
22i/9D2D/P1fU6kHhGA1ekYB2j+zoXF2iF/CiLy+bV9xs6d/b6BaqjnMK3REG4cTt4G/WwaX4SOt
EoYak/XuXkXlWKAV2l9Sn23U0xhjAjhpYfCTXJztKIW4iWKKdcn+j0VwI+kj4p26GKGeIC/Uw3Bu
ZbEtvHTAwtkGRr5gfhcZu9rnSFJn9TJbNzHmgRfkIWn0Vu7DIYJaMJltm4BKTVBCO0DgrkviBvOg
uuAhnCB8tNrfSgllccm8e5Vo5RmaaVEdQ/6uj1luu9neZX5vBi5Y3hS/6mSLRxixP+EvPrdPsV55
hIRiT/e2QyGo/uhMQUomdD8TT/Khauwkt3hGJ2vOlBqzvFzkjoSpBwmABHxBqcKnO2qN2mKqXyeg
+rUBxGj2/YLghkb6DcKr967ieceifJ6twOeNXjH7ULjwciL356Z7ntmgn8bhB+orHkX+k0Pm9bzb
bfhw3hXlCG83Rl2utLHyfpNWc6pJhUMCFFHS2b+M0JhiCEOEeady9d8iYmRRuuf/ssR7hIICNcxP
MM6y5QxS6sgpn5h3wyew/8KnNlvEQCgsqwP4aguzPjXZp8mO0D9zZooP/t18oCg3A1rcfs1CTZ6w
k/uY3wksRmLQcXjaybyT64h/hwTaEUZskl4N/xxLa86Jt+SEIWI00GK6zcUuUIW5ejYUcE3vSXub
8gxHdvkazMjDyK7gDvep6Mp0OMSujk8V1Te0DZvSd1jUG68aRnbtc8/OsIfnQi6Wp2g4ykpWKDz/
n1oWO4+aVwEHLtBd/Y+c/yWWibSp/p2EnNZU7GsT0N1bp4pksEB4FYjGxwFaA9MXH5R+wFZQPHWG
3hMUdnmosY7k94bj7/0uFQjh2h92q2CZESpyumC3njcluvOnu4Y+5VHg/aygrL3u4aratU+FHpF5
Z12tVZImG0g0eIjC0aFz8seJQEZ5C7Fqzg/BsnCqEx4mpIqY5OuO/OdmTbO5nONkO9pz7Xktlpew
a+QUqyxo2P5LokIn8j8cN0A3Lmx1UW7GjH65LBi/GYKwezj1CxYRdPuQ91QDx2CkXhW3GcVYMVVK
I7Vtpln8Dqs2y5yrO9NHB4O11v6bMV8kA3SstUi5mkjUjPSlGokbaZlxHDlgEYDo/7lBU2PSX2tL
eJ++OEUjPztMEgwMXxOeDMdCzkxh1UZpuNKCZbDeDlYIwpdOvsyk9G5JJ0KL/twh9DwJw0mXoTr7
Lds56Jx/nLEzvxiF2BSZKpCVXe6lTFk6VHiuQh9Zgw5AAzzQRKwXfa0XcsDfeal+Wztc6AQwm+ew
13vB52c4bUazJpmy8gN4PJQ/lZ03Qkz4wjVGpmfFtSxg7MKW48rxLF5tIbTrY+qkeygoZPZ0I7lb
ufD5Kb5fymmjP1mhQF5pE6exftUcpOB+6ghZgpmQxNjfhT2jUVPPHy8HGClh1XAC4VIIx12nUD+z
CsNWMrT0ybhBwfWxjiMhvrseVOUiGqFGK9tOywvSHgyhOzUttuqoIXvThq1nz6MZOp2dY0ubFXbI
sq3aEltYa8VXL1a1a0zhA+hz+XSJHcNjnl1bGE1dLeQcMr/uWmdl2iSPgViWdskNILSn3R6HTOhG
M77vDxSzGxGRwTFA7JlfZUIGKw8b2ikY6Jhk5PLX52eff3IQuo+RDLOeUHsvrvfLYTvHy1N8QIqg
OfxWW4BDPFDu9M3ERFX8SEwYnMeLyr+FpA2YwUzAz2pcMHoaLwMUwjxg9wbbECkY/Kos3pwkwR+6
fFIwKI653U3SF5PaTXsEprETJPj8NU0qIakNtmMn0cl6N7/UzPvf7PgLmdTa3NumX7o41dOCvizD
wFZ7B7Y6JhuRATVocY4EUhnVcHvnhHsaAGL3zQz1VObBdGjF31uAL+/fFanMU8cHShI78Ck6nsfA
bHC1oMitrCgPbNE/Voe8XEfdS/Voo63/UbYy6i/ds5C5R/j343y6ZvxI06RHGS4AEJ+xel5+CsRi
TrAilEU3e5NfnEzbWhE1QXog1VLwEWv7IPT+xIroh1/w/3jNkuD8QOaTHqOkwPGT/G0DuYZBCloX
e+nDteFzBAzZ1opxf5bTwAmogjtcjPB+09832ZjNIZhXebWiV5Up07WQYe/+0t005Bg6GTvV+ENm
00F832IEbV1ZpCx/9o0wyiN10n6Q/ZuLnUzO/xtBh9bjqbuhJX2jTa6kNFXe6C+aIad/VgWH3OMt
rmzOGp+HBJbSWwMXn+WYkxTcm2SZ73whw36atV/0FRIeXGRf2Z8RS34dDsyr7nZ+k7qAB3VsJfLv
vWiwAs3il4NdIqf+mvOMle+XdGhFpN1MlvHvTmw+GsSHUHM+FXhGxJ2vRvAJl2naZ18XongEAhYt
9VQkSsC+NtfdFOicybr6uewKonVOMd7KziBHarNiCB6CHXH+9QTc5nxo3wItMfc0MdcA+N7RCHcg
J0fWT2p4GISzNJajvO1IbjSbCXysuXuLpqnErzsiskLgEIrFv8ILqOb13jeo1VcfHU4WtgyHlC63
+rdw4VRdovYKqhL2WKAmBEE0h2/+5OKdOgPAgSgLNrzOrBPKEjyxd6pREg1qcLQFgXAB+39xPVi1
QRSOZeeNzExFn14daO7o85WgIQfke0Mx8oOYqnsbTegCR1EgTIok3ApoqV4la95zwDorUZwJTogS
2nGiXUYbFYnFpa/cve4LGr2GuMwx4MAt9z5WPDNhnzvYwPPkIm5eVW/TOqQoruziIVcA7z36zw5F
SLOiEmD6nziW0RUo3P1NeIl6KNANrwigkJfxQF2ppLikmvGtV+TRSA5S5hA8gg8LLKHDTQE9n1QK
/JerOqZbnvpUMRFvnFXAoR+ZeBFsGSaxTt6tqh9CkVpmLhXv7nsokCXSbEr0uAeIncjk1xVtn4Pz
GQcGfuTIGDHT23K7RqQiSMsdIs9dNxXkYgJ6HShHpNlFm6W8WmdGdSNzqzfixs5iI9/00ptAszvj
F8+YAO8wl4muxs6F73bwQeEGShoR7uQsE+qlRETkwzpfySykYsUcmNgk2yM50eNxq8EbttVykvEw
tOeOCX7jUMtARNkt56ZxPQvvcIgxEUCH5rF+7yHlMk6PruhOcV/edxbwrLehJqthB6XKhxjbT8Gg
ow11Y+VlCk8RalwyUKdX+Avl17aO8+vpcwrLgm/SeGQ3Tp+WOqXc3PhnRYUYNbOmRwU70El6/Hlm
QU4nTFL/E+eRHH/CbYPjMLczelhYEDOBoAShTbuFnpWHtNeVHvAHls7JmwPn69MkjW97iU+YOtxs
5UumPTxCRTVYnae98id+0SdwFK80J/+a0MrtsfgYYN7YjoXmmdNPSNji8ANiGhRP3fETrowTMgfT
EgxLKR+ZXPdRau332Vg1IjssK7ID7++qc19CQFwL9kzynUKpZlvxc44uCA+1sRrMAadVzYMbZS8/
UWAbdgQ5ORndE8I7WCxYE39Y6xlGOIcF9uIVV6/6VQ2qgKGhrp8XBvw7wP1sdw59EKbI/Ss9gqJ3
hj7qnSxbHEeyo5WHmJqJudeamZZdC154i2h6XP3E718aEFqVcgpwmBM8gzWpu8KnitiD9NgeSu1N
dlYw96ZBQbbKp0XQ5qOxIksQ9OelJ+o5IdaR59yAZ+yTn3JlUUZqMsEoQjL4IQIfe2ZGnPnkwFht
VofdcK2s+SS0C7LTha/RyefGzHc4CTIVs5lza8GWWz9Ylc74Krs86YQfD29MXEzUrhonMcQdFHL0
jmqEiJ8LR/3tLPFfZk0kOWuFJ4z5AcH/h+Wd5QiXSFkBsT/rwaKDfq0M99HlN9bP4anFfqpalotM
SB49clWsuyT8DepyAU7AkwfZtb31CLXasSI2anLsy6JWjlFHLcWgXC9wESgZkM29rxa0vUpb9pUg
KixT4nsEUS7OovhFB4CviOrFHrzDgj08vRe9Pl877JJgaNz7aZU9wQAkhv5XpsOPcoDCjf6WxU/i
iUO+sioBk049OQqgdExTAQTBp7kIzFLPpTTh60clFgbM9NRGSUZv01jYbKKhjoCz3LUICVH/rvYD
uUYg2rBuoUYA+k6KGU1vEOKXFFiJYQlpLo/R7bqHE+B2DReVNBz5XsYn6YKAzQ+HS2ODp8H8xDnx
BOQcu6x/kmUSYcWxXtynosFAx6o5HTSdTKUUvZq3iwkxnHKmVlLQNVuXaNSGTKWdVaGpq6pxGNOh
mcoe8xgf+bmBO9QgxiUsFzmX6kX7Hw6xoiX33WENuIXi42U3lbROOdBvDXxBA1EmYD1UPReGmyMQ
2LcJ82BekCAybbvnzpKkQ/eCLzFY2K7JQjDrVdQw05Q+a4OvoePXb0VsYPSIudCWPBclcQR/PXLX
zjCA6ZPhepj32R2JRoNfSSMB1n9VEk1h4RgwUOI4hpfLFBeSCOTcXpYVfdf3HJmI/gPLwUsmfjbX
p+UHlCDUVhJGVbluvOb0bHeT5oqyyRvJ38LHhgCBkFaV9Z7PN2p31chg+brxDunasv2+f/xs6sxY
JWPpZ7gnmuyFsOtwJk+ng8gyR59DMMouUs5v/Ut/MHBmghcnLwfPYTc7AxOILjO8QeMkkRTZN+xL
K7pWHgX9uh0+SJ5wBRCTYB9i3mPsQmoo3JP/zg8GO2sVYZg0vKczCKJgA/N6ZBNHFPD+Ds4GGpWo
/xq6HumF1L0tf8VxHaZ80bh5gv015+i9TkQ1ytJqCjURqPLzMEvc+eeAOt9vomnMBxT0WPEAV/58
UQ4Mr3a3vUUXL1zmBVc/7TQU7bCqQsvR+bKLUlWy6xDn3U738tzl9rLGrDgm3y2RhqPaEXUfswJm
Oet8Lj6RJ49bcZjKOtdsS94a4W65kDtqx3xx4NfGrqQKmDVxdvZ56RmEtDwbK5+507vzEaBWWySq
SNTFZKIynxTRCUumgkeaPA2Jr6pseK/t713iPszZTGFqKEqffUDIccile3Apr67AqFCb2eKrjr5b
2bi6uJgoErcO1fctmrZVafX66TITGnHPT+jMhjWu/e+HD1CP1pnY3Rsf3gQ6lieXpZrnViQ4q0nk
WrR8aphbecA5cXL3IUNLR46yEUWATTqKqAKVMQFWvXR9X+RqYdzyZAHGAcxzOBbuRZfcGlLyXng4
8MNkgpAkOoPkuQpayK+OL2OEX5djvZKrnxkbUBY5N0ujy0KqFmtSf9KqlS562t0DzrWTRmi4GSUe
NUNj0dWY5g7kZDymXBll1HfSXomFG1989BZ9qAME5wVHUyMf5i0IvxM4Z8z3g/F5w5AS/8Y7q15p
OLVrAG2tLCtNE1WVGRhQnftBcBZaq+4OYrbACsuy6s3QJA5+uiiN2VzobAT9YMq8H4u5zOgt7ZBl
CNMq7clI/ffqg+XS1+as+qK9aGwLJv9PZna5ORGZyLIzrp2hT5isYiGvehf1fCtjISpxJJcT8xcl
bXo2icjFG+l9LceZZpcIUcjigFqlwjym8bgeLNpT/Oj9OcaxKJ+q3Qlq/ajwa6pqj679oa3/kKvq
wrpDDtg0DDsXZEfNfjAKWuZ+7RomcZEoxztktM/cC5Kgz0kEnTEpfO8rn0NrjM+akv/pl6pOBXJE
19NtW/V0hIyBN8NMxt+eqE6tiwEJIHvUyVRJoah6lUz1K/ANvyHROAYml0kAztoNy7sF+kjy8Tp5
/Jf2KkZ+/7ZrQMYDPEJ5c/bmmuanhUrDtqBfWdelfd67DfwOBp+d509Tk+5n5rUwbIgrDrYN2jW0
a9Xzjp4wRJae9fxiEIt3QxSDZjAIx2NnzS5vObsbB2XJV/uGGtDmJalkmFMgCVOLWLr6nuHj77fM
QExe3GgTCtXIRTmmX4gLeF90NJpS/pP4cCFaDiK+Ls68dJM7wQEU4yR29PMLtkIPpTr2xYOSosQG
cQ6v6vKgOU3M0jNZFCn5rdmj804HmpSrOpsX2+hichW0yqCLcmF1lVV7EpR6rohTdfIeFGWuW+ox
z23towlFBHZMf2HyyNcMWTdy5a1c+VEUtF6V2cE8KLtMo3q+Y/kOkJft9hzZ+lMqAAZh027Vth/b
bIDAg+Ssh5LsdWaGAouiXscc87OMyspBREfblgUxrc7QgjtL8NLLLp+l0ZQN+0uW38tvPkX2rBLS
W1N49KrrArIA+QCOC5bPeRMihjpGy6lzHMLjtkeUCfa6u3cQu9sDb/U9S2Ws5WTq9vyl//vQoi/Y
KE2jTOMjhamRW0KWcZ07iMwtEouyAYQbmCGgobmGrTb6DRqBKO47loOxG7bmbiFpGoQWz3Vm8puo
saXjjf295hRPQXn6ZRmXXY2WTXHefYcRsdm0bokbgX/Kk0nopNtgwGaZbs7RXQ+eiQbDlkw0qer3
r/goa+XVStzRFqUI+QW9RLBYtkBC4LmMal0izUAhKROcsR3c254fVdRVryv+TqWLyNyyL9yhAVrf
dEe0r7ljCEjI6SFBNveTqU0RkBPn4iW6QcSdo36DHsxv6l0Z29cAiYJneM0HEV4I0BCQnZ0MH+Wc
A5qL1DfNKks8/yuPtCm/TFi7EA9OGwPXSK4PlPs0NOoxj5AH0sr8yQjrwWoUSxs4lfhGVvjxt8AF
+bfkCqFqJCdD+gfo+V2OlMfYvOk4/aK3el4wWhi7rDC85SkxPfxo1h/RNSzpikQUu+cq8y6xpyow
xk5aqN1yumx1i2Tq/hmdOoJj33Ps1OM6DPuwfntyu/acvhuTs882wNBvZnpMyMizmK4lR0cxabc3
HHsLurcbW1r8zC7jCgFkvp0x8Co3GD+KYI9Kng5SCkwIoIWi082fuh6VqLA1GgT/hbqexZqmFnUv
OZsgWKu+o1PKvkbkxvPct+eF06sql34BHo47fVXceB6MCI66sELL6dqXgKe920Tp6Ms2+TBBYTKt
zOiNUwovxm25h9KqN2TiqdkMuwI+zzbb47drzsBXkw4J3Hm5iLNzLhVGhdsy8dUlkhSKeuDAwqR0
akH1CG6IM28N+tVbrn2EX2LBJHeOrf2uFOZROBEH/x1gWDq/ZNGLDsUSDzMu/SNj6w/zDe77XVob
9gcElLoUw/8/CkVAqvC0/z0C3G6cTlaMIevEwcCxHIR1NzpDGvcHVQ3ez9ekTQoT8c3/Bej3qRIw
a0I0ceKtXE6z9zgYfyNA+v2wPA+7Ud1zj9sKgxtjZ9VMb9y9HajFjJeJssYESp8InqRy5VgrXrBi
YwQ9jC3oK2rEb37R071RsIijrarptYbBAvSuFb7YmDe3krN2cK0uAfOhLRBKo/cU3bQnRLHgzXke
EY5Ydf5PE6mBYyhXgvosttkG9T73TpG5RCWBX0zM5DbFQIECfdnACgGjTso2uX8ySU85iORq4Lb8
90oAgUpTOuVhHFSKTWOvSxeeMIJ2jWyRjvPMc6JeK5h6IA3RhmEzBTmTuKx8e4vGTDTJGEDwFke3
RvQe+0lWDrT/U6p8oYa3axAfwmz4reI0A7yoEAAllYnQLQiIqrJ3L2X5FLz63uvK7t/rqrPlmIkT
mvvBkcm/ash1Nkc2KWArdVyO5DR0b88JfUaCEzJ/t8qZtHAkhCanVRW5DHxSlWIAKP+TgX02tPAJ
wVgDpOo7rpXUdmeitwRCdLJa04jpt2qG4e0UvheSjVzqCHFvnnl4eO4aPvfoCTR96Ufx17xsFtnk
5kfzzsYNXcEXhsJ9sUke8+TKei6xYelkcA5J0li1ffKJqh4VmR8c+TzU2g6lf0pCmEhef07WQ3fz
bwSWYpk4lk2v0V3YALFbj0t3WyaYhX9C052ARjU7gIASuwplitHUoxT2zirqvEzfjBlReHMBLSDK
ryisGQnxpglIAIHaP9t2SAVQ8I9VbSBwJ9MZri00eUqO0mIZujO/OQkLN0NJEsCSNK9eLM4U+Vze
cgIRlyxXAEN57Zk+RtTy7TBm4suQRZ6ZnfCmpm2OnSLTpZICBILP4Zf54cFxDfY00iTkuyjIzGzL
Om3TGzWHCht4AYsndH8zB54ReDXIZQE0SngDiTqqZ6fb1kLntLDB0cnu11C3w20iqiiOfBejm64p
nNBipdaYxNW7MXrwKqKXG6T+dENON9gztPBsxn+wGaRxAtLc4O93ROYw9VZB4ltbInOsoQKy14hc
xwhkX2If/eSN4VZJulAsVa3bKS2GBlwZlSLZOUr/ARyRsEiJwWP12ijHmiRbYx4fduucwFyNX1mB
zg4eH6pPJm3gwrXX5lNzjrYI5D2pvHRzjAwkEYbDYQC8pbZ5FGqOCAeI2AgtUplQWYuRMXQB1RjJ
8YH9i/BUePRraSy8ZmUBZbl7RoGIgRkL1R66xdy4JNFCcRhRCwFtWhAdsX5wVFKsZpwUnf+w/jaa
ISKn3t63TfRmo62otQvpNaz/a48zzZAVI0jGz8FmtdNpJCZQdhui9KYODMHAKc+K7G/XkzWZfddS
uBPDj621I3SXxxVt/zh3rKyygXS5pfJbj/kuqNvqXCRj4+wX5yUSHzz1sxm6G2weeD/fPuUDPZ4T
xXK73twYRcgafnw3bmAWV6BDu5cjQQg8aFBog77+u5e7sro4QuJLBmOMm+PEsWpN4UGhVAlM5v3S
06y4tMP2yAbwIlB9CIWkfACm41Xn7mp4z9nauopVeqlFoh1FyFM6RELy15///16Jyhvv5UsNUQCa
9JH9UxbeHnE16NaEaK2ETg01zR+pGtdnFV6BD0QMdHeKEnTQiFXiuQviEMt8JSWUtE9BvxaKZD32
Kxz9b11lOoeHVfPzSbF+YpczTwKFvaZYKkRlC0c/+N1OY9WrqDOrmrV3kHlG0x0V/TvCFQv5Mr99
Z09kbyVff0HvCacm6vk/dmxwm9wPlJEXlrrDVGs0DpTSviaeRRm93m2qOjQ7c/KRUxDxy3ejhPqs
ZilIlRmN/Wu0J/3OI6kCqCnCS+COKDDh8SimpLXrEJ4QZ0pAPujJQ68edtl1gTGD2mpalGgNb7Wk
hbQuVt++M7QDttCUGSo5TOkhhbw7rs25ZNiZAHjyRGC9gcqv0PjyZsBRILbvPBvMaVEaEOJlibyL
9p6dmq5rRptrUfFr/ZP0JKeOMh+1MGIH/dl6yi2V1aMAkgMODpDDXrPjSAXmj8O6nzAJZFFvNGUi
2/w6wM3WnvqLit6S+sPR5foQsSyrjIfD/br0M/IrEcc1R0rCLPI18vH72EnzN8dBCLZXbbznC+oI
/37Ezbcu4TXaY8XY1dLzva5i+ScYHqrSx9ftF34dnHZYUEYrM6fKJQ4ytq2ccZXTblAlsZ0W5Tgp
hRboiAWz6Rgudf4v2ZqO0IMhHXK5mmiUkhotRbtUiiK4m52OhR1/3yk+vczb3L64gH71fFZIIVb2
z9XGwngeV4LCXONfXdD8ThbTEbOiQfJmm7DCKenm+gCsctLGkhGd3LIOF5vBozcYNL+oUeYF4Pxk
3TBg7n5OncJOy7MBvJySjlUsJOMU6ZY9X9y3KtP1GgXjFWMmPD3hy5Sh9Lw5WfFmyc3ZyJ34Z7wO
UNHTWFLssULuHDHoJ2g/Dng5JqJzEJznCGdN3afPVFS3+d2Maiz7v1KCDhUhfi3DMK3345Jotkmb
H70tUu+toTRs++yE/Lc75XV5d0y0pW6KeBH8m4hP2a3UoaspbTG3wiWRED1vTgZZeoC6oM9c3xOv
qM94451O+8qqHVUzhbH2LonbVP6l7bB8u9B8p0i8+gaCW0Rt8tVn9zqglxU8m9v/DHI7h77z+ybX
Bk0133lveUP5g7BOWlg4WjHbc1MMabjOo4+YYKNWaVjasrZoSOib19rEXO/wlWb6/KXPsFiSV29E
yZ01uj84kUUt1Owo5pfo3TsF3wU1ljAu2utMnwiq6CPhkdQZOM0yC1ijAGGvmTTT/JRwsxotO8XB
/eUB7Q0Fqh3YlfRNVf2PiRQZBJRNFwwv54vtyDaEatMCwuMFkGm4syyl1GbHh9BxarCpemFIetmO
ldgYpevvmrqsE9bnevZ46MrzonbGrKvwmoeV9ashdIWvnB2Q29EK4a5IFB9yww15/EvdtP4rW/Sg
cYMHUq9lUj+EK4070ZvHBCPrGPaHFiWUXiDV7TK1mbpU79qtJyWbhV1uRZo0AJYX+HBc4YX7T+JZ
zcjZurIPucrdkuMHRzIPFgJqqVh7DDhlN6ZvARVBFRUkrcqIlMH+OqQGVa5bIUHgwa9ZdFDzvdSm
NG45ceRRS4HA5KAtywIYDHe3U4xSvq64dAk8KaIg4l159wgcTl1+hpJZ2r0HcQQOcpXhcO+7nm1J
ZYXIYJT1wVVeQ/EgY7N9wgfXfbMkW3VjwznI2c2FZLB6diXWpNOxCIsg9yksDpEOg/439ArYgV7O
dWp9CrqpXVvybVMV0pkwMMzsrh348255fBpkgbQdcRG9X/tAGWxJ0Co9RZiTZFyInfknCIcx78RB
kfb2ZQcWYmy71Wh7/Kx0BgkcQbawpt0/2tO/d/1ZiGcdiQ2FidVYJ2AOAv1mkB4cvg0Y4a5vTTaT
2m+iNUOILtnTr20rBVEB7oy1A/Pz0+8rBXAb86oJkG859OmaBXZ8r8UXmoYQeDnKzyrYg+p+1oPa
BaHXbQncyVDz4NrVZPdtczHbWC1AHYsrm4j6GnrQsKjjPjN8FfyS31I9RXdHU9yLVz7e6qO5P+zT
QHYIYZsqAtf1ZQBOy0bkZeXe9HC9uJ0BIfIGFa9w7+WRvzSfUCfc5Ag1p59qVEQFoPT7WP197Mme
vcytlVMBghOak3Omh7vL/IXFH1+ZRXgwhK5pTfR8I3IWYfZ2DlCIqlA0i3Aqk1XLFdOuaFCaeUMg
htXTP5XGA0McCBqqscIcB9wE5ELJcpttYh2fmOIP5sYC0N23bwsrNxrHuGN0+++qxn/im/qDnEeq
XVlhsUhpoHW4p3tgqIYwLRAY5HoWA4QFDHj8Q+tNpthfGZ+CUsbi9L4K65oLUy6RPOP/ooQYrHv4
7kIz2WI1HD1vo5W8fsQn5Fsh+R4972cX2uai6EEGNW5DMWsygXRaa4jrGXnHjm/PoUGy+0jr53qm
4VQmzJWVUGWn98TyTftUJa83ZcgfOP+3T/fO/WFU395FxUYhlIaKbMhAOzHe9a59jzyMghq/mPue
WX5v8K3EVWLVi4+iviITCJoLvTMIyWK8cYFF5QdW+MBnyEgNXvoV42s6jxoCofHoB/HIq25cwZgW
JZN3RERz/WrqkTLjB/fHHbpHgCFa+HLFvmkgmK8stQAKgrx4XpfnXSi5PdYl2fJTPjJjCjnB+aWj
lb3UrvkxmM1tjzJ9xCtHuw6SmZxI12/lv+RbF3ibK5a1lQlBVJ/4GSR3GyGnhylxuf6DoZRzEitH
x2BKMy+87D7ziVBa6sa1mvP5vJdKoOuMxYph2mNcOdG8ZcSQMLXHYQ5OiXvhPOILqmEPpYCSsdXU
xNR7wNVPmEbEQuFbyQRKHeMqpORseKANUsJ+8gBhX8njhL6Z5lWW++zWDMV5w/sZfB51exUGQI5l
7NC9V1Bkr4IfQidhQbb1qJlEmHG1p2TtDbHkJjiQ8ymj1D3G1UG8ghHzP0xliiVAJxpvilSsUSCC
SMWbPx4EyZubY/pVE4/+PDLYkNQDsSwwlxdeZfrPvVkrtNGBq5AaZOma7fuO6Clm5KeiuxeSewRY
ncAnpInj6SwhKW0ZV+Tr4BgwOpP97DyB3QYo0kuDrFSx7XKtLDscIkm4cJEDg2qI5UCvL1BcDwTE
yNif90HPW8oA0zNauO5DZqcogEbQOQZepKg8UZM3ta5LEh9c7CBMNaCTIWIArRcbnZjQk8tJFjFz
kbME5QgQrPw+SpPAugLMJnYe9knZgFY8K65qACClL40YNUvDa2jZ/y5cRGwWCx14iOO9MoAYsxiF
Z6qMWa65/ER9vK+zlmv2d4fPsyj96xA+ovep1JahKTw1F9f/8Jlu8tbvBD3JBgj+1QBzq/lYEXYt
6GePgYfO4wsYJrLfiIzc2DJgoCBOsZFz4EplJmsnaaiY5g9cwweMPLAAfSnMTnyO3tpBaBzwHAWi
x3dTxEzKnxnfrKWY51erdR+aVO1pUXMT0L8SZn13HUslAIGgal/Jhgor47xu5bUd8u3bJ1TtFycy
nqfS2Qnq44qtNn10df123eiXAsMdLx1N1XHFR1X6nFRMDL+aKJ04aHieXYg02yXEkocTLVIS2HRv
t7wYS2EWetjevpd+3K3U+JruWTfi29TvlRlodXV7+p68F7OofJliB/kKxHTwfx/cmIF1L/Z0h9aa
rwuHDYO+9mBTjEHxRCS7dMiMjVqDlEp+O9kZvPqM6uA1udoXWsVJXDzYLmul0mj7Gvxsw1TME7Kc
vEZzeVVWJBexxZYo8k6QG729gVWW6h99Efd4MgDmpapAoMB9RVbJfkRQdoG58qlwuaLrMXnJN04H
vk0m6ze3J8fsw+nPfntGhRZMp76kndCNAoD1SVEIzb8SA9vn6Ha2tJUQYn5+EULsNDS0cBlIKsWb
aov0qizoxpM/oYZT0smGAjJp4TqLMwlVXLpWkyCpFY/GyCWCRY/Z7iY87l6WU3J2FV05e1GRwOnf
YETkMM0x0ju5ar+vNpgVTaHz6fuUabQ1K1CYC3DbNys9xuW3jX6/Up3MyQ1W/KLShf4oXR1XdZxk
DATQznOGSv4ghPSMOjzlynbNhRvFENzsjyQCZdAV4Jhta1VIfrMR8E2/5EvkaDz7e/82pZ8cP0jK
xVbtRjOSsCNe6d4IxZT7ChAmtOcEeNpIJO1P3/7bI3iED3hu0DkQHats58N18kgL0c57Jc4AvqOq
kuQpT6Z/Ruv5Qxz960Xzvl5fHO8wphHpJIoLQLHbols5RNLq7cEfDHfAetkBOUIXP1jRnxuDlr/L
jcBk1egjE2AZUdAqungJv/2/GzPbz8jGLgBJHCUPHbJw7XPvXk+nfC3a5MP7JY1daLv9Iix9f9av
c1AeBgKerp5eNfw5mxhjOMkgHqaCXoNCK95+nieEIo7y0P+oAbXtNng34vBTYBdzE7TcCifWoXON
4adTHbK669GPxwjJlAjsgPnOa6g/fI2gDeD/a07+7qVm3Tf3tE/TPyBsmZn/2Mu1S6W2Hx8s5yCM
bL4k7Sz2py/tUwVuLt9HYqJArjG7nmCEna5rmuQtAMueV+FtH7xP11e07UjwA0KG+zgBG54fSn8U
mn2hTxzaJUBquOZL70yz4WqzYh05q3oO8HVLVvB+444bE7Rjk/MOtj/RdeCVZRtzoVp9OvdQVruL
3GgiCdigfc55V+imV9faKfLPgW8eZBkMdUnSW9XDDX+Kv6L2y1+28Tu5napNP+rrF25kuBZzkHFl
TvPkt0AFR+A82rFn4ip3YlvC0pGnFI5V4DSepiwJBRBhmHj9fKYTYIBR/LodMhSqZ2q2+fjGftrc
0GGCUdPMVgiV94SaozDfhtq5qdlpPeAtWMyj2rueQaisCmupm3R1xgczk8HTdTsvKWCuZfbpTsdD
20Lev2EkeR5IfHmJKqmtOehapOUJ6y9tiddNVW8ixryQ/lrNM/NzuxW3qVBDzWwF1X77pmjzLwb0
WVeU5U88PytPwuqQK2taoKzVjrWT/6J5t8XunzT8AiFdcDMUFHnfnpmfdnDMhqxqEBxwVHjTNl7w
PMxIjzgTMCiA5ykNqE9JrpZrxQjXKoT4kesPPHwZRQjj+0QcuAbien8kraVFgmZvl27wl4V8ld8t
KZKnON+6Dle0/nAab46sgmtuzD3cbT4MQT6ucKMfcmnBSuf+HWS5NsQqJyF+oi713GuReFXFuTJ3
ee4KdHNMceniLoIzTUCDqD4HlN33+VuB5d+rOI6PuSrapHna0d+JKniBlZ96oFKeFrEkLgz/maek
8brqjwmdVziwu5HS7LxfCCYy9YLSQAdHx+7svDtWgBtC2TtHqFNjDxIvwu4Rq5CDCJGVAU440L7G
f66nVKQQzuZbYVW+mrtuCb94qKDXngxu8zY/ka4vZVmOy7AE3oal82gs87EGEZqZKR5OrcNAw1tv
R2rXQP8vQxnyq6TA2K2Cr4TACaIxryg+71QeZkdGHMrC4EMOkZiXcpP9ZjEPEnHagQspvyO/J/Ak
R4BJL8lwZsKcJvZBDRQtb++F6mL3Fm0Y2YHh4movyIZTUL32Z7Ztb0nOWaiCUtwOALmBrr6lVGZm
rstJHK19ero2M0UAuL4N978z2ULm2ehwUvpc1KVy+bJZpXmF6r9uQoslZO2X9InUYBXN0O8kS3/p
/mNia23szzSDDFspyvgpCp5lYoYE7B5LYuFUtE3z7HWts8ItGa+mLr9VIk8LdCMKTj9LlfGmkhCe
OVla7ouFP9Yj4tgvchvT5QWD6dByLvVEEATHhhhLypvyT6hQPojpMCb1Hv9z2sseH7+ny8C7bwjK
XSI3jc4DYJeVmAX+DWPsCrIaA9QtMK47k7qIKdcXJBInDf89FDOrQGJRqKN7uQAFPDx5njt3eFu3
RupGG0VfaCUO5RPh3ufNvWuap5tqnx5IT2lYUoreDerjyzrkqRwo3+YlRcu288Yp/XOtRjUUNWBB
VmVtVDCxmBwlGbDUceRc3Uu2VEPE2/ihzhQ6BMAKxMIQ5m9b80qJARAxAdoQyFu+js6MV1LZmZ/t
QjBwZzP74Zxh8vDxl0GF3uqMw6SypivBaYappIgGvOwdzmRBW9wetmSJqSRQANBDW6MzttR3k7QM
5k+qr6ZsOAW90jYsmV7VZEHNNW2schsLSDbHuXqL8CuycJvQ9oVknDd0sKccaH4C1K9xLiFrRr+X
/lJkDrvFyO5Xwf9/Snn9nDR5/oM1uFV6eugduF0hyjMJ9fYJCT8qxTDptu7cR2JwNpNkVLLfX381
zox9w4MC+bhA5FJ4W4l0oPCSCMjTGT7UrVkzers+PIV2sZH3bMTHUXVkIuvLKRxQKsVhkwy31u+Z
pO/PeUovZUgtcHGxZVvF5+KS/jDRnf5cl+1jL194udpklVQ3ikJNnoUy/k6GX1uqhYPSz5XY0gr4
aVVEnPPuzqo16UCl7PFkCMl7+5tEs3MXevibcviYZEZ0Hj2poUoPCFqm3mQ7w7nT1sBgYSfSMeQj
ed7teEemswUF9tE86AFVPpJ9RTZdDfG8FdBkhGls0NNrUb2FUGm9xGnF0ZKusECnMXGSZGdmyQvd
wooCU2cpgwS8poE7BN/W6NGLW4JdlnQwOhwehoE1Eqw7AG3q4cK/YWiGYKOc5RkYWKr4WecYwtND
VmBmyStGZYe7sQisxPJYsJYEyrzFCfiGfSEIvN2PKYGRnK7mCi+Z4iJBUGKgxwLqNm+kl4xZUOZi
lYXYZqLzi524HPoEE8UwOE+ME+AUKEZpAb6PmhSd+i0xSexBMibx+4ga8oKM3awLT31L/SI92/Fe
hmkucrKEsoeaQmnpzw4zO+frgWqlg9vsYHlxVo1J5IdSUPRvhOP4aT9AS1NoKrcplGQ9TjS/iddY
dreGQP3PwbO05ksf5plx6fpTv8ypoCTnpqlTtgBC9mfppptiM+/PP5r+vE9oXh6T492JFqxpq0yg
QukZHdv+aKqW5saG9qDmHeZgIqbxQ8jFO1NBtMkJjAwj5DsOlEil4ZrpUv9trhNPNILvZqf/0Bsj
7ZX8tjIhLUV3PdGpUiF7CaCP/5WK90zwt+ZzBTiIDHc3sm4A0d60YKhAY+LOrkjhKwg/Xpelx0f1
OToQ/U4Dz/H0bUAN2FG7wKaZaapL54ARQMEO7AbT+fr17dGDHAdCalA08GCepSkXanayvOZ/hC5M
DtxV2cYcx0WtHhUzRXh1vCje9pgipGR+MQA0bnLPGqHVU1iIoYaLGJGA2eVLLGPza7f5iUE57fui
K09UX+x4zyqqVjWLRIf2pe393Kzm3iYM8AO3c/NDFvKRnNbgbO3DVfGFGhFjOh9gw8347VtqeNTB
S7VSiXKrwkQNWqKbyeby3lj3StG7AgwJPuR9qncAEnIcEKlL9pWdKqbUZUlSS0dG70Gla6NhDv44
8Q7Z/OMzBH8h55nUOiuhwzb0C6MluZyI2F7eyC+jf9PPdNe3lQgsAaAU8esjXOr/3s4Q6fOZTWuG
frsY8XcBtz2cgRsMFfNc8MNazUbmjBCa7DRLoD4R5aQn2WDPzab8teuah5z3u1tIfaoriYyG29tB
H1NhS8EiOm6DVk/P6jm+BX3F17utDL2b15Gzf4yw9bNdcLpOUNNDX7wyI/u/9K5juuqYjBST5c+b
vhmK1QDzCUCh9dWFWnrSBm0qtpXc+Q2H6hod/IYX/nTByL3YgH8onxkC1bB8EsIxx6Im/xCY6fvg
6gc3yrrZrSicBwN7JjlW/xP5wbaTyo/QBqywKI30Kl8XcdhV5O/B9H9RkDgbjifQxgzig+q/QGw/
67IxZHy7EfY1rCgFiyfcL+BDBElV32CNI++5zGU8Y3UedzxQtq9QLLxPBh17sldckxC+3WsvYzzY
xG+iW8kV4ecmm4jil9bmAc1xk9Yem2QOw6JzU1dwjlBwlLXDM1SNPYJNBiSaV6Cn4L9e6D+1pSel
dOPXm3qs9pw5L2dAor+LJsSezhjqWQlcloP0owFPgqarBjkYs4axCxXNAUi+vzwCbbnyXLv7f4Qz
zOMi0TQmvPOpA6rmTA08W38rFzgJXxKnbvyLa6rx1gtABPEXmK39GpU3Cg9EMSCe11GzwmE0UUMD
voWZlgOdbwTtK7c8EfkJ61cXFmcHU2X159B8uU0H5bNMoj1RHFa1LWl9+xPsbFJOaqe0KugOoS1d
W3fuVqJqo0dAgjWd48HiX0HmJd4oy19gAhcbzyQPtlO6JWQDjtcoRnHlqR4YEA+mouE+xk9wgeV9
mbr6NwzesVVlqxzygcsUvIdKkStYhHYO3SwNlmTH97MJmzkFQ8P3WCIvC7r4sH5ly1h8k2yWEpBz
bXpter0Y8x9zQP49ShAyujHzmTpA06wtyGzzL1XAhmQcEZs5iKd6nGjZOK3UoKP+Y8mPx40mKc5C
zDmHrutCx1U4U7MJDWQfFGq2qCikLXBMPZLj/q4Ms8ea0iBIb2iP5Y5fMhehgIiDeQ5xSrtSiOXn
SE2PPn4RjR3dRrtzYq4LIm3wmu6+odxJxjNgGdwwL6culNv12jc+3zBwrvXMPZGb8LGqzR1XutRQ
/f8xNC/1EaYVA9muTrnq5MEixcRxR9gHB1OniWbc5ALmR0cDr4d5Et3ktFrNso3zwGfD5veTLPaU
GJajsyvzBCixsJl3BosMjdnLRPGlWVfWEnrCSe10+24vkigOocEomC1J+fnsE5hc41FdirjMq0cj
tkR9Bp0+OuGAwoBohjWWVTtmK6tbWGq1Hc87NOM7fbf8Njs11hJ516iVtABjV6Zz7alnYU6O8mtA
o268rMn8BXcyLiNI2vBUGbloC8A4iAHo28yaPi25P8Ap703vv+j7sGRpXfMUbtUcpsskJ9jVt2sh
GkeW4QGPbmhIpysQRZFr2C9J9IbYIPTB/VJZq5f0g63oP088vDJbP7XNbXw1InRbohbTiZAABTQP
NA/IfHpYXQ0bvj6hT/hDJp08Ll+XZGYau9KrZPZ7xEfY8LD/T6azeoWNIu6tcLa4FRelLHgoWwLq
2eOmml5Q7SuOHK4zLe9+fbWHC8xdg4sZaF2EXtHhbmIPOPCaqxZ3OHs0CBWjpB7AXcEB36wpgi3j
LPSuUIpXCyAii3vHb6wOtmhpSixDiDwApraj16WDNfU8t+7XJBkpKx1A8SSBRFlgFb/Qr8ipcAq7
CjYzht8PWV4XoSzucRCr05tlGmRHLVH/enX8E0oT6/LB/A9cB8djLSILUGZjJm0rLwdxCRVTGFk5
CZsTNzjadnqd/nZ0rNiJ8zVpOth/oEjrGZg2TW7vfFGpfNR7I9AmiBswwVuHOctuN7J2x45dwdd1
HX7CmQVepYrnfzVgBa5LaMVOKFZhG91+8Cvy4ZtbWcmUC86Il14I74+xjjTyPHyP2OfCEWErWyoz
fRxo/yj7G2bLCdyAwWJ5VaLHbnk2bFi5zls3JDXDdty8kdnxN90SD//A0+uruYQ2wZOXphfFaPvb
GXdmasq06xXbcxYMKs/K2dJhAPe3aquP6fOfZy8g5VcKN56Azz7fnkrDy+hD1o0RMtuga5UbUUc7
hfCnwCm0YiKY0TkrGXy794W/9yOHdc2C8gD671qPZh0uqQ/dbPMkTD2upF5U/A6S7Nxi7wHGJAFY
NcZf61Y918vqCiEdTBVOSg2AZ2zBMOwqxs6kDz+xpwspQ7z1ckRGCC+Gkx7/VK2+v46jzg8iC273
khWJ07KRNcs7B46PZE5yFE+NETkDtH9+13G8FX2ANCKIvLix1NdZrGHhP3yduZiC+1DJjBaW+TKW
NuaiVDRV/k+oUkHJyWya0AFA7U8Nz5H+110Ao12ADqjZeqFdAx179wUdQmR6jJExrLP2OBw3z0Ln
LmXIyqNtgR+OG5cP1rtUtqNr+7SNg516Wnb3g1IYUet4+fjZ1zf/96SPe3/uL0QN5Ofi626c0pjj
tcAYPip5qkXDdGqiv3SK8j329aVwHgr+8oGQBPCz96//4fSEQzskH0icvXrODUBwWY1af7gecTwZ
ZohoO81saSYaNWaD4GDPbGUYTS8M/BKtTnsZ64JjZTb/UDspFaxACJd5WDB/4ZbxlojjvIYEfy1x
pMg9jyjQOzzEk2PgLCmv0nrBqCN8iIDSnUUw0AKEPpm755kXXcYgXWZrEKAKqq2vO75H85K/2L0o
T6fBevIdUg8g2sgpuL/c3W32hmn7feu3OyEMVm7877jl8VsJBzE/2mnXSiP9RjxMU2T/pAKTeJ1Q
GoNJ30TdQcupvoQpqPHrbZ9TOy/w4FziPefQbtro54+4NsJj206ECc3F37JsiHpNX7Q+Rl+L+AD2
JPs2mw6urO1SZ2tGJPoG58NSYZbraDkzQ5ftZr32wQQwhn7r3yyYWZKEE1HSUA1kTcYQ9QSzL9B4
ijPc+eXZwyN6HUVpe6x7TrqeJoriwvzr5MGXgZ3aDdllBL0vl+JGnm1F+VNihU9S3DPzVdjNsVQb
Ry3b5pH2L5dqbUIWlZVxK+2FB6DKJgSQyZ5p4QMvaDG2X7YP0HXQEDy4G/PBIgYw1Xe+IEAs9TvR
WILVGdRA6eW6SAIsEOj6F16WpJZ5pH/SAaMkcY8xtV6bkjrjmbx7s5u8X3asdYk8bssjEga3zMr+
8sX57+wYa+D0RzDmgbfKE4tmhp4CFws5AtpOIkFFJnkRENn9JrA08nHv54Eb6F1590zczrFvqp8a
HOfijqazJDc6zJ0p7pX3eE2/KYM3+orCrRnI1/pThIjBsxckgpXq5KFj57AJWdSRRe+9I7+CNcm4
ocKo9hkC+FAHwHdzAU85BHoQsAgENvYhCt+UWqU+bTTtXlY9BYRsdufzLgpP45K/IH7OSEqqJXEr
chu4/8C1VoIdyR9Wm69sTTBl9I70z6+AvhjQRL9XvGB6llODNJsOCOLNrVs5GZmqIc16qN2uydZr
hn/fSHc6W3ZpbjtsJJH4bu/swkaVHdG8CGcqQc8zKjThyGPvwoLkj+vsEmaWBHIVBcrNhTBw5M3a
AzANBKDqGzi5FkWCmAWlViNTar3kbqFQiNxmnupAXqTtx40ukkIs376/5XvR4aMl6h2ML/feouSH
62m2jsEkISZ+lXUn9jd9TMHwua4kiymti74mCMLdByPNV2wk0ZtsBPdWD1xF/PgAzZ4ZFk4OsQ1r
5T37Lo2Z1WtzxuvHxKFc31adIFuIa6wdD3naEIfwX26cem2NwG52hPj0L9fsgSTl1W5upTrXXHhw
CSSttjYdbnKXad/DB97Z5EpYUedqrhropKaTTY83GvJQDHvmboiXS1uzZAGpTdvVDEkYgcyaIASG
QewzsFnN0msmK78x85RIF9M94OEyNQh5J9wNhCKBwhs1v4AbimuRFQlIFy2LAeYp41+5Tb7BHrLY
ywUuLaEmG8LxtM6bBwjMgUPzKQ2o1gE2kM34lQMivYViShzPT4zZO67MuTYPYC7yA0eugjZutBL5
xiCguJ7OOIiIM8cZO8NBWg0j3/0uczEsCuQLVuUppGS+Dqj40sOwbRashqAhPls3lrB/OTN/gdur
97k/KigMDCHWqc8Peb+AJcrowCVnt4nykk192Hzs79o4ZN9YBSp5k5Po8SSLGV2FiiRP8DgMLaUb
3ysMPZZWJfjUEF6fc8gRFKpMX5h4oTptemX4a1VgKQSKBFU7Z2u1oK+yWFUSz0bQdzoPcsLnnzMk
tg/TdHjj49wzP31QVpYDjgFQyC+G9QQMaUMSBDSOWucXB1i5IGIQ8JH5E4rJt+G69Wh6vA0ZLl4V
3UhJ2Saeil6MeHzU8opsVfoAusYmAcqMdEXt9QfstzsZsc7zXBOLF4f7YzYgj5beIsrqLf2gVcEC
f6DU44yVeBKktuq53deL+gCrcFAaWRcnW2lvUkz+pkLsbW2dTa1e05+eoBMORTMESbKgFSD3vdk5
P10ydBRa/7gLYlpa0DZUUN57Ln+9n85hUFeiTMK+cXg5ynsQNEdjVT+SHWWM/EHHnbwJt3R9nchP
WgpiS9wsBR3DY/dqKTMmegOzIo410MYDQta6VElLFtyvSQhXYBFBYE322HHQU2eKPDcCJySXyofV
x4GZMzF/4/YYSJ3AUydvTsTYCDz7/hdPSMZYsgUOssnE3F0KlNvtGmyowgyUkerGkoWh3Wh4PL+t
sOVQpt4VkyGt5XjVXQPCrHbzQ/1igPrqa79zN1+k6JT4NROUl2kTIn/QY9DFvwIFq0l2HEY1gjRU
BamyiIkmHr9B0L5TrvNxMKTSB4PQaswnsPzwYPTZmFgFzX68B9KhyPWn+KxuC/DoxlONFvDmgPmf
iFmrrbgliXg/BlAxx9LzzQ7ZkEh+WpFjdcqG9eR8CmZWIPE2Jy5dEsxv1HLtUzyWp62wXSVYVSFT
udXTIpGs1pZe4xcLP98P/58tzZsiYToC8D+E5RxzenrTgjGLtEuaFFffNhTMdOXTywhiNagoRlZQ
6yGbpiUic9lXTXu1mzOIy4dcibNcImwMujJ9uHZzhNjZeqnVlWEAoBnDGem41zBoX4C+4q2umRjC
7vfZl1LOMkzh0mozvHR2MpN2PZZoYQYR8l984Lb0ZKSC8s/TUDIBGS6/z1c68+CMWhUPPf4oJKip
NaLnBgnKILdpxhAtzFwW6ZmEwobDqY0e5m8F4+Hjwp1Rwl5I13RTJRTJvQxkE9iD/2Ueu+jkSXFF
/B6w1bh+OotSZ+K0nHSNllccXuZOJHhQTGMHHk7WbFhgRE60Ndn1TaURF/gc28rk1WO0i0O4zWI2
wsmiFoZ9LzcSfo2bvh4DkykypzWMvHadtUI5S5zwLilkXsoL+a8P3+PLqsK0ysAIBHwGeoQX8EG+
6+1IO9n5inFXSdvrPnri4qLpU0iRpzZzc+ImOxZF5WjH+oXbV5gJt1aTJlt9iw1isX2qfTBvXBJ1
h/jpn5dATESsuPgBDI24wpJHQO+GDyN6o3QTKKH0lozhPb4Ge+gsCvLwSGod+tctjmBvtOoBaDct
Jv21kXiACIkAQES+H06dDpx63L6ypYLU8NTXnZqLy1WTFZipKrWbljBsX9JMxdd4zGinJSnzgLac
/499URF+uEDgo48KMNntX0TImQ0y9RaTqcbMTkXJFLmZ3IkcR0J2iamyz40W6LKm89kcvkyNgug6
CbSWTUV3pSUvU6f4OtfFc+byOZ6fWLad494564EVub5oBFwabtcjiKW1t8LanpGpEbf7o44msH1C
rHksbgHFQHtaVjyFK28wKKX4Vng/1cXnw6KO+YRaFl0T1qhZIUs/Saw13fwqpiwcdipFhEukM/1m
AiDa1/b/MXAB4Brdx0T7CT52nuuHmDjzt7vnhZdTCbZxxi/q/JJU6YgKaMZ1D+5zu/m5Q3+rxEj5
/e3/Zo48OklGOvLRKO6Qo/X2Ll/FfzrtrAQc+myM1sl5SNGKi2SXUKRZnFKeI9Qc1PKbrbKGppV1
2uEvVRe/V4db/QOjSKdLw0l/gNVQ3yET9EkT16wehC6J4WcV7anF5lxL4V7njC8IwmpOHpS4Kxl+
xt3v8ZXz+7FuLi1O9CVjj05dRPvmqxGxKH27xysPHXpq3Luc03ANEvI3WuzyyAAha4wLsnghIKTZ
kNEMQjorYQPaI2y29LUK+g9UtVS95OmOhF3QD2o9Oo23szxKtyRcSkY1SCJJF1biDHwmWQGpJkEV
2lVdB4ikSXJkII+utJGUvWiD3qHm/lGgCg5n0DAo9vvtW7CEQPAitowIRoln/RVetniUGRjA4CMa
NS4sqeZbWE3MnA1f0A2yNCHe5SDhXd/URa7fiFSjRjqu/PldDzohe//4uOcFSDaOTMbveoT+jxXW
na8i9DmmKq6ZdXVbPn1Rn4N9MUi8GOPwhoVmKEsFKbJtiPj77iOftrLZLpHTB/Cv72RE/+N+XGer
ImkDrvQAMh8KYnOoea7deMEEk4dzcoxt6VN4/Urb6XxhaBKVOA+Fd+cnGYT818OysMNqXUrmUmnQ
sSz7UL7AHC6VZVbSGEusTGhgR1eDjkO0TukmaEUKLqfqnYDBn8xW+GrVqHDUcMLhG/kN/Lmi3WGN
2w1OWI1VP9mb1vv0Rxhdbu2F6H25/ZjGzZGyfMqdowj72NzvPfQ5k9Cq1emIoCAzyTWfJdYlmSca
VKQ1YkNleHvVvxjngnZr4/Kww6SLt52Z5JGnnWfUsfByXEjWG4slWVjswa+N31FKR8sHQ5Gld78A
6qp+8B8Ps1lGCoR6GdujfJN683p8Rp+lQbBLygEwK8WHWDcJK9wXiSluIZrvmgZpzFvyaTC96dP6
8H/mOR62Yr37fjfU9hzP2yFpuC1R8pnzWrhNANMchKV1Gb/jHBxEdP38OIJvkNShWJ6xLsMYFY3r
wCVfoga5yw85+PVlpa7c6GmRNwmrfksYlemlCRUoebc6t9XpvRDKBH4Kkh8Ntn7tuyO+g1YZitWZ
QxpVY0a1NfXvODsuOVZ6CR+KnbQLTqlQeA9gTQ+3MuuhiVJPhQeoJwjp4VyKW2X/vIPrLml+lBcN
SpurgTIrHIoNwoKZ9VGjqf3FXPRcCTseau01++X+KDPVf6biY2oSSOOEbDGHHY+bCiZyrOJ0qePJ
4+SnWgdoxXhGsjQM6zdniHgpnQtQ5Ny/KajNf1ZGnt6dt9mt8wQUYUX0+Ok8a3H2yUIXDxtzXP1U
GJg4vCnKXuGmJv0Jo1zlJnUekBIgJgBaZjghjzJO4umVnYx9skyI7R8ldg9s73QMpZWPzBhQG+Ku
JQ6kPX7OyTxGFpgX6sp3DO16Nvn+QunOyx3ozYAQ0fgUhve20hW1jC5xVDNEPsxfSJhIFewJM8Q/
Jiwz2peUYbo7HwCQ8/m+uRnVSpQ5ZzFv3zcCNIQ0kHXNuIqFkQSrfz1U4bRfObY4XFQ2glPXETdT
4H7nXY9vHXFc1+7wUMAEhr1dxdsK+WRHT3JPP0X1K07kqGMCbhwX/iPeoaNf6wZaVqxrgvV167xD
I3m+bMNXVwIvYRoREv2NlEc+EEs3VokMrgU+NNcEi3xKO0eLCUEDd8hFdtJ5tGIaCzPDVRkPwnRW
WOeIfVlsBgcOG5dLIYh+yqlLMKdAA2UAtBc5AO+tbU67sOSveSl73Dxf80JFqG8da7v6m0xjI/eS
mn8sDEIiWge/osH3DFsljpP3W+/PxHlaue/erm5iR68r/q3URTvackuOMN/OiBv+FB5iTwN3KJj2
MZdZ6cxd/cfohkCBagd/eCXlAkWBEYJvFv8Fvqdjqe7/gUNGXJ3DtJHsyWJGIRVNeP9eFvtjSQrH
6ldlo581UDlC7fxC/HD0kZJZscH0pVcwLAtzADeaS8YovtxbjWaOp900s7KdNaf2pdUfnIqBWKkK
TFlOTDJ0z7CE2lem6eg05UwPd0ZHin0DuFJokmrPt1E9U3BA/XXwdqaazBRuxHN1u/p76+ay11hX
nMapWbH2AbN5n1kCueRhJfM/WSG3XLYUXBdORdUIV9wMeS6hO8jBZk6JJV19t8uSsENhHW6L4JlK
Bl2g3gfjLP2Fdw/PHtxJn8apdymc+I48x7XMbIWaesUOljji0ttIRTaTTRHG1fIb5qrYJsfVwSYT
TsS2o+Md206VhKxXuCsuHkEKUQKZdN9EVhCFjMv2AiUk5p4zynvcG51dVoDqhUnnsoWHYwV8bbln
aN9CSgyGA296lLuI4RBBCi8PdcqSuhzMbe5zLHkz1PU+9+fw5r6DZvWL4WqinpQC3Rn/AlQQtu/K
CdNB/STQ52XMaZeCllQbNPqRY110o0p8g8PurwC0Py3hwFcIFzHNy6tIEYNtnDT3LPG9H96FyrrU
tc1nCXmk3m2179qI/WgZwNG+FlkU4b3U2itXL7rfH5k3z5GDUG6oRzAc7+lxgM8EIJ+vr/gFdn4w
zpvQ0+eTMUy+bZzkMeNRury7+iT07UvcB4sUfEfBHNXswkM1RLQ749LIBODG8Ym7Odvrj1957t0q
WHLDOOaR2wtw3gcKjrB/UUMm1Rzf8M7X/bpnEJAOQR8mPgLGZkNBWAyeWVJja1WB5kNp/53j38jK
s3+6v8whdzR4lUmfKFnT7fNTXWB7PVkm00W7AmiObAjo2NO4azDc74u/bYzvPfgjCEhpCNj0wSPd
aiBvbtfERXTq02rW+QGWVrWsR9nyvC0xyUYx9iumMsKPeTYCIL6Mu1rjbXv16+94LglvzIn7oQBV
xgr2g9SwHHHUT3ck0kgWD4r6bjTTOUwETFM5GrhBqmF8kQKwiDYttK6JsQ68XuPhTKzxO7CV+Y0f
6MZMX68aOTEWE1ADU0nj74PIRGtONp3I2yeIjBj3Yt6rv1NuGsZ9U6uxeNjnkYKAfV8HB+WxBW4V
CVzZYwpUXSP2jAgdLld1t4S2Z4TVPgVpav3ZtT+NR+JKVcIH5yneE3IsiYgO0qrmrNA4JCDSNo+p
DP+s8O0M90ZmdtkFlTHCGWGko+rMSg+loFZh4/512/j4ZGSwvmkrpuvD0ybDrmosF+MPQ1x5+IgR
deZsT3HjMEBxGI9lDUwgHEAHeDFJmFhLzN6qLA+s9XINWfe8Fpfw8kUKGFwRbh8AI3kP/Q0pM7DF
hq2Ni1ouGN7GcjxH9TfBrjoBOV9JTvmg7Hr2w1SK2hTnSPkG/6L9eoJTvyr6lraAQ+er1y07RsBD
c9vYiURPtVutYs3mEk/TKJ8aK8+E5ZHQdoYZf/cAV+FhELBRxI0yO1E1jufqH4/2o0kDJY2Ex2Qt
OxilYGBGd90i26go1noUtPh7RX0i9PVe4W12kbzvfQNOVPExYiHPBMnqihO/h4udXCjbpjOeqpsw
DliaidmS3EPPP1+7tiBbYeU+C2DrIgIOfF0aFZbotAeqXR37VdO1eNViQGYOZGUU3A6IU/5iX8tU
bnFM4yOsdvKwQoqwzPi1m7U6SsZcWBsFmcIBRi6XEPpDtlt2VKA/9gKTi0wuD4vWUICluHEocW96
tPaWKXNo9fZJvKC6esGwgJ29ncH91koWXdQ6k1YA8tkZWgt/ZpCfLiohKyxyKWWagVwlPNu0i8d4
qn6KpIzoq2NlKaXbsmlvDO7BLl3gqvBozD4t8GSPK6GwVCoMt6MqoPP7UcEA7QZ9V9vVdK7QmVNa
vPxYSsd2DzgvO+BxwqLkHer7aus3BLaYQ7qRxMJ+lCNX2txjM6ONL3DUKSc4ooHSSLzjqHAk9ur3
W8XiPZ6mCfnmcjngtPdUafGOA6eHYyJu5OtNyzjAWkUpUcSZmFyRc+dMWnwYJjcl5bRXE7vjROPA
qIUi9qM2mTVZ5mpbiyY4plqpVRqrQwBCYE8byTgcnsbNb7uBmEFJHA8A5p99dOQHINoELuobyL3r
e/XAVmlLFOQ66x4aaNnK5ESmzc7wbWxah3zwLiOcBbsLVeYxzAO72AviRRPMhA25lJtuYqIVWIkT
Jgg1lbU9oMchyO7tfL3GKy+bw40aAe673JYhRZVdLqHKhgASx48qtRNBv7Or3IBa9xYSMGLCc/3+
rzFkOJfQ5KtLwQpvxg+6VX7Hfa3q1Iawevmc2hXYDozQlTTHZabvuNvf6Ji42M4PVcSBc5UNQXTb
LY2ILR2zyzA3IbUtHDD4T4ukRL9FAvF4zoR+adzc7wbGmAH7OMecQF5Ylqgv1QswvOgJr9wPc1lU
KXMlbAzAugnMCbYfujcSXRALiXsr4fccx5qVDrdFdSta5VFpw25HW7rP9HL+zqdRl0IK4gwqlRnM
hvWAFRlqlz73gCwUi1UkXCV3ZAX8UpGHgQh8DE+R1rGaAX9CwxsnomQ2twMPwJtBfKTROY5/7i3g
E1QXPEwD7Cl7VB/XlHht21NDAezOTOuoXcFcthGW/sHYwrGUfIE+MZvOPdIAQe96M10QbC0KSNFh
g9b175diJjUCgwpe9n+667OeB/olpOEx9utnaV7W6jBdBE4+xFNmTQAvA6Wlq7KEyZhiXhyAxHsP
0O8cSvJ49mFjHeAtuu/nhf97FSrtaF+Hf98UlcMW//t4XRcQsCdm2kQcTAw0Lv2woRvnEIZwZPNA
5varAE+MYYS5Iy4lFQs8ChsvfW6MZeYD29sz6SxY/1PnMUJX682CIxP+FZ+qL6F+ely0tTzTb6uO
5JjvVzf+cW/T5hwYdXv7L+ABLfpZnr+RJVgdfPh5rVhzSuh/TbtSvwYkpvrl5tME8cwF0WOFVjz6
KSgoF/k58IytJanQsmRznhwhprRp97pkvXLBRA8FV3OJnoVmPdGoU0RH03nE9PgH7hM+eHtisXY1
pHnrAALL1wtxEPfYSLeID4OVTDKXSDhJdpimQIxKEUstHctPq+6BU+7bJXWlZmlfAC3sG9WL0xZc
y3sIhikXJJOEkoTOm9xij4wXvTef2RIsO9aRLTyIlSQTiLbP7fZR0eTc7/Isl3yXKtJiLTTDBEFN
kFwJmMUCddrvqgFU0VwpA+3Dmw47LVvL3KW1yZo042+K0IwFvnovniplhDPpYDCN1u8P3ytD6JGb
Ai5WB5a+bIATC3hSGqZ1FWkf75I0ms04QnW62J2xMXh+a8JOAyW+Ey2BZ1t58QdRj6Jtb1yLLFGv
Ys0fhfRppfJjwxyJ23VFR2oMoBAlpMRRksKOroKU9aefy089EhxslfCb+Oi6OtNwZvotL2nbe8FL
V1sPm0rDON1G4RCOkTJ/SZ4uUIpkUhJ/8HGX9QmwBUObQYcrS27lJCPt6adukq0Hnc3pTYlXNVI7
XjsRDjgO2usyIXGo28WThvDPetn8H5EIGb6FGlC8+1i4WyFDixcIVMJ98pH6fhBOQGFjv9ROhuQj
KC28AVMX5rDPjEKHr75qpzxmoMmwG4NMd7Euh4COpi0N8a68Qpx5G6jwN0MvnZ7grbdgL6JQhbmu
QZbn4MVmG+MdfdczDt4ftuscWTSfwaBH2R/8WwdJckqs2symdpEvfoXD1/MgHnsawV1vriGv7vXL
sdQXk4NmzYwDm7PmmSM0wBzYN/n97Q9bUSo8wcGKMNOG8dbnFG6Ef/eRVPiae4YK0dGIGMp3AUaN
SMdvYcq4OGxcLpbaroEgQ28xslVE4Lwqui5hNls6dGQmHM5vvLg2v2DjHXO09f3RV3hY21BPbRz0
VeFUTCmRuhf1QBUvIPFNeTizmR5/H1nLPbBnFdVBvzGALLMNiYaw2QRkb3H22EqqGhhMBgzxjI+f
VGAb43FIc4G2qQ5Cl9ueppo6TNR4FtMluVK5oKg+5MK0t7bWzLB5bD0ozsDFDIkAmcETprVRCI0d
9SNtUkZ+J/GR5NHTxxX6RFClcNl5c5vDzdPmI4C462ykKsv+WtVw0jzmbB+y1KlYFjLa9OmqEQrM
1hrZed/oLTNjVCM5aIu1IWqlXi+xZmb2reRmLCzV0SvpAF4VFLie63De3A+vOlnzoR6mLOR7+5c2
rLu8lzuN/5m7zyTQfJctZDcubWeT3tkRd4+jHcpPz9YeNMrlsGFbqxgyTVAr/It6bMKHikMvUBip
YjxVkma/zVeG4BaalZmaPw9jWkhWv+ATZk5vv2hqGy8rEwr5IbtjC7hY2lP2K5F0np6mfQw8+6O8
4KMwmYSKyQh5UzJFhjQs0vgyZmQm13zxXE0g2m7nBk4AdqI9UE+x3AxmRBo/N8yLpYH2YBoW1Hks
KHWbzn+TMfxNyW29RfkIpzDKD4U81Uirrnkh4lPicP4maiykrFcpefpuOKD2mGD8LgyZHImwNx4C
rNCcVWizIucs2acqclESsaUKgFnVrTczC6V/XXNE/7g1CxT/VZou/V99klX1vYVtCvGGdt55zaCC
v4kTFXhWhqoCGx8h3vpEolriM6IwXBNMZ7YtNroIBmEeKB9Y2mD5TukptGlo8gdyLbksJIDMBzFM
rjpczyx0jfYFwkNUYf9aO+/wdqP5lZrWEIK6TgFT8G+dV3iCtQX8WI15Z144lE1Tr7f5AofZi1Zh
0Cjkmmg5a9UXTMOVaLcb3e88v/b08txEewXKgQrvoOy0wjhu4hzy9haoTGTsKnKfU8Nd6+W3PHBm
fWk1giwOnHzKWzLS6ydBORp4jeT6+zLKhVH+F0XgsHLU1hTDmYNGuA4539btEIGUcPNgmCgIajlM
dybz3EvTNzyyD23q6zMWP+ILrkQXSvgRxj6NRpYUv64NmMzTTChy8mNCLeODaNI4BYHtx5GJgBUp
MME4FvOiPJS5ZF/2lFCVJi23giZpEL2hfgSVU1OznPwxxBaSULq7ig3SQesiOr9U9I0PY5wSKPL1
ELxg3zhakFpMRWN7/M28RkOLQEp5jzFiKq8zrNxqv4gD8LnxOTM4qTiihZiS5XlOqOVcB0erML2A
Bn51ywkiy7pdDygL7i8SyvQvSFRQzjMXkcknwGpNbX6KDeAJQSYu0B30PAE6EQmfXsNEpLtkIu4t
p17+l0vX5gvjTZ5bizbD7xF8e3ouwlryMEvECc5Igzszm9fWlVGvNUT7gO3otfYBGe+9a798DcV7
1eN4UdRAwFNM3ze9Ig1gmaz/cp/xAIaqC1SGRGKZF81bA5MC2xFt2h4g+6Y+8RN5ognja237x1of
h4njb9rUIYzr139wQtIyGcN6ILgy23ENelyENReJp6CC3HDXer3sIFaLLb6ynEQal4HQbg4GazBw
ZoNGMjfhUovpB6LlSalepagQluE3qGEOwcVyzOPcLNmz0vdPSsLRAEYa4Dt1mBG6jvG1JdxEzwKf
o2k9geN5fhbzEdXUr6jXDMPa+g4VhU4CS7TY5CA7SkBPKrn4HFJjs31JEAi+9QYXpZu6QZqqsCEt
peFVCESj1ngQRgQ3QshF1cFHuHDpk6Zu2SdFbyxKFVp2Zt2B0dQKJGfxquOkVbIvrpsJaGnm4GOK
/p31vNsjNeZvI8Mq2lRAdr4BzvnprjsMANwDzeXydgj9DMIOTHhCL+8u7HfWzwOxCWhee6K5bK6y
x5LpID8qc1f6U4rzhgzwE/SpavFPVUYILjC/q+UDsLGJoeCR1l/3eJS1Ft4n/f5huGvDKWyD2jZl
fm4Ni7bfeyK8yB3AboKlrPE48EeTBGxupomw4fB9irgG9eiCLQu7nCaUTgUrkqU0d2EbFziGVEfO
UYIIFYGfeyzggEmiPlxKbiQ5vQcpsHvr5CcxGOcN2ZbKUOXjq8aZFWKnR1ErRj/1WG4OrVhCaq9D
5lxOGzkhODkRGgEz7zV8KIVFISooBUUzIKydXC8kTv2QdGkjojUMGwfY2z00dGPCLgvCg5ee4GId
nRDWU8kzmYNvJ2ExBogxB+aYYYnSE286TC+r/dS0C0WRGBgW0Mz0gGkwwwpA4R6siztqkoBC9JV8
xiza9DncAwmS8ehu9K+g6gsJ2lhd975gw07zFtbPtpoWhategZc+PWxl+xGp0CR2Ko320FnEMEgn
BkVCAS2aelhjMLZFOw5kSRKYX7VouRqLvVgP+ermhYlnB/9BJpf+I+ioGryxaONoSYDahArdmTuE
o98Tcx9UMIl7ntFfT2nmMksA694TZyN0jVS56iK1r8AOzn/rt8VO9XUOzx1L/5SXqXun27q4CuWN
RL0LKFBKDFtx88djUHwEKGKT84PVeh99plMuC6/bhfAdLpqKLFuLrKucV+Cd6VnLvHnhZyKrvLHi
rnMRxmvmcP9CCursIzb3dmTzJaxTttWH1bFSGUtdme4ic3fxwLJdvW4dtYuC9KrtT3+62r+h88B0
Hv1uJeXtKsqmATPuaMDTgXDcpT8aZn0ww6Xw12i3eS5BwbdzgWSbyn/Rr/xnqfKKHp3Hq9fjemYG
XU3hT3otq/ytZ35MD5rn6M7YHfbbQLC+7025cRmEqO0RM7jZd7LCtINZwfirN1f6sPetDoMIo1fo
VFLXyFHFr9ZjU/8BZvRx6VAKPynH12JnASqFlJWrTfbr2GtiBqoKQXT9JIPKWOd5R1lkezdybohR
j4ob8o784EyFOVhYo+iqxQZVY0k9cpsMwAsoeT0K1lJbkdsKxlZV++D1xNjTOfflKW05SsFvu6bL
te0fiBCxI6ju8zQS03OAlqDjvp6exMNDBwhVrdDeCa44/8a1AMXlTTH50P9u4GPdYf/UXfHo+VU6
qFnb++wH65UZsTZ1e1Az1u34Bjx6Nkjp6sMCMiCuYogcYIsmIDJEyUW8hAhsaATmtzJCEUgisa23
28f3ktcvnKALoBnO3PtQRFJNVFLxsvmPMz2QKXmQrEQ8uQ7KJ49AH/OMiXzSIG5tyGSkpyoyzLbi
/OTs2it/WkFwHFKP3mrAnOgrywXYCUU409mmiWWaE1SSljZnP7Ix5HCEGlcwAywRWNqsCV9o6wj/
gMfvcJ0Ycc0WwaCBo2sAMK8N+WpXTnBPzNdiwQApy1I2chy/KXW0k+R2e46vYpKrh5RV/uGrGKCY
V3RNlA6D+QekJjA19lcaFYZOPmpQzAU51X5ZxqPmTyw4yQSKD37YoQmoOyAuSo5BVJ7k6HhbbQ1T
sMQS3oxy2uWSYrFDT2bgN3Pf7q+xVvFBiuV2+qU+LbzWCLVqFri5fKG5c7b7MfmWM0LONy291XQF
OMYwV593Ro8kOQyYXI13ua14uDAOou6fz7BF+gA8++A6SjXD+rF1vSulx/e3nVh8kwqgdITB/gW9
RU/TIW4IQEQVVQOcOXcQcMP7ogVAqjF75RwZMvL2pb2h8Cs304rTuhudO6eAIV3mtFgc5JvtrDVO
8ASSchsR4oTjcIkHDjQEz7mV51AKWuPdYLa6Kw0zz/8Bf7Meje8sg+TE2lgIyykF7n4UNWVI7366
9obODZsc+lMo2GxUuWAoKbX4nQKSB28zV/IyF5LsPME5jY3oMI8AtaH2pF8YIw4YuZCXouvyHmHl
5CK+mQmEA5+kOjYl1C+bvHyj/zwDC0v7lUxVRwcV+QCfLdrw/lPHDe7n/2bsVUaKY5KjUj30ZmjH
aNDHpjHVlLXd0fmpmMaZ2/CoxTfEzm+M4f/H6n5Gw9S73XUu6nOARxIbjaz5z35ldcfTGZGYlhLH
NoRXLKmBBvyI84OMervxAUshNs0RXvnYf9GrLw/7mVqvOH8QXHlpiyqand5Aq+zLTDE1PpViUdgw
Ct7wrFNKfMmux5Kw2oCD3R2Hp7RaaBNVBVAtC/6eh1nBPmIJ548iu1UWkBKK1c5Ii6/MTb8tAaAt
nKB++P1sYPfbhSxlpMcWg5O27iuASEDvdGX1wltOr1hhGdNgitB19XJBgyQjs0hIYUafU0NElKZJ
cZYLNGbfTCjvDUqLGKDySn6EIw+2BJBAynI7ztIzTrIpyqWgoIXrFhN5zzocGspgZGY4ETw2cN8b
wIu/WZmmJSofjrYQEtUnHY9HeFlqeqpyfx4Bm/vgq1r1klqajpJ6EU5hbBAix5k0bmOzptkI5VhY
pGfCJquj7GaSwFGBEdBpdtv+L5vwGrfaDLqU6IUtSiMJKcVo+v+eb7a6SQl6JgbcnVNajFtGVB2b
WYagMkztf4gtdctkeWsnSESkxlP8cWgI+Iufdb1N5NYG875CQbQSGPqR+a3UY14jI16OQqsmFoIb
YFqUhO+4etlxUl0GfVCban2lDozyiAPTMzIdyNoO/L6VjiXieDk7LDGi4K7WkBYb1XPyTf6cONbs
xpR0UHr+VhIub1B3Z0NJe0zvQ4EuxF5XW0wvDgNlKtUnMCze0jwoC63uH3PxS+HCAEs1dmb0PKWC
6MHUGup77MYLUD8rCY0TPXNB4Mb7ZZHEO5HbdjT4fnsQzKgzxU3a+b2v+2Rri2xUO+J2fIDzZhA4
hOKIi3afKaklH630hRdahscMD+X0hiKqXzMSgtWpBpFXB/fYhM6BBciIys1Bv7qMZ07QL3ArDzQd
WhMwh1p8n4lzyJsQWopT5U9nyLWHiWduy8Jle8V/vifPojui3fWBBW6aMC1Y+YGEEHheB0t+HENs
zwI3Kg4ajsNAarp6styRY3QpI2G87AIxylQbrOOyIYWUzLM5E9cWuxpnka2OAqGhE5BaKTs3V51e
p/PBckMrnIwElHonPJJfUg3Q5ePuTtujsn4xi01h/jQRgXXGOnA8y02WOD9jhILy53/EiMsXIlkw
1MTVT6Fh2ho9B1e9RcH/u3KQBME92zYN85DJZwMiW6blMcIyWKjumefXm9Q7M1LyVVbW+WeGXXyI
SsdjN1Zqzwq3VukKprITkO/U5hKZCZppoLdU4gtWo2P6nfNw7V7veg8LjT19hhi13Qg2VeWy1R4s
WqtVm7HTjX+W8qv3i76hlYXofaCDt/s9aJJUt6THQf14fOaFyCOhb+SI2ITBsydEd5AlkPGWxXb6
4ynbNwSxoUpg6TLvI12wbU4FYm27G8eQw0IE5vs+muSQlZCoNdUy1KcF0JV5RygsTvPRwNbw1jKq
RjYKuv70AyosNcbxhm74L3rLB68G5ZX/UN7f8sDK8tVFLDsN8iaWj/DHJgVBEfH/yQ1OEAzYhFq+
F/d44vW1YgpX++BKMGWYSWMiBHuzX4oJB420H6QANNVnrLJh5YK+JC+xR2NzbOXIY8CMv/wo7xEo
yr4l38+3VlQ4RPtELzWlrk2+vnn/RhHwUBi6iPYYx6tOI6/DPYM4bvQoAA2tef/9UMmocob+bP8v
+sqsBxdIp0GMlK/LMSiOulW2wSemJEsY5PjyurJRwFozk0vZ7fh//YwHQENO2FuvOFC3EDHS9Z2o
Bkj17VNUK3fY0UJT3INB1Kpq3ulGQtiLhaDrI9A0TOOmRp7ot0ROXrD4iSfCad/NQiIfVEwcmOZH
vMQutcihuNTeEKtwW7db6wmT+tmjCRL1xv2+CHtrdPHD5IHBG8rn6xVvdB1X6lH6ULv6/t4KAGqO
qidDx2BusRPL+fm66iV1R9Y0YluKrihYLQoQFPgDh0xJelRuHN9ZKSERdHWTBGpvpRAjYJgn6Z3M
3VFQRIX3MszcjgKXn4ttyznwSCB2v7P+MDkpYRo7KINE86t7+ViBm4NnO2IzUJUk89HYvN5+7CTD
Y/6DBL3KEm6QTVqThWQmY4TGOKbn0xIRW++APYPoQsSm2DFxYi7/qu4hvgScr2nbsosMLNyP1fo0
dzorjw4KxDQZgboZH21qGVaq2CSfWgcABpZalr4V66NTNKOc7GcfP60yldYcNkJ/o9ziaYU6whIC
3FY0d7/t8MlLLspfbDzZQAB/eOLmWs2idcEGrtUcML49LtRCUAEYYSuzIEOkG+aBczT9ezaMLOAy
o9uNP0QdXSc9x1iOPgKMoMySMUvVpin6wSenqVBd/0pxPXMoVMS8fOdEkMECZQlFjgHCiaBNQkNW
xBQLcLjciih2b/raEf2oLmMgd2FDz/q5yz6T8EJNgAOhqpgLUsdEC/iZvaXT+gus8/gjG0Islbkq
Jg528jKHz54TXVlhBYkyl7L21JkIPeDoltkXhKh02dN6fWw7fDHDgbkrjt7bTLXLClipRBQXargp
68xMMuhW0q7Hf/EGOX6i1dNJrhroeyGrCsazdwxqqMuWwEDjmHtL0UUdMsoehsu8NgmThUq9UK1J
ioewnrXC+vqeXDp5lPmMGIPTSow4DCHlajMUJ8mOOrC/dnFCBufzkjBaDXBM+ralYoMmaIqdeiUq
EbJOkxfNgiPR4dAKnWMNY4vEpK2OmeHdwmUsgdpRAmh0bbJglV6PiHwjuFnnNWBNOtV/LN2ENFO5
vhuwbc8Skb5H5nrsIYi+PaFLwWhwW8oq/dsvBzbgIojpAzlwlf3DII9HPmFdg7T8Eh91W9AMV3g5
33fBDTQg5zVkkHhd8nQBov2YFUNtZLEwBtH7GHf/8sbwx2A/8zVxXAfTBtr0AZcJ2i7pC5Icpa0u
UepGfPpJJpyEMuMJLkiTmAJDEuAyGYbOMFh+UT5VMc0xdRsyhFhWiTSpIivOIFO3z9Dlzzkkq+aL
wFSDukh7+FSOlfaEqKxaUo/ojZjusaqUusaQi+7d0JZFcCSB+3aWUMnQuM+Oyf4DHH14vCFj0mEi
nOCrv3QeSjcpBNX6y9Y2XmEXS0R0AA6pCsdV69TIg07ATB/x0rr8I5vXKNWSFsxFM/JWDA1kdhnz
fMHdJJw48xuorIXkvZdu6D954z6ciqIBlepjNCXBHxL0ZP38yrq3de6jmP2PPt5Qu9iCE/EfbCC9
6GB+438nzIoVGZVSU/fKCwGuNhHVzYh9VodzBoHN4idEMCiQwiVpdkrRsm8fg7VeWrjKqZU9XeWc
yQfsZyjXn53hA7ffq5ADvX6mXm5xE0gIFiZc/YPl2m/oGufJ6CI/nE4yeiwIjbcoooJYRBoVYiBZ
2pc8bny2n9Jo+xugU5A3KiEwwh0wEgxWYZpw5jSfUq+hh1LaBOoKzHRrZAl4Y1HVQeGS46rtmlPp
K4OYUaJnUSebpLbJlapDQxWlD+WOUnySYq8tBeXCo4HhsOe42DwYhSWfRE/+2ishy+Sk/yLby/KV
E3tLwnhQr8YdmcQ4Tu3f0kak517ecGXgQJoj7yFwh0FelIr5jFK5f6QuMEc/UgWnDcTDfHUDVCr5
OQsfy524spajVKacFJ5n+s2Fp1Cd1Uxm6tP5e6lfQk4THN5s6RSvVCsMkTNBBUV7uSeUObLg6EZp
+iRLWotz7CtxQa7IgiaPIjqbLp87bjJYxkp3hel3juwByKIlK/Ai7LIa2qyE+mjvvhDJpf+XQY6l
mNn9G30P1ysFbgTO7utYEc5jepUAOT8EQkhctgAnRgv1aGkAZ+xBMwovhMzknjGRHMW6CGMqh3Vw
1+onrSE2OL2gAqjkzWCxI2js8LbOSXlc1REAKgCjA+XIt2te576kxmXyBsqvkA7e7TVvz6mwRBc2
VRlzw2APJdzQHqSaBAohFOsPTdCnz03vgsE7a4td54lnYwMyhQgKvZdHUhAyNXs1W0FRMi8tsi1R
ZQs6IuyQjr02l92efOCDBXpfLOAYPPHsUxntVfTrsSH5Sl9B7GFKVhEwAJLlh/aFj4nWZ2M4WpjF
q3uE3kmiDoZkmfKvj5gSBWNS7VlaAqby1akYDxxpApa3pA2qMNBtNDYlc0epBh3h281NUcKZIdiz
BFeSTpM6YoZwvKJQ4RHDc3nA4J/R3Uwcyzv+GzPN2fa3JGzSrzOb0wN5fJMOC0eYViKsectMnx3e
LxHs8re/YUXtaQB+7LcaoZe5Hhj91NLtPM1Q1xGWV/oSP0IwgVgOQzgn0huUNCsgic/UaUVqMZ3S
2NwX4Xn0I6K5Xd2qqpANgLEOuiLWyyqN3jvhJe8ErfhoyeT7xK6FE0SpI0aJokcGSqLFe/ZWQ05m
kZK+IjjFoIumH1nc9nJoCik6Yfk7gZyhXnO6SvTFCEQ0649qMCOrqzTDkTReriJYbKBqzKZz/oAE
RknGB8r6AVJdFtd/BDN/GMkzk1saEDYB6OnV9L4iXdoXXzcvwx6Wa/LHxbzMn2LQesnL2lG8S8EY
byWzX/e8d2TKoa4FmNLTZcsk+T2NUntT6ue5vkg8aCCBJqV14QBLZBL9GiPZ0XeeewEs0FGpWTAq
MtrLltcFVBPH6jCRIrwZq0fiVADT+Bq83j2bHSN4elVZWMhO44jbbM0xcfaJEKEIUhmygTLlCDGm
VFSEg2c8M5xkjCHyI7hNf3H9PAMclyaO1JWtQOVtrnh7IRwGt6MAhkXLcbclwL5ZWmvTeqPML+TP
kafAEKDKTyW8Tb/w5P6UewjS/o+TrYa1WfEyGvVGL+kjye5B+Y8gvqTfzksxgt3khLJ8V2MdnAbO
UZOhYr7UyW539YD6Zj65uHNs0XtEqDj806p8L175IRwby1k+aCTd1GMuwuicZrxci8NnDZz/tMXE
lGTSf7aOQ+muBV+NEWcKCzJzFbmBgR39ItGmo+OkRUGlPFP6PMfI6VswWsQrCSsIDTDVh4u8AzW6
eMqO4YZF2jpBRVAAj66nTboU8JiaKK7FLLqJUdrvpqOLMySIzzn7wcbhW2JNRPds+uOed5u9pMhV
HP2V97cO8nBPyAF9Bl9bgCdoROwg5PWxkSAXkl/laREt5TaEfiJoxXJcXi2IhO3AVguY33ZoRsf1
9FetdCuai1NIIun7JH1AnZ9pFm4BaDHisqfghSDtD0P92QpihnahWS18ZV3iOMgWym+lOaeY6DGf
ymEOiC5ZV8ambm1PuT1kJatFyHW+bR3qRgKNVK0tj23cbIA7eSEDTKC9ghMYEY97EN53M1jLc/VC
Ru1PO2NEdBJifZ88bk0BQWrtBODK80FxychlquPXEUupXG3VqqYDVBUZC5JFx13w3Kqk8uSK590V
vQR7uw8ABdegPq8LmWSBWLC52IimuQ6Aeb5YSL/walZTXojL5VomtegVZq6xHEQX7kBCwsJZJLgy
rTeMMiKGwFpe6LD7VTEHmHTu4RmCJgraf67CHoW0ppyVxJ5pK6csF2UIdn4hykyRDhr5BoKSFbJ0
y11IkPnlQ9eH7w3oNntOu0cR0NI39TZBMAjHGjEvRntFmOUEj3HSz/QFV59TWN0uGER2BegfLFI7
tvQ8DJsIkf0bE7c5vk1D3zD1lZi9thuioykcXAx+n/Zj1DLVrzkaEuEz3SQ18FFOvxG9mmT9EKJN
WnYBk2Hlvob73Kg2iK7RVcb5lyfaL+Kn3eYEmoVmw4CR57MzjCsH80eZmWeiTJbZ42q47YRkgp0F
gvTGJJ/y/6NsUNLcheINFdiMtlHawDjMMc74AXAkC577e90jC+fyRMnbrjTJyLI35NxnNpuiP9sY
pN0q2W3tMLQrHaoS3QPE37Vkox8Og8Sl2F75yty7ck1qQT8EXt7ogwQHOQVCAxpkuPs5d4I0sOJo
72+LznRRqAAfuco2B5rL+hXgVBgTfAmoMMck5fg2wG0cCzjcuiR31ZnOMUZCgmaMjZVgZqkX87Ca
C9U2a+X2pyV4IIdlB9Sqho5rdF+iRaFhCvlymK/h0sOwRi+pLPC04wbwvfJZhn6sEcA4R/Uioz1n
Pma5cd6CQ1DPqJo8MJU7W6fzjd6R6rU6jFtR3nghwfRQWdQk+cbuFE08ba2XVU9+PsN7KAo8HNaM
Ju6r6NgqDQ90lunCr8f9xYwCCbecDQ99AvJk9Q8XaG4COaG/jACiFTs9icsgEoWiiDDXWcZt7s21
9u0m8hPNHA9ZYnq7MZuHm/GGJEHt9Hm43gWf9Vusz2yaQAbnTALBcg3SErnOScrRmCTP9tfpnAw5
Bw23vPEgkiSJr6hHYMhDDPsdSFKF/DEjyj1dxC1NKNtuWDSKiV8xKZtzu+kYW4jW45U8Uz/2T/wk
U51ZuuWfRQrm4TmnsK6dTn2G67+angpMF1kXMd8sPQFJmee84oNO5zswpwnzNNui7dx8f/3Qo2k6
TY+johisDvjf3hNdyAyRsgocZHI1CEuDaIcF8yQKqiG2QWbTdFs+mYPJcGENNVHLMgJXhFi3s1eu
EgoYYFMrLtajCHOOpE3zptAETmZxCkoQnKoi2o+YbxY5GPpyQJbQw+tM8+PctOTZfFdT809BdqfG
mMjopIknL4hI+cQyaYzSWzJTjPa+q61MV807Q0ciAcX2/5kN2KnYWy1bqMwzJgZJsbB5Cu7r80Ai
Hjl5FACGiPMVvVY90hDJFgPSxWONaxnh8l+vmaxw8YZqF4t7DS2CcIRLr3fVXds+BJ6aV31vqHZp
4TdGNL+Na20gRTRzHIoOseu0b89I7QwbR1yfAPFxqt/KjTnomaI8guNI0iTyhKsw1M1w9GhZQkO0
lEc/JVZQu7Xjpm2pgdYEEeu4fAAvLUmZJheNxU/qU2wctBYUEAe0hvHmaYETHULP2VAQanzR94uS
tVG0G9aWefIBgLidc91n3B1jjqWNOvv6bxNKhGPxdv4aaGOZnqNjIBjPsu0FyHivGWDoei6/RNKP
mlRpbq9CVUAlJd1U+rtSu/smGru3qKCkLxbxthdj1oNDxqIW3WQvdc+bs5gPWCvNaFtSit49FUDj
WyzGE2UCAO7vW6pS/sd8YlpUecpgDzJZQgVk9prQt+OW/5+RqAePIzdNRBu27Ly+OAPEpHHWHZGM
rrZnz7QGZwwuDcJTH9zUpDlmuczkW1POshqfJeZzhwejbjOF6GfCP3GpNdIbJLxZaYE5O09ZeBfw
+RlgA+Aq7Lf99YCTYZboeKdkXcqFpCc3FZIj5zi6u9SWfxmKm8auB7bPFGf5Nu95p3vS7LRt8MDK
vxG7BsqnisChZ7KFoEL/cv7P5V1g0QjeIMQO7rSKmSGzBc7gvxNwwMLgK3pYRP3R3JvFeF7sIB3m
tdL0zlkc3BQ28yKKPUauYXlJQ4u4M2mQ5NFI4J3UxZC44HvWppFdW2iiMXEWaqYxxZRb0jlJsUSF
IYsMuB4LSiRgY3ZUZ4LlwBG88bukKhJ9swJ92imxYjdnrxB8nEkR/wq4MOuBUt5O6Xr08rOjEFPr
6WNaXG9ledRjXyNPB17DdlFUcOnyAUMbbsYCrQBR8SkAjaazmxu5qNxmRTKvltzo0lKxKAh00JZv
L2Ssj8rWRGcBNIFwma10kGq8Dp1XiRzc2GlBpF4JVBqJ+2JmMRGy8yw2yj/RpAMGS+AxUNaM/dl+
y2g+MRGSbIoFPy2UmboLLX9WsLXpkwu5Zsj0ZhQBcZ4jFXFKTJu2xuo3mchy08QhMpET9cdrHptO
1X5VUuKbpUqMBsQL9pzJmjrYDNaMaqMXnIIeAE6qolTsvnErmBLkV/rfDEfYuFvpbYnmcEEB2itU
wPVFJEc2m9FzO2wBTGeIu93/yQrf9UkB00S5FU+8OfMdQHBASUHKvZZeUom8y9/JlnrfJtWJu4d+
5Z9HPtZbkVJvvu+1XR0+Car9dXBzjeESsmsTEUyKHuap21S84ZHqQjL77Wyf18pH2RirX3k+Kw3u
guX7soOt4kXqnVNZIbcCztAoQkL53HqAYVKKQEP/cTfzVtaAy/6bGXjZw2UQg55+mMHD2OhJ7qFw
YD+EoZ/5qnMJAtldIx6PL75fM0Eneln0odIPLnYma7oJv30dGC4t9ghvysmc6nAhYgAKlHuDR63f
tePwxidxKGyEf0JJ4f8HdsLNZu70AYDjGwBq2KdgpYJZYQ+HryUrxHfErpyZcaECF3OoXE5TWpAj
pTzrlVi+mg3wJUsFFyrAYFwNTiJGrgvrJEF/0vePXwIu7ei3WqkpbKge0p4cHYMnT5/ot5auQBmS
V3jcrieF0F6STme+ue80vTENJoJVd0Mpu8EyP8uBdVXje253xkLhX3yNSgASBjGt4ic52BSkfJgU
3rBpXRFw7xUTSGkK6UfLfER8MTxqWpZ19AVp58oK9NzZmZ+7TsmQq/eXbUu93xPyHOlfCbIGTtP/
mQrly7CbvFZ/uwOJunbFnw4VEifcAJycsnZ9OpsljRAos12kwvfz2mHCSiSe4rUd+F7F8EqQGDL0
g04lCZxjNcSi3bY1C7Xmc64KwUGbSbvBjTWp0bBRnqRqMuUWQyQKHh1JwZ/v/MJyaWIuJA8xhkk0
5lRjTxQ1shYsNFACLbXwMzHJYe4K+wrCOyHVEi1Jpt7D9ZxzlunpRnQyeWq46gVkMB05lnCrvNx1
Xc8l/QwGrTWcS5fV6lM4Jz7VG3ZH4itO6nwhdbwtbXqA6iOxMSkTLri5fjtAcLhSDNg7mEtj5dkn
teycPW5i+pGhfH0X5UGGNx4UhibCtZAViWsAsiNbT0EelAd/juCTueGcKJTnYaxELtc2kb3wPkrv
RdsgtRHpu07HQO8oZjIjczoqbIyJey6mlvy9cB3vE/oqXq/olhu9dgvNeQplD7walPA5U4Q7eoPk
lgdyYfmJloB34TreSWiAKeEgzbyr2zyzGgCb0BY4K9JY/pW8S7w8hA9A9nrCe6wbmDKq/h7hLN/j
WOCBd6OpEjsvDmaXm1VNZNdQXZQRKEym/CFbCaHPttE9HwzEHTZ0ZeZ0y14BXcRTTNAPPIdo+pow
PcGRRkV0TluNDd/mbfATzMBV3btyArASrdB/fexRP6Hpw20/4//xdNjpERuUWg155hE9Qnnr+Blr
sx0FXbbHQzgto8VRICUzhWK0blazh7bujNvwK4qQXzNKNvShWVAPvXvvgr0OahI8+5j/BmYwlNXv
TlYc8HORhUxARmLfGb0BkPHICCb8t6hrYk/iarzBa8KAHNYc8sGOfKEuIqnMd/PiEHxjlkEKajlA
7jH+k3+B1yj0A5EwcZtAzGOTFksdIuHbNrMQEcZMl/gadjIzri27yk1bKN8/DuRXoDw6EfRPVbQH
m5ftDLpgxbi68WKFNuta8qbIGPxZsSV+q7Fjc724vT5q22NotcoWuM2J0TcxxUhSOsYkXnO7LVJ8
7Fz3KSuVFMQuEZOkXXHtvEQ0WZUPHoh8l1Fx6Roy1s1Iqx4bYOMICPBxDXYb2RjdFLqi+1FmnGRO
aDk84QyuM+4R50YfLZAVS7enlEcurJtrFeOIQJQibabFgGegGTvVOLNTWVwHDGpvE5qhxMLLpGvx
/0/c7msNHe9ePMcNlx4n85JqgMa2LBPEu4nr7ilQRv7+mu3BJPf92D0GXkgHul/4m2CNgXWSlLET
4O15UtK7Zn4H9Yii+axBXhDBGw5mw78DWuDnP17LcGKsWv55USrIyZQ1LJOPHJA7PlOmaGCNjZ4O
7urqyn9jAzhZV8x3MgK66kz6vZFLBp3huZU02ud8y4VWgqZkqiEFdSGnNbHKFbIu+eUMwztJ3OVa
ZFZX6FH8fHeNnyaAtWkw9SLxCQDsm6VHEIt+UK14+ceT4coXLBIdGk2tEoSyaajkOZmzeRLW8HtW
36NhpoA/DAH0q6b9/RTOvJYpM8x0CF8JVNR1WseSe1uKiwDVIQLOyoBUONX3dE1OgbNi++Dz+jo6
GwX/Lmydm0GlxE1OylZu3wv8jtaUqGEVprYN35Ab45+MJHpYIlXfTfX0bQ2sF7oB7vhItM2b1L9V
RGK5nyfJ64BsOnogebeoD2ouXBwIlQpVYnOp4Y6CAYJTVZY2Ti+4iBkqh/AmhnwdEs4WAFms+P53
w9i0kfmOxC/D0N+2PSUd+b86ekv12L4MVZdYLrChKR2EW4kIW3S0N5tySYn3Q8uBn2e+JwXvYshR
7p5nICznmdQFDDQAda1xmIpnv7cO+LMyi4pPHVESvpawUQzsdCUkjUhbGzrRjzWyQpr2ohHnWcQE
iipVP5t3EVsuXpr+HeLHPuDpztmhVl2Uy2ZK3f6nner4jb6ytkRUWT2ZWR42zs0652BZN3kpZreE
O/UYX+sIcdHOSBqOvWMm+7o75I8g0TTNGCifXryHqAdyUzun6AJRLqApB98MFL9l6PUn7xsAx0fM
4e1m2XszlGfjAwyi8F/k9dpZFvSnlGiRb0tQnh4hcDMK7PJnjWmWyG8ExwizOW0e9qrf7emfWotU
WvXAcagnSm7FUARRRBAQDsBdIIywlb2KvIS4PX6ccaV6RLTBx3ougPLEiNfGVMoZwD2nZ0SN/YNY
EEVBaGao6HeHLNDR4DNFtYojE4I9y9fWzepNWvE6QgXac9UtUEBLWh1w4thvvtiGleyDX2OAanDg
yzbFXlD2m1widZTparbvmOxVfx46rvO+NUXXFqRwaElEM0wkaf1HnV8FuN/045+/L1BARA5pobsV
k0c87prX+d7YfLBC1osQiZZTUst1xfKqcD+dYP6kK/c2puaMXYP161MQjYwnpRJAs0RSlKgj2h2a
eBDx1wcYCW8CiJ2z7QUPcGBpim8VlAxwrY6hz1AJMSr9gJJ5Ncw0a3IikHJH3VA/8CN3bl44A6Tr
TzXxzCtSVB/hjNQT/+46q0y++8VgsLs2JGAZkusqEY1e9ll4ki7fpIuhsai5RDO+q8mujwT1lhug
Zt8pLNPInjmRbQ2mzmP565ceLlA71s9x4OKUs1jzO0GZNGIMcTzi1CTQwqJxgQWG8Hygid/fqqFi
FYnBfATK6mIVlGwkPZpxdE1DZ0+NlO3Av478nVvXcwd3frc+mK8K31860ysOmEFivy9ITzxycFVJ
iWNeq/Axo9+tQym7Ph4HD5qrtE25CdzJe8dCsmPmtEA2GETMOlYrjRepDwJm3O3xgT6ECLsAOXhr
0peqk5k87Kg+wtasgZ6o61aULUxMbstvAq3TVVAs/Rk1Onq8NpJAhurCjgJLYC3PzNUaAMIuvPmG
DoqvWVLnPD1AXGJnyzVex0yUZN04B0FhXAZ403SgPywNSLaCpaRuuuz1DFw3k86fAyJ71G4ubkM8
6FkoybNdOkmC0A3Ush/eCH+zItQObt4vm7J2YpgBT0rpFSgytkn6799IgPao2TLYAWxfCI/AJ/GB
FOfpLXw3K1VL1SiLzcp3RoyypLTycRCBwvI6FCrfK8ye5VhlytgXXRt+c2UnmDUbakttdhrQF+cw
XXbLMj/VpzIUDZnlCvAPzPDcNtV7lFD6ylT/0Bx7UPFBDFOq6xp/frRl2cDdB8aIvJRWabMgatUg
c3Bbrp+z/x71FmS3tA9uKB8k4C72Z5MQeIu53bzaB1OvtM5wtLuOb+T1BOPk8EN6xyS1nKafsecC
0zZaGHFZmadSrsJ3jxrzTtGkArEegimDHkWAq0JgMgMpNrHH1MuQdHEB++xktwQ746huch2ZbW0q
GT/1n6HdTVW7iXV5cGEWjaM18gGbM1ZIbCcmwqTVzf096MKsEpOKQUq7FNNXyFAc1JtZY8nK+r4y
wXbHtok6uWCieU+CM434FI+fcNZaquFLnMK79FW29lmz/LWMKkEas52KgKiteErYnqvrX1G1baEA
qxXBkHRwnD6b9SUBAwyNg8vd+MnDBZJCHvvz3unHhDySbBO9TBFYd4ka1luwQuhmD9TzwurQ45E2
Rv9pRhyCtBk3KF9JFMzzcAMOXxVitOWwPVelAE+oImsb+DPJ6XepbKJudyCoyR5LRfDJ0BX5qKfF
VxDb1ven042Grv8eO7KQ69Ro4pt8+KcYumcHjJUIOQmtMhql9SF7gIFU7gQ1aKZcqvk9Mf17Q7SI
Sg8fdRcaascvbYmBCdf7WMkFywkMAL1ZHZHBXkhG8zkdSsnh6ct//6RlsTnnY8fi8y0/O1sNtX6O
iOhKghfL6OwUWje+qvxadTkNtyS6ussBgowEZ2yunLyfuQ5E58vUIJ/bCDyuguGzMe7XeTGiA1c9
lz+CUEQkEUrRvOt2I+CvulCw0b3I7TT45q8o++aT7UTCzvp9asLDxmVjBga7cAUxQcgfQbCTBjjJ
3mV6PKvp4prc8K5nIMaHDLD1mmjBHau8Ixxzbio72qHhA0KoBB5u9clJYisAqubDCq/HxJyqEbCW
Q7rpgvVCm6JHSJq45tPekbqT/x53FH9+XByx0wgLgkpDMFTcDPPkDsDHT9spN4LCuMBSnHtCsp2N
/ImQksGueHjTiFATqhnJhUjjxYND3ZdZiZopYAnmmi36WVI3mrJARuWKAV6CH7nzFkMdVNjeDIbL
u/hEo9z71g0rtA4DFdiwKR9LY4PYrN5CbRg39kvE5GkmBSLsQx0J4kXLJaRQHqu+KgfpRj5G3mrK
k26k2Vjzbn/OFfy2c+UvzB5tq3SHCUnEe27RF/yj/KDIm7pqKcSE9XDMsip9mUVXdL1ZuXfoI6Ta
Kv4LP8cDIxNczqtgB3NUk0t2VLq/P6XUAPB6XH7hWEHDRqea5cPv9kx4p4flpH9oGGMHsAeNVpi/
z3UUv8c4IY9NEwqiWNB6/v3yN4U+rpycCS3AkOV3rqo7M7hYR17HbAU4dfs/tlUuCBTQWHqC+aYy
x6TST1R0/SUKxVpZhIFK1K5i4kLdv3slMXdlC9YtrBskorwqut9BtLGF8n35N2OO3UoP99sNTGv3
Yvuwt1Jyfvj+VFhudFlvkGDJHXzzJakzu6WwGLiq5RtJJB5DPZNg9Y/pKWU3tAmwAZs0WlyFK6HK
mC6TwWYZSc3OYkyy6sjOAwX5TnW4435q9Guf4IcDyVyQ8/gVUE3SqNFebnaKQtoM7BvMRY4Gub1u
FPOrswiJT+tEVBK4KJzV/6J2Ycyk3CRIgrqqCoKtgivJ0AILXIXNeyzuPYeufBVRhHn6PPiOFvEl
WTgrSLb6RsBs6H9WueRoyHWXQKm9BjTYDTTbHnAxkQOekSJ1cVfK9IAYu4kz5Tqm5GRdI6B5gEgM
0lCUs4Bf4Xj6rXiGcvW/ydcOkxxVcjvbqvUpJ9LQzy3Kog43AYDIO4s1HQKFb/0K/XqW08Rnaa2p
VDc1LnbzIU7VUADdcAhaF3n008UBj3ZOAQijFqV4+dNhhjCqN9i6EfVLX/0mgm96ampA3mLr8028
L6FAJpAKF4wE53oeU5IROSsIlE12JknfUOinkPYnj/IFCBRMDpSdniZz2d0Zk88DKJuOaPzB9COx
k9APS0bAq6rqdwhmDjKBsKz/ikj2+mTD4FjEsyolyIEiClKVxyGzqBxOKJhFwjay+we9HhCMKwbe
xcrSAjyMKxj8U2yvc+wbBpi99T7L/xavIQwXYYRP6bIpgCoqvf5o6kOOKZkRI8IDu1yNwZu7fYw5
O4SmnaZ/Nx/uoy8Cr4jecaZBy2yKl5bDgTOWpYtLMxlDWsoYk81/eIBYbBK74VnrVPbTpUvqILO4
bHOY9RiGPiv77MhfGgfxo/15W5MhW7/1M0bXgiNNVmt0z1jzISYW6kwInU9EoI9COBnZ/2bQG0iZ
vKaFxA0z73dojCd5w3ij0TGQXDNOlT3D2vEol+GSkaEmjSj7CwBu9I0Ll/MD+lURMNgXRrv2s2eh
gKWpciVJA9YHbjLKq2DRKt47xzs4DMyJZKDmR9yIJ488hQlHOBCgEja1c7pDzoRfOPYzB83/0JfL
EQs2O5cm1sLpcOG0rpXUd4zrkunA80Wgibvh4X/lmhW7T+lks/7WLIvla2DT3AsBPMvplh1w2dhD
wuG51qAFJuTEIALVFKFNmcbjPzjBbKqZ1YWSXDmYIgiEAinBtlINfazYlrbveCQNWxo1s4wa+4v7
Cw7BGdbwT3s0iUcn6D/Oa84yi5r7BoiwbNVJ2/F6mCz89ngD+Z6t2edWmq/m14/nV9PaOLvnZel7
ceiOqsA3c7PY/PqtEIlogYthbQ0zzVvEy3Vw8B7rdKDrSfXJriFe0iOTHanxhSOldDLtVplPW46f
OwEG8JEit2Nd/SOwFNcuTtmv63IYQbendqIBklErtcqwpRIfWO/iJCCHdByDYwjB4l8ntZP8Rwyy
Wr0WquVGYGhcD/yshsEPRHkHh6ak6WWiqlImuHtElY7QE2NnfP98t0dt6e+1s+vlmVVJaGiG2hSB
c0mhQMzij5aX3DAEfrTxPouKuh/y1ydBN2Xc96sgomQ67BUaiil247QtRM93Jw4+wysVwpR4B60n
itOFEc8WNuysLOd9UvBwCq/8tgH+59TdSfzMhp/xqeEbeckSOUmTMJUYtkNezOnNKkqM7VlOaavF
nRouUwFfWBGpRvf11NLz+KQ9I7UJwnJZWH4ViD99HHRyYc3gdGLxSCUJA01GtUb6OI1qiVCYT9B2
KwNYi1bkPn004L375bPKF3fZAKO9jt72iG2ucqO1dEADvVwV+a8nvCTwv8TRBO42FX92EwIX0iND
Uje36U+il1C0v6OMA2f+mOO7vrLpvHG/IloFx00YyIhang+RY1H6tI3/p0z7nWxbOgtVs4B1xVOb
9q7npT8FpAZyzyqRGZuJmxa3/NxbPw2qrS5OpDRwxC0MMla1Q3pPAKhGa/Ft166s8hH3xU6dyJJR
Svf6BDtFS4a3kGOnOPu4JRdL5p7smKRmRBlzyPlN+SktNg/aTozNae202J8aX4OnZQETsPPhuRWh
u5mTcowoxUEyRzz3DzJpVVS7v8KOu6bZ8Xz/oWER36T5zQdBzWegRGa9E35DytovHfunFysn1QPi
wRbGVNKXhCMlkAgzqbse/73EeJChGk4vUcxSsffvWfkQOyhJb8E9UFyWfFrPr7SeU8Gdw59STZdV
gBFhk2rbntwf1eupgLMQreYcXZWoxGWUrgNfkBOI4msEJWGUQQlSWXnD1mebaTsRIYqUsx/A/snx
1BuBtVTR7gKL//LsBcDJtxh0mIsbzxbjaRROqdkI0/0WsnFYdaRdMnzz/0gGvRIP8hLXgcKea8eD
/qtRDlRliw64bGfJYEjNCHoarUlechQfli7moKWc3IQ1Qq630I+z4pFWroHznaekpy+D68kda68x
sv7cC8DXCUN0JP6EbSZuKr9JwEvCraILDQa6PcfZKu3fz1tbJmgb3kjcObzVg9iKZOhJjetHqp2F
8YfHHlZST6uxlxPoc3lAWxpjJbAH4u9ZIMLkCFO44LH01ol8c3VnjBZYVRi2TKLROLsWc/5CFoqW
NqCtsVnjerV83ItjSSyglK3Q2UltXzY4C5TYoQej66shTlWGAMcN2RDQnyok8KUMc7lOIJ9Kihbp
rgmQC1Xx9ZgGlcmHgsp/WXr/tq6Zq2MvS9YKEV1uFOJH+nuc5lR3CB76bLCcemq3tnXnIzwXeeGh
ZlHmKjr0pD6apXYrcxWUX6Wy7zfgtQ1nIaYjJS4dy+6RPqpc+YXHE0y8siJLBM6T0h2FbH/hTmVZ
Z99LgPhUe1tlimlKUc7WWo1TiEY2UEIQjmXm0LVgGCgTG7BHthnCnjDsfrSAOQzn+LlKNoc5z6fk
ORamYvXcZs85x8g85MVdffs3730rL7rNxBcLD156QE6iOPuGyPCVwjebnfLio21ndjX3/L0Ezj7P
QpyVD5J9PVwJDVGw+uohp8ULMrC4nj/g4RooigWHrfUJ3EOg3EyIRcG3aQc1w1KJTdbh4GuQV5vK
HGnZEF2ROtUpitxVz89Q+VFGu+KCm1ObVeyYSjr2ZXOqLgAGhJHJJflsVYrm/wkm0r5ZPOAOylHI
5WvZ0UeW+jpjWE0Kz4LNTontTLQbCwr2LIs1DiC82pkzoZX5AltHYk5+VvTrBGhalCo7/ISbZYSz
j3EFSB6X2QcTaBkzfs60EbOzBWMr4HW91RGLU3Yo30sgjHokto3sMSVZmniHYJeqn9BV9RAOtPcv
RXKcxUPC9FU2GwmNaYPphSpwfNSDgF+YRlVuQJ728aMXGj36OJFa6CVP0CT/o4dbjgXrtuvVuvsQ
YTIeiDKwu3BxuBS6DKnZCkADSj62dl+goNPBsRwsEhl1aPXhsM12Ecc+AOwbjE9Bg4UcZWZg3teG
/K+lTZXuOeVm6KGAuGL8sIIdUJ3rDviNb2Mc6G1zzIZLtOwceo5DEEoDCL3ua1gOPYayjzXdzcVi
lFoSj6iwu/45OvS++7JX+wXAVQf61kJ4tA1KlsmAlfrkaqMR9WxHt1hYwlfcq5frmXW+y/vJBqbI
kF8mLtjjCijTzRbpQ8Zgon0JfJWDDT5KEzG4LgMrAcD6IWj2CDNNv6zwDCpYdWlYF2joNei67Dbu
I/JGpyw/WgcbVDJbyDdR0Kxc42v5C9pYVcm1txMHOrIvnAhVr3n0gEJ6RGeF1Fk1VuZ51PC89aBv
LwSMjn4j3sFDohH7/e1pVbkoPX9l9wTCfPV96yEAbJUF3jQnrSu79Zy5Nbjqzp/PLVmfo53S5nWC
YqNeaP99QVTIMiliM0SqnyvpLsfFOUUxGKbhBPqS2NE0iv/JIw04nB3zc9YjIhlK3yVPsA6o2khr
Ts/aE/jlysqIJTh0wR1lLjGBD3vhvIKDlj2mXOnCyPgisCt54W15eFOSDKysxGPBibKzZ8h+aKWM
iM+OLUyYANSmh/SZy42mc7OjlXSH2a31iyG8+chGygHLBXEF+tajH01Qt7P01udeV44oGJJnekzb
/Aj/jPU1pUdeKQm8pXvBx7cumKErYQptYkcVeh3tNWUl+j89dsPcrNKcayfWKNzq4+M2S02niCV5
YpuZLpHRhGlryrL8W44RsCNc+ZY4y2V8zgbjBnwObHWDtUzGwADzBtULOlB6tz8tii+KsEblvTIp
Y2GroKTd36w3Yw2e4OK4oc7/YEpUsoj1x1aFPzCWFOvNhSoTt5ZC21LIVkJ6KoJCl2vn2+r6NC81
RkuyUd/DSbGA5KYknVNoWqkHaYcAaIQUznHfa4CJxTsXNtAmkrWoFhYHGyX5EQJ5NsNxOE+vAjzU
YUw40AiNRTNy9qlvtb6BvO4o/wFaJcwcPs53ADTjii9Hz1h5Tm0MVRKQ+iXcn62eF9ugsqvfHT2/
3UGS9pQHvQ83H2PiKETOTKKFmbW3xvih5mDiciHbXkQWdtI/3YrqkoMibldukEmaUXNdulmBt0R9
jXRf1RicXATbIypgBXfQBvolUK1j1ljS2XYglkd4/eCyh+Ol39cam1N3sQPI6uey5gBaZ5crrNzv
3N2TwmjA8wOaw/kTJdBRrH/GwxWpB9nQe7DhSSWnAm6vk7u+TvyfVcnwGCibPLlXSgBYwrJCb7HH
yifsUv+mfssMbrfgOjDvx9px1ya0mVrZYxIiASsl7aIAlrzkWIP7jImuc8neMesmCAQma53UXf7R
oK1EpfiSLkKajrj0sGIcEWnVHh7W7umHak+HRFJKpPKzf3ftfrwZ7bOY7Jp1X0YY/av8z6UjGXEG
S9q8hw0CriNnMMpsgSI5zCY+BhpD8JLhWYE5cvOOJHXPS4CNZ/VJFGk4fRfUVC4g8B0p79BvwM5c
od+0fETnYlvlpultEXS5WGdFo0Y0kziG71r1JhPKRLHrw2vzpFCFpaMts/pefVbOsNB0bVo7gLDX
5XNkjbwYn0tLtzC6+/Tbnc8vNSLE+G7s5USk/lg1c56DlPLgjTjftu9p4okwyBc0tmop10D4rbNj
kdCyN2nHS3xlzdoqi7eitaZ7SK+Ekg8LoBAqeC9f7rII6BhxH2Stlvv3s0cvdVdCFdo37Yy0ZMun
UE4Y5wHowt/kFS52zhfhUuvN5VBmpiPY/+tYCbJSSQt2VBVcLQubcB0vKZKJRqq3dFZxR8ht2RMW
ZA8hXjjTYgulCLylf8WYE7B6Z2tT/jYWB4D4MD9TUB/hzLywXGBpSjfAm6eXgsgsBhkcIOEkK715
2osiF/ZrimXshMEap0GQ3nCHhnSXY45Xczp+jQS7tkSl3HYt7sZjIp1LXRlZCmiF/YJG3OikSE0h
ztOS1QVimWI5Wi5BT3TRImR6X1r8Z1JVPMGwZwNoG6c2N3tk6+mCqA/15SV9bgfwdQCWQmYA4CUU
gO3KWnIitZzhAEn8reZ0Mo+Ml5bphFcV4vSrXGiARM+jhnJXDLHKwBz9lpU4tC2SOVQx5gIlX8zR
cal9xdYKTLTOAnuaj8nWlclnSzk/GrOMsjt+ouEKBthGmX17PMAVvxfvEGJsc+WTS8GmJUEhhfUU
y4zGlczKCZP1Jdnz5cBwITsX2pN+V9Habn9qIrz/PSEFmmAuq1hLJZXPO/qLOvMbxnCmweEbXcVZ
yHHQL8ipSe7FyRBOEvYGrsdBg/x17IOCztOtF0CUXUMhGGAgQFw+6zYb8cGldyzPTDUdC/JR4bVZ
SXy7b/VBGVP5fwRJNi9MPLRzWuvHFRRqJ5whP4NgK47VlK2Y0Iu7FyZLjGuClXZ/Z1c3Rc1V2VOs
jjxyWgDXC3DLaJiSroBguqSY2Y8RdkLP2EnYKDIDmXk3LcpbJKuv5OSSxXWxroe6QGVkPTo7QmQH
uqNPDxw1g6EqfSwYr3FaJfrH73M4pRCUMuxHgAwrLydHluNFBwOAH33c/60Vre6YsO8xsWTuUmuH
uljX1God1JA/wcZYHZYsPiJ4unMVdSMyKwCgam/eMJ0bQ5SCaKanUzz2RoewO4jMqADXwk1X59ha
rTYpiGupG/MGXKxFAwfzmMow4/eYk03M4eEQC3Qs/SljoDn4/Q949bqPNdsDHBTpEIeFqPtCmXMl
9kfyEQyUnSUjel6CmbIMI337SDJkL9pQkaw8D1Vh5Q8+2qsbtfA10aFiizmyPI288wpWDDJbffpi
C78OIfoz5J+frIUpYz2SveWKeHwUccB9up5faWDLJ/P3BVTEiUh0rzWS1OX6zqmF6lBjDUZAns57
wRUGjuzz6khtq+5yOeGW14cP/XEPQ6CQuAY7w4QWTdj1/xxd2D+xqnAhrqIq+e4LJSxR2hprlmoV
SSmlqN462GBqb6u8XkAM38NPqg0kJgy7Prjwc3rMwMakZTTvZ0+OUbI+lIFhkKd0+MYLwugLwAc1
5LRAWVA13FkCUL3HDRO3djx5YrKMehPiI+/AwXsJwxn4DyCgp0hRhfijBDeQjHzWZ/U6Fx3gZzQ8
6YDIaqc2cwyco6/rTK/IKMyp46mbR2pbrbCkXRycZyOLFOkYGGfWDUpxh85xEIvPjM5uOFhDopgi
qBb2t3C0O4MpVZdR9d6io33BqpwBbnj7yvrXV/VmhGx5rrRpH8PtPz0aPTQ2+xWwcwm+Y9zEIbX0
cQijckfif7Eg4hj3fCgPxQ2Khx6gAxVHuur+Fogwfmx8O6aQh8npWEyk2uorVYK2HbfJeRI07yGm
U7jcick4X9IrehxkaQn58O2ry2q888rc83Ms2Hct4y6wu2qXQbxp/7niWSm86lmdXXHGOhw1gM+n
QoWVeV23yv7RCN787oHBIAra+9Ji3tMrXfb4jU57BJjrxZ4eXfnq7Qh6jDcur+8UyzWOAkgWdyEW
Xb235u9FTj8Xe/cFU6aXqjBYqW/kSDwDF2JY+j0ND4+d0GzsXFMoOw4+EU1u4vGqybX7WMltS/77
uYDWO/DlswForZoJo3tGVRDSc6Ua42PYhAdp7YGv102nK88QyAa5pCvqJ0ZLyX1zGg0huGwNnzDD
HIli6swhrzlBY+evw+B8fUMMmaGlK3BBiNIx2T7+MpERJ/vaImPgq47N9ea6tricg887PjN29WGl
NbUGmXQrWqYJIBVaQ4iKruxr6HK1KGrChi+QQJ367r/A55g0J1qz5bFuaK1ge63NjG+iY6Yfdp+9
wSmmnpmcAcrKGqBZiPZCO6+r6bzzxmZa0d6ymqPRYH5rnoMI/F+KLI0u/kPlaWhMFafD5vYeucCg
h9+SbfSaY+NpCDX+nfBPQuSY2rQyjH8M7gcc7IVAGKAGxFfoZR4M5bSHnOV+TsRWfQ9ByF/xrglA
0maULC0czOMQcznHtg1B9uWNS7iiT3GTw4nClmOpLGDDdaejL/+Hq/8JZ4lwButSkRDPI0Uy002T
mdGUzhmoz/5lUt0Ry7X/ZyeUaUOjJbMvP4ucX2a+UxgFyCOkv7rUZARbn2uj8oO7DG9zGbUm1dzJ
BYI9MObRY6UlH+oixqQ+XF0d1eAMKWAeG2HtkBk+fJE/CO1H0q0vTRkVGk1kRit1rz9fHagEtELp
aWVHo8/ZCcloYtcIM9eQqlXJxPm0huKSJ61Ed9e6rJi9D9EQhYcjGCEXh1slat6XoggdiVDA+ZC+
bmjU/DKS2pSecsRHg9Dnm6xaE46+RoNreqkKzJ0+IpryzF4ViafjvJR1xu7ScRro0O/WaWq7qN7P
4k4yyor7l6Xbp4c+KRGz/4kWJH6WBee0hmjrf9pZ67VfX0B6s8eoluHJAzSxf+1/z1bHA6L8ufLF
PI3om79eOS7115bpiGwa3/h6f0yOs54GgruND5lRsiBvoiCKN/JOktk4pmZr9UcsF+XGs71/DNG/
YhAJyxtvM6CB6iHDyBSss5EaDWwraL+pyeZwJFgVL9qPDmv6REe9CPxvc33hOGipG1K+6X0xNMwP
uxu088C910zrfuwnfAxckElid3uctnBKxGk0p5jUvX8vyFm9V73v59R2nePwx/EGTGDbeV8Zgirb
jy3/B2v3/BJrfxhrCvOTOoJP2hNoQ1OJiwacbHTApJJoYBwjicfUZftYc91Z3vqsQUYzNlKy3fii
a0IeRWKLntGBsOhaPYAX0Re0WKPzgEA69PxGcArZt1+MKRzWPHuG8SB6ffplW+17W66zYKWTqecj
2zXAzFk/vYaFYSPZAo+RUJgGFgwx1Ndj+g3YFpwgw4dhkqsxHBms3jintmPtzkb4hzkd7yUqiRPu
mAlXuGTZR5IwMFbvXzORE433a0ExVLqTgNg4BqNTVZcn0nDXbCMvQLISFhwsik/tVGHXh6L0dCX1
eFtazcc6WtIFMkNmpwLjT2AvA8nABrx0/BeLsLQ8IhUHgzYyiLDlTFtvfp1PmfQj0Hk80JD9Gqqb
VTSSxNXczVLVUkl291u/Xo27ygnqXF6A0lmicI/KztYcWYxunDQY/P9H96k89oRrXfwzoCzhlK9O
0jJPzixCkCOJmvAeRCLKPWDIp4lUbcWbsX+zGbvU3cderjERiatufvFaVSe+wT/WgxWzCCJWFvra
CYnSvf1gSRTqUo2J3FUIRv+b5IP/sMP2l4av80J/qHyV0VaqEi/0IU6nmOzpc+oR8i/FliP3LNNu
vHjMkGquciF9gfqUi70/a7smVTWyt9qkx6tfMJXb/bInusc5jOdL4Uq4ZyIhrtyemf6jYU6iiQY6
nlGioeBAwWcqtTrz27lt+8+cl392s7kDiTllDMfEG1+85ByYiALBwHRAXkxHvzUk9cn4BpP5hrCx
2r9tFEf0mMkb0Q5Gl6mOy/C/8MmLZWKZQfBl+aUQjUYvpYXaQV8qiCSQuVb9s69bW7QhUjMAyqwX
PHHymIIE38aKK7TPZKkscUNNcyf1Qr+kEkWafxQQlb3key6skd1DaF//rrDPrW8nWGL7UsPCqvo2
pfRNwPP49+GFvRwk6vnPlWMwTCpRn+Ta+61w1CYLAx9k4ApYRT+8W0UpBazjPmfhHfLaZjGuJs7v
F4R6z4KozlF7W4eIoAWZ1PfVQZHbXT7f6/7PaOFpqBydA9LrMKqA23gpRdUX8qVWScEgpAcLSvS7
LcEscSisQsXQmoNI9EcnLsbjRfcyA7vziEQ/9OgD/amIn6FWbsSlGTIuzBYOxvodiI5hdtq5chzc
iARFTyIb+wPh+bTf1aQt4yO9tsWEZBlCmDa3jximNrrfTmV5pQhDMiHpQCBYOoezLxgm74xMGN0X
Xro5rl4D3LDUsD6kCwwQbzsubSbfhZzQ+c2mbK8ZBCg9hz8dR6L8qIdOErMCt2vEI6gj4fhdca4w
dsQAvws8x1HXUbD2brKu4JlZIWGCZuwdGRBIY3Lp8g31INPCJdbP//j3DznqVy7oDiszVN8VKLrG
o0wCf/zJtnxWfSU5rdhwZq8qfB8D3GNAh163nBOoYs2bdLAP/4uG6lMoOjjbTO1rsxbDGT9oD71g
49d2BWvFfNvQQyySKUbkgYYzNuby8kqAQzouVBZUggLhhgFxLE0sPh0nNmpu5Gj6XcEjNZvMDdwC
L8YxE2/G6VEgrOQVFvqfeaOVpDbrDkDP9+IKXcPqyG+EsJJHwlyy8OJYuo6MPkkTSOqkYZSM41v0
5AGvOCd2zx+tMf0jUmEaYVQtlZxiYFUO1JJM6kWT/S8FIVfDsLATb/RwEivx6aper3L4SWVboF2c
HTKJRzRFjZmsLfTmwAUniRbs+g4mmxSOCB2Rh3/VXjirMj+ypq/gTTOEzGzapJTm4ApHCNJAyBS5
K7yWVz0pU2JdnCWwG3tzGDYfLTbPlToXQzmFKnenbWHFOfhA4wRbe38U81nYwDTTlyzTHnu15e4N
AfqnLEarrH4mKUvMG08lJwZHuKKqYjAPcSBM1QYEfHmWG1gg3a7k9RJHEgOtdEHDxhWanrBcdKRQ
Nw7tEDWVLv7eP6EKDkqc4S4avBZojp0eqfDzLRTzmduSDH9ceqBMgKjNEtk9AG0GV4O+Q6XOw4Yg
kjQUChfqbJvioTF9BVml4IGdC4WFxUFtBstcjjToTGqARnNH4gfTgQLJ4ZDbxpWd6eoTLCGd8Fjj
Bt+S1jPNizIaOixGwwHRSAHT3BnLuUJTmkxm3KVhxkLFIWo9uZFhiNKJjz0Eo+LOst4e9DOxy8WT
iFg7L2kUr6ofiTVc6fJtQ+Dwgqh1GkiHT+d8HKJh+0BjR6g6c16BSyKQo5JdQ+tm3l3Fst5WhCE7
ociZ5j6mg8Ju1/PfNhKUeZSDHinNxudKgR+w4H4TPDPWCvu19YYFe1x7tZKGXj/gEdSTZuQsUstC
WsqY/Rk3cfLLIdQjyZ6AkWDxJ7NHBsvucsY9BxWoZ4zs/lhMawF1lRCdBeDedKXp7txrfpILlf/b
PQKsHHyGv13r+uzGl7LXMBnlSB00pGwC9hjK/9AqscEJfczR5WsMTniMpJ0ejfipBeAUpgaMDst0
CY7ygOROHbql7qK9w/yJIotTDTL0NfY0biOZ5i2OaJeq8d67wXj+rPDAHD2fWg5p5+1jWUrVVb2n
T+Jv7ViN4xEnM2TLKeFs5Pt+QJ8cyOBAjWq0Hl9fwHGOe+tII2bK0WWl2N0IhC70z8TCFsxhTrNg
wYeV5n4ZA7urPCdnv1kbnjR2rxsotgLqlHLkY69haQJu643JbEfgyQbnIKDN+b/fpjPMzTVSqxJB
6l2Fd+LElvh/xKb2t84vjKyMg8ycvRt+6ktqWHgWliq8D938noITbaQYWQIIGEcm1FrD+PZC6QnV
N57+Mb6PJgWe2MorrUdEl+zzU46jFOKtBiXSeZ+HyJS7K2GGqY37XaoWIAOPW0R0rRM72np7+0SM
yMYuv445b+ct9zDMQrBYXnj2nflW8fThBoZYYUUpjhHc+0Aze6RR0s4fAGUQoAc507HBM7dXormv
ggtI7klUb9+UsFek8SVyqBCIfknbxwt0BBScIsPQ9CVKKtnSsXs3pkCi4afzL4HKFYpBL1geL+Fr
thma+CBB+AcUIaWvBgW493nd9nv3g/dRN1vkvrNOG/BSE4jY1LomopaYUJ/EKig9kegCJ6sPSNmY
82qOfhm7o4xjaExdPVnRUeNaOYR2YN/nz0OSP5AifvRxa/9/gyjhXGfGbnUyiNUyLyuuudWv9Aec
FcJfMsogXq3BUVxcn/BE9IMFE/VbHiHdaiuqoadnPd4UZi0Lslq3/4FTpMRjsDM2/vDEgmI8pcPC
G6CSShUaBfj2g8fOyilaUN5NowjzBmtxcYeXnZ5oq/eGyGq8F0DBSjtgvHypZjqsIGcJKHBplctI
uDjNo0QmAzfIlWGJuMHejum5j9D/Rarmkms+NSMjwW8wjOhuWTWszExaUujlN5lJBEytUA4AZspS
Xmy9D0WL9jVk0ZeVO6lj7XVO87vN5FE6vpB5jWBdP/AoQtL2zT+QjPFM1halYHoAo0RuLVHxMs7Q
u61mgl14R4C+HbrrlY85uo+cX9RJAdx1/Jn3YsYlSaOINj9MsqfQ1N2xTTrgJtSgarKDzbesDWl4
dc/Ro8uI9U/mYiFSsm11WfQq9g7a0Nm3+krfJy0xYv5WxqXjrXUlroWcaCAf3elaQhlTH2xVHQl3
qva3PyFthYmbu5HWmIjLY5p7NR32nMLztOO1vGu5WhEonPLrQj9eZ+TooYHqWSHrBwjaYtH6VY2l
KnXG4U3LP9aJvldXABKnm1K3Zm+MdRaV4OXN3msVKDAjjH6CRJ6dEPjbHfzjP0uabRfdqzH4HYUX
GUGJ2fub6wkpPuJWQoxrMVLZ94NqI44yUrEabLWRHGBKp3PDB/xubniorCLAYM6vI523/KPpNDJa
RIbllItOQRZ5AplL47CeNWR/R5aaxFFmbiP8zFk9DW5a8TLig9Hd74a9Qx//qM3THNkze0ulwnQE
fH8Ml4yYfsSMGKlBC/kiUtQa0l/fZC8t+dta/pivvacI2eyJe+/VicudCnWibq5WSmKfMv3TnwZt
oNYIirKQIpH/k1QXgGEBqCi6MpB8tIB8g60Znaec/3WkMOCXgSBUpP4Wz3rKv1Qg0+ipAtWRFTGH
EAVwZqMeQYaHoDwWd2Moj0BvLx/bDyqiw3ZEE9WzOzAcLQ8rjO7L9ae724cy2e4mjYtmx5FS/bw2
1n49iyzeqqEFGEYrDkawrXOPHCkgYgQzOa8qkfLCY64JSqrUC/m50BknIeuWx9H5iwpWZcIUwRGP
kukvs8YVpKeuuBaJznf5MGDxvQZ3Glz0nc7SK4MDfvyXYH+ZsSW1QKhZJIOK6AO0H6b5MdkbDXq4
+uXO0/xLrMAM1QvlJYZkUNB/lEtTZwXVqkVEY4q1SpUERynzA69YfUYVPymqyN0KyyxfwmHrf0CT
7nA8swaGuOJU3ONi6SDpmbS8a7Z6ooMN2LfcmUw/mvNQUQXmbn7JfnJ0nQhFCfqvkmH+U1vEPdGV
a99JpY7HUYkuhOdsJ6+oV91uqpU1ah1UMvUxtvlhHuop9jgDaveQcZCWtwkqw/43Qdd9dzh6J65/
/lDPepLo7+CDK5zwAZiJ/S1X8fPp/YlUKUu7F2Z56qg+l2+y4u/Vyh2dGLX3YLbxba1sh2HlpkEc
hCHh4AYEMifx3PXzRMxXaclLgXDXs3AZFfotXPZOXaI/woRiwsluHlM7ZvZI6DNdHtq2aDMYbfGt
6lSpMJmT0OIrCu3TmpLYcBJ3mJaiLhjRcaAXQGljg9uqlxLk2rIY1+vyejAqd/IHDPQCHpOVdTnJ
aSE3prpTeSbXqNHww2Z+8VfWcu/SYVWT00Tdtl5HM5McIpOMo3LMLhR+3eVa7R2N971KrUaQLR/R
KIlKG83ARqE4JGfsUjsDM1qh3f7VnyQOa7Q7dm9V8DvNi+Yg6vb44CPwdyzxRuzEJ/5B9Pq/3lqk
PYGEKNUJARmvdQ6f6BzoAXQ7K+esfc2e9dqgjosdpuHHAEfpsPp2jp72fB16/Qzq+PRWiX1ehxz2
UqXscmchiHplUoRShDiHwCKx2mvtJDjEiyLvvS+1AXyRSu4EI0zP2akJRwkDUphWwvmQRLh/FNbi
/wWcj87RK0m3TBW7AM29jP6sd3LXof3L7sj2Yyxzk2inFs6iDqXyRIMAOnaiNAuv9ae+Z+5yJN39
VA1HWZxZkPDegTeVB86kXAkDWi0Lv0DKT4oTWfA7W4ETs6dCer/swE07XA06vUVH4cbcKRECjciJ
NFSDpZ8ZjrkEedEyv1J1Nv0PZlOLceWm3lckpPVpR+Ma6yED3EP3dX/ZC2MoaFVao+/rOIXrx/fW
tZHC0IQuqKscdwRvymGcVK9bzBbsODignC4dOvjc7xAD1iSr+gQS5etzbP1En4QgSklsaJ4Tt3QE
eyIGlp08q8bk9sr6/8bEf4+TWCyfNHYsTC9utrorFZ4Px3Hf+raZUkbLyHs1RZ2fIVTxyF3xr+TK
qto6IT2iK05XUAJWZaOYwy6Br8IT6C5GDWjHTdhaX5PmHQYVD9ic5FRivJ2VWNWINAs3sLifABSp
O6fZecigXeR7k2rmjoFcCBQXwtfHUHrZnaqlHqT7mr7quhO/N4wp+gT0zY1G8rZythusvNZhu019
3OaKnEw6p4hWaLgpFT2cRDpTfpUU1CIKy7GT9eiRZ0tf+3YyWxjh+MUa0HTMiyu7eBxhmfl2BRb+
3GWWFtv0umAIfKPQ9/XoFHfHEfXqEM4tD1zWVkNntRgTxXbgU3x/izEhGWOJpuAnxC3zt109HFI7
yLCKBXTSuwZXMs2mVZ8hmPfDMkVS0D8+/RwND2JFc7nqJEBqlEVpRtSf9Qi4KjjH8zitNtF3ET3+
CVS8NYblKw5hQ0RQ+JQ9g4pJmQt9Pf0fXGqSgsf06IO5qzX56Ja1QKq0ysnO1EfauaNjfsoFQD+l
okK9gUPz+jnmcn14T3znioaYZT5ZVchqrwt2Vw4zslaxkl8PA/aZRS7CgXkVd9YZZ3FotocJfxFm
Yp00SpZUiycg3Yw2D0pEpNloMVCXDzNP4SMPws8jM7UIB79zFxRob8Nwf1G4SxZmQKZt8zAIEBNr
khWYkMdgef1uqeR+7t4lXubAidoS/uNmX4MMUKyes3OwxF/gd4mFDydn2RbtDdR0xZgcQldnaJS+
tGcJP6L1fPkMJFagFPngQJ5ufR8ZJ3OF2CRET8PR2t7yMjyX4T/sfRRHU7XRfJawCQlMh/12BJAp
TvVyK/KztdgIc2XIMPv4vy0y+QUyIUysp15HHMa5Uun4421mZzNpkoax6mT3RA/vmdj9J132KNYp
twY13dMhW0FPBHj6PxUCKZTVIuodxEeYdvqT+6AoiCgH3mV2kBWBJ7eMrHFuBI8ScCvKD05zhR/m
EyhWV1ISsqL/JicdZkbKPOlpZxEZcEJ3/143zOiJ1HBzBn+F/N7WYAl1JvOAblqYR+tcnvyVbKey
mI5AiZuoc5S75R5JCErTQXLbXl/sXOzYhc93HnKnMW9WDDrF8xx1qLPMsziMUlHzINfnk0maVdeU
O0bU7TrkrB+LakYb7caR+XRuUJSvZQOKwKCQJifv3MlIOjgkjYfluz+eRWeQyE8kkmngY9w6mhnq
U8N/fG5pa3OScROfuOtXMkGo8EHYPn8l6pMoOruEBuBpXvw4+MevhDmFDh2f7BJYv8cCtyqLXgN+
eidbq1yuN1ccr0HbZwa5FjrI5g0BV5MnIBaoxYnok3cKWkS9Y+4RjKmgePDaOtXfhH1ps6ANEdj4
k8ZBtw/Dom61BJghuYhNYoL6aQCdR+39u1GT7U0vDuw6OUgbspbsHupo92MDhs6k+w+jn8DoutVk
CFq0GPod2pONT7fx18/uRn1rhm2NKmgJdLGOPAKL+UglTzzJYqosjp01zwwLDtNuCEMJGCY52qgT
1aT91dtV5zFycxBIY6P+c4h3zDcmidXs/EHEhcPp0zfrvsqpFMSNlTeXoq4r0jdcdZ34klUrj0Gx
Mt6i2R2gxu5pUV+u1oHvCM0EqWmByLfMUeXIO5/s4noPpipSbFAgQNtiMW9ireD+qOqBYlybUtDE
GRe1NRaXt7sL/QqflEvhdHBxMJqkd46re4CeXK5eE50jXKv5OOPTQpo0aitAdmL/EJEX/UJlj+q8
l/a5FTG9Uxr1t07Gajfy0m9fZZ7pQz0j3Jmh9iET8K3Hr54GVJ3/9B/7Vm6bimBlREuMzshuS8ha
Rk+qZwERDY1FX+NB/rKqY1FsVsq0KxhWXWLLaKG1Zi5gFMUH8XvjXGH69ptBbPym0F3E9QqsrkLK
5VXsyQx/vldKK0rLy8MfJ/OrNggeA3gWhPEl2OYkMbws1gWmZYJGyrlDlaFM74ANLWlsUzj+tl1a
NiRuCqj0FBOVwTeMZK2LQM4HeQ6QRE5vQqIO5j69MhQNxXF638sKmXO9bbNTosdq6n3MbPVlvRsF
BepOIl5Wgr6i05fzDA+WuNDsdcJ2tIqCyb4WHlnD7l6LuYsfNfFhQeRAWdBMwMx7nNqEYhlxAG9D
R9ByPdgpg1HIR7iymJtFa8TZMi/eB+wHsJt1i1UnQL9LFIdZ4B6NQRTp21iCtytZQdopv8xn0xGn
6OEPRYClloqNOwsmvmbrR0wl/0OXFroA8gcDczXc3lkzl2zuis2eOG6fzhXBPCxxlWGkBH32UX6F
NqZXFXcXRDZGs9XIOcWd31gXO8xWDIpLLLzt1wksWwF1g4jV7OjSqJHu4q564GQf/H99ICMobKiy
hYSDpU9vscBUIIb5YV3rpw3BKU9e5LEgXsppiQM546Jdquo6wlCBsyuVimo/ip7pdtJwjPJ5YiU5
merIbadM3FszxLcj656rmROkHKHTeUn8u3UaCqtIzSKzXJaRzpRhCVvfHFIcTWgrJMr5THu7hI/3
xIJ8TVKtqJtJ+yFXhtxIu815fIZdi9tycoBL6iRrcTnbEZee50dochyNHb7mDJvbw5+c0AOv7S6N
6HtRv10t3hflJNf0EXtVd+OJZ8RpyfL+V7VKaPLFgVH9K4Kyw+jrx40HClXZa66jYQHggqUetKVm
bQpL3NHFdO6RLz6dk1sTYOpfcA90AEYSAz7J/zdhrohe9HVuj2WWcDuOhfrd7yeIlK/DTJY4ChPX
/3K+2jb45uTnONQF2G3GjZsSK05BW8ksPH/mSHLub+W1rFELVMerLJVMM7K3W+PrNcx5Qo0EHIcc
//Exo8kzabJruMR9ldg4LVjMtMNoGARSGQjm/64XsUZrqZk33uipM2WbosXQJFnfg0OfeGs+9ixt
8l+Nc2zdo1bAGxvm+mXAGJ02YT4ElNmo/7nE2AQdM032MJIX6LOYduDLxFhswfwlku54clSA3lLm
GA6wVyCpidoXhmqzF5PGRrWjNsXw0GVrwS/DzGv02JuWIOw84Ypge1jmlsYDSc8TyKKfn1X2lYZQ
W4d0ETfzAshgqLvOUNrAt0SN0eORztOTHUU4D8HP7xN+tKlPKpW38aV7ceDWHO+SqPvue9HrkgTk
nnccKDkdAy7F71MtqDeqFC3IbtMYMtb7XzOTRgMjNVXryd4jfFpWEI5e0DT5i4YpgAWmrH9mv7K9
UH90o50FJy/RGtqfe060bVOzojs+lChZQgP3WwiHoQD2/Fv8DwwcCuY18GFybi1zXO/DH4dGpF1C
xw75Rs8rcdLHX1LMQRZGl3CGxCVu+yrt8A4F+yCwbchfrGxzx7NNSXesDglrHu/vhdfaUYN2pVYP
6UJqnyBNcNWt/Rhqu/gxIP4XcpQtCoc+mHE0sm8DsvN4428G1KLNFcXLsR1l0Hm4CLwwpvi6QTnK
KigLaEPGtEKwq25k2K6rdv3NRORiEvo/Ja75OPZo81qZ1Qvnu6yctL8n8M3uveo2Fcxfh17VlJPK
/1tLYJFlZBeM31IN0PdnLwXdXldOvzQP77N1GFDgGyydS4mHG8zJ3EO92DIITK4XE1qzRdmi+kxj
xiOOFQ6WVmlsYFtdqa9ljFWK3WxWdFbnrXsTsQdETvXajl+nSGUxPm6B+ZN946BqpSZJfmA6JaMD
5e9CjXz+w4im6nIpgwXg5j8g8GKWtLN/vUfJBak3zsfKdDOeu9K7mPN/96EFFFjrrD6GiqtCYW+x
4rSnCCePw4vXApwQRTWAlC+3I620/j/Y3wn2YqWlAwrU+9GEHOm0UTHnCC2PKBMyYvGrBmFA+swC
taXwaSPylPiQLEVeJ5sJQ7q0XFrx+HJ9AERZZNuTWInL7jPPFZZf7FrU5ZID7ukv4YyHYWbyMVyh
usnpJXDbSJFDDb4AooEEblcC1f/0EVOVExhpDEPZ8TmoJ2ZEUxMfU6rkEUmvkrDgQpGmxaYqNMIp
TBGyf2ssjMvSm6gbGXm7fqJWHQRI8q+5UJc13X78VkP0YSAedDTeSV3zY6hMylHr4iWBdMp/PQ36
XZ5kGKnYrEH4XTdTZsONSkmNSGpX9mDw0qvNNCRJJ5mao37e00bTguOPfoPlL/grvXQ7EMIZQU2b
gw5MY0UVKQP/jV5Hv6nv41h6moIvpExmvN4tfgCheLMa9Fu80r4Algi+f5B8J6f1MDf0kWTgDokv
dCc1WFDZ0KUkiiaLLAoLkihFIWAXwGnoISu/ISjYj3l/28lSIMB34WEXVdVvJJkK5rm6WK5tkpbV
LU7ZkbI9smyxQpbZZPwOo/z9Jn+iM48bGMkpWaz02YAO487gQqkHS0SGNeHMAtSG2BlG+iwG60Uj
6dbCvEdSfMXYQ0M9yGpy6gXEQfNJq56w5DWW2Leof4IGOgf4smG6feljRr5oEEWcM5YLm6reVVLI
AlqvbNruUINPZ25eCLxxLwyD6BKw0w+tLmu2KSa8kbcHwXB0y4KLIr1lrznvpBtNTEhCxTTec6bx
McLfJJ3Jo1Tj2MxHIZychYb+OebUauhK2MOhsn073uqLW8hm5c0YWO4yZq4w3IW3m5jMRDbCD4sV
m8Qu++jXphMMtGWlqRcT/rg7nMKrq+YslQXy63/xg3VaZkcFQdJJbf8M4770g435T/paJvIrLThr
4oo3BvQx9Zd8J2E8s393GTpt58LOB2l65D1OhKhS6d3t+yvabFeOwv71JtrtNOnPdSs/hk/kAkHx
zsk84k0fidHZobi5kR8D8jEVeCFT7lwj4LEOcDPM+sherJNew6voM1cVdyWrcXZXoTaFXMlIYtbq
YbDFldozyXuG6CVjHTmnxmStsw/l3Hl0K95CBoFkGWK1hZ80YslapcJmPiw8Y5CtnPC9mx9T+gMq
RjrZHRTyQJoZEb+ewbLsb3a/6QoijFjtF2D3ZCCKkglUQsFClreBh/f+j8OT3UR0nmzIsXn4BBaE
QdR2PRZ4rbRFiJWJ6lgHqeDZaSX1xwT4yc4zGFInwH57rS37tgJ4twpOWQX/Ijw06fFn/6NEHzvE
aLIpcdmLT35Trln3HZZ+ubQ4uxdOH44jLvplJtKdgNUUOK3lyzrehJ1IUDRvquIkrI5clQs8SDtw
5LQNZniNHY8eXjIx0j9VA7lIUiJ6rle+SQhJ975+49TNRbqBSHAoZQkWR8gph/4vZLXEvQpxIVNq
Tln6pasamwJpRkFowmqjTZ9IVg9atiSQamhWgNeJqSA7nTAX6owcbdvzLrfv0HvG1e8ACQ0T0Y6z
oipUMfnot68aV4kdcPZgdD74eT3qvH1AfnJw1KXiAPwgp3qpsmjJe0A1mK1/T4c6rxeT2r450bOV
dTaMGMjInl5Y2Wso5LpwuSXmyCxdUVLPljrrv+KQVBqf7jzHDV4/hH12gw4adI9aFMe8ZvW9qa08
Z4JOAJS1oS00VPFCEt8bHdzYRadpHe4EAR1/XLeJ7A/eSKP6w97vUPvJLcEfxtzlkr2M4ttNIGw6
XYJf3SDNQ3rD+GbfZ9VMaBrkHoXbLPpjmtrmIH/+pePBKU2DhdEY2hHHdc8fTuhDAJ219oVfuxwk
L8Peywcoa5LYOgxBqdYquKxA9vDlilq9Skrfvb9qOyuU1EDzWOEH0WnYwvbxptKv90KrodgW+FCh
ePVyTnCWsTF20mEhUP42GxrqFrry/O/6hMwW+hPjrh9iUeuNF/ARrRwhMvrtMqy1cntAxqyLz63L
FFFR+2kfsLQPARsWnv0GhBy+resSCah5bDL+rrb2WwFvop6eCZQRIHonVJasdTFyoHsRP0K9SK+E
3+/lW4zzWuSwmTK0ceqamJifBYlqjzjCZ+2m9tLxhAT3egvgq3875V3tv/YXQKjUhGW2YdpAen+n
gagJLmhpRZe3NlZC0EmRZoLRRSeVo+DQprUatVGHYclQp9d691WG0WH9H4duPQnUmqZ9R2YJ+yDq
pf6EvsCBp63aG7uARjufzPwWwkO1xdup+26g5Qqatlawu2WSbR7icHIEU/uvfcqhmNVGHm1sCmqH
MqINcGnCTc4RlgwlcD9OE44T9iCmftipYQHZf8GX24hiIZj4L7mOYKb9HIS9AFUDLqi0tFH0K48Y
P1tuUfqhTmn/KsNbdygA9CW6jxPdrB6i91EQPchX5FLjB5T9jv/B/kILUIfG1wytxcpdz7RY/wq2
pGKjRoDuxFYNW0FHATZTOe7X2d4zrk0utNEvSFDOjKH1/xQO2SuLXHdJPKdzEvFECcwkeQddaN9H
Kd6PVfJnyf3USF2uWjbROAx/21YP3RhIsIrVSVibQ3wVX6dYjRCv45LJTUqlBQlZdaciQ86N5LPQ
wVk1rt7jr2tVJPB8x4IK/np4GABglff1PoZRPbUECyRiJ2Fgj9717OaDe7PE07ObEpkLNbwTtPjA
Ya4S4X9JSsi5X8OKbw/kZS2gwnCDg1gxryFVr27cUAy/RlEgCYhN8nxu0LNrE99Fo9JOEk2VoL6C
NUssoptrVT9aAj+Et6bs1/JSfGp9xZ1nsaqPU7eSw777b8w8UX881WjkGfhf+baXxS32kFvxs+Lk
XlwSW4Fgv11/jSd3uT9RJh9FnDj3bNcamAy50VCxVXhhlTDjmB5UlU6dSZWKGDS8F7F5bL8cmxcc
faXF+HSOxq+Gcv5j83zL3/lcD1bxmplbwFbanEWYlkMK8hJbXzvcDbh96bGXEyuoXxf9WtXBDSQq
49gcz5aYu96PKxrka/LjCk8xQbzdUcEuHeK2oepcOVohIAvAO5lHJlSOR62K6OiyiS70yilDJCNY
cJeJIpCpGJ8iYndrRo9giULAfiiICLMh6eD62JENwmPhlEZgCBWp+LfunLN8kuYr3lK9Ru9/ADeD
ARZoCTgYUFo7dYv+PGz5qcvRNnfj4uyMwUZyD63iqPfnRlvixsoJ1KG3Dd3YUqaEvxwrWeOhaQgv
HMJjuFyZX/689+OF7yEge+oREQzSW/MLJmwExamUq1yZSCnKFCsyTVpgBu8xx5Y9+Q5yfLSRkZh3
4IO8BuoyWc1DSX9C5WINyNVW+dR6FZdpsKcYggh3byIV7bwAvPmoMT7nqCQWpP3vAvim2zsBe93x
8f06sjnl0iAPqlNqx+OqqI+4XdyFGqlMCGf9mWZ5s8S1H7ZXs2bTZqD7as3JrxKx/gdfkg9vN3PZ
aSh8RR+8/ZEN18JQP6dbEDGgWomo54Hjign9/Rk5ZEh/c7oY1kpy1rjgwhpYp5T+OtZQ5Vef9jRi
EeHKDM3rlD/wItEJZvXwdqYDyhfX00+y9HEFP7aGAgki/p1qh0oALP60nIrBqNnEOCZMbjLSGj7R
Sjj4u9I2kY3Mn509t9nc8nblBMfA8f/Jy6smSTKnILeblDe35B/inuFkrZ5UdsFvyG7zNRSE3gfP
p9YDcxW10Rq11QlnDSPFKC6PEbhEt8g39U+Jeqh3Nn2uufl8qis//1udFPuXZbY4SNXwmpcWj7sM
M/OsiQat4MgENUwgF3bS1x/9tUvObD1Mhqpi2McmKNkdLJS0ftviPoUR2KDcNTc+2o0n2Fud/dQq
2/0/jfFS/BrZTsO4ovI/T+qMeVqdWqBLbGdpnyxhdEDDf1a/x5wSyiT3GzxBgJqxPVHb5oEtfYnt
tdj6yMnXe4yon4++olqAn+Weh7gK3Mn4ChSzzKYRrP2bBmPvylCNXEKMWotxP7I7IML6jToY+8ez
upkNqcOP/bN5PVZBXeu1xaX7dMKM4PA73tF1V+S8WbfdxtrFt2/Qju8tVKxkqKBX7Cq2bX/faWSP
OMQpv8Ejzzx+7mOoCihtkxpOz8jxdKuTdiwnQFecnl0qM/HoheeNztBUiEKa51YtEvMgOtCWxfTS
9l3nKpqSfay/0ajSXkXeQijeK8MgIPaj8ggncG4jwTvCPxWjQ6KQipeYfkF8YDrrKiH1V42BKzcg
1shL/YLN4mO5lDZLv8CXk2tGHHa1RGAXNgP7yJ9U8JeQm9JzYaEFTSvnP/b9amoxMHNKg6b40VJS
QAKlaEdclRggrN8KtE2xWJOmhsnnMgRTqjobsR62q5kXsojj/ByeUYemHwEdmOb4ksj3tdesqLhz
1lyE3ZposbrS2591yzaCmZD6Mu9m5yrgIUa6mrLGKAYuxr1ApytFvF30/EbElGvgRXYFOSwD8tdJ
ijznjw5y72XmJcHGHtUxOkcLoosJM0PYB0kmTMFYUTks7AZQepbrK5HSiTuiLoFmIFEPmEn0yrSz
wwRbBx2kvrbXVvB0pvR81KbNLRuUJmOwJRIjcoI7lZ+2x4ytoe1iisz1zoyV/suVm2DfR4fedABf
IW/ppp0FwlOV2PBWtAwQJn65UbdlnbWypsc7zf1/a+9lj7Yq5HZwTjBtX6wlT/5MZjmKkXqw9k3N
IeiBeRBaDNWjsmVR6REeHn6UlzPq5rBBpkmO7MYfMxoJ7uRDeBBCjohnVt4GUnxv7j6rcNOdk/pI
gRM4zvg3vhXs3oVZzUNoHR8bXG79+1oySfPxIh9Eakn7zZUaCEUhSdteCDpsHEvEnPLtfE6mquO7
jN3w4nTJ2m+sv3re4yduS9t4PlWpQ6B+hysYol8PIHDZzUCXckxIRR7PZ6KBpziOp0LUpzxrMWkf
sr0bFx8i+FzgVTku1OE9X9/T+aXQACTnZDQg4dxcnrR8HCbLCV3UoRTiBjM1jKxX+axOzDYVWr8z
3VdQvKAVmwI3P+vVzZNMT1b7AOpZYE7I6DTQdkzlPrVTdneV1mQPv0/z+s9dv7TYL3FQp2GUAD6b
XWVzYYRMRgnOYR/V5R5Kx0fuvXjcGVzisoEjHOTAZYuiRq6FQBcSs+cn3ZGMI0J5Uyh6lmplWp+j
BnJ17fnwUApOQ+CN3uV3kVRpvjcfYd3/g3v1iquQn9VUSGmTaOtSXuljvR7o/Gi+c0hQPRah831U
MlWabBQOHl0evEy3W1BQDBv2oQtEqrqiyeE0kxFJ4v0zJB1unX3FIFx1/aBJSLsZxWaPDL9H6B5P
tcUJQEexfat0VIYWigYG2X4W5lyH0vU/waAY/in1WlCxBs4Guq/k1ZiA+HAIw3MQ0PWH3ZevYW3L
h/FyNJSge+JLK3mlmxOmDAeObJmTkUc9P+pm4H2AAD6HoWWjiPGupggXlw8Jcl8W649yvCOGsb6R
ka5gBTGDSB7bOJNzQt91Cx0DNh6b9PNKWjTCX+GOahBPhzZ/e0xkUvQJ96pqWOaB+HG2QKXPzHiY
sCE/xjFbgPkjZMnhOfgRDih5ba9przyhHomz5af+bpE3Z/4Monuiq5zBfG2iuNodPEtXnsF1OU0I
GsEX/XULob4Yjv/h0PZVpFJ25GldYQmgHeWRpoAMV87hpIVGbSzLooCz1jsDZtEf6qHl/8e28w0k
6SMBWpZWEvdg1zK1CvUBzSiPpoNr8aNqdf0IFpSK54uiWFu7C+Q3CgM2m5e2Kqq57E2vSUtea7H3
dzsc3meoALqsi8dyabW4IB8uItHHiRN0fxM/6iyvL1jTrKmj6J8EpLPAUiNBVzN3Gg5BxHY3zp8d
oq7o0gxd4OroPJFAwVRl1FOdP3/ZXsu+3pJ6Z1v1Z0dBZJq9ieHmUyiH/DoiqbLOGkOLcq/pkQZ9
zybwezLibezj+aV/OPnNLg8yyKGDMV2eZJ2wZuT/ruhzTUYbbSJXNJAfWMpSSn97S73n8hgMkWl6
tnwbyK9/UuakEt546nwDvuVD0Lfgjj2tJMQ7qq3jDLfV+Rek/I46ZBibDbxWjJl2tXSCFUhJDNtj
jZcDnh1wEfdNd2TL2aiFhhSrap00apsKgFmQ/WazNpphV19xwRtc1pIvQTjqnoQbfDHxc4e+dKE6
7w0Rk6tIkTfjUW+pVcVVC8lvg9Mb/g8x5t/Ql2T4p0Zcxn7kn2s3xHiOU2Gh4V2M63PVQZChOHEi
JifbbYm454tqfsvseofAaLLmvp2p1UqKR6LhOUtyNGMTnFH1AcuS1985a/VQo5c0W8EdnkqhY4mu
wmoTY9ACbO70E6MGh6NtBGyW1NsyPLSnRxJuVAElwwhTz4C3MnYkfgO7QgPjXkcNiSvwVe1VkATe
zfKlcxWk0UcDzEa+XbxYzx9YPMfdT+zIHhQV/tIcukSkcm8DI4nUArgDEZcTm3p/LIl3di47C/yN
ANW8vTYfIw//2CkQ/WIBjk2v2EZ4qw3hI6t5XH8BmlDEN9P2Wn4NWO83x3YIL+VoVCbQ+5P03KuR
UZRS5Iy6W1E8OANjlEcWRpweNOzeVr7Nw2YJFDY8vMW0ie7NhhX9S3hZWCV0Efs2vaVSZ6mVL8+9
Pa7n4uvz29vzdU0JnHzjy2MC8b/D8ncLIQJAzA2wO1lWduEMDcu68h2bJ/8JcjpiWBjjvWQUByyr
8/L8bZm7Xaeaxdm9aLEmOZqIRlamK6unZEa1NY/zj6Bibw9woLQ2bmeo1QlgaqIH7KqnhcTOkLgw
xVzetiQflhmky9u3tGx6DKl35GFBqabS4c8xWeTH2+bFqmGq+ghTsYuGcg61yUoZ9IiCyy2rLtXV
s2EvNWlEaGfgwwusQi1DzGZk9cED8d6kwxQJvSwM3w2zuTJeSgm0ZyLu0RYi6Es1J+HZBrbOLItP
b8MHSRuu9hoQZ9rt07vZv1e28VcBHoGgLMU7XTPI2dZYH/JoXWsz3ACdyDfMN4BYKmkMVAX2Dxf/
KFPkOfOeJXrOFpxOeU5m60oY4yx/Um8QFGio+rOLRx4MY4pepbrTxw3nwGENapkY7FcjMFsn1cIW
8PgeE1+rwuUhF/SHoxQVSNMCPfnm4cC0x/cqBFofKGqwpiGwkuZVBbpA4HD3k85GFlSJvOvsTm+a
oWl6+KHgHu9T1Rdu7+8ZyQczg2UVJLRJUJkIhVfcx4OSy+ZTz8zV3uWNUpx9ndyWk+SyaH5QHAfE
5yd7hJQpdQ/4awkw2kAS4Go5YPuZwRMvpWbp8gTGEaIzMhxdjw+q2GZDTk3c5TXVSDH0aUjGtgrj
tTFxKBjL2kQ+rFO8el6ovj4AmhHWFvG08MWTOSxDlFIE4nWeoJO1/2j5Q9NK3/mv5Md3GGV/15iK
KwWSrW260vGlBmM5wanL4u7yBDs5B/4bH8aTAg/vsJpDhYpiEdDrttrQUbAUVI6DHhfDF+6j/IYK
xAYQsw2/W6MUIdYktVuBN8UvjXjLpGQrFaU1cj9p0jI2Gz5KkafYD76ISI3jNzaAV2E52J07ElfN
lKQQ1sBWIRTfF7Cbn1q/kceNkw6I6wDrDPYZYq1Q+4CV6XT7Pf/GNMOZnGnNM08W1w1P6wMQY9yu
MpcICWdmHX7X6SlVrIxbw6B0hHU0RfEs7ekfNFts6N9Me9YNaGwnRtscnKsRJtRsBKGRSZx7L+dB
2S/VgTNyNCDqFBAJNvSjfFUan4g7gnqd9LwxPxWTKZD21cVrogl0QssxA2rgXDtn4wMNy3u31wrN
rCmxG90Tutirn94z01HQzrBli/ua/J6AC7E3anwl2AIPigrfrZLrAD1T7+3/u5nXXg4oAqvZpRhw
KPVMK6p2BADDWktmPEFNqLmu+WLhpEk+wy8yKEd2GPF8NPx2K/5W2gXcSExxrYLdjzmVDQGKqnjM
jyYczLmtwM0smtEFFNMv7VReoTQsJjCROtzbnUez+FA6uDKGAcXLwF0ut48hCPKuaFeD4ycyYExu
3pH/kGK8RSet3ew8jlfEMwfESSYOnw1kMbEac14pXXbBJG/SJs0y7Znjs7NORUhV5mjNyQ+0bK18
6XZKC2+FEPK6WESf2TYq9q1aeZ3AVsK2/ZfNUU0VUWr4JikN/d3138sNzYLiYFDVUBfdjV2bZKYC
zn0UwePbKRkZZhjib71QVg69uCX6WKLonSyjxyio7WkfPasQJV7tnKM2OyADLalJF1OJC9hrhRy1
ZlaL7ZM+YcZ2ka3euCqSZgvFlDfbaf0iOzDtRN7+1mTMMF/rXUOs9ZTnMFkEBwVf594LGO4iTIwO
RYwtvRLxktXQh/MRasalAvM4vk2U5jeGJVBORVQ5nbsjkXcChiQMcf021NFhSPlq1ckazGZ6qqB3
HIUuqeGYvZZ635869eZEfBZapQdu2Mwt95YZpOOSh1HIqLTCemf7QlycskPYHX9EkHphI7IHa8IL
M2aAetFyxJORVimUzJbao6yL00JiXB66W8Yqr2iO0evjVKV4ZDDyxeggVFMxkItO+nd3qNtIvoCU
8xAwkfkgljGwihOBQwQXaUgKLqv1pkRdOshcUSRea3ZqKiRI/3tsOhKHM9e8RD1JapWfj07EZTFH
DI7xSvWWHVLF76xytw13/S+aQD5ikD/tTgrpoajNFJbBfZUvknCKitPTxxQHI6GaaAOTJDFLmb2U
RM9F8lME0DZuie+8e15Xw8/216lJyrWA7WeIEwb4ZeH5snMB1Sxjieml5G5VZGYN5hXI+rKzB85p
jLSCyiCh2CrNDduDHKrPMc/2KlDvOmR4vMEIZhYqjHJDmZqLv4KrbQvSP+omzBruBb5wE7vf4sWf
v2fHY26PSdwQPpmkGeMRd1bP7kwsfHNqowQl14fq0CllmGRQRcUuq2rwy1q7aaCaB10C3WdrXZyG
LdzJqHDsm9dYwT5Xs7XfWHx7AMDriR8vIAzrUjIcwfdcwzsiL52gMX2DcjFbKdsnZ8p2I4U45aho
VI/Xl/1jsaV2lFz+uHTn1J2RajZ02U7YhiWBTn/aAF+gZ5JMtwLScjS5wUBJ/6fDQzwHbVm5S6o2
j/x+cqBAwTWwNJz72g7ix/u2TRDfR9r8MuD/ZI2sIjC6GQCcFjyvbXK6elTgY5opbAKLlHoseQas
ohPVxyiPwbdpCiL9Us6ZG1tsOg9kntXfmsnyMBUsQ0yn6YMPzjG7V3DtIricb3lXNzY7XLScW+0H
gtuFmwzmCeUwDCWZjmRyDViYJTRP7gKaBvA7IDlYJcKvsG+WjATQ6RUY+3uNzC4s2fFS+KqDizfC
WwGh/yWeZK/5gHhO+pck3b4i3mwb34nrIb3ThRvnJEYDpf/i6nWLHBvrzkzNPeel4iBLK3esE2Ln
NF4e5YgicqKhiIj2ifr5+eFeQuNW3dAT5k1K1Xh5yKMnPM2YB4d5CuSI/+Ycg3YMKLWzWUrxJWRA
9UJh4AfPYpGd3uKqzl4k6aauQwGebbF4KyfN7b8/4ivdZfc3s85d6zoQkv21chBfodRd60w49pH3
Im8ZJA+/yr7BmZzMFo8mSmDUGfDKJBDFdnFppHEVSWOpuI49Ma1cSFE+T9hLNHugIwriaQQ12nmZ
4YXKZVkJFLZdackL2RcLt3wK2IfwB0wfREr9HGDphHI8L04c8/GOO/MnRrCKCVuk0iRT6IKTthpQ
jsH8reJZxXVP+s63hcoZPPIsRRm7ey375JsjWbWCIioMSa1frPObfB0bKdWXaABLu6hP3+1OoVN6
2pVoS5QczpWCremHKhnz/fYpfZBjhjnezHwZrZHjNipRSBGTxQWNzHolrOuUu1P5DxnrzPa3Sesi
w0wQdv9Q/RjBdDDMzU+aVXpW8YmxeA8Siv8tZFEEN/6PgdCBwgxz8s4BoEAEh2OPETUloj+8wNai
1hhpvTPHAQURYbkEt+u/Ec+DM8z7yiDBYTJvJuTw9C49JvgHmoLsLtZSXWlvyNdwxVGP6zkxnb78
UC2qSdi/vyiwy62dKYtoB6gz3FDp6pisUSY3EwCpCGF+N1aPD/MNoC+7aaDNzaq+PqsjcO2uBFrh
7xJxvJJ8ngxpt6ZTtTSPhY9e9O0jUJgjVN9vPLwH6z2x0LCA0gn6NDNQxuLv3ooe5rVKRdMVtzyG
35dNw/Mi2bWN0EPH01uBX7YP3nLcHQS4XpnK7m6Mgd2Bh1T+Kpz0bzhoPmWUlbZyyuzfrWF9XclH
u3mAN7gy/xdOkJRZmTNDK0T0KssaBvXcUXn6cFU+qhVad+DZRsUo9lT6chV0nwtIHL/ox5js0fOe
kTE14qi6EILmC7wyDxlY/IPbgRyqYYIhYc0oy/isELdXM2pDSizK1LMhJA43Y3LN9cgdBbO6BVSr
HqITDV3BlCquRDMPbinOiLfa7HnCViUui+HQkCgTbcuEma8PYL3VUjhFNjnNYxym/RlrIASj5IOd
hw+Mluakt94zP9unRd+21lZPcljeKFNi5yhkHsz/kOVo14rrjqQwzhSeMnd2mrIgKz/WAzKiGCUa
ra/j/5rr1ya/Wudwg/aya8sfhHPNdrxm8rC5fFVnZuX7dEXym9ige3IgFSlCSxydOTkHsI0e+Am3
IJ9g1mxWuajNwXTKMJWY2t/xv1LKnmXInmbCPGdUinnnKWSxulATJwGDCqzKNdFYm3BvqFrPl2sa
TPmJh1NraRWB59V0gahcczLNdEG0JCXkcsOlkhFBjdcOk4gtSemKZEWoOoBe9gmr892yZgLUFOMp
p8mKFuNQ1RqtjSZ3cX75wsxSv93fDYPBycxRsY1XxaMesqBe1lc/VLTVfbylU6JaY1EAeEc9gji/
82/VQUovfQ+rXcyIz2Qz/57y86DBHWsF0AmV1xCEir9oQE31s+i9MEtReXKkuqSNEOCKWEdil42m
hMpsneAUzDMObicic3F/4FK0Doi30vtlC97dvQwdCtHZ4SPXZUn/rXuClZI1DFWEaD9uMxwLRc8M
ONl9Q/eYaaBjVzKWAMdlkpugQJVNbQOyMmvbFFM6rdfWmY3LfMdRr5/ljbZbM7ry0jZFLbJrCbuc
86oq60od9tp+AitnjSsSEnphXmzhFb41WcP0g9HpND01aGXipLcBkKnRw3Qtq2wmHRLKNZFKbLlJ
3pewbRyNw4Weklz2b6GIRiE3sgT9PV4heeFxXYQV2RE0ShrtbkgG1QzDNvlI+OMxguqzoCyCAf53
mcMPCgMIoXJmym/WY5pOWgFsrAhePhB6SZgP/i6VsM9kjn+kO2t6PX3kv1qJd3B1Wgwc552o3Ezr
QAdGaAcwZGwQm8RIY1i/PCqno8cooPoEzTxKHCFK58zNrdPQIKwk2LycJyCNkGMwb10wUSbI5JfD
4d16pKKWLi6BOuIlhKWLvSpyoCbiG+yyQG1OJnJUxxuiaIma95sI+ae9rDj5T+FctQJ4R2p6R9k/
xkCB039GVx9UblpdXRNC74VcBovKYaUNNjGFV9mSMbIeK6wZWqB48t3oKXefEqDtx3Np+evL+VGP
a6nLIfpstxosc2Xdin86ZGKsPNPPWvRth8KoZW3HUB+zTO8ElR3bLC7weU3SVy7geod9pd9gCfqm
w1zzCO0g29EjpsI/l+YZ0IXF6oCZoQeiHzSLlRhwjvXzYiggk23tDk8B3kzkw2bsUImvw+SYGklZ
xybydRebEOnhsPSpPG4BZfEDONv+5tzpSvmkfbImmB2WSXwdbtHoP5QKT27yZuIezgg1+9uBlq/W
ocfNAZeMxU6m+xtBJMjeUwajmPdsRzCDAx7fnwGlcyQPUDJjUjtwqcHYXcdH6tnJ/KZf17iVjNnX
phlUhW65ccK+dcpB9OznJz2+YwUmuJypcSFceUcpBwclXd5e6kw5E3Q1paYCjiNsCZ4+ATj/EYOW
d3+kWbSMnOfbNGEYfNLtiMXxDkLxnU5B8chCYninkZsGbRVCV0gpQ1bv012r5itAM0M/AFFoR2wc
XM4F3Pf3Yv/EeS9BuAru0tyEzU+r9bnmgd4U3Dbb2ub5VX/ldXbq9SeNO9YL9rYlEYn5VvexoryC
uiOcLH6zcxPyD12UW7miqG109f+p/l/GT8u9ee+dOoPzJZUXXHsDYLkyrXAjIFyou2wf3cSTSPoq
Fq/4dF0Qo+fD848WSMyONMj+0aqc9IgcMs/iRtT5LmN3AO0BurgDu7asw7kmZ++eEpnQzmlUIW0s
VTsj8WSraJvknoQC1DU3KNj9k0+g4lq5YSp63bnUkvUVUwb+rZ3t4IiSAiKxBFFYEEs3BV2V72Lf
lpPLXgVUCdomhD7lHDl7BxAzMY4B/YXkUgG/fLD/RV768l6zq2TWnR3SPnUw1q6xx6HBDMABunws
ATuqIUvoN0ftIZuT5k3ddJmU9DmZ0WtMSjvZcIy0xUX2y98QBdQmugFNKRA6kMQhWeOjJLAurtRu
SPizZwNrDtqO+Iy0BsVER3/2hm5d4Vwng0/8EMXuicH4KunxD/ZvZMhb1LN8zlC8KdNyA6QjHuTE
L/qpHVK7rudJW0OAtg00roHFYnN35e2mvPg31DzxwRilbijqhvVP9DSz2zeyRC5O9vpvReQoANaZ
qb5txBRu0JW1u+Ver0RUt5ZVcsI3sdq4otRwvAIJAAZQ4VNZoGffTXEIyA76jv4SILjKX51x0Z3h
UhDPHSiv3uLleTVUmjMozXqZEXPQ4kZ9Rp5BgC+v5kjM0pzFy1XBmwmlCYbpFdsI0bklid+iD8w8
1UMhz4LmnbcHXv+qrv5ldTCS/zDRqS720P5z/kB+fPY4LSuKW0G8aAALYgyJT1QdLLSUdYyn2hRj
IVBLksUdJnaWt5vlre+CWdqPkcn8LrTazN5k4CWi+39QsgjRX3SeFiM4r/gnGKkwVEMyPpqciK2w
FZF+g5CsGJ8u6Bixnvx7kUZJNJEIekxgCXCbenW9GmQ6sKSA18CuATIPI9eeffz4NxK/h03fTesJ
FJzBidWAz8f4ZCpLz3JlcvHkV6GLpRObs2cjODDn85/NSI2zJc5L1Vbj3ddiBjeM/TBssDs+d0av
ycqoBImUA/DaI5r3Pa37b6ohnaXB5BlRmhivJ0rUj7gvwRmIuaT+QzyhW+y8IGGplX2XP3I1iWET
W9+9v0r3ODFQ32Zl/k31VQiULNRwgvSRD1YNQYzIVT8y7gF96zN7xykelqBZ21Xh5YXtZMQfBGfV
zjV0/peEEHFPprDU3tqKcLIww++xqQKv8ops0nw3FTxAZva9t39DEX+yxYmkSKIOYhEMRyZSz2r6
TvXMdxuG6L2KGbEEyHds8pc54HmXqoM/Ozy/wo4M1RE7l4g14y0uroV7NUMrJ7H1yjO+NVtF7OYO
9ldw0B94MBsixFfcUK25eHGzPvN51ll5gxlqhxLPQTkRH9RHhzPHbLLmHzZ1tSdRUNpT4T1qwVzQ
d0Mnl8IfKZnO0fZeaHWhZ9wBen3fCeO4YKdDYjdyWPgJMOX4gs2Sb2dom9AqxSaib4GVs2VmroAW
NhIgphdQrjST2+jMlq06rABt5Cxsf2nkNAHUJJpf5NNNbmXdCZKjMHmJvB7y/8e4QiUAGgOhP0Mt
ytnUrJaAnt5l5PICS/d7OVd5RGG9KeLppnTBo5ynyK5QBL1hDpKWPWCLWTfjIasQwGa3tbKBZM4J
aB7suma8Lt8GpSIBMQGohOoFKqy5hw7dBNyQ+6Pa67w5k3Pqc4Ti5iYpaAlJx2yR5ZZAMyfUUbJu
9yT+fKogUDtRh3erNBnArtcu6Ds9t5tkL7Y9nVOfqfR9lzHJRWBq4t5K6cYc8eMRVc5Bjg8ZwW3y
H9vkC/irRSHDxnwXucr5bSUxvZ+Wdipb/i1TXUqmUPV7ve1/OBP1ajqUpLdBXjtub52YaHiWLo8E
1NmCzjNsav3QAqqvxrN7+x+J54qjW0dAe7LAODLiKTH/7Rofu9mKR3YGCwwMA5JiOamSHNJmQHBU
GkSrl1Pg5IhRLW/DWNaWgbYtEecqq+VW4a9Du4L/ov6FR/KjjYJJw9CnthKzUWMQ/ypkWz56Jo/F
28G0Gw9rM/paAI5n0xEkq7DbZ1iwMBftM/4eHom+X6rgd6kgGtXVlvwOv9Puw5XE1TjhdVsi/OYd
SVtWlWc8RJPHd1e2Mv67/1CAnCEAGggM8v6zU/sIkTg8REcPO211HyVg02mbK2QsA39jTVurFjCG
n1U/MV6qMHb2BkRUKGmYkjdg6S/F45MWTVehhWbYs7mP3IqF2CKSPM+3iN95kbP90feYImGJ1Al8
L25fd6L9G8ygZ/o8w7GZ965Q9XS1qNFxB6vblES+7MXWZWyoA7KnPsr+TF7NiEdi5eDHQ9hg8JWA
L5vXwS7pSFPjNJ7FLn+UspOpLx8bjiJEtWof5Uwqa7YtNUZfbT7TfefMwO5gTWd5JNPAea3XXHQ5
Q1x4TBAPRlTdQ39RAzGGGpOtdBHjEQ6+ya3iCGhJUojmZ+Ahs7QerdBTbZmmPdJ6/uTFgIo/visB
L7m4ohRRBFruenaGj/iq7GbZaSJZ9gEkiCOZDIUq0X8aaS4Yq7iUaZlKZiom36/OPwIElQnWkexc
H8ssx2RksaoWbErj/LFIob/wSOO1L/hucEMc4CrIjGoIAgWN9WvZ3RtbFlrmFWulbHGcIrVVD7JA
46+eDFIJZl6L28USihPDoyLhZp2avpdjp4j0aXlqIRUPerhfo5HgxU5CmmtP7S4/MigYCkfjwvyp
CNnEupfsdcyKH6jxjZuFnnLxNDdXIkQpNz3srfsHHN+T/mt/7GqOo3w1JroqsjwA8lpHZX+1zIQO
QVsPxqVff4MkW81yBaaJ/KIkmKpyOSLNws3DceZtCoDtxl2JyeFBDftzMJ/yHnK7A1CADIUc7Nh8
LjGkrK25dL3kzYRe4JQIfjzBS0OrmIGkbgKeOZxwwrJdXjQZLmH4UuNpJnwfZauMTYZ7ns9o/I6b
7d29qKggK9WXS/F3jxDm0ZMsZJ6BdyBLB0JtpCQBjLrUWqA4s4ffRet8+9NlMccx5iYzO/4+vD7M
aeM1rF8IYJg9kF/9TTTHtabI7krxLn/wKC2kr1T/ZucLJfbhlfDXzH4BZo2ZKAks4NH7Sqsy1OYB
YqQbmPaidR3YPQ88NZn0ypBFeGAZr9i+h/BdL3uInHgmOgxhAo5D9RtI28oyr2HdoscQEUiimasc
GGIN+iXTyvybrBHz0/VY6T0qZi51pY3s/kgQk8+u6vhEnJr/X4RnE2IfpSBJbQkzNM2xXZ8gfkzl
h6h8ce/S7UKnmv/6ePk2ZATrSq4W1bQUS/zIMSAxpETV+BRMZIv3Btf0mNAsZujHDfIvox4U5D97
7yMPs4P+1J0WBYGZFkSs0UjwwsUIl0DSU8R+wOU41JaZvdMrbvKoYW3prNi+twTZ2uQW8Veo2Jm+
r2jKlHN9E3HJocSUtqDVN6CrpCORrrQ+1Rm1BHkU6sJJujZrc0l8l2+O5TEpc2J26saQmhePZbWL
jM7pqMOHJ5iMS/uujQrO+vxGcj280y8F/XfkAHvbV0714+pFKDHuCQAHx+sXaenzaMiTPCOCBWR5
UGeFoTamhf7g+7njB9ndJLTmNK/7+I/pR3iXETl4ztDwETGd+lpy21YATwJdOY5orL4AA8Ohpspx
fOVYRTaTIQCa3bi5d4tDjND9Ci5ns29N99XHQSwfeJU1XD4nn2L4iNVRL2jlQ5GffEPHYTOgnwOC
rDA5f6uafijhl9J8YZte8X4sSaCw5PuFaHsO0/ZbN9uBIjtJ4hzGkTRHjmz02ef2P/fDYFuKkdbl
TsIoe9h/GWjvSK+SkKdh4QhEtIlzicw4Bwm1EkMh3Z0XywFUMhiluxE5CveC38AtZFOwEJ0E24Fm
TcS/sInp1jxUNCYhQfaG1sr7dKmkKO+bsabRvVrk+5pKL0UlZhRJjx/gALG4lDrBoCDLIHAMn+1J
b3SOlCsnGE7zUwaUUnEWC34pSuQMbUjKDE1XoPeAA9jf7BPUDhX3vI+r1ZivJTAOKktKLRn9XUfr
TEh9Th4T8TF4TmxPPOlmaJ06L/1ozqJPeitO65iqpGb8mnkQAZT1uJ5Ww8yimEb5Wc0IH2NQnEAc
b67d2kqgAcnUvg6JIFJ7N8kF/WpSKBUi5rrhmAc+OVx7oETGC2RoLT2mZ6ndVo4kIv1jzCd8DY/o
8k8NEaIZ4iJpcEMmSdtMIKbM3F+pkqH1Q/721hZSHH8Pk1YMgbpvwoVkVS+0/SLEFvOTaxC9UCAj
E4acol8RlReY7D/J8cIV5nli9Y8kXJHaGkQHB3FZkTA/ryZxjL1jsasP3HYA+/VcaSOMbETGbTSf
5RkAFjFAgeNiq7w4q4GTJ7hCyVRMFn7j//8wgpEiHVp61gzdjaCTOmFzXhUlXPIf5BGI6zrSxnq6
21j2XsVG5MUaUyPrFherkp5nTp0pyYpVkEYjhjB0/VKK+DnZ6m5acndy6UbigjdEUjOvVQUOnlf1
5zLFr5V7c4cXoDsAFQNPTnDNp9M6EtqRbno7f7w2oAqVtG1qb+NuS6kJogb+AaxU9+dqjpFO1my1
tyXlW8ezBkWGdfziY6gf0AAs1EHRu2ooDut6wK592arm8X8l/czIVeLuCJRfGsEbN+gPJkXcEl+E
1q9w03A1sGF9fcx17+Y5a227cO15EPr//NImgkuCUgpZX5C2YalAy6D2hxCKrN+f1vjQWrxDWmsE
UtMZtOnKIGIelaTHtWNxZtfFvCAaHCgsAKO/Xra+7TF3vG3S8o0Ip5sT38I98s17u5dx3QoE3sei
Y81Ja7u+7ImWmxoiORWzZN7MyaBkMzyG+1ETx38F3vONzppSD/QFLlVtoGeAtP+dQhlliMkKFmbv
EHkMSa8hHivibmL5RbNsKib9rkts/0cxsDNyauQFPmqvo9c+MBtH2/7kX5DJYngfG2gh710wt5aW
ww9jecS76pPPgqkAFqQL/paY1rIfdXuKbuZsz9+KBYj1Df8t31agQACIEBAdvSgdIgEWAGsUwm5P
KSGJ6eUSaaBxFHIFfdFAvRJTVPNk2PNjSy+P8mdm7/k6w9yzfls/Xwz27PJJMArcjlG738tVqgZ+
Vi4kQT2gd/qAE1K5b5eOPUADHHzbThq8N1+3/182cxfNQIBFIP/gwuWM0cfVFrFKwijMx+VjrXBg
/PJ+uTQuo4R/UfjDiA9HxSG98ei66FbjiOkxbrL2ldhEdghAMdpe+XGeCjsSKL8E0LjYq/1cuoqE
P9zJdquE5DxglWuA6Er1ESQQqMT+g8ONk81BHg6eA5PCR2ITEXvDvXpcWP85FbuBiKZ1B+9sLd+/
E4WHHZ5cEKXo0Jtbv6MCzN7LKOFPKob0DZHrghNhr332vXdDa/gXa89NwC6SoLx3e/STzVSlTKeT
ddYuP2JLeOgNu6NV3SmQaZhQHmss7zU4YZce+Pp3O5irI60MnDMfIR7DxFVoz14iRPADLR3o0+KB
H/Cfr6wc6VEqG7114DN0mImEsIX0Yads51M3ywnq3EYykgzblhdQg5NoPBRVskDyI00TwhAq3g2r
n2NkTm8hGfTQ83ZknNa9UMsoDNihP/jm5P/NPtR1EGTEcYGny2GhBYR45hKwbsJpWsyWpE3z2lM6
ZRJ4MmY9GXkdtuV1n0YMxxL9USwgWVFlbuQkh9M4s2q4mO28uogKtDxwfdluTDlnEEGs0I5B2M81
mBNgKcmJkPnSnn56YcvP9Vwi81yq0GWEC3LLg5Sz0lbl9X2vcVLfedM15JZO7F9sWKIChc+nO0Vn
IJc7v3wwLbMCtw4rUvPeXNxFm3zF1Q1Q+7fmt4xtd71LdHeyMyFmLxplznKubY89LlmrIsydhpW4
sJDssNPGKamNv8iKu97S2uSwjniWFl6jXE/Xq4e0fv5CFdd6I+1pXijooCfzWi82Dn77W6sS80AU
TI93A9YL4KanvO7+PTazmHBy18h8VLpYNDJactaB9aCM0Cj2u8U4qzk3kGVNlXOTeTlGyjD9mGRR
u/1LVxkKJIuDktCCZzLiEeKBjfdXCl1A74HmKhKhLkux3PXNK9wh5DwiqVNgP2SLYG/P3QJS1I+R
8bl8ATmIuxIruZzDi36bixyOjVjIOGmFFQF4mqpV8YRA4zZHBhIzEtayqet/APyCL1W64HhGYR3f
ovBRBf7gSP2SzF3+iN8xYoocvk0xyJ0UV8JXrSWg9Zs2U2m7Gxt5RMLE46u5X4tmrB4HEIMv506J
4XN8BNDXWM5opyEKnhv4J1NAnTyWzQknYkWb7AEhSk6XAToKAEQaUQLfXuLCdZ0vwLS+E/U6n5Ik
dz7B07CCFJK99JPS2zFhlC4zILwX6K30LVWa6yPjrmuNSWbJBzbGDz4I9Zlk00xvihp7n/ozCQlD
K+Pq1R1C5HTf5LdfjQrrDmZ66yFa9foqfB6teArgfF/78myRl9cavNgVxDDOVAE0UT1GNSXZPpXM
Q7s40TN2cfrJCgCifX11BachGzVYeQRdZLRx/Ivrbz7SKUHylTai3JRvVTW898mU8TPmJfTf7TgE
1EMmuUDevbXs4dan8Qu/wRMegPeA766dF+LT/1ocYUxPtd/Nu8fNe5QESotECo7cO6OCyRWPdYkk
NSVKNYA0qmyV4JvFuUrLk5oXrbrv1nkK/2SzgSQ+CdOf7pD6HxPkMxbdbeKxtO2QaRZ+8lfuJ5Iu
LeAYZIOhP8UZ7fi0e9vrAN/CCvjsTWNh3ncwH07pG1xF1YDgpQjlPDBaEG6PwZsJvEsnhW+p5Xfc
QIX/h4GsjBtMBgrpDeHLrU5HeH9Scvg736KqqeA2Sp4rqdAjoSjmPSJrxj3aOKhUkjsFlAEDbXOQ
vmiFqtZX3NgyDRIediH6G4PzNS+4fhALl3RB+QSbQgscQanCGz4fkH6Tg+wBXU8h6NEtbpO8CHSc
HrRm1Nv/UKHvy0N3GojFqS50GiYmuxS8n1zrwMWie6KoWTFy0ZsFH+ByG8u+O7kbqJH0a2M2+5m3
R4c9hDhqRjl3to3OZpTEo1Aon0EGKoGhNWYu54bZQIThC65is3wn2mTCG0BB4T50vvIi8Qk/XZvM
LCFWU8Hj5hJRekjx2pLuFTA7IgDPZdN55PmJbvyLhYqUm2EstFV4Jj0x9fVHOKc9t1wzozs5PRtN
Jh4ezyKLBpX7SSg4+pjRes7YF+ipsPqUjsY9CsmIV42nr3u+vI2BAWIyYBEOCVognWDRCxpZ1rlH
/ImzG3cbyaDycHfxHKIl/jQsG13KAze23k4Loc3CwKuqgqILMqkYXw6JgPbzqj+1UwJrhgwV3Yp7
gCGAOdjzzznEyPPxux79xtkwdRuQa5NbBhVi0zKSKBXwvqq3F2cQVKImGJEpM6IpBUQsKY5INGQy
Qw0TzlzJW1ozAlF83TUa70d+xgtyOdV1vvdENZNaDeD3gVRTZII4IBr8ZWcUcqmLRnAFnrG3gx9m
UrNfLqaykl8+DW+caTd8CL+0cUsfQEEx8w/mysGAzTQ1G3oBKWG2Ua6BkRkeDYL102aPizvE3xEy
bmx7+sX4WQEGVK4LEix7njtS7BRimNuLxfAuD8lm9XS/UEJUI442j3UdLGuE5D5CDDovkOl2QdxG
UKMJP6z5ltiwa3dUwWN2l71oH+uWjn4EwvmM3AEN3X5gSkHgYItksbVG0XlSfudR2T5+CWcJPdnW
qcuiVluOL3u+jPPBzI0kJAW9oJhm94qUx+gJMV28946Pi5J2vKM7MihR6vDzLEVsptQQTGdbWUBe
ra7kpZWh3gW6vUx0sZ6IcrhwlhhdObl5DITpdXhRy9NOduJSp9xQBcRxSoZhIfe7njkPSFlstAlT
B77gIfBpmdvS6+pc47vHxFJnKHxYTIq/CAcHYEX8TnKeWzPlrgT8wuQCAI8nr6U8ls/zs2xC7yei
sUs/2l63oxBSIllxaEg3G1ueROARV2RnIx8r8cl2NRmyeTNsGy2NDF0lMK3042+TjxLR/GJW0enV
iYExPrQ286Kz/g415gXZBnWGvrQm6simusYTEa8mbJyjxA/8/VwU2I4W0VTjbvyhGMsq8hxtW4tL
KuF9XKGfHB/0few6ltTEN24l0MR2VB7XrSb86Hve7EvVGOv9NpQodpyQnxku7QmJIS8ZpFmWubeg
kTp3kBO8G9xxzmUx6yHCG2mivTCBCo+D7NRiTS+dJfM477RBTW9+6msX5BpHuKTzvBTjthisZF54
NeTjn3VRT1vuVPEbI611ABAWKvBX8tXK7fk6jUyNXleD847CdfTyHTRfKyd7plHf4OJ66jlnRpnU
oj0yOMTIJRASgO9Dm6ZrqWhl4StYk5qFEAHLbUwBNQo50MbvSpNfvZskYtSzNlQkCCiyLCdIzgB9
TyKIcWnmJXWIWBDCHCH1srOPNndASeISV29UOowHiUDMyP7J0RCHZOIPec1SSCKFo1T84I01inuD
dXMBnRCF03R+ZBorYLEKTdtbJbFR+7Ztda54XtpozqCm9xbeIKgP8VjDies143dfQnrelnFEqKiZ
7hQfe4aoNciEXiY98jmgckCvWdHH9yhTKZLlog/D+paM7qUs+jRbqfLU/QmZHugX5g/vGcWkzqsx
VPcZXkvWAOOnq4nB/wIg0kIWXkyPA8caEwIK1z0ENJiIQdLAZdcu+CwlDUkD5OuMY+KyyIKAxa7V
66Rt8VTn724NsdUgN+JgwFYmWnHrcNwA5KIRYSEunjcwspkXD0HPqAQy9ApMet3bsJ0GaS9GQr3m
8U1Jiyh008Xi8g2KMjjk5h8BJA+OYLlZLIo4QhZyxXycraH6kwZrE++exqDW6lB1bKoBjuYjXsV5
Xh54Ls/hVj0bl5muJfFw/6wSu3erTID3aKFo3T8qpvlSpuV0Rd2+nh+CaC24CP9gPvArGF+S6wSl
hNirYKNnTESF1/stzWBQ0YZlDnZkvNxKYrI3/gT97RpIaOsd1TNBvAu4vVPzFDTNqi9OBxvr1tMB
lIWkRfCBJPZnybz4XVTDVqpaylGU63TFnXVqojGDvtKwyBN28IxyNgXef5a9RrzEHruEFun0gZw+
uwRmmA+TaGkqk+2/abg+SLkscXT7x2BzdcSEsRZq2GjTmb4Tm3eWg9JR1tvgDL30tv6ZEaFGaiOe
4JOs39fxCOrQze/SWAUt81pOIduJ78RjorBPMy3KN4jb3HhyNzNMtSgS+zVTjh6dVEVZ6/g7Ps5O
uWN04SV/5KHxoRvVfbOjcOAxs3NCLvehqlTz2J33Iv5q6KJ3tTeYIp3hFbS+e+mMH5P6ZSoeCgCZ
UeUaOlLxo5O9l8gdFE5HtV8RKdTvAilrsqEx4IGnun47lS3cv0GdTxwlAZWL5V4FT5Kl+mL7jQ1b
toB9RFM2BDTPXYIeVxUm7FNolsAKjqp7G43SyD6HQuSYAv40pdx3O6//J+hvncMRWUEqZmImwDHH
cHj4pz1CC/ZZWZAH6RWZM0fnu5iMTu/OLq7X4EOxNYaLoiUd7CVYj4cE9+FMckdcVqbH8eXAfXyX
Br5wXkuZCz8JtlwY4WNPZjyqm/XQ5zK+5rxOT2gfjC9lJol2ezqPqlx25qcGCI9t5g8B0USNBRkp
muI1xR97MuG/gsBbC7vxx9k8UMfh6kk9kwW9Ksj7Z9dXT/FcJtHPeU7NOFEtjVv3u4HQVlupOvBP
lUypl254gf4XRnmh7nAYsWPbqd/Gv6iGSpnuJutMZ+O5KubI9oe4YnkwHn+EBuDmAInIN7xM47xy
A44TUNSJEbH29pGjg8JspIfU1PR/dHy4tf5CyEvac6KfV/FbJpj8qfDqLZesJzJy+oricCdmmifR
bjbMuIudPFkiFYFSKwpcskM7Cy9Wf9LI1JDUwDbhzPCNcJR9gxZD+xzAosrq3GYbnZw33dhsj6ly
0qAXFkrF5LGOvBRm4SM3Lep62xEn/D8PGzxmgeqPBtlJtt9tsbY95jYb55ur6AFQ6Gl906KWO0VE
9Dfu0cFKPBO0pX/gz1tUCH8RXw812EhRb9Ks8hQUVoT2KM1EGxC+QiyU2dX0DfDKTIIOrUO7IONa
YphT7QWxqlznXEHQLp8olhTNpNwt7GlEzoRuV/xunKTMGLGbxq5uegLZfpbwF9kFmhXXSl68BTmp
xFaIVUmQF2KuZr3W48H9/5knDlTu/NaUfirHNorwu9XV9ugPdNs4OBamj8ho7WFYCj/MAhFg2spA
NRoWrXXK6tJizIOqZQMsrKYkgRAZe/jnSH9iSPxhX2ZtHZ0MGC+tWtGluUguNL23IOlvtHZXce6L
5Rt/bBJ7n6ytDPe4tQMIRpUpPCWEfY39ZNuOA0zrZQXbh/DLJTny5iisjOOdSJ/ByGS2m8sk7zii
0Bfzlp+RguSlpV5QaC87u55BqPT6D4H2PMbKJAtuQLJGs3HdupMtfgauBOUjKOU9H0HUY8ntgATR
vJBqgi7ac+TCGxFxFDdyTg22A1nFvP7KR4HBczzX4wXP8E34sAqyKgm9Z/h2avwNDuOOnSxD7aNK
oUp4WZOVVVn7483CSr0lBXMl43eVkDNSeStwvWyR89g9rYPe2m31mMKGfQJ1VZL0e2BaW3f8U34n
mi+YVeJ/KVXgI8lEUT9PPRt2ldE8oqgh2dh+9YncMxDrq5JVc/s03s1OpfYHeIDzcqmRMXq1PG0l
//a4QOeQqaZYpwrdFzofEQ+gyvP2HALZ9gJ5jZYnyyszc7JKpVHmQtns/yCFz1zvX0JyKfsmcFov
Cw3QdAHJAUB5EEjIOcAmIAl3Pq+5Erh2DBOEPw15eLNMgFDwpPkOPlhSwxuyhPyd6Hv6mp0BbBJn
qhxaWzULTt5uSIlQWmaEkQV3qczn3T2ko3hSAMRdsNzPytmIxU9/B+nLy6Z8uLPXcA8IMFnTnNoJ
yYw8ezX/gDvffi+nenQN+XLxi37SuneZF8jn0TU396i5vHzl7qklaQ+rua78NFSDIxvjOlb8hhhR
NvOfw5TFTGyUJW/EHwS2UedZB5nyjHCUUpyA0Oylab7clpF1GTEvsPCmpDUvAuhrY2RzBS6J9r/4
pB7Du2aldCkeScJyY39fYpxu07Q1rAeJDJa8UYucCgb4Ip9GY5Z7EZQoK3bQtrD4c7PLDjgkFDUj
lGrlbOXFAU5f0ZQkkqA3UhJ2eJQ5CMw4yNAlfr1pT6FU0UeYAX0095vHeW3xPqbmCgQaIu+YUBgA
gHV6W6D8pqMHf6ds1AhxaPowaJIAyc+FTUvn/nXoU/CubaLRLLHfMwT+/oUfuHEvKk+OWiazPw3i
SZR/NnVYFzeRwuZN8jyqnfAJblZPowyYxNKG0EI+FB+VHzIlwDyWOOnl73U7U6ANSceat6zvUnEf
uMUZrPmDEdcwk75NRX0D0mcSDBcvYAO5QYE8ZVGZJMMyqjHCdQot/11LquyqEvRPoKeF4iko2MBZ
OjXzZeAejTrj3QkqYS8DmRywbPbtVKBytIMtPLSJ++U/t9jHU/tHNBbVTEuBKXuf2KXwlJhGsFtq
z/uUhWV2hinXw33Niox3O5+U8RB1AfPB6YFAnwzgXASGSgL9PMqzETUQuUIDsqtAh/V42iiTSMRC
uYqDELvWe7IpRRBehEuAOCoLxe3M7Gxvmgz1az+830NwiD2EZkfoBfnR7QgEfNBIRPIlf4es/IzW
AeH5/r8c6yBKURXFbzEG6DqyjXzV0KcR+yC++0emE0ke3Cx/NM2j9+Q0OtwuCVF+2GsNI/LA1J0i
p2tYat5cSJKusu7sbx3ZWyn6mEzzIitCKgOV1gyShyfl0FAtHS6tKpsGrKN9/Bb6fjqaNXdyA0UT
1PHjEpvIOiHKe1mCbv7mRR6QgNwGqLNK4czQgILhWABoMYm4ft3jeESwOvH5ZbRJdCnbamfI0EHN
NjoxWllXK0dc4KpkN2UXzf2BcGYR3OcTZoV8ORvxoVp7EP+m16KwVZ1Qos46Nl0t8J54IxHUFkvW
myURV8CaTxu8I9HNcMUffEy9clxrFChtFI64jX7On+aZ1vx6j3alWeTDbjEDAFD7wM+jg93stpCh
6CL+DAvpbhSyKjFQq8mDeqIrvZL+esGPI3m3QQ/ZcA/zXnBIQiyZncdjh6HcgalQigjwn/nWoR6n
Y6JwTPF8MaLvG5g39ECjFIvR9/a7X4hA4Q2WdbQr60CMYBuWZYdOmkggwbU/5VpxVDH8zNB3243P
oKHYCKg4KpzAV8folj0NXNXfm8veCKQuUZlU2zh3JnYiY/uhRVIMaq4gmdA4n9nu28rvDoM4lZMi
LpNrUt2JLnCHu7QlhfT1NNwNsXotkWdGFmtVVLssznnpxFQDJYpiKtEHhaJo9VQ+G7kYCy4HPtf9
idhsPesHp82Ag+sYHyY3tQ01Vl5oRwSF0/Ga5a4rduoH+lbHvpAA0ZsM/24VpqhDnP8omOqMA4I/
duqcBcRDl28CmUWeu1xOKNXTF1GaTjDPQ8EvQQ9zvcKu/fRleMhfTAth5E4uJ5R2ce+Y24SA0LMq
nsu0CQS+j1SB4v1xEifKHsoD+pAlOxP+ynhHvScuINqLspsPsNKkR/aNhi1+X/06uulxQHIYLxW4
G9LX+BQY2DUU5ZRXbQfUJH4IiR09g7ZIga2kOCA9iEl1DKR+IYl4wcEYp7Ww75XtGvPKZvRGKKQf
N4nZfl0GDAg0zy/xrIy8N9pmVuRVAAuaqLeMs9Ht6S+oyqyq9M46l5saPvQHSwq1ELUs09qymIFz
HoyyQ02OFYwa+yW+1auw+B6G9xqlCtmJwtHkMCpSeJc97lWf4jyBP4RvYG8MHxZqTvf1uFLlTjGY
87/CbMEELWULlrsQwMmwmXhX71AXIgcJ8WR/PIVej+imdt9AgvrvJHIkvwHjg48qivDHJnyE4IYv
3a7K1Z6JUS50mLikquBZWIXXgVLBziB3AmgLBZAyLPy8mTReR2qfro+N10hqZLTuf8dWSGhxpplk
iqFDha0Tpf6Lhe0aBGtnObNABw9jNswZPSGsuj/5TwhChXwGY5l1jtrHCB4DeOsB2l1wmIVm3O3h
c9Rzg8gjwKDJnIUQY2pkCfmq5aO6KLIyRyieyQS50BLeTd0PDZLTuT23D3A2xND/ErO9ZBsDPxC5
qY1Nn4kgFPbU5k38j8D2j7pkyOpQuJi3aYcCCYGq0bqVqcWUGsv69L8hxuBcmysN16/Pk9vpbpHi
w8zaw8UELMLF8vfz+ZL8ir6nZ5/lVzUAHrdlB4p7SsVk0zBEsC5BB7lCXsDN/eeJa5FcnrFlDHvQ
XNLdHMV3jFvx5hTfArIOtDEcOdTDJux47R3qj9j9PsO7mAoWjx9cSd6aiSH4e4tQEFc0Y2BxyuiC
llEmNed+885jBNQ0jHxlEWKgi5OWUITaloQW0p5mjsyuQ5x0g+HeREdqHoPEY5unDCeDGnVmJKB4
OU2uoinCDlVv3T6SqrpqltHHM4p+v9MvJ/DqdZ6MsNQlRJCU6ldJqrN/+yte8x7jZWpTjgpY8p2f
xVA2+onR03/0mOSWqDhC4d4GD/W1aiDkLRQaTVbrsW2hBJ+l0hs8QReXKsPzp7ipyzmOPAjLo8vY
dQa0qBF5BQmoaxjNdqJQwpLLgyCmvRQ4mVJfX+m3IWnP1S2TnRulMEW39IDJ2AKQmke1h1GUaoda
KmkweywA+Pyh4sIM0M6z2a/1SV00nR7TxZd2AQWde3fZ4MeOXxelC14bW3UM4q8xHzTWZtWAm0/+
od/7qn0zSTj0TrSQ9q/viGWLtHAurMMLlfNhFoAd3Z13vRPZxFVEqzvSdgndhnfQYa62iW9vH22Y
njp1iA2fG4KdRbLT/vlqKgGqaTliDSVLIzkHrUA7mIYx1GBmA8HQ0Oi5cXzGDLDiofOXrO9I7hN8
ncYbwD8SD+Sw10WHzjMUxAJp2fWwznd08vfuj1Bh3lVqGwuDLkd+33z/jDaM2ablUJY5ihrr4ot7
+/EcPIbvIDCwWX+iI47M7kahMvU03YNYkggCHWo4FGkeBF4+j7LMMhtM3Q3xDA5MK2p87J3X1P+R
/djNbR2K3f2OZqGV9OE/gco/VpHhBBX9GhnipAyVwuc6i8bP1oPJRFuxmJ9N4FlTXBnbZ5k4qruZ
m1va0UoXogL1RChHGLeh0nnDumVX3rW1y/8akZdwQ994KfNb5oVhtBCeKHtth6JYMSbky9JMLrTQ
hokuYL9OZ3hI/exZht5+eBcPUuIYEoDIi+/iRAkKzJJiJTMx7tpJa4leEUUdvfJ5Ze7ygg8fG2lM
VytKqzCYpRnxZTIah5uXYqG/vZr2a1qYQQaye7Lbtnxjc65UVU4bIs9DdUHFqTIQ9dpqprYY9xW9
dtQjiOjw39oSDOptWgQS1QGm0ZXDuw1mehOF7brVYddsCbblsED83musNRVQ5SDdrvpveYpIVNnN
CN7q12uODlN1g54fyttHgpw8saXOr5P47Z2mzGJ7V0oXMOQ7MoOAIZrAyZeXnr+A75X3nr7HdIPL
noihY7rKqhrEjiA8vf2Ia65oUGZY9M0Qf68BzM/Be6y+uE/pp4yRVaqBQJBKm1qZYkAJelBnTt52
KV3nztik/MivGw1zkN9Iy6k9eJcdAFJfJvWVG+5V5qeKbbf3tlN1TtvwFtbuPtmWnMVWl7r4ZD6I
X5ohBlTD1Pr8M1kQ2KuC6JOlPW7FRbfU4tk/kvbqUYn3KPxOAFQTjWQaYJujHeMwKvWwiY3e/6lL
UZdEKiXIpeYwsRy8GrLzAT43ZyY7BQ8g5sq/NwZ0pekbXN7TF6XB7twqRuUkelx1E20rZSPKIBEx
jlp+ysVY2jHnETRMaeArZ8LQ5B/hFdJG7RSSuXZ3zExmoMakMnwa6cmZuJuCYRVBrEtsg1ia1Mpi
X2BHytbP2vpKEajFNP12rhrggJetOOOBOtma1Usg2rg7uWLUbg8FNmsJs817uE6U5g6xCLOpqOp9
n2XTeOiD52xwOqdg0fiEoUB/QxkzQf76POh9D0BGyAIUttyAS+8Ic9O3z7KlqOSPStZOsmThu7hM
vDmXnGwJSmE8Go9/tmfX04EIROFPC/2mdSq/GHaPc8uzBvyKvtcfJga4BsgT0hK2SOC2T0DwoQQT
TrMYQiQfnsnZ/OBSuT/1UQPU0HXE7u/kHOzY7evbX+Q4z1V0pR3AkZSCwKGshH+c0ZF5QLwm7whd
12V9/JPstURHuqWJPGAcxDczONpqErNeaGnJH7PrDQTTbT675CWIbBYECkHuhRjOr2Wzr6zVEcJW
te4+uV+8tDvvJ515emLOKYlXpGXmsWahy3TTUk3KMCUgIQ4IfZnAMluQXW6mn0AEFa8Gbd1gsGB+
tqhSmQhwsbsAUK6mW/PjbYnnVJikc/FYUjeZNHt7O1E2FXx+JXdgP67/0bnFgXwMECYztk+8mrMp
ZLUeUvakgKIm0vm2rnmXtD871Yny3NHnJptwe14v3EP6esPcGCVfmI8RPmoffQQLfL+92mTNnRAA
0iDGJKAYfagXrbjfC8nGyVZNoPGtMoqNHH0nnvO0gJZMDCjn1rFPNvM88kybKrlHskOrXCbcdD/g
n9vieHilM/MvbrVXSSYdNFhzupqDTejPLNjmuEgquBl0NWMs14BXwRGZ7nDRfYKpDYel0qZtYh0a
3FBFPariZD55bj39ooAnPhdZiqUGknW2BiHbGf72lTVlWqmCOlwrh+pkRLircYt+bYidoEMjV29i
pKIF5G0goGwWnDGSDor6aQSjhX/3mOReERVdobNoVnLu6zpdyl9VHz9gTzQAKFRbyBPVLEZbs8D0
dltcPjkIoN49L77qwiyMd4NbvRU5TYTrsUkthnxEzgrZtQAY/XT11jKLkBZBayjvzvPOJAT6fziv
bFy2ElBA89lrZiYayOoQrYbair4dSQVrJamOHU9FUFz1YWayab8itlAi583y/BfIpO0vniPiflXr
MsyvPQWLOobuXFQXPfjbp96e4H40DWxokEulXO4JKulGuReddjLe+zMrRjOvNTQ06rkeNgxg/1xF
SJF6g/R/XTfveFBHmajEN5NUCrDrhqJ90TS3O4x1iDVxQy5nDXKHW8PggsUGBl53AEUffYE9LT0V
PtYsb6ahF20KZYfEurq/hKDj/mfQvcqzMehJihiRcMt+SGRgNcgOyKS86ZwfL6af6B+56bte4vUj
Za3XmUWc/TdDDEBfUvmHz4o9XZPxFqQ/8qP/HwXUp+HhOssgJGub1Bl5e3HPrLTU0mcCZn8XJFQw
qvHJMwkM93WC90LLjGnqDlfiAQ25lYSm8q42JktQ2pl1ggRIiuNTIDUnpAzuKeqd79/GHdFU0z6b
gfoQbqx6iBFLL2ah5LE1A0Q+fXfINa0/0+W7zc4PzhNlCkJD/w/nMJRJ9Jd4uP2kqND3WONmgevm
daDieTsIB0k6ciqIBWVfNWRcg6qjoENUGpgRRSDSeuWXjQ6dZtxNMBfKLzBfbskwYmJIUu+t1S/i
7EqgL4Xees2aNOHukl3l+sJJKOGU5ofiaaItsOPs1oiy11FkbACOsk1jiesDXyOkAngXtagl0f8s
KMooqwTahaaU0Sx+0qI1j/q7pwrh9wjPWr2hDHXnJsLogsuu4cOqawlSY/qSsJWLAMsooq8Lg86u
agNlA9oZGYBJvHSwH9PmqJkrb4zbwJiz8YlusCOI19UM0HlNSaeqJNtmu4RX/hTawRB8rYZjEde9
eehdxZXn6nWuBV86+ERlgFWqddq9RfNy4EIB8olZF4NqAL0pI0Z0K/YzcAcnACKWZ6PuoTalpKx0
jafDW5KPx4ZfL1e5BMMhwHPQYTylTNTArjkjkJG5PC0OP9xIxfBOjDgSw0InvU5nhXK1x8OJFDI6
Nv1oifQ83rTGbgO8jZfxVWTyWvU1SRD4GXWL+KLUZel9D0k/7ORTRAKxGmkjf3+QpIrl84k8ezvr
PbeGzw7J2yLiHVABmjCawedeCfq586JBs52j1YHo1Lh95eBa4fGDtWTax8j0n6hk27EhegQX1vRE
kGcQIk/zjQV3GFRFvqGiTLSIVPe+AdsifQOp6W1a2ds72Mtvm6KPvL7o59/r8R92CShZ5uHSnnVc
4Ny7MCAjqHzBUha+9aGFyJftIYMIjKDjjuBUTijqxDo/wywHpAgClIr7D5pBH0QcZMzOgZgfhvmX
4heQiJIC+s3GgUm0OnnSiIFOh+bSNhRSYLDs4h1tAdaA+2h3NildA1hnBpQYC7GygDcd59whfX/3
07eROzxOFQEKoFItPHp9N1z6ueylqczPng8wq3PFaeCvi1Qqsi94OH6FM1iCT3XBmX/1U9q6xJi1
UQEn1pEXrqLUtZp9L6wFM1gfCs9/oiZnv2UF3WVNcMh63eJjBCIPNWPcHycszkb3FBOfkH+QBgTF
Vk/hCuFc3ON7M5lOKfzpUr6c3lBkZQBquQZCZ1V8h+HCCfg8m0l768HRi6CyynHcnP9WNgVFEe71
lCmFaG3uKe8CssdHQXvQiZ0owAdgvjsJ7SF8ajiGUMyWsWYNO8A4wi/WhAuL86XDtF88f+9nNZ0P
/iQrs2P6J7iAj8ajAl3WhZ2xrVjmI873xrStVDxaLJszySrf0VJOCNZp9X8QkyWwO+Absb9DPssf
uQ9Eh5Z0HOxoUFo9ziQl3FgNKazby+qZMPHuwORTKF8N2gcCfom1cI7vGKn5NsJdCxp+UP8oUOn1
EpzNrRVPLvx6ZHt8DMxbexCtrNfG+RacaNGrTtiypzw2d6yHcjDGmhNLayfLRb0e1BfYzSjJKT1F
J+hCVCvhpjTa8pqJfhHbD6wbBgwOPla+fK9bIpmQXv7+erR19IJagEDUA7/CSDSjV4eHYMXjVFYU
yOx9X9g9+3UfyJTcyiuKD624ow4aba6EFqGq34lhhCJ8gpmyInbG2nIYQV862r1rwJNJsR49MenR
9Gc4X1Pq29GNwxKJDCfYDJlFZ2Xoo3zXS5bhd3T9shc6D1biiIfo2Q33/rARykWmeaYmJ1XqpVe0
QXgL3ga697tD8N5aVRIXLaVw5ZIm7tfp7YSMZcmzSUJriH2vvjOVo2VOCZl1UZLBwV/SBZO9NAOw
gQDJ/iZOpzWaBzvSzQ7Xxp8B/OpMFTUg2N5PvEEUeylR5mzZ9q8h1QYGcPfvMdWmQvs1Y7qmg/rn
l3JVe6PYl0TgsFeqjEYfKpXxi2DsYvh5ItxEes4FT97uOvkqKTAFEuyCq8n2kmPb3EL9w7SvaWzn
FHE7ZeuBpRCso3/R993Z1DV9Oh1SRKfUYGQ7qQ/xUHoOMVgryNchOEyAz/1HzRXOQq5ny+kShpBd
ZtIlctoiAacrw/1Xoi2n/1gGauGI9QDTWnPjTYPH94q6J1kk+zOGrub6pyuDV0lzTqOaAWev+XF1
0gInsqKCC+M7Pskvl7csS3oI8iz2b3ujRRsXlCy/1TTA6OshPXZDIzQ+Wcqtb5ExViB/N5M89I0I
Obb0nwA9tobPr1gPVkKYjf4/5luZlywj7XLgS+NQP2FkpYT+EyypKA1MLqMQ6mGy77X2SbuXsqgP
NpIhDjSDIlOl3KBAx+MvhU4Vltc6oK7Je3UnbGEu43HCuigIovZIgPDXPDtw4AGRNHA7CarGrTG3
X82Rg3I3DBIx6JDfbL+WYiq8cnEleuHZxkzWZDa4wNJvP1TfSzqNfXIckVY/yuYm42kkrB18gzjy
g0wbsKi9EUnEqUuPxTy7KxY6+u0MZNVnpVf0Gwjvi75I2z08Ts0wluYEV1QYN15DUL6TaFME/pne
WAF28DRYNLcK/6HjZMxDzwsXEhH1ci0KNBQl49xTbPpj7DcPVkmLcNiOM9F1CkG+cYsk7lFl/V2g
n5qspGenkSdkZnjCohXm8RVj8Ez3vzhm9Hxp47whdXBexXSdxM21w3O01HC8tG9/Hui1LcF0Dca9
4EEnmGYjiPwxZR7pUXuQYfGHa9qbrmIZuLSxhRLBVQvRlq+w6PaN3p5Wizoh29VMtQkCBy7TS9dG
s0E+uReVmTPE1YnI/eZ/3rxXM1+99AZ81ez3HkZ0RjthBUGVa3w3J6Q1QIwmX0GkJYUPOo8Dg133
niF9uHmsYRAMCQD5URWA41BVyKlzalatT3nHp56UAD4iNADNb14xT81CVgaHGVQB7OyG7vME0qC4
Dftw2VotNaxR0SRCY+mpudY8//KK0JEsHhqM+G62bMH22eJloqi9jKfKazpaZIZ9dCw2Uuql8p/Q
zDutGUbvr66sAWVpcdkl2YpQMiOxDR2er6UYPGcYq5i8FNu6soDXOr/0hhfeD4H140/3y304LcWG
z5uBW2fwPYkbCgi8P9ElP/+JqTcP+hKFL5UieQ0GLr1ESAcXyeInaEVUfkSZgk2bg+1zez3BSKqG
U3wgMZlo4+WpHKo23hFGBGPvFqYVd/tTRA4dbzvIJC0waa2RSi3cJltZ3GJsibc2V0Hu+j0jYFS1
nQI214hCBwIpEoB0BDsaUIxYIzCqPXrZDQZlpEu9IxFBB2c4UC5hfrVmnwmr84ZiCAjeOhkMzQqu
M17Qe+E9jsDFp/0iI/fQ1acSUYzXTa0y2vc5yWrE4zmXbCFqnVGBhL055QcC7orS1ywkup/HEncD
gcgXUAOt+paOGvJ9f/jw2iI0+1/m2OSVAfADCyx0+451IzToNHes/71Xttr5kN2SwzitcyIk68Zz
qBlWLNFN9DAZBKEySHkhh/uibWxvxbUbs2FDJgSf7P2BeVLq0DgqRPrZaSMPKA+c3B5sDhqNlT4R
/OyoPptfC0oix7TNzEEqTeobI8Uz8RNA7LQUO4rF8ljb6KRek3Af83tCHcIDCoPdLWUJCONeRHCW
6D6++C3FVkCOzgsiroFtNqgjYhYIvRELZQxnFFER/UIbvjqaZV4sIQ9waCO0y4p7RlwGC7hQBR1l
MCzLjWg3uoAd7TQnJkqEcUYijXIL3RHXxr4yjrPHWrOx7sXUBqS07N7rRus0upsQQ2kgUjGY2861
jWyVKIzLWvdqaLGu85hD2KR1SuNYK/2noIIELnkjHO+9z/nofn/HFFET7qKWghmpMiyr1X9765Dk
alouT/Z2ry7qcT45biC2egLac27RgdlV8qQxrr/Sl4pNNhcdNPKvLlfqi2Ogr+EjscDgl5Tgq1e3
YUv/LmIFw9mDopxkDE/fDVrqpEpbW41jpslEkuV7PXQDAkn4HZvPRaf+6FeJufKqqUlj8sk47FEx
/Msml+X+1jkvcy06wCzKR/Wj9d15rSG6Lv6jVjUgtj7raPjhOdHl7vn4iqIxUb/K4bZ4mRprIQZF
5aVBrFYRwBGoaEmJPBiuFJF4eDexL4PgEkZi1TgKg9PBZ/qTO1cPTpn7X9e3I8+0k39GBNLEn5HL
EMz1mcuEwH/WWOwcXNRsf101VxKpQTNmuMd4yGbqMkqXp5KpTLOMgkvRehDSunGU1UN3XU80Lmbo
/iTTjVP1PEEwUk5/9JIsd74sHnHUDNmahyOMuSWD/iMCP2vfDwfaiI18bd6i5edT0VVpLtSNpNIQ
UKktA4F2+1/CT6eo5NtNh+UbcyLtULixinzT4/I9HNLQJ50AEOZmPXu/tUDRBP8nnob5y5E10e7o
xwjmuDweuvO/U0cSevWj6EzCTC8MHjF0/Ujkow/3Cd8k/bV2TrQoOgtxZvQrZH7Ofd11Swh3uFUj
knVtFYNs7iIWcZiiRjTJ532a8OGsWBKFWR9nh2yWZv0oeLpDy0KQqyHYSmfUBtW/VXNw0HIRXF6m
gz/+u1a3EDgIGiPw46paC+P7I+8KJAD92VZtWYknOk9IiNVQHPkkG6vEAFIf6HHuFt+WIlvmS6od
5hdnWfkKVjPrBuO9zoncz7BE/heTt2qSi3iQzwnlrjYIyAMGWcH66jpXkQHD4pW0i3DS4XQ8MWey
I0a8nuJm8KnIRiU39TmbFOW76qhE4EZd9Z8zY27Gg/gSwQ5hROXE43WnaYxApLUYU+JDGlR2PQi2
c50F16czpz4L5m+GAuavWMLbyDnLn3eUg71cnLflCD+NajgXDgUOfh/YKreAhIg0AyrSdDQlSvyR
zQsKSQ/ehCIyfjTAkjZI1s7iD0J9fYv9CG3IVEVgZtq7qPlkdb6Ao7Ggbbp4PUqbV4k3INaPztuP
rTS0Sg6aQjHiqXmnd3q8g5QE/riJDPqapJktGMTB1RxHCXOewh0Ch2qKfB+OQAUolQ56kis7cY0i
ECLFd+UZPz8aMl6oqga5jbaMzyfJhHZQmR3KcRER5pcpgjcZ6DjqMazLmvSXx3DOnFbpVo+7y7rv
b+haoMvLCZrCKBy+epa9CGuSTFaqrYV8eMmqy261RBCCZp5vr1Vh37S2qvj8NkGFk//SIayj0MbM
3z7IKaMJ1SeSNSBL4BPsIhCu8WH9DY0hPT06xpk5aw0WVlSC4mqLf9K160nZFi1CLJsBXap4KhVb
7kEyopLR4Ju/R4TcjvHXXq9NU76jJcKwypb5W1L7UiKihay8OaBDbKGJUMrp3au3ig7rn3vp74C3
HZbpDix6AC/p2IFPaTrdLHZDWeEVbMUXzlpECZwLz6TtT1DA9drxSfStRlT6dSpdcBHlT45Wg/Cq
avOhgJkLxjjCzzhXZFJ3YWBkJXeKFFALX+I3aJ5bHWG5sGoyWg7oTkDIOy89RSpMI+ZCpwGVsMtF
spR/o8kttpcSFhNlWBTKWCPXzgjIQK1PSDfGCbZ27AqUhaKJhfzPYK6Szk3t7f4usOQ5INQABY3e
vSzJ0qc876Ws9VrhWEVwtecNgepXtENSzp9L8FvW0o+hkOifGLhRI7GpkOrpVULfZ8YvLXuayzUT
9s8vWzrrJ5OvfL0SVGr/pu3paTzexUVYpmmihwWPR6vqivp7Wn/7UvsdTvxCOorFS8NqXSNOqXmW
+S72JiDi6I9DE5Mkpgk9KJe+NoK405ie929DPWB5KD/9nc0RtS1Cav8MB0ucMXCDS045Be+IY+/C
p1dq0KPlk4pb4s6yNbZXjOzZHCfxKtoHG+yvMFAUAwyZWg69TBbmVoWanC2tEWOsCO5FPG41AQl6
4J0GJdCb3gNOXXRYkcmj+TjURRtHRyB/LMq/CglXhYCBv1Vw/9063lF3f1xZtD9DFV2Bv2mFAWtg
S1hPvLeukcwpK7uVhbKn2dHdzYq4XPWgNk+bhyFUjQIPd5gVkQqn54cK8mdQBIw2ZpRA9LTI9+4Y
J+8+E4Ym0VbD1tu4Jn2yT7S5H2xuD8oXsGcO6UkkFgpSEhaAcV4oIkppZWuit+/FKqICkpFb8lkP
InV7jTvBGHdHmH91wk5ZIxbgQx6e1edc69c5XwyNl5WX7MyCQBrS6dGqrh/aXJ8bi3sBzDuo0gMW
K1woZ9ytOIxGaLKDk78eG/BufZKDTd7ntUE55OQuHAB8OePEQMCEmIfbrheyVvpHsbLs5HbxYgax
YabzZ2M5N424ajd0crx1xmVIANj4DhEdMyUdVEP8mUfLtOF7orBIysXVPYqckT6RR3NjtOTC3uie
hhyLPQM2ScGvmtap8HfEt9wn5qJvXnz5ZoBgBVen8RlafHJRkfLlzCu2t/ozikabW7oDtAlacuff
DGQdF2N+i3KKwsRNssT3duqYz4LnjDvQg6TUj0YleTmF+uFhjWo4wMI9+rzvjDPeLj+Wiy43eJld
UbWPjNk2Ak9OFy5iQfn3XNMAwJfmlFPwao4ALz27Fyfh96q5SahpSFV1+/NL+O3aMiFAmK2hs/i0
DDYfexCjap2Ul91jJmN2yduOzKIv5h8iCV3LWjozPjifFli/MqnCJVzxOlVCtmGF026mDAtcyIyX
jgYYOjaADzImVV0zGhdgZ3wWSOCG6F2g19zJ7XugnGmUhSLvAkbLaSkAnKDmE4riKe27Rdnda2vr
8Vgrr+UHl+tN8WRhejgfwq62evrhhpanoYWVv0bfwSg9xqxB1E7ei7szOU2idomRhGnRYYAf5VMU
N+ixR8xqVCi6EiYT1bWW816aI3uOveUsAuEQ2fbZMTEMw/NIKMxml1u09fm26kDs9i2rX3JySHVN
yFIEyKREChJl7gmqtTFu2s0gxLWK8cVg1WYt8EvkUzqtaYKPqFabR9wpUPc0Np+yT9gC/WzNQNIq
cdnCiWlKAKeKaku3U5NaQ/rEy+vb1lzGOsgVWuWh0/mrUSNDKOszgDh2famcyUSyX9fddSOk7ymP
9o9akmZEpmoF5Ya+txs/5iEVf0GZfznpxf/RkOCYk/Cp9e2ic0rarZqEBXLSfb8a2dCiRmf0EAGC
ZFnFKvSArLfT+NOiLNbRLNCc6H/00ClRvsqGUQ7swbvDAZwyAHd6V255VQ1SZwW4ezL22DH8JjHQ
UD/DBprD4Uo/oqNlLLOm5K4VKDxojPJcmRILfl9rFttTPfeMT8ycTt10NysOWIVagkwG6EfHo8Rw
BZ0xZHEfNp3e7HH7D9lw/GqjEznfk0QaLUuXxhpFR1MHJKFQql+3mH4B9BW0ECUHZPKZkDrDyxn1
/Dk/Py1fWlioytWENrkd8WMquz43w1Gd6HEJbVNYzMxMd8QBx+l0bm56HSG6jjHjzZDM9elXpSuV
c3XiHff7ByFSCXklAsx17FkQvAStD0L3/sj8FW8wE4XHGAJ5r2mVFSI68w/iuT08dHqZRmw7X9nm
sWQGFLAVmjxHIVwqA3KF26RE1xa7y6eEp2a17W7k1DuR38m97E0evV3Pfc6PLDlLeVi2YVSx/OuK
+jMc2f75V0EVQRflisG94zd9KSyu/jupS5XiAS3MnMrjWTxb1/X95yytBZZ3SU8WNLK7t/cxZmZm
OEOe4cvuAzFmXf6zSkkqgRMv81Cqe+HSvnSH/Ol8h6W86fDNCG7MGLKhsehC7K6n7wQkWcqm5EJL
PlqzC5ustafeQlsC/zHN+m2THzmH7bQA2Ta3eb0lzNv4S90tq4gFDo0117TIFpiTVrAI9ZwMWHiN
U96QPCX4VJ4acZcOm1XfjuufBqm9CDKkwozpK3uCObQvuiaR92xSVYpPflN/V+xzEpUk79KM0OLV
CgQ5XKGGgRShGIF30dIRNvMAnR2s4eDq0XakJd/ZiBb8paZ6k4cdXBzKgim8861yPjXEx11eudR1
bWcLIJq8SgjS7ms9gYEj2YdCsvdbbnOcya7fDOfgFFhwIUylY94qIjaJnK8caO9Om41x1/6B+KlX
By+1cEF5RqDzE7bIip8yedFTv7CgcOWmnFeyL8oRmgre4Ltw/tGWwF0I+mntyrc1uf4Aeu8lRbMe
7o1vfWVYHlfwDLEHni/vJp37Dd2S9AgdV6vqNebKhDyQf7+pIp4qmZPqnFOP6ai6Mx0GQ1luKXPh
Y5toGdFFzKRv3uPparGnLj7lGqK8GjjZJnHm5u6Ql4Goc6/3fjoZVGgemP292/RGkJHDKBIC+mxR
WH6L4RpVFvaC3bfyzlYPeRxaoIkMmKSBAvluli/uwjU3sUk1IzG9I2mEb7qQ6vofqG1kM4a3etvl
Ncr9wurKDq7t1SrWTNRM7bZm0/ItNEedH/nhdkZM0e3pCdb+3KLF+CTErluz/Ip/bd1kLBgG7paN
PD/Qk/3lhFdHWGPSV3aH+PAQmuyko43tbj3sREIm+a7iVcOlFrnxlUCEGUe2VKxgyMLRkxQwak3D
PIls3E7zplKHNjdgTd6vbdUWKQVmh35H4whwUoOnSHJmzKEJ/9kTfxUAxddsMDXAs0+2i3DIc/I2
Ny1/x8bYfEvY4ibxuXQ50UfLVctdpnwTtn83Xd2ORi+qwOiP/I7AxhQzCWovqgMOmVXgVmal52YY
IBx0MwenWiH4NEjX7nTgNn5YBkLmScXWlPALZuvmv5bkUDksXW3BhFmK1qC7K3QmA/qoUyQU7QZD
Fd9YDL+fCKmSO6GR3ZtaQ3rxtzKMaa298NltMw9qQ57dXPjZk4C7M4qc4X+S2ApmvciWpct2hWCJ
9m/jYQWiPdIbR1zaGPtrbz3yVlpWq5iZRFKYdURhchTptOaUj/ButKgRrpXx/CWViixFcjUDqr9g
A9x21d402dSi17MP+YbBVSVmwTfDKcjt4X5jzfuY0kmNCgUiWVplFYyqGvQ0jRaODQ7tCMnJSXHR
S1uolzykUjOecT9+DolSdHrbGQU6idVv1nZQhZZMEa4mmPqFpIqIIzs/BzVIBT6eKz7k3WT/t7rG
HaUb9v1swZmUdyU70HF2XSHcZc57DAMJDzgJ5vZJkbDbFfxvwWeZ+sgRx3pQaptLyHnYBi+5nmdt
Ut+Uwu6SsCKxJMQgV6TTJp3v09fEU/+i+gvmheIztcBt8mfO3/auIsb3H/1cYnMIG9E/IbCV/tUj
U7hGJPMTZh92uQXcuHPPL9qSQjY9bw2puyaHmEcTmzt4/M+cF0GASX7fufSxnBgyfwCwmesXoIX1
9nJYmjK34hea9Lp1h2BLJpoPHLp21dSdwGjZB6aZXVNElsADANOV81G3H7nUOYcuStvhiBrk2Nxz
nb0ySFCF11vD0R1GjdU3jHfWNmtbIAfkZ2wdEI/cZzSlxu2hCmmWyFCuDiAjpEVX+Q7vkiJTAkUl
2IhgJW32shzxd5s+/z6N+2Wd/XLThe/E7LnnRm3oCGGI8EYwzqv3bRDZv1kxMearOKCinj/xt/V9
S+jvCROYL9NfOq8IzSWFQ+OqYkUK1URstAs1NJzYhvQw16KOKSWaDa7tAlsXERucTrYIfE5K+Iow
opy2EfcA49SDQN0TKZ3FSAoizY2lNNZUVQ/n/xAd/XXiIFMiCDZsdzf6dknh5daCfWfjO5/rdug5
PaaZ8J9RfaEk7bVJnZ4LWrK3Pollh70w6PDXo8hfueTUhUOCo5C1rIaIvBa5KGtPzMh8lIPOO6AV
yGNjO5eujG9zos6IERVczAPBDdugvzSU8nuXGmRJGXX515Pgz2rFXghZ9D0OvKzSbbxd2NL/wKqE
EK0UcOl9yYLFAKm+DVUDTPpqu9/+goS4yP8i6TPRWiqq0/vevg28brPYcSSvX+dLPE7zpQaCU+6c
jWHNsajGN3YOYqqt8w67Hjan3lCtOEjubHMA1Oaezusetu/fXs7wLGv0N6UtJBbSc4JkJK0utRfs
j1aQZ420u3PkE84vJ27x4lB98D770S508oInQMt83he+ct1acCFpMKX7TyNZAXWegbBYOhdLN71h
PanlMmNxZlN1/ok8Ch87QdGqdGAaDCxgE5Fh0cyDCdSSEsyZwuKYIz0lB5LYdPsfCWxA1J8DA3M4
BQ3MSi82V6Ms39UZ7Rj3SzbM9tdAJO4FwmiaF6S3nwbjQvQlygPuBwmLXIqjEBXN3nyKp1MMp7EH
f0U7+T2lvb8phzvr1LMgvqQiVN+SS7ZLe6sct53Ekc2gAbJOOzBjZcfVnpaNPOELeN91JOxixYlF
dCjVcuKC2VaLPSnLaR24wEtMK5pu3Xydgjg5lx6ZvKQsilFSD4IHsEtu8+awQkrdBbjZTH+GKOpf
5lGeuKTyhvQtQA7nvxyp+PacWGmzB1e85VF0aYUWrt+KWNkLK/G89Wj8l+ZzMdjS8iwihZHiG67U
sNW/lyVkGsqT/BudjAXS83tiCDvKnLdXRkDKpt53kI+POEYCjODthQhDnYOpDiAQr9wPrMwh6fwB
Sl0ov6cL6tbm2FyeWqkHhMIQLd/RtlsZM7bIlNyvgcORxZKzy9vMnoiV1mKuJvAiLHxDxLOoCjYl
nIoIFgob3h8PxMsaQVb/4IZX/9eb0pPPW55x5skOoLZJvkR2oyPh2NES9JYFESvN02yXM2q9230r
c9IrlwbdwFtISwA2BP+2ZCdvy1U3GLKu5fWXjH7N8/0d9WLWfByDWDZ6l/LpIA3cVvPypRmClETk
SLklQF7MMOk0RSxYjLPZAElq6v0wvf8zQwKqcy/4LmfUBcLonuM3YOyYzY2yCGXFvT1p7hVEyVTU
WIg8YTAI2LInGKXnDMJ8t5lbDt2DZhMjCzwEd3yogiK/xZ21HAUgNox/NkBczcPaNo5zCTu0oKxN
Y3pAE3KJnKHLRArnR/Tzw5EqlDq3T/UYq0+UcKuY9jorODdi6Ux9gCTjvcEKHnCeTIEn73uL0aZe
9e2NHNAf0Uth+N8lvcE3a/QhequVMhdJMTKYG6+DGFAqNNbgMunLEfCFSUjtYk24Yo2DBmGHOeOM
Dh1jbMrJIqCeqHQNMr7SbvibhiFD2f+IRaAcqM+hfOVmWSKT7y4CIumB4dU3oE4xJgrzrS/T6tWr
dRxpz09A6+r56PNH9h0E4Bsf0TEYNtJWUHhVTSAPquYuRIFTSjz6T1H7BseJqF710wPW+rpnRRBM
JybGgu3VkD4DlUxs28TK4vibmX1GsNBqWrcz4BAvLlmC/T+yShpJAXKNfEIegwX+y3j0Hy6UpqQ9
yvoxYg4iurE8r9qtAZEl293ITdppVSiS3y/HjV9RFQR2eLUi0L0k+C4fX6osjYbS6x3rVrTXdMW1
jLBR1Kf7JVhb0M3NH+MY6Uxa/GSILdRyN/TPr3thnVG6VL7g8qV8Y53AQzIcrZT9gWIsOafNBNth
Px/ga4PKaAqyQ604jPT2QigoAWGNBxUFZrGCD5Ci9fmfwALWmn34g6IpM9DF20u7UkREECeQra/O
IwafETQrJDaz2xNp8qPYbM5PMsOIihXpjVYI5eo1Nwktb6NP0L8P9tDCc0rzcJo6WWczMe3syHWt
jmDjJ3bbmvIFfUdsnAj5llpBcY3xJaxS/fRw2+zY/TLS8OPyPJD9gt5GzgngdcstkyEYr6unVCgJ
nHG39oJm8aupwfJn1nHqOLXalrzQctNJ/ut7iAUtPWBrtCvvpbDSY57r907AE6PsidO+Ke9/BnAb
f++PTs+XpqJnHeitYqLEe2t7qmtWqIHpimVUZ5kVSOCjOH6O208F7e5hRKNLMrl1lHToT5hYHuG4
nNugvXm7zKn7UuEOzwxo9G33VS1F879vRYlBduvLAOIkUN1Ejb0Xf/q7Yk1JEQ3BuzwsDgjRTSAE
Huxxl3Bw++OoajIiex/62acWgoeLLrzM2s0yKgkpK8khwm/tyWJFPbSaWWu8RPpyNXAJlL1pWDNK
LBOVkjHaS4wKV4pQZsEokOtSYe85EX4eCfNcajB47v+YAkznHYv6ZktlJALHo58jRKAlfmGDsZgW
UxbGZFCUXPInP7sNYlhtx3ftZHVtiJcrlCoTcclch/46Xe7QG83ilLNaP+CX2JTar9ez64BS49gT
4tTm8fzy46KFVtmew4VGWOYz3WVy1bodv8tVnv0up84Hxv5cW/EDEK9nBWXKcy68UG+88vsFbw/s
AhRzdWy6rLRAU5ElxCg91a5kHdgOb19CHJkWZAOClULEN9kAI3QKhI32J1NuRkwbnleVoWzeI2ef
Z3JQZ6MXM/kXu3jiYBVuWSkOAXckugFbMvIFtjGX0WlenMAiyBtI8lwCvzRlk1cPlyteRs4uMk+i
dPTA6p1nvkiigkvGjS5rmD2+RLdhMgWXgI5fBFEFjvxCh3C5GCXBiqpCVlqX4HdimPJstG4ep7YG
HYh8xflYtVUdQNzH7hw2Us3JLHOjWU4Tv+EzBnyXPPTKoaVea1vwf/zzzem01UjV+RfhRZaMrPnL
cl717gCzkBtQZvZgCv8SMGNGJJaKdRM3zLkv3o+ZDpYVIhgagHBV0vBlmfRRTDgaqwzevJAxCquP
IuZig4/Nd3XIw2cF8P2+4P9evH9JhxDUPt4xYxaCLxoTxeNIuiQEVJGe7sg8i0PQ4MUm9k5CZLEZ
2YQ+CEHPONjarTa42yONY97oairbxEnioxrLGUKuUWbQA8OAMCgI3e91BbHme+xbG0dwv0y/ZRrk
2xfDP0ssJRd1ICFDAoOfBiFEa7w7uT7x4AnxdsJ5XH9zFVbSQUq4L/gBm5h6277tRVVaGuG/3Tf4
JS3BqNvldDCFREOSBXBVQ5lyrdchTP7rkDpPTBeKNsRJNnokrHXdtkW+EFcQ9roB2gQYYGPIQoQd
e4KAQ+ljERMfXLbtC4IoqiTKTL08y6GG01hAn21pgeXoNH0cXenTBk9ApmTtRKcGshYUhzqPHu3C
dkhcC68RxBxt7YuNnVLc2+zzFTq8jbiwSmTLQuOs7L2alSqLn0sKl9EBNjdRUJoncztKbVaDKxIY
R/qPcoaUI7m7pzOHsUhSClNCGZUOv/bDjWU5rBBQYdIQnLjNIbWZWeYKFbUbyDauQNzAKWO9vuNf
p2E4QRMgzzSJQ4EKiorS9Kt5GbskmLrjuW8uh3fty098MogSYgTGWOOAgK0bNiHjtprOQhyxFO5n
UUicu6l7U5Zot1yyb4tS4adFlhC7lNUJkqViWM784MCoyJByczlQwFHZSfJJRtBjNfFFZNTrVD1C
c6zl2IYEpwOhPfR6raQdOIhA547vcb5sipN3Gc00grBK4JLiV2IhR/WR18d/MUAycwpVehi/q+th
W6dmN7dfCbSweKnzVInOsTR9KjgiVY5ZAjz/e76big5BGpwAnUVUvPtT3SglTVagqjUXyM7zu8QL
0BF589dwCzoRgeDcfgVAAtoTncm2WYmQYRNQYAn/nvd+WwdyUUM/c5DGIbHjiadw0GRfLCtiA6xA
7nduo1Zn3KB6wsExCZBxHi5yNu3m4z4ntZXuISUrwAyo57PC+ZHtNio3H2yInsPpP3xxRCmDy4OZ
GhnRo2lIh2Jr5GdIlObbv/IuixHwj45Fr56AWWfQvJy+S8hH3UXJ922iPUxCQwCmNm9BxD0s5L2B
v/LzeYUHlhuL5od+qyZYWdyvn29C6fF5vI67Omv32Tfm4nNDalMHSWUXfjrMYKT3LAmq+6rmyPCg
p7LHDrCyQSzg5IO59hMwVLt9d4odc8v3F0iVcTK6OPPye2wpMgse3Xmm1kz8lt9CnJATOSKA2R3g
+UUBZ4jSayW/nlucbTpDkTMGPjDS8MsDowkHawy498pvDpI2kjE7UcSi+eG9naD1Pd3WFKyscAgZ
x1YwiREO3vxtBaogUemWPq5sgTUnYcFAWlll7Arlb8R7jZPUyNc0Z/F8eFz+VO9lCTsfyz7Nc8Kk
R51/TWGdLY3A4tgQl2RKU8xQbpwwcElLxMfypkNuSS5yZsK8ffeFYyBn2pAIP1hWhrJkyx3mLnAp
Tjc3u63vhcEDSf03QRrMHFpdNLC9LF1X/03UVMnZ74wldu8H21u6XDNu8fZ/xOCP2vJik3Im1ok7
p2z577scJFUbNFScuhZYBhVWUEZGzGKnAXlbcUUaD9aeNDUoVbdIoQ5JFe1uVZtN7s64hws+s6QW
cemOkjlh+FUJpia9zewdUxrY8fclvK75DnG+za9GfKbxf8ryYYRF2J44mfP/UtEyd94vmJPt3HOo
55EYAkb0XYuZg0YIguZ5DeCSSyd489yFVsXH26gZU86Gs+27CXe6SDKR1sLKq86oJQHnvRd1gFGA
JWJsKNxJHDoc7gunAuGgTv4qfc23ZZr49B5uIaEcrW0UClC4/h9ycHUcaTKoFDt5bzIZwtIF8ZWH
pKftZHQpba61P0K8oz8/BdSVBLDGeUGqRpG1fObA3kEDIbKpD+KAIVOPe3M33VURd9X8YQZoceL3
uoa6br6KgxMufE5JHyPpEvlI4OhOd0/MshZgLYTNSF7NSfcyhy3TZOjVE7EOOwz2DbLewj3H1Fwk
C19TEKavSKh56pcBwMz6euUeX6yPJmcC0uidDZx1DsnIUR3q2GD48n4jxpJx0bVL8JRnIsgmpv+P
ztVigA0lV8WJLjTeRRir55cUTCrdHDOAF+wUicqtxXb9U66CToaMmAbJ8/Jbw6wrnVXL28CxfLfT
KDJIsRUR2xup2MqEBfo6r1TG02rO99NgkD3uE2AzhykRXKOnJNNDp5uRbQdHQ54iqgfp7hHXmV3w
0u/DbcxbtQO/h5HtBgmhArPEytj6dnmf6ZSTrWEuAFTuesQmkcriZaK/6ZbGQCscaPSW9a2hqTGN
C6NMfIpvKxn4ysLnZOmzSepYHFZCE7+IhyMO0jP8bkRWlCGYEg+Yo4VJHRuXqX3dK8+NgfPN5IYS
nVJtgZ+6iDrsKyS2wSWY3Tc/aXOOB2/2WGWHwRI66F6EaqpzwUsyqxX/yzRTI0uvBUpeaTi7Z6kg
kLHH92AjE9Jb4J8IwBagZ0TyBsYJWCpf9uIP0+Q4nX0yhYTbK0cturxajiwUyXOBn1w/+sMO6R6q
Ya1snwSYfBvd3bX3akBc9mlMn9YMakLU6WK4KFAgoshnM+7/FiNROC8WYJg/gJEEo41fekmcx7/Y
rQWeojAPAsRNAaXzQGSWljtDUzzSdQqvYYMBOktOVy7YVND35XNMjD+S6b4/q3YHrlYKiW0TqhGS
awydReBZPKMzL1fwX82b1TodQpJmq7dF2udorlbGGPoNCaUa3gXcXR73xrj/I0HD+1eUVG3xeSVP
RNCkWm+HEDRTjc9xzBiRHlSshm1QhcUTin2qZ0DiOrw92OXfCugYSRkv914ngiqLd7Jf3lczW96c
dfdy/yiwFAMJT+yfvj2GvLOQllYq8HxO+jY8vbhdaIn6UCI2XEgdCLqom0rOXs/dzPk+xDKNO9br
yOlUZkbLXMbAQHhADCrEJzzua7rsRwiYCNqc+rZ3pNK7j/jew/jkNmoYNiEvSG10THNhBngcB5mU
YUwIWh47MLMCowagMDl1HfEnJewGIXyx7rRgEm2nXW1fJZslX8xK6BsuoPIk0JR0TEKXJJ0zVELG
FtvQgMIiD0XHzEL4Yo6GHqUVtqGhukAvmc28pnrz8ZquANX7Y3meq88ElsDsALcyfSmjm73T3Ejc
ryypCYyz+Y5h86HAZOvu+g/3E0iiIickwoMs+CDwq277JeqB+NXzYGQEwRDSQwu1AP7/fuH97DV8
oDm/xJOupZ3Rx5+rCVALPnMBzkTDoH39LM2kHMa4RChwlw33GpRPWLV2wiU3IHcy7Z/ggqtwfCnN
aIHNK6j5ssZgiwTmHq49Cy+6L75yhS5EzfJaa5WJDEQSra8rHkNx7TAIx1vzSZO9sezATAaLUwKe
/hmaMNK6w7+ibW/ccE+phoR5T2GLTeSa9ntUBqGhNyGlLU+6JbvpwXErWJevLi1y07UZ2K10Cz4u
L62p6Kj1F9hoMec3zB9qknWQYf2okfkY7E3K7iWqpiyI3K5yRWUYgab5xwOHmtCgPy94b4JgE+dG
g9yZxovZtZ99OQXsDs9SyOwbSWOI1Gl/DdttIGfwJRnFg+TePADuCKctkkjot+ehql0IdQjLT/N3
UXVoYP0rA4z/7HJ8x2bLxLTRLKuKdZm5xV37PGD6NrohKcVlzQ7Quyv1gk3E4QrvD6aZXaqVWUOE
nt71Q0cnH3f2b57Ok8Y6Alp9M2QUuGGgQiMpiRcPfOfHJHg1VMMipnZ8lrNTJNO+FDvq48kq0KSn
IDEt6PXLq7IGLfpS/Kixy18UMSYtfxV6j8MSNDuD7njYi2yKY7WaIHSTZFaZo1uKrSDCmY5SvFLi
W7lbgP5Sv/uyRDfqxYe89b9eFr92WBYpw/lK/shtyK2Gl1CX+dI2wNFT+4bHwHUywJNvvroa7nD+
SxE89p51zBg+6lk0uf2ovw9a+W2XjN4naIlBch8Iv5NjTPJXjd7K5FLPJBoEJDr/xUM+7aWD0smi
XPBMP/kW9844bHSTbvWr0+2SNUIdaJYd4xa7x/5j4eDBXuINUeR1r4xQqbu0n+LzdzoMf9oIC01g
tcn/zWAhG94EkL2NDP/ENx6elGevCUmz7nfFvBNtgkaE3S7QAyyNtb/d3ScTTXaO3l37/F5G3Nod
CK3aGY4bGoXttfwt/7Uji0jvMmdnzreMuLYtHc+3YCE7W4/zcfxHk7u7/FXuCxSvmbHpyyVxhDtY
tkpA6pHJIgspuCB8M5oGarLHWW6Jrus4u0wJ1wW7OUgvUAs9/tgmi2U4DIogROHmgistCRuhx1az
Jrp/9CbXLB/WC0qaOtP8ZYGGqsAMIKKbZE2M+LwwqgAVcVaHd0FUPOunRm32bMHYDVNIil8ieAmm
sBU3Hjhw7RETeJ7Whv8sXccLt3SBESFOsiRJ6i/b4+Kk59eJnmts8oEt1d//4V9HBbxwJu95Hnaw
kO5Z0yHyTMPxAd2yGQGKSs0ZVMxf8Usu1PaZBGVWucHy3qwCJCC8V/g/AaVPTB2NwnZ8B7LZkbKM
NNyxqMprS7m4B66apy3G66fA2rPp6jM6wPreAEJ0VaYcFm0p1Khdp+sgDnUvIjEEwhoW6aSI5SCj
dNUWH0dA8wVuWF12R9nrkrNCIsd2HkhQAn4ncTsQ6s4DZKxhkbcN009M235ufs2Lxngi/EYC6jNP
SbDaecL/j8y6cqe2ns826Y/7QNuOuKCt70MuIcpTUDyam/IBKku8bZZXEZhVoCfnjB/pRZOxsL9n
AcL0uo9a9M7zKpqh30wBnYRHIsgsfGm6Rbvs46nXtNqRpFwQJjN/Ba/bHIZB5KD1+CXKHERMJIAC
q745voDmIoC3z/8AzwgBPetYD/S2wdkV1fNk1K+7i2E6vKGPpV8v2dVrf0Fcjl1epc327ssqdCx7
30jBnuDJiYXfQmsEryTFdApVM5kgjoGqLSro3Q1v6lJ9vHLvWa3V4n/Hlp17izUXgadofA5+Vxfw
c7meKngTtYK2EkCj0jH6jJ2bbyD4qsv8RzqPvO9kbM99+uccSbZe/w10qadHVmgP3g/IBNhs2Ug3
BefPx2QyBP2sHrrQ7PiFgAuMWeCLVUwhr3MMBW/MApMnYYYR0kGPjZNOs+tFDa2ldcNEccXMVmwp
yzBb1qUE11QhNGcfkPf1gR/N2tAgRwIC+3tvxxhG25mqpcDUj74y9b+t67m/9m1dAyJ7bo6vkYv3
1lUdVELLDqHZG8qKxG8Y6eWXPXVqcoY1qZuuUZ4zae2yPbGkM9x89CqkC2WudS8n8sx1D2cDYtj9
rSeXfCmsU+GpxhDiRzbFaxk80JpVScJbrFVSHm97+/CgVI0CO8VahC4YxIIGqyr1oASiNus8Zwlk
ep9trUY+2YRaa7+OFzS3JRbQM9/1SCM4vxz+Wt9PZBNyrHkJm9ySyUmL/FJswNJPzihr1MqWaybn
0GrH+4WGCnfTtwsLukYb7ZCmy8C9GT66iCcJS/IQ1ZtAuB528GRGUox9Pj5qAB5f8n5asfVzheoy
B/49ffOCfxzguyS7J51YfAbI+OwHSAce0D11FkoOWaOe6941Nmfi1Py9U7IaZMv/XO88u6iyWW9U
AIxGsOKwxLWTN6kAOfaLIlo0MzPh/bqc54YMKAL82j7IA9HOyBrYkIBbeDZDQU1Yxwnwej90wD4P
NJgFWPeLD0D6Z5x6BnWaQBavopQjPgyw2zaQKdrHyJLDWtGG4XPXeEwFrQsu3rFOG+NX/rXOUd/G
gbj1AbMFhHky8104GEAY9qaJtY70yXlasOxFbS4QuoT+McK4U5cQjG0FK5ePFbhfF7piHg23zVyI
c37Psqvq/yxg1Mt+Jq6d8LTkBIc5pDmfH8SFvyP4JvPZFf+HmLu3hpgMbMR4C9e9tirPGJx6N/P7
iLhJLNqdX8HNJgc2ostiZEHGcwY/TWeW7ic9bB1hbOpZd4q+K2FW6UvZwgzdgVed9EQ2YZaVGqcw
gLo+FYrGuxEdEH5NgQS3r3Mu8HFRn0SfJ7boMF7CI31kUkVWLsKdSYyNvM4V0kaEmFnL29onw4om
uDoqg149aJdFifVKtJU2xEyzqMN1rp3BfJh6K3S+mQg9xhxwKo75uI0ZVUQriCuCee9Hns3+nA9x
qQ5zYuBWhOiCylByczinAcv5PqBDr9CEmXu7PhYFAatruh5eCZ8FRbXyKnj36oPnlWoSMBXh2ks3
ygLM0JV+55P2URqo6e7JmKf8vOeepSgbBNkxko5C/r7alcaBT3Z6R38Y8uHmByorN4hMgBnZpwrt
PupWpB5neMi/XpAvz9bN+gL0rYwJkc294gcR8CPo0wOo4CMPZqK1yI6EvKfUIGBkZ2sKRw7G2YCC
yCDz13HW8a8hqCX9m/6BCRNG7MNNcA6DboU1IA+BG99ecP7NBZmh0kMJ/RCMw1lB338bXoJJJkpe
FWpR+nR6AU0SfzNmZfy5Y8XD25AxvuiQyVqdV8WWnABPesHo0xc1uCcPIlWp7OJ/C4QfH6tkhpvF
TPl2sr3kJF1N0UZGnGaFxoj6VG6X7sAMGDl4ASCpIN9ypTBsjjouDgtvzfRnLJ4k7rRbYZseQxut
8RUzALeeEJT0w0dk6xNmoAOT+buadmgra+ksbkbqiO39zGbk+jpCDlQSn9A+JAZeIZmOdp3SOJqs
+j2uEVQfXD8jPy5BMGaGqquYjFNYOQVIQLoUrg4oDHILd/I8DL/x1ZeF54lZF3vGdnmTKU6JFWCJ
Ch1ItSIaF0wpZuO1xxuPdDJTqiZdITH7tTl3jhTA52Uva/xg68UZ87N1otHKddA4CcoYFD7jRDlj
23c6DqPxr0n/mGhg80dog+HxSZQg3qaMrIRa37GTUsG9RnmBQbOUiHLpMpAHMUOeiuvERgmylH1J
aHFey25zSeHudRpzBj+mOx/wK7McjakfjIWQeJx0L55xpOcK5U/WacjB0DZoT2Bav5N6+Rjw0O9J
J0yQSRttjNkZozocXSZ8rNb7PTLYuKqFoF38P5J3ASvnCii5v/WAYF1zz2+eP+23yZ6XtOT1pYSD
IA33mTQrVBoKcfNyWSya1e0SOaWaFiIhcjtDrW8/nubeFxr4Zo6iOCtdEnFA5pnoKV/b82kpcTcx
QKCc0bXRz+U6CanEdY+sBU6a6uOkgKc0/kijF9CD60LMte2Xi/pPgzwiDgBS4wORTN/egMeh2j9K
jEI7uKbDeL1kc9N+i7WlrUyZntHCJC+OnJfzHELIPmU8XEBCGe6EfOs9HM3yBLZGsf5R7bm58Sxu
goP/Y83gW2caFANdItx6tAnAbMFMjPnBXxmuH8m75bKlUHWc+ZlOZXMVbyZvwDPBkB0+eDyC/7oe
eBzyt/EBxBla8vyN4swZhYyf3Z4e4ZobnT5gkxtdUo0BB+c2KNyfXeW2Fpgt1P+AulkEFjqVz/53
XlAkq90fccPtsnu+1becaeOUFYy0I7vKBWBJn0mWdqWVFCAiO7HFEUOpg73Lk+aDNIigOp1b6Pau
caCuXk/yh0GotLvf2xzvQBkkIFd9h97t691mGCY/0V8coWZGdnJJi/5SBKZ2Xgf44BAsLMe9gitg
yA/VwNb6g8pVznIgXAX++FE0iusRxefw7TSSMBa94jY5N6gTP9F1xaBY76d5H/xuIQ0FIXf2UiWk
Zg8HdBAwoaDlNvFxEZ+LUmTo/lENGHmWrXzBweTUi5HoqFWlkMm3aGl/dPAGsUsBBNO3Z7e8Wt69
FgpLIOHuoO+z/i1/cRXJeEFRkYW+lidManrGwIRWfxb4xZ/Am35XN3BJKBasbRhz7T5bvM1tAZJ+
MlGytDKbJiEeUMDKw0gGJeRQapTOZpneGWYlQLo4DKRdsAvj4RvVKDPjz3mXzcFvCsx24Cgm62/8
wzFqUb/BYV7YKyZLH0IAQduMsWP/IcavLKVdnpxChFZGNGse13mxELmW4PUlPp/0adQrjg6o19mR
sTVSHVdFN8Q9tWkt40s11kplPRnmr6oeUAE0QD8vNEezoV8T//+Ai9Pti75su8N88t06XDQRNYbQ
PDvo6so3QsbiJG0GrfQVJu3bvMWzW4Xx1oCutVvcpbGDawSXHfYYsd8rZSeQn0oHFMDgx8HFCNyV
0OVjj5PkUd3bmqAA5z8/hQhgSmeWUYvwSavrRzYDY0fR6dRDiaJdtKwvLiwq4mG2hmetU5T1Fga9
YxJCGFzZI/s4QjMOu/xWQsgqmL2NEYvETEr5WrAw0Ra/nGIn748zjYA91600acU6zG58eefP9izj
CWfScXTEQIQWyimiwlHyyGHwRNaA9GsH8WQAmsjCIN8cLxtoRFXrTP6bcWvt6uwx3FzJVBgN5ERc
47fMNJPxjqyaVxLIrhtJRtoY33sxaUC9yAVl4xYenEnPmT6El2Zr30CEK8RrJDZlzAxC4N8RJZ4y
kLzyviuq2NUw/f2Te0aG1xUNuviQ1X/eKEGF5wjYFQnvtbwEqDH80lu7m/Mf0RVMzLIvjoEuzjD2
1PcQDEXsIQH58AFjM1D8oTzeCFk219JyVGqyLBUyHCbfOBTh0PM7D7enQuvEPrTKy64uOa4nlT8C
pA5zEHX0Dvv1TZ3awm6Ilfwgh8o7er0zY20ulWPmj/aggGUWU9OI2q7QZYP/d+nYKgpmheTacIxa
08j19vlCf0so8c6UhQ9deQVpMpz0rKFZWTRt9Uvwfs+7fIa+yfyf7ZL3NdKn2ZVCNlCjBxrd1cdV
D4qFtTs/A5DprYClRi0tJ/IhqlkxZRsRu9LRO0HMx9Y4gDoiRM1iBClgddyp54b1uaY+k39BZC9r
8FR5V4wvaY1f1KOdZbG0W2LYvX6Dg6ixzSF2ypRNRyormFFBg3I6MwtatF6RAJvZkrWXSTjTik0U
REhJVzuVUGZ/iiv7N4iwmWzrH9k5aYC15tvL2hP2In9h1C5Rh83MdjBfjmxVdfrrW33lp8vlI0Ea
XosAp2bGzN4mUkOCprF1lQJbZSX0Q5UGJyJeVMAsLqOV9vAle6u1+r1oVx/LW7RknMIqKMd4X1Un
VdVLkHGo1HECnOpSo5jjtGs3oJojl3bD+yyII+W1RYc6Yr0fKu918lZFUIiFqGkIkqUe2OAkrQCY
VzU48ymPmn0Hv8FhTJJ77WNiv5Q8pjohhmh1ILKcix1+3n+ibaLAbQtSub+vmZqF3uU5DA7nBy/E
6Mn+AVxwECGywr+A//K0VqszfpNVV1m6A0KHy+hkGigCnrYN0oNheoNe+wb5uAof8DhiHWiTLd7w
/ftPsdBI0tm1VbuB3e8+gKziNlAXif2rLHApIFLICK113R9So6A09S+JzzTp0RN4XSOebBbNng9e
qUbAlx4Iy1K+74wxrp9udrPK7wc72uyQN6qmxKlDZHJpSaXyLUkHNZ8zp1ASJMk0dTBurJ4ZOlbB
zM1JiUfRtkQGLXKOHbAb0TOnrqCvSv1UIRe/C2TxgEaqxO2BNfOe5tUTvIKaHad4zccnXtvG6C8W
BUpFjsfrM2XdHrMBRsy5FSnKl0ElxlOYVojsBysfAM8nSVARDdO2Ar4i0ch52TT7hZnneelQ1Jn9
wEVzl1k8VFBV+08h9Af1ms5BNosy/uH9eJnuNkv8Ps+4YiiueGQYb3R+JXVKpTGVeZ8POlOEP5Co
tdLEMkAeyVSXbIV7c+8PHYQa8hgQdjcnb5LAZdoYu8QH72vh2O8kxRCFolOgyBtywnPKlZlZig3h
DyBOad6mT3Wz6H4bcfyYVImTcMZ2cyq04AxZzsc7UTB+Z2rntboMRJlzYqVX1p3U6VRzK3XcO16u
X28XWh3TE/HK7MiSSyfS1KWhU695W8qqSWD54HNKw6381TzXDLd8X8XtwxhFZ1+vql1nL+4wni5a
UJJfkXvOZ2A2vBhotlBRng4gCzfP5Yst989nZimeAROvcKOObs0jys/+qpoPLW5zTamz4UJvhXDU
GDx8m+fYEOUHRXvytNjNo5c3x+bKJq7tZdlaFGy9qaEZQxY01n03MOcwW1hpHG3KU2nVQFo5N3N+
VkEsxUTUeQ+CprL0ps+A3OI4bab7EitayzeQ27y7Hz4TsjBabjHsxeRppgf7diIdUkSoXAJbmnl0
BusSliHcuH5UWV0xj7+Gj89Tg9f5/oZnXIv9a1g8Btt3+/KDgYNDoPdjOX1h99voT3HkTUd8nQEf
K5ugSKzOSO11a7tol7zFZCM5CwHjMbynSUYtmuITzZ0I+fCZ1EQYTg6aSC23b3vOVlKjqhPPtS+T
toeCb4Sj1HJ+/WxdruD+sAk4fZ1caC7RHBZBaO1O4KfmPV2Otqve8Lyaf/DClo6qvViUmNx7jCGx
Sk9iBYwQu6vxyT6Qkc0XJEXWXqL+MMYQDBBgYgGWvCOoslpmV4Mm/Ct+lrgLsR3gYvzrs/ZueREz
KfK/nKjjH4Fc7GzxVOsv5t3JfrmVqXsT/GybxyCa8NLvYH7BCPqwkgk10H3MDYTJa1LTlIoGbkPm
8lBUr1BV7qFkV1W5quVP/l2AcwOsWXQsszih0T8AVpd+OB7fUgpTUFDe6ZCmLzg0iTj+K8+CuD8a
z+2op7bKd476E1DrDmy391UlLZEicSrTq9FKeiPD0Mp/4G0tnKMk9ZDh/83moCQ1viJ8OvZZSVew
K01roHYPlnjslfjBtXjYmuyESWikdMPngKA5uA8ij3VPnycOsVrZqydn+1VGZTZ+BOPH/dbKzjKv
yzykKefrtDIhmlMWscoyRCWtbuy+q+hq0rDqXBXRH1yFkLNK6Yf1Be3n3VjZh/pZ/iLvleBQode5
haN4UoeLe7sn8nNc7VBhPwbW5slD8Nr2pVfcaFh5WrH4JVvEsDSBXV7ElTdFDx75x0Ue9wEiFO/u
xGM022Mn5pSXHPJ2P3V7LmHMb4VdI6vl8lhbVoLuWxsfgowcabcRkGETHhnagwal2wskhoVSSC1b
lx1Id34ComOS7N6r2APNKOshy+OXeuLDwCEPJbuhBkUPdOuq+lLnMMikyBWQw03ND1puOJF1mu1S
Pb17c7qW6LygUlg3Z8KZg4W5WWG4xIxqWiVDCds4nBZOV7yP+u8b02/WF4rIcJI0SHtAVcSwgFfl
Lo7a+FWu5BpKMYVJicsDHZXtuRMpJ5zh/bscN/Neb5RBCfhq7oNzw52HdK7+4EyB3/V6U8o5jCY4
abZh68tZ4ZGf0b41qZA2h6pPBA2ezrFuh7z6rxY6e5Tph5ZJ6H/gv0wPdUApEtdUncZ5Kw+XPQNl
Tc8mEcpr+8co8m4KcpUoQJ94B62VboWKOQNAHEGMMZ9uusOqrgYngIfW9brTxjwmLrpFKRgdgoMI
ErbPqcolgCgGzMstUYyWufbDvTM0NsFI9AbwPmUN4H3KfOSZVtEBnZqlEMz1WpgDU2cAgqt5PfFA
rcMQkqMBTd59giB1ZgXXCi9ZL7oykIGnz562HX6F4OJ0WfajL3MGkqk9uUQagvyZn5P3JIaMfRDu
+S2YjeDMdYa3+ur5vPP+cXsCgKKaoobXlICryZig2AQoaa6r9nJNoKsh4CZGIC95ijcHEYP1DWBm
vWEJlQVzPedWcnA2rkflIsozAdsp4p5cJvdY35SxKEHhj5bVeLr8nK4crJxlS5FSrdbfPyb80WQ5
gcqWVj39cUZW2rPsKIGr0Bosq2nlqe5rXfIuMUaIv9rnxbEYlntz6vZ7Diq4WT/27hI5v0fiNete
ptFJj1nYFikpEi9+1htyAQid8cSUrcB5fSoNx9Apb8FR+7weo76bU257aULboeDuqU8YCvAi4u8K
r7E2casVKDLOpQb26v7q1foRiM2vlLeelrWKCgn+TkW//6Hu3KOR8CA62pBTb7GbdTbeyEMb0LZ1
7AfV7E2Cp1WdJ41JLbdonu/z8WwVFcRaafXn4xHSGMgVZSDm1w492paOfJLzYMhI6HIZ+cqKYcgo
WoGEDfF8R+Z613CGA7U/uWo43a3QnKO+UYzW4S0dgeeweB/Y6zz60vsM1+gcPLHbAyHFNZTMIpdW
hFy6NPRaq3LIe2L87CJX0Bix8W+eNa1Idi5IRgsEZR45l5QFThnugAlnYSpKPbk86cFkNI1IFWK9
3o0LLbT1rLtloB5SpndW2eREMPdVVpQmS4NMaDZJZrzGcsmhnghKsxRBmIba5qpJcAVh5MPOxOOd
cM37BUG7Wt5jjwavxZNqoSqqL6oKGGT+oAns3PFAxQnZSOSfkh55VpCGO3uxOjF+EgFbQsj6wdV2
ee8u+0YrUs599SmIMb2l1Pg44FjX2f8Vcxa+J+/p8ePX/Sp0vbS5c3YXHhVF79cDuqbw1jWnPjRV
cezZ9Kn8YOwmOfG0g2QgQrzMNCNtOzQif7nKtUXI5zg9mC80TjIVkMnWeQvUzI2bKqv8qt2syevc
ORDYHj/EcZMu67amGoUL+/DgYhZ7mlCf2Mnl25M7YAzdRC0ygio/qb7R8Lo5CvXdwNDJEqwRz+v8
PBHVt8dkG6TYhCtcL3005CQNNlc9SmgvmpDZ5DQT9w3Va6IYzNwx0WJspZB3JoYCOd+FLs8eybeK
+MMs0MPf/MhmCXs6Fdrm8hdaTD3fRfD0oU5koe8AImjjSLpDlhsOU+VfO1INXP0Ik6sbZkD2bHfl
ixxslb+oVRNR6AWlmMefQlpwmnXhYqBjkbPK7jgiwuasKlcRYlR5MwnW1tkDJO6qTUrT6502Dezs
n1lMsfh/BXX9D/irzaqI/Z4c6ER8IgoGUDEUiNKL8PZjmBDPIiR2MtgPmdvkp+Tp+4s5viqPeFQZ
5n/xx/Letn1qoaJBqo4q8YGaNcj+MRUVJjxVf+E000fqJHS7gzz9lCdowOpFZyOLEV5Sz8HtFuQ0
IJuOrU1sCnvBH8EyuNcLrXeTcYxC40ooRheKS4D0fQDJYLdFP8Rff7imc+6w9Jyz0zk4d37Lq39G
Qn1FmJRsqSUlqa0lSoHja/9B3uzdtYh4MWurkGaJBkX92UFvLNnrQC7urDrSYmDdAzeWEilB7TW4
jrw0ZvSROcpxmSxfstg7h3zWO62Tw1RvMsFapgaKro9Z7DVIY5FcKnpyjztfl5KM2WqWI8gJmMqY
6n5d5B84+V/zihL4oDhOR2/t77ms4k0hZ88JWGUFjEinRtTM/+WF0EtipErxiSwCkVwyiHUK8Bmb
I9R8kroJBFIiG2dqqlv/R4lr/mqYt6sSivnnDhdBOKQ1QAv/7JAAFlM3xji7GdiGTxQwO5mSZL7D
lDpK64fiLe02U4oUZrzcSZ7r49E7olIUQPJjDYnVYIhnw2zyEmUwbPwgQiJi2rjPsLHU9/YL3qKl
7tMA6Uy3KXy3GZHfIiF+7g9heKGGwJ3xYK+Tlzuu11BDaHrsyXyxP4lEk6fMIceIAPX3LmFkhVE+
wkDgmwxXgKLL7DL2z0x3gSpul+qXKXiKBy+6oe6zIuTYE1WcDYDsIHfdV43VEvCzCBIA2aMxOPrU
C4OJGFFH2oeNBLcVIIWRRXUei5nfVc3lIFtdf122HR++yZaDWH6jCeyAB+RYEwymMPf3s8kIqin1
JbwkaPid8+GSaTOk7z76wHgltpJrNdupqcoCd2UiG0O85ABRLYrevOUfDvazqJqfIM4vjEevEVts
5rH6no+IxRJ70NPlQEuuVHnRMS/Ac+fniXCdcobZzd7YZzDVLskOxStTPoiWl6cVKtADAaJ1qMu2
fcd2ij8zIv/6RmR0wFXYf2Htnk85R410OOSAHJwPt9rWW6I+mvwev7/TJtX/ZqSZz1uzXkwWpt+1
dEwIphR2vNRZK/njIMHEfKzQtfh0m1SxKRd2aX5k5mGmwt9XbG3eakC5YE3WbU5xPjSnLVvCMrur
ENDgIWdidltIJvMdXS73KOCHmir9xy8W7Mhd/XHhOsgfCldwOtYkFO0jP6jSb2xvYrESIaSw5Qpn
3fQ+CCmklCUp+gEZmj5CduyH71ioXYtWBCrRMOlzLyqYrNQ6NY2aHW18knPV6Cv+29Drb7aPqFJ4
YWiTk8ratYsIwv7kbqfDqLcln6XOf3x2MWFKU1W//z9qahSm2Cja14Vgci/QipY1d3gqFd5+l1gz
fYfpmi+StOzLEoCUGR1mortL4EIMjoSvHTwPBJySIOrKnpymHaIeAt0u83smqD9sXzCLLy6ANPqc
MpTZ/CI8AeCZm1tplkVoju0uToStA7ZdYNJhPOmRxBH/g7Q0LJ5JS26sH1YeO68nwMnFzlomAj30
vmFr4vZOBDCTn0QdhK4nEnbrNCjCFDf9A4ZhMPiZsfJi4DPixfmzElrsKL9uNv4s96atFDQVKq4G
Z7V/sPmr+KzLMRY9ZmsiiNiblgHuexVegCpsCHZTQAJI9yR822kR8tfcDQiFMjupGFRMo/k3O9GM
qM59KE22TdpjEkkCD3p/RIQcWAkizMkr7FJXdWBVb0bfBjWYU7dh0LA9pz2+yd6xJmPt+2BJdNwC
IWoMiS3E4QZdVBdRoU6bi9R8FIiO15sUUmXhaRU2W5D/kQQxPsaNdhihV2AKBObN0oepC5FEootH
r+zljE2kWbrxKu+QlD6Nowe2fbEJvkQWBVAU24EPV9HbRAoPv7RvOaiXGi3Xrakpe9wvtOAmgW71
Q8XSaEbY8DR5U/5vnnaBLYBknHg5VGj0KT4k3vX4FmYm2WU11Oee04bCgLAlJnvGcneHbwNyOk3i
4IBJt58VA1E6XY1n5+9FRRkE/OI531jHMP8AfRRuI7lzGQTgONHJb/8hmNITGbXZPjJ4nTE56V8J
z/irLC9QpBTeqDr0c4WaObLyEqZwaWMcHtkikXa7dyIjEAX4DDbxV7ZnIGJiwrL3ceSO7M8G7PQ2
aqOSibfLQVP7F16Y9AD7VhgogcJUoNykCBHAvGXVzVnyxGppqRMmdGgL/lYThzbmNEwCOzJzmd3F
KeN8ZBdrRaXlVGC9n5vQCcyS1XG0jc2YmAbphUkRXyvHWy0c5UbHmyQs2uPvAVk8+x5/vBYBNa9R
Bo41CB15hHVmimBObdX8T+uQsoRS/068ZmAJ5ABIP5hZwqkzdSnSucGa1WFbpMpnE8ppzaglH4h/
Bpd8BJjgN/f/AqLHWnFqJl3vBLMFnkvmd9uGeQYMsNrD/PG6eYws/WCzWanRj4GyKIth26mQwx1k
6vkuk+L+tXKSAcgypBBQz4g/CUrIZ4yXxsVAInpIvBVxL218kZviryZTiZu1j0X+5Q94G23YYqcV
ZQOX/82trG4sklmjfG5LPRYpYvi2Vhfj2AShRFPEILgS4sUAYI8xgDGBq/KdTKMV4Vr9JoFxo7Qk
tV//6JIRr4nErsCHx5/KrY/fFtf4+k1pMyH1u9iJnHWPf8+dsTGcj6wnNjZAZqoofDJd9RHyk73e
f6LrfpyPPT/f64Jhzmg9/Q9P0YDR2Aa4Oio/fzi5/U9M7f0gQ1URgxjbGNX48OEf8Y20A7Tj6C8h
WJHvSJa54fzqjVY/XAG39rAX5XE82bJrm2citBJ/0P4+tIVQGjx0NuxcTHS9/LGtWx3j4EWVlFHX
z8sIYrSx32Qs78dWekY8X0XyKqJdSTnkvpNzXXp8Le4tL2OeR3SUp6zczso/jyNKlCUBCWZtafO9
53IV0ScaRt3Bh+8IOsLzp5OMBdUSukO87GnrFMKUFPdEE1hfLXdxoVdL4o9MtyV5IFYe5HtaoGxh
y0k80Kak+0FXm7GM5C+Y4cS8ATwZMKlrBzwHq4Kdy1zYEcih2TgvL2lDqA16hbbEbo1MAm4bN+sm
TjQDrOA/0LDlT/2Q+uMldbu15OVDboW325ApNncwHvMBJZXHVWZANb4Qj7LHPr/1EWOndlbKUELB
FN7gnlF0dPzjnVJ7qyJM1cCpDzzCq7J8RkbnANErXNOToNyb4zkkYd8pn2u70JT4FMuYELJ12iaR
dyTsSecJtSXbC7wO0l8IE7kIAKZ6MTZE/uwjLk6B0J/2Y0swJp8EhxHRnGeegxTRhiu1/DbrGdm2
62+2mo8UTvwP/96PC/qtyb5iMyOnhZ8n5MMfV+N+pvyZ1ZJiYaAgvGux76oxg7VIajpmFhITwYEz
k/IZa6HU3JBxdwi2w7eQ4RmV3lurV9DXSUsR/4OEsOE8mlFHAJE/XqXEpQMEwp8ZHBBIvIr6MJfI
AO1ktLaszLTdPougObopSktvfppzZWzwj8SIOPWI7E4ID5o5XFuwNkWnkYtVSHph1k+ogVeYzi5I
5jGq2d71k7Uk7iTmC7IBcDOUWQTcSxvvyhpBPSNm7HeT4TLW0bo4ClVFaAQ1aYdEWK8MKR7rzi6p
cdkNeyvLWqzWwfNSaIWr7R7dnnM7+0sDw9cAA7s9GeBsM95WOoISRc0MX1i0bY1DInP9RDPVCNcm
6eec09gJOi2iLpV+s7afZLlv9X6Njzj2nW97/sYu81urUCIavfQcN2HREn77Bfs2XI3Uix5rNtb7
R6mG5y4nObPwIP0IS0CZ4quzVrl1zjENJsrejPml7qfwNq20o1dSBXKP1sYQ2nVNkAoPpT9wYlET
RjpyNoGiXBYNrBCmecL+A/7Tdxhd78AOrEcGjXTyMeAHQTE8l1sMO1fwczUWFNHL6ZLG3q+3IaRg
9VeVyNn29AiqE+p7X0k6u8+49nIXSeKk6bwGJiXshJHO8cuszFQQMZbgmT15NMYCnOC4Y2zZxUj6
9hykuosiO2IXH+H9DKBfXJbssxI8ESA6Zm0T9HAUvdvF5SpyNALxhQdlRqk3T8t/IBkpAiG8r3xJ
BSi+XCm46JAR5ZdkbnOzoc1vlmTpUMcG0+8A+6S9jDw5FgZeDod/wYCGly4bGX9uFhhbAhtZ2WpP
IOFc8ORBG4q7WufFJ83MVqoamEDxvL4TNDOXnACg+kYogvwp3UFF+H07ewoUbiPrBIcEm2vrAZAv
vw6Fn0cDhlSmbhUZd4LkPaVxRKv/ydxYj3X1SoVlOflMqhbewB2xQseTrTPPZlQ+Vn0TmJ2zhmZd
OhYYPVu1glXpEn+W7MMD+l7xC8KPmPCTAS+g9HPN2t4J1D5CK9HOodyRqOm081l86BuLTpVdBkL3
nxQFg3ltAW3qkLlxHU5E78oLUb5xl2KOdNuzYzWVq11ZBMEklsgA2SBYZzve1iakYKfjAcs1Ac0W
itLX1X9kOR43625+9k2WjosMxlCZK/PPb3rn4eSUdt+SAkag0L5UNfNpc/rWrSFwrNkHilt1B8qX
Q1o+9g91mDmt+u0QFUkqIfXwkFs9u1WEzNQw2XyXgcb5Pf58gQOn83eaBuBnn8paN4QgR69MNY+n
NcNoiUQ+JQz4xwXFukl/ioys45APODt/qz/KBDKZIiWz99U3/44ZauseP6GX6Y2GZ11thBLoa0D5
khJPlZF+fNPDzjPEZkVaUK8z5mtdWzxfcpbJuZ6jHp2ZS8WDYowPBbZuxxQ5qOWOtS+TzbLyPtbr
sI0TZGYKURTFuAS0fegV0MwZlt/qKAl8vELS/+JuieZQKlfyL3NhycXg8pOzg6V5iue3XSDvuYl/
TF9UvKF1vEJlxuAAUqp/N9P6CTXwu3pHVnETQKokF6Cw2yOcFgwN9nAG5WGy0VLfxnvHjuj+FbfW
JXmK7aAMZp9+GCtArZA43Njgq89b5ei8lhXxI8L67GoUVQyqfTH2RKQFQZbZsrOB+9S8BzKq2vve
QMG77HMv4ab7RjBjNiqo57mzVXgJK41GLBwm4tkaKbPrMCJ7UqJL4xVJyiPls9R+LA8y+FtILDFu
Mj/O2KtwF9oB8G4TpIDx7FpStHo4E+0x/jqBGZQF3fpyhKYWEiOAvdmV9OuVn4WHNGWI53f9OVv1
mK0TVsKpCbYXFWTdH/W6SzyjdFKeRDvFMRmDzfFJbg74UkHfAqUW4bny25/9eTuh6EImdOfuQ0R6
kUH2X00JJxFkuDSQmkYfWcX1rGuh92tIdV4TnC/5QscJoCdekQPhy538xXo7mUBJUOsyvWMnHs8c
jM/ECYiVj41SWibMY7OQt7y7X6dG7FDR4laH2ALnVsJKWW1o2P5my5V139DulPQ59QEc6H7KGR0s
OD7dLHZPXXyOAmJKrE5a9zSAj+YwZUMWk5SNbHpPKw0oNEKH1L+1XcgzksBqsDJO8XpVS2uvo2v6
D/08XNY7yqiQNELojTW2b6J3TiABo2gzYR1zoxqgzQt6Wszo234T4Pm3XmdnV1uv5hwasYBdB7iM
1B4Di/J6ybQH2iwcDIb9blT/95zxZ7rTNypBOz83uHFiNJjAmnOWkREXe38yLY+ihiOKkwktzyea
3rPb0gEuO8a1JAzhjeK1XQorfrlCy6dsoxRfE8BEZDuGKN9/8R4m3u9dyHNi9Ezn8mf7zKdntNVp
zqeBvoX+fo7V+NUOKtpBQLoZo2Yf0ltL1B4urgMexvH/1MNSCIh1tUt15IkKEJ1H+wPNrre5hxN9
K6301Q0VHOOHRVRne+dz58817KNaRfBCBhAcZAmlQojqGSQi9iLl9Sg8scbGVCMpb+6/y7oJKFmu
ha5Qbl3hQ1G7zALDDQRozZMLriOoQKnT+DuUsPeEqaHsyflwsYimaD1ETBqJMkPPEVfwcVsJIZKj
Ex3D7OQb9Gr/PGvqrR5XcztBKKuas6pn+daClVY4ICHl4ltC1zK0Dkk7VbyimmVT1jHuPgVuZw2u
LeKp0phmeTm/flrY3oll6ie03zsx+uOlbteCbD7N95Iis7o+7LMh/PHcpApWgRt7scVBYafUTfl2
XhkfqBS7RUlDeyOef9OdterY0gCqINiYeF7fd4n2rdDdBI9jdRlziZHutLaN7TqiPhnlCk1N8eY2
+dPAHxBwdWTbh/eqc/jWXiNAUcNpRO3l1zmYcNpW9JVnqTU+7NYFn4LLN9vqd8bi8ukv/2E8pgcX
mGv5OqOBhhs/6bb0eUV+I2UDirDCGZQcaLEZ4EMkCFWEz5eRzbR7fCXJhqfoTVE/4okUxxf9XzGK
1jbKi64W6+SFWvHCVPYlmJTcIlvhMMsc3QkGc6f5OD7B2DFQ4/wb+ZTNuE6H72uEq9Ia2N9WSaGs
ef7AhQ/X8x0UYq2dSg392YMKMv5JrDFdfv7/GtKPswGvBOyVx2qEwmLfnbo2BE0UgMmZDk3EphKa
euDHusBxhy6vqCTi4QBE+ujqlRBjQU78VljHiJfK9axqqyc7/TGUNx+JTwCVJuAHHTipLXnm98sg
tv+SUU7qiQ+4WoTNhO0J9erlAzsb17F6AUa9rlKuLfrvIJdSVAcJ5OnQ7SWFlsENZ8ZZe7o/0vLc
LurVD4LhdJv5eQ7/FliQpE1x/dwmCwtcsaofLUUl0OHUFWRbbs+2DgdaoUdmbuS3hxtlrAW7+vrh
gHJNSsgYwIKfralDHliyzXtghW6Bjt3EZ8KQ1ftIVf2PvugyqkwrpPKOIdJrBo9xPAkZE489aq1l
YgMdx51/uogMecGQH46hseHgBjfzjlzk5B6d4y2+T3nASnKfBi6eutqrCRbc0k00K7BM2qaWRedU
dhv3uGaovskSr1NF45zexCiawfu1MukJCfVI33P4PVrcbrQUYY+Didiv/+SCHDHBIUz9hwuQ+qBy
vZIX+sDDiZ25Z5gNCziunOWmRSs10rAxttOkgTfx4qrqukCLwGHeN1hXEAhgoU8bO0Z7XrFye5wB
8qt4t8GJ0sgxhNH5hedOBGVQag05o8TjSMbB6Egy6FB06ntmoboQcT5L+fn2E9kLRkZ0T7TahI5x
diuaVPBV4ShmKotVddsWUVedRk+giBWjcVXEQAIfPBt+wu41JczWdcxmxO/gK8/izuTjwl6ygAjt
tIzVebhp/1nRM8lMcEZLOpjBvEVO0sllPTli5qVOZ++6VcHqv9LrMna/MvIGnXG6m/FFBgYjy4Qh
aopTX4SH/79ER/b1axrke2kxF6llPUoZ4bQoNmyukkOe+V3+p+Fd6U7PZAVII6f0U0ZckFhTRz5T
O2SOL8woqYzuxvLoY4FUI+Zhhl3PPYvyCDZPS8uWiOaJjJhB5+q6o0ewYJ4uDhmSOhVOtyOv/X6R
qcfywmMPm9fuyt5Fl01CG/SsW9/Rupndv9eko0NSl+n9ixDJBsVFKy9LtRVb94uxCPOFca11cWhw
59RTrvPd8HAo4oVFr4fdNQPXHM7c9Mz0FVrWV6widfrTo4r2Jr9ZVV4+G7nFN15m32zeyUqp1dz2
+2Ap1CtHwXu/zt2LOot3d8x+RE/2QGVZrD+SO1Wdz9oKS28T2dOqo6i60W71oIruhziAZsZlj/lI
lRUCq6R8K/24l03AFZffVtWUqvs7Sx+hdEDykT9FhbOKsJVaOFLMNzcNYneMqYa8UPCkUnqmrqqE
Otf22Ehg7oIM3nNMYHf8/XS5xgEnrlHvjS9zNa0x8lyaDXNJj5t6vzIASwNNqcX8X984Dl2WiP5M
fCLAfQRW45ZHGZwhz6T7+I+FiQ9HxwTGwFCd99hK2XnROhtQrLrG9zJ6pZEkWT2qyf3nZbaJ8JRf
YeneDY/B6q0iznqz8n1LLPBjaUeJCfB3tPtx5aIg26cgkh9ImllDTrL4bB1n0jJZOW8xZHDDC49O
uBljbFECzGdyXU5tEz84IlbgGQC9wm1huaU5pb6tmAvVSIuioWbCEVuDZZGJrIE55LIj9ivBoSnu
lp5ZL+BJ8VAatL6R1RfVYzfXmvX8F2elMLRXDSc2xlt0OT6xxPh5C0tXHOwYgrZsqPymB1vprrFp
fYQk/VCVPujyREaiqBU3lDMYsD49ffLyuZCCqlY1p2wZYBqz3jyT0jUaIpWBw/RxFpPdynwJwKrU
E153r5ZRcUi3XiETKOW9l16CjBWhOIFwEv/jwPRBK58hQ/LaJz5u9XssVK2nAzwyu/c+hzfLW5Xh
16FGzUB42T7/EWUz+ArLWKEY3hm8LLkgFW0QimG/Eqp8zOJHO1lpIJssjVIrlV71Fc/izQu9/N35
vLxGccmiWJZpFLmOYkvrOBX4wmmNf/DLTCZX5A1DoPhIum/hL0vWdyTVvdD/8pAjgDWI0eKbLb/5
T7ongSHaB5otaRd9UWqpY8CnaRevH1J0MVPqHQLXRiKwSmwsL+MSyAr+VhMpc6s0ede76+8SqOyk
M8J3qmyd//majDmqVtaQQ/cdove4hHkQZzJ1kher3UPj2raZRSOJtRyWm+0KTNX2x7sR+xLaVOqN
tO4VcFD+c9QSonR3IkWSrxWKvaUYnWp1yvlGgwtFUJi41TtlnpUatBJq81gVyOS0qHpRrTlGgAKE
h6RKNkPafbIoTMpD2ugwRGxxD29jo//z0mUfhMeXBx4jpAKoKAi5repcQRJrilvC2ii9WLtpHeF+
XdfptI6u6qQ02UoLlw8GvjYSbBbetoSqBfDTTmScd4p53OPDr3P5AhGwGOzw5Vjd9xAEC5rAFzey
m56GjMS7Cs9gP7MWmQUpogboyJFMzz8tEIrFZMWfP8izyDj4IICmFZ43bcllJjc3ULH5WViZEi7Y
61Rm5ypXowyPNchpat0ghK8rI7NZmqzQgvZ0ks1e9Ij20q4des5JiAUu1hzgpoXNW0Zvij+VzufX
ea1vjcHTGq9RaaT7AKz/tquoPrrwGSuOn28kZT5IuGfMAZIOw8VtQQwtD8wyrTznsk0pUbEm7buh
EYJhpAJ04afOTzdjBVpHv24+PUKa7KMVZ2QQkMYel/Ayq73sNuIkWXO5LqNhYapOqDq/ybvHsT7v
y8THlqPMJ2mBWas5txV0rf/W1dkHJoX75Iu7MAlvbKQfmCmBTFGbmbc4z2PMU5Ft2J3SklJAiuKg
2KpTwAhyiPMEzjugHDevhve+lI/MKzdCuqD25WbxopAkL29Da2ITF9uJ/wKhLfdjrJsnHpn8FLow
yfS1UGAgR13lT2CZbp1tVzRl78uc5xS2L+vHivg7fxE8sBcBWh2Vt/758PQoG+X8va0IY7fKz+vk
nKDjTb/NReNCcDvrjOBSf6/MnfjUkMOidhnfRWbm/aQyQrfE4hUGGBP3X8wL5udrgfysqn5y8u8l
GnB0XCIcBCuZ++HEZC6qE3dsi7RCOxGE1lxgp7qoyK3YZpfCFVFPuhP5IUthiieo5kIRtzE4jhi0
n6kqPw3FT2yCDP7K1216ShUrzwmx2S8EHV0IbMgfHSL/SLrIB7v78fgGZF0ZdmK8K0QTFiijyhnK
M2VlAPQrksBgOsnwyD8M4FJuB57ThrTxQiX3s6ArHS7nt/8xsXIxTFbGrSrN/MmxbMQkJPsHcZBU
ZDI5K5IC+TRKJy5RgvpyiHWykLoiFh001V4v5Tgsh6F8MNLLDPJgSPgiT9tNbOBcOa5TXafD4z6l
OjnCmjJguMOQjoK0GeCdNizDvo0z7Ms0aZwLhDDkGOMgjRn8+88rEjRjMHMH6KMcLfWnYBxgXUI9
qa+8zvTscOLZlPEwrJuDJnkZrszs4+4EDE9rlh/ZVRDwNaoyrhOvjsfejI5sH+607p3rEBXudyjp
5dIJpIHwU4uC51isBfHlRLplwKo46npSHkTft+j4aAu30kz6+cSfA41Me3IfjeOzUmZ6eEhspSCA
pJzBIIo/2EXL51ktqAQJ7VnnYtU8VlkZrMYF6+y2XCtqYdmlpgWt7cg4P49BSs0tXpBeWWip/I4x
VxHpwnIvY/Qsz4Mg1+Roes3ARv+0jjJo+r+K9F9pg7hbximR6VUpxI9Ujmj+OByDQqQAA4aBwTCm
X7KmiPms2Hfrp4XqMQEWBJV/aakBA9nmkV6HF6/kqlS89ZVe46R+3nboUzXfpzNv7NvAawNJ1y2z
FvzCwuUtrtdmZkr5/lKncq5+lCsTQiiisyheu2+mVxXhQyjIRMqkEzTy8XN5m1kkQUJHufY4K3Bq
L4Q49ahH9z9WemSxQgErbdSr1H1DTwlZPfAk6RD/wfY2erFenEabDO8RXVa49MnuHF3l6BtDooh4
ZxSBuMc972R72feC3MI01+132FOnKB6z933YJT5RvptdAj7m7lGTJ3rZ548boWNOmy29GcykXhIL
7rD3C+SC7xsyGiCnYkPQ9B7rdXao38CJSS+Mt4cZyzBKxlcFGnTfqh6xhOYn4bIa/b08rHrH0YtS
JPlzH6SNo1tG7SdR7lQTIgjeUv5/8hYrOpPCcp+fGfgdq+aw2ft7pq2xd6DVaUkjX2/oe+kAqIp3
cnTw4bmCCMToOxGr+89rXnxgf4QgMzHz2OxQcjh0y3v+fpPwCQbRjWws4Hvq1Fm86nZwcL2Y9FDI
EqdfyIQWyC/1omjYyPKSc+8nPlNxOeRxZahsjSue5a4S0lbMbSx7CCFbpf54s61Axe9vZ312TBSG
a1T4DP8g+mIF1ncP9GI7n+Feyguj8Lxc5rm7O/CWULnXukj3hD3SlBSnUuG2c1OpiKel/ZO+v4/d
0JNKrxS5hJO6sUjMhtE88JZdvuMIpwR8/y/gj4C5hbeURlilV7IG5uOwD03LTaHFTyFfrpaBa5pT
V30HD9KuJA7FBgckU+O6+SK/AF6qqfXPKvIwYhreqBLO3n7zIiAlHTIHWZYS1mhWZADas8H4cZxU
fkpwVqhM1N5pV9oEpRHahMDE/4Zkl20k02Ci+KsveAsNRq5r0KPrLpWY45cEXEdMTbs0joqa+Pgx
CIBEUiIdeWU77Ml5SSWg7NU+qC5YlKEy6FJEE2OXCsQPuELCvu3/8nKP8ZeS0QSWzP/MO19pWpOF
NBgacCl8DI08Wf+MLdKPK298Zg+azA+h8YOwpf1yeXw4DTokelFTq6dRPOex7/56oq/lrH/g38Wl
VhlqQywE96Bp+dTXdsQoS6jqncohFCDWCClGLx4UPaKnoe8GU49zIZ8yoFk85YbBoaimHglu0LIj
CIhFPX2XhLLSBnAZcsfYdZWaRCuoeMPsE9i1AQYpSxiev31KY2omY2n+f1Y8LvBwFZfdRtVSFGTe
Z2ks5jKz+v+ZWw6aMKsnuCW5FQVhQS557/uQD6jdlmzKFQp5mfAvK0uAtmlrlmaLLrCna2kPU/5m
qwubzJCVT8pK1GPTBQ7HJ+Ds4O00zHgubrJGJ+3HgYLSATNerPgNQ4oyXhDAcGOV7SVWNziXpL9W
xHod8z5cZVViMojjuB35u5GwBj1KwDLEFz+FE4WXZeUKNH/fd2Gvn7V6+BDtay4Ojns5ccnC1eu4
5X94oBikVs1Rll7nST+LrpSpCvOXKex7htZOcUPnywg+F2E74DigI3Mx3ZPAvr6Lnbg8eZrYlWnK
ZwQ/bcOakcuGgDbL6+n1vmzevMxh8kTf79MU8eM+VGVNv3BLXmbtP3z+pBxg0VkNohqvPabJP6hV
rjZrXZz4nNLyLXIBLIN5T/atmRVvxi6CqLQbS+PbAHqNKBqBAaj1doHQ4OjRUX/I5Nv8He/aZDgQ
jCWNkv3XRtatFO9F0gWnq36Z0uEjHeAHNWiV2b1vR5psT2PpIw2DeCTQApWVmqUbEkP3ZolCGO0E
8qByfN2oqkw9TyrdTbSzML0MY5z3oqtBUC6ej+Ds1cWDBy5hMCb8bZscxbrP/lm8L4/5YoC/v8el
FnyW2+JfwWXEc41nI0duaCzM33vobxzrOJ9kiRLci/k+hfnhtacWnnnjVPOR8G4YGDmsIdPEv07R
kqE5yhnTBIud8U56rWVMcLVURnbozEyceETtlzHuGzPIxlk8um7rb80gS961J7tS5Z8Av80CSxqA
RfPlcsgdPweJE2LC9VyDmbUMChwl3Sy61vFTxU2wsb56GhzRLJ7aJdPPbhSCAiDNbqmQsQV/E30T
fhBR5scQTF9jDJ9eeDEm9XJ1nPriZvKDd7FJ/Et35d5U9GW1/WAcEW/7TjP85ZnelO6JUmeNfzaJ
cuqCtSYlzHpBbLeqb4Z8kF7s2vokqMoX1bN9mDH/ov1x5GrCIBjmF7r+xhyhuPnQizAPCJ5r8Mzj
k6flYUvQFrmMFQ6bZq04bZOrFDq1N9pZIPCiKm1d3DdHsQ+FAMpNg/iJEbm6b8Rtsv6+OVLTrC5J
nQbZ2U8KToy3JBdza+2ql2hEwPlYegxijVzEBuAK0Rf+uns1j6VaUoPDkY5q4w7mlKBDU67TEB1+
t4ckFAG5vmz/OsME2b8i7m9LX26d0JMZOIfFLADWjxVsxnj/82EAITe0H1NsTDYN3vVXkFPWTKnU
Lmv4w++cMJbbgorqKBU1o6QjiKeAFDHZRheVI/acZs0E7oD/fHK5ICmEvp6ZWlc0feMs+GnTO083
/NXyocblODEpix35HfncG4a/Wtr+C2Q/4TGW/CoT7HPD6Kj55/5hyulLIwzx1RdR/24V+W2K3FIP
EASIusyg0VXCRwtfgNWpw9ONdtWrzRgXOKZLn0G+NTEld7pLlLhf28y57kR7z88xVvIB6ySj3SJ4
+sqloymV1wlZen1bx+1fwM8A0w03h+nmcEF/uFmqIXRGgx0ZJmr9mMmbxeXZH+LlChAMJFnFQDWe
8bMiAzBeleApbL9Nx5sllbpEAhWkkyTi3pRWrUyqQZAXZO7zm7aMUd3EMIeKrv1MuCZ7u8Rny2Yk
+jlvrBXw1hUJOOTEHYpcjGk3a5p51WshN0/uMPefjsYHgYLsxmQLVsvYcOced2XM8YUcQA4U4I9G
RZNog13PlaTBFyGt6iGu1zyjH8d1f5F7i+zfL1mH0zyhKcc4NRxrT8LqyL4oBWe71BZivAf/j/Ng
gj0kTAZxr4Cyutjvyt3EdeyVpU0XAl8/7UYhtvSdGcVyOcwlTOlq66Hv302zXQUzzMPtrMW1GnO+
qNdnUTa6/zBUXr4PFjLsUKgMgCfTjij7c7BXEYvZw2fQQjrF0q6lLSi7QnP7aDBZL8rGyHmAz+8c
Db9x7SAxvRHwA27drB82xKF/mOHCuhVs8yUC//1YyM/KY/jL/8Ox8+2QWECJkdrQNG6IQLugsWM/
M3zcusNhqbuTmzWcl/zelAuYSniYzY39vd1CThq3VRXcsdz5ZNGW5s3yqBmobp1k+pS1rWEhVtr7
yPpyOr7kHooP4xg6Kwg6X53BYtdzWVYvJmZRqmBBeugE1orkajqeU2GCzmJCyRfm9mXSVQNUsQ+2
+e+oLQFLEYfhx3lrqR8PHAlvSLPqLpsTbyT/L+zK/BrjmOoyMG263oHZ+Zjl0nx2Z8Dpi9Y+0sio
5cd1bCgCwQSQmPTr1mzdFK1N6anrV6yv1xiZHyHUA1K4t2mFuiNf4JJ9YsGq01f5W5Mtl0d/zdMx
oh4KhcDl6qi02y0gbShSuw4vCaE67v3WRM3gE1iFBj1xRp31IvGVKzDFDgVE+cGQcNF74ECmOv8b
cITbZ6+40xe1YBLIa/2a/Ts9GX+y9cyBxEw2atJsHYb5gbh5R5JQrN/GCA7LI4g2aL6QWkZOenlO
So94keNg8YnH0qilp2J80+FUacMWouUAO3TDAG6LiAQ89UN4lp1nmcx84k0RUelkYewV76/1Ue6V
Di+jhFqtz0jTL2qpTOMEWJwUg4SlL5tqCFXAbdtMOC5P9K1hnSIaZaNvmuumXpStBmqYX52uI3Qx
3jZ6jxAFYOG5LgAIpNSGAP74iaOeaCn9Q7bVct1B548JYGyWMxdlmGMB0f20aT4AMfb0YKV7u0LF
JDinPTzrNJOc/3pxvrfdZ2ekKyJi7aVpKYqsIZ8ZQTGs8wKSPVaCABEofmC6cfbX/yvtj4PkDEn5
EvUsDtQ0bbZmzNN/kmw5IAW8O99Ol+6/6oyT9HsgP2zjD7p0UPf6wqY83r+N55aFeVAUPzEy6G0e
yhSjNXNJFdl8wQ+qIlyTTgsmhhxV3jhee8WW5RiseTpcxRfGg47bmJw9DnILhdjDD2IO/UY2F1Qp
JdDBRgBE1SS1LJOL93dUTFU+rouH92ut2iVWb4FTKFjIpN1oi0QuPlHos49ide2ZZLRHL82rONSM
rbKOEsfAhd0gq8DLhjmTw/PYoCg4HdHubjDCIS0ezrI+FqYGpFGCgaPZwmwaq92gUg4aE71wRnvu
QsVxsSQrggmqrWNQanfeXtEsQ+g7RbvXhLAzBj+/dOtjXdmAaqF2oCvKuyMlBpLt8PMc/Ct48ark
zqcW6U+O9XmFMeGon4hQM/NP8A/ZJLjhqk5O9Za57wZ3L+Gui+5ZTw6danmF4LrEhhDeP8Mq44BB
pGH1YYfeab8WzUo3MpiRITaVAcnjvnan1Ezt4NFiG3pxSOT02nG2Rf+gMpj3PgfdW87fb988+mr4
zpA89gkmAWxFC9jjnbvWZwGxJ6ZM5B6iv8Asw99zwd1qPP6weS90CWaUB57wklZvWA9C+uLypnR/
wNep7hXb5qsU5wBsyH740/jfuYTwQsanBPcawrrE/GZ2c/DPGeEoeCTPB7X33zc95U7kTTMsDTdH
Rkt2Nqt9AU8dc+Mfsxv12/We2H8fohNuTqLXDIgsy/Pzk3iYAcuEUODpjGEIJB1w3UEsBxQLVxp/
2kcBYeJHXTf8Puvj9tYrcw/nu1uK2jYEzOFg5cb3C4yX2AVH7tIWHHz9cumyan9Ihz166AvdWBa5
CrZJkPxfuBdjySNFOi3kF1na4mgzLG6TpyNK/EbFmerpa9sah684zosLu1GTlY0vbp6KeULd7zD8
PNrobhPUAOghO492Tx/7W9wvmYucOMYeTNx9tK5X+6rIg15eGjSMx2gga7pr2gwVAncypyWkd1NW
RIw5mtc+rbOCPguMkYVSXyCXH5x755RgXQz4HdQFHAvjwIviiuxEDTP+PfVpRXn0mSbDgPbZmXaM
DejEYG2SP+A2oWpKUBF31HWoa6lFP50CZ4DltKMYLAZYB5hMuaIkcLhqOcL8mlVpm75eD2BTcGB7
KiSru5b7Izremkvid0kQkC0+c/ZqO9MhGyuDVwkgpemeMTqfhrAReznIYR064Rx43+sctiC+pgb7
Yp1M80a/8encVX9zbMdIQQa2CN3LrBUvPIAwOR6T0O2NDrxGqnOOO9jhHrezN4UR1Ien02D9fwUj
Du+7F6N2zAf20VhgDq5bE1GaLlf/B4qBi2HG67C9tCvTFQ64SQx2YXFbuN4BpcyYQu0nMV85k1hs
Q0R4Jzgi89Q/SivwbBYR2NGt/zV5E2FClQOeZ8ODPVoFOzImVzG+X/VQFD2dk4o5M7+FLjSP21z3
GQOaPsndJSaqigLtAhdKUAzUYL76BC8mWpwM+Cm615HhaLwToUN74SOm4vY28ImDbAaQ/l6sZuDO
yREzfvAR6trEbn/ILHXpnz8gB1d78ycl4nnw0oyEPesuGVM/K+0E5wm6WAHdtmOVXJpIRW2ggT3L
lAWrEqjg+PPNSpi87HJ9EX8w6w80L/GL/Jr1+xgToJTWqxv6lanw9rFlSKL9Kt95oDF91CHA5RN/
xzFzOf/uaO8JnORuPFS6a6rcmr2tUIyW9W9HtZIWosg/MsGuPwf6J8WPCPkviKwc3hgF/473UwQb
llRGllpgOMTy9RIicSArYs3bsj39ea7HGzpFaeboXuE1kb0u5do3yqeTqmhIZk2fa3NIHuJSVQR3
Z3FYPOf1AKAQxETeHlNfRQYwGfBZJydewccUB3aLXPG5YTCVWcq2cZw2b9OAN/6P4br54o9U03Zu
1F3C4le5J8moHL3j6inxWHH6KzoS4Eno65HLjl7boOzUAJ1gRJOeBCMC01yBjyTKa/Uo686VxIVq
KxGGlXGyCi6X8dNiFWpwPDxQHzOFxrdSgF6lIFlmoGD8JH0iXyVfEA+S1hxMAPc8LMkFaOrV5nQ/
v9SJyyJC7V5L2WCO0yIJ4xII2CnBAfKUT8PML2Vw3E7VaLSRk8/aJen+PRHUVg1ABahQ9vIUPiww
DHhkGIoDPXIRRPiM1qltUCm+4CcN871IicQe29uQhS4n0yNvHIYxPLvRwo3ZXNGGufj1XI36N/1c
4WW5VCxYHuuT5rgMtXXdS1EhgBuUzYTFJ/1FAskNYMteEfOyHwUrdSmwkwYFpUgAwyyv6QF9JQoU
w5vbxjdjFkduP0pZ55G0OU043krC8p8Q9hCjaoU1Ao5kx9wtDi5G6VkFplqxoLxDG9AEhHo90Dnr
3k2nUfSXa/99cry81NTwRoyjTz/iTFwY1d5b+oTZZl5JveGDDpsWb6TPJMyWx7ImlzZ2EQ+f0qyi
ghdOSkN9xPE/XXVHwGuj2BMOTtnDAHlE61K9tAigMoMQbpXxQUCSXdy498SGZjsiEQc1u0oIuXum
A5ryk3ILGl5DbzVgJkFsRzRZAm6Q7EyWMmKgi1QNf/P/lA0isuqXJUiP111mJIm644c9bBU6JlR7
btWlCG3Xnj9arJ98LseepCfBk1yBNqhs+4y+S1+tq67uYR2yAkHDsIqOXwmAye8yolsoHz5ycpir
Au9+4pHIq6lW+9NcWJnaovcG8W4ebQSg14y0gKbWhW+Snlv90FIQ7H8KACEBc5h8sF+UNXBaOwez
CIiXkcy1OJguFBjyeEP++yWNX6Dxg1o5EoBY+tkxizQ9yM5AVeIIJD8ASbXxbO1/OHVXilsAngan
noEi9uH4N1kpTPnMDEaTUen64vrKC+3SvKB/rcNvHdL9bkdkPUGCCVgQf/sMhkVgoerSbHoaYdal
IrJBb87HeKoG6j+iZQF27YEunR9RXOMzwACLfkuEfRyeqGhjOR+dvYXWtFS31sNPjN59l2pW7sQj
+3HsgXG/U+OVWFaUnbfPZ3fUy/mUZGOxlSRaEfa95+ZmXs0QySnRrV+AROIZSroGmSYAluKiLdj9
oJqnaWaStJkKfDBsElOiljGLopnYY9WkKyCOFaJqWlMETNLz7xIRAQwSfqG/UKslLIUDCecvjFf1
qg5vMU5FiPqW8S9GKtpjf64stWx47VCcZa9jjORL5Jl5eFEK4gu7NlX45zKnq5JtWdhnxMvjUxHq
BiLiu3p5I1EKfmMKJ/7zKcN6jba3Oo/hVP8Y6yg7k5GBEDqzfxvwouahQeHMILNnW+QlNj0acvjm
b2yDXNvOPya4LDz5NgONN/j+2K6vvnrRGvUZFzRZR2/ExiE0k/ZSRKlCt376uqt410AQruiV4/qA
Y6gzWSs7/oMEtsgfXaj48G8Ex0H+YxbJnB6Imeu3lBvOxwvdETyzeMukrdF3l65UOmd63nneHdFf
ewHYDc4GNjNZj2rtaDaMf/ldIdAc2KUL4TQws88M1k5qj18u+icPsupTDmE+qyp/SCT+zqRcrEDN
f7fxzW2DZw3yg69wdhfN5PhSlP0bNrMyCF5QcKl1ExcxqJ9FBZOfkqdRLqJCqcbJqItdalvh1p6C
EZhYaiFJIymXzPMRTHB5rjua8W2LW/L+6CJSHl9YtfRmmwmt+Ufl7hQ3JWRtcW7sO0IZfBXGwlmX
f4t1aZp/q/2JEX1a9JfL759ieYt9k4asfmOYXUHIUBXyLvnLSHqzc/8Tb9n85coL4JI7I6nZotRu
uijCGCz40RGLlxqsTX7bBsknc/k99XX4wxkYnAdPWiI1YBq50CptMACSJ3Dkcq4xBYUx/+E0/poT
2MKjKvKhCo3WkKL1P9t56e98pY7QPdMtEzcGz6B9+SjB7SHKtkPU2tgDQMc4z4axSr/XL/JsA0J0
EZs+CoR2MM8uNqc6y91Gr/82+sG7QEmKCN5UMUXaqRhSMdnKxAmyKjRl/H99CzbHczN883CTnRPI
5ZklvKsRY1nG3+jrEI9MB0gujhEocR4Z1HHwPyIM7DwWM57Zqo5/kx5zVRhhiuIY413CKDuqcz1M
guh9azaoow4z4aSrLIZ0IJuicJfnjkEN0ACH6niHftHNQhyq7jtjKUh6p1xeudkiu9l11/sfCRqv
fEVkMMSMLL5QRUAKg3SfoICXcy+FvNJylr4gEo7+m1vNutmQzGhvzIk5mg0WJv2+ZeTshaBrC16T
/bkXXgi1oMAVCEwV7kR1pEiKBQYm11Pn06bHjgWr3m9PYOJZCQawgXuIfdQ/wySvMRNGViyaqzQ8
OJYaoIk9iYhWfnM56KwQzUBSMffAIQBS77D1tyurMOdxKOvKeAjVo4H4xFMVC6pCJwCq4NrbT1g/
7GZbvgjYgSqtZmPKTYcTqEtN343yP5GtKIL31ux+NsOgqkTRDJI3hNcveZr36euEw4YpyW7NORbD
5LLaxnToR89cyp3qzMwU1bEULlw4KeWl09PHmnVQsl7y2Y5u8IkuTiOCaxwJskaFUYKQijMZIB9C
YvgU9rgtkj7Gffk0C50qjuj8UefbdJqy3fOs5EVpkgfDLfbpCnRzTr/PUD8s5akgr3vYW4LV8gy0
CxYf1lU+ex7G9rzGKX+eE/omBTgXW7/L6e/mswambmweqGR4mnqGnfxj4gQDZTFo18OyoaqGH1K1
CMnN5H/8uRI9DNO5Tl52+E8TaMmCG0GspxclU6tBPAAj/6odvzWrMmJs8QmVkM6DNhMZ1gsj5gtt
ef/160J9/9wAEsdLjwTC8ke07mwqNnhAd6ghjLbwsp3Gh9t8dqPV6SLFq38xGUcAh1vX0n5z4DKI
jvgnl2znXaA2UGsvr2i1BcLYDSDxWNXA9eVzzXsf/BeRFashJefAq/ms1EE2NAh08W+4CRbe9cV+
CCg5EMZFwN6jnac1m/r2QGXphuAoNVUSPf+77oM80VPkqVhdSOJNirbjh5oD7cIGY2p4rqtVeQHR
myfrk4Bq9PoVl1xHgAeeFS6DkW4IVuAXCm6PbmL7TzXdhOh2OsWTnwYZH0dszcmKCQPBIdc90qe9
XRhnkjbfgqimkcQ5Gh+E9ZFvZYN1pfvPTixt2hT/CgQ2a5ll+KpdV0YDwE1oVbz7P19vBEU80hLD
ONGJFQ5dsHlpaAlAXiH6JV5Pnh5bqgfnEzyOfNGTX4cek+eIo547OAC3AUaAvqmCcBvky2ZcNfmP
0Q3DEQUOyk585kywmrWY5s8hLQK/bGnz/IZOd+Ed7VPrruDxxMX+8Cos8ZyttRt9qSJaEcSrgQWC
ZhGA87wQMrn+MvbLQnljiauRvojaiPJBcRYz/N4UxOWnMHm5o+zQkbQS+1XIAxnvXsPSB+aS7EQ4
Smjs+Ae18sEKpYs6SNbFLZePR0qSFqrIfXOsgpQDT+yiyLU1MUViFuvfhJPRSeLJW1qMk0LvBF9h
Dab/njSNvq7S9O+Ez7T1GRXm4kKGha6M5qsCu8B3m+1f7/Cc/UhgyiZeepfxLWuCWvqFB9CCoh5r
7Ob3TuKpBAgJtzmwdFaLauHEilYKAqAEDbGPChTYPCdmA0bHMh9xzw+oDkiX5LdWa+hQocdXsf+l
b2UOPnHjOhfmV6Ud70QSRX2Ji3nL24b1srf30jnBhlG74HLQEwONGwbtPNStvBKDGN9f5MLCtWc/
uhW/QRRNc0XnONLVlhMSpnIq+RkLRjCWOgWzdjqX1/MiCAAsU0itPuR2c9yraXmAAyUNiflNVGhh
7TJzFoNA9XHkYce7wVr9EM5kVmaFSeT6rEuT68I3w1yj5PQfg1WbSM/e7dXS4oPqUPbAERoB57vd
5RopF6vGVWSk+ioncYyYrYdrcG4rtbsFk48qwrqO8kxNgeZjfuqXI88Qwk7JIOwv3HXh/IO5qVKV
bovF+3e/8w9ehK0BWczoSIcm3KA9XOCCopBig8dAWSVs/yikWtWsincbKgacxUJUeYo/1/x1nvQv
g2ka9x4ZkmKMf6HVw7fwcoIA6BS4JrIxXqPjAW1V0Z6Ut/vIpbV320Qsh32iVSb6teGWtdMwBAl4
HM8JlnFufgNlPs1e1o+HM38mAk3LK04/erkIhU3U1f3BOvFmaGHFzCbFM7KeInWhTji4q4ozrfmx
VIEBoYeg8lTyU2oZ+YVzfJNxrB0HgO5jP1MRBKs4w3Rgm5IGDepUhWsjOjCNKw03/3MrFmoGVI2R
HOrZ0OrlxSd/RJom/c1TPgBRSzyCsvDGqp52CDdWz38dbLczFSEAtco00fXYG8DiNzYi4dUpWpT2
Wjy3ULhNQHGUvAAqUVChduqkvCmgzXvQ1KEEWdpZYQVl+NJ9jxJGzP8wLY9a6g3eXYChDWYekSjP
zjQ5Dydtxq1w19qtbKFJnVt1gLNB/G15GtkJk2+cIKZWQSeiMoWxRDJ/4am1Mhg+JIU5vo4dJ7IW
Lon2dMPYYHFSJfJIYiPI88Ftntg2EsCTgnv/anrDRnvYXwRdyuos32f+nH+j5MV17WbeYk8XTmNn
rVsQJ/OSst5FTeAZU39lpYmjr5l//JyKWUUY/L4wv8M+O8DXbptFk/6jWqucQkP1rzRonrlWbhhg
pDAySOqr65eIr/vaC30IqWRLMsJBJGd3EPK07EIi0mnR59RTzSVYgFiYuUxyXKlPRD7v651Qqthm
Cs/jk14PKJRlLajYdBcJ4DrGDfrKCkiUbFkPVEarVJ29mq5m13exP3GF2Ur8cTO9kzs00eU9NAVC
dFtZVtrbacWoq/qwBTPIkMG465yoyLDQrHUjEOXGj+N8LxDgBwUSRZbbcw/UmpRJckSj3Du5+Epn
KUNxZWgo05Y2E057kMe/UVbn8pxv1LurVA0gzjRLQVY9229ag8E6fGgnOv/8Z5AcNSQmL0fSBgYV
qL2T8CBgmgPtEIfgEABR9nOfzU3nMaE+V683y6m5SM/qp0krIhe/5fUt0/FIBxw1fpWuxp4EWaGT
krNAEGtBPgKWE65rq89oXMFwVxDU1F8fCfPhJC5gi9mLuuJ6226MMP1YbyMStu+v+XOIDX6J5n6+
auIp1GUm82zBv8egY6p9kE+Xo+RLRWXOjN+FP6SRVkEePB/osm7Fg3Q7Mu0LEtY7vt9tcXuCr+uo
X14rIZo+2PZMLw0qnqLu2QQlwX3xpDW4BMd5bC/TTmpTQUm/lQsmneTjThevya4jMYvZQOrrx8zW
6AZp8lBUi0Xsmuqo/GcwrgHtSlKdFiktlaBPWC+aAbTmWr+8kBJODz8HYV4c5qsvxSABVF6liJWe
G/QsWSC91kStVcVjoZ+oIDGjqgFgHMxmgM8JQQPaxLGh5wRZ5lMtP9JvesbOaJJtgEq7T0teR11K
2Bp8KTk7kJO1d1obG98H6f+y9E5xpFmUQE1/uqWnq/yjdQp4cUZFD3JhMXq4YWXiu/XTuQzfcFl9
gVn8FzubgCDqCcj1XBctRpbe69j8LVJxb4uQuw+R76bd6dTIyDFR2gzxS7ptTiQHqUcakchSdBw7
eFzmgP67C4howUe0jWZWMvYBGOX8Y6dAn3NjqoXNo/gIDtPYvv6+GqSuLo236vGWOU3vjU1HUmX5
WXDeIC2XZgfuPg92eWSl/EmaqXeBEwr6iFlR+Dyzc6PMcTmX0O2PVjRnuv+HWs8WtSd9Btee2wPp
36Aa7+Sq7Jgwl7X4NQq1JijCv5cCrwlxaN3I5tSpuRMOYrGo/GvbQzNN0LtmHiXQnQRXEdSxuNms
FfJDP6/1Qd9CYQvV3vjrYL1T6PfdLDPZv7KCptZVKElRmRx/+CpNhydXDF77+PhGWPBDmyHjbBla
fr7tHsyBDlQqCPx4tiDpREQVrrh3AJatC/H9gXjXCjbR4QacrgHPHuMEXgeTndWmGrQYzRuUjuWi
qJEsUIK9oNfJFedA/8xaj1MeA3LnapHFDStQ6NAKtvJDuS1jKSjDYM+J1sQt/uW8igIHRIPz4c7d
ZyIDRCHhw+fERdIcygoMFPD+g2mdLi/6RJni4kKBvpnzj8DirMbIThS+ZnAIrenxkpLugGiWTKO5
MidiuLw+PttnsOMd9USw2hleXO2GteI9OIf1a7JvK2NIseVBRX2aVZ+pMxyj/i5CHSDLkNYHpKWq
nHzuh0KC1/9ev7ZtEACPk6P0bUEQtKCA43r/UIKmsp2XY3E7BLwto/wZNTNkfRhEaMp8e5LPk0gP
LPczZvxe0cbRm+ST+tEz55FQu6T2D0d9XR7dkHrHH2xJ0mC352GdIr6/P96FrnvegMmguBJmnhAp
903OuniTfvrnXOvGJHBK4JyvYMRg2N9pz7uc7JNZSl6TMS7wdY+Iw9i/sdH7liINAtwzTw+FLvXs
PFGafnOVlbNEmLKkO7xR0B8VZCYmwpSCwjpxNXWFRnnfgJoikW1R2EBgtozCSq03/pZHki0v75xZ
ewhzk3C2LM2Mt3sMl4RFU6uTkTpnmNpei7GUioAOBV2DrBG7TrfnPJh2JbjnK0NEZ5BM1ukZz3Z3
Hl32Y9nV1OsQEhfcY23lhT209SEFDfHZ/gvfwS9eaNS+BvhV41gtr5CADca+kpYz7Zl0wVF16v8+
xBNmoEDbDAVyU+MNKxz9N7dmLQZQfhkEEfcwYXMo7KEASfRqLS7S4X0qzR/jV80637FTw5m5QZN5
CiEizxGQqfZJp1RJjo30vSu9B0M9LBMg5vSqmWNu9R8U71WDOPpqQUe5NVCqyUhkBJH4p8rPG/Z0
NEcZJS5jFNSwjxURmH4IO9XpUhnV5Z0+2yj/kYpl2/BXsDsOsH3QKXyBmzQwubFJvaHA31CbFQVG
WpxKbvk9eb3Q/Gehvg5btU8N8Zw+F8CwoJhmcjAr2Bhvl3D1AmevsRT3V0FID38xLB1W7gRO2fxD
3QdmdD+gQhE1brDXNh6aQ5ziB8qgQc7MsGjYJ/PFzQrnvHUdUwSz0R+H9uZ84e8EQ0iqs8oIhHqc
31F0qk29gD99DLXggfqQXTKCqpBqdQqm/mxPNdkEYQdKloQrQ/xNPzGPjjSaQF/PRFhlyQIw6li3
5OWCa9qTLDCNclDzsrrwiK3hzoARTWxHSMyObjMSPsJKgvP2iFGNZtnwN3U5q59MgPkTtVhStsM4
7ytkbXCm7QjuO5I09OcuYIkcK40Sdg5FfFVMzpqJfMWp27Tye2ci+u0fipLWKoueSIWOMpIm6Sk7
176fyzlWXEmnC2iFj4ojKEPD6e/6BxFrBjYepdmiWdbeYhREAa/3oJPXZ1BQosxmfpokB1dT7oUT
Xz4U1gpdw1YRF75hQrnC4F5m2gSJS8GQEzSq2LdDGl9ihFeKC6WAa1Xkd41LXclROXx6/GUuZCKU
WE48+TEnT7KXdMouJexXs5xo6nUMig1eP04JC2ykp5XilK9isV3YCDnOPapkfbdY4S/hQURd+Kd9
amJ9FJ7lZGm16K6Ev04VyjnCPLwD244iUXDDgU04HIz26R1cXQ3kSiwkTRvelj/Xd+/KRpZ0yWEx
H7LJzlU1/OGc3oNvps/z2r511x8jGxxn7nfUgbPXdW9czXlcte1HJYDlA+3wKedxhpPotwcNWVe7
AsR0ziXLMWKRj9rs7Z5gzXuS0Jo3lM7yD8+RNyyVEx80OhY8iDEfS3AwdhPR+0OnsJugcWCUnSt7
8lBHgcoNUc4h+C5I6Y6Hk0dxLuyi55Vt10PWaqkzyVyu8w+qz8sXwJZYEdQKx+PCJZDJu3RcOIzZ
FtCAqf89lXw/XxEO6qC9T0gQlDFOikMQIh8wcXSR6pQTBJ6DgpfplQx03q9boMxATksYAE/fFg2L
vL1ZXVt8Ha4Zp2227sRpxGPOQi2wpAU9DymoNrngYGctcKYxJrmwJjIU0oCigAXzpyHFa3GuqZMR
QpWcgODtTdDhZPulTTtDirB6O+dT6Um3F4CsRW6ZZhe2Vn0SMHtIwSeQZtiAb1aendBW+bVBbvXu
lP8XVexL88hPSYaV2uO+xtSPYL6NO5frk25jXuAAIGcyP0xWmZW2CP6OWR0/fR4U8J+nNNUfxX/H
klCHLwPwRa8x+racoG50rttLSwW0PgaihB60Q13fikEXkS6Sa6UGPHm7L6/x9ySmy2zPk3EW6uYE
ktQVQ3KUcYvkvOx7fnfnfcmG7n/RSG7KPC0OfOOBx/cVDpsp+dilJMttonRFY1jMYuKYctCHHKUk
BgIjLEmi8jtGFG9qPAcYTh6hdjWdljwveTwQ3KWZ0mXoexyrdfk5LkF7Zffa31hl0PddrrRczOgM
N7fvnjRWvgkJvGzaA3nfwMATh7Bx0ltlvGcl6W7ZhHIrAbhwfreAUIdc2IIktb4gaD1MzyFU5Kxs
ryQy++txN25dC5d+HjdnNFIB2WvssXhk78oYRYDFyXBqok0rt+z2q6CCqAL/sdiWANYyO/A/O6FG
u2oLqTQFKLcYE6jAC1k+/7ZQYKVnfZNs3xoE8CqPcbeQ5jjsm/vOcfFCViQ4HCMTZDYH1L5t1Xnr
W10oBjYIz9sa9pVTbTnu+hqdl5c2URd2zqDJUkLZM06Zl8ld4uujxnjUimE+3RreOz4ROtCaGhNu
1X83SK8eg9SLGae+eiLQUOTT3QpMEQw5oPf1HUThxeT+GH7Rsui1jpzbz49CJSDImUE0AXFKwHJd
sofNhYd9jyD+BzoPbn0CChHnPyT84dyhkx6cUE53okJTT0QH1cX/ng3hwWmyp2D6602RpqfDkDez
u75dKwiBR2n8iJROtyqTarjqKNShjJd68q+iZ3xAeqFUAzM6KsV1WtSk87iaP9d9GdIJAxoPBaii
5tRwruzjcV5yqGitPglkrAGphLwobeyj4lIs7ZailC9K2HzRJo0m5cz2Y3YaCGeFU6vEhOiXxqAl
rqVVsvR4/0vnAnig7LszfBwbaQQOtFA4oRqQdVspTWsquTXHa6AL7afSx8cMYn49mv6wF7UHCXpY
0W5aqMO06eBjZw2BXS1cikHvV7MrqfvKIiJcwjs6kvJfuZVM8y1zakuyhQRORD6b7qJ/1VUdi8QX
aKsv9bto5G0NQyG2Q6pAkjn1Az/kLj/LYuITSUwxOJe/x4IOGriKKS7DLUG8AU32CjxSxwMK1t/X
63cvQaBJyoRM3t3/5wzhaXGg2AmRmLTbMFx6pw9/O3tvNPJYXRwYzMjMrGMSUAmbMoe26oKkfmRR
yvMfTaHBAwaikPmfGgq/2HRo7m/VEGVmLkBdjxFzvLxS4ByuUCbCmYUoqJHmK0OzFfRNasC9Dvm2
LbHYBy1lFXn3kaU1H0OLCxeiTW68le6t5nsuT96cOT525WCV+4al7TSnCpffi0dbfcm4+YQK56ib
9P63JWnpC/x5GovsJtWDw9NtTIkDwfT/nGfjxAXV3yZAdJ+tajOE3wUMg7FQ94lzENwkxW+aGwqO
qVvyld973IplK+u2IH4/u/izsHvhrJzCKoxkCzvaARfXA8/uKyG5H9Y1PR8THMeIeI2pL+vr/WGi
C9afwYM3xhjGGZVrcT1LhHPbGCwtmapefA9nSWLClooO1LI4OJUXfZg5+P8tC49y9Dx4bgLYwRJT
9abWsGhyq++oy8nyyZ4gtTC068j18UAqDNC0axr2Ea+Sb2VSmwhAxuPzIeaX7Ymmx/epVukpXulR
NTRsBilCCfedp7fM17MbvHNqAmGV61ewmXpL4waL0pjTscdowDEqQzG44qdEepNGwZKu5kCCvlae
jFtUQ8K2ac0P6jydWY9qcgD+SiyDlEliCWca/bj4xGa5kwfZ1JjqLvC9TocCgrVrBnQsqnq6aWji
o0xr/OMoqZ4mfZv2WDPy+gL/oLWX4EA8mDoejFXc9az1fwgoNsWzGu8er2Ye8musCDBv2/VbcuP8
IcKXOaU2zV0czxlt/+e4ichq7tz5OXxyTE2tQWBfN+pZsMaTSpCgyw7s01dDDRW9if9DdHNWD2kQ
SROx2WpHAjM/vBiE+5p5QM8Z2eWzR1DonpLt1WFcXaL8xs26i1Rz/05HosDP/uchZBasZYxW8TUe
HgFu7S4TNNf09cg6B41T/8v6EF2Q46minqxGw6Y0YC6CK7EFVUn7HEtEj37HUGcz8IeOuh8EGWp2
K9rWCg6mx9Yav0X7YoM8FWmvkqwl2LQ/tn/5Pyf5KjJh/3TM2s1hsERSTRq/eM14OI4K2q+r7g2Y
jAwh5MGNoPtghOmgom683tt+59C6xy8tMLD91ScHyyBV2JazUbDTwtaTZsj/SEtNmqCSnsJ06vQv
0yZu5DDaBKXcn5pliBqjByII8pS9AWzwPZEVdtdvJcSZ4B5PF1WXILOA6h+mkprMlSE6e7TCIoFz
jZ6XguBa8BRCzKzQj3jDU/80vkWZRqrvL8dnlU97Tr/g53KjLmRpFyWkr+1QUt8scVk0A9U0ybt4
mVfok4s2F+WfJ1Khha1Kcpz8qKpWzc1Y9cMlh+A3LHckVPxY1okGv3ZCFubUXoXEpINwCv5Sj1mF
CacUzph5l7CLc1ysMBKQx9a/HpuUaKXSmKE5yZo+BT1C8wZTNPDx4kLXmeTN6uOONsGFBDLnRSuc
R7kaSTsNXZEmPgW+KkBV+f3FHMW2RwwG90EhvRVpbxzstcbQVy6l2E0CoBGetAOU7iP/0pWBcGyH
nF5dN8FRmIZkavL8agzqB7VkMM81nqFnMmmodm3sgxeSf3VOmmPIXDRBfPuURR6e2ivFvFqFbfH9
DYxs6jYO6q8+qq3azwklW0YkUfuz9z4VrHMIOdSwO6pxH4IEkQJoZWNh/0FRn2p+BwldzMAu7VJe
SmmJElXlj6nOHNO1OYcthrOU8hiN+XQMfxWSXfGqkZ91KqCt0szacbAwHXEqUOkUQOF9WhA6/2JZ
rZCTcRZMQ0ZCWxZ5yqf7MynwI82R1Zm4PGzftiVa+p6Dlxhn7pvYEb+5hm088M7MzNXL4ffyje/C
6WW8AM11LuoyPaNU7zXcAQL4rqd61E3YaDgDpj4nnk9e50GoG/SIlQIM2tMhG92//c+uBUutTJoG
6g3BJ2ZuGerk8gEV/4mt53Etzz/Hkmlp50X8tDzl4pp+KXevjL9efVsB1s+m0XHnB47lQnUBbTby
7vPkhEjUqkE5RvC4zKcCY+wiaCN5RtWFWwFvy4kI+zZ1nWU6rKpDHPMwg0I1hHEMgT6slhGyCKDj
tZcvXyrw/b6T9zIjNJzLyaymiKe5ZRyZzKZhvwe4Gh9Fyei0lCW+u0U8xo7nafaudqH2JULCAJT0
LZ/Cst9X/k+zEWCWtH5RHxIL9I0QlDNP13yJ0FuuiXfNVwK6wdsPThbPgFlrWCmm4FG1dox/Cbfb
6AvvjisD+/EJX2vNrFf3De1nOQOE/kaXhcXofC+HZxU4ou7wDxGECtw9VbfUzDTxkt5YFcwVIUpq
aHNQGLI6QA7jXP0p6rF3j/gnRqINsm2T0yJ1uol4NA4PBmrbRf99E0i3K08LRrW8kMrGMMV9BKUf
G2C0WYPMNQIiPGYJesuA4iL0AuFkQYci9kTZQsftn2yzYEy+juhfuEuiIahCn4ZO1vwa433rHZYm
n3NOQjfvhMdqqfz8LbGuysg6xf25Be3OZ0ZGf46goP/8z6IE7kSg6d2z73ZFRmp+hvpE7elADzys
0+RJWWv1yTB1yKSPz0HKQrJK2ZDj2x0xb9jGwRce3owwE46woCUAG2v6ELuc7i2UkozB2D1yBIJG
B+hXGa8AGBmT+GXoDv29c4aQLA8XIdGwqMkzBvfeZFHbx0Dm4KLR5SjMG9CUW9wG/2DassUsGN03
lRt4IDWjBt/Y7jCQPm5br9cOngk9x0mKFxbmpTaeeMDCcwaLWnOqXZxfMRRCrPlBLKqcPPAY+swP
vU2wDh+P+KdGzcnZJs+8Nfkua7m2CYzDOhHsMqF34iRMStaabiGYAXckCVv7sar4vxG0KzZUIDYR
KRPbmNLoNrNBstmRnbZUxv0CYVumM9vNdxOgIV3s2Wy2x6DzYWgjbdGPOPYTbz8sLb+7pQuIREmK
BLpz/fDVcKbbFTYm9TLy6Jx+SR897FX6kBNobEiNn8bxsQEYvKgwyiRbnECuDMX3uQ8tnyVmHKMv
1Z7UnvBQfUoyh0GpHj5ov31A8AYF3FRAivsqjOOJqxwgRIr+75QM19T+Ql9ALhI5yDKsn9+JguhQ
HN/RVCZyae0yU9QXeazxnzXUZFMh0GoYJwZ140sYx2P0eG677qVA9/QLcw80RBFTb6wSAzyaAHZ0
IsQFmBD4tX1uQiOUo/jJZ5o582uvS3x83GzVTCSiQlfuuuBjJYIW+iCw8mhU7d+YaFfFvudjgSlW
mvwNcXth1k3GDwwwVmTgu8nteod5Y7IuN1cfyzptw/cks9T3t1029MQ/xE2uOd3wJk23TlZOwYgb
x2LrCBs0WZZTPf1xnNdayI4KlCYooMlRmWy+U2WvwPY3lolSyKAUSJg8LMVjBFPJdyXvIVlJNQCh
tEI0OUa6OqEtQXVV4590iuk3r6xh5epGmru0rNpB0Zt5juliMBMnd7D4QNq83EXjTI4XYVd74O5Z
xLLAxrYc8iQV8S8ZlractmNU89lL5J15r4FAuht+SJyI553GsN8fEN3VwvuqRAA95btW1DS6GsTB
IDWhWapvle4nGwj1GTFUE7sKTcXWMrloq2d6FTRthvv2rTdJKqI/vo4Df7+0f/z4zGSDNQjA8229
zWgQjT3Xnw1LkmS81CFdSJqUKNmqFmxrxIhYVPrJWs3Ci+sAGvvNWr8JKNzl79qlxCDFNpTqpuOT
dCGy7GfELkdYMn1rcew/Lem/BQBB5JwSmZT4gqQyfCS4yqb/MTPYA0vhNu1IUD9x/HJVDPphqrqB
rn3AlCxsEq+OQ/IcTSzu+k2JA9AdDZj/bJSz3NaLxggBvAu5KisDQiskFf0qvIfDMYEJaNdMDsO2
dfD7bczImo8rO1sGDkugEYmS1OzTm9BfQy4jUcp3G+EIXi/8r8ezB0NXfNXK6swn2+lUhd7ZND4l
S0WBJw9UtzUkTmDJ5cvp7CKmTLr+180Uj6GG0irEFlId8udQgMTBAB8P2FvlFLLGbeR/jrUK2rzA
gogOjdLMCZOGaF8XBeNtYsnm8OkKFRhGTfN8efl2y5RLwY9HQpZH4hiHPZZvAmhhaYz8W37FjNY1
Owcxga+EVx3MiAt02nZ6DwwcA0NanMl4LwS6YtR34SNJgERwoco36+5IUbUHBWrHa1iYS5xC/G4Y
Z3MQorUkvWPESeqZGEFbi/EWXYheU3CIil57ZHKAwUj1q83sJC3GYRlYQt7BHr4Q3cvTr0gL0IHd
eKC2/k3kWpYs7UZtZQXTHlmB9T68J+2fL1jdF05rJvkGy70lwXqG1LTYhaLyyJGQ4OO1gUN+g4du
CUE7qaJ3Vnl7sCYgfQvBLjnHNKkqeUHRebODNJX4snETYJVMdQjSGmfYpeEij7u3v54PYIOStomn
ONelmkAVfKwq46Mozt2+pB0CwxyIL8Erqi/m1JcRoxkfV+zIn/KCHJqsLGegjrXXMG8xLNmJnaFw
GyUDRHf2AS/ET2DxuOd30CzcLt4UOKLcVQLBQmaWqJfneUKFtnWXERmnYLc6ILY5UICmNV0UZCfw
H5FQ1CmqB4TAn7N9qkYgoWzl4q2WaYT0q698xLceYZp5jZsRzyRuNkP3dK9x9ZQGIMNIJGg/o1M4
hh7mYKiT1cYAZxdu+nBFuylZt4Hjl6pgtiidFG9hvydE2olvQB4SUtqzurZQPaR3i34P+f+Cy/oP
kG3Hu17m/Ouy+AsGurLzKq59BeH2HXVy+dqS5RDI8lEEHDD/mrbh2MGrbzH9yu9BWkHvdU88kbmN
kWdR25+iLEaH8PDJkhPsJMJ/v/D1ypJqkU34V9lxgzi4o7eIXSe7JxTGVTjCmxD6oaLO583G2AM/
ylSUUP1v8U6vCclgAOdtjrCkbisOLjHJLDDaDHSIlFYixH27yBI3GbU5iKO1oSZRjZZwCoWU3QnO
1+GWEB/eWLSDu+d1iENonm2qlAzhpmtlpGGNzSLHg8IgBBJ3ya/FH/9mtuH7xfZsDxkFJWtTnYSt
glrggD7/sGT6bJfTpmJPhttHGmoYstdJUC9p8fpHryu3xenGqAE2Ka8flqyBrwH0Tv3sF4yhr0ZU
K4D9ryhfeBT3QcOtA+zbhIsNNgB7SIj82IUOyqMeOfrVmd4aUt2//3N2w8gntUs0Y+hOh+T9nloH
G7PnqoBWFXncd4qI30RsngvSEzVAZK6HxFKwVlS/V38tN47Vg4mzp5s6+rRYH4l5jJ+K+PCET/LD
57XIL683FNJF2cxVgV+sh+Fycl5ZqaIxXs9ySDGi380jnl+o1DU8JbpM2IpGAIPy/5sHTGynvX8v
fShk41q/Sf2W8k1cioy4tHo3t0yaGOrNe1YxVpzDzMDBU82CSYXkQq5IGfKhHTHUSeYB7h4MMVkq
UORDJbX7q92K6cVWIX8R3dVG9XrKyy+mxrKAPtaCkMGuzR7PRagailm9LQtJ4FTqWAAQ4kh0GTlB
DjSJQLS7PcM3JsgRiqSobldZoPj5s1BDPKOfVaei4lLetA+7ks9Qylb+w40gV3x2tdXMay2920h4
QibZdjJ44JA1InPSySs9fYLoax2JqsVpyVPRp6oYw4+7okgSqsNpXnQ/l6RB6yHQ2SajIUlZaJ+J
zgU/acp8cV1iuYxEJENhTzhFPihzXly1owVxZZMSq5PKlk8go0KTYftY12bV1JrUXddEOVWeXtm8
j77YHOQl2aeT3uJQEBHup2DuUAkYC6itNKtnNc+2Gm9EOT23zF+tiAka3Ixxn5Ak0OuSRbZQ/UFV
tK17obqfP9VmiNTNEilf0us7atwcjd98iD33+Tn0v5rZB71B+b5uzBLPqVhMavS5P3eZzCHg8tQi
7nFPgR1WLlAW7p4uHANM1K2C4bIutC5BeOt+I6aoFNZRo0OxNpYZcZF/ozCIdU6UdyW4wE4sfhfw
4FqV4G2OczMyxA5l2WVTzyaeqD7iFyptdYZWMysSh4XQskpLbysxPTye24NCKwAvIZVezu1HgzZm
ag9/bW7cJt1gvREflx9wzpYxAMWvTj49jYjKMAoCydVXQATbed/4I4kaZurAeWQ+wJ/sVUl4Q+7s
dW1NllylbDIIU3H8R/FcB3LT/e4FF6G4x3RIC3v4bT5woBZnjjuYHWKvEcwAVJjtdpPinSx06MSq
15MNxoJVaRFXbXB4Tz9oCq5Xq6PGLyZ2rhITeUTvgMJ3NRzfXpCsztTy3ci5pKG1Jsa0AUd0VKyi
sF2Z8oMzCTpbCIU6G5AJUfTuV3XSZcwg5D8pKap3sC2h+SJ8wYXWZGlQAeH7uheHr7HU5OYmrjTc
gJ2jv+De0xjBB/Kf6mXUYjqdgB5ELakqPGbWqlbphl4ZBPwRmS2TcvMh3zLXFjNwgZ1tyj+dOsMI
g5h/BXVO/I2GleQQqzz9jFhVJfT9TJ3SjyXvIMXqFT/xHvF2Mz8Ph0p75MwH8l67mgbdaL+v2qqC
orsQvEPacWiIKwa19kalTYnbshjbAlTM3ZAf7ir67tdoaM7biizckq4msxgFR8F9vzzuWXf3FPtG
/7Dn0Nwz0qrusNpPtJd0pItOi6yM+1AoLo88HCYhGrN8CGQ2+A3yqlQcoDKY3iL5JI/l0KJFMCjk
WReg7xSoLfLS9uvRnmPYVz3D7fA22TIC8iEViG0Va4rRPpUKfg+lr2S4he6O8Wb9jCoGtL+iFi8/
Se11bpyxBPcI5aJOJ/ybzPaBJzWcK30V2xaL5Ha7/FWjuaEBSvfqa234qzloj9bXMLCJTyX6UxuW
8SqpBCtRpTLddAgLBEGmKn5SA8BqpaA23IfUwqdixWv+pFp3604imkwP+2Wx48ITq6A6lZkV+rZM
QXq7mNlEWd/Tdr+SmgG334mEC2/6eq/yK6/p3LdFwB/FivSdr2AzO0zG93D47bhzCP4AxB7V7Jyc
1MG3GPuU/N8xrYgd//Ra40HeemVOSC2JXPw2GVC6DNnn7VQ2KmgyD4YQ7/LEm1z8fGPDlOGm1syo
ExVV2Jxnz7CrOuWPz3DX4tZOxo7lnh+BlH47xH8H19huZ7IdMKp20/8aqNAr14SDeOZ5dpwKiHdB
ktzE/9sp6f9P4Wnje7KTbzuTTmHK1QEbR1FP38yWwdY/ZhC/SMl/EXl6jQZP0uHX+S9e4mnZP0TD
B6pgqTk1yImdGtDBnj3v8u8LpVpTG+COaYuId0SfgJPUFvQM55x0SSy2lYB7AKAvLiKx0DQC+3Ds
Tx6BDMjSF0dpjw8gLsbdYuirJuQJXGPIcfZik8Il7BG2ekVlnC2B/zBktMk+jn21Wan54VNrSfDZ
zuAhjynn82WgPQK9Z2/aHIHU4KJmJXh7uwT+szGC3Dsezb/QwkMYvBGMELO+I7btmfyNCRjZofpF
Fhz/3ZKEY3/OTLgWIpUX8AnAG6vJa62xBR/8UCLCvj06nidgt+prK7tD1Jsih5Aj/3h+zkPTY/aC
NCu/vva4Gk6Cwlcn0yHnnmaGzZ3sc3unaEuE1WUvSbTfeyf3A4G1J6+SoE7aU/x3appMlnuOwyIh
jb3eXe5+5A/BFUCx6yjEej5ziwcz60DFDXSOn4rjiyIxSJUPn6iZp131hluj9rYhURXcvTCzLzCI
5dxZIoXt5+hD+snbjAa21Shp7rohZY/DM9kSlHUM4lgeaf8lGb45X0quvdvypIsh3RlZcu7m1mUf
lxmJr1rW5R1aX3Wbd2TZfTo+g04EP3VzcdrUzWdqrVAa+d/f9+MFQEhRHqhHTbu0olQ3hjFzRKBZ
H3M8OuEt7dQrrhew159H8fpur6lOFskHEeRrsd/jUgJd5mDOtAV4ylZoBqE1OSf6XACZt/aq0Prv
nm6+yEW2x/RZbLdbQlz+DBCFyNNYr1CHzjJl8ncn8eAIu5Jnum/CZEhJ0eU1h9OoNQPNnzZ6h1sX
iQudZEZdsvl31kzWwzFKcdLJIFKGllKwd7UhcKcJmIlSx3zN/LklV/jx8a7cxP9C8HhqbZYiMu94
IEqbzGC6wsktCCnKV77fMBZKnzT53s/wsFg0FpYKx5lszvip5LETWpgLIbQ/pDbZnBd1QxiGvVRX
mR/gxWNUGXXvS8OzZ8LvmK4EN/n7KgxWC7HqlRCFROLdQDJqb+9PSr0/l1PtWvCOzN5dPHJfXQtt
r4nd9NzJ8h5m/ftwu1Z4w8idm7JPf74+YiT27bMPpJ94g40rDn4+o23KLPDV8OktvWMHcplOAjyO
nosdpBIQd+s8RBK410ZOB/iA97yesxyL7pgB3bZ47aX7LUjwt2tkGFQ6qfg6EvuwB09eAGdz+y+0
4zXWBCc++r+yR65JBVmAYlUVAN/4NNrrcqiMWQJn4lTvLtqEm5cyWwdHVhREUs3PONbqTdDsSj7T
sqePGpipsUVi0sR09gFdlwbzaDfEWDxpfvdmlxwyrXMzi9STH271Jz1152EGryliyT8cgVdx0UYB
cKMm52e+QrgiGU3ouOJ2ugl4EojV7jCxENMW2X/sScIa8H6ERwQ/TQHdjN6sh2nvuvRxAIPdKNwc
fkNQ1t0hp0aQYWiP6bvad7mbXuMqFJc3LEW+TY6GH+DTJ6/Ox76t4hfhaYbBzW1Qm39T1Xy1lM1y
Z2l/IEA7LHsVzCZl/e98TmFfqJT0KZJOaVoqQtO6H4Ia2dc0/omkYBqXZeyVYdXucY1cPWv+9BlE
Vm4WY8RNBbKW4RNpgtuc4Tev1DHRSswp591TQ5WvLirA8GqamHjyR2IsxgpQ7ykyLGPkaafYBGOQ
1HZC4VKQKT+eK37k6pucqj6aFqTvZ+9USJHOTgvoXhkQ4uqnsvXfc0Gka5GClClfMJkXX1rgAslq
oLD6xLcfEYoCXbwQdb0YDD/aC1fz3QLXzqERp2SDAycWpMNEdOtTXMLImn5QjZJM7Dio0rApQw1c
X5Ol2dVwEkgAGp9MMMCUnH6+AIYib1sA/zQr+jgSilyaQOgzbO6bhAzsBwmAwFXSSiE5OrVj2GzZ
ZGxfgE+MGszjA9LtyKiRxB2ZS0JyzxEJTd5ojD86g07gw/E0oddDpEEPVCM5m0lJc+sWDKCP7bBg
U5ZmfrA5AkJpESWq0oPsuNmhC8X/HagO8/Iug5icWVBrgJygK9LpmOwB6tGEsNkohlGPEcmdUnQK
XPERSjqzcdzTbnXXzu26fSVu2zZOdh6Oc/MHb87yKpGRDiJa37R8RifuPC+5rPLgA+flDTbx2lIz
Hx73bX9KxDCPVHVYun5x8rUuwdUrAAylXeTgXjdvMHzhq8NYPEPqKc6RuUSzF0cQYKMFHYB135Iq
0ZAdKYM/IDYbIo6UZaaNc8CClwqrci69CDtZigXQIKPhiFHj5497cXwzTkOxSKnpVHFCk5w+L82c
Mn7J3oVSD62VMcvAq/38LQLNn0USNJAt3oSThc8yexS3+DHP2jXqy6lZollSTzfPKpwRfpSDNa8N
Y0oYCS2WOrkz8EM2P+83gdMmN7M1Xq9cL90g5/pZZ1I51Y+88IlzmF6u54HD84z+1T5g69dHWUpK
JAb5izI5QrFqGHGz7D3YSanUfZ+fLX5/7/0xYxh/qTncifdJv8Q3Q8heQnnB021dEjuDfdG+wh+k
//PeTs1gcVZHvYul9uxkI5/WcfwyrIYLtgw9/N5EN55/tcQPRuHAo1NogfCZO7zH9fp5jeaSt/Ou
QZiwrU6GEzCPuweZEWlLvsEYFF53dZkNIHtv8M9MEL/OJsVkSpZKBHjOY8Q/22VEzBVIGl+BnhYU
ES0HU7811zkMmS8Op0DuL0x1K+USmP3a+Af1xoRpOkE+lQlFTTNrmPZDgdIPH023FsXegBp2j5M5
AfD3XFr0A54kbN7P4JeglaAPTD1YA72h2iSkBbSLVQ6NPLOGX1KgzyqyJGqJA7LZGQz22iW278LS
fuvZ0mGAvGGFJ3WW2dUbep/garM501WTHsqzPbUeAr7Fu0pPhPSOTLmCs2sX35d1RFdnDFfWbZNx
fwYPNlIWnZts6zhIXuBnIoiGaF8hz5gpJIHAJ7ygvzHkuB6db7mVl0Y3St0Nkai8tO9cPlN96ICx
FA70prwYZ9DEh9DSyg1g897qv/1v+52ZfjM6bzfu7BIS3okd+/ceBzfoaCkwTE0oAvtEfGXkvUT3
aa8FrJLtyr1hQ7t01ODg24xUJ0oTEjMe3DwikWV35uOD+r4jCSu3v08x91uzBbAIHjYsYHXMbN7e
GyO8wq2IvwdeZ2ms7HMgk0gFtiyMLd4I1LERG0R9Sgs8lJyeMNcgVzGrp7IhC+m/u/PHW+w9h5v9
HONmxF7wHnWXZkSjKAVfL5Vr8z/cJeTnn7PjpTpXQDQIha401JM+cQjkPK4Qro49LN5dn7xJyuWT
qFRouTJspXU12I1lAPAaAuQHfWwDHTzOafJxjlAW+uLCQtBGYRjDs6bMxyS2H/KMSulqCmCuEDGa
Vq7xxR+UPNRPT7ocU6vK4r8H+wN/ZOMVXC1qdnXlUQmC5xUU7NHyeJDZAAz16+G2B+Is5hhjtfir
AP1A+45ECNN6HAdxYaPglsF2nlr5a7+TLlSR48Wgyv3hddRBxhQQuXlQQiBK1gMVDCGyntYkyIkN
veeEt5ybz67nYkMW70uy8BfzgzoBVX0bZbNlR1GwWHSfcI4aeJc8JrXiSAXjNh0SOmAkKNYRDp06
qRidlrK1/xbXjRt+ccoWEr5DqEaq68lqhkt5WbwGN3AVncAQlwBe5P0WZ5cYhrNF/mKI3tjK0zZ7
SmBAtkbpEI24YrquRVCOVQ/7R2F6BM1CDPt4/7VjEl4SdA/ukXZSVsqvQlNVhaGAgjOk/Rf2B3Iw
VuECVdMdmFoC9eBPQLMsYd+oBMly+kpoAEzOgwtbS0WGB7O5W9NMW/udGsqezDcXf5tqHqvPalEF
Gd1E7knHEcOX12h3m8hlVEN+txMDCpvIMp+eLb94HGomrmZmJDYalXVgbVXNO7feoZHBCcglrOLo
Hn/xmcw+C9X0qHbEn1toZ7sSGuj2PAWpBpahq4U+Bggc/CUsf+Uv7UuiQ9HGLuD4+0WaTC3sRwtI
jQbRaO/ZsQ4jcKEdRk+SppcMO3iyOuo3uhJmxaLpcyepr62OT08vga8cTTzzKsj17hilO3fB7tYQ
riIuiX7JHDp/e2n9LpFz1e6zGOdgEyhrPD7XZ05gc7BFdum6S9Gz63oOhyTbhtyc3ASas+QYZplM
ZMeOKc2IH427iE8NYT5S4aFtl03xuG1cBF2f1sKV3cMqT+BpdrZlSgWOUJV4vwg5VgVQFlJ+rZY5
9bV97sGWM8RMXSaDuTmCLVXkD0EbF2NmT0MPYhOPT8SjW2cTsV6KH4iNmMpYxHQ0Sy+wrZiBjdbv
+9mAFxuCJ5hwVt2CBy8UmzOMcw3c9PfY22ab6MRBChY24ji2BLADpvKL1Lyv6ifCBei7EvP26LLM
ULqUPKZXNzWOXf3kH4kQXjXkwmpfQ0jKLK8GK4nH+DhPQVqdFaXV+qjAVj1CD16f5UMfmGr+kvZ9
mz5Prma1rs7rKA5iqhU4TqH1a/ld28iv4yJn4JtTTQcSlfLjVnaJl2sEfy41A1IUxFjfdt14Q+ql
LQsOV5SpRfdoR1yOEhdLZ3u7RDaJwVcFoEpq9XDsoeoSfHn4Ojx7jkonBw/9GPRG/YVj9HoYRcig
z9OptEThe/owJz59/SHTHzJmKk9cmnLIyZd9A6l4qoqj89ui2AtqDvRGGWuyK+WGaMLYBZfdQ0Zv
/bQ8GiSOZwhedeeyxm0w6V9k1nRpHCieA1HlYvkTgFXEejyjnOGynprLhPJYz6dpdr7qBJwuCizs
6TaA0d0S5ZxjFMkAcHS2M9lbOY1g8sSjbPDaXNz8PFsoxV1onBz5i6/7uMlsyDqSmb461LjTK9jR
w2iO2tOhHUKuRAFTY46gM9F/s+pxN8EJSMxrEbuzERFT3MUWrveBjTREsFCHziY0N8u4VYUg+kgu
mW/P24ndBF5iyFqRvsQ7/1DswAPpkfOXp+ppABUOhBAicjLooOtz4HjlGqlg8ib9vviKr/SlvU9b
wOpl5NYTB4qpzP988SRga6iKE+SFPuQx7rI/mF0GO9FqekvZH3ySe3oXsNafs2bD1HnhwT3fXl/d
MqaPaLwRIUtSg/amcJS42EeFHvwThvNKJao1WhSuWO/dg8hmQTAthT84R0MZltFyaxSHbhoFA7lb
PiX+08Ey2fRV+ZFeuGw4Ot+nXPxp9zafEcDhrz2XnqTHcDK8PbyDQnvaw4YhM4zHuMRZoOwiT4V3
BFxBYqZPbaWRXNIZp8iaKUylL6WZ+opHkxlo3fg4J1dVHUJJIsEvhsOeMX+RXt1Sf/qL6f69x3f9
MYbEkNPIwn4rW849tVaqkJ2sj0duzOJxKze0e269XNdnKgKvdHTG0dz8ZHe0rZjrcMUYvTeItFVT
Dn2RFxGXKT3+ehlQ1Nj2IswcxTjdbzReVWjt9T51p95WgHhLXHDmhCpEKGU9emhbvi74W6JFIia0
qOii9qVSUbDSn3pTMdMNXi60yNJrZjU6EVtaq1+4nx7hWD2vWAp/IPqsyAqriB8F9my+dtLc2MOn
yI+En/WlKqB+YMy6joeRh/sUAInVC/73GL1O0Pz+rUy1klBVJ1/OUh4CyZR/qFPovWtBDvbO27CK
S/8qxKWUu1vJJTXg7BLTLlGZY/FkjTf0SLzJ8QRjSzwnndhUyP3CMjiB/gRX0/oiO1o+XqYcwFJe
uzuGRsOKn3ChpBt6Z9oZcJ9HQCe/pJ8NPJ55arV2IlKdExLeJpNC9JKsoXbHksudeUnM3G9d+aQE
xh2ydvYjE7EmqKAH6BIwg8Cgk+ZzwnpSD3DvPGG5+Y7niGYVLeXM/6KTYwsZOe7vuWVvus03jQY9
h3zO0ctv/1/Pu0MsDVZZVnaD+QpFeFwyR64v7kD4eGBop4bi9HIRYv81D7JBx+lEONH5Z0axND3X
k3uqy7He/Klje07aqiIvUezjizhdYEauCjtw8mB47SU7Vk2oio1IcymXqTVYYp4vD0/Wpx3gbs7f
0PvBwdXRACcvH8VTKdhVWGCXsK9T23waoZ2a0NBUdn7+Bymz0vyBxKIOog3MVvSg3pdAijLY2mNL
uw5ikDfUvpaKPQXKXN9xgufWqLwixO2XzmEmJk1o9d8NvpRqdQk6bAU2vDtov9ZL3l+0nlgbZZD7
LBk/AG9rASq6Vytv6Kf4LdceyWZPkfetSMoZicOT2MkN1gVSae5CxbFyjLr4vQEsySPySoVjmrkZ
JiY8VEtLFXUxKnsPL5d0VfpL70f1VSWR8B/nY4VrqsHIUaj90er/p4Xv35suW9USZj2e96T7aC+7
g2drxkv7RN+ZugI368MQ282kZOXthWdog5Y0W46KviHJDwRZGAwC1pPdG6p4BZxFUbPqm/h9Q7y5
nbJNjgLKZ+sNcqsoYbEGIPIJt8PqKK6vVucQyzCAh9Od+EsiD884asIWRTtbbFBEY1BCmA9zOd9F
WNadSC+P5ROZDlD7mLjWscvME74f64oT3mi+sGEi1S3v97mLmlIOSu3P/d9kKvFfXQdfrPGMZAU9
0kRk9WsqGzGHABTbF0F5LBiL9xtsNbo1oT3TWeUn1Y8FAo5qqybs5O/5xbMDe3g6s1SGVoJtsTqp
8tvmXFHapcEO/8dANY0k0ccscJHumXtDxQZXW3wGItK2aYj9xPogz2M9xoMH50YHxCYqKqUbVc4/
usNvYxndhMvgeAAQVrwFWJUCepnom2OcQhUMTJ1V9eDyx8PsXnCcbUM/WM12+9j1KqKnnSJ+jduR
Lpc9fOAaP+Txqac1zUhpvPbsxW1F+tuCZW6jNMx3SVjRadYFv+4lk5is8PTg+iQDSszWqbcw1ync
nZ38hhe/b//mLNT0tOIVng5sQhWm+kNl80p/ZURXCl7d1x286u8dPComtWk9NwC7SemFjHjEndQJ
1eTslCmVho8jCrjCt1hUjbr5G3uH+oQpZBlM+1fLvFjmxw9Sc9hkpSRx7bNMhhLTxaOgzDNYvuoO
0fWbTGDYL2ENKw9Kj1F9xKQZb/D2hNJDMAmZm0Xoy2tLyOnMclrlOmbywBLb461BUMLr82uTZI1e
DAPyFjpWSJJ2vAYzzH6CLhSotsXWrliIpaUKYG7vzrGrd3a1JjA4x1Lbpq+GHJgeFyTaBeAZGDV+
F9e/vom4eNTNz0GAuV+lzKL4srwcAiteE5xLV9oFvBHAKZUtnZ2vWBu+7K8Ndg8WMBaaycRZsrwu
qXd82nAnoR8mR79mGwzQaUjiJRGFENEcabAK4bKaEgaZhLsKOrl593dyjqBvydZeQ+DS7fPAInRM
tRiIaaTnxpC3WwcK9Sf6kV3MbZB5gBplnBePROdbzMRRk0i94621Ly9fJ97kb0m31HtSlzqS1SQl
DZn+HzE+wAv00jdjjsGf7qSeqoWVZF4DMtnpAMd9i85fB/t9IHCc2yKuX8kr5i8D0/qFL2WDsbT1
gm8AYX4A+IRH/dhp6eKLuWDPER1P/P0H0l5zTE6avUiWYZ9IiNJobpVkj3mfqPqF75fZonvpKHD5
KZcRxoyCpyOasimuTEZTtfLmMt/un2clwbFcDUwSWDfD4849AgZONYaVhzhggGfOsUmDZRJ7ONoz
cmEjxtTNePqNgtzO9gCYoIeeh16LkOR2mg6LY7LssYHdN0grLFP19oBMF3hJJ2MgBj294k4hVJV1
HQQQzslCz+CXWRtYCTg01FGehrqOHzycccEdbxMjSofbnjZsn34M/2xpZBUQSaUcnMp1MI4GuZ/i
KhhXny2izSgippy0xjpZLGQQ0A5X9OikI73BcxmMlwM/igcsxXnZ2n7AOB5srLNogIde04cCQFvd
GGfV6aSeYQZFaYavKWgE1CMo0lLGWddkQ3bofyHA0xN2gScTwaY1npC8JJ3H5GRWkkzGUG4oqf+m
PHsBmb6xP6OalTfUQ6WfB5RFDmTZCTW37AxyIyWomuJF7n/8ZkiR7+C4Y3ZQgUcGQsriXHfbYbDt
n0TQ2baRtMY5IWsQwwPnalYeBeXzV0ZbA/BLgi/V6b/9pZyM9Hfh2HZM34tgyGELCaWwh27KOZvJ
XKveqZ4u2j/cMl9CBS7mqYo9Gu7yeYSS8bkYGbaCSxRlFe1g1qfMKrFMx010BPZn5Q2VBUR3KUAE
tcGTsFM4sXGWGDomVDO0s51d0kZrYVG53KLFxo6ZU+kNFfLw83Pl/j+x4vZtPTfFwLjzxpkoIqP7
BtP7FUSOgVnlxe7G47+sJbhRjl2cBODkDLxaR3rvAETaOC1qCsW85v6SxdrdrdgJzfp8Ee9RWEnp
BHFHz4mY9jcU/StCkCutG2CAvvWHPlrsIe/rDoyiAp50aaqrwPak1ffO0RGdL/Gezsj3Swn7USgH
K0wuOhHT3DXys4liZu+y6IrltO+CP9lC/AD/haoM5wuSImJvTB3zUx7g12VzCTSgvLhwd+nQA0RW
IafjEJ3JXXgyLLvgXlQR0LGR4fnxmv47Sr14HVyuaEXpp9Lrzsux7lDcEK2er0SHy0malYIYKnB3
V+HedFoHvRYbpOs15BlG2SZZv1flExd1FyI0CCkz7S0MUWYx7ZS7Pdomjp+CjZ3neiA3fALt5jl7
/VcmBMxzx4H0S78WDBjGYlha0T9LgUMS55diCGc5kunYoQ5AqaUbl+pJKpYOyz/T4Wnl2yiEjIHC
RcIgAMjeN+w0ik5CXB6oV9KcqlFlXjBKwnVGxb22AMJowCJBJXBZROCKZRlhsrMFJ94Sgi/kZdsG
KiDDkXj4Mr6OqpEgif2+tzNGuitmkQunUa671B/VuOrll61MwdrPeiSC8M8b6Nb2ymB3S3hmBXSI
pJqJ+S622aoDnu7xhEZAm31HVXw3B44+PH65WjMB3O8iplloEU++6DvWIi8iSydrZpd2NE409TA4
JKNhrbSjgyP9wubywmloErX1L+mcF4Z193y0It1FIQEF/NtH4wWCnV0vmCXQTRfeR+Ln5IqQLMAR
PToUj0VxaI0exZM8Hp8rN2NH9lYZQiGbgC5S6AB4HsGfHljEv2VXfaVO8hS/BecaTh4moh469rYx
EvP5Islt8ZibAgAlvcTc7ImvNyxRW4Ewq/p+29oaMUVH7YYj8yENWIDTrgM/JnQLm9vFPFsD3bqn
3jET9m04FOaDuulF//feHMg4eFqZu3mxik0FS0mC0JBoKRRuVjKBk8dKXfBtnhWCkxa9fUQ1JEdG
5nf4EkcaLEoCDtXcVmlKMtNRtRNJ3qa8N1CY4bMImYj+dIpOUD7w3RT8TH112JGQ12mVkCQUBMXs
F/Dn9/Njxdjy5omg/V3fpp96/xfEseLakj7NzZu3qYtYrnYBIPED+J8PyzXZEOqFfFjIx/a7etU7
BNNwgk0LaiS8qGo3Fxg1oZP/wqKqlmk6pL5Qp9jQNJV5TgXB6XltQo4I0wAwZ1w+kTGB4mHt6CGL
ZGZEUgtOZ7+bmEYhykOh5oQ69ubLEWsTiqz18ETno3Yk/hvcjlRGculQR8TcUHlziwCNaopO9Leg
vCTKOEZxiAZT9eFNHboqRRq/tBL31dQ1SLHCdXpV/0upcXccspJSG9bgoNboJw4idgN6dBGqzMTL
pwYsFYAhne4+KhVu8eMR/DPL/byghGA7T8+soh+2lzkM+mHFSm3FLV1rKls2zY3oiK2UKa/iDmyU
drbThOjPXPlQrCZb0KLpUrbuXpaRQ2/TCvHfFOuBQYmGousyfmOD3Qblz/v5h5aIHK2qUUSdIyOL
xCn72YAUzQZB3u5flcTu7R9+Xps0CPf37e+w6Kc+eyxETDf2MXIMEJ5noMjtBuQfhc4hjE8i4rvM
J2gDdSPMOke+f6klaEvVTG/Oa9QC5Tx9dZsd9pFZrH0RhP/KNYVc9giIWi2IgoA6FERWm+V/2+ZH
dVFK1SQxpn2V6w+WzjdS9Sbouwd9yMenHQz9o4z8423zIyii/dr3RBiO0yAeIZpZK/AN+FJk1Xik
ZDLJlo4XFNy26buX6k4OMXh9Sr7KK3VrsLr2bvC7XCN9HTjC+QsfP6S8vEq6tgI7QNSPYud1JchG
Wk2KYQjn4FxW5RxmTcApsGSaNRCLbx7+G1Np2Rg0B7oWxb+aJHW9MeMr8e/jpsShI+dosJNgIIF9
1u74+0BJYcQ5/pkEDmnQgHkusA9Hzt0ORqh8ku4QKvj1NtOKctx7AEyKaQpYxJte+zROdCIIg9p6
ODDpF1Vr+A//RxniciszqTuvM8tHHESJ2CzQ54Xlw/3sexmi2Bi2M7JXWfyM3z1q7CoNi8R3j5uf
vFkldsEHVEUP2YH/MwBBjnTZxRcNmjpOA/XRfMFkJNRClP9+YJA/orb8sUYf/IPMu+E4pexNAddl
38fkhk20kIKnDwnvND1oRs77eE5C4JSnbNuzzdlf+3uz5tJ2BpUFlUR6Ji/jv3AtbPYhMHRqoBSd
ON9qSTXK4pTiRNo0RcMK6VLN7wfRBRWIXqp9HsxwZCI/ZPGikHx1/beR3eGGYBzJjeNOaEwQzzRr
XUHpBAq4O7j6/GiDFHjyf1F0rcj89A+CowdDumjbZ6fhoDIf98WpzXO2O6g/TRt0wbRjjbwD9xTd
5mSUcamspb2p0PYQRlHjgCxNdKJjspYtQMcLwAfMl8KwUoETFelKtcuA8hnzvp0X0I2JD/KgE08e
hN88GoqXvtLg9URbrHzgx82xUnTgT9XCAiIp8LNsO0K94Q1cGFg4a8Ve+bopH1TJFbvUXgt9u5sz
y6HFMrOmgOESdpiY5mzgYlEsMj0Xiu8kieo9NqZJ2M/x1bP5Dp3PuYPnpG8BigqObNBm18NGlJFz
7/aJtTSR3dD8Us4vtxofN3q9Iw1vKoLCR3cu98l+y9MyxTNKG65/LRuaM8rj2c6/UmCh0QVehZhv
RvEY8WUu6DVeIjcxEorOD8q3d7oK/KHU0ZGqM3NqWYQjRyIciWq+v9meUToD1zRp0xMAEINYjae0
NSyn18WpefTftyY6FtzA+HfqFtHdKbOI6e3fUDbOrD4b7cgDa5nM+WW8T6PwY2LxqEGFRC9NTxtX
Dg/u6nfOvZR7GJvWwRf0BvSB/iqHvEzC7w+TJi1CPK4VJpPrzFHAmiyIPd7ZSZjE9w9aAgEkgTQ+
giCSLCNdg5uqdBoA+MVNcBLOhsCsKkuwxWtGLqOFcLyoV9cHhYmmKoKthWRC72/JJz1WSFDLLCTr
SiXm67LZCRmo+a8lUpgV8CIb2aYdRwHovwl6E2gN84zslWlvLOJpOvyfQNXXXd4pdJwzLJyKNiX9
yWGOKikJ/x1XwdXJ2CIq3B5BDRkOJbwAXVRR8IO2atN9YkSEKZ4ldtxrb1HDm0nkuYWoghWfcthU
Uru7IMBgrU62DLHyfCgYphvyW1kRPIfjg5TacryjXBTw0b/a7ZBREhS08mpcX9K+puYG6pQURMrW
us1ODXCmRbEeYADPerMoc83rXWSTjCPnbCv5h5YYAL5gg9L3bLiELCb6JduwHxzZUzBxn6BKmaLs
UWPLeF/j/opHgXI6yJpX+P/aJ4AX9ryaT300DpZrekiC7u9V8Wrnrkudru7T7q1GaScjaajApzlG
SxhBoxVbERERrCiziRq2QKxjxVu9fxt5fmp1QI1twR6oMbqmuWM6waHLUSxrpXeHTdN1e+expGsV
plx5m+VyEHXZx5D7AuOMUOjo38OiHQlC2qVod7ZkXCjS/iSWFvzXyzLpCLHehidLN33lQd4eZlgU
dw6zlrlDalVkDTP3IrBdwY5L9kTpq1DJAF6g0dWUM8uCqI5K7Z7FD6l2T8udDZI/elooyg7lIAbD
KYKVK3kMVYt7EQEk9SH0srJQP6WW098vuMFTJyTf+I/GP4DbnbnRNshjI9Eky/GrxlfTdpbyKrL6
TZnYl29lhGrm5EH4IX2RIiohjJrm7zQHMZ3i7s0tWuNd79crV20Ccw+eIrjCEmZQsHFecFUt/R4l
kGf0U7tRLkg+eYswDGm6E2n2ZNSX5HWyopt3RUDhnZKydTYip/kICjl4rgfQTcRwaOVuBjD84B7i
YM3MCwB1I701/NH6pNzmRF4X/X0Zht0rO8eLIqufMlGEkJuGVXxxThdtaKR5gogtZQAB+kY04b5x
ZdY8vkC3HGrfjyEWHNa5LVlcx2U9am1GgNEnayVDwtYNma3gkrl0SXmzTUrAISwTFzQDGy1uyEg9
hPFVt7S/Hf82q8boZI4/xsjTFbprm+svy6evWacsuuQHW4YnqKLVpCehmwKSrXgwqV3KvpYi+rol
b9gY/K6bk3bt2b09F4OhU0XNVmL/WIHBWpyya3KxBP2Pk0zpltOmZT3oEivgoJfTdxMFrpX/tsNO
JNcO+8EgDh5/BNmD7FaW7hUcijtw5jySeQkmwXcNB9G0goNQEGa+/3bKbMsTfWau8eNsIia+S4Xk
zV/w/N73L4KOYwzOYbjrbjdDlhK+tQfDsm2ACNj17VuNTOYeptMP0HMEz6YjuKfBe1Ff6aRcnHTQ
bGn0fmdYv01XXni3H4/49u/F5b7971TSh+TLr9hYMy6rGyoBmVVhXHT6OA9wXr1bogbxTE2a0Jb/
kQ8m6HfQ+AaCudDrWPWPVpXzhVQeVxmmbQH5aFm9DFOGn/LylE69bnI/C+FktCaY6qpg4mzE4Ukb
rHYIPwtuPPaZsP4g3ebhJTZ1Gveh+IWPJLXIl/K0xQSSoKiNGFi9q8geXTCkkiz8K/rxDUuo6LWj
5hJHFXIqKA/eGXhEHkFZlEHH1dwAL25G6+vKjc213v9dDqxUGUMJuCM/YH9li/9n23OzYqYtg2dp
jQQGZBh1b16HDXZwRhiGnQQ9VRHjanhzrXjPmP4e/apG42ShlFcMUnoGQ182KUO/fmDHfGn6pfSe
Qm6DN5qlY8Z0p8rXZOSljahM5/+3ypKP9CuPIMLVAa7tRXPFaPv14ist91B0lxxE7j/M2crmJ3dw
gn0DItG234ZuE/q/bxSwoOrXYYYVhj07qc0orR98TCPVf5bEj66wz5PnrzOwOO4bLHlzHCfmnH1O
/9JCd/+5WPdXo+aJK7cXBSMBoYVMoZCPoS18kFPUOvfqLgitljpb0vJR/5M5owagU2K2V3LyNQOX
JLziOLRw4zcJlCF0qfnrCTWiWTiX4Xo7wBdnal/jx9/LR1qiUf1T7m0OUiiq0hHPgZoO0i/T4CVJ
PSYg3w5a+mS43cicDKkjPk8JJvtlluKdOdVNyhc85uek4HiSr03XRuw6PLkLvIQm7TB4Y5aJILbj
u4cqAixRpOJmq2J8eC8RSlK4KlRoP6MmO+j7/TvaeaLI4khQWLZR3TZuEEPE+A/YlQGNCMcJSF/6
fYaZwYYNu3LT9RWp7LlPX98RLEQpIEEXzSfFPXSTZCwQk2EgSBG7YTIfwJQuU6d9LHWJOjVxIXNi
JvJJxlo7B8NNaqc/sCi4hSFZzvvSrZaQ+aR4mcY0c6BCEbiV0bKFHA2dZjMZ4UR4DSHJ6QdqxhJB
UFTn1wU0Q9JtDCizjvrP6h/3arDa+X3U4ysbk0aBK1xM+aG7MuM9DR4LgovFb+Ce+KbK/aF44v7N
b+y6Mb2wWFqJBwcZ7ffNNlvqqqKvIOurjeg98BZxd1rsR5Ef9wfeb+7kmLlywXfnkCA7z8/kqQgA
tBmL+NXiAaoZXPcdp/eRJsoFInUVNWdZqPnv8j+TLn9pPUVATKA97ihorX8qtM+YSAaH9B3vnNpr
HHKMKbGo5PSrWTrSrTLbTcbD8lvgJIvrzzYGmC8bKko3IIhsB4dtnDc3L8I+Y1lvvZ2DscudNGOI
HuGpsa3YlVteW9e587pzTvXl5GQAvR72dnbOcaypk/+6CGb8AEsbwc3JtlX7tLd3E0dXE36Q4JXu
6cNPR2vXFL4JKoc62INhckNcCLUt9o90ykcA/LF2KVywy0I3FxW3V0SbQ+04iFvUFSCFiqDP51SV
AhStALSzsilsbXRxD7pBnYtKZLEQocroqd4lhBwcdwI/NDp6ewrFCEt0D8a8xDKmIWk+Gs0rbJAZ
wSBHOqGeIa816By2BcDgc54S8B1/RxfuymiL6SPWvHU3zyILX6PP1SkqbFYe375FChDYUsa1f2b4
391KHlXHwAlM7SB7zNjvCQ6EDmIZWCKmjlXL1P1sqounWzm9oyGQij/Kb78+aVIqPwFsEm0k2Bbd
CrJEkgtpZ2FsnD0UAndlQZn87PvxjZhcYfAOn5RHuB+NjOwVI29RKira6sPypaNPYylY96aEYYpB
5Jc5v+pPh1/EW48GAYonYcNwfuAlEapsfqvSwdhGUxzpeIR0fO4cW2+SvzbUhmfPuUlSs/PLNiaX
rA4JxhYh5YIkP4LvwdmUO+FpDJEbnviS3O32QpK3dXkMNTv03nwGWXE1dE2sTC/3P/rSjjB+GpHw
jCCsn3AJudPRjOFyHaihjGEPHS38aTUJKhUQo+ZjlmkfpkcKUW40NfHkhgKitNk7ZFErLXwCVE/l
euNh12azVtXw4CCpxhOre9Hgza88HDULnfGL8XgHrI6l3kal0vDSX1TFwrI8pH37YEh9/4twjlSO
hII19pRDTiC6OqaLJv4MTiV7w3vD1LpRTg493/zxtLBTbIGmX9DeotzijIDta3JA3Jv2ohrs4QKt
Nyntc/CnTT7+8+oX43uMyAeN46qhAZWvO/GuFS8uZNb/8vbsSWuBHqkaV6zfItawmtXbhHUxoBgP
igmJXHZVYifaz5GhO8Co+Hpd75Mt6FRPm+ZdeK8ZNf7NExU+2WISpnUcoWZ0Y5aOwnXPmR+tGMZ1
zqXwpGUlxtP9wTAH4NfD7l9pACCyHzTaXRpmJ2U5emAziyb6Ua1wS8T8GZJI11indTmzwObso1AY
CSe3KsvugPTAM5qySlZzx6X/4xUrDEBmGVhklfbMTnUUg2qr+H5TmxgUV4C3SZB8mXrNsAuOUAEF
xFfWc8Uwl/g+XKEbRX+iOLWsNjeUobB5WBOY4o++OnHU9GNhWrV5RHV7Rj/x3a99wpbwHv5uAnOE
BtmGgr4nKVQ5tOROrxeqQzGTysBPJ1FkMzj8/oyt8fruvSgfJf5aBiAinyWuWLmoCFsmN8DAZpee
+3mjKE+dKuXXd0s2kBy+p3LI91M+99doFAgA0e4vQuIBTXVwSYYMW1NlIKkJKVNH0b/Jhsb7F5f4
d0FO+lVrZ0MBvkC7SgoVPxcgGPlPwJaN59TS555TQkx2f1obsrVuVNTksFHR7AoNFRc8tAdDLR+m
eDGaKpkXXNe0F5/cgdGV0jWKa4MifFSYlUMO8LiVoh9EQZDbz+uHYcgjad33MmnWXfJGrnNwL2sK
JLe4PnUOHZWBGV1BFDZt4hr3mhYP3Lu+dgA6thup/lvzv5B2nR4ESdWKGlCG5bqWmvzavyPj6rzl
vYOi+rH00XoHPklXf/ioJm6nvTMfv43L5Mk9ji9DZasESMTfqx9MsrQpOhp++wXcJHFy0PMWbzhk
MzQ5xN+jZP95jtifzFZR8MMnyu5R1K4cGAiDk5LNbmT+BJuV7j5d3n8kRNHXRFLWpLAmDOu2aD4k
dWe6+Ax3+bJzO0Fxh32u9QN1ZedRZtPKRuRGJppaXCrq2LHHxm/83bPM7RYw2pPgm/M7gq+5ptY2
ylj/CNIOEVNl/nrQLj9iPRDQg5wtciy/oxF2F0triL96I26dFODYWQoeJPB28o0//bCgMluzGT+t
yn/o4H6OQwqApr9WcMiF9e2firKSa1gSHsTg5HtNlRg5QszIsv/dfq7oeQ47XkpwrLW898Nj+jO2
HKM6war2HfxPk8rBiDaKUKK7T0RBX0PFH4c0Czf6TWQvIZWA7h5bhT/08hCS2oMTVnGLEcSr4yDd
RHnkI6s1bilcmxD0mojmH180kF/KurwtwtkTFysSXhjkBPLvjuvZ2oT4qXgl63ylBF1WJfTOicL/
EN2Ma3PWtLnz4qk2ycDdXq6JahAkCHxsrUjeoif/gHKMu/JT8V36mc9VaHVR624r88swlDTDqkbM
WFLpaVVDTbHuvNGlfu30ZAXaVsmttkDbrmZmkUXtjxhY5RHPohPhklG069BULA+ITxnfNqqeKwXp
decatkAp6XP1mO2uK30aqWjSrrANmPOuneIlMh/VA1v/5/J4bT2Oa5gm15jFkQl3l3ZCJP4uSONI
vyzHwfZ3tyfKcpOEfJuDwUgAvkpAqYVBxxdrDCbL5dPknNIfZvl1oqn2CbDjPyztLfGY1RQacWzD
p+hpoJlSBKco1q5ut3C8fdtuF8ePiLQj1/3XiDkQofrgKSKN84mLImi9LXtwRcTi24dXVSQL3eUo
vdFPmXtS4025QjWpdoiccoZsHAydJ1v6mH0zqnBglA4lPW5SN8MTs3VUnhXjs+WPtbf4U8I1Ofen
5z8h0Yxcns+zPP5+t1djGpAryLV0pyO0BEOnRhake/Pp1QsqevVQdgU4fj2iMpBQ1zOVsl5C1U4f
tcBT9AdUiP9QiKWatP3ji1K1eLfk5MzbOWBU9ZWNOaG7Y8M933oy1642+4JpXGOFY1XOJCYDvpTC
1i6TWnLitQnxtSh6cyatClkMeRH2lKOXystJKkO6cq5JgRLaRxQo+rlcRv6WU84n4f6e+2Shej5T
RQ6lWqjW3Gj0wulxhpunJ1IWlOvX6GBdfgzHjw8OA5infSSly1UjQtmswrkZ16NHVitirIA4UJES
AUYJcDvDj1HFsOqto/K1jjYvoGNXdiS00AWaeL0YUbmoKS/xfKRVROC2ow4SRdxMk1nqxUYDLBZw
q1etjNkeQGLdNeJFPzHfD34HqhTkthQAyBGkhyHSmYGX87pqhex2n8F9qWSCkRu2YPPNrWle8tk9
3l59bvJwD/jWP3OC24rB7SiaMPEsL3UbDUaW4aq20T9ldCGltQvca4NF5IUmRNyiXJ7swp+EWXmL
qsuBo5Y7eKEqyvBUgvai4uEos/Q0EY1OVUiBeQj8TYhUeDA+XmwqskgVQwyDlRCj1lDHqv3/+md5
e/v3n07/I7mryMRAy2uvy6FneXi1OoZHmF0EuyNF4zr5gjw2t+Y7ZmWukdt4Y//xo9yBrO0AgEQw
kvL5QYaerUGd9S58sZKQzepb7tKGkzKkgYffInC7VVTO8cv37DgzweoU8Fen4ThQiJmZpdJN45Oj
6qAtS1eCxrykta5pTUziu7X+hV6GTNc04FvOQ8B3wEtY+j1929vdcJuWinUO+0Z/BuG/LWRodwF6
QrgbErZ8tEPDMoZ8gP1NIcT1A2r3JIFtbDh8pdBLeYegiNnVOEg2MgPjQoUbtWpRbbQ3zPV0VQnY
LHLBnO2dAnShkBsWL2vDNDEkUZnTeD3X+dF3yxM5owUhy0HT4X10fIbrSGLyjasj4I/ap8hhCieH
2b0ClMahaUDHZpNAlXp1DANhxibGbCmzWVMe14iBq6snzMDh/5cr7b0KB+GPQHDZSUoZx6/83v1Z
047n00GZTGwhd0Gb7gS7PXmrrkXcK9Co1eGKOoImaokP1daKpup5YP7kA++PDKtb4i8j9xHd7J8t
CVzDKCgjTDllKNcQ1Cz+Ud4GdzfOrqX4WMJffjZ8PZmRpxr6XKkhtWlSTmlq1M5q20ba7XvoAD7c
gvQvDy2Vd3mahDHp64JO1O+LNbRZkmdmdX4uKWEI7N9+l2qG8CNoDoPH0fpez5SYNLniI3vggUyL
8KD936IO+OhmzTMGH8iH9YMA9PRT2RYfkM8zNkojyTzcRmYQrCIEjEik2Xc3AVXZ+FkpkVItBTsW
chGd6VRD1Jz8gf7uU6xC3pKAbSfFKJ5NWXyzp/MdzhjqICUNEfm2bwZTwKC8v3YhuyyU5CM5aOVb
ZB1kFs/UPTIWU7+fHsFShQw8Pnd0HsV3H9jBVh1dni3wDkRj7iIAbrU+wHuwCxhwI1abUM0EAjeU
g251SOnJBTBv8WpLxgqWPMtTXbyx3vuYnW4nVqHGCEULoUMJUScaWvF7FXuHfy66O75hpE9m64eb
lxf+jzoL+3+8SskD78/yH6uPTQjFBs+dJwq/2G3NKctr27oDUm8vwOh73KQbs7wn8lTnSlFz6JwD
iJCyym4qEkUw0X1GJ7tBWOI9xa1l54icecXOTdQSpWNtmcUR/0j6cbu0OL2mMxQxd9eLL1yzi+W5
HLLnm2i9kGm+buzhmqUPeNua/I9gsngFm/LFYeDMG1nPG9yib79sqyHyRfh9u0JXEE69+djgmLFp
k8Fpj8Q5/qwjg+pglryZGMzu0164oe7qYzjC098T21lN4pEQBFi9pW1QKHIMnESBf7TKLCABY46c
MyH/6MQ0En5tQzr/K7ve2b+eVOhQ/a8WmGXNnFM84y3YQqaQZxrkNKsyaQEYsLG0KHwhy0gnlo4F
soBXztls1gcWMKcqgDpmH3n1jPJdR5wd93xIVkCBOHKz7UKJU/Yf1rfw46/F+mMTmkE+RqPUPYSN
32Iqzq9KSjmGGs6Zgcs8bNBIe7UdrnzYFeT00jlu+ziAd8G13KV5s5r5e6JfLhTmR4he92mIkvP5
N3xgVXfdjNiHfN6Z/HzVbOwXoWJsMfdZNZyjiOyHw3kNInBhyymc/ztEBC26cxf12jp3P/IHTzum
sHpajVAwYg7aaSu6gGEI5oU2d+7wTVgqvzk1qZbXhQb0HypWOzSHVfZ6oU3/KMxmdbumFlXS/QY5
35yHpGWXKehM5/1IuoKdCFR4jo9ZW1epcCqIoi5UNF8yzDYIPkKdLUqoAyi8exdQ0pdqEVPS5/Cz
1SUmfPZHCMCalkmhbTYDrC8yVMzjBA6GY0HcRm0QBS/i3gRBIrfAavIrwON43n7VeuVDgSyPJF6z
XmotWp55KIbV9tAyq4Oy+ytXv9ru2yPUkgtsiVmI4je6C9+NdSynud5NBIzavjSeCE98GaiLD4sC
4YQ0Uaz5GEC0fHW040/n/j6SQF4Afy4GYvu2mKUm7bfMhDN+rcixQq5mCouEQqnbUZ2J50Rolr9H
QIT4kG8dV2499OTPqpfWykzUj9UBQ/2DsXLtfqKkbB624lsS2FKlXtYuQLgMp5VT7my9SJ480lmR
pGZZ2NBJsUQp3x76UVT8PKPR8SQR3y5jB45S9zodGH6HjCIHl+wtMR3S/smUqI9EokEr/p/a6Byy
n/zbL63V3g2L/dBJAOKml00DU9/OwLGypaDp3slYiazooGJ/huJSPOt42Ysnve+o9kR2Yxflhgp/
oUVFzb+Oj+z7zRlwmipGUAPH/TILZqBnKK9TNX1c1Q2A1kvqcYA7jDfEBxOhmSHZOjoHmBPKt5mg
lnxCyj/eEENLQEQsTUlvo9/Ii56UgsCLzhAfqjeYXQ/EKRj2OLlIh1W+3sgWuEsMFJzBPCLGg6g8
wXVwZ+OZ/uVbLClEZ6sdMxBZaayvUpG3bbyLXX8eWbMAIcMV9nHzjHe1twqSQznXzAByr+wO/fr2
BEP8tLa+8oB+gFnOwT9avrdV6sruhv+9vrR1crbrkameHoT9wxHFvedojJVcZS1fxs9mZuOBbTo0
75RoUfCFRnGE8zQUyKZEnrHWrlMS4uysRi6eJQIzCyD2Jp79KHKgzFntQiFSZ+2Y1e2bECOj+7+6
kIYX5/6vzmIL/BhktQ0x2b0j9sOaES2LhgHON5Pq8s3gEmn2tZq8nwDCo67uCqnCIaskv7NyBS6Y
wQ2qzJXSVYx0ZYvDHsDS0sIEVm0Gu1OCjuuJ9izWHvOtRwO9WbTipJUmYPUtWS+HTy5GhIXYXFaW
omB+6drra2DA7kP53ivlougM95Ny+fZuiUMNdi17OIcqKNFz+cUNtXpuW20npwJWQjxgiMsMksHc
31RML9yv+zCiVki9rGAwN/h7366IK3MBbx0nmajappS7Wf9RaPLre5ghidPnoOoPHwxb9wcWQ5oa
P4xgP5Q2ieIuD5tSHvhzyAh/S4VBxL1HTBLF4HOp+h/8NOr3iKMe17DAzCCCDQl5FrIQgVYC0tzV
saNwispoxxscqg2l7WbZ6b0cE+KGb/xjk3RDMGVsOFWOpFQIRv1Mr+nFXV6AsK/Jk0tyotn/RGHl
+2ckBkVc8JCXbHdD/We+hUBj63RuIfw9OL/UrybNZv73ajeILEUNSKh+mTIERvpDCfxe07DmpwDP
ArteunLY9fVyMciUE7EvjRkixdc1GPnGQUNtQQazG24ajT3BWysEXFtzSy86Ri7dDCpn9HuzVS27
gak6rs8M8OG6DVqWLtE5ontOspcM/CwCWVATiQ/5ILBcj3u5ZNNhTOGsbeUSxc0+b309YZanleJK
3T8GUmVZqhUwIyv4IpyQimyOd9RQNVbjksV0XIaunHKqAmSujK1Cda8vgMklbK8YK/QAFdNbn0Vn
hmnzrZIh+1AFods5G8zS+2xpr7914gJ9TSc0YKAsFyV/CvIHpdx0xSbmneCZDJgSjxNVaszU3bgV
Pui2OSV8PBDH4PbfGQoo+Avk25H+g3YS13fdboZMmuRfCIjRDQFXfMJ+3NIAX/CVuzDUqJSj1PG9
tR1Bzm/VqcGJcsJeUFeSIy1+AKOGY4QMno0xmKmNnC1oWnyThC6R1WnaEBXirFjDJcVWbHFbSC/V
tex0hJujiHB/f6eG7EPZX+5AkgP1kuuzOR+9IRR7/qt4WL0B2yloOUt94xdlVkYVz5+6TOZNGmuC
FIvt4+6pOxDoJ0lCGbVMnjMXEWMl7FyyGOxo5dC6+nPfHW23vfc92zzypnx4uk1MosdhnE23t+TP
EKy2octm0jv+ScmvDEqknRPOeV/8RKCgie/C2+MKNT3WnJK0eJFn0Zxa6XJQ6aq61vIwJxwXYqaD
QKCfGLLNnYHo2cEkqvgcfV480M8/iSU9qK+ryitEdxTPbNSbskVLLvOhFOEf/sQAFsh+v56EZZdX
S/OCIp7PLJ85CRMcK8oZ1iBn38lCAO79Pt9zj7mDWJ3Jrb+tAjn+Tpi0EAGOX7BrHDLmJWEVZaOy
cVgCCvs0nwMI5E+I4JLKcmBCoUxSmuxSR3AtNK7SP6fNd/B/bUDDWMfuJnfHED4ks5r4E3uNhJjN
DqN6g2MzxEAyLDEC5VKCVhGNqJ1YviITjefE7NFzNR7EabmBJDhK+/gHoY8wa9NXtdrc5DUg442a
0YK2hfRBxDQUQ/dw7n4V1EX6Gqo3VNxfgwd5aozpUTBBrfbjXXp1ZXe3KadzUMvQYLypc4B9B3vm
iVaDuff4mK6DA1efceQgvOSr93pCsIJfkWCNQ9Z3/oe+J8izXYcSeG3yDmR6NOoXzDEiZj6beXG1
HCT4VfOHXt5jOT3KZhVi211T09mjf9pM3wHtITyn4TShY/XTw0U4+H0EuTU6wNvCOlOwOhXc5LmB
eK9e0caBRb4ljIWIURaKtCKVe72bRy3DNR4nvBKOjnTjYx21Yw6XhNsIwTiH3ATf2SQmDHb4Av2t
irkbJYVT24gXLg8E3r2uye6Nco07tNxeS2hF0cufjIGDGi2LKujU6XkbTUb2caYqfioZAH59gwmM
jp7vw8R+Q5w4ehaL0z3aj8PlBNSLnqO/MyfgZBqljmSbHO7vpzBp/HrlJbdEFbvRz21/c8iuOfs1
8/u3XbEGrkDjgFzKZHLH80CfMUu+4A7hxk3Jul4LBLiaWGm2A80PJ3uixh8Mc8x3fCN2/uuaop6D
hbNDJCSc/oZq4wgjKvqBxtrR2Hzz/Csg3qSKy1weOhGtSzKBNneJVncBnIDOmDqeLh6GILb3yKzs
HQz/iN9KXFWX5xqJkgPJzfrcjPobfk0gKHyDQZzXHAW9Z+5Y06RbLFdXEocapQWGVWNra+KiTQ6H
JUBqzsU/mD/CjrjEQXXc5RYRkDb18Wj8jOvpp9FKB9U51wBHT06kxW2EaKFa3H5jCAbf9zW0QIx5
Oo1G99r+1yIcoCXhHY95eajSxRUhRRHqEHHX7jMJabY/W6suq+8kVUX09+Xq1isJjeA+upXVu11P
h1e+5V+YEVfsK/TKVTEO3lJqXZ6ZvhP9iya4tsfJf7zpwSjrk+ddSlmaXQGG0+CuF4Ys0KXuEizn
XL5IV502htkjGyKGT+kg2euJ+a7PBb6jveshNPvMHSuxfr2tWFwVPPMFl2uqQVaV48pc0NIW7sJ9
NDUg+PZ8EAzbFzkkUjsjdEdqEklJfcHu407/4aeiiwmzQ5NKwffmuJ6vM5CugXexfchruyvR5+1n
+B6CW0kfS+FKnwi/jpjdTKQyNcMZavDOlx1/bcMQzLCTbi2NA4hnCA9PVre+BmySyZ0MKXJNHXRi
kd1biCzxF7oDOafJoq84PIs2yhwRxvu5I+hrlXMzGyjJrkmnYbzwj1+0bK+fkY1YVFBdwM+50ia7
+aNotwR1tpvXHGD4YqgktNzi5r1MCdCLSCUAsS2NMCuGs+A/27BWBsDLP+DDZ94kvVOwA8eTPsRb
2g0JUu6U3HV2iuAuMkOEZTGrW2lTxos8MQ/gns5ByBOtm9PPTGqr8TlK7YVBRJ8y7kBuwMTpR8GW
s1lA6dTPdwO5l1ai2CdUQ811oY8970FhAB6rwnHjrWKePfQuEfMgGIricKzsksnvNJ1xT2qAbbUB
oyt4DmujrdU7o58ALpzfkZRuD7y7MqX3ItTSrOEsZZd4mvHJnEYCcM6UDnftRrFBARpzpvxUn06x
Rc0zoc7BxBKgXmAPxCMiUrIui46w81wn/tfQk3APkd+WExfcBWxmgzAjP/HHFqIuJ6Qs56flHy92
Flop1Ph4PcAFyxweuPw5Wh2xXRyxv8IgqB4fuE3u27jZ4NG4zaWX7iaftnDU1lj4Bw4VTgGpm1g4
YnsSNk39nvmumecWfZCQAijpxNO51QgV9yiG7Ciig3H2P5KbVId7MFtcgVatsqHJCnuw6jhCwymK
PJiFWHJBWJdyRvc/klz1QLg7hLVtTA9MxPP10UKTQR04SlMHvgZalOj6BFzqYOsf0eRex29ElKLL
/SETQkbvaCQh99/uNBRz6Clw76753vV3O4zzs61qXyNjJZaTdntDRllQvrop/4g07QJn14FfvQ6l
x7Q2qLT5379Jqj7i/Jabj3Z5NxAZOLslymQjIioWSL9xDHLETt+/oZGNJT4/dGOiyKp31W2xZpTD
a9nbuSkjB6M6syucgDNoilsBcCGhsjVES/EB+E7FgO/ZlSsYHoYFWO5SIEe2V03X6fU9rBXrJYQn
RjTNx2xqIZ7ygxxwCmXLbzqK6gII6GjIyc9AdM13AhDX+XCuQrnIsAiQ2pfGSZm0c69bYTgyFkSS
6OeeEllBLKlzqiI7H2K9NDuPC/7it0Ke79t34cp9hy3FXdMcwIyAtJ2Y5IWNFHU/58YQ1Fh7sVGH
4K6Yq2DSapi3c+e+KPd/8Rt8Bk43uwR/5mG8q4vKg0i6KcrHqE3NVPPJ9N5ZDN2NxU5uHXRxNsDy
IzTleKCSOQjxj0cXxq2Rd64XbqIYD0w7O9t6mbf8Y6Lk9HRCkJVZ0iMdqH9kFFMiyfOdw0lVZcz2
Bf8DcRdMiVp1BQCn6oktY/9C+lsTyJ6zPs+pJZOKeSBed8S+VEDoAr9/Jmzv3Z7Uf/tIAOOTukSR
EoIy07ixRAcFoDhNt3y+ta3pMoO9iIyzfZkxSMl+sa/9ujLl/uPj9HXZpqKIW1V1+PoWc8dR/Qby
S8Uv81QKUQs9hHxf2BOcyYw/c7bLIIuxzQm3BUUea46n3kfuF/IUX4He0gYj7aiQqVx3XXh5y2Kz
f5MncI71M3/eoE47t6c7fhR9X8+eKtzRW7e13BYwYIEVJPOXmI7e6c1mHW76sjjaPXvgBFqg5D6b
/j7LDzv5+fuh/xL97uCJvyM696AUFuVEk/qEg8SjtSQEJ3CsmlL0GED+jwj2PByQV0+Wkd0HRFbn
FcZf6gNv28ClMQ9f+rQC8VU8ScUJpmk5fbp/LS4j2kJ2x+mqpAFu9K3FEy941h8TMDG1vFsw/Ygs
ZoqSH/FNGXiprCR6e/VXVvfxVpHN/0s5VXxaZfyhGQkcKRFMQyWHLJl5vmEhKcs5hU8EtGzc6GXM
5RA+IdWnAwCeYBAxj9raBpoRJBuI58ysU+wvYuKz5uziGmmzTxVt4nBOk31n2uTwwYVHJ0KvTto3
lu0U7WYgCGxmu0vFfNDtrbzsJARnY8TnVfgoKEBLB6yd9JNHjZjAbD/a3xJv3f4h9yfz0YOyFczb
B6OzJHDGy1hLHgH8wVTF97ni7b+PoUY6wfuXoAJwmxgPHq5IeGYdd2KP6frLJEqI4xZ+2l+/4sT4
tH0tYS7y2pjNiQoe7GUrr80YTpydZ72K71dwhmCK9ZuAnNncXcNpQ7kiiwKq5rQA5JFkPKXHuvF3
Zo7R15u1hniji4e7sgX+Ki+6jXRBn+XVNFWDyKjNAAZ+ya3hSSLUqnVCoO4j0mq++qy6bXhA32y7
Y0wJzI2gwp49uIpa5np+lz9Tbw5FNaW44I0jM3dkp53uVZuSgWbc2WFHYixBXsoxkWEfsje+4w+d
IgrwKjiD6g8tSa7e7zmDgzbWOxgSTdXKHruTo9rvG+sJ5+bwpP0x004XNswBjbEHt6/31PCWOhb9
7CYIvBNRVW3pkDAukzyyT5Xo7xtTy7916lLWmvognzpUhJoBifmMC70z51118v20S1sLj2Moa/2g
CZCB8+OPRZtVtm65F2lviXryApBXwKL0pQT+RLQa6xZ5P/7swcT9f5Fw3x6r+wxjtlXx0wl/OZng
4eXuymDspxVO/dVvQU/jyKxcB2lU/E4MfgxtmyktC9gq+DLggitD0DwrYFHkOko1nQNbPV182dhH
GZERY/8ulUNiy0jB8spwqYR947MvoDlqp37tQqiyi4kI6bdAghq4f1yjGiBkn5lOzTmCrbJ/PqJC
vLKn/WZRjn384ideiQ95aSHCCDDaJ9kOsb1gbSSRhrKGXq9EzXZ0JxVkgKHxdr+s7wbClSf+d2AS
40WN5X1goAPqh3T8tCf67h/foJ5+yHQwRW1Z+P3zH1S9pHFoud93sIlJNgiX0JEdC7Ngx8l/jd32
tkIqr6OGLFUbkygZowxxianrkHBpVfWrI0ocf6UIwgdQX84Y0gogYjJO4ber6NUcAclAg992X9qh
miZFAbeuSlJBPNCPvXGjc8D8uhfsGha4EfwF21Cx/YdvPfvIjuRDcR1LiykOx5HMWSRqRXs9OX7g
4zUVqTxGRZSMeXLlEiNrbCDILvrP1gEBiEzAqQCaRaCeXXUNOdEb1I/g9iYDQIm3wmWKmiduv03y
/q1oF1YNJj7wDReiZpBdKf4iu+q/EPabxfMIvuoNgRmZTyTr9jP8UL+hus51vYD5eMPmFl2EofgC
Vz0/p9sAw5fiGTEnb346KIfx7l23gDmFZNENYnCobeg5f27aGRBFP8VacgjpQEnqN2FWyJTs5cWu
Yt2YUQdLMdk730HEugwLED3YnYTjLRW8H+H4aTGMr/VxqhrUX0uezfhk3W1PC/Z3rLk/CmZkpahj
VADzQed4n/xJyIBiOahFJyD3xZuFDfeRaGkAt6LfYT1YpGIX/W2stF/UJEZaeH3AaPsIIasbBc+t
36s/aPguu/mIx+zKDpdlrbbwy9UPvq/1NL3NzMrO5M0v9OGsaPz3CShuvZI6x7gqeC0vPGyYJU7M
Lb1u2olUYlw5PDzUEvYv/Sn7mWRuqZEsUNHnjQFuJ2HfnTvkMFInxKUi5MPa5vgGCDdf9bAlu5XQ
vI1Q9vamSMUDFRnoxX7b0x00+oZEVMUOfrO76XXd58gcoq7rxTWHtdtdm6is0CLHzMDhf3rzESqq
TyDJkhy3qrfSb+BkwJnwornc0WDmKr2zYYsQYdKFL4bqfayEQEBZa1lDlcbkdj1u3IfptFbKC/BE
MAColx/OX5wZKIuLSa9VoBEvSwLMxBjzqUBdqiuEh1KphIjfl0KUblK1mqT++uquBSykLIXkmLfy
m3r9r5MmeaKi6HysnwWsmCTBfjuFDamsfuAkZhhfD889qkjiRoiQPzvrW32xWom9+sOp77uPtDBa
xLS0Th3lZkoTl0RqjaocHjuJwdCQNUtXtBZsdLlwg17AUmjMdRtbO1Rab8NBUW+tSKzGWQ3OpEpd
wzmpT8PSsbmuBzS5h1rI0X5DRph6UcwOGDdyUSI7+BOtdFyl2XvM76BX4bgjq1jrce/7DbJ+uwnA
ir1fabXaQoBv2N2EzdVIsFE/VXRSRHaMjrb5p5ww1g1rZzJyUsfbRTuedRDUIf0FVKf2IBHuiqqk
Y5xD49Qzx+zcemKbsn6FU+VRGOXdvOh7nMWD5x1ZeJk8/35SVV64e6avE2lfDOoMonn2+M8d+7eX
gnnRLwaviJwsDq90QDuIGKCfGJ7XtdXRfCnZyyGJ/1ywL6FFnQGIVdYdqHcUfC4UeOl0myC6TdnG
L5ObMG/dNwiiHSUp3bjdzqliJ+XqBfBpRUmslOc1x4Us6dch8oygI/8C0ZnLViqyFTCF7ygsM/JX
WenrJPS4kBcE/lKYwtDQKe0qtMstoZO3HEVqatlhSQMX8AUb4BnHhHVKKzi8E+EyGEU/RQXr2fH/
JcVeAlUE73b38tJEHEzFowKb1t9imBUBq8xCMG8t7LtydMIDL2yv7omSDaaeJDn21Xk3ANPwrGAv
+H4zSQ/agbAUqWVAJ2Ayiapb56Iwi/QSdC2Bsgz0pBK5G4YRSYz4poCAcikLfpS5Uavg1vIbs0vS
W25zEkBS7LqGf8ePJ6rVhQ7veFtPpBwRuZQSvkEZ3H/eXDUhOLreS6H13VJsxwXLoh9Y1Ktvxp6I
z3bU+rlFguO9izHfoQ9gAAdV/tZzSvKuowF/vVO/SSy+Z5h4hItweRYx/Sm2pHm/QM96EuhNwNvd
+GjNNkc3dATIo1OUtooYPVn67lhlIdDjZqK4xKzC5bveOkC1NjnAFPcSL7Wg7Mmzm+jj3tZd4fyt
bfIY1R2pQrFTbn9aBQAn3Fo+fiSytDTCxH8lra7tjJd+uIQR3AlSPxsps6Muu5SEQoNja1XApS8I
jzWA7zzVBpMh9Lu7e4AedjOTyes2s0T2uymdPULHbzbOIVZ7uNcuo4a4wj56jG3k0+PPfmbRpUHj
QCJ4rbKYwsYyKslBegyfVVTwOvIkkL67CwgXsdmH2VPZRT0Q1Vt2xDrTfGUd/ALU5uHa95b7p+b5
yQoqC3uc5OJ8VtOfDHX7n5cW6/Ral+RDQH8OlmKewu0dKy2kPBvMLPJ/lyHAEfk2poVzqhQY2O+h
KboAONITLSDobnXOh5JJ1WqlKFln6/bhHKovHC94fXkV8gr/0wdF+p6mn3rks8Zf1pAoTwn+qzGF
j466mfQjvpI0oX3tPHCXMy6wCfRLSkeGbE6/0sZpJXu1RjxmUgGd1HdRyaqO0U7f2qeF4ke521nJ
A7eV1JskX0yUpcrV/bLAXmzL7JCUYPpPDD828HUa6N0yNQzlBQlbQq1+G1lwQcLqoFgoYKB0EY+k
k0Ud+oiOIsvUENB2fQeCteqSC4xgiOhz15oKBBZwhg3XDYOMdtCAkuD9sAUPwhBCrbTAlDFgFERY
llyE368xYBTqRsSHEbVIu8oPra61PPsAyTrYzv5oaubgWBOiisDTnI7ng+xHl0RTDgi9vV3lTbWL
0Ke2+KAEoCemsKAIATMwyXD1aDC2BOd+thHG1keGJqb+6XKrcCuPzKU7E5AMjknm1/ItUg3MGt8h
HgpBTQ/dTSANM+qnvTGl+m+glfPn4jsZ0D0blHDhx1gQgseBrLpWJnaWAjfTBvAiCm7pTFLvvhhD
KUT/YzimMeNouJpSYob+7yhiqFoAFnTS13ta56dmrtBoP/9h/b3do5XzhDe/sakzZIv2lWworZ+Z
7Zo6qmgrP5DFuC8flHqYCC2wD+UwY4UkHCvHwaNFc6nkl0qtJzwbs2ET+Ylzc5yXxhaU0wJAyH+d
mwU+LlfA3posiFNn8h3RV/hCGauqNoA861Pc4fE9YWseumCViiE7+ohHXN7eGGvZOFOxFksS0HkS
96jjMxETmWYKaJth3W+GDV/2K20WmlYjwbW/4LrczDOpazlSsD0cE5K2PrdA8zgiCCyjMFrzWg/v
R39E709WicPgclwkZWpayDo0PDDY/5O+KaR7+6L4XODSooYYTy00T4GvppWs+Ji/GKnCqCVDlGyr
tCAhM9oKJFTKVpVmfrlukkxotpzH38AcfN9iJ9qNyS4Ycm9/bwVWD1nVq+lHylCSHlG9oQSmIeD6
+Lzd89YYB7THiKU8gJuDsL6muovW2pg5Z6PHCessoPFmZbN33GEoRl74gKTjM9CfvVOScc7Hseiy
nGARFqRMIqu1ueWM1nCil5MgwHcBvSU57FBFqY7gWwlZFjTw4jEwsEjGWUz/vC1lQOF07wALVDeH
ani9IpvUKk8yFCQvHl84bKapynK/0E9G8CJHFx97zPrStaP3HW1NM45vIBd6gOJw4msgfE6+DLvf
AnPf49WJVViXPmTjmJHEl4iH5kdhGhFG0JoGNsdXmQCjEDx7OLv+scgS5fddJ7wwuR2ssCINW9jW
c1FO58lnaYt6wSVXhKXcb2seF9hayaQL1KugNC44hDc3snnZ3tkOqSL3thkHA8VNlgBbgEyCqV0a
kH8H1bGFRqpjIzJQnYA2QYdanzgcvGhYZMnm9tO2lIRdMyMy6mn3Mxn9EmO3XWKnChG9u5214H7m
P6X3gteU2x6vbS+uo6Y/5TXOau5t/BTcJnlMR8k3QpF8rFxlzxlrTbKI2CVHffd9/g1VyHo7Nzq/
Jb2pS/fehLsaw4H09zVE75I46r+FqPwCD83jhezpSYxTcJ6W8A1vdzxkrhBhaxtBodW00jz0CDR3
OFPVmvWLimod0ZD0ACE3qdRhKEV+s6Xtt4Fn5QusESVxoeWo+2OBJ0K2pjdxA9jnm5k/WcmiXyQh
lzvBKfGdMDBHrshSY/EydQvEUA1ZoFVVIxkUog/V2FjtVXmlj1m6h0QQjmtEopnfL+OLGbpH2oS1
yeSCmvUK1JrPoE4V4Q7Uaxo1YkFs5MkTir1/36uG4u2bCtRMh3ZnqCR554YnODiPZacIuFlMuyKA
c7klGBZLzD6nYfhMPGliICQ/peLzgAewp3PV5t9VbSL6oJrjpoGJsoXpl2LW4QBPr4bnacLsyBrX
6lrml03qzOWpyUSPaB+sCATpN4eEm7CnHXAZuhk8swvveoG3BbzB85kaVrXw035pWe5m6FBnxtW5
IxyzW2eEwF7y5i8ujIE57AMe4Ky0+HgL9NRD6pxGjgIkNiQf3rorKAD1VLNdlRUd2Q7XbfNttkEE
aAGUpvlbNMC/Y+rc+BVDoyiOk63x3LK9CyKLWhyXkVce/4w0e8qYtf6IUiuhFkrgz5/An23GnXdr
7qwQpXRWvBIXf+gUmikyWa5NsuQrKbXYXmaE2YpdsOrumlULyrlzxsVR2kU4gguNNDl4pbT82pge
28QOsTGiOY5VTVedXEM2mc1y7zSH2/GbRHXAJFGwrg1idUXsQdvRriVBW7GhSvT/1i2JIiYG/rfE
UFp2k71Y8HRJiZJo5sXAA3uWo9il6Rcp8vGGTCCRVz08p3paSi6SV6f8Yue8AHfVXfGbVPTqpLlH
gypblSPCV9A65HQn/je2RHcGxc0toJ8yecFH3WFRs5iMnfM8PJYjxfIueuSyppBtFnjskMKVPyKz
TMoXEFARCnYzHnXDwah09qzZyILudDw4arccLmTjoaHhJQPpf5/RntjLK+vwF2SJ0ne1YuBmi/V3
tjLIxeKzj6uJOjHCJYqFHkREFt5nsH5VaI9U5h4eEZeMtrzE+oPjSS5/N7ug1d68lsp5PfRPSxbO
9JgLLqqAZJ/8+khwPeOETP62S5lRsqUfi+84dHofXqTKyN+KJ106Cy4JshaD5aBwmZiGROYCbXz/
LCdT5+/B3MSTCQxMjk2bZDrmt9vxfJOEC8q8Iyh6H+d6Akiv8KZs4Qk4NaGU3HI2Y5E7Qki7PKa4
9ezVJVeuzyLgr3/DGhstjgQukzKNhJKtmqFZANeXsi98cRoULqf+cQaQFiBFDDUquu4a2vTCmKlJ
fqw9Uo9qGoGHcdWrt3ECDa/CPaB49u74Bi+wJcpA/niWZKaJHhUR0m4z8uPQUf72NAZsBz7g3BB2
DAGTbVwgYHxfZOJV4wlEELt8fcp+bAcmMJ7jOupKjgqtIxvFP/C8GIT5+fGj8veB9zDyhFRNLbB5
YDw/05dm18L4QpdzGEItzah+mHTKmIntFHEtkPAuMzl8sYhQReeSBS8LlWyGKPlsyspYrpagYrTp
hwitrtXNpAodFjwYb79HXzyilRyzxbZdAsE9afI0rRMuXYx+Upy6s08Zl8tI7YULXQRsracekFdr
Zsl0RE6g4MjgQRTJ1JoF/W88aoJkl3xW+aMfYSHD0zmAOVlUTSKfDyy+4c7GJ7H+JUqO0iehP/uM
iGpaxeWxrttVD+MqPf0qiOWsPRZq+QmMxUBn9OPVuwCKxDPRg/Ip94UEiWEVjwFPOXTJ8NG12Ebl
UL558t5HlBpUb5akRDMNIdSpp+oWKHGtpTl64jEo8gTDFLH9+bSDGKJzDmjWex28/NRcA5XNDwOY
6k+NbJUtSkl3qQDRSImUD10fRqjM9cvydd2kkaR+97OKNl7S+hDQHPrvfWFO4hHMBcpoGgT+a6CZ
9Cj/+KUptx0DdIBYoMPvxNBtdygqJ71vGLsCNt+wPXjTq39DSo0dCoOql3OoHtZXhlTLiZswv92u
4cEi6w+4caqLyJRrK8prBB/QjkB/jRE3rpBOhd55lmUQpJDeweLRNw8PuHP4dSaBiiv80JMt62K/
CpyvZnjG/P6GW93tiAgP7WXwDEtcUKn/REvzDcfIygh0y+/m6GDrNK+fz2x2cveQrkUMxoVWTnHW
lx8ay/7CT8zmfda+LNGg/u2h3mSHhOMbFFO8cQ9HRYeMUyV5rylBZQmwNNuPmPC5cEuQwUfSDyAo
ade+/CajxUZ6UIjNpHq//6lqeyuKS0NvB/X22RadkLHwGuUbih6LPHTh32fuOcW3tZes0PQ4wc+U
q5m2Q1+bJ0FgkuAAZg9b49Pz7+aXmDeupGEHUanmz61FUJoeBwQp3EnxVczEL7RW3W2RbiYZe93K
8NiA6FegfQXkW/mu5gZQx1Eh06Ke900ZGdtPoWMEWmmz/rWQwNDXWw3+mB5EGElfj5TlYQVZOVg/
pmi+WdiJMKxKZNsmIDM9ZN//cD5UCp1oIOzaGX0Scv8kDGuHFsCv+fpGewxOsQ63zC67Ah4oMcbc
lslL7MOAgh9TDQYeN2mJSJEwWnk5+Yi352UrHMfajUYwUMSh8KVBrIUfVAcrlHnVovvRIk1731KD
ZfuSUZhZS/wR3R+vw7ISoeoqfBNcTbQjsdI24Xbp72zuXYvKZ8DSsP9dYCLpFwR6pwiA/D19FV8G
A2pLomIgpBQWFds8jLlpE9A2mKjoun6UuNYlGu6oaJq8512cRVKnQmE4x7X+9xIikz8yhIMNst+c
bpKKMCqCwqzSdV+Kn1hg/YXjIOZ8VAzOW1DoNSC51vtrFptIwrRkvmLf/wYp4iaGpE78bgNqIysJ
RaN+y/WW9BRheOj4snl7sXHqDGZ7MXX7hVjI4eaVDdPRufZybu1RWoYYgsB7Ts7izI9kIV/5ZZEa
D1wxp4yYGIG4Fm3UPIvDm1NbDVTrv8kh155vsprfu2rpLE6Xgat+p1Q7ruxPdAYyb/cj8mJGDtGy
OwyusPUquWOluU0IF/pLAl6F0PSesrVVcjcnAz54dtgsguKkwBNC7vDVmm7RSwJuZJ6Y1Fmp7RNQ
UDAjgjwBY6jgYm412CnnHkEfbpi9ed/3Vt02ZkYAgykG8CGvNrTQh/JRmc33DcV9GHL2QoOn5h0s
kTYwjKNqFiIIiWAzkN6700ajcGDtqTMbaHYiJHGE0+QLbk2KlGgYIzx3bSKGDYAG3cXdipLgRmOU
h5LOcbJnel+HvbKMjYUMtf/kPmH8TPcbIVsf3ETcbGIQDJs1f9iSXNciD8/DEKFeMnDKWrCy/RjP
GdJH6TdRgJdnS5qw+7ZLdMyxbmyKVAAknH6LwVcAKOoD0n/3I66O/cS3tzH+WXw1jqAFaxODY5nz
mZNhKhER5LHNhf4kWhgxZ9GB91751PnT4j4Pjyyvcv9fdyFGA5qUkVGJTDvhq865xTZt8XI1dbqW
Oohd1AQpcBGRcX88UztGLTNGNhkawMMO3xWe2yXua3n/NN5djjOGBOdmSDalQMD08R3TYarAPEYu
13bDhC5s2rQH+bbuMW6Anevsg149ZJmIhlGhVTmTh3CvJAvMNQHxz9ECqRPBaS4j7p6abH4QzZZn
W1Hj9yTl6TnRGIy0NiRkRCpQptXU4QenLt72yYt9HHuzgiK/Nr2/2X6pBGrNy+IWVF4kSsgF0uSU
dkYMS7hcqXPQ4MZVaul8btyAGcvCpJStjy6+IP6mwWwN+a1z+Uwvlaj0mW8t7D+HAKZBnFX+iTnM
UKWLQA/R6eDgC1sE6KCuX6EFRBcrNMiecn+nm1E4UXRUgsmq9PoesoSERSnKwVLGjbbHeWGcbl7Z
a/NpflkFF+i6CTiz7Ro5KZAKb1hGDSirEJvsmCUnHMOVLR5L+0B3aHJsgISWrYjMsPomG6lNccvm
o2ryDvEgOsEj2fUC/xij3Zm3PJ+pGXX0GsSruFXkUpPQODgctmXmImFU0a6Z40ODvzzC9pUdVNvZ
dm4szzHVrnLBYbrufITg9LOBHFQOb8gwHxyYHx6mvEPBXSk2TeaL81HEW3AlxnWOlxmMdX9GYR2K
VBfla9Fn6G+GFY02IIu2lOZ1IfiNKaQgXiWA2ZdwG1HJDZldOnYYZ7zyvqWFuy+gUA7vZzxmzPOp
ngXW6PGe2JMDcjgX5Ep81a/QZZqwqMSk1v2ccXwG2C/KCCSlDyPuxTEfL0NOqvILnkCtosbsDZKE
V2ALrlVp9CLc7aE/9CgexwrgoqSpPJhIv3GA6WH31HiKzWjRA8SjO/WoZZwxowZQUEZDp4ZV+6aP
K5fNpHUkS9WUgSMTnnLBK9IZERe6UiLImWWr39dC52XG8BVUWIeolwimObq/bKmbP+UA+kBON77F
85J92J7CiYQTMgiGwQInbuMIhUCHgTCAMse2xNeVVWHKvaMpS47bOGLI7Mjv+oJVlO55jBCwWi+C
ifnBA+dLQiZWQt5xpnKcEoxG7my9TWig0rvAd9r4m1RjXLXcAqW2JclvYJCxauiJmhOftHFpguTc
vwCVKzfiFPn0wog0jMu7BGuMIr54qrmakcdcOboRa/5GY+OOqvJ+s+tsT46MxoktCJ1+/f8OGmun
ZCUaZXWM2WsNcgiblflUy5VWOBoBMi9Vle6IUyENQlfEKQ1bKKScv+7efETnP9seCqRh/Bc4wiVG
SodgABddK/KnR4riao2NgnhOAEXPKkX3Ct+9ZPyHt3eT9Z7liNmMgiRfpJhvWGK4A7+MPylCNeQd
OOb2m4grQuqjB08wlVs5OtckwPUFFU8RvIJgB+rkLmNfApH9pnxiux+CihEX4Smrb0zSPMzw1yHi
PHVKC8OT/jKP1BxsGFQ8sNi7FuDP/TsU/lQuoxkCldzCFzxkFrrFD1DfEYDKW1ua21K21PqkBwMf
FrcUwtgG3BbgePcu/pOAbtZm6n4acHjhxSId97cOwXU7kuMRmN1+I6X9pW61HjwxEVaVwPW66rBw
pxaXpOdIWGHBdUCNGzPEhe9RxRMymMpNbvEWtIIFmJ8t51k7uWHo4yavQDhbdepNvnzYbUv1vYHy
GHrtzh+um6HuHtYR4CFXtRoua/S8bGePtwW9N8Idqu83moO0Sw2q7PudjCU6l4UB/ngbBAvLNC2L
uINVkugL52rJUoOaegQUelINLKAq9lSyVi90ZDyF+I9eot0ptK9sMgg0kViRN7uRH2bQnf5lE89Y
hiswNaeiH5ikyL7J7T39wBlStQnybe2yGJBDc6nabcKpUenqL0ILOOFmpnq92gba91hlS0J7UCU+
PfwoesoQ3iuHRj0L+5NEGVYXyNG8vj/2us/wH6pPi+zeIGHzgxjCN4h9QadPUBr9v0BPQwLc5t9M
NKiPYgrjSzHN0RKdryVN2kSGcqh1xe3IQqWj2cPjT68xocCuc5W+BUBN2umynjaw/A6/1cAFgz7W
UY436C+kvlrCcRnJOveOXAZhfB6l7czghknFo4Om2VuXWA1GKDwPdFR4lio5wyuzP2N0EXCg12cI
fsamSsb64XNxtTBIRt7slWh+nqsBgfCraMpbjFyAHrdbpDucjGHKupQnrk2myuZj+/r805OzzQgq
D4JhKmWiLTRKFEubOUocS1jYPC980yCClS4AMF8fQpUy413c/fvXZt/alzWqN4anz/nZG2VEJCLO
rl+fWc1CM9sbB3qnYIPGan8Bgfljqf3CTC1C5A5dqZuc6S+wJKYJXGC6VR1aQEOZcIl3be3b1NHS
2Qc+bElPTTCdWFYr5HeHZz4QHjL6gJQaAKtY9qz7BDrjgsCwPeTgyQWDUS9k5b4Nk1Rveyr1zrgX
Q1TDCAkbr+b+g4S81YmpjVVQFSNATf5Fg4j+M68Nkp6G+XN/ArrqnZ5YPB4PsZearY4CzFjk+QJ3
HYksnXtrc+mKR9JC4a2KT+QS8DdCSSwL/SZiPvOeXjHV+OFS9nfiSSFzB8mEGiuzpe+8Wcbq4jK2
4VHq9TSxCP9uU+QkVFwxcpoLUFrwpJCod+ZtgjVHTczEpKsM08PL3byfbJbq3IVX3t3BpHzfKcHd
MrWau/af1wR4ov+JgW4FGhQT+Luas8eitOo6IewDFqWjsU3boXhYg0aaSrFSTvyRSEzVE1lOvNUg
RRXOsJCiF3uNi+83zxmhVdfcH3Vw2tS8YY09eQEtrCcd1aFrc/TuOTq/Lh2tfUQQoaFEj2LBs4Rj
9C9f5TBt8YykME5bOiDnb8U52WobfLobeiapoj8JtZYyZACLs8CJbytyBCcWq+orA0+XuAckjaRF
24VGf+5EuW48jtL+d7vt9M20q6ReFBZKbhQWlmVAz7sjTSqd3UsiqoxCUTLjLCQ8TWLac1B1N76O
fh4kJtcA9uXUhJQuoC/P9xUXwJlqFZo1XfV8VLECS99JknelTrERj7KXdr/U527skRV3emkRvRFX
NfZzblI3oW3rHiflRVRQbiRiHlNPFy/2k6JxxsK3dqiio2nZyYfhjrkgk/audUaEKija9ZhneSqr
goTHtyMMEJhYgSOGt/TXhwA7D2uUHi7W/CxOeNqqHBSYxZsrloUb3+5VoTGZLOeSOWTlRIz3q2RR
qmlhaejkeLFQAhprfTLSmTUrg2udyMQ+IU5PttAcKtCCapKM/KvJJdelh3RUuQpkzaHo8SOoORnV
gn9wtTjw6eLv40udjXQ2Btr6v4kD48iOF55RbQ6JodBaLbLZbf1aCKjimY74fLiYkXWM3PmHGmJp
HOSAGFB+RSnH7poY6+j2mXYmznEVUyag+bhe0T0l8Ns0Lesun+mucd/a4Q0XOPnOKUqU65Uzm9He
USV/6JRssBOVFVwncBBCIFNGVtSlcEaDWMIaj7ZEfb2WC91/fBAHncgfyTCfct6vmlPivzpNRTJ1
qXP+SSxuIcgb1cgVHs1fe55wfH3TomuACSH/qy0efp0oByuqtd+b+RYVp1cToLXacOqunjVoR75H
V8tRMilMNid2VPYN4V5V0nEPyDtxzMHqmxqZfmmILLs/t7UdcPcd4JyAXlel6i+XglMfLc7AX/ej
xGs4H0pzFhoJHI+a1yV5JV+YCPr96X/Y2xhHtm0MmiTrnwo+BGBFXUNKCLGRxgnwXDJj5hMQza1G
rdQBsN/4Bg/yB+D4l5Z6zMhgQEudE5fgISgAnVnAXCOZwW3zJnHXC3lLUuTikpozY5USIwujkDTX
VZS1JKyUYjeaBaYZO07qmnxStL+Wegv/ZirzMpwXu6Sz/ooqNQeB4rrbGE2bzxJNcrObTROjxMZI
dbGf+EjcpFRFazxMYRzRCKDkP2KDuhQqGhqUlAjb/iEDHVHpj2ARccbcV5wVo5TXPkKzDVEK/Vsx
qCmfql2Z274oX8W2rkArzMVcdz2aP1W4ky8gPYILRZp9dY+w3cAjrRiYi2H+eqbIOKXvpi2QQRve
2lR5Jont1Ga+NjzfzYT09P6WOB0Gsh7DqYfHYcJd/uni3EUSNUEnZZVrhIE885zyqhO2pdRZmw5w
YMW/Wiap59wiYNPA4Duylg8qAHz9v10lUEhOCdiuQZg/XTI5FLhs5iBI7oLBiF/TJD9o9JKlUeEw
3mqMAo8Z9HhxEk5lxa8IRYQQyj/TIOVXmCY/l2z1Q0T/Zd80SJKehWCJa9QIwR2anjrXiOx/k1IK
yG6odR4OTn3zmZm5b0rumD0HZJ49PS0uFnkynKOQpoCDHdm6NFbQBO2iz5ZlFyrTudJGYlwcok9f
HJyE8YI6ZDrGpwNAYjB4e01Ve0Xtm4j0df0oIv7IRZe0GnCah5lPSfHFCsF7y8/6JHtVJKQCArAV
sb1LRfYalFWdMl8TArgCG8DtfAerWpDsaJUaaz4dbYXhhxgilmOPlR2RNK+gkjgX3yB6YrmaPMKG
Ahhg5OY2vKbknTxwp1vHVGNvv3GUhwqObW7VCaqI7+DGh3dFPTA+c6rZe0r2UaSMjRHnXQbgGjQp
Lozq4NtMoormVAcm/Be9iJ/NiZBvqo0YogJApeXMsX3/KMBZhGpj7I65nDi/fV7PTwaxtlxqIb1z
HZFb+WlRM4CO3Z95b7qVIXzLsVJmUYTjGqm+VGi/Nmp2hjKr4ICMb9E/zb+U2K1lTT7JRZaAmuep
tzxGzM/Iwp9yL6by79J4awS+FfzdyjGb9xCLHUKuOE0eJi++0AS74eoE436VFyfsqyh5TNmDC9L3
H+beRSKmtJy1ONiwYl/6jaStoNgEHa7S19CEeOw6wVliMzgXcdzzf2TaLhw55o6RLQcmmhuoaOaf
Eu4a098N4kkTl84Np7/b8rGZjsjmW9TaLZTisvHDHut35IPJcvfWyDjb3abBrnlbce4UrEk/4Zq8
Qf9/MJ57br9932JBrZYzVWp3L1TbA1mKqlLvrcEUhbU2Nrpm7bwV+LAeuYOFLPTyJ1Pm93WdYhfm
Sg9Y+jFoWtj7vZibt2wEIAwd9hJFAKVOJDPYyK8ygRCaYhk6ba4mOqQGFyBUQddU/pUKA8Xfr5Me
rTNPqrgA1EdaqGFQN6tuRxP/ig28PapljtLW+nS77yXsLfpdOXR9c6f97HwRKT+lDoikSP6RKdqJ
pFkIcf2WePFMIxs8kTD9dQB9Dmc4t/rI4IXjqts/4ZJlu5eZdZXofhje+slNzL5rBt4gbgiRuvTJ
2rcLGOAUgTTpZJbinegcvxDD91ZBZVCjgeu1LNJ8ulA1CltT7qgasdT+AxkwsVL3RLCZnNPTfzsw
nyJwLWJP5tPCDTmYrx9qloUxEpYyS6vVIbenGqTWcrjRas8DWzYSuC05NTDrC6qQhddx6tucRbVM
1KhV7N7ObowcxxJdM0wPRxXTzYUCC8zq5m8OnGqH7D1Os3B1f00jw48ylz/NUTDP/WQjYuw1NDzB
yNFYDgHxPZeAtJISH/CeAuOGJL5Z3CDxNAbSb2LoztGTaRG3hL83CKeqo7R8lUBQkbXXmZp+1NOv
kbCrm2erN1cbvre72bihEnzWRhutueUI1hbo1oOTT6WFTcm9TbnptfSt7PLPljCJ++UrVIcJt8Yh
2jGCBQeqmFJGTghCNAVm9f50AiYRY1JsO4EZ+zQsbBFE5HzoIXGnuys8Ee8+Ad8Ok8HqRzswI0+W
6UvNTXYWs+2e8MrGW+ITuoPjxOlMtimGMk3J9vitNsDxHG73vuTeiXojgvivemVC4T99h5qeaZOe
1px3JM0SAAREYf+IHNVFR2nUADLx7MWiEkLLmxyd27IfagPMfZe66WJCOPG7TeuRNTJxtGQ8zHvb
j/DoQMJ1yVYdKHeITmoYUmFJeMH0YwdASlHvyTO1/uFmoPG1hNRdfNHJCc3hWhBce8GmcEz386Uf
NCC8u/4QoC5a1MIdg2DZIVciD0wTk4zTDazRi2ra/QdbTR1fOd0gBlABAkLrSlT4gFnUc9BOv2eo
yK/y7CX5Hht2TrIo0mrjUQG/1T4MHOn0iDceN6yYQGI7ZjaWFrWV7BxeC22Z0U9FBzQOVO6WXmdj
PSy3pQIjw+PCJsnb2cd8/mdY03h0i3JK/wQ2O+y/hF/mfUwOt/viP70lnZL+ehoC3irvk7y8Z2AZ
GFCeeuvEdKkbV4CtVl+3DHxGEPv8qS6mP/1XR4pVqPosaB1rsCpNyOnxzHwkncncI8cqDX+3FT+c
Kh78frZCG8zr/KBEKcbsvl2EKzsTJa5F2JzZYDdu8Ml+KmayUqdCfXDD5Nrh57GPwdXo1nFGmRVZ
M6g0mcUSYCw0ZQrxVqbHLQWDscwxtCv7A10wqJxCjiF6PVOl280IMXy40qoSr36onnvM5yzgEFOC
QStUwOXrv8wv1YoqENHEkwLrMESEFgfXEyA3MCZSuP0QoCMwhRzadcab8MOk1OEfZ8rOqb79ErzG
4z4gVCICwOTRP2C/YOiu4CiG6YPAIyH0Lbv7UBAmP+j6XEtYM3fbDE+sg2SDkkhldh1oxL5h+p8y
MZiEmCBzAYdy4VzDx7aGUDnrjPusrkfZxFuno5C18tzKKOr3GAVhJbNqmDe8hdQoK7/n/8BRwFXA
AduDRcV8ydhmcpoGgiyrkXcNibMLXBUss4KMpJmz4n2RAw7DfrnoBqdQgHmQJeFx70shSJP5E48e
PMNb2GNcUieR/xBFEMi3CnLqdmmEJnWJkeS/l6yQzGKl6tZRX4lP912ecnKiM94c9JV8Fm8YkB4S
DZiWqhLf8iEFkPFJQ2CpaGxZxIYWvxqLiPF+2DoR7+2D/Zh6GdJnmeq3bcJpcQP2u70L0b2afhuV
ckvLxRoo6Tu1ZE/9WdvT4GJRlRHdRCR0UNxvQ+P5Q8XC42/6M1RA2Q98eInuKNJknzw5xLu20wOO
EtBvtuIHz90h5XHbJ6JgVoz25HGykLB36T5y3AV/jETNZQ8CR4xw4QNuViTUUyhpjzPEKRWCx6jO
t4WlkFJGPuxsLl/iO6fgZg+N9t/v6eGM5JBV0j88WWG/PlJJdfyCo/qHbcX4+MOM8F51HgWbPnOW
4DbGYrvDphA4Y7wwalHT1yLWJPnN2t0Qgcc/bCMnwU3d3/9U3SCkBhzPxDifTl1TD5KbZFZ+2KZb
InGnkKEfF/rsWv9ZiR668muZtS/zWlfSefk6l2AJFM1N7HmnuFfVC7t+cpHosOgrK3bf1E1BR+3h
zi4pMOfeXzlrNnH3aaU33v1vdaGQxQGp2GsENYUZu0yPWeVOyhxd3SU+V2YGOWpBNDDjJcOh3dIQ
voAITqp0V8OSCS90SQZ2KBBFXfR0Ub5siNr2mYc3ZG54iUE5JbP220g6cNO3anzVRh32exexxZ3e
zUs4slvu6eroAFy/T40QvMm1h5piS7GOL40rnlPCfMWQf2VP5s3gxd+y4rWr4+Yr4cM+gTT07OsH
8FgVktEFGKtRR8wKN7+fViAYI0VsRP/W5yaUqCdB5nb48hKrBEtxz+KDX66qp1t2y/bDKMNQ/87F
+hMRbMtgNePb1QMgBhDGoZyufZ3wpNFPqOEmHI9pV6kcq7tdguyOTkjVtuelAg4gBYOqLxBpCAAt
j8CuylkAlMiNOtD8y9JWNP69BqzvUIpyQJ36kY7t+hI/AVBoHzwspG9VidMjRo2Qj+qzSBDdMYHC
KnV1O9BhAfJJgKPO4R/n71ttBEamcwu2Ti5Kws+Nyr3UN2sWl08kGoyJJ7P4KN9BvUHuFPzYp42M
sTaHVN794RH1LaqR1DBb458lIiDTRBDwlelkAHXI/oDpxV1FC24+tQpVGZkk9Jt3fff/U2iqVORz
3KITNBvTl+GE0oKs6MEOLTTvUZSQqSGduApVDW3Z9WNTmesCaKgCTiSSzVdXHJ5uw1nJbUoEZndZ
n1RndD0aBvMN/Nfr2tk08c8vrDR8ZFvNZzWQqn2RBBsR2iwlV1XAzbBtX/DHPzWaQC42wHj9ifOh
5d3oavNv62FuDH7Lj+ttPgln1+8pUXfa3OPMzoBTpi9UMd1zMo8qTTchfR4/xt0Inb27+AeaUM6O
98hkKaQIHgfGtWQBgKs+91BvnnnQKkKTP6iWCAfmeYJa82Sd4gZsgaXhUbJ7P5gOx5MfL9C7mS2v
6l7vqeFdvfw+KM9eXzikepXIkCZ5Hdfp657MWiIqeUYbNOWfFtlwpGVUksN9DqyuE1GtSIrYfn5E
RxNt6OykaV+XYR2kj49iDD/3hqvWbz3SREPFwOdXFim4vVf8cq4ug81taSHxuRxYum+Pv9s/2XBz
O38+R9T31GSg6s2sOVhivFV1VSI77cZ2EQUNQ1lC7Dh0sgpj0W0xeFIgWhhOEmvGFGVw1FI1KLhX
dAUrajFtAIBjYKa7OzSp6PFKJ9TfANmEMr84UbYtQFO3FY/GQi+kWRa7KsSY8CrCPzDBGqi1RiL1
9m0WZrXygRsApNGLT2uIQVCQj3O29az9WAXaZ/vpuTNc03T12RXcszebfEFi2Z80IFHTmbObWA7Z
OvwuvSySAPnmvuUlgVttcb1UM7uPEeTKC/9XxqaNOo3bHKUBH/ww4D2PXb5pgSm6hDZKac34TJSI
UAtGgRKFnOdYfUdA5TzqWAE9VrBLwqM0zT+23QFmaS7jyfac1h2eiVH1h3S1xhi3eu/T6KLGzpcu
3xNbZeHcWqy5nfpbeMJzczLFaL0rvN/tzw2s/bvPw46htJcQMM1VhffFYaVw2WZNkqUDpc6a5GoX
44meaeRXvrXfCQ9aGtVz/64z1h876ZGP9KcrwWg95Pf/OkizCnaVt2hMd2kemB3tb4KleM32FHQz
4t2Ys5u1QybIfiW3qGl4d1wLyae7iKT+MunBcuKuW/ojlLCLc1y4WBqRxnK1xHHarjamCdKg9g8F
bHsC/5YrceGTfv2e4kQvTe2WYLyqg7F7m6/Ny7OJ2WIAK+TmwQMzKT0MOFNQZZR3gHn+u1K/ABdJ
aSLbEXWvfdeVen4/jrpRlce2kD8/FolswTRFo0YIlTVR/KRIsfQg6JNsPXg6wfRdtT4j80Noc5Fv
gq/Qiopv/nS/PCbP1zR+3NHITK1BaEMWUAV8XCG96wfb10T0N9R4HSUzvmzP9i1XxJwkr2XY1VT+
ycAzj5wOSTYAiH0Fzzrfp6QBmFObBI8vZ+sWaE9koczvCmPDEX1h96F58J17Xj6wuWW6BdIViy/x
gRIpE0O1SnGYlg0GQe5NW8bZlPzjXRuStZAfnPj6WkA+Q/VRPh717T+BOKtyDcsLgwIew19UHJx+
881QVDNuszVrFXSgfvCJkKjzlf88LPgPT9H1XUDWRSvITAbwQMcshkkN3uKSTr8UTi/sxNU7QN71
dfqu9/QEhhhluGLq40UGTSsFCpdLakr40pVQqTkPXVUZ6rBOQsjbsPxOmk2a73FyTWfPbVAtC4Pm
fZJN4Cz6OfmaPPFvlOM0H5b3vmZOpA/2YqYDzTy5oJgMGtcg9XjOxTBa++tE4oL4r+aAn5ixWDLT
4f8yRgLbSSxfojg61jq0i1EvOOXyZxd3Dh6EH4/rZTZzpVRJ4Z80bpnmEF/mWE9s8AVvJ5HO3TXY
nBOiqxJQNkzjd/uP/ofyyXQzJ7dXk06hkarVFTQ+Jv6Qdb1Fm9hfM+Y9jqdTh2PESZKLWWKHHDZ+
uCUhBAEhfZlCGJGI/3tH9GWUi5la+fyImRBsYfhdFW/1RAXT7T757MGSHMaoe5m9uxmBBJdIt5Lz
NyrN/TDng/TXcmeS37uB9bLrPkMn4twaObmdt9gdrvGptMyTt2y2NjGvqUiRG+DAQC+RpnV/NrUt
fdptGjLhyzLQO2A9+aJ9inVLFrat1blp5TIxFqVp71LwJC6BkcwJziVHJAWQSm6ddD+51+7U3Ocx
ODHoqc622C+dWmmIiZhUmv8XHCyN+0LffbM5fSffFieYO3X9L5Cq5PSfBGfXRhkCwKx6Po3fOTXp
Mg9gXLxMREEoe6uOQeA9pzdfUU3LIiqfGpeFvu6TMmKODjqscGkIwAXnQBZDrrKP1Uan0FrU1fAp
GLCuWbz2wo9dyi7vDDu2vpoY8nBcAmIsQnMPdgSEuKXMflfoKSgy7SdssWSK6pH+RSjkI4QkBcyC
rSTkVyAwBiChzEK8hCvXPgbBFjDlxKzh2vyg32NvHoPFQN1sJ4cS4BHhUijS5Qqvmxv4r1JVu9YO
Jr92Rc+JtorSpnqw7PtkyeIhobBDe6abGUU+yl5GgAAFColJa6SIhXpZ0WOHUQJSFYxXd0UfSrLZ
+UoNfr1yOSfsJxDHMYtm89UZ6vW8nVmGDBKh2PTbhOzC/h0Zviv9tqWw7qm5W5+075bi/S/ypch1
I+OwLZRwFEb7YqE0p1eD8vlwaPDoA1KIfzYsuljR8rpS14mczzAsjkHarznw/Rx9ALWoJ4i7GOAT
zYYUdd07P9SCiwk+E+DweuTjNTTW5CNkGOMH6o2jofFJbcMN2pUKChSdC/wvpNw9ZEZFFgU+J+ZW
y9uJJS3zvJFvrfVCnNvmZRez17YPrfYI9gdSy92JguzNuh6EAwmqaDeBkOZvemLgw/XGd+PfyNQj
7Wd1EURriyzozbbsMqkEW1OQSLAu8wQHgXNF2SFwgTZ+J5lqAo9fb+Y9gcvH7+FgolwYIAeJ4p9r
E/yKA4r/NMnWDWiOsWa8IaNyHqLJMfOJF/DSKvgkQYNxmwSGttABeEpsjnbIkyx1m8Fesk3zyNVX
TvqD9ULV90Upxps/ZT5fRRTOoQfKyPLtQbWr3f7DlXFGN0ZTu7zvLkUD1ld0gAhE64mK0kifIM01
2eulpQNoIQE2V1XAuKfJANM3A2J9vXoGmEcUsvqPHraGLmA8g3H7zxr041uieiww0FydrA5n1C0s
ac1rPy/tmnjdyMIW+Rb6pec4KgVuqd8kSeoQEHouP2kTQW8zJ+GbVVwcXTbs4zlASXBjonz+D6Yr
zy40hqks+iz1mPgdVWBNRRE/U8M+uxKbdDnI4xkHyVJCpdqrfEQIiunz0J+yS0Oipj88J8bb1hjL
UXrrGAT2JhDytvBeIS6I+fYF059J63GTqx7kEJnpS+GjByhW8VoAN+J02WBN8NOzdl2GHsCkqL1z
EKjD5yyqfHBqeh8t5CLtdR0cDShSt7WJziZ7yaKMWUsEPGOAuD5a/wxJoSKk8jhl6cEuCSLbn+kj
6eR18NTRl2JFAq/ODyXunGoskhggCsWqFOz5Mg0m7hmtrfu4uRbBta1B31n2vykK4ZC24h2RPgn6
XNxCXlG0sOBe1xUTC2RRw+PzRo3sbezPoIykyv8et2B7Cn1y9tqHP4PPXDkCVRBorhjp9KlAmopa
zHrGr2RikLdEHEyeE80nw07W9BYs1T4BV4l81bgzl7i0L0btnSY+dhaPAfkSgHyHqW4WVyj9g8Fv
hn42ZAau3RFGT/BBK7Vg7Q0xbeR4Z/RBye8ljQ+luTwxqJRCLIMRbM2tW3uzf0vCyn2gnwwJuBrn
zTVtlyMcK7XL51D+RwkDmKdfQYOTozlpUeCtUEVGvr4ElTDJf1lsXkSTKXEhLRuo4M7hvQBEd8op
TiHfO5GPv3Tsm8A0jm81zYy+kLJbzfZKwSXpzDm4buCT4VYwMsiMIreU4SpVyt69wSCj9Tf0bSgo
em7T1SrHqHTQnIR4m7ioPterSKZMxLeSdeBNcCZ+R7X0LIpwSMm5HVw4bwI42hKt1rxWfPJCHwl4
jff/T4rc/5qSE39tPY3ytlg1lOc4e4OXR/Er27gI5whI/JllFCf3iLWABsh7Ufyc/WAh1TIxBc4E
sW72Bo6IFWsjwOvSq6i1rDdNeDBvyZJdK1uG6W3lN6Na7wEL8LtRpG2hfJPhhfxnFraRbxU53eb7
Ar9OWbDh/bWqP0u41xV5y0PkaWOe7hkVIUosT9pRAExUDLDK/QF0a5Aa3RWd+2MV7N9H9bL5DSXE
ojXO7fJwxElLUkt3EYE/oEG4qYno0wczPZri1PaCnuFt/9nAo0PqxpR1dhas7ORzO/Bd4Fxjw+1l
lKNNinuh/CWKVyUB3qCi6X38LOmi40I3JLK2Ax/lMjZxLcQ1s0845AHmEPQKl7flL8XJa091V+X3
lsD/iHs//UB258SESIqTqeDtVgLnUPG1Gxrz8jWAYtnOizsa5Ygp472UuKbAiRsBWet0dI/yrDe+
HsHHrvkpqd2pnBIPBnyyLZ5HdwUSUHkvd1ED6S3OILMy0vPpSlHn+HxhfgZrvSf5PLuOlnnokoWE
OAjisdtqISJLZZ7mM8cyKjp0k+r2lqvn902q3A03luZJ4TI0ctpgHF/cnz07lyvE4anjacOpQlZF
U6luyvlYd+Rr1yhHLnLXvPnAt1hej10rRfUBAzAWEwAe4u/qHZM5mVapxWoXtRd/QmS+Gt1CiL50
TN9FhBtyiSpCz5oeaP/bckerWOzQxK6/3njZdFQa6PrlbkxaOvPu5J2AvM75KFBZXYsYy8dAvnUh
cu/mabUrstQooM7WYmWIaypy8L3ucWTEYGM7ogfjd2tJEPOlVabu0q0egPnz9NKxF4X+5ZMeBYkb
+YbcdQqTDkGf0rzC6twiWzNDLoDsh3eGG7+TFWW/HNIRJNK+oCE2SoJNo7Y/37+na5yjnc/HeWVk
/apSOoxDlTRXYxdtiaWGliqm/+Hr7C+KQqAPFlvlonMFwHWBM2uHRKSlBSQbBVipBmwTsDCjwmvZ
5EE2vQdamL7eJFIUxO1aEqpzq6WM103ouneb2aFQWRVF2IwcU17ZJm2uma/5HA1sUz7sXORoUenX
lJORWIaBDMq3moPD0GpN6sjaswYPEnEB9cUqvOfOyb5Dkwt/myDzs9kJhGFtAAw43jCEW1MzqWDO
Za1FW+y5hNczS+sk1LATRafHJ3HyfmCq+MNHdoc+OkhL8FFn6RdCZlIZ/f05oSvgFFJ0nF0j3avY
Nxn46A0sM9Tbrd4sr3Ajynl43eUjSN2DahMzPE5ktE993FlSsJMCClM+JXv8O8pc7oT2GfgoUmQI
MeFjmTPKLn6mn2WTHc3wcm8UmbwffdD1/yGAadKeM2DzdtWumZkom9VkuO5RwD3dhutQf8lIuWsb
cRMXZ8S0eVagRNHaEH/rYuRhBCLytnDcYe7fnKnh/oDwKbptc3pOwEbL0JJ2lYKqbFQcD0+Y/mEi
yxmswOkle+4+qxHvx1b6FclIafy/nqEXR88RJZFCmXDqvqDYA8cbrH5+3P9LSvW9YeZZJyIy5MRo
1W90dJ7Xu/VTOOlhhlDtiy6vpPequuQDFkrWbPF0ipcvRrmog532oCcsWd7UBjrwlv6MYDZZAJ6j
+gCuzDt62Q6VBO0Nmvti5HNgeCYCM02q0dRMCP5Xlzna9ZzUyE97xckACd254W7TD7X7eOjTtl2w
sY7GQ+EFomBu+zCYtfYBHfF+MxZTlytuM46ZtmL8R2c9C8XsTj6UW9O6ylSuzKrLWbaexqW7wJK7
xS3gFgQPLapqcxvYxziL9KzloaWpPCcuC3Tv8TYurafKfphJYpR/UyqFQzAM8YwgvVF9S/yPhcB1
bb318eM2mJ1zX1V+pilLrTpIdNNjdAB+BVUxBifTyYp5lir6PLjnjnP7kFgVAtj3U5lDbsEO0K8c
0FWzBW8QZmRypcRP+V4PV3oCkRlElrI6BAfsSZTarrIOjgbmEjMAwAoCR/MxL2NJVnIgOKbAwCBL
c3bgP3X7b2jTKrMygTXGYv8ehDQgjYzu+scpYefhn42/1/7vtisbawtEOjJbPYg6efAf+u6BiRJs
Ohv3awQ8YRCQJ6QvVU5llZNgNlKqYeKcrVlD2gYuBH8vWmby4vPNaglvrS6TleWHHTrULMyTks6e
1iNxMmbNHdhdqBea9Ecor/nJSDijw00Y7Q0BL3f86b2cJDeU5AuWzA90ZGufpT5EQ0qhp1jKuPju
4eGlvipKpG8ZzgXXWTDklt8kxt45BA4j2putVw7fVMQ8F/Ys2V30x8Sew6s/pKAsj0W93rOSGLU5
yg5Kze19A59znRcEM6EmyLV+Gbrm0YeiBUJc+I0zdxfjzX91S2FuhCq1x/sy4l123Z9PQfYuGABc
Bqsa4ZMo/BamWLMxrHOQruzWztPlvX69lxH9vQQEhqgHIbRsllygIXi9qiUbZWhRibhK9Rck7/f2
AWNQ4gTq/BcA5vGpy4uhf2Pu4lUSCyEDtwFY2eyG+n9XPWinp50fmAhjkHdvfxAIO0ANVOHXECro
VfeKCzjw0lZfXvtpsAqwqlAPEi4V1hFjLJYQnvvQnu73S7yzJsenAx8Pt+ZjuV5/BPo3nDkNNmPc
T0++b+ieYlw1b5BW26rNxeh5M0n9zjrzUUMRQVNE406sGZphPcBoWEZOgkKzTNY7rONu0aSyEkO/
1v2Gwz3ciIOBaJsvnrtl1A2HfJ2A7b4bhiXAfFZAcejpZjGCOIRpHG/UyRxaCzLiksUdmhIXqKHJ
stcL+7CuO9Aax0AbhtJXSPz5fHbRBVSVZQHVxvdm6W/xrF9JpKUMqzKcJnht2nprus65t2I9GCeO
AUebfC4YCCCeVFPSTXW4fkmxL+R+BrBts9KeYm9hvR1D9lebxpcvrVIHetj0qOpTJaiHFOnAeouB
TTsYtLjvn4NxUHGaH+DtfBDBpA+czCgEnpgDICHFhJuYhhLkwNLaMau8jzN4HRrK91ictAS+bJcq
uVTQGC8jyoWvReczRLSCAvRj/7iXpygHroyXMlQH5Bx61uDfdl8wC8RZhj1t8l9H55AQkYFnC5uc
wfik0Ac27SFHnS5iwintRzR/faZNRJAVLGOdI0gLqk566OSbHhA3NKAQz/gVX+Nk2Xfc1GwynuoK
y5UjLEr1Q7UFv4KEwnMIzAWahTZEhUfcoOQ5/xDoYuBfKrhv9phdfqEwhPX3sZw7A5TyCqHfhgBG
WROm62xtO5zs71ncQAQhYN2aFU3Rtvxe3J5Hlmz8Rqih5UBvlVpCl2roZlp7cn/7dsyRsEdLaUs2
1ZqSJQkTSFW9CajtYMP9k5VTgIbRwcwyY0y+N7UX5D80bJz4oqgbbZ2DkEA5W//nN/HPedBazM2z
FUFBAhmsF7SG+D73+5Q9JCstmV/DBprO4N2L3vZBRHk6xaOB/CpB97tPGwmGe061DsTofndjMfWK
1oG6H+EytN4TDmzdkLNWWy1Jf2+7q1oWfKqIdP6mdhZtq0ZfBBMvA8YbHXpgAZ4OaZV9ueKuSsKr
V31SAyXQ9YSDnUklHcGzu0U77CI5tpIa3QiXVIr+1gPkziLHhJlCRaBvVI/Wp3Btlbj84IOCREaN
+C65gs5j+iug7PQOnkpcjtH6owRF6x3d8DR8CO2ya19FtfT2EQhhP9UG2xEllSAZkyqhWWCnx/a8
obLwz/B9wC9C2usyZP0ZyIbVRaXNIxwrXWO7o4YXlI1P3yb77BScXknXE1AUXN8BBjA2mTwmhFVK
X0NaZaDexxVNYaf+oDLYJC8Tepsvz+2zEevi/FNKHwzX57Zxmk7DkNZ6HJq4dbMoqsqgMd1/PVtg
P+qb3XkTihh0VUm8/WVAH3DsDiQv8uxCabpZQ64NGoCRAE1Xqa3zMHtgRhUo9emNOTSBkrSBPyHr
jt1IUjSjo81gu+UCqG9KIjwdcBe8R8nNKSCfAm+Bak4G5LbiKSjIU7OnVuESqmBic277E/o6ixga
uTWOEa3Jr/mPNAzj5ppxMTzjr1Leoh6UbYxM2mHkmfxpNH4OlDqvAmRFiJkp0W+Y62ZdzhVvf+00
fTKAIe78zB1hsBiGLdu9iHf4fUtdz+0xcygX/SfIrfY/GEdP0ccgR2n5xkmJTQlXGCea0FaFYh4p
XX4KLcapYDHfQ6W1KjkNiukoa2lcH+gXloFsUgXweqTaEtBK7ybnjRM6Xek5PbNznwg3lTp+adij
Wb+i9jk6odHVWkCj/d8VMcFUzwh+v7nUHsTamwtGu5rxvzxhjwXegRybrhxo9j2NOkd3MDOQE92G
UuRA/MJshglq3yLGoQlMeqeWpamgkzOcE7vPl6GhfDVKyX1ToMsXOiSzoP3Qoz3SxzBOAP32Dmhy
Sdxy63nQ6F4lFvmPRH9fvuoANljVOm4+x0m5+hIBYGA6I+vBsLCMQ0A0PdPcwUxXkCAVR+c2naW0
2itmMAVHQRdX0wR9q7EIaL1q5lhovzdnrCWINDvhNWT4tFV+5GPfkvXX1jKJ3MC8H3tRED9s5QNL
OivEFIbP0i2N0eMkTpnwc7MiKWGJPtjeTV8IpbOGPksWya52m58Red1R7ll11NjpqsvRmFpenwsI
WUwiYqYj4jjIfhGSuj314EjY7uufHR94Ilpupe1F9PCFQcRdEoeFmsHCUuwX88UOU4W0kT4txkO5
1B3fd+QmFNrhnSM3hM8PU7vJ9xMGKTy9kACD56DOl5Vj0ygL7vXVPQrszJd9R2bGTtZEzsYrIfJF
/PCK5iLTKyBKwex+c3Wiq6m8K70PRPvbIJHXEhDPNomZ/80sWQmDqybVOobNCl57SNgRNAPSl6iE
iyzWPE0mxs12BzITxlFDd0dv1PkeK9yEHH4e477vOURTVny7anCnXt9cZCMqh95IfwYV/Cx/RLKd
iMEwA1pk7N+VMoJ6lr+6mnmYGSSR4f5lDR8XwM5fLJ/vbQsZNUm6ztHZSHwoOvy9xtpmcdad8xLD
H3qr/A83crVjWyoUDMzed+1Z0tyazmJKQXdSI9F3cmqk9iSQV7s09o+NClQsBrESUPY4WUE7tTLo
hEQ1oH6ApVNXSAh8dsKTr7LqolS/AUnLrigsTSbIf/cfvjc83TvAKfZNyGEyUOizSJnVvZTc1E3q
14+bPdAoM4UKe9MnuCLhKCXQ7NufTe5ezcVrqWPye9vtgpWcnBQbKw3p27Pr8O55uz5ARD/XCQVT
CKSRjc5D/PdJHyMj/jXd9Q+PV4zHoaSuMoB3YFIDCuxCZEF/Dz4w+Lrtgnua6i/G9eUoHIu6npsC
BCus3wq2EY3CkGvsAq3/RdkF9dp/aaLurPS/rIj37meh1VTMEbmFjQuihMC82L2dhDS7MEMrPtOP
bP3OQ2ovVgCYkyc2a+UtDEFs4jiVaFFbK1fp2SK2mPGE2eHowIG1hhKSskVMN5Y5HowlVA0KxG0r
4c7VF8tfFbpY8/Emf9uFpcXlq/E0oQns18jPf3ymjZgxN36XG5NempyGDZGQjoH6i/PVgquma51e
oJnnkMRh63LkjW+rro+zt4qIHeRlMsCYkQZjz/Uq67PPHw7GUKJjyAX+1OtZWNaSOUtxbxcXVxh/
EJfXBsH4KSEI0LCcKJnBf9eFPSAuE/4ALzKIWH+HoQ/Ikv0fbwozs8sB7iVIEWaBMYM0ZuE1Gd3P
1QhuLb07YBG35mqm/TObALEYlVCYDsSKBRzZH6Wb0BqmXspy4/ZIYc5K4+cRL+7pYhM5yZtHNszT
18RRl/8P5u0iITvpVEtVp0ie0hfHPFjPDIRASNPVGZKJq8KBM/burs9/OE5folW6m9FqjSSlibpz
oXLQdi8CCnVyPdUCn2MvipxuK698C7wy1QmSdGx5JQmoKe5LmnE7Ho5QE7Q1/zI+ICWYJf089+DQ
lgCyrgWXQSP5J1tRF5kWfiGX/FZu7FJiFJwZgvEKzosegcuZGOZs9mldwOSWIcax1+bpgsvoa3W+
CPCHc+EozTbaigfdboA5fb8C3GTjyEY4fzidI+Kn8blZFknTdasG66rB3T3O+Tu0pLHxKZQTGlmZ
vPg9wFhxXztH6IzdNmlrOFYQ6XmBIA5knf4AOgA/06eKaUoTkBGtm0vq8tME/qFIrylnwHe7NMHW
NOzvWnJIiO0BWCY4otEdx97gd2XMhN6vOSQixEUyp7KQmbGbooVMnCoKIZMYTUqL7jc3wJHMXnJ9
Xi/2q/7T74lGFhtGplo0D53VRXqRfgctSfBen6hmF2m6Bi5vpuqWsvFZ9cVglmXpMKZ7ECnS0U93
CSYZEpItTnkxCIrXlhcuhcd15/yR/MVrQSOn0A0T20npV317P7z3rZVRiuxdTUx0+an9pYghq15b
DFIOw/8TaWecqskYBuIU/QBPj/tXvna0UhhoZ+ulgMtBCBH8fFeo2oYrc9UQX9eQ+8NfjI5ZEjpj
rF8FzlsU1SqSD6SFfVeyirzV0c0Z8W6uIcwzNKeghrKsQywTs97/0ABHbozmXulAm7AXv1ZafxXA
RHOgJd+MsTm4JX/kSyVqqYgjde/rY0X2xjRjsBwq+plmAYOHLKyqidoT9C54Hk1HDaMUffrVQvPs
T6CKrzgNlPlN8NucuMxcvIvLdEOX0zYNA7ctKp3tB1NhdwYlhjVR3CgRJ5JdJI0InpqnBv1+7XM6
PDgRKuVNXeBLlRGKt0MKBSTcYZ3+0W/1UoX/MwYGjz0J4Bh7V5A0LJMd8sRGJ3Bth+gj4egpxW4x
dzwr+r1USsotyILBxlusTB2ZnsR5oP90gWvzEWBBm8fKmkS7Vslc3rU5SlOBXJEir/6amsbGLNEr
ob7itYnKyzVFn0ZEs+s37j/aAfbwkMMkwsMppBAMchz8ZU/UCzg2nzWw3XePqgWa9djcBObz+AXz
sc3WK3DOETmoiAHv82locWaC26mAC38IYBm8cRL8m8iZ6PNkej1Fqh6UxDzNuEJWoUxyfW9bgslF
F2z7cRXk48GfiVizsgi8NXo28uqLF3J3eVl3c/R6+1gOmoz3Gio5JsxO71nlgDJh8PbPdxuVvuDd
OUi+I66BsNOasnyII/t084+ie95ewcRmn9lUXOB3z4g8PpX4Qp3iLEnLYMyfwgHVnRYrXjMNupYe
dJYZQD8aKsl/KUFGIZb3ifiAIGgh6TZJlpp+jslEyA1VLma74toc540dy6O6qpVKqTuGwGLwRUW7
9EZd35D/y16oaHTn5Ws4ce+hWCqO3nCuIMOeh1pYNDWwBVxkBqAxId+82cWhRgccJ6fwSIcy46W9
g2NYWXj/cf0dF5mK4wl1HIzFNijYh7cySAkXbgv0UkisA+DyGW+gr4WxNL186Kqh5CIg6WQ0HEbz
6rNdGc8Dt0kFJ/bxv5xvJdSsfvJjCwJi/51BZVIrWApIIk+4ufdUtrlr1flshqp5kMVYF/hJPxXR
FTtf9Hn7hMdnxeXBEydRaXh6xSDlRKhRRUOFNnB2vaeUv9QWGgofPeGbaJZRxR/x9iElJSuL+G44
eL5uZ1XehY9OPACDHGWWX+PnMsQjLAcU22HziZbIYHKQNT7t/6ps/BGf5aOVC8BSz4qB+CTJheca
Qj4Yk3eTMIBDyfe8JZVeybZt8H2uUtFt1haV6ZZsgYVIXXM9fUKoCPRQgqPSWh9c/SnvHq05iA0c
KTO6whJtt8/lMN0Eoe3mFF8xPtc8miwcMpnIo2i8Hqj8layNhqIC8Uk2zcik4ZAvJkpLM9uOFiUI
5V7R2tGfm5ZRH0PPAG8Ip79SdNj+rpQHgh8QgzwXpmgiaz1L54TEclD2+9/f7qHiPx3x6zyevLc4
/94whJWjHsLiPehJOXSVMb1JAu5vpIgTWvw5MIVJVez65GxBOulzyKz1/kWcAP+4ggZUE7NSHBPt
fNRvBX0/IZKAv6sR3ny3c7eQYIeHI8P/zLbSjUw6TFj4/IzvwM9TcTVt19Y7X1N/xPMNeNwEqw/y
lKY12mnT4j9nNTb+n4g/0QEvLi4m8GGIGiYSAsDGh5lt2GRD0abHjaBRs90MLPjItXkMcWbDR+bG
gKDFoRRWPMCh40n9AOEavPOUERIdfZjThdAlJ3QadVUNEG+ixxND2NFMKAItAAHSzOJASgLZ67Cj
UguXW9iTEkl++25pv4jAYY12nd0rrb3glu8WzkUK0dpBk3LDM0L5nLGfitvCZAdSWnBkxaj/Gmfy
1hcPva5OyEUzjO4V4piEw4Sfd7vmrcPgx1eoMl+iKwnpfU1XEO4NExR/PtsR4lYMzW76KzsSOG2K
Gb8lGA/qQBSzdwTRmGzl5PpN9dqOcmVUGbM/6OLMCC1ow4CgDFLzIUO9tvLcl+ABu9Q4Pr5m9aTc
Ro+wCcvakN+LcfSJbp8KTpw72CGOU8ooVkIoD+AaQTxjy301yix2YiOPLAoHZ6TqMEraGOxmynjF
Mj/a+wxwnKHayiTHdknmEK3upU7YIRg2W+JuAS1mQrnoWVG4+Kal09GyTX+M9fODMKjrwL/jecV2
XtBn2PwFzMb/I8ll/p8swp12S8dy6sNBN3gwCtv+yD+ib8PsL4+QzkPI00p1ynA6qGkK2+073ZFA
wHM0s5Sjm0vavZVEccvvwCUrIwJVfPA7q7efHppD1PKKcrjzAfZX4cFHr2LOx1TMIMbka0L6F9m1
c+e+F2eaBeMRkX+Cfxm1ProolVLQ3UwzS6fSUqQsTRn0vkygwc5Gbdn+HEN9cJN+gbBGweTCF8S3
PlasdNFJYd3fbCC/j6cK8129977ELEY8+eUtf12NNdWFSW0FfcaHbcSdkmaFEQrMBEvNeZWbwLt+
islD81WQzpaJLEKCrk7IKzPMwqnt94mYmm9nH3uVcHqKuEm7Td2dr+6LyUQrCT8n9p9CNAwj+NIU
VH9OSS0utF/acKoI0soHKtOPsFYGaGPGYgWnJhYjJeM71NX/zBoApbOAh0skOI9mNOiIlhtnYuOc
AvLb/uph9hGqV0vTUyTL2V3EaMZ6KSgmPzjzoZVbf9e0FVCqeEEX51i5QbvMwmGRhWwBtcplnC+M
WWM0AfZFToTRQ2QcetvrkGoAS1qIds7fiRtfFAI0X6QI191xxVkxhU2u2utJcQi0uB2LbLw5S+Vx
GcIrSOSutUPrwxA8kXE/vL0LSjul04girhp/+FYEK/Hk0ZTzeBLoMdpmAXf2rqOns6xiwbFCq4GU
8xdWXy8h12HmnuF75GcJI3U4EtUQF2AC5OjhdyznOsdAOZ8kSjTLdZk/VQZfikuEer6i7DwZdjey
Kr/auT6slpy9Dz2rPcwI7xa5h3vtLCVipAEB4uzEJq24IEzSTXUZe0AdMZfZUyCgGQn+xgpIHLHd
8FknzSpQr9ZN373yhfD1UcZu4H98AC404U/U2ow7MU9ddsrNapGxC95BGR0yxCnbT7s5s5ldkxAB
LOcDVv5lApM8bnar/M2SQ/Lxelagf9xhOQWtKvtYIVj0jxVkRs2zZMNMIIuCwyO5QPQeNA8AWooA
plD4difao90KTegJ84QN4pniYwjqcDizYOTZ2roAYN0Su5cmcBMhpyMaAJm/KP3RE/IoI3QILNGn
9CgT2Oso/r7eLX3opI+FFxnnsIGEoG3SmSFCKaZPEyI2osS590PChp4znCBbfpKmjR54jzip9Qay
5rjq4AkDJq7uMLAfKf8BvtbVQ7T/szxLdymv/6rHbtjc7q2piK4FT327qEVqgffd7QBHncqkGkKC
Iukam196xYsKkR7psjIAV1sU3gaeZABUZkBBngyLImqRx+YLkrgQyEPEtx29p1hvy1pKJY0SI2mm
TzTfBMtCUKqhSQha9/VfJMbbA0g1d+F9sKT9pyZulgAg/5lezASTYYrRyPHS7wdEeVoLRWO6gACG
gZ2UtTou18Gr1+gpYJ6QCQi20Ys1cHeHjCQiLjFxBJpQfUj5yZO9TNBK8tD3npm/QlIH5XBtOW3c
k/jz+ztaC7MaIm5PGieuHVqPNIBDcGCuV56yG1F6tuc/h3nYUNIpdCWxTVBRnH8YLes/PqCOTnBQ
5N+u2Os9ZOMCvT0CS/elQ4R/S743AiGPMvrUw3fZ6rk03MVZ3woDI2iJXmQqKbVSpr/hJ9zm1UOs
Ef/5bpA9G2T6PY8euodRKLWhV2o1qAo0SF8XItyH+uzR+DoqFx06ESmEY5dSh59OIsk7KvPZp//j
Ig7UziXuW3jl/vKIO0jTwKW34u0wPEw/wouYeqKSvMwmApwu9ajodNudnSGYuzjaX4RqvjTPdQY4
Ubv75fCm9pkvtJ/OKVZNkmv2xkludW/2aaNIGkN2m4X9or4tjgPYSHtFryqhdik3JQaJBheMen9m
D/tc9fcb0pZKDhgGRE/LFNQ/M5sB+q8LmqwcGP8KH5vkCXKHfeJyUL2HUbJVaQR1hwZjAcpTRFws
g0nAhyly4wU9w4P4qJ/FKHqIPefNypL+ecm5QXIumkixqTVgNbBUE5By561b/QxWfZ2zi+cHxES9
GmXByIshlTXNRSi1fVzPctyM+0lMC/TpKn1ABqrkCxUo9D8fGMTEYgBI7cKRP25OCX05243P5hkS
sTNevFkstkp19pOdAfxIZ1EpYLjriTQP81d2fgVLuT6Ulk4MbNQ6rlEXcKfxvX/MbzTZT2dMl9wH
Jm07JGRJs5uo+8l4URA05jnkWYesCrNomeFIfL50kVtVPOzICOXAcmFrwpDvP1rskwK0iYChKf58
qi9nK9Al7oSHj+ksWe6PbMWkN3ra2ANCYhJh2e2jX+PJ3lKpocgoaohiNhIWWg2SK4rgOoGr5kRA
iRivSaLfwURUicOhK1Qs5XReA8Oo682r4Bxtqv3X+QzwPzxnkGuKBZbBbX339niNFXYzt/1QMhi1
2PxjZ5Q9pxAj9MVtbUWa6LewiFt8QueN5Q0ZYrtdhL8acPyRD8PHhV+Vm+9tepIu50T6fiFOoTzP
jOVE/tnth05/Nb6svbmX48LOhMdoT401ZhlHI54K0rwH80Cv148mAdKTDcox/jc2SMsM3LjiQpbF
W3vt2dZV3fhQuAjmgcgguW+Y7PmL803oYgz38MJ/oak4SUEyUYpaOkA8Y8Y9uF1/xFMIWgEkkVfx
6ny4b0K2t7A9Vlp8XQNNy10lzeGL2E2JXYKM8FFfAurw2OYebpSDyd3EefRvskcDuONI1qzsxXla
bnJ7Ha5FdjQOzBWxF21OGGOmQc/nbhLPqEUlCKZm4+G8ppr7JcRHInnu5UFKqX0uKiLvFY1jtawJ
E7fsnW/M4NBRbcDlYKDqgaj31hRcQyI/f2TspPOXwEupuxrP48N7TZD7+VkH/a0BZdxZSFwTgZS2
4RVl1156PZmgCh+0ABCZ1cGyTcDrI4fMLUrY574Q+5c2R+dgM1tLQQwtPN3VFeNmPb+eI6BVnM85
arZOqd9sFIQChUJwtxvnCLusDhQpSpAgBMtIxovmdECTXRPmm2rYMfZz1lrtH0D1gpsA9YEBXA/M
pntwNE92YitTuJyG+aomsHYPSzli4oRws8RE0AFRcrwWvHpL/Si9W93mnzdE2Lkvn+wZ95+uH7go
nogVRpQ53uLoQy9+WtNZVvRJpLgC8p57RxgXx8+e1P6ZUN9rkgdmOrhYM4rR4AxutOkoctSRL/yN
iqwa3d2GA2Se7vSUlRgYhoY3yCoCNDsNRNiKZHbzGOaZqGu2arr4S/F6qnxt85dOwHmU5GxFS0hv
+Ir25oskht3BNq1cvJRoBg6LcLardQ8zmYOm/ElCmYFo2M4iyhHkP/YlI5UWDvC6ZSXAPHlCab1i
rctD5mTdkJhluYdvIs44NXqMXbydud4Z2wjx/CXJhDu8qaSKbFrDeSn5mqTorltVS+F/w1CP6p9R
bTO+vlsnkx7yngk3BjzVLoyQ5zK7T/dL4mehIpUqk+Q7zc8SY7xKgUOX8ps6+zCyujFqP1PuTEEM
CeNM3meAaYdO2tatY8wMIWsd+/2zOyimImkUq2LaBX2EKQIsi/ZExjHPNR/aR+Ge89GyrWVPrkPe
5Ez9y5Mdhvx6ZLh/w8rFdUnVuYzzypCjGd9sS5S6ruIW0UwLw0tNZ+QjvB2XflZijzSH/WF1owMQ
X5C+sdN3JRlYMpSrIM5w3dNUz9iNOuiXc8PFegUGy/XmetmTiDTS1YC6yKHSGGdRYL1SiDBOMR2w
r8bNjUyNn8go72iPfgDql5mafSTPz0TCDXhkgSN3MTkq555krIPwm1bwlqyxb7gOkANWtPx9rRIq
alCInkUIpUIuXGBTtq3FJNPT5oNmUcqy7+ztoZxifBvp8+rJyAzDQ6oBm+Ha8LRxlHMpIE0LXnxX
RbdVKQCcim6GI6SlnlzVrOz0mjexd2zjuflJgom+q8D2aDrsUmJFuAvb8cNFgcBwlXyXJksG59Gj
aEDqA5Ky7ugbbkoriZ1VbGI0yG9FL/DpF/l6rfbcX9DZeYECnhoFBxkx6lTBj7brQy20+6PGIJjJ
/6wVOvqWFBm4DJKzB05LIczk5+kvGZYLOBGIgMTOH1RmZ46qpPiG1VUbNUAl7M3E8gSEX3eu+6/L
6XRJll23wfZKbBB2T01TYH3iRr3iC0DhAooNFLdktJH2RP9XDsPxngnBSGUgymYm/JD4zyKm2etZ
2TfGI5TBtNssRrLd5g1jwtD5otpgXgAAfN8SfJ7rsGOulDeSZT3L9pKaUVujr0HCmcOB3iQzIUnL
wfncV2u5jBX6Iq7EM62VH3i0eoPU+C11piiXNfV9dC6mUYxQ1aJkhDINBwQI3ofBK16dnKR8LGyU
v0Ow5eKx2uDnJ/VxaQ36ykU6InUWvEdUA8mvqNjd57X4WcBG4G2rmqe5wJ8OgaQ1k90aiUwvkcBM
JmTXDClVOWInFWigbD0husi7AxbyW8j1n3BAwFXNdHXISjbdHN8szX/sL3AZn6RPHbDFo+R0hE8q
2iRE4EHuHJ5Po9f0vvEg4czBSlWDTbeg33r7CLFfWC3oy+11HRL1rgkbik4kbyHdKU5qeoaLSn3u
lssBmr/knAZydhCb6LsnawRwPIWGdF5inYCXxWA2HeWQGK6rULou8Ywpts2Bko4TvYN/Kfpxgqdu
9yQJqGT36/SncJjm3rPB8u1fnTvAaPMhzF1BiR2bGjt5gFlDiFAAlg7PCumgZlKciYh+lp4Mh4p1
RIdsfHmjmb07C6ZCTyEaNHZnd85fwJ/mzxKjgqzVL7+Ti0smflVs3AdyYTRjIo0qoSpI0GBc7e8P
/lWo6aV5azq4krKPCKqhSU0vN+zL8sLJOCQ84gF8zX0CBGqW5t3JZgIm3/+kVVyYCI2fkSN/thHf
xLElQljWX3KAOzH+3lUVd+o/JFnGIzGMYoOlPQFEs9iTfVaXP47NN622QfCxHr5CsdARfjnYw8FO
w0K42GBtkk4K9DSIrcGPDHnD6BevMYG/PNVAHzaPi2qeioNzhL+HZ900TBs7D87ngMxYULVHfFxB
MkRe8xwZhNsGmF3NU83oUCDBoMZuVRfnmDZMydditB2DcwbUj/IrynmVfqmlcJ20/erAmBhR3orD
AclWb0UntDRpiOnx3U+cGCQkCFtEsLas1GLr1ZirJwNwgQ8VTRUsewoxyUL0I2VRpnCeYxagHo0H
aKq6FKDOH2jKpAlW6cXR28yieomGFLg3XeaF0j2mvhWiWUobDxJy01CcP3Pa68RYgYmVEKl0xIRy
5ahTTMeJhr7kmnmsqIq3rD/jgwtu9mcHFPr2NZFAc073qVcjXAnjbshQT/bSKnPS57XDXxdZffP4
uNLE76lTX97j/VqmFpcl3jaMJRYGmxGjIqWoKL3+ZlOzk6jKI4SU2wLAYTMKwzqW/8T27S+amk6m
nGO4ylJONAOxhDlv6Zzy7Iz5Cn02qKjzH09VVwfByBGYbIywl5ceF/qp9JQHGmIAw+wUJa4vQM5/
28QN2Mysc5TuXZhuoMuJnY8LFLSxsOLjT9S1mgBcDT4ZclJ6lfLwIw6ACgoD/kRmShuXMUpEHoib
mKbvTt2nzqd7Dua/gMHsN8Hyybg2zXFfS5X5wYAKVeKTLucRBgItzHsgF0hY2gHQ8VYtlTpOKAE9
i8pGhvtqztIL+tvNgVNOliqHx5CJVj94Ji1oJEoJ2rw74aWgUqsEVa8FxgFb7FHK+2F1w4gCE8JD
LQwuJdfTRQAIJdkwHA5aWJc05qUz0uFG2a94B2awHoXwehD221I59Pl7jvf0pLCx5qx+3rCvLUs8
DFKIycCcAFFHSznOxow077riMo2Wuox5GvQw3OqfdQW7OsQ7BJNJY/rt2r3Eu2LBR5x0wskJbscr
aLz7h6uj99/AqjVVhdnwU9V+F12z31t3aN7C0Begs7Wq+iSbSZhSxbHQ2+sdq8PQpRXwYUoDiRY7
bfrAnsyLKead2E63kH1FTYTYyXx6r8rsmwvC2ov8Q/I1EwZt+sApHgub/XiODjBjKjD+BN39j6Cc
R/GPJoFfo5U9M2I7zJzAACsShn/cQGuPMIbo5Y6wr1nY8wPBph66A9zNJBfYGQepmxDIUZ+XMJVv
mtyyPGGIRsw3V4zWkJSB6Ckd4IHiQ167IZvw5cLTVtFM4Uvx/KVmVMCBCJyUDDqy/HSRnaZy3fMH
Lr6Tuu95lCTbNv1yLnW6dwC3iu7anKw0HCadgk0Tktp+2U8VXtoRnrPPfy0AeN66yvrRpy8cCnx+
qS6WplYO6bSAZ4Wy9nUoxN02ZTSHWJ+Uuc5R76r9q7Wh3YjT9Fv+/oYnTl5X7pBjZ4wCIhj7WoOa
NMmbrBmWZFfQ7TjLV5RCyMhDV9O3UWv7w1qXXNfJrTCht2a35vDvLaBOvl3G1nq7txhOtDleE404
Tei8Tmt0Oc5DTB62DNLdWRXPbT0OUcKJ2IVoqCIFTAxv10iw5q6e7p5FRLrSwP/bdWd7UREaQ9so
Yhr7rHVZTEgKPVSFDFOblpmUypnrYnwMEFcMZrgVSYzF1kQPAjKUb9PnP6p/59fij832rwE7es/x
UbuqaFqgUj2WDeutHpSBkZk+1jvmArhTDYn3IzRccnf1k1iOKuR4BwmS8YxjZ2vfiaSHERZ1TOXY
L1dFQuRPwwHCKWgdc3WzxWysMGPMs7TooWyr50jSLLFNipKwM55B1isiKvRN4JB887SzhtzUaXf/
JvZ3DSOf4BLi5QWpDQ0Va+TnDeRxfZevHUcnQRUmHFQiENep3o3zUcMpBZiuEZJNcehYqNvO918X
n7Y4dfg5xnU4+IboSc0aGe+CvlcCbxjKxknNdUh9RjRi5u/2nzljg7eX4J9XOPUEMtOFxnDR3l3p
qR9XjFnrUa3VbxBOixQMN7nf9oItwP8HEIDYIwHzDsB/G1uvsN15BCLHZ59D5Y4R+afgjYHN6DQJ
gd9pNU8UnZjBXWiSkNZWcYP2H/ZDj/bJgjMAGEoNPtHDHkd6vIKP6dfEEGs/sA43zSsLQyuwlmj5
Yj1Zqrze8y4+M8ieF4NTPFs+ufHcfgeoVC/Jex9F4miXy8eWYLh01H1xu7ugMu1hQ4HAKS+Jjfh3
/iUJ8t+18+SSVnjpNgxl+A2grCfggyn9x/IKvXVlCfIhXSUbStMQD5iSt3yR4xuv5aiXSiYKQbBd
3c/9du9TxVprfseghDObI4NG5zOlErm0lMCQ/j4s4egusrs21TYoploNd7LhVfmwbTpIkd0nOGC8
PVbBQhDMXVj4ep2uo+uCDE6spyd/WNdRL4dGMMlnd0R2wCyQyVrovmbom6Od2W+QmHbHGCJ+YZRS
QrkvWhaXAelC+GrvGndnqPcRPQnMu3SlkHpTXe1J4rQrM5zulez2nGAv7zX26dxBVx2svzPoGXF+
Es+wT8VpWJhjjOB6GpFz2nugSd9HY5eegzO6ndR79vJ9yUc45Fco/10FMULziYkJvZLpVWOUUp6n
I+DKznKBlSdH93xQEU/HM3neHTxtYuqjA2bkOqwtef4a8Tp9/nSGZB2vSXbSz1L+vnS2ht7H0jVQ
+whNJKz4N+lpL6878qYGSwibjQagW8RZ5MP953E4mNktZcKFZX4QKY/kv1qhdDxx6ToJpWIPn8sI
S4iRvnzoacPS4Acs4kioSny9AFRmjSEamYc7l7Oaieb348hvILh0IMCbAJKE1N4MZYSEe4UTATEF
c+BQUkF/LsTm3H05zEVwAwm+cpVIQsYKwumIm0qGI+t8zHdyL/mQmspg9y6h2N2YzfikCokXFz7V
dLit/8ZoU6N6OP5Xb/VbpCGXjuHHYQ6X3PqfdCEua2TkNU6yi/MPCmu2B0Xnh7+4BbJP6Soze3aZ
xD97LFCv3q42vPe+YXg3FIStL+0Uoo0B8w8+05ICn5UnCYyQ9in8fezmtiGtxEAuuORt34yXPP/L
g8AqLl4bduFMvijaTU08c6rGz7xmmneeFuSBIaUIoXgY2npIWeoCDckEZiaXEB3bu2C+h3DJeoYE
xE3e2fI3F2JFUeWz0isWqCxnl1NoGaWh++VXqnM0rBNmQes5ufkqnhIUpNHv5nz11jJ8H1/p7Lv+
64vx27xqk/x+Bum59Gs43QNQWZZAHr0HqfNl+n1VGi2ZwfMlLge2GXQpRw/cmvLEdIfvLUp54Zo8
mpVIf/QtGvuY6dWYS1C6+JcR+iVewn1+LJC7TOmnGLmubLhZAfKLylS6f25vlC0dQBdO1m3lJz1k
GdrcwnGHH3x24SLRYT4MSc4oML6PqU8AZi0Hf8LWztbka/Az1B1N0XRuDhT3jKOwEZ08inuzyw2E
0B1/MSgZwyBCdX6fkfHIYj74BiYMBYRgMxWVa9o9Ml8hCpiGnZJCwo52SZZuZzACL4PbH82t54x6
5s8ZTCUiTKvt5VzkDUKAoyGQSzw+cqtsuH2Wgur/xmm87ph03lw3aCbR9DC996B6YL8Jns6iHUHg
9gOlUJ90cA7FXxhjOZe1SgwGcOE68komIzALsL/3E7RsXqPzdGR0hL3y5ODlzUzSUcPdXogVSu26
UdTT8MEmPCr1vKNG+RXd7v77BvL8L4eVo4bi1MocYgtnf9TeZqvta4K6Opa/m5MjLh7Ci9ysr7Es
nwX7biFN8pDJ6ZegnLXCxcd3zyCy9aTIV0fVsQ4eZCyJbB2K+Tyhdf78VXuIXi3Eh2mQSRkPu0T7
b5g8+ONR11vcjqVw9LZrN6kH8LYoysn+DVHA1/SSSdQAtNNwdiCHz9sNx/8WslW+sMyqtweV5327
jazecHliB73DcI9X1fl/wz39yVq3Te+6/dhpIdbNTMOtLjRd7tQs1tnpcWEkE30iR49iOo3TA7ua
RqgEB18AWtKTHAYIDZ648upb8b9RbvQibHoAQkauD8GSJ/gh2oaAsnCmi4C7iqQSbDgFPvsmHyBb
cSoOartBQZaRt9YLmo3KVadyvUVMkT7lmyYNCjwOIHX3bY689vYJMUl2Ql+yVtf9+cJSVYzj/Sfr
6Ky/N7RG1VeDqCl6DOj/xp3fdwVvdcwSGP6GDRBijgi1WM3d0UHXj1EE7HVjRZ+aqp4s29pmxIp4
eXCs8nNebJIOJ5eNYfVxhFBmHcG80OUSAUrVSJ8V7zIYKBeG/fgpQHmQJtsew4slmwFhPO4YokdR
MFNkxL/jPSPB13O0b8oooWASgFWO2o573XZdSnx3EScNdXXXrnSt2S1dGKB1HTTTNm3SHIG4u9Xd
6TwvpVXqTMhmEKhupj0isQEl/zd/Kk49f3Tsq7CBcvnKmOcbrr0k2ruB5iZFXLi2Kq2UBi+Tl3qo
gSIesQSWRpuUWeYw4ehThfxG6iWyjDpAyJJd7VURCCHLTGz5yDDvisKqhit4opxb+DFKU9lFBydc
6aAc6Z21qyhjyuGulnscdLaWXE6KUJW1LYV0rfqS4dwbLwPn28oqISMJjg/Mz3VS4l7ngl0PRUqw
TWi/PsGZZ2QPS4Ra33g41QC5xRylOEw60LWgBAhOYA6YbN46gHkY8TveIwoW41nepMsSZY7LmKnD
Khhw8+uJmdnrwDVPrLtujcyF1e6edKugMAVRXN9+viJduBK947bpWbjYecmKgesG6jsIj5sMbxJy
2oy9OB6h23REJAoyZ0FQ9q1m3HwfgmNCjpblhf56ZhOBaBUtYQLy2/YJ4lt7Azh1FdwEsU7qFk+M
zwhY26AqAa6G/oJXGv39DsbVH4cla6t3sDGJRSWl+pmfRjVPby0hANi9982Me4fB8b9tNDysphwO
Ui7AnL8ylHtYabhGSoLWXN+e1RMhX3ieiUM52Tc7j8wW/aCZAlMRI+yF/vac1BBEfa543AjbwdSl
zl408ATSLG5kqyNcMPyRyHQu3+009pEgjWqLQBWzIlQepXIv/47I4PpF1Y2kcwCK5SG2YbIpvOgj
TW4GIQXdG1509qWh3ObiapMf5FV1t/Jef0fqTbA1NMEr42dymGhbYhj/pLi4IsFwGBG82ntWv8/i
qDWlo5FpI6QoBkXnSfpwPb593eE11h6lPWLzO9TXZcEa+DBmWNk9OUJ9YJ/piUdERBkq8eeOx41x
v6tDfgajSvyYE7DRygDmFGKDMR89HBzKh3yHrwG7nkwjHUFlsuc970PeDGEaCyC4qwH8NkWjFrXK
YSbn2Bts+TlNx+N3lBoaoIjy5OAf73LMmG1LoDHKIMAzN/nnHpfBvi58Ksu3hGuqH2cnUkOELKx9
yiMjofHirrFzfNIwn4FBV/Vkmhg0LRfRy7zEL8zNb6resR6fq6UN0uCUdvsvlkUX9JXTo2bKXmkb
GfMmtlgONUjTu8oPmuoVSpZMJG4WPRgJR799aHi7VXQpJRqwVi6COxceezTL9Hm80APBZn3UewnE
FShozPeEOnNdGhX1bC+4qQvE4RdczgXPj3PEbh3rSEKGGlWwTDta+sUB8bvcjJZfO2ZDbZYt4dir
5BYlgyNP3Tb8wm2HNbUDcNznzEN11CHuCUgeTbTRp0nBSg7FcaceeltHmnRDKjziunJZ5DkHMY/A
8jqsvmwevp5ozGDHO0AKukoXY7TpHgo+LntfqkY44rWnhmsX5ootyq6Yu35sh7kbOwveS/jHQVv6
s1kKj3Sq9rHt7nl4cjN583LqDrW4sCitu7kmSZ+FJ23pWiquA1lT4By/MSiUFyPQLTBHa6I1VNLg
7sIhfo+5/3PRIl9EnvdDwtAWqafwtzbV3vd3S6zymKVm452QjH5UNJ2Y4akqXxdy/Ivw/B7ONVXq
MWKVb9RgUjzVgLAdxmsGYDEwsznsd9JC/8h6Pnh5+CS6HTMzdsz7PpCAP3hcZJAy9xEXtqVh5Pub
Dbbt+04HzROKAnwQbQ28ZcRWtBIdyuG95j4pwLEpWX3+dLJ3KWITWBNf4SQXeERsLt3D9hB4NqlH
c+2HS0c3qnoQuo3wh0/bfQ1umDiJ2K+Clloid7Q6yuz2SfPmqE9lYOAqrHvXZnhhdY5Fat3iWYUE
erPKR6ZCIwmuTjUNfjL5iUZnsfKYvCg6KCPWY7RzmJCx5rq/AaUtgjUdLJPVTCUmIqnliHv+tLIt
cqfekfFx3DagWdSVe/r+9x0WMaMywmuyBUVHEnNl47ZKeW38+Sep+0CB599ScCivkKxzHk9h2jHJ
pOglNhZcypTFCus5++afdrRF+yiKhYhNCqHlvlQLN2/EpbSpsSfjJ7O7GGO1qCjzbI08ysd7olmo
/lNllYbDxI8i5Y/6WMNvJ+lHpM5s82DoUXSInwIppDEEhMOm/HD+PT6YaMLsCdc4OR5Oo9Rt9a31
CSTD1r/eqsF47EUDn/IyIQY351njct1a//CQQ1rGi5iGMo5Ca1EpN1UnvJZ+VliVUA+gSnoxiFE3
DPgzU3+NF7nQIxM/WhazaiU04Ym1fnJiyHHPoomJQPnyarB4p4fBTNTTGipc5yoe6x1XQkUt9uyK
dh+J/9qoVpzaWMdCTWRLdGwVt7A8MAbDi6VQTfnLNT1VPmdILHffeCHUh7M7089LrH9DJkQXXDmv
iZHVAeYrIzdnRvE9+2/AFbK7DC1vyEHf9vHlffga5oxapfRDPJUWBGznsdo4wXuDzjMWfnBR4vXS
btzq6Yu8a0bZ0XmGFeQ/BEW66MCCpdwweSey1pYcXe9+XQCF2dx66Yni6AchQJ0M4FNQk6DiqQxQ
F96vNwaisQ5X+Q/Pt0KXpwqEDcjV6KHYqhHMCzT5gpwwKfVT//EyGlX8bNGFtI650xnbQioPVOfo
xvl4N71nmGH2JGQKpiHD4VngVBfAVJBDy65OXpnidAe3urLK2ppvKFSJ86fB3Ps8sw814RpH+30p
ujwWXrFVyAsEjanj18xB5P36GUaZ6kpM9hN2+BLqP6tUH/ZFJDfsCRnzIQW/tnmUBiwMzph/hFec
1rEyrEBOdb6m9cOyte8rNGAi4X0tctNVcnBqaLN/xWiRNFnk7NoRlaWiYYX+IZ4144vBMXCdbAq0
/kvOUCjA+cTiooYbxm7odq5tMadQNKM/QOkaJmJCovA+9rh41no6WCBgu+eT6TRQHYvjQjgEddh4
8yaGskdiWfegMG9QMcFgFJDXm5RVQEB/jZM129qQWbJNrX2981AE66twvGI4ZSg2K0hzGJJcVW0/
VOwhOWi0y5L5jitJ42wXfYZaEc6dIkZl9r0yWK/w+Wl1ImjXsf+kfykoQt5vj7VQyUm6uEGpp8v8
vwWttygmBAifCnKmEQyPPhDMfS45S6jHvXDf5OslPvUUXCt6dkRlH607ZY5HyV0wu77NFGzKMBjk
cbcXqdm1QPzsgRqJJHWnhP6IHQewl9r/dAJR1Ayo3C9yiE0DzdAMe47l7Bxx56e8Dovc36vI+hlw
xM9hXRLt+tgT3ndc8Gp4N/cLgKRxLkcrRLciIxhgG/zWK1p8dkLAV5vcWnLqxAisXMMGDiEeSSbX
CH7FcXsrEnzq8T2uLDaWQBEOXTqypMLMA+rfq7iUVxPVVoeP7Q1gIFsIm3r0IC9HSFzrKzl8/Z82
4k5VarqlB0Y7TGgGoZzGWT5+oB4N1+6LI1++Ezk72MPgz5syFUbiTJUx5Gt4E6KBt7evMOPcoIIT
ibuUCHkNySSHfjsc6aECzBazm7mpi7TzTKWaEiX7nCDGxqmnofmrtt+CQiozCW5AZS61EE4JyBAW
Xiv9WCd3buwAE1lpR/B4TcTz+dBcIlQDXCw86yFKPolh1n4Q2akA9GAVFB/xyCoFYOl5AQKpLLyG
pL1sWvpUPnMhsaAD6yLkWdPvT8LU3q7bH8Dy0leOAmLsv+2XZCfXPDWx3aWMBuwgvfMOqbDKLQw7
H1xbJG21uSigPPzYFsZW2DGWk5BXCkhD9xNDhSo/LTtPGykKaT+3Cf/BUbsw/fHP7W4FU/5leeIs
+TxxgD8iaaky/E0hkfo12EerHECg4jCKNg0z+PbTO7DQSqZWWgKFLmbdUDZOAU2fpUj6c0l7rR2+
k/HGibt+8Prd0sybwaqSYCHCM83UvFoG7q8vr5qhqLsoZaV38InS+4YFnmIHzKtOXOFwBg5WWLyW
dIWNKG61YnLJa9g3jBV2H57sv5cNxjorIOd1KRK/6rJLTXk/m92UqeXfwgXRbmfqhuTtSVXp7D3F
HD7jmBjpBEBr/0rIwjxpjbfpPl5F2R13o60lEURS7o/xNZrxSEHmgNHJ5emQbqoki+qUBso6eJpe
vFwpgFHbErfFtFoQSIG1E7UN5H5F6+zt+FV5UCnnIfrZC4liqbtsAjo0ydRyhNv5SIF4xwZ9mgEC
VLyp27r4OrkAiFHrJLYwBAg+dixD9tSpa0Tl18oP4TZ+RcOHbNTDs76gxmrpzdxGZDp+OpsA+9iy
TjBfOu1QhgGYzvLLYhRIF7wu2p+Sw/wVEeqrfzZ2kFQ/Ug0zhZk/IUsO8tCwGFKBZ+HoIQ73Yobg
lM1KZwS+ltvAfnA4eIsuv+ThDRXslzNikzBW1ImNnzzb92xe6ZJDPCgfscVy+fjbio43tJOCYvKG
i+kaVCmc3SRrviVy0qR8BF+9Fx5stdI8jRHIpPu9qIVQ1A3bInEsEomxQef1EO2v+G09Wfw7lgfG
cRkw3hWvFUnTh++cD798hwlsFsw079Ep/hFSvOucUQuM9GnKCaE/TL6bOjvKHk+tHl+n9NkQlZn0
utohmHoBC6vJr+2Bjhpc/mjBAvH3y/wcixzViMth7EWHSu2fzGQVoXdnNMoefOy2RfaK2umVKPTK
oPaVeLbdFsBX8r11mgG7S96DwPYFUT32LvSTRAPKQCUJg5LIRjlvtcYrGAi++j9agrXOi53qRSPo
nOb3kGREv1mhfRcMtttlA5Fcu2L+eVgqZBZCByYlTlIzU3e9G6MPLL9GRn+iD4EYZcBoK1L+PfuB
Nwew1It94W7MwR0O22+v5rksDmbz3S7NJszlcGIdtZ+dqhDuiehDSnrXbLZwudykI7/7EpraiXxJ
SlqYFTjETSVhQFcLv4dAXZ4Kdw84j1sgDjH/ruN9RpJAUYXp5eEzIvdH0tnqJFCEentaB5eFbvim
Bqj1wr+qXc99Gt/KZyFXqu59waVTOl9ooHQyPztdN5sQ8P986Q2bPBhUt0AuYEeDjoO4RvbcfjmZ
MvuI/JthmfmV+etYibKfiB/mcy8XOG5sgDVobq/P2haZSOM7VHfM/C5omJhG/05v2RUVwBoEkzze
Od5x3FGXT70122tR0+vTDXOB10Lbz0NS5bufDuFZjncXuEyBnpeMtJvObvsvaGMS1+1JNSRwXHLH
Mucoqk5/5E0GKOsHTsjltLxFDgtxeua4upyAg8RrF3T3dKv+PYv7tketudwsSCruAXU1AhlwKDI3
cR7wSLFXwQHIQiJseARGXZi/jr4AKt2ydcFg6QRJtFcusl5pDVp6sl4p8aL9LzimzoiBYLfNPpeA
NfDcBPYu4otWQYHhAVXEJI0SLSnEu9FPIXjQB/XnSJnH8XCI9mS0rqGtORdgUxbbI95tEdJcju11
b7gsc68+R5bzOtfpflUISGuvecLtVyqfl2Wywdt4pSz0DrWzN2DxM2X8wrZt5waTFkKCiZqTwfb+
6w2D4ruvjQIrH1r4nU+EiYBZIAcPhtW3o9NYgj9jfzkR9E7uQDTMR4UFBz1VLTsPNFCOpzHo+qiY
2GNJWbiY+ZF7d4cwKsQDDIGIKAqyD3lvfrdhHRE3uFazilwL8A+p8SE6wxZGL5B8ChgsECy4l6zP
AwDWDZJexRn7GRB3uwx14AsMgLqTKLYk8AutwrnDD15jYW091Z8gFrr/DpVSU64Fmdf2JFdREtFE
CbpyjvpCKH+FXJ2FyOAf58yJCA7vbh2Fn98scV/uHFKFb4Pj93Jp5Mv0ISDq8BTtpboqo4KPf4G9
ZbWfLeiG7vUs6q4rMGVH0om9mMvB9TP2hOTdGFdIkyFQg1RL/n1JAuw6NcVrIkIDK3zzCNZs1vcL
2H5UxkRGwmkzoUBOyZ6296dr35vMeqa1iA5XGgZL0vP5TK4lZLiDvV2I6974LeUl0LI71yBB62no
hw+n4eNs9nKhBpBz45dqOrKpy2KWpknJS77SWp08NWKzTZcOxqrnTpvi+J6gjwV6EKXrI/BJ2XtY
Qxv/BQtE3jTT9RerrjVWFnxwOV5DMi9bv7EArJweZJihi68dwRiHErjk+GxcrGU0rS6yKAkxbUEN
MWlpXq8DOvPTGfadZ73hY4b267UkB1fcxoIXJ+8C/ydwsVpwrlNsepcBzjYurJuohwWKq+49T01/
t/FKH3U+o9QtWHioN8kTn12jk7cVHcQl+dIckeCYSNqbbuMebz6iKeJacI5REouUeX7yUIFogKSa
Ym3Re4P2yPjyCzrV3G3WXnmHWpuDUaueasLd6yBzRrJ6Gtx43v0a6VZKJyEGhVG2dQ1s0BUFqw0e
YhIBcJycECwWOhpN2qT6jFS3TdCIb/sua7+gpsNgSch45Wt1cWCOuvoiD7UilQFfoMnTTpQvSbC2
TQBeZEUYgPf4B8WjwIfIbkLTxTe7BkhdGhXKoQ6FUcw5uwkBXFKNZT/ca443TvauZuNgBRX1ELab
gKDdW0LMpohAmOUH9NIgaHfztnQy9wdw3CxU1XMazuGk1qAFKVSMcfV7nBbXad1lP0k9MjDpOy0f
EJL4mF/EiiYSWvdr5Ows6jyzVYhwXwQH1IWQbEmdBl+W+rc7N3yC9LuJgbS8lBWXaaDJgPAGASm2
BplIfU2ZmkfH5EXFobo5q47skklK67ubVrIh9P0CnZCHyqV5z8Wjsu/RlhxynPtxsnCUeoBngXJ0
dPnIYsSPVFFIbyf9A43NekL0zXEoOaUq5oIJGciOI3GyuzTQM8Mxbz0tY48yVr9F5VlgKvuYxABH
DBuaqjlVFztnefkk5XBA8XD/Ae/PsZ3Exa8qpPQsBRHnkaOxdo+FxL3ZGNo1q+qHkG3tc/dC8cmt
4AWuTG/7Bq0hhRjPZIjYS45JKEaBTTOjtLVziKkla4Qf1fQa2AycEzaNTuRyQ2zvNPx/ayUXjWy3
iKaPrYqONdCbn2z/ASTsWQtizWnw3hGafC41J4rNS4Klfzy2t7zoUdmCSeSmmnqorvF+G+nlaMNf
5p2FdL/WrM5tu/uvFknoeCniv7TM+QOw4nQ0nceIcuUlWvwyEKrbfnTARLy5fqJ0pHsTTbRjVcA1
spCIeheLe1iy7iV/A2pikV8aztivhxKEM2CDPn61We4R+VeQVw+e/jGQ02vosPuRLY0jU9jjglnR
PyzaHPxH7UHervVHk9QLIZviHiY3v52R33w8Q2n4oX6pTeMDZW0Wq90dh5T3huu7HDQO9kTaR5Qo
HzLRiSykFnZ63mNzPuT1Y0I1GZ+bALApWJ2ucK6LrW3iblQh+bDdFGOrO4UgOUPwYTNqZ51GljwI
2kLlwFNARY8dcKgV2hIM8/94OcOpMmEQtrANYtmknodn0udbMaDusVsQVuJ/fnB80TaptmDZIyxy
TqAVp+qCS7X9yfO9vpu8g2VX+DeGoJGTVkpuUb0eelcmNV8deyERqGrtIlpq/ajQeMtKYez7Fjg8
ZQkUbbjVoVwq856VltiaOGlIcTUyRaWXiZlyuiFEP3LeJ8IssyjgwGMNB25NMSsSbhYctBDZnA86
FpsRX8sc6HM3STOm4ChsVrROTFJsPX0/kZwufFg3lowAzIQwPQo3HVxLCIvSlD/vK51GI2IBjtNv
CpHAGlBe+MGmozFlUEpgckrMMkQipOIt+0j7+1TooVxrQpBUVF+8oiO4mtv5BR/Dn9DjTd0i3jQv
T+QrO9LWBPRjJ8UppKv1rmGTKXEw3wx8dmAly1NVt8xYHsHa7Qq6JTwRiHrfhumUDpnTSkrJ5GMJ
v682GtHKm+igEVfXC/qjS+Ihgm40p4a8MJdawZsJK2MSg6CIbfDOpMIp4RQJuNfz5k8RDOw4q17n
czkaJKlBOHQEDWvfgt/xyfE4j+JHuKGKmAvwyqNXw79utf149R+kT1YNWJctGFU6y27GKarKgDuS
e2GvjAHDr5CQHGsXOF/JCzbvS/uyhI13FEcswCmdM417CPsvfFfop+12NGrgzDFlXFV0AiDakUUM
UccHMaCgHV/JG99y9/63YlPCeSsatd13JudkcAfciI2GXRY3sB8wYXQpY8pDjmoDixoB00AMORhj
AoCf9op3ivxCNrjuscGJSdCbIfR9I3iLPERcpgCoXvb5nn/TqmUJORd7CtPJncvkrLpHJCgdLjl+
ze6kArDJLiSpI3h07FQVAVOPrqCgRlB7mGZigMiAElxmXEvLqy/UKFJkvoBHDoxcdW/2hfUMGszw
24bQ+dfDuPrJyiPj86HKhBd2ZqcWygKfBGLoRlJjknfZKPi2axqQbjJEJDOOgOYUNbHH1FPj/7uV
wDe3+ijhwsGGotqZW0pHCfzBzMaQAoFtAHFdTZaY8YkRddBTOXurJtRDmZO9Cai4J+iQeIx1quzM
8c0tYhwujFtq2zKk8Xr7uYQgpE3hdGhgKe9eEbVTGmM2BldLFWuuhlhLQjpyNyRbE4se4kFnJvts
E8XF2HFlON7jgK/jOejUgnq/SX7t5aaucYXYOdzfH73wQZtqJHLWU8uLhUWW1nDb22c8hF3DTfLm
K7bEKtZyiZGDA+qLyb+yo2Hmc9alqzmXdRpAeW/LsQ1lq3ow9eoV/mKez0hrth3p3OZN5cYySY1I
lmHs1eNHEPANh/nViVv11aD0LDk4IHlL/iJJrmBFaEZuTrurFlea3VurJnH79XOcrStZQFgcjYYX
3H1v52jvperkD7xEwhFIvs087hKCPUh1u4VJL2TW4L+ULco2L95mDYCucM/U2nveMrlFzh2F7vOi
ZsleIpy2R37jmCGruQv5fDkiY3xibjZFq67QUQEUrTSIigqWWFNpkGj9niyrgd7B1Ji/n0ovZJuv
C7l26bxQZhRswvYgiLMCapBuopv58+kARgaXHtZRrhMWwhhOhnp50q8IQM1vF90Gz0WfHR+iPqAR
yrWSAYDy46bf4I1DN6Dfx+SLhH71m68GA3FcxhlU1EqRrvGFG//C958u6ExAC04Yi/G8bXQNDtqH
exM+GSbCQjYxKseM3iIJ99TKEtWaZS9NFTRQWcWCZJ5AZ4s9l8mvjw2MT8xXpWya12X82TJOVMrb
PEBIIqgzY1vnenzc1EfjPOQzxidTcY9xsbdrLZbROn1Mrv2f84rGmH4jrCoAxI4o2EIYGzhIEACQ
OVNCAmX4C8naXEJd4uVjrQ7OOADKIp5cg9HQubWnSc7O+DccIx5SjkUb1kPvKj+nITTgACWUoPya
PvLDadWkzlX/0U2RehK1coSHuuChXpvigmWrIk1Arqj/vcRI7nKV/UEp6CbzIPOv8gblNOL8i0bb
inSXrNiI/LWd5Up22Z3mn5uU6zrTfCz+xgTY8QKgwwoppECEF/sRC9pI5PgeuKWd50MarVPuqwDS
UXt85IrzAUSAZY+TPOcm6A+P1LzHUdIlCa96nShmjTZnKwGhgtXliS0cAhzvutrIldYIZKxXWcJm
ztyZmHqaipZH7kf5z4jFgcHY132vY8je/XD8cJ8g44e/80q2E91YeQeqpK/i7koHMSUW0Qr0+2V+
c6V7BGe2OmZL9Tr77h76MlEHy6MdzmVBqae0L5kxW5cKe3kEVNG+LGUxkpk4BP1CqBAceUCPTloE
mwUT5+d6lpiMjJGYl5/xfFKwT+tNo+ChbVP4JpGtx8f2VhaoLm0r6ldZ/DVzPdWRsi8rlBZsv1aB
O8BSmlJbL2e8D7bPFpQs02HVlq6QziDedFanyX2BDWazXrIXfI0GvAqJJ/inUQIYWUi88MUbbQ73
eTmhfRTrxRHmOn0e1NaEPoUHtcShzfkb0e63LE1cjudKNjVK2Hde0fmnge4f3T6M9RsKgqTD6JtR
W9kycGn3Gtvr0SVZj7XiabCUd2ldYcfWLCT/7TUImlsZdjfNU+K7WGYegt04/HHn/GvX41mzj2KB
XUGfeWbd/v2Ytdxko7TUf6kMwH47QfEySZur7eCgUB52P3QL+ChjdmduTam3BMPw2fAPX6/DEv4Z
Uf7e3in5Z2huYARHuTbMgEIhLeJdB+TTJ1OwulL6C+G+g94ReCd6+Xt+WJqLhamHek80FtLjs2D3
uI+E2Q/utaFe4TnbpHeptpKYNGzKkErPGQYwZ7iZid13C6JR8VFoGxnQfSH4vvPe3HJL9WpX6xtG
DbpFQC8JTS+AV7AhEWF68rYLL8O/5HgF6DOJ7ux3VbYABFYpukOSEFazliU+i43y49M5w3ElK00Z
/s/Pi2rfNL5nl247f9SJxwgGXrH8My6nvu2iAud/J5wraQsZpRTeLtub/8UE8var+nOfrLW6mEf2
Yj4FlryPMJgtOb815GnILKXrsxR86UVHxc6ixC948b+D0gIkF8gO4/g+eLHQ9DVt8Z6THtFwnAgT
Q0MITBL8S/4wB/E832WI40NqFiIrZqRvzgNivlg0ZQWLueNL7ADKTCo07H1vQ8xpCcJMsXW96we1
HbdVeGS5X85dJG4il7FanycqSrM0128YtfDpwNLDrVJtC1JgEboHdF0+FjhkFZBFlU7GEyTYXPS3
rjQHjuwznq+sNoyNqU+yaYTb9eY7GcYQ+SEURvHnnpEtVj2Ov29wU9LoLUDK0xppSmVFUnU/q6PU
N1DMoBFW358TFcwHZZBHvc5i26f6nk6eCuBDXIV1ZxXKzRfiGv/70SgJerXRMRxrFpkb6zquE9Lw
I9PK5pEtIJQlLu59UrOFYZLNAY4xePNEcXGOp0Lo7uSS7nILlGdC+jnyvt5vApIUDb5348D0TPIo
DK/OPnnPvqgdgVtviB+e57exDTQT/IGymb3E2kii5s5soX9CBWwM+EdETgZ2q8y/4+E3BKFBQ/Bz
N2Lcap7mOGvBgvS0Pp+fsPvTpP8IYxmHXhHKEk+ImNucZ8rh6vzJlvEj9NxSyyENQx4u3sv1ZAoL
pYUIprTGPfM6JvEEUQqktAJMkUYqsIwYr7IsUaNKnSvUdyWkJW6hiak8HQi2hxSR8K5PJAZTSMUB
KM5j17QMHP6Z/xj8Q3jcM9YvWCVEvl83zseaAQUbjSVVT3Gp54qXf0/ZY8Jmn0vou8ZY7+U7NIwy
BKt/eZpRktE2OFzXR0Kzu83O7ApRME2plmh2V+Z3RcLt/Tf03Su3BDPAMauL48VHKLOq7hXiaVTv
w84f9yQhfJjrF2GrgUa3GWnon2tXL0csbJPe/OL6hhXjkHHqGIMNuGPj/wkFDJ0CMXikbzo5C3We
EHko4KJ+UuYKULOBGezkYccBCYBhc37jdByf+vmGRa6fhBuIa42sWcUcNp+oaN5P0pZwTZwFDP9M
VmRzK8t6CSermihxAY5489ARlH5gykrV6RQqUgSgtIWGkqH9Fznks7ND0d7Kt8FqNCnCgaQD5WC4
pp3N8aG/WrjWd98SEON6ZatdVYtbGm0IE25h/m4rJmWYSLfP9Rfx8Em8ZM2BjmRq2/KYrmCmnLHy
RB4YgGeQx5Sp+mpWE7Bn29QI0yhay9cQeUAuf7LZzCwcb4lLJP5CUs+NtQRRD0t1EUasEsOGQT5F
RH13XqTH+ae+XM8FI6RtRwUPktEOD9+0cS+lfol2A9jTO80IUuQtsvcGUP/SVNHT/koan5E377nW
lK4+cPykt+Z7fvS42pu3IVzihpfFgXIywX5p3bD0RO1j99Q8Ke3r9zJRKYFspvyxA3Wx8Eim3lwp
mC3OURlFC2KK2RtdG7Ksgp/+gc+bNV55xVLfZEtRoHlgSPSbJ5ef5lenLq1HmKNjiZpzjgwMpH2N
mrvgbtJp9GnFSbKxl2PmHocybbQoaa+B2+Puw/7c0P/gsMKlgOnhyyhg3SRwa3plejEDuilEd1zo
HicM91q09z8qLO467fnVhpWF3oa1pe7e4DkpprQci7mihSB7cJFnPNLWTT1upCZ2KCzTuyF0fnX0
eTt3BToZPJtI3qCuMKP0Vg08pUAbCgL7FTz+CoCCJ2Gv3wHxfbmCeLY6I4TMYYiroxzGf+czDEoM
cunp2IJklQMvvvsNxWcmvn7ohtMJ1aJ2UtHvDxiAMWrgudv2cKEn3bNj4D/uhq/n3Hoam3EVFaJ9
ru6Con9rWIH5O3I80PWtV9PQB28IWU9LJ+n/W431d6C2tD2Iadg2ciEBdCRSbGMMsWD9QrJCEJTE
nOUhZSDM2oLW2uWO++QJ+RS1QTXPvTVZEPVeRLVecNQzg2DRSVLW7/VeJ0LZTFWRXmf0GT5xtfD0
dd7YS80mEg9psRlkNAjBgGZEWuaMBR5dHZPmh+htEpOrO1wuDBoe6QPV7yON9iNmHOEp3ul8zy5j
aveHX4c8TLZBLb0AptZBbchTMjdaJ6qVkv1gOuecn7oxk2EExaX2wAFmD2RNidxURZPoKGNLmwj9
3M6JILderKJrT30bL2pRt+umDYN/Vnq0oggkfnbKbbLHE37veUpT8pzNuzhUwplHrO8U5DfmUhRn
uTG7FuoVCxavpvy5vBWebauRDBAUWIkLdpHKX+yF7ppz7seA6qANajaHdK0Zql6AJRRFcQ761dtE
5ordiOPM89opE8MXmmC1oDet2t3/Sfpayph19r8C6/iImFhkhtVTaFUzyctG00kbdSRu9v+4HBE8
JjMI05KrSuKJFQ/iIMgUfFF6YvAdzBoQhg3TNO0UgbgskSWWecBIJinbvpBzILfjVwX0P8RfAhaz
gtf7sGMPnYiIPpiIWhin72ZnR50Pnfxg7lI40VTl9op/KdzVEOV6FbEetfQHKX4qq+ZRtILDs7RL
JDdR7frwxmoaSExydeU1aZ4M+ImwyUmGd9KFoQlBHlHtKbBlMW4IMv2+W2iTmDqsPnCX21uHSx9B
LJMsJG+jicTmT83LLEJFoNHot2I/qnw+CyzrbnKK+1jgxL1EXu3A06zujoUQ2mBxl3opxZiKEvXV
taOkXJWkIAZSSmcsMjraiNbZqIFY8/dTiH22GELtW+lW4BVkHaRzPibToIgs4XUQO/PLuXUxsXQA
t2oEihhqKfvFzxESpxIV2C3bYgeAwpFXYXFaKFx+8MPUqpSojPGZcl57mi7iDr5FZedGJxw4T7dB
WP0fOoc0MRsmUHJj06vMTPQlKCjCaQlJfXKhF0mvyUrtrRE161Io/y1FaoWmdjVrfhD/UChVQUNn
lbWLvgFUgK7Dt8QGZYco4VUQkqKYyR3iBEY3q52ysdsiQUZdsqiWMtJSMXc6d/4wvZeC1y9bdLIM
JMdu5dyPK1rNy6WOw9bTKZtEv/+dNFqgxntHc1Owtj8QSHQRwcGReYcqTxvuUIihtMjN9McwDn7B
6yIXJxwTUpmGzxwLoWwJFsUZNe0tvCce1QDUy4jWOLeSFyF5AodIm69r+C+h+41IioHdfzSDK3/5
jGAA8eaKDdA2K4V7zDmaZvVv7xkVCW9yV/Kvyq6EidJps+E8LpVn9gqSjYMh1iz5Vqe5zwGJwpiN
Ma2HdIuvmTKFg9s0dvd3c778Sqb6Oco8TMxv3zoOR3D5+Y7MNlQTyrum9fRb98mcowZ7+LvfJVEs
aIX93p2estzz8vsemDV4BS6Vlzw7moEZ+xPAfVQ/QZ89AC25Zsz8/ks+Emac+WENqlzl9iCnBQy5
1yi03seg171YOgPhl64Hl1bUehUfEUKqQXMUb/MhlXTUEKxQYIo5We/Lsx2dpuqznr5ccd6ojzrJ
n5qzJjLxZSM73Q52qf/A09L01gCvbpJfB6fiI+D3rMpp++/T0ntX0dZgk8nO0BXsDZ+Dc7A74fQu
jTue5od2vL6NtxnjBFbJCyOAjPxi0kIZPEhvQ8ERQVBRlYCZdI/tIahtKjyAdAv20UPpm0o440+/
+i0DAeJQMSOmdy4nUIVOkEvz4fBJ4lybsFhzNOUsYzWB7stgWjQJ3sZ3ghMaUgxuV9lJA+RTKh7J
VEsUk4gVuclwgu9KiNnI/GelBB376Lza24lHYtvlA7ZcSvCVKIOsR1Hp2SMI/xUu85gU/HZ8Sfwv
rI5CJF57cKQRtNwOXvciJIi6oSka+ccUyxLV0FZa/pc/ZgpcNmUVjTUsexkRMUJ3yi34c9iVuUgu
D+Fr3FSGhfrmxfCoZ9PjYycx8EsF9V5JLo0CVDzQ18rfsLjRSnf2MBeGAoiG4DHsxmB1kM3r29Ze
EcvrD4ZdvU/+TBdvbNtH1MEGMBsXO3oOaaPf4n47HvJVShXJd3aTfc0vY/Hx57kj1W3jRTQGC2cd
qmDHzYwgUmqrGH2pG338lw0Ozgl2uBhhecV23O8tXhsBemkvo3P8ccKVcyS4FFu+rHeTe8e658ba
ZgDuamfA1MqGhNO327sL/OVdvh4hCqViY6yHCy/qc7xORbykXWeFxIesnxTHxtjP1DUyNeYlsS0w
Wr25cyLtMzn11PsYQWFajfUhM1gYO8FDs9mTeWcjYHhFhMqZI2KbJYGjIIT50504zPqrh3nse5qa
7nEXt4F9S4ljuJsNEEFkeLhG8lmroJAo9ytKUaYrTZudm6Qcsm4j7TjMNY02b2RedJdqtfxGjbML
GdMBgvydK1SEvc/Y20kcODHJutFv7JunnhMFzQDjlIRBPrd4DlEs9gpOoD9u/RjBa/U+ONWgDh9y
fYEgYZM+ZQ0haR13/XTft6UUdsLpaU5Nt+0pPGUgVuRvZTwCM1QP5bCbBFAb8leuU2KpSXqHZ20d
XDnGHublAgjupOPrHpsvjuwYxlHaPk0oaWuB8dXGTGG/WY3jnpgITTqZ+f83TFyCjkiTw5775QoR
gW7r2XGBqQsZIt/pl9VgVvKsWvfDbHr30oaMZ7oLuygLiIGE3Aa9u4tlNYp20LBrM0Lq++zqwoHS
c/wBJd5by/jKcwH6gDT0ds2IBpeINwp6oTDIdBsQR8cibpDkipeR7vZ+kHXuNo0Fpfdo1WSfen4S
mvf26F97EWZ9QN4zc/BNRNBM6V1x5aqeNpAuYLkXjrlSJsKwF9wfNzrfRvY/jpRayzB/BMueN/eK
10i9SVyq0CIXhOTD305dCD3d8cMk7awTLQ0+Sz/lJT/zmlnPwHtoc6bn/c4m2oBahC4RwbnPieTa
itAVqToQNuITEKwz4cUBT7JLJLKVRRjxHek1yHeC8I3IjEUGP7hF0RW8VuBww/U8mYfUFW/kLc1t
CgrPZ5s7obwSRh4bXrM7sf+m1nHSIray9/+/Rqwg6NR53HLjH/tKqyPEpUx/9sz5XQzJUrCrDaVy
/ovDZJSIj/1/FmxXyrd5uIvxzOFWdBMFQsdi7LN/zlEwwNgzLd/x1GyyIahaMTU8FFl4u48TDIuq
2cu+/ZIbVhZDSD7uOcI1AfQm7riWerq6SsxGbTY6VN8nHncQGySP5mmo57Bx0DPQw7cfbvlpEw6u
9U/hFhXjVWdz88aW62VfXIozVuvLtb/hn1gyrgtfPPZCkAhELc6hnJ6L8BYMqbwCnL9sb+t1ZJ7h
4c2LHe4pXz9najr+s52w8G8LZveN14HdOG27JRyUDHj/2EmMOFAxi18OeIDlM/ub1Y/RxDkWgfu8
LSFRINypUDPjOBYipQr88YIiAQd0X04mkiSqYfrklVwHiN2TKFF7JNJKdOGT/qZz581J9K0EPJPj
TIVAGFmMoHKtyg7tld1KTw20diuhxkazSU3GlZuSVD0cxxbG/ZfxZs9yuomxUa763GabNCavdSZT
PtsprqsyXK9kBURtYjgWrJPIeLxOgBk0vrZ8FBJqK/WVVGsVqpKUaPVZNbMD35lcxt+KV3oGdV/F
oRhwyAtcsMmddWkaJbZIJasiIGqH7qMUiVvBFS0ozrk0CC0lDBEE79y6AU/fagCtx1OyCZ+zZKwx
2AfxKu4hMEYEvawVPjDdMyxK/amK7eZa5rQay8211NlhWWb16EOS7Zkj5L5BAfW9g4N/S+JqiIxJ
0yFNvJ04DEvQyIQ8aILrlhp/+Eqbf6A//dB0zDaGEymXZA0h+QZRQnD/Wp8scFn1WhZdpAFILwHl
JK2Sndd/eL9dU3mQmzQM0yeZs13seKn9NOUJvbARlkT7fG8vQb4frpHmATWp1DZIkwLZvI3W8kY5
pvhLWr/Eig42SZVoq3xSSXCwIM6i+sGmBW+/fRGXdKFzYuOPONDRiksn/tpEXSOAzySfvFl9+SJp
5WbCMhqT7LsLB0Lqqkx1JUS4nkXkzfEJ597P3RAy4NBDqF6xMsBO35cbOWM/P7RsijkMp+4PSbUK
i1+u8trvidF1xFH7u8ZYc0bu1EBTsFLey7tPwvS6HOjWWCXuox4UjL0siN/xDpr52WRsNxOTZ7Yv
/abcT7uA1FE2QjmbmBlSBExBMwWMU8jDDHYMP9K0FySOFiwDGX1Go5nOBMDBdGXBEWTEYjgtCovV
5yM3NB2IpekGzrEwVeDXMR0xwm34ujTznsyoLxBXG0ctgVPETC94S6IhMSzvKS1kRNfxk65HD6Z2
e+ujzkUqKgQfibjhYcp0XspkEWd5Oz5ZQmDd3aRhnkiKsnEpQbc2g7wAuehNqZc0V5Z6uZiuqxVa
/AeoWH12eu1V0zZX3+uRjFRNJlt42LYTVi43AVc5/fLQyS+g+WpiBL2U71x7zEsb0EBtNTAtykJB
AqgxjQzlQy5SjJjAq/Lb9OZre6sqPE1hd8wmWru+o02wAp4SO3EmtY6sxVUxtqefFcyqYgFCylyc
vA2/NWDeYrhceEgKT8Pe3yKrJO+lg8AGcA1XtgvsAy1GerKbSe70pPVzQPalGACgFZV6Oe8A47bv
HvPs/23tVUNBxNxaPWUiDv+N2EVqlolVFXJSroEEHC5GY9Zb8b2EmWdpUC+0Z417u+WITnKeIZWm
Bf80pjCINKH4K9+i5tGRK2AuK/pWZvLGMeZSUYQy5t+nbvCm90K+tac6SWmy0lotmWw3N+wFpsFs
/R8PwxHaZnp37qeeEMzAW/MiE9olwsFa8UN+Gmt2vo4/nY2RrkkwWEbGHYK8eGiN9FFvK93U5mps
sJXeJj23qsOeeq7ukiQfFpCxxmu8fTvKbsix8a38xzTDEuyjXlskeybNRFpwCTC6gvkBX3G0pg6B
wcrcYK6et5zz1VyM/pjTML4pEN/dueyhsJ/Kpk0F6U5t2NAzArqVhdW5pWNi+okGu4EumOqfsuZC
LbQ6wNUxzHk/YoSEpUU4yMFom+BFM2nix+D7I/wS747HSMmpb5Y446BWek9bPts04h6z2o2qAUnh
uj2NpO5v93iM9Co2e4ZkkDHii1bDEqS1/j54wAluLIOdfNrh26vGe7n+/1kDt+Mk1eZqAfqN285m
K666i2X0IPsCNW/DwLUd40lf5LA0ZTI1Cw8TGYX1Nf/gvS+kBBhpjnYCLYSc/DsRf5TZzHHdMs3e
vn1jUHXoxf5eD2SGIu2p67bvbdULFaQQHvvXAsGNyFm+TIqVNyWIJIIkpPUs0tTRoT7UWK41bpvW
ia1nMyexj0YygyKXk841tjQU4HDRIF9LEsC0OKSYAcY8lwsRPTNoCITpORzl/QR9piSR0DOzkmMk
QwbUUWfc5rrPjbho9zCGOlQIBhdU5whmyGnVl68AalirdcQG8h5WrKMkmgDbwbRRDfWU9f40IaBw
S4ABqPWVY3nffq4cPCyJVoVvruZRHUcCv1ekWncEV5cYkITgaXPH0ylw5OrHIhk+D9Fd23qL/bJG
eVM89U6ci/HZDGU9mtLK/+uz6LzkanDLfm+Bu2LcsMx14pQKhwly6c2D+i8+HCAfB6y+HuEgEadq
mSpQ3ijDEa82XsvXS8HvJn9ULnZBEHrABy6hAfdjP0YifR3lfG7mZ/bdVH/ThKjyzIs7BjwDNYkA
8EDURAbgkwbJlGR6VBavaJOGF3KUJVW3IyzNR8mJZw09s8zOQ3cc5/TYWNNALRSEN1eDozQK085I
GL6eEbdh8P2rm/qjWrKYwyPpXHAUF8z0w58JukeAAttiwUsBJy0KQFx9/UnzAri5+PQbEJAoVfds
Lr/i3jlQu2vZrXr/V4jl1b7lSDPKKVMxCVw2kyajAcKDJ4UPCHcbTtOXs9mJJXggI8r2Ulb4JwrJ
R860/OLD63bQIQelstIXpPxR9OAUQ6uOT+s62a0lNWYGZ9y5+g03nNiurmF/ulqMmik7LczLUg9X
h8y8dSP/buk49BFSNrn0cfnk5x4AUhbrklNXc9zRoH5HUbJpz095kiI+6/6DkGvPZPmYMsvCmbil
ppuJn5LC4lNNazaWcX3wnwezMLqj1dfSfyDszDmb14eNn4EPGGzZCxU02XyiEMOgru0wK8WaCS/F
aeb4L2q4GoT6+rPB2gdXA5Gy0BzuWHFVcz0qTPoYpKV//My+CldXOBZoNqYKE2QpY4slSsjzi/Gg
uwpwA7hZZZEKfKv2bGGKo8t6l1EuMzs/bz7hb29siijihxL50eNsTT3F7Dyq40K8ybDdKEOqtaPX
+XxfDPQb2dELYwJ5ooBM+LYRHaudmoNfr7sryXcBLgAMfZ6LQNxxldKgChdFFfqZRdluRFjUi6Ms
y+pFm33QTzakn/yX0yOnPIo2g2eIjBhtNRe3FxxqeQOnouR6HCbxTHeHtO7Gw9frfLCwZ9MD9C0E
LkK8HxmkqOcetY9bG2a4u9p9CPr/tGRKq4lz+hNXQtX6Za9hZzMfxce1vFjlOsRMve/1JGFY66Dr
GNSc+IbBBz6WwK29f2I0tr8zbLcBkumb0vo/x/0ySgCzCRVF2sCTq/5y3Wie2nDNDci6HyP7axO0
T2bKEzWUe0fyuVDfujCkMMOGBc8vZ81AJeOC0EA6bcHiQSnCx/FQ4OSNipdc+iRh/gSBIcci85kO
sdGZgCTUgLj4CPNhiS0UpWQQHHQRzO7bLbBu5ac8zxKOEGlPh1dMcNs2wtBedr6FcDnPIo7WDQsz
F97oHts8ovDsURqbU4ERBRszyX3wvdWjzvnN5/nhkFD/OzC04f0mFoVtlCQedTP6k4cXnV/xAALH
a/oXDAmL660MPsDtf+HSVIhObkLcdz30ZXzHyNUmoKNB/43IzXL95c6/Br4bdAHFgTNDgFeXC4YH
YLHCt4QfilafRW8h1WpYEGSzE5cnSalCZMqfq+pbBygNIIb3taAhTF7MrCN6XqV8vN8eeBqji8cv
AnYdLP6tyQScdv8CngLI1J16xPdc96s53AJCrRym3E1BSR7pVZvXEyeoccprdaLDx7HYzFRlc3FO
wnQkVwO4CoD+HABAGhD5YQgTV/SVpEd3KP9sIDiPmPXCW7D/JYlefKFWKDjUBe+5pTUfSaX5L+jm
XTD0E3i1p6cvJ0pjc4Ym5hBV3eoNU8O8PDGPMZggoH+1e+foyDRjc0U5u2eO5YzrAElE5zbFmWhQ
5FN4ZqmeJmV+Z10aqC1uvj4bbfTkdjo0p/AF/CSmxCSKWA1avMrN5lo5CMrOt4E1nmGQHMXOBVOw
RG50taflCHZRjAt3aSfWf6k54ukgNhpr5R6H1lj3klOQUjMUORFUF5snMcH+WEdXjcKpkpknR9Mo
VlI3WEXOZB15849wNmIkoN8YzEj6MHNkL95acbFeHQEieyd7Ct3xfZbAiDp2RHpDP3aX51E2Fpok
TvnGGk1HQAqd9hyOFqHYELZ2l74VcBQYVFlMgSvagVwvsanLucG1wAmAdq6x7SytHbhRNzrICAri
h/PRCLtkqft1FmNW8MWRvMsy2D7XR5/CFlMz4ixj62/hIngB8u63OZadD0IeWDfIOASdvEzZSPpd
QKVEsmhJ+D1lNEEyAFbkWkGtw65yfosW5i9L+rmr5ePWUa+4ayq4j/3rkRtL2jlVWNll7odueSSY
fYmFlq+dY2UMsoOmWjC3yZX8MrCAWvWkuRf7ckXCGPkkIV95n8QEjNAz/E4nl+WmjgJtkdCYxLIz
89Gy0d3ZTN48fW0CfzHdZRjTirxW7/3oD3yp60m93QNikdmKvfrfDtdYFAdo0LoCy3hyB41OlxAU
dVKsppXrivhdr/zg1U1/yZxjOxUv+kTkMhycDVL/0AX2fO/l+AU6pEw7R0ItvXeEUxQanKiyFuuP
f+PY5hIgNaLU/truX9E+y4lOFpM7tCpsDJuSMs9EdvP7a+T7/ZCtdpdZgvp084K/NDb/5FS9yC27
pb/5aFggf7ud6HAranu3Pwvh+hjoPL04fInh7yPOspE10YVTV+BoEnMIYg+R9XSSQvJBbmMbLpYu
k+FB2RtPNZETaKFh5FASeAj60xmoaEcqDRH5BN83Fr2QHlolmBSAYsT5OZjctAo/5kIFU35SKdgj
Gb0+JAII/t/RYHsD7nTASOLCRbZH49H6xXfLcdWlpq1THCVyUN9U5yVtUWhrjo52R71DVJnz1aaD
6zYGj1QWkH2O1LU1a5gDRC/xmNkkUcXmYYdC/tVuSB+vzFqeI4qKb4PDQgCJdOr+kiQjE2h9bYy8
YNTgVquJ/k7DMmnOiXwgKqsipiBenDQisB5JMb89QmhVMDraYWZmNWmvKgHz/gwgOyfJX4ouIbkM
kzfhtdM0vpuCbkYkmTfw2/yI5QZtFlVCmflFRo5Vqklh0273futilEvQTN2Kw/wSJ1xIDNnsCVh5
o2HkHNDSBFtS3ClaVkuujnq0CvsJu43c4msrAhGwsx6uGgOtlScS8+mtjVXicN9h7P6V/7wUtxxm
JFDiNwPBgGfBkchq6SzkREn0m+dDq2+DgpmlbkZyTIRy63Fe6fHuB9aM8BHtX0FrwA3gaSNtx6bi
i3C85HOZYzJ2GOBO5MChaA99JLgW8Ggh6mwxlWGc3//ozA4HNuH6AqJPuz3a0nzEHZmYfiO2VVx0
sn2mK4iTgW61siiRoRO8iIgnfvRi5Lw8vQiyDxyfsmCC//MIMZn6YBIcLVxBnVljUwDpyotBXIc5
QDtUol1atnWBi9+gfEMrk72e/MWDfNxOvTKhbeauQOsun4G2oHXFSp0TQlNc69ds+HbtLMEqdM1+
KmxZF3nwRy7n5xpEhu05CioRElA2CVg/mgdTiaXhV0QGQQ8DDrS1U2HB1+PWhcB0zGPPCxVAJxaQ
ZIXjRNOGBjomauJn6i7t80tJFa8dfPO8cB6i14A532wKroLFesUmx+gw5VV8nFoeyN6aqcwxCdSI
umVRL2yGKg193J9ajP+tzii5ywLf0sbiHRi7IE4YoUEm3iiDdpf03ElcNRSmmOWp2yObQI+1LbYM
HjanDdvQF+KWitvbVf1eA1/CNHv2xDdQ+Wpw0yaHzm3C7WryAwhRV8Jf0VNg1p+Peb8tXVofEhIb
2NsUrMjHkjPrYNn97ozD42Ozi9qyCcFFpEDlUWkPpemeEYrSYmpCVFnjEg5jcI/k+wWIefE6oIc0
mmgQoSEmA1p7DdizWn/wf96ffQo/5DdhkTHz3RChpg456PlpBRwj5vBtNc8e9QB2HBWYb114xyj2
bLex32tQ1TlMgkxjSnXHy6b+JNkGMTg+xtgBksLWfEdEEMdmxXJZTtOAv5O3jl+fmYPSd56Zg3W/
RIBcxySU2WvsPZy7Vo6ch0Qg0j+6S0GC3BGtlevHX5ZuZs/Ws03VyEjYwDPsk0U3Wz4+cOuW3fP9
BNmOpXd4NorrgNHjeeOPEJKj86ZlcbI0xu8xFLowoNAxaL9MxBTduZcdBwKCZAud9nw1pqXslz3j
R5JdWVFazbHA+xQBmmdRI3gz9CcvrIoMTBVs9pEK4omCa+6nlv+MwlzCg2lGYaqTKTgcdkQTRxl2
m0O3rW3MfT8Mg4UM9XuNc8UAemD6viQfes3oJySoiZ+FQbCaDMh07dI/tAUdd38aWYYC5SXhVX+d
9LY/Sv9bh3JLNYQiEy/IWxv8+BjlkSVhr4gUVHG2VHVEpld/W67NUbme/GvyugAqFE0WdQxvOPQY
agKfF9jcpoM3wMY/PRAuUZSgWXF+ed0qpS8OQWXCWgVvkfi2eSCwMvMPRSn0e/BymQ4ZZLFeBKQO
bHrx7Edy6nL9TC7Xpa8UDeE2PogiFR6rwHV0/o3/yBtECdlvTUSk9pmpq0aEPYY3ub+pkeFsOJg5
vHJKMk8ODKB6DjARHS5qs/gKQO/pPfMeC7AILIln4Ws82fUl56EguHOX7BmrLn9M6yU/qV11vQC6
cWVazREOV8zok4IKxEhfPaT1YN4MUIGTu6FglCJpXEpsWgBlYrbiWhrKNr0EDEj0qprmSCjg3zNx
rjrLjaD8bcM7EOe7G6lU5dixOlZyt08X2Lnhg8orw+qo+KAUaJx5qQrHaFjtjB5Q7gr6secnqa3J
1v99mWIZ8nXitS1lY9Qu1t+hqCk28dSxDxTmkVTAIAcNRmYCHdPJE8QqT301aDTmx9UK/EaJBeDV
wR+L9We4BjMLfj5mJF5hR5hx/MizCrr3EM18V9b5CYR0WpoY7rXgBA/wKIl2LAY5eO1adzCiZt0i
kk+7vaM+UhEV1ew8RlOeWxm84IWzmLJBT6YmMuPVB5UEq+0r0BrVT7Ynz7egbMoldrQwf7VSIxtO
jXZ/5GUo+oTQiWbI3Rp2Tzk5VbnLjUZ+Wov5wlcmjsyH8iNzWrovQEOeI0E/XK+9H9vfxBPI6Oko
9/fULbSaVYJvxUREOmn/oZfVN7DDJt2E9dklXe1jujVhjGZAw/nIvtmD/Agw0x7tAcEwovzeCHEM
JoHHjtuLKYv9NELk1zCUWoLECj+Gz62nwyWdAZ4VbrTldS9nQoYfMN0Z9que2RbRTuN4gniwGTzi
H5georiHDm/Cl2nYs0PecvXmFUw0oRAHVF1zcQtYiEFzni7JJLGMfRnHcHLJF9GGpVjEWn68PAf7
rM8JjK967yenT9pcogJ1t3Br9ktOGQx6w5jOs3ViZm524VdWow3o9C/TddKl1DGNC+rds7BLnj1L
/swFNoX2Uvx+gMnRtG552twkAe5jcC/e2c9fg4HmFt60QuPhkFDtBRcI57Swd2FQIG7/YnnwhZz+
vRCv4/gqkaUrVBovumfWoElckSXgBCUNeLsZg2MNw46n1+UvSuA0CRoRnsYNbZbM1J67WTcBwU47
tx5zT+oiJyhC7XKSH3lABBTR/9zDlz+98p+BCrPBLx2/ZqgIXOumPOYOPdaM41qTYZ2+r3Gi7l2Q
9cQ+8J7w0FKYCHz/4CyopJGRMPN9YAREM/6/Yz/eBUS60nGi6nqn5GfjXL0WHVjImUhALJAwB/b9
ky0DQo5PZJB2WJr1+SCyoQdxdy369HU9SswwqYWWO5eaWtH5gtJo+9/MjKt5wCJwICQaCuQYSurS
c309kf0V87IDvoWRnUSichDAYZp2erq36TcV9QfzihaPlyPyYpTAQSENv9upZwZYKUVQtj1zFdG4
6ULc21eS1VRTCJy4/hJv+g/JM5dvqdqUSy90Ws3mHN+MtrV28H+rypMJLDenN68t+v7U3Ri2op2C
srEXDcuw/78nUGlm/yCF6rzJNv+A1fGDsuRgqRssAia+a/gSyzSq7ObDgMgrpXrN797BTv6ab44a
dxBltFYtr6iJWmYmX+ud2io97SqTO7vDXqqND8uM7H4M/j1MxXicZEXrCuMBWyfVu0WwVRnVNT4l
EyzVUeGvoI4BMGg1HFSCkKL7LHUhhGiA5atbqKZ4HAcbYn8+TL5KlR9BEO4Q6odLS6LZofQAzx3Q
1vZlB+4fQc0ALstKf2o1nNZZUWhpE/6nlBhHlet2MAVSpS7gMrKEkbl2PD1e1YAfGqxs/GJgBmaZ
CuwAi16J7wZ3iMmTFlRxrduwN4nlATfRLdisXJ1fbhlOKkB3IMnIusz0ywuLuDSqRJwRxyy6gEHa
7+HKhHU2w/aLLu9R4cGuYgTk2EWc+POkr4A8oLsTtSbRbZD0rJzg00iqF/6MlrvvnodtCVLJDtVj
IPmP3N3uoqgpHO+si+2jXH5yNUokzqYDFrwVGFm7k/yPr/AkMda7OvGzcTEMwWozK9JeMYRe/RXp
ZczqrLijcKodWgFuHhv+x4ESyiUcf2D4LaRYQGanofFK5uec/5nUEy8gzLlD87MP8vfSiIr9PG8V
LcDFUpBUdbYKPU4dYhkccRBhfrLtE+algzIRiKt7EbKTHr8Yk12Q5y7huqYI3uLBzTaqzkf0AO2C
Yhvb3ofmzGF+dh29clZ99IWfcao7DsIYqECaFWV7gLoT48KNucj3IvtGyOgOBTivCid8JAWqAhrV
mHmiEdxL+s2YefBRm3eoCe831VNnAsMQ9+Z1qqQAKirLRDFFKsrhug6p/zJvAaL+e/IT59x9jX88
n3z7jth7GFaDQt2qEtJNbzqwAbVpMvNPMDT7NAGaceqgzxrJRaHDTupfEHbarffBkY9SJUEbS75I
CmFVhB0sCt5hqy7XI/mszKvv12iuYve7qYieUEiDWh5gXmcfzsJ12EZNDc6d4Yzz0bkZkUSUQ0TZ
tzFsAvHVUrTnMy+ulImCsQNnmzqPESDB8Z1F/T9tK656vSGgofFbSzclTLIVBuNgH3c7Qf6nry5+
X+qzAMryOKkZb4jU0smdO6X/QCaLbxT5qed1VHviNCVbl0bQ64OPOZ1iE0Ds7AlUrjxnOnt1DE7j
GCtaOEsbNS6J6mNHFXEsXjS8O6gp65bB2PpXz7XSoCSMsXa/jWKBIUp1yqiHQ3h6x5i7gNnuifRg
PiPLbsDohJ7rvZ0v4FUwOs0hL3SJiPxYZH3vXKekPkjPuXeGHdcfz4hrp1fUIbg47y8j64Nyy0yS
GBCLz4N/25+3xb/cVp6YbKgawHoJ9F/ICq1shHmr24rjgceCn7Vnvsn0tFuaYe2zbJmbU2/MKvwt
QIw/F9iUj3HL0URgPkrBcc3p9YzoHcsYWTbadvY8kj9lfbZmUxUpDJk4W0TfIDkh50iFJnafQoiR
/9msJUHJKOqu2xnHWHVxovsFr2viNJVFl7/lqOnSWmTnnw1bJ+IkVSIrPYzKZfyfWeJnBnaXjnnh
4gaWu5PwfSu3c7nu1DbVmiMOKC5Z5OjAHlKBc69CCO7AmixzYtllkckjXsvgl06twlmMxGHv2/Ra
ktWJvQEjhSaB8rsEMnWCrMb6jhmn2aMSPHWpdTBGgM3hXcOarTUAAe5ip2lCqjv1pz9viXMR0sBu
99rEcz5zagTagK5rlMCwsDKNIVBX33/XLQBVItnLVUnD5q9apuJeB6oDwQfqh7dgRrE1S8IOTRLQ
208q0/hg3/kUhz6QB+DNVCoJJGVPlMg2fLqcaxig2uxP+8fvIDFPglESB8IcQo2SXIOANLSL7LLm
0Erve7TYpBG0fhreYI15UYleOenyp1Pez8X2rdtNNCMydFFt6Qnbjj1Pf6y+ZEfDgUpaK8tVOQ6U
TQKS2yiSOoivKTTSLs19ZLlf5yIzFl2FZe/6a/klRm/iFj+GphRyZF2PKauzjsLwrewTnzBMMNu5
kszKzhm9YQNLnutNMsUOD9W8jhhXcOi/tmCeRFJyeXHKRC8pf4OFkVFfLUci8If/1L5cwWjXRx2B
KAwRpNFWnZqippJSgIkNAnRZbK6YIitU3uwzFKTiKrA38pls+PUGrfAtJ355+cQ7NL1xkvsvu/99
9vvkGcQ/OTf1irAO1HAMm4KUa4FRs+FWihc1gs2iC+HkiYVg41/aH009LaszdSng2O804QNXMSr3
Zir2AFqxGCSqdLP0KJnVT424z9YtyXyGZkC+g2Q68rD2BQcn1N7OOclxLcu3S9Oqz46VFFh23dup
x2qUWnX8s/zX8PyZLUQb7YDOuEByXyeclJbKt9Y2gqS1/YMgccvygDeys7o57mmXbxPzuXjEj2Zg
Yvs9MhEZbYOvYuQYfWraRpIB/noG369KzJ7gmNFW4Wzo2JOWriMmMYRxjjhT/dPFUeL3o742qQ1p
Mxgs5rjED1AkLbpEv6ppZ2pt9glcaD8GHJg6nMXqzuFc9g8mK0SR2ZkQDrF6VnDsO0YY+O+ldVWZ
sl5zyKp83Pv9LFafzxOjJKY4t6bLzwA3prdydUu9LT2DvD7ICEfPqpUcOp/Dn50kzilfhsc3baHH
rwuE3QyDRCDlEEH+ZYWyrUPy7lwQJq7A5ZxTETuZQOz8tmF0BZX6HfzwFfom2+bGV0Fa8H33JOsh
7j66YlMrCNI40mgM+0yc9H8e6iQRUonJ6V+RLctqfILtdz/3x5obESe8XwX5znWv7nlR9eNiVuOI
7qQmOLlClu1qOGLeHlSwKjFZnsQX3D2j1YEPCydOTuEObFJgtwSfvHNxoCfm6/rU7eQMTWgNkxbx
Fr5l/uhsUZGFsAZd06vMKGp39omF433BX5cvrDTWOFkvQ7EOL7d3v8VZIKWK+wLKwxondMG4KN88
mYYYfHVUhF26k3bgOKjpzchsPAYrOdVpgAWNeZadsg9kgJI7ntAmszQP9gDa6GcaYYW544exLTAd
ZuM2+d8duUzezTR6O6P7f/YCv3RFH+l2WjspPGqiY3fxIYjti5Dmk4YXOMjim03KZaN+8wLhkXAu
Ymw1aRSWqj+0RWd9yF8NRUUpwS2NZBTJ13YNNtXabPQEnoFsVYFuNaIGwukH85e/xPZJsX5yY1kv
a0YvmYMplFbsBsrr4nMgF3dpvIH3FlIYqjS4bVnI9fWWQ8+kYr+/FbmqOPL6tsP7NzhN/lxkpm5q
0AQO4j7M2JF1xXNadjLmTPw+TWZOfbS8YcEAiGkwa1ts/S2f3W85eMyKuGaL7eqcIJPcifnxWtyR
BUDLHQxlfaIgsBBwx921tyNpNb9wrNQcAz64c9xXWVw8ozODJY8M4V4/HEWlv3QkKjZJMK0VOGSC
oSkIKLE6NpsiYcMWkT+yogtmzGZHG+/ZXzdlgXtwrq9wvE8AXj+/4sLgiOGZabj9fPs8NHztZO4V
nV5DHvSWsWNXiJzKPSeGRKOaLUQtw7suA5QRIquCTlB3YenqiPICTjspyf38lox9AyT0rMZ5Ulj+
32IM1irSPZ2TNbxB4L79XWcLfy4X6xNwVoDGx6BprePduNPbC+P1F6CXa4erTumtLDKPQSZegXoe
d4IGLKlW7DcIFAaWVxs7vU1C+4uGvLcVkEF/i7vXXmw0i1PpShcKOYfVzcANo9PtrySMxCyuAR/r
DIg2Iv2HGXxiWUi8tfORgz4EmyA53AMA4EgrXN7StCzlyNcdWaSHqeUuEHmastDVPUWFXnLGYdhb
lDBvw76z10Vay1khSaYmqDpTQCPqIabAEHmM8M/Xsin84H04IubqhTDETVgzwHCEs3CksIosfDpI
FxTs4qzg+ZRJ5lUzjIcyJVSZ9gXjsZxhNpVt4u6QMhwA14WkQUAcgv/bWAZe+kK5hLRTEIikrZWy
qs1jJYSgwcIbD4KnX+BwqdPE2+GkeyObvNlg8vmHy4SgaxhTpb8Lk2ICt2Q6iv+EnXqDT57J51bg
uBs3DjEFjKAUgzkLw+Y9k7yzhyxy/bEXzxGVthPVl9qNCf8D5gq99d0mmPrHuw8MI1bAApb1EWdc
9VIyJGf7HV9nMT1ugTVEWRLI61SZDJGCnY02K7zxRVyMUffjKCwkRK5/efDLKhbn/qkKAKIm0/ya
8Qv0oKSryg/c5ue4tlbsthzEJmrm8f2fF6Y9cMar8CmGvlPVQ9AiYwJF1f23uaEVdVh5m0Cevtf4
xJ+f3dKtBIrMAG3eSFFw8/5p0mgQAi1k7HnV3kQcHqRMp5JOqmDKOOQFkBD/vCjZ1fbY9UTLbrC+
Z68J/72QcKiOmpfsCvu0GLkgQpRk8CABe3wpioAFwcYxhh9kkyyUkvg8KN/dUZ6d/xTDzFxesoOh
0nCmpmIQOUR5pGycxosPlJo1SRtRYnSQK/BE4M34E4ycU12eob4Nsy7dN+7nE92HU7BJBaTtzihz
tkH+whTpApTcDpGDluaD0rEa7lfz6OgOWRWZsh6kj4PwDUIcT+kDoEAYNr5zX8vNZukBoi3tHYsc
Wd6qfMIp6bBxupHkwf9QLMGp0QpzNOL9Sjya0ERvAissaRBd3bg6NV2Z5xxdKXExh9rTXqQ61/e6
Pksa2sa3yTB/ppXvfKktGgDOMxx4O4BCPu132sEfeV503BtUDckqzFOP3RumXf+Pk+uyNoZRIXoM
gdzmJbcuNl70xQppx+J2HzPfZJ9ye4t2PeN7rRnoMHB+ikXN5NIlwXXMrMnBuq2JhnjeOhfgnCBr
Bz1cTJaI522xDhTJQsmCs7d7ohh2W6tqgzghPf3BDH5+LirqpmW/HO14efKfBMnZrhkrn/HXqBRJ
lEtYQCUkymslb6NnXeo6m0WEl3zmIj08BIVV75Brko2FjmaawMJ9Hj0ywuIdqfM0FWfEqNGCYrmh
QzMD5/J39DP44/i5Su8JW0U3q1KAZNl9AXLDQyKAIyvUvjnCdccIuSjT+RkXQU/E3eSTV23/LkzZ
wXvtZ5FTcodkIxFMjU5wHeIABHh2a7+V52muM5TZDEZmPKZsfSMLs2IwyRNmeuni0NfRFhkjJIl5
l2br+5axzWawYmy1SjnGxD7blsPZhEDyfPZRIaQJAoxDDQIvMl6k6FUEKgBDqqDpuxiOMyz4N+/D
plhGKh5m0dz10EvB+QkIF4BY6S6Scdzjft8K9BVp2+Qht0mFBp+TfQZmiocUyEZLqC9yPbg8jMmr
2uFA7HMU8th6BrhkM6leQrqjEuxOOi61Fuxt6vEDLSlpkhrKqIgh8WGXHCU2MOJpVEeQc3hurbU1
VcsJC/A9UkzSpL/vIpVLU3zD7XJ5yGvDKROPTA8oMVsoJMxEKpUuMWpl6/aL9r7ApuoTiq57JPlI
oQyHsroqSVEI/44enqaWbd5RC/2XjjoxDBaEOgBt2UUb5w4zY22ww3ybH8qFXpwlkYXqsQIJpQtr
vTygk/0qs5LmNDskS+YQFptP01YeZUzqSsbLGNz86hk3BEoB017z67Ior50hCZy1izDvz8OSchFs
eCRNd0tK/AEcA8dCTTFSmwcy62SVwX6S0AgAllu2bPNBErEarRug4fi/WNxB9mbQVgc2fpS6Qxnd
PfkAFRoZPByuXiFwgzA9VgNZnSKZBmzLqfTgUdVeN1cNJCAXF4BuXK4D42RYuZrCzPeM3LhrydsU
L860HVbZxA/phK7dLKTcAlsbsrBq+SzgZECPPu/4BvhIwPnoFc3evsO8Z+mZZNipeb+A7mJD6zn0
fvgoaYtR7LWMgD3QAC6nYCzlHPL6w/sGuDvW13RT9R6P+5J8EGCiWmphvRKfocvQxR4fVXc7m9Tb
LxY3WrEOCGRAiCpfB3paboDTv0vGL79N2gEIKgA6wPxEMzyoU5/3GMLwCCxs1pfx54G6lzsLC5K2
saJ7DEi5VmLzPeKHJeU2/IYdceUI0s+KXm0UfYqCzOePKA37Hpbsv6RvFj/h48X9GIdHvaSCJFM9
RjJqDLKeso0FlAxLzkH3SKs87r9dWDVVs7GtILk+w+bQHiEZ9l6L4hV4Zgn8Rj7DH4E5dBNBGhAN
3MJG4pFnWOGefq4NhEpzswL/bW7o3sqiyO3OXBT9SzMMlb1gJwsGzhei/x6tBhwI5UyQHb7wNbAM
YOfEp4Xmfr6lNgOtnsxXQldf1zx0pl/AGnRAGu8BWx34vNcFSDEIlpcYZaJodK9PlTRfW748kNPt
vuf09s7o1QcYvfW46BkB8pIAM04fqJxLuAvqjFPokvWEZj3FNvqvJ4E3fyqxWdldiddXAyvcEMQk
do+BVy/SKjwJfw9ITgSW9N7PxJSHnhaBHGRPbja1O7KnrWH9MC50bMbOZTiu9MPyBENRY6Kranag
UA6XH98k7+Y2ypKR6MkUH6GSxXME8E7i0ZIMONnibmb0wJPJ8JvaMpABlY1u4X2BmcvrcvIuVGGi
8ARl3+3t0lAnZhx9L2jas6YGp1FxRbc+P2t385PQC3FRjCuG7fRa8hmc/5s7CrLQc9zVacRD749l
lmWGJ0HWM1gsT6dUwDuYbjYyPBV21L3riIiMp6FCjNgZlQKVhU0ehEkHedajeqcCVTx3ed9/2Uch
U8s/7AOdhGaDNv/tuCIKNx/gozBopqxcQptdZ3WwIN/BGU0Pxm7UeuHYAxNZdRIR/vm+ZXd04klz
0uqt8aCy+966TyXGmIVIUwbeZxngLOepxk+5gHTuknR3afqZFGsy2hDIMlp0JW64onCU4+xjjWn+
faXVuffICOsLBfh5WuMm9/KgFr7flqcR8snMELOA1RDIIX4RE7XxTsvruXs4xABPQ9oZYUZo/ktt
9inKiJOodpCHI2XmCNVSeSh5Uk7T9Ogq2L0NDycADREH6TBQssBmALzNP+iJkm04rJuyhDYF2lgS
OtoZyBDsF6B5gzZYN8J6U1g6IPplF2DvBfFkLrrpIBW986EgvnSLxChI/6cp2M/+cVFsm1sN3J89
LP2Jfj5F9xXg3wsQIQUHP0BcYiPx3VbIHPhuEylqtnCnmTMndL/piK69sqh/M0c8Oz7o+7eZdmzx
oD1vve2EitFYofCM5miz4VqfJ2DGGfM2AUrBAcqzoBfm7OHskNiQisAktob7mLiXjdZv4uW92Kp9
eOzPv9P8JLlFzMu16g1y5SNOOW9C/AmtNsxk9h82PLd2e3WYytIfhyerId8cEzlWYYXlAgcwefpM
W80drqFBMsO12rEyItmipxiY59Zd9JzBmJfERj+FxsIBK+AUhsJWnn9AvWW0MILO9SvxMtZQnsiN
XUNWISSMvIsuJ8kAZVA8MRf0cvwOw7b39vuBlXY/apqZwPAwc/sVb9YXMXTg3+F/MIWPx8i0ZYDT
4CqhfKuaIhSTRnP3TxgV9Uioewm/96V9IEHFUMuBp3OeIcgyS1gZ9+w5/m3g1toYwvyXgbTVWsk2
FVApO9iJsFMEAcCgWUL7KsUITN8r9a1mUBI0wOFHKpnpgIf1hHIXbtit1Uqx5mq+J5UE/BR49Lwr
CNl21JMsPWvX6X1etYIwfXEVeJRj+hxjdhYHDY5udlqeNas/BgmhWEUR2nffoTcLNQuRNX9oWhlH
UKECvJ6kgeId1c/RzEFgYNG4JsjGiRJIw2vj64RWwwd7LBgr94szeQ0CCFBCebEVUbRIVxZ8ODEq
CmGUD0NI7QN3imq8jzZ6TUNzucWlgMSOh70d3ZS9Y2TgjpsP0oJ5swdaWRvWZCNz2jrljOBYmjtu
3eyelsv4bm3v0005ifJYu5CDNv/VKjwLUtxdLk4nyHNalHQhQ3N2ZdZKq3a8vLDfo3Q1SffN5H1o
VPXBGp2GkEB1aUHKELSobD+dpJ0CxO1oEC1wGPdXzxWaWpDQEN+UbM9t3+hRYUXgeVYdftA1PBfe
IIHaWA+k32unt2+AJWKmQMqpu0OEfpKAUNvK35+Kl5jl8VE1IfTQslhpkrSUlmz7JsExGc+JlZaM
Sy9AZNp4ePct2HC9F8Z/BqW9aw4bDDduDMioljxlXDRX43C9+TnaMcuyDpYquTGkXxl9OXaRIJfN
2FUZzZdq9QGfW4Z+RsdlggfjrEEF38nSrXz2wUXJZqq6Ucd9yVGkJ6DAQhkqjTndeSC6i8HuYhJ5
vLKMzO6FC8+BrkAwZJYyTNY7gi6SFm1S1WuoT0sz10XA0E0dUGy3nXI3zEd7fx2Ccq/XIB6d3RUf
OZZWtYcCQZdhx8ilA+5OGMmnHTxTmZ5y4CA4a1xpNIncbIzA5jzSs694N2qaHOnxodihFnZWtoGa
6+PifFwiJ765h6GBQd8J518uwocjxcJ/N0ah8JSg1NYcu9kTM6jN7ulOTfP8eV2TuC0WCZBWCcwU
3X2P8Wq6lnx+a0FXXk7HTTwa1EsRxvEdB9G1mCljIxUIZwQoCgErYwIlwaJtb66fGUEIAHNDnRZu
euEb3qbIZzZQH1YJ3HEnmCdX0m4zY+34FeWrrAM86fTOWQfCzH/5NmnsS9fXgSGAFLdAKbPG2qLL
ZHDgB+37/I8AenXGsruwre6ZM2dOZPHhMMtr8H1sEHrl2IbHM0nQX5kLhdofHapivC+DC3U0Iczp
RWe7zA0SWk6tT+r2MZSplESaOyrAZfxkco356ZFWa/pbsxkqKQoYGszYA4iw5p3/eOXsrmkeAlnI
KeWi/zoC449ACxKFqG8higkmiD5aEiMJjjpa6jJDW7MF9i89Snufg//U002KugjGep5olIIJSNZ7
TgKdlwxBuWFfCkZVThCYN0/wIaLHXxhtE+5+Cd0JIHWQFPX43xS1vW4zH6u3OwYfl7c9SObvEeiy
5xT9HUblt2HPfXbDZL8fASLNbgmbzD+uyYte0+g60JaqNqhLXwiWo2Tyz+VnznUynccRKOp2EAMa
FjFOzd2BUUFW6VueMiqsf/s/CJ9i1L/K6wMV1Lvwiaq75EbOh0LIUks6WYvk5XUenWNz+zHXEl9S
DV63JgVtpDEltdIuybnevHpCGlslK1Bka9kd+tO45HwAJLyYcdaweIlfr55gjvju+94h/LNLAVMT
i8BLoC0yE1CXZJ5EexP5mOjgrKOVsb2kfuZOYBSk9e1Nxma5ezg7dxWtCPNU4b54AxJZN2YkpJxk
IgJ101iWoTvIJwGe6TiaQqIiKnv5RaI+o/xgienk1C9NL3N1ny3qy5OdLJ8P6xeDXoCoFvpPt2zj
X0udjPsPzGGvHcFdq0OpBtrrgqDD1F4BYCmaX9COyje9hK19ajT1aDN5rgFwHL5FurTxgHmyIGqL
rB+f8mUPqrqjgnzXQYDQVlvfdBV64J+awChIaD0VWdQzQeT4ZN4aTZtI3SsY6JOGSHEGSupI/r2L
FpCrH0sRNJ8rhhs33PDvB4lSxCYiWFSswl5uioCH+g+1a8W1CutX8E5yDEp0p8MqJqFjE3VQ7CuY
nXoJ7D+eEw1c3D3Fssyq06Vul31XHxLpealv/x5gxiWUDhbOz5Jrs08MBqOGklC5zGUPuEHZBZFI
R5/E7Gwt1BObVNeBGTg9G8agUP5icpkJG024BIQjxPoKiWQSWDUGzyk6nquiHrKJU1tROTQ4mNmd
YRoiwTRp/g2LOy5dhi3+Cuw6tBp+BAhZhm5xsW4pQyy+rx6D2TdEIvH+AklLF1jZfcWqlbsl+HX4
5VdzdMWXMs17h/5/hijNwlpqoaxZs0J4pQA30NnP9rai7D3xNHhO0IUij7ox6tSKMB6/Y0zGoKB9
szNivIi2F1ktedHRnkSJO0ZJfCZdKSSn28tqbAD1YWLnB31AQNZio+wcUuEBDmIpFzg7XXP0oI28
fy0RjwGxVuAaGE+TMDoAWvKLWKBMG7TzThZK2opmox5IRYo59noizlWl3txGMzOQNP/8AP0QvoDw
Y3bx+ncIDXz9ZhLYwi3cDoUlZ6Snz1ep7jEZX2Sk7VnmUOY6ytFRqRCqg05VmQsL550LHOvVzcK9
Y3YN2lte+8/FdtpYCxahIKBV975jeIXoGrLfrDncN6LACx1A10+dsTlpQZsPmtPzdQfFqTKNRxHt
PFPIX027VbKA7VK6hd/DZKh8HzIxQaXOJDUwiAlEU0uEEX8LDaxNYzX1PN5Mi67ruYDiP6lriNQB
x6RtE9S6/zI3hp9UonKzNXKS5OU0ADJMYsqBf7vzfpFQnEwiYbVN8s2dAKSu5r+wrmIWhLBcHQjm
fB7dK7FnvcRu4m3sViYm61I+0rXr81CqDv39TgmiTpcNR1RLj0TqXKDrRlJZRiGgS+czkhv5MqQt
Mf03/mh/2BLg+51ordAZTlossJZt4inOLRyGXp0orOh4ZTaokv4Qo7HFHym0oTIivex/2Jy58ilf
k2xpfdmXcB/MIwoOvZXWrFkQbuyCbp+VrJPj2j6v9pOBS4jN8pxbLNTFUlFUYfMvs3uuZS7kGPdk
dbeKKXU/W41hAk2zKx7pZKyS8zsnTuvfRiX9w7OeFhPBYIRzbKnOeDyKl5TaT2Swtzir28o0162o
cRgCWlnbLraLkOs3XQ8Cj3xmxCXVOxpdztzSrBo0qOCckQY+rsovmeA8JUZDD4BD2TGD2cNBrMbG
zUA69Cv5jhgGpTgdOUH+jfAohui14ylcnVNESkHpIQQkqATAaFAqFxdfURZiTw+X43DBlIRp2DY/
xlovIahuOcXoQ38oBqMxDhC1BWr5fCwTxxF5ZLheHesuykvbFKWe8wT+xcPswICvOWxC6w0TJ/od
XFiOttMEC35zhT+cx8ar3vVjx6qt/R1EpfHA8uTHqTM7oGpNvGYOajoQ9/vow8Pni+QHVDf1Mk2f
m5Zm89I6isyWmKVf5YlJEFnIt6TasvFL8j6CwQ3essAk5mRdlKROTaclCMbJBOAi1ZUatCdkZ0mB
X48bzCZX807FxpWN3wapCacbyD3ylJLXpg0M+LosrL7e56i0b7t9TZJe4GYwLSxC1/Ct9BAAUtao
L2rotfZGE5hmnAOhmmIu3jtYplauW5mkM+pjsVmZXrN95bW3h5dS/nx3n97OZ9dTz93EnxAKM94u
RcD8FIspl8LzCFZiif8Q7JRkavaw4qylV70x9WfB3u4SL8nTRdJFnvlq3OKq/KAbSIaOH9YpM/9I
k5WfYwuGQZ+zI3YHTXoC1hUKAl/OkEZbILA1dAhOqWh26whMci1V+w6ROGG0A4Nqi8Qdu5ldyOxq
lPsWTRFlKmoWG5bkC/HIfgBKOKkOwYaKOZdheDiVoJxULrGdj5H0GMgrUYC/5n4c2XIZdY+Q4yCQ
ePKKhSLkYd3akRs6bWEw1AaCf0B/2paGXDvA3/rZzNUUiJllMa/1g5EY4A6D+SJ6firzCKAXLJKx
mvzmCdqyHfM6HPeQuMtf0ffUVDKzMEUkyhJOH3oiSw/h5jDX7VToAjmunv9X+XIQdNDdETgDBPk3
5Ae6hphMVi+OoHgRlddd82fDwNPVR52OnarM36jhtDWWHl7Es4unuW5xzNIxxoPNIRuQGTYG4SSP
4uTlS1eiuxrTn98aKQ0ZaIufjiyS+Dwt0Noy03DpBhqdtu+jjR8XaSj5p+lNtnDGIFbL2Bnza1x/
m3fI5NhBp8TK2Usv2J31mjBqjU4FY6l/mTjrszJkCwWGUVHpXZrfmJKlMZPuUYN5fvqOhPJqbIJG
o6cKlp4Hjj2SCvmeIiJX3QWd/XmO7c4XgdUUI9P33zJtkrjqChVxQTSe08sMfHDxOvtp+5FNhSfM
hBrVVehKdeeHKj6htxzqTj5LlgkKKU6eUWZk9Uidmsc/WIkfGlEel4Tb+t1OClYc3d2o6ESjiSJA
Ih1xt1Fmn16peUA2zy791hpfCJq5WJPlRtm0EDJ0gMo2KAD05f48iCi9AW56MFVTDrc3bsiEGiwA
pZWBv/LfH9uRaFxZnVpVn3qBW4bhlV6nvU9IlaewDrO+eVHMaw5hdug/+SO6BPPMh0TQnBv8l8r1
YWUi/pKux8dST8pG4WzNZQPM0CHv99DHM1Bz2SocUrtYjxMBDOmlqEq8NDWhCtesWuwsYwIwUJ/j
3x3RCNeclqZtmZcT1bY3Y9vZ/AsVEpGmDYXfi0GAUJ73/vkWL4SwijV+gqr5szc6zvd+eVubLpa6
yZV1ZIMbIMwepV5F0KTp5SDSb8OEHeRlkGFXaDGINAI4CIaR7xMwHXYADSts9zvi/DNHRXlWl46M
WYpGGxILGkkGo0sXxovA/5DP5gQVAxAqQtK+EsPDBnqDo2YulVulcDU4SLOqO1eh/gsXSE/G120o
K79Y8FUiQF4Ir+aepNZUOY4r+4Zsxe1Z7Sp9taYIKh03Q44wEj2Jdj106aFtRePnxnJVtGZYAKLO
td7amvcbX0xOtBmWBy7kXy+XN/tTDZABuDE+7Jl66zNdRgJJ66i8R3kFGpoiIypNnMJeahGGwmCF
4O9Kt+00wggotINnQUSB0c+oHnbh/Us95CYmDP7fSsrqvBhK4HBVcAoZO84rDjjJEL10cfnaGFj6
CHw/VC3Q9t5VTCjBIDZjG7AosazVBMlaGrJAgEAD8rPNe9ib8VLCe+2t3DXjIzER2Etd89AYX3x2
EbyVslsZGLj+KHpk6N8h+ADOWQtYXyvZ3P+uad4bFCdRlzsL5gMuo0ZfEPMo/80kYOAe+g7y/hNG
mPOVXTCjne3m1Fiprth2aUxG8z3LfSF7XVBuWGM5RiO1yF5Szk/Cn7oLFZ61UrUFF6yACqr8UgUJ
AY4/2hbT+kZoYX1ICyjitqbP/W4OYZJHne5KXLsYPpvcjnkif8Es7AFFJHuzEwPi1CiyKoX4bFqI
Ao9pFKAF2y+Ch+Osv0zLJYXYzVLoDhZ6mDKofpYiXZPtYNghEFZln9AFkqtl9Exes/q+x8jaaW6s
8z6TQOS/qeyogb2xEvJlvkw9Q40XloygbHWsoxoZgqm3rp2N2Iq8N2HxJHMi4wPUOLyBnQyDdvXm
9a/GJNRvp0ZCA66HxGf0EmeiSew1578JSTO23sYTr2IgZKJpY17zZf7jYjc4byuHrHvaQo2A+hqw
BlMhSamvdW9o4Eel/kfbMnjtNBviBPrnU2Y+7iaCYpK4wiZO7aguN35s0RtLtb3lCzgpqpwn1zs9
Y7V3eOqDb9VOGGHEpwSOYgat2NNC9BDgjTmhmngtOajg1i/v1istuighohVxGkE64xpXOLxabP0O
HQOsf2StRENKs0BzdQApTtZ45WS6vWu00XReBzF2qQdGFEgDhMw0LolkrGUopea3LR+gI4WLKxYK
2PhfQilC4a/KQNXRGDZd5D8WHfn/JswYnDgCZArK4mr4Btpha/wAmd1vNqx6Bsdm5XSLegFmBidU
09+NvHgljZmYzLS3Vl9OCdGqjDo9pc2maVRrpRAi/CKBNrIJ+jN6tjrKTQMIcQ25u4opN/3TC5MH
b797zEcrMUZklxoFmtkgCQ4H9ytjH3Tq7sI5XtlMyaxUQUuPPviGTRuhNd3dmjOxfgERbRUItCKc
6DhVNMmvyHudIKTUefdiQtD4UbTdXiS7oRMKtVgs6tZwGmws1YzWtflGyYt94RRt9JA+qQSF8ctm
0YHMJfnUgIqvVKpxgNJ6ZlWEn4w05AagKJODDZYoeIWf7LTv4xuD6+AJxgCboxfyMt4FZztN5zNx
8ylZmoH+YIz7XwKhCF1gVGhp8C0niBGrhWCjDvpU6IJ7ZuZ9Y90hX49eyz+Rgkr9Whh0yR/4oBNg
EteIKANqGvB0UTYrNu1iE5Nz58skWogMhNGnIzJ8DteRn5P6225EqBaGAD9xbW8QYqkwKDNQytxa
a50/HxtMTbtHMx9B2ACC2JZLtSFIOltQQHKl1h1o7RqFnJ+3xwfslni/mob2oWvX/ylNMHw9gnyp
tUIrniagBdZh7cFr/XDic2SLHyfy7XwzLXsDwhF/6Ne+luaWbNYQBbjMa/uRCf5GxbG8/9Bn7bVt
+oPeAMNjI9vAkeyxbLU9LG4YAZDLWqgesMeXa/rxFkB7vF5T+kTHnkacQqNHCfm518LZMuo+AqJT
A++KhazZTUc0OJMUnXMN29DgOLVlnbOt4wQWLsKjtavX3tQYzQMzO8izlwNsIM9HDwmKgzbOf7JH
zsJZKp62Ro6XzRSxNzuGUNjKrD2gWnjkZi/tVczo21tz+dQH5OBXz2RGOljndq8VyA4cQHotzNN2
rE3qnw4146NGypHHB3+RmWIlJqmFghQAf8FmP6vZP6vn5ZXKKsH1jHvWYWltl75QSRy8Fj+UO0O7
83z2WlGviR7ZUT4VuuSqAWOZj8X/TAUhzHM2Nk+bb0A9vWk91Il5lqKfLdPb85RQ1MGZO7H3Egrw
Wbh2iRsTtRpdk0NPTzO80fUaVxbtuDpDbjeZCRo+mssDEqUeVrmXQCZ2+2tWV2Rz1aJHJ188HWCl
1nCSbjdshL6xVuTa7Xnmn0PowjnCr+YVq/A/xJDpqNmOjE57V00x4hMbUDqV5xZhwfWxcRVJ8shy
JMdeMvF9ZUaQBNPPsJwdlkDOGzwLAaTmP06E/7DClwT85+ynoDCNKk+6k4UW91vmX+edcLLB5lkg
UhSEag7k6T7QKRwGg9t3MlCOzfy8xbQ4GVn4giPLowpGggZGt1FlilG1LCY4y1cEP8wJj1XClQIP
6W2iCQIm0a389eTAIiD6noat4ZcHTs8Zkh4AnhUTAuyLHFnoIOLyIui838nLKe9gl/zNuvX9ZswL
OdHf7azlRVz7O+U1dkCVVlVajaw+jeCyFgARUG2zBtdtZCWwEGhbk5KniEIRx38L49en+raBsdYt
xEaIsQkJmXfN1Hpm38a2XgUF2BMRU45GyAbFqHOAYKbRpxiMmE3SyBuC/8VAkgoC4TKSpWfMauKi
4GUOA/Ndq+QFlldDFnvnZNYqMKVMR/v/ls9b9dpXqI3JFqy3h9guiyx1hqoIzEy3ZXzEeGN5QJ8J
+jGtfm4Ap1qBeI6pmrTKVmCddxWZsjC3Bm1w2ABGXaWzZHMrokCrGN7ZJmqfqCdiOhTTFu2ko4BX
SoMdmjroN5/D5b2oE3deZCVOEDJ8c6gqAtGopgRA1nMQD6RMEI0GeH1JH7pK3yYCGQQeOtTSukgn
HNKglt627ya5C4buDxjSe1W6dBd7TTIfKF1S1CRz472n/hpCawT+Z3V9i9KfmoqyV3mgFhkIl71p
hZEaz5CtvP/SnGIoViGZtj58CAkl4/JYvURUCFzUbojn6t3EjpSoDZ3bFRQqxy6bu5bmf8ks96ur
QbmMKVj33yh6F3wY341DLyKOZX1sovGemLL0tb0dHAfE4EW5LBIBRIFI5Dc9G7nOmdUVis+rkEj5
W52mG7FImBL7aRZeNcbJYb0HsfxC7KOs+ptsZZuVmo4W8lEuJrXtsBlTEjBqpymhXNs0Bbt2VlsT
pq6Orf2ctJZQ/DQQKTuKwrd+YtfNp2F09HtXULJKR+nAePj/mIcbZvaavSGno0F3DuHN1B3IrNqB
1vs1n6AF+b+3MN+14wmJqcS3sxXD+jerVteqV2vBleARXRD5phY9acSHIU0kdJt8+sgRRMY30NP3
NifGsmIb3EV4n0R5AaZL0iD5HUAgqIvJcFUTPs/QF4HcXcZeNinIlERVroK53fIri3w9yVZo6ca2
6bmXYclMnrkBDhtgmqYan2kjYcdD6xhkdaxCsRy2LLR2slkKlOPJ3kO5o2Mj3jlussalSyB7ePXV
HRa+FjGYKPUJrwd+evn/mq3OegVznjzcjqNOpo9hZC2/GoDNqPi2AvK/DQ1QkVrf1QCXHaChnEdh
8n0Ay4fpx1fmp7WxQP7s7IRpWI2rp4fgbD92hk8l0zLUz9ALwkCOcgqdVbMhX99skA+PuXgTFZ1c
6BDv7Avmqlq66l6DyMYci92xcg99K0Hrsy4FlLerAW3bpEQUaCZqbsoB1iVjcLl66cAP5HGBKoQG
qxvmjxXRI24AljY/XVjuIumMM6IhvwmLXp4v1gqzC+p2HQ1C74m6bkNB08mb2TkiDEvenLFezmqA
we4rSGzMnV1xg9444jpRzynpDPbaXSkC8pQOmuK6ho2nPTdQx90UN3veujgNpiCAK0q7RjmEy0qk
lXDgirxYJcUH2XDbfkYoHj4hfaNiToN+EysMNm5VcDH/vqDzRqYEwnA7mC7EZO7kFOVwkiFwfD2U
278zvAWoikgw+Tfr2p/+/qPMhbAhhQWiqLaBvvE8X+ElLzU28A6DyAec0Ie0jT4Gayswso8RtuXT
R2Cx3nREGxZ6lFHtNm8FDhXzc0D+87rzET1flc+6PsCAHDyXOjps6t5ukk7oUSOTiKtkcEOmbEWk
hxBvVANUCAlpeQN5TikIN657LeJ0m6U6IOBSjArbmzSHd6yL8WVPRKXEz2sF4ltHQh8m5R0fpwoO
7mmELyGz6L9KLDIKUa5nB8gigPiUo9++gRnF+8pCAGpe6gRVLyQKxcDa0ciz5Ilb09+tRBC1gqlY
8pKIcznCxkCH50M8g406wkaUXPEW8hN72O9N6ap2d0+aZvcZPWOvXX3HJPVBOfpu823P3BzS/LG4
Zl4mjvyV1PHyFfDysQtWxpDieajhUt45CWcNIEHodpXyLmFdCDyooDvXbOShWiK37bg3h5hThe4O
UXw5XsRGIZtbYsNzVqUrhNEMhcK89ewBJExQzRsN7YPKP+fjyLRTsk6mAoop8uDPrMj2YBp8ngrR
BJQTJistuAr4aHzblD7PggNfNt282bokOrqs3IN7b+AFrrTvCOQWoKeh2EuH5cPu/KT0hQLpAiqA
E7eVzRxgSb3pvTduc9Iw+VaX5wwsFMrfUMnESgdVc8ENGYyYu16q5bG1a6SMyUdFXfhB2EHc9WAF
J3wFG74qbNUQmnLP+KCOyIJv6vfgZxQTUh6UEg6qPIg+VnPSp7mjA+2N/BpYxwfV1ZSJvBrX3D11
0J2rnYW/10MP0p0v4JbfF/5A16FoW/8czjgQws5bUx/bV+pMamxWAAk4GvtjgyBOC/ecveQ1VVTO
OMfgc/PJKo/qz7NXZ4hd9lVxIyJhZ3ovllnPEVqVnXFsphIJNNJ/Cr/BiwtZoFJnfjTwjYRAmA1A
IGLQdQIPoFGCVYYgX3Dd0lQk1sNuKx6FKrYm1OustTg4pGE43VPw0qtqA7Z5c31ZzHa4EeSg9o74
CGqXZ+d8Fh2fmP6SAscXzPWw7O9QUluH5zpT4pNbLGuAIMAzZPgsfPmcALeq6xxIKNs5YJDCmbX8
YZPXbsD/QkbsOOFH1J+LSsb5cK11YBJ+noUF25ohCqgqSCf6JbmTEwqNeHl9uUUdxV0eRsh2OTUc
pq0ZjW4VTXZTjdbPQB8reFyt/o4xFP92uSKg0qmnQ6f/oSgvT6YmEmWhpYjqNEtN4H3JjshHe4E6
qWrQ0GiL5eGH3YjKdKT1BTOd5omZWF/MQ51uTnfRsk0oWg/gkOKSE0KpJBn5+RpmCCMme+3Q5k/i
HDfcu1km6PMz7ABT25ewNP0BcbP+oQnhhEcsvj/N6uohPxOwZq8VvjWTPJ0ybCSZNsF4VcEK+vis
5FqAJ/nuRY83haqFSk2gRjsSbG40NFtooKD6Q2RGZ6LxAsHptIYf7ON7GPm8OHgG7DxC7/iB23MX
3dHHcCn8SyyqTBKFuqERyL73G/IAG2+tpIK3x9Ug937V9F/h+Mx1JXfTeVhaSsyNtv0oRa0ZAxZz
S6UGVKicjTgLouCjOOt7lKD5QTV6bWnxHtIPq9Z1h8AoPBJMcX2KkYrnOjbXB4b1Ap1wzSljjuYl
UOpSTu6KXy9hwd0QGAs8RcsPkw4e+xONIabVec3wFBjhddrnXkRQepPpE2AGMlchIttk0a3Lwbsx
8zLa20Akd07VcmqQLB0LxwpMa1ZxYPu3KHQt+q071JO4F2Nd4k5GBJiyVAFnNArix7ChPsBDcO/+
tPiPJV3zYd35AuRLe+NkINOKkWlcmN2b3/C6TB7Uxf/J/FbUDD/ck25Nqo2GDSr3dgxsSG+u74Oy
8Ns0gz+PZ7L0W7k3dSvozZPyLdU6YSVNNp53rpJ/naVpwLCQVGXSjxJx25dW9gH6ljvjxs77nke7
Nv4hMmCFxYhYBT69N/buS+M98dPeEGub1t1Kt0x0gQMxKR68NfvAu0M6K1b0/f5hDaUTFRH0Kg0D
sa2J5jWH6qk3lbgXmjxAkspZ0qRLOPxalBx67wW2wRIFveteBRUxZWcnTmX9v0K1dyAYT8rH6aQW
3dFJJz6BKM6plZPDv4UFqbgWiho03kNku/eP6yRusZzWnu5KCXvI1TsuabASwZnJvPI77wZs4oQG
j9euVmGWmI9OXwIEoSnWP4Ob4Nd09chLtJpcWTL1T6EsYqyEv5tyOOo40t+3lLyl4SJXFgyFwxTf
/9dPuqIn5ak0Rw5qJFZGgmntZm57OirIITxw9uhLiTt37CXK2BniMwC9DR5PXW5flNMAjmARO0XY
sKXGrUfJ3E+vuFpMx5XcJDuTmZVi0APx8PF9pmyvb78+gY9ppCcI9fa0VbystPZBiTw+2vd9ur+S
9aOaftc+HdNIyd8S4776TWKTrO4I4DT1vM+EByg7q+C75zfQ68Ptfkl0OXJiCygVKyrL4DavedpM
DLC7Vms+/6UfAuuygs7L8QvU6OGS5eZZv3N1m+13WN1AV2Uw6oMuM9q1+/3A+/Q9yRlUFTywb690
KrJW39FwA6foDDVc567WnNCfMYymCykhcgfHLYeJK9TBYmb7S3ZmG+mz6dR/aroHdNwITf1Nv7pV
MZ7WVe5axx74UuwiwLHnvy5FJbDzTJJqI/ZrnWNl78ATpwS0cBRZ1PChy8ZhgA+HfapjR2AIXMef
LWwfylaXpDRkOZJyzV1jKROS6eMEZPzhL1k/qwkn/Tsjcr9naQ1TJqGFUx/bULE4d1q4+pdebD4Y
TNA8xGYtVoPoRz7FKDvC76OzNnaCfKRcWKjYYzFy6Ve+SVvYEdYAdxoleP6GOSMHeYUp8Lg6e5c7
6Gputmyh9KZm4cFUHJYaF1pa7Xj3woZIEfkjlF3SggVNi+Zeb6a2/r2h2ewbNYCClV1A+E1sQvrW
mQ+5Em1hW7L4epMWhvQ7fxoBA0rTrSSO0aRXGVUlqFV38Lcwfbu/jziY3NQno8LLRWY62GVBOc5f
X7ezKsXHIjJcww3olgSHZMm7tCnERMrwrSJrIIFavPirgof2nOW6d6qVTcyx5/L8212255eKvy9a
Kwjris3hppjbGMSqQNRpN/2huyPydTrF0MUQK3Mwjy8F67sUlbE5zI+AFrlUhqJNkbeyuwoRZZue
ev5LlEE02g7vMeaIR98WT0E81CU/ugmaLoDsjL0oD+D7DlDB7jp7mrv6Y9K8wyWqLQyuQiNV4ium
5ODEDHTFN5tA40kFW9JdRCc8Cm+ebzyqWBepGH9+ugkZRS/EaB/5QCaTEHW4WxjEiEQ0E8HXKvom
Gbxr8CYorP+1N1/MmvRSKCk0O3R2e0v7JmxKFfH28Uzi8ms1AQLRm+4VeCr523aS8BtyAwAXFYeU
ckWfC5bDQOrDfb0Qn3zFq6U7NMYB3KHatCIZN1AJ8fbAQSQSvHuEcIU7zAfyrasgBeZENsuelS/X
QnKxhHyGakzGHItZFCdnCeRG+0QSItA0vFrbdLIwmUHKXERVXFigW793KwUspNfdRaodXMATHle1
2y/+svhvXVb4fzEvLNlX9sGlwBjxVy0wIs/RPRsqqHh1LNAly9qDX7aEhoO0sAQx9h3i0BPq9nTs
cPEvyH9TwsQ3ARl/GgCMA5TdL9X7ddHFUDGi84EmgRtcXhJQmO6aeL1czj/5/BwMWcH0kXc2KJMA
TaikLXGBZamu9MJJfctldDx92EErJLPDuOYu42RhwPO3ESwYrExYJyzWnUxwI6qkW7+zf8zrpMTW
pK+/wD/8S6Jd4uF7t6H9aaky7D9PKwN2WzpprIGpiHMkO/sgdJTRgDMHsPl4iy97u66ziRjscfSw
QYe1Ezx5JTZJkhQQu9EcG6Fr0vff9v/FitJxz3rYna6IxikBcgboFSLKkvkHQvNtZApXbwCGBxWz
pxfpiUEFOervbF0RWZ+fDHO1PE8guVvYx4me4uNGidvDJPXPFAMF4Hd9jioa7es7XTaVzleMPK8Z
uH/R8TvrJVb1j74klzaiFToyeZaUGooSql3OEh16BBwoPfHmu85OdJCOa41FeOtN5rRmzuS9kkc6
iGkIeGcEJGK+t3UYzQNuKi4fLLfBFhVWBsmV56Za3YTOd5bKnzvwjmJB+xjbuNUSOVLcqQjk+z9l
dNRl8TaPvDQN6CSnvxMvY6SeIgiK6qpl3OVi9idlac5Z5lHlHyKAYwjoFw1+wnqaeUO8KsoDw3FR
vADddb3Fpmo06oxm6ZQJ1kdVThB4bvhKnV7umjbqxg6RYI9NWfmozhtv05IeSXZh+AGQfrvPL0lK
Lm9etdx/95cTaoMuh/SR+iT3J6CnVoF/BFMNWMmXbwyV5cVE10KGTmAy5pEjxr6Yp2n9684IJlPQ
K7pykydRIp3WS4Y+MVaE9if1jN23U+V2TscZSNAiep7fYK9Tblh8nT80NCo0pitjsiJyUx1DXjic
wgn1KOJnU0b7ctN331+NO4F9sFkoKBaSx3G/ZsOeR7diDATiAj9lTjDV4swRuJWV2lZu506fcpwK
21cY9sNABRTTcT2LwCjIxqlZVmF0sU16uK8FeQdBSviL+/0TarwaBOpMwBGQZd6JpHWhRIbIas69
DRMZT/1nPhT4KA1BCE+1Olf5DQmrrYNF2DhrLfc1zP8/dT0YtnG+/BbsADVF1Qebx0TAh0Ktz19B
GziZUQN+w6ap8aB0+TV6SnxjWsKb+iDyYpANbGSQoPFDvryJLBekYFjy732LxbOlelOM3q9Dh2Pr
yoYBmeCtYmnr1Y52RxWSt2YYJRbpP+svD20dsBTlpemjKlnbIK/KlN3wuLQ9fwFddRYFPe1LwYcF
Kwmx1UMtqVwd8LRso8NhHL58n1JMX64w1NdgrbN0QPKvuSsQqW9RLtELCEv7QKZ7zjWgPYBHUese
2NAfFDOiuveFfc+xqlayITVesc9hWPGf3WvzniC/TbTwS0+wgYmmw9+qg5DFtE0fXX/4gHY3rJi2
urVQctXW15E5N44rtjZFXkcnYnhMHgAfz9l7q9ryWey4aRsAed7I1viwGCQK9uEFstuOzY8HEdpe
2XEGdvDpMA2hFOQSkjb4JmTbcjquafHA1bAT9sTp0iE6O+a3rE7nRX+SMrQZjaj1XNfgDxooMlNe
38+AlNnBVqGrotEERWUHvyvVqndFlSobsqIb8h2AqlJfozpYeUUyjR6LEbJB9t3PKjsmJB+qhSUR
/m1CsCxdj9NHMfA3zsFuGjZ83fIAjz15tceoFRbDm4OLv5NrubOVYlxNaG8Mno2v+kmNOkaStnIZ
zBQRphQnPogkMX4m6LbK/z9Lb+1FaDg055U+gcb4+pWSSVBiNFhRvK9Ale4xtuUAwLRcqaft48et
3EqwOqeDyEB8J31NAPgaUviP7Lhiy/85yX3z4t35N+Rla2MlqaYi7fwGHIBICey+JpwAjR+Q1TBX
yU16sff/Po/NEpEPvOoOodPgjWApVe0lUd7G1Q3EqCTndYK63kw9WLI57X0/5+9cHoMj7WEPSIel
Cf7v7QYkmhNv9an+/+vQepWpjw4rbapT7t80KCamBS+c8zDd4jushRKKTlNjGNJ/GphxbnT+3jy7
bCnHMJapxA4AN4dkaF1272Yon1VHyvtC6WukOBUgaKvZTQzFbqLMlfKFIAsQNJhWkmiH29KxUKho
r7DmCcRYvFblvGLKJ80/bJhQtEJrZlc2LJJ8mp5ObJPRkFmfd92qOX77w18Gc8RIcr6LhRMhTIVn
zpNAOQbWDIvy9kdtTzpknd6D2S/s3GR938N9r4mDSI6exAdIulqcZFRpQ6RjaNqe+eDf/enkbX0+
s8HZAjbtQKAukA9AS1Y6I0QMPZezrztszvCHQjmq0G2VdC01PrltGkgta4vmGOfp5sHllB+m1q9s
rclZcmVMBIkADlNVcy4ArhssdfMwrPpBh4e1i0CCLG7nZnsbC8zPQ24G/N+nz34MXbeLssfmRgv8
Yt/N7+V0DaZ7sXCMSZ35pFL1trVSLlZ5xbDmQvVMlr0IswWKRKT7EjEQCFo5wP7pPgEiKx0QChdm
ASdfQf6FYfI4m4jZkKQxJBJuLb9RriHffZXyl6RWfaQj4GJ86IyIdd7LThylPA4G7dNi1GT9YZHD
xPvQtOnWz7I7dSY0Z1yOiLPbLqiVxghUhOLgcnJW8Sl3Kj/P7JR5np77VHpi7o8keiUXH5Csr4Mi
R6OtefZcWfkXZLvkRA5BV5Jlg3qAqf2MvW0e4KI06BrKqDGPSY17dlznvdvSE1nMwnzwamWBC/eR
vuj1SLH+EFk/wxmQocZrecLrx/6q9MwtZU8abHXyiL1SYFRM8vvKBHSSWMPzEdgxnyZPLm2X4ItQ
4oiMePHo99m2CkTXrFpBSlDvAwpd1o458DAVswwOTb+1L+FMTFJPLB/r3WlwC2gVITbQqtkgacbG
hKPbp3z/M1okp9mdjqC4DlRdD883z0DsWj4RCr7Nfl26ppfbFAhOR/+aJ4+GTUHRCNt2kkrXckJ1
FCWk9Ap6bV5MpXNfEL4cUWnGOY45wvj1gBCy1o+4EG/C9iWYAi6JjR2agDUMWiZmssQ+GmfOIiOD
bQUNd8xp8bL3GwBVpmfT/MP9jLC26SwPJwRqz9G808Nvr79HFVYWHQ86/FJe+ITD3czZG0VchLkA
oFKRJNOG/qOtAovKJ1JgcKEsp9Un/dY5lqZJjWkS7zTbbooQCMXCxG9WsJaXhRVjLXyTFFYQnEGY
uDmprQ7GsaT1hs7dNvC9hyB7HpDSKJbuUGPS4OCj0JiqohBanXtxwsnZFOKSMhQagjtS07beuZUh
YW43wrw4DECs49YkxicVOw977d8OSDskYUzvn1Qqc1d3H978vU6P1uA0+eo+BWT7iAGeRa/b2d3p
sN69Y872uLcUU5VJoEjPUQS435hxrANHEZhUfb18gnesX0Py4iHKTiRNjLV4wBQr0IQbOGr2Vkmd
qTP3jp+a3mVx4RJLb6PqQAEzaqCf0/z9FDbJolr6QTpLNpcJg5ax0NH5gBWb70yHLMbOCaM5O09d
pksZZcyw7lTTSq7aZibUfNGVSxc0MHw4hAQ+mxCa5HOQbml2ne+bQmNKmHtrFPlcAKsdM9+nXurg
yuOctKnxFVhQbu1NboTKPhrfsbg8C/s2Po46cToqE+JQtDcXkcmSSV4FQajNMRSNbEYCh42qR+Pq
S5/ken9ZeHJExrrW2XTQZB9UdR7AVSCXwIobzLZjH2rmUYO3E8pqAV6OTtM69i+MVqG0jYx7sCEW
S8Ob7tL4Mg/HyttOHYT5utFXW6FisyPj/vM46+sYRwedzrJm0RGbFSAbynQSUcyZQCw123wYHVDf
cqeUreHaG32qBG6+ZvcgrqtKdBFu5c8+ZVXa33SeVU2S/xKY7G3VdTe6yrh/0EAvVmTyyZT+vD6V
bwMtzjTXKIRDu0zk5NuDhNs7DS5sL2KAH/lv1qLjDtf6f4pqSytNIXh3XdVM6eJWLYFgnlQZEOtE
0UDUho2Fv+KxrB/KJyIvTgJxca/M7tcLeNCKzXtp7NKgQg89vgOmYF32VJMvxr/iNRKbTbeWYsrv
j7/ix7eoOA24tkNb6I+vGxDhdi4phY0yfSlG5MnT1IhoS4fYqJSwy4+FQw2PRI18MvErKL8sY7vo
1bB/x7DjgP6syqIxNdYP77Jc+MFo7EFb7dJVFHRkFlBLfVEbWc1n32jxqb+hc6UXRhOeA/zrsCJS
PKsqLts0F7L/5bC4+8Atj+hxj7i7Cgg1jI/waGq+P0t1EdwmPzuwCPDd3sgCZ24zVQs9okovKTzU
ntJ8UTr9xLSeBPFqcIR6Fk65Xs4n8ss3wndf33To3NA2u+I9V5YZitw/2Ur05WBnd1XBtH9XUGcQ
Hz3t+QETxdcbVwdIMtzqWE4V+AdxlGmXcaGeko6xyhan0THxOJScQYYbN/grzaymTMaO1OAo88kl
j6W/8j5xYxa/0/p9uOyRx2dNFv5Ok5HrDHH/l4mUnnRLV1hFXfo+lxOsjTAKSGmWb+Rgyg7D5SAp
ATKWJ/G77svffBaSL3OT0OWeInR2IfOD2vH9HISWKyu/z82fnvWK8Kp8MDONe0AVxUfFwYK+6p/P
TPclxrVlof49AP6HF0uLc0L4/PQSBQNAioF444DN1I25zwmfMQizWn/pyoNvIRT9AKHakHwsqopR
cc8TGUASW9ZzM5DbGMcMBXhQ5TBl0BNpYRhtr9wsTofMiXymQn2zmqThWY/89t/aGS1eWB7m6opH
obqpDFxPEARPFMiESuuS41hPldpM92gFR3zjiwN+Zng4K/Dm39VfNWIbIUob1U4jz9rCL6CcSwsq
BlVeUGKWqf3jJ3YnO0WaYfDyN1gr8UP/nLqSNwlOvdltMQOvotGtDQK85xNHtAWsMuyiePcC+U/B
UeufWrCg0DxeK4BjncRjF2IvIWI2xv4lqONL99C26C/QmgWj5KJzfqGl6iJ+ZioX6IIkTT5ZvdwD
XgqdXHzdoMRJ9eoCuNUe0x8Xn01JDLDdAV4AVB1E9qYfzI6G+STIlsyv2pmK+2kFgpw/mwhBrrNE
afP6PPzIjEP43AE3eEEbzGzv2+7ODuTiVK5eptvhktlknmgr1Z9lY6WC+AGblNWY2Z7L6R65obHW
GyZ5V/rrtaHQZ6DIRd7bDaYhn3GDnaqkMAOj71rVD1EeLLl6i+CX4xUkqU/FmCQtb5P+5N8ZSBEE
rlcKb5VSvVwCGQVp0YeY3yiB+k5zplVWZPSDehgdawwgeUvnwvKGXJumdu+GWN+rZGucnammXltH
WAn3VsIOGbuYDyDynKiefoMeSbwQSyYvAfKUZ+OFdCJb1751O/u2mK3uPwF6M9UxqLAlAbCvOBBy
4KA+pthaQ2IprX8TrBhF5A36gW11p5tkGR5MTn08xDyabfgWC+SJmywP56DlFBcExnc1rNI5kCac
p1U3QkdklT01qb2nQM6Sx6cI44topjKetHvravDlWCn04Z11uV0nRrfCTnknn8ofaVBb8JetdZTV
i0UfEgjf3biVYWUzNh6ySp+Yl4UaXV/bVsX+CEw2JWhHt3u7sKoUCzxPTPe/nVFd56jN8Cae/bGY
nXnenvyirQloY9qEOA3f2++/Dyk8LSsXT72cDm99cbidxegUCh7hshZGvurk0mTKO19WC3gEZc2l
5X6F0vNgEo5okG2ol/K6vn+UHkaYf5UuNeC5vxjr2eZ+7glXDxYIiVXWwWf5h07yGiLf+6v4wCSG
6INHW/AvFZP/5V45xpXQvn3PG79RoaS6tUX2DtH3BbrcJgpWGlqzAlqqwr2aU3LyCYkalGyDspTD
5/7m0bCRfGdcHMEFGUACk/QlDofqflTWrd0wOvIV31GXIFOJEfyIeh0NePljfyWuhnMoBrkFeLef
yawPxMt7MODgjN2XLvMaCGZsPYU0cNr6FsVzfNpPap4NzxuaTENDMnb8f4OQuL7n4QSBeL452D+5
Ijcygehjwg9Y3O8f9Ru/McYanKlZ7V+DLP5iV/oN2jC6JnAc3O9C+zr0Cc8fmRA//SFSEIaxAihI
5Vc0GfU4c6jsYXWKHi+FSFlSHG2oa3rx5dTCrqJiQbRbRAPvCSFy7e4npA1nzI8nF/BWCMsfy2We
xghMBHII7zaaSAK258rj26tYpb2RC3EON7ZNrjRRdSYr7AKr9yyuSoDobwUHqpHDrLmpVBzgCQp+
hnLeJOvJs+zrujXc9TnrnTxTRWi2eUuDsAULplQQSJ01GJwo+l/wquKyCVoxAHx8/24MHAhL1pez
oK76C5vqswz6eihLVswGfPrJupHnWkCLlnEPsmVbSF5yZMvRCn3ucBWwvmOyRWfjwmSbiy3+4wdu
MtIuo+YAjYDzoXByEs/fKoNxPIW5R+aoRQblI8jP7gI4VUoUI8R/bfrA53jvwBI+Vb/XnRNLdiTl
mL6OcxAzGmLju0OR3I6GBomhCeI/i1PXIZnlb81mQmOkIOqudnjBufEnJrRVnPAf7N52XIVvWcXO
7tcdKRQ/gSDMS+QW6VJ+nj++bV38Y0gbLJ5q9bEdmFkofqpE8ZJnPZNVfcCZqw6rCKT7wgtmZCHJ
crKhPwWsp3ydEM2vtQ7oqaYbDl8GDCMI6OZcKtdBEhuDINdvlrtQR6EbYC6nEEOrs/CJhOOsRitc
j9ikUDwv/0wVJCTPi93NuX6gD20XbdPUfYyPn9UyjFjASbGJHsCDJy46UWNSBbnG2NRPccXavR2X
kMuNbDQFjdd/1M3iBXzhNpv/9/ujjwJvRY+BGmV+LbLHN8vpJYmjbVePbwYvi9GhK96ZcwPe3HKz
Q5dZ+ivmdhBtVJR5tYaLIbfYq2i5S6qfM9kYsBd7EPCX/4T42dEEqo5uLXA3QmDv4slWEi5YevHG
ph8ytCuvHYBQcwdyUckRye+eJafcy5hM5ZxIkUdz2v0X6DzombOS8EkCeeV/2idpRRPEyfO081XT
HIm2MDMRDIr5BzVykfc1CcIV3g5/UpKkdpl/qe/HUZR4pC57UDbe/bK7WT7HVr+19td3nbkBbZGw
6oA+hVOaK5ooxyQSTs9ip0noI3IC86XOlN40YS6+SM+WU0IWz2NuRZ9nu+MIR4CupVD1ta+5xlSm
Tx0CC/vu7SqvbnFHEl098YTcWUMhwD2VQUgG+pv/8sQjlP6ZBB3BFgJPXVzXa4XGKcIfOVyWVMG0
QjTXvRNzZ6cgycSOdO3XPp+Y9JaQb6vuT8Y7cBQMnKMvup70KWUBql8N4bfx1KbG3w5+A7AdipKG
9zrqpi0JVH8BM2Lws6YYGYbdmb+3bNPHtJGgo7kyaHT8fU0x/cuRw+9cFex0y15HqBDrXlGVwBJm
xSUT0L6Fmm6N+hkKzU4ZLF7k6cUoLzfpbCHZgsPiFyq0MwN0Ozsddg6qjazbiDMNT98nGV0xUUPa
niutv9m2Sj7EmUOJ25uUDbKnVPig/R5sgnABQRt0cExZchYuamq/f4P2z8Qp6j4RURnLyqpCMhJL
lXMKmeSJs4TlGzcOcXD8HRWbv9agyxHeN8Z8DUG23zkAJg9Cy7m1zJTLyE+mED/yK8RVTn3hxfaM
R/JORCLacG6x5tE8cKsCeP1GjEtYpUNziTkr70czzIdJs4/mS9BuPf0bY/9IWxiRanFnQMglVCFu
SdVQLclZMkA5Wjx04qWguczdqPkOXyZeUWUcFfgt/eBhzHewII8HE2hO1Dpl94IIWclxtYHhUMy4
moJNPNRfMix7xqmiYmxoAouSAzl9pRpN4lGf050xGOCpy7FLisyUryVAnp5mdiz5DVHE3RJrIVGE
7AtYjHq/l8yvdliUE0Wd9e3ft/62q0uQr6yusRT6/SSFQyRPWtKjTMJ9fAYvjXKQlWAZMjaMst5o
HEt7iaKdvZtYBknm9apztWUvo6562yeGNZdgs/ZRwFPTsGjpssVFo/mrcBMaEwWv74lKqYlzmV0K
BSCpFZFKr8TT0i4jSyJEhPphmNnjdzzcsGYNENy8kKCKcg/QSbswlbN5nDXjbvWYZ7y8Pc3YhdgU
UCvJ2XvzIyov3caXgfGlL1yC4vitE43JxvNtytytaQ9fCJwR1Jg6OQocTY/fsJ0yWHwJd3eRsDEN
azgTWPDKrPAM+pnkgQAt+DuKWXQFloAalRx9Rkis4iwaP3FDroh+0chNiOcLetynDP3d+0Rg2j7G
WsuiAhgdtywFpmPSnmjlcbdaYoHDS+Gyk7Qh8IfSEhDydWOxNnx2bazcdLIpfRu789TTaOoiDiYi
mdicVRlQeoncfo5wVChN7iFLTBEMC5vPYclP3PgeA1kO9fZtzx2FOWn/rMwXvBQwfAxfSqLRwmGC
Q3M5KlDdBCpHv5S/exY4W0iBT8DNJVU/VuLl4vTtN+oI7qZWzPUi68kSWblRJB8bYjn+BQMdttHv
e4+zEZY7xj7aekBu6X6eDhaSO8EPSXxZLZ7Valo/Ud07VF4p3D2UwWZ8ebGgyjPyv07lDH54JUjy
XzEDQCoMfunWJ1WMyHIl/88WbE7U+vh49M/KhmctQSdRbxHEJ7tpS0t+TTNwjSoU8ia68+OOpwvc
y6wqnCewDzyhrQjD3XOjFVyr4QUNgEl8FojT+f7Yb6iA8mVQ4m9hskpyuMf6uKhjKZcVPmicigAF
PuQahvty9ADauTu0+bN9HJAekELD3subbDvlqxPkIZzcHi1k9Wd7m860rh7u/N4yznLGTc8JvwDu
npcHXaoItuGhDNoInWq7YRnL7t9ahk6W/kBgk9fG8dBclUGR+xJukH3LI/CVSUSaMeyBXPJTlUch
hd30DksUOn2/Z5sF2UzvqkbCI9bZkMx8RNRjnE+g2+NiJaXUdFEDmEsv31Ov9iseWPLinE6sglzz
vO+iAZ7XO1AE24ZnnyTtTV6wKRC3zHum6wDgsU6UaS9wHSI/Ehdks6ywFosH+0tJTosEHt6kJ6jU
ID2OV3jiYs9rt8whShISN+2lOCmtVt+i0WHYIRJsQBua+1Y005UGmG/k5BF4LsUg51E3TJGPPL0U
3eTdhCxFqmE08PiFNBVj9G9yJvz9MJfKOz1h7Jfwpg24Ke2Z8cwDrQD8ntZb6rmNI/yQnCebzvbo
D1mMNgMlyxi6SQ32pM9lt9MOOKyEtLP1Nxdbd21bZWMtvVi4N0caVJOog8yX3l6D7dhNfkdyq4/M
vigJtOTEnHHSofsyM1tgu0nUn/pZ0CZpHp77dXj8ZPfSo0V4Wfw0oSInRDpeGu4BcN46RR3bIsHR
LiO2HB+8l02XuynEvL0xOfXJmLaVoqQxxJPM6eZLfisFVck2Qis+oJ9LPb/B98Nv7HS2jahXRu9N
Ix+AMTre0tcCy1P+f0BVC7+431R4ENemdR7KUUZB/0pMD6gKlrKGAgnOgjqT5rkjw2tWVZ3uXahQ
56CfdYnWNq9kUY9Kpn0/31eat+XPKi8KoMmBm/jA0mGpvCxMQlQ12BgV9qDCw0tgYllkdVFWOSZy
W9yY/fA2IxAi4B+rx0PmGbVbYHHiRgSgxB/f14l4A/0TrWQ3bA2BqCU0nmMEHPXvSFFa9o4xvzC9
ZLJlgLOfTwBOMmU8PncGIRPz/oiZueSojtWtKpNnqQ71ITMdcLmwIR4pwSU1NaGoFxnsh6zUkXcJ
RzuRkPhPcvHf3haTpAoZyZWHWPRWCXFnGN/cNb2UesGlK6hcicmyfGWLiHO3HpXLTQOLAOoH4m8u
+06CjecGkVzQIMzVVbq/1dbNdDK1K7Olk4n5+T4DvWxhEgsGMjRQxbkpvv0zwX99f4UTb/5fO3lQ
evlnhEn8o3mXUqR0igU5L4ePuibsgBjHpzxUqshLXW65dZbl1TCBVPosDEUEkmNAT79D6B5kI5G6
20qCR97jvDLj9NxoSTQXtgrx4GzYOui8FkYlN2ZvOBP3g+lxHBtecqdruScJuvJqyMKGV9gL35Tu
AzCR1oNkE60Os3dHcoZNItB/42nWGZzgzNaz3+IXYdart7fLn1JaK3GaLONOPJDPXLC1ohN3APGe
x6PYbxsMUrRC6NMn/D1QLjR3pBl+C3gXn4KTHoSldwjV/fPBorgZIapabzaAzdrjMOXOkB1WQUgN
yVmzQkz2ZgTPEoq6cZp9hIPSblj6XX+W2yjZLY8VjqgASqVKcYi7651BqXDx5LgQtJhrbvPRQ9dw
CnB8kaGQaufM/ckjNL+Q9xOqyXIE/Vf3e0kkthZDCU8CbnS0kDArMFl2q3KXyWNmX3NdZf5UBER+
EJIqCdE/Xx178okTsMgTIB9NIVikz+T4rA7xNgyWv+f/PrRpeXoo/8J9tFHcG+7fp3evwqGo0O6s
CJasrBqoXpb/tSGLNGgFwg/MY/mZuBJ3zMqxcqOyAMaREeLfza6vVEzFlrpru0bsDjmnaLbeR6+O
b8x9hwOVydg203NBiZrxgiP2/EGa2zyasdRjCnanXDjwaDkkK9BhJvihHPCAWNkxO9cisvmOMRJn
Kd/bX6TBLVEbIM4Rh4xD4qbjs0EvzGS71vzrYhoCp7ESgLBv0FENx0M0hWc2dPv1XCGkZrdPIE8I
70Uxa3pB0nsxlbbRL10jKugQYuaMCuzHkKxzXMNgKTxG8GapSCTAPghxB67PIfYHYthz+m1oRyKc
r5PKkdhvOK/aXu5tgkfJGAYDvKvgIGcgeMnISKwPhLqTLcQfZTs2um6CuZ8pIf+n+VDqI/wLecb/
qaH3oKdFfgkLduLtiyk35IPZop92hDiAWXFlx9G+WkxZ+K9w0/T7y+Yc/6MEHOhfiVY8nPA1N8OQ
yaBDn0dTO2mFpweF/2CL7Er+HLpYRoZyJmOLqQ6dZ8gGnmUiImEpkjkePYHD7k5/6WOItlcIIwiR
rJH52xqDLhybtpv0+jJCIALquyDb7xKyOjL9hD3a9OavAO0jC1c+0v9nC1/PfHBKeTKuXLMlWfnM
8igIrv2qISVZJBi+kLL7ncLsSH+Qd3HTcwvZtMf2xiOjKt4qLHq8lfoYHypsdc5nH4/w110ymB82
keG4FK10xEaxwLoTJwrNpXP7EIl6obqaYQLuUXwfS3Knpt15z9HX5OfDUZI4KONkj7tEQvKS76XU
y9PmOGqoTEGmAMRfJSjlPpiZ5lpDiGQc2quAl8LbABEdDcZpOCbF/a9dDZ7nVsGNdmo5tPm24+av
ce8wW0arUjDByoeOj3Ljzgz6geLQernwxGsXIcqqoIn2IzHGpySjiWT3SXx4C0VCvEZJebjbcus6
yourQHviM1MJOOA8Ch+ImAxZICWe2d/0SH8r2FVH3GIlYLeuSpOwRBESabOYIjUD6UconpenD21w
0KaUO2R30QpWYBj+QkW/KjxmQy0wyfDEK2uKjHLaAciBcPcNanBoJrjKMsnlU8BekCRX81WuGbt1
fkWK2QiMgz1N8aQUUvBjvBKz47JMSgEWW4kz/TJgKCVdzJLEF/ZyuoOcHioUOPN06DX6SXBGU+JW
t1ZxzZT/emHri1fiERGd5sOkq82idOz8PfXHMtLJ7Uv1Wuyx4c37m1630aaYgTqfqonNWuUz+xDP
5FbQVyNijL26Xu3sXxTtJqvGVEqRzTsT7Sdk/6zM0AWQmCzNx4V6I79GdqZglYauAL+gm6VhyOhb
6W27MV6Qj3l8Q7KInNUVwhOSE7SmEr7wDlLv5z4UbgsmCEQd/i2ZHCpnKKn9JqvCaBZscfyacaMQ
Hvp133q8T+rrFrKGXKaudKJ4vKVLIk1VweTiPHvu7rwgLA3/xBVrn0Ox0G7sF7AxJ+M6AVhDPvL8
d45XBi13xy0vaV+sl6nI1aEIFinxc4WEXPOe3Fcy/tBehfZdXEUkjD0X46ibChYjJVjH8SxJ6jZ0
euDiwA6LNIBOfOhYsdJPRaM2MBdpb6GT/Hz1ZnUsEr26tQK7ySkZRwufCbPphJtkbU4MH+bMP9GQ
SRr4Ml6kz5vzP6aY+/w0UHTNo7gq4m29Lhb0ViMtWXQ8lLoWK5kMPHzVzUAGRtRSPiF5hn2LR0S/
RBXS1ZsWG8ZIlf/mq+WbTa9njZVAwdDQJtJ5bK5TPmxhNPGKsYEnqK7B3NiU6nZzd1Dm20r0k6sT
reWx+VCJSOjrdbJmCIxJZhonxFG4IV6sRye2daf+jEvC0mbMJWp8v5V2b2BdLE2++ZC32UG99/Zq
gnRuGO3dsFSQBTtDVHsgQ4peJxJAlOsBeIEsQmgdhnQwCroPtOc4wb6crckEBUFCCDikUtZ1vdz8
BYI3Pp8wcca5Jo2SpRje3LSwg6Ehe/IEILWR9ZH08l3M4UeVh76o4Dfep2akP4EAaPTnfj7rgJ1j
/ZqOwNxpA5bxr6JA/zypUaUkm2goiFxSjI6BWL+Fg1hqP5LikomdsDOSUF1vrz12rovEy/dB9NzD
4PcbKOkdjgv493QfUZQFyN9eNUPNfOhZ6QDiMGUleDeoT+iXYmE/OIO+ZfQRsAFH5oVExt7CVtfd
/A95315uPDiSDq8txJK4LwM8398r/+RV3C5H1G3m4GVi6qVlmuxOnP2dGCHdnzYL+bUTA1KFT9zk
/VjxomPab1TakoGNbaqcze0QUw+TJKHcY34zrsPXZ8huULq8tE2KbXDxXcr6/R3eMG7wKCHkerBH
ltcl8lcSWQz10o81ivOQ+oaROADQnsK/KaMiB8stW6A9UNQLLlmZPTlCRekLO+OgH78QGzruEMrM
+OGGuNKkvPcCLNILbRNOG5Z0maY/4FPn5jxS1UQrNbPPvpr248g4AI1Z+QCw2KhQ3M+H+mpFoH7k
+JD+6kTAoX7WdRm9DNH6mvjoHua8dkapKplNa5eAGhwVj//Uywbte3fJzlVMGCshm7p57CdosqGc
rgSf2klQa/bFdzOnxL8yHHokILeoLDN9rPNEdEn4FO3PDy5UinfDyzow9FNkRFfDBhrTCFKUDNiU
dYAFLIL5D9vGO1awt2OEGrFbjqQO986CPK/CPzlnYElM5RcsWNKd0jRS3ZvzTSG/H7UDnLewG8Or
GsTNilvlrsxaKidzZRLuqr3mIOixoCTqy1P4vlQGnUCEurR9nb3tNvvgqt2ylEZjnxGnyjiXoKBf
Zjpe5tpN+DuvZWROJq7GQTQ9syw4RqkpYgecJpBL79Ao2IKjNYrBSwyhjy9Reih07yS3v7D7k83h
E0dtZsV6mjX+0oAc9YZFuzZB0/sT5Quktc/1mf3Na+2pbDr+bHULS8L4HEF8s6XIuwB8FA/+yhKJ
VC+BHvEUwis/jBmzY71wqCgo/mwUBjoQpzlpGf56HIVC+RBme9jwNlmXXNImGT5vPi5Gm0UUaW54
gOh21S0583f/tB3PN1q+AD7Luo0BiwPM9+RenGUipXw9vr/h3mYjJQt7Od4Xl+wtdL4mvCldEuse
MzuAqgOWZWiIroKimYrhwxN/nJPRmpcxUo1E7oBO8JjjNWsHR4Sdfxdg/OUJm3jk/JhfWhYEVxkG
gYF9ZiKjv6LrsAYxZ/PfjXA8VrS+AnLWuRGw8yl6UAeuAL8MU7+NCDE2Arux/OUvcDc9qbMcHJdS
7xkwWGj3YwofmNjIWi/0l9tqAIjiNT7K0L214E2Zp+hflRdfUv1INQ1M75XpO7z3o1R+ykCLmAn2
i81cmtk73l2VovQRBOXfL+BVxQRVD9SoE0/tTQy819LtLX16pMnOdgDOnjJvnTGxc0zdAkQ4067B
9y/RR4eqfD3fTj0orJdXQzK5oE6vS1KQ6yE6YgHd5rQ9wVbcnXgLHYeUgqXVTOdv8TP81pf//56/
IQvHdZUzQNLiAT8lCxmEhpUJ/dgQTLsmo72vAXqjBkMD5bD1hHj07akjNfQLOvHC+hDKWX1Kp35+
GfzAidiJBEtKXx1+t7OqK9qgJPrsmC2wb/Z/ygm+D88qq3aCgU3qliEL3X5x7U2T6jWk2vQRwxnn
FJkTPcg87Jb6edIj6XgRYuqOBo89q73Za71J0fubx8nkdypORgZkaZLuqBSZcQx6aEyeD5u7OmLH
AFVMlTe2wSTkGuPGib5Pg+QYmCstR9fOn9ER/gNF+oKSZ7HWcXvHYYMZ69HtWxjcgohvrW1xykBJ
5q24Yyw8i9sRVl2sdA0vEJ5a2dYneyiHLSWvLN7qLt8zpWXKVz0BOmG3zQrfDZt0h3sdRzZfTJ1X
R999cET3DSczHfujqVAW2hp5CsNbJCh7VDPzsys35UN9OYfQxM07KIgL/jSpt49QsFVXHEio+XpH
+gooWOlIYkU7+lla7keaq9m8TkJd1itixO7QBjWbDOv4dAB0GIAapphhUfgE19Fcvs5M2jcEPQdS
W6Vosp3q+XCulnDDtkmzAYL3r7ZrR7fd8T/eeOCbRy1NpAIhp2EmEHBln8W1rT3SnOh1vnWpBIVy
sFkRLAjAAFq68n8+VHvaINmY5HW2yHXObardrqXYhwh3I7rY1KUXVFTqFMIa537Avn05nRr5ZZAe
RFICfjOuhN3u7D1801i16AgswkoIwxwIHAaN2Xx5m44irZNMjPsmEp0KFcgY1cHHf0nMH7/6UK+P
vBmnND3Ps010A1JZ4cA+uj4TVIO297meZJDl/KBdaeqdeO79iSyqX0rRcrdCxxX6FnnL23lHojO1
DwjcG1h06jgRAqv1ztMDmFIq6E21gIqgC69N+Eu3nENtMFVk59G1tX2LSIVfrH/MD/7MJdqxkxMf
jyztaQEy+cE8YwbjwnsqSgEiVReObuufEsMw7Jcrtt0K+LR0XAcJ/cwYl20Uu9jy0tAW2KLN2l33
EPHSNZSxJyPJOgf6Qgreyt/quHEysX1Q4WMKw7BlEE4kZvYZMlPaSrycnQAqWYy6Dqww44anhbor
pPtxc9OH/keDVd3khrtZrtk9pc1GicncmV068R1Bx6uD1qYCGnsO3Xt7ybJW6K8r18BWgiczfYTj
Btn8UezIZvUtbMR0/pYlkFc9dBK2ZhmrjtE1LZxmD36/FcC3l3UkLWj9yegko3051VTc/ezYLqi0
y5bJ+Q4cQzDHlPQ+u34J7TlCbZHjZKrw6NCHwMCq6gjWNQtoctqTQnJmcBwtr0TjZeBwneSk5Ox0
VYezom3gJL0FX+kn+x3EFJN1Ei1fNKQ6opXgBwQrJwkGLh/GFlV5XnoS3vpRMl8bq/7Yas0vy9Sh
G6n6tPWR51RgaQxmYRPPq1RC3d52l3oPwHgrIGbExAdHGHrZkLo8XuUpGnVH1DpAy+XGH2SrOoVE
5VZIIOle89RurdD/YCMEIRg0D5jw98ccJ7FzAYkxcQEWTiZOuguZca386deDyGlLZkiA7GOGM6K/
tWpRhyc1QUr4Ij3PaYlWhrjnhpTojM7xG/3SGmXNviI1vTinmTGTV+G7IcggtnzqMOgn4WYsI+Ux
uXcc6ild4DGUOGPXw76ZSwS71R6+NfVWQr3wP7ZF8jOyVG91qVyaL0Fyp6nvIxoIH6jX/TBYZwXC
pluwRWmrbxygIWtBoA6/tb3CkQvRnqEBMhEOJmvPcU6mSqvxGYz6n93LPiQ+h8YltQ4df+XhED0B
wLQXSS86i/ax6XFJ26P/ycyfiXbcGTCZyXHVVZ2Ab/5+RgB+WBRp5iPzP3v0pVg8yve8PC8R8Wk0
vNgXJAUr4atwPi5GNRXkYY5i5YgKsQFpItC90ZKStrFYLFIqu17+l8JwFPGLjzseQBRsjiTYMpgd
NHF+Wgd7SADnEPLX5OuZvhlGqVbKy/UoQVac7gPNd07vsbv/f3EdHPHjhsXqoPN+TpyRm9m1FVie
T5jswHYphMps/EdQ/KN6PzXF+CFlewbvSGkzniC8X6YCW4zpcOSwNzMCfwVLws7eNO7nlUV/S0bR
4bCbFLuUO94vkbkOU9MPkoXbBR5p0W7bvvfuTGU3yjJVtwoM51ldjHXUoAf1qR8lCO7HZWeaSb24
+cyOtEAYryVLmn8wvRuvg7j2yJ4rkVH3iIR0F9CfshB43EPZnwa4HSsOYhh7BY3HRsA6GVQgMiEd
Hd4BH9HPc3yNEKsPaD56hPcrg5PxLPrIt7s5UMNPGOEMc82buQXhIK4f7sssNtfLJ4Hr1funPeMS
F1WOSA4ZtulXM0WgTz4XPVbIy5st3jz0Oa1Nx7XITztCm2FGdz5yD1pa8jETv0IIy0l3WbugV+5K
HPpVCxL1xXnrVITdJYZ7EAqev1prHEpULR03Bk+IIwWM6m8Ba5wKkG9Z3hrVnuqMxCXRVi4zp7TP
JwCM/Rtz+9RwWF80DyRhyw61R3azDK7EhUKRRcn9NsvacbG+2vI4Mphs+0WLAJmMZf7crGOm72Wt
gjh8EZz5VTvK+5I2V3YAOFWsQ9x9uAW+SJwmrE/fTD08iaDlp1KfNFOdoRr+VJvkiKd6e2Ye3dRn
xiHpYP5BEj3XYbNboJLyzcP+86MIz2BoRQuu/PPWgeO17lppmF/MbrtyJzwOffzkXNHPmv/juqgm
8nLX8f6DbQIRuS7GRNQaJgifu0qoI9KxckHiGAk3Ed3wyPTFcdFFF04PHcq9xRuRE1gMhS0n3G4U
qnEHmAVb6QcphQ/tAhoRRXI0tgR3uHT3w1ayXf8Q2owB78WpOTlpud+IBYgBZVeea30Ty6d9rOum
2fQ6L+4tbcdODv3lXJDNLKNof/OUyaCz/yLAsKcuXQhBhFPNKSStXZReaWJgQeoWIxWasmq+DJUC
isjnAHhPLipKmqiXOct2LZWvhjwomrgiBBsbxqSJ2Hn3jsPedmC1YxXLVgsdXmZuJfZSdKjzYxpj
mf6g1D5bk7afupFCc36VbNPQ6m093HRZqkHcOCh4/4XbVeIq4ZBQnHWbla/7jcF/INAkCrI/GqBh
A/Jo/SSWA7mml64OWI6Q/QZJZLysVFXcu62zeXBZtsfNdLVNA+OslRWbnVLeuBt55H1SLMb8tnUh
PTrm+9aBz4YvZu2TeASYiMBFMuoIxd6AuDq7hRzPKOckSYztqVBYtr6zuyD5Iex5H3D3YFUFzXxl
9LTQJmdskxg4n9U43XvZ7jwDOZD1eDeECZHH+sXijyc/Zvfdd8weO5UB/F5lgCQUDPuTbHVF87N1
3S6SNZcqU/bZofTpfN726PK8KT0TrelRccFnydNyM/IgLCq6ugWY11+13oz5fCqRKFeyipCELL8l
5cg/Lb9USsMMSV2AwzmF98tesUrG3D+ifI48DQispR4lkbDXzeyTOwtDxBT4sJXvvKxhNsdE30Yg
uN4PEB7QQHKteywuldgA1Pn2n9GUcyS0pG1iJDNG3a4xSwoyWgPhm0ZjoG7TcDA7mZ6SCUhSGk6B
od4pzGuTytBxKtbe0nav7I3KGd/3xyaPp1vH4qRit+BEqkS4ReZYkvsaiFhz8da/4kiQKDV6Kxw6
MwXCSAuDpvujdkmY+d2VpzIXwxERY9N56d34C0Lk6MEsDDSOrA3RXw8K9o9CJOMsKkkwkbxIRgQA
isiFdHxtIgIzjOvvk/D+lrH0mIobZ2qpSAbvS88fVx3G5qc9tnNoeLENQ7ofBlwBMr9+z5vDkzQS
tHOGwpnsxZC7ztpTn6gyZ9zcSWABezRlM+AsB/7XGBtjnphrdKwujTQMpvR3UbgGpNe3iAdKEEx+
Lk/i9lwquPxcC+c8Bq1kB5I/DFKeRaHciY+oX5h22WkrVTXZowBm3E5re0q70ADwbRm64/wKimG9
rD8Q+Ot9F/MZ1q1D/JZ5IKKEefMjSxJvCiptsjdGRZ4h2y+eJHUcbBlVmLb9lqtdXrF/4xYNH9CU
Y2Doo5fG5WfgThg+6TXJR6n5h4vBh26fQScrEKxbfVAGAFGd90EvthgUlMCZF8A0WKVITLENyRSw
AJP2tfJC7AOCbQmJRFPOF5WEJGA5GhYXcuUQf4KxZK6p64+pNRo00rpeXoZ+Ori46VimeW63uNGH
LhFPdy1LpW4kwhh757Pm7J8245dmBnHttxm5iKEXgX8RR9VXZpNUusJeyCvPmvMq9EMP5jnAl1VV
TNPog6sSz13iTWRxy8PWn5yVi9YVerDGJO+j0bftsMtzHstq0H+Knp8fW3SlY2FuIQeCcoIhO4kg
EbHlX3IllHyiuAQzvclHwua+rMr/KhQX/Guv6T7lF3V4itXHBVH+sRBFI4r5ewPrcNaHDQauF7JF
nesy99fTLsYPirGD4iald7VjBzR9fUP7tBtrYxBIEesNS6Z/G7Gjts/+KE8/0ckwJor7AEcBVjfq
5q+KhqXLdAGQfNE1dwZwg53ejpJFwgzof27I4T7Ygn6sU1MjApoxK9lAxJXuGGgcihYdmSr3SfTj
suzQO6iudYUpBP/D5ptvXPaFO8mjp3Br+Zr8xSEFJyA4H4YUJcrM4eT9wsijrsuYUchAd9gQ13a0
sZ5xXACUKJMTihadDLKv/UmfDhqu39Dw9b7NESRjEA6iTANpOSZM6YSwHkbHYupyFhVbSyzH3l4G
6lBe6dRClsvKsxe51Oo2xl80c37XpCVKpXZbn/R+0QLuPWWjFwZuB1brgvxpd+59ZBwGhutO+hIp
0sD3UYbv42pqd6c1d/XzZKy9ZC0SwSK4ira50w8imYrYiVKu6gbazbvT/80tkE0hH+W1oFO5KJ03
ZUu0gjKcY0Ht58bVppyIec++rFV2eGSw2V8co4JWWHmUuTV6nsyBFtov8RfR39GEplvsaRHsGeYJ
ASLSSDbcJFZQ/pzAnLct6njr0c/4OL/3yBlKe9ogspIYziWYnWqO9Q2TZ9Me6B8OM76hLZ6h1+GH
8JsWqT+fBnryig9rbagp5/8HtZ1BneiBFcJRWA6UE8B8uHVZ9UDdSO9wuNJoRID2wtkw4q5gjmyn
E39rKcbGe80VVR6rryVgucWeUYdrPdsmOcWPqgaXxzWdK69ET/CLmbH2w7X6Pq16z8kw77mlsGmv
1vFwq16H8V3aU9UoZ6b8M+zZw1/pQ7DsqDUOrjJ5Y9IlyyaW7HDIL4oueeTTm6KVvzeqBxsSag4Q
N+K+Nnb+r+k0LeEVurEbS35yMcddJUBddBprMvRrwGF8/NwvAxPVwGKIasbUG2sB3G/U3rod+X5w
C3btlzPUrxx28Kk9IvhpRZgReX8swOlegSw59NjIjlyGV7f166zIiPRZ/gBRIBiIBYzJhUzN/Tbh
0V8XVSbhu1HlxUUIy7phdKyW9KUpmuzdGVPDIiJGgwkeYL9b7VQhK0VTyYmzz4oQ3fRmQ2qM1Eso
6Y6yJMW4Ml178fCol2+D0hLOHzQU5fRf10ww5Geacn89CwZCeiXLg0x6p9zNHuZjDJQJPwyoLkhW
TsD6um1S6tWUrMo7RAlhBHpG0th4U/F9W55xg17Bv24/Dafk0P6KRH184nzvMg6Kp8HxSNhLWaiN
MRS9eYjrwis2Iya4hR2YfHhTTvD4QYJqxhmUdzusSJRI4hBhZwzh7CGNI4tQnRM/EIWpt61/RXa2
rmXw8/4yUsxsyfVmvOIv77XEUyYYpjYPpJPhEv/ehWoAvapQAPirgIZDVKcNfFtdt4jqDDh20fMv
WFa3mH3sxHv6vhybupbmcDOe9UcfBjkwUqFAETt4wdueXxP0gcYErp9PBiqudUWW1BDx1y0RJPJT
R2G40PZC+YMi47JmUsLWfI+Ix9V+z8tyOylOk0uNMoxmflAJm5kfBDVuB5x6NC1fKQVBYbScGqHJ
LQ3+Hz5py7wxaqJTps52CHDStQdxpt71jVTQO7Qus11b5VoBR248xxphu8xxLoKpfanhZj16qfYC
XiMZQeezJ4q4GA/+YIGioj8xDzM/2vYLfkY4sHR4Pra/lGAidFq0Cr+suEGRyr70G+LU8+zFpyto
0RGR/ErMmZuAHjECcBaUAOqzFdAdsRbWlnRE+Q011RDhX4BmyDaWjiw4GqE7NAVRl0D3OY1DIqBm
lG6o2Rih+yU0ZygLaCxOiFs5lRPvyDxFTFQ+LH341qWCCavwgK0/R1pkS6UeEKzIg95ybufRoQ6L
5WywiAGfjXXOy5aFdbNiKH+RS/II7CdeO7/akWkkAnIHPk4piH37s8MzJElWqMIHRQs/PRscIOuO
ddFPZ2gPN72YoSioDFYChmQ4nbr6GoXE+Ev7wnxlRS3RLlCESCF0Ecf1WR1jQBMHl9/Wqrm5dvVp
sQvlZ/KfY6KFAgHpxv5d4yjDndTBu93nV2KDVDEbHMZesqDZmxd7zoiJ1Cbaqfirl9oNS6T2eoAp
nvoMhq4itdIH5s2j6ladzGQneEk6Q+ttFXHj5TPSFkuZdBBzedeAjSFYtKPPeLgs4Rys0JckDkLN
uqQPUkt4yAzECwl8CjWoBLH3KiH9zzmfhVn4grMijm/duMsB5OB21hWluCwVe7mb+YHIRQv8CIAR
sM7QAJVB9rYCFSb7u5kioHib+XC/ovMur7hAakkGqSad/6/7QPEpi9IEmx7dRC9hXYRLRw3uxPjd
L0oDdvCCUtf9D+BYBUL+jSWHL4rZBUdOIyWoiTsoOa4nDN6Fvzjk8ZHk793vrsijTpdmr8AQSFq3
1bWe04FZ702lvLKkYjCoyALu6YdkbqQF1+KoxK9byPsNGToh0rq8dN5L6ARwG7zAYPOd0ecTx8/z
WX/2wxqGpw3Jmt0R2JRqONh99ZdKfDxzUgUEbPYrCRze8uEWkJRO7faJBl5FYdMAhI/Zj31jULEp
3DVdIGcYxOu9XgOFIiSCvpzmz2w6OwaGDvLyD+J9OzWcrum/T6aqaUVlDdUla88VfLviIwlfZ4tM
mFKyVI4sX8LmbhfQkiOfxVSRHzPzlfmsEzAKtvWn+/7n34myHwzmcpxood1xkcq0PQWnCT6JkRIt
OaOByze63XQkhaL8VGj7epkDXuTIYyTbpYOOZZhxMRwZY72B7jGguLaW3v+YxJ/8OOagrlJHItFa
PJon1Uq3XwOKkYl020bwVfD+ezZtaeC2L3u/FCRf+R5ekZ8vaiAy+IVuG3zI/ddXMlNZ9yz171jC
/1YopG4MphUZCZnQ89zv9HKBFoplayeTGCXBAylnTOmPBXvVEtUQzmFuONpY+gpQdl2AVbJ95y+/
oHV2eVH9LdtF2LdtKggEPBr19aC5pDM5x/SJ0jqRMw6K6kTLC6E9esWz3aX5tTU9M/R2x5x+krqo
zH8CqYPsi9FMTQuT73ukRabeEdGqmldhXoVcU3VuuAcqBsaZlmalnKwYLWe3HpIOJkUkpRJKV3Or
UwvypjqNxIoU6lrn8dGaIgstiATduYE/kS9zJ1dVB+wFt5NDk0c/pp7lG06ZTQe2FsKSn9doMfRL
VlTLepYXw5fJMXHcGEQIlaHja6UHhQxwGVKcPpjEAcxIuiz+idYFh2ZzJhTSp0Lyy7semtM3SuEI
pQQAbcuvHkGRQogmzzZ166unbO/BRngVaG8aEQs+bCqTTaEKTQFw4GzqbDeqd3/ITr9t2hTN3Ysi
EOJ9cX65CRLiMa5cKasOtY1ASXG0xZFjetWpZCbR7BxjRY9bmZnyBIAylUMLAZc1j6APZtnZ567F
M4Nh/Kbckd8eDmLleeg9NasM613lFMtX8hmlWCXsBTbl/7HOI88SlRFe1Ne0ub23VenZ5lbTq9pn
bzhIfhtf51D6x2n+zBMip8tHmiolqqbTIoUJPJln4dNx7IUgnYDrj4buTOtqDEoc5pP/KeR+UyXX
8dxmZC150CkOoOLXgvjmXKcAVcjafGB5+NOi2ZoIfZJoQLDQEaDNH1cvmcedYXQnXDQQnXLq8jgP
TZxXLlPWr5FZpG0O3KsZfz3OQfx5Yjhd23cbWgjaZoccSsH0WGuthAhD4L9LSf2TiHBmx5E9yXYu
eV/SLppnTHBerU+CHD7zvvqct2ALjoiOBTG0tnSCTfFzHn841XsJmiKVqpdH7KqsQ8BhlMYIuufd
rVtfwvRhkwkMUn0XW52GZ+KDhNV8vSa9+r/i2zG4XaIxfFKeoJjvL48rH3RaqWEJZ29f3TozurwJ
X5AWKQVV0XZ5HHu+9rLx2XVjxdPpxh4Q/eCUQ4SqMAaZ2gSXcHmB/BiaVW7ZUer+5HBNNpq4QeP9
GT6lG1aspLDAMFlkeQYgqpd++rqeoqsnNSdy70H5uaC8S9xN4J56kLYjZ9+36RUsitvR4LD8zsso
M0RCPzkpMc1nZjatpON8R6UHtEWQ1G+Tay+XXb8Rn5jPzR5pjxg8h2zxhjBptoHeDZjZ5uEtkNj6
RVz8/egPnzv0/hlanVd+1JS0ZUM8vxZ3zEGj8KGQahz9qondv7MBHdyGgOiDi7BtwgIuj9fH7GeQ
N4NCRPu30PLhgn4NxgiMO+AVXRCeJntq7QCLpin7PyaLdlEkjU/E3vT4MIZklyBh15LD+dXeGs1r
qnGXp2+gQOBI/w09TmLMtlqxHmo10Hj7kew53eX12ETnIucyhtuMtfvqsYKPgnXld7J5pysc7Fiq
tqHBKFKu9rIG1KfY17R1YVL/Q+O2/2cLKuvQ4h3rMEQav7qMMaW1AZuzptws+LRWbJbIjuGiQsdN
XcEtjc5ffX+3W91K1uCQ2Q55iRTxP2CJV3kcXKYMXEZ2VXgPtUmH1zwC8FbrdZpbpjFlT/KDznwo
aoR/x0iHa1g/3WxJMlKifxUuiDPvMif4qqsItDtfXGhtG8sgL2THkdqhb0zBFgMjArNZSWO9id2Q
H8PJlrzncEJeOYKv0O4tLnRbu3VLH5u2v2V5QDPrswdVyO75mM0vv8At3QWfpi9wyB565L5sBsMZ
sLGBWO6TKfFIYrOVUD8ze5tEyYcXZnqRDubDc+fzjblPrEQ13m5oxuOU9rpinZol1XxM3eJLfZ4i
o/pOWtFSbiTtPHwlfFx45A9oKz0KXgLi+tLXDeH2hRf9MPmECflC5EO7iMxWUMGtHunbjfS0Gx10
qAKDUhnFFl98PEsD8sTBd6y7cQ9iBunxlb5V1V44/kULTVY5koDQRMDXotsn5zSTMbPmgbF+T/bi
36nOOMYtdoUwtpO41RZMc0YmjMsYtQ6EEQGuSCl4nLKzktnO+ZuQj6Sacb67Scrciykl1FaQXBdi
e2ThmWOxMKofbV4YQX/1xEtv+iYM1YAK7Jpvx2s5VbKhRNpzP0QLzrW4sNeQ05TyoJ9UkOupHrU5
+PhXO+//i6MwtAcfIbcsvy6TzSff/xZVC0Iscylv5rt/h7amsYDkzXjOMl6DBPiqeEGt5Y63oAws
C8mvftXufqL9CZv9XiT2eudCk9ogYIgPsLoKquTEVqtpBkLPvq23z5AU2Rk3Tyi9L5TAJOQXH81W
NQidDeD+Dzs0ec0XD2a2VCDQs/d1fp8DLav+lPIhlXD35/q+j+Ml5/wIIz/JVOKxGyclnXXsQbDp
kaDpZPE0rerHA7nI56PoKxP4UqmPrSuse7JOcrnuPgpT6jRfkaaBkfjydjxpJ3GJUojpPuZ2PkKX
Q0OQpErK2qF9IFrb9hDBMHsQtKqnD6Dej6hEUmk4wK53C1kNuwvY4W4QRqFW3zLCZkRFrDS4ROri
fZEawE/8EBxbJhPIpPhsrj7LAxKswFwfCsxJewBozQrvb26HvkabfNyw63kftqoE62y3H0k/VRIt
GVW9Sh7eHsH8D/ehIsJSYoMXTlzowIXUjtkQxipdDN795T9P1CSEculji9YSmQbxIlGxsFbTVuZ5
nXfTPwtmSecZTKfFrWlqngqcUxf0rczlLrmrQGBDKkOjN+c+0N1f2Ell4V48iX6ow9M8oHIu6Cpv
zKM3wzzk2mnBw3LtM3ifb9bOftqwcTeauDnO647px3CuD4JdRu3i9JJRyYG+n6M0jvOmVuQYO9ea
I/vVpC6ZuHLwwQ8cNjdLUUY3lORXXnZ2zKBFLlYyPwy/ZSjNfUjwK9skdhua3lb3TivK9Ia4/xgY
P0IQLZdpG+oTupbUTYl4eP9+/bY/DtSHs+2HmLnM/j3uc2G35er9TZSxOxpNac6eouwDt56NIoS+
7KipDOVNHha2jOuJTY0Pib6/jX1lbs9N5NrVo8ggfepdi7jIw/FsO/RYE8YkWABwC6NvqBfnM2yM
aoQB+Pjmr3e5CBw/x3n4dQz2PrEhFVn3+TAuESnqsiMIXkOLlsuTrbvSoa9LeJgC6j/E2fL46caf
Rrropxbnmn4XhYTQ9Y7jOmWgMwPuVrbnD0BMGOFS3wUWfOH+YI8BKDC35JhIwubDdxREPjVVpAXz
kK8/x/XMxc8TGfiVabEavreB6phG7fDPXCNcQYwat29jHSDj/VS9tbx+CyU0MlzlZWZlTNkAyPhh
OyYb+pOXr3Kwo5l19Mc4KEKWzlpsMLR/FiorqgqWn5dPHUF7f8CIp/7OgcwVU9HBXPjMDYJ+9K7h
WFFErU4movD6yZ0wEzSV1hvcWV8VTRuImGJr6USGlnSDR55yE+yJ8PbIPFXXgzWHKYULw9Hg/n5w
oycjJotDlHTVD59aF9QqJv8prGkMX12A5NQNuRBJyTM2lBTUwBwkQMyYeOvlRRirLLbHOO9BR7ar
cKJO4OxI/1g8Tf69BrKRY0FilRQlbJFot3Z+SsLmXUf4wUIk1FxEJ7ZPbRJudQDBS0oia7/12frL
VxAFbff4oF0/YyZ78J/gg81mTqKwYQ/O7VFxL4hL7yFBi0J8YEuTWCGwe+dN5lV7wF6NA5SQHu4L
/s5OUw10yfoowXUkqMpyh4ijIKi8r1jPlDuLUHeDB2/QaKD/CQ7UBLfXVC5Hc8p07lPBbPMGOe2u
5Q4u1BNxQLE1GPcTjFZSD8KOfYBboDsaY23aXzfbU5wY8QRldb0miHZYUbVR+udyAu6wlbLMrRUm
6lC8q0TPDbBV1uhNFEd0grXBaSm71GupM/jrkQ2SvDuYG4HKpF3vazFjeh4ljY5vxq1EnGRFgH0H
EEAmaOpy5F6sNWdKA5UUnRzztBAIbpD3oTVmd2Sx0GfuReEWiD/hghGl4ivZWMZfj81Y7C/kX1gI
sX3WDYptB8xWcw99qw2pi0P5SH+nRwdJbj3sM/IhqMUGIjbgsG/RGxthI3PdNeIiFya9P4xymGtt
0LHxRN+znAqubpClfO4sj3IhmhIT+HsI7Gh7g6T1QHK0uigFXzdcCusljg7iLKiA688PNGAKn9Gh
Sp9yXeL25mBHNCzuGbOg1xrzxkz3IoiV1LgPolombaB/WXUT6sLTn4uVD3s0lucGWo2X3NTLRYDS
u8hS142v3Wu9niYWW8mAqBIktQGRuG9KrMnnZn8GOwEqogBr9eF7/8UEHCUc8COV770sNdNK2Y3Y
dUYg4l2Bvf4f+NxI682BIxQadY+y8wVUoBScZ0pN1KM9FIVClem+zjy9FaSeMoOKKQ/+yu7sV6W6
R0anKxniiWsG0/V22BYEEr1xOnMJBew0ebYqjF+fxDtPcdwJuEhX+jz6GfKcDvaNyeTzQrit4RwX
ZqUkufdLwK2joWYt69zWwaXOJXkDE0cLJiVMmC+1NUt57ij2tyGUvyo4aTWq7kM0AWSmRL94BH5B
I9VPmdx0yuSQo3BvKzl9DFVn7WXLeJyS+GhVxAbOPy9+z+CfxvzPAkIIy0+NimLuC/a7YaE3peWK
OqAeWqOvxe6jaCcfTVKnqbyCu5s+VyLeBVwm5Xfh8ZnepFiUvWblj2GZBJZm5GaScVo9bg58PTE7
iWXCP/w8MrKWJNmfUjPx3A8wo+hT4f4HWXx03VJae4ErljBfc+aYu+EsvinM+UWhik+0l7mKwi62
xdhx/nX7jWgsCi4U3n2Cuib2gxrOFIZ+/LwpAk5qH6K6JG60REPmIDrBlnB6AqBk/ZpjUsuI1ECo
wLtutuz3SPky3zGGYHdv74SXtb6BVONWLqu1cXgxYj3traBPpQBYpIYRlXa0GhrOjaQgaAswFQAU
xgtM/V1I9lwmWC1Vux6Y+LhO3DhbapImNVVTtQkHWvLccPKcvOXSJtlOOmTsnTLDIcM4qMg7oy3M
fm3V9sxfJPklDriX34Htxjfuu7sG7QCnhu6WY6ZLIbHJCX+/nkQSqMrWoc9lOp5DUrpRpouJ0WrJ
vZAX8iwJyO5Dbd9bB9ME0RS8HEg+2jM9T/6Sy1wvmqF56fY8tE/WJ8VnhZM52SPFwLycKuFdvnMK
kTDijeFZxPPlItFVMlH1RAqn8hrfDvV/oj/bKn3lfzVt3z3f/iPOdAa5b5hCMc68wXq0vyzjL8oY
vU5yp69JH5lmWa3FUFZ2Q928H/IUXV+RNK+07D80VdfZ/X+iaNS9jCB6l7eWLC3yZvLuhU5126hT
4xJ3b3Ly7qqDfo2zosiNMaI5JLy35Xdt9c7jJfmBcb1JsBi98SCa4lKpnFhi/jrv+DPoPH3FHkr2
asADPYYDmTVw3lHB7FXtyXB68GTFBrdWY1oQQxT6cIAdKUD5o8uaU/BfBHMS/OpszJrMnHkOq2x4
8IAyIQAMbmmfteXV+1VuKgUENR1Re73nT/oSteMySGUqs84iSblCz6MZbRobytfV/FFh6S23RBO7
nU+9tQHjfCDHBqqWR3BkUPH4Uc8mWxDxi7IafkjaRsDWA8UT9oG4/tcx17hKQZ5HLEksggurRYlb
+LsREtJykuCCQOuaXI2z9j+kqVaW0bWLk8sC5TXA4yLttZlzVjYoAqQ3rkGItBZUrFM80KT1dqg3
Tw2NydBePXgadjQZWn138xau9quUgUdLQr5l5Ux02VF+yvFDFuqZrCJCCJ1Le+LeXPiVt8nb1zXx
Po1CTmKgfFtyqZrHR79YNYn1+3MuvHrfV7LSZnAPlhKGnb/D2rPZ4RXR5EKO6K2m6lY/KVgXk/it
g47mc6zmbcvfH+MeMtoZx2tfg8zT6cXPBxpDBab1hqEczLzSJMjFTMMuIi9sBpdm00+2IgRlhM42
Q7bbF/TxrYgStNXCC7Ydb88Zbz2+5+7yznhgxa7XmxIo2u+6YHSshytEj/Vsu1g/I2rzSRIH0MvG
KIl2IFH8CxihkxM0LM5VKPUj6b36UnOLEQ37c6uu+YuPvT6PlSqd0EYnhb82ZWQpEAphz2nxC7L7
xkL3BgnYVzan/VDsGOqwkAhXgkHA/Rg0Yb28w8GGK7zk9DNSiSpm+vPwu4YoKEqwVMzOxlVP67zO
n4utIGn5C3SGerBcmC6ZJ3cbW1I18GMcsuivWyir/iecpFl3o/r76h4ZbdsUP2qEa1UUpm2/9Zit
f7DibqQfPw2xMworAUsPNDedI7H/3wBgkQG+XGu0S4j3rIpBy9arf65Cv1a3sDhDLzejTIkVFrZ/
ekytNlH8aTRDgUFw5eOVZTcKpV2MxRuzUzEsDuD69eNQINTC7Ff02DmdyiSuQ5/IYKwXmKa4rzsQ
uixrvgo0k5D/2rKhnL/7n5nN4/AL0exJ9+aLGg+6DOhmFtK0cUIkl2dEboZ4vu0cKjNITYba40cA
Qwxh8g2rstAHAMNTFjArWzuMraeKFjaW2Fn88Ui5SyyxDwQGVAVw56phxA6qtlCwbLeabqrEsCDk
a4N0qIMXACj2a6QkqrYrOHSPOtOqXujSWVTmoFvv+3Dc3qpV51HIEhxO0LLJ56htYQkBvK0XRuRH
VSQ9h6k00YlNCxdDJ/Y1lsj9z1gmDGfnE1DJRVf2iJtFV2WQbETwb02qfG87la+02FkzOfEbaFBO
ATApJc9hvHrksB/2sdCJ3+mbq3quUXRX1XZJG7xagmxWdDbLvCLaVq7q9aWXYLSQGf/izOzkjp6o
XC3JlTup8nnYt3En6cA7vuyJRiaAi31+5iKNOe1kfb3KBfo8491lx6zz2IkQIahe5n97+c2Kku6g
RQbAuwYYw5M0kSN0Gm195hYkKafrfCaEVI5TbOA/2fFn2hCL/SLEWUbvd89Mc++gJi8o1ILpCudS
0X0ztdiczS9l0dWDUhp/WhE143C/JUo5EAYxWj6oAVcQ2MrcP1E8K16v2wZx3hlbLXpFB+dtdOf5
lJGUV+WxSSz0vPczgsZZAz8a4eb6QPGxyrNffS6qQXnIhk9cOSjE1R9TS7oaq9ftWkTv8G+Tsh3T
4BJAMvESzT9k0mTZ0zaAF8qbJ64orcMU6EmZThm1HubW6Ix19tGnIz8JLYawLgAku68G0YJ3bkSk
FoymxR0+AtA9EvntkC34AgZ7wXPNBxBJ5tfun42P+OyvMKYpHLzXZd8qHekt697MD3TO+qv4etLp
KwrqQW1TqAk0Di8GhSW6j7ecurbr/hTC6SvCmhjckTRBO0tR5lEKGiYl4Eg8MAO5IDzSHQWZavIA
kv+itH81V/G5CXT5bBcSdd6U5LKalJMJxA148c1Z0swGz1F2NeBoThgiV6kr7hpVKLycnVafNF9x
GXbidApTrF7GZ3M3PiqXxmFPZvDHnY2slz99RxGKaaooIWCz4pLZ/SXRkUhTYr3J1mRkpZB9ICR+
lXPUfGSykBRJlvpF2cj+jdWTroUS/FJKUy3sgCZiCI3u+Wu7YA2vCIJiqrbYrAI8OXOx/0vK5ym+
ZpKjpLQf4TSAXGjmn5OKW9s+PmCmy62H8Bim7UAAH/8tqA2j/dIyYjpt8GUYJ1kn8hbA5W0/LQ4Z
j2EZe1vzLr02XrG/+0p6mHnnfelcWJNe523zD9D+Qzfc14aCl4uLfkIjI1hyHs7s/ZjCQjkB2Cjz
7WrZ/WmVryx1o2kW4k4aYqPZJOO/2puwnUNmt423a+Bo8q0+sTbQ41yM2vu8iSmnNtLT9Y2GDSWl
Szuz5RdxAhl+GCibRCQ+YuLrwhN0sXvYMdETBZeaysefM/jwSOR4uSSLCmkVyrq1vbPan+JEDH/J
nlVTNo6FDt2XoTV30KlzMer1iiXJEOyNXG/cm9Vu6kB6rd0shFFsH0ZtQfooOFtCCy5SQTg3CP5k
vCzWXmvsclCJzd5joL0EKqNkqoCV0LQH5u6Nqvun3GPQ3fFYP93QQ8UW4aY2e2PdJu+qxjhtq2ro
pLWODQRK88zoVOCIf38tHmeRBigamllAPZJ8D0ppvscLZmVPtJt+R5TyP1BwrC7LyLD7MJpcjPr8
Pf2feYDQoGPXAl7TrI0lcea00M1bXehO8IkPXsN86Xxyzkh+iv0PpqWHK6eoaFFbPyf24PZcXg19
nX04HY0I1rU1AlvNLPHViN6ytRQf48OsHHlJoYA/ym5j2v4+//sxAI/8e9qSqco5yjFPp2BsmJUT
yLRhC3vQcmsTXehrCCnN1Kl/U2Pxjg6zKWEFZ93vp/qDA7PzDzTKUHpGmE/L281Vv2Jh510KifDt
HwoIoTetptyiWmNybcnsXu2vAPTr42DGCC/P86r0CMopSdkKNCCRr0jsmCRyswwAX1bBG2KvYHe6
VfLbaskKGLIPm5uaW+8jZ3cNiev8XL0n9CjYv7TZMHCZD2tk8d5haW1x2uQGoh0adpYYv7wITr8U
46A0BLL6UXs/ZccxRJd+Ppd3N634iRupS92t37VYmCdid7rmy7TENe5pBLo5fS9ewk1FwuQjT5E8
b2EZr9Vw7zmfQk2BHj1be28Ss6DPx1VEZ8tSQyERgw0RVGyCSp8Xu0H+25uWU5kDTmQp0i/y1GKa
1YrYkdsxzxnv5s432AuujomcPXOPobBKGqZJC3BT+j1BRSbo0P5jLV6/CYNs3A8SBffh5i6GIHzR
DlrhdSe9bvrTXmS/z2jTcYbLYDMfi48XCG51Kws1rON/zBn/8LAmCmwxgR84Fd2go3ClRTi76/K+
EOQCfPTpkTpGFOpqpJvErXnrrArbVvLSSAFhAZUP4DleDr3e5MWNn1DnClOfGOxUqH4Rvore26fo
rfPGI3UxAOwEQhqKa1jb9aE5KVYnGdp/7cBPenQi2ahI7ESBj119cAPxQKYkI7KZBc/9el4yx4S1
zyY/InOl0jyDVSRuIr1fL2TSCsuDQR/muxMgEF3IDz1U7S5za+08U1ieG8dfSxACXwEk44tgL3Sf
vBARh1qydp43Rn1p1zYZ4j13HYlZcU0cwlDWQCt8EnFLcByGDWtKYV11BvRIAmJ5uxmu3uUFTFT4
b1MeGiRWvo2TWO6mEbG8YO4KjC5eagk5xjZKqftd/TXKt9d4D3eWtSLXDrDwiCv+Af8X6qjdX1z6
iI3BRHk8AxSf5DNAeE344ta/Ci28L7yFyhtrml4F0JvDk8SWJt57qgtxJcQP8Ld79F/pn9omx/CA
vwjy0Iu/zeGoXFCSxZjlXylLXD/Xaq6A5P618upVMrBrgWH/wtI6k9wCcBI9299TZdhFlD848a2e
mtWVGYh8IrJ9r3yFZeB3jNWpn24jSuNWgXUuNS03NUkP8ewPVqmXo98BkG1VdMiasd5jndzRkdwt
BK5LxA1drYkeXbEzGs8lJDtkQHG4CVObgujDb+Tc0fnFu3Nn7+Cj4Cs2edFdjRWRHGeFGSI0rTz0
JQCfb3M5K+xsQJL5rgBy8oV9dGnapCMuDzg6d7jliG0ui19/zfKYV+JEzedB+j4yRcjy7nz41vPm
nyJPtFY5Jddq1f9U0B4K2xjqssI+4Nv5XyNJXvSwf+kCaMeKj82MwM74h/NOoeGgDjDwExNlBYGn
/XPBjDKI0eNRxEFPVfDMUDsGXv41dTEL1dN+rxqLhqhzTHlETvxBL3NWwCk/aBHACasWCIMDbV9W
o3RziaeMRlSGK32qmOl1niYpuLp0AuC7wjeHQ2FUk/jLEA5KniSz/cRgpWoCH0Zr+Qwa1etDI+Ir
XnyEiinpDNLVplMSQbVoCsOsMzRN2b2DDtODNJdSlpw0HKx9GV+ewjIb4RwCHDIGJVVM2C1ymoI9
hf0LCEXcszF4RBfv1ZaBxBsmYAdIT+pDq3CQvQhgBJXyPWQnF1ONydNTkdicUmkAE7obhv3zfqhV
WEuwwPSKSvTQwbu9u53Zpdz88nkBWyDafjPBJy8f5xKBC5ZIvPPOtmmMcS+iS+YbjERq2ciyhFNX
AlI3s4leXKevsBcvbRVXpDT0mLxuBbGhphbtXIAtYZIxzb9xfkZeV2qzE/HOZDGVGov3CBMQ5K8c
LKXMqVleQWpl2AGWlbCfLMr1lzt1MEj4dikvJOhABZYQwwQPOI+06iQo54FZFvFaivtmHiSRwKHr
/16VmXssTJKib1u4DTrPS0dpzrh0Auf1p+9NhhY3fIA0uRg6OG8cCTGcJ4XB6DZmjezxwIffOf1o
gx3fXgBJEsumoUpM9U8noZt/9HOdjg+37K9tmxoir/8CcfNI/LdQ6tiOTaP6poVjG9/gKqbC7GMP
6zncHjJC6k6OD/zI3lmsqzuZr84IvYWw6Y/QEGbM7FWBQ4etmf+IMfk45VSoZY1TspkcbkMYDMP5
MVFXz9R7TmpS8kXDkMRy5DUjfKWf/OS1yc6H8QXEhf+7OX1UAuI3nIO3gxZHNTxn/kA9qQZQsaHF
9JvLM2vyCGjVXw53I6+uopNqAwZJ1Hn65VfeferzvFv/Z+NvZV8ZRYMMspSySkMLfqr5wf+GDc5A
g+XvYiwyJmnUqVh+VNkyR5na3YYsC1x4JT8OWT2TTk3lGWhe+PPI4KDr51Qy3GVcMDqDf/ZDC0fw
rh/jL5m34M8sD0pSNChNQObHRSUBCXDCq/SibT03m8DP0f8scL5uVfW9Tt6FIzx0QI7Y3b3n2DP1
dCVW2kkZ1mifjYpPlys/km57VmYa4mgkHevuG3ORqpYd/bA1zzmZxAkorUS/7K5ujtdntF206VZm
2MycwcszOQ8JOS6FJqz8buRETru7JUfW8O8WmxSlGfRZ8rF1HcmvU0pGNtrhE5Z1c5qvhxj7CgJj
sR2wiGCMzfTUOp+DtgFNHE6eWrdPRBJy5DvbCSHE3fyGAFPZM3c72ZI/k8/kOoUxFYOcm/NSSq9E
rK1CoyQDqB0cTT4AzgPNPs7UwXh4S8uxPME3YhGUDjrnjIDFsb/DfWVUPEOoWEX8TF0noftpzEAo
Mt12RN1S52bhRTGvcMmiJJUWX1GF0Cc58GKPEyPlYcEWYkOGpFmOpNUBJaBJ+RWQvSCABQtyUJeQ
tW/XTC5DUFoIoJTieT/6ExtNPSQPaYwcGji8lLwQx1SYi8SeBa14D7A0gQ0tAqPaty0ID5oP87Xd
Yb3oJvPVGlNaGDGz8y5vRlokE/KU5lLcQVZpr0y5OdojmQpB91pW4Kywxoae/KoYSi1CWU3unWPv
0hoKNnUaz57m4cDmy/DhnruvpBS/QT9RkqsKGEyJjjeoBmPTYv8QEh4E68z1qbxzhsanz/aoXLxk
1piOROGHQVnzPmkxYMDSko5jix29gWr6lkeCIHtniQYGs9zLkzq1Uhfm80yXe7e3BeD0Jlhwiqkz
36fYVd2CCPkVEdecrDn8LNQaIpCUszR4+/l5pe4mGBCQQ6cS1YBRAsik+HcYERsfR84zp87ZR43z
XZr+L2poXDfZPI4eoNs5BmtLvZS4wZ1nq6yIZN4JtKHMrBVyoAuli6bGW3N3nQsPt3nmAyJY+6fw
T15+Nf78K6AeQcfLRUFugRU6PQSOPVkrhhlyUUB1GxePvR/55r2YpL34Qaw7w7mBKrdiNoC1Fagt
7Aa0caaYhyapKZuJwhANM14DwMwxysK+6qmvftf8IqRpco5CDFzBCIoTLaRI3y+ZZ/7hLzmXKacI
TJs7Ja82D6BV30dOkDrrz9Nqs383QKo2+msxNTP3f/7k5i4o/uqGwFxfQJUhETBVZvB6CG6tX8q9
oszKOvoiQdeVH2Acno+Le/89lD2uA7Xr7Ri0bTtgw7iNyUACm4BPlHRbZg5fiu8BKtvDu/VJN2+V
JzCnUoR82BKuteF3+iQCm2IWaAMdFSveQ3JkMRC1yIcBMj9D1kbI9vY4DesXH5KJqFWmKF7Sk0Yg
5PV16SVU95dx/nSDZX0nHXegJuE/MO10C3mUck/GvqRPdb84iGJs7OrUM1bQSR0G67KziTkm4UUh
KsMeLn8Od5BqRkLVS5+nO/FgoUUVecZnSXTMPuUvTPsqmAqM5y7Xcl0fTa5Lqy36guNWvPfbMGFB
ZaZ6v5lJ1gohWSxLfN/1jAsD1Z2RfTNg+qSb4qHMf/LSitUxVZJxx/UJ2OP2uulHyp9PSViWtaiO
Nr7vXsVQQcFVphgccMHyEqE980ouCHc3BEB0zaB6SMOglnjLhPIj4UOG6EqTp3BAm/qK+2hviHps
d7vyl6qFzE1bNKYo3io7Ba+FgqXvA8lQwrmPjlZxbXmIy3yJgVpzrDc8qgjRyzKvZOXVOrjVRdsC
KmDJcNMTozUmc4On25Dc2Olem1huPARNLufBAdkapJBW1YvM1wO5/ORAWcHAO5cIkvF7xQvAsgNo
dusYxWfPjVaW0xw5T8aQPxOGkfrjoawM0IUHI9lYhmuK7JKk4kwBMDD3MPNXTSS2WmYJuAvmfMum
1qzfY2pgSNYhT8BnnJafkuQKvXfKExI3ivLIs8HzuNeIH+WkGSZ7QONdzJcDuUy7NHec7V8mYjap
bO3hCgjC5T4WV/k4xitOIE9OI6oQWwPrXbPmScq2tEEIy2pmUVw04hxrBnuuzzA7xga7EWC+HoSy
AwwJpncDuBke2Ypj7R8aQ6Xs6wfAwmggZ8hTWoPR7JhIIprTLVvUr3wzpJZsolvZvsh7wSkYmtwm
fVGwBEJQRndg8AWQoNv/ZLUaL4gYq2yrlMUstxCu15bvWmvaUIggMwRhdgjwVOI5Y/2zk5OGORuo
z6mcJGSmgHdc7Vj8iKcKdy5K7S/VeWO47gWzkXin4bENvtom29487UJmPH+rDpYaSpnjNaCcTe2U
d5ls/DEXcnbpGeqQhVQ25dN5wrYe/RG5Nb6gDNzeP3jpUZaLwIP1GTJDXZd28DaLgBfpbdNN3u08
Ua3F48WY+b3v0yWaD/HJs6CouLXBYDfiE4GRUk4SvNcy9evhm4AJnZPKaR5u/ypnEqLyo1s4GTG+
KJkHUmhcrM7rOVdhu/syZbThS8zZQtjnpcBZC7nmnViP+CiAmQmEWhhERTFu783YVoCld6E6NsMm
G/339XgIbWggjgQFqsecwZWseJjnG6Ot207y5oP4RX6w0CZR5fKYbsttRUZSObZbjXcT6D3w4kaH
rt6ZEoBjzKXOcMSSczTMtQRpRCzUHWrDPuvpWOLbUldaPNfW2OB91f5ub3I/UZBkg0FpNfnT5tx3
F6E+OKyxELqGLfBVyGZPZQAYQDiZhDha8N+dvwVEJSUDFXZi78m7ypdjDTPnmKjhXmK/WdqksOxB
34A6TeHxSuaxvc/ijF+utSaJKCfBu5fUdryOySNWmJ3Sq0a5UkjJvyGWx8axQLDjKZWyEB9afMOE
HYMsfhcrCTBLbXTE2jnxoQUKMcSskCudCL2lK81sm82S9gHzmKoXVYthPHBIQd8puMygeCv+TX0c
zQc1lGMa8eBv8hdyFu1ADRRh5/pl1ZjE7DV0yaNMLDwQXrUTAdpH17H/z3ZhYdQJJZLPVJQhi1AC
5F4dSygPEXqDpBD0b0yOy5a8OLn/5IB1J+fnsc45ShdaTVaS/dDNmRLe9mBu1tsXq/sl6M91/z9U
GXC30y6KNykGdi9ux+25hOY7RrbYRDhq1s+QyoIdlz8BbTYYSsk3ClRlnsQLBSiTc+Q33+Rl+d4h
lKahGQcx8DvqpuoCIpZEa4DGsuuHB60Q+c2Dmpbph4mLPtlgSsEeu1vnZ/tdKMlFITTOYDwNFtIe
5HaQc8y6AFuLGL3TpV8CKz65/U1o6uvEZbuUYEhMUUuBPC7Nl2MPFKZmJxwcEPDJ0JKi2ljVUE8I
OYx0Z3mTWQ8z+M97JAJY35auFBAB597wMSqocF/cyyHDH1tDTVgTnENR1+D7IN00tSJo1JsvkN9c
ekyTIdGL0Rm487IFXDnTiNcl3qX6KkjtftzTWcJ/D27VCc6WqQENWtMPH15fRwpoXvHx9uqWnVMG
AbD5PUXbBYuBdtBlIchxBVIlKhSiQh0CjRkFkiIqP5RGOQbq9RR2Z3mN3gWiqCEbiz8BAwr8GyaQ
XjmZE1Vx5AFQBs1fah4Q8YPST6A+cTcZA0OLox8iFcSy6Il+wpPDdrvyfzcEGf6re0FitDr8dPaC
wG/zngdzd2vXU4h7iGlnUsAdfJ315yU2xDpm+XK8Yy8CjgHs4hjjLbdrBE5nfubCIA8B5E1i/MLE
S7X3lLXVHsH4G36Loy6Nh+yO26Za1tOpCJlZKO4YRbxsjhrhTC1TfhWODtWzeMut67hd9fDrPQ1P
3xGA4rQn58lcFSz2n6Crli43mw6LGNGYVllpKA5CAmu6hgQ6iRUJpEqdOgmzU+J5EltmoZjgxUSj
hmqXdcMtLbu0ljYtma15VUZcDiPriNBQXP4HkDXfUnjK6IL3mpqeR5gxfQ0JTDWU94YtLyhEc63K
SVinug5XwcAP99WZd8YGP9d8chik21HFAFA7C9FrNKCoPTYAgicJpovCcFNRh7QIy3mBky3Z5EYO
Nn/IoJCJTsEXnks4zDxNy2YcOp/025YRtkj55Uz+vLtOg4ye4vx6ts5AgTzp7digFTCXCrz9+38v
ntrhRnqhVA2uGvaW4caixuhyZ+3rVI6i2pMxhBV3LczBMRMR0k2uXzPvOuWc47SpGjBMj0sRs/3H
pyzBgP2fZlxbj84ejFi344/OKr0kxHblEgOjuTSgIbt1goSTrbnh0hZe9BCbWOO5DlhDSV5TTNOR
YauF2QhQmyMDSxk7SIMOVvOc0BuHxy5MaM1SqUbJc55/omoGd4bNZZU1eBpA0PKVvI+zot7Fc17g
ezfAdV5b4kRKf0BDzqAlsNZqk7MgP5c/IzyZOAXFNf8hOEANRX6L7PifA0xkdodWjPOuNNGPt5z1
r9s9gvBpexnIOcHoSCOii61sUs1PLc8t78DuPMWjh5DVB3TUs4wSNXwBwpE85i/VnkGdetDKYcDS
MwkUwzOqWK3XVuQ+dhMbHckhnNBwVpkQO5niLJq/Vf3xXYTbVO00fAuWChGfFLSSAC1oJ3h5xwsg
Zv9j0GqrV5cgTYj8/qPl8OPCqOwrjJlPUoxp2HgVN4L/cdN6E3zhFLKQOU8352mYmgwNvq5cs4BY
LnQNXFvHcHfi2eRS1G5/8kzCmwwRALpOXI0V1aAbM91m4HE3tUvwIy0mT7Fv52bZckZ4QIYcvgWC
OvjXCDtlsn0WOdt+zK4CHybwhVMkf0+AGTj863iewIzpQCIFTt8t6TKcwzh09SBCOu62PndIMxm8
HQTNl2NeJMg1aKD80tT0d9mPyDI+qiob/1A1kN+TugUNuGjdwGIxQybVF+b4RldpsyDmAkRTMi/y
QTld/1kqbD5gd8DeLDqd5lcaXSBENizLXaUG5OtiA6PNmBBEM1/L72JQY/PGv/Q5XjBlRcnhfE8/
UvGpqWDjvicdZLFdeUC9x2JzbxM1Vo0pQMHy2Z3lt593IxZv7ddNWJcvjMw2TPE8PGEhB181jNCo
cdkRBS/yrHHxnjDxxhtoFVsH6E4ZcKR0bT7n+gAMP/0iIuQuGNB0VxuuoxWuY/6t5L91O9b+YA01
6laEoKPcfM5gqC9YCB5BEmT88z0kDVkuxqTTbqLfg0np/QI5KbVX/q7nJu4t45g4vWJMQsCDYcPn
ehRNDfbmmsFoTaJb1rEypfpOt8tu3N9JZVWvos0RFR6Ics1OO+P/xRSe/GHu9xHVb0zxS4KgLpd4
cXzA2htPHrLiBbTEgMI9tJItWbRLq3lJtWFrNo/vkc6xAtZJ5XMLURHOCMh+nQfSZydZ2gDaQont
nPDMfSC4lTg8Eiujp/IXh6gOpSHO8iQSgs7O+pZV2qG1ouVU2PUSPH3frPfV0vXfyS5QPSdETW8c
R/hIE2TrXJorEi+IJzwX6qfoCedxI6Qk/O51ptxwG7YlDhfFi9H1utwNxak/LJh+sHMYWR3GP1V2
E6j4Y1cCOUTIaPKmDVwCRud7F1NrpEa+ADX8g86LnjNQKpL38UZ09Ipasyu647/0hty6K8SXTawO
UOftqWcv+SQaed3M5R7Q6Bx5Xc0EQl7CEKlOC4yKjoYfMZ9+SLhwRwflLVL6csChTiFvs3P78cks
xh3NeVguoxDCD8BC00Wl4gKkhPeVWo8QREBcZ4g117kK19Bo9i78Pj4OOA+49jAsMhS6wjEpxh9g
7q6zc5exXqNXUVWyeDOLuyetFAPnLRzKlVovotl4J1kPDs/WeQ161w4TLmt7BQT2pNRiAv/c4DdF
aeoU3PSkUvMHlHUtZOtLQmWyMUTPz2VbpJ8Patvz6B7H7nkqf2BRl0GZiE7PIa8V2ds2vuLmp7Jc
3GKMVuOtlTak6yGpVdxl4ahRESjxR7SJotvhwr9K2IcP/luM+sX93Zft+0atnoZl/F+m4vAZKeg6
jWDvBP3NCysI+C9iUGuyDSnWq3djbFokacQSoHEU0z3Vp8pDkfY///9y4IDCWsW7XM/vjZ0Pw9tG
WWnvB6i4PML3wEfoVKTllsmLQb89uut+Y0c9e22z2XT6UDHIDULu8wBdXpEXmBQEwqnzPI2/m6kw
G82ycTiv185WUBvcm5IsdopHaJ1SEIFGe6EgGWK0xq8QrUtRv3eBLJcyQLgQv8EWAFEhv8mMowKi
gmIwKcV2AASxmT4m4dV6hzkzsHjcfGsz7reKIAzCs3KxmVuEkHuP9ePm5LbbsFElyDVao485KTf4
rULdMYMEFrCst3fLYuhiIYG59gKuPr3DGuh4S+HKMVzJ9wAO6ymUcoieW7ZmEb/ROnIxpgj8tXx5
1mX46AANRfhDRyG3O3PahrhU5CYS14yVDClMuuaSSzBiY7alJCj1DVIk6+QzJTFKd5nCv4qwGQxs
375RV/rhT0DZET85KCUIsLO+6EfxVOGwyd4iDltHb4+6K2dfKIDPF5qkvTSSPoUYMwMubaJaz5/C
NdIPJIdkU+MBHYQ8VPNp62Y9676bJlz3U1MPKBDwoCBz1rS9ivYsHOZtY2lL64PYX+vJbd8wEkZP
FoPdyF1OmAF8nr+4xjsxfkpENOm89p8H22K91mcZxG5A2wT8+zTAyW6j2ZmXbPXxOSZlEvX9pWP3
35hHpZCGyxxp6Jc3RhRmcDgzEu6zCJ+zBUZ0/cA15+7DJG23wWXXhHkgx2T+97rHwgd0ZH2dhrh/
D0XMh1qdrJ+3Kb4xW4G+0KdxW3JELm9KpIOKuH/gxuHWo+P2R0jdHHJCAcFTGWrIGeulwoc2L1gP
K6glNHKrcvOGeMhIgggKSWheZCbasdjZDaEXmsdoWPByjh0viTFlVPeK2WUYdt6WvLSfLy94gXIZ
Wk8DQfahXvzXMQuBwKGuin+XwtTc+TR6SBtnoudfiGTtkHXiO8i2FLKF7KjG/VFztpkgvRQc6aXF
f03p1CW/CS6AVjJHDO/6d3DBtFms5bzAijtlGNwyqB9HEGQ+OY5mDw6DRmpqL5V1r2NnYTPtCVG2
lBJ8KzIpwqAyoSSGAN0Weaj2s7lA5a+W0q/uxWRPPCOulIY5GQUNXIzULBRFCqMzk3/F5BCaN9id
5eQ+WmzUtFdET/8l4r9HBleSdR1QchRXeFhUe2n0+LCXhxHkC21U367xlduOOXEL70JfmAfvCJuD
5LIeDvgn7vkzfv/XvvaqMca4cRNW+FN5tW6Wdv3Fj50c9aKFhwQJSE7ID05vWe6cWnruUdQDmcZp
Z36+WvmxxSYh/TAzA7Jal+hQtOI/WtaXm0PUcKz+wBOBe3zk3FrNToBUJcoOIvGUO+D5KOKx/zGB
4h4E2B8pJ2vnf7vgDy1OBki0pKMUPSkEoOkSYt//2EQXIiFq+aTzpQjzzyn/KiKzRavivfAb+t3P
BLxwxJfAo0rEzaPH/gjWjf/vOAzM1gJVMyzaYIDOCC9l308gLgRrk++GmkGTbEasTRYjLhGRLRLk
Bl49QGX09JSgG0YsIB90X/tqwLsr85blwqWETCZtNx1g6W3mwSY9g1SBNTkrG3v2Zz7ldU6lb9bB
szkJsw5xiVWHJ/KL+BtM0sP43S3lZ0pyRV0zIxIi7surQzktJ4nzeFdua5oS8lD65wceB0tuxEYD
xOT+hJp+hX9cu6Y47KvoxspOxaWmu2JdecpEM2SYkTURT20Kg6LY1HkLdsU7ZsEOvAuCkUt/iScV
OjrEaGvSzdPrOJaRdECQSsP6NVlK9HJnVr3RuO3jRAAQrrXy2uHgVWOp0w5EkBpA+v7fFNhWEAeH
SZ68+VrlEApMvyf/grqpVj7fn3jIC6nqV8+yl5xTj/fH+k5BLLMRDhJUslF559F83sqdZbuh8JqD
MsZRXHbo6qS0hirRoqICNDygWsYVKPqGJL32WhOZ8avmSURkC2yFzLimkWVqfhNWAtX5XiCk/2O1
23x8IlBiiN9DtAxPi+WHh4N0kCpBnRjdveNaGz16xOtbzmlGrsITYeEeK8tZJv7QyveVBdr3kKqv
bd91ZJNdzKu0G39I/9NjiCzf4GfzSMwItV91A08Aw1NIj9JdHiK1psORvsVO1RrnuRVIoh6xFfE4
fbe6l/G4G5d62b0oNseWi4Shv+a455hSdg4hvm0u00BHWbjSWuEro4Km8NauZV1lP70hKLrAueJj
odnKGP4aaBOiubHebCZebZ+nLROZDb03ZL2UbGDE34bq3ECJ0yii1K8Prz6keTJ2XKRkmDP+iI+c
K8ranPbHCg9spTfleS+yjFGPb9qtcK+aKe7DQEMKTBoMtoq/wyfcBac/Aba08eZMfvKix8bGejJE
EJiw1YszHU9ZRqL1G6gLaOsCWK/vvivsOErlbecxuiuW4z0Ts17jGph3y1v45WL7JBKV0onkx7iS
XvYZ3SGvTDJoimRDtOGTycxvnEVo6IJLV8ckIZMtsbsoboDH0XZKHMxubCZa5nE3Mg9sN9j4F/CB
wLvJTmSvkGdRqTNJwSblINyAbSO1zoUxcAWZUYWqqAYbmg7ACR/gnVBgNlzAU8u0WBQkEfGBy+BW
YhUjRV9EGqGDhnjiOlLMUjX9QmFouSBsbSbbUrou0oeSOz5DdNHn3ZtCCVDEtFVxVEYcO/I2I2pQ
ajPIDpI2YlBbFdEC15LTaUs0MLaQBC54SHbXu/kkvO0+hq0wzh1Li87Y5SFw38XFygny8MOuiUfN
0dWP0yHToGwJ/uf3QSEdEqGISYRc7FzVlUYwGKemFTWDmPbstsJdgwsLkM45oYCZbT7M2hpfH1Ll
P1QHa5ZI0oONwPgT5TyHnXhPCfw7zw+O5nb5EfCv4AkyTqD36Zfdmckg+9pZtHJ2uc3H207J4EXn
tCx5HoR0/z7qsHCQbnYG43u2g23/qLJqKS+ddw52MuZFQSUhEjdWibVHfbiRQ2zGsIjIJ5N8B+Db
ZML9g7t1r9bSILEUePRwM9oNUX9k1H4Ze/jNZ6jYAJAf0UmnTk+IRwcOEYZ9PKKrEJrenGX9CMjU
9fasw3+qk0BhRnuARSQRph2pI9lKP3ZKq1g+7j1PIATVbG+Ms85JinIhu8bpGVjSIRdcUuDJ1AZr
mIT2IPC1400io0jM85KMGgdM8ymQLDI7ZlBUGhzJb5/G+3TYQwC76cT+dYwusa4qe8jj3KnWaiXW
OkivoAyrQtWgJnCV+uqBt1iC7hYgGDfnpxDXBs+lw/ci5HPYlIMirvkLmd5cIxc9/KkXwYt3Pq5Q
f7fX0R7tHLgCLOvGXw9JErIhmKrD5egrk7EJCSey1r6PxOp2ChUEQVraaic3aISo4SgScItXynbD
p9wVuZev9QylFn3MayIxjdSxqLPmlOa5wtgSPhK+BZiQ4gDYXg5KNpXD0yOFG9DedzcxudQMOCZ4
OaXa6wR90IWeVXKAcwWwSrdbHrcTM4DmpWNzsv08mkFb+ZYLFg7Swq380ZU3Z4vi+VUBoqf/pFjC
kthRrhx52zD7YYLw8TSbhJWrRKEyXthcwQubM84dhdjBj5isw+OE5n2TolhAt5jPOEHj25z+TSoU
cACIFz7/maXPFqunlQzQVgsVKArh5YtidgmHOfgwMS2P4Rm6sp5CHfp0Ja7V6SdZalZ09YvLKAcl
aTv1dNJps16F8+hWtoL2In/8ETVWWsRmNKyRYBVsQXH2sXHR+goLuIH31B9LceoEPTp/YFDMSLmw
bkyTJeFoVHEHYxH5EiV7Z8btKRYfDPp9lyP2DLG5rTPtz+Bre4iSQZN8RbMHusFaB2EZyx1KWQnD
LwZHpV3dBiGMYGSoxcDmytRF3lkXQ3UoNfWVnQ3iGTB7001+AAEO3hNv/VqRb9gLGWwI6NZMTNWq
QjwQOgUFlYGzGtoNPnG9kJDyDS+fMXbgMDJlHJfCtzwWxP+gxvC0713Cg1uHPGE6hetI8gZXXTrY
kL2+SBwcoFBP7SgJIrKR3MsVtb4QRbGvxwVAJN2/dyKaI5gx65lM1iB2zCM97uvfoIK7AtVEbiX5
/Y51+VJUCWi2JVUJjJbFjayqNnlCTorLRU+tx30XhDNkw6OjugKqgEwUpMH2Kkd+OlqY3qmbt5sj
CONJhqWM63in3oNJIzGAPTIZfXx1wYf7f1S3Y60cGWMV9cReajTRCklZjcp4OPFCFR2KslG5rR48
DIpFvYmKEQskRd/UoLmKKzhY63DuOLEVz/tRqxgRJiBV8whb8RD0oHajlpKp/qmYpeHxRtC8u/+s
dqWYc2fZp3QySPK0VuWSdhqrm/GbGLu0JhJPfQGwcaoVtw/5iYQiXL7b0az7qsL0iHICRwg/+M65
0k+7YKAylo094izZ0Tt0BHDkUL7maZgBpWajfJhQGmcytlW4veMwux43gIoBmqQts/ReMaSlh2T3
a5/djSEGdjYRBsqrkpIAcoj3smy4JBd5bEXEdcoYc8ZMDwH8dO7/yPa69bs4gqhuvyJHN1ljjZoi
XlQV/4X4uQJmwakSFNVxniCAQUrqOnHORmQzsuzfOC0wNkR207zDHhY8OWsDwMIU49Y4VVMO0ScE
iPkWQuzJflpEKn030sP5p00SSbxA2hlTzLrFQq0u5BHvan+Rsl3AFCCtlvtGarF9X3nOIi2pBilE
NWpbDpV4eJjeNhb8eKQWRUq6hDkIojBqGNTHUYs1MRkPFOurMnGji0F306alRnOoi4XD1zQ5c15q
1A8nW0qe8JrjVW0amljQ/zNJxB46AUDE5TIBbCbDZa18fS0x+mhggwuf3ZoXTIQFlSI/rL1nLxsp
4w3OHyWaWDt+kzr5XfEeyeXhCK4j096SpCC7FKmQxLN71Ab9z5sKQWgmlDGZLJLjway2Dnz9upQL
edjQSjs2qYPz4iOeDqvFraycWXloqjf4SKDScy8Se9cAP8HoN84MImC7jXz70k7j2O+7bBFwJDde
WqGQXzgwTBGYAP0JRWpZ4rdCiEc8Id3QUwOtfNdpMA4ZrKSA9wR1dSXoBASldPT6ssxJVPjLhQ8V
sBPb/VCgiQHX0pvO3GDochJTityYskx4o0C7TZWGUvqNV4LlZRT6k358UHGiM+E6dvnAVo7sWeCA
xdGGcWvJoTchk0lpWiKTnMAzKvBbOJRJkZfZmaCPJL/tec8iiPsTPfrhPwC+NDbFEvAcpG6UvsN/
1qvZ+N/8BFAa7rwrDUvgg92S5bhbDYVWEnI4FV49WTRSc+zUxBXaLvXmSbte4qOJ64715wG46opd
lW4rVijrCRvndrvhPIqMMkCeo8e4kIEJrCcq5ggIGh3qgnfYNf+fbeHj1w0GRcd361DlQALF+l+L
r+Xqe4rZFuA0mRQMxegWEC14o6+Bt+lLeEMefahdRTXsrSa2V14YUgd9HF6p08tb7PW6blX3IAS5
tJV5gsxqlvrXlviXOZDPKnAXqEYSKrK7eDNJfo3xZgv9jqXwIx4CKGLqYtmdnR5OIc02pWqMCpfc
IMB5CZme4eC9zPkf52cH5GAgXEKDIomG0BBYkBMadeHlVGlTdp10HMyBUt7QqjtDELHCNd7XWxQk
LHEtNF09RH7Lxf5QuPrC6FPVYHgHqVTO6ck7Jje+THYoaIQuIWFS1y9PwadbfZF1ryZrI4b6tFGz
B5v+wQbY62t1N04O7YERVLcCeCxG/EiU/RJrJGsDmGz6G/VuEgi9LT6Oq7KNktTXY6oqRmx44eQn
nWayJW/noZ+APRn+mHMVhUyejMVZdAOKMFh49Horq8pw/ASEtlLK69t+xhwpx4jGFwVyqIP+hr2D
V6Ld/ewEgLBXlZOgvaA/IkgZZ3aqMDY9LYQGKV6N9Kta8s/hIEb5spkUrRQ7ivXN9GUFbN5xMW86
hdbsuMAcoWISwTEfo1h0N1NtNlaYJ1LbRMFuJfh0bRQwweaWqKbcYDkSRDFt3jts/2o+ftXqEKTy
iga5saAlPCnDeE3U+I+x3vmnwUPNmQLJVaS9LVKnQtMlAzVqGKta7dE6YYrKW0yENbuMoiK6BUHC
CqkQnmbwin3obsnTY9ZRVNCAO6zwdQ8PajHw1fhd9MrAk4Rx3f3/uAJTtBTPc2TGmatoVjJiR+g8
w+tbN5swZnwmWUXoYD3wvroNlAvNw0lEmUZ2aOyvGBL0WfumoqSbefv/WWsohaGMr9kmOVUymND1
nfHVXbKZblWqtc/1dIRkxT44A5rdTTGaLZKb0NC36duXeDYm8W8RD7PSHJFOfu9+y9tBjr+RNk1/
wWwEzxLcwTTJXg26CPYCb58KLsMbVTLzG1Hqriwf+OXW/ZTCN22SJajcKpgyzHdDYkFweCf3ngbG
/E/4tnCWSFSafO76Qli3L2/N4RpSMPNocufr3PgG0lbDaMb/f0UGFSkSMBhNKz47PXF+6Q14c01z
Sp7oF4SpWUfGMg8ly5Ol3JTh4F8aLZm4h6v41BuV4QrcUG76OKA2g0jFYxpjrRHTKWcY2rul1OpL
38+LGXfHI5drDIjgkN4lS4jy+4SfghuILEFhqJISj4q2TWF/6obEOKy04EEEUU6xRpd0XYfjbnXE
e3HSMekaHK90MkBTZQLPqiwCz5x8pyTyaXvUkaidmxMnCzPeszwzXyFzCsgZhkp7eU1xoyUs6pms
A0gMZSEOH7vlR7hCVtA2tiGFuLODUjSzO0CUgQZIu3oBgZKWoxEtzGUWjJWAw3eGnK69fR/pS/nw
S2bieDJei2TwQvmtHFclt4qcX5aRj2WVfYZKQ71qVrSZMgCkEJM9Phc3xtgcc5BQNWuTo3FzG8Mo
CShhPCObhEp0w1mbFvZ0NMfe2Fq6x/TynYYnXGgafQ0RuuAAbP0rBLpZtgIkFFxLPUTtvQuL+bPB
NeHvw5e+AACfF5LplQQWiw77WGKSxGWFXpkJOJGaBjkjnYkkGQZ3P3lrwEsD9XEw/QUfQTFIs3gb
i0tBdMYzU8uULSkKD7rTVrNAhZl9pv+xVpTJm4tRMh495PMQIzFpK7eAHtu4fM8+UnenQWa/nzqs
H6HMXJfaShLd7aEgo5jYB+mVN9HErbmvCZKOyo9GcLMjW9Iv/CYwf4twCXiDTkDAkqQBaW0VqXkI
YZr1pa+XG2HAXXKVNjEru7vEBwM7ToVsCsPhCw7Ny883ZqBCKhJ3EwcfLcZe0I2QWK48kEDKA3wk
sPH3TtaWCeZ0SvNhU5it9k5lxWccElEyioomnO6/9Lom/CelZhXlBFK6Nd0v7CbNmaBceX5klxdZ
xLJXHxDOtyb/2j4waQBcsSDUEl7YoAKObh9K3su3e7ObL8QxKfzxG1iV1ptme04hpiR4pul6a15p
OE0PtzjzdNYb6rKCRpBUsM0tdwmb/h4J38yLufX0ZEM7i4CJeOe8BcDPf7t4T3mNBZBhClLzxgLx
2iwUhju7+BIY1Z/y3TOYmjDgBYKp5D8/X/ajleyghDZGDlJEfCTMTTu0q7bu01/1T2GUUdyvFtGY
lYN/7ufbx9errTBopGm1tDqowOhVdyqxJIAMnUmrL24Vs8RS9kZtfQx/K/2wCAy/U2HGRz+RgxrS
12t3HflNIvev20tVcGhfGCyQQNvlfji2SwmUsq+jeBNyum8p+0K4Bv4e1Y/HSu0IjzUumVKigSyv
2bSWO5bEv2joBZQSEPeTRAFabMZSJT61xwoOxISGJTOGQuI/iLocrmIIAnYB2W0e96SudhM938a1
Aztbtd8ubvwtuIWAS2k4DG1Pt2wAug9sSgz0aT/fEppAUOqUwjA/0SqNN6OMCzAtuKHFF72EXqWc
uMbADOymQQYOmK5A+ITWNsjgD5jwDLIueOJgskA9mM37vgJMhBhE+oW/VMWvdAMTWjEWHdoYXhIG
hE/lm/qGT9OPvsXg/42jZsfXiVi6p5VXsrPSDiwLdXZUtp06sO42UGsMzSamStBDg8gE0sIOqOoo
QCqDpmbERScFVpsxrJEwbrnst4b8yUtVaIVDikNdW5V6kWYX/m8HHRimBM8EPzbzx1H9O471bAzw
5CfKWME5hCqm69ys7jbGI2AsqrI2j3uEqaFtZgShBb3y47s3dw2VYvW0bBVwhkHC/3FqInBIMlHi
JU9FqPxAIcCzUGMNxmh+ywblnrplfm3LwHUUnVEA05w8y0ngmyK9V33hOb753AQGLe+Ct4LK4SOV
wDC6w0RG/0sAhdNHqNjceZwueR0o6/MzE0TlkrNIJG+yY6nptZkaF19p+dEnyrYX9YeXw2DGsi/5
XmjXmCTpN1NdPWWCFXwdznQ/Sip616Pg9UPHQO8PTlz7MQKjcGW1F2LwMg1GBj8zK2SKaqEKPBKl
woL67D6xjI345GTGKl/ODMYhh4J9C2U4i4LjCJnO5ooH4Rf5M0mgFkB4T632uYFQN70PKY6PK/Eg
npervtVtmc7QyRduTusu4LFWMiBtPplQbxL+6FEOe7WzSdrlaehQVjSiYBEn6FLurr4K8OW9ZQDd
Ge++5XIdEJLPxrL414w695NHdYZ8C6w9eH96yo7kbQYlNRVStqM5kaMSK79L8gfUhyOlr7izMv9v
cSA7hXNxuB+ERGmEDF2GUvgsHYKS0yfpn640WngiKt70E79ciBvDM0S4+2XGiRwdBnEoO/qfQLvU
32cS0B1V3lXCKgRK/z8xUdnu4clPwj/8RfF+CV6oral9zj0Lgnui7HBFTOuNuvLOtP61mThCe2Nx
TJt4klMEAqlFbbjfLKIEHydcNQlbI/uo7e3g0tXkhPYXaiQOy85KdEcDf599XVtkds2GtG5DGJzn
qlruBNVd9I8AmCO6CyLkPCWAhVIoMT3oXrzqIrIUjPRhN4cJ2ZXcY5D0gHfGuZdQ4Dad75juTscq
RgNp7jAjQdLox36K3xc9wgeB0JmiwfqCBAHpjE9Ur/gbrestL32fLsYbiA6MKSfDz6lv3bX/8pmi
746ioREpIT6MQyRn7rhKp0vI3eFulD8D0hj7OywgMbXi59W2aOSUSJ0XxAR0oFZWn0qWumVtW3tu
aJm0ATuWWZQ2AMFEPnjJJkoGj176gY2mizzIfTswd43xRfAMVlXledJmGdR5vceVFSqKEK+EFqWk
Y++zUIPyx5Mn+a0f4u+o4xmY5E5bj4OplhPZd+iP5G7YD5v30ekWwR3nTpIbHVpbjrNDI9hUgjVU
ZFnVcFVMJBL+Lc9vquS9MhRdBWKQg0WuXfjaPWXI13OFqbQELNkPMJ9Y1ETRH7E3Y352z/oXP1dl
EFBErqgLIBdWWA8X+BRVXVdH4ZxudpMa2+E6s6JnxqH5XndqwpJFa87GkNWtvZVa5vEijf0TCbGV
td9LRGt8fBUUQAMmH5T93pwJTzMNohF2Wnz7hC8jbWYsEXFhIzh62aD2RXGOxjnYgLCpb5Q6E/fV
Onpbn0JjEAZ5NjraaXbUk34uJI2zKyqOzi2jbYf2XOEPyj8O1BiVkC4//u1wsR3UOaSXZ28iYIyA
VDNR+JZsT/HOs4u6EsnlNjRhSwEVSRrDwOMiGC6yoy7k9swYmRHrIw57IyFBwgp/iMbjLCHaGPHE
XDLOY6hqjFRMgWPdiMEfRRBtAVwvmCEzrBPiNB1P3fTIvDTce/XBXK++YEoAXmOvWGoc7VWqzyrC
w58kPJJl8givyVWMQFG4ObZcfDaBwMQRkFwX4UQFzTWEkd68a8HD8H/1NDPcmRqNsVYrX+Uh+O07
FVLyl7T+HqZyDid1xGyaIX+vaHxUiy/fJ0OhJm89KPGWowl3cljUDTKxeKY7PoXc+3d5+zspAi1b
aEl6Yl8jx0JU3+ssRvdHG0qFZDzJHSUpiFITSCHeYIW98UW+XrzZYqJXWb/5TiVqw44HId/+NlJh
ZYZkAniiRbXZgCZPfUBbPMlioTjLNIA1B/6S5NqaDO6W1Fz6HmZkgDpuGMgOGR7dtGxCtsQ7X1+r
HSGl511fPBo2H026j1xjzte6hQ+BDe2O5ZTVdjgdnHE65RfKezKj6plXIo42oHvWudWLy5SmqSjN
exaWspKZEg0v3sZLWfxcg8CnvBaVAtBDVufb67IfhKShAFhypMu+d80WW0+EgifBO9xg94FLTbgq
lKe+DBchmrTkRl8DsG3I/yQf3/5/OMP1VMSTqEf3qSW4EfyP/tAnKA/Kfbw0n9hFeiO1k31Wxs/H
wqxhBqahZi48dM2Bo75wcnKjdqI7wR6u7w1HXru6lX9oG88dHjM4JM42IlpkxdZkcbTnlZevqn2D
yxCiAK/f2tba19CmC0OKcZ9qbEUuPYmLtlDpBxxP0/7zVCf5rMV5noGw55QlPujaAjIZ6hLuwWxP
2wGJOBSzbu6wXLGbnNWYh7ACsVERb0B1RKmlVU/Fyn2P3yfUYQySMiGgMuj2BIL6Kz1VXhjJhb83
ZOYufBKSLTLumy5f5GXXz/e0uTiX/lypBqvz9HYbfPLCaOx3mylG61O8dzuRT8/ZqhhZzx/LTOTl
KvEbKwNkYsyCr/JirWicyMJJAbHODP4k5kkub195OTCU1sNsz0s9/WNBRdaW3oMhSiRxiqFiB3/4
KcyyFKOiAIw5c070US+dA4kNqRwo0obyzcA5z/fWvld9h1vFC/KKwt6812mVmYhAwoGnB8Lzk+2J
HhnNV/8Q9sZRk98uiLght00XONyWm7ZiibWyvxZa0Q1DIU4Ny2Gxr92oJ3dCGev0Zfm4mQaI/ydt
A4tP4zqaP3r5lmwcITGY1XHxHRzWud8QMPlY7es9/V0UY06qgCfMV1n+G5qcIMWlStv6ka+TRJuZ
KNfgAvxc68MP4cSLwNks2tSD1G5SFa469XLX4+r60d/JqFrgJ1yrM0hC3SVfx2/sfGjPfOWlkXJI
D4jqQscROJLjeFj8JIJDCzSGx9y9gqibxqYQ+FTVSuYJqB9yFTqle/dVKsJZ+1BoGi8W2kct6lhY
W3aniESB7egtX4KNxhdnD0iXEy9+09rlh7c1nGbTaEA7YjkwXJBypbTTA9UeUMIZUykf5H+MRwME
5dDR48lxkG8YZ2IlEGDgNxXQjp7fh30cdBVlZm7l/uA8AdBuudOLKbTpbjSpt7SdOtghQqTJOKAN
DAwzPGayUhr5+TIqNmkPErttnYOcxTgI1B7ZrYWAspKU6tnmRAdY1CAUvjE3P/FFbrTLUZ1u8b2p
d1vyAI5gPycqD4veZoKRLU/b3ir//5u+AfbOQGfq9AAeq5oh1oPFaosFwtjRZjSamA+QFpcOLy7p
CMUMYTQ9F9TK4m/4IG7Be4Gi13l+20BN+8NPZ6Ji5n4WCt27BLWFR57rdIEhlFzzoGQR1ppVwpQg
wTYt7NvqY9fGFdHfGmn94L9RF/+2oHKFJKqxr7qhPt4zUF90vxD02tm4v9+n9LhS9h/dy6Pad/T5
d5YK/hEveC/oQH6r8CT5s5DNOmbo8lrvqF24brxlqAyhPg55/cUjz9Y8wMkbU2rNVAryyQUHZf6g
EJdHrrEJca7jKa/AV+qVXHMyFeV46DeNj9CHSEdic5XCL7qXeSnx8T9v5Kg/zdGn+RPkT+8Fq/Vh
HbCoCA9R5hWaIZbzOTYtQlQi7jCikHCEqUpZefSakiYhXtT8li09O9RXNTZoFu/Ekb1acP3M1MUk
5mcDfDzHssKEl4DUpFRYGLtNjPmVI3aClM8fn8QwWUDcggpIhnOVfjBzD5k9ELERBdRUJYcjLwP+
whDaA1xMv0KOPvRFmu0sNNjwOJENG/FzjJLByZj29N2ROFbFXBLt7NzJw4N+m5qUg3RP4vAJgS4K
jGyf22rxTsmkb5NYP4pPwBtJndMzF9Kklr5zMvQv2vMjb6H1qFVqKSMWOc6DR6SlZ+AKjl9o5b11
fNFj6xL5iz0Fn6uWWR5XNgJrwTnepwTwo2vTc0JrAQS5VBcKJeJ/ZlknGFQRY6S7vCcUXXzwT6xF
2auZbPJAkctKgl8umDoFeq3r/OXbxlqEvymold3h3Uvcm7+qArd/hieLdmlqksXVKKOeBQZnhhUQ
xBcKM/YA4r/DZndaGPEOlPBEuV6dBqI/ibil8Nqym4T82KXU+gvm5nD7rMrylq7ZZYg4wfRoK/VX
LR0yg2VWkR8Q2sJKHBqSkPLALAEJW+uuuA3IqL4n9V6X4orHKgdrk2e2kpyraffct+EShyfPZqTx
8EJcw/aYdic8D0X63fJZrKgh4LLQfy3G+Uiow9kggctVavlJq20/l8hYVJiVn53/qywZRhezsdbO
WqlJc+PmyVOH6j7LN3nT+KZ8+P6MC1/XE1/mcYcBrxprs/xvdnIGNBxWovUzvkfpvCcdCZRo5hkU
dfg4A8pgoKalL37VVIm68uEb910QWQVh+5Dt8BMLYYEJnbiBaMUruxv0yvF1lzLLtmZh7teSQuum
R/ZX8UXfatgRTEn+cTMHLnpv6eePNL/Gyk3KuY6AW+bOph1fvEYxt/GR7i9NuS591PsXMn8sW9HC
Xebt9P5An+E4n6lGhbGfRURDLFzEmFZ31Ow4Ng6aBMkWRUH4YTGC5v+ef7LjhKM8cthRiKXkiH5C
uEGUFfFjGDnmpcXYUyNN1bsQr/VfXs1DMZu77LUPJrT/FIu+3HF01i4J/pdhYxK6/bIC7n19sK0V
HXve7WeA30IzhawUpXsMp/kNUrpMp0I2gsWVD0k2nJzc/TFyCZAaTYcwHjaoqQLX+t8bPIO3M4B7
CyP0x+zLKVhVbCBWSanRGi1243bcLvmxpTb92QV7cPuyM4AQfYS6SAiy7LS1O/VVaqE0OH3YSlas
g7fjFqgrh5yMSAzDiMpev+4w3ryxTCfTG77sqc6a+lDD91cLaVDdbnxtCQQFXE/eEH5TXfkb8vm7
mc0XG9Jt4RXjfjyC7xjLqiEHaWP/jn9CfKfXwobfJ/K45Al4NEbxQ3Ikcpt0KIvhRItQgELjdA2b
ADgovy1HXj08SLkNXdMokO+7z73HSIoaJLKbhgaUgKOwBez1U+7lAdc6I6nuXy6HR+gwpyDwruvE
FI2TTmluq+upLl8ZIKepgwKqAs9oluV3efhkXBmVWJxkSZnEorb9Y/l79QrHSMzYkSTuZUr4Wiut
9+PpVishYlwamI3x7Gtf6fVUZ9gWb4XTYxwmV75kd7kLtxerJ8xQu0RZe7Xb3jdfhRita5MMg2oP
q+DAS7OUz+Em+3JU/J4qVngoek+eNg3z3ypZ1GmaB78mkSKLNbOLuDTFF3uHloAzUv55ayRRFJcV
wMStiO9EUVUwO2fmMJVvTn9DP/u+oMLgS6d8NUtK3f5YbSRJRKNcIEXmNceuP1PvhQI5fT5s7m5u
g3zDHVXdhrEgNejVuoDVmIWNKlibcZxRqhVa74WhCGmfRK514lHnK2Ap92KF3obnV/LjPJvae1w9
NezDCDyu3A1258X7q+ewUJghzD3eC3226g/z5iVnKmgUnWK5aAtPZhQxlzBgzP7BT5d89xxC3lpk
EisMup969GHCMbcxUP5pUeEh3PRTym98zgGez8JOeV8dspoS047ZL46D3jHXq70+ToCFl5O1AMLY
6vhSbBkBmoqJVCbP7QXFu+HtKAKalA+on6oplMJ4v6aRhFTeXy/SCVS6GfPUya/K8bjvUwyaXObz
FiAelve+TCSfUSwFjN/otI6Qg3EbNAr1MqaH2aOSxkMYlm6yIuzDXMh+xWcf3v5qEmvZ34FpORgO
Cn8Jugb1sX9TlH/Zdtf8o0djj4p6jlpwqlEpg0Gp14qo6F3pcFWlIhyigsuXhPZ8pQWYBILSqZ1U
fvqe2keKe/9oJFXVSydjkNiZt4D9BcauKpgsbYC8qHRjDstoBVrAyXD3KTTGQd+ueTYrVBpm/7FA
kGjyhvEwGfdZfpovg/qlBQxuLOWg/fvbW4w+o7Fara5C06fiH3ZzxIjXgyvXXRjJDaJN3ZZx7MHB
tsa2rn0xD/S9Jd1lBvFwsufmLL+Ejo+nSNhIfugtFJAK6e6JQDWXQXUPrt2kSRLSY/zisCxJ26zh
rAG3inNU2+dhDBJN2WMDcQ/Ha703EkpneyvtTAxaEgFuBZBf3cWo5JvuFZSjJFmHdkMGkOp5stbs
i5MJ8qnywvQGtngrcpSb0ckb4qKZDUFfxsLTFJ3kYp2aX26EKPImgboHEMQuO4hyEwS2hOzc4pVh
CwomCsYwtUr4N76+yzMZE3/N+TEbQ73SaNfJTxLcKEU9xQo2on7Oc3zOb51yPTkBGWa72XcBtgrv
pdmQzvkkqtxuziHc++xBlG0VsjpI8WmadspHk2m+Wrvr8buDFDwISqUhghZcgek2Zy9BVNh0agbP
3CURDV5+7ANZjO7CdvsB5A71Ddsx6kiLMho2NBit58lpNAqNl5X+f+V6OO+LyJ8h22m9diey6iwJ
gOCe5BU0dUjUvzWAJuZ4HGeFWmpsXOY0t0uN158nPYG2x51KDZCDVeP6Hp6HZAU1tmYRxSMVvC79
Uge9Br6P/YwMRd1KW6HKgSUqsTOV7YTAOVSgVTfE/kkMU3KEwoGi+UhVDOgDTjyr3z/AvTIaLAaV
6QGRHypmxI8qIYToI7j++DcJJuKSd0Nb2qnTTfBQVAQtrkuMHhiSfaleBAXYuZzrCBc+GFZVWsBP
3t+M9A4/K+nxk2F/eOhAvzoa21Y0xuii5T4kiMavvHMbCxvdphiIuM2Skabr2PmfkR96VRTLQNy5
JOyfBN6i2nqRUE2qW/FxNRgcbR0YrZR31guU70iokxPrBMcyxRFaYrDAeyab+owB4q2lrvT1QVny
eCtrGbjeDXaFZkH/uDrMkk3uzDDP157Hwma8ZSbt1Ll4e6n0EDC4dywZ0brUj9Svwd63A9l8epES
kOnXeMANTzH8La0uyG07tkwfylTQv3sXggVVxya+DDin/f6L+YGmTwHIEAEprg43OvqpNw0XW4hK
Ygdd30VAddaFT95VUPVKMc+NgJxkRO/zJtGv+Y8Ec9dFDdwZaYB90p2be5mh56MCKoPi6o2AxmiR
Yr64Bd/x94CTqUCbCrpuJOHLaluyyr0T/vmrnxS7PlSQYZc5dRR5vD2ZT+dv9K/IlJkoK6M3xgJ2
CMNeEQoPXgxPB9LcIdQvMSIA2S770eLkpEeAT1jQUIapM/wmcIkLqmk0GSWvn/ILrsRzt2lCrMgY
vGnq43oeIprFrnpjILfLyEnjXgVrjtIIYyvHJZcuzPa0iIZiZU1QCtME781PGDFsZG83/TnMuoOa
5f3erEWhTeDp2OvoVnrNp2PIp0Ed9zUWjaa6zxCAQ+ehvf4ssl8KxYUsfIEPQw2vB6KOOWwVA2X4
ORUS/JhZtj/eSC8LGj0cJlQ/beyP6g94h3379MI2TzfWgG4/hf0e43MXIikuSY7nKqGklMAKRkfX
5hwZHgmF5viUdQhX7dvO/8/Aau72d+8LvnrCZTfxR3s5D+277CuOdqyXgxctjzKo4k7kV1nGGeTY
xu1InD7d4nrj2TNq45ZdWOlvR7PQTz5U5iQzQCZM2YxXYYwUIsVek2+LaKzVmMDi6XhgRwhQpuEI
8xeMxfk4RdVYeujdc++wPI5PLcyPXOEq9mn3hiNEoOukS5BJ6lpWdGskUpXXDc+z93RJLW/+mr5t
1rF/4b49Nsqo3VNy+K/x+2caiql4WRe6esJompDpGIIBwmznFfg6xiXl/Hda1LpF2chIoyqEdLT4
u6Xx3tO0otAPYUZ0PP4dbIRlaEkuJyQ/Q5kMLK040jhRliorBwztBglTFfsfBh3nuZsAewiokRpA
6Mt6Uw6aX0gmi3oUGugq0kGkeM9nQmBb3bThMWXEcWZd2FO7tfAT+gg7bcVXrd0p1/YU4b6ljtJz
tzMOKjshEMp4hNetJr6FEqLudDGTupGeGTc5R5aElQuErIGDMk469YUtR/6O3VQI9HTLaoWxNUSa
ktWKXRCB4xpjF57huN+FHT00FLCMGYB5NzeXtmfEd9PUUGcmgfFueW1IPQcX/kqmu+FUizxLyFJo
d1i5IZWaPevWU+q7fmjvxAhF0ZKj5v4N6vzjTPUnR9idOHfjvWlcdkKGwD8OAU6FLd8dNW7KLx9m
3+PCEoT4pNywur/hjvNEdR3iCMROeJy8rxIXdtBSEODV2YPIIgPvxoL1aDEbyREBsAWY2LG5t50X
62EIyhElEPjF7nKFYpV4er2mV+r6Ur/JP3fSzoHnq14fdZMMMy7/wcYiIJjqLlZstNHRxQMoC3DG
1DI1/2XQuj4TzfD/o9Eyf90kkxC63nPCjhC+s/qtOgMkcTKtLW/nkeDgeb0F4Xms3AxFqNxJY2Kv
uY7YG0md1F7zmpavl15n2i+FcfV0CCPYDzUB/92dELrCAP/PZieiX8xAYDELVSiKNKRGNIe+40Ed
B5zlg/hhSHfd1H+azCwICeB4GTJvEYGW6LKqICcVaF5n/v23D5dIbvBES957ea7zSb7M0LVIkv0J
mtfFFd1hdh6j9usnandW5weP1zOeetzzTqf/6gHc7T7V9Ki2ZgbKXHFD0mySOFLxe7y4aPQ4TXS4
xO5oc8sZQ3wPGSJhrBUe3xiwfso/WoZtEjqTD/sBmzoL3sPm3CywOyi5ck6HK9w1BxMNRRvxKbuI
DE4xEEoPgGUh4bzj+v+1+HIcq1DPf6TjFca3hn08X02KlsXCTI2pSIZP3aZacHpNydhvUxG7ZtvW
br0E3zp3jLG1hp2byTv7fd/K/EE9zIRB/YPj3mEO5487vux7i6EpyvKdIO0thgpWAh/+TU11Wz1R
0FPvbqzOo57HXd6ZdosLVrG8wCgQ84xm/jjtXW6GmcuseKT+ZaxBULV7Cj+uZFDCM2Mqoj8CQ9Jb
J2UINuPhgkIJQGU8B+Yk9rGaGJjRIVxI4dH67yNuloi2B5GEp8VLmrERFlZRB98vakcXDyC2ScoH
f8SQAwh6cfmyS3PArwyXiY1P6eB7koSSUsUw1h5/tpmdcYk/oFWt7uREF2fDHkhrY9z4ctoyBi+O
Ye2cX9u6FiecaS0LQszDu9C4g2ZwKcvy6XAidQ8jJvWe1lQxd9SgkTnXPlZtIe4Zvbd+SkxKGikk
U9D/7+bsIbkzGi8tDToyQiWwFsJaFFegD7WlVOpctoGtvEUMtuzO7svrebZOpqaQJAUHqlD0Vnwi
/7SkHpwSPZet9i7LdY0gpmuWti5zdHG1oRHISdH90uDhTKfsHYDY+TDjIUf86hasmy3mYdRhl3SY
3JKqIA4F5He9u/lknoK60DgGneluyBR7+4eWguxpeR9ztzKU8GyR5dT7jdj9fNwmx4K9mRGHTvG2
xlurbjufpy/0/wY4PnuohTKWjTYphaJm5DCEADlVG5g6rT+e/m7POlFOWamX/nLzEKfzkb3SjtE+
u2JiP7k7SAY+tE5AAebcumdfdQqWxfHrdrZp3lwW1vFPaVaCH3IR+icOvQlJy5mOVpnaoMSnRR/N
TD4Oun9aFLn2xZLsxlZxQJvr+TMadEfF7GHB9LDPRUQejM5t9H6Qi94V7DulGlBCvd9smxwb/eqS
SNMEo9rYDsEsWQtfwTZlviQJoqI6n/DwDnBkSZVIdsrSKbB1/cf/uPZlunfRajxIQMJP7KoU/sAb
hfpZ7ZBAmuOAYiONj4wtC/PPFAq6nty9mI2JrT5H3axVTUgyPL+WF+pSinzh0+9Pec2exchz0h8A
EJXk6wAJ7+9B8lLsRZZ+ze6LNRhh66epUZFzGz8aZHZOaEreER0qoDLj8CucKPE4orEtuN02hFZa
AWb1KvJ02IXn/Zhy11rGkvC1la3VsAVLEZJwOL2GbCMjyZsUHFeWCfvPkXN1HcslqwFvQbCcrvKr
lABXSTEXCIAAaz8/QjrBUfpNjjqO4qv+MiZzTFWe5SNYjiATq45S5ftaXf53cH+MsdA7XN8UfxnE
XGCjbmsu4g+kq5skgxOMw8B9CRjIDBDBTNrd8lhoZkvNmz0m0E6AfwxXZ11a5Yjp6VqUV5VKbsr1
2HbQRDmQGhm0D2de7p3W+eJmcqe3W4y4JcmA4BD5Hgdh2TlXNJgZ2x5zQPL72IcHZzIoy5b0yNzN
QDPoB1+u6NbU3NY/oCXTqb6zCNoFf7f+PgvqoX1JQGBnJrdVba5yRZQnxlsYIRY69BZ6KWFkbeHP
AVnyJaY3MZ7SNyWTeltvwmNT6OS5inSjjaXn854M6Be51iN8bP1RD4z3NPv8/566yWv3rec5vkel
drNJaD064nqSvYkAcSYKGJYLfl/yWrxOEmWdnT8doaL8+SB/MwjKltHp8HlpODWOlJNKCjqhHUI5
C2zJI9IWq98NGR7RqpCmRDCBwYM9mwoe1cX2+SxyR0sWo3HO0EHkYIpIYJY/CYmwiMLtgM5mUunX
aRGku/COSnK5YMdG/+QiW4D1TbisMb7KcnR944l9R+hEcCJCQvfuuyBCOJ03pC+o45kaMHSBfDmB
xLXYj0cSCPkffrZ2svFH3t90MBONSWqcVsll4/Mz4fqT5eS3qDtiWCuKu8+ao5eNvDCj5xjTzzvv
jGtUtC0ooWmfdqd8NbGuVkTGUrxj/cTbrs+OPT/KKWp8ErsAJO5fuIqo7dGOi6BrNF3JKf2iG+Dj
bpxjzGjvIpmkM4d26QXG1se9LtQYX9m2vpfMVosiwbgoHJBV1QYUI3UgK+dhOl/e6DjQ9jKqp86P
CJDXWaC9Wm+G412vTuZs+4AbGsq7PzODFSghcxVbqoKdLJMK4hw2bv0+6zwKqQ/g7cVCVMCpzpBW
3S/LOoqz+roiZMM1fH2kEIEeYJhoM6qRGGp1jukQFO28T54dQ0hvnZ4JtsIvHIROvd93HK94foPk
dMM+cHYBZclzWXUDHJ7Hb6Et9ho59Kpqc5z1MJh6imSbgoAyL4RyULo8nxvkjDshAkxS4BEmWFE+
vJAX9Y9+hTeQYmZSf6voQ60Jy1ZAg1LvPsAQanzol7FBjLst26Yr2oybgXzxakNx+Lyd6M2w5Pz1
Qlwa6UugfnpfgJ1ew521AysnVlUxsUtyOH1zcNf2DTFoKOnmxutvHJyqMnBBJlKVyJ7fqRWtC80s
Z0EV7dk0iMEfXeSTvCp4ogE8rSwWUkKVfDXxCzZcCJoW76HJ9uAgvuct9oqvm5mI3iXMROkDvYOl
GdbaN1Wf0xZDTk2FcusbluWQgAw7eTcyRZZs8UADc3glCTNtuaf+Ibj9Aqwqtxz0UeibJjW6oXQY
j0jBUsipjD2ESosL/4D9aCwguA0yVV0ETd1FdEbsPazkbpmsC0PTcA9bZLznB8gFkmMu89I8vd1X
karOhRrhhX/6QNyjY+FFszctsHEZXobdDAhfEinQmBGBUL35En9pZiBjzgdrLQxJZCNtQWwD3Ekh
a355KAsn6t3j7iJyMisusrABEjl+8MIxNxHnzmF/xWVl/DCGzTe6tgEpR90Pf31GKX3isfuZEi7E
OOSFVf4miurSGqkExCSQrT635kAGwuBuAv/gn55jphLQqvmQxJeoCPP5zQRzFNKHAJRNKUsFLNJB
rMTfCw5LDLMl/rX4ry1fjGhED2iLMyytQWkL5Oy8aDOmwSY5Ut8Y5iT/1LhMx/je/5FSlzyR7X9X
ist6pl0nV5+WlJttGkXrOUCJKqyENEGXrfSMO3UiJChJEAtGylheJ/Rgor2PYZ0UbGLlCMfOj026
nLiNdW+0Yp7R+0IA0P/XJmMMNFaNiUBaGH7zrZn463o7EqucnhXUB+VBVTeyhX7PFY1dYWTe0Nwx
oIlpmo+gt6X2pC60zZWzy83mI4MfmOmKMzJ+fhvjPZgeYX76QRqlz8AzODwkR5I5lSRP4JPsJdOL
BWOeBaGIEkiZBEiwWp34nT9EcjIGSM00rx5zYghna/aVyQANjieFl5+3hQiHRC5rPsYdAktELccQ
ob84FbHvR5tAeRKuJYODCQN08WK5uzIqY/MuYkAeFRF61SlakSbxfpzJ94vgwLuHB69quSyjFV4d
fTS96nsxQtdhLwFHNOoGZgesoP7D8V9w5wK8NVhlCGQEMW3pDNuC969A88tuebSSSYR6RfED9J92
qsGtXuZekaGkwTgtoNEEeg2IewzgeugOC7H1bh7IgnuS4+yg1pFGXskltjnN8KXcRTaVthcRI3DN
M4auSkKmEV7pJAsij+Wno7Ua4ZefmBORFoBd33Sx0D7YUfOGYUN7AmF9ErmShG2NLaUd0nb3cIB+
tzXezLPvIE4/2wZBMobSyAmrnoVn1nKh0216ZqLYM6LOA3xS3itXJslvWMM8V/HWYxufrc54NMkK
oVh/lCo1vS8mIoxvDkrJFBHGgw68qJBs3vY3Dq50QuVAtBSvLKHk93962s6Od7EQZBeIz3jVaLlO
LcCzgX1C+EDVyUSM0nruIs0kYdzLnnLyPa1k5CQx+oj1Q6+HBCFlz4oH5KqKa1BoOf5YFpydER3d
+/W24fQzGSvmIPc6ekMWRUm0g2+QLpEmoqv/kWX0NKEMVF67ih84CR/husnmvxKXYGTitz95G1F8
MkbVlQ26XhVYOPio6pTp9R8aJWQgaxOKzatLFijItEds4U46tTkRVlqZOOwcvhbuxg0hEdQKjJSl
WUhw0L/IOm3LiwBZlKhoWeiAJqDI+hSx0AlW5LaVsyTjj3xWSUoAmWFfH3rg69F9mZEpa4vCfWVi
i5+R3pOEyU0mgljm7rrEKDOoJoOCCUY6yYsFo1nR+1xK7EAowackPb9kU0Popt925rwtLSktfKZw
AMDfCIUO4IAmLOGqmyeO5VHV6AiJjV4t3R28Z9L6us8gGPU2VPQxuEyiFDRaFYwtoVhYukv7kgcj
7SQ16mRLZcypmZuKUqtMAxWkSOL0lmQirwEcOhjWQBEME3PG29M00Hto0mEJNoMTkWD9In7m4Wgb
aqReLXJByzWsFBc7NLXYJQqogrZ5R/lEj+YFP7xf0mkDNExo9yrBeatGZ936AfFKOajwS6R2AJvu
OymJZ9b2Lgu2m2L1k8Djxn22FPfPx2iDsfWvKaRpA0CSuXD/UJo6x69V+7HEBwgGazcCCL0V3MwT
96tGmuyQqLQmE5hDPGFFaiLT9yXljMGLMKJREFhSmkXIH5wg8wvckjbpoknUFfp6dG8wwTM4rEDm
HGPFopsirndUAtEesSIvHULAzGKESLdp8BjuxWXGUVuhdYWbNPuZIxiGJsB3fdp9Akuthdke9Dkk
2xapiBhiXKOSle4EO5mx6UFbP74is174wFSiR44S0woFGhyFyFdC7pJvqI6bsE+LL4MKbjN7srjT
5ZDye+DBa87hmTrNIezek6+jfRhbQyMe3dhh3KTKvfZuBNvV5F372EArx9eeaqlALjEaTumw5iKd
vJPyu7v7YB/TbE6NnqWSf7SHvzBImkf6oLli+qxwNXZ0GI86yxi0Y8f3LhDDHrUt7QmOUfjCbaDV
oMLCQVcEEOzs9APtLu8lpUpaUNoQPiNpb6NIC9mAh13xqJZrQlhJVL7vHDlgqa1apK6Os9Ljst/R
cTiVfrU1usGM6TXAd1YO4U0zfzhnt4vze510WsItpmjPgb+cIorco87lFVGsa5n1F15n1FxSecaA
2rDXBFfUp/JzuZOLcOz7YnTdyMXcD7d9uVC0Vod3J1GTAwY8Qok2zj2srLFyd+aAWOHLuLOoFsNT
TVnaG+JLa0nkHnm02F6o99V29lRqTzvGM+qAqrb+b/yi24CkY2/I0Ia6fHswmihUj6p+rJZKkl+E
M4M212+2Ew9e0vX3pBDrJi5mytDmKUBk21lSZe+97hhU2IxbyaZvd/bO/sIw8zToEe9JCxFM1lZg
2m4iNXhoK0dl7Xi/waeXrXWkGXcws8X00XjXpD7YqSMAPV+COqKNn2KTTAhfneBLy/2uwGT96NIr
9AagARPkhJRvwQbbw1uZy7pj/K2wuJTUb6G/JR7uvIocDNy1+2od6P9RKzUeFGqYap+bHl6dSBsb
/FTzC4Wtu6T+KJDiMjiov8C9UcynI6SjKfEaCo12npZeXzi7fYKAbgJdbGsFHPQVAjgTlkyNZft8
9YMiWYqTvkv+u29GjSqTe+RsO8ChxF6WIverG8BhRCGfWDfCo+Wf6e0NkkghtcJmye/QWJ5ivNTN
aDwWY8iqXexpaQ+8HU2N3YDZXX271XUr4F2diGYMW7JCXGVxRRxDf3O+1a3qY//CsX5kfRWe4x8U
CyRB3l6/kpvvKkuq3jfbAKZIG3k4Kfzdg4EaTcFyTBL6Eb7YlzRcaXB72CH82mxKFn1D0GHTRfTu
MqDSKyVeJnc/wvs96VBkwA9YCHntYu7Ryje5ToVNlktb+nO5/RAQBfn/U9ZZ140yvq8F4lP6zilk
IiRIiEUmfEJziFowSy+94rIh9LAL0ycxWVEZ39Faln1B/En1OqBb7KL5bUtPG51/NUmjSPg9PZA0
f/ffhxe5rijd55vyR+bIiu8iGr147FRrnRP9E9q1v5FYBdcNVrKCbG5wNz0KCSSVX3cRoUGiptMT
kwAqPeMEE9ovtNiLpC4uZd/VF4XXq9IE/85tVPoGA6sVXUGMcHp0FfQbOFo7yLYi+JRPbrlJTzoA
POikFV9FuoEUbJz9YhJnCxv3IcnWEesEdsTsDxI9AjcSYwJsz6lQQfoNOeZOppzknKpi+Mefw38D
H8sOCu0UIkT/K6lSXLfJheys3inKJ8P5j7CO8hw1VvtC9al7qhiUE89XCzANbbHhBvYQghItTKsi
cwqBi47WbJQ/BK7hZd2+dEZyuvcc/lit6bknNsbkKEYN2GS5MG2e11BDCSMhGVVzX+vUUBKOKjQK
yEpMxcwM1DovoCuenrdQC0IAwBloJ32xdso00pVAq4AAOzhDLaLmD9R1g7UFeMhUdWxvCul6ezVJ
+xp/dOdjKZ36KKkFb7iQ0Obk64mSGmL38dABfnkoJO27OKh3II872wBj8MZwRxrvUlHlLQt1BkzK
2E9fuANMmnW/iOUfABeCDxZwEmlULUaYsUv697e8ppDZfsm/FUwayfldjBFX5cAN2QbJNaXMO5Qh
vR2MnuO6W8aI3gMIOtd8O8ukP722q22nJsgBOesL8oX80Kl7rg07Q6joSAmyepnO8iPpQ8PWYE5/
nHJg4SwnAeg+PURNKI4JKpaR5Twi2zU4iQ1+vZLPQSewhMGH29bj9+6TfE+GHyqwhAUxKWhSSnHe
hXagNSXWYsWPhTvIwRK4htuXUFyVcZ7bKsxSMqzShbjjcq3GXmC5nHnRqL/mOBrSWArdfUktrCgv
6J0SkZI6X+oz5FpkhkF/nzGkq5gdgZScBQvvqGBiyTBO2XnSK7sjHW9Z2GlS9fH/Fq8Y5VvoJNu6
ew6KMME0Ft/bEsUKjkzQI+XGboLr9vUGHqMKQ5wYZWo48nkPaxSv+Vb+ThOEzTxkIr+MrkiKvbIp
A4qqC/wFiFcaKDPVvYi+dUOVQbGJhg98qUs4jtdHuHLzRm2ZY4wgRjdJpRb+B+ZXwms9H0HwLxF8
uSBhkyIpiJ3tw7BJstdx/6efwktFc/PqNIKSGoePGZp5CIqoeIEDiVcJ2mEkrHqBbTj2f6w3QCz7
nq3Oy0DjO0zlkPcHkAnoYkCIYk7C4ZGw3RnxrS010PYZHp9m5jUAqS3xBTA/KATS44kGteOmMxZX
3/d80bZYpvIpQZbL0QrvILqvAnmNAs9jmONZqrtLnAr4ivNn0zbBuduDaNyC0N09Iy0WsoYNTkXN
H6GDwoutHl64VA71KngUuD1wnPGmWGmrT0TwbCeWtyNP3EY6TqqGwBA5JyuSAXbpFtxlPnDZ9wCx
iFys4GoTxk64peYj1yGgoYQ5Rlancqba39E7C2tbBBnIZxu9z9Yi/zFQZ4eDyLCeE17+qq9xV0Fy
Kk/K0nD97MMO511TuvLKoDBXfuNZ1Za5OwqcAD2XNnXUooxRMfAYfxSQV0vonSfpCMCa+NinmdmH
LX2TySWqVkJ8Xfno9aWwDvs2shuEosRUlfccRXOE3vLJ5u4gQon/Uymh81cu4Kf4d6Orvhi7Y4Ey
mPYl9/NMW2rvpsIq0aVC9uDL9MZKNHlPsFn9Tb1JLFXCIDswOH0oBz2F2j5y9FTwBCZ6ZKInsTs+
n0YbNpJzmbH4FFeMjK5LLzur93B+gFZ8VGbCj70mOvWLir6P+26lujoMD+157fG28BaSwjPY1lrI
eS5bI76uRGyilgpB2lnlBOeIVaRZ4a3YrFHf6GkJjQo001/Ec0b3d7lukHnSX7LV4UYPevXOQMNB
3aM+PwSC5CWcB2AbPE9HZ/7SlgizJbPe/8suyrW7Of1k28Fxl3Ts3XoGbkZ7am5WtgKQ/cmtIAeR
t95f0wv98mzeuEWvaD2wdwZLbDU7id9aglpiuxv1HgHaty+fIkOEBthZup4lRT9F8fUVxyYD6LE3
ak/XsdDLckKwX0O/i3wLAaDUFzfKiIAz6jYItxkSX4vw9978CWunuWTvLfWwmJqUJhQhDjwnUdi+
6L8trrPPYkeluMaXiUIEeG0vGJKjBc2OU9Z9nm0hk0oFxYKEbh7UfeTUX2dkYsFFpOe+L2VUVowQ
lgQtNGTEUIT6rGF7orEyiyQPWuYUPfIv/LKtu2NWrtNx8Z+JqucqiBlwDmVNTQyfVL+qNCQxjFa0
X4IdPDe/PvV9L75+qJJkWqPyQuWOkRTHI25x4njcJfwz+HtN6lUGe4RVgJgvtZrHWEBq20b7wH5R
9l7rxNMK5eOBDpCu3tvX2sMpnyacgUj5TG1aHFzLBZ1DRxgAdT5ijP4S++o/Cig5WLxZTFt/4hdM
QcEP8UOPx8Wd8VTWQ1jE5cfeqwlcK7anPcHgfVuzsF3eOmdNUIQwx/vSUkOlg47jOLyVmirekfxd
vzg0I2/O4Mj+UZ89HjR3PAV284pdOXIyRfl5QRE709AFXhi0gJex888v/i+9s0zuEjBQ52PKcnX1
fS4SvGftTfz3jmq09y4rMY/ivLMph9ontpDnRomncg8MGRMSWNdtY6UWj2S2B6QC9TWqAYVtLiMC
tGWZHUmnw15dZDD1ej9tm+5A9GFVjQ7WgtL7P8egesSUF+PF3f88k6NhvCcY5zv9yUUWQ+IATGaC
9gseOmac0nTSpuwIa8mJgp2nAH9YdIFIM8ip3oyx1wX8/evQkwKmRm2r7NZ9NOghzs0s/treKTOD
NVlelaQuQjwqtLm2mB48cpOQqO21Ec3EL7FXJnwlxuxYYevKfgxKlxNrMZSPbICUl1c2g+hYmphT
yF9BqEIxwgzQbDPrQ1Pv6M6plA9kuwlLR3ToAryS/h8Dc+Rb1zWr8q5K2pTFgBPhd94/wnTNwCuE
+BVYHA+RmXaGyRVvSfU9f4Yz2cGzcy+zqC2voulmHh7XnKENoVjVNZUcBO4L9LRIL+8Y2sK1Icvb
XHa1mR1LR8aqm3MoRI4NuzZAYhHac10QoyxmdAMtfLUfLwb4dF2bl52/pyF3FS4HpjUjY0XIUNEt
EN91bvEExxUtjvt/VzB8BH6epTiWj9OvbvmQITqNV20Z7vqKipw3DuwQMDc29+pDBR8W63vV4qeB
HK7ZW8rM43+K850Iac+1TtZD9nJi7I2i1dV64yVeqvitPGO8lKqYtLQsYfzTZaKtVmMFsiqZ7Jnj
cigtxJWiMYmz9hmucyLLaU4R8uWsmkkANYONyEmEZYGvKEr83DWZv7w23nsy8GtCQGzzPtG6LQqP
BuALdIy2a6ymy7U38Yi1w/SmoNNe8tUKQmPppCnE2ORpRbQXTPbbSYzN0/ER31IXqbL9maYNXVzx
CqzZ6H+AthQGf/7gzg7Xl7E2E0lgmluq5DogZ2KceT3Zfepy8kfYCjWJ8ytuavHyHgp64C/vgNEk
cLrz+evgkGTo1KZbv+V9f4jcxkAfuimV32V6c3puKxhmIBW30q4J4/6kmFO/txIvhafKd5FohVKj
YXAhOZhKNrKqcCSgsvaPjsgV8hO3g6gw2Qcm4wMEvzdoXallSCJaQoRGaaEIix8MAzbuzbib/CU2
9WYNSbQsZN+KqacBye+mWqzTnlrxfZ83oSVXQXbK8buYizEUIixfl5zlONcLwdw0dt4nHo2/qJB0
rqy4Wxhs5Wigbua2ndgMqtVWhh9ervTc89KPS4UKUzEziC48/WEsGQHc/c/lL5wxUbfTDKuzuHM3
tGWh+lPQKcw2Mw5T/qf/r9raVilGGz2gfIy0mublczSDhsCob2CXNGJo/7pldqrhjRNNmXRAGKzD
5eTSI6cTlhalVDVW2E+LlcujVyERL+2RNDt5yQaZmxF2THsaJ4uh7L0IIQnatYu7XQBRvFdGVCtp
q3uYst0KnZ02g8ZJCzT3FPQaqLKTkDkCjR7OThFYzDXtmM/gz5Lx7n5vx99hSbKnFa5+ATjXaiFm
2oJ/B0bZkIDbhl3I0MJXlEPnHKjGqdcZeCSLgju4pyFUsMToW6YoGrUt1YSH5kwMfl0uTyH4JU1o
58OOZCuA3SPqiYKwUyFNe2cwGiGug0WL9aWw/oln1q9HmHfBlFV7zGnz3Zu485STzhlXTBfxKAz+
H3034is9tYcO9QU22gRzJepYFrzjCN7rtwpYrePg2p7GsUsE7FFo8nTfOvQbsWY5ArXyviwq5rP/
GckUHg0SPNng14rCrJ0zsanZIoFpzFJwIv9Azxv/rjAU2G5eQLjPfs4KsEVznyJvZ4B8oG8fsEMl
6hadOR5pi1551xjhthFC2Nt64Xq2CniuvAVraFjSPsc0kPuxY/hxWT6cuc1aJshBhimLnMaRSD1i
zvkohdcCGscBm3Op/9DRrNpm6NVRFrMmesHJT7xzb9oaNnYMIZhtcu086dkdH2neUpqH0ICVpQMC
d8tMo0FUUvZpaIk4NR0ITsTgUWx6Is5Bz2N3T+BONIpeLAwroqfxbqyKRtrrC83ouA1f+l90YYNB
W7YUqh3DqNqKY9wuw1AKmZ0SQngSAGwThRV8r49ALpvR322oTwkjjRZidF8dvZfGlQNQ+r3xwprm
qeMTQEkjX+1Exv4ynuKKdOHzknBWWUtWb/H+tywXZ/SMiZHlmZks8PnM1COCblfoOrw/ezklOmL5
9ZnIA8XVWyLvKRlErff5ayyNLE0Aa8jcYCrqWQfs0weIeGnTZ9gNFgnaPDHKQh77gu390/6txfrt
VkMWSvF5hM2voq2uyA1Z3Qyyv95P1fUxcQcVT/9myEPs/nQsdrKa4pvvL+Cn90aElcuHznYdWyYL
Zyc706iS66AJ/4G/+9dssGA4SPAfgrVrXRwyRQpImn0YoiyKsyOdarxEQj7NcpIXLjiKI3ZAiQBF
y0eChZvnPCgAeT0s42IhMmgN0bZtEqXi3TS/I1POlkGIwlBmmQO1eXeLLikOk3D/vZuG46x+4ypW
yNy/V6J0RzGN/aPOx3mg+F743VoHZ0hjaYSFbVZ6pZ0PO/IENTCSg6dbRtT+CrGxpNLnFpAt3w0d
UpjfJQTbbtk+MXnhmIVI4w6nVPqnU8FxPXu+39b8/IdMgniyUiNMTEjjHZYBpJTgw4POD4s0O8v/
vKtFGcvHaldcVV6ORHSioSdd+AL33FPWXspWHP/rFqu4+f5IPS8kaVdw243sDbOwJw5DaJsTcePt
gBH7yjHSSHnR6pzjK4jYSgTrPg5aiL4d3vp5MmF4UBEjumZ9ZxmmRvhH/UEqdaSnToYD3nwWSbNG
FAcF76RxznpT7MYiKvDlNJoYBXt1ad9FNS/6lBRazLWmsdY1bfWuA8bEx0o1U/c5RYi2nnnyp69m
5SR+eeLLYNaDtSuyjRUV0TpJy/GSqZevLhcYEhFxks4NISY/Iu3tEGIe4xalj92MIrrfWSvuIU98
7tiPbBJ/2Ic72UOtgFKV29ZlaHe/e2RNsbn6m0C1p5fAWVtu4Ya1++dh2FkXEIuzc/XSt2bUcYEo
WYDQ3lVYE+0U+m1kcS6W2XYCNz6o0UPp5fMA2vNS1x+kcHCUQ3z57J2uqzTiSTwPOFuDjt7B7owA
EbIAZY3jFJITTnvXrrckQ5AGN8t9MFf9TsLLJ70SGxegiQfhlEg29Qc47GEQ/6bfKNi2e4AdqAQ5
guXM/FTkKrYVKzT5PG4MTYrdyIOjGuvW4xsut3RG508Z/RbD4YAUmpIunDGmCabrRKxQ7sDLKr3K
1mIeN0a3+JCTjihcKx51LBc9GJd5UjZ4MPDfMObz0gfXqagP0/KnZQn+HOWBwbHHyfI5Tp9oGld3
LJNEd6iQPfk+1QYihkdTyWgFOgKwrRLD31QBn4Th03aszWsWJTH9K5zivYwfc6FVNEJPj9VjA7QO
0A/E19S22Qm4A1IXRMQV/X/WcV+S0Gcu6aKWuwMWoQHr9rj3GSkQpFviL8gNQuoBHQbD9GY9zTwB
S4RL93EBRxsLPNaKbdKEUSt5cgMalXDYzxP/x0VjOTY6+VFHieFGQsKCaBWnZRetvmS6vxCuC7kt
S9/IgiBo7uUpA468IDahubrSGfo2Avxu0SrkeHXORbAHGerjbMdK6l+QL0KtHEzwcrcCgcCFtzct
/z/fGiEKh5RY/xR04aq8r3IrMXEsJFiR16KzyuMWutGYn2t1OfhS17GD8WPIE5DRCDtX0OBj0u1b
w2fXcgG69ZlxEl2DT2CDQLP5+8bHWpeuzd8lqALSOwnCl/DfwoKfkFETquG3HdxaAHPohnbIF3Oa
/dOpvf5w+dBo39bEljoYqZzs5ImcWac62WtXM/h0C5EuGyCaZXf2SkJFZd1Us70IsglAyTcHYc5A
zY17HThMaUt6AE+XrK+TceWiq0H+FlUfC7BAzxnb0eB7DRWJ3SPLun9pHno+/hChbrXMVoB3K/8I
9JOwPLzHL4cj6fk9CRFIJqZupEygJhZUzghd9jNw4wp/zBnFRjDVu/vx2Uj0j+x63pHFec8ur4nb
B9EVACD+uKgZ1VlXhFtrw02ts71Ok6Opnbzla3cIy73pJandFzutsoh+bEJiOCZQ921l0BTIK7X9
KEDtFYmhuMidFtFs153do5CwtBuAi/bZvXw4L8kWZwlmmCtB9DL5ne5jl1jKYXQlEfl3aIiFNSC5
BUxiNIBg0TOhV01SsVVP9YFx8z7h5mGxtsiE89jT99BfuKBQ+4tn0lowIv5s93kkFi+LYDynoVa2
7WEfYdW9EoRLdgbLPzAxgnQjxOL7EDdD3pApdXfQgBdTrN+Se80MO13f7KNb5sgd24OqI+fZeLeO
pjLk7yJ1A3iMHQIowJqeovX4X4Be1un8dx6i/kviTLld5sti8TJ3e7KfIi+C35MsWMtvJvEXcjS9
E7TpoBkIqyzKlckqwMgXBEFffoPfVpHid+0I6b/wxxhVttGL5Dvf4PF0Fdm4VMpEHHBad9RFOrEQ
lJkWfEcpLVc471H4zJQJQ0Y/21wRXFZ8WjXQO+l9h0/fBRvajSeOA0P4YAKiXIsEzEYY1QCzc5E4
W09jSdJ1qNBFriFcEFUcoh64uvqyXMlEL4Hf/DLO+3cRE4HyFQSH9ILHNDwmyYyVSyBwuD1qbzN9
3ZF4+VmN/quVuerkiYYc4oM/Yyu1V1+ZHrfHl8yKfeRAPnjUeuEg+TvcVLvCsovmx+yaX5VO+ONh
RW/BjQ4IMoADOsH77Q5Ar1Te9vi5BtGO5jBJtnCjrST0WYtgAc2jP1DSviKozIAAT0eqZ35EmQZE
B36Um6HY5+YlOc+0hFBAZYg0wVVdZsQIudUApDUTzK76LpNI4+kU8KiGYB9OkO58vQfX5r6cUBBI
MI74OtNTpIVhcndVMT2oy6KgK5DqeKEeBJwAxnpWAAtLzdxjkX3ijiR9j7xzxeSv8E+LV+VIjhN6
ULaQXTkSTdWfNIL6w7hZEe8KQ09k7KT6EhR9zVJ9VqzxqouLdZeplU3BcxsPwW9YGxzbVlP6wrkX
QXKVpbrWtkDcYMD6MwJ6cIS+XEnpusp/3X2E/z/0HSx70+6SpVnhbBqS5xZw1Bs3eWOSB9W61USm
R5DdjKVte2Fylc8x5FTHzuysKMSLTmKyUgYgWEoE05BaX8cX/Ku+6KlV/txeCJKUnMcE5EEJUSQX
jd1IRbeRGqULe+00UcHgCPpL/gy5km6HNBDsyAJBFb5AsF8JDElx+X/8XoI5O4Vr1fOFFfXmol07
6S1/6gQy4IyavSRudIOz9lYp4HdrM8e0lVqVkPuAMm8kkoOYAlzwgFMq/WdR1MzjPIUvhbiyCxxL
j/PiCeoIZTrBv6Fl5DlGmhSro+ptkyfCNGiDNvxB8dZ/CPcWoh/3yfN4BhPHE1jfJJY18mp3DE+P
TjBUWfFIjn8OXBPWcn4ctz9SamVXrL5Rs8uVyK91zZRBqPOgGW4F7huxxRD5vyixiMagPvQ/cwIK
JjmzLgW0OuX8dE0fL6wpO/qj6NUIbeo5vzRm5Lg4mz5qWA9NLFTraGFTWvojZg+jIw6fAMiNJuad
U4T2u4Nk6cs3pB1wWytYob2H4cXN1G8oEgztKrM6YF/t5gcf7PUWtML0YVKgUH/v7rdvp09wLsSM
tNps6azzviLp9PHtv7mlF+kfp4TdmM/ZZYrUmYc1cqtqMa2iMWVTUzx2LjPW/U2soZDMwOiRItf5
+TYxggF9rRRbZCqAE49MlSl5BRF0H79/wNw+Oo3J9RQPd2gYhUyE6MRKtuQK0zpSIeef3t1axMZ9
D+yP+1DB1FBVvkH6MvMR8/FOXa5M+H9TbBzyfyM5nmh3OK2S587PrscnoUBzDifps+K0D4qyofcU
FdxRFqyQiMU33suwAOY0gvtSla5GUn31yE4BkxqTqou5SSt3x062aaWX+dVmYFW4e7nxBHuiIYpt
gCueYX//9VBir4Y4x/5L2f+pXEWaMN9JZ0TfFR0qaoC0xNzE0o+Y1ZM96+omMTxvtAhuCvTquSp1
lMkKq4napJdyxLIou65rOw9H14UqnPz0kL8h4J1TB5vhjb7lFpwXRIOYDmpM9w3cQf1ffh1BLk4H
XelyrjQT4pN6bjQmeUrtL2+ANZWNmAe1VgINjTb/exfCWB0bJic4EUMBNXTKP/xpYyk2G05NNCiN
guVQqskDTHSlmwxM6k18ffXiGCzB+WycpoPocnz2V223TBaGm4TWQpl3ynSnzNOVZqm1aj808Fsd
+i49HakVhOmDsf8d4TzBiZ851/clapMPXJAMo2gE7L2DorjJLQ0lWC9Qri5SngtxFaCeu5WFlelg
jXW2lF3lNVeD5U4SLYIlzqygUjM8BZqLiW4UIOR/1ltXUwDN+khVDM8ZPTU79xLpoQBihiBfCOEX
d1q2rliwDT+pzkLrvpC2rbXCivH3zOVkVYP4/5z1y87uMWrDy6O0qXijf9iK50cQ6y6Qzl6aaHKo
Lbv9w4q6F4+MhEfmmFG+WcAwEHaHNj8j1+WHV9JDwt/nkVgaLlXYT9WzaZQ5nnvTcy5jqfboZuaK
e6TkBhH72I9rtSJifJs622IwATAN8LLYWcxhqTEPzw1ZtearhbLRUn3fkT9EqqTqejMMy8sQx/E9
UeRXyoUg4IcE1vcn0k2dFQUSqddcAMKI9SbpDcYINTZ7f5Nj5FbQ270AmP+loYQcCFN1qVMj3j7t
JGubVQOXx4HpiG256K5CbYWCbqQgc12ko7mRhCpFEUuAEDsOk5Kj6YKdj9mgWa2q6V9anq2y/E3b
R+PUH82/bJmEQLa04bpycZ0Xhbo4rWAEVU741KVl+1/RExHs1aSC4t/QZ3emyT7rHASSSBzvZnsh
Np7dd88PJWzMGwgNrNm1uGpCLu3ah6vJtcLbHoAaJ4xpWT+8mSqCQXp00ZO0xdnclp18JFj3nPZ6
g3lECXaFnJp0wFWsBKuaqcXFNvuvgS3NvQ7wzKL7B4hlQwZi8Jl8y6upPyUM168v6zhe91PbbgoC
rQKcG09Z3pmSl9pnVnZmFta0NttZ2qdA5ViR5pIpnkHfWBZSIWGeETjkr1h5VM1kTR3q29pPBPyh
BKw1jz55yxa2nSE8mIdSYAHJ/6ZizcUcvVbJQcjboDZOZS072eGGHPeCF0UQ++REJTx3rru/+dNS
Am5rtv54gsHhLm+CZY/nB5HrXPEK3EUS2PSCIQB565PBZviWFMUUknUcXme1+qcQDQbME7DIMjFN
mJOxm1n0sEPrrzrvOT9RUUjJ9683TMBAKvIFXwuiJ1mmD/eXqDd7rv7CmY26W6bVyRn9uQn9/kfM
Xj/b5nuJnGEnkTYwYIA+8cyA7QgoS09kp6PepRdigIdxmOV6tU2aJFEMwAwq4oA714iw2LOa0NGP
/sl8sgDtyf3UXupH+i2ipm7vZ2n+YrGlEYVMGLIxVX+KEWFLG7FtczWFvrPkzR+BzkrPKUiSCKgg
FAKA06Wz7ipdfL4btjogT1J+y5kpA/Uq4oBICLPF3T4DEOz9yI5r++c9Nn+/UZS/oyiQBLfMP7fy
WDEzofZH7YIXC5V5Taqm0KFwyrhouz2PheFRP+tKM4a9yDzNP1b60yQVwkC2MpBGa0xqBbqXheic
OQTDrEcNhm2QyD63IpL4CtkwX2MXJYXqusapo0Yvdfbf25N1IdphXQK0m3d7EconcyI5eTsu22mH
EjhkK8LrZ3fogQ3/R3lEVIF9L7qobEjMSduqIihlKzP3nXIuUJrxRvXVUio5uGyfdnTDiKl+kuFD
zZZazsWgWqNes4KUAr4z1/VW5eP2K+ZYPZqwQwRxgZlxkFPkItcfpdsnPPJMkh/U/zmRqy6j0kRR
by2YOPPs4FQwA8NzzeupTnHLyWAkrsltNv5bKVqiuZgiyz7dPQ1zOxx99whZuEBS25Q64Ghu8dbY
ooXkFyobeDbPdCvyoCko+d7y37YG2NUImKOeWogqA4XZZY4Zq9mdsu/wWuzbZ8/83IApnj+zT0dc
qfkuLdpSnyRJm2McWMcukaqGvWx+X7VHFQ0ceXeiXb75TxHtsgMzJpIo/iN5x0ivdkBLEKdzqLfL
Ton89edBASABLyHPG/LuruFPGY01OHZJ8fjQ2iGUJO1JLxU9flVUKeHLKba75T3rq8T5yZYDUlCR
C1BgRuW096+OhIt0chBBXwk0AUxPfme4iP4cvbutiaD9jkgM+voGomatpWiwzbr3b8jHQlS0uISD
ht2iN2Kt/TKbY4tkNJdQPIyRBZc4NSLJ0JR/cjXgXgJQYMyBE0OYNCpcS2agfxtUy3bun241Se1T
9icDdQ4Xb1tDuIZH5vaZjZ1TiHTE+1y+VDHGbOH2PEWFaeqNOaJXSuN5f0lCo3yMGlnpXNym5EmS
35ZrJzFG7M7uQeD56K7QvLCBKDFMSd6b2NCGyssAJ/FHfL0QtOIiQFzAcXdT1W0RvuIadgO/POlV
6EgVGZczaByKbT2CD/+U7rKazpfgO9Mguot8TcNcZcCeUVKyyNlxhRX01vrkN9swXsGzQX1+CD7h
d2wyYtLF0hvHvvQcX5seUbeNbMGWFHVLKD8sAG1MMh/U8SvDnWIbvqKZjCLude+Oj8TYRoaLU3sH
rT8ITs5Tc8wY2HvanLVunB6o7uZX/5ijVIWg6snK31k4j7v5JkINfvMb0D9M05SB0GW1Opm0l2cI
Pzkg/oDcSpLPBtkwCWwERvzZBpEOEh38he2CQYG4XpGt3j9lF8hwTUi+qZtQdyDwLrNfts5hOSC3
aCJs6rfnm+A4y6sdI/dvsOLvTX0hIlnlYnPxairipXDUc/uT/fhBKFGrrLBDt1GupO0F3FiDBA8e
oeDw/rhFi+roCjS0Uyni8yhXOMqgeth0e0U9EQnAVnL8/CrUBcpK2jJEUYeoTyh3Pb4bJYeaS/6H
Wqe0m3VeEUjXuKOnMSsdAzh/dEHiNpvYj1RAeqYoX2+6CSgkzfw8tzuNm2LuCgb/cnVfDg/W02bC
5SvU8M8geiCVE3z7mH3I/t3yITx9sGCbb49QWu3GlRB9yu9HPAzhP2sKkJga/uH8RJl+6TOYN3Gv
egpm2KDiR7nm1MXj6Da+i2g7rwfHg+Yud45ojJ/RjfpF0hx3hdPnQ04WuLvCe+d7F2iY1H2rLmk+
St4uVRDH/Fq6MRnZs7OdJuI69uvWdDpicnGecYQI7tiD++k9TBtbFNyO9bE1kUaGixTBsz+cTzjf
BumqX07wTw5EuzWW3UdXKAkJ9y6hqkuBQmN05TMY0X+by5cEsq3+nQY9xnHcLs23qad8mnzAdsaP
8Ayer/NMMO0NL93AUc7+hVBE+ONeLnD+1opnsYyRMXEtmamU+agn8r+/Xky1RbFpI4aiQYJDeugP
NbGVz2VTI4GU5932wr9zVNQjTPx5AMDqAVH2CtYhx9iGHkFkiEr7lRFOnLyQWK0cIGabClqwUHOA
aLfBTWkUdJZHfg9lJPJ+4Xtn1nrpTjtzb35i/gJqjPTViRYJqDfVBL4N3TbkFsH3frTWw9UXuFzw
te7dKxijjIC667IZ4gBXcabnZKrAS/WVoLtiY+Gbv50CvA3C3wryCkRl8jtFLGV0ei8X00sryj4e
W6uj6HMhbHFfLhAa1r26UlUmNATT/GlD6fIAhJel3syHwcK14PxiuiaEf/qSmiaLwdW1zl3X7Crm
nOpLWdNmgB/QEXalrdjqe7z91UG3ei2MCHypKZfLGhZQ+Ppjv9Q4cq7kKr+qmxW3NoYKNaB8ml86
q4OlxXs/gTSpUZz76fVJIcyk+k/HJoSU6Hxhrqcd3AZhpEtmBEi4vWn5sH6xSw5vFvPwY6KlQQ/h
Uz5vt3jhz8qH7s3PraRAq+G0McLY7Q9kp7XtmLCZME/Bmmh+Y/ECWHC6By8k2qJytobxtZyVOCOA
0Uhy2+S7Zfz75BNUVa6PxmlSxwRVmfes61dMXVUj2Ob4v3vjVOlvq4duVAIn1Kn0wsGtzF2w5Oz3
wmLfpVKKz45wSQPlfBCFBMk0UkgPaVF6rd8bE0TjYz5+s3n/KZpfqxO55iQat4DWJZlfJK4zMXBX
p0t49oBk+9+fOsV+IyfJfDET+KiV911mrQHPp6IuNK5QYD26NulNNNiRoxxdSiMqy2xeyO681DK3
IEqRl7dISWeaadvT2/tJ8fgpgFmc3M3Qz7mXyuKgNGGqEWup1xtdBMcAPjABZvmCBpsJbLQQ5o36
Hib/xoTJmA2YMsZCPU/R/g8AThV7q5exd0CZxDsp4lvjB0JmjPnYh6HQajZHqDf+Ue5Xl612NqR8
EbMlQjQQNKieRGehZzhbLxMNWVgz933xnYCbccAb07o9mX657j32Qua6tlXlDZIOA6b5JzAmVuWP
t3ZwBxZl5ImKnumFMsqhl8p4DzgGjLC8UkuHwYKq0vQ2Xup+E0BmADkebOIiNhptv/PC6zcxa4J/
LxFI+WAA6Vx4hnLIadmT2SY686wcP73FLyPnNRPVhYrA3No7tAdvv8VUKagd8YD8MFEFr0fRmHkl
7lTRugdI36MBDZDpMM/t/NTnC66/La21bP3NeFJTL0HwgyN5tbvMkOdhynIMEXa6PGtvWfkzw669
AWDGEIZ6BLepDPT+tofJljMQfdPzDl1WmZfhdOScZaVslPYRHpQgmv6lx2M+sf/wJSfT7zEX6fno
QjIIeppbcjhI5ZuD8z6lIpLQmIfBXdYzGkUtSgDY5N1LZXQDchoFF/0Ytgp1GwTXL4ts0u/tS/OL
NI40t8nyet6XIjd6ZaDqIOZc28DD09K7koQYPuHKxpbVTPLQFMDN3ArSXFmlLXe2F6DGIE+8Ly1m
LO9zdM/x4QjyFTYABRJ1twzBx6POQVYQIfGDKuUv895AYilWQkIZ1I26f/00CxuJJcICB1D4bu34
8uxMUzhEYlcIG/8XLLfkiQrr1I3ohYhlILcMPiWa9mKUkESzi2C6trwPP+UttdC1gpv6rRD7Vjhx
xAUVYQ8tbCTOZ2+nYr0QV7KHZ5rCm/SWDkcnO/uvrLvLDiqL+Gz0k6qIjxZgWasTgJKoWqtAiDPz
0Nl0p/XDvQopCCmfjj6V4eFHx+umvgSgyoBE+UdRuV3LwMa1AH/SFLce1OkhEy7b5QzZrv0PpPlf
i2Dx9CREVXz3hwT9yONtJv7QcupLnUb87OFVdksdXrqAM4zsXcz+3hQNGX5syGUSHlsjX9EDFjTa
l057OyBw/2xW9tc5ACJV1NX2hG9Ty+wGFKlsM1aZemrxOQZAmf85brUEp1PuoELbLJgkUjGhTSjG
mcC+IvuwzUjrMcYnIYqSJQeuPDxzS5I8vGvdgdAXIAjUw6S3HMa3gtvgOgjYLHnNXwufaj1AGcBh
xuVP6Wl7pL4ZE//duD3vNnxjYup8/+WddvY1+JE8mK3wEax+L0tC9435vbcaTfbxXeLePquXJvkf
QqfrgJYZlxamzprtVib1irqjN2cJQ6XLVJGea/JmgNa68RNFxj+UXBfzXX705sVHvesKFuNitxOF
7FqXIGch7amqIRR599b+7vxnJ77Ij5+QJaSueChtxWKlAAqwffws7TBY1FIGWE4A4Dh7mN0trZz+
wNSJr5CCMaJZnPTa+7uH6p0mrof2cmc4U8SlcMtkD+b8V6lCdRQjddOVpxziIyD7kOo/czLxj+lm
r8cpyS6EDMG23iQ4Wh4CYeI3S7TM+hWen0/ncsKMtQP3FLnzpvLYj9vHLj+tLCkhx2jRYU2pLhDa
yIjBd2lWTrb8rGXWOcwKHwfmcaLTSdGkd4n9ogNjVxWcAvCXzTn4J1WcxufZl6ANAJ8YgOghE3ih
lGPUB+1rFebC848WJPfVoah77PlZ3VBwIJGBzgFlF1kdyeDrd+Rsiy3tiIm4rPkdIilUXN9TC7So
58lZrr26VWfl0As8oqSbp0xS6aTTe5Wko3c2Kd8sJIIvTE2EceP5M1G8bhHxphuTfcidPJFcQ5vb
mqbSQp+XgOHDA497iCiSCPSrDSW6BHZy/UKCravYGLylNc87cczhdqCFrPSsg7VvJFdb9Z+Q/1rK
hT7tzZ9FGQmE08mSznOFDP+d9MHubQdHfPudCQowUEES2GYzi6h9UeRQlB6JG/fElulaykYqth2B
Qs6Ez23P+D7ZKTHUhe2hPbuq5mpj9xRnK27IfPx+/XsLtJy8WgMIggmw+pSupB5LCoGrklbagBAe
UGFFqk3kJSsDnuF9UiyGDQVB4KeUqTYPJxJ7bVXE2acfEg143vIudyAjy+WQZHuT8zQksbdz0x0R
j6vYx6kQQ9axrEYtpOfP3wLZnQgnAab5qu4fpTrpDjVc0bJLKn8cmYS/hr85fhfU4meb3rhfJvcC
UgLMpcW5bovxLsApYT9K+wbha9hl6ri3JGKq+YdvQBcgdgjjYW5l/ih7XyUPYR/wZzynUz2L0RFY
NtBKicL09bdtAclhrT8DeLXxGokMyHrBeKWtfla4KB7n7LdIhisZbGvpaOPQ1P3qVumq/YKJ0nTi
0WPHVJVffnNxHodHg/LUpVMi0Cqvxau6quXhccnvfJKjZqPlYbePiha+LTU5DRqq39MEnnYdY4if
/D2YY4e17WygD6Txv5fAPEuHU70t4H3iHjYeb/bNPr4P1s0Hs2OLGgXRW1Z8IfGCG9tIIBYgEVqp
ew4seLJ0nkdXsgpSAkMaurt5HAdmuMkOw8S3zbWOvCv4j9BGtM+jrawJBtr0WaCJJiaAt4507ZAG
L+w9sjIpX66tcZLxx5Kiz5jUPVyvPOwQx1uh8EYvdpkiEtY6drnpo1fBzD051y9UHbx1oQsQgNBj
PTdL+q3eDJpomFbMlhF8mEoZd5dIqSOGwqoV/kNVcYEQFvX5eaKod1Jij6+iHSERLAaxF5SIpKi/
TtxE3ylhYo63eDO/dnnoo1uytVgY1/FHG53qJOWXR7Q0rmwByZ0w5+tRsTcBhG3NBYxOMtFdP3hS
mKeZOtaca2Smx9v4VergcTruFm7Nhpph+xUTYnGm98IktXLTX21VSgLxcDErc5a5U3ByTn4UhAs0
i0wbcGhviBZ2T4blQZagIzKMHa4ZuAMiFYsM2IwCgghXCIU3/7OC4/m2Qg3FBHeggfas1i17cXzv
qXM/+ed0Rnx8tkqsJh/HXPI+gCXsE1Ae6XFOhfgQ+WnkV2uQn2xMgS1i4WOVFrTscTiV6RO2XwQg
tdrUQ7z9gmzBiYPiw1cfK3X8kzXPO0gtkfDWG7x3lmC85HtLEmTYyy2AJkfPLqOK1NxZ9sZI114n
WJZGVLIUjtvIp7mY1dZIBKdl65ubZxXPWAorUY3QVh8wrYk77JQSx5C2h1mSRPavfL/khCKJKAfx
E6bAHleE+aNROf0r/JlB3BB/xf7Oad32x1sFFWgOZLg83XHOOlHOnWf3Mw8M0JuW5XjQIbEVv/vW
OgNQQ1spr2UGKjzVHbCZhqO9HSOPU7Aob7REnbGbcQcdvLikb0XZYnEqPrf/mGk4PfWNjAvXxbIh
UkgYidVd+GHJSvQBxn7BrgO0aKFI9YmPHH6jImn/l+eLZV4KU7VRp4xdKCWQ0xMUXiZ38STev8rH
CHfXGHpEs4hrdKO4mlCBVgSqFZMuZ4jPsgzGkztfWJ1B32OKqYq5lh5BsSaWLL8zvPMpjjp1jUV4
KRaAXgkohxgZdfq+ki663uLygBub6ON4z3c9H71hB4jGSYg1joP/UyrkvEYgkmEoO0sSuwWqlnHH
TL20UiVIeLAWplIR7o9hVqK/0dQoMdqR0dzgaBFfKhlJj5MEqA3gAy1lO1QRAAlA3knmNsmGmblh
aF76g7tNJDGGBZ6Ai/xlPV9jG3shETDJytfflNLZqhzGoT5CCdL0hkeMurymbhFpEEd9Q2nbyY9g
IHAU0nTrvsb2Ibe38R7tfg23rcdo1P1czOYQinxfDMta1QoXnzdkyLRvvxPz7pr3EpAJNdfmvB+8
FU1rOgPmFR7WjGYKuWCSdAoEemgTIvsCliXO+Ru+eZTmWZKpVt4Bts68FfGzCxTIHpQ6k0gLqRQB
GkmrZpaTx3vBlvviVXPsIedfEr/RQ/qF6tL1uXZAmVZ6vmPGQpMTARRi8P1Z9l8XXgQEjAo7jiC1
qvIXcoHizXRrGBW9OoyaiX+t9kuxL2ua78LAb7I+2k25lcbdiMgZ09BjDg1Y2CzO7K6LuXelbtfu
tBk/rvA19YNAvrWF4kBRYZUyjPqfZ5CDFi+nvPwPUBcf4yI5SSrOBZnNk+7JW5bNHinfqbrzYn+U
FEz0mclMwzS1sT2ZHBL+jho8wkY0L0Tw+ftJhLwsYB/QE0F8Kwpgj/xg9VFgd98oYxInzO+IgJXp
9dNX7Lzigt7S+UsLmklkHtlEsvNPuGtqVeOqdwEuBu32AhOYe3fbpdOP2KlO9fCKxJbJy9pOlbxC
NvBSOAwEb2ktA6r5ygV/O3YMJb60rj9xKxwrOgIvF9Vont2VMc22xwNElxq7YIWyuHG4QnSW5+84
iJz5J+TCq8X6c/yAlEPAeYl7QSLu9NcKnhtv+T1rVmzo9zoGwICiDGP6IkahHT9QoJM3AEDigRw0
4xFAx5M9JlzEjx6emI6ib6bB5CK8wz7dbyPqmSjAU6mpDjperPzQ0qlaeVGtrGXZ/GiTWYN8Vhpz
LiizAOCAgXGQB6k5tQQp89met6PnQ44G6vEbHOOhbTMv7B/ZTDjs0iMlQSNS5Z8wBV/lDp7H86B/
ZPoVt7Z0EtooqUXXNYwTIxjjxHEe6rMQF6+TYYPmDaJ7P9DSMK8o3uCdCvimJsQS7PdSJ/lJTVqA
RKTAXpHTHchlaxWtN1CXGCsg3UvglNmryzHMSAsws6ozpl3GIeD2lu9elViPdu78gpgnNrtkMxBJ
rTsq699zqu9YFGvvuBB1sKnwuHxhTwAWD4XtwU6x+j5tjaMeQve9LcGBedIhQhVwsbW7io6/d/UB
aoCrAiek+M2DCTJB7XP+cO6VUFbuN7sgiAWOtf4Evflv+JFp96UiOfbhtjjAlhDavFhDf/GngFUe
hdrG7QNDlNFkD90ZDcM7cEaLmha9+fNyAI/AXm25MmSi5+lUzPa/00Z+6lomMDyOAr0z8c1ad0sv
mvi0N2dCjPbbGfdlsQH2i++EROrsFlvIKrPMeIlIp3TLPX4s7ZmACl8cU5OMP/kWRs9Bj1lWy+tJ
FbiR6w4YRUylHVQEbjoVDIov+p2Ea0tdkPOaLTv+gInbzS8Eh9T96QUHjQECE/r9HfNtrBxeRW//
4oujX7XGPQ5jO/vQnpijZ8gbHScRhQ3WOPyL0eiBDG/7wnJmM0obQqeemKZIXsRh99NFBCRLHlQd
V+O1oal5GYKR/1bikuAMhQfmKZdGZw5x2Yk9jkipd93PyonREuqTped4AbJVO3tfDvKLkRK03MDE
1bilIdMBMGELO/5FN7xPUaoNT3DRL9q0lcjkzFYBS/26vftuc1sW5kkypOG/Q7ah12OvEKtiANId
pTmF6vVm2/IQI2iwPfxCAHMDVoAP3wBf/Uhp4qyEYs78CXcP3jBTU9wsw56vo2VEZPmIx9rYGHjd
sDi680rGdZ+MHw9oM/zJXmqSH8a10RmzaGVGjw3D1+6aI/UgRItn+H/0v9lNpvpBAvE3oIXbGGkF
bHspMcUhQWl6GyeJfVjpdDFfOmL6ed773rFxE5vatDa7uRkVoySlFDjYaNALCnGuJjxXLjdBriTs
RPra5AzmqxbU2qj2I27KxvjV+WVEHq4jym1foMw+oLh24P8jrSaPJ3hzLhPNZ7N8WEMe7guOSQ9y
6iYTpAxqaJxOJZdW+lmDs/4n7Awv5WTlhE97Gne0mlNgAT+ZUeB9s6Jqd5Wt+hXHJYdFI4xGCmam
F8aPsMopimOZ9hRFmMgoQhRKuAwleGDC989adZvhOpoCm/whXjGZ/5HZn9aeFG3EYHOKqdBepShh
RL0lQDwLJ4XVLVBOv/pSodZvMqh45AnmoeyaJBF/7NdBiYGm70j2hQRp6pIGaXtzPv0pG3PkFYd8
WC53uqi0yCKVaAiE7i8w3QarQVl4I0KWeh6qIGHX5nOm8KZZB4fAirKPBRdSGgOCO1dvXxQfMxaz
aLTt1M2pxv1NKo62tn3qZ29fXCYdRtZilZhwQGOM5dJy7OnpZJf5kiLHoXBcHw1ICZt0E8hEtWDl
dEAk8Vob6i26oFuu6ahFXuJomILhV7/gpCkp5A2zeJXm4zDYcVeogNRasBmpqa/spk0c02Hxu9v2
j+g08IFcs/vcYzpU9WTjqokuXfP7YqurH4sSYdF6dCWkKwv3JG/tS3Gmjb+H+hTD5SjBDipGSxok
U7OOkoQdaD2Hgkd0oMgVudiKG2Gu8gJ6AJw1vGYU3+W2O16KqX5pIxU5NxgKJehWSAykXaKpSP+I
CUP5nwgFtbeEqWYd3HZV05HNvGzGd3Q6BnpYe2NPa+tw/vf0B+0PjMoSz3SuuyvFpoSgzGTr5ihn
WYW2faB5WLznHFf9StX0/n7fMRyFw5FrQcRP3Q1NlAujeY2Jg63WRYOZHlUVLGzo6nJuBcSydDi/
QO8q3Eu6DLcnDHR70atdnOwqL+UVTE1IYOg13QeoghoKZvQ3rVo1sMuEpRdYxX6GPR+4ERhTWnqf
//wnbsGj8GpbjYdCGpYc7ZvYo8Ez+kkiLBVdev5sWZ41tKT+zpkeiYLUCOYeCU5Aqvj0+AySbw8P
XQAYOKy5AxeqvTY181rsPwMsDPJT6sc+Muij5j5LB01mwRZFiCBrrrHr28KMh/cpupAfsphlk8Ay
XA+f01wG73Qrl2Z64Z7afCHIwr2AaE9uoBdpL1cyBUjv1XcQRQkA8IyyHTFGp3L5fFI0dCse8gv2
y3pFqBswOhMm3o8xReI7iCOFkW6zUuHE+Z1/EqZKWhxbhhGF+6gRZDEGgpv31xxT8rdbIdrHO6AE
HSmE2Iy0dddorlfrjt67OQw2DrcBls7GH1WzjhDBAr1HljK1KbzLa1nDjO+0jisvD04tAh/0KQWs
VjIX6xPKp6KeMX5mnnxFG+u9+YQLh0/fPv+09F2xmL1UlJ4p6uoSL5QEnBJgWmZIEQk54cBiIaDz
80nfOZznFwqI214m03wzG+0tRN9Y7ZiECjW4r5KLampETZ01r0TS/PJJZVziv3i7jvbYs2RFrfRb
ZApZ7gs+S4LNDIWz6YjHc3Aa3w00RgmNE5KyhCK0ft4a6x9fFWPwjVy9uH2sQ1d0RhyXXgAu3eq9
7TE86ebp4cS36QUYm2QlstVXD3v1fzPRBFcyLkwRzJ6e6aHaGrE51sDHcHaHAqtyLUyEPI0aC8DQ
yGbKCq9OyTG1ESv7VlA3s1fr4xe31Gbe+jKuPuUJcyfbcn6rvZFfP5zK1pTUZv5G4aMeuq4rcj7L
to5w42CTQ4kYS4mUr2WQqJG+r2WTb/dyDPIqOEppZqx2PycmGLDoQiXHSN6dI6ec31L4x6do+Jj8
npNge2tEj9Q/qcTr2ws9QMLTvrq5ISZ97IZz53SlfZXCIDx4BUwDeSIAH4SxbVRUNepPWA+UoLmk
lfg6n7mALKfqzLLqDlTvLkoxDvuDBChmxxfmS6TMa/EGseUxOGAKDIv2TBwhtYhzR4XWS1CWyFd8
Yief2yyPWZBxghcK6aSKa6+3JPd+4nHXG9Z9CfAHJgYVfjkSGh6SwoErnMfB5uNuvzyvb+49Bi/O
Jf2BXyyXmxCDooiYv3Lmwd//N89JUsk4HAjgpi9ExHZ6ZoLjNYVK1qXtR8jygHsED54TwyxJ5E1j
tLDImXadKk/FYCoz5knvC8xVxwHsuirAJorIjz+2wpHjbWv5lDAAjh1mBwd33aGAEZFWqtpUSvPc
gP57eHuIRNSOGlU3X2aTOjYPNMiZfyHP3SdR8za9+ZjICkEEE9fibZ/CtGNuSITt8XSvx9ibUqBp
+T7DJW4624Win/oKnZtwEZA/+Y7BLbRcmj3SZzqBjFkWEls0mw29UsaLAQCTfn9qbbD3vx8TvynH
W8geTD7qvYCL0MxvboqHhcvW99PZCRnNmj0Tm170PkNjCGvdkqpw6P6LPt7S5e9nADAtTIJ1TBvi
GDLh7U9Fxig8xajP/gR6fu2CfWOKQ5plFe1zl21KutvqWpxjQBDjRpgYhuNyFnulEemAPhXPFFdr
2Zw9wlRQeHaIl4khkwfdwVQMgdQgcgfsS/vG4kpbQE/FubE6RJYo4jiaJsHLgOGoFTMizC1VReZ8
3oi0bxrbdUCAfj2spkhtVX634M+8lmSWxQxNvd1t+V/FCdq44DPubwQyi85gZ3JkAmwKEAdb5wOk
giuNs50cy/c8jeDZTIYqF4YKnxHCATJ6vmEqRN0EfLbkcVjR0hnPlL4ks6/syOtH7cCbD/v0VRNR
uMwSPCJfw9cIOrWF3qkZNbyLj6SICwJhpQT/zHnUUMRTQ7rdKHyisYwMC+1v62HRR+zxuarvN5eg
t/HYZIUIEn4MEy7m2nh3bvM5Z6LhrQrlTOtEtYjKNhbGrJK2sNajk9l8UpVlRQUNEmeKXpGXSMWo
V93/QL8t+qCKEDZdJM6tDhFib2sePZyZ4IlaAYBHOPRR4CjnNdeE6mLe/nRNCpdAk6C+2uZekjjg
3I/gNmsWTzQUMxeuQvl3J0poJBYVNxwHP4F6n8FfO76cZkrbf5ttQFad+FKetuGs/xUE2w3ZSDyK
S5YkhVZ8Yn/SoPTHkTvYRSSHIdQan/aPvDKnzJWJ2hIKSqg/0zVLKS2S7S86U3AFerpCq3TXjjEj
VNmfNVr84qgrr7jdeQUsfCoDz1Li+ecwQZZQlVr8XZbviOQrN6lz+kc4IAccW9xDWDLXNsXdU5xX
tK6MBYAoQL/z+YndeK9YcaBkFORR1nfN9J9eszv623VxXA5B4LUknz1Qz9R+n9yQL17BWriV7B1h
acrJqi5y8wPGonBFk5oP/pOKbDYD2BbSI5OauVMx3gx3yTksRbuhMysoEMRt6+FkoRNPvi7B43ji
aRcfXd1F3SUIyMW9rI8wU8/g/h1mVyP7V4GBGMHJdhTn3N/mhqYalo3QjUiN0L6/0OWGw2ZzPJta
b/WX3/KQALd8nSvz4Qs2+6NcoHOQY794bJAacmIrlXMW8EIFVMap6GvFrO+qapEADtVTLowKZu27
lFWEl5XpqOZzlee6iyrC1apQp0eQBhcoiHpGT2NfBL68EClIv3Zyl4S72CBfjsUoyDtCh1DgjYgQ
3/mdiV6dgJBm4D+uGWSfWR8rS1AexHDQR8RK/W5Pp+mUowy+MUf7ZOnpsxc6PqwufwnLnxu2eEgq
DLcCYTsjHP6OomMZhE6GJHjQVdpaO/iHUQYqQVkVASjQ770nbpZw+Yy6y3uO9wEitd1DJknPTGBF
c5sYP0KeaiPOAFdkCPlsNfQv67MDrB0FDa8mbRcHILHoSmAnG5+F3WZQYq5PSujWIdiyd1B9UdUM
sOrXLwAJecxfAOTdmoCQmzwkyhruSD6LqhCaBimfVnIUP4NkwAl/sdxTOkHjgKUjgsSrwQB7+Pl6
XgsaerCmTfJRWDWnRHTjnEiUTIDk/bHnbNabq6bAb/lm1eezDxTPiqBDWcNlKHwUXTEoD3xLvfwk
HWqK548M2TX5SK4L9aoo4I69JrHxO0GQrEG37RtpDXpGDSjfYIlxdzUBnqHpF6pNm1CnHc7NBEuK
Sew1BjdV1l4A8KO1zrpVKQNvO2y5v+PI37BwFISzmvO58LsvW1fVn4TMb7RzgNzc78Q/vF7OVvqf
6Pja+KOO/Jws6shOREc9tMtzPqwMvWm0tMgAz7WuLDelrYtyQLNDufHf6O4J1G4tDNs0ShGFPyDR
HlSG91jZCVkVheSqQi6fdI9RsmtSuaWm3MDeSRDaN7s8Xcb5c4TGvHLJZC/E1RUix93hPJe80dNo
NMPDZAkBme46fm9XBW6cl7dOsARvTAd2NotubRZtJWIP+6crjEznSi/7tJepr/kI2Flvm9FhWiUP
mlAEyWy/PYU0A/HV5Eilx0mqg42WgHpURh/X10NRmSQtHzp+/mZHrcnToa1LBT5wVCS0mm5S7U8G
P+s2HDCAYtQ4DntGWHQfpkSf9SoOX5S2xUz8lswlXqYFDLZ8q7bBcdNKSj6F1+rPWsjJeNH0W0zK
6klI0uzd/1SVCj3heRXvhBeSmL6fomU0x0vUlXqOpjdG7iwXTV12dvC5DxAC6gNaSleBNFVSyzqQ
v06nH+7O7Td80swWvQDZcHiyh5wuXfjBiDHVAUHyZnGKAR/ankUHixuvm8g9QGyD9iIY+DS/UFKT
OEJYg1IVWs6NAtU+zZY+ay7I6rRTEjCsFBkYxXAzYnJ0Dkoba1qvnOk9iHD+8FGHG0n5QToNvd8F
Ex1iaGwIdgwWPo/StHzrEItquy5Wc3D1euoltcYzjimHrdaUAczwLuizBd2fACLBPGWBo1o/6PJF
9Eac5Vi2+x02Q4Xz1caTXZdYoCb7NNyowhMBK5zia6Vj7k4WNadRXf8Xz/rKw4Omu2bqkSPk/0ks
YEduFYbz8ZVcleYZ2wuAeADm/RlcaMNHJpvqqm+lj+pR1Nk076z48BWiOX5hWRzcRNzhjQv/65jW
KE8VePfI0aeUupyWHrSrKinvUtPPPP5oHiXvOfDje6S+csQ0RraRPSq0yzW0K4oJe0SE3M/MfE1S
5DXDimYy7enc4YHH6lBV9HR/Aw5JDC2jYBeAm4xdeF2vg/sv16AJ04CannY/SUcz13AIoaFf4f/Y
L2oNlQSrbpfMq7+cZdbhzuLbIhUJBuwfY5Zcg2RrV5NUQMy8e4MeU2GbHJJLdPn2YMGouaAXOoyx
EhPLpi9hsuWtyM2lL43onQkdQCHGfXiTP/0gtDTvJ6V6t3o3uv5Mj7wVWRZ3qwZCgYKGEwE2Cstw
VkMxb6Ow+6OoSMu6ValhB2oZQJI8kYdjKoH1skspuX8hgp8NOUH2APEjYJpqZj359MEF/3Xc/ynm
8Yh3vLMOKFE/itK22Ka/L0O/u8yyd7JaB79ki00uG8RRL7bln2tS6AveCu5YtwuYqRQaUAlEE5rH
F+QPLBb6RU6QD1zHCd9U45yXp2ujUPuS2gYlEA88adBRLMoXuJzEabRZV5VBdG8jKG+Mj0bQ4rIi
nbpqVkg2ea/7gpkSBK4WvEzlALUCocqn47MUDlyOYzeqAISaMbyLO6ZBu7y3mY6tPm6od8ufPord
LLY7BJhJtnIlT35C39rH/3HZY3wk1PyWX6SeFlnsVu1p1WBTgvfQovFJxa/2gB3XUxTsp+7Y/hTK
fAIu8cxdFeiO/ETrgnhEUJSjSzC7l3GAsgwGUI1dZRb/SfRQOvJX+m+3dcZc5RBJ+eW5Vjy++dnq
InrzDJiCbjFM/sTKfzQ3yvHZOrRFvQrMueYriRxiKdcP+d/Wlr31CApdkCnIbutedf58kzntxoL9
DOziOOsLlkhtkReOmsjfyVAUWFpnXyZFXs21CuRZ2MSS7meO0Bq2RR1R8LaPxzIHvYTRRvTtCJBo
MHjX1XWcpm4JEaFUgsAv6WbCHruy8rsIkwqJGoOpyNLrnLnTnI50chGYiD5EeU92lF9uBf+pkXND
L27xbkw9niY8ZH1o+m7WTbdxgyL/K7b72NK6K1lW29ngIe+lnclmjZsSor0WvN5GrqJ//5M2fZ6q
c4r4Tz4lLZfEljGp1Xgoxo3AfRMqKhB1PSU9WGCtsh/YV1lHpqy4Sge40noVPDjKtdtqT1p27LvZ
kBM8e77ptU+/irPFrnQD0ruAxRXSXxHs0iAs0zHDp1xKRt/Dr+y4AVTW/QBSUieFfldzg+3uqBZG
5pjPPGb0JtvUjgaIfa9qmVUoKPkXvSp8buUyDtvGXrNr8Q8e+LcSA2U/I/JFRpMxkozqENd+uO7Q
pNKjDy71uSI5JrhMx7V1hKgUOWOhkSQpcGrbhN2cfo04GLnR/eB++hgIbgcc5zt9Z1Q8vfAk0sTX
6wGBeofQSgVETC+qjao8I4JNPM8gFvzn2dC2J83LpHPm9lXV+KRZGzoHY4JHDbdc/8jSxUhTP3P1
EZx8/K0/Y/gGljAOK6b36vWEhmzgW/wPfKfDU3a2MpgSSTv1ep9+QWebrk8/39NE82OVe19eKKBV
bB+r2MZWR1uTT/bK4IQqBNcRL2+8p4yhmul6AjVFipIUQdCnDwIqWa1yxKyWEMlBMhHNMMJ+Y3J/
YUqy/tTATBhlp3uzcD7Fom1MFEhi5MheZ11Rv3nx2pGWa3hXarOFUjb5DxRnBDXAG79H380Kixtu
M8J5gRZ+V5nQnDThDd3Sx4jNZ1PIyiRFXjyBQcFSVHAk+eYVgYymCOYQavDofh9FaONcoamkHpbL
fUNOSlNfqytgvnGUOn5HK/asCm5IwjVuJtVJq3KR3/txysKyddJXqYNFks0IDmjVZllS5qS5sxC/
w6UthH0ugJrqxlmRYHg+SWBN5BUdlMbNJZRCEVlTNnCYs56eCuuHlsX8tdLYjE61G+P978uALSD9
ZAJmbd2ml5hEj6mZoxnFsSUjcBP2fjGsO4MuJG8zXIzLg9P2H7bCs/mMFoTcPSOQJtSIw0/3LKXQ
p6PsMvLzKpLGuOx7O7a45+yWX9W+oyzHqZPdAc14gY+OHxv5wJgh73Ssx749iJsy/EathEIxY3A/
taeoWjYLj7S+4VaPxEg+Nz06zmUTC1MtPSnjWwRsqFOX1wvzruRCAWj0OMqSJdQrfDkVn86tmf3b
c90eZ+kMwGQcpqYbWTri8bSfmI0CNNNTb46WwiI6gUKaNabTOE+Ahl56VTRKkU41GQTzzMpeD1ZL
a0GSteP8HunQTZ5SCuyERDQ70bIEJXmEDYHRmCCIsiWAC51KvxSs6ISJAXuhx8TSe7QBDYAd4chu
1YmcQDNqJ4jxBG8nSt1wmLKbqAxfbR+ZuG1YyjYW004UKUkf3KJu/0Iwrp7j5q2T/AEaFEZvT2Cx
tNgILehMFXTCYibEdnSdu6ECl3izqSggeTm5gOrT2FKfuIDhZ2Gxvq5ZM6qyAEOPgrMuVXlG23gY
sxLkuDWRGkWWlfbV8NInLjk4qP3qMX3pTreCV5XpmqwSTd4a2FNSosF8DBSqvfoUE6raIMQeN++E
okIwlNN5sfESiIcRY/KPTHjJ9ffEHnO+fuoBQ6WEwQiK9itPPJWzkQ8xDefG+dsdAkjuz+GhWEjQ
zkvewEqew7X817aHsdR4h6XLlRDClRbkaxGnbSbPTaVoLcQYQht78JZMYQp1PNELC1DgbDIQacd+
0uSjo0cUSTHkakxMh9iMO3kfplgebZTdMSzUqYzP956q8qTNsFIgxd5gVDwjV6ei7jTZA5ehkqs2
wFA+IqrK1Tazmb2x52BU6Z0CeksZ4dPY7N9GkO8D36aAuYUimvVXOa2fAH3NXH0Ixdy2Wm/jdoCI
gBK3ce4N7wLv6mWdc0uLchYzGzdrhPLFzxKfv5DBADQP5AdoTo0I4fFj5m3jBEeSJ6A3uT1q39jE
rffU3UTn/LF/4Yt98khwIBH0bNaJ2QjIoHH4Xi7/CJC2kkzrHd9+Ho7tmG8vOgbKVHY0W19LodNj
Vi45dJH4YdZEiDHOxE6iq6yq3d0tRLUtRV3/4T5nQZK6qFTyh6ipGl6VZoi62NAjtBE22GVrHqVw
7Sut99pwbszG6o3ibeBkPt2zgdK6Yq5a3ihm0l/qsQ/Hc1k3vjEa0P3HJY7oTFVaCYoxyPtQ7KHu
g/Bezh5mDLovZrkXshrS+iqGlzEzt0yP2aF3vx/08YZiHxJbC/4Ul3h+LLn5TX2m3iY8GV2J1Mh+
AbYhA0CZcc08nDF51Jz797xDHn600TEo1AMltZtisqR/Y9CzubrFNT+2EpcNbmaZQmRyJEWEDFYv
RqbdjmtOdKgRlD/+XoMV9VpbcI9D1d8SXMpGLcXVDsxIp3L5kGlhZHki4GgaGmCG35njglpJa4q8
UwGflxASxyTdirJVVhAkLqWE+Gu9+Qwn3vKQ8Iv0gsL6/864IPwqUtNa8px1UfyI1NOGGhkf16e8
HzNVtE5ZBvTJ0BTzxJNC1pcO27VFyUjZJKfOLj1fvKPwoNSfRnWnpbiR/vxgQwfBWd+hgIYjmdz5
EC5x8MWBJ7Wj/itIR6dilOqDn060ssVDOcqWfZCKN2elT9yNcHGFgM3wS0kaHjb31hvc2TRy7H6h
Ni0/bH01QvOfrVwJVhL+VaIEHRuMQkXNVaiIHZVdv6bzISeDffomXl0wfIyK37bstGVruCQ2puBr
NBhW/RsyjmgKp0jIsSAZaghrLn+Y8pz8p45xtQ0JwSnMmqvPFPbEt1UT8Yij6c9d6cSvfC4gjQRB
/AlnYODSNRLx6oUOzfmRGl4UthKyWD7vIvNnkr1WNyar6ky5/xyTALxpM/sqaXM6a9T9bahBddNm
b0dK0y3nOLHcmUBhXxu1iqndnOhl+P+lQ/T7D0j7CphgZZEWbIK5PUSeuIYZXee/+MVlE22xGC+g
Tam19kDxLJzNfF9ViXMkz/KHux0mFE66Z3m12h6Bl8Oc4Ybr3L44ksbwsGcVwbiofJ9Q5IztNeAG
xOpr6Gf6R72eNgK3CQMK7kIwuu95K+3v7IvVfmuwXJCH+xECiwDaiKNqb7G8MKYa7iT6xk/75jRp
2RrGXwZaa7GK1hBkjVqP0cRqTpzFsXbz2TIJCSsV/kYiOGX4TaYsmlH/qBkKIsYOu3UFuSSzQhs0
u6IEYNaGeeBQ/qbznHrqf7ZgSuBynuBTI6JyDxNOTO4cBgbuPzVy8sCgn4+X3mwzm/w5PtxRdM8p
YFdKJL99jPjHE0hCyFE4YENqTMIdWZTisVxVU5vWb2EWg7zgYdtz2oc+OpBOIf5RWPPDrodxrZdD
of7NpSuO289dZVttkMkBKZJjpUso7S/+bXuqTB4auW0xeHpaKpLzE9LHr8FKW24Wm/jMZmNxrRfq
rHasEGfGdZi2FN8c/6ay+vWKQB9Ak+dXEd7PFXIdo4UrorOaYwB+oBo2ox7t+42iaO7EP/Xw4G6C
6jHxGbQvBe/tZ1CDgCui7hZhYkq7aTgX56sEHFwIgHuVuYlPD3C2sZyxzfg9w5idr/jRlhf7yUFF
XCSUiWvGzZl3EBR5+dy/byeFV5g/Q+RAA5C2ni0/nkjklO7Mj6iwnyFIa27Rs4CzuqPtaldGwMtI
Kdnpvu48/ziQBu1uRg4N2vwnpNRQKIjobL+nOOYYLPZrbc/VFTN5QUEGJlKSF3LXf8wC66I6EeEE
zTcf6TANVaPyMq4Tw8MN0G/5J69dBUGIfhQGENvuK7Rl+SGOmdgJkVmdeUJDT3hcae253I7pTbJL
AdN6VsYlKKv6/EEb8NjBdzzaDc0OAEH7C+KnBFYMp+L8DZYlwE6MPRRBsbrwua6UmJbcw5SfVc0W
dpsRTAdMFnSZk7+V+qjQOjrX6adyMiZYyCWcdlIO37ewcXyGQLMMhDY7+zkhXPbHDnT9QfUiAj2Y
Spgdof6AxDp3v2wiuibz29mwOo4JAvZa5SKCJqQd36yVfmmAGIiSyAHENOz+gPkcK+8a4MJqRC7I
jCO7vAW/dUnYbDSAjYfVHNQp70g3MWqPLq0/tiHMHJ7iNlEjMo5Dq5HLxI05ph0GNdUD74c4LZ/e
wmu7pZxOQnRBlad9dM2W2H96I+hpM6bD51n4nctCI0y2u7m47Tfv3OMIlN7mQYn960fvOlHC297X
fmps2iUV0RHh+J8mH7ZXW142eCNbpkRgcIGFR5XWvZRZq2mkvLJ4eoMfDxBu9orEJVNvfa/LwepB
OwZZ4f/1RTCpvQS0Gt+60Wx+NU0e9zmb8vkQJ3kc4g4ba42H8LifMtht4M2V4VjbFU+YA5ENcleG
94ah4z5pgXgtsrt/I7AIDo0+yN0QD79OR15SFBQDf4wGtMueIyIexn3DV91wPM9XczX3TFchKt9E
WxjkROaLzdTqcsezne8x2ZNH4XC/wRuliCMu6xV+zOmMdu8T+Mchzu9SvgRwFo2FRF02Vmd0DwiS
V6GFQ1wFfCwPlGDDTM7p3KXIwoFzmSstOf2K0XJgJV8KMdrrI9rftDeingVjEo5tjcegUTXv45l5
4cpqOwgguT6aVIpxeWl1uUxPISBFM0QZggkIyHya0QpADFqpekGJ6LCXhpdMp309N1Fl1gO3UD1I
AXi5hEiiDwNm+p/CGqOlm6vpSCl/sJjXHpXdXIhISEHOhdOQno/ynfuJl1RU5zaLYvGr5f4SIbRC
zlkS2zvzENBmF6kfxecPfGCAl3NLQlBzSYgxn/V3JTLy5HRTkIJW+y4AFwLoZY/+5IonAVh/f4ww
L7Jv7fC25p94YI1ZVzPo9UE1tp+a+mIQV1yrRhiYVz6zyK5DppU1YkJdH7CgczSQghJNRXvuUdW0
MXCnM5HPZY7Wn50WjaGPHld7RBAgzUHGtMJC4vCiC7L2SWd+4XjJrQMXEsNNxh9RC4yVownCCRBR
M4TcuQALO/QG922dQTNAQAmiWwGn19s0HCI+Xkam/3AeTxypUNTs3ZaMPQE9h0bpRvS1Jb27viyW
Mw4Ba5fP953+vJ5cAxUBEpJYIk170uKr2DX0Cf+XwXjam+gr9s2T85oKvJETjsa4bQKmhmdAfSfb
Vh5Why6Te7/VuqaLZ8/XHz6hjb40EM9p8I8uokMuX1n1EdJZAuasFcT65+GqVO3QsTXcXGocccR8
i5tsAWJSgq/JtWIn6EYtWsJdp1NKYhwgRuHSDfMlaUmYRJjUCaBWjWHym4v7dwWIpJak8+ksIFv8
x22d38HNDqU5mCCJeqyTvyg3mv/H7egC7Iy4BKmTt0wlKZ0T3hZhwigBZ7jrmKMOfKBwFZ8I+N19
uXUel0qFfj5g4Z5rjEY3x0vi843OVoZQtW/9mCbnFHYqoJyZTZingSM6puhdyH5Zwjihu3w0owy4
dK/uNXuY6Yg8G23ndjSGQdmPfKIIx8hNiCDHeLbBSXufNWWmaOiE8v6YarFdZQEbEcM8WeRH0vb5
ucIOE3DoZk41/8PRjPXd5t/gIF2jqniW3owmsrgvhOrNxidcLcBI7tAN5HrOvq2ZzvZ9j0inCJGI
bve1aMeyTrEFJ1m5LsJHQ1f+5M1S+XauerId3Jm/+sSYKu02QhnfgOu2qeEKVRxH5yNZQEcKg7cg
jFeg1xqHkoudAZTeRbApIo4nUFrvQMvac4kFQpF7TBmAm7V2IdW0RkKiyJqz6OAFzNooGH9bEZLO
xJglnJSpqC8aLvXRrYcn3pnCyhYS/MzGWnj1jjT5x6XuuvKfpg2i21eoTDv+c660zXq/oUHLgM+9
FDUPjgnVZtKxrNQSgMn6dIJ6zKXAHf1sTCxRiuA0VDLDYqsidXhEFvkkioyVb8HoW0FHEJilY5Ps
hoYJVnT3N3Gfv0xfvAc7vudqdrzF7xCkJGqVO1FlTm/E5RB14Q8bJfkSj8F3HEjVyMKMzfUB8sq0
HZIm/6zeb3JS0oYyXdM2xSNnEf/rDAvxofn1YBTEm+NugbVrCQeMsLATOZLrIAv6ko4c4Wgz68SL
/QJMbq/KhwvMaC/kQ1sBjc52NUg9X+xZNKx5/q2Ej+3OahmG8/QuzjHPhY9DYJaBsV3wfFl07Ibk
li60VHNtGIK0iKf8vi+E3pftNZp+9hidRQ20SqIArr4UCxUpBvkxtqdevAuqy8vFWlJIUwnkN4gl
YtyTSDW5xqqReH4gFr18+oTUyTLtxnYlf+/et4qvVsrfGPgY2T4vGymoPB5R7DmDivYdMA3HJyVs
JVVYX276EbcRhh7PfHpjx/BuL/yxzA4SdZlXIZt+oZvwFEvm0WN+RSYs/0rO112gr7s5++JFtslo
fuE0jZBNPXiknqwmoMDFXKl0qQfH7qLYlet/VNj4KUhQooJq4hUpq0ewlXEiVxhuBdjnVjpZ9EHB
FEHdBiRviW/Xxc3nUpaGJDduASt9779Gaujzpku3S/25zFg498tF40EQLa6hF2kBFikyNIJTlmSS
XcIQ36yLHh6o1cS9S94rk/60PiZiGTqfNnRESnq3/dojaXQhCIqLvyBzHIedPCjbqNlwlj48AAfv
5ML7dQkqt+5fJoW+U6q/B6vfhoxj3i3aNxvxit8RMcW7OhLb6U4FAMQ3qQxjB/igNZ0lApi0rPWY
gcBVUiOSMRnuCyRhalcxSQKq4o4dZJeKuCCUqSazoUdWWsnDXDcmBmAfRJgkX09Z9f/SKu5w1w5z
5Z3y/ONk8LaFUnMyII/cMlI+YhZh/16NOMFaCTCBKg0haJGop8+I5X5VammhDxu1szzWUTL4Ps7c
scs8kUN0QLWlhEGYZrNCKjl62i+fYWXr4ivVbc1EMEWXI0DpjRE5PCZ+PK+e8/RZHQqXEoaCoT2j
qWno+NgIOyOO0LLkaJryhxvA5pmB3zB9ELFw1xDTQd4Gti0NNHGjhBG7u68dVTu+KWXo/PeUzCVX
M93pn9nPQmUjShfyfrVbPAzDx4c7dnJ6x/SiNxZIKWHBAY1hIMebj2hSwcK03YChTM2GhgUB+eqj
33eY0POd1iH/TGS1fmrAAwihzUnTNkXtayldjbKIiSpYUiCwaGkfVrFzHfrc0w6ETykFfRpDBIXx
Ok3CBgFCS2VVsnnW9GVsvSX0MJC+PG3P9NLJIbyb4YO5cQMRn5Mgmbj6huQfxGOta+/FYbu5YmnY
GVVlh2osBUCo2y/I35BiddQAP/ffFaz9E21Fa3cteyyXiEPVbXjW5AkeArA7Dgzq6ev95aNXpBvy
qIjiUYG3thgYwg60zqSfj8mmhLsrBmSC/PBc6gV8v3xM0Zl5lY3Tj6HmOjsPlqYLyRw4bygbpU5F
PqHSDKRuxUWpNIKCT3r8FJtv+lm7/Pshws0GADSZCX6tBwa+Fi/H91qNHRQ1o1KZlqCAEZ7jAKCH
gXaqpJ4CbZBgERWIIva5/z0rgH5AP489oSRadNDIy3bbwWa89MCAGRl0cjcCe85fCr1SUj4XCuqW
vmQiH9yFQLhCmpadL1bl3xkTWaNFxDvTvKp//ElXmackkaJyNJwlnl/qgrnCEW/Hrd0PxRHf4+Ia
uYX7V/Y1EXMuNbFmsZZdJWWD6erv+3ZmOV37UgrpIP75RTJVcJkXWNcIDJbcdPlT8P9pGqxhOO4s
tE/qfQ5PGU0SdvqsCXe++yuVKQdfrHIfzNnwy/wz8gwH95n73b41p+gEv3JSw5SyUuvwY7L02nJA
zO4hYjL1eOimLWnSEdWMSL/N3QjoyVw1bqwyfhY3N6xN7kKCAgzjpQOJgA/wBcaRvbwWfJLt5v0A
3p0Kk/0gBI2k7VeQRLhZAddNncmnHVTO81RwFjasa6UWUMJh9ej9xlqBTzLs1f7Ry0K+0ipE4HMp
naK2Avjt7wYQBX0zMHPXvI6WDfyMPRUeQyP/sc4ArL8G5jOEzo7OXnIXu3s2asISVap64iWwDxF5
ZCtF5f/KhGvEVv8I0bAcLYoWM0kLOP8XxQ1t1XQ/RCpZDdmNpzkW+jxsc/6FJwxOjZTiyWt7DWdw
Z//YKeYfV7O+AyPoEl9M/iSbxqts7BQ1ha05CDjGrCOQ2/UN28uU2iVchM1GBxGn786Gh2i4iR1k
T0Z0BUOetb3R2JYDQLRp0FahmXR6DM3mAhjQTF7iXj7P2LgOwUDQUe9jU2O5VEjtoOpgrXU2LzKb
3k2109m3I6sMm1T3uhL+lcTTONNshMXaOPuB7ir0RwXtNNDXtPIP87FAPDDnC3vcAZn928uyccKA
901msU/JFvRyEcULPLPYRwZzZDlHPp7yR0V8SEU9Kc73F/IuLaY5bB5epM4We9rL5eMwNvK2upnD
UVZwhJE0aDOhVE/I7Pi+bO1TPo+oGsH9iMhlH7SxKoTZrQAyC07jgiKx4U8lz+bAlr5gQYHYbqFi
zbvwSeRNRh9Bq+n8XApa3G5pnb2zp9wMWy3FJcfQkUwZE2Srxka9bhk2PspBTKZAAkyM7hUjELhU
8v8aC8IWer3cDh4Jv4pbE2X2MXJ4o4flVCv7EzMRhW60Cc6xtUcesSJvXYA8vw1ubEOHydkFpFSo
zNe5CLHkb//qtd98l4Xi/5AvgvrVJk20pJHiDp/ng7gc7yLel4tM7ZVeynSVLtou+u2EFhYYZO+G
gTbfKT1gSwRO9BHgSJvqf1e1AYpR7eRmssbq0GosmnlIivp7dPwat74977peOqNNpOGiN+tl9Bjz
+tI8lVkPPoz7TNHwSD5QO2X3ekHEB3tvbx2EI+ZriUy3cViBHwXv//0Y1RCNhXXsfd8aS/4SJ2zu
CTJhihlyhp0ckDtSxnbL1tbhi4jPzq1+Z0QZ5o+try18rzQisdE2RJU4PN79WyI+NRInbJwZkEh5
ySLJVrCRxO/S1DWwLo2tlKn6/DHIzS79x9P2g1g8oXl5Q/gP2vK6KM9W2CxIwJ9fDPVYx7ieVK7S
eakuNzn9bTsOOcSJyyQ0TUSpS8oy2zfb/0GvdhUUV6MoPXVRPiljy09IKq5IOJWUtC6NwgEvLcwa
s4sMcDh85wT9V6gqv1W8fFuzA/SqgWQYQC1wkKO4RGvO9smtHxBza54g7KWKN7bsUPo2G9s/zv+7
REWApgCDDLycqJXSB8UnYbMJRXE+dtWgrZgjbgGgNYILv5mg/HOOKmofA4W5/iWC4v007lPwbsUk
Sm8kyZxASi2wYln/Ane7OFCI8wyCvDZH2FyUcA+APFdrReUQGMJma9iht70fpNc4cIGD9OfSezTb
HmrbXUlRXl6jT60rISpfC7PueeiJUEUU3ZvNh8H3XGAhY+0BvIMFrRFqEoAyWg097+I05iNDQDML
UrwgTXxQZ8BssiAAYCjgBcDZLyLlXvYMM0dSc6/IEGNbiWg+/oEPJKOM2SANBNrtvy3r4Vs+ctTQ
iN0KeT9+VsQvsl0biqjZIB5Sh9Wj86kdQPibD2R43AdYYzttx60k0e0YiBYqAOl7AmvriNOhC00v
6F3XujpDeHZpGj45zDDEQ1Ih7DDXy6CeHvfaSUzMLYZDzzbQTtZjGnb3JwEFPfiUl7R+3lXhgR6r
DXcZCAvtZe6gMi8qH4GwCOsMqddYS++4c0Q5Cvx1+9oEj8UvejXHANHdZ/5Qju/xHATAGzhNZDge
xK4Z0BwZP6ynF8jPw6mGnUIgoOqCB96rrofpQ2egGmPEOtFywbS/G42eCkRnbJOBkcAzKg2RU5UO
oedVDX45j1KYgGquvY4wMO+64UPTEQNezmdJifIau+YeeCAyrPeTM1Q/OY+LQcXbg0PJdEEEvKwa
raOL+M+T/U28wjBXDWJcs1hD6+cLqUbuLiR9R4bJXfBpfiP8Mnet7UjKRK6r8JZr4abAmXjt4Joz
m9CreSPZb7QIyIf8ZZFhQLfwVMZVTU9WZtTTz3eJEvF2T1dtPDyFx+K4vfkDjSs0PRmv3iDAiq/K
ZJQOm9yM9Ai+fHQc4SS/TaqEHjIvrR+I++vv80fRa13Bz2N3qpqflbzn2ZUroUCmQrFQWOwbWnQu
Nj+TJ5iDXBZo9jSQjLTpen3/LSkx2ihvfoTaVyI5kCohBz11y+OLZz3ByRS7Ng34VZsRyELIF/yW
KpWOvMEIOCipBc7HraibKBHQ/k4xYfZwN+ayPDwUM6/FG7cqHztnX58bdYLmVWtz9JdShZcR+2My
V9EJ9Ht5dxlMp5X8i/P0P78Qe1JuVYEyrvykUfeh6ujcicRHk3FPc2aG77oUapkocqtXvMJDigKz
is78YtHhbeTyWy8wcIcXP/PZhMReKClYOFdwFbgn3VKuKza6MqczfWQoEeZc1KirDywKbz6XzE67
UHfoDy13VvSobp2EnbZ/Ygr+Qdy84sIZACZH+JhHbeTgq1aONPEJfCwQHRrPeI9BAoh2BG1yf/67
HiZ6Q3SE3EB1Z9C8vAJ/D0ZKS869lUdgvptqw1SZ576MRLtYtsklxELbh5yovqV4r7tpvbp4tZzJ
Txqk2zGwFzXOG6r9ukVmA7yokjJKRxe7H7ycgVba/+LCOwpeM9rv5kYH4ivRLMz3WWWaiYwCu9ak
i0c3KRAC/3u2Wq5VXDKO/TXW0le7KUoOUWOmNY9YmPfOfytODZUDBr2Bk3W/wmtu0bjig+HvjDUW
5WuMoew5Dm4MFInyEW7SvXCVXCW6xlwxBi2KHH+FStM010hFJqFAwo+3WzGjp4Zg3H5zmKdBeHUF
5n2EsnMloFFabzAyOyIba8DSThG+0bv+NeetGCsMADWGt4NQAj37LWcHcAXUay9+pPpi2ycbyzSB
KBJRcmJ0sy9Kj8L1OXMRZgQi2zl25qSKMsAUmrQDyVNWEOzQoimPpJq3NEqpZ9EblSU1N0uSrXIk
EvbGikeoPcc27ByDO/j93ZmY9W6sgez8XlVdC0Q+G37RfS9HHoY+d35jP0eKo4/M7NlZD+O325ii
7q8cskNkj/N9fJUpHDjuthqHL1BhQ6iK+mvtuCbzUnLyt1oKE6TBysHoMLCFykZvwyTqkKhoxMFg
p9HLcje+zebq9tB+nEvwb83ATR/gBU1S06TSbzs7WdHPQ49kHsfvP4gHB9LvPZINOU3OtJp5KlWH
2hy+GQVqj6tjQpfyh1y4Lz+4cwYXPyn45U+MAQ78QWq0QTaQMIL2UchuWKnSn+gi8icEL2Fg+/mR
JiaKNeNSBV2MgeGhmqfm1RQ4grjcBsODFp88T6xsG/OkRJRs200vixvZ3uNLCTla0j326UOZWGC+
Gznt+SWn0bJ660al8wmr3idNfpCf+p7Kw5Pqqy3eYFYNIvrsBTAiJvqnqEx5R0iSm1wt9hrrBMH5
ejMywosn6V327HVYgIuvn1UqmQ16Wb+yNnX1DO3k3dLesHoDLg+9jE6wHxB1o4eUMLmpwpKLBI1j
DfvQHdM/5aRQ2t1HcanadDWi3hVQGTvDzZysOKqZCMAsIMpUbnEsP6VmMRZKF4/KOe+qARO8sk67
igmV1PWSpGjhYZVTO2LFCk4WHdBDJx4wMoU46ODJ5aSVB1/FUYqf0KkPSd+QE50FzuMwM6pld2ir
GwtyYwwCNWj8vOezh3lVjVYmZKwL3x7Be4lGWl8/ltsso+aXww6ka8Z5mW1c/CxGYW5AnuVfCbS6
lTJ07JmU123oKPAF0yAcgzhxsW9GDh5v7oXXSHQs4BUXuXd/72eoxbMzhzFobrk4tiutb9TiDICG
NrT3x2JDTF91FJQUEZB8mFf+q96wD191rHM0/K23Ntk5Up9sJWRhJyKp2Q5ctu+j9BWLN8pyf6zG
MEdLPhNfcFXcU4fMBiA0MBSrCMPnvnv6+OqAvMVhWtnGnEbE+G2w0GhAgKB/1uNgnMLPH4Hn7s/F
aNrMaVrqTQ+9L9K3VBchtSXfo6WrV05KUF6ZOX1q7D6Jxt/zkhBFt8VnoJR2sW0GxohYN0euRkYY
mqu26RIg0kWOYELWT+V0MMu4Y0PUpYHnJiX0GQq/JR6IMMoUFrN/sfpQE8ZXmM5KMK9eMexL+kNf
Llh8L3JPxBDjbGkNzdfCfDm8lZAqovLmeOipXnqlfxqCMZiUxl5jpMaMixnuRnzUPhLy1VRdFHN1
49SRIKPDaOBy4qc0TTmUlcKBm7CPMl1kiKAx0YbDiglx/382FiolLcRocLleC/GtVfp/to427l3C
OyYGs18Pme8s9Iz4iQB6RcKoCwiRQZKqeRrE3FFs6jRETCK2cNO0c3CgjSndkltrymXDbnz4y1cW
/hX09g+bXSDtH12JZ/hG9zxb9OIcD6kdviyl6lSkY/U2A7zZlfYzWEKpZkuddbCZgkjZnmTAPhaZ
Jqo6ze4RhmaP+DehM7W9MzbwvwCAUUaHsUMEKXrCjCfEiylcO5A0M+b+hzwucMOEykaVkHChjFt+
SqdZ8cRBKBbjn3aN0Co9N9VMJMgjvMwS8jZsoPvwx/eNtiEgmvAKRo+m+x6S/fgoqlWokhfRQNZo
Jq1Q4z46gh6niIF575/a+HlgDjOVnDV0pcHrvDE7vlcwpUHwzkxt6G0GtFdv5HUt18c/2RKQI18N
31HCcgUO8tERYv9gvvuuR9M8cHOQCCygxgoPbHRE9oKG5F+Pw5Hrp+md6wc6zSv/5rhjt0IvreJ8
sDP0j3HLb15SIjDQ75H8Ej5CZGE+X8O0MguC7o5tlAQqXhboKHaRGjjqSy+GL4BFUbDE+q/oAZwv
DymIwabZiHopSSOtj3jv+IGkSnOYCRNNupQrY9II7CyKylP+kLuN5IOfgfCJl6wQLBmyPaBu7GiJ
uiryb5mbRtGD90FKmzzSXsUAF1aveQ9UGGyCy/4ijOysUayfuEnWt09cnGTU+l3aWjmuo2w9kkab
Nu1hw3ivki+rwSA1btr50sRJnUtbDOlOm27S38kS7WUT7LgBooyeZnvFzHYd3JnWPVtu5WH0yNtM
pl1s779gz6+Ao9O3/+thEkhn+CR7itktQNmVD/hJWsShIwI/pCm86IgXU7oVO+rwFGS4j1pSxiAQ
BKhzk8weH1NsHRGn3Vl/hdi9KCUN7X36++snnX95mUw3esmJMjjMWRmqgJxEC76NBzn2GYxIVnAo
yOcovNJF7jXahhvjuP1l7iT/jSnhBn9bzy5Mp9jJAwapP/3OTdMjMHn9SnIE2yGOqlNiru//BcZW
WjPFYAxiYLVzKTq9Cd8XmCCn3cqankq5bgFucXOrINJe0EVeScrVMTe1RLDrjH7i3ip3geEpoaVR
KPwkyr89GsRVYfu0Ys8nBfh1wUqdbw+UCT3yp1K8Wsg8oBgti/O5MuFjX+uJvvi8bX8CpnRuWXbP
y4SfaFyii5RIIQ4Ju/jTsLpNayeshuwtsL0oNNyAL2iSGLY/rq9hS9ILGK8SF0DQt4FW7L5hIvQv
Y/KTvi9liCX6Oe3lH2oOmq4VE0JazNPudRLv1dCmyQDAzJpvBBYPGOmjl8rmnrlChD/e92nVkYJs
QG6wV6pyVv6osfy347ZNjLnLGgK3sZohqQ+aZ74pLi3x9+ZiUPAlfk9zopng69TkXgOYy3a87F8T
AQljs4YRfE3EFPjNVHIdplYwDiaJ/iCNDmjQCcsQyIsn11ohu5HS99Z41IK91woI4gCuVaahjCta
EvIptePxo2FcDNHLsyMubMnqhzDHm0lndtJrinwpxPfphdLhTQ2+czsQPxB5ikzJawcPSuPUloFb
Qved+QgTxofqXOT1mud6AMbb3C2LN98qGBRwSa6avzU7vRoNRkcErH87efGUv8DTRdpaBh6zHCZP
vJO4KhK0z0xEJ4RYPMVXfYRp97Wh/S9vHGiMWIJ8NMrkm1c0AO7HoQWh4ZuW3uje5/b2ClbhK5WB
WRIBBWOcADxKeW7H8LH6Gw5KDeJu6nogRZA/p0M5i0i/v6Q1KB7Ef7ar6kV3uQF5EABi9zP1AIIg
2yZC4HMrNYckm4HrLkoxkKjoNCtOSoTrKF0iO7SSwS9b6l+SITrQAaAevdvU9r4qctRu4xRJAT9v
sKYe7DHagMYMHoiobc+wexnDwmg+eL52GDJbXEgcKI7CxS3+CGkYkzkDPedYtynZGbWypLe0gcbC
RndgcE00tderbYNmlAM5DlaXqYIbCB6L3HiybGObMI6BuCxsK6KipS0C2OtCozxywlpoVIFDkZPA
eEm+cB84cb+E7YkBIVUAItUoPqqMUdEwvaRP7krfkt9tVyrAtFfW4ovMj5BzTA80HfNftH+Ov9Lc
KPdhQBrd+RT3yM8QDx4rK/PuJ3lnUQMNJ81QfROc+8nhZuHk1uX5bvNWRJSwQ2oOD8RyJdqQIr+c
dGvVG8GTcPV+Xjwq2Ytzs+CifU4HS2tKvv2dYShqqHNL8advc60nMmN04GEc1XGtxQzrr0y+V0kJ
hM/zhFi9FvNJq0Xuu6l+R/w89+Xe3OBJ+xyJCGMJfPqaMKIq1oKcOhL7VkXeDgYEhUIgj0MlJ2di
SNc0G9a6O/SNbQH6Yj/7JFsl+Otyk43pqE/qs3PPKTX3iHdlkwkz3GO6Y8lELCEBb8YXrvQWTaVX
J/LaqzJDYTwZAxZpvY5XAMXK+gk25lHsf6PgRRcbDHW/x44vcz96KdAZ9P7WzHEgBD5RNnt42apX
8jKot07GHt5H9W3X5Levi+VD2NZhXXQ9DE94PKnOirsRaKrLem/7LADF3i8wrNS6C7dexF+9ijX9
zUzRS4qhDnpR8MrDGOGflRxCenAdZKGZEhpEeJreEiZWRB7TYnF4+ZwvM7Mjt99+MNSXt7RkhrF5
5fUlkxo6Ezjtf9pQ2md9iSOp/+wU8E6Fthn1BqZqi9WGK5evZ4pDffzB2nPSV9FPYYgiQaHVMhTa
4mMvMYTx/V2xIppyULbCdk6s0XZ7Pn+7b6nRxDdf1mm+A8QNAM9V0YUA12Oj87c2ic8Fh5cCrzIc
EZ39KmWDodifZyHDXSTup8ZxtGNfk/yk5Zi3u4hzfQf9p8oW59mg/2STJWpYTHZTmxVnSjcZkLs/
nOdAYX5xznCnBEh197KHs4XT/s7KWrEgtbWvqVfaXolvBBI5astiAVGn30mqhZjnnl9w+11cLZsg
hqX/tVQPsG/J9lzzIJC169h3mme0JTQa9ONbuLHdro9Yfxhkxw5A1+ExChawXTNHwSMAtY319g53
8B4BgNvho9gF1B6NyFjf0huCTAPI7ik+lB+hqg1nBlHPAE1vGnWjn1r2yht+uKF2rIj8f0meiLGY
j+jh1jyhA+BYG7Y7q/rWPYfOndjqyVwLTU6hcWQ7RMBOoww+5xR2mOOC4Q/dFP8VgE1drZpQ9jfz
PA8/HF+88RIWD9TDwoDbmI9PIsXCHWdv8rcT/Zze1cK3xR8RFmenhTxRW6UnUn1qE9Vq6X6ZjyVy
gg2XaC70qww1HZzvGe9gAofMCowYQdANeLdEU6h6MU98bcq83cRDrCkoGEkY6+BmQPMhGG/aLaBI
CCC/BFKfPYSuTAMo3aXCajsw0v3O1UUP0tdKGSvUoJnvNMQVQmFo32+ZHz/ONOjfAGPwJMXhuwbV
NK1E24B6n/i/DIS8ens6Z3OaCm5fq2IV792x3AxfSWOsOntS0dNLFL+mv1o30ApyC3EadDx5CogK
ZN9akEua4XyWAS7lrW4P1herdOdRCaxPXhkz8PC44wv7Sy0h4OkmF41iHyO/3fsUzg441Oipp4mm
vOUhjXBMR6OrF0Rb0OLvuYm1pygByO0XHb8GfQUOQkBoCo/NvfqG/Z4E1Zcpp2rkOXRAK/THa/Yx
9mJ16UerNqwrwfjHbPiavqaN4NtDq3ev5kntWgqNWvAedU5ZikJjGjK0Q80wDpyZgwKRDAVPj0hB
CX1myVKqC/lw7FrrCZLdLV1CwNNeAQpDfmevTi4zcQDy3mLugpdEDpfv/W3HnSUdb4G4A6jshOZg
W131ZCdBhDHG0OWVY52PHYv6eVqrkzgGaTOeSaS814qkKTg1Yt3OVe7qHFG53UeMdIk+xvj1nI3I
d5Nm9jYI3Aoiw1gUwKKxRnGjTl7Cut5FdS40rRUaq+odEbRTlS3jnm/NpTT4GyZCKOFGVEn3WNvH
SopORHIn12fOx9/pOWF2UC5GBw9hq5YdJS6efKY13pOqGj7jksT7MABDg+xzwu1ZmBR6Z+r6lEmr
g88wLiLxqCnMzlGz9FFYB7fJ8BqLYptEDMdqDRAb+9ZWU10lDLdrgW4Q1+/hCtxx3e/lxQgHRCT5
qHhJBYxTzm56fhEVf1E95VEDCxb2VYAiADeRR/AcIbIkZMsoe8z+gKkBRW4AW8K6VgDBEjGsa4yK
9njPlp7QoJ6U8D8IlrnIgPI2OhAEHAXQtsXSco05YYeCJrwWveOeAxNJ3MlVo/A4YXPVtZebPtlg
sCkG111GdSAj+AiQgN5Pd4mHOprI/KW/2bh4qHl4QQgCOmGCOntIusbXCABzZCD0kLDFHT9PH0Uv
dHWXrcv7pmwT77Wk+ImKoQuLxB5rzNo0Gi2a9vJyJnIRK975g76D/nNoGXIyRG1KNlt05NB+RZGV
ue5PYq70bZomGyEqsPzbMEdPnzsKb2pDRrTcDP9r9XKBnSq6YPhGZUAkHDG4f5jrol53sPkKOChA
EqeuNwIGD8sXt5diwNja48+GCFj6agZRRJWCuElfdI0TVnNr7v2LEDH9n+yTe7+HNupkSBRiEKB1
80/TfwUN1Pg/MbCOljQSLTJm2VCHRjX4VTnrtk3j8xiNhJpCxKQHqX4qAql0su9faWlk/qMT5ZJK
4ilg9/dKPAvb4WZRPkPX8iwDTOfuPDAv60eiUmP+OE7rE/HshKFrOmIbyiHB68Ab0KmfRrOciQ40
371TLf2B8SEa6Zwlvmsnecr9CPaMmdyBGLrYlufvfsyVcYU9PW2q1yPiWyIPBA4YV0zQchOSewPz
RWMTh/imX5Jfp4IiOgdV6uxYtsYczc1qe2vg44NT5wPbzLZ77LHJFc4ohmxu24E05HUNhVJ1cLoM
K0Sx5aJQZ7vtjAWQCIsTfbHYfZ2EO6XHcAH/Y37yyvIjsH5YurmiJwgk91sM/w4fvyxyPc1aINd5
pfWh+DWWquIvykdKJZnF7rr7lAQZHPstxjHqAAX9/ZhKiG7yY14EXEniAEDc0Nyzly4s3EhswkfJ
wNc1MhYwafi/CO1kt60Vrxn5oeZF84U/v+6it3taUL5nRKZA32VlMJSYijrx6QxDx4ZK8TdHf8io
9zrTNeg1+94hnpBp63JZrYhtVSdLrWf90o2eFJ7k4gPCd1+vF0gzZ/8SrXFt+wHNsMITPKHF17PM
W6KI8vmtxtEDl8SUWm7xOH762LwVVnvFW+dPOHmhdRx72YUQcLAW84w/uO+7VAIKggWdqe6kc6a7
/dA53dE0+Lpgi+YkP3AXMViK30r1BSeiQbik+2g/ANrBrZo0oimhU3rhJO0bwwki5xtwi0XZ2ytU
3KY4Q8RsGJ6dqjrXMKR2ldcT5siRo2XkiRfL/njqjRZCareBVqBNGAMWGAnbudSIq3tPmqV2CArD
w4N6JJ4EcOxyZuhxDZa+28N4fcQa4qj/F9sog4OpgbGdwhKrkD+jH9dva9c+JreW+4N/ytVgPWHH
sooNd3Jb164cNfXRz/f/gbVkEI5Va7Hv71bVO5iJjXz1wRXR5aYKs0cht4wyGvDf/1xAH15nPuHM
0RNOkx6S+NQzvxqKDIYx2flvlT295mHKRmt43/EePba7vneMGjp2qg0GHocp02qrPz9GWpzTpLVj
l7G9y93j6Tq2Xwhpt27yO6V0jRi8JTk4ceqngYbeP6mVj7kPkHlm1Sb7DV34WlqZpSIEYE7dmREA
MjqdS1RZWncs6heaN6IBkGeFAZD8k7df3xhGZUuZHlkH6EtjFTm7ihx+Ofv/eYIpHe2yr64pEtSd
V1rv3xCOEdYzn3+AlhmZ60BUoOOUoWbCVLfkxUqjtsWq7ZXz4kAvyhyOzUHAwdcpWsgjV+TRvOA5
OKHaiGV5LNTFQzVZiKElg2tfEcU9w6vrkdCU+CsfoNRGVgtoq2+/LKEhfyd9lVDjNbRyOtKdXNJz
5drQ7NEVMUJarhatVw9B5B8j1vK+fVsAMlTmBNj5C9/QqL/ATUlrXqZAQHvQ67DLbYnB2A0sOK99
aEMCRh3jzGTBEpHb6so1eUVfJ/oIRNtuvQUM8W+v7kGpwMTg3Eb7lk/py9hs/fwmFtWjEPEd3nre
v7sl5v6ThKrrAk2kP/4Hhj2g0cnh8QAyBs5H/InF2NFwAALWtMNLaG1YklnbXT3x/AX6PuEJ7VDp
CuyM3AT1ATVLYxsbOA7TX0AGCm74nwlW/OFGj3veEdIYwLU5rqgVZacg1A21/sEgnX4sI4ovAnux
49ikImkgZbyjeXrhGMquwRI36eECEZYWzyvZeKnvboWoUXf/lAG/AW0UMJugQJ4MlFv3omHeCS8C
DiuGar+ZrsxCFuOz7hrUXxg1k4cItulaNuM1DolbNxP8yAmW3HrNHQvK0z1C6wHhfEaQ2AXEI7k7
cH3DRwgQ16lryBYA2Kvl0GHWhG42X89O2Y05lx7Kxd3i7OUs7YNDZ4w5RvDaDfp/opr6LuXpClJr
W6HbtfZKUcGadj7QcKfESEdFHtQk5ZGutrdM4BXs2jwJS4iSk6UOxK42RWf5q2/7jRQJdNyz+JPv
vZpcI4100EImYbmwksQqxXyh8Dhzmbp/+lRyVjb9w2Pr5HFy0zM9bNM6+FTcJDrYuyeofoQu3xdm
6Ql41yJreB5wXRzAN1SoFyCbZODXQ5tiH0wSV7Qu/jZJrPd1EH5+SlWSEyAz4rlh0h0gW6fhggis
4n4JWEAb8s1rVZ7uIgxs5LUovV15zUBaGzXpxah5/I39b6AiYfhoshrcqYtp+rfXRrZqYndho9Y3
Ym+wgR/IRjeU6ekCXxgkI/zFAsK3Mt/JJ7x+46Is9PNlvMm8Ed2daf5KCfm91j+ySGJiLsJXcqJb
++T8inKELf4bwyBVqq3AuiyvVPjTKYJlXirmh7uHm1ZslzBBVSVg5Stmd/a7XW04yXDCS2s1812q
FEsOk8ZBZOwoj939cjwUcIAXr2/HTDdd+/BePxd9V5Z7D5Fo7WyvI5+gpqjGq4K2nFVlRJJ/KAMC
JvyhVF0z1CYLium0yaC9saE/krbCZfxfmXY7EFdEqM9fYaZyjJPTNrwOYgEjdaVNJBl0chLJmgHi
aJN76umE7x/oRKxsppxnY3d+eMUW3lJieZ8HKviCPipqbNo/lv/Le5fQsK5qzVIXy9pP3jRUnU51
kgikimBiL3cSZAT4D40FuI9frY+n5fnivQArYBhWqH32N1lrYvYvttK9gzSVghWZ0qYYDtIglitX
4DnL5uAAut4In6EL6egiAb+0+KmkXK6gattIlXC9oyaht6roHM+1oU6C/G9jOkOunnrH71UIMkrw
WQlPJTZRYVY8sbcQa4XdtVBFNsYWfchv3aj+VtW+OCtYC9T2Vj+966Tt7hWSvCR5JP7f0zYc1oG2
nBhmb2d83yHsfNJJ8AjXXvjttgPU8g66d24aVVxy5FmJBUSaFuUNweJkCFY7aZdQkapfZfX7TERB
OKx9vpc1244Kt8tZjcxkLW63zulHgoJI0qcPQtP3Vjws9KDQowj2KHJGr7laEkakEPM1EtO7bJmT
MYgYHuXidIF/xnhxyNGgHGGXHqhj7sAR1Bee5Ig9tV1/+l8FWGAyludYjeYoI4IrUtZRJBEE4cKc
t660/eFghZcxn+tpntmVnIS/cmS6rwbZQxaWK3YwWvDx3FGovkBQTAZdLto3fGDzfp0JSiEL/sez
pfWTCPNKk7SynGW8inMw77K2E0gEvVwTwIrM6qcKORjDpPteMeWz10bN0PPEYbE+hWmW1DtmXTpf
bBjhfvafCStzxaeIrRHblnBuApJk1wV36po7x14nC5vaWweB5787dNF1PEPgDf0lfUewqDW52dhI
uRwRQRyRzRvpuyZAofjyE59281sj3I9PKSeryUTwIJmHzjDS6+ypMLWNDVIba4EapIDs/EHIDJPF
l3GP71f1nX9SnMUuDudCcmimKKBI2iu3aXGnve/S9JV1G6TtwzGH6D4tJiTWuaT56s5ANeuvWoAh
MOUxUmYeUPM1IbIHoRKfE6Tp8PjAvdwZGFzInavDvWaZk/Boa/FZE4GeWzSgARI9v6o1CKIrHRxt
mfdxMBzHzkI65dCO3za/9TyG6oKXWbBxnL+H7+HZSWJpVB1vRX1SYFlkORswr9Fg33GV466f9uP+
685zLLyrQ+EZDOQCu6elUTThETVF1UmsH6CberCmP+F+5RJGt8ro4k/RP8RzaZKadPhlxL9ye68W
+Z9ePskJSQCin2Isefxs5utV0ZXjR0PDeDnuBPM7COPy5lM3gj3YxKtZ2RjNG/tRZCCrzOiUJUQf
xaRRF8K6JaHdf9i82PMXNeoDfZXwI6iEvKzT9yC3L76KbLCPmSXdd7uHvS4R2Ggoqs1MGIn9Bulp
08WccBc5qKpYWNkd/NDRNQceVfxnS4zS5VHVZvan7m2C8kbyZtf5t3usge6wVjIMBCqxNMtKOVd6
5FSHcm5AsSs0emzB3hQa/+c4SEY8thU5M9/Fdqkda8Szlsu80DPdGSKDNoQICP9EHwcWQ5eCvNR1
5Ni7vQVHVzWvjUsUcs3mGXAHKdxlI7VoYq8YApbJPB4sbO6K88Mhhmk6Nwf1bFJn5uUrAfrkI9ey
qB/19L0gN7IL2RVqGMd0bs/EMrLk30E7c0IxWsbl+5AcoN4vB6c5+7E4EEHCmXw6D6++acMnVkCb
A263gWDbw+u70CdQnZqjXekKbJyFESSQq71PlcdEM+Lbht7STMzEiPgPupP1mW0NrgzDihrKDx7O
fCGmZ7Y56ngqEq6gedLM2SR7rMhbXHHhjKookBmBPhDVRaoii227w5cdlMiB5jis/aVKOj7mxiqc
ahLPbkzufV+UpB0oqfWHkjoYoTAq1figabuGtXU6Vwej3l85gXtCFLwZgZscE1hC3I91CmNb6aPZ
P5lpCkkwWiixmKp51X+pmAb+lHC6P18NpfYPyu9G4puYtjNLjWPCykiLmcs3kR3Zu9XFWoZlNBQ8
yidgM0OzI6w9jWL7iFixUeqJod08DiE3Bla1XfW34qzHMg41hfbL8QAntOa4WXK46ut+oCQ78NKO
qINoAjBsWJMbUN/rPVkvBCFhB498869lSwMqpsPJmqJYsH7iImcUaQIZZ9DPFMD0nMXO+RfPqwnD
iTy9a1tqZnGTKajFhii/qURy+do9J/DILERF4AxFyeJzlvsWRh4DUFACFpog2uxdSu+YuqUvfwMZ
4FtLAXTAsw6nrGlHAZsaMnpdrFyxkTufBvOigFumoW2SnE+DQlqf2dALhu5o/1i/K9cCinskewvI
QWeHnQA5VvKFc1PTANgkH88hJ4a9sV+FEOoPdqKGvakkx/1H0zyAdi90aBer7D0BIK3l1JPoRPpf
qZL0sK67kE0lVtSPy3MpOmX98hvkGyoiSZc11NoNwFwHVwwEfntYmS8PfLarWT4ycDFdgQ8mxjIb
dQlAlXtfe7EnMzXCSTi2cM+o4muux8JkigCeJiT/i1QTID4tJmtbTfxMKBpDXHe6eaKmoKzglbnM
wAfDed1t9EUb6q/JERpMCyLtkqjmV/z8J5hCx3I7muWmOGgYCApii1vVrlMcKcHlesPqr4vUmj3D
UXiO4qUG14DISuMnAWUfmmETvyYrgbs0ixU7bc56AfNMLEdqfQOLOyIAsi8uzj/y6gCrne46F9KH
DQg+y9MJssXmLzVZO/Cn9EyxeA3BkR6C7+2yN4+0Gsl6dMNSLFEkiE3p5zhduUic5y7KyXHJBMvN
23+RWNyKUS8AVIYJPY5W2wImp/lHgLikBEgrJ3wqU7dMIVyVKlETvu41nUPyVWzYhegCn8638giZ
dAxR86iJ0S1BP/AmIjfHBofAHJnjDoguRAkUUIqe0yLzXmFdmGMuUeR0x0wekInHaZuoF9fZQNnx
prxWiBmJFZM+vKHnT9XkYoKGhckXp03sv7AEPwPNa5hUpNCh/PmLVJ1SK/Xj+9GMsWUvMKzOhaAo
vUiL77eoyyIQ+w+iWBAv7dn1Wz9qn+m+L3eFPvJbgx6zGoDs3jSekNY9/ASWGZoOMAmKw0mqcEDZ
bkHqBl7vey/Pq8xIiwu+ssw7+XXcJigex/vH4jZ8Lh4FJ5W0PUIX3buLaH9zpp/1P6d2yWpLScaS
+uQeUF9h4+Ax6vJh//22FUNyfEx9ryqpTKcz6OMqm/AmgvbpWSlE9WN3I61DUX6XSfvorAwZQ8So
0YDdtsyjaf8ZJxmQOxnmr2EwjJ0UF5Ctse0F7aalXPeqcSDmVU8HxivAZOKkghkkYb5r4zktc5Z3
msKxJWtSll2GrsnqFqbKWZqlnYw27y5qxh7Rj1qmYUf3HKTdhl7joEUPUvEZxb3evJBOTOznGJu5
GRCsEcyjI6nHO9sZ653yVZZaJ0DHtoRw2Nx3vEcEv7ylwRZOqMfI/WHYRLg4hdEPaPbcsuudu/yp
K5FxUJ5Ryc1Q4Kiiqf2oiY69fvGmURhIgQEuW3KJSoXho9bHIU6amqRpDXLUCCTMSf+RdKt+0WHo
Rd7KIBYLwcLM5AcBRLY9ZKka6MlZpFZEpH4h60D9j/BfhDHKdtdl4SBbKDKuAX5J5rXLvvTyYNrH
mcVNqVEuWuDn488fnOJSnpznlOhRVlBSSqw41JprnYof0NYbiVFeoopr6/MfGBOLPD/yEK/wtkjU
q7MqtZKDPgo2CInoa8pPijVrBbP18k6+ikbFouDVUDP1xHa8CcLFEUuShHDa14qAvbIyV4D/XkH+
abfiMMt14VYsP4jGi/ugraVM0DdSvzNmIjdtmILdmjmtybc7cIsNbxHO+0rVdTH4p+rvg/VKVMnG
XsW3NbvyTbiF9mooJxfFGM5MXdEB+jcaSXhcbMPNlLNkekGIQqzQnyjr9UeLXWtIcv90xdPCYKer
31CYt0KvdM9AVrjsmlzWuPgWlwsooljQNrWtexumKyzuJy9bm9slqZzZjk/MQNOke7MfsT7W54Qy
yjb2/TWb7LYwsQB65BrIe2pSMleDxtfz6gu4abEqtS5lhcFPsM/JiJPuznRppM5crM0eGWeUtEEa
QIC3291eizC3UWvMDtLxImkmegb0GF4T1I+4MgnQjQJd+T08mBoJF+PeLRh743Eu/+X8C/JyJQ0a
TKAdqTvYz3I/pV9vyA0+QvdWTtgaLouSTAV8XLY+t9W+XsQJ63sH9XIsucogqFlP6lOH9msGk7Ec
zVXKQLdNkrUS51iyT/OpdP/vu/rn2//krRmadrSBHFsPYK7pKg3Y6FzkzTC0w1Y/9W05syc8/981
wTOgR1NvQ8HigNl4mewMd7YnHMDwJyrTgb+/3sZNErGGmXcyAzYX1viAvJ90uigI2LRHlr8Zw228
E/j07SLWV5PsYBuqJwic4WWIG/XLo0qU5vhxCdkUwL4R6Xx3r8gIOsnvwRfYSzgE37QgYfhsqg3Y
cWkAiG5We87R8DzNC2Jo9ATa04rT/RRT+f4fi67Xk/UQOOm6jeTKT0xAt44G+MzkBibMq8LlQQU2
FN5WB/jLiZBU9RlZSapYdDk14CdKVuDKuTrszU7BCrkzOwXFFZjmhYFHE/KYXNmK/K1URHhlSbcH
fCNpXadPpvAomfaPloJGSNBcAm9c8xi4gFpysvnLjIvcCVsmYmujaalAcszSlpIn3PZMAnU7MYqT
t29KL2HocpvIH+rmAD+U7UgxeKgl0nkmGe093mnZVm2mrTMoCaS/LyD/kxjbaA7jOIGD4S+4fLYw
uy/VblI/UkUOAqeAQSKI15DSsbCqELmq1qfZ5YpZZ3v1DNZPsIuuwKSVZ6AlBjbP5CJ3zrr2BvGQ
A6/yOpTN9hG2YrgcjebmSrahFp2GETxRHnMo5jx8XR7VbE50XVBnJbgr/XvHbK+eAyQh30fVpKJE
u66dRlTa3qBd2aZ/LcsSj/vquPALKwXepaD99hLOMra20g8V3OiNu2kTnpsJjvhBuFbxHU4tQSv3
BHR3SaQJaNnFg/w7iYw6v/+tgm2ohWE/hAAPk4d6W0ODxa2aNQf9RaPLaEpOqRAdmUWLfIULC9vL
SF8H+1Vv9KjL8no4YiYool9Kg/Hde+u99+QfKn9aoMuVI3vm4ZzMv4PkHevlofCENw5O7zN5zyAV
MRJ2tVE4wgsqGY4gRbcmkAEPTkSd2pSSY6Lyw6YDFQ6mBeSmm7UeuvePTiPJmZ1wfnBdcxEMLYLp
jGcKEPgD0PznDtizemObA0ntFdaJL0hyZWJjIQWRISehKMSw3KTLWwKrLY3yFdwcNw5DZfGubkaM
jzxUHFU2WJbWyvcu8SnV57MRZOn3XqdqW21fteGgKzAlryYUOLs3Fkah2Z4Y9SlTOZLx+K57BLlc
M1btV1AKtNHEVUOEw2Rie/HpjY1oaD2daSTMOSbmc/BxyCdLPR3QH7l2DVDbSArfDH24afobpdo0
i/SbCuNbDDgHMP4W0JAzrFg+EEqFPcO74tpNKf8fEGTdCB8bPHnYq89olKXJrjqshygxFJe7F4w0
VK+779yRkMNgREc7N11EekiqlwhhozPzvOUHv1ncYHcBU1bvXEw+8tOnEunJXBStACXOIJMOu/H3
HEMx5IrmbZX2hakRVzZ7kwALG0+QPvHvmpEyUy1DztDLnRlWhz+6daQTCdsRDeqsj3m8TO/DL/bP
Y7CR/UiDrFSg4178TslKnX7eKcalS6MfKPEEVGMfTnka39X7ZqhLdAadGFmRZjtzCF0gi2Gx3jp1
Pkpn5ITu1+mmXVNd4qcWob+DlMuOOZXu97BA0wjETViYLp4WXqVxzQxhx6TVVYN924+os+uihzHa
t7jTfQeOgfg/+lRv7/s9yDpRvguFKUYYG0Tq/BJZuWyyS+VcqLWDIMJw52e62E2oa11pOUM2nvjt
9hIYFEUvPrMFjMrwvg12Vjxi9Jw5hWvF4B/+9Wuq5SsXewiu+C3E5+beJQw222SucQVk/ITvy0r3
kyIAWJGy0WWG6C0xIc6Ae7EYTHL0vIOJhSXLJKlnQotPbAgU7wZu/BeiKM+XbgnR1fBOQJ2i2TCq
F1Z1G/enDdT8Q4iA4YHyLnGRGMY9427l6M10EpbhA12IQRmoT4j7Di/n3jw1PNplIAS4lLvvqFGh
N+RACJIxDUTR4/qSbqzmpafhm2ogXRlD2szBK/n5ShpgDYjm9MiseLwMQv8Thd3azU5DgTG6lJVG
kEKvOYwhUYgGiToq/s1lxLNWAuVplGSwaevS0XRWouNMt9Y3fV209pChE5u/nf3otc9HodrPo1ck
wXIHVyNL3r8URzQYX85jRs4RWSySGKXpOBEd5ZzYke/xyeBzjtB4M4o0qKFC20ZJEimkb+iRC0z1
R26gjlGDnE+FIHVImK/JFOscwOuxo3/ZOckE18NGQ0BiLmlOeHk8UaUFDfsqcc3rksEevi27moI2
/O1gl8j2SoFPQ87Mu9WhHdshFCIcMcQMEJ0U5hoAUOB5E30F/nGnWB/skgtQhwDQEXVI3ppkqI8U
HY0zuru3lHSUH8yPYy3arVFXwaGsrY9ZRznqWIL7/d/eNUMToBDcxNQ6KE0YvZl7jBXaG9hTRih4
zjRo3FqYFux3iQu8sLorK0FPoqIb23vOXdvmLxuOc+jOVmQcpvhTzmpWMVcnHDMWDvYmScHDGTSA
NjX8hF91FG9aMJA2m+UPK19kKnklkt0/0DhU0Lxtql0xQiVJu+4YUEV4KTfh8eUf3D3E0OYIXGxF
FcP+V4vGTAcRjaocwcKN4mbUwqBG9EKRyMZXtMb6HuWEK4/CV3hm8gp7gpZ1uDmW4GZqXvejjyIR
y/KMUYvZe4kZh0QMdEpiN7Jy7r2Naj39CqlFeqFfRlKS7i7ASlXEWfS7GMBCXp8Ga0nrIJyicdxP
VzNPoQUH+lKtDQNDCLzc2xY5QOiNP32lW49iEHNcTT8pFQmOCVIPA1BJ4d7qmu/x3En6ks5wFyVQ
NqbyaYC2jpZzIj0SoIV4cQHgTbs7HNk2Dmd2a/n6OEUHgwENg9tkUD6neLnRV2XgyThEmWbsdLYV
uiYAVDr0B/GiCxzNwD4XyIDYmQqkBGLGrcIBhzwJvoW6erhlVyXUaSKKEghnCyANpakbg57UWq3G
JMOTDaiJSkYg+t4hBENLHorI2RlbR1JCw0jkonv/zau7N6wqz/ZbEIbu5P1Y6WGLpFxMyq3uJbYs
bB85l5DVqTxcDTj0/8RV3I4gJCM6oVSu+bZzd4Lyx/SDOOx1nxAo8LLBuExcDE0115gdSOg1Ry9J
gHdLsqsF2blzMW16VccdatiuOtimCBQ1EaQ/orjZY7Kfzqj2lDCDKeYTHpYwyol8N1yuRXVXwOrj
zuU+bBB7XF4971XGQMVtAVFvRH52F19Vwqju3pgBZAMfqibbFbPtmP2QBdIbO1Fn7cqVcq+1ARPh
2ek8DqltZsxvgyzcSr6O1Y0gq5Wd44RZ+PHxYLbT37vQWFLB7v7rSQ3k/rCSrh112pMy9guRrKLO
vHbis6kdlBwXLIlNgNweo85uz5RLg1idy1d5LpL+aR+L54xtgd7VmmgiF3aukSUcR3mYFulQ52uz
84ZbvEFIzSvcyXAMQ0yiq+Jv3zXVtNqINyBCfbZ+y9Ih8xlJ7ShTZXP1wTJv/pR8dS4uvGrTxLA2
ziJKpWnZ+mACN6W7ZuFNxH/TZGcaL+OmAFc1jGgfN+brSbmgRUXaDlqU1VJECoHf+D2mpHyJsjL4
+wJApAfgcoS+q9xVlSQWEHlZwZdz2gUfCTlzPiQBSyUsOVNPe5b07XcuQxiU5kUeMefV/GF7ELsh
AaFXmy0UUfFoMfdGNt9nNGQBLoi2GvB8IIKhMXPCSKQjVV6mdnf+aehSugt3ZWs5djX2oFDftaaa
zWRbWkHYuaHam4txq/jev1qXn1PCdqCPH62IPehmFoPYtfXSWfbv0cRkJt+MzmfZ0u4BPuLcEUxd
A7q86uz6j69O/zVChfiN88ZTdd9Robem8yNcZKFyy0cZ+Vkv1nwfOuy31/8CCkUYJlPji33oREHI
8lJnb+AxsJ3vSOgFHeeWX1TJw8eI4MFlPI43goutiZe0ufM+UZJ6b+bhsB+dlBkaMdt1pvfhaln/
g7iednoFzrc4VC0kNbpiZAXAMCFhEfHGIXKpQkhTGyfQMr+t9/s6DPGF50CcE4ddavSB0dr6M/es
4q5W4mRFA0XkB1Zb6WyrUT6Qufrr4bzh6ohXV8N3X3MXf0mqNZmvWcAiqMjpFUirc4reFWD8nmKS
FwqSc99+ioutJ4C3MbVS64WV0ht/Hwt662bKFzntuqKGC9iyMiu/suhA5U5iq0gse/OuC2o/BLpY
Vv6TSomvKa9L3ADcnbq5npeLcrw0VgLYEAvFRhO8aFMgSR8XXS8mP68/oLs6YcZXbXKMya1wSNkf
M//+H3+h02yPNrCDhNAINZAAq10421jDq61vtGvHUzc8AM1Yb3fO7V2yEnzu3CMDPX6oV83TrvMF
yP+9T1wPWi+3tyzrCE488AGUSAxq4U3Fn+1eNVRJnP41w7yRCT+Sj0SmPaD9dyqt0aG0MIUejH31
DNeqIbuekbfCikr7aNXY+Tark61kTuozbkyChtuto+vKbzVXYWUIcqO7hwAZKMXF8YjQOAzTPiGK
cOHtdBTy4Sv30/KIvSliXFszp6YJJRi7yM4UvkUVV6GIdlQOVY8DP8jypCyJ0Mi+F+PAo6QoIbI2
S6VRphSicOGnciwWbp3l1iOxX41wrMzMg5apTJSRSvxJz6T3eVCCTfO9nuuWZI7UsgWgGzZeE3Mm
9CRODiWQkpr4ei4G2Uj9QZbA8Ki9wbF4yZ+NylQNimMXoOlopV9WdW1rDtSoJMplrP0Ro8BdLUhT
fkJHy1nafLpvZ8w3xzHaGKBkmafAXt5dAJI4h46Ifqom+JCY8pMbxp4IT6sUWdIUyJBrg1fOJ2iO
WxJbKkEqzVOnShOXy7I3/PCd3gIYgZZPMxl8HpWMh2tL1wJvX2O9TP2gvECh5un+vlW7MUTHJrdD
E7mNmYX7AnRMZ4oP1jh4Q1Wf+idIAR8CS/IJarYSdNSkmBizS5qlqUt+zDJ5EpiKXiTizi7yn9ah
u9KD2OT5wJwUWpulgcWG/JlIcrQ1joKZZKR6osBdk2WHb3vqaAZ6w4McbtJB75eX38FxOirjr0JK
J83213ZRsGNNo754bJw3xEC+5m6BNw4cgybuAP5L10DcGKdjqdwfRCCoYs+6T1uyKg3Ub8+P+Lm4
sqJ6Pp6qtza4ezjDoTYt9MB37G2wDavtdyPJe5WuWlYS4NKk24pNv/4zo4j0XZcBMRLU3+xlQQH/
UpM9VtJTZQk71JlqFUNbTwI6i+FmjZhrdz1zM+w2ixoDP1HmB9iZT6qjTAP8IZsaYT2kPVtufw0B
8rA4PB/9eLobuh5QEE9Fy3G1ZVByLGB3QnGLQ5p1IdgjvFshQuqxkCMNxA3jinHve/A5eR5HkwZE
PyUr4EfhaC/nKcueMFXjynXiH2kkpUrzhzklUcC3gUpL9YbPlbGWqLbRVkGkdTOdfmm7bUGG9Fg1
TlOy2kid5Ik07XzwFo4O9nVEI2zb+ygOID0vvK18+smrxLFdnI3wN8mEr25LN+FfZuNMmuCfTnmd
zj28wsMunv5ei724Jd1hmEaVESrrwzTbsOHEt5KcO8MKdcn30bkuvdu6ltkzeg+ZpMh48CWpFGD7
BRAm3iPxWMeoOotAprfAlHQCm3Upcgza0scYmZkrCRJSjyTHBllHpjr5hIrCTrKJdlX/6w4Ls+lE
cqvUmMB+2vNoIjEWuv1cv+uvErnHA7WOfmkOIheagfMO6Tp3I61lGE+76rzj0HqzH2GI2Sjx1Bpv
dzG5ROa5PufYJsMzDdwjf8NfvEwLnZHvE+/65OqxseOg1hYGcc+bRHiY6m5h/1kclW0ezYx2dM9T
2ZWrrvyhed3Ot2q+eH4yv0x7dnIb0Vv8DWAiMfEvoYZLQxxHQ+t3y/J5g0XJf8FIEemh9EG7tjJk
pw3JEtGHXLottC8Sf8S2cf3qzmfKDoOmbu+fDOyZ+d+zlb9EQji3DmyVlc02SN/MAQnj2OpXDTKn
k3RqOCidD+4lJwb44K9jZGo0+EE+pIMotz89FQ0tSZsDCi6BUegasflCdDtqAblohJIyofTnLbzR
GkHsJPHaDPFgCbS+Ugix4ZLApweNH9kQYJ63X+0v2Ij/ANGIo57r/N4MULDX9sr6seNovhyzmgul
+udCYeuWXQyiHfgEJDdo4IjOPhFkhsHRToGWYdG9vnsoxXhVVxp3t4tVfM5jWyH7Tg23EG3KzEi9
WfnUQ3zeCmExGAD6/ZPfrgJ5TuOxZVcVF7DymLZ091TiRmrVEYVoQIyubEa6ms6ExrqbN/iKfK6j
zPb6Zl0tpSF3CU3Oe2oCBYr+KkAj1P/NZCw/E4rpq22gPJWQNcOkYdJ/8RFbciPR2Rg4kllT3fDP
NJds82AJrfyjddX8f3BlfVvCaz5OQR9TN89kMqVPfiP5xGRFcccENZEFtILFO7pFfmkb/pnO9oLS
WNDkZ4AVslu8zSHzi9JTMvm54Sp71Ax1CAdVoFENRmSUbdaxDokoUmwEq+2ho/fxyaqyTUmfNuBf
dF+/evvo/iQ0K1nNMPcAwqPVVEKBA/leILT9+fpWpLAv+xnybsAOVT8Fj8xzUEinz6OElI53dw6z
uEB8+XfqLqw8M1ui7d9OQNjamw3Ov74Doswqsc+2E4Lrp9vDxsuxktYA+UBvg8CIaRCWBhXTwnsK
C539pVJLFG4WMxSyDhRym3jhC/IwnURld0KvAjJPuizTE4LpjloKjI0LDEURKuPOq/tNRs/iIgQl
59ta8wgS/8xG2ZxiGDwUctDKN5yNkpJQaMo6o9Gkd5OePeXHfi3g39X97VmdP6HCUt8ZRFNEZ4Mv
BxdEWq4zldPCD9oCdf0wiAtDV0lHR00iFh3MJsnK7/KqLOFmnqa16P+kUHTenFEotV3FvR+eRVwD
36I3M+eFDdGZYjckpFjplWONUl5m91rUbzS0e/56WGnJo2wPRR+B90UlSPOy+4YI8Cy0Y6Wtb5eb
E5nfLY6ZIzomRr27bKYE28NnPbOCQ1fqHGPtQQa370AopQa/ntV12hV1FeM6nHo2AmLJEZVB3GQQ
5mALEhDG2gqr40RtpWACjmrfOP6cXpSZ28KiwLFeWh7/JNxzrr8cUY62ZSSt5w8QvjuuZmwrmWyG
Kf7uWLEX3wB/suV/hB6zc5gtFmimNeW7leu5bWyjcNd27lONUPHHZsYCODc5n8Oa9jOppV4SUv5W
6I8dvx+RNbZsRRROB/d6GC4FPEhq79O3Jqu3MHWTzYdm4jfH6SA0BS/JmpctSE++EkoJhkdFxFRU
rsXym8TuM3eiB8GR3yKZRFzXst9JBZLjZgJC4GRoQILQouXOYnK4w78VEkMjMHZ1STbzRhdkhGJg
HyCGuW7StO5QknuuyGn4eoDULFy+9CyjVoHe6G/Bbm94AUWZ2CBRCcjtwf2halWk6dvBPuVtNAnJ
1pnXnaYA4483vpkQ99kTRsMdbvikNFvjxes4zB1nSR/eKbzJ51BAsX1L3spB3JEKiqxymSj/fXeq
e16oxYtqAGD+Qr1t6YCZTURVLfGfoD8tmsPtjvSGotzxACqNwrYKvKimh94wNfBSbTAPRmrZ9tJb
s365/LViW/GsuaKGaYFtS2o58+QbNDNv9Lcbnt0GSMIgBzlQ7UH3HrHlFuzU9K3eNw/Wku6Ok90F
vS7vQ+8VHEuCEpmDE7TniRDaGnw5Hd/GftXfCvsI/5CiPfj7AaSPuQ8DaAM0UhlDWybIt+i+29nj
WSJPdQ67pAvyXJVQIVDFEVCPVm0ibw8NWOBABD/6u2Q12Vs+lnb+JzxGHp1bJtLDH5iEquEkkzxH
yiw97trzygxUgs1UEir4bc7k1/ZHZC95yxOlAAbBmaRn3qTfSg8O5mqcu/Vw17l5TUXWMqs9zDHf
OQLb3HupvX/XNx6q/O6mH9ekmGyLLfJOk7hDhIbOdQ6jF7/666UMK5ZCsb3zh3QXHmlTdixMEA2l
6Z0r23XCjoFM4qYG0NxRT+7Iwus08CNB4C2R2KHLTrO3NJaq2HCPveTavIm+cmLa3cBJh4oF1XHS
eK1BXdvq3ebhdVu6DlhSzvBpGu/D4HN/KgU3eJLOfZqsYNIs1MRnMyA7C0vegrKqwEej61VgcKJ6
SqcgQ7ZH53OWTaucJWfYLXOENKymsh5mpDqfDgRyzepOHrFxzv57lDAUFjPPpkzjcLt4dO8TAIZw
5FEvE2XWpgfTlnO4f2lMvF41Syrba7NwJZqEaT3Qo/whVy5dk4T6h+jYyeSXnDnsdDv1V5AbedBe
ief77KUzZ440tdIlXxRk8l+hkwEe0iygOlChbaRdgNDQRRMRdCHkZbSP13stt2CouFoF7LT0QYk7
4P0SYfczRQ9Z05HGeuUf7Zuh9OGJPhmE0bRT8gaTKyVOBiBfw51KwgEeg/wiskzxMtPV5tsmF/+D
n2a6WLO0bDWRtiHvStitrCKgVvluxxyFZDdQSapOdU3fRoJdzvhqQMFwOZHgP1XDUmZcmO/cvKC/
rX90KxMPYEoaA4jc5XwBYpeQY37nJn7nww4wBQarsyZ3k9ESb4YOJRxleD34UKoXSjg4LPyji3SA
7XXQ1MB6MkxWi4dVse7jzgHg9Om0439u/BmKSV/On0IVspVzAkk3JSqFnSFzNU1uuwXW43LnhfTU
gP2QXUdycUli/r3htwaMmMtYH2gARh2O6A9huEd0aeQe8BqD39jnH76ztiESxr204zyYGCsOYaCy
PtLuFl76Ysgj+d45i3NDv93Jnm5ROJPpC1krW11kZPh3yuV1Z6tpVLUfysN83y7siGiicdfPGoS4
lurUbopkB4AAmGL/CP9HxNwtlVSoy7FnSMUYhrftSivy9GFp0cBLsBgumCCq8yXWaFGgxqJSGvHX
Zr01hgnJcCKcSJKk0QaaxxHxK9H6r8uePYyezxKUs/zPK/ZVoBvBucpLyLfPYCj1iJ84R6pt+g36
tPEgQdb8SAXQLOOrT+ycA3BMY3o0GMC0Zd/rBDqDmWtXLFOIY2WSDdK1rKVB6nY7qv4HCQGbndWP
Y3FjoZS/ywHkukHqb6XedC6C1EM0/ZsYTzYeamhdRpF2CyfNrgFgsI0VvagCZ4LFku6QxzbsSXb8
JDXqYKIIiRZfDrpjPM5Y9jQmpa1zTaH2KxNMecwQzv/shtdKPJ//iVP9VAgulWeLzfG83koAWZVP
scNk2J37JxEY87BIFj67Zf4dlUvEpnEve0kpSKDhWNGOfQGjZ/wMiTrMdhWIE7tn2EHVzmssrDQ3
Bd66fWqAns9xfgS2VOO25aHtkiFzgnsopRfu1C11maBBNGm1hnNAsgFRVoWn9UyY4/OY0HoovrHB
7FI8/NzsdB2w7jAcP/NKhQZP7BqriPUpdStj7fACK/YnIX+ReGDPmFpgZRZrvXX2T3yjzG48O0QO
1/MURI5ok2ShZWH2hA1p75v9YNplgyhiJYAIPnk55G3QvjZ0YZ8rfdXx/5zL/kQiQzY7NztibMNa
U7vykjhCdpd1k8l2TMH7BP+EMIsDyLDyl/LMBJHceQBVuacrEeAixLzKmyBJhMEP5wnTggxLFEPR
dq4tBE+rPjGEMzeliATOaRpmanirWJPstj7ij4P8v94yq4kzPQ3iWQS/EGWp75C/X5JRErKbhpOM
s8h9SplFGf4cS4IYwMww9EORD/19elb79BOsciocuRYyv4Pa3FXkdZCylUvJJTSfJjepGtcGGySs
MRMKkS1uopvj+kwleZ6PQGFPiK6fgKtHNlEr2A7/vhAxlhC1So5KWDHUWv/CPJhB80VmghzkLoFT
e6wqV5Wesk/i2rpRUYbzgWU+g1BsCe+dp8raqybN8nVXceZDjYE+GqdGMtS3ZPhGbUEYNf7TXSgN
DrdAsoV1EDXGeaL7pJzFB7EZdJW+ULjN7p0KAUXVZHtfXS/LGzdxUegxI/d+eFfqnITO6NcKRIh9
hb60+qL2A12v6WCNQq84SAGPsjRViojW4Ix79APdJdNUMWXFN3xW5FYocHkeru7BQsznOBMOnB8S
JlKz7xVf7TzgKQijZFej6colG9Vxte2hEo8ZoBi6eDH16XVMZOlYuFbm8XZ+x3iLIT7hfNt61V/9
rdsOyWJj9ZBrwcM9Ui8Xk5RpEbeqD/JjSAi0CC0DY79vxfAdu7xm8FflYCVuMLju04TdFV1ffULa
ZOWNu9teu3LIjL8i1fqadnFtQdiLkdSBTY5q7pinE/+vUOdIbTzTz9Ab7XOWg/Va0KAzXE3RiQNK
2QeD0O6FcK7IbkHkvB3cM1dTyGOc/n20zdVYawBkNT0jrV1T4/XWmmj93RI8p2+UcmdA25GQZxcM
QVPPl1oN3wefmEFyNjt/6efiE2//nQjVz/MT1vq6s6Br1AvTEDdtCbH6vWEqWlDxHdyDRIoRi7Ab
LYA7w+8jhlCQn3dTZVWXa121I13VUd1m6uOsBOgmDal2ohGsucL0gSboqArS/mTzv//T01ZKaPhg
NlKSgZ2MFavv5p9W8XciGFu59S/aeQL+CvZiGyS/YCSbQq4vaY9pY236zvv7j2COFakiu4yQhnoe
V/ySKKBZZ+YIhXIbim7W5K7tZ/mtqrqAI+okFd7qnBwTTINxIeE4TzeKXA3mwm+F2fFufLqL5CRd
GEk/O21j1W9x0dKrtPEv4ZFxg4mKMfr4MtygdRe+WOBwtMjYP/fpqWAAwxgcJu+Pl+rLdoHfMxNL
nunODN86drVcRjlviVTdfigkKavwroX2Uapl+DQUdCjhptbVvvhhkyd362wOql83f5HnZw4ewblN
pfFd7uA4R+gZy0eMgebSKiy9mFhw47JCcMt6UGofQWay8uvt8pGhgkpeQ97RI0Ig3l2XbQc+N/0A
z96BzNQo3XV/EazBb/uxpmCf42R91RNXJDMQUpL0qdiWuBtJwRka0Z/isYXiV6eRAR8tq2YF69vM
zAsEXqQ+KBFjmd3D0eDWQYLw0+nkRD2wlPINDKQuU+fPzJOb/0iNI68unPKCtMzxP65eam55j6Bs
2Atn69DpK1QSYJnNvPESfiUGv0Kqr9f+Wt3TjCWzS7Hsiy5ddJJcdq6ZQeb8DKIffNzv4cO3BNP8
MBhWBzRSQY6kRG5WvcxYT2AuJbw4uvinfltPiP2kMqpWXQwo4BNCVacL3cXZQkR+7dJRe1XFmeyH
S2eFI2DRSNF3ufvRcPfwviSiVwqc/BNSAHV2ZaYtFeN2K+i+9m3qus4PE8aGMfB2V8n2Ylepftzc
XcGwHn1pLTtzzN8yf7eci023bYuZyr3PiS4913/7xcgQmcR9ScJkeJ7teuSFOnHI9PatqQ7wLUu2
pVTSlnXbNWWWKTwOykUs5Xs4uTciuSB1mM6zYhZWjChT3WmYGCDITcbJs1CuZ2nZhkobX94deKVQ
bjd2grEQoyKujao1/kzKTZ2LMKffbOW+UY+FhlwP5/cAglON9unpGe9BOUOxQhfEWkUTvRftoWT8
qnT6zychdI/hvDsZalLinMtGfiKwJNx/1EcM9nI2p97jBkyTgdCrdA26iCXQnptjUcsGPNgwrO1p
vucbVd5wpYhVwcYMeMH0EBfG/kSlXLQDFZF2GCwxVtU+vGCisf4PKekS//PQg+uouNalFhkB1pIp
CEEsAJGhzYgglI8nCnnMqYxiknaTbDQePY/L5QaPJQU01ANh87FMnMyUjpdnOymaTQokAg+yUanZ
pUktvbb0dt2PCThBncWU3IPoNnNstikfWSkW+89+WWZeEwyFtKHzAH0yfta3PfZyqDHr4FuWj1qT
sJaCxzP0XGG6SqhyhSTsWf24a3miMpaqY+M0+OWuY0w8LvVq982wAJXwtOiu1L43v7LqngHkxSWr
pA0oNLAtvOVfzFXspQlPcibuAoP2zTO5owEy2FaK9G1u28mMRrhSgRb4KO08jnHFlcGMYOm5mciG
fXz/h4Z3EjNUz1LScSZ6Ab3ZHJX6XUf8zkypQZOBp7FodzwkEIE028GKmiaSzHTgTmg/u5BFwFEE
/+OpnJb3mnzbr9P0mG5AODu8covO3OiXRR7b0fUrXcw35vHHEq2oRzWhtYT8a8ZatS9wzyVHQIWF
1JmDyUM+OO/vYRnXxhUtbaiFcDMb3IjheKJmSAU+45c4bFA4fGjLofz7jFj+X6Sz6bI7YAmloIjZ
b33JonYTyUymPQIZKH4Nw6V04mk/YeS6LMWrD76+dkq9rm+H1uNiMTYBFCOB+iYfKFTvASLuv2TM
oIryuIxxOh4bmKmsOi9byIp2IG+VnO0M81VRZdA5gchndf16XZoDpMq6+4w89RWfxFb7oleas2DM
z5gpQ+hagJKDNZBXNMeWBnRnIlgkN1Cp8EUw6JbYvcYOxlYVSYbI8eu2CerpHXLgn39rNZ+d01nl
RNwvEonSDKCa+3mp/IylsXOFJn9exJt2Cgl1lN15cqGNCNtgpkr9MueFERuCFofXCz+M2imR8dXs
0I7DdAa/CI9w5FMiFWSzfmPVGBMTfnLirBeqwCXOXrPfTgoCOiNFtGy0o0EuqpaNX6l+YBOJh6IP
EFWyHMIelC9erkbD56jaFwl5prIjc2t8mKkxfAYBN3qaEVPnrFrlDqwSPjRb6vwLfnL2NOkstgCl
5qXe6vi8sfcPmAPa5PF5xRUNEHgvkhgusNtXvH3Mv9xBFNCIxB4ITibeMvveAcgOlVZB/gJV8uph
xiDi7glpuUrqBZdrqF7jhfNyJ3vBTk7obdl1jUCuv/wDVYbBAL8PrwBG9rP9I3iRv/28Z9S7n3Y9
AWJK1LrDu+cndhQ82SLOX+h4bRGxfSImE2uGhGrAvlj5xxy+gZVxRyFXYvUxlXoerYZD8Qd1S/O3
YGqqNQKNf4irfvGlPvdgSl1vWFIC3GwVaO8F0+SquRNF0onpTtcjd70VY4jWg4hwvbm58fdhPm/w
lJO/6ZfpZnlcch+G4nypiyjrPpaHoWoseesmHWvCGl6455oY+U/VtTmb25djHu+Vr9en9fu0VhWH
lt2S5EYfSB47RQqwzTaKGBuVkrQ7KGPR9+6JHlMnZiro7qjv2rUU8TFWG0qgzqE/eLi4nvSkzFD0
R/LqKpmoxr0QfBUCzqab5o5+8f2DcFpLL3RqNYwaHOBbpCaJ+Hr1LMIX9AtQ6M0bhU4aKFX++t/5
SSl7S61pI8WP93KaV5crPcjTkXKU3aIQ/6cYOLjcJpJnCRyzpKidNXLVPnWZ6AjFxlPN9eLb4HOy
Kh5Jj0UigrBVE6pTODYA1QKg+bB0uPosyIGnAhtccMDLPRrcuJSWA++ozgHZgc4sXFx2MRlW/yP5
EdfMJ7zPUjVvCvcXgDYQgzePqxPN5fkN5fnpOhnVRbb6XtecIfbg1uTsZvq5TTv+bSPFjrHc/OVl
O1HgkUceUXaMmu0zhffNIDqRTLQOG8Y7VyQOOZkQJwNhtcOuGlGS+28AL3wEHhk0fLtn6IoScwgY
KNDWtoaLCC/4XAQarc+s0qg2BL/dWx1mDh4B7q2FVU1tRhcCzwl3yB/Oadcn78zCEMX7LzyiciB4
deXtC3GcIbU+zRbB6qhTLcrLC4xYbYr35gOA1ZP46o5ZtAlWhiFgyhXPQvs/cVl9cjQ8vMXLDxfS
wiajlzffJNLB9NbWhYBCiKgBGz+dEMG7ZbxdL2hXBq1eGkgGDwobAu3XjTZXx/jKfAMxYOi3YJYV
2HVXEgqC8UJMR2p/3I+SUvt1MAW3mo/xlg9JWZg/FOXltNyfRJlga6/MYBQXc7JXsqlHYM+PVGoU
6MmRUoHgX1f5DtV79VnprbYqNw/XUGX6TGzgUY2AeEOSYzU9qjVcCflgvygyZncHB8M48cWsQb4t
jkf5LQkaPuv8BJQPqdFbfBm+P9UObNdxwUcXqd+VVHCSiM8iJ+XMYlogoe5DroJGsC7AhzYSS/t0
585F0TsuewB5WU8XJWJIcjbMWmiGfyX5MKdQt+vO8sIxLEfmbKv1DiBs4DMqHvWtETJJ9JcLSgKj
sp7UnPQkbRt6ew+DycHBW7pxC7ao7BAaoQmINE8mVfYdf5T7Ufk0XS4Thty3y39t3zhyC539scaF
DGhBC0OMtFKrpY5eCI/OtxTNIHwn+ei4i9DUF74KpP0/urqJfr4+HtTfVKx0y+0ULpU0uDnjohkC
YtolSlEQTn6xYrmo9Y7bTkDVWtxiXpYFfvO+L9rN72rDwMzwYETYdPZYWMA4IGx3lIF4fYSueq9Y
9zHmcYFo0Hlb+EjbM6YNeISsLEimdoR/9jQhSZJJhT3vx91PI1639VMkdf00wD9ZZkqZ4MEJOUNS
DooqgtSc3D/CRPzV5ussbuk8nvwDShxgCGx3ksyA6uUk8r2Elpwj6vyNVa67ltO6w8aKwrhqHSLh
3xVCAQgl1J4G3y7UFW0P6xtiQL6Fb1pmpkCwvp/Jr84a/IXwa+m1sxuV+GI2oIX1w+mLpJoM9158
+RwJgZ8xg2aF7Ty+6iygtgKCQQ0ITYfg0fq63VpsVytS9cqE2lDyTx5uGJ/di/Jqp7+ZXpe651Xb
ILAoNfDLDtl18/nMDWuDmxKqc3dXgfmRGH7zlED1yqEvHYBv6y04EE87mdKK8Zswv5ISqv9/HOTd
EvzLaY0x/0C97dpbhShZqELldcOoLRd4hg8BYiakCGnWZtOGo0MAETOmEt1Hq1eZ+h+M9Ny+Hn5J
Q16EMbtCbGcJ3TG67kGANmI/cnJ4ME0EIaPn2zN1EwHxe+24XNqJ/3qQRP17aK3+XCF1ImQdZCx1
CvWX6VmVuRW+d5RRju7kuGHpRifVGMjvJCJAr9ezozgbDSODSOKhZRRC0DBInGIBZw8jsUFaY3ux
PbXcaQP+jC4bdtWSJ590jW65LT4+59Vzc8la1hqJWvthx+wFJOf+Uv7u0IFzNBwYk5cuOJfbzWB+
DZ59O2EX3s1zW0lMmPnPPBvYLXijOA2j+BdgZtIlWtBCmwC42oYMQYlIMKH1rO+NKgZpYvFJmlcP
B87yAinP04OGzq0mOGkDQ46nUKvFqagtkzSeqoBSMCU61txv634UyXpluK/kTjYNPTjaIoPGZeZ9
a5HRWsDTwztpkEZoFOeXsTbYZyqpI248lR7BGARBVrCsvRXI3z6IklYizAai+K61IJYtlOakk6sh
Yqv9D/mZl6IGE7Mq2N1We0saYBL0wUs+f3jdxM5CZwL0blJrSbPdWMwLe+HbTcsvA0Lkeap+9DQ8
dLHFFcM+uirUjYATJxj9Df/eZoriUtOvHusgd/2kz/YG8+6iJkNR6+KPSGXn8JOvdt3el//H8dyn
ZCwlr6mjdNJWVFSTJ6q5wO6RwCT9bJhXT6tFDa633SFx8kNQ68dOOzTjFvBf7uP7zOL7Cy67eqKG
PGVJe//xteEEsc7FSULT5SsP9+q+stC8PGBWiqlOs6/bYnItknUMs8z4LqlB48j3nwriKUXKLwhs
Kih4f4ZN6mKXdpTfZukys6+BhUPZttX/JLIFWzmvH1QACBpUhfV1twE8GwR9T2HtnG9Gsv8EsYcJ
s4IW2XvBSCXhxT026VMUrkpOzPVpdnQzIThDqS/9FRLZ2coZGeZt+wBhc84SVt2S9wX/9uXacBU7
axUvXFKU+457saiJRQxnILgfHRHrY33zTUnoLxmuOrDZUaaeorVLxQLl0bYFIosY0ChfQAg/HF/M
x+hM/PYGjPKgqV7AwVv3ZswR1EYJw9h0BpjOeYg26y4DEPwfuRhyr6XvLv5Bj6sz8F7cTKX+XYLJ
n5PaUyG/KmPLIs8r39w6uphsNJDCa0JaKjTBeXM1GSvHhSycODerN/TM7FypI+8lhhuerXL5BYKm
/d+vJD9wHowKDB7GOLifPv6UXNWMY+FDRWdJ6CfwD2K3aW4PkBO+kIJ25PqmwhYOQX1q6CkE/p8e
IduUWRWAT5S3GC0pAX2r5zvSpWcULuVz98aCeuNtSXWbWZFgoJEu3VRigzrl5NUXXrCZTT2gCosW
QdOih94yMryj2ISV8hb1s2MOBZlSURgkI3zUQ4zG7LNPvrhuePs9vtFuxF5G8DVsT8WeViHPME+6
Uc9mR1tBN3mPwtMErGSNqCV7Ey8gu/hNPlmx7xM587K+XOF4ajRDA6jxEOq1XJcacaAvkiDq6Cfc
r7EarNL7BfE87w1j8tT4ST+RyfBhgrPud635KUdnF3cZErRcDHrPg67yMUfcRQpPGOgtGbzz67zy
PFEuFAKtkmUe7WM60ESJdDBO1XRDhlDTf9G7xLVtx8P4WMAVIvLM4MIkXURFLARgD+tufZsiu6Fe
OXblSqbpew5/k2tMZofxwmL2/nKfrUAW6YYib8qLo3KmJcSuoPcseP7KKIB8fxJIIYgJKSIQZcXO
mF2zehLy/BaOMrMppAPZVH8mZJmAmfBAzkrl9iMXwwe4/P6js0EPFJRtl88aX8dZH76IIEB+TLDH
M3VE1QHIwDs+iKSvTV+l1t5jsY6h1orrTUAK/o9MAdaUaReAmvirhi5GikWyKct/+nuvZ+IsJrqM
bEyL3+bvGq9zqbGxrFaK5txG0tTePTnJBdbEsyxdFlWY9ksvDR05tv+YvOrQf6LUdJc2O23HlLeE
SDuLRnmjylQb6+GL59Wa8RKzb+Nr3qDjE2W4g5jqG2tVTaVa4daDZYusWYPlWKjXPy+ZAcIxgu3t
Q57YajJP/Dy40TDghS1Wp8TsDuqLJLH4MFJskMahlQzASQ+EDH1cFgHMGI32NdlziiKOYgjL1AjB
KP7Q2bYSWbpuaEB9AVXAk5puAYnTxuxPyIBL+Cn7J3OkNZaYnBBNM5loxxkCdMU3v2rsWj7Fkvgw
uL48lWRcADDBwVIs7Ln1FDAKGO9lTKtRdE2Xob+nnvney407FCicybj2+LBg0tl2dbH+5jXwbGeR
8TN1G0Dez0eIWBSsVg+IuMIzCC+6U1zJ8t9YSHOO+1bhXRzviwrckCsCPt4HxalqV2GquTUbhM5c
Gn32Lt6c0G2F/P9ONnNZVQPlMGcROm/l7CTHwpLP5b1VZ3OsViO9hPFRwAdU7YDw6XtS8cOof0uA
gXJgN++2blrvoAyNs5OBIIwIKAJj/wcU5ygF6rkRqmXIVhCeNwbz+S5GSMcjKuxCogaYCFCggPL/
2/lNiSqrT7gk+hdnOOiY54ujC5nRgKf2VAyLNVdR5HTxj2s1GQzcMCAHQgZS9Sydc+7KJ291lgR4
557mqJY1Q6qKE7+gvFJC++/ENzQYFvhrbGr2RW0XicbIYpCkkNH8GU0Y7SHLEM0hfytfAN30L5am
f9hZ5Q6+Db57VLPpn6sv078v7zsVuvh1O7T/eUyXJ6n4wzVuUQ1QO2bWpNrI08kDcxd56Fnt/Xb0
FPDV3fdiNQ7RvFEpnutidj2mJLJ1jL40bk1CCjPZxEGTfYimK6Hxvc4LMdb+ogWzcpJbgVJEuv32
YtalPRZooRDnlZb95HWSye/uVmUvyfrW4KWLAVlktN9yALJEx7eILjDRoI/sV4v5OtepBgoS7ChB
eyBGE2xaIz1MWSDF6E83OQchUh5KnzxP7y1mkZks11LDW99mzCj09c0q2MzZt/LR5byLq4bpEchA
8S3twgeuzYJwqC/M1yWm/FQCmvVOGuHlqzBkHiBD+V3qcg9pxvPTBVYFFv36HUnXPQVU8TzuVWQW
SgDHd1c8G7oyzycGVID04cC8jp63tKJTHslV7Oo2WnP8axMrUQauAjmEe5whqYcENDr8TJ62S3nb
qAv8+C6hzPNw5KUfDs7BH199N6XsB/NYg6e+rqGaVkcmEeC0I/2zgjcqny4FyGxD208ba6EzU+6n
JPqJOwptOrB9yT0BlgiR9VllQAq0BBkGnrNnx8mRRCqH5L2YN+LR5G0z2t4yYl449KIPSXUadTTX
7ooErExyJGl4B/vCYsbMUAGX8R7c0p1lN1EzGAPsV0x/8wmAtBe+DQYSCxrU2uAL4fsg416HHJTZ
r4UmBUfNqboX97f1c/BWvmfOC9OfRZqGzXXEhXYPZAFpLwA/qT3dLiT3rgBVhBoWRqxN38/vr5gy
cZuqvjepd+1e4a/t1NNesG03a+ozdR1u9HEaXVQO92IUcN0GwCF1FRUAd1++KDBpnzHFqMDq30ui
yITGD3b1BHXx/AB1SWD0VMyG+JavlB05Kd8j/SZsXOwPZiPEoZ7XPzp3k4BcOLvWxJm65cUglQnQ
xu33TbftAoNKSBbhJgSmWSRb+tyi79LSDMl8nDBRhsfrltbSHhf3j4EdaFK/937sfyzCJUB6JXYS
/Xfmgi6x1LiJXUmy2MlLyQkoRZiyg5lrwlZdTECi9cMqWoelh6N4LLazj//c6imT+C83oxtwvwQa
ukun2qpIeAnjhfuV9TpQYse3m4tjAguKGia0MoBVUbsH18v98QZEp3FD8RcxbDW92j42p2n6bW1e
SB2N4nHdMlxvCIXmxLgpiH3fSIw/jFvZEewEBBoDJIZQENKCIYkjjAGAc8yLkqZewt1Z9PEifNoO
8sqYmaQgyEYZxmJqb08b1A0Lw+yJpSPPLnUmAwF6UlJPkJG+AqJUyV7MkO3QQZyF3M/WylCnSDCR
EYWcbF4pUCKoIu9h8+1C9vlRwuDDWa8MnoGbsw1V914KVX8+M5hLo6l7cMmkQjR7APakM+IsADRE
MO5zdj/DGqTqKoW8knkI0Mz3h8ifMvXLyZtwdtH46o23gtRUj58Mxamy1bSWgnZm642bkEaRHyOf
vddw52jYXFLIfpGQOmK6dXBNb4gSUZ2mNvoHSmEab1lCsBDg10/DM75gKO7sz0yvBBb2OhFLS6p0
ei6eVyOe8/cqaquUZOR7fZSAmi3Te4udesN36ynztmopqLDPolEdPLEk+CIxVSdC4orusa2isYWh
r5gkL3UStxA6rKfCaGmXyoW7yV4UjsC8K3+AFszC3fg2PFTKpS+NXvxruAJGCygkPWNysseIWjlt
SHMa8wRh8eEzw6z0CksDhhy+UnDD2A6PX/4zMufHtQR7kYnn16ml7RIdqwVrFFeHqH/EcMEXa97l
Iuh+nn+JVG0eiGPFqGbCEtlcvg5hZ+D5nHwPniI2sRbhfAQnzV4kvyelq14ihsn4dbFq4U8uGXFd
mQtNOtnNnmx4xKv9r3h6rWy3Z2R4KGefVAx+UthJn+i4V93DDq7iGubECSfYiEyr1x5OYjlFLJqS
QAiVobYBHhYbkJsSPa0+Sz2v1pKIRg0yqkz5HHMcL1JxYnxDu/Cour6FvEelmOWZc5SYoU1UfhQU
04JaWVvAu/tDTiWh59PGt2b55RM0r5mLT72nIkRQjX6i+l5zUOtM65CmMO4X+s1z71ucUGHiwUii
/urr+2KtnndZsPnnif2GM5lSzlT4ffaeW+gW0WyuCwG/2crKWD35FAHfhiN0iqKBxdBrLLNbEMw3
oacOKwDotKGP3RIKwd+6DudBy8wiRdUq6z2FtHNAghgre4zhqUr6iLpRucKiKtO/jUTpAGnqoKci
ytBL+VvAqaVv0vKrZdUAzpyC5FKAzehR9jbvN+301GBKqhZ/tn/lz3f9ehgsBW9j6FbdKP1aDPVS
7upzD+6VUqY4I5g/Fc8ewh+Zzw8aMFFOrmkRjv+MHpErVA/gP5zW06JbKAwfeHshPA3IuzQw/NsI
kQsErH8SyUlNoXX0MZ+DHl2xK955oW+jw1aS9y6WoYALffoBRJTSPfA1Qe4rUuscYRM08QZr/UNX
etmbARIqP9oszDV6jdib1bwdME4MhO5+BHOSXuCSQOGAGqZmFvZht1/yClX0bEYWg7Sv6wdpfQ44
wkHMzvNFrs+/AlwPiKmHzZUfvrAUEAfKJuYh0MvUt0/KxSRLFMviMi0MwTj72j1mv4tMQVXkDbLQ
v8m//aG21cSgQiqiRpVb1sgm9Z0XYzZm8vX94fl8JYKoUBLNkY0JyGcVmoHRah2c4yVhi7gtKzoV
HbtameyC8WCw8xM7LjL/5OoFpJ7YArYIMLCOBt89WW0a89GvzM9aB2OGC6lSUeh4E2plKLheMgyq
RV0+TSGRXxIc0reXoWXFkHHnXpvRuF7q1ukHlO/OCaC3TO/l5YZkkaR3qZ8MwBOSa+Nkc6GqsJlj
7Xh+KIRS8UiWz2oXeU+IphM8nQhJttRo9sKSk2oZhS4LJJtAJ+qZfdYMMEWdPLwCgRxQyGDQUKs7
/Yhlnyyf0RGvdr+oOo4DIDU4UDWmvWjcbTrAR7lBl8jTyl80ZK9ElI+5beKkhCE4zVzZhKsLqI27
WA6thUKfLiYBvPfeqCFRtTqAUEm2y3prbW2EDHLF2b6C5DA1h3rQQXru3vaawjm362bLH6k8Qefd
12Y9FX9Tg23tdxP+U8+Xd/RB1Iah98D5qByW7K1BO76mXIGFN0ykIULc1s5GDAlTarZgeseh9Kqj
iTDwe1U7mObv6/gixO4XBmiYF0kx17yuwkCYbyW7ikbpBlHEqLLPsPNMa+m7XJqBKxw5+E+/Rpy3
A502mjwNuuVPNh1JQF0kXsw91hPvcV9u/PtI0z8c42TcO83rwPIwzFgf2NNCe9kKUem9g06BBTZV
YWKhU4Zkpr5zTPtD2dv2tF2xNCbZG94z0WA2SiozM3N4V+p01ElsxhnoJC3PLh4CBPX2UeX0GuGY
EalmK/I7xSPAqgnOBrxFy24wjkfXE4u5cvzDc1shjo666utR1SSp7Cpkriry1BcVDDcydzKPqI6P
6SFlG/0UVyS1vLEdM6HjjJorahVIU1Soa57l1kCRkTiDA5QkCwWZGwNYfW/L4ajZM3EiFLKelTPu
YY1WlBkC7sWeBxh436CBIw+eVob2B1imlhY2hQXCPwO6RGu5XE/geIoiaDXpRSgBkoAjMdXxn8uY
DmsdTaz/H53QIuzPYJdrRC5PiOtEFftYsNUEz4e8RIkAz8ev3729ELsIcR2QBMYD3rM3Ab51X7JM
I1eSbQHNEmxCgpJ2HET3yLHWZItkteJsJmhgytxuEUzFvBTMPvg0ONFysJDvrj0+3obj1qSIK2QR
iFLAvf3lyqu8MRAsepobWCV+m8mI6VG+Uxr7KWKbO/rhVqo4WGbjMYZTk/LbGO7dm+V9ybt7Elul
z8oQHbS1oDH/BU2ozyEcpZJMoZoVf9iChJP/cBGssf9FNPFs6ylI7aeTMUa2RhVOlxjYdT/Y1vsI
GGQRIr6FYfsRaaqfjL4mpH/znmX+PeHONVNKKEaWPP5kBhlGbox6lMR1B9Pgnrew09+glGV6sHRv
0lRq1fqZVQZAcHjaJMgUhXBU52/NbgNh47s/vo29gRslwjeW6vZresESHSgAWpoHtYcecLE2PBsy
7xRX7JwfyFSf7PPy5cHxp+/mASwQA+KO0EHOENbzkT6AwBM3L7M0QnZ2o+ruVust2+LZNHuODikt
uDyS0c9Nu5UUttlwm+mM51ES2rmFnd+t3PDjAfeBkLPq6pfvAuMhlMSRUNivBsMLD8FnVJBU4lCD
Sz2t4Ecr7cTXEQpCxrwKhPqsF7dplNKdZKhgI4cVu0mCpIlbx8YjlPA990HMvwljGcdReteMx7zf
/0q4GOwEscBqmGsOjqZ1/8yfuXdn1l8Ebl4oraZxJwAiIhW2aYE0gwTzd/h/sVe7CUY8YbgUCRot
zCerQwIQ34qHB01KdYpJ8Q1fM6vshHYqfeoTUCtPUYYKeZmeEu0ZlISr5xVYeGRSpi8EEN404BJT
MKlgX1rYh7lksLy5+SAUCoBGpZqbxTjtR1NrMdGc34PTQBvum6h3Vi6wG0yn0TqPmvrWu4D7uxwH
QMsrPFLd+phqip1V07aRBUCuM+M96e1UU+h2FraGC8jjrfYMKVZ7h6MKyvKKIQ7GDrzeokH9P7lC
PXd8tQvA7hN5PiW7lWXxA2alKvkqyucu2BtlDETrH+0nIJnxRXMTEXZmdhIjI6ZG/XnAmJRQVBHr
hGXy6b+e1V5BeKDrp2lJ8yYwqM4ZSIKFzioefdaqmwZPni3CcIRID6BiEYc/y6YvM3qaLt8DaYkd
glIDnXKPZaZKfaQW38t/5aEhAbVnCimXDLL7zHui02YfMAE9/agZ2i8Re5BWtliDTUnqyFSqTk8n
7aD6xo0PXNIE5agsl5bmVJfwtAzMCDzDxgOhiP7FC1Bepz2JhLDf0TdJDGncYSV0vQIn0vV4t+wR
aao3tRN+ukoDamXJs7BnR+kh0tq/GaomVSrTVRslCOATwfPYIUogQ+r4EmQvJFVyd9VXRLXczD8/
ijeKuP8lGV7y4nLNE0poExA8xlxG2Wa7hbfi2YU5x26jAgQG7SWEe2H3Q19xvjI5N1wQgdw485zA
8rhic0+ejo4drcRyvPDYhCLXEbNZzBjAtDsPviHlMxwHgI+5lJ/mhPaWzXEchCbHgnM85aZwrVto
y/gnhWujDDOLV1XOyB7tJuZfRnscdG6isVWehdurz/IR/6pQ/WkI0S98g+ytFBXulxO2xjcCOj5v
eX7R5BQKKwGAftS9RpzmDUJ+QFeWzspPvNSSw4S4SyOL8aMMOJ+OQu4PM2QIAaGz13hIdde/ypyT
BpngoLiqZ+9HYq6jbKbk70II598URAwT9aWSVnYfHfUjtO2wwkDbMjy9aIxNJpPaYoI0VjCORO0J
m1a+3XvkUKFDs3oMvtQ4Rl3JdW5Ozo8LfbPzGGke7TCRS1lejNUaV0AZdXv7WlmAlpK1/OYk1EBm
V/ZnQ3FHUvkgJa0BPrzVTh90MgUZIlZp7J4019POjIf/AbEc/EGuY6nq5xkNAXzacx9TMuTyKmXG
8wuVo6vJp+79Zr/XTL2/I2QWkLB6x8rfM4N/MGwdUyST+OUsp42bjFdj50i2KjM9aCyk7J4e3U24
f7pMqYIrdW2pT8Dg5fIxXEspYuHWZpvIB7XhNFT0szqZgu5WbUkn78MUrF2rxL5opiYm1c77G2UA
p1YJxJ0zzUgh9YWTsKc42MDh9sGBJ17xTEjgimyp4HsY5RI+PL8wraL+G08TieTKCCumNuNm00xH
x5NO+LFmvAfpZfeYGfKZSRh9d2ZThKRDMlbdQX5GpIKa4/CdHWRtlDmLas2DcKklsiTrk3v0utG2
Qq3HSkV3V47zATVvvkiCWlAWcPZ0ZjGHQ/FG7lu354JB1/CV2hSboNMtfIlXUI3D6DmAajpTDArL
3MgKnjfVcAgLSdwA26F290bLlFQDEibPMflWAt6KqhgUiBMrwIC/8XEDwIElPuTeD0jxpQp2v6Ms
EKlL6QRUMm+1hFKKoL3iubOSa087fMznb/epitTQ2FFdlaLPPpXha8MIu0aYIj/S7nBVK9oT2eiP
KV6+jwaaklg3Oi5S/mXztK5et9mWp0+wHK577hmVG4pHlP5e0DMAUJPXe8Pb7CDForLYZ1uHffEb
xDXYXVmWFiQD+Ykefq40O3hHoNwe0r9ojZAsuVAuUx8vLkRILKOBhuMzLskD8brMG0EIdQhFyyCC
/6PPYw9aoHXmnKeMTtvq8sMry+D9lrlRoxCI0lJ4vCrjlGmBgNXOJggLpb6j8/RLWp/91folfjJY
/iD4woxxb1nOAUZa2dHCmUk4RsvuZcZ3d5Gb8Tck406+6exGZ1Y8WgwmpyxvzWCjuL8zikenqT+I
MNOJyqNTsw81valxjNhSc1P/TU4+u7TrXkKvxTalbYP0dP6YNAvkhu9+XiAP3pQXlOXF+1yPjIZg
BtZHzyraUMtqsOmnbw0PZyDBWOZM1OijgVsm3jWB8txKIPuXWZLoZI1DswDfgN1DHggvnZN6x8Ru
2AlCHors/ogaDdWP2oftHlUqbXDE0BmGd40SRcbA5H36szqo3A1JEfcbsSuvbFAgZHIk1RC4Oeah
KK3E5jEceZxjtrzmbiDkdosQHQ08J2OD6gMMxchWXlswONN3ZQGhqjaZEkcT7rk6emzmNAc+Le9v
d3B1WJ2NtoSqu7lA6NOt0dhBlF2y+6NAiQzrnjZcMglr+cnOAgnF5M29bA6zwfWBnJmbehECaz+h
Z3I89xVoj5rDrYm77JmVgL821BrRr//pNPk3wACYQU2v2O8nrY3AepcUdIqrl+QOc+zZQxGbdwYV
jVOVbEpFoSnjrA6y5hx2I844iR62azwFkxMkeUX8JUVTzNTARhGg7qkzzYp9Ox1owuYUHUdT8YnX
44sLnaM5un0bQe7yHParVmy9tnYpzTNZGs/18d/ueipmDm2TIsAEO4ujdqv7rjCEdZJr1qDyYAti
jROkPMjA4D+X8e8ITDOaO5ytp3xFciDzIJ0gDOYFz0zCdlXTX2R91zsBMhelSi9wAU4/tIBvwTD0
iVl3M4RKUTo1+/C59Qylibs4wHk6lvL0QfL/Via0rwNwEOATciROQAqNUWkX9hlyl/vpjYKeRKkK
oHRKDhbKFMsyecerigvr/+EFDOYM65Ru21WWcb10aOsyzntAbN1Xiu6f5zIKav2Q/GLGHuRel8tL
RORTReOG2gOlFv3jOh+XfLR512QxKvzreiReRMRF/NiR5mTEG7vkYHwz9TSb+rh99fbBboXaKkkN
JWbjQ99kzTXuUsoYLHhSGEsoxIg4paF46IfRfU5j2JVSkgzjhQEnYKQIkydXp7RqlNczRESyiEf/
gK3XtOBrbPDdOiG7MISkCxhXjMLK/pbGXeanZreFw+8KAR3hjeMyUeFpPxy9ZptgwySKtkc6Vd6Z
eLRPq4MrwHLT+SEb5To+TqhNWbcPTPgOn44zpZ10WSF5aXxZL7x+4DfSd6diFms7e02PJbZ34obZ
W8/rLZB9+fNqqFtPN+QSTVEv0lZvEDOJ0fxU90dxpsmnOhRIbN13XCioRHHn3Ki3zywQ/E4WSR/7
98CNx0OWwcHRqRYZU4uSM3Z414Irm0wuh0zobagQ1ggzdc8JGX2nv6Pftwe6AFVKKSqK/iE6Kdkg
dxeI1xxQUX2JPT/+HJYq2Cy7xhnhsecKnwU19VaU/SZVBNI/3g0v5EmBAecbj4PGCtP2A/xdBP8M
VqkeVA01SUp9AA6ImjFLZplw8/N3hIkn3xrIJ87beMn4WHdY8LHFAX0y5riiUu5gZaVOpWosKAop
X6Vyxfkt32jZYKYYVrmtCK3OKfGSzz2195wsUJxcPiGEE1N6O/YQG4xy5b5MUI8z5uYHa/2FAR8L
ozzNiRSEUeCbH0vRsXiwIqPaF9KiCifGvbBD28WIAfFofTjyfidgbRC+SsSc6GF0dYnG1kgp5DwM
9iSHw2Tve/5NUjV8byhYsGW8lNUbCLlF2TUcV1fkWPdil4VUAefv5opibcyqyzZ3LK7D76khE44x
qiuFrRigFJuYqsAHjSis3YWtau4vUPYyOFq9VABsxhOLsEarZz95+CYCuzADV6iKqHYUZlzS9Y94
czQ/alLn8QIMAdr45xH7oVkMfeDadW4vYUhBYXI7hA1ycyzX8RaQWxnNKJeuXXXATygXILP0Tthv
g22DC9uxwmI5/RhZojltMUsdQddC3yQ+eOl4RISJg3ZPpPpu8fLO2ZP4VUitqiwVUP52MkvuyrF1
DcHRGIrPpNK47GKNquK6yazu9NlyI9mZkQ01nwqI2QU0rSz+nqcb9J/cEztdENXEQY8REfa5rC4E
Gwbp8dIXWbg07F+gITRh4WnuGfcf03fRniWaXQdhPRwmAnpwpvGdg7LPY/xbQFjQgV4W0nCgEMch
2Ym58gKMNw3IXwejrMY8Yab6GR0bNH+i0PaFafe6fWIVh86F4eTFxA5cJSSS6VKyNT4BNlW0dfXO
Q9ThVJWOt14e1zI70rCKvoZ1Za/QFczxjpqqJ+e03YaNAwnWRC1LSLIUES8MyQdpHiwoLOsW2ykP
Aqgp67FPEYiUk1Fc7fK0UZcNzjVKpN1B1LqIjFzaY3lgbjTI+SdoRW4f/rwMFo8yYFaG4t1jzLYq
70JqcWz6w7eIv2nKd3UmwCLzLDt/mDRLM8W3V6MZG6nSPRiVIsuJnGLV4YR94fmp176oCz9F2cCO
tB8nHL7XWO4DBzSnC7xPna3PzLdoVcd8QIcVYvWDLIP2IpwxiLrnAozd1PSXkMAyyeUlhFVy0Enm
Wt+2felhbcm8A1Xb+WHuMdRPsNTthoKiwMQ11698Hf65lRyE5COU2AoAerqATUkMZorHrt9EUAF6
F91jjaAY2DCtjCREAGgsU7vGVUhZfMKur2gcpWu8ILnTl3scHMSyzbAIt3+0+Bokq/ZmKdBGm8nv
/BLc653Q7qEeS/KdBS962ke+CjJmDLLoBXQfyJOn4KThvOIEZ+OgsX27HL9aoYOwyM6cIqMWD+Ci
BnsIGvNxWkwhkJ86hO6RMlUrJxfpl+Zs8VT2K50FZ5CPPA0lUNE3QuXMBFYFwa6PT1V7hRlA+2KK
I+OlQgyL/9m8tpK/LK6ged1fg0A/rBZpk5kvMRGOHo3ioQ8Ia1/TD1m5vyyjTAH7puTyUN2kRrSh
2ReOU7sriHIyH0k1oo0SIa8dhBgnNpMBcrQFAlw9ORABhFs13rJa/5pycyOwuWxvw43Q6NwqUNYX
jWFAV7Y8/cM9BoM3pn0YtNx2c1jPXC0kVMuULx+prLDHA27Y270w4rAs0IOuMzokNxcZanJBH1Oc
opoxPa278U16nwlySewJ557MAjPenF5vEgHS72A5nVqCKCQdIRmagDrplInURnZRDB6YiFrPy0vP
Svn5AyupbkI42lkLd50YyTyWzvFinn0hlktsjREl+V2Kwmsy6wJGULSWX8vuoIw3AbzKJpJ5B5CH
taxEzwKffRoua/S7Ka5lZo03GuI26ONz4VNASloyJYhEB1M7LSP8rdbV9lHEKS5z+VpJyO68SD0h
j3+tcHfdo5t7J0p8Ty8rWpjevRwbGGTO4isJZobZlNw44yg/cYWk/gSORf9kXNn+tWPZU8WETVeE
u+ku9EHCfW9zizL18bVl1QKTWXSZ2iYqCVI7IgapcrhIK+Q6v9Hh787a+9IU9YUDHeqY2BKNvWDU
7WRmRHMaNfBwu0s97fDQACKH0JBT84GF6eBlbXYO9kldRPiPHxjATDtAeBQPLEpe1H2lAYMZhuIl
YzyoB3wstmhX+URdMBZzJIS03SA3RUVGIIqYOvFPg/q5Y9aHKaoG+rvwaXcm90OR/OsPh42ynWq/
OZqVu9h02Y+P7lgdjbT8B0PnTiyLP12f0yuzrKXVFzEO+ZGkPqi5igdr15EOsQp63Yj79ua8xF5g
oDetnFVrbaBcaEYztGIo1QzxGwE88nMrRzK2i7hmkbeumJT2vf9rA6U5b1s7oxYrpEW7akx9QfvF
X9+WOu0ycchAkPEXANdNEofZaNJaQp+fbCvEos+/ptHAopvBXBnkMAm5dAbRzCxB1HkB4I7u6aGM
Rph4WxtS05lbrMjaZOVudf6xYl8jdHHS5L6jlGkW2bPDZfLgmJMemuhAWXUaAc+petIWeCQ/Wu5d
4ajWUDZOAXAAVt+WmsnSerKGG+wK+CwpTIZ47gIZDJd4JhgJSpfruEcUJkWIbmbSN/NOkuBKt4VP
CaNw3O4twJm6kyFx7CiSldXqHGer6WW4Jx2jKRCC9yPhLY3YD8UHSSXNHx76T3p2z96GWG1G5QBD
DmSbJHLaE7DWX6V2ifkrKukEYjglSjQ/77yvsCNyoS/om+NRQkpj6sTZqsbY6rYxUbrjao4yLcxw
FkoWQh8/ujErSF7iq6V+UdhMRQAZJ6VHpiBwC4k9ZDj1AnoSNcKcLt1D+TWk6KjCc4xeReaGmfNj
UTyGl4u80d31Q2/PtwSXmt/Gq233nIvS2iuwUgx2kPQKTAdpnRUMr4SPMua92ZlpkQAeqmNX0w4N
PCXUKeG9aPpsHmUFiekkUhLID1LHpxJYR2b2vyNLoIvVAYH+LhHOiI0Wogo/x/V1jQjytYkPWgeY
V0gI5fq3kAC2AvPTUpMPOhEZJOreTED6lEiPOieqXz2e5jpb4nMu07syWNWpvKJeKgzy8GpUsUG7
tBB7AwcF1OyljXVXdpWFZ0waw1VxrC8ornAzv+Tj+0iwNgKIJUmwIdtuargzw0qO2qnncGsQu8x0
X3pfm4F8ab5eAGT9Lck4qVvK5WfXAkRGnunSRAhUNI0dW1uS7DyaY0TSTJJe/wr7t2PiQUfplDFB
SkiWJts7+bsl3QiHmHyG5VbhuPbGUF3CHELRrIKcY6wWAC3rMOmPzInN8w/tjw5vxsQc63HzH2qC
FEUBqapvwo9C5dCdZP1uJnDytSkU6liV0QxY9zElWf02aqBEeJL0ClvxBFasMGC1Wl2xCxlBJX+x
eA/HxNKtirzpISac9z1uxbDrGNSXbbqt5I4iqDfJxa7Tg9gWOPxamO8biRjnQr/ZYoO3hHGfb6Lk
dBgYjRhtf3wwKwz1B21cIWhP6XcfTN7l7i7OybSUz7A7UlsbYSmt+4ZUTzU1ca2KeNBqiC61NiW9
ZSkMUU84kkqmY4XPjy7mYx3ZMAxOiRrsezMI3uprRNFkLtvrA4PbJlxRaG5WfXH2iQqp/Yk/ZJUl
i3O5513X9q2FuG6nCNgJ2dRfMC6RUk8J5VJrwbnDrPROO/Nh8sStSqmh+2oweBqB75LGpjZBkLZo
1T0Dty3iIvuTI2PTXFQMsiGd/ZNaqxFN+D1VxptSFFSazoMrdE7GK/Y8ZMYzYlgmCu0Fy1MM3FT9
8YujAMalqGMaVjVajn6LFHkj6FEFC8l5+eNomnbKT1vTWI4lFWm5GGg8TnguV/sFkNq7xyC3q7mz
bmIdv/3uCczsH97megWolIJtFOmW7BZMNf4n5t1CKDdAtwajOIWOvMJ7H4sB149ZgYgobKa1w9E0
r76Uw/Y4Mx2LNWzZ+r/OxkoSDs6S4K3YFApbJnqiK3fDqyXPL6/ev5BdQEBFB3XD7vxUMYlqXCYy
CNRyo118t4hjk21AQRvmBjKXsjK19QILy1W26+1po87G6aODpaM9Vl1JfJmIrPVTIPQRJ9SOeQ02
BG1WQnkBHWNKz8KeMW5orCfqvCHEQIv1XLvkvYUnT9jyZ1WBS2LIac6bZlkCLrggsGer01g4GqAv
QOkKEztAKVW+sIF19ND9M8o7TC9f3QyIjJi1Q+54m1EjIBwAzWE53B3VZkCJBKycVAe/40q9hUkN
zzbpXmNmR55MaNXUlGa/ZH9QsD9gx4U5oBU//jOzAbRA78FozBxjHJnpgYdva3smJsvMfan+pRsy
0OiOSyqym44DTs2ArYm/dBwkUaWMi8uE1Ww9TgyzKROMtFXPEcko+dUNnK4I1z4symsDcGi11QRW
sUDnrarDVnp5d5YWpdI2O1/2DRfqSnDbWKiozJmYYTEXMhsd0L1TTlKtMzKplhNUHtIP00VSp07m
Tbg1c+7B4fRu3zWMpMC6oiqYJd1Jypw/C3GHCtWK459jmkUm6Gf82+fJZCwGKi2TUHlc7wcN+Lec
bmBzYhNagritLpXAQwuUh2IC6KXBPSkp6IwKIU0vrqPkbRtmZftLdn5LYlb2ZlgwZXaThhe98E6B
ssY+IJa3/p1mdeTp1ePv3QHQ8Wl1HdZIz+da11tmQYKmL8a+Zlu5IEz1n+gTspioYKg1dJGyba/D
Ayyltx/sn2ZkovL02VX269Avn/cfTvsUVnCdLQdRgSPaOlHgJRDnE5LZcasnA36tMAq3jRj6ZRM0
fQAlCwEf7VPXxahRuYMPScMDIRtxdFgmVLczoZQDWqTl89i/PaJj3vXvOaCYfgs//Z83Q1+4JZJn
DqbPN23rTXbxM3SYITEMGliL6fWupRjBBv5NljK4dYWpdAlYBhZ5Z2UQbOYG8Mp+uUSeZYMGaDHo
s57lxsx75zEwDivuQImrViwWFeCDwK2wSdiYtna5voyRhh3aBvP7leCuZcy86QpOUvPCMrGMucZ/
OFREb9ZVEtoSryt9G51UXZIofpU4OrHYbHivsET4rXLdw8jRxIcFCcTML4s0q7zz5fZyvmDubP4B
QJFVGFDbTO/PGJfY96pPFyiU//U/Gm+zhfRl9nmcTffZt2sxtl1kR2yPSatu/+5WFL7ia70eshLC
FbDPqU4WmPko8e/47C+YNjUmmy41fM5k31tZLntz2JMi6LgyU8dlzoVH6JeEbbzbJEMLnVGNdFSO
6aSN9DjTEHzq2YwrdRsSBfiDLQ5yj16GptkzFbDeGQQ61EGhmRdgLT4l23i0IOlMGnoYVa74jsRa
NNxhsaTl8C5C6KMQ2zusGC+yPmCiDOuiphQ7Z4Psm9jiM0um3mURojYgpL20dQcuaUzFYELtP/+9
V7RMBppEyZibtKhZa84Zmmd1pdo9omKAd37okUIQIBxJWjKgmKJsK55aLkxQCz114AI9JW56Hf31
2kO7Q04w5C7I1f+u6/bo8fWMBS8Sm9bD5tMhlGHtNlve0zRIH2LDSO3bQY7aMOiHQxVgj4f5PXs1
ferGJo4KDMza0+YmRs8ZXtaceF0tNYzNw9F76BLdwqMn6zTcP+CUmveX5xquU+l3AQ2bu7Tk1L8r
82bt4FQW65kt+m6HX3ZV3Sz3fxnHrQH85kkMwsAekgcTtWGp0OphJQRClZvwEU+PABk63uD3hxFT
86APi6GUfrUrReSoxiO+2RnBY8Lh8c7YSAKotso0ESNYzG3n5EBuVuRteBbft1x+br4NSG29Xy2O
/BRXBQWxJeqYGgcCmXYhIX4tcPO9BCT9H7z+RD5psdilCPVVbvFApZ5sCTq+QjJdTf9syzfhUduY
lqgjj+XKAJ+4RU6775ynuhd6JEs2eLsn/IRTEnda1Z2DvuuBV61frVVOfiR2fTmkDSNy3VN+KjJj
bFt8VxZ1ZC6yjufD7TaolzktYPSpBtB0yh9AXljqo4ZgyWK7OQ5C5tdJ+AegvrgmVpN3MhsrvEn7
nlz+lhKLWQQEUgMIQo3MR2bjNoAHlQ6Y4Il/Xo6ry1KBLPsBta84L1SL+97BrucLV9o0rMVAFWmq
5Z41znCGkPvCxN8thUuQqRkP+YgVPtGtWiXOLpd6hQ96ODT9T1GP7IlPvf1sOZWYUkQRY4kXZcxE
2uAsFwNOrdiHXsTe/39yNP/aLuSYDH8a4D/TJgFVB4z6RObYYM1qc6uWiwL+VrVByVJ/hon0DFib
VMWGoXr5NBYwr1TOmBnZMF2B4SYkra/0u25ZpPmWhmvQsiQbCI6GYBHeGVOKJJZNX0Nhlmjm4AIG
dWKDMFyWls5a4+llpJJLq1E4cWCb9sZE0+FpdLBRAQLauU3GIAHQiL7S4tpm/pF3jWlaZkM09Reg
469q7aDZMb/G/qC8tafZ3J4AY5FON3ENH9Eu7K9ijD/B92WbYGU2/gyVC2nA5juq1vWevMCc1SkF
lOk37EicLRa5AYAiEdvmQKbho7eGll0EN+Fo8pF6hTBIIy52cYKQhegwwH/zsC0Jk9X1StxjMDi2
JnW18W4sDei6UOuV84sYja5OB1CVQ/lp11ucJ978r1MaMw+QH9ZlZJdAjcO4Liugw/EVvuI4MAO/
q+d3QKWgoWPWd44MSLexlzOI0PKdwEaJkiCPHGH7SlYmELUeE4JlmgmiFoXwrzK5YHwezW7MvbJV
/4x9vw9OeH5OjJMQff5TfRFU9Y64/L5TjXsZ9RZzbHU0I5jUqI3i0FbCWkSz6LCN7K/NQvykOWp/
XadqZ/vPS9nz468NUOvNdlRUle/uIKjx9jtKVm/c/xQTJpr6f0HEkrkEzI0yQ5j8KHqlSBopToge
gD4/mWS8zs7t14MZ7t3U73mrDcqsBIIkoz6VlqNc9kic6xwkf0oz8SCWb+YlEgf/GY66yVPZkrJI
RLk6iSw7yG0Mnr4tW/AjFUlgVQ75Ado5Rc6JPebNpqOHwvuJs6yeu6XykSAZibmxu5gOosj1qmfT
sa9qnCou3IVB3MWHlRARJ8itWlOqw5BQH94AvSO2x8LDZpp8Bw93mlupy/aA+mbCFhmOqY94ZTAE
jrQqP/8e1QZGka5jmxuCMlyCGsL48lx5R9WI3Ws52RBejkpRqswEbVjSLbsVNK3ycZT3hI0qLYL1
i3PjJTHYFD+r49vmmn+HSsWmWA8GduiPIZ8Pq4Rj6qh54RNLhrpm0aU7qOQZWENYT7z5kYI3f9Nb
n3u6axc2id1MluJvgIUoVwDeM4VGHjVtUX2rMbDvgdg3lDk/uAwbQqMafdWYRUA/StHnPIuWfTfY
qQ4U/hulgW4TFMXWmeoIjh+gjrWThF9xrDX6nqR9eh+A8bPe+mfdDBty6itFgplMQstcH73nGfHb
+7MjFUlLwWaJ3ohVCyeEZAzWejmzRGLgkNWm4yrC+DPthcU+zwajKi2bBcBxrTgIt7e1A4rYAt7B
hHkDy312ZGQ2EisYLvv1W+s/eM7YEc4BZ0mKhrn70dKrdcewYuUsXjae/tsIvzHfgQWMdqZRm4Gm
iPuIqeVOuOP6djafNIBWd30Odld4LBB14wuwkvmoew99xABpInFL7Rc7gPKVNii/x/kG9qGidbMU
hCi1B04x4zUf3uYpjVe7QgSqjm21h0n61n8wEGkCqByl/mslZ0+/8BhofgmMB8yuh5wATZ+4FxsP
63Zm6uUr9btkGD1bABdAEgjlKPkOZTfR+rhbKVH2bUzElX4buaAVFhOb0YZpp0OMKHkxqfXRzhSS
Kbreu4gezL3jXoVzKsJHOWd0NUFSmg3PDBmx14ZJdF8HSi7N6eJcC1SkaP/Hl3xs7bi9shwhHYgc
ugLns1ynVop+Inm/uicCcsKklfZ5OKTCWcEI/oISVN/oAQAbsNVFY0Z3261s5x75ZkNptFerIBC/
KeIQpbrgWt1b/GLtT1naNHMdb/0bC7WXptJwph+QmVWcShk0Jrx9AkIwPLIpJ5Nc1a4TWVjJ2fJR
YjY+U3aQrMdxrtrdfcttwxGYLfVXu3FzhDEDo6NS3oS7VllxC3gGvaye0zrfTEQd8YW5WI6U5WvR
CKTWke/b8jZVnPKNIm+7gD1oT3XCO7QSK+LO1emfVV1VwcXOjU0OHbCaF9BeD41NJI8NTOTJJQeP
GqtpWPYtgvIdaDSRsC7a82s9AdDcs3U9az/mKohJc0EPWOv/YzwPVYHCc3T2NAPNvY0tsCO1gUF8
URyJxFM2o8D7zUz1hP7W2GUqKaHwdpRF2feRo31kPQP3gRUXqlk2oOsl6vWcOURiGX5O0rRf9yBv
iFYV8pp8HKploMNvtkbLRz3e3yLDL+61yh8Bey4a5He82JvVGTMAmdIdt7ISRCgOt3qEl9Zm6uNH
fzRsZqMuaBClbdZLsRteeP2eURGdmLRhUSXD7X8YHfX1Xi7WdNRW/4GB4/x/fEcEfff5Uq033PYl
E5M6qe1SsAzU09cDBgkwWYr8Rx1qSWL1dymHI2R0MbRfdGjT+A4k3BxNgONOe5RoLTG91F8aeWW4
aw7Ycukz7FrPfgInvt/ijJ/UFtmBF+vmhJlrJoueubfPAJ9BDvgvJ1A9l/xd1hnPl5iROr/jWwPv
exYN/wpwSGn14hLml6DcLIR6fquJ35dDa7uMrWpHs0OI4QeEMZfD44AHCzgiZoAV1czm4jO3zUlN
NGoXeNn+52xR5d/pWjl+2UJYRpo7w5DQD/pQ2gkBYd7O6kCFKigMteCndBBTYptMwf5osxVO+5RS
518E6YADhYoWNaw8sAwKH92y1GS7vb/oWNqgnVqE/wMgskkvEumOGsAjdAEVDZp61rNSzdDpLfXJ
Vns8JrIfLo5YQfeghDJa+LJjAEgAcpdoFO1Hz3KqSVe4e2b+m72peDF5vm7e3VcZKyB8Ei8p1yjo
niZFbeowV8YWBcaD3+qr26EEEiCmuguLvhElc8S7wD1JuHbWt8NDpJCc+HBmCragqi8Iu5g3Nmps
WMFQDSU9aO/PoYyGrfF6EN1bAFu/b2BHoLm9/LM1A0zqK2ps6DYkRWXMzL8mj5nptXMJBD23+ekv
rUfA6kZ02NAKi12HRwEzu3NK74Cn9zZkHKZZgnB2ETxv1jKp2b2gMY91WwdPEPny1qiFr9i+BtI+
Vh8RildHTv8NvMoRoCI1rmlxSIsKg8O/HlzfeSAs2SvaNPovtxIRhZUHKzawGoxok7AYDS8PVVza
W3QZ/1WVP9mY+pXg4kdFKDkOqBjtSwagp43SHF/iGMnZpbK2foxZ8IAZUaRyeo/xaSygGQcn5qbi
R6sSk7w1z8wfgsbDUHdttIGK0JIleoD7mXOo6PMY+xMsrz7QA646GQVtlewT+aiUOG5Rsb//9JAV
y3kpe5/zOu3tV/4U+gMKnyBNl1Ctmreuei0HnCg8tuW28JwuexfrqyLMJl7BsnOmWwL5wKz1pZIT
QgxFCCAZlUKeoubOS3TaJO5kmfuGrK2N7DYkSS78rE2NkYeUKrzhvoVJxWX81I0a9YMvpZFfdRGk
HS5AVyllottE7PXBxZw4GT9MluJ/IF2Fh4uggU0evQiUYbF3AqbKU6TEbZeRJ2NM2XSazz2fluvA
0+yjGJ0JzsRSty/PJecLyXsiTCcPEngvFBQEbo6jJBMa1YlcJR5HjW/bkWXCikk6gTYRVdNICtYl
h53G/SIFx3R2NmTFKjsGYsvcTCm9NcuJ06TxU0SZdQaYzpTmEtcWsAeGGWej5Z0zmXLkRdv5p0u6
82N3UBUzOuzus6b+DDNHidwNn70VR6qM0RZJMOYmNotQ2+FPFGqX5KMI19Gy2lIy+bBDia/9f7sj
VUVn+whfJGHHkPm8MqfqLmXqEukvAcrjg3a3E+LpkzhJL3Lt8SoHjAC8t0Fb5PdhCbu7Sk5rxU9R
5VHEcatzC+kc0D1JgrZDpF9V8TCM2aIPk2zIiC0WJE3Jv1u7CnxKwW1JooQmLEvhK2opnDluB8d0
CdzNNiBs95ogp1+iuT4n+SquaDI9RpbyZSKhZf0eWHi4Oe8yHOWPXxBEHjckifZ3FCC3Nper03aE
nDQT+IHUbIbI3ogxhT8tPuB6rK7WSAVHytn+IkqFO3vBzWwo8BtCCikoGybfLrPF9E/M4uGwhUlH
ilKR1o47QPF5B4JDatQ2mVvOLWf0DeqpIZ28SrV/JFM5vIT4aobQKjZJcnu0waNkqysmSOIXDKXk
2URoWH9SJhiLoNIdS7T6iwqm4F8JS9oK4wnNeV2QV7lMiwX2SsYSKesnD0IygmXPueRt/F9t6x7+
ejIKNlOlJrCWPHv4DHIORwK2cUqvACSoc5Ax7yX2s1viUhtNsGThXlpcBb+RY7aABlKwNypgJ6j8
D//i2g4bQQuU1c7liUuoqTjk/Fm8WZy5s6eIjSR6NR4sF/HIbvQGyxYswdIQaGIP6LZEv59jE6Y+
gYqoGB+7wqbsjEXM0fllQ3kM82gjw4QKio1RH39LVorLbNS9uneSkeIHBiF6xjEu6a4jysweNhtX
XCtkfxha+/Tu7aIy7dy1yt5sSKlQygjZ/ZO15TLhqpeL08izRSnHQfusZaJHn5/9E4wmNY/9XV6U
QKwCQPl3KxtfmlrEkJ2FEQGRP9RXR3NRQvQobcImLaxENjB1LoAiA7JzRruLC/cPekx9v3IVr6L4
JPxrpZS3+FL+YgWRQBnm3oq8Np1VZlKmP1oRRJtdxL6MH0WbCKQ89CnjXZ2gWADJNPG/e22bpyfE
EtvI1O2nNqDVdXX/jrES+nytmyd6RdQ/ljal8PLlV0YXrCk/xWfHCxqJMzSaK18h19UXHszIWo/u
oEB4foEUNw5GPLavR8gSC2ZPxG1SJ3nuyhdTwY3pPD5coQ3743WNUyJpzLgfHm8hCffT2R3IHKYr
mY0ZUDHyWTA2B4tEqo9lG1MtUTA18aalfoVMjz9jCh7WRjSA3E1YJ2MLTkDeED7cEbz1GFyfSkEx
WD8HfQ2tK8Fur+bio/AckljiSwmD4rGjaZJEC6TNTLJ7XHop6/nRYus2yLue6IttgWAb+5N0yvEs
jUi/8X7AmtWV+u2Co1eXA0xEO78urbiMLkRJl92GkgAvEWjk5C4ALbH4nam1jOYxMpE4UUcp8TAO
Fq52dyhWLAwd4TXOUeLGb+2zGIcFDMf2Te56NRrH7TxVJTq0kjtCzIEwv1FJA465RnEyDd7tu2Eb
LX2pJjT4Mf9T5MwFY3x2XXazCRYgSFUGvwJtnjLh/rlzWxjyCl1BwDM9sd67a7wZP/HanKrJJHV0
pVKa+MXW8qtNqjJbK4o6JKSH05EhrsFUMTSIOqA9ZAgl5z63IjpUygNmise5ACPBaTjxegS2S0rr
kVcQd/XopvcoSoPV/seKM5VfOiIBSFZ9qSi0PrbTywtODHv0PSGAY37qKKoSz8uQ/Xrju0593tmt
eAKTW56dt2Pw1s1j2gywweufVAAvnfEUytc5s8QeQMCoNUunUUd0iMGwp5fLmD9x124SHqpMCTvJ
D3m8C8iDx7juQSznIMeRBcZSPYoODPSCKJ9RhOJEBEV6v8U4o3c7Ctrx0OMl9v+UfiJWF0e25iH8
gQ6vgYgbX2w7dNHVzEOdbpfZKbwc6NYn42/akheF2aPesz71dBKLFi6JBO7/ExcH2fa4fETzeXbR
cd8iW3XAFfSSqJiEhIsvzOZibk+p80qQahpKwza/jjBKLCp3pTzq4jRBnkg23rdypPZD1RVOkAJv
+Q6i2W467GjYbejDiGrdQJEMZqRBv0yUffFe5+Ahe3WKiU/OAbrjOyb15fYfuJTryYdo7QdMeGWK
pJHvpade7Wy7RQrUlig1CBOaJ7ww76BU/Lip57anQ6pgKVBxrgXMzZyidK09NHBOCI5asQ0fZ64X
DgSJdK8Eq7eMMo7pdHAczEodsZJxFHFbwHtF+/K0W4a0pltkRe8abjsbSFxfLo81RX/WmUFJC5kN
haRC415TbU06wwZcFRZSLwqR7bhhaBGtvGTKXpXFjyN8J1RMgNisEN3PoFyRG6mXwAPvqW2yKBe+
k7f/rjZYULxKITWwOqLNmkm/HJq+MvFDSZJf5PYIddw5VVbia+JWZFWor+aaffSS6o1tYMurx4tl
nWMNmJciEf5TcE/j5oF8Y7xoKcq1Fqd1CmoePEzP+blPQ4WA73g1bD9a9ONAxs24MSI4rLwCdn5s
+DNAk+R8SKJkV7YilYFNgfAaev5VwrZYUPtzJpplTp1JiVGeTijg8lIlV6br16qA0y59NaS66ND0
/cHT8Zce/pULHb27nQx4i1J0/3WKQP5LoVoxlpbIe1d9OxiIr33Esncr1EkEvVTxR+VmcmcweTyx
AxHXJbDYMcTdfWW3NnfoHrwMbay2P62SUOsHwNk/AnuTn7+fIq7qLczgqe6k+FIvAhyzWSB/hykK
QJ/4dtF0ikSOgGGq0OZBTh9KkGEpWjYpgTV7ER8IYhjVAu2BZP/62gipHWJH6DVszt5USqVEZrCZ
pG4AO04DCa/0WBYo7qAn6LVI2Pz6qzjOo3KuBbATTaPjXkLU3H/K75nHVS6jKEX2bmtUYGi8dfHu
XLqH1LXz+zI+SxKBhcK0gw/JwoTlPexT1xqWeZYSBRVAXz/JL+q6agJQoA3mVJGzMsJx5mk0KiMs
doy8Yg4XK22KPZNfkJbFxaOBQQvQt+wUU2+iou/3poIS77iMA+dxWKvsbnIicxkf8WyRIgn/vVmk
RcGrrEKb7FEKAVyU2YoW2BvKRIJnnLrRzLScBkyosYpoPqNlhvsJhU3UaLpOrXxy0tLmFZLa7j+V
r08VLkjzcFQUTmsIlQFPLF9yC+LLH6jL4lLInWbCe7qe8WNgsTAikMNbgXyBawe4S0yM42NIPyQ5
GJbflSyO5dToW9cGlP+S7aMrdmLpX0+J3FGVLi6JblDIoCs23dxFiQR0YZHhXotQqr2pDpzB+Nb4
gvqaken3rk6IhTL/U0wV78IiWnvciZ1P2GX/8aq49N3ZSsL1QWdtG8gOaMdNnPq028lN3B5de7dt
BiOhvGG7hWe0D0mjbi9EsN4B3QEBfNIUULyBhhD5qwIe9hcS8vpJrMU556M9nO6tS8HYgc5XxhIx
PWdxcAh6xnLCseJU0VxPTY2En5U5K025XAWc0ukaZOMNKScphKHnXe2HScuNAej994fnhurMOMCG
xxGMiTP65+yrtvN6BtHUqKwoPRGV2Q2c5RWcFPWDOW2EWCcya36OqNtTGfH/G8dHkSw9gk8pa2n6
1QlrW3NJTzF1NOLxSVr2SMGvy0OCnxIueTsIM0BOce0gpl4PipfbgfCoiQcKZ5LoTJtAEiy7fDWW
DpWWNz4tGIlY2zE7v+TLpswYBQ9fdmOvk5MgSmG+JWfLcJyphIQrkqByZcaHlnAHhS7vYjdHGWJi
e5cF5HaZKs+1SU2yI3zLg0a2Ozv52LgBDDv1I5ZGlnL4fHYc48OnbyZ3cOzjnDXyyCkHT9ZcSxni
bG/dVz59QDSXtlcAcekVjMYn7UDyppi4sGhdLwodktb+BIhIz91IzR2MFsMHgBQm5n16C692/PKN
EN0QXBosqGnxuvx45XY5kEEK1sP1gYdholV5TVg3dOirE7PdSisO05ZDxG2qW67hvmTgvY1EvaES
QHx6ei8eX3jzpcWAlhd/338ECMKV22qe5VjGD670TiLIsmsGiNd3Mfay1Zkn6tjtfscBJDFUq5KZ
l3kq/fK+7MU0ofPjI+E/nGRT5zwlCJLvc8BFfAEi6Jzr7+exB+kpA8mQ7LF1rfkxG4B5xw7eKlCi
TbVvp4ax+QmuBn7+Re+Ddqm/xI7C+7+lK07vrJS/ghaMNFAPblk9FKmIux2aH0vCMAxLK8NAKT+u
SciMZiIO5GHaoJRPkOmjH7nFv/yPEsY2gxR1s6tVty5v1rvYbisjCblOCd8iZLbCzWExyLf7amdf
sSPvhrBs3hkp8pTxBeqcWOjQR3SmnvDOMODabah+rveqCqWufpdXDBL40Eh5kPKjpUbQLrJbjw/K
cvdp844z4Z0lUnwqcjUpwpsfMchqAGrJPI4kUSUbpJPxxHEwLOM8rBFJcInxQ0vjIBSKvc6/sg+R
ggRENqRklcSMstkfN7e8vyuPnlhKPiEP17XlzERm0Rmq3G5dr8sbVbF5YZQdIPjp06KqOzf8iehO
bCFTh1z+OqdZWnx/FoaDIIpITaRtXD6Jr217fSRVVKmTW6nkq0V5BuRDIUzdwQQakAw0orTkUgEJ
CeBpnuBp/Si3qezOgka9X0MAWzo2gVzbZ+aOPhR8nSXtT9ZdotPNrwwjqUzMYvy244N3r8gvKEi2
ZBjv7iDSfYWslscuLvGd43CaP7TQyRAbkq9bSAz3kKBRNzXQEb3RuV9z5g6IYfm87QhaM3Dp8gNZ
RRegNRHyT8bfoqLee4sqGif9LpnUrIRBJY2gbtsQYcYcIIe+Q7G+7zpBxVjseTUwMpENTLBROmNF
E/tIb2I0ca2ppGbEnzeUnLIj4KpH/6FyIIYp0miHerA4/J4fMVpNFeevB1W08bLvpvzPUW9tAjpQ
kDZ7RsGcp7bxWuhP1DI+OWtXSMad3rCtrGpFOhqZyLiNR+pUVsCS+hoCJeMuyJqCDz4aZ0Bg8Q7n
M8ioLoVhN9czBLSjiRpUK/AJPaABdDSzGdKEc34InOGyHqt07pnEbDKZZ34+C7yMEtzw+1nQBDwG
JUCsLQagUK6PA3sEFozdil7/8muQD4xoEaBD843d3VVlbcxck631PxbtSyX/gER4XodSqunRKrfk
OssjjEN8dXd/sJb8S9OLpLfoThKrlu+vfcbX7//1AWUJOoc+loSYpnyeslf8YUxMs3zVqBqqtlQG
5WIf/8JCVm7iOV6ZrlXK2LuMZ7aDIpz+06l0elGxYkrCX5prRN8Rl7kxW92EHyL22HAidSAn8JXc
U1NENQZNnb0jJQAjDD+IAnYJzu5srz4kTcXfJM27XBfN0Lb+3/RxVlPiLHM7Hanc66BbaNSO9gpD
/5dYa9m9W9LLFLmzMDIeE5KNs3/kq8fE5VlpQc+GCOvJrfq6mMgmuGfXTDgWB7ne8OCpqyeZdYcO
Qz5pkWgS0n9Ez47AemMGJwRKNsd/KemgqL0LkwnWuuaVP6UzsJWuJ6QlrD2yhPJDV6aUzfWmUE2/
egABiHf7tPTt69rXgyI8IkEFAbqA4u7dYHISkiVU9AKY+JVxf6lGcwHw0C3HPIVehQlpmHrzMaA8
c7dmDPnK4h6M2ZfbD5e6ple9F+KA+Td7Io85af16+5n6jSH1R9T9OVZeG2J+6idEbGPxNY5RmYrK
TLeuWbWDBvFsaUAB+P+EQuavu6CKatWvi42a02GhrVgwFlhc9+lvmWjc6KtaZfzs5N5oDt49CpSs
AiZq/vFEcbI6d5tjRLPeKc03C/jFthpaVozDNKCF+KfjsUC8DnOwdA1EK2Li9fV0ddrG/v3Hyogn
bUaEs2Wm3w/6I/yTStFwRbfNiZPWoaeucLOGAPocWeClXe90yVaq8QWkZX52h/R9E6ZP4dGZF3PY
kcSpxftoQnlb5sPVJbOd/l6RyBcMlvLfatBuQMxe07o2uXWnYJYto0N9jqjLF/YU8/ZhAxaoFHCX
+a/3aiqvHEOJ6RprtG+nZAYevSqdDZehN32Ijj/QZt0YSfTIpMpJdj1riwVfeQ/SSxv6ICgVR7+f
qoxfs2WTsmsn5EaDmtFK4WN0ucQQPEfvhcjU5vso9BTcfudhyzX/czIJPcI2M+gk11uPzFZjhhtm
+HtEfoqkwnzUUv0yiteaOXABadjn6NtW8vtvfSIBHuEKesI/nVTgcGv4Xc/2MeXL3aF6kgpTjn+i
sZ/JpCUJD69c/cyhoV0jFmTdy+RxUWA5mdxcD7ehMN9SFBfBT7oorE0/LQLfiL53Wdvq/caTcDIB
UruXbvsL83dfFJXZkwBHYfHXGVEfAagEa1rz6K9pOQTLrTsv00ID1ejl7SZHnffW/cO7AzI3dFo0
2EOdWtjwnF/3zUoqIl2aWscVIqfeqXY9qhJoOBtXdJQ7ceqCI3c0G069EkuYlNHns5r6HkGSdSxp
shlfJvycmz2ZXRcPxFbNeobLn9fWW3jzcaEW39mQEOczfGQrJPZG//u713591YB5XVFwgHchV5js
xvueWFk0waCLALfvEULcKoncg39kmLX2Vslgw8V/7MskbE5R2OTMpcx//nSKjrD+X6Ry1VyglZkI
mk930eZXEZTbhIP12dqe3YG6YgeyGrY/qglUl+l6urmSeI7vpxrZ791i7oqGrc/aKOKZURSwFIOS
Fr+9r1f/MEV9tp+ufxDYETOtCdpBrLJ4//VujCWkOqeWK2Al+uLiwl/fKpk4GoZWzbAW03oN7ZRk
3KikMMqwaDoZnihTNaZ/oMxgh8ICyMlEmPALDeC30UtovQaDETGhI04MOIoLoCazsPCG1sFUd88P
5yoIv46yRroJb0+gPVi74Sielm+S4nLiOGGB3ykPRtTsGZrqRcZZNzJFAUdeoJK4Kbc06EDniqz/
Ayiv/OJeW8lMyMT5NORHdMzOm4KARH3wJX64qfYIh0hgd/iBbzRrO/iC7N7tSmsYSYgAyS/eCg+D
332ASiqQhTvLSOWo6/4vw5pOykdg35WYrg3zRGkIZ6MHPuQWhrlvCfRLiZPSR716aNvDYY3M7Yqx
eHFr0YT4gQsBVKg8KtaaWN0dVtQnR98ddfQOegX3xMT8Rx90rPL9aUnin9q5f9gIYo8Vub36rC4o
2VVZG9nIevtUaBH9yn1eGLWJ/9w+Ypc/s8jd6QWBKuHEtBvlq64FmwUIk/W12GZl/TbkykAClilc
C9HraxNiXvs3kl9piCiaN9ZY3vva/Jc8em1V7aSEy8w3EYwgGzT9450bKEqLi7olymr/7P+UfE+c
C1kbhnRfolhmjn7MYZgFRwMlVvKqWtMGDVPX2sW5nCB05SrKtZ8o02Phx/Fe/Sqf9fcjUPiE7D9a
kmCUPIGhhCIh4v12jeFo/OilY0vi4mJb418UhY6aCR/JODWyjWpSP2vppTK6wWeY9R0CGfmCeWcf
0+HnQRa8nVySHsyxi0m/mhSNE/aFpjOsiylr33UOP1MxkpO+wOVzC1HVSxgZes8+1UnKHLl4Wrww
i/pxUn1MrlAnAD3d6C81DrlkY+haJ5qY+V4TOLXIQASdLN+URBaJY4GzZ1Zg262tIxFmJAct2be7
wQro5QKHaMVrrDMcpAbE3qPtVyE6BIst3u01wPB+DAg7jieCQ4yvjyTLxkKnXKnCGy+KWJdP+U4K
dmC7g5elI0EiIgIaNxXiN6/cPt0UH7nCUrnDU1aLKmWiQgeELNpzPIPPYoZy6QogDlX8l7diaQlF
jccbkaAbS20Tk1QvIH4rvPkeahKOggS1aeoIsgEUU7bRnhSqaQcZsF0gnuLHj/pWbKPWTjdlB32V
mOakX91+mskPqP2/RE1DcH64HBtaaQf8sHaGGRblMZI4wC0rZeMSe6E6IdYxs5+qAJTcwsSt6AiA
g2MACcdw4uxaIN9lV6ofLHnicW6Cur47xcREoJx6TRdaUxyJqJQyP8W22OF7OCcKwpjsf5WEuQK+
G/W4Oac8KdmCGXgVzeRPFNV1zTEKN3yX8bjYRC+xxE9cNVtGsgv7Blg8JXTY2kAck1VnlNRH7WE1
ioFQx3w0ySuhMszkSN3eTgU79q6b1hFFY/9kA2UB3A7u3CLMnuje+P5A51r9LWWhBOCIDznOpvNQ
lD0goDatUTJ52n4MLMtBDQeDTicJb3/q+w+KvC9kxXGp22V5S7lbp2p4/5sUocZqCiT+k6YVecFB
6y2zyeR4ZeI0cRp8YP41NdMi4QMCig/GWRV3mEiREyTXfSyMZRyi/QtLLCBvaroIHlj0ahL2Lryo
hIgTfNqwhP+IcHW7e5wBMoXGu/RUOi+195inI3jn8YWjK+fxBjD/Xc9hCabW06CtzcXCqP3AccZT
rw+RkvZ0rjjfaFmlgBCGDSFfpm6ms1XWNk/j2WZ8GDZdAcQ5POa/0r/QBEl+1ZK+HvOnfeGa0jQX
VhlS8WkNzaERyjvLFBnLnx/V++o+wick/Qr/V3bSeiPWKhtqCrrClw0j/iIlyXXhQ8jGpQf4Hwh6
/V1LCIQq/K8CIq036bm3/DmXTW1fTPrwOFkCMMUbit36HxTRCTwEEgvP2ghY++JgXj7n6v252xdS
PB2Zrn96mw6OgnUxomARVKEsOCPxIr9rx+dUmGMUVtN+uCQlr0rImDYuplRQVXUaZbLWy2mYxgYN
AcPPQf9UkEIWO5U0pzlcBEHgmeq4I6Nc4zMTqqs4nXi05n3lDXpIsyKkY5zsTUqWqovinxYp2eiE
I1mf8eeCr7zrHT9RaYifPg29ntnwioJeGofJHZwGU7wuHQuyPHR/UvvWCjNcHNfZD0byISMUbJay
DJCqvLd64pfTzFb3C7C8wVRTWC61rrLMeKeXhhEn6M+yrlXjtLrBnjQNGWYZDAi3OAD3GRJdiRyT
wR3HNcVcZ8CABHRy3Lj2CcyIxu/zy+Tcbq7e6wJLT8bpFzcrvQMoIsDu6ofY+N9isejMw+oAvB9t
YF9foWX2BNwdDAZeYKcqyrBfWjn4+uPuKfTA+JUhE3qZCqFIYQLG69BdzGyQF9IWJInhb9jdoJIY
M8fopGvGwv8sTcRxFUMm67lYjuNynNytc8VOL5QSP/u8nQ4dHWfZ9ULnaVnB8+ZfFjh47299behE
M/oZ9Y14OloIppRUc4Mbc58x22JBUhQmh1pbGY7uAgFzoaAloMiBz/ZAYnQZ7nCkLuht5+d9hqB5
lVkHxYpAGl6rplg12HxQvos3tRh7j1zUiZA1evUsRR36JoRjezzXkAGso0wXJWAPtCfw4OlUFYMn
gDYcE1tjaPTNNUso5DZrrMwXoy7NlBN9e2GePXNwHBtIviAOs9VuM/utQqSYLMSXiEp8eH8YeFEK
Kj29YAkjfw05Nsod+TCVybYV2hC175K9XAT+KZxJ0pMOVvsu9K7SmBCZqhgf0wwW4qq1g3dfcpVr
zYYZJ0Y5kgc5GiPp/Qc7E/cA5x1BS1j1OP3n1/eTiLzLZEuzJ8dKKFJ5prXGvThJ6Xhwjwnj7m06
HAn+3lQy4WJeGQn3uuCN5RVOewLA9LLH8lCkQtxdxP5CRVWMWla/dU4w3nvB6muaarafpx3c0TpY
aJInAmkkYppQod1+2yR09khJct+DTun663Mo9P+0YZAfDRx8/nIQ0qQR1kWgOP/I45ZI3+1ec1ew
AEWa9sXiJlV2QDphyH8yd4+Dw/BR/oQtzAxsj7/iRG9mBX1l2VJUE4n4bzVLQHQgauCzTp1brtO6
t5JAqzA1lerr4KrP4yST1bupcCP/2SXvUcAfFzSeUDBikn/T2XWaQrXfw2JRuYD7l16u6iiKAsnD
HRtbzV3XDhSpaJ8h+plBM5/i+QXnO7cx21sgJ7C/oEuPxX0oh6ozBFYL7ODGJiHFWIPtPh76t05A
TfrvAMbTe3oko6D5jLkEcgrSfgIpuW+j5JdDiyUx1ktI94GDXWw/RBdNpuhww8isZEwXajcgVAS5
7eRYNljWXQHnAy7kQqyoHvvLdhFwGWnTVWFQsyWaBCsLwoxrZmeDUAnuz+Gtmc4L6bgWLnlP9qMr
EG0h8Xkusv/PXpbhnJ5WoWNxs2YW5Uo3b8tiVTg+eucBkADZiXfMm6vCjTrMRrGil7cFX6w+BJ3z
hZQFXpJ1zfCXf6YPk4HA3FiQtgcVidRu5enOTlaeZaf/Q8ChKc+lJM21Y6/24zV7Sw2f6f9wBMyu
4FyQXHLwyQ0xkWFGyVfE3o+B35+DSlnGC1nNsndMyXE/tlcEHpOnTFaTEoB3NFC9AG4saZLRLbYb
k5jHKYVbQILGNatgsT4l0DOYqb5ISoSV1T7idBXKQhVIQ9BXNrEGHu21c0yBJXDX4/HD5daAmJsw
bMqzzdv4FzE7y0giAGQM3m1F24Wg6dL+mhW90tF4fVvsb7XCFpUUIG9HxC042g/NaQX6v7O6RME/
IeyiiFGc7P5kghy/Yf3DJe1PhLFVGmZ9/h5Go6XOpC96yKyuYj0KDLaI2wVdrqgN1Gerzy5ZKNCH
0byk/xr8nnQdRppb/mEUa73dUlzUzHVH3uDK4HkFzBwGqoJsMqnTM+Am5bBnmstkk0BMJjVWUotE
fClBEKK+edGcMHXKL/Ph1uo5y7lX9cs1mGMi2PFDp5AghhePidZ6SzGPFz5fSPBDXDWG85fUVJOr
nfBgizSPbx/xH0GH+JTruPf+lHa+Y8A0q9DV8zEN9OneQBKkisXrxyAiaxkLLvzRTzgYRjYSNucG
1sOe1tWrKmLLU0sriUgLTHfDGBK1Q4rvp2lvu+JAPzCcNEC/g2QfvTyqF5bv5w0uNfhh8cJ5e357
1dGFjsjtrGzeya7mxzMr3asTo2X2X69PJEU3gBPHbclBPaV0++J6SRGlmQsslfzBrJop4mQHl/cr
LGkjDKpcqV2Z2AUoPeiraYIaJfLMJJiCN2/VBP5TRO+rh+jsTj+KhWcZsYF8QElJn5Ak7rFzSjHW
elOL1PgdUR4i1EgvHL1AkTh4uGM1IwCGdeLcqQbbASBbwODCmXgKuCMzxMSa0GoZ05dSqmLFG6q4
Ka6VMhUv4yHDAnumBfZV8Ap5QLdds8b+p3UVMHlFZIFmAo0YdMMB3EJGbYlZJqk4iJQx59G2ANth
n5X39YDnrJN/W8JXJ0zud9P/HzX4fh2DawgzWWzzFWjsaIpWab9yf7AS04nNmXI9J51rUvmlUo6n
RE5dUPZcloXbQ5Rqhy+hAtMioHdMUwJuLOPAj69V+I0UMOrDJBRzUQxWBoBy26hi1SwH9aAUJ6AW
QyK+9cxX8Y6rGOJYKj+Kbube8EJKIE0NwaoMKEL7XS1lSOF92KgMqwPlZMf0fb2iaoXIanICJyrO
Hm6AqWSX0lqjJ+u5UYPLbjZvydPQjv9vs8/o+BTpAdlFbTreu6YWK1d/S0sE8DwZxs9ERbw1lgiD
KRZX9YxxihWgUccwQQcltzsiULuDe894VbQoZ5Z/44mEexbxce2P8LKAFttl9jF4/oQW1ol/WdBW
dj2zEpUENFKSu4lNbletZfJydim5WKZm8hb9D51c+d2EHO76W4Z8wPJCg3dtgoAEQ4j3WB+jOp+k
aK340L5HsX0PBjAV+XBr1QiKsFVowgDPgP+5Qd+a+jqv+uYs7PMsQiZPqgA+ze6zr9UHiFsg8FtE
jTP4B/jeRTOce0/9YzzuW9jpjUMbiMuaynPedjk5pA5mZOivGyYrSnw7yz8p8TV1JMMaIVHK9zFw
RUdQqAMa+9kFIINy2DbTnQAYuQCbLBWLozG4kfWLckGfRhXwfhxpFnPmXtX3uvKqlrXuByO2zsw8
MIlRo8/ynzAI0A7Fg7AuZ6DmXocCpyHOAyxrFT5GS5o0YnGN/5AyZYMnZdH6obZzAO1R5Zq67/Kk
RS2mgpFlTM8bLVyhc6gpDXHldZqzr9iHWO4nR3JvXc6vaggJs61XDDhlMd0+ZX4qp9qlrh61vmxA
X3vbJJiVljLi0e6INshrznf6gjnPA5D6+WvC+CUINoMjlBi4aRHtMFxqHSSfiNevSSZ1Ymzghm86
MHEzEFaLXS9asOcREOmrJUBzJy9BvphztFBdrOsd5b194PSfKDQMi19FI++GAXUvtvhGTtBZh8N8
RBWOUnGohbmzLL340rBmByfEO9j/44+cAkJ/4MmTf1of0NsQSYn0J7n/wwbDYZ8ydOnE24XolohZ
+4AhuD6MdcQQoU1U/l7IiEb5rI4j3JhKNMIA4rA77NgnxzHvfxMhgdNFp+G2BWYxvo0QEPwOvycA
iZoApsaM+cz0GXTrJsanK2L1Cshhe5YCy+C33T3gOvhZqcWPKbBejvd6UJLXZh1jShKbKTvT4HC0
lgzwJ97TqhyVRLCd47sWEEAq6hj8rrXfh1djz7efrCx9PLA8JHmOLgejN9w1GcAGrkb9leI3EOSz
IYullWbPxaE3L8ULYyDO3bl/5DSe3Tiuwi/lI/Ro5khr8GqOEqk2f9aBbgV+/6M1BhM6jLW19x0U
EnmizCN+jo5b7fJoNSGl+vx8lX8AjLJtbOF/HQunlmkDfQl2viDIMTGlOWlsJeoNueksg8RxVvM8
4z3SdnenacKwbOd0+Cv7aOAXXSke+1WbROoHfaFYOKbcuw0I4eXLM7T9i1eUP930UR+dQsRKE2ku
+N95vvzhqBsLxnX2A/Vgo4g67WU0l665Wz1FYWmXzWV9HfTRGUmON0LNsC/wuqTroJBGwcYZt3+M
AMDjNV4e4PYSIqbodBTawWcqwrN2DkQQ1a/EfMRTeXNfGcfpRpHU07rkOsW36dhwXJ/iV4sJYGKI
v1//FAzURaIhbbqCnlaSf26e/FeQVEiXKTS5ZiWo3Ea35IxgF3+H2aIfCeCnIDr6JAiwuLULzsCn
1nJiCXEz+aH9dI11rwPbyDtvz+A4x44apYR8F0nPVDxU1gukN4ZxNdCBmvsFUNWmbGMxVNglRwiz
he+5zjMkLiCOwlYFntdWm5UUzdKYvzsSiDbwE9e47x+j+jODt6dl7FqrNexYtFnq6aATpBEwRPVm
InHRHofZi/s3IU38o8e3nOUAuEKtrg17GabogzrBCPwrnxIa/jF8VS/PXcVUHP6sLUbe5e18Stjq
vBw5qNM9IDmpp5o9SWWmynuGmdzkMdIXQSoWTuy6uzazfcXQS89gxNNgpFPz8HWx7EMx6a4au3Oe
xNvYy+VgDsAGwE/lz+yCXS852f363/LNfWDJ3ti6HP9BlDqbI29gWZWVd9lzMVVf4I4INqdevbVU
rXu06iEJCrcW24t56udykT2D+YWRV3jAyMKwooYVIYfrCflVAh3xuKqGKQHR4I42ORAG/92O+wCU
GMmWdGFMLG/54rV5IaF+eXHqUXctGpqlxVfeYQFpBTMj4UZnvMVLOTglgtkbK6u8Etl4bpw0J+5i
HP5g5TdZe23IbFtty+sNMTyQV41jPYW5dfHgazGp8OIDapU49XIV2rw6/vv5gV0zUpuebg7TkYky
ZJiFAjZtvdcqtzVBk0zkDi6InOoTyPEXsIfVMdGq4rPXi3m9Xk5LuF+W0MhP5VRtdq09frzX+iYQ
dhHgx6XpFgq5VVa63Xb5hQwY75Uk615Yy4QdtpJWbXiQW0gA3Go4dRsDfaNnhQJ4uFzxp8rDXlv3
+y/k+AHUzS6ZbehjJOKSW8+6OUQ+gq+ygmw6ydMATmCAD5IPT+thcKLBltTuw0OuNZMtaA6SSupN
b9rpov5AOvjIZk5sl06Jag8vMBTHhw+OJPJRAAgUV0EwLgYKgRfV6IncxKuFsbdv5rBvhH1U3/ia
/5/0EF1lsLRMysMQI3kCzRT5Uj5bq3vOjCV2ElYRmpHUpUQmUzdg7tPuCNK0n8uPng4koUb4XKlm
fIr/o4RbO+PCTgTquFUrcCwHsTK145vg0C88Xyok7RTrIBtvKguyrJtsNqFbegFfYGIIlPqJIDPM
Xd5sNHxo8e5OXRLRTOjhcymh0U4VzKoxguQkSLTj84c3OkIk2OTBnOa8CgY/dwjV25FaoaYxuT+0
27gVQdzJaonxkHXvYGBPb1PAq8tdNHvieO3CVKcbHG1FFklRP6c9qt1N3H19ah3LrkZohx6KGfa2
Uc6sij5V0ZAulWJKdLIkFK74ASer+EG5GOPc4sUAfKCPZa9+vQWsuFlwTyoh10WsPsCPY19VUXRg
lBZKtyS73dUEFpEXz+kK8akLbj5a3JRMeZQIkpbhCi0IGNRSnjT7Df+MN+kxCNKNa8iwkaldfGym
cp5ler00No3xTwBkqL0OBTjSaifURtL5AQW4ZLAEs2EBWh8XOnPIy+f86eLos0MJTrutPG7qdjI/
ADiENqbd/+++8bZ2XsEs2WRij98Tqk7CeBnGpmyTwRymYGiwwLO+NZui+8lhGFzTxksKCBKppPP0
jbrZsCVRTy+tU784uEyZHnxow9IYNjxHhlggzAmHojl1+j/KFgiVuaLLaCXlwQC+JTGv6xsTVzyf
lNgvOxYN8J5gW8oBi8mEdPbMObuPJewOMSDif32lNB64b0lPr4vtk7g+2hl6wCWT5ryU8jp4ArHl
nVmsSwH+0Yfcbn6hnjgaIXm1gxcvmvxwIbhe2iB5rUkfzrJ5PAqb3+vBsHhtwqvDLBhhzj3QoIwa
J68zE1ztzslNejS35Z5J66Sn7M67/OGwyLlcVgQY5W22JOlePZiHdADeON1lyzDO+sy7pFa4UfVI
4dFB7sKA6RC407Bn5OgfwpJfL/CrhtnzDXbG33ey0cMYyRCZP5w3WyGrt6nPxoEDAdW7sypuG4Dk
yaexgZvKPzMoau8VZ8CJuUR74NJKgif5vWtjE+g7sdi3aqg8n4wZfPw7sRbq/61swc39OdA6yASY
J7gX4eZc/rYpP47tbf2A582xuY15salDJfayctCTmXRD8Hdvpvr/p8PW7e4HJzKXLrxbBelwi/HE
fKumwx8XAnguEwXTw/kZ8ic1os6WnBfXVmhr+vUh3M4+T/yekmaxAmcfRBCiu/vbox6WTv/vH2eG
AKf9jKlhKegzhnvcigIh0f/0YHyuAehX1WJqGKxjxASilC1agheKaQhbG3dByKWS+hmXPaMEtHXv
Mm2j6rqMO7Zfas9dpQgQ9nJUsneHe8XQAMK1LnfXieRq1x2TVTkbOWp8LJB2VdqwlpNr/CgZZOFW
aNqzgdQJmxqE4oWAyOsFn9memlRNh2QNmqpJjhGXlTrwaoYC/5B1JUT37pkWFuV/TryRSo+5u/br
0lEl3Ht6GZdkKXZUw/+J/TSCTe8LYjML5qmS9/ztUoxNAuyyJir6siZZgGALHtUXECoG8ssjwswf
hVaSLf7K34lhTowlykkVq889haCJucMvUb4y6s5t/qGOca0rXso9DfnQzUyxEh6hFNjCDJgnLElf
YaeH0CKZKEE5A8VghEtlUFlL7xz9IzSaXOzpHdGSYmfG1Pcaoh03M5lV060bU/CDKb2I/j7hHXn6
ds7USinVIYRCYpjTFz+rFonXxZqdEXHZF9DkYfycJGIwogGmrRJAN3243Oy7q7HRzJZyrfHOE5ch
80WJ7/HVHYdTgoewHTkD6y4je9O+hohNklVkEYrJ10vJ5w7FXJHi9PkuHl8qrxmmFEsdqoysUxVr
yBxO6glYw3JFwuunJ/QouPDOvtz+CL1gSPkMy66Q5ELIKfsunK2Mh9Ffw+lSGKzmXQxglgAhUAUA
PV1o69HcAWLMBr/Y2a8GVkCyBmg1uIiCDA0xCf2niR7Ybd62bBcXBC1lAldYBhzJszW4ZmZo7YWq
XRDz8jXkg84hG2xVU/50HyS3D8eraIoEZOdVUcMAosaJg1mLU5maw2b3LtMzA+rl36x/mrXdm+9S
Zv9bNXdNM3792XrFggsixuI4tQsoGsDJ8NDodSUxIIh3Kd+djL1CEIbc1NJv/DowNWUMVvihBONT
I/zSPOtUAwMChYsH4OHCcpfeHarKgTk1VLp4dEw3PCXxzaYmkSaXZkHpJie9gk3QG7dEbfE2KDV/
xovs/4O+3Qbx3kijVaBvvO+XL2jYablycMxvo/a3+6lVCkU0HCR2Vij8AX37C0CA3/QxlSDCi09S
0rB7v62n3WhS0jbeVVt9WpA1R8Xz+dQNkVOED7i2wTMFjXWX85NDIB9g2ywkPs0I535pd1n5G2z7
6vnrFr0W9AaZ+EGCEUDv20m9MAyaRGfgmzpdMRZcXOhsiual/KJwiRh98hzNylQIwVMWbS7WfgMn
LND4OsW7rswarn7bOcaFnh1s0qmYV5fJZ69ZNyzatUNQNY4YASS3CgCfCKWBZdv7xK0Ytna2BcbJ
i7wpu1QyyVHI8i+L6EJ6KN04fK+3H9nC4hpD4bR5LJoJKuQ9/y0wt4I6NfKy7WLbwYHLE9W/v2vj
neuUJ9I7pALN3D/9sN8xMZMuNb2LQtxeB9tLtXyKPDoVmE5QwWZhchZrEA9stwG6Gfwk8dq84yTg
yaKTdrT0ERbWBgoIChHM0j8rD181a56iaSRMxm7+Podx2oOrqsXluEVeOuKRdFiE/dpbOrSr8+Xe
nOsc5gDUjGtgpH1sPxHVo3F4G+sH+wtuNNWBz/xzpTL8rmtEx398ebKsSny70fjY2peccc3bRjiT
IpPV9RDmkYwui9iSO1Xiw1yB4JuUGqbCYR2nDpZSZOzPpKf3v7cwK2KFtRMw16ODdsJIEmprH0wh
IKMbtQULuO5P9qnZHcw81f2IHvdytOv2c+pyR3T1PlQjarxbxSg63Vb6Yi/B6o8NqEJFe0p8NS7j
5OzcRLag1Yx9ge/twFluRlRXNQ3EmJFQTkT3yTGxiYdF9yZCaRDAIdxsYfW+VD7NBX8y9nNlBIWR
0/d8zI68CcwyGu3YEUjYPCexN5A7Z6UaQCv6q02AqRrxGN0+kWwheUPh7Zuz8/k7JRgsEm7DdPx+
rTn5RnBz7Y1zvrqDs+W+6CccVYaYiVdnOPVPl2ZnHyvFI8BPhjNDqjY+H9RgC30IYohuyo6NncFD
nSZpBwlURbuplS5YhJl931WIU9rz7uXK6QXi01TU022gd9gPVwRZKkbeUuxSNpDrbxkcSt2/WlwX
OYWCU1c9BB1dAtVk8Voe00bui8rm/QlHiDmzpp1YMobJF3bzaxn2sJQXOHpPrX+f6Jk0cOcLK4rd
ReVbF+NIcZhjJx79fe5OWk2maOxIU+OO7G+dAJlyx6yZWxC+cFt63qQrQiUGwdCEzxJJfcPNXZsK
riRS6324/9f3AOAQWHXR0riXIKxrmj+jFZeh9Oytjz45seSrC4iI5bYuBUkPC5dggtSFybC+mjej
Q6kPQEXKDM/fOsJmyx3Y+xq/7CkHRhiYw6d0i5kDwaKUh9NsZNLp5ESgIIljL+nRRWMkBOYD8v6M
dN/oBkmaVUu+y/wfntZt4BPHo5LDCxINzifzay0555+nrrglqW746uAHiBDlOaO3N3UUXk/hX/Bn
Snl/TGeVAVD1MDEE7iluPICpJzO89ojczVWWxO16LGjT5Hrx+hEkwKFu6u0xDYbCN6lltDLjmj9b
msDPU7gxl4ZKuewoR7+1tJngZYKhtVSFO7zKNHrl9oyMOqDGULBsOk0dmEXQOpfdYHO4YgXV5DYJ
hXmXyrRs0O/u30vcCOB6hr08xu0g9H/Vh6fW2lQxDnx+ni66TWe0yNJIKNY+jXJycMEii7MQEWNs
LmHu1ZG+f241TNvYuJhuSCgclCqtwAXloiVG3Ca/MOd4fw/NGfFRRvT8uJL0NE4J7voWU5edGgtd
oErKVkrVyqkTqGCM3t1yJ24ZaoRlOBdOU70xYfLaCuPtJtDGqR7d+5Ia0AUBuY8aO/PIKvis0sOs
6ueCusSBmWQGwSFZa3ZJUpp+UtwB7arlV1UIokW6le3mUiGgkFrt/sylJG3hDDTcgS1Z5Sw5vZ9Z
1EUGCHZxdh2GTC1/9nxORhWi9bF9ldj/ppTYdeODio1Uns6g8pF6kJ18x/D6Z1RJOaOTtz0iU/W8
vPeUxXIuxQPr63uFdjl3cHnJlIDdwg0u3QcANTk4UyMvlWg+KEfVV+G1vZgjZjs0iiF9/C2S/SKS
EAKC4vt94aJ38MYXwsGM9nSuEQOa+PROCBQjVw5MuGq7UeNjKTiljI0gjsKEyTKCoiMnXyrGUt4r
Jrr4uFzqJxdAaCQfj/ALpsIhYj/bZ+jhIg6VIAgWXLVwrW6fGAB4PPqYYFRSyvIW2qmaZZ0/DrSM
ZZvgKXhErmi4pMnF59MkpognsrcJwi8Bk7W+mPMT5yENfawe0KNw6FJAm/mnaG+8iArrGVPvYp9U
eDczRHGgSFkn94NaTlCLek1JWmWASBW60qhxUnG+Teh5n8NtsWqoIoFVz+cUl0RshZPE2xWvtR9P
ATGkOStATazjmpcuMFK+FaUcOMBpayWSgbUrMVBlZCtAYPd7dgfg+gf/XBQ/AZAy1CnV55Yk42Or
30N4MEu4Tw2TnecJVnoTh198j16jzFj5NkpPw6NCAzGTThyUwlQATdWvnqEQTTrd4AS2dxKES1ss
Z9Vre2sEHu48NvjzBxLiXU7Qgr2Ky9pwhc0GfzZgRH4IjCUeZv4Dab7GfnQwP/nXTdqqCfA7GmQS
fN9Z1I8/5RBdJRESdGobrvTy8awOi7yrawZ+WAT5+rog/J/+NLHl33rjArKFBvAmtPKZLIkfoE6R
p/pPLynFBKK1t5GeJMrKBrv/EENk/7oiotX8ONZDE78MZIucOE+NLv5kGlNL0pZ6jvU+cuW6hIbV
qWH7hA464P/zFIUhM/fKtKzR00wRZ4NDE6ONuolbCBQ7+V3bStYgQae6zHRg2542xgB0sHj2FEZe
A4GIluEldJVQKbxJ6lHpGAkI6nay7mTdZHfLzHhKuIFwUEHDd77aMV3Y+W89eH9TdpTOd5XVcOQF
58EdrcRvAfgAmaDtz19ypoCxrQlAyvkO/rNsygMplxt4lclrpCwFb1kXnUezMnStYIQ8vl29hZLP
49TUoNDdRWS+fTQ67iPjx+2QSfA0YrLi+C5xFQx8uuFFKlx822OxF4r/oBlt9bpzxXXdb0/Ng6uH
WBjuRLK1LQN+b6dmbVpgL/9u/YM7uBq7nkwvyH1GTHyj0KG6ED92JftqrxBX3Dhw4WT9hfFXcdUg
p6vn12owIe0EvLzVorOYX8Bu128lqCrHQ6nNZnW3s/nh4MfAiKKFx950AZeuxrkFbkCx+6OcLEbe
8xUFXBnCM+s2owwaa1MQZS4ntn5cSEEAshVQgyrLvURH/KASsVIaKzvLK0FLHNDXOfJC+zw1w1km
W+3lJxNHc3hO/x4xL1z8kR75egkIiaFUzHgknXQSIkGjSbOxwZ8wuQpuhONsWrBiLMih7clsv33S
rs3PkSuJM461zcWB5lKQTtqOBCjODxwL9BFxCnSvQ/lxl+FKiuSUptBDaiW+JDQM5qnPrZX+/Oiv
/VyoxihMe/0UU9Q6my2AEoj5DvP1otRuSoJdTfHfv7/f0lwLenodAjjPOxZMmE7OXi9I8Vv89Yvc
jwpHSRLo4FgRqbp4ojTvQ990sc+ILJQhpuI6wBthFsxSavio3sstk7RmNwWHSD3MtQKoufLoHtfF
nepmGyIILZV34YPIWSVWrVLY649mjR+qHnkc4PB6xDdfZRosbvratkfmGTsOPZI+08isBdvkT8y1
E/pfJF92UryBD6LBokoP8HHAaBr/KdFkz8hTSp9cdpX6ieFXszYxqNp2gNoqXIoJk0q+XJu3yZq+
HsvUKD81MNnX4QxSo2/ErInU2JzMA7yhuSvZ2NanBuBACXLA+89VMHq9/DG9w6IIplw7nvvwxSpq
W7HJ509OFQVM931o6EQyJhLOdHEJEbCkd+CTFC2+gXlBzd2hHusDEivz8HvKvqfNCNJqhJmZwElQ
+FssOMMX7B7YbNJTtWZLc74pbhEdcOolt1pZBLRo6vaS2VYw0FFuv7b7zxo+Z9eVXGjnitNsscy8
f6m9tK1QxLgaHxPkugBptejxGzj/rwSpjkLfXvr/4giQ6u227Dshq6IZNo9EM886rjlrkemOCr8x
qfusJEAZeThfcqWJffnTL2icSCHbchoLzdqWf0/QYnGiaaBOyHYb+n5LWtbUPhACmRZHTAxeGJou
j0Zzz6186WOPzsVKbAX014HtuelZSuH0XBSDtzejPw2vDLm48k43FXg3TTA1JONyuMhpVlz4iKPM
8oFsFYoxxHPqU1XlH9qUYfxOweBKRyq2VFGwDj4ZJzVEVzHXS1hzkWyoJ5mTvY9y8dkm6xUnxKXJ
1DFosLizuzozv8cZTl6PKv4YKTw2DygQz7tu05pprgScWzXPBpQ6PUx7fMk8rRqd2x/na1rS5+wD
/pj9XBMAoXNwgnsYuK50NS/xfaji0e3NoqBxNHsQxp/6YPgIYyd1TmY41h43gdq140Kwbp4d5MFp
NA05hc+PPV8y/hSrjsh/CRQNJ+BQg8jNyCbhiM98xsa+dmSSbncTQyQJ5Vph0WOcA/W8MO5e+UJD
R/aWBts8cXzOBPkT7ewknmirgePSJpWOaBSJK4j59WrMbC70TQOZPVaGrDMzmkHgOIWF2pk1Hsza
/jXufjuk1utDUGcYNl+fTjO2HI4PetnXDGFTenBXCxlOSg5kER2B9YIt7vPTxR3V9M4GxIKrnECt
yHnDnUwbiGzc7pu93KsoUWXMETV2hIwjIoDD9xMizVKg7KZqvqxnjWaYZ2q+rnpTijqh1zzJv7iH
Sh9W7MZUeAJ9oi17tMuqxKUNuZGrp9jClmGKAICKwThEmWGxXIiDtQZkFI5gUqODHrkaSrI5x+gj
RXH/3GXKx0adVz6WFSfJwlx4NlZkUY5Flg6A+MBCRV2pUs0TIL90PYrLKRbMJTfTtkvM5eVjoFCv
nWlCirzzkejrQLR9rYjh1YR3TX9ZeDeryWnKoZdHx7OIC5UYV0DJxK99VF4GW+ku7KfSTUusZgdc
QkWYXj7iunz25drNalELFzjRahs+qKAo/kRrHoqCbZUx6TRX3X9j0L9DyDkdOQ9wWWZxkimYpysD
iIs/26x9MxJ3tu+EMCm6h5tb9DCOvNdL87sPQd0GQsZFrfRgVywd5uzLS4DFNuYbIcr/4sBLmzsd
Arq9KMtQ6+aAf+CjhNfQeQfoeU5/tpQgrwqlBqfr4ev+LteaM7Se1tv7Vz8KcfFjsBOK8cr+bSUj
7oWZEmP46xBLHovv4zZVSa7p92+gXYpRaDFOQr2sIW1jdOrccLWeCkUNKCGTCnn/XdjdZQ7d+hcV
k0dcCN9SSx/jA0yZJBVN/fiPf5oVEJ3+bPO8OUFnwtOjw5r159xyNlia7PVZxABrQ51GcallNf+W
yPvU85t72Ypeq2LtDQsUfwfJrnpsmjruvq2OJpBum866W6NyHC6nEJ0jN6WzAbNqMZvLi0nPIUaQ
ctErZYKyklXzC9+WQhOQ1cStVReaBjqrM7AZSThkKhLZeY6a6oAranfeN2rgttV5zCcDWZhVgBpc
zxv59z3KGwx2jAqoKCTRQ+OzbabjzILwoPbQPl/MMufuZ+KT5zpqXYI8aOOg1Dv9aJiveI5vp6jL
FBWOUnDGvIR1jkE6GmFK8U0igwqPJLuvr3jX0VqPXfedJ+IGduQi+DbsPyVai1jtKDvN5ok2sQHL
qTpkC5L8SuXuKXdUW5jUW8sLlXfJ0YG1NNoesSEmSyl78rBtcYTPXqYAF+y0DAPh65x3OYtXMARx
xi9J2eTqrjGMkcYSIHz7cZu0dH9CjdaPHBXPl9hEvZry8428i6ZmyXBafzRwj6+OVRzccPv4QQ6I
5O3NzxHlg/fOCo1W8gzJRqDbUniuLZXHzrupCmVl+45fU1i7xJWLu3WQ6Ce/m3mwP1KW1DTMkwpp
5E1s+AORwFfztdKSssBJSIBwCaneIgOXB3DRlE6aXFdJBbO5IBoBO+MDIXWkFkOpTZkt3tF/uj6t
u6R1j1B+ghC1+3tvUQCBns4ulNBlteHOKDM3zuqw1x1puK97hUdFxi3dSOV7aPT4R0UjqxDoBEMJ
W1gZls8lozLwqJZCZOvBFUdmNt9nB+qY7+xrDxW0Qqz1SfZEzdguA0MKRrBdCKIaA7nIU8o4xrhg
PlJafg5IJKd7Oo2rw1EkazsPGeHLbLU6M/oAC2Q5eSzOI4QY06qhoAthCtqOxxRPme3kQHE9GAzr
voA2AwlJ1aCM3fO21ubeRRll+CP7flay6O2DcZMQgwJZ6+OdrmsG1P9ABpsM76eODvDP5zonJy/a
ylqn8PbVBwb+j4c7IXQqaQSQPy2TzugFOdjbWzJF2kpQhgCoA/AbED2XlQ3zr4PrVkz9tbtXGequ
zpdIFy7P8INdO9ReIsVw1rUghsNyg+sCTfct2o5N/A5dE8T6aYOaJkWdLFyFHPBRAMvOTUN2AQ4L
9E9I4izCcDbot2kXj9IPwc0uj7ZEsuKxHBfB9SzDQeoK5uL7YiOSr1DtSK979ztKS2HkPg1DaZNG
iBRpluLKxy3P6n8Lr8W+Urv8Z0M9mAJKrA49ruuqOUDKHBLQft2QdFwF3C00nmwmtF1MGunyh+dX
Rql2dKlTQfNaF9DvNGvMakBX3nnNrjrKnhFConP+8092JQNSXzOn6nJV1ssHpNK/4sRFKhlWHrCC
B2mdPLkM2o6D7xLiFwEqHToIEF2fDbKhguCL82D1dVDTib5ncpYYOK8fKGW3QzOi6wBlwcfnZoTE
znbyZ+SrD4phkKp1jh/5HyEnFDM/1MdtM0mfhggIEanSL2ku/npnxxWy83su5QBixkzqwjJi8lwT
N83Z4CcgIW11uKYZ5EujbRHYJALNTp3BYkWaZo8Cy3hvYXfFuzmrahx+lEBulvNZPvupxj3URYvR
sfoKtEyKJl6RnABWHRxESZyCv5VHPQGi0gcDLwZsWmfMssFeP7GJuFQeVBDK2j10PzLoWpPjdohO
BckGsQ6ni4DWVzGkUyoiGlMdfngoEQCYpTKLyGgHG5TnkSu3/1M6NYNrdqXQasJPQCwx0aehk4NL
oHMyhjvS0Owp0zqlDdYE4iVJp2cBB8k9DJ9oCo7viMcnYd1hmS/ltWkEUgvG8ORdNAzcAWDdsQxH
P11CRYctqJ7hMTn2SCGHfCFjmUYVmVBKDUGhhJa6nFED7mD1q/CFYwq9MrJPB0MYJimGZm41zoF8
HzRwtaGENpYCge8VZdLoExzCbzJ6cmYaad+sDRVLQO+fQ5QCsSlBj52uY6HCUtbkMzDfcK6VMLIc
Z9Z4Mdltoe5w/UW3he9M84eqcsZ4nipVbFac5BOJ3ahho2Mn0VW3y4yNMlqEFWb1qO+sidn9hdYT
9wu3lCjvCTJ9BcpA9CYqDZY9CDknukHjq0SMiHG/Hhf3O3wFfRvwReJfunLoc1JfepAfkEKlxghZ
ohG1s+zH/7vnPithtWV2kOzOxCjB618LtXZ+gC54ziHauaC6FHJD98hQvUe2w6bNZsGIL6X7tE2f
T+V7Uo/vdVAXxAk3DBe0fHgr7+1tfNG65dk61jPlB8aunRKYDNe6cnOWT3TGDHqbbxJ9xOig9cnY
ZVktQn85fdaXLKUXjBx47ZoF6lmB4AB6YsnDPQHYjHVkTAoXYF6aDI7190U9PReTf5djQLTjzLlX
40hBote5aQgGlAAjHBS+rNtxT0SfE6d2t8qlNF205yvJ7eT1RIvWr6r19Zjeofv7WGo4H4HN8udX
3JQKNNQDsqNzix280bRHT59fMMPqbc8cWCEi/hytxP/AlReOXTais84zxlwk7PGsIJOzUxhn0z/n
4dG5ylJG4VFV60uV23m68yrj0PPrf1v7IE/Jax8S4JQr52K6ZEmLaqhrFfxKZgEcmVZkIE8a3KLW
79VNfF9zQSGvmOHzqKc/oxDUbnQzXlnJUMszx3gsecrU2LRvvvMvjYh0Bt/Rwz/pZnyTLFbNM44t
nONWBCeEjSbEb+iSrojSCQH3aNbZoCWU1rb4DKn4by2u3dxDSWmH/cJxwfP67MGJK5o/j7HQOGSd
sw6m9+2oSxkr1xsRJC4cmvhyS0xCDrcVJh0rWBG6ErumwUd+ZhYN92RVPqA8SnWvcTjEbaec2kaQ
58YHcnpPXz3Q0WMS6lY/8OG1kiHV1tNdgcspKF5Iv27ZLkzOs+Uki4jYbQI/9I1D3c7hpMEAXUyu
lrL9af62QHoLgfW5wkmaGNPRaUCnzB28dDtqNq+8tvuN00XXLYDCdHkKFvW8LkCS1XAJmOTU30zn
3F0PIIIm2F1bxq07STAmeJLzHRcnD2U2KiAvNM/u/oD2jmCQOWb91xENNyE+Z3R+Zh1E+T4YIf2x
3aBIoBqEUJjHHQuM6/AyC7DXWfJQk6EYdrojdUS0FjT6W1HhbYvopLCTlUWvqyUVsEhtj6VthfLW
HaPPVsXWGeAmeI9mxgND9o70Vm++pik0mNE5jyEgZ7xsu6y4AJwven35wqGQ6Tj5PT7xc6KgOqX9
hFi8vbF9bwkaG30hLMYDOdbb342g1GgX6POajjzZyO7DUqYvmMgj69X9qYqkmDBJCNW0o7GaEjus
u1buXjky7NeZgkBAKY0QNDEoG5Xbo/ozSbLSEKv1MRqq/GhPBHdt1+PB1f42qXjwWL9L6C9UZHT0
wgepWonfsuD63ajx3W5XsUs9EkySfC2ZMT1IQGkS3SzVxY7RMQv95UyeWIr6q3/rxevvx5YONdoN
vWJHl3X+3JyF9Q23QP8G4WJRVnQ6CDGD1Fs5HtLsFREx/qX2GLyNrRcZxuJEGCWmKKD+jq4iLdq1
9mRxyW6n3/b0xWUYnv3ILXYvDhvblclE3JSPLFSuL6DCG3gI1q1kLuPgM4uKee5jKaRbH6IBktXq
4nXD5OzrtwsAMSKK5NT3UCpJIjHhW1Eo57zcB0Eu2TIY9xyTYlfcIDGa9oeB0+onK/LFMJlWdl5F
UzYvgOXKoWRlquOO7HvJmMIxB0tZocV+BPsc8rE1sB4pKLANsHxJ2PJ/DOt2odiAOa5KTzkyw35L
r15HHLb8xvWH+xVUvWGCcso6Zat/Ukud1UjMVUY1Czwfbl7+0gjZd4YiozkNv/z4tbByf38aVU1z
qZyHnf0bOSKUV74qB2iquPP/oW2gPbRT0o2QoHVszJtkGkK/PhVj6uaJPTk24Z/IgOX2rKxu03lW
dlqeD1BmA15Ay/YBWW67I2nf35GqKbpDQQLOx+QAzYkoq7rFg7Yx63CFbdJsW3UEwQI1GVG32G/T
E1zutHyGYvrDGmB4ckxFv87C8JQm3272cCSppH/k7u1XRPP+LS4QV/aoT8x2XFnS1cPiEx1P5GYF
n0f1/gBSAsxB/T2rLSC9600sCaC6ufO3n3Xsx80VnjlCZEJzXTkxJuP4OXkc1MdoJYMTc0oVwZL5
1CPnF4vKK1akM9NK6QGJTOBkqN5QCANpguUIXP5wbo9fi4gV1gPhXGoiyhRmWov5xd2TZH5T+GsF
dTgBdm4wScogk782bQa0rh+GcYjRdpnZzGrYfqaTM/CFHWEPz5A2PqnF5YjtBT4FGXPGAmFwuvRi
tWLPhJj4UxwmPxgi8d9+U7R15Rqt+8CK1UzFj2P71bF/geReUcICEl/LUi7IktRNIx4LGYIs/xUc
6O9dGN/rUxv3gPLDkb896fj2O+Ou6naEmnpBQgY8Eqstr7fgpJo7siW4a0JNoDXg+1isf32mXh8h
K/6rk8qISGBcDRQrYJLKsyE0KWVgL+yRUgCrZBFz0bq6RnKZq7pWTCP9U/FYz3X+slORfPCnM6O7
UbaYODokqF+9j4XswejgXwi3u76GJrqM6FjISP27Cv/xoohD0BmxM8Z172HYgiD1CyUE4HhkJ+uP
HyFKGTKtOvR29XihYYlVVha+dTeLBUcNsz/yTfAdebeO046bci7Rl6BTdUA6bIvt5M9Ga7hLpkC0
PkM20ZxUug1ydICHddq0Lx7ovwwQn5QCZiEDT9IuWA3iY7hCFa21WcKHEZYGIFmp+i9J2h+vT10k
ZA6DM6TVTh+amqZ0OgiTb1XuErLJ4jS75LINHqXBgTPCQ+kp1RAVQQIB63BLOh3t5uLewu+Ct2Cc
Tc8nkksbSZ547HilzhWLSm545kRiPzggferGtwwcwinRGL5m3zkCCLUdf1+/2KSmIoSSxSrknSqQ
GLVzSySVE+iXPPuAO0lXzmBBKfaBk+XiivMV8kNMfFg5L/cglZoRphR1GWvMduoO2gXajhbryCnm
mXyIk68C2LdKmqMr2xAdw2hLfMkPbSuSFBE25qABPartZH+SNtiRylzP6b3xTVG6yMpccmD0Een6
z36lPnRcjS88asJ36NaXMqEjNiUqIo32OWoWN5yiGjy2Wb9yjxCAZ9wCsK5HAvR3yDtd1dMq4i01
UIO7btHcyr+eeRTptAXaZ+whh5rCKEe+EBpkdlfmy5ypf0gQJqodR/QFpJYxSmw8LV6NmHRbUfnQ
1AmpSg9Q3wO6ZpOu2pLGQ3qrRZofWXe2NhVRlJCW1yB+t4lLAhveTrsIafrvEFG1/9bUgQVqew5J
W7uLcY9tBd3qEspnViag1N18payCMj2CNUB+wIdAKA0kOdl2JqFU30oC7PP8Ax5A969uzU4Rd9Xt
VqCZ2jJ9/E3CBiPvpGSeqLv3IGKPeIFqN2F1W9GVB6tqJ5A3nxsPqxdE/nOA8zSvZc2alHV5kgXO
8S9urg/2zxJp/9wD5ANEYDAnrf6OZmm8cxc2qGdW1+qxAj5qxkReCE7SujSyr2F3jrVaAkCELML9
aYAJdVfSgsGNYioGq80vVrtuwCyfRxKno+bvKPtOFevzxKkG61RjD+iQf/NL4KII+nUZUqqMqS1C
Ois/AtSaVoYglApc9PfJfY+bvFfm40TLRhW2l0R+GzI9MBmE1uCdekY6cOClQ5ICqJuz7oa4CuS7
xHEtMgQhUS386fbfcnDnEJIzI7XRM91qFzveMulRbL02DN8FgaittxQ98DkDTrQAjxYGM5esIxEq
zyG2B7ED9xuYOLgRzWvBsa9FJlDvJTtWOLhIVUBcfcjdbX7kBf/GdA6rBjvZhKZCXNC0T584KEDx
4S+SEYiI0MaQUxunplFx2y6SLfszJtHXK5bPZSUq7Yq7N5OZ4yiDJTGK4CIrATFAC9UqpVpwqyNN
2B4uYZozKwuyNULT4cbq4Kh+2qW4SjlQIjX6ZLfVy9czKW5Aq1Q0UMkX+whlZaKTFGYucXEHynYV
DxOVmxz49J9cFUdBiVfgBNNavWC4sXse+rM0Gh8latIp98lxlpX7xi4beDeAYeyRLOs4rNKozf/x
NioDulLriQqtopE86brEMTCG+LWAJa6BhAeAZOWX81Jsm7+KuyI+Wh2w+WRfyD5HuQgR/KdOzoDp
FkiCa3QfwV8P3oEXj8v82NSBUH3QN17IgLEle0MopZArj4Yg6Q7EO1uxzQ+6TXck42PBoFf24Ah8
Xlr6xeR9maUox8vB3/+H2mk9EjfO9H2RkalGt1Fm6Ra33tkj7dSTpc8DcYrrroyziyUonoICMw6s
SU5WvgdWWfajQIi3SQOo0poCzAVpjLHOJ498C+uFLGKCySTQZV1iEI8cpCGW1m5QK+kDfhRHZtUL
TNozJ1g2MnbnrZ/9GnhA4+H/YW/H1Ryq36Ce36SS9RnqCI2QBrpHkQDBorW7xKbSHXtsKt7tCEbV
DU491TAxFlScI3Bux/ogJ9Uo5W4xRiayBd/12Lg744Djn86+r1DzHIGYMofr3Z/fESER3aZl0+om
09xSd1L9c9PtMsi/ThcKp0o3sVlK1P9rG5Yoy894ZuF3RR5cikJWzngxCOqv+l6fMwPz5QQf4WtQ
JAFni/P8bGnHE0GOjbKfykqQsBOKr208SqreiUixNG5Z7QlqODmL+rjEJ4CuPIVg7oziW1YG2xhn
IiM7HeprmaUcaiZ55G+WPl0cmLZdCqFzbxUMggqJajrB+VXCOWhTjCrEzahPcmhpw6NNtbn2h1/m
SofvPCkYfPYBvA8MAeMDWQcd4H7Kr4Q3mCWZ9yIxcHzFT3lB+DESdGOYX7ZWwQrevjnYKKfeDvGY
xbSI9e4u5G+dAAXwkmfJTc9RQUdmwQM4uyt/XIxZY9o2rbaI7D9ZmONqcF3fU0VYnZ1hUkfu933i
BvoWh9TfQsA0KX/H/kdmjodh3EqroVlmmewOS6yONSBsyIonXlUYwQgdQ9//j0U7y8S2GO9PMa6i
7dMeG7AiiwQ2mIxkT01q48Eh7iztkrHRD6eJFD8sxu+IhK+za4+MvPDkLICO6oE3W26MQyUJlyvX
b9c8ifMorV3IiKE5v7cVVn5JD4+y7/WDSzvIxT+uGZRWhn73uYaIaQjmjF8599+SPDLAf3dDT5h0
ZMwId9VPPxp+GnoDYlccgseh54JbCRp7dsOfgu1YXj8W8cB6CSXH+zPhZ+/KvHJSGslnh0op/nIY
JWj1dL/05LBPThJ3ePJikbugB+beofHPRRTOJQ+pbd2bcPolrIRiXsAxmvp6pMTu8hJHfW1OhhHJ
D02E5bIt/eyEz6C+r0hQkxoCAlMyeo67RlMDdOZaY4t8JBbzOkXCxorFHxr/8ZxyGMhbPfS7mzgg
kzoUI8NKcLlBbi1gW3CjG7kZHGT9HfKpBa/ZE9QayCeGjd0qapaYACu2SSjiEMEv+IhJm88EEKuj
cf5yPY9dI02klAq1wEFa76e0c0+8lCe/o33x7H6/TpU4UMjLiL2xO2669DC3vulAR2YkQlfAoU2Q
Nea0qeCFtUsO1x/iOMzzPwTKldJt7vJKshjjnnqOPoE7sIjocHr0w7qduK5ARXcpGAKVR8bhhvw4
4cIAohaZ3V1vfIgPO6LscxwQ0CFfwFNXkt0MTRg5hu3+lccb1Zz1JB2/6JG/FYxPCfl600oebI6e
qqPcSTt1tNDswZ68KbALoTfiEb+kTULGYIaE8nvY5y6FhCD3toMQUlJlD+ErVljLHXfx4JvLPgG7
aoxf77mZsDd6k/tcBKNBIt7mBVvU9IfC2Lg8q2odbyWtvpqXRPsqvDNbdhio9EvQIYtFNryZt3xD
9o/o2EcYCFi9xmL+uwIMnc13WArZbIgbqv+4GLB3oOTbJ1nhgmZhR7jgThes0mfTOvtJS2r+4rku
pUzYDhhI6A0lSgO8AOjRkaa0w6w6UObnUp9UNvbvZ1AVLm9LzF7DGiuLrYsG7bcvR09H/98sFS+3
saaHDUWZWy4WN4xl49/BU79tHZ12sO2mDQXNh7ZtTh5J3EMcy45UXIG/ZGri0+0B6JsPV7jggK0x
foxPxBw0lZDwQRxeeuQjU3KC8HCepAh0rvtUG7remXweEvCEDI1+d2jKhFg5Gt5Nu/dIkMx3IQU/
ojmGTsHpAMQhZtfzQ3NZXAsrhNyYYABKX2VrECf2nnkGlbkF8/sENl/nHF+/M2/2hOjjwLH+AZ8M
kDBFfbyZeGHoD78ueICMPXrkevATasXZlk1qTqVRKKN5qT294r1XU2QQ7bNVCLfIObSNPSMV5lJF
JpJddmFmtz259aGJ26ShwLSV8GMg69YIZRAnx+tJUl1G8qvhrVBMuzzoxjML4b7SpGYzd3+aoNfu
7myX/g3pukakInpIEipbhXK9+3OofXn+8Cw9iR/DRdXS71e5IRneaqncRg9n3xcSwUKyNqbyLUuM
ZLvvpY2oMMpnqep3ii4j46x0s2sH0bMgeK8gkEMNDMwo+b9l0VJ+qdQGt2lXsJa2QpecJkhp4q9v
P7CrhcPTvjBZB5jtLBIZTiYlJTbrlYBOJHNRHWT3hGR/WuRqQu4mVJE+bDcQaHdJ+ng/aqpY4qLV
qbRAe77FPdUYKGduFjA8oy/M9c5MPN74zRiIAQ+/jxX72FnEA14fCUnb+MQRG6XHHfY4VE+KZ0XB
ibg+rscP2Oh5sSj964iXvWfEEt6BNRylGw1YYFNsnesdedBxAZBrVnMgG/M4qCJb6d9rflQNiU1K
PfoSDvqjKaYXe6dLSrAPr/L3FimQYjHi9JVPgkpozMD8hCb54UpFW0j3KfdyyXheI8L+IIeAHUTP
6fYTGaoeWytipaxOsdUiPvnMinbGKMIF+MBIBTF1Ss+2y7LrhaYFHwdQLBH3bosgZ5HkW6HxujoT
eoiIhqTJ3D64Yr0C6VUEjTCtEm/atCSKpWLAiqkTQEJ/PHqY2q/fOcY/Xj4pIPJs0uMaXQH9CG7+
fe1q7GM/1Y1oShDp4Asdi+mZKKLTJ4X3suZLGbUY/CKv28MLLTIJny07m8uYZUPejcn482wU53sg
oqByU7jNzg9CIqvdCb+l92L4wV2OJIcOKWrR4hcc4agTbzgSi1pisFG2rto1nQP4WdnFRZXUmozy
0HrtqvGOFUzmD8QlCcn3kTMjRSZbqOYdylY7e3wVfRGMjdH0FyAbGQoQ1l9HQRnPV26+SUSPpE8I
8edN5jkmcs92159TUAXvSFH68pXw5+w1WBlu8X6Pf0jwq8Yd2vbKNUXwO2zmIVpeKg8wG19nuRS1
APi1eNqU04aBvovIBgPFOQ1MfDJjEphqKcfHPTAraesx0BNkmIq6u91Xu+zkts0ckfSY96FQg47/
8WuI3V5M83WAtM2yTZ71OjESycBbi391QJQsQy3v/eJJmQX4QxoIgVksrflZhW1/V5M4e9ykAa6m
e7AOkOLjm9PzE2iygtS+OnSpD/h2xYHLcldSBYtH58xmfoHX3e3rUQvXJR9tUWHfWDp0EQe8va9w
I7wiIKFcwAyZg/B/iu7Jt90WbY1PobAI5Rz8v0rREr05Hk1fNoONe19ep4GIJPxHwS0QqPCBi9Rz
4g74xNtTTWH7g0l2kTfX0x5JPSGcXJkVLXWqOdqmnmaUB8P0Q/PqI1jWkFxHzu4EtH28LO6nSkFZ
K6U92TWgn2fwiHSfsIGacHqFiUVBy9LxLKuuS9e1eXD3rE93dx5+WL7VtGFuM2zwBdYWwaB7vNnP
DD0yc7YL906ulmFsXjRQRisP3pfyvEYEHNV0rkTiFih+pOIWiPBSjXHeo9irikOxeJUAQ3jiwD+Q
KYSKzQZKLTwIFrsJVaVlb2B4ESN9WgIaUhzI1nzWHYcmjHuBPREWrGgA1CmQ0VBsl6aDpRFmiqCE
YwgIBRKAI+mY+1h4IbIfqM0QPOYPAOCb7T7G1cAkBIaz64Fe2mykOrgLH4bUlEqnvOpbfXnYT9sU
flOkssnBYVTvSdcXMx+Wq76iV9zwjtQqk+g7a+aY3cdHX923JqF1YEG6Y/iaNX/eN7puTzeuYSrF
XE5Oz1Uj/4SJ+HB90iTzDIejvLZqhVpeZ1x2ZeLeFZ2u2PVOgGjNbyKqt3vKFg0xf6A6b+4rjvFf
A6kFdHTtPp7pzuN2xbzVmyxwFwzaRaziu7ixWnuLMbPQVD/eVA39B/JIGj54Ib0xQ0nmlT+F6gEQ
OXj6jnhFnxkV8lJgko42U6jbtmdqNWi/ZPoqZQOTXsQ0OQkFPlgyooxBnm+YaOqCG5BTOCo2jb+U
L8s0+KXo5yEsDoShbzUUjb5p1lca2alP4FJJkhYqSSOv4Hrtsnn3pirr4F1b3qRwEQhObBmK6X81
1Y5VOKpEJe41Pgq5ILFbTa2PFHZ7BkK8+N3cEH/+qW8WJWKqEIRGKKRpSB5F1XQUgg6Y1Nhp96GB
yNtt+HCv9MttcwJgZXcgC9P3fyJ7GWG1wI1zP0s+/gCBJLm5vA2gOmpar6lVn86t09Kw0FDzsw/W
3uuevM40nipFptivX3IFRD8mtUWdkmUxx7tBWZ2LmAKv5dcBJPPaFA0zbUhdX73ioelM5kGzWJXJ
nFD9UHJ/5jJQtO1s6TFmI6b/PuZmB54NhkXz/0aof/NF5nNSlDvMt8KSvAE/2hBerZpTpAjfrkrp
AtCaXM0EFT+YiwhocEGLPa7+rkDIuAQNoLurYVjgNIBAmHED2QqDicz9OyvMVlMMHzeiA91kpl3M
24t7qvhbFse9wVEdjKndUDqOjoHuKEMj9xpOePgpwEq9w1GgWujYHf76twCIapIgCv/Zh9LGEfrR
MBF76TIzJKjNx1XRPT0Jgp34YS5uwJJJHs6ShWVhA9arEnXfFmpk1q4S+DGt4w127f3khcYt7VOn
LEKUVwaCzPzQWpIUbKWEbUWMbq5LCwZRhY2j49A9Nv2Z0vXtILz5hYNiBPjsUUZk5JmDBkdMNU24
sT4NLR5mk4RerKT326o71wPEjhqCikrvNaAKJx5k49e1Y6jXYI48qEfYeDvcu4bP/+Hh4yPy3Yn4
1BD5apPeFoWLVNVn/PUVxe/+k4gMfMBHwDRW4quo2M4sVwFj2X7ooXriSUWXGutNMW6sC7pbZMVZ
il8ttXp1GDbHVAzoC52ptA0+5WZpMyiazciTVr1zyhr5hwQ4L+rYisrqYvWg27ajXmINaj1XqGdx
4x+DRT0U7FX7phSXPNxD8yoVH/r803SIS5E+6C8MzCls6+o3p8jxUtKRogGXjF8+ivuyOYz4Jgh8
BCKGCnyGUygtSJBPIBbiRKnrUHQy+UnkXCKhZyXw8xrkkyzB+QmXtpGGCLIJRkg7RY1d+0JPdw57
qmxK6EU4DvdSmTJUIss0B1R9J5h3BJmuUuSxNutNq8Ew4O7C4Ef4IaRxpT+nSPom9K6ZM+xuM/cA
3KO1KhZad2RguzJKAGQhuJwqW6uUyqjSoXrAA6xUuKcz41udv5uN8HSW/68BrqU06EtNll7vVNH6
+bkHSMlQpHaaR6lkzY0zjVuGoqDLUpO7pbQLupF4Vrko1dOwKbSSMeppWVj3DA0VaSq1nLMOZFTI
nvMFSILFbA7wsJbbxb6mwKY91KpWtbJd1Bwj/YwOFSBgHNfbMKL0KMJUvZzfMCa8TxxMvwEgW8nl
j1UtaM5Y5LY25r7sM/z6r5UqkJkbmHL6DNPww34eporurZAEVCbO46vW6Zn8v2DalpqGSwVOwNGC
PfZHxF7JpPEJ+d0rndxlEBCsjwQQHuA8DgJsXXXlj5mtua4cWQjRDyJZYtRzMzkzHL3FXJX4vfUG
e76qnN19ld5OJWklUVdHseWIG628ciej52XgCwJSWQASiKfbvZjw5FsVm3fUHkHgNaZjdFrTvq9v
oTv6jkiwbiggilwmSdmLgKMhgTQ+s7559lSsPjCqc+oBifsx84Peei8+ICf5eKybe4oesjv7zDAU
GqFXCljvHAsfCiKxzNQYoNlq5SVZXu6FgP7i/zLj1x8SyWDteRlenZN9F4TLcVg+SkSG+ZzeET+U
pT6FFTdtRYQ5CHTWlqYeU2RyhUShRuJkSpe7Z2vSVGSWs8UaeU1dfLBjRGKJ3WItNKVaa9Tnq9Gi
Pa5CWFujn7J+rN57NMdqJ/J9ua0zky6COCLmmsAPOG97jK74YeWwk3448seX3yOaZUY9ICfQ/is9
/0awpfb0VrwKa/engYEU0IuwJ8cH/UxBDCBbPWmKI2LoEAaob8//uJtLzL9B3p0dcI0HumlnS4el
fgr3N8tJKDzt6XdcU3ra04BYRiRu3TsXYxDQtQ6t5R0PmwooPyCSbhru5HPQRutIhmVLM0ErAM40
s+lMpBWCqdPU/ab/KLDLEPrhxrj8fLTrgcTOrWN4dn0v5rW00hX99ukIFpcJpAS1DSELlZRgMg9t
bxRXOhss21XbqtClIKbP190LnZHSmFZIwQi8w61pssxlz5xbcqLrVDEikvrmLPFHp47A6xsJ5uUw
wTUNT5n7ZCXzrvr6TZVCn13sT1trhYvqZQxuraJNvvYoAO450/g2iXx+w8js/oAbkOqzjqpNZxd9
qyAe1qZwWFbmrY04AsN+RbyUs2et4HFq6CCE0U71ZjOq9xrkGwqIOz5fhEd3mssp/R19kO/hnz1c
AzBuzFU/9qp52w8/3PgGjwzsgIl77ROl3vRnbBCZut9uJEShksPaTf6BXmPePnFSBMudP116PUk/
60cGFYgaqTAGo07DgpdsN/jByv/E2O/qIdthn+BmNxAza2gdXkpkzNR9QBYViwzULuzdQoIFys+l
3MNwNMCmFVYnqJCEh3M4ShmG3DUAfixK4Cdsf0E69X4zJYinKsUzzUwGQkaCnSfar3oRJg33GWxp
fnzTNYlQ5jq7wUobKjX2l2GPadAGECSwLsah9Enz8/aylRNvb8+ZU0wRKYlqbmypnpFEZozPXoOB
Hhm5LNE6qkzIrtk29wehK77JqCYMSNOVarbCWETHTNX492/vsR/zvYRpv2Qr9VIed56419n22J00
xTY0MjeIcB9qN/Xx0bHb34FXxAPC1HNB0jTTPXBRl5Ql+qk8LWDPtbxzCbesoRlNP6JJLE3I9QkK
uZobn9jJ1fvGLpqoJrWm1fU269MIZS9g008prWoLGGtG0FO9hubcQhpCIy9v2olhMeGEoD6hgpVo
Gmzx7drSh3bLmVMTV27U0Apzcn06cjSRGD6qiNjkKzoL4XZrgN2cOid97wRIa0hARsxi+Ag12SZi
cMQBghS6nMolVvoiljwsCwV75NePRVJgIjSMUOw4h0yKECWm9K6UQT59YE0sG778wPLXTn+fmoU7
5Bk2Q8Fv7xp0d8ArH6j5GbvmOJ54W2E6UIA5jm0QvysotCzmh2ft6FyioOU4ZdCrGcIDyXJ+hoLX
r279uTkWUSLZdJvJ+0krWtPeia3aBGQMDRBWfpLc9pZQ05DLiuCIxY1Jii3WZk9jm8nVfE3ZMvAf
vT72ICqspxoViPekQhctKC6d+51CS25aYTjqPzuD0fWOeqiYmAX09pLObIbZaDXa/eZD50dqYqXE
zBsVH7h3k6MZDvaIgJ17T7kS2n0Y9yiEs3Qylbzi2t+6HVBtc0jNkBqhLagSA+2r2yjYSpuKVj7V
jDaRpIjAvYqbcOFIW060zjch35DH26OpNs0EEBi8FNlIOZdCBp08P7vcYHmnUY6kFJceHVwR1PzY
8HJH0yqG/ScQvw+fj62T8N0MFUQlMiVmLvVMq7yj3azHRSnKAZOiRXoptPBdc5AAf8Yy/yL9rJyO
LYj5mBERMCDsi+WIwOLw1uc6KswHVRxwk2Yxp5DRPJaT4LZ89rXCJmjugHzef8/AGuqSz3pUZx7k
k4M3sqbDa+6BzFw5TqxKabeBlwUxw50hnLjq1wH2dMWug9ZcJlNpToWQyHWNbgeY1kDvMT/VjeF9
GldZLVDwfjDE+IWgODzAXQvsfxyQncqoJDagqmB5HO0g6rguyrBbBmhK6QyLE4fRjj/f77Gc5jmF
mIm0vKwpKE/uLSQcG32/KzjugneeM2KUar1+20CE6s9BhvvlTa8xNSKY18tcFKghZcNohX7rWdE2
gFjSGCeKh4QaOW0afmYZcNM30tbYRdGq5o7pLv/xuTCKjGTqlUYxV+s9WG30AKY3i2zJyxucazQZ
jpkMN8XhiWdccnR+ZIbP+975rj0u4gpTxeZW/37Liu7cVZZfQXcXHC7cMhuT3n7TbLVSYUiv8jIG
tU1cixNYXjagobbJL8TQPrS8jTLqX+e2UynbE4iQOJ3004KMAX8q/T/NDq6XNmc22NtyWMB3AY+b
6PctsCn0V4xxDllJoeB/HOQVcMd85c+6AFptIwChNgAy5CcUYUwICPrd4knlLvIG69wA1lMSuvPt
qjRoQJ5CGJtSEEu7Tme6g1eQwdgYz3ODj62ryZ5IMvTcMCSHt0qAUABGZy+XPLDAW12Po0y6SCo5
NkoSh5R+wMkEX5PRn/eXUxBX8YqpxEUTiIa3vZDa6fUjdrVeln2D6Itt6amXs8I680zLM/MWRlRO
FVjsbx5KsnenygsqNqn+NiZfM+TNuRMPmgjtrM14UDgCBDt1QUh4eB/5pRPjDsAKXLXFO5MUhKYV
gsPciISVjj5yrT8/JLoLzrRcfYD4lZU0se+bBls4QcWdHo4Zp58veQXsZdadJk9DzelXttgLIvR0
Q/uhJ6/cO2bJ2xYMA/eKgnEWiqODUBy99EsqSPYKz+dVOY4U5qJp+HS4kTZAsnwFuq5HUYJVLu6K
AHSS+YW/GzkKyyRb6s0ZA5uYDWd3T89nkg9Jo7Lw1I6kfkA+mHXQSTYWwXONWIK+szeE2SvUTARl
iwQOFY3NWMiXUuSg6b9D3LlM2wCDMA1HKY+9C39U9RUOC+3k6yvaU1jQPvvKDZhf9W4TcRSqJE1V
uSW+dUsVntYGjEkoXSW+JQ7jsNBivRXWTj4xeFsl8/pseoYTMeQ0CXWeB7GXjrvBbz+vM9srGY4q
tpnYeGkZGDOVIaBWLVj+r59zc4lAEFT2mS9Wp54uiGJ9157gGkKzCFeQzwuaARec1ZktaBzwH8hI
U50TdvSVwSp1F/C+C0bb8GVeXzeHaGW3AKGfqkscLew8ouWLvmVbD/r0ooPi64/4hrCdLCtjRm0e
9xd24/l4qfO9TLtdWETi4O5AXBIfBWiYVo4ZQsDYEzFxI+tnCGp1T8FEBWPJxenLrQp4xPyoKXfp
qHlE1EpNzcv2dCRT3UurYIv+ja/vr9K15bkEQK0Jjk93M0Zj15v7ZbAnfEIZ1iVGv5RAEVbqmPDV
HsXdTS+p5NQNN+oXcOKbqu/MNzA/QZ3naReDcd5sjla8d+74RAJOlfV71RYbsEhJLoXX4VaPJd22
4yj1U5BKygRbSGFVornaoBraAoWsYe79UI1pMWOpqxAI2Qc1Ol8/cylOhN6KwKtGJ6ZzQsqRgmqi
3Ki01Cwq1+3T1wUKfI5NEhErJkJPA03flCF6FfLCquPcoqkDKmhbfhfj0auRyZYaPY+ENatWg0/W
pKHQJXm4L1PPjh+4B9NgJ3auoNn9U+BvkXtvJjvnEFUS9Ky/oMaE86tKka4RTsQv+/fHFrVBpXI/
9bp4j5wRFREERQ8xm4jAzLx+eMq7UTAGIyXMHzBSrk0bc5TnE5+ni1sLQVl2stvK2ldyHNOg0XKO
O7pXwSdRxX0XIOxhxB6I6zPrZBYigGYg7vrPHcGpuHYwsa6yUoTfRbBRUs6IEs5T7wcC8qnYE+E9
9FHbm5Z2fgO5X7DH+lUjCx5SmLygqSRifZ38NnLxM/dL0csoNS2WP/m5KSOLnJe6ZxCdH5PpZpyi
ZLqgJQECJn3zG32NUGi7OS/xY5zMgQ2/mnYbbBPzLzX70HGLUUr3WybVQ7mo2Dgye7edCpuBh+8U
jCL238mewBoEz/O/yGq8K+6LgEjp1LyXcoKpkENhfwxSqQLlJOSGKL8W4ENB/rsCmFLc+mDTUDJ4
fv2k/YL4V9A+yKp/xFdrN/6Df87wZIbTJ41ua6AHrmkr1FpHzdzZ3mJxfcsETUveRtPQ79CNeRXt
+uCmUfja5zDd2t+NaEHPjunRWWMV03OspnFSAI1CpbH4xpjHVvhv64GLo7XD7ETbhl2DF0AygSoU
ZZVJl5JZad/hBQP0bEcQYBMcU9bqj1Jnl4MzbQdnuYbauVa+j9TUbm0iHkUXyNgicGl6siehQauG
0aVELKBQ0L37dm/1gNCTUo0N2Hd8NzDfPZe2HbabJBTnvR4mwQDCI/1JMQ8MJv36x7APkGUVL1w0
OtqCnP6EcqqeRZdEiP/cFu/712yk9jfhjorF1JiVVMONJ/KB+pbfQBxix1ETYBFXfbFNGbTANSYn
1MrtcoG2EReyvIsruBA/cdZBlLq7JWDOzMiEap6vyKxby8wLIm7kBPQQC1yYIExZ1Jxx8r5ot9JV
bZe0+mEMNDxJPIfE4lGHvBhVr9pPMkNIhMGDjzD3hp1gCGGHW8CT+dyd6icR2mRlh0X9n7yXzMoL
ycsvTWH4NhJ3ju3x+9HVU3NkARcxrAhpNhC/kErru5m4CC/VqsymAmmwALQ/0qNQI2jsrjz/eLla
0bhU9txpH+RBRSobvH2TRuYDk4P3Ytbjyyxt+zKk8jhPFHvCeCz/46QrSRcjqiyfEXZ8A28WeQQQ
xc3B6jI6za/UPrS2YIUCGiB/LA5zOMtD9Q9gw+4RAv0HsRlKaVDvOEuaAabMf3kfkvs/X4en5T/N
2sbA1gAJie0/pCXYYtamQdiJOMRGE8x5IaGDXHPxQBEWBqVIuGqRhozOxV8vWQXP9/2qENbzUGQa
tGclbeiElKLZduKZgXFx+5MvxSIP8W7ZppnH3lMdTludWKF9a0MfrKI1mWwd+bRy1ANeVgn+HabL
/JK+F9EUyEA37j9U3KZNkfuJBVppetk1Xwbq9a9X+iTTjtFj5dKILoV2iLwm8L+qOlx+hryK3Q/7
11hf4AqSppqkRSwRb0t5hrtlTIPhH6bbswYvq1DGJp/eYxf1fdPSeGlnOV9dOBFj5cevGp3yQo0Z
gD7klv9/fHxw81E/cr2LCLcfie8OtOz9Emuw6xZQXDDSJADtdLtSw6r4G18Y4Jh9wvPo7O8jnRi/
9qiMh350ajV+OFq2+ZHG9z8OWORIulSvrbhpT2VcVrCvSeVDwTNvdleZBGyC/byW+0psBFoE+VSn
KK/WXXsZPzyFIDhwTgEANxFLrZBAxmQ3yM4uIOyjcKJqdzo3GKAvHcKKQU+t78nm63xJXhqm2/d4
1CcfZBgVr7iGZCvzftJtSqct7WzncDhBkNzRSxDpYqSYOXohjkklaffYGkhfMTIEWpASmGze+dgU
rq6Cu78Hu5oQ7FaGQtfxK/KF0CMNKOoK12K18n6SRt9hGczmoR15boHLSR6hQw0VYu1Rej1uJFsW
JcHS4MqwXX5PdPUZufySmS+nfXdodeAAwZL7Mc3tPf/3GSuTbdjk56PU+eH+ndC211aSQEbnDsTa
nQkRV0M8RLC53jjcTic43L5TjpWAih0fUSatDo2ZtmHHFV/8OTIrpYEoxUYXm9OkNEQXG0TVfS+N
ojeS0nBCsVX0WzrBc7OXULsrieqaVv3nJQL3oH6C6NRZdtRlS7vJG4Z2yMAepY02ZkpeP5rpzNTD
4TbnL0FQBvKNaH8ANYbyGvhTZ/Qds8GN7rz+T9nyrS5tippxcph+gZ/I4PFOhoRt1o3NA4FWx7Sg
rhDLYvPYYhvuqJFRKk0W5LUfOsXL6cRarRH53GleMlWjS19lYg1/RzNYrdIvE3fdBapNmVZTIwwA
rauum1fIqnkJd5b6S844soZ4bQux3INSL+2yIL8oHOAOcQmZQe8V8OlJeADyYCA3qHgbYTLskP2n
4E8TJ8oAv+3WEeRDIqmIaqxXegS+VeAye2eFZNVLJDh4C/AxvVw0/Wd0a+rE91PjevhrY1EKmvoO
y+B0BtyhDaw8xejjKGAG18ybPfWTJU4KyTV4ysUjcEAzVdj/MY9XMnewlVxV/58y50s+Lvks+qi8
otL++398lJdLx815l1Di3nlIGw4NRqI6Cf/kri6+WhpfMpcJ9ESZM7NDhvKFkphO2hTawGH/0VX0
u51GcUcnpa3+tfKvbQ1E5VjdNAoKZiTeihlc4mbQ+z7Jf0FkbR8UC70891DetY1GO5n15ZbHgJTW
IXrrUGKuciWFziFd6pwE8MoivQADMDF2BbQpo7DEHal/8WEpPPFxTvpcvsDcgV83WOIEpa2rcreF
FNvxrsoEnQIaHEOR4oWqHLRUy8hYLuwq6n1kRH1LWJ7SFPBuPuTz6CyGUwfeFfQdYblDwu1O8dGm
NqTs0RMm0UQJ/diHPqCBwkmXeE3QV7Yp0zhlrtDIQwxVnPpxqv7C94122XXRLeRz+k6fpJ+G2BVH
5UsPt7JbZ6oLeVKIkILx1Zm1R7WSLzFc4rGlVXXjtLrbMmATiA3rLWE77i3DtODJSIGpPbkla/Yx
xcjwX/OKnrQOEUEKNyh+/mlqtwz1pTcWuM1cXmxZDJNBIrBcNfkHkv19CTtce8K4VaZtX5o5oLdp
VKmgRUE7ScYUuKm3tstAVKL1eaTaqA4BK2+vJlCIHD5DS/cCN5aL0zrJOE4tdiWi4W8V5L/SJtkW
sDRtmwWUbbidWyv6LNoYP5n4FRsYEbMIGLqEn7PA3YI9VbuK8PPBnmDTZjBxvV1Lem8z8tEPTeDy
eLWNMpTFrJtElCNzdAjQoY8yZDSUBPkIo2hdhMMfyyQavb8yeZyxA+aC8/GwmC0Vl4OhXAJ4itcC
e7vAf5xhRKwVvKnyKDD1vfdBiwkpX3tjhoaxnbQH8CVGNF6FxcMcNpljtCu+O5htcEYX6O2qcBz4
jXQaTMuPbx0QNjTx320Z3p6H/or57NuPmxEpA4uwmi+FuWPD+eRmbrVwpA2821l2mxyuEhKPZ9wI
phIhPxBTRXpE+XWRxD9CtoE/bGkYZ9IJoNoudBr4R0Q5VMd3erDj3O9Hjwm+/0yVNuv091VJbk+z
aZghNcurnR997XZc+9tVqbXg4/UQl2hFCC/3EsmdLYyKptfkHpX/iFwGxCc8FQ7SzZMLR+hKg84K
6AWKvNaGUL4zLHFbPWOpiOtGKGYbDbLp2jUJ4TvurGLEaGt5zgUVFSYjuBcTZ2RGET5/pNOQjdF4
LQfakcjs19XP4V1teCnVH+btXt9i6aPoHlDl33HizutLRqP7pfe+TugRFBF966IJRpU5bDkkPEBE
kxTHXl3pM8I8/1/JisHke5GKPn+dzGQ375P/z35FGcCfkKMFGY1NMUCYoSW/NZVAqCzo82SrIRxM
dHo2DsyePEoXJ8o+qnSPHdNQh7Rn7wc3vEmibYeYpx3NfMzpOU+sQKoYVNGDYP3XTiZ0fZ1gXJu8
y/08XfaApLeqvArLEZCkD4FE2NzANOvurh6TRZCTLi2sI8aqK6SToWJHA8vYVuVm3/+0IETKHgiu
YPFf8UJT1qnSKCS5MSzElaUsGPpCHqBHp0H6Vs+Zv7/6nmxqWKheZJyE9RfNaIOl+4bLnZmsA5UE
/kXnAdf1yLq1naw5KQ9b9anlE839ZBISYGlsmGFnnl3eetC+qXPt0pV7akNP24eeYm5eh0nMIp8s
jLA8go3CxdlxHUfPTtBfsGKMLVClezfdeEaSO8Db/iJG72kJNCIrFVMo4QkXDGKQdr0h01THuGj7
mEOyeDBAwNGcTXg8udtes96gRxrnsLdiFNk0A2OMiX3BXGW8iaCj+Uo/KSozx/eppuZieiRLh+qv
Xetr+0ZE+c0lEM7ePBevHotpOaNNCGsp3j+U2lSMlvEiQVtXniZh6RApC86sNOIjt5Ws1ewrBu7O
ev+OZtMz1iVvMrM8cXN6ztz3WfroGoZRI6hDl5FnootQi7XQiJ4P/jB3S8uJdSpWPHXwGzwBB+O7
pnNXSjucCDXtX9omyiD1+mjGE2Uc1JmYuSUnne+VKG1NVOygqLtiBL/ZpGxL77Fh2YjH+trnb+sa
XQ2hiI8ud5FjtZff676JW57Zy/KNzdQ1jFg/VA9JaVPlP1Kx2kC5wO71dDABc1rEGn2/TjgkBzLu
71dQAtH54D4bObVR7+w77XMDtTexCg+LrW/gi+57RC+iazlCdHmxMY8Pp1fCJKCt3PgYhmrEAs8E
K5kblU74P21tE0J4xzAv18ppb/0AuD9wF/+kzei7wFep1c6pb6ytznE83V8WKwpgQgZFolIT9oWg
Z8Eq1fH9OVB+RPa0EqLO8wU8Wtjml9JWIXapPXevfiMS5zd2xgXi8YN0jhsU/Xx50FuTEaMONHIj
KSpXV5RkJ1xoBrRW3TwsQ+Wt8fYnmBEasKDS9AyIn139K3atET3YGYJCIoPUJPvbOsYqV1vd3rXK
UkIiLJ7eTagvX9PNJdVXXeDQANKosAKXNMhh6NkBInqfcecnVN23fMxGbO6r5oEUo//JLtuv08zQ
yNIg2tL8tGUT6le6ZqWk4vQ5ejd7gSwrQ0jyZH33z5sPqwdVJvB7GRN7bT4XwYGfiX/FTeTVGFVE
DPG8sV0Ak3dOax2PYPs0+/kFLZMSNPIrbQymav+J0HEm9EjPaoI4PsYxm5dkHcDy7LZ08lDqrh2I
rBnQ7xzgg4PkuFNXJA7SKKTWFlFfdkP98KwYgVTj4N+LLyK1lb2sx+rbqWuVBkDbRh6BQ9H8PA0Z
u7ka+e3PsrS8LFQuNqJ5wVMtxHsiSO8nYiOHHKKc0sxDeFu6S2DZa29eFeO4qH9phm/7iNBnXG8m
8xLVJ/c0Nra2nnXQWkiSSB2x4OKsfMcobO+YYz03/ad5PZTXPKUcQAutNUapE6pltp7aKAWalzYA
AeDFxI9Gys6dYT7iqVfPCXjCptZGvaBG+uXJkNoBh0w1jNS1bcU60ymy643Qu5+Ee5jf81VQYr4m
rfumf29lMmV16iIaKYuyxCJftHHuZY3IuP4I4DbY9Q8z+LF2lrOBzUtgLruO/oLKeJhlBTNYY2NS
Y37PgOJ/0Btn4WObG2+ckNyxZDx7jzLR9LPoxQk3vF3v4G0TVDY+u7vI4W3FdOjcPhVkGmtjJJBn
T6R2nzySNjjxX3Entd37N7jCTM3UgHrO/LPjo+fqh8L8HXwFQ90cefsxJfa3g7J/hzTVZ2Fv40g/
pjRKvtbvysIQKtqkP1VVnDjC71W2ZwU31Ep8PvuRgF84b0GlUabxc4+DhEdKyYsh0DGaud687BtQ
jkJrfTs+YbkiWfuhQ+VQKgGbxdhkzfHK1bQaJoF9NrzBakFU1NpTdEr6ITWk7XPTEES3Nw65Fk4o
YTHHbssH3ECKO0Ewoxj2YqMz0MnQbd/30PMR6TxwQplo6zpMMYETt7gGnSgz1TyB7e/7Sx84rU01
y+O0BIPhUyFyH/2mm5f+yY3hKJdeD8ymDw+Q48n8Ets2dzktrYmmTq0Fy2GhfVbiLIhP32VHrJmA
3mb9VXrps1X46RyKx6IHFzh3YcYXCgKGzmOVDOiTZwZpiRfyPNmdc6GWHluQvcsSY17RLymorenC
UQXLA2tD2ajBpNYBnjGpJnxsDFUECj/K0JVx3maVBvlCzSBBxKp+xW5mz9B+C0lAhXniwL707Yc2
nZB5IBz257K9RwRWJXy6PNVo2qmbENVhiSqVD6P1qCWFCp44KMkgKt9qEVd0xgMtkwK2bsOQdwZg
ny/GHoHJAe/PlzkR5H8C4YpTqDwRRRTM04sp6ELSAjbetCWIrD3+6/rsu2aQfbkhkt1vGoC2SOmK
UVG7TOpNsm7O4B59aHlVwS2tcRSekdK24cCcNeSDAJ5RRBUavt6VXhPAd3CnOZN/YoY6QT1RHvRJ
bQg7+o1Hbxywe1gCC9wIcCoAr4G9PQNOKNVzi65P2ud3Kpuzm+IFqtaNEkIXP7e80dMi19L+UsY0
b+TyLRqEV/hDJw1ECRpWS7kwZ+0HBOAwUmeXWL78aVhNj102QZuNC8LEnwPJVz/iNXaJ1PNDKW0M
P3tTHAmLV4Lcp+pyagJx6LFic1U1cHi8ffWpvHk/PRzslnMKCgvchbzDi5f9refagoQ/4BtyDuXe
qptTx+zYJT6kxMkF+K4R90XQkMfB0vmcjO9vlPkD4QggVGUtgQtpYoVZSI9NxNeIbK5Orwf9FMCt
1rzeSdbo1jp3LtoQELrtpd386cOErs18ZnE1Un/czv979ZGXARtT5YH6l3wb7u9g5WufO9mrBduE
Ryhsff2XVxZxfb4WbPLl4Fg243RkRgomTsZ8M9J78nxPdJSQJDtHCt6z2DTi8xKnz+aH31bo6FP4
E/E+icu9fZTTcJ4xfPE15RX2etFxu9TypW8wnC1oNeiV6ZTKmoaHqFl/zHaYZm2hkj/J9ZJ6neqT
se7PEjtxCL7+zTJnjK/ed5S/vcrMg/1nZUEl7OyMzEbGhHk5fJuAKZdt1z3N+bmPv7tGJ9sktg1m
HNkeFrARLoLsBQ13gKmLAg5UeeBvwKGuCAuv7AQBBuhRow4lKVHEBAWUO4WAoAa/WHZlJVO/duM3
/O3o6kGlA7aL1UBzsRpPbTeLyx5RjFSPWyi75wjBBSzyTP6/imXLB6iQt6WcdZmBKSODaBSIAlkm
Jnc+rqQNmCrR0BywJYbOi0anaBTNC6NjRLWKV0//7uEPL+/NRK2CoKMFkBoOjK9rclTzBdPSU1sG
aOV7yOMwsTNZSffHldB6zAFgd8g/o3ncZjZ+RllDGxgwWjPJvj0P5g3yq1vT89sFTCFqYjQwaMKb
8PeqHK4hRBQmapP6qlvWCH0oupmnkkf+SLxysFf/ptBxM7PtsVaqjAcVxRhVCQbcAy7b/t6KhBRy
TFFbggwubhguRNYZOKlDbeG+hz3eWK6dPaV8TfAu/gr8GSQUgfmpFNK3fdWUfyiZrGB/Egi+yGSG
Pk4HaH2O4s5zkS9K8E2e/TNPUF0S+S5pB0mMLxf1Hm/pJxVQMroJIMGZbUigYbxkL8hebs74iFEt
s6nJQeTNXd+rpfCTKR+aRMM+Der5RyllQ9j/RW0D1WcytITVEPLurELP0Sj3aXqki5zfyN8XeWPR
Zx4nRNaafJYm7/RuSY/yZut2j3PYcgJhN0d+PG2mP1QtsQ3cRklxJg24/RRqQ8J56TN4uTdpzKyk
pbfQKNSYDRnI+TH0J/yEEwL13xjDn6Oe9ZSaiRXlBbMglGEDIrWO7116axgqTGodPUgyY36l/xyw
camOOn0hMQl6Evsv2qP52VGQ43Y/3CjaW8LzyCT/fg/dGJRJg4TMU1sk7zB/oKZmXrRx2a2wZFoq
kdQjESpKjmekImRFpJI5gC7Bmc//OKPhEeFayX7+g42SU3p1mvOMY7pIo1VAE4DZry+YL1Q90icl
Z+0qbipQnGeXYJYX6qEfTVowLPc0zm7MHhF1qUQ46R3HK/kfGhB5CXV5XE42qb2QjCs0PVjEw1kV
U3hwnGuuIWIHF3azmiZeweoZIVIUAN7GyBzzE8C88AnIzMwYiQtp6M43Zbd/XbwRw2uFQ3nPL7T6
mVdc+ZqIgUA/NoBgsNuKM/qIG9kg9RJSDJzCOSenFYYfCt4yR0LtYfbDba8kKiNeeipE7sZdFUgZ
BWZmgKuGssJHu/kT0kRUblsNpbqPGnbwXShnUkvgbQo48QxcICwMBhf2uh/VQ9ek+EDk74EufC0Q
jxRxFxcqkne64hCUkT5Hb08vxhKRYvtwnPSM/tlg4mgEIDRBg5iUjVdagtNYr+Yp4E0p232jUvlu
2Ppi/ybM2ekxuXF5HmvNbi74yq0P5qgNYAWTh/zw1rX44V9v9L3un4g+QmYvCdjAIvD6RVF135UQ
PH8g5c2p84xxw9oXEdtZI0vFl5b/Av/Q1AwTULVpJgWd4Gjf03C4OxZKfzivnexdo3BzLn8sWXgu
tKWdnj85CRq4bVeNIqWzXuRtTfPF9z8AOX0VdqRYQlSvuKyz6l0r/hRpEi03v3kzk+1S7zFgBWVc
RSD4abNAHPotHJTUqYNwmKA0ni8plBgc/FXWd4880ivdQB82Z4p86/ShFHFJ9bkzB/dWekjUJA3z
9iHOp8bw1VqQfgh2POqI+VcouZNDJ/P0j1hBB9vtVi7hztlOs31c/JgoLSimkg+WKv71hL0TfvWK
8OQyA2PPXnj/q2E4DwPS+4jkX3eKQdzoP1533BCUqPkZOPWt2zsPvYLd8224zuA7chiE117fICNi
jNIHPmKP+hmbWoEIxxDwBsOU6e5HS8ASuCi8hEbiITPFe/DhTsNrWC08kpNfv9mNUPm4vf1KrDvB
Awq/osTY0kXZX+tPhFeHeR9Td4dQgp7RL2fxJIPGNqyyYM+4GirF0ZzT+i5+Qq9vgWFRdbD8tJni
55b4y/5UsoX8zvO1SM5MemoZpdAZvGJgNQa6yRA8JbQ5/QG+X8NNqYNAoBNxUi9sRHA1nOLAlfdl
hukXOfOE2PH8c6koAdKwwVxN4W4ZpLaGeo20HeaZYUr4JaAyTVAXlFNhnS6UcUiOYx0ScTbAEecV
VLRVRxa/ZcWM5YnbC+ngPyOheJ+haOjdL1ZV4Fwr/47psX/8zaLGZPHbVLe2EziRwCj4/uGkdZ2f
tkKa0qaWkJGAmE3WN2hkgpnaocbuUv4EAI7NB1p1RxnZi/UB3s7mOgkxWSqy7zxGY4P74uPCNqe0
ywqImqe1pVPREwd4MCra92DYVul7YndEPBGyyjRPeEisTZijgEhlj9C4LND+G8Y5NNJCvD8suEbI
Dowoc98uEV4zgsZGk+EGb3cxwhYIQ1/4tD/bUMopG7n52zmVs3sMQjHtJChx4lTiYM96qxMylcML
+9Wc+fh5BZykDJkE6iqrqOkjMuC+wRUPBmZOnBsLutWO6qkXIEdLEvJS3ja/CU1vZJ8rVxSHin1q
pWJRPUO8thNtOz7JRFZdONBF/JvZ1tOoXPWzJKDxQOz3sRFaWsTq0g2DWzHRuBxdM+HqnG5GM3KQ
r6/wbLC5ysd9iPde3dhxKlOd0IgX8hvEsyYrb9e2dKU32ctYjglwLFaZEDbreOgpQkP2MJR0zH9i
nAwkF7mU78V/DCHq5mI/Nmc7dHR4eH83l5nzS1a6Upwu4Lt+2+ykJNmstLPTdmhYLT5uXFEpeZft
8F0lUEso1YKpxCDMECrMaA/2bmckeiEO8y+m27L0OjX64Zh9ooHBQLwLWMC+QjdyIDrhHnOVe6Qg
izqAvZILS9H1zHYCu5jYPSY3RG41T+d1lDlo8NNsw+FTZZQhkts800Kf06mJ0oPXQ5H8083KBLLw
racG0Y2QAq52Bi6fkBn5uqVd7c02FxMNY35Mfo4GvseIeBOFGlK1Uux73u0DZLldfqaW5wkyJ8xu
xr/pksjOBnr7jLunWMjp2CFlkCdd2mURoHq0A4VAx1jGrhxCqk9jyfEZmKRoRwUSy2EkBQ6jTIoJ
c9mwMxFeds3mQWu9z/F1EjUMN7iVny4jOfY6LuIpukRkEUafctT/631gvDemLCq44l9rJTJKCYye
Dmrggo+t22AVYt/WCSvHwcx1Y9gpFEmeG5byxFfRLuKHAYaQo1B3og8uOdgW1Cet+iF7ajTmlc7l
kYevbjRcQz8I+FZaoqaGhusZ8Qy6djm9AjISNxphPsYz0PKmN2QIDaIxIFw7ljBYG1tsSEaj/lAm
rtuT3KhWGvZHQ/kIr5XYDMRAFRuSdIYi+E9dR470Kcnhyo5QfQHJL8kLn9y1v48K1Goc7gSayNcJ
qSIX74rm54sQA2vi09bFMIN2RM4HWLXFDZYgYK3bHzw81hc4qu31R9jU4kZGiTwWLSyHjcH2QPG+
0ivQcbipYlwaQDOI2t2FVMIycDojX/ZlujCX9Dm7ROsHKjkJsmvCWAbtEVACLmfk8DyvKOLFly+1
GzNpoFEQciWFM3Gd1FyPtFXLecS/5sQ+xxBdj0w7COPi33Gmweoz5YpqxpLUM9o4QOShPLzuqg8l
dy5fBb49vGEAfXv2Idc9xbZmRHFRAqBWRTohOFb67/oX+pBd5LaMplYoraqUOPFH100YN6BOLdZE
j49ErUp23iGb94aL/L5Amf9YggDWFmIrKCzQYWYy8ydqnNc7XIDWLYDJz3jqV4/htaRvBkWC7RLG
RwaHebYS+Kfkaa33NXa1u7xQtgq3HoBsDoURA8nXescb75B5WImJaJPTCnqP8qnfDQ+bBFbZOaSZ
a+azobHGsTVwrIq1Ti9numnu809D0Bs08T1s9jH3wSzGUR0U88PXnIY+t9yPgfz4JslubpUNFNzC
i4C5mFDlnkp1B0aAkgNij3c6C7JaNnQKptAm0FDQjLJkGodlNu8w1UVaepB0tCBiAtcUvbtH6bme
32Q4vZE7h4eyhZQEXIFlMYUQjDHiHhZygPmP64X7lJL6Ml/iq6BHHjXp6iliDlAhJMU/D2v8SX3O
OQzVkYsa+5B2biTPkkJ/Qxk3shBGnvMm4qW1S7wm1y4y1ASMAtFtiz4NCdjNZvCf0d+x2ePva8DI
LteN2bFiRSdDWrlREl4NtjMSQ7V1jYakZwXJmc1DATWBiU++s3GAhI7qhmvVZ91NbpmXzBip2tjK
7nmhPv5VY9eoJd3kLi/WQB9lf96iRCb6dmiWzSTmHNnDD0HWCYsnyQVg7zcL4JJ7BuGdsNtHn14z
VXyrMvkRNwo/LB/zgxHZjEnBlv+xAucwaf+cknMXfywTohyGGyQ7CLjSOw40WPFlQdNRiAbo6Noz
X1h0sCTPSkykM1WRmXEXo+I5TyWXTcWoBRNdUWBEGdcNXZblePhV370/SqbZw5QmnLUG9T0acE4T
aDQ1owMXiOtHp+XN41j20qGr3x9Srbfwt0NvyFUfK/xxvnj5NiXwZzdSusYi/upwGP4gD/OW0RwG
zfMtP+Iv90UZ3LkLeHpgVnCjdHFKtMISgLgUVriCzvkmeNgxEclSi/PBdv+5No0DrBVgaHT6qOtC
7aKQqf3BW52MX7KTj0QrlEcbPq1qtMcAF3z2iuvGZMBZRETpCQXAw6bhUwbH/qtr67pvjTZCgeJ9
bkEVRH1NkkKw4p7bqLznEBi0w8+U0q/j6goeWnJukPpQ0oESWMlUMzq3fwBX39hWXSYDWRZe9k8e
sOdpl5iRYfmFGrpYc+0rFODUuq1VjPYIB7PNQi7mdG8aWS2TwQyfzfGTGy4f2zED8Cpw9Sf8Fpwb
YLBmJ88gmxgku9nIwoZGVdAFOXjYyCiHVhhrxmuZKS06GDPrVEedqrB5VUE2MGkiOuMCNN8H9990
kibmugrWOslbIozolQWJqZbJisKQqs/1eZvHDUD7hAHtT+3cJWQNkEE9NrkUq2dumtQpYlnR6bfh
wbzs4FtYZNHSarooy9u3ocnL4P6ry7tUJDz+9Wi8KGYJWgyq20Lo9bsMMhewaw5G6YzGZTw6mJlQ
90QV/Zq92mSd77GHTygltgVqCjXe3syN2/nezo2U6I5u3iwVQfpZJLtakaDflD1jisfCEB/4zP9G
NelDNddsxX1Y+e4Lud917fWiH3pBbR0yELUeKJtjQjv0ERgjgfo+yPcGRFyGIgytiS0aM+SHdBFI
XfsEpHdVXulE2sU+fIuzOpFLxf8g6Hi4SHM3Cj/cUtPitEuadfTEpjlOtWH4VVoo9fBTyw8lsujy
ZBzGfV5VF7zi0SqaUzxNBFNE4a02J4WzVWGX5gnBXAGwYlgUT/PrUEoEPqjYDrAseQO27DFsqkFn
USWn9qLeww1deAQVaMFIY151CH57BdJfl2FqZj779hrWhths+3dvc8YYEuONJvSfN/2DHnCQF+pH
f36zWKVlg+y3rBgxA5ypzZMDRz2x4Za1Y310mxZ7FQf0Zor2DVNG7+iypx6NotI4m6vIVHj6lhyI
mlMbUGXyxGWLhxSJH3FPt6XmhnhVVXFu8l3jmNbVXsMTxC3brhYz7TqLr11p+hPyBbr7ko1voPvW
jFoPesX/xi5r/HW7Rku9A4EjfBb6actgvuFOAIFzk46iDIbfsTdLKcOAaLdpJdOobnTaVfleVqMP
zLrJ8XxdMzQJ5gF2LHJKXBSuFJ1nu4N/ayckZHz0b9qB6kYvBTotP+6nZiFPYJM6rhNQ5VGOnVSX
Y5HXEVgE8lKVKSbM7A9WgleZoBnbStuE2DGZgg0mCDr2DjEZ27FdxngenufnyB6+hGrB1Khy5ILr
8hgIjY9pOLLsq0GDRRRbAJ7sklktrVrhoQk3mjGApjWMcRpTkWT9Q9mgDE3dx5Nmx7roNbsClBpa
gMq2JysdxFY4efZubp4I/5HTn+Mqyajfg2rLG1EgHrswTSZhnTbPpdIf7NsXe9LXfVEmfij7a+Hw
o43pBHIG1KFHsl2RQUIqMGzmoPSSEj7qnvqNsYlJIo8MGm76jrzdbV/2LG086EJZ5Cgxs9E+I/Fo
nGweX5wqnMr8YBhvV6Ag/B9CK1iDNNM0y6vBkOSTaJxC+QUjU5yIWDmVrqa87bkVzjZTIv11bUbV
yvSI0W5kGFCv16yozpI7XURW26/cQ+t3h2+/V6fZyijWCbB08i3h8pNxo07TGG+zWMQIUhyF5c/1
GPWi8dgnB/3c+/A3drHQcVBt0MAMEapR7M9uMrQ5sg4dlmxEBozJaDsEiloorIxmE1KXowk1Utok
OXyJ6/d+Fv5oKwCWM3BnqBLb2GHwZMxLGirkCOhwled2oQLYU8iKHnzrTmcg4EfpAURua1NS0LKV
qYp4nZKXxb6SWJR7J4NXKZrTvOnxSY83HZcnvFU7h7SRTvA0+FCfGI7kabRCi9KQsG68LewU3Jh8
pj06QBHxmDlfpxZiW5AtxvCIKluMC31K5w17c0j/Vop2/uACb86R0w4ihBBqJcAsly4e1yRFAwfB
UW//eMWlpWGxrYu6g/htpOx14IR7Vk/U9pYM10tSB3A4+DOZeldzC01V7CLv1sXoCiSBAB3RHsvZ
Z6oOaIhZ7zRHy/Q1+6mQLSoo6TQaxWGdEXM4gtcsYi7ligW0P8/hky68cP/Yz5HGOz3EHLRc4/+t
EwJepc15PDPhgrznCwF9g+wzN3BHjPrNOeNAbRQ4D3cQ/bIeSGK2MQvhRTwLArb/TjPRTBnydZda
m92Aa2qMH7xIu149CpFNouk3waxDxaLw/rp+2wmQi90OPFUKysOzWTRWeeAyiT2riTKgyIcKqs+x
gUvG8fFV0Xgi41JxFc6SyUyrEv8hJqvzlGpRdYCZcYvyHNdoaOqpsRtkGkoMkRM0+lPTuYIpOr8U
k7BLv9f+uVR9uGtyyLX3B8rEOwCrtodYgb6K0S4jWMkqy/3wF+oi/HcPJRZ0N99Qu5HrB0WC/JLw
abeEPfe0NxjFUmQ4uOSJIgd4+OJKFa1a8YQ1XVGVBbJ8/r8Vk1A6NoQCybXQi8upXjKogTOxl8cl
RnCt88UhLexZRyrJ9jFm1gwElalnOJE4FKW4jTL4OAi7A0EajrORtvkjCLiF78BBobKbfWsOenUB
QlEfhD4YK1+3TwFpyfR1v2QP0fllRFGv2+fNoFDKm2q9v34/qqCpRzz/H1RnIZDW/ItuBa5Rp5I+
7I54pFbLxuSW5QuvBy9BhSWBlozYF9P/ekAY0HHHHGKU8n2knij0tknslkHe5zcc0m4RcEFEQNx8
J1tzZSOVFYx8N4m/HGGhp+mqq/S0FxxkwuHUE3TyU5zBW/Zq1zzFP2neWIdO1lKy7kuRBc2TEXuC
NnCuXp7ErJ6U2ac8L32iuQsNfxcQQY/UzE9M2osy5hDRjoOAx7hliXvNFF4x19RupfY2nzyhBaid
DUNU2G62TavrHwYAyvjnkqcZ6hVIr+Xs+Ue9uEeajf+WLlh+oFRYpW28ZtoWhHHn1QPYykOxJYBx
xJpD4m/HC/Sc8SfaUaayYxMQlyiTbNyyuQ2jBazHAl1pROfYcY1zyai3Zo3dywwzv9J5GJ9qUT9x
EKExwYKK+KaZXOEsIb1Y5Obv1p2ipX51TemJ8kqxdiRojHmj3O9xu4f5RIJ9+YWwOCfYj5dAs7Ye
eB8H6HVLwB9sm2qAEahytOxJRU0Dow4GecU71PS2x/8m3xMmIrOJPbtHwa4F2/oPw15ujfiXNP5p
myAM+PEGQiBkIaWZhoh6zPRHkli0FFTOD+vGTh9WMFkWIIyqNXChOwC/eOHp3ttbKROnjnHkILj7
/rIxRfqY2Rf5olwCANHmcQFJIxX0Z2yqSQwzMTZHnPbrUGP2kxp/eVjiSU1Hej0y+oFuoKQoU5DK
OF3J5DZSxVNXx5OAenwqws7oHX9Yiak9gooiznmGDS6S8TJpH7RrA+FO6jDXxy3Nkj6SqLCHtVlN
6NGjklpWfB8DbClAAtwblzdTQbRtmxs/NN9QHfDULN8YwUo+8/6YQA2RYBwJFDvAkDQF6RoTGhVw
Hf0ZBG2aKkCzyJV0+jec8iCm3SC5nVuIurfcSP489yJ+balbatOIanAEWsCZROlpeFZG1j8nAc8D
n1Zq5ngRWjN1eSGxh2oS6qtpqp4kRS8a8yfAmhjMdkmO5AL+eN5/hEEqAFVSs3If9ew8etdVJme/
xC2zc75ke9Td/ZZHvPxYkdOsZkAR3c9/c2Cooj3PAXCIw6lfwkyni0ZhUwulWiI6yRm5O/g5AOuL
Scw1FJlMswVGYCkCBm2/PgQg3Q7fsGks1yCRUYYn536RVv0PCxKHUEUwJNtHs7x2bIZecPdNohv+
PYYFsJK4zU5yh8DbxcwQImapQ6qVve98NwFIDeErxrhlOgtRxZ95GE++yNPf8eDH64DoP7gaez1M
1zWmB80cZF9znMPMNjr0/yD88nzuXb//VSzoYesBizZ9nCZ13lBb7C802uTqFDYqbBwIKI5P0avf
T+k21HCC/pic5cYUctd6XNwWHQ/+MdTs7Se8lHXLRE7Vd/tL8t+sBE3mqtuWMssAIT7ujd/B/UdW
KxxFkTri/bb+CIceiSb6bTcZotbLbD11IsTS5xuGIWw/9DvIaDPhXCT6CxlyJSr46aSRSS72kPKt
qOcSiA3FoLPrA+g0QV3lZeSYiWnUH9dzvQVjYi3RXl8sgtZkOpNI1Di19eGwkbGT6zlFIsn2A7Zx
p2EiBeP056aAeVX8y0c8UIP67fET+NeNXac7rfMpUtKrFK0oKm0wtFoyN31GrqGWZ57XllmwPZkb
eM8hAx1T/bCYPBYoYTUQTZvEF1LotHlPW675tc3AhtvP/d653X3z/9O2Y67h+MDN69AS4YcSUA2K
XRTlQN4SETXA2p4fyq9T2FsG5ngA0Ux1qb6PX+uFxWt2A4OW0Y8tss0PPW3D+zVTvb0Va2roLI2I
D/bgpO60Cg/QkEj8V6wpURT0Qftc/O5fSqBFKEbHaHodbWhbbBUbssQ5rxZZwlKdp3D8gmygGgKq
48HyS7kXVLIf2gPEwmdFX/LA9ZDPfNaK600/h8aJE53FLtaII73/3Xhav5evLr1w3ZdYYzbWk04E
3CLqwseeEJNaNQRqUyRcOSist4n3/rcfqoxplHBlmwqltLmL2hSZP3XIp1XPnkerrkr98G0AT9/Q
YHfzRf7SIeUZuTJ/K1MPR+XPzft2CA5RjRkWBksMsCOqRrX5EXh0UjvT3dyTy2uJZdiFPBhLHLvx
m9sI6t4TB0RkS3uD4s8oVLGwy5KpKzn9izAI7De3Ki/qXnBShVKrtAm0PuYNyMb3IHf6EwA8/Xbh
H1x5T+yLgDSOg7Fv6h8Q7ukDXqAXbZsux4DMHZwR8O4TM92cDSkYSh9i5SG9WyDPbVDjZ9jFAVyL
rupMgeYqf1UI555G86MEwOHyqTf3OaakUWWaR6Ysh8ztoogxZHvFJC6dhkhnZVRVNeXRkUmEslMh
p5nW46xA2GNtEcK6MgPrAQviaGxnzBvxbM036XjE3WXGfTCOIeHfy7Q9B8ZckFKc6Ef+c8Ss5WI7
uLDJYb5Vz5oAlgvsIBeFk0qPzS2nS9eoNtr+n97IZA48UbpxzAcJ/qPTssJeJgWDc4EcrqnZUNmi
VekfKUAT+FTIcCsySLUpyobNw96H66GtCe6F+Hbbbo5bCmM0E1F1wmqgkfZI7JY2nfWNNAVxxy98
gsY7qg8C4+6QKyopk1NWLvie05RusACBsdGyjU5oE+x1zrUL/LVYi+WBirw/auz3AXLzBz5I8Bix
uMNQo9aLE5BVVkw4UNna9cFUpqqpScW5Z/hjXfgkQosJFWgnJr2JkwLErkE/jq9UXvR4L8mEx4g0
W6QNGcbH9y+UaWG9EAfmEYA+bERHMFD/DXPy5fKoz82TxIStlfFhVN3bDW7jxle62VywIMzQoieb
QUND2ygjqFbwHv5pBMkV/qZrkRP7pfm01lwhDlGNmf978QTNuLkp8oiZtvGVpZsWxnFNocdLVuQF
J9NI6VEtuhSazwouNgyH6EbldeE1fgPEddFAAfImrJ47j+xHlHqoRVv4Rd30TcyCvvFzyXoX7i8Z
Jmjp/C7Si16X55MYngRu+RpUDPXIbdkj+4a2YxqRou75Bq8ehT1XLNzNzkCW5Cfb6G3jFvk5qVTh
+dEL1Qen/2vPeEKOaVPM6ipHU22Y/rN2ytwQyAR7X/5+vuw8Ue/vHEAZIKEE1MxWTlqkhNnTH/pq
BP2L/xoG8PAPB9iMk3bciSkvmsTaPlhBUUnZz3EV2U+vy/LNWOaA1btP29Tn5IA2Z9s77THqrhTm
usBOarN6PFc1wrdpB2DyF28e/zcfsAN/LQAlvBsTvJ2Gt0HKi+BF8inU8s98DXHNyOSV6GV3XlF9
bRIlGD9sIzJYVgApYfnBddL7kK6iJdqUDi6HgL0gE8hdGl/gMNkp8oUXY3RaVQsPyeic+tJ7taXT
W1F9RWIEuaHT+QU/3dCoOpif/HyG9Dv5+KbaqBE6V2yWRwGiOpUUSU22NmkmPOJv+GFoKm8lmS8X
FEKZysCWye54T7pbqz3NQm5mmHJk1nfcLqb4fYmHBy8TnjhYXLt8MzCqrVEbUCtb6HKHAgaB31ML
7XliX3tL2wf1tqby4M0bWp3IJ+db6Y/qRKQAPW/Hwon9hNBdJCxiwRkjVHHIp2kay4zpTIo05fUG
Z0fTTKTrmin1nf25ORv85QcHZ6kFkmylWH+Dhe5m2ame1I7aJRISaJUeokyvb0MEKgdP24l4pMep
4ThIu0pRTDBIa5M4VpaSCO4rs7DveE89nRPjDQ1GCsv1IxiKLhAtPFaQuKxz6fY7o2gonezWMHY2
RJuDR+H8oafiojdUx7PWz29ghf5vsbO/446xDYhK6CxOMovjLLaMPf4Syqjr2yc0/Q0I/cHP24V7
oaEaEUmJAqiiCDKl1y9GA39bPgqEAnIiik7VrOubSnyczYt3I9IctrOnRl/HqlKKzzMYWcdixOtA
mvWoibUrIL25SxxAcy6QqGouxFKHogHcFYIu4q/S0m6PJYqGH4wbgsH1NQmnM64jPnOU9A/f+Hdu
57G9G6SA7kOyMz8R2kzalCvdlJaC0JWWkoJbMQJGmjBGxLIgW2sBVToW4BjlZf5ubUFQU5brnijR
dUNxuo09ypWXWBGxf0PcufXWrf5BkLF2f1MMzX6ZhzQSN4WdJ9DrHRg/MALLlXi5NnYvyZnsehBM
8b8XmxmFhe4jHnXYUUge9w45tEyvwZ+gntRRBSfJaxSOI69dEPDW0LGghzJNO0Oj9cgPMs28lC+4
BwVfNTdr0cRQdGPkT69f1YI59Ch+iLHarmHFcmaFPL9zBeBoguipUw/XP0HYSkN92p7PFJvSCGzP
8ELHlB0etcCazcEIiRia0GipT+jCjOw8+KPOhNgr+duEMa2VdhXXULXw9P8L/NZDrzaWip6v0rbJ
TZ9u3KrdVX2+Xw8cujDhOjA+fjcxM9eOazfBUjr2m7MN2OAthGKH0DlUI5dkJ4WCsop81xV2z7RL
mCNJc9QK31CWOON1lGrl/pSPPzSllsD2XkOWJ7xWadiNh9I4sWFTjO0J4W6RvbnhYZPPPo1xmzsW
jAH9YfJlT0aBrWEl7H7hECyulg45SPSbh62GRWxbLJEL/NVh0zvUbQpK692zsfv4WDyFEWXzLdwx
CJbKiCdr8/6snOLW5EY9CfOh/wgi5I0YGC9jmQ+0xkrKoCUOjypgtuq5gV4tcKERfgxf05DlaE2w
FcH3O6kiIW2MDSnmBrT7TLLTfMdDJ1hwsZcyAfhqPE4Cm0/QpmjbE0hAPtqdQS47NQ9DMCfdt2hW
2PuhQQDuMlASaZ8HQzbSN2fky92WnknzemMvYp0uQgEdvHuWS5HyE+3XKbUqYmqc91Em/eV3MnWU
5+wQ+4qp4CdafqgwwsQqPJ4UDINkvG2xKJ6WC6+4Amj7Prn3YgUu5t/AQauLtHNssyi5al3Ewf06
WLakRi6Pf1yff4Zfk5ntBiYJrugC0Txl/FUIuNnA3mCYz+XnurvP1AmDKrn9VYe85ikR2FZKCtvm
w9BQSZcp0IXT+k8EOzkdoxFslJogPAJULSzpqCfVDgahayB9XLOu1pChVQFJ23SBY3dGLKoGeUsL
1UAmCdv7WP5CRiyis1WuVKdSePZUyEssHEfRiiPFn4GWWC7DLbuHAdG6DEURPdLtgMfGGHAoY9OY
ln4lmQwImg7IRm0nS9lq8dTh3HO6DCohENqOF0AvJuHLdzPVNpDkhaJoHefCgQ8YWII+/TlhXM2s
MyOnmpRb0ggxng3gxKU/QOAL6W/l8VOPUF32nsL1Se4CDxeE0HdeKtZ2zWQZN4p1EgRuLQtvvv9j
JQuhBP01q46Xs78MCi5NOuKiWXRtrcTx1XquQWZONcEYQO7XCdMkkh41Hf7VUFAAdn0lTaHYtn/k
Vwc/SHovgNYwKLvKXyr34qwbNo3McOs2eDz2GC2cJD5iLq/SpwASFM3wf78VFKoRze3HHDCmfSmE
3W6U5B1tVCN4HZul+eh6O9DEzv2j7FU0KkZTh7HGwy3LqvhSoLEZWEFW98QwHPmNl8kYB0vwltaQ
847euqYgKYyJbEI0rnmOBVC+EXAM6rK2apjsjrKpzFQA1+VBUNqBAxnQ977bw9ltc+PFaJGvi7Y7
h5+sm1H/Si7PnjQosUW0aAp8dmdBw/Y4nZ2wGsbRqsL0EZLtq5XQZaOuVtDDZku2RyN3jVNaglY/
4H6X9nAc0WfvSWbzTqKWgQokmwCV00pJU2CdpS51DjxDj9mYy+/RVdIQ0GSnjxJ4SRiovvniySBE
mrN1+d0khXuGSoSY5hhZ6yu9Dodag8d4gc5b29zcZhn9Dql8oRArFAcqMba7vq3c0qU9ZKgkp4nt
732zArX05hy76ixtzU4R3skMw5EbySdhGGUsA6q93R6ZaRYR6GvfLx6ifavYq5h7BaZ/JAdB4rt2
3CAKXg85RWbpkJ9OrPkCm+TcEjpMjJMkwpF6Le9EAo2VC8qDIl38z5HuBdNZLihR0uJC7Np3ZWVp
aaLVdw7/ih6lUQsIAwibMCzKVa9/ILW6LkP66I9kkjPDQ3RKsj0v+18oUoT7jWWE+SW2Mtb1igym
ein5KUiHbyh3Y/UE7iCTMpYX2O5G1DgZ8DBYZalLRI1XGtB0jDUGPWnciMOHrJ9iETK5/FX6HZrd
ZkIHxJSqQOP4V1iEehaJ9xsgGLdp/8K07+8yBtMoc4IHQNioJJJIDgI2jhJdzriO78d20h41qP3e
9KVBxl0+KXsBCA8uhjayTt+ztrMeXvNpplOFNoFxBDf7IWaKmTkZ2cHwCPsAuE6MBvcHX2HydYYg
c2QkGHjAACnu8s3D0nciSzBGjpknCKIs9C/F17SuVeCDqjlOeDFlEZU5fK0xxsvQsgG6TTOqsa/g
3rnePgEERmwWBZMIO7caxz7KuvJ+dkb8iW5nlr/oZUhhYz3Za81aKZiynv73GZn/vN1CtnUdssXA
yP5aOQqIjq/KyT8hovB7Rmz7ly84ZRbiy8QRJcq2SYcsmCBu1M/0UGGDkmuEcHeEE/3hWmQXv8e4
tHDFpu8z62C5tOc2MyCivGrIqmKOXfncm1r/0qpBC04LLR9QT4S3JPRQRuY3IuU2FlQEzNQbJhgY
pSzXjLk9l+psSGaDpF8mRCpJRiseY+sE2M764EW7ugt7XanVGMkEDxLZIMWI2pqzjVhP2y3TiNYo
4RkuP1HfbZeINLFyhcvjkhUbW7U3pimPboruE96bDJK59aD3sMQbN5MggGRtmYhE2hkPCu2P1KtV
1gVSuVEZbUgkYWbnWkB5ELecQwbYWTn63Yb9X7+SKgeNucJ4jiATCnLq7H2c1yfszU5ZIQw97Seo
3rBSqFppf62vjOZCsm4eZpnj07bU8wues99MCqbNjfHIb25mBG0u/17zdaktxC3adENWf7NpWdpE
xFpKZcq1lfTXzOgOiOrOKESByD0CLEbIp9jAvk3/JFtsZX0L3D0uD3eZWN5Y6UoUW70EciQB6R2n
cBkqlcoP6IF0dCBSjOeOS7KLEv0iDB5rxLR5AbhkIH/C67Zm+HtZWXNyyg2c1JF7vUuJl7NuZtA7
SCTdBuio09fjPG5ecRzUw/h27rdyakftfbcYa9KxrqBfhas35llvx+N6zCV9AFdQFwWMIc+qTgdK
NDmyCVZtClYK1PViWQfOwf4jp5VcimQgy4qhT3iV4CuiqXtWH2aGtQTDTltcJ9ZBxZRy0xH0Gptk
67OvxRPvo9vd/wtnJ0k5bObJ/EfwS9M/sJnQr6FXXruJNaM4y2pdYgmzlV0pfH0UEzSANUITL4k7
wGlyHQY/J09JRJbdUS6aeMCZqvEn8hsfHFm8mAMFj73GIIL1UDgcZvbYRiNwdLfSNyb3iiGd6TuW
CGk+GbWRuR8kMpAIwxRAPuixJXeLR7i4YGx7ppG8Qq1XjZWU3V+paNoJ7Kc/WHcRCTruTypAYt8J
enx5V9poMJUN33t7SYBVaUXjAwTAzsG1KxBPvH3D1k/0u1HJsLzbR50v/Ds+8N3yEk4v6zSLVf9I
r9PZ4unmvVLY7iIb5sUOP1bP0iL20lAzq9l/ZrBndIdKdmaX4hYgzZBX/KYWOGKyQmS/cUzT9x5P
qvKsOcqmBPdcKLXunLBfYsLZnX7iuY2NMnxbgtGTQqxJ5x2qUk6tzR/26scKqi2laTnWIzAIKmYz
TeN7NV4cdZNaSOuUu+sUjiMuWtICtBU2VAfc6AoGtoVVjoZdM9d5TL4pHuqnWLEdNEVImtL9u/YO
4xNbDW2KWe3Oj10Cz0z+QsrF7MSpL3mDRgY2ywj57TFuS9ECPQ9D5z9kF6ts0A78P1prTkO5c6Eo
CfAPdPB3UDqrXsTqB5TBCo4Pe/vggcXBZWAwtGpX/iCUEFrUDE4m8BAY9xPTv6Af/2nftYNTFist
YtwhAaimV+cHLxAPSXv9nnuPq5W3Pr143L8mcgRYaADou81XqJB3DTs4XbMrTGzKjFZB94FvFgFV
LbFJy58x6agur0UzpYQqpvQDQh9kNdiRY1LT0HkKag8VejD7AN249C2BRBYzOs+DWV6bbMKUX2Iy
G8bfdcQJ6gmZvgTcMGaxW1JvVNGg2DOk+frLyG71NWW3eOW9fJb7EmPDCvYiJWBTZlyz6ZGqwz9M
efX/DyjPyI5UJcIexl7Q7nJeYslXqdssMn6k7MWSDbfo/6kd4ZClCLZM0hRQH36O8VG26D5sjpWd
Y5Lv9R8b9nR5YPrXAnOE3Hc7c5gAeD1KUPlbqLMIIR1j1EoJJjPUkPEofybvcK14Jl5Egz2zOQom
VEejOIeY4PcaoNcsw4E7W42J9m1q44QplbF/9Izy3GRwuAy4RBRfqY3NlGOaMvzPh/WesmRpVn0A
NskQBW8uCIAeEDgn53CAtglBgYIgiBdVUC4iVKa6K9ZqDdrOd2ZQd0RhZiERMEHiwBXGE0txhwhf
lg3Sj39hNTJjtTDaIVrwZa5tIx0F9W+aXivoZM9lMT8lKLQ3lNMpcpI2sCy66Ju5vPyL6JZYnCfp
e7GrLIfHZHjWL9FY9kEhJvZBi84rPJpUlFs1nZzcnvav3PWgF6A2MIkUet6KAFjvD1608Nf9v71j
Z8vaIR9Rn9s035oPjQJjEUoBU/Nmgcz45lOJzpumULv0/uicnHfYDLVmFjf3lmRlASj45cfMIi/S
5zcAxlbuayyBEDJh7LYRUpm7eI7FBtzQElKos7CWTTkaswNAJl4RZdz0qzl1PsEnL7FWizH+cCnN
bkWu9e2tsSTRD0EmwbrevVMy0xzhSi/3/pLCFxIxnNpFxu0PqDcBUnmJd80bTOV0IUoe1v4otWpn
JJIfluqBvGbKOEi4e0h2a7zEgEE+B+t9ZFO839qW2k2+isuDbGfypUn97ehwggc4fDHNrh2CsYGR
w3eNr6CRGZ78+5HLvaDBJD7BrRSI/h9wLRbrpHiU0NCJTRiv2EnrENXCfb/6ppLuPMRbUtGJ67ZZ
taPE4NfryAVa3poMEh9t8++wJjPUdiBWMBHZnmLwJldPZLSsOsygBEwpqOlDb1syH8xKsHWdFTos
5eSH3BI6luGHD9WqS4qVyZr8tUJMzPVxnGZMa588j0oIXxRF8u2yPPSvhZgQ7kgRmM5LlIszaOSs
Ey2tZcO5XYulstdp0WS6AEF6A67ibcV4wg6bDEPBnmOYWeTc25cPCcCDo1oWybat57rhijGMclHL
3hRo5vSkWO0FqiX9Nc+WB4wEREs/J/mq6x3cTuYYaaznX0MQDXUaognwrGuMjL6C/Rhn/F+Ha4m9
k4SI/F8E0Sl9O5ngpSPl0JaapZk+a+nsdUEAiZk2Bx1qKrAHIX+Ut/rmPlScxxMFj2fac1TSsKhe
Z0G0ewectXjCdEcagGXwR3slAZh84J2/w4Qm54p3hmMiBvjtPpcV/vIIKf75xqFzHZa5UrO2p3R9
WdnStZRB0+YFpIc3O21uwogEJ6Rv9ELtOfPFX2fUQddUhPLEZBX6Ybqw4gWCplTzzhs9w1QvCzAK
2v9nlcJ8sUzMQUZgowMJF4P7jAd35MqF6U+Hn8GGj4dOHAbBPl16sTnDPOO0PcSkSfFqdDnEygE4
AYDy8TT45e1TC9g3oKAzcZO487JO5QaJxIx6t8CWLDentvsaXnAH3Fk3EbP2HABmgkNv9u84pJ1Q
vZZHu+ehQiFHfQmGGyaLeNAFCJ//nXt0Zqvsde2iUUj7eU5Pg00khRK/0mIg5VBmiuEIavCcXHGR
Fo+fRGo2uf6bT7fcUGilY2PXz9wCpOYEo0pWn3FDtRTYYhhySu7K2hE7mW63hUDkEfxcKTP9iP+l
cOC2pj0GwzqHWTM/BD8zSl1+Ef44EGpwlFiqpb5LYsO4q8nQtwXdm8GiBnux8MnINySpR2Fylhen
9hgKTuTYdXDO01BLmj3S0EDGZjjXo7+v4B7KcZ4gmBZ4O5gp4l+jUl+24RhQ7uXQoIEVLfprl16k
4Tb5IYkzhGy+sBM6knRRQPlxudJ22/Ks6BJrGQlAMtXVIzMaOam3pn2yPgyVe80Bqr7T/c3fy5wC
HRgW5M0TJpuggDv9Rk8uGIeGQR5mduVj/3MT3sCmzmaiKJ9GfJ5dPc+gkUNZy1Gg03LLNsD8ECJq
wTiU2GAEOGd9VFh05B4itpazBuxCGlf43wQPLVAMfwG7+lO8eZFtFnzV35CET34DAmGK/33qePVl
3Sa2Ln4iZRe80YBbCv7v+xG+6V6dLNMiD96OkC9eW2EEwFVK0+5O5mSfrUn/3oyA3DnfvcBcNsYk
BR5kIOjMWlPSEm1TG8QKbJ/gYKGKhUQxoMW6CewI8uSlFX3x2pSb4aL50bsRrUncEttF59WBiN1X
MHH+s2mAGMmpwqoVVLcBZiU0ZJpc9CRjyPQvp3m2qjL+/WWOi4tnO0iT94qvV4H5FDF5yBt3rA/y
4p2TSpnHCltwVZ2uVe+Kr9RJOE7WaA8kKMuHS0HxmTMRtFGQf1f0TGgK8tQSxLTZ2VY/xbd2OTt6
re2gwqmO28yhc3KoRD5l9zdYjiqaS+iTsjiROKO/X3FCyomJEH1DLQuW40jhfD/M89BylX7HJ7Wb
2TgOwUcNURORRTdiiXTYhZnotU+uCOXyAPfa/kEPj6hlkSijSBejeclO24cvOWd0dx785I8SYLBB
32fdu8N1NwdnGSi/88ktFtCq3xNs+GGqofjSHm0/C/9o8RQBVQKnqGOFDKle4z6q2QKT//ZzqzpD
alcupGcTOHsvaFpjlaRxt+Pl9+7ct4fkIXHVVYmbaCS0Zg0t3YJC0ZqxI1a/yS1zCociV18MzLk6
9ReBU4a42A1P6TugKr5RK3B1IfFdzbB+Iq7IenciyEywixbl48NmBbkTx+UvOj0Rd3yco0IJEaJw
FhlYx55eNFGkaFR9X97VA+x1wtdX2Z3U8Ifp+aZOiF7xs5NRn20aa/Ia8uXZRq3k/Leoan73RZ3e
J0GazNY9Rj5PgZoFuXDzlUJ7jKNDpbAQehRym5949E3bVaKKAw/ZB/6pTNR0TOJcT0Vy5NY5TLDq
pYwoMe8fSr5Rux53Eh8AOcQkVmhZZZbFI0TXsckB+8U/vcZs7XOlaXdYFtOalB6muKsEbVYXLp2Z
6J3aIJG9dPcWt9NWU52JPV5P951ZdMGI8N7I4BAo9tlxaIsT3fBGO87yn1+K3tBnZmPP2dkhjEZu
tlZ+jEfSfztSKc4nqTbQMgoY7GsqYQqF8Spc04bOV7MOCRKB/vq3jBtaeZg1dru+wDLDoPDpMVgL
hRlue2WvXM+b4a/jUjETKz9WIGqRmnbiOt+5lefZ77La/f9AFU8Ach5d7U4N6NvmymJ1i8iEHSTR
yI6+OgafFni5n4Eqe3Rv4aB9Du5bnbIoO7qpQoVqLXDB5oJzaZ55yopNzbpnw7Kn6jJYTY3NA7iq
dj32p7eBgVweLjBYMLb5rWhYQb9v3zQUg7Pp9sDMP1z5KcptCZOClLHfuYqyoA3OfnzunVUFNoaK
qhD8XqCKdjqAP08inbfpOAtT7IzK5L5NvB5Ubdp4DIhZ9PnZDcIhgATz5w8u08oBSTqZWoL8gbTt
/fGavfoWup3MYneJ5HamxPklfbnqXNc7sGccKhXiqJxzVNJESfkEiO4kPa2KiNhyiL/lRo1baSF0
LqN5xg/udL5JUjNrKo8dVBSnZb/6/lg9mS8fqCHYbxtN2MT6sbROSqWq33pubDAPYZkBrNB9qzU4
hwXv1AeuE46IkXjClxMhB2v8VHV16zVH4mjvBMXQglOxZlBZ1ahcDmJpEWfUmV7+RfJLGWnuGbR5
1ic+kxEXAOxHRriit83n39UMiGaForGNEaXRrjVc5HwhekvxXTFKbjwpBl3fMu2l+TP/HB15OD+o
gK3xsCFge6OYgI1EbHJ11wm++C5eA214ftALPjvFBTuf5AaROJ97mrS626UdVKGoYfHgYp6DwJlT
cGI0/nGwPQYQmkZFu0yCZFM3Nml3akuPMIdKYEXIojCREOYWOATkoAMXhN0WEEm+DHwm+rgX+vLJ
qGqYErCVoN1caGyeXyvrFT9TPssHMMiDkDHhb7Y9BA6cQuzNXrtx3H8M5bSVsoTprQIIUTWCAH6D
CZZP/ULHHZGpMGGJI/w0RKRHNR+WmmofC9BgoLwIZvot5AmuC6c2aw+fq+1tZ4eBVMdOi7+oI0WF
pMcc0to/AExhDIIB2mnbpf1dnLKstt+cLhiQwsPpNRCVxGMB8AVsI/dxSLdkofcUGZAh8YR12KRI
ZU1RtYzcPcA/5BE6iIwUd+2E3SriVcD2gX5KLVN5abwElp+v11SAs+yQGjKNxAMpG00m1ql2/9KN
lvJx8Eo0Dc6xlybEbdftZw4L8tN3Dtl7uJPFhmcax55FGzV3dPsFsdnfDckOL1r+bJTJ+u9WHmhl
bjmx9AK6MQw1WBe0mPs5/dYesfbODIoWNoB0NYPZery32AuBKOA7nv6O9EZbZ8Dbq0qtFGkkrnBO
UCtr/WbO1BbZ3TpkJLk432Hoq4WWY2u7peBeat7jqPiOkyzif5KRL6GfpHSvNRCUtcB8+ehEXosr
8dxE7TpJ7Au8bKxplKJs8EVRtJcTSG7OkjD9Fj1A8F20u/b5lGrl0XjZWOIxCASaGEaba0C8owa9
Jisv7dzI/oRV3WFqXGVzdbhtGKvbcwB/1oW11YfXFgQgfXJlBkH20/ZGbV2EiO7XpQIjcKtE8FBc
ixS9JwGuTmWBSUsHt6SBGkSNSzXpVXs3Qqy9prpGLF+Nea7dRZbgE3J6lCKCIqDU79dvJ26Zs8lT
OlZQESuUyeSoUjyoptpGTi95Jbc9IwNsCCJj40AGQwoPCCe3w/S+L6ig+R2vpk96BBOpGuSwcZ9V
Zu6+cWGTZkaFsVF6zaZXPHuPyD4mNDd9i/CqZvouFjgojx3gRySTHTtCSXduQI+Q9orV47Bny5oy
/v6+ngYXBN5AkjX8qMbOrpZZKiPy3ukZvSryFtTrKtVoxuv7Xw71+j09klnkiz4pT88x6rm8qRS0
0uDAk8wEtYcBxShIFB3pFe9f3kmJG5WBzsxKFpyUAjLmz9KMez2f2DNV1QZ3/9Tp4kVlVp4BtSZw
2rscWzz6eQ4ek1lYY0QktwIg+dQw1eB0x0YQMUC94jFGP33yj3N4502nJX3fQZdjJYVlcwwGiLUN
jrZ3gQgJIDzXbamtgcEOy8g0tXFPPURL2jX6EYwVaGyHadnVge+zlyNHo4qc+vIzz99EZmdb/KtL
xz5avpDYGzAVTFleqYVeNDK4TOuZaJkKu1cp35QJa3wmCd4VrEWRMPZhALxW705zn1XMwXjjy/G6
uvTcO2uP08Zn6kSolZpdv+tGU+ZZydGosc5+s3VB/qSNhRKlqCkVjEODAStWDCpLKdEMXs1zxAGs
8WOnuAgRONeYYulhHVHfC30oiFhvZHU1j6MpUNk7Vqf9eLTUYzkVG0wvhRHUV6qPrcHhFztPil10
1rbbIVdcHHRA1ppiZNeKQzocKGAIof4nDN7Byzzm4TaejTn/KqKeYLGMeyBK/47lAw01nNGywj7U
pPFxv0sNY3/8yZiw6eN8aRHZm9o2JZOkYkejmvPHchzuHcZD8d5Nr1Cs/t+qs0AZERLhQ/3Uzm+L
P5Kv2C/j5LhPBTUhVzR6NWrW9K3Nmy5UNvk384+e1Kx30FVpUY2UEEZJpB23wakIjJHwPMsely86
lMvyf7JlpMVuZlJC5EzFB9AbFHafeS11qSb+voa78C7ubam2Jf28qlWMn4arpchZvkiS0Np2fqpY
EDw6eXaBNs7uqVqtg6TDrpaCIhtecl8xOh8ZNoaXoftR3jmwgI0rJroqfPWAxey5VZxCiy8y94yT
HVr2Qf/go5N7zWra7delZS8DKWXdHFQPy0xFJ3s9CukmV0wnSEuhqALXhiHuearl4UJYKOGvR6j6
82TlYZoV/HMHZOwhC3u4Hz6NY0i9M1ufWW6s7jvtTnnuTsQc+r/8dK4BP3LfwMLvmSUnn9JZBZm0
P7BFDI0oSDDlAJRCTXNJHdygejwviiuTqQvOQ8MPQhQONoQLyIjH5o1MP/pjC6SmqXrxkQSnf0/i
3830E/iH2bVMt8DGVfOR92ZNHeKUz74bU9Y50tocX1IXEz/Q+dNtb5QMpW/+0Mrt28baW3FrDP/l
925sxgtg7POCiMeD4/b1iqO4ZFgmVUJ3IGdCgSc19DWuiVeB/xsknCF7kWcGOF0l/y36LTEQVzjz
45ghR7/SQ3SGoS80e2VrHIqbsloVhISvELQRNFac4g5fRHjtLL9awwKQ6eN2uASKCZVcGzA3o7oc
fJAyBSe4eTRgtL0mPs+dzBgRkBLmXy/IZCsnnV6jns4SgkbZp9D5BiNMlLM7O1Vr8AFjjHaETr0G
zbbQStXZPU7TLG+jpf5WBBiT69Hu/ynAkSEEZw4El1jwd6unCKvDVk9oeRZXaZ9N2LHF03MasLAK
tbR+T5kpVG4yWcFo8JMIohgYPh8tLtyFm2SdlAOw1Qj5iQBi2GJShgzjDpGSVYM2Qqmgp8YC21mD
v+9Lyz+X/Ie/EXALDzjaOvNmAYse5KER3BRYCUkWvHeaa765SxfPPiU4hH1ghiY7b3HrvXq4nLcu
7lrAkZ2cYNGTh034KTmUZnHPDsm+S7M/GitGSuVudLNBwAyJfV0k9HYqpTVumnrjarxau80CsaOk
x0L6qlfBsvcmagZcBhKyqZEzymp9GFtWa84JiyCwxFLdRcXSwOXKzBREChXHRm+YR4t45U/K7SVk
xwIqqoy+iixQUUZxrk/MyvHeKcUwhDHA7TsXEvdUHvbn7yfqlkHcSwMot3ttXaLyomvfzYG0gc5n
uI612eJk1KhzVX5+W7vPlGlm94pXewjwxI+138IGMFusrOMCLvlYvapXZ7/iy1L6qZJN34z8OnL0
R1cN51RcAwcXgXwo3S0PmLmIpjrh5XP3kLhzgcd0fHHihpRUdT5yLSkQCYkC20rRXgKOYYVuuMhZ
PMSmKG2DvreFwc/nsqTNBLrBJao3gAC6MEctUu0QfQU8r9aRKqd/BwcBAEOQENySzBFA/hven8d1
ENmDdlr84MGfdCEa7SV98Clbdcvm1OX2xs1EeR0WKwF5YD+D5KVzDECNTNuhpRWR4O3Rm0bf0Y3o
b7hS40zFH3F9XFMf7vbjCeL+xSrZNHkNCrIzMENIumw6dhEMKibGJ90DdeemgqFCOyLZTtz70Neh
7YTnlSsik+HS30DDyGFd4k4Vg1FFWcFs1/XjrATqTeNIqwsZBgfpOoiTnOvhONb9bUoBFBuyXrEp
rPex5Q6AV58mVHG7LvK0GdkgfnmnTT47WRCcU+yxDOxrZukvbrva6glclgIUnjQf+Aa5Ngq2K/LR
JekHIk4MefdlFVc8Ezi3jbldhWa5GxrwtFT0RORZXFrZwjejACKp+mO6dG62jJ0U18WGJ7FUqYet
KMY/vm9Ed8LIi08Toc+izB2rHyAANjJo17jDBHmi0tk3BxmIto3XkJ8wV9QpsXj7OMCVHa0i2NwU
KrjsHz78Rk0nvneIX1IdIw2N+Qe6SszwA4s/f2+ApZNJcYbjESmTG5FW2bGuPq+fHyU0nxvHMOzQ
XE+jCEqwc5aO4GxvXjjPSEsyB+iRD1iBKUHJ909lY3+hv2ken5DePMsJJWaD38Ooa6YXhjtp7IeI
XKLV89uhaPmzU0Jo4JyhAuWzc2p8GfBpzwolhxXThrI3cGvXk3PYx4JZhrDS2Sge3gq86laME4tf
LIph4OhtkR9PKCrV8sxS6jKZodhxCgJBVYF6DM6VWu5UF+6s8RmA99rZ+eF2btw7vVQRFcjc5sDa
7TX9wRvGFU9wVwiU/D/s9W3ymub2n6XwRJV5DN2zh1ltq/VLP8anugJi6QpnPZ9bz5YPlobrvWKF
qB2EHZ8sJZIAIiJl5jiCGpKGeOC4tPVClDR0igpNY4aEgIorVI/pFGB+UXaisR/ohJWqTyN7Mido
hl+KNyjxtT8mgegSxWujseZ6/plJyXIrB897g881a9Lg0E1/DV99QzD+tTiK7vmFY+Bp5ii+PDGp
r5jJMbKZ84DVtiKpDW2mGclC7EbO+lZgij02zXItyU/Iwy/vq7coGjjMDsf4jNxGy9Kzhn3LskCr
ApFZtRwWfeiP0jUA0OqgGMnQyl1MUttJOr5wbkM7zzSj4iliBRz4fMztkYKI8SL82QwaG6eKnIlN
1kWYHFbsLgvC3PngLzu1JjVLOIcdrkCQzLXugNzAzG1Czq03YGyJKZB1mnsA5PzMZd9OMyiOWW+B
Lhz1zCaZV2GcB0o55yiR9WrbRbtAUMJJuCtf2/mLpizblQpjhMg008dMPolx+7QtBo3G80MFzNnq
v9Yq2LoB0LSOU6YItuWGkX/fkSNj7snEGEUFz48SS9VgzeGeon12j3wYCC4c7H/ekRgIf2EB4db9
ucwcmv+elALjivYFNLrh3wTQ+Bu0f8H5IHmLHDUUeq2h1HtiDD3UKdCzeBu0X1eTeqwSm7A71Nnt
kLEywDahs8PR6V+NeHOwIOJc6KaacKGBItOC6YPyOMpTCDiEKJyyj3Pt0T7ryP/tEM1pl2gRAVXN
wBqJ3MNbdPtz0AHoyj78quIRbye0AI40Fk+PBs9O5zw3/PRgHnNf+Gtmg1ugfaG4G/fevQDGA2E9
nFjv7s42+3JhGvmqs1Eli5JLfCVGNpBeed9ndXwTpRTqtQVcBgC5FA6Z8V8LuPzZQ0keXuIaDSKR
T9aTSkEnbO4ypWYghPOZlLuEpsAUvm6M3uo1vPXAHvLHcfCt/t8MuV40mAjbdzn0KV9/Uz60XrPS
A+AnyeZ4ObnX0OhIa94wKUNuunrT5AastuJVgBUfUflnA1kLGTrjFFqFpWZDuVH8hIqlJv8HvDFp
ZhxjUnMd0g12BAzV7s11xNv/nzPkvbpq0AtRIl1l9jT2dAlTMEaWhjnKQgt/GJta+IR5S8W3wVvr
QBf4bHHKJruYx5RiuFHrqlpP25EIJgG/CefYjP3JeIyjYLG5bMJ7eRJ5x/b1bOcbuDmLtclWpVKF
Nqo/JZaWlXO2KVu5xUGyP4hO76oQuECcYVvuT0INF6MZzl4p0GDCymjR1aoNsU+Vq1ki8/0PPjyg
qsjPH9y2+IGkKsX+XqhcUNWh7SbIpyby0PpBMP1fEOfkBHoQgswKkivQCeMEhekO/Ivy7V9rY0Er
YrNbXAk73yWCQ7KdfACeHYyMDrwOiB7JzUqiVphmTCKmZ1yc+CzRqdNzKZhBaHfsASQLHZFKNfKQ
IgKWz7Hvz7vHYjchxoKUozCgY6AucETbNIg07QR0D8cU3amqNaHGCD620tHy45AqKEy7Irngvt5I
xxvACGlvD0sKpinPQHVwnIUCkDcG2w9+e/UKKksKIBf9srVsHtBTGjG7i/kVdPsoi/ms8LBi0xbT
UMt7vOgOfRbtvek/xE+Eqxb1PYHs3LNR4vqahRhEqjMgCPlIue3u+nyU5x4LJ44HtpBfuWL5hJFz
bb06pbAPMyeY9nYmwDyj8KbolmDXvYITaKw4ce8mabJ034x7n3wkJlu/7xcLjQ1x81b1/uRH1/F2
b3DFG+QCkYR9BLYmdomTmCvW8js+KGTZVFXRyqlROebT3v5qx5gnPako0bUdtXoittMh8wHPvV5B
MrLXbJ7q4HU2QU8c5OBq3fK3XtxBHFKAY+s+Dj8S1mPmRIqD3QY9nCO4nUm1Pt5oGb+2kdangFg0
KoibKR1FNdOWop1Z9LMYuFmIjGsfJXWqKPMvgg6Rt7NJu0Pb7nHrRWtRcVemuLjhd/Fw/cizI0Rv
8C1WhhlrhIIpSrdDh7oD6DAuLplvhMzBlvdFvndLAdqyFAYp/daRqGAuXzfN5q/ni6QTYLzy16of
v8GiM7W7xC0PfhACKb0Mxm+eidmaoIyXJmKm1dAKyHRbUj42TRSJmsVlchkNjqwr8EcCCAfGe2N5
bsw5fTK9eDJVJcBpYfT3Nt0xACp0lAEHTBMlCy82sf8+CdSO6Nr/AmHuelqdrmlMMmllIvLtvHQT
86q1h0G9k8NMxQADjNNF0gU7uufGzBOB1GSL3Qz7dAJMcgMNhckTpTpjtIQDUNd8TCuo4uptdgXs
neLRLZBdsBNQ7k8GQxvHuBhgW7DUW6YJEncDpZw0rxpN7AJMq7F+022tA8cqvqjvWvSBjif+wFKK
MYQLdvYC+SpJqSGV4Q2+NazcoMl4bx9Cn4oeN6QzXYLNDVceKYYe+KUIz+vfX6xRdCvRFyAS2UNu
eLlLnDAqNniF8tjHij6Zd4yKen+BovepL3fV8aj82mM8l+Bhe3ZwBnfrYohiqflUue2RD00Lptk6
h2GmXlgK+cISANcgawCmqI4SEEWlYnzzxX/VIwws+mtqWFIxXkoT7uUSU8XysIBxrclS3l3//lA4
3EibyYNODP3rAun6d4aiZ70dOeX+utVwBxL6y7Y5TQLc7PxHoLLtVzSvuUFdUPhVzfEVI4LnLSF6
QpKLC+fNlP3lzlLaH3qjnCxr14Mt1F5vJhzvQSRlVmdtLXsbTb9liGiosSGeTrd3HnOt4Bvjd71S
by8guKxujkLyw0GClJiLOO0zyCQoI7unSaaAN7rI9J+fWg7r5CybYi6g+X+XRSR7hGP93f94DCmF
mm8f6uS0Tx0lsQbAxOTd7dGVTceJAjuMwPgq8bN3QpSCE4pSA/TnaPGXNt/YcFV9/zIxIs7q/Tnn
XZI08vp9tQWfea8l6mqHe8jpAVgABs0vPntAatvoGlRes+u8YUB4aIp1r4sFfpC4l1fcnKXwdMzt
ppxeB1RRAp0qb+9Uy5DU0SuXeSQ3GOPM+TWsp1T3mMjTZcJ5FHaJ4hkGy+qO5ZSWGQ8lnnIiWBYX
K0VZ8jB7mUedl9YCK7bZurIsgeoflW4YmShzJdsItqGJn/VocH09wSYYzfThWu3jRgWwl4mzuVZz
2/aYFVQftVcxj+LvRAufa8dvTC4F5I7ZhcPsBowAhb2AXPDgID0IVbcpMDwS1/Ig/ho/JMsM8PE9
qN1wRojRdDdtrhutTNrh7Jq3Cibw2ExzCs6VZ3nIi896999giYWzhcynnmVw3y+8wHF5r73xNGfQ
vDqL3/spWaPCPWJG1KMbr759uixhLFnigrV5WZjB76NwX1baqhElJ8dA7uOXnhZzL16NcsNDlF5d
HgWliQKRRORBL1H8HkkhE4UolUl5zIdu+Ap7r9V1iBwb5afZVZ4o3k1cATzYAs+YsUDLlnqKIb+B
HpoPVqkB7XVAcV1hZTEFnNP7EMfJX4MjdrjcKEyMFBcPUFnNN+mZa5xSjUdiC5scY885eeMIAJ6L
YUpS3wLIptvC1JCg865pdKgCaUDXON/obKImZpT4h4+9UuU9pogN55wQK/LiWZjrC7+NYgLlaEvJ
m2HWhn6FQwn0ZLXHcZuZ52iOJsJ4DLqiqbe2MyHc2HVSFkqbs1bxmKBkxhbCAZ0oeVW0VFsW2zzG
bNOAXupCglVoV6f30EK6fPrWyzrDdGhQQDwIKZQHF8Y8v5MpkoUESH6Q7NierhljTRrM5y0OWVOu
HQ+CRvPJH9f5fEdIRQrkKvuXzwZeuht7nkCwZr1HTD6DvxHwxVYMUlvwNUKxl6Xj9GiWmXaH3E2m
vhrvZ/lMKTYjcumXqM/UznpCsJOwOeCMoUVmiGzRqdPem3022nO4EPsKJTpRjCuNlgnQg/pfeEYJ
ZaQfZHJA+u/Ullg18e+WxoXSPhg1ubKlaNIBCwkIwKTPdJpHcQGVuN3PzFS/mjZDekopS6f1Uk9o
9NQ3n1owT/lw/qVbG0eUSFh664ErHIsDTBFE1GXDcwc6jX9qKgWR5kXlod5LPXKF6CZloUNzBjPy
Q0ipP+lqh9QB9tQW4PtHrmFaSSuETq0JzQ1iZBeNoaCEY5szfimdKbBYASXZeD5nzwjwjRlacIzg
ubHPOo6AMk8PM3pO119KUVQgAoushL0PNx4+KMQiq9ZIg00r09FZ8+L0//3Ea/SXiTuE0qwaNi+F
73Durk/QBcyGOuEY0cwA6E0l6jSx0ij4eyuG8gpCB0vSBvfpDKPYClNJ+aoP8PFVUc2gIn1MWXuE
xYyJgW3ojHdSH0077n//pjoscdtt+4xdC4n3XFOeo2dQE6/NXAYm3kEU/tQLzJHSh6j1exvFyxvz
P1SAJofpK/pjURtqiJIY3q8C/CckATcfglISo43/pVZkKcCZWtY2EDt29pnUpp2Sk5Go5bIF0TwO
rBLdcQ4HEY9O4PfQ9ifE+hmU3Fi7A/gx0Lr3LMK+Ixa8uSUv9wFtHJkz5i5PGL9ji72T/C5TkYEX
zMJimDuH/Gl89KTxaEDS01oULZ0MzhXXdQJFY294ZYRfh8b5mlTfPzssdYaTPgc83q8ASlh0vN2N
rJ64Ro6n7XMOa8IyR7d70XfzOS4Ixxk8Id9Wh1wLBrt7fUTCe28rIifNUbDiti7HUp3eSW5lgkml
xszGleeoeSKFw58meLUd7HdH3eRwOOwcuRgZ0nwyJL1ES3uygkY5oOttQ0UyiWgcKCdLg8FtlEkS
UcOVXYqAVAY7wperC9Du/8fngzMB15OLpaZTtkgZ9EZKRQGxDDRYA+UkMVzGRrfpQaWTJSMSU9I/
lv4LwJpy4PTxgSsRNp3MkHbWwWK1wUnC10vC5QSKxDRfSF92SlHeO72hH1eAKyPOC1vDbWF0pQz6
IPrQtTq1Oku2GQQPJ57vjVt7UDV/3L7wugkg6GZqhnNj+K7ob+4JTOGsPsIuULHvGaKWeN+5L0Gq
k0ItHYcfDbo1WxOUeydFusCrkEvyKNSSlx8BnxuJT+M9uAN7eJwoNd/t0NJUZpP2tcp3snP9kDsq
ChkCn7wYJzfrBXOYjLxxK2ZyFcKzEBRpzeZNpxpiQK4nMTrms2F72mfHtC4bMKd6Y/9kKIXG2M1I
HdeGyJdJWWkZyujdWdspr6AdZSQj7Ld59CSrDCxfHRT7RTQgvr8acy3ey/zUnBBHBpFLkAhLctX+
VW/FnScsfbSk+zW+dLYYZAPtWaPhGy2kb7QULVtqypiWK9ZFkaoj+dR3MlG88bNZ9ZKviie4qWH5
FxL66+MjklaJ95pvMI26EKt21nBoB5yK0MFBf1rPPEH0rvq7gmO1C+Ak7VcGVpuB7qF/L4NfkA/Y
aOeAqrAtwrNV8Ts/kelX5JuIzCb1SAfoHW3HeQaVf/SOxNIKyMiEJ5Wxnhuu6UHvUJYVpEXK2hKk
ylGoGBPw6/Nh9oJdaFK1GHXT0wDyeHOpuWs2B/mFYWjaD1ueF9VK2ZGN1xbDgFej1wzADpMNy/bz
tfbG/3g/C0fIwW4W0NV+Zy5qPpmZIf7dbgrjsX8V7zIlLfMjX5LGR3KAYx3lZwD++pJ9RUiJbIpj
c4J9Dszu65wNWVM1ne//2oDjYYrtwSjKx/h5ISYq8+TJxT3q07XOSMk+sEIQSznpr7ZzNiCVLuPx
5a0/aoORzNaIQmGPxITXCHEe1B1uHv+86SiWnuJnVd8auZLD2x5vVPwXT1OcMJKCddThYj+4hQmX
Ql2m815ww4fgMikjLTYAInGc70pJBJBq8UPTg6LSS9rOY7d76vCIoCj4BfGzICR9b6ZyUSBur+BJ
CXQNv5ylcbDiL91iuKuLAt0JzVcpxB/VwpwtcKi9h3yQZVv+cib8HAcPn0qIkupD6lnLPMMnZ/7O
COZTSZY89LV/zwsImCi2KcMEEUMnyN1rQ8xgZDlwFGsGCDigdSgAxnd4nRjtem/5gxwtrJxBojOX
bLIKMLZnh0ZmXlk4/n+08IKF6NBPSTtjMyRhnYmHA8InHZS3qqoL7aMLuaN5iMxRJyMyDTmg0lqg
sxin1bAn1QI1sU45TE2pjtFehwKzw/UmaAF3hiRnGvOgoPSEcOe6ZOZMR1xb2bjJ284WKOK6XCEc
S3HTWzAo+7202KiiveXHl64ERDEcr4++GhvGoW8+24KPDKIrxQA5sqVzyL+G9WSCFpmkUsl1Eb9v
Ws0lAyAm/u32xQcnVfzTaC+oXpqA0ajX6AcM/blEy/kR3kpctWAvuom6docUBQGq1J0U2HUgO0pe
870CvMP9PamtLq+bok9QKLDrTiUChadB/2L1IkLhYxAUVewcn+2LW38HBBpNb/hYKBOKmUXTvhW9
o5pI30NaP2s4xDhhV2uWAXwjhKVGNLQzJLDQEyokjwWadaq478b/Sj/sZsFCX+puOgq6sZBVNW2F
hW84fSXULSkHVtvj2UVga2ggief5EIb8yjzQl5FznBWKtThHFUTb8SyFQpfnPgvTSLMYD3jeKr6b
nbWKneFXpHzQmjwbZzg/KMkuOPNz5y5P/x0LUumAq7OTAsMCJuJap5cKeRkohgmeH6ySepzD9Qu4
DPqytnnjkpKVEANG5Swi+jUWH+zXtJyk9lKlqQ309/fV0gP2zjeyf7g/u57PMn9jUwri1ticksSf
bOlhaFRYzTnUJIp8JrKCSuVR6B+EjULaOoJruFKDO2VMGr6wFGvFnsNEvZ0f7QBsLnBaXE3TM3va
CKSmtlgb95XLNfTuUwDFPGvbZ+NFMny+YhQDZeq042BfbWkrWXAue4R7kUorMPLfGrTJTWtQYvgL
rugqetO4kRX+oHBXMZCl9MbNEkwPma8iwIJmWarzgGMbSZH7PTXEZPRQ/P638D73I3S6x5psBuW7
+MIVIW0CYsEqHD6z9z6y7yNjqW3TN6mcV+p5/DELvvarrCZcIcHH48r1sEK1uU+7zdzjluD06KPs
XaSdbivI131vCM6I/1O2QmoEh2h/QxXayfveRWjKRdpv3NZrZft7msTsOGVvKsrsNq4UNb1bwS7n
KoPpjfo2NG7VChcMlT0rCwszUH0N+r68dldVT2hFeXmpS7bpvY9keog2AoEZhbwIZMo2YmfpkP6d
sY81hVUute/4cvjPRovuj7kPnQAY6+4K+ZZ6+RFPmRRHDeah0OhDfmXejyX1RNr2d8B40t3IAM8P
2Wuqo2fMQLhZB8eM61/2+K5JjOqsEqcNjhdsq1lo727U+vLAumWUBGB+YIIDjF4OIyVhqodQsAD1
/tgZGs8Y629KtSd+dwR1w9o4ZIkv258+0LYHIwKO1G78QAG/yoXlhkN/YzTp7GiDbEX90RC5QZeQ
xT3FUHq2pbLIJuBBRN+dMVgBzA+gA+mwwkXFw6NcPerDXXPRF5JRs/YukAzA1kIkXIbCX3XgRmcb
7ZS6xeteyzLcOviw6HP3erJOPWCRTBnw3ez59gOC9ne2gdAooSPSYH9ZN2N7h3Gqklx8RIF1+vli
PhzrlBqtd4gy/+reGh7yohP2gw2EfrxudjM2U+PsQzgBVw4pid6ue3SjUW+zPZm3m8NustntIrXK
/BeypvfjQS89+s7M8ME5IEjEDxrTi+Qbaznz0qj0BbdaoeTMf9Xm2ZkNcdvsNNiAsu8yBQXG6PjT
tgpXzQhXffAG/nOs6GpellwBEkdgIyzcpalSa+U4e93JmcqlCikbPOXz/A9Cue8sC6OCGa2YHKT/
BqhLLxVv1Wo2BYw+eKt1qz4TBsMU8+p28GXOJp41TYla63abFVrQ16w6xIfYo+eZnlgGHGUzd9fG
ut0er6TVYjYg5jiemgxDXA2MGfNpXHpYupu4FV834xN+g7LqFGokuL5PAoceknMPqMFG6CK3idYL
XyVDH8GUQthDxEVXBnLqHrpGoncVKaH+RjB1xKIzfFG8Ejp2IX2ESEkBiw8AZMOZpoXPqOCOTLNw
uQmGu8HZS6XlK6E+7o5v8irak1YdYrqodh9v6dQ4GG0rjbhLnOcmCszs6P/Nw5Bo+ivJZZp8koT6
XI4m6bgGUrraSEZ/bTBOX3pHSxwTNdlbX0QoSOuVZPdKwYi3dVqwlXHLPHSss97Zniy6k/gyd8lL
g/QNWfZeZzjFdbJVR82+lfgR2m3SJb1fWlyRfqGBm8sjc4Gs7+dc0u9M0gCGK/O2kbEZ0sPIFDZe
MMX7mIGhK+V5mFAF+p9ckF3sPoc4303sVUkzF9+4hzGo6JUd807u9ng2EqDvQIGsXCf6Zr1zKoMm
tgmVE3foEKqp3U5ICnXuXf6XnC2+6xGJNxmAP+PvnadaX79wR/qXzP36uV+DARMtOCXeCgypseLp
pViflvUeFLC/njjBqFBvOHdACpp8r8GpDTlhQ5hPdg8IqXi1B0zUReQU10722gX6470jqZxdbXzG
rwFsKzci/N7hs/glCine/Nx1WHNMGmMbvUvR3BFRkW5NaVGNnpOsYX01QjgvtTHrDWVFo0dShkWS
x0oGOQmmcib12TGSkZTgBI/enXzg/YVMzIptmNy7oRU5DDIZm+eEeRslokiOmkZopOUHOHDRSoyX
3zUEZFYD32IDl5/j8g8n83gkdCTQJ5ARPmb1frikLypN2pBNxpQHLOznRO/7qKzHhU2vBMdLL49K
WdKLYh0E+llvopbH3pQvZ3ZMyPwXFqNULiLweYz4YQYF0KaSV1oojTEr4y9mjvRa6SCDwJ/oaQj2
gxTVk0IeIQSIZQrAqXoKdQLp+Lscxi8TW+1XdvSjALstfMlGXDAEMFX1VZOuM6YGeelmmF2zpwnp
9NDPRzftGN9liroaMjmUE3APLTjUiC/kTHGQCRXWmxYw4uGjW9x1mHnNotMaqHbow2DivR5L8KrQ
9EBaQdRE+n0OOckjqHFbIOUSvNworBTZs+dyAsRM2qrMAh2T+goIHoGidSVLXMwjjQN024kdODeH
QwFY6wR9XOywoJJuTJWBmCMAuYg2Vd+Co0RmW27G+38e6TxmoHLl86w7TkxXPl8IBzXT/xn5xWNT
hiDWyabI0mlWovOQ2Fhw45c2akg9C/f1qVfSAcQ56A1UTeJIMwEf83qSwOPYZfxaQO7taTsSkHCb
dfmH8JxkOBI10raxp/Cvm2/HOIBwtR0jMxg87P8Y1/UuZ+bMc2tJiSO4nUPU5JHClqN0wzA5r+dL
p9S5Pj1CEnGk/dx8gGt7ofh+37JrAMSFsqQWupY6dVbwY/PnXQIBRTV/+aIO+DGCGJf0Tts8TUU3
A0hsTNF+9YB1DUTxLnoii/mb4/lqkmltMFRHVmU9KdAcUD3V8lIaEGm2yu+SlbgLxgq5pAy1whcu
ADBP8cTm92Zc2zSK/7/7LyF3PV8vME9bTlCfcZQe1HBMSGQLMnMSXC33YVr2X8Ka+EGmFDUwg9gx
29GJhNRx79Vdae0kDXOi9i8cZKAiSf93ItG30XaPfnKYaZ0pl3kTCnXjzGQPl0PFBSpcLp8gLI3N
FzXpUedXQlMRxMrbS02j9Jng2oSL4//CIFb0comY2FerjLQU0Rjn/WfhBO6s3kCC/XA2of5nKHmX
NZsVG4do58mTCu/gN8HBfy9cEwp4IUag1kW0kXGLGxUNWCRVBhHtS5LOv5fsMeq6iVsTVyVKnyc/
im3rmMUMR93IaYq/4jyKiUEAHE2iCMn0yflOOodN3UnVxBUsCUf/Nj0fSboeoybfsZKcPCISaOkW
m2At1qKQj7NbutODjLdbfSiX5IZKptebKSHg3d/yaQMVFdfltxGU0qrvQlLx9CuAi6J0rn0Ju7tu
NcJ5eZx5ASkGGtafVwz6vF/c5MZG/dS5gWV6e+KgjMHRdsm9CHsy8ewLq1p1lkVOTc30iWuJAftL
XXtRhTBiJlGmzwbduTgnwJHTxETiwRY3khfYPCBTtB3KO21gayGO3TKHLNMNZOvcYVIdcg3ApHFy
nQt1GSRwxD+04U8n88scGnXyTWkkxYT6gC4ylkKmHygWNH+BuPbELiVwyMgJA+I7Lvy5H0SdigIk
s19q/6rMOST6Av5zCuUXvka4Xv/Q2LBipzs3DoMuWxLEgPv8GCW2m8VpS9c3oCV79z83Aupp2uJB
IGW2EvjTiehML32+2ynhrsGhnLSDW0NBWBYS5yC74KtSNapY2jopiGrTpqiSIL2uWDzOmLM4hPYn
L1sz7xeksqlV0lloeJcH6glMuBReUWrEY9SO2cZlg6W7AQ8z7giw4oz57USmVN7AMt9da6BmuCqy
gGoksxxt4llCF1NLmH4IBAvtJ0KEH5N2Nwu+bf6G9GZROiFeqzlz8xVa50X5j/FKYM4IK99Bi0JI
hO1I7MXS7EsEf2VAGJm09g6cBlsUoCqcQGT4+5ch6Bm1eXT4E3HxXXRynefTXJgv8gyHSg5DL0nr
gVcPPy+hIyJxNdwKGTzVA9fQqjMYtLsuuqIfAVjZwkB+enNYcVVLe2m3AgPgDMEAepBn15crplIx
UGJ6bPJRpkWKTRvwIbZ78koJkBiMYZtX/Jw2Y0ZS3kwnwYynhCQVmTclA2BRNKetVKLkfVsj+vQq
fYafQRdUkiA66DUtw+RM+3JOAd9qt1pUDCS/UdRL/lRE5yfOH/x2VzlNjlK77cxPeyAA4Rpqnw98
2eZbiV4S383SA2fWWJnSh0z1sCFu0B+hPXRsWMF4HQF6A4gFmoxtcJo/CDRPeswULs/vvgf+SGwF
22U6oLNEvVhU6F8aiP9wf8Zs2lajT5b3T7p8YgZE02QzhvNR6Bidn7jTA4+ciXnBG09JKoDLER3D
cdrUJdOFVB47pXUh3zdi7Vht0NBRRZ+3f8ENDQCsknCs4Xp7Any4cGzB7wSEZZD6Q2QMOLdd9F5R
CMuNsB847ttmGIKjb8JlENx6kFwC2Xu8c+6p3Y1hiHYVVK1tCx+LS/xvbDivvXpV48eMmA7sv5HF
RmG7RR4CMXcSzF1H58nxgW6JtL98SZR1yQrhM++TVvjvSMm0goxkRwZG3hk4UO4C95aE/5ynI4uc
s44X5hYK+RnXCCWPw8oqu/EnkTqtD1/BxZpixG8NBVPECMdJI9hKaJwD0A6hRoaOwtUHDiHDOSJa
nNwL9DpuHip0MsTixTzf4JLd/Hfl1gaOwsD9E0LNUK8p6rZdSz5AHfHcPotJrm3+b9oheVQorZSS
ayQUsIcbQjWKDMAHA2IEAe53qKTacpAr43TjxAFiiuYhy6CMrKjkfGOclqDHuszwFQFhfqkxWRPg
WdUe5J7ewhBmLdYtM2HEyygisJWOCJLs5v+nF9vkAJokwmzrrREBqo+qbwC4kkGyf8/uxd4YEJuT
q9ZaC/3vp0X3A8k/QfHbSEyKdbvQMHeqqxDAOeaCPenZI4ZGSMT/vpsxZYH8qTMOGyYbStTtfP63
0AdnITj1I0x7EJG03uZStmBY65HxV4E1jJRtxTm0oalPafq0P8reBg2Ol0+ART1LLVvmmYxMbNUw
jRPQZ5bGly3/fBxG7Gh7HM4WYEz6ZK1B6poWw9zXT/Blhf3+Z4eq4oBotuutJvPrzxzNKLZm/sJV
5P47GUN71MI2pw7CfqTqp2ic2lpHRWk2Y6ZcVISR/XU34FbL5aqI8N9qQj11w964X3Same2xr26G
+Nc9ESIOabAqjN5mZ4b6WogPjStU97AyksagGCUA7GB2sn6HnMI9afM+0b0O/vqE9wfOltTqkLcg
sCN6KxeRSV8PyQGy0/tOwRF5/bk49gTlHG1VFQgtiifKZjmtD9oY1GXYUsP56Y2Zb06SMe/rz1px
t9Eiseyo3JzOzC42BA2qYYL/cCM97tOqcoQmKmcPp03j/rco0u62MTg7PMJsyoFEfjeULU5wja37
hC0kd3StQqLQ4go1MVh0xIH+DwSe7yzgkOPlYZ4kOhh5rFoYFhbXBwOYpVVZR5P+KGmXiyWHGPoj
s5dl1yUb8MThGNHnT0YvD/PkGV9BSzyMqjS6EjPTisiiqOCmiPeOXbm0Oo7ElXOkarBLe3Z3FUhR
D2cYhCl8IHW/gojIUnkLVYsYGPX9NOUd2+smW2WiB/mYpaGmcuxGkqkGsSxRqN/G64Do7o/XQwtp
ajnoCceAc3FYKWqB79lQbNacEgVugyEAwSguHShLLV6r/rinFh4rIsmf923qLFl3JRWMZff/zCtH
EhSo+k3HEvN8Jdip6dSI9ri+gq1b8cXi62tfwtsqQ4yOYkUCTxkj2TqE4DksIkKyv9hfhrbLG47n
s7sWA2CGD5Fbnam0Dl6UtNpgLgX/pCImKAmztahLB6ZI7nMlo/MHNKXIW0MYRxWfMAakIPV0PLEn
XjGCqsKth3uw4b+L+C/kceIFeMbm1AEbGQrmEgrglsQYCpVYrZWMvbUW0UgKEKDp35EncFcaHaad
QyvDoc9E2u9KMrkzIPXIOByQIpLiOI2wO8T/v/ROGaZ2GrKblSsKdeEHtYDWVqStSzCa/PUpwO7R
APDt2vz5WzMz6xf0LcTzsgzgYy+NchgMj6HcQQu7Ksb6lc1pnBwLb0E6Z5dSCSsvVfezYu5DfOQ+
85AQfmdgqfp6xZJWqDo+euSP4DxOt4yHDss1x3Ucmp3CKckCRT/wexx1akSsWVbbrhdilZpVE1wy
j7m9Ky5Ne9e67t1CE7LOVPCp8IZWdGt4kod/8EDevEM+CwwsnP+5ZqkIYAGnRui/QNkaWHmgtQid
Iu1AmGG6Siz2zLabw8H458s4LqVBC2oQopsGu30J1Tbuh1G5bXyJ7s/ad+QIGvcYmXG7Enmocuwl
HBHWEfOJ1qAhSWQqV1ijky/2Qh1eHvu197PJ61cjs/37uFMSO20+GWtlAipZPcyioe729yNYfn03
/Aba7J129U5Sm1SDQXNwU/cWNMwo39F6pDqWjXGH0N4ZvrRLaN+sEkit4FsL3ZRW13HIHSeqmMp0
teG6++iXmOC5FYreFNfT/EwtGSJSWcra4KR/iMt771IAKzHfuFvO766KrACcPsUeYwNQbInGwLeY
XmHHOwkxA/pZ0VUq3fnvJnKHHDus5umuIvwznrQ3uxUyGfxpMoBJfi4SWH6u+vGy9XJb7hhZ3nWk
acA3kUnp7wh1UM7aU6onVXMqQ8Md51BcuvvuhNP0FhdfmMFFJ9qmANflQfSw7FX45KD0w7inMZFK
G3/eoX+ghJ3RBwc8lArL8s1WoyzRWdKDadpt50ZWlBHiKZpLo/N0oRx+xCtVJJLOKdYhACN8wOcH
A6isvidW9etls5CHqyYJ87589+NSliwWYbLPIljTkC77n/2cyXFgjk1W7355edvESCR4YnwLzFV+
eQghzUqpNo/vviBWs2/+MIdgu3hanOIZ+H3eHKAbMRIViXn0H4t2vWyzGTXurDO1K/pf9ttFqK/q
40G2l0wJJ5DXx4c3AXhIvLd8AmOdoaSHcbUr1l6/6ni+QLS4s0u9bWY57N8KVIhLvje9ZRtT41oC
4/cB6HPqbeCs9TyTSGEmaBW6LYdWdEgGN9zHT3dl/Uxxg2Dfz+i8i657TkQtfx0c4jOHfk/5Kqvz
LayA5lzaBHuIzd62XBbMaQiJFfvSnoQBoWWaUawl3ZLtcgQThbGl75FRpJFVVktAfU9i84y4yqZL
bipKT9wquJgQz0X4Cw1Szb50w2pm9h6svp3qHtrU0HYAZBlwhzJk1HmeONIBgACQmWxioNe0tBFK
inX87eImN0sa8E2+hnyRhGpAntYzk6A7mXtVAUjGbVCH0RODcnC+McAD3o2VUgdaKazqBFq7uWDo
WKCfe/nViKZNQ7O9UOQF8eUwRdG+FfKMGAq3Tza0a8xbURHLF2807bLdBV/eHlKcgrwDKx8rU24b
QvP4OHLealYeYg8dh9Y7YMM15JgeT2G+LX3XwNWWV1IEko3lLQhQ/wnNhdpPXILq5VqVRiSkjxuZ
U1NINmkJFTmBZcjjR1YYq3MMzUy1hIxmmFMt8twUFPmpCvf+TzWd+DgNBLCz9eNZRDjoyq//xj9I
LfjyctFGJviPJm55aVVVBePp+EdTHTGo1hbQSOg4OXaENfKL7DG/uOmeGir6EtNnN3rfE2kdxmE0
wx1aGdlVX5eVIbsaTMjR2KT2wNplf/U7Bh4UKcGAGq68UzXs2OVf5G1KnWwaL6xgBGY2yCYTfMwM
wTu6v+9X/ofYwkNABrk4qWsK57RAwk91WIwnma5aYqHD2pD9vrP6M3V6fJUENaChlJRUU+mJybDL
uBa4BN9iqtCuD67g/xrnrzpUEbBTjxNQWPo2u8SzFMCo5jHDeygFQTf23NkO7kU0MjeOnyLfBKvg
xijYimIeAYjc93GTeiQ4iuddrthaZkxVqxLMWm6JYgP5B7eVKBkCVOHN67qyqNUK7x14kjrEgJxq
AkQ48Tuq8AFf4dA+lP9FNu/LkeFd4C0jTCeS5oOE4vXf7ZpFtqBo8twIka1nisJDhSlKStw5MkLL
K/KIfYwTFCEoQDZAILW7GSdW3rxB5Kv69vlEVSEIgZrbkEdVX6Hjfp7RvQZbqKrByD8pvHD22lrl
j6KZmx4XpDVaD8Xs8Y7x9Uats3T9bbqHDkOG2emjfwgWJi/OAhQlp5p0kAa+WIJ/dVzkq9IuFw02
5WXyD06saVklEvc2A/Aa697ZdytygjXxdZbcJueWjVA38B2GeDD7mQvQ0LifocwyHKyVLwO2KKRH
L3W+t/GMKOY2xNBobfxjxrGkX2y7w5ROn8SYlD/Y0n7OIXoDiAKIMxHphug37bFglW9JE5m/WcOP
yQvyTm+lhUNfQsKyUtfy6zVJOvC/u8RN2evPC6jk+u8p0VP7vggDh8ru9YJ5NnsDl2kspZe/oBdR
fftN2ndTNpeZwLLyCAnxb4dkuhxu69EINmgxai47ClHT+TdBUqOsYV78StlXRMonSRogNyCivtI3
o1dvlVqk9dOSjKrlyHBAiLPk6XWfZj4XwiokANmWwJVUuIAr6+0H9SEiEgguFmYubM9pTMu1yo8V
X8hJsU43RDfIW56hmytsIWqrLMWRSr33CEhI2y7D1Uc9Ee2sC604/QmbK7MZrJoT5R+u/4Au5Vgh
WCeirmMPw9apbA2OocNMGp9BEG636RxxcvDCA4h6Tn5A7RlnTsXMEpuJHU4PApUKOv5ETISfR1VL
npgm8y9yX9SKd3/ZbYo0M6oINByMQBRtkna1JgmnM1rBsFO0feZ7QMK5ZluFqKQf/2i/nOGPpWjD
DbQGE7HEZhp7cuzqDdOOqgRXBquZoYWxILswiJzL12Vf3YXDvRpmPYXM3ZLo37RKJ2D1UCvIiztm
T1+r8YrLa+Z/NzZlptTt4uguyw73DxixyFgDpnB9VttpAwEVyplL3wxfH0SKXvoe5G+TqD+k8pIv
hvw0YsUfwVgzLZwOY/AOACU69AFm35jGYnhwotO4J0ZE/Di9tPlp22Q4U0AvZDaTYrfJXBqPYtT4
TAyP8U8V5BHO4K22qTWXyxZ9igtHROsOYkxkwFUmshekKpvpfb4vsMZHneceCWMzM08fD2PrZPDb
gUeLJbTYV04m3baCMVwZeliFjsvKn+lYVqz6UTQQj2Tmeg0nTcjbJ/l4fMXYaTIO7z/01fN8KGro
lrhVW71RoXbHEa+7o7/Ce/9Y0bBjNRZkgq8Vb+p5Z25AntnmtokdStGP6B2dkfbxYTE9Aok45USq
zoFGHhiKQdKXsOA9ZwmPCrdipq5F7QLZV/0CxaByiKbJzLNUzcNZTW16EsmGcwsuHChbFaPkiwft
RI3WgYDVk2Tds6oiGfdzrvSQFcWZD7tsMHTNfsSXBjCWZ7o0zxa8YleNZdTcfVLkMV9M7SGIxPHl
Z4paZ+RAwe0NGZhyznBms4WpE7CyL/Ii6bprEgmBOv5wvkCcBUx+v+jzGR23WRxCXXIXFKVQOOjG
8bTSGAF1y/cr1NTOku/wQD5zRuF0U9wvC0XEA4i/dBGYjaHJVjK4e4YXpzGuiA3kz23kOreZOt4k
5pb8u8+LEA6nOSZw9fQ63jIpfS+5/JngFXZd8ehQdimxdRwbJXtLldMvleTnqe0qKhxPa9Rmz8yx
P8Rc6cBo0zNuJJAyQ+gsBwcscj8InbyZPJiOQ/4TjnDtbRL0mSw0wstoyBOTielJ2q1JUdLPnH4V
uEDn+a0ugOMdkyGRVXj+mlJX3eH0w+qElCbySQ/lFcQ2uhsGWZPAGYBWIgbZZ4TIEUFXJs5L0XZ0
4Smkslqq8StuBa6+im+TLk+2X4lxlZB4Qd0I1xAV4kd4a1lcF25CIHhVIJJN6LqVWKf3F2Ppgemg
7W2CVvwH1gfZLEXt0Q9yJbGi1rHzs8lyqqQDpYWu3xru+V11cb1ASAKv7CH38YOt74UHK+wdwScP
eX2qwZRSFnncBJ4rX9HLU+gcgbicXkSy17Rmg1QlRVNKhCXBAaElKvptgBLrySnV2rwHA++KS8zP
WRfDEI2PBktDwXwiwRy9/C/LBZU//ow0aGxYS7RD3be7id6pTB+heCyYGMEDrUgR56iIO/8zkPx7
B9KDx2anSFnzXpepyLyfLIqvJbhw64mT0su3HWjOu9xYDmxoLB8pVX7mUaER9XHB4V9V1XzKcTy7
s7vExVEl+QZWFVJaqUZ8J4cTJQ62MzZuC78kej8cpNHxFJUPGHiCw1avMs2MM8GGTAlAtrdeOeNP
CNXb6FmR/zywj0H6H/FOsRH9OyMU4JS4YsSwEq8SA28QqXJzsog20D8GwVQVTJMeqj3euUkJqDCu
0zfDWiaSd4Vxlr/SYopx6ZT/XR4TpMbLMtboipHPBSVUZW80lakA4wt1OR+GBljRbaFjaAxAX7O3
MwzGhTWuUfUD1yicp9CeS8EE1j4N/omgG7cDjy1LUPxziiglikh9GxKrR7PhY1XaAi4RW709rK8s
vFF22S0AollLUr8lhimsEo4VPaSlhz4Uoe/y3GxiJxt7Ftw1hOI6sDo6hC52KUJqtjQmLkCiqTKy
yiidhYrm9+A56exP+5DguJ90uPQwnB3fKGCVVErip7C58VtMvXxezXxClXceZFIqYShhQIyn5Pid
3hk2ZbjeXCUF/O7uEzATMc5MX0znWOl7syThs5SnX32nLYna6oYpjjEGyxXp+zY2I8F1Hy7K02D2
lg2OpmGk0RFlb3/z1cb2OoIkojNrL8XdiXDyrZkOnDIsI2jInWozMVguu8ABSKLrRJCX5SacX/BQ
gA4hblH6rVHfYLUD8+A3J4RhpccFy5sN/t2SLLeMtMauLSuZgO3FqyNVAbuKt3uFBJXNTdB0SWTc
pcP6Hyzau02eusGaxTZGYVpVjnLOeIst5rxamroFcqjKd5qr+KdXlt2fRIPfMs9SRQf6SjkiYKu6
/gOCOpb8lA43xr+HxFn5THPeD7vtAbVvApOY6MLrAp1Hv28J1jJaG2Rs3QGrLVun7eWiKcsASPkz
c1/bImycx9cB9grhEul2WL7oWG2Rf/4ZwLJ26KFzE30k0XiOvVP9ZZvyysKxzfObB3sSRdAzttzS
5rsqJsVvRorw3DendpV0RrCTe1Krt4y2TDI6kL7RWzM1cIiMZSAXCx5U4LGwSqdL7RXqPDdkX7H6
kXdB7hxkZ/X8gPwWyxq+aggkAbo3kbuOPeUEoYrB0xuEgsjoeC0m6csD1Y0s7H5zGwAvYN5G2GqG
XWHvypZlrR+k8Khgk5irF90HE6gWAIB3EXLx4O1Cm7/FQhKbr1FWLPS3RZ6mSzuHu3iHTlbtxjDk
T/1It8UyKGw2qOowmbkEWGvbBe2KPnoAThgK2HbsqL5UCQPyV2bbSmHFB8xfVG0fUFaVev5wtGgG
BSMrrr1ivYUkoJ2JHOE7G8HmWoKE11xvPQs2Wiz+PysffMEhOXn+64Vn7F3P2aEYNCQF26btok5h
ySZdYjidTCIPpPtMX9c8p50Rd5YVHGJ2MUFH9A1jREHq8zvl092ro+ykM/HwCc0/vclzyY69baeU
x+rZks0wOvjzFzXN+qEg5fIOv8UuqY4g0gfOqyAQuJmx+HubDGJyvHyDgIycJ3oI42CSEnxoNRUu
t3EUMVtioDhzm6tnVYVW3ynoPdHybR8FkXCpW6NF56M0w0A+1L5mxbX1/T3GQdi4elFWHoW3Mgud
Cdm77l78DAk1wFtBU/OU3azL2wHFhY47lGhbQn2OPgDlXhF4NAqZ/Yx2lrqw84/8lKaGvJ+V6+1m
KTULGfZOI+nsP+pfOgRGziDJHDMHi1DdftOrMfoiABLqMq2P9/r73GwRfv0vrlTAqifwpMpj8oqz
NQHapQKeLtSTLl6ka5aPU05e6vZOzbgaZGBs3wl4bLKyPO5ZOxLdGOEXOvfLDuTevo7LGqjsrW1t
OThUsAZM/zMytJS9U7gDXW59IVuQqNpoNhWa2j2tbCmY8fv0R+TuBxA7mNJkN2G91j1RO+YdMoKA
gHNDPMpu3vJDXp+fKgUaFp98PZHUIsR96ntA+hCttQr2FODqGoGtC2eFwoekOdMwvXmhUEk9S1hC
nuHp5gWQrsbDQyddVURBcEdLX+HugNExJraDzh5yo0YHQtNWRWk5o5p18G8M7VuwJqmgOPz+rU5q
KOBVCPBEkYqIDM3eYv/zKQ9E+wHOOZRetks0z6zckmXxAG7BAIkP4RtLAY5u5Clmuz4moRri42nK
IkxVehHV0OBKhGcy+4/ItlO3N3bdnYcSvslMTquGeRdLCbNmuq8Pe9owatf66XCvIohBK1XTDXVk
T4OSoqXyVTnki9DLhmKk2tlR68KAGG3t/IrihA1niGa6k4qv+InUS4nJ/i04GDm4ChcPeMCp6ew9
69kCci4GqVwfLzBbnMVqmPxCIovKNThPtW8UZ83i6wfkM+s7/p+yiR1BZ5Uy1qX3m5eCzSvfgd7F
+WVcKBmC+lHgOpESOc47JbUVyL5KEp3KpHfiYocj1RWklf1NzZtMyOZRhG94/5aEi369ekvpaZ7h
RTgDtnjPRUD9UraihrW0mTbQDYlItPbUYxQv/Q+PHsiu7fD4myVoEK1al2mNFWMah/X54gi+hvv8
IpReR1J5RQGdo8E1Q1TIgTJknyENdGthBMt6AtiUG9jjk8d5S92iK0fJIqnPwQSqY01OTnBq7EqQ
wTiACWXxpHlmmNSyv2H8JIMV/VSj8eo1Nq6vcumPR42lwgtCtOhBpU8si8RC5E1gfkKTXqX2Y/H9
POctXWiO28X/Pzmt/uRl4oNx3syAnCMdAAOSS4DDBXrK8MKFKSrg50rjQQWy5DxsnozsYzzI+zXH
RmhSbZJEAL4iFOqEUvSVdOgaps78HFhVDxl7hupL6RoSYse7BSmtxFPFiL/1ZdblQdy/HFcCoO1F
ebpVqtGK1kBculTQhnAnE03fzJ5mBM6yOVHDF+E0QClJcsRri+rJ4pVSeYEJ2ZEoSaFKo9S8bDTQ
8DB3aSKmffajJ4jSDG8cCIZNf1P3cSPmw5A2JHKm4zjPb34jSNHmOv+K8VmnHfRI0Nvx5QF3X96s
gY89KKerLYPBomjPNlJUcwunUbvr0/js2q7Tx6AaAuVwT5C2HxDXaHV7dpSykASteBM7iE7xgJwa
cC/ZY2oJlZ4hV/Vd647yVMSgIXgv2eWsm91gU4+lH52+floW4mQMjhuG9jc+JCcgFm9fqv3/8xpK
xr8vaQ8ZOpTm2/o9S+7uEAFc0yJu4WAxeC5aUYDAqw4TICmkIodeB6/8khkru8vr06cmdShJ1wLO
97OFhwltylu+TuzXZwLsOS6Tj9g/pXEE5FRAU/bOG+Bgq+zIT1AsXXBci58Q2LVPt5obxbiu+bvL
ukrYqXn2dzSdTCSUGnsdmQ28S91IziRTydeJzUJI6oSfc4Z0G8eFFTqbkLgmDlsxYkPvw+g3VIGr
oO/FKqBuxqbu7mnesQ+ZuLH9DH6F812WzPl6wBHayyrJo5/PpSalTHxNKkAqBXlOGX5Kz5Q2pUga
3GWiXUVOX6Rt6cIqXH3bAHTSDzOeBcbI55IHXp6eBSi6RXY7DjH2iOJtbOzd/pUIxI+LdeFWJ2bq
9Vzypg8aTlUt6qjYwDoS3Zu9gfRuNUAxLH4D14nPeLBJ2FWmoLuTCc+cb1SxddNgfTI1jwymblUI
KYLeoZoYz8TLu0X4SjF0YXYKdVdp9vXvw55Uz5iPfPYkHB1EOUxNiZMdnwNw1Anb83nxMWXZRzEa
59tqI2R/QuQHX15Bd2l3/dirBS2Rc5EnwTLJCDmPeY6DpBZrfbx7x0CP2FQMc7OqOcKLyUdUH5Xv
naxSJ5xIGLuhS5JGau3b6xzu1C8DD8oGSYOweIzVFgqyNX7uocbwnCtUubxXgmX4HMdv9LgSruqb
UiJ+YCmyfeEVvce4AlqN6+o5Zs09nuCmFVx10/Pc8sOG3LQ2pkohCjm1YvHkRI+KaTT5S7z/4Glp
jwrsWCx8fp57LxwVwcwqzZNZ79EjK4Tieohz/u+xEAAi4TRgCk8s2Dxsr2U9XLz/Zfpzzw3G9xaj
dbWF5hZWsbyE9Mdg0OeUluFz6BuiyZQPX4cxQhkVWkLI7WK6lDUB4/jiFAgK0gWmalwVNTDRZJVY
XUjTs+S5ZYxOCth+wL3oru0tzd5tZNWDh2bfWo94av5frAMTdiSUe0Hla/ZUshDUL6hNr8Q34QhR
eRKpM2Vz2dl7bKFvOzsrnrQZZMUo1Wo24tU4Sf3zlrXCEtxfbO4FJn54smPyOVEuw6FaeTGIvxf4
zm7wlqKGiAAQASMHr5dHzFZMlPHe2JGU76iC4xLhaa5FDfhk82RqhZVm5VnPwSu4nuxG37vwTPua
e9b9ALPxwzJW0zLsO0FihO/dGKIbQELfiqPlagsiwC9KSqpc/NHHFHq0kGVRLI0ORocEF6sKwpCs
dj/qL/oNorvlL6C/Ga19c+E3vpuGGK9SIiGsZfBivpCqYk0PFlu1ZQncYrjV04VspfC9F79V3kHY
Y/QGaD4qzRQrEMkPdi2cv747RgUqik8gDctn2xWpJVjnfHdQLX3u97wpMv4vdNVdGdhjf48fSXH6
FnD5RnFAt9Qdf+L23KZz0/f++XxW4pv3WocVktUtpWX3DQ/BtSPLtAhj3PdI2ErhA0aD3e8CFr49
gNmxqw53O5wRO3S+a5PUKGwqz1vjq52a3jZyIpDoTKQLdTz0MKObi03EIWF35PeYrLMVjc8FMF8T
0JpJoo1i9LsHU9LzfAGeUh0i3cTmBvIHDbOlcSnvWiMIngbc+/2qbml3hpYIq18wBUD+XsE5Yb3a
LbL0w8u2dsConyRzfg/vHitqEIaJUJnbMsOYIcOvdkAOFxQsHb8/XiDQGPB5IC2Sp0hrwX0qQTfW
ThXwWfBJYbMRJn7LECmRJIzSWuIlO2jaFGiG8h36ZU+YTK5jUGKjObnAn3M0ub0N6hdB+UZR4Trj
S658BNXRHgdD7EV82+W0YzKn7Q0519D2EE9qcDxFUporXAXovXynHe+C3SkvDwUaH7lQfmaf7z4A
zpmQBsw1opuUz07KrKV8PTJqy5jYzgRx13rj0sFHrz1SNlLpmPSHmukFNIuGprwNcEdeS4HmJdBI
L4UqSuuV58I1C/jvAU0OkTj1GtReuoJSyLW4rRof/X+r9e/+20Bqtq8rmzV7ajnMbOz2JnarH6DR
xP0tfJfr3/aVsmIzPZiK6qdc3PEgqY5virbuQ89Xrr04iMYUmMa9EH2nXVu+8cLhJLRQEp487yyc
HyAYy7J+BptZ/r8utgSO8gJvr4TlPYK3f2h2Qri8xU4LgYfNLFpOE77lNVLtZ4L59TUFDalPn7Ga
ubLjZ+BdthTMORT2mVSIl1AKcKpAkQrcQd4Csg8D/KdragyCvQX6FMBTi9d3ucILHwmfbxSYM+Vv
z7IasaqrWKpn++PBmZMUflH7g9xvehem7hyMFVIRLQuBp/WzMGUI0RdT42hTO5Vy/H2anCUB7XnR
IpuQ4KtBajitMzYv82pA8vxLmmgKyvY2IsZ4ZJraIKsgjCmM9xzP02RGIc4I60z7IuK3JPEpfOWo
VOLWo+uxaBtBjhoacgH9KtZtbm7/zRarj2sOO//bfzZZjGCi0ArVHxLFSTaizb0J1RlSSDza2Q3u
hEVhTmE1hmg8xGaqdB9DJDeEhbozTzJo+MnbKQiqF+lClPEW6PpeKZyqjWRWXQwsSflY1eaRwP8z
uIFGkOAd10naD0MEMhmys6dUEuhnN+stTT5B7Z+AwmQ8WxV7JN3z8dixE0pQABzQPm3vjPWaeIA+
qBjaCTk9mTzG2YGpi1baooC7xJXwnMmpXQe70m0zZ/5iHhzwKXlcITkXM6E76KdL3iXM6bU1rTZL
ZKmTYkD1+gHLrbOdXdYbp5cWvnyMPdIJFCff82S4Do9DDdRejO8xURwhO+QASrfV8ahZAuxCVYdh
//SmcCuc0ad3PwsaW+ARrPPcg1w6GJqfMZooBk7V3eVaNA57J7F3hHmf8y3yLE0Z8m1/DyDDP55Z
ESeLnWjdP8Fiv6SCXnTGP7rtCo1sxlgLFdf6wU85bSZnosTp8g3SGnOo3ndF6U1mNI8aZv3QVHeh
It8S1O0A1xe1Hu3Mxw028u5gj/0NPcwOzYLGNHBOqkknWQKlX0yljC3e+wWMhkeIE9mQeFqujT92
JEXSzHwtC5SQ6uvnhE6Ktuunnql/oQS7hjwlKJkKDbitnLtNCIYAJuBA4613KgjYMKWZLegFSt5H
aMrbTdrWNanw8HQjtXASdxP6lE+ynrR+vAke1HfaWhyU2/PlSZHt53jydE9CGy+8ilEAUhajERJP
//83LTYMoQVu2cddYMrCd6Dk+x2LBtfWqV/RqdoLgLY1AVsFaobpPq0FbfMU3lEfurdt5UwDzqSJ
bDmOEs6iSpCBRYxz977hlhvpE1VgAgv4igaf5tdUt9xoqekRVyOsCVN5Mx9LeYOr7wq4K4uPtMm+
N4nR2LXBbL8PN+H9ZQatrytuw4SPwhxuNyrwnSpt/oZe54fHa1iLajAZ/yFgrocuLzzGEC4mgeYx
xT7pUgcJ9aUQXkilFRgug3iAVi3ODx3Ixj54sHi6Iqe059e78UoD1CVfBNbmcxCW6hjKdvcYqqF+
sJR+Ul2EmQwjiQPuvjfQ/bAG+3zES0sutAKwjgnXvFl5X/8lJonvT/ZyKdJ1KlEIcxASDkmHsET6
NAm9jW5k7vPu0adnnKnoZeeJmlt6WyjzQhIBvvhRVl5KgQVjRjcXJhzYQJ4NLgfZgTCCdEBaS5vu
mHWMfRHrZ4hBFPO9Ae33kg5B1O2aQesd3BCcg+ydmnQsE5cok1QS4KnsxDbikCWOLBP0a2HB2F4X
g9DzmWXdooTmBGiN7tSrd1c+xTJelD3MQVlZ4rSnmkIf3XMfJsmEvtfTZychZTtzr6gLz8tnapMt
t3CU43UnRue5RKix8ZHDqZvCTFQ8KkChWRoevN4o+c7w5KLWi0vmI7/RRfAs5KXd2j/mQhv+QViO
49NCwqNkcTPVgFzRKpuKgL50PBCRm0LXIUCqqYoPCJlRrK3YJ4VRGNh0hA1KDHmYKU+Zvmb7qU7N
hZMW4DYJy0Tiz/o9D4hQd+9ao+c0ynfiWZyh9tMJmBFAIoCl5AkxMS7o//b1qTrrKCqEY9f3/B70
pJQxI3r/IxlUU6k4X7UpiafdMYOw76mX+f+2xfvElWBQAeebiI68+KA+8Ob0wabYBB4Uk/M2sa4U
oiVIszYimMtZ9F6n7hHO4RiDre6K0PRNVHLXuI0ZV/bV4cP+UHRh1xWNV7AooNrr0d9B+b6RA+pc
fDLUfISU7E3CUkH0nkwtakJrsoijSoR16RzXYP9gH944NdG01+rL0fSvQvpSQeZvZMYDhSn47jF4
KPOYnmVJBkbxhzUVhuE0cS8F1rVaT9jNdeSQyWyxN8FyjX1a14ZKC7rM5t5OkCYc1PRrkJ/gwYwV
lCrckD3QHL1SOc6jygPTENp59rPCGfDXnrrEqquBO2mA4HVlxThpQp44kRPi8icR/hRdDZ2z3eTq
WfztRY3mGtQUX1KQPb4EZY4Tj3XhP2uTMkYOiPlpokbjamJC4c7kgxbEIsdauPBhMDUq/rutCmVT
D8jLyv3xzWMatWhIwaa9lwYtglatdUdPoLCkxLg1nDMLCkI7YPIxaU2k2yKa+DqvwCbpngCc4iwO
LehVhzwNibA8BwTTgg9kYiSsLTGoGTLw8OQ+p/nV+R5IFdCoVHj50sH3C9SS7uKxtlXD6Vt/IXDx
jCM+Ko4CIi6FhaDB787calfYTbPsLnfje/q1kL9yDoG3s73Nb/A2+LFs1KA8EIjfXt/gb4abyWEb
E9dxJQHlkkddR+422Jn95oU2xO1BnaP8Nvw4yJy781hFFOXnUE7xLilBvRZbEZ2xsCX3j7tR4QOW
Sk/SO7kLHY3P+59sHYt3FV9GENogWqxlN4QhZRQO5bqb36WckWTB4gCHmxK+j7f+uejp5e7fvVMC
Pcjg0ZPN9BibazdOOXLA5MKKe3phjhJ368D/jCVYbZs2+m4mVwYRXKb2OInU7xmIxNgiUr8C9E69
51J2JxMicGfbbc/BjyQ51Bw6AwP2HRx8bnCe6zfcFVBkkztFUEg0C5lwnqbG9BYERqDcO8n21/hg
to3mClHcXoDBapjA0JduyJ7nt0sCQxyc45c8+JqBAkADWesPFH50S0zifUtsh5VD0y/ckOUFWEi5
RmmB6TafwZFnsapRFUN7tq0+rdG4y8JLxin+zMlsj9xvADzCX0OpSGpGnTRwmFKvPDzktJ3MdNy4
StxPYgLleWy0LTXKRgXJMpppGcw/VUuzckDsSrY3ZBd35aGG91fzwh1NQE1SXA87EkN6hhA/N9+S
1hz2Z6SifUxre0qvMPIWatxySV7/zjJRt2S4ozxMbiV71eQ/ZbrvynVnF5x9g8SKLjKcCBSQdcQ0
bGv9UzejSLkOtH+wXAbwzVNVzQHdIuG8FNn5gOmoPPSUpovqG/uPgZ/53pX59ThRtxuvVVjwp8lF
LmNu8K/qJTzdF+q4nhmvdHVu8lz4nanBm/8PsxcapQ9Mt5REZX/QL1nnwsRxxENcURnGMg7vz1E3
BfG0VqVepGAQ4U8KEc55ZfsKCVQ1p5Z6ToiBU8wxm6Beawgw2P8AIVPHpXQ1DlqiAeUpv+WCws4U
gYnQushO8Ta1wi9nvXeSo2MkDlwCt/W5xiW+lR73hMHZX2KedOVQSwlc9CZ5MkTglUWsJFqsFiwk
D8SH220AXIQh+wIYc5lImABn6KsO6E55Bz+bQgIJbrPyjtPpqnnSPQKIXaw8N1uvN0bitCKBtE2Q
ZOCWi3DCTyMhy9M+4roSUF5z4bzyUHUJ0926QRbMdlJrbJylYAxDUpOr9xSVwtxyZgrpkULKDy+o
kP5AKzSZXpziDRxsJUEG5Ts5/oX/um+L+/A+ENi4r6/WBJtnW1VBSGsv2l3QYpV2+H44T+cnFWFa
C8kmqyiz+2tEC+2bJ6GVi3ksxaVPAhtQDt76DA+etM+kG/V3LX9OgpHFdpBzm6ZMvatlCzh2A0ir
QgFBWeBo07TXLkcnthDFNYYRgltvExJZ6JtFkKxOMIcPjs4+C4bGRAyLXFW2vXXNchEMzH3u6HZE
q8pjfqlyn1Ke/8qq8+iqdPORbboLIxRDsuQriiC9zCoC9H7IYuBKjUBO9NV2z0/ECfjA0qNXm2AB
vJV599ECcaoIQtvD9Lb5pRiUMqjdtaqlr0wlnhiXXUIBQF3a3KbrmzmNQQwTgYERxWbqO9DnT8+u
dPp/DAJrIWVLF+AFObe1C51rh7nuc+CdZ4m4+BZ3mlZqZqSlrGDe2vhTMkkxtehpbqGK5z25HIn+
Y2lEiWM+pn+6X1jHr08cqhgObwP/Lv12cA32tgCJiEziRtwt6+LDGKAwiFRwnFC1HrmZwTSRkPy5
MAOVT1DDFfBWQNItCnWEAucGLIjwGJ8EO8wEXu3QY1ow0rnaieGUxRbuOtgwVAlc6PpWXgpwWutt
sLjuQJpKuWWIuCbhy0jScgRXGvtLmMm42X1U0+sBJaLsdE0Gk6BNegpWHZjguELWqTC50mHhm/EQ
CyJNXJcPh1Iwm+qz2LrNIyepJudA4cNGovwo1ZOy8MeV7fZU5yvXl8OkMfoSexbp/xjNvlxRbazy
8dRlVKJ/sGSEpYWoaZ328mfFAMsNcBjGCf5y+8FusURY4DRkAlcZS76cZOkHnOxs+beO0tBlYkRF
RNuDeeDOWEq60AUW7vkLNGKdLNsKiY8DCwR/FrjZn2ra9m6vdcI2IXgc3Mb6UxsTjXtd1QDeLi4G
Y8JmL+cW1HzMktD8giNipapnMAl8f2QWqINL6VHa9Jxcl15bl7kq/Y6zE2iWBWqimbc3jzjmduD9
leVyo7ESHclmyzTRhvOkuoqjgQiVO8pzBm0Hp0+LZvIZLgq2MBfYIYy9m0EgjVSvoKq+7cbMGkSr
P8GzwIwpotwZLG7T1d+XyXxdUqRU1hrs+w6/NqgZK2BIXv24TVu3TNyFEzbZrRIkOXQGZd2/w66u
fLzSgY8L6dOPYsVZJptUSagW+c79VR27zlDDj1fUZmk/RsJ8jj35YvFLXfobq4z9aNbGd7DQ5mCn
526qbU9QCZiahWWPrHOjUsYBOxXkSgiaQuAJqPIFEBgwb+83EFt+3/7jmPXGmd2ZBnL7V9N27m25
ItKNcSzNsKO+8NJKhvWegBPCo+smECI1mjF+SL2JTMfR+AZG7oQhXcxkF0/KcUBd1Vj7HnDywrCA
g6gGh7EiCBau/eXNCNvmcumStb2CFHeMU5wXa6UWyTLgnIazh/SiuPQ20k4RlcMICr7JmVtuZsNG
Vh3A2k0A9VxAq8jOs4bVHCddwnZmRf6n49SSSIAtJm+gn2dkW0gD5pT0p9ajcHSaM3apZBJERaIi
Be6rKALntCUw2JtS62R79h18vwReRQoG9umn4A2TsOrmvVIsGYB61XJDwq5v3a5NzoB5w05sYx0M
pjqkcYTEF93KnhRjzhCn1FIHE7Ol5MqpFnJtcwcs9LFcysMU3Crq9If9SV3ofujCeza3SKiCARFW
2qDbYn5R+x1Q5AuHyYFmqdfnFNf2JmbItc35cJ93ZA/f9sN6HDC5jE2sR2H5tg1PHN8o2YfY6A9f
tHA7oIZnodsdijyAS7XmHTmSXDmM1KwyXZXCU41hS1fj9iwMZf9jmEmiUpy5h9+eQkZe6x6N/0YC
4gZ6ulkT6Lc7A7K0x+EmeWstkMblBReS1NxyHkK009OexPtbl3VXSUo4n3a+8yhCyuDy2UixArI2
ZMxPT9TBz95Hc02+/7SjBaRE5aGi3vGXXNY1jJc243js9YlR9a04uBU6J6XemLiYn5//szau3kp9
xxQ8d0v2+ja6aR5qtvesUtGBYsmpReJUUUR7GdrcmsEyAKQFxWB5gd/ZtkjAAaFl/+2RLakJUukf
6MUt1UlDyNfYi6Xltw4BRA+GOrun99l2WD54/3xNb7syzYF64NAvj+z4K0ceLGvZfJ1KF5IQAyi3
L+HCwShhX1Z6oq/AO0qVI0b6+j9GL5eiYNbM7fKGc9Es8W2oExk5DF97xCdH+mpDZXWWkArBytDO
7qL7AdeR1Z3scTcsy9VXHMXvdrbEXS2wciRwa82ctKdcBckQNRQ3yloVRdXgsvEbMITeUDKkNVoP
VjL92hOsgsVWF0eqKE4oXSLlYyJ/XbXxYPx/qW36cfS0J//lG3FA6mR7vR08df2NZBypx19B47wh
UM0hU+NQBkZSuuF+Xs0ykHd7jYe7Os8+jB2e3WpHntrp376viZ98rAMt5TxyDwoWoKW3/0rOr/Q5
n2EMS4T2qIaEkK9E2lzbPdlHJEUonvSnswi5/2Tmb5+mtHj1qyJHghst/jmp40ORkGK7XgE7GnpH
RxZOx8fOXYa/oFfG0Uxp//OWUnoAhLVUWmXY5wQjM25wvegcrGqQFAfrofjUuLoUsNNPdHPyE3VF
FH1zh+k6j5Q7qEKzvGj3Af9ykFUj3NIBeKPoe6rYVLO9dfSv2mG0OSBwRFlRsXX+VcTDytV8/cOX
iJd6FMPkrt90XU70vMqF67f960iJA1OjywBojjTaUZ1VII0j9qSBq0t9RV00+S4WYGTbEM5NuTTO
1yMGnS8ZEkf+jQZ7/eUUb7IqLFvWQsq5UOzLAlioA5jQBctYlNut7AfXpglQeIf3rX0GQzY4CzBp
qBmb1FWa5gZlWf1XY2lY1l8IA/VSzs8ZuUrB4ZORnbIAAnMooPHrHHBsuNkJ0w/JZhAtgMD2A4Xi
iscNe8hD3lxE8ln1nlPm9chEhC6h1/jCW2jFq+hM1/us5Ek+Au3ZTDm1WF2y5FiRFYycKGK9PmEX
xMVAhVA3HxVIvMs3W/30JtXv6NRMIO1iNnj5x/KLb52gaFSCuYeG9vo7pdZ5y5BkhO5bSgW1rJ2t
7WRRSdCD+LymDH5Yd4zYsAJa4+6AeZEUHH0wddaQfUNfl32XkVkxUYjuhpbYJD+hHBAwNWjbf8QT
pi7nkHcbE0H8hg8xt9lxuETuYuO6DmFjviu6HK4iePC2AMJ0hK/HoQrckmDaKmU5QKNN1TjCPmA4
B/AKAeZyPNhdMsYu3Y6BPPbODCZB3JN3BjdcLHvIzBiMy5Nb1KdJcPusafqwn5mkVi13ARUje1QS
WPMFkbcPAVZ2nW2upfL8AZINQk3leCOkz2fEWbRQturP+94/VLvNW6oUf6BnzCPZcDfJNQTbg09g
DLwlQjSnZ89WEdQTMOZwOLIsQa4c+u1DLIQhzlAnOLT/oZ8sdTEpp7ZnM3x6XTgo1ZrFWl2ddkW8
I9zE01rPs8xRiTUD0VDmxEsm/+OCLknxaAZa70oGFcLzHk8mh7CiFLYOYfCBJPwIpqK+IifeB/T8
BurWY22k6/+pBxl73aydxRKRT7OHT9D9n8JSp0BT4hstlVqbyIqkPfI/KaJbe16EQCMDYcKANM+X
aknJaXLaQJQH4hnAwlsz5/I3d1Ip1QFfL6N74/p/34HqhmXx4i3VsG8Bhd1LkmdHRQqHgnkzMcvt
7nKJcSneJCnT0LWm4gy/kQvAebZl8r+J0m/Zin47UQw0p9voAVeJcMp8FWiCzkWkU3c7Z3A3FPA6
xzzY576KDxlCsmPXtu5bWpmrJGU52SNhy3Wwr2+6UANv7Ge7SlfPkeObixSd7h2UEYd4q4S0dsJi
KI3igPdiju4vanbx8OiMerm9Vclda7OInex7FjBSt++VlDgMN8quNX6JemtmU8qjnWDpxL8kR8HC
rDpKImgD2MZDlgTY4OyFHkVqJcOBEPKNFlqJpVfDMH9Wvx8eOd5UZLFIez5+2mPi/fd1mQYgIzZi
Rl0oP3MjR/rtEo6Kt94ZHXXD1tw8COMiNLMsqP2cegMir0dioR4oHl7TeNfy0fO1q8Rqvvz4SsCV
gRJ0Vyt2OPVMZxrPUF8Zuo4y44SFIuDKQv4XRPzyPzAwxBlzLWyBBV8mO+qQ3hzjfbowOzUYsl5A
Zkwejj1hmmTbCnEAurgr3lhtgA+H66WEF5RR5gKxjdTayO1qJ/OmfrSYHR8PtF9sKDaTvaaUV8jg
tSpff+wOzXQVsxd9vehEBWzxolcadyi0AVMg5y4KRc0sX9lrPQw8Z3ehRefUJ1mC1of2/ofvxbqP
Go30H2LTpTAtr0VYGNfJn3UtyDs1cCKK6x64xkbIDD4Cm7gpAPmxbrIsHgpKhkj8ZaDoCUkdPY48
qnggjki5kfbd3k48qTIOyHVTv77Eaiip/7SxesSTsoRZYbu7FO1rJClFAN+q5U7J+XX4WRxAg0Wv
I0qQkCFwKus78do1zGgWpQPA54kzR8FC5fOYey/Pq2Yp2yjEnirtPlYlSwXn4ixHFHd3aau+aABo
bp6SqJZuXiT3y4VnGRGfEOsssA1vBAljRIOekT7B4chWzTZMMLnGWyCji4DjAwzb/Yc41Ldq2Jmo
nyFW9YRKbvWlTHpH3dXFS4rFOkdY1NdUjIRBQ327/lEr1+8YvNYSiP0s51+q7zU5Nc8pKqHjjvcN
Jwy6KTEcaJzrpgkhTAHFfnUKQG1titohv6dHfJtsTtbKWXb2BDec7uyYZc+v8Y3EeA+vSfHuV6fB
mmfJD/yoky39DhwRbugtj7lMnmALKOfJrBa8Tjl5l2g6cR2Mp9VFCK+YBXQJ5AeLu3suuJ6YdMOR
FOQjTQsP59ZMWD4R0gn/PfZ0Bu5P5+FjfcHRq5Xckb+hKzHp6qd9UYbXmcVB6Xuf81M/GEJp9Up5
Bx3g+e0noScQXImaZAYHhkkLYwdWHLlMKfPrjc10iqTu0rmF1ewrYJEQKAtt+OEgcoqRYb0Yi3z5
tiONgCYYcLV51ThHGQDAqAHfdxPLJbxDO66dZmYFY9FwHgnB8xHVWkYJmTTELmXdW3joWvvuCjtP
Zlz5BGb75YQ4VRUNa2l4CUncJzqivDvOjtqb6nCdLioo7Zp3kXI+7V284shCi8cLpfivXXDmM47h
bbfWMAJrqu4CX2u3YsgIF5EFpSid1D3MhQkR+36WTTI54ofP5S4udZtho87DTZ7PVq2D1O+LHOv2
GfNePW78OVJKAGlvxxEwFHFRQc38xCaoGHZDQGl6H1BCxKrqfGPPgCONi3xGeXya7go2zmJluzRP
I/LUH7LWL4Pyz9Lazwvc9t+uXi70oxUhTUL2fYLKHT4kw7HtGXWm+VKgI5XQ8YZsesFu8BxiB1y4
PXChBUnaXwoBxwpByOWhPcISBkC4AhXUylvb3X+K745xMJzou6I8fh8A/j/39M7nXdjAaPunLxzY
sPPPYkbgTfVnekwW8kp33CLWtflQtBokxYPZUWYM9CexLf/wlrvcnwWEwjQsR6o65ykK10wZelQc
P/XKb9u5FMwMslFGxuVaSLd7Qu0+dliXD2heSHHTRToLjrRrzLGUo+fWZxiIdq4108IQ6iDi1kHh
Gt+yqFtVjtx1fviLcpT2ZM0y7X9K6nHdVIccVhZh2cco9RETHMQtNpLTy1XWmTQJ4Q4krcMwM2nn
yWKEEa2wSpiguY7h8FTGMg6ziTZQOfliEforqeZcQXXEn+V9zRytTfB2SS0nI8FAZwEU0Spkk/qF
YK90SLIbNJAvr5Z8e4hz5cVzqqvt8Cen2/BKSg1NVNwr25Jg10QVsEkrB6lCmuicTCjuFWiQBEXv
sFQopW6bpyf0KB1Yi9lL3zrBWg099iofbzFCKzD/qcA4PFtFFZQcmNZdT2KXqWD50PW0fZaMUwFk
pGqDcaol1NxJa05dUNrhEfYQ0QKdLk350EBrIEis6ytf21Zn/nhGYSySd23Lqd8ychU6amRmNzNv
aefvuWTRZyl4IgnOiDi+2oCIKRW+MPwzVhWPDMTrzkuQ3vEHNEn1LTEOfRmosWcb/QmLMp8Lpvzp
AOquf3+ikxxKsI/7gfeUUZnAkZklZ9v762lOA+BHHxgvgSG5vBzqgh0s0iwJMIydipQ5yhSPvFBj
mXZ42CFRTxYs78WkcwaZgJLZW8LcszpGkULtX4Ls/5U8+H/zx0hj/q60qeQJR6NHA1dmVBlsm+C0
qn5W66gfReRAu9DKzG1RWACYpEoMkYqV8CnSru+87Z2i4Iqlzfcy17HFgkC2FqX02aVC67sF99Ef
hFVgKs3ghA5hmDik8ciK/EZHypzg/PmWWs0XqvsXD+l7lh1znYFpU7HgK0gqPIvU+mJPBqoUdu3u
JWWrv8AnGUS015+5Ykza6QMGo6RQ30zWu4yuE0iHFO5HYiof5dprU8CV3vdSqauqe3f+YFT0USw/
727n7CKJUNTsWYYuoEndcdeLicyrgVSO5/i3zIHaE0GHOCj+WhJYLBGsNQZe5WTOVGudLjroHIgm
mkxrUHU5k7soROlhI0CRwihNz1eknhAFgopp5Dc0qkEt+4/XQpQqyPhlnq+Rw81lXR6y2nlyLJew
ea8dYPPP1xagsklbgVOCBNNCTOcM46C0KgJ6JltDnNfDQOIoevh5vXhlFHd7JyyJPuzCesxxxIBY
gKXSm9tigsqfq0Cl8R4LplTKexSqWbAhm7PIz7DpIoxlF3LbYK5W07OTCj5xKIGOLNQwH+12JRXl
cBl/TsgknuTyonjE1xgBPi1JlTmR1ZdjBPh7vmhbIp5P2Ian4adSEZo1bSvVckZkQ+RVvoJsNysL
SdA6yyiLW7F38mb/G9usq4hfJwKAvr6x7r3ejSmF3vCynJRFodh9QD6VIBP///9w3HwNdh3rthtQ
ahBSRvfCsJAkUsIi3QRv9H2Ri3ygMiD1HDWbcqPdS8L2OCwhlk4kepo0IJ0l7TRVKbiQRy22GW7I
2fEEuiTpBdSNZA5OiQ+p42mVJDqnPN/DNKDVE7HM6Xb3VAj+fNQDmk56E+VPVApdkHWRBHqBIiTF
4Et7+X5rHh9VtQ+qNykbXV2Xbm8cR1w5Oscn1XnmN81SLP6cNfUr6LCluBi9b3dusFEYbTsovYKh
D896J6A+Z3i+0EA6+hu1TBF+1cgC8RNN1Auw/5aCEC6nQJEvkg1wn9Bnasnf/CtTfp0o55g79rcW
zqcUvjzipxweUdZAmvBWlg/7JXk0eQJ7QdfcFQnyevPxjzQgDY0Q0YHVbI0aioRD+3LyjztVdxOl
Ty3BKPCiOdjk6+rrLFWcDThc4Y9GuBDynS3pU0JNJFregbJKKshHnhD8ssyKjk9ziv1bIfIVAygF
uBLgLlA2niws9fmkrmoUVNzM7sQt2CnkD5y4LPP9Y6lqxXCqJ10e9by91Ubzoz3zW6MWTJMGZ3Ls
8k4KTNiritxSVgSTj1e5B/HFQGb6iPBdFbh7cQKlCYLIuEn8ZQ+f+K/hwwb5FG/LiuqUT3l8jYpt
Gliy5FLRsvnTomVsiGugClAaUQEsHcg5DSd7S8jBBH+rQ3VKrtP9P7WzsTQNbBnNAUdp90Qxt4UX
lGJZ+T2ngzYk2TBY8sXkAeU3g1FcanQjSJ13Xz42ranJVovSYws6Jgu2Dmfmnpq55N3NkhmAob+x
QBVCRXG4h0usln7JgE9FeqEeleJCjZRpcIfK4jHsLZ9KGuGcA6wUAa1J9LWcjQbiU7f8jl2wPJyF
xAehU1mcPxN3p1PJ4Xp6TZhe7BB9cO0fREa+Ki260bKIFAxAZjPEExjGJkaGMBVCrS5s3yuejD3M
EiCS5O+g7f51CJYst8qfabFIOtwIkaGMkFpwnpdZdH/E3vienyx4kwHJeNpreJUZv7NwJ8vTwP5w
va+X5iKUtSoQTPXZeLyGH+IaCUXEnJuPyCVoa1AUYIkFzQFd8MiXWZGWjyKFYfH29qHNgN8M30SB
BTU/QQ/Fn5Mc8i0kOVH9pMznzPzSIB7HSnSMTou4r8uNYHxUfYhPlhHkJOBnRPhxZl8BJQrj+Z1T
75qQG9s23heF50x5DdJth1KVJWJ5eS89CxhssEFzSfnAsJ9KzLYNDWz8evaSKEFRFWPpuMRo7zy1
lL5nWvAkrW/YXqhPBnShe9bgKRR/5Y0lnYzt9Jksjc1wo/lOiAB60pBxRNFBgCRvQBdB8/WamZ77
l0lZx/77chn9wVrAhb8xEc8NwzSTtN6YcBEd1Mx2TIAqPfFJNxamcrUlWCN5WI13E7S9WOtBPlFb
gERMQ+/heD4q7dek6oKjeYBjoR+iEDEZQTNA/p1458o/LFCBfCVkdv0wKRnVsk8S91eMEAIfEXlD
J9sIoFXsEYifOOl7oTpSEbH/P/SfTpSgu84uk7fMsp5wZtw9MLOxkoKBaPXeNiAH45qSYrx3IcpE
1XdzTSFqzjtJqROHMJFkzVWy8/OaZDfusWaivWxHtsHXodppqEU8UMwOGPit70BTQXxq3JDWf5+b
cxC6TkZPaTFiLeNh1FU2elnANGS9ugU9sbOyTtOktGd5+mYnDd3XnfAecLzCEg+RpJBAsFun/JvD
Lw3Amotp/0pLdlEqO/niYokaWQEiy4amZwWBWeSRMdVMwcgjuUnikoO5BbNPEUQxwuqbpLj63jhj
LXLRHbx1LbHvbEBH9Cxg7nrVd4SAwsun8k7oFVD4u5IUtSdS+2r5kM2PCu3qOW2grRdvFLMDX4Xo
7SdMxgjcsrZQhyxIzmuSoqH6C5c2YbBIVVmhfjoIHoPWa8I9yeWPBrlE2+hwszS2RHP8ywptpHBQ
pATbNeBKvj04W7b44wVNjTNg8PKBrShPnHYmMKu5j4xBAMDbiSL3SzMw9p/XjTNnJZZSo3Y9bF06
Vde9CdDhfyr95C1H9mLVBsZtepwmol3uAXcyQRS/uRKxN17eF/yW6/GRq3tSLu6YQUQLvkmgf3Gs
+L/2dOghgYyFHCbR0ztGqf/AYQYAsFmY0ZuGhNs0GDAmg36CKOeM6uwdcfVe2kwbxslFK8geTVGS
P/t89rJlFyzmrXoC+5M6YTOxgDGxm6Wvry2allr47EkBXxUvAlZvFrlj375XOu6a9ijuVti5Nk+C
UsvyjmQxBQoXIKx6rZz1QPBJTva+RJR4jUuX6UvfX7E+AAWUu+GYRdXdZPQtaBfNJ4S1wtD9r2Sz
UU7R4ZtbV2ncjyr7kO5VPzgL4gu+HrVvtluvhGRMQ9AQKNPuUj4zVlf4SJtYVZqrPpqv086hVEAx
ILSJoM93GloKNDqzWrIYlJ8zaeMNVTg8dI85LEv3T0IMocgHYnl9xioHTWIZMiiF0OFdorDX/E1S
e0N8piEloaRacqEF/glM4+20z0MEkr2WQMlFBdJcVGcRXJP6kYFAlnaVe+zTQ/tUtSzvpp5/QGEA
3hH7eB9fNrCvTvTFHRNhvyGoDO56fmGnRPwJNb+9p+MN2fqLq2t+rWyXJKIu1BPCT818rmsw2iKd
coYy1rV+F2+UDQf/Ci9smrj64pb4rmMiQNeiwI3koLks37A90qRJnhclkHF9S9sxqgX823m6veYx
n1cPib8XjiX7UGUB1F/ndcgZ4IMzHcMyLUEWuVBXrS/c3l99m07yVzLl6ejGZvsKW9yvZbU+rNa+
ebsll5oZDju1UOsBUFKH/3nOGR0PA5hRLSLmo+a6YQMIRAm3VpCSJjB8lUMjKU9bFeUTbLm2svXc
duL8PYF/CosHXeE0eI33cTDZRFhP5Ny+eZ+IIfxJ/csL1SMawd1TfPYDwnsYE0Zc1fzgFba4WkAY
K0bF0olBzaPZaGQE9PzLrV+h3mfI+yWyo7HeGNeH/vMsl1EMv8NRjeQ2pY1rtaAzLHNiznj0vNoC
smmRdP65EwtMZDwm9JmaYuoIXLwXidijE+R9av8Zvt27abjq4UNWuYqhanYQKk8h7NPTzWzVJ7eY
I3uOD2JlB8QIWuYJv3v2HNs4KBrgtZ4EgsJOi1ygAZZZN9hJ1+qOPYMROzh5Wb582I6tDY8BqwdV
0sgiHsxulKEgQlOZRH0ipqdLHKf7GxF6ND9NQi7G/K6d1/WXwuwpYKYrzEBoi6BCVtpA11Bl85b4
FdfsCPrsJoQYsh+VleSysM4ppnPotvTGZJb5ZHIgG77oeKkzLK5v0BX7N65BOdd4QDQM22VLYx0l
6cGs6ikQ42wgY+UDRnxrzXlarAWXsPpKP9At9w6UUGCDtaLLNAiuoRuqzkV5L2O3X3oXH4TpM8v7
kjmx7PbVuRCrtu9BDhqaJp+1wXfyWsL6CTH2EP4HIuzncSkOYH34ucdciyJLuB2Bu2hJanPyqNa5
KAmG4wkl1QJSr9sC8KrU1EALVRWqXJm0V2YPi8xgkE4g0YCCACdEbMSe6NDY1Pbu6prC4JxOfW7J
Po5a0wszhqtLkviIfId43MY6XPR4pGGU+m8voiWG6T3kYUuIjP7u7JTWKdcyep0yF1FCCobWY6zu
5nCAOqBRJpfQdbamCK2DzTFKdF0/ta8FwgmLplcytEW4VA2WEelOdlYS9NkyPR9ZAN8h7npghKqO
wDkJnHr53ynhvc403Dbz7tJ78mT0bwXZtXdPxASEeRKAWSzkYA/7QpXxQnY9CY0yAa/KDYU4awmQ
FqiiuK0hzf4WUFY/FOcCuDRYjAv706YtMYVXVisn0FGUS950buh8Cyc3HyhS5GsXOgTBSiITq6Sg
cuvt6nj9OfeGQrfCp9cuSfFFQ35poaVZJLXaNyckcd5BWLGZh6HThn/0USMFyNbrIjOlfw1bZ8Z2
CPoPYYLfjbYXOKldp5E1Hdh3L80C9KCnAbyeOsCkCXGOeioWrQo1C+0fdDIic8bsOqH3spGuFB1V
XPDVIdUFK+Tual6shmgY4na3UCfybcIvYRfbu/VPJ3bucQopyeczzStXRUuNS77AGzAjpZ+D4YYI
yLaRHlWk6htH3rJC/imit2aBtm44Y3l6yZc6e65yEjkLZrf87CI3SsxdeISecK/u5Fid4X+gNdau
mfwIuAoB6tlq177BZbLSBOtXcoFTfdwR2h/KH3dekZKe6SQXxngumglpeN88sPj5FLCQVdNBLA2j
YS+8AMn4r1REfFwdO/JAVfvhOXrNwByoTM320yatl7bFZHTvlC97ASfUvtjjyNBs4K17mfWKYm+l
iv0OxtRKZl604wRVH+lXv0vXeCfKcFDkbccmEdVSgHBtZaDKKeDozaKpthBQsTxsjEMxnRf0qkUh
IAhrYv+NFwVFnS7qo5w4jEzUKukIH/Kn7JWeuGkQ2M/LgqWScD9MFIwfKZR1NuQCdRKElnxulT3r
QVU5h+L6xpypWpno2IVeFqkiMSXUWwLPhzxhxEZB23Cp/A9sOXsE36yz/ufKy8TXc4sHgialUOOI
aSaUvYBcHN+5TA1zKi7FkKhADt9sgBpjD8YSBN9G2uDLRM9r03A7RfewwMdgsDY5VrHD6s84iyps
bVu2hTL8JnCnJP/wgcoq2/sjAFZZh9jX9/lVOFq74O50w1MUITdUBddxpR3bf/TgiA/xTkCRYVir
BXSZ7ZIuAHiNJFpdWSCoSFBiPN5vGG6ElkBEm7E+vm1MriWXeyu+Sex1JrWKckKwCmT/BAL1MifF
OloqRjyIFnONXwyrGC7/fci4W8VNL24A2A40g0EZ25+PxE12xv8pHVZ93CR4to5XleWeXy638wMW
VycJNqw8GYQOljOD1KMGCil6lcIzruPt+3Ze7lePN2O2DJOammf3rA1+4INg7POEQYsYZ6ciVwv0
AUFZuqJ61sY5AKHSweILIU8tN1mcER55adCT05+EZ5fzeuTcOXKuyjGc6aPE5SSLH9adiEMS5XPk
jya6ZhTV/BK66XeYXOZOzgzX4ot7CAnTar0gZAvF5hh8YW+8YeUqhix2DRzR9izjbV1LJRgnhct3
lS8KvVt4Kg7LMJvXMn42+05klvyaPAWrQYTrz9gBiXs8sTYNCxinkM9ktCyYHu2skqV9lmUif6WZ
eZe7Io34aHOMfkOGX93elrmJVhN5vmx3f1qbyDQLNp0kxwK/ktHADY/7Jfc+xhyATwj/cH3CgqWq
u7Wh7YgbnvH0Tujb07vlgJVTuf+7PMEnpbbWeBDVWgIg/wDnNLe61Fq2Ru47tvKLZJOWMySFJOGH
eC+illbm5GBh4Li6Gs9bOS+TLpD+ITaZvWsu81n0gMJ0rS+kNBz6qzNSAiYSGJgmFC6NZ6d0iXhd
vNB5offoF5ghNB5tCXli578fpXKW5aPnLUuTImDh0Ga2DsvZ7cp0Y5vZOj+lOW8BPfoCDrxHNpTM
V8BXVymPP5cD9fFFGqyGvbaLmevVp66Pd9h0tTkXmGCRu4rZwcQ1yhFxtTQYFz5ZBkizMAovkqux
mwype0v1086LkaRdF8VVCKgKtvBJUVpAO34EIO/A0fMvn1q0xZ6uYVNGP6uLALDPfGDsTnDGEBcq
GI2FPSYn4Na1rZdcvqtydT3N5aWfVKUOO8y4QQOnts/aOC+QpCDjoK98HlHhyrUWfYf6RVj3iUPT
XJJJKhSPEDjxHnMO2m9Az1NSjal9eYIwTNCSU7j3Gy2OVwP7p+RVbbf47CBErKJRr6UXX0I//3GT
+NZ0lZbHt3Rtic2dkdCukSwP2rqeovjH9FWd+1AQ8GmM0xlBfdDV5JX1DvbgR/LT4MMJwByskrVe
hILNPIiwrtf4OIZicyMgP34gRfSKYFacKrfsflxrMdSTVx9KiOZ1Q7j41g3lrxenQ02lK91qgM+d
uN5vQnkkxjp3fqwMiQ8L0cOvYTthVI2FoL3DqWzh/qxEka2sculRvrIpOMtPw6L4r6u9dsikzVpp
ykehegudxfmGl+Tk1KD8SBk6vsFCtkQZWTiMDVQ0sP8KRtKsPMaF1oict0JAOtsUtjVyiniafDNX
FOZ+qPxPOTEHtJGxnLDiIE7iXJUbsaVKVSpu3KtIo207g/qV2hbh2oCmtiBbGUNNrEsxytcZafO/
rdlqEefU/Mc5tBW5jIaD8zS9xePzsaNRGTjSvrRqp1BIODRI12mGU07KZiinkxn+dGRle/VDxnpz
3mhgLLolsi4izfieKu5J4ZR+OcbExCzGqg97OCVjrIQGd0rc9BkRoaBoEmRih28K3m5fT8yV7523
MGDTziheLNxckB8xZRaRzC+hSz+KwAKxhYwh+5/XFsnAsjW7hXV0hOTV8fhENuZkayIB2/nreJCa
4Jy06GQ4e6UVwvIz0FkfLa4yPLKi1JjzhbgWiHUUlKKFu/Hr+5Vg0pPJ3dsmt45jA6Q1FDiOf+tY
Zank0axpZR+FSKYsknNbtXLtmQnD+DjCdIrBUPFzVHZlV0m/ZSVNDYwEwwlBYh/5pY/XNSiiMImC
LTEPznzZRkrjUbnmXOlFrr7FaqXr1kIv7MXzHfURN2coaeM0g3boK/jJEKn1HqW7Nil7037kuhlP
k3L+dCOMVW1W0Xs+6zvYfIpBULTcvoiYoFi79OPcGKHByRriX5uSxdSMxAip8HQX/Z8rDD2Y+p5W
rGeoSuQzAmqQMdN52s4vVDGxGKqWLxIVrB7TXRCzpA12WPWap17+RzLx4AgYlESjdxKcRVlEZXmS
7KeV4jvgB9TH7Hjmwqv6BYlMBWQk080O36Fm3BuR/shZ+wzAX4n0rj63ktXyhzKKIsa8GsPEGBvw
Nk/e+gORqBnMTLkTCcqxYHZ6zIWZ4Uzkv6FsnVYwMI/rV19IMX3Qnzn82eBNOehDDXx0maZIU7jX
L0t7ILG31k5OFptkeKas+xcCFLH2D03fHrOpXIfEOuNfPwklx+RDsaImRlbNkSX6zA02cmgAy055
PGUSIkP//4GqtS3gPUP5KY3kke/uuc8iGZYCQpfwitq01nnbY7lTtkSdxvkwmu3goQxV9KPPATHP
ObwWfP3qXVd06yZ5QqC9MSJc4Zelep8npiV4vw6vdcDMozs1Pzs6qGAhEvVFI+a1tPLJiZSaEMbq
2AfP+MOxGmCwEtfFYgwg3/Hy39d5e/BAqXwp7hSCItInyTPWbBlM0AQOROpbhKjiaMvLveuj/2Fz
A/VE3CFsQtuyC/GIzkYtgG3ghudeJA79Ty1pDQqUFCGoXCK72v+7kFjmUq3Lw4tFeJOb1iQSmcPK
9E5UPC3bIfOVeVFbOezqZ6QDJ6DfRV1oRKmPNuePu6Kxi9/IN3n/bRLSw8sMqQuTjtJ+SkJHQwKM
RL9mIsy0F2yhGjWZJ6h5IrtnWlBI0kZONcQMlOiG7Vlv9IucgoUeIcjkCQgXXFpagCojhjSNtvBa
bOGbkzwNf6qI7h0vLzav72ldMrUtH3J7/VaHz+/Kc18ZSsk5YhlN6ecFRQ6Aq9i2eM6LtPZsegcP
B9tjTc4L4V9Dy3DQLeDprwI5xXPv6ICuKIk24C72HjfCmBeUXSgGspysi1c9aLqs/rL8F3V7JNNS
tzZznI3DxcUjwOkFpgHvBLV2itWOFP7aJ3JNUySSys6TwQD8TP0DO4VsQxgozcZhvFu0ObavUSn3
Sviy8bPZ4/2VqhpuvpoqiluCbSgSBEkSVhKtGugYhfh1rtPPi2bNVBM9k8t4mm/0/5pgG9+0WBqa
dwvGkR9ch0dYaaREQmZC12LV4e1kWe4Np2mBNvE7o0lVCnyasQmAfnsLE51J9Wh8vNZjCOK+HRrb
3mYUw/YuWHpoyN4q3ALoiF7qFV9aLF3d6uZpJVRNX31hzvkZ1HOkc+9owrjSEcnnAI6wgWVhc35G
fHhya2Z0wcSbV6zBqsgnZVlCN9xO2dcQ72UxlGS6ZxQhQsXchpPi0yNNT7Tid6Mj0RfJCbucyf5g
4ixS5v1HR7NgaNpFHIxy9M10ee0rVX1Xz1mPR8zqCBRd1NKxpxNseiUq61w50cgbubQVJxa7nnQr
W8M4H2Mzxdi4BvyqQcpTmhXbUbWHK1Bdm6z11R48eETDwvaF9vpykXd8+Z+MS0B2UFURVhnIQLRJ
B+SYAD7tq7PBGW85qsRpnWhWitS1bcnqFRojjxn4xWl8TSqUpYuWuowGg0bTwqS9JPDwBH7Vs2OP
hlDdlRLgca4s1Lpd6ERzeh34vbzuS/njP/31kF2Y6HavTx2GS7KCScTRD4JC9u9aOt+jWVEyVm19
yKEv55+52Kv+hW2Etgx1Nyo5AcKULex16uTSsG75zWcQBCkdHbNq/7Rc5Gol3iMafafuITFflkky
1l7NTPlvhmmyH72JA6XsbhQK3EVm97i9RVPrn5wR4JHMSpI985bKPlZJFdtn7w3dUjiAvZkhqE+B
/5HAO+KtMBhr47dl0n7Y3cX92ucO4sQgHhFSfnt5wQ25n6nz3ul8aKEp9csg7Bc5p2FK5VIKDhfs
BlYNFqCQ0oS3uqTpNhozb+Ea5eCRsbqoPUKsduLFFmT/hL8XXkpQ+BwyE+wmSEUqQktW/UB6kNt8
oLBr9e/w9XqckuISW98QmPanJY/4HQlH4pVACteYNpKW1cyH/OtjPThxX0rSQq15BoaOmFE9BhmG
yYAcapunhbUQ17t53wYCMeWp2ahHNvkwLBYCUDUKq5BePi1QpdJ7uKa3mfCpLEuPdpB/wgCD8OVM
MS9mJiAwEcfgDMy/OpU0E6FfL21b5a6n+3ECasnWYNbS0UiHf4rQshAKzK23tI5tLwkkCnBLjYp1
NsYZlXoC3fGJd98KkuaL8Aee/Y9oETjrTPvduATV3J6xx/LY+m2Mmp9sNbvJDKrazVYGfMZWAsK3
pnlZOoerlBVvI5OsVP9drWl4S73hWKDlLiEfF9v01Njq1sfI7Fk1w5CTbj3s2l9jK8gESlYNmu60
YC+oa3969ZBv1GDdfBK94MOYVs/orY/hJgzBSDWoZWbL4/3K993+W4pZVa15/X+f2dHV4yKzY5UC
KlP9ej0qd2Py3oj/N1QIv5QAoRMQU7ftZg6uPQMtyFm6y61Jku7tkvxckE53PSDysZnjwWtG1EjT
C/7WyVYHcNUjynOkRBx5lTtQi1THLljfSB6m2DqlN1IOMY2QS4Xby8Ro5tr24C4+bQ0Zs0tXdZnY
kGdWPxvOMGX6HkadnPd6AD3FwyhmybSJz/NugwTMOpNcsYk4xxVMol3CvkH/MyJlkOeDRuxpmKU4
WB7i/1GFa8uHMPJcCCMfd/z/+K0sfW1nl8MX0sGg06WWD5I9VkdkVfBpjjTG5JWFktbl+O97KHFC
EJ8WrNr+bytqpUaDOaQFIfFV8aX5k0v7fC/DHdvFGVPeJQdxFC57Enz/lJ7jeLvqDTrJQAr0i7jP
tSA/neJ72g/H10KMVNg5rKKbyuWnxRm6vzVRzI3ENRY5KriYabnKgkmVYipfNoeT6MCJz2DQ4hpl
XIg4y0bMlqY9BnHczZ4GfClB3OXH3fZyC722Kt9Qn2C9+cLbadkp/ZUwC4FSaDQBWiGg1xPpkVMH
O1vxLKTmuW28/vuaThBbb3mPSnVtF/uMKb3bG8lM+iby38Miy3d5GFbDy6A4w2E5UsJI5lailVCz
9lQLZA9hSxGxOU/8Bt17NLt7JqnIjGjUu7qloPd8nU1KrPEX34opR4Z6Yk0XwfbjIvLu27x16msW
ylXsHJmWHCNZ77X4xyCpxVxhdDK9lIfcznY/aE64DSQXTy24Avzlpcd1RNROgz8qoPQqwZb6f5tn
GNi6j8UAcZkCybOMaER+W5CJ6rncbZ64zQOl99cA1xHN1y0K5l/DW4u0i87euRfooqUOz0hVmfED
HL5uNuySkqReAxyOA+wNZSuy235wnI/4lhLXr9isnEOD8BpBv9ReWpJbU1IsV+88ArMvuPdVJj8K
e6vLynMQtv69wMNxv1kxvYbjI7+fMOfSEEfH7afTekHpV9l/9GXAtZkpH1WhKRfh+1RmNLxjBfkL
0ShYJTn021hL1AGIBbxWBnFPnTzs6DCSZ35oFjUVfhB37nx3VZF6JdwvjvNsEQXSyylxrl/VWNJj
GgbRkMbcyTgMeWFV5usQ+J140m8QQHpwQWIazc8hr8qSkTGbIuh7WGWwJ/rABJ5rACdV6JLDeLOJ
SZS1uSqxwS8wIMys1fTq5ugXZhQ6MJEnUkYSYWar7PPVEOQV0InvTssPuV5qfH3hkzKdWczmBf/L
d7jWm9fcPUyznr4LIWaGF8ptj/kocg1skBCPMp3oL0UjXQkQc6lMedxGDqCRXr/fOrG53hhzwqxY
dGIwNjXo0usOfc/7PTT1P6W/dlJW/TZ7otMvkp4CHLsg0vZ7q1kKkMAYRrWwmPHAoc98btQf2q6+
85Az3731HKaAXEwKcejQvgqvqs8x8Swwh82ViTANYIryCrmYNKgU4ekH7eVJ1mwuI4+dcmpqAMaK
DVyxw2K6RYpetASZwBCZZrSUZ+TnhoyL1Z5hRzEtoiQFXWMS9AaC+AVZqawggjq6w0A44qe4xJka
bzvDSfXAZG5OCABCjfsbAKqQzqWZ5a/R3H93mrT4fBQ/2Fhvbfpj/EXHNwoOP7sxLtA7OWcS/CYw
LekX5XLXopVWhKMYmmkIF+T7vMjrUIZxcJWGaUcXTvN3RGevzelBgxLc5LwfYReaQsDn8zI3Tvlx
TT0FiufRA8r0ySF/WgQEtASyk5LdcO3acAnAhu8D+/mNPVdQOhGJitH3qdxjx4zqKIUBkR5uA3y4
8iF817pWGotIKfO7jXlFUTEkThIU9eCE9mAcws2sjDtPH/gF++NbgHtCLbvbLmGSbNSX4SDSlwQQ
8SR8Wn+TYPjLPlaWuYTSxV4u2qpDvTFKDtL6LI6qeKF5FD4CYXnbBn+TG9sdeHZ8bfk24kGHDMk+
BZVWe1yYQngkbWXmYjlP5ZhfbPd0SH34whjvazp1lQ30vKy7rIBicJTEJPppYmawcj/aPZUbLbkO
FRT8R66IekjUzj30gWCa6+LJ/Cm0Zh87tiwlI1C0AE86UntPBhCGY29jhCGBQ6BVh7pksqDIKASH
75aHACpEPXCPf7Hd8K98ksrigE5nVQKBx9fySUZEgyi/ZURAlPlAcBdyoG2bYUT6MPZaWtrlEIaO
DYk1XFZ8ci8N9cZSqahJHIG1iuJYKwVIkvAzTXepmh/A4F0104wVV/JswfX+Po1/Tvjze1zQ/RIt
GLqaVZMcKFqg18rze1BmPYFHmA1MFVq3eEWX2AEOJMcea4h9zIlmapIMCM7qDhqzmJQPf+ouEafe
nBXqMZ7H5kRYMuYUhNIjDZe2YMtl/BU2sUosYR9vHfqWfXqmV3A6/RbZgLB1ole+F7bdnDejYd+7
5QVtYi8g69S6rbW7XgeDm13o6pDlDtPfytBDWzr0q038O4MuwOWGv8TjP9KIrhsPXbfiHsGS2Rot
68nuFCMjRt0BHsqSQIMq7l7RWWjPXoIqz2a4xW8/mbBPj2rhrST4p+w3E0yn6i0ylKcYBsXECg8G
CZJE9QWsqe+b5xplEcr3Gye+qhzZgDi7sNBL//vGcKngFGyPhJxjOC2ixMeOHvwfyeqIByuNgbrM
F9jhJafhZGw5oEP+5L+6f6tNrzSkttwrhT4306I3yzZAOGN4XPQPtpVMzpvGTSCnYe4vuhSjHuOi
bjHFxs+/6w7n/49pWD2pEqyvJsIwLfV5CQS313DQJV9OnNHP2bqDd5/6dn8Aqf9O8IVv5I2vz6Vm
1940SdYvAS2fuhFygDC6MlZHW+gzf4GWO8g3vLfbRebZ3xXKAV+5+dNhDG/xLNF616RZ3lH8PY9o
2PygqNJ4xH8VbTAii1bMWgs7cJRi96E2GtxPU/OwmqniuQhAGQcUy42mhxJs4v3hVe+TGNmNvfc2
PDutIDlmHzD4yJEzJVYa3racoGB1UJQyK1i7Zeepahi/njJp0GZl2VoeP09mAVv5Ks3NYbZGtet4
K4/B3OCT7gDoP8xyDQcpQ0JFazxqdBl87+PtgEvpq9yYhDcKAmHquvveEcEn03AIqmvg78W0rRzl
a/gVJKTBOHAtk0a4dHaS0QLrR93s7gPYSszXCR/WHoRynLG7hhgIMAhKhZoQhEM2yAFgwlbHKMOX
u2PiRFnQaRHnofnoOB6nFjcKH8R1wgmoGiA3E7BTH1OQbcXJ2Onzb0smV7sQNo26a9EaVebu7/g/
vTYEboEWU3CU8EKk0JueFhiUHNkxkAoPjTzZct8vnk5KKR7ceaGehfbtWQOxcambefhF95z7KHBs
FhIWvOVYiCc0FnJtC2JRy240CG3Q8liCB334rZBvLDMmlABsHf2rrtI+JNELcMI7fCq9j6r3i2NI
gYd82JSYyqzksuILZDEse+x1SCFHIRsOc1GSKg0MPkebSpqahDXKTt+g5GusRtxADvXgMTSNs2b3
SnnTIMShZmWf17NG9iUBFZsHKK3T7ACq62PIbBu6ReRSekBab3kgU70w6ZleeMpQbrW/GV3b5Iel
oY8Awfu9CTvlDl06nqVlvlFGD7LOWp337WwjoZhBQ6y3p9TenjGs8ZoYIQJkWwq373ggu0ca2vZI
gSZI1uWy9iYhDTIy/zo79IObx45vGzJAlYvcVYs9IdcIMt9ftcRVfGgVVmO897rjUmDp7ayQUNk3
aHD6KB1TIdcp3wVEnXlz6PY3kHntjWGTXfu/7NPDcqGlbbUY7UVak4HOar00lTiXONVmkDOD5g1+
Lya/r9RzUWlZ8RBljEPVROu8faSfyKMU5Q9ecNyDcAYC48S950TbyLVSwr1+fvQFoiseGxEBF5kv
ReXeCsaGtUA8djv43dDJi42F1BgzAop4PF3vplRdXiyRRKWVvn6I+U86w16+jAz4+bs59uQk+TbH
UOYiwtbYcz17E76ZaRzPOVOpnYDhDO5d6JT8UNYmB1lTf0gmYy9wsnWhLQvlmtMMYfvjsHHympIh
LegIm+MN99eAvaSGzUxpl09Vl1fa4qXivHnwpN0Ij0mXWO8yknvSxazzMDJRiPxblY7lbw8OTQ2j
j1whwKUl9FPH0a8XAaHDYhvEitWA6Y//aM8QWWI/++Xpwc9af62cqa25vkR2lCeHE/XkcfAqJCM9
PjvD4aMk/vdF1wfp1ZhNqp2JirysxzeLU1xK23Wl+gnJK6jxERSYzkxXBHIat7XSYiSTJVzIl2dR
dJYrN4bQZUZtfIaYSXjOLPSz2cInZbsQ18S2mAQddnZJGUcDpkBlPyEPmy3jKd7F0lGsViFgMX/o
mHtdeu5hNAgj8w7QYviXnnmBP+EHNsGRVvl7KBfZHGLqsuwrjNb3FONxb0IeHdoqS17tLdEVMZCI
t4cXP80QBmf90qxXLUFprSdIqDMveLnGfmTFQQOehqWWKwVx7L4ud/EtjxHP0IHFHVb/qvAMq7D3
gHKGkeMzMCemirWpbg5K9LNDqPhYQsc0IPvoRvog/HrdDdicqrLtmNWvSh36XuVPLsN/qMdr+QlI
ERoEBRG5jVe4Ii4y6Nm0RfiFvldRTvstVPUKHh1zFZCk23U8WIGl2Jo92rdtc92gPKZT39W1iaQh
kWJaTw+ZUqnjTeuEu1UMTHdZgJGjUEKoOZ6QGsLCZtxNExNV6aPtwI6MitE8Ts7mJDY90EwdIeQY
mW2Sj1vITscCjBz3astslfx3z5zF/nx/euHqnPl0xBl6XuBwNcK5jiacRwghGap14Nm4ceclf1f/
eM1fPNTZd05GGa//MTeX5v0iTDoUbUgwYKwSp9E2aHhDtCj2gA1bMggRVTG9Uf50otQtq6BItmiR
PFiWKsF7313xYgGpbk2Yqrv9r0f3vS9PDfJRfoIOptiP6EGICT7znyeW/T1Pgz1sdGGOMcKW/Rsd
VackM9s5uGW+7JxzYDaKWm8rCoAC7RRh54VIBFggPcuLB6VogAWMGtalXun8m98iyLastZzaQwBa
reoLu2JaZ9BeF5s/MafgbvhUSKdVFbLKwfvU5GACleHsL2lsMnYKAGnWPGKjANFEKfRNwquwaKsQ
RS6/KZOkE404ztrgVP0cCTxNj7F5nydR86G2/1sp8YQMykQmn9TML3h7cANjQ78tOqawz+cdCEI/
R8KLue54EbJReLyRv7OaesBQc7coeC13TtTLDBcx3LglZsT3Ux2H24Ubl7O5Ba8jSOrmB5S+XzD6
nta7sZOvrAJp8uASntATS9c8l/AghnRu7mj2TuyM4ySFVZwj8hMQolf5MSdJw2SnV3fF5CSWjQHk
s+PwOw4YTLtSd7xsvmejn4Dmeog8gd8XxHrw2XkgWA5e48TsjZC93IGFiC1c4jIHoyyvY5aZnhQF
SBiQ9c3aGQAtcqgpxtcdsMrPd6a5AFKzWcE7+xUbh9mkVT5rEp9ulX6AfK2oNvpd6H74BGlZryyH
QlpqJEeYymwjq4r6g7ElPaA0pOTfb3MsZWvfM+3um7pv8MttwPODLKcAn+2G4XX/goivwMuzbL3K
0ThETC+wRsgOHcQoAtfxvlfOfXh/Gi8pXj44VseFlGuFwpj2cHoYyBazOnsFFDtLicZ2MTUI8mXg
TPzhDLYyCmxa6m3xPkms2KwrUK4yB7CNSvw22ULKacYhKnwviazoRaMY9AAhusKljhBa88BpYd5E
iq54X1wlcr88KEUuHMRhAaVGGNVcIlyWqz15ad3WT0j4dbJVSiTUmsQ49A7+UMrgAh28d0daDaqw
5EgiRa4F+yOr9u0tbsorHxfgaa57z2V1RvptPJHqT5oqZ+v86X9plcTHogNtdxHqCwUcP1DIW35i
717Gq8I7Byb8E61FKKkSt6+N6TgbF6dWypXN0xEDoKg6C/msDyKuUfxUKaGsp3r2FFQwzwcEvmZI
kd/mJPly4B+0wUT18opm1zC5UmPWkU4ibMB5zKn0E+E1bH5iznaB+FqU5ZKgn9nV+VAMIExHVH9P
tXTULPdPr7YIrwiOt2qAJ0U9jlgEZXdWtDnVewVa8R1/DpyVGA+sLVmyt3CJOg8Kz9xmhx+NeQfK
dXyvfB0nnlfi+3ZXLz36vkM5XGI371Fo3qx1qLx0JZLOSZWs+KUsWuHQBTy+UwlUzlfI5CygfSob
xt0g21QcyQqGT66DH73Me6K9B+xd8GLIPRmM3/6YuElyV6D0l6wvB5hSfCltGW4h3CJFXSzWWhTL
6i3Q9nH5D2BHJzArQ+87Jc3UtM6D9akiBp8glgtkfx3v2s3MdfcJwUELU23LPG8dkmldodMnrM9+
ep3BnS7sC/5dJSOxT43C+g3Gb0EF5R/Pl2F2n6d6dO+FIJc3qGsn00bXuya8PV3JG72yR7LiLsW3
nFzsV4NV7oXFUkSTYFGeHHAYpteH8nN1g7mVcs3eCpH0Cuu+0rP+u9bQp+B/a3hsIog7YuXNGwyv
/0ZJARz0SwchjyIsShmJBgR6D34pp3M7mcb94UX/SqD9/pJbSAXAMdFmv4sIAS9CXHG9IFmVjs2s
cSkCuwcxTJesws7LtkQp2fP19h2WUGrOajnJ5slaT/JjKyeyCU/ahVWft8nI9qJcvHTYmkYhD+yk
UjQpc3OwCpNohSHMSlo3CYKDb3gPDSHl3br++srhoPbMFM8MqG7H8xjfXC3+nY0yyJFdi3n/cwXI
aYrSY7C/eOTsOF0KpnbR6s40WWRYA9skST1o+LC86XbUsmWVYKB0ydWw/WrTMphspV7LrDjGT6cX
qytgZezBCbEYNbpryegGsNvJj5c33kEEJ6mmafy5XbFzoj2zgVXVdcX8V7kXL+src5+Z3GdJQvNZ
kb6sSiGz6/bLxeTIlTLDas/AEdwbSMyCFYAIbMgDBQhHXhMqvYzgGnh+d8s2rLMe5ar8mRXTbTnj
avHaWyrTYrWcto+MWq1tjN0CEjMEHNQhM8KwN/ZlQ9GEtpQGnnnDBj3D5sF8JZyfb+BRX265aiQL
xisau1ZWTTGz/EyBShNXd5RHlRa+vOGiguBVRuk2r/OEQpMmxsavEgXyDDIVY7+JZUWE3O8SyfjW
Hlztz+4XAX0Ht8Zgdgot8Idt7O74Vv2430t3gc1XFv1jge4+SzbQoTzGBWcQPTGpgO1nazbahnjr
aSwSfxmxgMF9HEta8swigmfQGudfYxyaLcPXT/SL5dd5idBWphdAuKnFq2uxroRHnh/Pb6qhiBEe
cqVboyg/r+8uItNCWe4VvRsloJ6VHaGUBVqtGDioHaqcDblK9p1urts9zT1N5X2EaVpohiWPCu9S
Xj1Boq/RFYuNR6LO4ma933QP8CJFasGNQK6FJPtlusQn70INkxwa8p0s05EnNOi7xemn1HQ5CANa
B/oCho8w2jiMlTm1uMvCtNmu90KszKkXYQeVD66tSeQUoarHSOJMX71kr3b8ZShWRhRG/cZtBFk9
bChWsflL//ukW92UYluqpSeIvomkzWx7DMiwq8hW/E3k0H7+M2A5BZsBeGqvR1nxCauHuP2+nfmw
Y4scQHsY4SVgb7IrhN5BQ9mqHdbB3e8jiC7d2BXIfg/gttICuKgnOLJ8oY8uQYAe+HOinw97BX1s
kH33GYxuZcDToQQE9ZSu7QklpfTvx6LUJf0JqX7qiJubXPliQpLsom0YAjWTszFZgmg2UAaa17mX
CiuWc4EbiDRgh76ZxcwExes91322nsNcZUTzLpAwjrhkzIFaTobwKbowCjGipnxbfVIFYKOo6Pho
wVQkwvUGu8/Nu0HOSmb4J/DBeRrYmTi4+v0+KLfHNpCGngxbMTVuXh9Hyox9mLXpltV94LJA6+33
YTu81j4HJL8mNOtDq4gYMwvMbnnIv28ldU2FCbFBnB83EFeG5LJv79QSMwC1CcPLtZGk2TIRfODf
yqa4RPsDXPWp87BrieUbzYG/t5crkMyaXbvnPznzbr1l/ZTSYYc4pMdAjvPrYzFTh1ilWJq7KPX/
/x6GnhSvm445rSK2R8MA/7qHQhvJW4/zoRouYWaLh+3JC1rVWGJNj3i1ME88fpYKvh1HBX30Hijz
fty0D5q1In6GUSh4OPp68eMvkFf2+NLFjVWbtbn8TZiVRZtfWXsb5ngM/+AY2PXUiCJTLC606MLq
kZZO3UUFgQDX+uDmOVcdIpocB68R3ldiDw6CdqNitPKtUKwVHAIG5AF62vbbZGq4sSyRm5CxdERH
wNjcVB7xcBFBtjbzDkHBL5As+0rLcZgOEa8oiHujDF3yXs2c2hH+nL9HZOPRVjDHt26e1gW4VjT9
Znuul8LbC4ktYZsXosJB2WD70L8kiHabvUKuwXcfkh4iiYxCV9/6zHunFlMnFBNaZd68qAB45sn4
4q6moVnBPvgJdyCpJmigIXk1aNKlDvsjuVb7n3smztWc1yoJdD1TRYtJkFiIRAACkyPLlPNkg28a
zE4XIL8DUkj8YsTyxpKxpJjDpF5RD/t+487QYkWbI8BEfh7B6o5mghIpIdxWbBxPfTL37OrK1m9p
1SlN5/ZL3JcIuBfzDSbGnAQ1aYZuaGc6IDpyEps6EQpc/bh2nr269Pez6MqJge1p/doo+0bIEwPD
cUCb+CP8JDb8bMnlcG8jJ0hXQ6wPrJoctHAk+xO8HhwXgjr1B1P5U7GoxEHgQWw8mkOgA0PejrkA
OhkBHrintECanLK1B8V7Ga5c6B9b6e0jYOsaHWejgNU5IeziQjmK43WRhcVS8vXXFLa7v0cHDP2V
9yNZvoZhreXd+gqzMmASnVmI8bPu/A6u3rJcHOHRoHAel6px8vftDKVYFLcYE0zrHu6n1BVyfFiv
cTppEh7slK7dKlNh0RhZkw4Ql7j8L8/VpRzKXafMoL2axIn6NOi3Q7smWt+QIzsq7CO/OTm3SBKm
QZtMS12kUm2BvOuedqUaEyNcVc2psX5jIJIF+XIgEvmBoMP7qzTsajeKHUq32I5/wbhfoBUd2ohc
pOzAedqzdLbj2vkGXxxWcNumiMkb/MEVy4BAG2Vep18DntZBf6IwDlHVzYLRwS3zLRQiXN3r3zeB
SClrUF+hwGMhMXsAjTONvWRGKWJ/bB7iSdt+XpyfKJuLx+qxTFKe2anIdkCIOBMnTqYnGDXSaC4F
pgacXWCUXZIQMsbqN2N0PY6YpS84zKknwhVbxAQRiUnHSCDbVG2ZFWmPidedO4m79uUdcMjLzLds
HgzvE2SFGAe+oErba2jbfZ1901cxpshtjC/bQLf7sqg8O3uc+nOSgB2akz3dSZxcx2IYDLiw1sSM
zX+6OOQGd+2B2rSxZRVdSzn7T2XqlH9NlUUdz0yOFDdS1UDh3YyczzxZTyrLoq0hi122ISPYFxSq
REg6rG9ktK4D1HDvGmoM0q1lchPXqJcopFBgeXTxoilFzRe1WrIn4t97ikFSyf9cOkTJf37Rt34o
O2SbL1AYuutZuaqdp1gdG/9UQOBSN4DGcB2yQsjUkIUYVDFD6i2rGVosOsEyu4JYdHp4KNabLRA2
fQRF0qbQQ8mHkVkm6/wBMmsmcRNkSk+tRQGcqHyNksJ2v5mFTGPcK/8aCnEF+u3cyKGrL/KBccLZ
Hy/V64XmG0YrSPNi8tyOZ8NF8IwNgXQ0NvHqT21F4yRcTr5bJ3FOBi5TRrpcOx8StcpejdjElGx0
8lN15+PoJhYBVGRkRBEZ2Smb182Y8iNb7I5mUctQfN7hHVraxic3B3G/zSjVl1PrfwEgnTnEqh5p
NBDTjsIAp0FK0R3Z9BGFjgEsc6ONsOi2vgcQ3Bn9bDd6AkGxO21q6KCG1zYAtaROqJG3n62hJA6E
5C/ctGAZ3ru0byLWDYw3KaFC3x8stE9I4rfbI+LFxgYXbS2g1RqLlSjgdfsgn0dV5LlAQ5WAhg6Z
kvaI4SGZ0SftSQl6U0wIdmo1vvOSK8WRUINjAo8/E/0LFLF9AceyTF7QXwXJfqGCe5hJmRy99qGm
ouJ+BK/VuRltynDwoIltUVVzaxJFSo5tQq7xcb+lAFKTiBicPCVRjLwu6MZxKgXCSO+qmDBINeYA
3a1Wx0JJLhLiEaxu4MxpaQ4xeXQPXGETPbHp0XV/UDYL2/1eFIj5tLXr2r8DhBqswSL8AFLoe+9n
5g0m3HrZaRJxF+kt8yatVuZ6Xgtj1mZ53BxETdL6qaSRytSZbXJFNcYemg18yTi6HRSisqKJTRIe
J2mDoCquWzXCOXT4ibNiycjkBI3A/FnWlkj3Pn4JGvdwYRhSb9epuz/wkQc4nnB9XqW6HoEHu/Qq
2ufMnL9EWXltChNMQfo9zzE50P6FBmedOOwtyOPlNrgfvDbXdf426QrOfRf5WlQ6XJZGGGAk9iki
RGdTRKEKbIg1mnR6IekC02NzFYU8WoQz/YPKIqsv5GbPUQpgKRSh1isbWLzFM3JZnb3sflsMcyu8
fBxs2N1yEIZtuJ9Zy3mO+L0XKzs50x7536tKalAPnD1o8CUraN2HbpQ1FrtksArongOitKt8iZUF
H63MrRS68/5VkPCCgcN7fQOOrcaXhCXvenrGiYm8co0OURgO19Y/JMTKuuUWSot1FBNH94kKH0GH
l7V+/htJonOQKx+AquHb71Sw7bu3pByB1NJan0wkJj/gmd0mmGwOp2GV+YJ/xWy2VcZuHtLTMAB5
lvlhgWR0q202X7RJ9c+aOyBIKLnJye1gfZEUb9Jw/s3LS49q1VDjer0Y8S1aYWlihWIYyKE0E4fr
GGeWxGuZAKfvp5XY4AgC4bcryBpFxxM1NGwMNuZiQ71Sv+vTlCBkSaQITK458NTERd0nSX/a/bGs
BMPgv3afRGtLZfWlj1ek3EbD9bSm2RF8v199Y8SSM3WetlK4yioHJJ5ItaPqEajsoZDPjF2K+Io7
Q+/IWhxMrSV7vHR/2SXZ46vrOwKScjsJ35ZNU7dKoYdpnAjwV6BZwXsxkYkBluKIvwXCzH7MPOkA
twmhlSD7OffOM/o5sTztCXwHQX9yYEfDWzQqdJtUBZ+t+hfM9uX9gSfSqJ7eihWJp/MknnvPgK26
49vu/4Ao4pC5zidGQkUTgcN8GmzRNLtZQijjbY3werJtqzfgHNsU6OkVhMziYpsrmMHt/G4A8HT+
bMWrVfhl76TmHdfBmRndHtzxTB+qT1uqMgJKZjnTfaUrxpj6bn6TWQBJsxaYZ99d5Lrk54fCsoAD
XFoa9O0otETaot3uU0N5P/7+cwxjtGNvop6bnscnjDf+9k0zY3RC7V5DHsRcRgzcEQJfzVH7HhMk
+6Zl05XJb7cI1ROREIeTFMH6bKH7Leeq8LrKF69o6KOzkOIa3rDNAFtCaN2KospELdF9AJNibOll
G3ONbtz+Vj2SRDqLm9PwnzbrIkXCuOErSOGCvNGZQI/7qlGe2OmgZWAolce6dUxmd4i1Mkocppfj
KZVDOVJhs8u8lytz2g7gbvUQcOIcEKl26Zikjnnf4aEWpkF5M6wZOiRgDlv0rn19eOgUvLsCcK6Y
TvvrwL+ARh4zoe3Ipb4XLzXjXPD/IOzkvQvLgnYunYJ00KrokBp67gu0KKPjh3pIKDJjsxIvlUrm
225X4/YSkejWqr2loFzbJMQdUTczdiiViANPlTmdyNU9SDGKSCoB40hK+3WRdiac7BMhaWfWIGtu
wklqJ1T6amSAIcAClORO/5Dy4K2b9SDtWU4yO95Qx1TUxN4UyveKc8zwcUHz4pEijqhI9jsqHE9I
napqtgfaY5kEOmMH3nWLw3TqicnXl3HK2pCGBh9ka355rTlka63JnFmzQWMfpeTZS/elG+KUl4JK
IMGQH8yDWjD0AHnr6mVOM0P2gwSS05VlLaoFwElx+Ri9zcwtbAX/17fc5P9xstLL2Ayck9+M1quM
HKpuQnq3RSMVKSYRLz8nt3w9UExG9xh7WvjP6WT53v35gigyRU/ro82nS9ORqcwnl9t3Q1H/0tHn
2O7NUcIiB72gxBAL8SuXciuh5EKm9zZqHUEoBHyjEwGSnSXqbc6bMxyQ05eKfdTj8JgRve/o+bfl
xygvqoF73YbOgENo7Qzj07w6ivBAJesIVyKLghZSi1pGiLJW8bW2RNbenCXpjzF2UsawLnxLEBE5
jWR8o7drgNt3Fn6qz4plFdTEY72y5w/dy5jcBHpOiQnCtypnfG9CUfvFd3mgCgQuj0OYhm7txfvO
FkE+i/cPOb7RmAlgpheLHPaRuWH5j1faLPXmwjxcgWBhdx8XEbGyzZLx4OahUxHgXJkOZ4ZLQojW
E/oR2cm/cuDlzMlj9qbLmh6j5h0P3KawJNgzuCRRja5e+IfsJPxw0PlmcVKQ/S7qqmmkX5Um1sQe
Z/G8yTUjnhQ3Xuc0c0bT0VKUx0Ltd3HtYgGPv4DYtBT3sIKyXnMMcOHxaeSkaTgAk/yQ2k02Pf1C
pdJo2EUoo7dPWMamoGP3iAL/tJlJpMflLSZEYPq+NWrBIuX66W2r9lZQWjurOk3pJj7MacmGp8uW
UbqfzXdclFjYVbGeVBQ5GIu032JGoruXsOf+dLZfPNeMakYjImrbslewgl0fxt5HTwNZ18k47bQ+
BaM3RKOl5frJ/03MCb3f1Yh9p5VOOHRfjGMdiXwpO6IRWlSPZkgCQ4wegnjvSfACBr51mCsAxSvV
kq/BAPAJaypdcZPDNehkJQMDOLZRgr9wUte6Y0la5ShmOV1FsE8Rje+rIBzruAykhho1GuzxCysS
jOCyeJyqao9h6mlCWKjBr0vxTprJjepPv4wLJ1zvoAaML9ma5LysPyrHyY+HbtFy3SpVDpWQtX1A
yUFqyIM86QDrOPiBM2HLtojagR4BNA+EVrm6cdAUu9UbZY0nf0k7jZitmgyDL2phf/0DnTc06iuk
Vi0BlsEQi2NStRG0Gvee8gbu2zKMJBP2ZiwevTaVYjoJi/tbefq6cjvKkMzaTFyNCFclj5QP/IK2
QmrQNp66JG9jopf7pTt7WEQr3L85fGBK2611Fhov8UyNVpilQly5Ml4pCyqf7tWj9BjJY87bpjtn
vRatZXdGKedvlc0taU/EsZX7wzzWs+7ZIWD42hYoAnYvsqknXQc3RANf6qSOWRBnRGy4eAAD6Wqu
C92SXRHvd2gATWVdYocVnv1VMZClCPgAlurGOgmnJH3A8XkfjTlgZIkvHrfhUXuHoetnTPKQsBzh
xNSUKA5q2wt8s6toZwI09JkqES5G/i8EaLFE8BwJBOJxZ7XnQTu50JD64GZAG5Uenp4DHXjnINAb
Zg0QcCTZ0VCe5tlFRDfuRoMscoDR3ZzPDYhxKAQ9Uzg24L1cBv6iwinARR01oSRXo5SlZceQMEr4
6gIY2kjunAHEdKI2GJzvEXVDN84akDymxRfhrA9xlQlsZHzCXw+89HkpCLTxsIW5q2APcnAt/5Aw
F1VWsE9xnjiWZKm9muqOUsvRPOR4CAz6MmMw0M0hZvyTE2UzXQankv5cbEWZPHTwggZ0rOP8jILI
yFKBoj6565rjuqQK9BGnzG0WhXbejP9mIup7nB7pny5+hZUQTSlaZ4p6buAe49Ng9ilHmGi4Gm0u
n0n3G+2lROy9Gh+kzj7BE7DgFNdXQQdIrPQi96squ0d1vW38ZvEBQs6x1PxRzaGyigmd0z4aJjS9
Nm1tjk2LdgY9CoILPBm9rAvEU1f8Fc/cWO5t2zA4akjBoa1JeEU613TnpoV7rfYmC4Dk3EL5yuUX
0Z2Km7FYzOcT3eyMMhF9dt+EU/De3I49BY8p2ifPa+FYeMa2ddXACru9nDrDbCMrP2lWjPPOTZDR
WiEEwoUoSui9/BpdzR2iaDTwX7Pq5b/1Ve5tAuJNio0xm0fDIdKo25tPCIKFoYCzZ95OAAmHlVuq
qLJPl6+5Gti9Osp/TQm3MFb89qrOL5TTClZ6FgyS6VNSiEydwQUkxkdwqjL8YHacTdInDoGoim11
O9OFphTNNdCZ6IYtDb4rdV1lP0WSKfca5KF66suhwQcduwePXZyb3B8yJz/NTOhULFNitTpRnDpe
pqd4AfwsgUqnCpW1YVjWw3n9vxd8BDKQnzrRs27rvmdtwo5HkSr2GW/9PGmAzBAf/qluLZ92j9Lx
L6QmLaKS+ohpuja4odZWGYeWPlsY/Hcfsvp45SqTeth2sbf88OX3IQg7hrme/wqqDjjFBOMb2McB
WbzfU/EMLpx1o7y3kstMIiPxMAN5kmR+mTGrRlR8/WwZElUrm4rugSMO01ujUACpHbzXsEV6v3Oc
KSQbKl2MbvNbyYexsrY7UYCu4cS87HxrX7MrFncVqVyY/oWy59g0i6aKhiwQyWa1nXeS2aKCQD6t
WJDVDafRUSLtf4y38heDANFr4QMaGFWA3uZCjCuc7GM4cigecDgRMxy/7UMbr9XKH3c/vX04rsrG
BbJmYJmzfqNHEFLYXr5Ezd8IGnHbMM7PwmqsT2Jymi8eUHNXKyEfx8r6Qt6iApkkG0kbefkv8nrW
hb76oZT4fIblMDmIoM9snYLNvdJxpyFXem0mTNgZrQGFdqaAIRG/ddohm5MNi8WJze8Yu3zERivp
toJLM/PM4qNJhcnK9Oq8DsPbUDonH2RzqYcsQlgA2GmchRlktA1x80oH4UWKDZx31xqetaEMs1w9
6hveuXG9uiFPgEzX7zPXLa+vt9BwH8OrEavGjfdlYZSRubYurXlKr82xIy5WGxRHjxXJaYZfURZE
5kyG4SX5hnVC5z1Yb9UjJj1yJXTgHvc+m73R4GyjHQWJXzFikyLX1tE9l0z4MkG/AoAMz59fv84Y
JxdU5ok7Ejn2NZmJ2Aq2wLRZhNHKwPyxzmqLMgfGdlhTngZ8E134QqSwOfVS4C32mgt7JXWAfs91
PJqXvQL4c6l4KmF+x84slguHfhusX8zb78DzsrEjGYrcTvKxvgpzbtpmAj+Q+DeUZFkbViwCHczs
4bIUbaSq5rmdel933m8IzX6BuR9Wcc1dvJ+i2AQ0N6ulZ9GLQ2YcB0DtfZfzgwA2svVHhSEFT7bo
AxqsXF/C+F0WYobV9ajYxuLNlkN3KYGxqajNIP3+uk3tZAAK1LCqCF1gJ4KWT+o4ZYO2pMRYLZ9x
IPgq0WpT0gOU1opHM5fTzIhL8sJnXc0pxihwj5D5NGBkrEtHO3n7tl1q/zgbAVyCx9b2z5YTYFwJ
XmV2aNFp4ra0CyknPPHsFSSopUhsynDbX8JhseSTIkF5cdaX+ydhmgkJFswiv3HFeqr7lVTdX2qb
LPx0x5z7MQclcxDSsCk0Hmnodl5MR7tGf54NCUgHvWLpmt5XOFc3hY0Gd2c3YhivL6j8jlMr1pkZ
6UFC5pOYF7vuUFhin2AcHCqbvdpLggQtasBXQjbGAp1cFQjBOohI5j3Q0GFYXQ4+l6owivEgKSLU
9Q1UMGMzJsY3sRSoG53K2Ul/HmSq+sPwhCvxB0rHuNj2yZGHWM0Pcizq3cgqgGzlXKIi17yl1Ieg
0Na+9GaP1psq3ZOhNtbod348qeMZ2GRW88WsGwY/CgkIUbbPQ6YPHsG+HzBZ6hcF1KNpzMbef7Mu
J38C9avq+Mt9w6fbGR0jUELUcdFcr1Y6YFTThGVGDyjRNdHYrDDMigNaP3QOqnNiouiTr0t3lsZV
U624Wuw1ELn52g1fzJ4BbXFC3eU1iQKtl4w9/3JYTvF5IKkgwLouxfSs7/41P+Ak5pTbPBejfh0F
tBAQKdRk7v2efkMbtFlJnIr0zAxX83hzuNa7MkTVSTEmyQwerQrYo5FicNLokXYx54499Xk1/CPD
ILLb9cqefalOVbtt1hpq1tzsf7KRFc9aiNmoifKL5UehcqNdCMEQfSDf89Fyv9/NYQEX/UWdaxWu
oZg57ncmVIhpA4JN4Zgx35Js729pS5sb6mq6AdT+XLLrtFnyKHkWpm8lLxPr6GQ8Cs7pZIipJlCm
zYKTXcs3Id9mUfydLw5zMRGc6XDSuVMBpCIdMUQQnBMV1/18lTL1d+WsRkKt2r+6FT/QZ1weCL4A
PjqYI1Aeel5u9daxbHpDgVGz1AnB055yz1tRn9WAPCfvOmyWHh3jsuFLfPDaysL2wL/zv+Y97gkn
hM4go01y70AcR2aKLXuikGAhCWdLoGzJtH7y1ixC513ym6LD7Vk4X7Y5e8Bq/toe0vuMmyEgFMzv
Pq1D7t7iVRkzdIdSbyoTPYtvyTMqI1pb/Z2CSaqYiscv1ID0hXHMURE9I7byWuJuXDxTrNQxY3gw
F6uWL+pMhQ456AOAViLl4Jwb6a+zQHjRkA3m/YC9Mq4Olyia45gkVVcUizy8XxHEQF20lI6VCC3Q
iTilZEVrED6W20apgV55pRuEumd8qsXQpePVLY5IYEs4nmKq1AGpnLAYvYQa0kXryu6Nbj1X+a+b
tD9LpF6iveiomQUjj7H+zMWTXzQZTJGANbgS8r4S17DNU604/tExwDyC5GB+9TqXuhsS6FfchjPe
DeHl4+aK93TVA6qilXkePSBXbioyrSlJagprEwrBrVizTS/sHTv1/jfGaAPer5KuupZGleL1WPVv
LNjGVBtJjrgryVGISyO/5zisiDVxVN/9EPHhD18zEORHMwPi5CcvJqzxeCN+obxEe4165LDQkejH
R2G2/KGRCzG9yTQ3dHwGS7YFJLC662hLd/lzFDhzv54dYqzQm/qLnmR794RYywchfBhbMJIB+H/I
VP5YgKZydacuyXMF5y8Dcoq5mREOxYchChvfTrLbjtsmTxcAX5aDRAopCGgHN0Vk0griemBFuqj+
AkzkRdeKBYmNoCVuGwF3Uz5PYamYUStr4kHyVRkzNNxoGvzUknq1y823W298/Sd3h/tdvR2ga3Ae
vk0J467f5KO7avrRc2hs97N5FID5nERXjXBKF+wBQnErXUtUsk8BzhtcWdvuihuzZ058L2GMD8CC
f9ho61cUmkPk8ODdlx4UMrmbYA7G72nYXhMUsIxwH2SsM+1Vp+CrxAZMiEwehrgFFMpfYLy7FHLh
0P/rz0UkDjJm3YyixDynYqhIlGSfUYNlqG5vns1io8VmWfdyfF1pYQaNU7v7waiwRMXiQpG+IqnM
tCmU5hlIs/q8UmaHhFPZUPLppGGsqDP90G/IxBtozj4Alg8OMTiZrwQoYNXANOBY9etRfMAiKoWB
/xC3QYQ8ka+iWHbWCYy53eoMc5c1SJZV0rihXnua6wWDdnYLQbJHhk5I2em+DRQwL4aw9QQsZN4W
2+NFiIyEL56T1RsBA/udV2jG1CySje7zUZnA4F8EJDcv6ab60v7tBaTIvFJvQEjDyZkbupw7dfhL
aLjCwnkJmrzFBlV1gCKaboXf9H20HiImNK1al39laAWAAf3GDJJmgnAzlyAMwSBcmlKuey7xCUPu
gQ6BURJVrlATrptN9P5lNUueZ6k83Cq/C2zIB8MpIad2bHVm/c8G6+U+buo+97WSI0uI2Vo5Z/Yt
8/01PEc6fJDGvbspre8KWs2bnz3/iuh8PNYt7NGeIxdbpROsg67zo83ZN4RM0CGGD7ZeC7YV5B/b
RMIuUJjAlNPzmmt7k/OlujXng6HPOH2kNDF5YgmE/8zu2TpKb04qu0360oI3sOdLTPcLv0DQ7Czz
OhpWrMcyrhJXCmHGxu4jpBzeR/biU2F/3qYyAFcg8NK/AcZsBY6OUyGUf8Z7XOURzZEWR2A28hBR
jMn8VLpNkH9ETDh4OJuInFNtrE7Vv6rtrwJaznPbwrUVY00gzqB1Zrr20URX6uEWac60dA350dRw
8izMlbFS6B2WhLfHYphB2mD9FEnbx2jeR9w1Sc7ZyYza/n5feVqz+KI7AYBcR+GEfcSEXxT4PunW
3nR/ZjgH0PrQPvrdLtXRatC/cfD9uRUvyckHrTSceydwe3w953mKAU97kOyRyqecvzGt4PfYI/ah
RtJEbd/liXZEVb8FLR4dDTH4IV6AyyyFSAuwdUQNyORlSI7ihGNUWDPVn6Z7npwqdQPAa9zYKIxY
yLSLc0ME1o8OlUXeNBl/2e2coYXx+ycsqNrE0jOhXwPemmUs2Ro5HA4j9iRM6D/PMNyj5Gcxzw+w
59pe+N8D0XXipMx7IVsOgXtjXiz7akiqRMktn08CrUjyZ5voPCAyjOwYlD+2Y4xJiw2kSxENFWYs
+1lTHYmVjDf3y8+PTvShtNNJEiesA5XA1zQijd1OK7yPg2BC+8hwDrh/RtgN+MRWzdQs2uhS0q/1
P0hN7XBMw7fflnVO8wt7FCIMyinKgiCveVxGeOsTFW3VvfNTHN9zLrBDI+fMKirVRVbswYXWyXg4
NO8ah7t5bhv/g5/Mbca7LTej/dktH/z1j3KqQHGyHBUHdBXgMTd03z6Z3k/v6KB72iOwv+lrc/si
mVjBU8DrbiRqWioWRC78kSld/aqV1TUid1M2GO4SLytgsVFOTMl8sa/lCWqZ0CRzXt83nXAWHN1A
ZFDFSmyumvtONOOhwb+hbjB6Pa8ol/OWbx0EOjk2vMneXwiQYRmtQHtegYK41Dh62CaO9jPsDfqu
od2NbZ//t3D05yD2TiturKK1tK63gOENlH2WN0RlkKRv96Ct9C3egB0uhTdyW3ub9zB/QVhrXLZm
dCNU3d5AjGERkOtdIiaSav3mGsfQbHAax/StWtoMuKVe2YwfbZYGvm5iqupZJygLcFJmxeHw5v/w
YwHuxn/pg2MUNSTz17hbIetnbTZCNSu6xjRcBg1q5ZDi3VOduu2HrROVWuzOVcMAqI+ZaNeHPotY
6nD5UWxIuUFOF22UJ5cDsy1jpnBwF4AOGvGMG94Qwf5FPONEIRnZGY7drDCMnbTCWFM4x+xAIRXP
UcGvKRp8/HtTE0zQLlxPn/dFmBuMNJDm7qWb6su6vJIpc67/4115Ntu5U9yVJOTdNe6xVKIChtMY
D78ArnwuuSd341nAAZZk99oLoMuOtfXViT/ofT1+M7pabqdx/Vk0DuYkL247J9+VjiApwRbmmAGS
vqjTGr+M0vGw4t3TUUDdfUsR0iKIs06sWRtJArrtfGPavWQ3Tx+r2SaGOSt0Ei9s0b0Lz1+Y++UW
uz3CsuLxwlYsHAYv6sk3LdZll1R5lRncTVSZFJktextmXdOiC62yHd/etr1sUwboTlSyLGSJqOwE
jNjlbQ3sHfLLCaGiy2sWaU010h8cuaQI9o9c7XPUEgGzkMYF5sZFRMMyIpLu0uLOF/u+YkpFhpjX
5zYYBbkDPInOIeDsy7SLfwjHpxMv1/8KJtkDvHpNr6u3rRIat7apfi/Vqt0Ia3bTJhMxdIGftdcM
ry2bimqhpAQog+XeUwTLH1DN+zJKoxzlVVNJ5V9aD85lQk0O3QLYsfrYQwg1IrlAA/XhyB2luPM4
cCyjkoBywRmBh/zQK/f9Y7z73RjmuHNTmn6R3bDEglo8yuGTqdSKEWfWsdAzyAnazDnGwGNTa5HX
c1pEjOqG+3gCTBIKObMYjfmIKoKPu8D8QUiVccEn80LXQWbNFgGP7fZSW5UoWBQuGHAUUl0dDc4T
/8YsdAMXZ8DHlXZiRBPwvtiXsNaBrB3raU0sKSHqi9/orenzXdyHKUfS+eh/i4Q9CajTN2POQxKR
TR+ssg3+KN5bklf3yclgk92oeFu5Yh+PDpaLnkVVDveCkF6fEKTBxZnlCr1JcUV5OsJokiJ17DiN
hnHLkcd5W7rvzunNkScGUqZ+pPahTd/7keC3raSeqqSGQNi77/ZJh6rMOFmd8IXffb/KXI/bY1Y2
dwvGiqZpSlLzJgR2MlcHqclElg+vR/KJ0Nx5o53jjxuOAi3XybVgAffoG/TbQHZSV8O/CNqChRAd
wIO0BZwW4koS/hMFOPfXvvIWXOf4HzaZkY2iCAlnGUUSAILok0SJxcpu3xj+WN5JSfCar+Humy6u
yFkaaLH0yjArOS/EGSyLLRsCgDnh4QKvGw+nRlXiRAwolRtidBFV4raPSRGy4ektKB9UuVeHjhFR
b//VDvGWkSUnNR8uwx63o4p9mPA4YZenIWLCbRISMKIusl1enxYv77PRKZX6i2UWpFZsMPT3uglW
OMbFe8Oreu14OTuxwQJpMozWp96vhSGlYEJIbzKs4EsV61J+1JKM4XxT0EyGgo9WWt48AXYcrT2M
EIWVcbjHKSHME9CTzqD1bHfq9WrIxnkO9QkDbHAfBO9Z4onslF6nVS7qBIiAYSlZWdE4mBKEyf3U
mqNQ79KtmUsU4VLzPqIZSNL9N7tTPmwNQR3YKI0gyT8BcB+KvME8RQ/9zeSA8h1/z2FWWFolBhKC
X3bChzmFPhazrRLb+s+eU8Ibi49VhiQyq3t1dYH61kLxIvdWLdKMHtMDDz31bibQS6iKmdXdNeJn
CsPf+F0QW7aQSwrlZ6KgnI/YslL0KCDim9J8utyjqoX3sqT8hBP7DywKP9w5EBjmvKoZ10nP1JMp
orKchDoZgxB88DotrXZuYYt+OVxNXsMc2X2EhgjK46BnSMa/ZSNBye8zgxBBhn3QI33x9/BoY9EU
0Oa2uxjUmLk8xvVIuItPKV9kCpUvGcc8pzxt4QkgpBPTTgZ/BCkY1LwBvVKxibgfKSq2TqndCbYz
wiCG5MCGmWJ7yxpnbSSNgwY/aLK4K8YTtM/rV16XwHVWth1bcaU98+l76Ck9JGXOi3+eCKnGOkcG
nrvk+q4kQttH2mTnpDP8WH0WwyUbSBEd2T8wNtAqEflJXnUjYcapf+wpXOhBuKInThZDWeBDc43f
Rpw8VpLQrrfavM8LXhT3gwhs++zt1b8YXCChR85NrhoK4eIoBBMb8Tk7nV6gnn5qdac6iA7XvCRT
mM3AXlB3KU0gIQ7scoZFZ4rydTQEQxeYRLvGmNFw5M//FedfHhIljyhaUiQJ9Y7y5re/vMfno+bh
35JYrTqTT+CiSqIjaPnV1gT96iKMUm75b/LfsUesC0eNRAoN7jHAQrtB6iWnTBLYmyyM2ktSH9FC
9O40l55WkwDDUawG2eDwJ+Y/N9K2phOe87Zgz9sAP1dmUA3zlzMtyoPZBMDNydZe1rW58J86BWnj
Emg5I/S7InVp6lmmiPC9kQYXHvrCgur2D26t9fEmCkCB29WCy23vHKVlybSLUrMS/Q2u04wDxqIV
0AhjRVr4BsERvKw7/29V0PpRkTpCeeJxXRKrkWCCVZYWLMMBqkBA0DVnchph0GHwgpwkqFLeFaXC
gnsj/sdqufCYs2Swd0V5qaf95jNAZqiufd3QJmZKFf0O4cPhKECPYi94yscYxB7rZQQqx8OM7Zpf
ARnEt46yQjeJjuUjWNmerENDefO/nCSMtjuLDJbMA1GVmlsmTF3slo1l8OMdgVcxfiz4zWu4ocNM
1IsXcBhkzbo2HFZaii+e8owBsTbFHJtZN4MyOvQJGRlI9sMEUQctMU4O7u38cfcsC/vRm9wQJowT
ktfKPIy48Vo3wcamgahx1ALOSlZO9PDVK03vIpi3izp03tOF7wlD+Y7fez3WsOihR2heMLbkwjcA
rZ89qZOXJWkOlrdbusm2no+3rwGDEzyPilCwpEzbSSyK8H+Phl9LC10EUCFd6e6lBvWQ0DQqcFwQ
648tnXDaTrXUfXXMzCBGsFo63mFWvJ8RyjH4LMXHD47DZk45LdFCFck46iq4SZgC0bKWkCUKuFR6
l4ITuM+nVjUZBIgql2wyK1b+q4ZuJ+Th0iA94cJwI4YRiCqJ7oDEogARi2JadI14ZD6CRNHZit93
88OC+Kj1jZcZGfRH/fDrwTx8er9H1lNY3phLXaD7JoRXYydNuiKsegErG9Soc9nXYVAbJOt5sofx
QsMssKOOn4GC/xpezudRapCsoh45Fh29CvZ/XFgPbldAPORC7jhGCIwbquq4l3Gf0PrqRZQq93gA
WZXq/vcm6/K0CpzkAC8GFwLKd5eS2fE7HEXcxcleiwJhkpSe9WFmzdnh6tWIYN96mPk6B0PTQF8M
OL9jMP234YDMxuhP4qVczonE70efRnroQZdfIM/MrRS6g+XAqdnzXdIVlRAyPBmjppqR+CM8a5Rb
7Z7YYE++8PORlvLMdXmF6ZmsABg/Uc7Q74yWH9ybvCBvUepXGzRcnHCuB/znYzcY9Uwxkw8msDgn
AsgmxB5C5bDYOtiJOi7hJWP3ctTVhOd5h+h+70bhzVD0CZqZ1pf51qvaHEtW1ndwubh9O0RqA/K/
7COKbpXP0vU/cIsqYXT+qJJfpaLv2rGQ3dwTeVrFcTtXHDsG1mpNKDILl9+7QZcbQjofBbkiTerN
I5PZA399s7b9mDpfP01FvXbx0HBG+Z5kyCwuiY2LKiBmEe/HPP5GzQ9jMME6eqXwPUUXY7JCgKyC
yH8QqtvaBGrxn2+iJuUOpGwr38RlHqwo+5lkKzfF840zz8btID+2QPHpMMLvZ1DUAHkxF4WG9HGT
ZKlgVlJuYc6QwPP9cxyk2NhvpMpbQ7Cq1kBreco3rgCNkjLk0/wxoNl5YOEUfHnOvVAAhnxtDTes
VTfDF7YOTtrvH5sDwG3QNzFqhJekYYBFLOnykGOFgwh5dbhzt7NuQwxOHnFgxC9zV27Sx3IrVAxS
7/OkipzPEkxQaLceRa8F8EZ0SZ7emnEh6Gj9Gf47cf6mKs09nFg/qlTnt0gPCY2ZX9njlCY4TOPd
QQiFFLNR1m0VULeO5hNvoZK5xpyxndBGPPi4vbJFoT8yV6Lb63ul9yN+6X9e7zZxE40mviRlFtwH
s3K5VtWNU1vZ0gCR9/+CzjvyNhq0solEteT0VrJkEhZtOPwuSpI7Dh5IjJX+Wku2M9f9If8QW6tK
jSzzvVZ5CT962SDxUM0ZZtHGkQjUuTCdch/EpZJpXEbnCMjH/SNQKU2fJK2FkrAalhHEqs13Vnt0
lz8LFzrblkL47IRa7ewMGWU2AKOGl0Huzt7+RfC1mLRmT9gqMffEco3Rs1ym+AiGbu/7mVg33y/N
PK0iHajH4HMlA+ba60r9IzCV1mqOYZ2MoOr3GxbPrdbJwlf3ak8A2qOVC5/jIbKfaZCRLa0hmh4C
7Qs1kXm2OzFMc7WZGNAX9RGusWGzKkFzOrQQjdth978Y5cCbZfcIwEPsD5aLP2haKV+LheD+OHqR
2FmJPDnobDr6TR2l8NWFBwsIYSfRcr5d/W4GCJfC1bqSx+Xvml4FVJnJXxwg3dGtheh2fYFNCdrz
B40DOAOKjCdoTo2Bjki4Ab7ZR7RcTtOipXrCpmdJZ7VqQmKZLqfLQIeDWzmq8amRb67/EQ4znH2a
HO7T0KjF1vpLa1v+L2RXk6ZXGQPhsHtuja57VUnpqq07fjaP3lXNIlKjjtaMQLofp9tan82cjZSH
eyIPccPThXk7/gnn3w6jX2c24+ezeqKVA03TaITMQq0Ag3DHZ//VP25zV/qPzPLDwPLckvf7mKg4
z3rAbSw2hKDXyf2LykEnLzI4YXyxxTWcg95vGGTDS0lljtauO9h91xuvBwl2KQMUw/Mradvmc/rU
OlHVfL+jhRuhuMtV+Ku6onS/o4afniWOs1cLOPZSFz4nwQ/l2JT6RzH1KK7FLF7vEqkr4nZHTaJx
6i+mwJi82SAghcLYqs1ALI3hXEm1n3+oX6I9U3c3q9sRXIyH9IH0XSVULAmr3nNfyTeMRqRUxV04
3jBT//+1DCmubBHTbYkNsdqdMMxdInSfbHJcvTWJR5GCMS2HfzRil6DxztjIBIDP3WUTObZUQpmr
kLPwI25cg0W9OVbauc8KEWc+MMzIGjdzfNmYO2w8BWL2weym9tWvfT8JDcFFUv2KcAbUlzZpqNDE
0Hfbqc6DYcpPPHSUUwlGyoU6OBHp30sfRyLGZbc7Nqs1KDJ1OkUq8E8ghqNpPwAWBTSSR94qyO7g
jEzzsbGBM80O8GqqRG5eBAMnDJCyfYxQ1DUis0AOlEtAmDM4jQsmAk3EHI1Gh6fQ4QgmNzNRWzMd
FWkyq82NzUdSXEXb76+x8A5OXrFqHsihRIJhU15kK+YQ+us8TZwDHlMtqeXrYnVfbdZYi7DiYJ69
qFEi89IFfc9Pr0nfv+88TN7gJFjeY6yMdOuKI6JPZSQphkKV7K/EsscMfJimJ/s3qt2TBdc5C64y
H6hf1Ca4HZbe+t8/pUUD/Zz987VgXiGiTdWy/JMmxyapofwud6ryhUWrhzKpBio950OhMYZXwJko
1YiOLd5Mw1CesA0oandJ2MLp3w2UzJr84XwmAdeFghZnM4J9WvTs6nC9ywRQ76pxo1uSE8WPZe7M
4dErzYkOaXTUx7LPy3tlWumD7qMWQvhEBaY1/zR1k8WNo71kwLQkQXoV9jc2p64LqCMxOb+4hIGW
iqXEBJb+uHguHERJbf1cHhBqDqGwraOLweJUdQYz3e29uobQiam4ezhCZmtrN768nD93n5r4onn8
OhCnBvD9SaESYbJQ0zBvLi2t/2dIHHmTj03hQi3Cgegt46NvaTMlBc3nnenAx2hDV1cHSgqe82I+
20QHiZr+K9HI6iEuCeANzCpWIWtvvbJDNHRIs6a2fJ2IigjkAiVEJW86LAFVsp1Z736BBIAJKO7W
UufgUyyu+GzmTq3aJRAmf4nmxuJV1UNiY0ubpgmSvXCj/nkwKkm2CeclqblrggZPfNiBQz6eq4hJ
V0xwntzxgFQQtfJnmeIDbSvPmxXoEXD2gvQ/Z3YLWlhYfI1lfCZd0o9aJHC9I7iDa/D6WXSlasqd
z0o8JzOFYFza0kGcOUZjkqAKWrRjuoPE3idiLqSiSScSLjAL6X6aPzZ8p6v2aj4OgXnf8fnsyL0g
K3x8YvM5ZjEtSYMW24Ev6PbM8a6oAKcVzAZpTB6KIDikU0UQJxLcBWtTX98UpB+kkL1SZJblq6Dc
tRbH2JjMaLb1jlBsAtKr+VEyuA7Jiyt67+ZUwWc4jAf2ty4P/H55VUea9Wiu5OUZ4T87iNMZeOh9
4ikl7RSGZM9lWLxb9DtX1tbfJahq08t1VCIGQ6P1B8gA3HJJdELJPQa/qrD/kN5V0yNNPMCHDOmw
IdgXeSiIzpkmxNawlbMWYK5RDVMHSofZKjePnDSbNDeegtGgF14+h0ir/XraPdJJGPb/txIHVxtt
vXAqBw9/40hlmtMIlqyFLNFS4dbQsT6zYrt4VKl9hLtUwvm3KNcqu56SqNREuhUCxMvNfcuZT/Fk
y8FDPdSvw2ad7ITABh5wyGs8Zfzu8izxJBWmPkKOXbtww05Y7UtSX5BJ0L/L3+zU2bv3K2AjGCgL
KEzEUCW9nPdaKr+8uyEnm1mcRydn5EqyE5UacYuriAWyqTB2CaC6g98V5sm8w/pspONEoOFpV1tc
etYbYbqblNLrNWy5bzRfN4qXt9xVwzoWXbd3IJ7sMMfS5vFgY3cxa2eKQF1kpDNRBr6HWRavKJJl
19MpLPwIflMzGK1LaXbhXw/Bi+eFI3a7XBgLFR8BdJ/kF7quJIj/j/SwrS2IFxpoS7rOz0vJJ9co
S50Kt+Ee48VDUEu1/Yx/N+M/Bq+A/TRHQItgvA+iiT1hpdteOSZAX26IcZ+Cw4p17Q5h+xuApKM5
vNDSftsl7XvsPTgRE1CBu92pUUmdTxtQ+sCOVHfYW1c4XJX8Pk8+N6sgIAXiIYsMJ1dezkSt8DMr
1Vl6vuV1h8Fz9KGOmSTd7pQcSouiDIpAZUUVoH7YRbaD+uSQOMZpYOxKbWHmJdrgu3NEPl5EfyqV
kIL+VVLtCyzB0nu826yecJC87Pru1xLA1U5BAsnZfBRb9c6xRHYgZfnr/F3fHOvSsGWa19Fmps1Y
1o74S1OYDqZv5zB9hORN7i9lCbYRFh+T2UiBU2d4xAkTalF0M+0p0DQtE2fQhArYESg9DGrlJNEn
z23BaKTv7rciF8T3uBQF0emaCchc9rHun3sfGEaPn8vq4z+zKcKLjlRYqF6IWba1VMhJQeCbC8Kv
3UNVh9G9XE7BnbVH/7P6xgIhMLNImQ8iw8QpL/+WFrrOlJZly7BnqoeCljFWhuVHtAkIMb7sYZo7
macQv3TqeHb9c3a+2qICAvJG4M1QT1ViIhP/46BLaVVBfUyHsyKvXg5h2wl/UjXKsqY4IsAG+QZf
kGnFdBJrNr43vjdAigBYR+29ipKp8XtHt6ne1PJBWOMOqckLcD+wGxid9z5AuLxVl6Y9sPJXLghx
PlxEYGdyjL+AKcgAw5mb4IluDdkwn+EPQMj2z2XmGGAvtySmtru6yqgC4T2RYv9+NSrMFR4sSnpt
VJ6+L1GKI/o1eDxUaouXofRh9DBTugHMiGi0riChMzAvfqB1knKnoq2Hp5JxVgUf7zTTYtcHxOXI
XNZliuFdvHSexZCA1NGly/X+vigjJ3Ydmx2BXlPI6VxRjnrKGYu2/m0JCNNXtBTK+Rsz84B6i388
MWQbvQx2xTHtZd+Hss6rICWQ5f2iPOz6CyO5ISjuI2Xe+wfJmPhabOaM2F/JSDlA9/pHReNjr3Yx
Q2F0PgWNi0kb0EkKNHS8D1nXjqL3pto6PUJM9hWnKD/GdD+0dZhSDZWpdmj3cklMB9rZylzoHEyj
IwEycnZJlz5LX/yn6Derun6mNUcPqw1yqj2xN59AMabapy/w9sO7pm4SmAr8+aUkxuMb/21dCSXj
inU+TrdqynVTuDxARM2d1fsrfYTwy4A7YXvmvN5cPivBrrqBz/5uwPRnUgj9+GDrAJVXyQm/VexL
yOg0Nteat/EIEZ5mdANmQbve76g3sv9y1Xj7K1rzxwcmA5b5ScX0zhiCuQZAgZLNSY85a86/d46w
KIr5wEgI5WMKH5luodMPwnUd8spoBfuT7xrObI5yGfW0jgxCkhPoDWH1AnVxV9L2kbmuz8HvFxGR
8h6kHRo9dicSoMUzMVMSAibGGeq9gZBOJ5QJYlXR0ZumwQzrD9EZlfl5+MPqJbn6HtIZbGPIN6Ns
9zPY9HATOyw4K5qwzm7oqIw2twEzVMoMHd8ZqyipFRTgUvx0vG/AjTFbmRgw60ua7elUDWsplKC5
6/H2U1vxQtJnIk1mz6EvOu4pVjEnQhti1DK7ePNct+sbWgktxC1uGGTsY7sffG5xmHOnGo8LEjmm
cyCyW+NJsg2OL1pTdeBG1WfKyKN+aWx1K7ZqSHW6p/9qH32MGK0/2MR70fzkeWlOubO7jUBLflGk
98lAwiaVcGEmq78/zm5C1CN/g4jLLAmUfEkAwb3Iu4kurmlQmIQfTuMK1bjdudWWiaja6E5ilvgg
h+xhG914N2Fp5kjnug8T1AKeFWFIRx5eHyNB22KIwGfU5zFnRzo8SZ6B4rmMqRv9slvN0ji1/jqI
xk8uhrfL3tPbkFTfch4snJBesRBtVExTn74s78r1b9lhoGiTtiXFzo3Ac3NPk0GbITSYeHmALE5l
GEYCUFDp0PVbFJj+R0FYkAMsIxd7eIXCM17BO1Qnd31c/ZZkJQL23ryaiNiVE3jwuJVdzhM7Ku6u
kocadNcC3BHzBFGUO/S7XY/6VKO0VaNymHHN5OwJSO0uempknimzAqvbiwMxiQmpbzYjyrk2Kc9R
+YOaL440byqu7gzaGGZwffinegNWx5BTVC89RwDWCl0hYwiTkAw83OfHn3+NoQWPjK6SnS00aT5X
68DHSelsDsxO/yF9xsEYy11mfPjctAtmeV8eGaPJpZ02Sq1+gEnFxh36D//H+hYdfNxvETC+ngHu
Ppx/kI5dliR66PDnDhyPKrHRFECKEW5JeWkKPjjMXmyvKA/3wYhRbidzronmTNLsCDTHarzEXqw6
SIKyKjIWlg3llVE5IAILKTYxJLsNP42rMT+ICoab/Tso3PKnH8iyz7assCZWSHmD3Fgiy8dpIB0H
OkYRwjrWSyIEvS+SHOEpl7oyywb8QnJCAh+wpjvfkTAfExMmw9HCdXZC+k0PfHN1AKtwBc0PFc70
gdr+zibs/6Fhw9VRvRwGokfaTA2qzZpO3bIU9KCkeEwr6rPnXM3CjRRatvbAIRa2Th9iTCV3oIG1
I6wFhBV9A22tk63fE6i61kbM8dnrVeipD0UYUiauyp1DvcoZ/3VOoe+/PPI9aV5Xcokn7wBIypJR
wl99GVS69wwZ8nZiqz7MWJV4xazQiKdvaLmfHWaGQLPssXo68cvEKwCENheHsvfk5+LlqNulVv6X
+MW/ajGDU5QVRjabhwYplRJW0KYzJbEqbpqndzMTKYZetdCVi/KhaxOzMqXTc/MfforEKYfsG6zS
A4zFYyMSftl6o4ubnvLCnBMBOlcgo5isHRyNSur7gaU43IdxZWoex44ZfOX48GK/Fv57GnTKzXSW
K235MHn3ZZoK1dcXGD84n/N3niIxaqI/vJ4EBkYj32bcBXdUJsbKtZ/7JV8NjJLKUqvJrp1n9JTF
G/eoAewG8Mi9k6QpCSfY/2Z0QU1qL1X34Now0fP32U+AnMNCnCp+0NA8AkBWQxFndgk25AICu/J6
tezalOpnm6vFex19zpsyStX7y6c/FxC4YZfWpPV8kmbJXL7AKLgGanDPYfNj4gdAXbq3+POW5FUF
0b9JJGn5GMI37LpH4p3kSBCDthFAA/O2d23h1nuWZF4/IniXgYTd70XQd63bSOhSheZgu/Pc5z8C
HHpvWdbu0g9Xz/ObQlcDimln08fGl8EGAMO1upEj63rajLQlB6L+pWXQ8oZPFArgupttzD2IX8IU
tIuqXyhBk6Iaa/rURF7pz7nw56QR1M1mKGU+/OuAaNuqM/knHDaAtAvk7pzfmRMgEo8oOXnCc4oH
Vwt9R1o4P5vvmKwbPxmyTeJRQ+psh4xa4wUmiqcymTPB3nT6ZbEHhe+5tZu3zbY+QrK0+6Effttm
71KrzO6ZUmR1KkSLESmjlmkvC4m8jOQIXl8ltEhlJfndf1RKYNCVGShIWcpd1vwvBWPG+JPlRBr7
f4dgyBWf0+YK3XdUIY9k5qyFRvK1FCvBOsbtMhnMsq0OKRxHhB7+EMvah+CgBf/sFgaNrmCnCr3d
67nedEOGbnIYVqAHYvIwYutcbO38l3H6NnsKoi5Vv6QQSwL+n0qURarUbEYVafxQTb8TW9RuIdQ/
8wibAVKDJCmiTH6aqlyEBFz/8VtVBacqKevTP4f9mrzlvE3sIu2IXUAeVJyh99Kjxq00H1lS8CYP
I40OZSRX56bCuKB8psPulDFZihBGYl61xDxGOHSR/knwVTcYOu03Ctkt66gfIY8fSlQmWh8B2LQ/
QDlATr5sJjVBkqK8/ySw6MQxAL3BXXqwBbaogBoxSV/gUflslI97EkfVVg4ow3xfQADTbVfUvtdR
XYrFAIc46zs+qRJl4k0D0BVwNGdIcG9TLjFD5HM9NKBtjKxoRB0jjc7ya0F6u15n+ZqbLI7oj3hH
P7hEe30xk4pOpbou2p5rsTcpMx34ecnCVaUUo1fEetNiJf/tFS5iyINNNo03SHAaPnCVcyzyW0BW
Lf/gbRoh8UjICLKBl0IxgEmerQ9dk7HmIwtJE6R5gDsaLxRMYd6tPuUkrCdpCTmNvn16E0jqFyct
YZ9WLkTQagTK/tJW1pcGTOUcWO6wYOVPb8teAQQl525HoFHaNqXTO3J94r6ZUC7fZCQGrP+rs9aD
eqINNwmpNqWkAgTanixiyCMH0WGeP7jHMeJMPfprzxHKdJtZ2qcmGRVvY2bTicI4rn6lL9vG2N1V
Z8wYdje/SwmLAMuQvbfPR31AADWw3oBQPn8Zf05rNSbS2gR6kpu4KuZV0ZP6Y9P5iGWz5n5lA7cS
sTJf99kWzpoYUq4ciHrezHF9nWk9RRDsYaeGLRAmD8j3/zs8WeAqamg6vunxS5WTAc9JPXYNME4Y
CEdXdPUbkIfdQOfeqhaMOfYwceP0trPVmHJiWaUEj1fNR8W1FT9r5rGRU9AEcARoo5W81AZ9Hv3o
XDdi95OTiAUUCCONmn8sqrtQKvorxySTWzqIVaDJUJT98NDUt+FlM8TC2LvuOZ/1Kqm/L3oWMhUq
cIxk5keqRWYkxhIXmGn3traQW/FJz8Wh0cB6KaXizwng+8K3IwR9PfU7esKwAL+gdzm20h+jbOSW
EMGWsgFMSWR5AFXrSXhRYAgzkDmksJHIFjVubtdjgxAeUIEi8YT0/m/744zM1M4kV5u3dtRS9isE
Z3KN3a/lt0GMRUY7Ulu21Ejwp3S8SfyasH8fZBvc1i5FcZVIz6a3Knnmw5YWpUvJwqC9ifW4Vnmx
RpHK/ld1c+/hpDULYUWpHek1pNkWUznKK1KPirB6D74bGKSMKgVy2alsbM8U7YUlC+LFWYx6d1ZA
X4T2G9ob0m1bU509LlAtZaUHPvUQGFM1ysXk48Rh0qGAtTrJDF1UJjqUnznfA6dUFnRVGIdS4DsM
5Y8ONDOOAR3QWHPoC1Kb4qEG7L7OKRVMTYT2v3Pj0wINRctFmVg7NtWpztIHgt/3gYHMmGWX5A9Z
n+0VoBErw9l10/6m73uOZOTa43FJJ0CsNDYAq9tuOB5nGaaoZ3LogAW4nH+wth2GgihRICg5R+TI
4Vayw8u68Zx60f9ZPAusqc+mR9py5hZtkdJtLHvc5sEu9hXejbWs6H0CnDZ87IgLDuirgCTReNFL
QF5KypXzNtgsEiiXW00+8mO4v2L702tVIKiTztVuAbAJp/XCKeR/5rMXedb2ge9AyyoS2V71rvi/
uc1bcnhNKpJHd4BtO/ymBrCzYXlYLfm/WLh65x8YkEQ2irqFJWlXq3u9eahFRbESeOtqCggmVMtI
iUswGfircckdswUzjLTPDs25vphM1qDvE7bW49VOqQO4e5Oh/xH05C2v2d+URV3x2ghJYKhb0qi+
qDHcJiY4y3nVVVkQTcNhoMsxKt/ffVPPC8Of57MbeTzlHtSbQ2Nf+lzKCdvA9xsMieOldjExlHyZ
VKqj71xNNmIx7Hkd32Lo2rPlLREEeGZyD1LBK0DAzmN03CFJxtqhHmolADPNdaF2NNRCSy9oZ/1E
MZfuwd8jd9ln9t7Mwg4sIrKAiSLUZ1JA2H9UIqYrqVFlZOZU/V6m06YCylztXuDLQqBVzBNdZO1B
41YAcV7sGWR4Io6Ktxq11kKQCw4bZSFjrrDdXA3twK7JMYyxcyMsrK0N9wKpGuOLCa6RXnVID3OF
tbM36Xw5ssTN7tl6tsrx0WL5+3NQ0+L7zCc3C94Eb9oHUU83gcvZ7S3hvQ1JdpL0xKdWu/jqD1b6
MK0MYR0Oy/vuNJMXFuydfOMxa2AFSL9lCyMoj6Qbp4YoGKlZ7tCF2Nurqor305U81FsmeoyYJf5B
uyh3Q6sLySFNnhZWzi/AxOXsL7MfGzr+vtUK5ES6SfjRcYnVFwwzfgn7lZEYOhlKF/nDpiXz4RF7
Xf+t9jupPZmMLe7zLSRqHKDek2Zb9SHoqddjwqpoRtUmekBx0SRApOiZdRnUTmLZ/cTv1YmkXFX1
+xy8yJAH9eFdErtNu2lJs8pR+a931DqIFdTUASxKp64cjWtFbyEXwJck4EJcjKX8ZCVgiH6nwbUS
nFplYIbqjYjoz72btrr+rfdsF3QEuCPdJj9cH7rs0rG8aww7h3HNemRqeZS8o8+MF5tWzrNwZtSb
f/1uOlYwjgatAXT2n9kmxd6A+mN4ow7qTbEbLo8sJ4EWtX5a0i6Y5o5SjVZSXRYD4XTFDP2poMD0
IifpYb8FxH5JUoMsaczCJVtesjR0HEK2ikEq8kRS0JSlsrxCMrD58TsdMjBHQrUbl1F73RFpWksC
x42GlmG3H/dsjShw9T+n0cMMjMJz3l+EyMwwvqMUU0JDkSr9q6bQ2xdH/Mv9s87SxSvYJZRGUWH2
fRU2ZGdSfyk6f5exZPvzcs8nWSEdPQSzwq1SLmhKNPr9IEfkMSxYxIrd2X+OTqMpssyEhCkbvvVw
tlDk96je9Qb1bkYK2xKRy5SVM7r+Xq2WTfpWikowvGPbRF7Lsz1DU1RSrAxoJf3OFBp52cVgAoSF
n/cCCxAYKNe5iFNc7bpR41tNxxgecK1z91nUHY5BDiz9SXVQjr/hGmu4rs9n26UzbMua0VQPmGzs
p/agG3+ljT7hypu/ShIDyR+5mfz8bzbyxwxGt1btgCULOfRskGa18UVZlPrIizq63Rx3ulrxBWSQ
fo2CRmWe39ucGGA7tuoYpA+0HxNJrYoYvV44+d5jvtbQXQN8rKdc3nFY6aaZ4L1oavM+xwaoTUD9
io5cxTeX9g6kvQFoEemjbDj/HB7eCK/E+WUpIqcqWfrk8dUY7y9jZ7l40Behi2XUHbKd0VTfqVNU
rN0hQitY9qARZHTljOhKEaDARnHRbRpYGF8QuVk9pUUTVEC3aE4l2U9P+QDJUEZbB3SsYOvf3Mb3
mOG4PQaHPiHWRvgErVsWZxA2ZXXwvFkYlXVFFFmcTLPkrIWN0z4ygvnf75WOp6DGTm5pJRAzkGfF
SCB51n5GQ2YRdEYzvFwGpc8g/k4AfMi8aM1uIDh2ei/TbClm5cdwFpUtQ7KLmhd/VZWe2TcZ2F+v
qLABLfa/19jDXPADAjo18ZpVpSOw6K5PrfPjUkjXKsXM53ytmkv91e8AIjuDA/AL3XRDKqF3a34Y
XPbqWnr6ncCwUrOUCgd+ChX+72f3I35Sk2imwQ+dne3T2/hjLGqEy8MBs/tKUVstdlRusiSbYuo3
9TrQ/xrcOWZYfeM6zexL3yLzGGqUdgX2QaBSpT2PlqdAFVLKI6D0O+m0+uToVu0rY4t7lrzvbMqW
6I8uYc9tBrxAgCcjB8+rML8ep1djWn+9If1rYIu9k+PQL1LQEUlWXx2YsgJXYJ+xFjr/UdcjvMg1
G7cFuMTexVrmC/QxjYNb3Su0L4gqPjrd38O6G79MGsiOV9dt6ajrEsdj5OMzHnMZ5uvwo9aiWmkL
WicNtseF13ANqn1mAMeqmQCfmM5hOQb+tKm16KE19qEb8XkD37iC3P+kCoat7mLjuueyfH8VCLoN
s/ojATfm2DZ9F1CmrT7pSQGczF0O5pMF9u1PuFFRbA8Gxc3GiKNZ0crW0ZyaTnYXOR54Dm06bJ+m
iPb2uQNnH2dWyQSheScfC/P/5WKZf6hy90VMxF4uYn93PPnLMfBG9ezw+M8GmzHO5EctM3Yo9bJ+
dMECC9Zt+uSBkrT6XJJ2Btad2V0czriSukUPEpGVS55J2UvHTAxY6EOqx3zVjXnex2BC7eY3ddck
3EouGvXtTYiWLDrl2hRFJtFNazPwsGI5n5nEil208FxmMb7g0yKmlq5Y45J9R6AqHuTkzK5lfC9p
lAH2Q7jneyN4Gd1u5CZwkIIUbVnoIrrJPeP+lxybZrLMyAsWKK9alETvUxQUSOWnvwLZnXuZd6yL
NLjPNLxOrvq+w3JuXgD0TsRJgQ3ILVp6+aIiFKSBo5WTwvh0mB12Xjkb6364n4H8iYDBLPMciFcZ
x2QHZoy9YwpID6o89EQs4zM7yKJXSG2mX2fL1RQrBfjj7UJcv8XlwxZJZ1Mx6vnLRB/xTtPz4x+U
vgERXp8OY1wdJP1q4Rwtx99aTVsVZAteVeq0NKlMx85sbz0BNpGPZisifoF0ieDvXwuLlY2dZQBu
lA2nZJM0UVSVGBug9lBRR64MRssLaig12QzfWuILJZw3pvq65iTW6kQDbiMP14EPGvobLC8quy5t
SBga68iGGSZhm3iJjO84OhJ7kmVFmOFkRPOKOJ2RU96Kqm/O1/0fvWFJyarqFv3iwPYGmZGdPNwA
tTWLRCgsO3wOmEk80Ve6baiRRo/i7z0edFvbczlBi4RmuoUZSuHDAuGia4Im8n61EuVEPegzeMbs
kYj3DTYhw7mUegtUi8vVLmTf7/4WOs+wnyYFOyjiJb16EBG4XS+m8GBVg1FtuAa1TQRJ7iPHejzi
/Uv4IAnF/4vH0FSIYuENWWGgy84VKP0PTAfzq8E+BBgsTR8jPV3/aGJtmRNj+ASeigTlZyVmxSnU
rjScScNaYlj6i6zqLDZ+3VQ4kMrkJuBQDxvk/cCDXTgL7qdCt1QVzUMxrZGe7BPNz/VJOJmpTUiQ
+eA6mOxj7riW72QbbFMqFR4GEZD/bdGyUKR3n5nF77N2UXo5NGnmR+awLN4HnBicAx9nRFzeh5zD
UTHE8gcBwgo38ReZECnwyrQl69icESqA3o1T+cb4Xy2yjXDe3btVOXc1IprxkUiGXW4AJIuiVZmd
DdYGwWODUlujCtzuXN0JU+kCA0zAl37A37lHz5GqZzc+s/YZoYGtNSrUhXmddYTpAMdDEO1rhvvQ
oH1218vZtmzly2RGfMqr0+NfgcyOsj3/DmL0YEPcVN2mXuzhDjwya7dRYpuv3vx1UlWs5DdUKKJJ
vvQHxaJi95K71WusJwjR+hGRHLK+08WV2+HFvXH4A0xrmPKIbp7shuiwuRnGGurhwWru7+H7NzJB
smwYyo3aSFflXx8hTzLumxRSktXl6WsiC8BLDfC9j0O/RvYsNsglQG1OD+kmo2qUfy4thsG6Skid
rgyyBvaXspQkFNvUO48V5VFN3nUk2stHVrnECRzQoTr9Lf4LeAheoWfNr5zZVCy06XH177thQslc
E84/4vicGHB++UdVU+Xkusux74qjwkU/Ln8UMYA2jqzppWxmcJ0/fv7EmbuO8ySWuoGNyc776XBt
5NUwAPHQ5m5lJa5i8YBpos8fZv5R/PJxeBpqMJEHuHhYtz/52LORh8jGhwECoV8MEY5DRxZK8vGj
PH9PqEL1ErRgqN0akCC3W2/YvQBO38EStRoQhbwfap1qrqxzkT2qCxemInY84NJsO+yrAyKj8svo
MXh5zTp1sd3I7HWIeUosUfnE4+jzNEALeegahVOlYsgtlEfK3OICL7ZMXl/e+bHdDWM1MedXelM2
EVO6aCAYGIcRbxSZCX667Xtm7n4HexUqVy88YvNVarP4CBNqgx0U49JEIvlqmFjhHtoM+7qGmQYJ
G5W7vviKF4m5201oSU65+reoycmKd7rejT2/jp2QBa3nQX7lHhCzimUx8InQqAl9WFTpYokFdrsR
7Mn6dA5ZFILi0swNBO3bpBxQsLuATGU1m3rqTKu6ATH8YJ20bpMLogr5ijXXiObkAoojhxGQtKmp
sfeBwJ01DGWPlaAjEb28GGkXq1cToJSDqDjV5CtWZKh3BfcBmtJ0wiv4/jtHhc/uOGeVbyhrUhef
0R658HjJYZybZEB1x9+oHkf1Q313b0CvMAGDEjKo7KTfX0VPZSk7gwkeqYWVUBfU8tYpBhOaczMH
kVub/1k11ywkubJLm2X413uEsWmkSLwevHGQ/zI3B3UC7cJC/HPHE+K4Wlv/IcLXgfbIJWLo+PNB
1p2CTKbxNV6qVDEoyAOu70gmi4GgqAqufOR2vkAmaWAm+2y3ZpHUdwqFIL+iMIAI7bdD/NKPMwnD
hBjMkcX2a/tx5GqBJqqYEZ3atfpP/zGWcPDSiHayrigSYygsUoeP6Ec+3VXHtlRFzzyY36tAh7lU
8iAulphMy5kgHHLKzRlBCc52PUGpqo/dfMwvupckv0C0zWAhvvJTU+DwFhCF3z3dzxg5a6PNSVAz
utcxU8Ach13k3D5F9Qd13LjgTqmHt1a9MWQjp8SX4HiZYUX3DoeJFbcaNSh3idUil69uGVSuBUMU
cmWww2N62hCZ3saTuB5oesUyyOWfyd/SefNrOcJHUHbEMr6Iml1O+KqlgAwlkPJnm3M1y3N2bpSW
hcej6w+N9t2YjQ+dtESX++L2XjtsycIYM1VRWxR+YRyp028n5m1pw6YEITbEfSKZ/1xnlR8qHNLr
RR5e3qCrBVw0DiXtSYZGk4oA9z/dy+KutmAcdzDXh9g9iDuL5exvg7LYKNy737Pc/lQ+Qze7gikZ
H39ygfAlHrN6y+1T/aPDQeko5t7DrBBfPUjCRzj0nCBBjN6GetUTUTkaXhCiLNlMK5hYfyLqGOHV
SZsuoahP6MZEehAnIakGyoHK7hwmorpbYJFtgsfVXCiv6POG5BnsRx8ZGj+Qp2GAqIXCoensHpRg
+S3FL9diAKt6A4izc4kbBFGR9OIBvr8QjOzNHOH2IvVHGHq5vExJPoi+jKb8Iu1LRPGRHGYzlVjx
xejVvumb+DgzqYttRCXHt/EaQo/fpucggj/6oaPjWjacKR3jtHjeSUYXGlC3PPp0HnGl51Xka+9v
KwiGiy++VnsvtmraMaG08sF/QIrbTQlsXZvdIdMMQgJi46bXoJBTI6z8cQUD5wLPnEQOkOnXlX6N
+U1OMxwB8VO9rAi5HpjnJ9Jqz09JGWo1IWu0TvC6iYbKT/Dd7aFXa+HSJj3QinwVPV3RhYc7NUuq
aau1BvOf8CfZmcovlJguoGlZHXgxQf9zZFpHZPvRIjtsFtLXtrft72OgbbKr0gAaxwVvoV/Mi3J0
jKiy3DJH5XOU43xSxAmBdW6i1WaEYRfq+IJ/QbDXnz1ogvns8+iWakaNk6ibHLzRBTn2X2ZI0PKn
LTLLKAIrtMBTE1E2iZORkhi9ymm16GkDv5Y5hUaRjzDIrnD0Nq7jixKvPyaNQBpJ6FCl4/u8Xbxu
E+WTy5ap/RKrRdB+c6fUf0bRSwV1BavhjTusB/n8wHRi6Ten/pgyxgjuDUpz118XhfU72d/drpDh
/xLG5BB78MkOiXp9ZleQKXQbLrs/0cQzD5NuBvF/c+FMnV1cxYgu9QB6V7P5H4uEoiFGbXP91j3W
64gmBAVKntJ3cyE4eAWNn8U29UNC/lXj8YqNi6wmjxDS2lWaWVX2eucgFwEmqLQNdpKAxvkYzahw
gJqqZ5C2HDpSs7MXaF9OGbZENkIMiFcoUrwdV8wmDewjSwnou5N1ik3dmbS7DITJi6ze6pkrfI5H
uCbh/AaX+Vzr0jEeNBuBzsi+LGJ7E/46fjuyRknAr0dan3xwTMGd9N3dtJSyzD5jxq+JILwRMiMM
xMRptmez11dg9K1WaiqJ5PWC6+mYe8zCdXDBXO1+iMMZnp60euHrqJlTYsnxo1mI/llnn4HjSOms
TNJIJBNpXwrKOrc97IThlKRrjjtJU3wxmxjqfmOBQAtxXo+vtkXRK/5pAVfCEkWR8NWLLP8PQYHu
wfLIKWeImxdI/tjy0snOTOq7D6sWih3yoToj6KhO1/P2wzgft4PMbP36vNohrWmR2+CBxzBg7mFv
OPVIbtk/zBbMHn3F1Y5ycMime+XkOthLBMONF0eMxqTVttf5yyPdAUGY/0JO19j+NdvKMuhxyzvF
JvLCbymzNdC3X7wc1KCusOzC4HaloYqgoEz6insDIAPrNN5Gm9patIGxEs+59+hvXuqbOXAUi/X7
u2d99i5R9/y9NELPpaaRsK85PQ4q2jy6p7Ac9/IWTZ4JLJCO4uL8A5K+2TdObs2XIO7uc0cEL+3q
4o1z9crzYd+eMwO/AlCOwFis+wXLJnHBoA3cf588TavN1xPzK+dTeHlJhaosr5oHCvtVEyzv2s90
zh2bpDevEt4vMD+00N/48YQOd6K+T+XHGH/4txS3Ck27RgVRJeRoUPiRUtAIDzinWLh0HHL6z0VU
Mi5lGCExSjdiNFT8VsQMjoyEBcwOr2niusraSn6mX0LLrZdXJE1JNYRFNuOW9426GHtkEB9XYc55
dmQG7ZV3+PJ0DLeiW3SwJwfwBJDPyMJ8aT7itf+tkXWMew0qV2vUyKWTKosbnUuzW/nP2gQSymwr
+irTX/aIBWdLxMdWaOWHWs0v53FnXvDmHRcnD+SWEsYq+5FncP6GJ8yYy/hiESf4VUCsFzztpZdE
Ip8EziDDcteFaJqCjApe7hRZ11jFNJijSnAApXd5FvLLRju1F4FNvX0coBHM+F6jxvX6bq6n+0Re
h9kQ8bji2ZuzEa39VapMdgFmy3BQAsi5NuHNe0kyiIrdZaW/uiYc4gjBGcSfwg4dicbbLveKhq45
3odePtXCwznWzd/tuYrvvL+LQcYXJwRM8OxQVPuR66dfeoQgxCHcAf7yhqLHpo5tE6hcPWBhmCHf
Ioo62b17IDwts2NGx9T+XaLLc9uga1niZ9WItL83rPqxGumTr8/VK0Hv1H0dMnbwO1PH9YiDdaVY
Vtz8HGqEkKVOTF0qZjaCwy7HRmX0PD0gnMXFF7a2FWBYreAb0c/puKZ6t2JYSXMSTEOzYc1k22vm
be46D4yMu8ypOv3pVXiKzI8xe0hSU2cTTa8qR36oAgFiSSjmbAu3euDzl0/yrzsEMPCyuRxaP2s6
WBtl5nM40zePXy6H7FJ1776nBTmYJiAiDh31B5EkRLNqF489I7tcYEOdGY8AWVoH60ClUXOypBRi
2oOQAOk6PuSu+ZiYF53PL6S5SXhwhIi2mLMgmcjP7ZuVg9sIQ9VcRbArewe4Oes/LHNjgcRmU6zC
bXuFq/+kPDGBNPa/9cTq/x4cstf+z68i8QaM5fI5vwJcGiIWJKUtDUJu9tK9C2avNfd4ro9vR7JM
/Zz7vRZUcllyx9VIt1zrJEAtCKW9LCGDE/+IexMAzr469iCIS3mZrBhRxaf1bCXK3OoDEzR0Ls9M
X+/XcM7vFzgJfSH3AdpNmdRbLUVXqCD3odCkGtakD3b35zB/CGtqG5v3pVONhB+XUp8qdLdnWGyt
dNq1JJIKx5OmydF0lcx7pYtzFbwiIyUj9ppcAOL6pVhGPxkoOkf4EyVVuaDQC6OqUwgcY5kPWxlb
pg8KjVsriW2qc2y+qWAIAkAgTWQwcyWI5TBvIj/Ss0a4kPFf1+n0RJ+YGIJuwcGYP3/8/VsLmmM+
fhrzd8GuKERYBFAICmqmJaZ5Nr1V++D823JPkuDe/zF6Y2yvdhUGD821k5qMnhK/DSPkasP3P/8Q
9YPeEvt2+1/JOiQ1YJAaJde0e82CAG7r6qnNHmB428utY4DDBWdp8ECsGSpVTf3iF2pJ0V5v/pbr
Q3GYwp4GUeFqUw8ezciTwHJMHmyvH9XqIycYLQr6WekwJnJzFtjlR66bwEM/r8CbJTCQjrqM/hiH
LxgQFO8tDqqtfs7MZS7s0YqTQOaElY8igle0FXMCCgi/DeriywOZM0Es7YDoWW5E/yP7LMW+dBhC
UMXbrIEXRNlNK3dJ0WH5CVci05zjSPXmvnu7ueOwju4rq2+l7RowkmC/JUiB/8WURenYSTtsJt9J
4UJiXzjV3B8msd508NPLt7VTp4TQierxw7PKNAm6f67ZQKbVTDCtBbQWdXjav/Q8RuZZ6vgYgGUO
4oJHVx8VzZm3FilWH4sicP+zi05bz5jwyuSs8kMNQE4XBOuSMawBNHPSrU94gAO+G22WH26V7f2M
ADCoO8uaAKU85TbX+egDyk05r6X8zWmGZRvzr22JhNECeqK00XD5GdvsqRPKFmKL6WN550Mpcz16
KldMElx2rcg0pvWoTf6qfkhB/zvlmTU0C8H/E6qzpaQ+MWc2eawsFXSOsoy604BZy4bnDNHa+tdU
UGBW4/roKbMMfy/TRIsy6lRuXM9b5NmFuVb/5rfLlzNKRb+jftTpDqtveLdzkpzrLekbOvTj5Ynh
Koo0hIREhEB6q5/XTQEoCGy5otDayLfs+8PE1lsnSDTfFlu2inPEeuv0YNz8vy8JGToutrTyaRuK
Ky9O+9sD6COWHKgfDu/vb+QwYVcIhZ2h9oalFKf8JluH2+hbVXrtED55R++tajb+on0Fp8RrJI6g
wSGGPhmWj8yrnM/EK1gyv7ICy1E/eCsJmDOxD962WxUNCUQ6LN9fhnb0o6ubAx4S33Vt2UlpYLUN
8g3ONkgag8h9kgDWkFdtEIMaH35NLhbeVg0NV9gBnMaiN3E7gq/DjjaiP8UkvcW7T9RlN+nXs5ez
EMDtk3O78wmsAaRP42+QN/y85AVN70oVk4qyQ1UJGpFzXUK7afdWyQoF0FSV1qmwIix7o1Wzd4n5
SUl0gNOSSo47HHgUf+LsdyC8pdROMnz1/CaE7UrUd9+penMLdWmSJqqgPbMYmCtyqYx108hiiNds
4nMkjGSs1dRkH6OC8GqI029MjB3zKvo8jOs6oiD6PoZ09qiBRqk2/GbuuLCpwruZLpcJKikqGVVO
rqD6EbmxjMqxhvRkuHTiC7TF0idXOjGb8gSVP5OakU7w1WLlIgIlLbmLj/qKm8QeZSRHmZvT0xbd
78SceDf9uYBw7kQreiklD1FxbSyUJGZbVEPDkwIu7HsFTH919CoVWYlg/whCee4btkligQQUysUw
TDvzXqPIrFqgYzVCmpb8iIOn1tI7YyzYMLTi38TwfMfKv62rVU2KCscIBTUl9jGcmT7QvHvCwar5
wg68TVIrTq9xxOxqkC1Fam5x+YGqsoe2eF9W5HeA2QF85YG2/11+clTI+8Baux3AMXR6/byt76xH
jmxo85kYHBMH+JDWHh4eyuClRsucC1tNhG5nNUn7EpzeMTBB0iKmE9MDIG6BE8cAelsnBt7nD4VU
VIR1Rk7jilGtOFRBDpGlVXvwyXvjjsQtL39MORGocnSbj8ks2XxXDIeMFyTQkd4XE7ri+8YBlcOW
+YtXlaJXhaaozj5RdcixSsXUarhN+BlQ6YAfIBM499AvPAsjXNg/nNymr7NrsdNGSIkAAUILy6pL
NDTaUD9ciSBmpSnWJ4u7X2kStITb0E1T5yQtK5S2KJR1G+Ax3N9gHNMK2+zkZAZ2yhv/2NnUnHTL
H8eBAnEREmK8B9/f0Mr8R+j+sZpnrKezYEEQmeZGBjU0vnYmRS22qHgk0axuaekpyGreSO+c+lQH
T+zWrbHCBCqDwEYSRbBKO8lY8mzuG96ZR3UhUNGWEQXbcaAwYYNDutf4k/q3g9JzAy9g9JVVzpCZ
g4J2PJ4ake2VwcZh5J2PYBW+a5MJKTf8OVR4LvIv4mhAOx0GA9Hvx+ueBtak4suSIpj8P4KMUY6J
iXNkRYrQMDPc1HE5+z7oKJJY0oV80+3zzZkPkfK4Msuu3aKyXfFVRlBgG7Lmf3W63YiMSVUUUH8f
icSSj/hmZvbfyz+bD7+KvmWzLLggdygElG9z2k3mBZqZNooKshOa4GfLD3b1pkd1X37/iJ7KTSID
dUMMJwx5HA0yJUgIQwhgzgF0Nuh6YkFvjZT9ympvvoOusbleL2Ft21uzZh03V6wvHoJxolsPbzOH
NHhxzlg/KEdNRxRIYiQb7f30P/Gm4E3UMASg6l1PUo5WBRLfg9E8YACvO95edvbg0z5P6aSMsQEz
INEhy8q9WX3Vxe1p5u/MoCo2qGtIK0HyLvxmKKXt63C3TDqxwfHsnCFQiRwD2A6T8bsrGFe7wC4t
f1u9emyQk+Ahs3xLCBukYUDxLGASKKVhbBRAy1lZMb0WxMGbZAJA26KPOB3eHVIqDHulPGxpzKO5
bVjJuzWkTKYSlfKYs3SayYHAq+fbg37bw++D3NS1xdXmH7mK6PwV+GYdXVJ3fOkx4TX/4EDp96Jc
AvK1f7cs9piiYRG56YrymFViBiQWyk29a6EatQabon3y55i8W7Fcd06CA3GT4P00Fsd3tpmPYrFf
W3Ff5E5rZkUzLjiomiHxKBKMbM4zgIpr/4J6NnSQRZpIz+zLv+ouRKHQ6VVQlaciMVEDMRV8HFc6
1QThNDb1Vj1uphvB3/LZ5DUjpZchMD10OxUZw3oEp45R66hqXJbUYl3byQYKlz1AdWPN5L43hOQA
VAIDqQ1uTRWT3QIvxPazauU2y6ysl8/WAS79N4FUSvyUmndZR9LEalIO2CcwZykGvnuVzjuV7opD
5ByE3x25ArrZcai32SR/D1QHXOIzqW7byLifZTj++O4Gs/13cZyBZomo2F6Vo27AuWWxEByR/4kj
QJGE6PYHxL1+3L8ZY5Cz6p6SRG0HZ2gW3Nyn/69zKS8+FR9adzrLnaHcpOTR84aUvslvtB6tl7ph
FbnK4eVAff5BxlkXRP2Z2esycoskiN5/yj5bvIZKTDBWtv+wFZGWHG/Xi4LZbWvWOfxeULcGGEnC
RBCSLkgWuKriaPMWRXqYbePTeFbuUdtV3BITzjTG6OkZfCv5CxWiqhZxfj31Az49Pp6CcydnEymo
P+lCeUXSHhwTgcuF/N8PcAdk2J4ZcjBnsE4YM+nCMvLL9LgsIT9/JWHGs+yihVbZkyYUPUBMjnAI
wy68nYOwAzPa9HehnzI5Oq/NS84+1G3N/a0/fxpmrwx5uB4pDj1z9VO7u7q3eqohnguNYQOrHDl0
wA8pEem6OTKjkSnPz8dF8x0wt9pW6+ntCWrEJR96ZLRLYX/fMQaM2TptGkwSM8bCgRBoGvu3eVvf
Yekco2G8K5DuS4TIATjO0PnbVfCWVL6SZ/BZ4mkLPUA1QlAsnpsLxzKIb6RdWslmWdoRu6jw6xZM
0JjAGHD5XgakinlOsk0k6Tt21rKxKqjR+9/iL64t+Lb4retLZ7mky0VdW1DxL2IhfXGo33p2eBzX
xphCP8wMZQRxKZtjw10De1qtS08NaMG9m5r86hsWG+2LLU6srMll82G+Jjx1TFdDC/hBnKNA650E
gaVcOC+8fHLc73lGdKFBYIzDvC8N2aM9w3MJT7dUM3sx8uBMf967N5U48nV30kykbHdv9ofxdSQL
20TlUL8b12qOSCCfMMS9Z+YNht6Ai/KUkrbqm9xaatj4Nq8vIRoRlHeYMwqK4vcMsSmFGfIJOFfy
Pwwn+iRy1ci0NZ5JPWfK3D2fIjdONdWnhVT+YvnFjn9JeaVL6a0HQVbOv3W+x/haSFNz3BHVbrtm
nQokuMYROaUmVdTFmIsoQvQVPT0rWuPYL7Y2FZO5m0LR78Le9lIlcYL67Y9x1CLxKk8pUADbk7mw
TwztRxhciSpnSCweSv6SzDUZzkNElOjBljogWltcxl+Vm/L/wD4bosfvKKw1FmRlUa+jZbkWFt5E
qt2Wm/SBLoq+9Z5Zm5dsGZ+FGNQU8DH2SvfVdwnHLo/RlMNcGdCmXctwxfaeZlyLQIZa7glsGctQ
fhlEnL2UvUErQQ9fKSBdCO74+luNz57nSbVuk7ybEKJCsKztaXxxqRzcfkem97ISkQDvCvBuEr+s
Ylb7dgAelAhSthDTm+R/EGAfx5k27+vDOk5L1TXM1VOx4WhY06iK8Wc+DyV0GubVT/Ng05eAPYzC
y8LqNh1r+cqqBLkFPQ93fer7+l94yyVwRx6Zo1VQj3PIpfEtvJ7Mnv6VsLmWNlJhw9YYhmisNJ1S
ME2ayIWXSPuF9wG2ks584C6X3keR9JKlDv8WJ4ig1yUd5TjzlKUez/zDpLpOt8pLgDcIl9kPzGMs
ZaW4OM2aJndOUt2fQPSqiifcuYhv7mN3Q6ywj9GJmr109DfJuMw6WyZdVqZ9ORrwHPkDv0519JL4
Jef3oPL2Kzf5lnw/aL70F9rVUQjqCwZmDaFweaqLNNGpbHT2LUkR89vOAHz7fgE6J+/KPF7dHF7l
FBR6NW0Dm6ieBV/2HYFJ9m+pC/SBSYeYxAMmNJdov6MZcHItKfP4QLBsxp6Om3t6iUba15zazYYM
rYpa8L10UnW3EyUcoiQONQcAV4kkWg9AFc04ubzlqWVTCqnbY4KKZOfmHdSKW0K4FS1h+b+HWT0f
0TgkD6rbnw7Y84+d3pPHIUojDr0XHiyyXz3qPTlzWCPke772JC82SlzGkVc11gOKJLCDnD2lADVD
7a6St+DgFJyPEFoWlrAJjEsBX+VDKanffb2bo5NVeuVogGblaOOtcpeneWt/iBtMJ/8Tl5omkf7c
uvCH75Epn9y232rHpqF3sQ0iIhIT0fWz6zQhfQsKPfaAdU49e3iuw32MnHNDrg+odJA0b5m6kjZh
l4QH/XwnZdpwJBzy713ay+VEZutsWDRLzDGrnyK+RXKo5MyAQrS8fUJNenroiDxY0WE2gJNiw67O
WmYW6J9cs+jzXz8AN1RX9zkzTfRQ1/g1hYvWgrdXGn8qujX6KHeUGblZj3UR+QmAV1lqEE9kKmFT
wLmedXAppcwetITLsqPdYBjHrt3jnY3r1bhccf7agLv+8hEpzV9zjNcstJTW8grydjDvJ3nm+3LA
XYJzq08LjR1cLDD1CgIXXOpbMpPvUQBXPu1lB8Sad6/sc+W5X8kadBcIJmdx25pPktgoukGSGPf0
3imAG2LZ2WEMvNqYCbAqxXyMQj0ttF3sWQp2ULXV1JQGlY0XGdVFHHjXhYHVWrKm7tI8dW9TQmMr
4D9feptF38MjwV/93Vh/iY70+j4VoNbaiS6ljbpqZNgJeSeAUNWYW4pMkH6Xq6N0QwJzNz5pvPlD
sV+uhh2ah1XK9t7GjOMma5VzA1uMwm3jADg32FCvYh4ducppnsPf4ldNmKXZOqKABhhc2SHqjRs1
yjhUQ02YJ4fGZX3uEjnx2zl7ORCcXKg7jjUOXGL3AxcXptMGoLGXOlC9eZBdQ/MxIkLcXc962S3v
XlJz6vO/o+vOuMuADfrdZTdKetLj1ZpeiFA3KWmvC0XJmn0Bhxl4PRFhMZOT0XJ9ChbwOsRGJ16t
Uciuck92fKRdAQdAC0jNUn/BFSnxU3m3Qsg/3VJ2MN4TgZWg8mHGqKFDZUDswCgvF+VWD2WIfYXN
ZZ9eAHYYZaPZCMM35dDPWcaDp3TyzZl0P+c7StdaSOO3DD+NiD7VQX0Sx6V4QOBqtqivps6oTtLA
WeMD4hZ6ksesvrcQTUMHj+thIT/0jvVDi5rOWeip9EEg0spoMDb9HQDbYkO4WFBd9O/AABKTDSgb
6dORxcw7K9KvaaRFuyv77c9wyFemnWCF7ry9nBX2iVPpQNE4KsK9Wq4M8csFgbmRup85EOOurmRs
iKCzCNj4IS+1bUw751AKnGr4YZebRvlOT44p5i0Rle4+Cg63bX8+lP2K6/uLvPgpQykv/rLHODxt
844UaQIUQOzMYItOo/O1GcYin75YJ0bKmtTuhKWnvI+U625zg8t6ZS9s2AfoudUU7pnLTiryYTyS
aCZHKUmv4C42oANQMt2QRe8TtXERqmsyarv5v78Aj7hYihLiqUoqvQkcbVOOPCi1KBIg7WFJhJ55
HW9lEKBsx08F2bfJtNKKraNeriiAYHkGLktVAIQb95MJNW3SFrX+e4JfiZCv95IZUSpmUDq2rUZL
CdbI2L7DJt1muRNfbt3bwI6jDlrx8PIDC6QHunOkwF+6IWnac7NzhtIFYqw2s0w+4HL7tXRnQL+y
39lyb5xKCR47P879GMuOI6cSjOryv/zhFa1ci9J87eIWWzT428uAchkO8BsFnSzzc7JrkoaZ5MmI
dGV0qRDCm8lQkXn2JevlbsXTUvAQX1Gtn3+tiUekGyGlCIzw2H2yu9P3yJMpQSGAXgOQ/ij20XTH
CfcyQYKLpKA5l0W+GspDh1cUlRn7/002I33EtiNuWZfHJBODChWqeHExfhMts8Mxw4GKJV+cU+KQ
FnNTJCEja6wY/y/juk9c6DsYPAdWgCIkv0f16JUhVynI+FqfwZCpKapl78i1zTB9/cvb2CkVQDi8
51nEvMLO9xKVE0wwHuVdC+ncWfPjRNls5sk6RnN9xxmm8V+DjNG/UWb/nypD2RRQBNBjOkVJlo2t
TN56laA04tZ/s3In35DqzgM8jZvktEbH7koj5yWRyUek5W8WTAOSHpAgHshZnKCu8+TDpNBtRtUM
uSIAsA2f0N9yYhEI7r+IOqlUxXnxsJc1BInkhiG03elg51Gl1o6+v1/BTSOdfOVl9LnE31fzJNcA
EdntfO+Mn+fjnz3Vpu/GpT8STWiQvjVejKdonVp2IiouFrmObhGAN9tgwoz0AF58kSy1qu/4c12X
AxeAY1c8m3MyxRLva4ndbmH+jXM2NLcQRBfdi7bZxdMKrRmIJMReJ/uxeKl6BKNKoPJWe6oJADRH
GzSqbGcWoGIr/GUp7vudZSJSNbuL4FOAxbwRdAWPedzR8cN0Cbh4x0hnTshHctjL88kfmp6a0Kfg
q7UDtdhbGc2bcs6L8J2BhNvzz1lHSglHatu1q9Vn3zePsvvjMbtxR0bHE1sF+umi65LKNzcXUTSq
Y+FyBrO61GmV0sWgK0Ous3OZMH4vKWQdqrJwEBtq+Kz8/XpxN2Ly+yTlWuJxGdetp4JQJKv5Aqah
vG2F+evCSRguGgUXE/xOqprNBo8TDP2lHaFVQa4DZ8K5IOvIsaPYfaWDSjrp381kTLaZJDLM43IH
NVjRa6ET6YKNxdC5j2ZL4E6gJnvjleBDKpURvZhV/LDQoJZQR4zB1ty0ETQMXsiS8b1NJgrwhgBa
rv5+0fXLHpE5pTN67cBXKBzqiT5eMrHtq/VMYl4TzVsdIQDc8wZQ+tvXAvAbkw8DqGG2iC6WivtI
Mq5iP4iFFRcd2VpnD2u7SjMP8riJqxFJAT6859yOroq9P1tgPRBVQF6fEfeHyy4Q3/sp3I26dtfG
oQsYTfcTRHfkUInlfyib0BMVP+GFhMBPGB9MdztN4IMcrGy4YJGwsStlNevGvEbVXFzCFUGftDjw
7A3QsZ1f5uA5FQeddmn9Xqqxy8xqjuB+ptcvrzODzj0J/3lYKtIK0vcZT74pjLTo1dufL9D7ahJ3
+01gu3iqLYLg+BQdm7uqLzglpM4Ae84FCTv/RszHdZ5fqC39ENo1SSKvWQYwzoOSeQ2itL9h4dCG
YMcetFOWlbFLq60X7s7ljcsoUXKBn0zoW9wnJGcnHmqwv0tWVZt4yqdbPgd7qIkaCjSsLuN5xe82
U38ijlEDCSXo2voxcwvSe5ciEgszWY1SXW9tGfKLTY0pqJOh9c4xgNogkb86mnGdzxzimoxxdRaj
Mp1lD0eE+jtalx5gnte/MpKP9FVbA/NQ00IillCSW3HW5HpswBelH3unOZIJK0vvnKQ3xl0LjERG
u5UQmwa2jHEKUiN5CoJ+w1mwW8eCm//qlTcqF+hCD4MWpDNQ6yFoV5XWgQy6F7/SLUQxwI+RyI7x
OOnnC01n5fdCcOVcfB3q6iGemh60ryAj9sXALGMqeCF7/osNj6a83hYI2t6H6xnahe7BdZoddLFn
rO7FR2QgcYoBY4cr/GFVkVbirO4ppqGnMhe6ItQ/DnsMj5mmA5+s/d5ojvhIgABi+qtFt6XbNmKH
9ejrm2HvJtwdLncbFOlKjmesep4YIcKou3Pnmt4XtAYYncjOoEvipMHnIjaqtQonBuf8e+cxlG9h
ulhUry3dWXTb/M/qIZx3M9MsxMDa9LNA8RiyNsK7Xwt/3E6SW+ujd/c8ICNsWZNk7/UMq6xxLUUY
Tw9oNDXhWaQH3XtMz2Ogzd4uxtib7ViKM4W/MqZiPsl2AhjIdOQue1nkOnWoIscka+Cjn2q5fEOo
93Jz1LizNNtsmDitqLFksr+uxFpJKc9GBxbIMDH4fcp9RCbom/RzWZiWsm4+Ui5xL/Aw9elUTyhH
N5IkF3DdWjJg3uMyMJcZx4BhCyzRnxoip1ruFrI+iFCPyAJ3cR1Rs/MArWHzgZlDY7MrEZymIkCR
D40zn9LqBPeVDiYYv++9fPoEwd/e5wyf53tecO0oeYj8qfJYr5tUfJWntbUOzUondjMTPNGWW/lU
CqRY+dza1hsp9Lrv33nP6DNxaYniHxSp9g2chAdqfyvlRX3NdqgEoDQ+b2g4AyoecZd2PVJq4Iqs
MN+lRMc4D/So9n/9LoimLWgNC7D8DGiL9lT+lCFXIb8wkP7PE/zl0gPP8ByFDXqr0dC2Go6J0s9Q
0+CJoKQXlQJ9LxKdv75Mh3kmxnzE+/WFObD4D87c+jF4j0AtlhkgoNvm8sEFsQt0kzMiURtBPs6m
mm3atwa6vmp+wgdOEkaaxYm3Jv9t8kjNVkEayKbN/nsPANqLn+FNK5SWj29soGvo7O6EmyGTi7RG
j0u08C2fcYOHErpj1cVmFvUtMUXefM9+ymA0zVwtOaACkw017+Ii/R+vViNCZVo54Y9DUCGDsq15
9q+bdfM5OfxXniYhse0AXx3fVDTu0IfiXYZi6zh8TsLuNbZlttaAqCBQJVnEglYC5Tkqd8NHb+tB
p6KXNQkjgUGlIoEMG+xxIeALbwaQ1SA7LT60wkNjRNctQQISzzTDox6kny1ags12VaPwRcvLgqex
Gfu1FW4ypcTgFKk1XwXucEyNLckGItNSyamvNYnoJ9e0Vy3xJfPb0CXoUUfE1UISU3v2pDgMgmG0
tQDdIxZHNRKIuxPqpj+ZQv6EMp5YO870xmTrY97n7rWF9JZfz733EdI7cUfPnVa/aihP6ErM8MkZ
7y2/Wk1eZEsLgJ0pghtGrtglsR5QHhuflaosNzCjBFO6/FUX1l2RU8xoUZFn9bumB9QHX7z3LVXT
l/NMzYa/wmzkAGnxKaRM1AoZlc/R3AkGOhPQs3uGEpadLnxDDNpc4WCTt/6EkRo6YoTJfHgm2pjr
aDVfyieEg2RYe+0jDxZquOo+JkGzM60HqtK0rwJ7yibTXFHtqcEgWkAKhDPl+uKQXf2mepvaKX7U
ZAREW6ApmaylrXGsggcWJztkaKgdPdILoQarsp/XZ9eyYUG+ry56aOj4w7pqxyCdDFR3eNovZ5XH
Ld5THMRW3ks0fosyr35XOP1iQqcZp8yWbLHymdHKoWuwwq6R2cEAkHP9qTLG6hLbv27Hkc4gp4L4
1STPcJh5I2bJzhZCgBP/XRRv3Z9A+L0azEKtIRDzUYO5Fi4du5M1F0UvfMfUHiPUKPtM11cC257m
Pw7sFw91agiXYHQs/YgZbUCh4nwzW3MmqvrA7tPIok3fl57YrMFSGjOHJCAU5Cm5pPa142jE75pi
q2/cb9vkkH2BoFse4ElAXZJkOMJbgmrbMbGcWUL2jWByAS/ntWKvlk6ECtFi3+kU1QybZ/+xbh9e
ckEQxonWD23Ze5gDV8qIMonvF5vYyhdqzAZReNb21Q3NoQ9RzJ1vElwY5SHYm2PXwIJX4xKl4whD
5u2orb5V6qiGouCOPkD1NfIcMQO0d4g+vhFakUykX/jdpc27nxY8SOxaZl7tttTmiJR1zS8m7bht
TFHfSt1gHA3oYRfCgJgiyG9wBraFhQ37lbWja8y934Qc3DAs4ugHt/lkL6PEgHlHb685W+iLvJd1
ZxB1aU1T8OkM1IRZ4dDiLls/mNWarzZIIZ5PTlEGrib7KbfiN839TrschB/xwFB257+BFvJwSb90
yvfR675iqcVRswYAIn3EAXUhaJs7uC16MzWisgLqYM6+YC+liYn1vkfQY9YtTUbYpdCGfbFTL6Vp
0yamG+SE8rCUKMmPSIPgKurq8mUjGSPPPy0x1L5YBxWCJyjY76QK3a2C4hRoya/yT1axiJNdTvcR
2fU7zIeiez2My4I5DoyiY8kZ8wTKzaREKm84SwroQkhef6IREctSiT1b+Wtqy7lNQBNqYieqIOy6
lOgQiO320Iij8PTS7jBI0eaBuyW27xNvLBfKlMzusp+TpwQSmxsKr0MNjaZVDJO0sf4LL8rHAuS8
2bGvGudSzrCM3XE9sPw3GcFYlnTTMEoOGso4juuEhDTFL7acQg6pX0V7a6q0Gh4+Q8MC4zkuzdeE
hERPft2TYh3ClUlM4eFT+DJ5xfgsHha0qjESb+ZXok7ZlcS6Rka3bcZPqkQB+LS1fqOdvfPqrW8w
VcWgQapxOBMrZKZdQUz/BdqStJ95o9uV0ku0zAfaCuedwXxU3Oa9QjMG2tWK2340vGYKb/SvUHSV
NH2gjl/QtrYsrS0oSsOBi9wZNIvAF+DqHP5RR5w9Kfc3zE5e8B2Pg6rbQRD5lO5LtuX/SYwKSGvU
XudeWhRJMBAWeG2Ebq8GqK0tSU65aC7e3ttlq5EzneM4DcfyAPj8dOzP9/yIWahua1NT9vuG5cKH
NZUjBAuBtz/tYWrieB17MaBAUE/hIgENkkktbcTNwNixYAWENTemwiWyLMtqu7onnmJDZ2LFS+7h
jezdO+lsHElJMCh/z3Sbvvx0VXPM8oUnjzsNszrq3FpSGrXFWuV5bw+6GFOls8ZtQyMcJfS2dVgV
VyRktjn3M7vIQ19SU9ZpHRVOy5s5mHMpgB5vzcaHHxcPPTQDhnJ7CiAPvNwmjAkzXhmLhLvSkr5g
OMtyRnF1PGB4zLPtYH/9M5eZSSgcMIyUeur++AXpq8Q0jy4wXM5lB5QqnyZr86VofTuthpqGP1iH
PusNeXSKRwj96/wCQgPywsUOQe5JWo72BZVtVpYhGQvWbu4Kz4bKMdmGGeCKLJhUrvgQMsqcUi3M
ev1Dnr0HQ1pED9fw8DZTvu8uQueWxOzuma5zQyOX9PKMDmNwW+KAJITbazwsmUIw0ydA64hFS55g
tU8U5EPLuYHpadNUAsytct5apyI3bKx17hKKlta2gBkqUcfNgwIAwRluA+h2wP4KrjRwQVCVmMQR
KHGl/8jevQhf43cKBR2I3m/i6PZrtQhG6UAgF8l8vI2QzpmBlOznhmlq4v4Q7RtekCJXcMZq837j
ejSys1pmp6hEd1nAshJA6qE3OsEf03dFDCm4gptORHh9YB7hNHlTzkGs10c0OxTcX7ZSQLGqij4y
3VN0qEwlik59ge6gNUFOFW+ZgJ90ZeNk/GEWe7uPbpGOY2nyBGcDgWXAoJWPnAKmbfeOeeKMwEOG
wzbqUU37Y/x4o1Lp6sTIjfeyiC6mWWRm3XAm15HWBySbuxwJD8c6Cmu1WELcXXXmxiuF2lzwe12I
bzTrJCrTsc5CUwhBIxjH79CqDzG5qZbLMz/W9KCOQ0eNlOOvCLG/5zgGZDBOMS+6RGHGrktPRGBH
zBls0VTs0+Ew0+64ZNHkJBvCuXppcAlaRxRxprVvkIkI53RoW0QqXXoDrf/WkGVTfndn8GGBBhWI
mVWeVwGxQlG5PW3RR0iaFfcQA9YVMiq/6Wq6l+9OkGyAqU67Ann3hkaKu4qvNxBMelO7DL3Cb57c
nzs6ru4ekunhVm4EAKgT7lgasAcujG/9PgcXm6RoduhqhRv8UIpL/erwUQMJajLwL8TQyFuT+d1W
MG3TVh6YIeSyCGQI5vNRNit1C46uMnImUgJW4bSG/wYdRvcZSsJU1UDxE8ACMEMiP0bcX6wGWMfQ
A7dUnWETadnCc6YJmjRoPG9x2+TW1VUuIrajHLAsmTIMtRZGFtBsNqtp/lFsFf9y50H3t67QVuSB
4rHpAFVtlVyeobVznz6zBETzx49OLVpY/zo9wwpumwyxNBSHGoanawNbwvVBSuxSBATcAWIhDdoG
ToB0+DvNfqJp5TOinK2BMr6WfuuduYCXn0XuaCwm5FI2fOTnB6zk1QL59722pslSlcrh/wildU0D
2ZcIjYMCfOPiK3HyQozcX9FvVEEy9+3RmhnYcJg2rS+CQU0Im3XSEqGH65cmZL/Hl8njA7fJ/IG2
JYBIgrKHNegiWAXtsj+QfmPd2jGDZ9NgD66+0h0NLuF+DPeqEs1zwDN5jxzsIAQDnbfaB+LrG/rg
WtNk2a+1OuSu48I//Yh3F7jTg5FMAr9jox5QkHAG8Ive3lf0B4qxYb3DZLZLykz+obKZXwOiL/kB
hs1Sj2IF1Q6O4FCr23UKbc9C6uG8RDcyRkJKwf7rET/UX0B69FMU1OC0UcjmdARMcMA2YEvz2nYu
XCz1vM+mXBlGmIU+5LuAo8clGKvfmYjeFlHxcfBrG9EpEarmYJ5UaUts1AFUGAiG6Okdg4skocSh
5A8jLv0dQavC46mL7aa4CZIcjpdlVnE5mAPF9NeV2OuvwNWoSc3B7JQ0UuZyZ5sUhhidco0woNPs
K2RKRRsiAAAoorGwyuCc8pYXPIYQZsrHjr2t25Wo3/m1gODFYDTmQhaOj7rTzLITtFch2cy3pXA8
ESwrEBYqZK5Ml+4V2TIMezPlDvi2Ru/uDWJEXkgQ9XePSq8irDZuG9s0wTXny+9BgMs65uuuRk4b
eiB1wgHk1aZ4mlACJ8TR4z81zjVjTdz6YUgCoZxwywCelWMnobJv3HOOv7bVO91GV91gqC9eINiQ
7H1WDNWPcPmiFVY/gt9c6IsCd3SI4v2SJ6fAc0cJ7awmY0E4aGJZ2sRGL9jCj7yAfyq1PvfbFU5w
n2+S1oRvMU747PTPbF0JvTMNInBccZT4wD6Dbkgkms9NX/CDvJS7nPdt7fkJ2zy8qFsTXrbjkUvU
cSWRW6j9wrJtAc4S4gCaRft4N1cJjZ1+603lWHdTE5qiCo3T5ynlooRgtLfEI15p5O/wCMQUFt9X
MVriQG7+g/v3qobP4BQjISbdSXyRVIBlgDov51XkHBpxF07MLN6hiZ49f30EpTjRB+KZzvKdVZ2h
4pSkp70/PiLZOoOCqDMwNdGhMCxOTawxKyJYEHNFglZb4qhPrfCseDFyzxFtDuUJT0pMFREvu1Lr
ZkRfIbKg3oTwhN1/n/JcLK87DjW2iK++VIDaumIbJbF2tMN2CKfTZ2xqLx44zQXb5OGrs7FIRb9c
/lVgF/y3RQiR9dtZxiHloP6UVdMwEIqLBB5NJQouWTud+Rwb5GJeMH8QK8c3rdya4Vn05hVE5/Y/
JUCsisNj2FLiLJxNEN8BT1hiy7pwOglSMPOZ5K7FgtF14zdhThmeYV3UD6E91LdCcTr8692RI1tN
XE13XoG3VQvU59q9aTOXdo71x9//9Tt17VAd7M29zIg4YCApWSY7haryOAgcXnLQ8YxrVPm3yvwu
jXZU9HBaD5CK4o7r7f1BgddwpGtN7OHTC+np4Xb34V+4BwBp7P23lmelcEaLlJmoQElHWzXVRC2P
92Eb2tb7a45clNe4e2331pCCR4TMlS/YLvCMlyHSBnVYT8DeF5vSnsRAIbvtERT4Cp16xCnrfZtO
j3XCsy0zjlzJrXtHAIyMwIrunqK4xpMdQ4tTOj2t6kRAut+ZTJox0JKQAN7NxID6rnmZO7Dc7Ot9
RQ4EKbjCl3TpBGzYdQG/4B0McnJjljinmXPRXd1vxzwRd/Y/ENOQl9gerjB1BkL/6r+yy/iWqHd3
TthuGpXRadOuNF8YGchYnaA/pN49E1cpej1Ruj3KBbxioMtUJdJfXmuKpgDw0dZEv79WQOruVg1r
F9ALKtrXwWrc79+5bVqHD5pgNAiaBORIUbzMyFhbi3mFSFwBt+PGi/65EBHoduNMLEVW65GOKJuA
+rGB37QBJJw0Ojf3G8Jv2Hby8T+B7G8hMiMl9wJKlG6wgZTVUs8+bLp8AhjymOxzrAB/znSlS/Ys
mAUx+jEUCtQLgOhWOb1RowB/xGVOXCXw7KoAbBu+l0XSoGe0OYLxG5M4BsGWHcQnRwm3e8Vhz67g
MotfsZtLuoAz6W2agLqLhvQ/HXSQIUEHLugUj2k9i87REcmpIG7V5JReTWm5IsPRgcyPj+vWSgR7
ZUy6djzn3N7h+11ZCMgXG1wxezRCfc30Sgpe3A6Hx5vX6vf0u/4cra3HbBpt0tlIEXiPntPJO87L
YN8lYNtdlJoQBdHIlQ4F/fk3lS5ljV5w8jaW5+Tt7OMht/sLFuq+5506VmkLbj6oe+tKdSro47UW
nhP2pP8FzRB/j2CXI41NWk/EbXOA8b/033N1bL1b5YPGXA6Oc5ST/y0ORDzOdpQQiBfK1/hb1cI6
GNuNTopuTBpNmc49vTNCIMkrBUu9N9+ClM3R+Ys/GFNNnGtz/KqltSj5LkMICvnE7BIt+bImV5oa
SPE6WwHvpsjaNCj/6k4O7hvkywE2zd1uRstzezeNZIgbJdkFXpS64clZ2cGjIrz6sjH/+gxXyYX0
fDzq1q2k9XuJBFaFvyyuwgLYD+lO4bCn9CBKbnAMAqYit/S6DHdai0eHQmiIkImdCNlii1L/Ji4L
IJq1njeV0ZrVYje+AN8cAJPrJ0q6wLjaJPKQOOGVlD4RJGyHXv0Y3fxml2JtNsWM/OHrTCjRcqVZ
pg/PCv9Ke9poHX0w49Rvdrmcgg0lZ5LYzgTj/Y/a9f2kfUhgyAUanECpyWtWfNbJpXcaLBDrwe6y
XlBRhoh2yj8Mzfckkj6CmfFq12lXLwBQ8FWKFcRTZb7PvHm039M4lbZTNazlei77FNq4xUMuzPhu
BStWrv0IAwZg86ZVT3uApSmA0QxmL2Uk+0XL+XTfXZ8susBRpKzfvSE0c5A9S9WCSWKltMbnxz7k
OBi0c1ciWNdA3+czWenTwIt/PdPyxIFoGEQIhULxLkcWdWvRdNbQgRX0U3JKcaXItSHl2fi8/7DY
iuprZ4BdN5pWB17Ly53pY9u7Y6O1MgkDURCAk0h/Qm2tDb6k7tT4ci/D1FzwD0E621TlFQB+LmfB
aGAapBR4a+bmieRS3d3pMtkbk8hN6ASGbTmhflgAMKxOTZJAprHZsce9kDCXwdFW7bepUX6IlLBa
V5lGXqxQE48zwqEJ/1hwFKJdVZtICMI226U0SDDovQQZHFygSmEkgPOY0JEn2BZovkKBJdQdFsel
2QLie/7fXRFr3STQ2u5tdXVKDlBgzzvtEZye+CEoJzjHBjU0NeTLAaUyMOUsdTM6iBmSOSxpqulG
8uuEGGaHX/dHVUs0qDNgA86sfSIX1YffGaqGlNb7bQBuUbEpQuI9xxXbsu1edEv7C7zTK4qkTwqE
QAAyd7oCWApQ8gw2e56oVZa2D2RnMlNz4X8r/6MQBOc05ux5cCKfX+1M5SJFVETJIJXOu7y1x1hs
eY3bb4gU/YYix2cPRSOF47d+V3jSQV7cNAQn3Y48eU+F52xGMWr+9ydN2gS6laXmtC1HIibwByKy
F4Rn1MOExIhqgwFGkyoeuTU6VopzV+93WVDa2s2EcS71wRdi9pDTfxkJAZjmWWnnXl8wB6jo5HGe
qUuG0ElLT3be+Q92fy0vH0zHNq1seHfm3xAF5OKXnC4Q4B4tSVtBSVWBVS7nLW+qUQ2Q6Jwogfha
Lno4eH8OC6YM1JvF3IDmZn3BCegBtpfWAqhVdxsjtTtHi6d6uClQY01Jh9orYBi235kob8r2JbNG
gtHDdRSXXba5QK57r9zXEmepe/ozjG+GpIOwNkXuxmACyxPCxCpiyaYcA+yZ6N55PyXUsJV9CTWd
PeNb8DfYbtSqAjTxtWLIZZD5kdjLcGuXWVkOCj2wRvHwNY8vpfGHFyj9hyYjysbiPuAP6HQwnpDm
tX6CbylIziV/ihIXVIJOfDMuVKi+bkjW5X9GMCbF8DWkbobcgwaa2/FQIWZKhDipIPOa4vK1EdNO
mTf7SP6FRfiJbMMMwoJ0xN/sNVWgtfZSVQiBReQJAKVgj4r0y+gehdIdE6wZGwtJNNRDutG4fcmX
uJ8yyT+yQpBuAfjAciWLr4nXl3HMV0oddcoebWhoQ3EjyzRBgKoPf3WJsZFYnFY1IrNCPbVfiYcy
yMKPTZCnMo1NT49cOZFFASPp1iGdTTvXZdFXzJQI9m76qdBlq4HdUHyzMqEdDA+f3SpIOHRWcpiW
fK+jjCQf+hPe75hMUvX9zdLDwG3pM4Q2EX8VIrk4TUpsRTVt0v3ik8Mzv19LzC32HRGKRSAk5+TI
6kArGR148CgRj+KjRzCsZ8ZG8cqFjiBMjaQccF0X9L8l2J5EecLQXHKMpOQDjwo7FeMnkGkjw2lR
QD7ZxmFbOgX/YckoPDtbCLKw0M0qEE0LMKn7tQyoqLR4+21p+vboMDZGJiDNo0q+OhOoyv8Jmz8I
6ITIzPDahkVI3HIEVkb6biQQFZLu2JRcNUbjaWta8+XBH9KMAx7W2CN3hJwuHVSyBKRg6lKoB3JY
jeEQH4ZXZsOzPrJOJXwnAyHfQiHwu2c19PEh/ZnZSMD2x67hX/XwnZO0bzHDj5dhkaiMuNpHOtKo
K4dXYymEDNDOs8J3MHdQ5temm89GHBRUFKs6e7vWN24VPWdMauEWRCkafG5U7rmWSodkE5Q/8cD+
TTJ0MnzEw04aHWCWi9V8Av64OPGyAX45MkgvT/dcZxiwm4WC3U2L961CmzYZqWpNt4Mn9Po9tVGC
dcfMh/zjA6XWzP2dAe8eA5U3Y/h41ixXFcgY23EiBLivzJVonMYRf2oygtoIKoSTsWAmt/xVgncy
uX+RsQoHW3GxffYfC76oiOhdxSziTmaZTdgOHY5L+k6fcQSWCSR8NIiTq1jyy9uPrjV1HVujjUa0
RMzZvTgrmANhDrG3sfm0aE3QxLcYVuRcHwDI5FXfnSJ/+JqgS0xqDGd/5cqE3rv1rmSsIOTkRn0w
O0OtAkqqrueOBiOOsoRokqRCZU09NG3yP012tqPLNB3eEEI5b6LkUC99fbl+XjbfQqPFKM1SNOXL
lIM9EUg0uLz33YvXNDLoIAwEgmccaDwXqqorgw9bnb5xFyKwHCCAOI+NP+S2mXni0KQyquSpQIOz
SwpedZpkXnySsOFVEhTAl+DWQn2r25wNIXgmkrWgYf0xaokVaqPgwASJuFavuT8Yszd4Dnypazkp
qNKETGrQmpF8Rc6sdREoH/O008xyH4Rty66ID9K+uC+IlGTzZxFN8dz2z2sDOm/vq/CdIiaAH2ll
TXOVYtBvPYrGLzSp2jyS1hVmxfdgS7Rkc4xE60f61H89SbzoSjfUJ9mm9e6Bp5iQBUCHnq9xgbo5
XsOO85IvR6kiVXH7wHWo0NG6YgpInzG5Avl5SQSsdRwFWEqIHfWn9dUoyB9T1roZaRMm7zzRecXt
+m4XCjFxV8Dgih87YhUhTxP/UUe4dJeFq4EO7WZGZ0OW4/F3KKHrQunO11983FyJHrX9P8INM+Jh
cpZUIR8byZDm/OD9ElT7gXPgwwAcrPK6xxRJZJUDyNiwlpR1oExCteOMqyT9Cr93761ydTV757Ga
LtcEZ+3zLHBVQ23f6CiMHF5V8WOoMnLayeX6gYD2OboR4xf3+JQvnpovgxzarLgQNrFrtdbTkLIm
jWvCEKq0UjhxVs09jXLSgP84eZB5sZb/PDTzotew4sAFN2GTZiaDRZvWlB1YB73xZe6JUS0NeEG0
NEL/NvQFb/zQOKDHWxEkHErY3C0GajsJeZKkaZeh0vLEUyJP+vHmYNqTstqX915RSfpj/ts5SEee
lYvUzg1JBVbRc1ostH1J6iMTmDAk2MaV1qRZ0gQKF6mZPQ7pTLWxqZ5AmYww/7FsRqGWMWFCTB0W
EiopeqmWMRLoX28CeHedUsILsX79YxfS8X7gpFgh7eNmhRpPzlRP8ltS1/tSXf0Ej3cuBj+WGjRN
P9HNCVgem8kVdoR7e18m89o7518qX7jusjYmluYwxsnU2LtdQDADD7KLEOYFWI3LER7yT6DyKnWe
LBunfI5fe+LxOaKkWHl5B9rVc69f6Kcr46Cz3xNmaaBTccj545xCG+KDPnfkEP9XfYC3QRZ/Vx0Z
LJCG9wRaquj8biyoIqXUUed4D07hMtw4A4XitJPVA91w1mkyb72BO5TB6ixJoEEiM763fGHDu2vZ
7DiyiqeY9AgBVYiZAZwJ29vx/4wazLBv5vgY1GmrZ7A+P4QIPIBjxi/bpCTM6KyTe5ctL+bW8VL9
f7bR9CB5appz0tMkYZ02qB4MDIqbtvrNFH6fOY4R50CJdtso287ytU/cvSTfAiXCUV5DXSCa0o/u
dSd+cLDsBE1fpwfJGv66jlGXWAgSLEGx4PbQUTsPCfklXbuYtd5qNij4qhCERN5vCHXElf805aoN
KjycwSEXq//TsGG/LXZIDn/RKz0RMUW4MY9CDnvsY2Pd3ichQiWpX+9t/QlRKNraAmogWVMLFxId
JMWI9i8qowNZ6Jd14e0FAoaHbxi0WAGlXPbkzuqppkujSFUzAvMXKK7MzUt9GNk+BoqE/r+0tL61
fziQeaIYorue/gUNb9E5Kr+UVjFzPkbEOJEQhVArXICVJZD8s90J6Qhfc71YMI4nH4NRxhZmyDLt
sxkdzXGieWE57oiU8y8/g0y4azOBUzFkqfKvrrzk5eqnTZmja1UfwDyYSytjS63v+45QIQmpZK73
KVHjlaVUPBoRt3OfnU3HF70R0vlX7IebSu2JZZC0nsgZco9sn7y1ncNTYaxjXMikKlFKTsEKOdvF
mFzrL1xaxwixYspIz+xXMGmwBzezc2kU7d8xHz+yzsf3ceGxyB6175zdm6vfV+LnqppyfLGEuF1T
IED3umT6uVgHLaJyup2G9qhFwqJADwZ3fcyvS1CxWITmuv4vD4R49AvZdMENLNDCURHP7rsL3Ink
tkbgAwDNog6u85HH8ySEkqjJql1xbF93bcghy/eumM7U0UQZzqgHgO2bABPkRgBUjWujFZZTOohQ
VJ1/G4Mq13VyhcVoJCxAXLuvlkrWDkw9HbpXZ4KHm6t+kbGgIUN1EPg08O1w73h3qJCHV/mxGF2O
pFuuoZ9Ligk675BqxWGZAKXpyiyce9BSD2J2cnnl+NZoI8qP+/ns7dTkqvQXGbh4he3YEa1B/Ciy
wQMAGP208dHfXS0rJGuNYusbV//UrpVuh24CNBIGfU4yBIUdfYFj63LkqC4fWn5mGpmHu64gP24z
MLCEr+JjVjvkdqxywjCsU2PinKA6iD/WdGCKMjH+HEj/q2kKGw4BPCMakEXctqWXwt1GwwBNxy+w
Q/cTZRpJsmYYKlR/tI41RFpbgPskCknXUefmMoFnlP/PfmdLm3jdYkMnwfsCJCIqSe8uyf2fMVw4
W/Nhio4rxIfIVxU860nlebbjQIlL8FTxNJ2bSAUBg5Fex4gjw70n0iXTHbbq1qoCtelUnIdWl7kl
c1bE/w3KAjQkPkgilMdJKZPqp98Saxe1+jaIsc8qgBedL/Vvlfny4LgwpGYG3+3I+HOwCIs1wiRp
+fhqzQhUiQY/MwaBWCUDkXiqiyAYL/1R8LlYLS81TSvNEVxbTGizUcS5I3cmaVaqKo930gSN5Dvq
6hFoWJvRxanEOcrN8m4TfnoFQDElQavUVt1o6zFbNRHoVjtr0fl4vMMFPSvzEGmQv/VE0JzzDA/S
UtyFU5w9OERWRm3KrSbY0NJUbwQJfg4E541/UacstoboyVHz4kVUNFXrfMKJB8bg89NWybte73um
ozMx7W3Clox+gFFnT8zZJxjG2qNTVg5imnrpfab6oNadAxsSDkbXXwOFFCE2OZqQi4i4TZq9Na27
QUSlfHNLferIRMD3OUl2oA3twJaL6o48H8lkNfuxCZzbKGFoAA+5R4ktqtxrFInGPAXVwdHZBoKL
jGydlHQUX3aOLa/+I7eUMO7VaRuM1KIH+vmCTLCQws4gNUFLLlC1s7gJxhItsBPhiKfsy4OGHCda
2O6k2f88deuyKIi7UyocWFjSI/2K+AIEc9OERDvkoHwEFoXskP+COC1keF2PlcaZr0tJUOjzUY0/
MSjuWOwj5N0wbtxA2Hqpy68q4kC2FT46PlT5b7aAl8NyKYEX2uT0eQkBrlj+M24LAqpgTxq7Oxtw
OS+FFGwBUqrikJBhov99RFti2km5S7MbnQwCWrtYywcTnVZFiBVp5pAwo4U2D2JockQw/R8pGLH3
kHg+v9vSgThkVOWED3wNhBecVyD9QPCxuBXiRmDES7/eBFviyL/5p2kq/uq0IL3wwfUklyMl7SP1
F6+Hi0YcYNvr4W3KhhmoU3V/JIRZHEj7RrHqI90uLAQNFOPHQlt03lZ0qPhPh0QaEYtyjT+Cqz2t
A3/JjLYBE96RxJRuHJLtE7j7/B1qNOSsj0lZBwr6IkN6+n8KWMybLsjUPGrQ6Ff9mCvOSv2ZpINX
6L6Ls9UCjosf72nLOK7InoNRDX+I2C8DDMYYI0wue9I0IZATUvboeP1uE87wkTgzVLu25MkWcu5j
1mFZreoHImp+Y3T2A05FqGkk/daVF2FHlPmHqS982JTFXVUFPsSr7fXkpQyl6PX2eXBjgaCDxt+8
NM9Y6AgXBAUGo6R0SwQwLC9TV9v6Yjmwqn3dCkavAEwvUVs0G+xpcrh85vvtS9nFzoh5G1bg2MWW
Yi3D7HH2ighQAogFcYmtB2wGoxLWWcat5cnyOgN7h0tyImtoydUAv8A/Msmguv8VJZXYbLEO12MO
pJszA3pKJG3b+Yc1/z3N/BsZ9JchcJzcsjQcDptlxQXmSAj9YcukDFIuQMpCvwL2BCqdo+d2HBlR
KLmww+RjWxbeJVhIN9ljaGrya+x4wn6P1AAksH2cLri/54Qevym/4Z988n5RlwE61UJlL8zaeR8n
FnEO1KyEokZfT15uJPsze4KPaud7p8T5VLjXBQ5foqdwYTiYmYdEZYi9AiNbASWJawTyhpcY6Fc/
ZalnJc/ceAqlZ+BD3F+ldz36xyJ2BtccTFmBOfWcrk+2BIyJmnhYVqU02A6QEb3cP7g7EdYBdhxL
RUG96EjEAXzVYK3ACZJggRbGUaCM9im9pCuhR41DU6dFuEc+ap75mElKGs8/qK8tUQh14OOEcZW0
EJMgOYn6RKvSr09rzyHgdZqb6xvvZ6UVZEyO4ukIZGphMVOnAzoXIt871AtCJzHZkKIFsjDWNGng
VswK6I2QpwxDOQsyvBjdLz1dgnCFEE5Pcli9JPlbPs+tCg8QXzvkbv2p6baBIyk6lcki7su8hyb6
/aBdePbjILbLYl8srtz8kUFJVln6wjM9dtTxPa8efEknnF5cQUoewWovFA/FLqzMRwRJjxhX42F4
DZUU16CuwFEGBFpemq5t3pHhHSDCXNWiYwyW0ROWU9lS2ts0zjKNyzplykrC6KkgQBzrkl/fky7N
WUB0xDwHmzL4i8838J/78lFvErktw5xKIA8FMYXsf01QDgI9V26N555PZcYk1Xmc1G1Utiaypa3e
bRgF6SphU7m7S6mdjXaJ6eqBBw7HRvWOmQluG7KwcMtTuUJ730E1I8QhhaIaisQxHgzfvK5u78Dz
WK9kkRmPMABz5cAyA9S4OhD8xwSabbLoAfBxb1X+qKP6K8EPLucb1gO0aQWbV8UjUR0IVHovuqc7
wvHPWLNEJLiBFO49h1GXMc1sRVHqtvJIDX/07iKbKLI1KYnLkQ6YhVPPSb2HWnyvZVe6yLUwnsAW
I1EoPtlV99G1MSjkV0ZbU2LoQpfupT1ykYFu6nV1tmxzjTWkaRF4C+jKc7eV57jF598Mqkv/7ROr
dqIzNmdH7+oAUHCPosc29ADpk/PT/NUtAcE9ffzlAK7XcrA50/q7VKEtWf6+DATilj9FwjLiEAhX
AStnGBGb3nagr3Kvi+FKszhqySPMRW6JmLl/nMZhPA89cvInOn+WaYy8zoxD11WgvEZ5u1NkrRdn
wBGbymbJQ0zzDN4dubZrFGbRlRePuXiv3+ZY0Os8sOwbAuHqVXVJAUX4pxlIbvX6zO5ECmTyFHMc
EQBMr+KAXgR2FI6qrnK/iZpFwLo2ABJ6l49mhR4AGAC+BKNke0bLLxcUXvciYBOkfWbZSHsIQUR3
gDAbvdlket7s6xo/x3S2wlNSq9bTiNj/xnIXXb8U7J/+OW3SVCsYNv414QKQBHG4CnWXWUxeidUc
tUrQsajwjcL2qPURgrHoCJgSTtXP/CBwC2PKE7PTTy+DedtqECSUBBO0h9sBqBGetRH2BdAf5dU5
bVyeWKQauoomMkZ2TBdcOOT4ce1UhdKSqYl1rUeBldp9q+QNVK7RQogAcnGeDsq8h43xD1nAQsEV
b6nWSAh+wcQzO0U3JmBOj7Xhq3x82k2GT6lwjSp4e0+KI1owf7LTUSPJVVDdS/vkrwCb7LmR4AjJ
bS3lV4hGGLC+hNlXwe5qJ2W8KR+vV0xYNyaXfXvNNRbMlroFNLT2+XvesiUiHi/nKM8lFglW6Yb/
HJ98nuiMMyW0HpKSQAnw9vQv/HA/ip+aC1cItJUOwtJZrVtCSjz9nsYIkoDd2wYRatn0yAUhaSb0
RQT8aCyyHyeTAACs/nmzUhTTQMvTYqJ2cV8AYcwgWl71wZuECa5RE4gmAK3O+Ux4LHas9DMH8QRP
SfT8Zu57cU3o37ZVAOwT7qO1zisIXAuGRbt/dBg2r5fqCcRgSQZDWJyNKHJCwL0aVRbQP0mEpps8
Q715syQHHKu5Bjuuhq0xwEiWVkN7UJrjnLdsFis4MqveaF9vZo3mmvlzPMQYpuCPkRVQLoBUwJ7t
njbtqA3c0PeCifjeDHaNrcxCcUQYYA2op5zjfDHaKy3PKwE2YZntoi7VRD3IWn0lAmAPX9Dc1ncq
s3Y+qzJQ8q5emiTqGLIXOPYBgBO+pL4nM2fTMHa6CVE7stFOoFk1cxTpv/R9k6OlMUB8hRm7xyiX
liDwIsmQ/IPJo7zGQ9zWI+1jb6hlP/RBCzDa0rBonjEGh/gd3OX4yyqa8PbEdBXmVYEcX+mP8HAs
xgEmW7WBGXAWh6s2JJSA4Gcb07FSRIuWwRC5ASLntqNrnJFVsYAqLl3FiDMXYYCUr/XTEPMMhYnV
rlsKKVc01nl6V6RaG7W+1AFgKoPRfx68bd2FyfpATbiZymA1+OxmQDmfKyeAqIPdICljCXEgdCE3
26W/2Ob49Ze4KL6FFG5QPl6FWGTcWZsDL+rdCciI0nwj7LuTr9WRDoOKYSnAPyZllBbGl9IM8F1V
2ZGixLolP3Rr+BrMrrCZn7z5e23AQq2oGVVOvo4gDOMPZEDL3fLwAstlazrrcGG7ky1lo+sMBL4M
PFPNQ6SxIrEeTgrnT+BPBB8o0fhV48AsoznLB7+GpdO6P8VtM7aF99IWnpJGsHQyBXuUu/AOm5s1
ZR1QYC9c46YecDlAxdRAvFafV+/cVk9fzJ5ZEDpf/X1Uf9He1b31MV/fWbhmXca6eR6UirAiK3gW
/b1zZ0xig6ZcY0OYmXmgRZcs7qQ7Rgzhk9oZ8UfH00QDLwOs7kJ+Iz6XJlNdkKR5YeY03ZlG8c6M
+vbHzHtI4aQmcVgHqs9aXkaUjqZuwVnvFuQHAlxDg2qbYee4Kfag6LfxYuuE7jo1pSajZCsmUbHN
u1kK89AnNGBL610AHi6dv2XrsXiOt/B0uqWpX8i8wOg4k818gCT3WeUpXqyzAckbHKij8cBwebnE
UOussl2a/Fbk85n7gdUVImSw/XrPjNI1Au1pKr7Mdi8UKDlHPlkUKc/p8fSPYPjphfwRrgY5x2Kn
P7q+eG9bMzmrr5WvLG1ASG0w5UEbsI+gXfIXEH/zTE5AD0YVF19rd7Y3QLEmKiwLH0htdJoL0lXY
yXedAfBcoeB2VbrzbgFJQ7ULoeq18RocKgmqnEo1wYv9kRWbCObDCwz/JMdFPUalP8YoW+zOh9NH
yv6NB23nsXh9qVsSQn1Nels1VXmfJ30DxjGME92TdGj2wmCYqoebjBA6Tg7OoxqZ8SFg1KyfeWc1
otJBSoeemGG99f15du1TmhTM5FWE3Mwb4SbYGWW9XQdE05/NoqDw0XCGhFgWuRJ0R8ZIK2IeLw4r
MEqcCWGjBTRG8obBV9WSZ9hYSWOnWJob26viazbXndfgpu4ohah9GVvntXXVwByS+ruk7dbCzl3O
LpuekyuqK0gFgS/p2YXUyWRZ3AjU5hkQqyjttCcdEqs/HXN1sqPInfXfz3YDaNNpAL3FeO6m/bqQ
DvhribyxqTUvq/JRc+n/w69hkJ/r2sUWinB3VzMbstZclxQL5b9xpQ+J8G/OepIW3oTdYkVCfJWZ
Rzz3Vof9DzBsEWiattXRCKqVAFyqHJ5c4tVSdbbEAOCrK6A3mS0BASiqqwkG8K11qLRDaxX2SEEf
lEvXaMGhghBEqSLH1DjRrbZD1E2vz7R6NnnoHM/lUfcCQmCXxTe1N5JYbnvgYzw1R6hyqe72rDKC
g+ahLSmepZ2wCHWbf2QAyVlhZPzlB8sbFAkczsNt5F53WQ7gqZgiNzRCDfKgOw2ql2HM4lnU5Hy6
rEYD2nHaGiogxR572wC3f0gCS3uGv0bLPfoqMEPQaoM2Bk7lkjRF+vySp8t5+XbhqyjNZQ154xGX
DLs9FOmD+sLE6efGv/uTCqX0lho76SbPjAJlMpVLpavCmn5ECjvedfkoQ630n0+4Yur+a6T6vd1f
RY6A1XwtkbFZr+W3woKVBeIFr810tBL/ZZUzc8BU47l1o1is60x2hksUWumj66ahpLHhZIYQOScx
dzrhf1ohWldMvWWMfSR9tXCWq2kgKc4VgmPkRp2mxc6EomLI2mk9k07MrKNrRprli25z63aNfwUJ
bb9ATjFlIFlt7hGsNET6lvbVWbRoJYac7jVN21bmR7D9Npaap9D1oL0aCdZ/sO5jMsxVqiJVwfTu
NF2Jk3Br/GB1DhT+SSOyEGZG60c3oHfti68/TL7fh15DpDemIHtTkAixkg06kzyRJ8YTfPqd1tNZ
I7IPyrJxWcLetBinXkHGEj64ofHPB/RFT5GXgTW3PlRW7v0OcP3Gdad86rz9Q9zAVPl4QhyK2eDF
NJHmqUhvkzBMZ+R3TamZWDLzYmJMm5mtyn6eU3Z+M7FHDsQaFt9m93xVQkKYl1g3SNw0RM4U8aQh
a6cH9qIzWuc1Nr3//h0a30caDmynXgI+zLIn3lLps9lE+yjmn2QlvaJqzxBH+/2b7qhGeECp1Jjw
UKjch5eZWMElJi0vV9e1mchs4QMNza54DXUa+2i00ZxUmxzItYqm/F/NN48ajhrTuA0UJ2SX0GuG
ZA9Q9R7Wjfa+lVZp/ABK15zLDnmTe/5UAg7PYuMVyePC2mn9ax6V2EWCTZmxgISnRt0CS4oVeN9V
OtPPWdPgB3Et7rhaEwxnipnpEJ3BuebVZQHwzs+U4Uw194cBrFv0aX8DRRnivi6gBifLI326I8Z4
qsJgPJV4F3xGZZxXjPMBYkRJB2bdfmlcLxJ2xjiOnfxzF8Kz0Ri+Wssbl1zRCnxlvhJPpCapmDOx
pl4WNahQ65FNZl36eEBWV6DVLK0hFbqGCivhNIGroL8moBjQPQalPNhyv8iiAppkoqNJLI+dO1Mq
Ud16LCVDJLnEZ/bsPIuPd+GUPH0TUx+rUx5GMR/qkPR6pkbwynBu45cafgWXGUSsbOqVUjkAPHq4
5UCYwz3ImVSPlxapmCnWWzE8pWL/zeBWFsM59XflcLpkKv4L9O3rPq5mUg9kTZc0mCUchYYi4yXB
RjZItXySezjAMI4YTOuMXLgClD7leaG1fNir5ULuuCLP7gKqNeGrN3BQ/CcrKOUwEkNtZ/FLlbiQ
ps8Qeo0BrKhCjntRbMWHR50a5dscAtUe95bPlxdf3C5ZWMCn3VQXGnGDvgOyJNXasX9l3sasLnTZ
hen9LmiaXuhHI/DVkZlYC5RXVWITAX6m19Rvjn9ATT2pflD3x67whfBJLRyfCUG8Gwo74iaY7LaC
1S7YHlCmYyCHZUgNmTSQrjyFxPYL4QT0iVMpfobm64V3uGvDvdwl4FI/PBGxWj/NLoM+S0F++Q4R
QvFiYXpk7yWDq8z7DNiRCz0S8x7SI66HdyQ02IrrMqjnZZm5VusC9z4y4REE0kuX7CPOP573oHLS
Cxr13BR3WBwsaFRORS5LUT7w/XzpIT3DtlWaveBHhPfqrD72b9gW3zUwcDI7tNs70ho1rsqjwIcq
rMGKOToczNuqTobjq1Xc4/59C5o72criQlc+4Ry+MOBAsKynuqEFmL/F/t8FUf/DH/6cG5ruIrBh
6oZ7DkHrAPdW8ry/DPnV/vMKYtq5Hs9dfD0//cDLt/RuB6iFNqmHqY9XEDh13uA0QJgRljHCWMJ9
1Zs6Y8EdwIJI60QN0J2R/FN0Nx0Zt9q40mqSChliNJpMD9u8MnaBGks8jLQCawDmvJjKsjnB/mz2
b5Iu00MR68nAHsPNu8A4cpKd1fMc2dVLNXOwIYbn4pS58t3jk+UYXdaIEFMrr8KvyA/R8CqlJmEy
3Ks95mrz3Tzn4iwhcST0hR1ze8OdZgqNnTWH4EdBuEcjEL8yeFCmeEzkgG1VKZAbfmu+mthAbwNM
Hiu0xSHLHxnZKMN50QMISFDZW1c161mlZmUKEMh4MzpW37DBxm+8NONNYhvZAFT/VRD2z86qn0/x
wbfkMgKmAb0UR9l7ZnHWvWQvtZ1wb/WEShVMIEqPTmGQRrsr8LFgW/o6y4u0fIOryTBKzKt0b5I6
1Urt1dkqb4XOnaddtSp/H2iw/YRlWkyQtRHoMeKny40DV9S1c0jtPJBne/EaFCnHZSYAE/epXAmE
ugcZa8DotHqoKFIQbUTdhFvqvPtdouBHZIt1O6oursGX+fFXnfWUYs2Q2B4HZaTe2QYbYnlnRQ/D
PFb9bFvReKfb5qptPUdA1dBDiUEjm3fqjkCmlNpbKoqT9wh1iTbuviUArR88JLqnQHGTKZCy+7AF
BfJk02P4GhRZlAkmd7efqTF5sACIZF2236rM+YYGq5tVsVyl1T4ekFn/+I0riOxsIErrhAuWJDST
2XRjJ3d5uY/elO9VH3zwGYlAMoROXXKiSxRhJwgD7iXce7tBo/X1Tp1tzCUYUNlw27kc2FyfKpof
zJ6jjXgangeq7lmojtgVq+wXneyMvKBabVcBUcY5A+PNEjCLNlq6AunWtf/AUqOpCCiMxZfq3qhE
QPUDnvOCva1V2jWVHkwmWBZaAI7V2bsr1ggi1RUOzjliDjgzvSA0zAJ8uU4ptnCw4Gvg7hHfuZTt
0h8snJdr3FqgvI2vgCb8VjHI501HKaEkyRYTFelN591po2c4ol7JlcMiIkrHQzr2xPUBKU2o2RqR
2W9fQ/DXPOy0/HkZVLOLxxmZE8g55ft2cItf8vzi3t1KEOQygZe4Y57vm49Y4rj7spQvOyJE62kQ
vpfN3YRDFgvOwvB398xEkmyDj4j8NuXh2H8FfrFEdkRzE8oqnARRRX9AaiYsIDp0XoN4r1YTTbAA
/WyURp1mIRB1occRNRZmaZXWkXsbIYAPDEkfpUPzhR544SZABCe0MASjD8FVO1dpqvjZFbitN7x4
+cuTakrWFBk9qSQLnwd4FYFwoU3675LDvdl8TxLmUark8k2VcHWMHzpJgcLZ4ppTxOd1UjuRMhUD
/l5IOwaePD2vgcZY2pKONx2ZLh+IuyQkMKwKZDrOhpx5kAtXfOkJsM7X3EGsrWa6iB99/V8SRswh
7MraZ1nIX2ZDkj51PzUC6jCIbrDi/pr+vIGfFimP+jbhLaMUqI0ymrr8gnmcCHtqollNFKBrdYuQ
FGRZQuqGKcfIMf6dV4Hg9uKzYppVKVsh2e+1RiNxmDu9CLdtLrmIM2o6sz+OLUHZFrTrGR2t0eL6
s21Iqv6WnbUHTkfRITE473Jwdq+ILQ14YNJUSvPIxdAD6PvxAfOwRovPfxmH55Tl6P1MYjTvF/gg
dcyWiQRyYtbTCrkIVJ44Lk6gJyKU+3SZNqAZvjDCmMdaptkUV7yzAqIX3EolpNpsJyAVYmSz4jgm
cVl04AjtbHJuZWFiQXKJQtL4kgk9s3Jft4fKvtD3X55eVeWMSGEEkhPuUKLjeZbgjzdkSdgXxHkF
PTMK/JU91QX/I+gFqvktGv5bl5kNbC7a4HxBJmUOEdxlR56pLIipnWmrDjprXzzSyvX6WAGnvsw7
w5zYHS9oYWjPuJcgnYXbD/B0r+1hn+m+CEBrsCZN0jDEZ6Q7AuaL0I2pBe+ACICSduVNQupB3w61
UjD12B2TiQ3/cv4QG65oDZXkjVp+aP9fgrkoEa7MJIlpI+j7n+yfysyfJNf2b8XYVeUAWwO9l/FU
9WxJ+0MkxQYKEqFclImxtrBH2pytITFzimgG3ARWpY4eQ7uJftR0VBh3vY8eMhvxM0IoN83N6fxR
DbNuZZWYvUqoQANOqNs4PITzDqO3XOO308MNNNmO6MuZkuthIvGmdPtYcXTeRRwqJ7SPMYmn9haS
P6RlagHtndVCM6wBhWA7/ZuAfbBwjeWYAso146fqBJQ8CtxI+jC5WWbdHDSiBrszJ2PCg4Rjz5FH
DVZeAVkQl74rvbW7JnO2zEpw1Xp0jALGy79YYfT63UERBgEOFYO7dxq/Co/Y3ytpIa/QdJOP+eWw
xPySPJ7SkGpv6P3um2GLYXgZeyRVMF8e+7BJEvunSQ6ns1umWDDk2peWaJBPa/I22g2tAKh10xlo
rC8mGUgaRq+b4lF6HtjLvH3/nDiFYKYdnEHciU6LBmatMUikr95dbJzDv0mRgKBjtsdJD4T57R2j
kCUPUTAGm01//R9CpCcwRSmFLnDC5aCqbGCcJzOU9PA52fi6bsQQpNpCElVvLb/l5xJycG/vd3W+
7cCcXYRSIm30OQFZ61dhr6pisls9snwlxlRA7QHCYZB6Q7qNKpbeuIcko9q8ArKMMDB4kD59hA6x
nu+ac3+DmN08OL4od4fxTUsaXEi0RhAiZm89nZfase+myPazDS2TVkbzsl2OOPW1qBZax8eHbjyY
w+K9JCynCG0mKbWyrP/XBlf0bINB90iXx/gaanXwjNhAn/ak1CVadA9xGZJ7sDuK9oVEBiPq2st2
F9VSYQF0hB+B/fQI9MJ38d9r9q9dND0+NMqWK4Fr9D2lfHUUbGE3luR0FKyS/ICgeEWiViycTcml
xNy/kPumQGJvtZxJABvnJDlkUUpI9II31dsP4muzC1Qic15FbdPq3s2CldPdkM1xWdZvBQzjRd9F
6IIIYknR0l3H7bnOnSk5mbSYH9vt20SsxsGbt/jas2RgqJQ18mG9Vk8ac/dEOxQQd+mv+X2nMrxF
euLYqMThgWK14IlL1TxErf0asWZYYWpdHWO9ez/qCdLOM5HCMNQhyn8qgYSbv+8+n7h1rPDBJFSI
VmlE9gEf/HaWhdNgpsQVdDFiTTTgbBpOnF0YQm75KcwW1671HCEIKrSCYk2VnDWLjeTYIQRh1yWM
Vjff5XK1SBfmJA/t/Eb2hEhgImxJRrluclEBZ7uIQSxmLBDf+VtXAwMr4KS1zC7DgD71DWk4cKM5
bM54w2MAgvA8RXC7llP8rsPCMypC82vLe97QkkinLEPZY5UlyeyJ5Nc9/+z/xyAncVg0TV+XGpx8
ikG7hZcC3U+EEIIgc0x/dGEGP3R6fyFoN5vaJnnzvNEI3CXlYj5v0H8BqSB1FBrLIR0N3bsXHcnm
CcncEyFDiyvdjChxGf/wQGkrGzvt/gsH0+OZj8K6HHDTF0ER7Cky3KwZV0jp/+WUXQM/Xu4TT0dl
t8SouS7yAYu1wFt/0+s4DdqA800/g2AIRvBy22gkisja3T8w8AFOOzqzEGW0sprXkiaCQGTGfV2h
gDlmkIk3uq4YkQ7uqYjESabkrC6XXki9UiJb8jNc6h10XNu/7ccZEU381zZtQlu2UIkn5Nm09ROv
7aXlceJRIYXDN+czDDjZ4Ua8xLE5fZmbFbrnxRN9XmkjDLG1T8AEwfQ8dsi/wQV485ZOOkEFbeOB
TF0nD8lzpjLKq25SJBG1EXAhrvDL86Vo4ppla4v3zyK+Kj48KoLjJOh0SYhemXbg8UvqA+n0yzdY
T73o7FvHd+73pepw9GWcuda/7ikRsDADpbk3seEWkcJCrWUOnAFt/n6VISYxcXq1AUGOTA5ni7ZA
W3osRRTG56NMCqMu93binOp9i1ZaVjfqY2KlE6WMxtHPhn+WlZ3zvEzLwveOCUkqWH9H5ycU+rPA
myJ0+UhmY1b6bkSau1yl7lcs10xsVfdVErwtm8qSgqvWG0inYgmOqrRFLhCNQnq8VhLxXreKgtHM
Fl78od8IzYcjwmlELO6ad/3Mwt3YLIYkEzFQCFrSMoO62YacKJEA/THpCJUG3y29sJcgzW49fw+w
L2J7UG3GeMVVT8nJLKWKBw3I3w61/FDKRa8kkDgggPG+my2SjbDkrc/s7uuVhngTqT89crOzLgVl
YNZ7mMxJp9psjhAo7p5hvDpGrUP21vs+3G1BnXc2vD9akfgRjhC6owpWNPaoutUuHRV8ON8lvBBU
JxfCuwePjq0PPCA1Vsoy2AwegJ82NDScc9BmiH/gqArYfDnIJP6pInicpVjfLbLqFAxjsqk59wpQ
mRINguy8fIOaXOXkG6p+ChTOEKeFEMeppmkQAKlTphuyiiHIO0C1lJHuhaOKa6fWX+3qqmUxMQ9u
66y/SAydDrHg9k7vuItz5QlP6InqBplmeikBoZmIT0qZYMmuY71JZVlyO2B67chRylO/clj4e77G
EJbti7H4M4xxmHjrMtW+kg+snk0s8j77uvklZRGUTznqCDOceb9NM6ZwQKzeH0V9CDlfBdQrMkEQ
HSTZHpunkgFw4cv4DuMsFmvHTGC/Qn2qkWZsr0ieqEu+2s4u1u0psSSvMhF8raRKEAbOuKN51vAb
iminytl+HQ6WiqWaJCvJDwu+yHWNP8PkJaj61G+IRK1WKq4JHsIqUWKDcjzRYfjVll36DAQfC+mR
l5z6mE8jhGLYLmx3CuF7AFhzr9DCEQC4CJTqiTX9p0PNMVukO/G12v/gxogKgcCgjp0w0pOeTTDc
7Loya44jamXtMGV3ikalAXGsdEfort1kfDzF/PE6jhPAIUduuX2W2G0qtbhHW61ZjPiLlC+PvyLf
Kyn+A/c5HW9qRy4U/iFCinhpsKvkaEwY4r4W7Y9DHwHQxW0zL2XEhd+KNRr2SkoPgvTzFVtl6X7O
YjcYdkS92hdyLr8kwGkL6oEfQcNcegoufuzfIYXWN6A9ODePo5/2nN77JqbIIOsih/gkPcJvK9NO
XON628Hl8ojUdx92aIysArEND6+tJjY+lPmPjby/iPoClx1Wm1OuA1kFgWlg6tu/WmuwZOfad2n1
aRv4SEU5zifJVCWaN0itMUNyICwyMGPxl81HadNHWColdsLST/OqUWQqpDMsDZ6stH7FlSY2KutS
kPdr2QE9Tx8Q2yqej3uNKpgw8oWOVZzvLx9xcNgKkERAAQ0tG6/ZH2YN6+TU1AvEsM8B3pMQmt4F
nWeviP9THtC4kDxFDAU5t6pP1YX9b487+s0iX1rOA8snsYsLh/bKWmclXXbUhcpDF9gORKtBYH+o
/MgjNcOoUKS5FdVqH2Gp3Ub0W1XT/trW8eTilJOJgts5fwfnPXpoQL+VRdNakkyz4ZaPxdogtETz
7CYZD5lMgcNVlJnCcZmrYrhOJeBK7rCvl52sbVlhSk+zoT/+lahKC7iVmAgtgSzS/2tESKWmolp/
tv3O3MNhrQDOojgvkQ6CRT5N2zZni6lPXSu9LVm9+Nu+plfRbmVczI2kwU64Gh+cjQWMusOg1XXR
abG4CdFr06/mCIXKBce6tQmFicmNRMWE3QXIcAy2ziPYuSSGOzuQPm/yTO8aSQz/Oz1lsdZlKo9v
XNR/UO7PDIr0vaRK0+S8PkYVs6yHSUl3Yzy26v5U1oEY+0sl/gnAG0WoW/yraGKZCINrdXB8CPWv
xWj+/CP/4I2PJp1iM3rO2aHAKCcX1acZzZrxtH8IKgS4bxj0EyQdlUxAn/ySdh87G29gxdjVTkdq
+ZFeSdppUT3FfBKUN2ilAhucjCXZ0r/qToNg1N1R6Xt2rG7xNr/dEXz84uIwjpB4O9OfLo9lTCEl
CWxf+Kbk6q14w/4MaB2XiW4UAG87AxCqjiSKoD3JidwN/ardY7a0PyucpAHRRr2IlY8d7APExCTM
WtDfF2Hx5fRuv6KqcX8vu7raZZM14SEKBF/6oBwl+/pu2zmDZt08LK2VJVD9edKdGsmxDNMPxIqQ
iX6c08G9OWJ9U+lR+4HLIwuSOlDBQ+la7W8v080RSCut8wIqaK0Q3Kmc3eLjUg+aCuoegK/gMk82
/2zKhA/iv3/xlTBHzXDhi7/kN/kns5Pov587l4KJ47cyem3fG+jvMEZgEXHcYs3HSHE+2S+8k6mu
UoXZNY5UN+vfR3yeYBt87K9FoDLzbZ5RoBbbzdISvS9rNJBYI+5kCheBDf+liwsZ1y+Tt1zDBmF3
NsgxoDHNQjeQviZ6X3zve7vvrbMbVq2IY3LxzbLL77rZL9LY1/x7ktftl+0oO/Hbob43c1GqYABv
SeJOHZVhipQT+49yvbDnEd1img90xf71p/+4txYrzZDI9DM5TtiScei5OlfB1dPLcr5xHfDRBZay
RV4hOG1IkaDcC8UVKRzqVWdZwvgmctZG3uGM1a6j969yazwZPrGt8Rvc8/10APIQ/BgSPRWcwPFs
aMQFCOMJm2AGKFFkGdMXRjQ8qHJlrs2izkdpCv42fU91mM14qirXIshy6/ypMh+KQmPpe5vRZNe+
coeViisOdiFKyyrNAVDt5jkOYKPKYm+fklKXQyOqWZw9y6C5/S9DvzwxsG63Ta1x4uF8zG7R+ZEc
d0YEdt3R8OOoph49FrkJhFf9v4dh4KQLy0VjI4XNnEz4zA14abyI4QcRYlS03WXaRgUx2Lk5voBg
XIPb6oI+DQ/RnqvN5cbNMT43sHELJQ93VW6VysDMdPDARO3rJdQh3Uf+VQLj+HQ3XCdoaSRA7LFg
aNow9yG32FzZMl3EpSHC9LhzP8WCX6C8ba6n9XsekyPfgbuthjpgvqxOqJ5w9cLAV1gm/xxlFcCt
p28dgIiMzzShzrhqBqfRCaXmOMv6nubkEasUC9FW/NG5la2c5IpUaMggq7EQV2gB3EWoOgB+FRzH
WR80iJD6v6ASAHu1FPPqT5U1G6eAjYojOdiMqlGcTi1QkTHPEPcE7SiDCtg2T9Z0kRG7sKy+r5yn
LMJk+NzVpUdAN2qvlUuJZDeoiUI9dAQSmiei1/aPJXj7LqNgL6VLNadMz0g4CTA3TCIY5A/orlc7
5RfVrLPwjqwvBDTJmUrU9eAV/e7ZNpkLOzKyHp8M9S2zG7QHS+Lc9/Wqm1FPOPCalHA9Nt5bb4uU
e5POSWrIjSS93b9DPCCq23zQ+sO1jYZlKgEIC3FcMWOhp7DTxy3mASJLD5gTcuuoHrpmjTm4U9yq
MeLjUtKouO/JO48luVFc9/jnbGxOdHLxmSWV89pB5J/UNWHdN+0YH97EAz54HVb4IJgUFItlCzU6
Jn7O+TWkqlqvaur+MJaILPq2qr9R+opgDJL1MdjAxzgNfbBfKI2rRl0NqRPwfKCZGLogwweNNut8
akNFNs++R8926lADsGSHeq2UDn+QWl2xj9zCYNG9QHCrvE+mNPP1HHpI4UWePIIghbbShHZbVEzP
eIhNdzrNoHEMlZRWZvKAVZJsGv5uJHmMwlH102Nhq2O6zhzWq6Doz6L8mLq1TEv6PVQYwNy/x0GG
+USl0rgsyjLg+VGl6DykpDzbiYbT+zHoFasDdN6qkzGhJVWAs85XusQhSLgQKFNamLLNRn0IU3IM
0Qaqr3rWAsMlJsITLPNYcH4GVHURb8HehinozwunQQbhR54nXKJdrEVu5khP6jWzTpJGDroiQdVW
oPFpaQLbzd7AK6plLykYG36Fr/i/50hJQQGcsq3w3sHjUnblfNizTUMcfXNWO/88XzlMWZlzVOCG
h3+YLKtX0YfGDrUOIdc+CgGWn3pEbk0gDFWtv6VnmdxrvAO6UmP5KZvGM5/+9JkiDBgNq6p6HNw2
W4WEatZsj5rQ6oPSsx3KtT9aDdXyohVfzX2c/2X+Sob5oC0DUdozsp3/RvG0S034jSYX+owG+BlJ
suroMUbKbqkYWHumdh/LkEM6vFzvb3MePs4yefeawgMiNXQSbvHw22qNOW8DFp6pDtx6Nm5jHBQI
E1sdwne47sfCFs0im1vRgfiz/XJ17tes/l7HQgIuWwtbm1RHPaF+xVxUo/0X6A9NTax4rruiGkxV
9c1kljGeexdscsUqbuvyFatSInDNzZoCEwIQTU5msb33zUr6q53ilvmZTsfTn3PyC1Ri+A8S+HXM
zpPWxwlGg47GEgi6wng8vgaDYQyUDoN0lAX8vMFnsyxRYT1vzP6XxgQN1ImGZUTL/AyX/TuOBLcO
z75LWT+GM8r6y4tSdCWvzC7bcjMBtHKrHwMtFogjcB62JtA9Ixr0lerwsJjFHaUw4DxysHSeHrYM
LO6HttRmolRrDGhX3Yu0/mMV3oVgUPSyLpIFWiBwO82TdeByaHcYfEnApGDfuJ1lZBC7EE5YD4Vw
8BbhhvMvFlXYAXy7S1fPhUeIABg4q9auj0qUwBfLsgr/xwiDJAgmKUymfwandatc5d3JWvjaazMQ
vGDeYzEHWCszRoVTmiWF5+1ZNw2Tj7wwcQUqoJHHOAviEiUKi+3vnWjFqOxvmV50MK7RVtR0idkL
3nhhRpSr5x7IvbNstSYf5doAWDMvM1ltZNRF+P1b7ltp+cfkSCUsY33/QtmRDQuDEl73wj3d9r6x
eUilXrpfvH/DanqNkDs+y1uMMCdr2L5ARtP28KGXfvH8K1WtfS+dCBFAKXZh1YsoOJHb+ZXEW5Nq
LaNk1qH08Wx4cHKD3SGZP/mq3ONeCUDboCfjsOt3DHEHCHHlsxvE3AJgUviovvH1kzwbJzAKmrdE
TVjouI/8AgAIDkmQHekJc59TDnq21AA/zIziwSSpVFwBv0Hl7fmz0SpU/g/FZxBM/liRp7Cc/AhK
SPGXZpjOUO9SyGNvf18ebd33RJrfEQ2s6FZ7FEU7B+jvGqfWG98BxqiTkL608FyE9TSmeJcs5EmP
1we2bYrQpscaVXhEKdxOEo1th4LT4EhaqvJW7gV4nOFe8/0KufpYZWm4IL4kZKR3bzQ7sQKSX/kF
v7nvAzc/isDyyCHXEXF4a+xsUbIudw5PWhk7CaWdNwurPc2vQmqM1VxOxlBa29FBn6WhtCG2Rfnt
vSLd2n/U6PBkIFaDAKcVkheVNjLcMkQzBJYFPHp0OAcZFxm4JLSVi9bDlXsSMIXqjgRE4TiYOyzf
UWPEEMAx3Fmlz2MpL7v0W2eDn0YySujSRseegp7MxEW19KdSf73H8E3UDToUkWzsSr5vY9KIB+Zs
gkVcRAKyCRa0xlPGdqdn1GQjP4Mzr+y+mGKGRFBAv2l+Czy78gfedP15enQ7yiPAJ/Hdv/NW+z2J
Z84C1k8w1tcw8MUIPLfTcgN/u0MuRiE5GUEAHEaa9tix0qxUvqScOt7Qhf49TG4fTWgofLap7k/b
r2rOSe3xfcN4gLnwSYxTZ+8fdbWiaRnN/oiIrABUo4tHfdXha1Q3/3ZqbEcSiBPurRMQWWC7VJui
W9CJEJFNa7Fv3Yd04YB2fpLlej5q/WvOAB/p5wPyZi8ejMdj+P4M658b5yMiFISAHATIydpJoOHi
JBrHQ7TDEstnuKoLqCfyZmkfRe3S4H68JBp9H/ou/Un/A8SnAMpRnIw96hLF4yeoU8lPXafOMZGo
/AjJIpE3kBG21GRfrvkTXNE5Or1AwKCOhZ9AtbPIkOmW0Zov1CnwniPDAEJ6vK0oTLfJ1gABkLl7
fG9Hss2otjtBIvnAcUxxI0siTnrbGNJaFOxLmUcQghroCsoAvU2kXb0/Pi9U8dzo8NseOWyPZ3J7
CuhKyq/wcEcFoV3dbyhYZs6+eSUlxImoiRiQPeX+S2FSCkBWGBEOHxG09qUPeiOaC9AfYqgXSd6b
oRKjvjUhoxHtnCCaCUxSdFYo24oRypDTmd5NGVKgW1qvh+AhwAhZdWQyhQkjIdC6iTOuBraAYNeP
OlukgPpB6nZAT4LIbfkcILnQddPVCrNcZD+iYPGLJnFtfaqw7paOPD0N6WE8Y87XpqSDHuW7wo64
75wxXmcvZ/X1psFs9a3+A9kBMOdQJOxBugI9gOv8dwjfai+/Azo8VSSnBO+w1U+rB/wCmICfMwfZ
q/OBRlV+4u5Fc2G49fG+PE0kcHXjxns1Rj2cck0Y7GADZKw/fnaNv3YGUaLjWRT52syNJi6XEQVX
1qogCI6n5gfW3Pd41jtdqqINpBO2NhRlD9ttYO8B6KuGbdMlUE0Y/6LeYiHcx9UpkQ9phiM7l841
tDYVCYXYptSm8pO/Pe07R57w9MjDa39V6YvkXoUAkRYJrtFiOWtLECtYeqJSdrv0KjOKZX2lb0yX
zMcpSuctLsyO0FNWgkDOzPSHPQLT/Hl8SmAGhwbXSFvSjWH+igBp/UyvptwY0dMOUOssGrNXAYl1
rrJhwMWHR8+kGyzGqvI9tcOwIeP3IDRIe3dmYrYizro/KRlo0DLrleTVLrRWu8em8GB/LvBAF+93
drQ4FbMq9sJr1WOnTcF0q9mT9XycY/n0mExQPrS6ntkmxUQPGX4zk+Wz6c1glct1sicIniWhe9fG
KIuH766D7BPjce4ZlY9w8vxWrMG4BivqcA1C5JAaq6meVD3JZfhaAShAoC4YlvKM3ofSwsleYXhH
wlJcrLaEUDQwqXa1IjBCe2G1WRMTVZpo9dBFWAMiHRti3hltyGjC4Mo2ZI5dn1f8WOtxaa2mZf9s
JVp53v3t5df0IHn2+CAJpvb5V7hDPSsTDrqscceJ7yShpCXLen8xFafQnQeFLIDl+4Fj+1OeZORd
knmKzE1c1T7op5U+WQkxk63y79kbV3H5mBYVGcKZdYgkEoUFKEA2o+W/UFadwlyziFe9cf1Y8+Xz
VSEryyOHSP9wyA1SIQqQBo6JG5cyeDqFxgJrsEiyXPmwi0c2gpSvWiOfqKr9O3VZ1qx/HRPmKsK5
PGWyFB9tSoYhjbkkCUi2oeY2fjPBhdWXp+VFcPtebPccwhk5UBQr7y9lGOzHgpPU2Xyq6Vhg3YDj
yDppwyaWj71XS5VxTXsrN+cfOkvkTfpi2TCojXINzeJld3p7I1i33gVPLG4yMVwMsgqDIkrL3O5H
pnENLV0qApEg9Wj4neuVGF9DdlY23Yo9vFKp+Jhbbrtbxq8N42Y6ZVSxhQU/5ETxwbTAPWKsViQj
WiI2u4ciH69UXnqQi7/Db6vi4tPDDUXcc+k+YjFxM9Pk8RoTPv30diDbpSHpiPffvtvqosVUa/RM
zfzcnbVBZ5SXyGJixLWQqXyalCJppjDzBwapWqZhw2dm1bnOQRsDwriFvDr+MYFOXFUEMY32I7RJ
iekZAimD8sKmm3eb1+e7oNEVnNvmPh2DEZ7YUR3eagGYp6h7SgWi6WjPdgUBR8RdeOc765CchCk0
3Ko/19wQbC1rPXXq9REU6ctdnVg/JZidsCX0cUkL+2zOZszWYmpSuUNU2Z2yFOtaYCgu6vGzxsb8
CptLPmTdp2rbusZeEubHKwfS3DQZe1ToSs1ZQNPPXwoT1eW7S6V1p07nTabA6rPvvWWUaXu7qTKV
Ng9KRcR6E1N7L0Lne0L2r3592D3MwwaHtsegzZ0Zxg47Zh/R8UD69FerFUHPQJ434ggopDE5kuLG
LjJhLIij7EKAQ9nXSyZRqZAF1VWDZ4NM31Gd8/IZFi+cwIgi/LBGynfve/g2zeMCNC7TYQDueb6Q
nPtdioSJBrZo61G2dOUu2lKnsfab1pu397VF1R7kF4UNioEKuzogfk6RR/JBmMVbZ+DOYESTMRC6
DFehDJbQVPuCuoqNrVGWLLkFqVcg6xf+ufrm8LDa5g567KSnro9ZE+1iCr/JOKjmsVfMEoR2HpWl
70MKQoANvDUSU6+0RY4TEHeycAusZ+DrC/Tn1zMhmx7P6aN98H7I9ocQHG+gy5dj0XTtrR9HYjsR
9k2pcLohIfKB1TNaTbXhCHrjMJJqLheyAkZbDNnfIY7VLf6vylZlOhldFUOTAqA2Ncu+ml/yYidG
AL1PPPQ8P44JabasauOINMqty74pwMaffm9CWUqSdBGIHAg6aoiJozFOs09hQdUintem8vT1BxqR
S0avl0+Gxlafj4HStyz3AkoSAt+XwB2mwn3Ih7sb2p1vCTMS6TUJXk+Aql7pLSWuXcZujMQ0iz0I
zdScLq+iDhtgpvM0W8xh1MNg/hje505tAnbO6KmUV6Lo4vaAou6KIeqvOngoYjVaiPhqF9xiqH1L
2vDp8lkICCgPyssHykwPoSFU5YE0zvt05m++jjqUrutdj+B9fC1OZlvaeqSk4eARSpsCJXTNSZUz
cFCqExIZT7ESgPgQJcpUe+NyCqE4R9ercVrY8gqTIiBFmaz9eXT1/2oHvgFGA9ZFbZwS4ipkoitt
iSYo1ftwzjuITMDMXqL1cenZKqLfEoyUWWz0q6LefbhM/Adpj4Vu9hWuie/KglqlOdFJRc/nxHh4
m+nS5m6ZVPkrNjVhvR/mTnK4SJh+cQEiIgSrLWYXTLRpqGv3aOUlw1WBHWg4kV6B8Vev1E6HH0K0
DQhdev20YSmQcAv/XJbHg5yma4/PTQKiYgmNTCxY33nIBSBxPHEqdkcE7JlQGHlCJMQpY8/8LohB
qTMy37TpeexCYXSXz+0bXYb7LmG/vCwXsSMaS1OGqM7eLxuJnppeGeWKgidQ+6o9G6ZAuLiUOPJF
HCFlQ1cg2bmhv1A8T7oO6jH8ilYG1AYBbOAEYQic0kUCEK2IB0v9d345pjl1ZI0TrMw6tYqKwEg4
j4hf++GM1epLCRp5QPA3q8iPAaKX6vvFyub8hDAQ7A0lUdGnR7Xamq/czhvFwSCmAgexV1j1Vwyx
ByOj/wtLMfcHA1Uv8WVGOPTxQrfQc5rO/rIWUeNGsn6w65LE2T24DFM0LmCbSkWo8tksL17ty8Hw
mR5Kwr8gvVeZnupPjDzgVKhwc74dsfCGdImIquN0u75YhYd+36h4Yf3AkET1eaFKUU4caHNyG0bO
BfrH5YagtiMdmRAx4HVBZmMzw/4YhON0S65PV0SiA5XDoWsEjb8e/tpZ41WbO5sT4dAxYSH9EfCQ
sO2ivke9+x2YOtZ1vslqvzeOvVEE5p5kopF0mvksEyYk+LwJoBqYDBexPHGY+yw6QPddaAXpoxB6
KcEcNzSAfK4dafYPv1MBG5X3SsEnIfW2Mhk36DpBui8ScprMoEg09CbzQJ3uECSkFGO+COnkXgca
PUpEb1mNKhQaxlRmaKLRiL3hkJ4UHl7/nl/I1HOVosBUvH+Zn40rQejsutX21BDZh35+HNkkeY0P
50p6IKQGC2vxoPPWc/tUdx63hPUguM0NKbwDmJc2ClXfrU0OskSmSAbE+b6AbHvzABLt+D/28IXG
oR7Y4wMM4Ziqyyi+oaraM+p0x9MRm1o3PgVNEwXdUeFvrbSFaNPKCzya7rjQ+/+hw0S25UosjnCh
P2Z//LKn9jH+/5Fnmh8czCExGJmN1cxY14QXTN8EVYTT3tHpfsgSc0YsmUTC5qIK+wC9WVUSE7UA
tiR/kcHYX3a+euTXIMdYz3ioV/xzFVL4ARIKxwWuSyRZrQmkLlutxm8ugPWSTS4P1UlnfOcLZnxd
3LsF41ls7dss4EalHq/FB7MJlLp+f1LE0dSsl30MGgMpencNi3Oc0iBbL588esilaFwEhC6TH4JJ
u0sp4hZM7H2mAOfsd2e71L5l9l64BuhcQ2HTxC3dFE0VfZAIcLjfsn9IC2XmlDiO6eKZO0i40B4D
VKrfLWL+/kEUqKdhN6ItMYScBbHhGzOVOf+QKdA+2JbrRNGdFurGzGIv4mnqsBVHMBrboIG9jqrq
URS5XVbaEQf+G10rkqW0tB5DBwY0fcdnJKesURMu5tB8IONmSvx4n6LeE9wwE/x8U+Uq50RIOSwe
UuFOjNQzy4TuhnNYKOJFcL0uczjdQpBLcGEGZ1FjYLo8Edqi1XeU2tLNdoOfhMt04WmQj7dSxREk
ON89DGuVIC/WQQ9+T1YRqKRSo4bbWsoXi6sYcsco2J4r03QJ5oyro7qwNO9BZBvH/X0Yd4HkVE9m
FlFVlwyvW1NZW2I7potfC01VtoHIRFDBL9FgSXilD1U3CJWSEc++dI0YKXjHSGugd9zIsHAvFNJ4
UZPRAT48UaFXpVr7Y96AWEIkSLgwy7JoqZaSocODs9rcfM+mJxltvnPc3VN06QvA5UJDiwWoyApD
+4I3YTfu5vQb+SZwKUTCdl3QJGGMzqa+F4BcSmOGJlmAeabX9AaPzGjPAqAdY/E3+V2spEBRN83L
5wW7+wv/y8/IuEyA/H2ALZ3o7wPuBdbH+mqVuy7Emh2y8tz9m5Pgrk+5/JVfA+fZeNMLs5EJZPhO
TS8Laakx1v77QPrDZOIxRqeKSmqpFsvyrYeNpugvziLYXCiqD6gHKCjLV2Sj/ouNSs+MskgCHpmF
0JEcEJdoEiLyPM+Uifk6A5+P8rzz3MdD3+5DMq6y8PjvqR64XXOoiFMZUkki2k9q9ypsEX3D/8zO
n4mDAmXTulWyvfT/IbMTPAjTdUfeiqipvH49LKjzjZox6ZRVi3Gt8NU61KwrL+Xbnb/LcmfZdE1q
kcklflvKszSoapISQwhcc5F4IPyOABNK8QvRaKK1m2HH3Dnvn0EXiliPgpcu3WgPUqvR9UIKne3B
YzYMKZ0FjTOFI9uI5jU/NIyMUbuBkd6H5o+28c6ldeP0iPoNoeyAcJpUYtqY+YqHHJZuKL9ZAHVt
pnwLCNBNaFoM1xf7bVYaambFGeOEls7UgcQ+UYxK1E3LQSa1HxqBxZZB127szzDUAoUTLGiitBWo
gl+QvoGX9QUlHyaLvjwD6hHWaQYnZ1KcSOJNUenPrX+/Y7QVtZjHie/X+Kb51soHXvXs+5HUDMBT
vlwEDxgZ2nZZ0u0x8pp0nQh1d2Hnv1OyZZdj+Auw9o3rgQPhKDGIIZhETIgw3CE5gyDk/Y+Rv/ZB
+43xvdTe+KQdSnoqovsnCQfuLGlQUvKoeasqCc1wPkL9Qo52jDCUDGZRNHwfBbAgvR6vMtPDMylp
VuI3TXmeULO1/JVwsM0r6cmefWI+RHPDnRYT9801tXfiXmkHH/E2kY9ZGDxnIo+ts2ep2MyIgIlC
6FNlYoZMrjlme+RqfMpxvm6AtlMOrKhXotEKg6cWkJAQeFCsVoKZTfFThjjMoxcBOA1XmJXskFlR
SBV6gTFUgUtpkGruG9HxmL42Ug5Jcoksgr2pkRKryAfpneBa4WsffElUmJbOGnvFWoRvoILIgJRc
vztikFStNHtC2dHj0UtEw7+IK4OpbKpwrVR73w3adZFBij+oUR/b1t+n5lkN2NKZdT1fE2qdcdeU
+ac6KiOzG7rbp9ZN2juRlFuDxPop1q91CSTh2mQHlpBjDCBqoxyWj1MdEXU+8eCp/HcQpYrdbMrK
kbI3Xwqm5+R3pJhhckzyeqXaMNcL4YhZcijCGy9LDIlkpXCTwF25516poURbBr/Q3HdzZ73TyMOo
CBEKceAWfBaOUDRxWSf3Vcz9leQMMc7wK7THi4TihbO6tf23pz6bj3muBTx0/LV7Ul9UZrfLnrRI
JRwy+v5zTFD1C8KBTQDHOuIe9zNv1tRnj4EMZZ5R0iYsE04zAO2WK8ywzqw9Szhqr4564ikUR0z3
VKJi262mUO/D7cXRrPXJPm4RYLjxDZznVDPS/8MrAIY5U/o8WI8yOYbq95a2z7aK3nUxK9i4aabV
jW109FRI2k4WyOPhG+ZzvtUXPweuKUxI1IG5tFjzI8FBvaCV/P+6ulUGN4Ln7u8Z4IMb42+3EZYn
b6oZpa38WBa09mBH4GJeRF1vUimeUfWAxlP+T73DRc5q5DqA+HIMQieo0f+5JCx86zs/JXehOJpY
k4sxNYRfjWM4ZzvIpx7V8QD2XdwZZjfv88NJ1cWqiXJD3V4JF+cDgiUPuKog42NJP8P/mPiiZ+HS
ysfK5mIolA9xZaCoQgJEqlsEzACRdq4IHrkuIgpYtfuj2veckqMdzxBFJ66MdPc7IfzGvaBjFGc0
Lfn/27WZjxKwv7pQcJBCLhWyeD4c7Z3KQxzKqREBYIZpMLGaJZ7xgjWZHq2s4CyeJatyP9JnYGEi
e6yzTn5dyzzivR4Cn9M4UR2Xpjj3E0PGneAamr7/bv6Qhf6ZEt8n3gPZKrCEyJpWmq/nWP8n2NXQ
nSZRVjbACUN30EDtf9jxya/eMHHfpLP1YAWYBhG98yp53CgGvPHVVGVZR8+lMtfZjZNcQbjnTr3v
aP/aHRfPzAsuI5jd1qvrIfGqHLVtqLJvCFbq+7mAeNxwhpmme93W+a6lI4/4TN/qJYTb1Mk5rdWd
e0cLfAssb1kacAc6R/cmCKSHT8Wz7sNBByDkdgHOXy5IUNJDoNohZlH7Rn18V1cqR2qTIAly+J6f
UWNm5nWF+adom0hxhPgYoIheNtFhjYJJfDpRrcMfj8tl+evKOAt70unKGRmkcSlzjRIa8MLkso5o
nqN9LUZJCtLkyS7SiE3V7AJayI8dVu43n7R+q6HKwPuKicCd6VbGqA3HYVDFgt4KkQ2yWSRLiVCx
GVPHfDF6c6ORdKX+wolDklO9rGb5ffjfSS50TWFVuT1wrAxo7wBBToOY90nHrC/KatQr8UOKVoX6
u91DtFSFQIJCILwvSewwUvQVXm7ZWc78vDSQOoyTZgUmrSI0KVHWA9PSoh2ai3c/DlLV8rSBMjaf
ShrZRB09kbxBlMjgWgVF2Q+sp/1n76YMLZUgvAzJ43JR8NVyPmKmznhK+6JKwT1IKYCKECIH1kF9
aLrsDTEfBW9QZ263fpGbtZnmNmyCjDioIGgmKJEtGGX3/8iXYMsdkPivYZb+tCKKn3EKc3CZbbF5
97usr103Mv1G9C4bDNmxT3gNJOLNBIn4hHwIVv3+v+yx54JZftnlVrp4rjDmFCgR0NTnDMhI8Qf1
HhV35oaCE/rLg5JCqZvwlSe17SQVPrdnHzTUEtatCjDJt4Hmg8IsxJjr7kJwKoD1Wc/ceRfoAjRR
Bdi4JSByRGDLAInkjJJUWOKRWdEzckCNoeAwN244Px7jHozo+HYdo3ss8ODHnF6pit3XoXTGvCX+
ViEHc8AQ9qwdRR/Yxzg6PjW4zTWDQ4VGyuDwCWU5i2n2XW23qcUzoFksQ8FuSnaIjHu7tifppyKO
9V6j0TAL6FT8hep9Mukz3jUXdPYAf/mHjKXy4RWVAAFol5CrefQQwCRjtKIV734rgf8xElIo8Zke
LDbwM809DEg7faWxUifnvjrarwJVj3lB1rlIV/3Lvpa2umrCvdz9+qFaY1zwsXKnt8h3n1A5a80m
dhUBCg9d7qkokOFIq/0UQMRhe8Zu3N7XmPx3vJHvXdjo4RHSMy53XrH3EufkKhdVdeSd5Xk/10dt
B0YgX4VRvsMV08nQnGODyoot7tIIp/6+NYiQ9JRm3Ch7i+FoaN1x1/rePfEqF7MvDWKnX1FNeiQH
NmkJnjjzoJ6o0w5iUu7NYOgOxarR7/+Ffn2BgJV2K28NeDWQ4HB+9WGCJzusni4pdeP50PCWBRge
53Eqm5A5nM6MmF/bfk2GVbWEMNdlw9Dr89ALyIp+/8m1HEC+oPmAVLjntSeJ/6wtbw6wLr+t3LZS
SzK1hKwsqCITUvRHd7G2+4cL3rJ21yFVf3AH5Efaq/wBlUbcA2yE1IOEn0u040ITBgeoAqKxQ+Le
ogsy5Fflz83RCn9lb906OFnKHwzjZxy6PpaFWWIweh0235kHUz1ADJxwveWyyizQuof1uefUXsQw
qKgNR5h3xwmURD70oP3NfmKKvAQigTts443xL8zPQlfFM73Oven+LKjjz3/AHMKl1Mi/V24dcqRh
dYu9U9Bt/cHQV8folnv8vBxYMoPl1zqwClGCSzKyjgKn1YNIMN9HNO5NlszBQJe6dKfcxHnA7F+2
gsZ4w+DgYzEu4ywmOsCuVy1gR9dE4dkNNOYh2qxKy82H9rmyZPH7uwypgFIt0A2x5zHRvWvNxDzm
6bKAsz0q8kxVi1pycxx+llCkEVZtAskrb3/DXVqZHyJz9ONluLaaB3ENjx7EpXULvV7Rw8vUpASv
BzVe0QV9f+WYRSjjuczb1UKsgQkLddqkHMZgUdL024P4ge+yx2tx9sruBTcVxn3T1XRqpNWABUme
saiuGXKK7KfmY5dydRcb7vLHsEqJivxCCqr+Ms29Ns32VBD3rmqn3a9HaXjg+XDVFtGPS7bwO0fu
l2hXtbXhdLei8zrKYdzx+/8/RcflGZvBlG3kslI4ALhNk5qMOvSx2vK/EmbhJ5RvBekyzO+QAI9t
OhmJHNoyEH1oX2lFEvVPSTaEF4N+9/DXYyhr9Hg1SDqlRJfQJiv6+wx4WpYWD5KbECs6nNKavr6x
KVeHoUG4hvFluUttDc3KYl5Iopu4t3y3PS3d3nfZDVwO92GNh4EyFq9F2p7G1EndwDdiS1BVIkDx
NMHswxRoZ8NVKC04BBEajdv9MTc6qDoHhEdshm7bVUFlRoCuKSLPI0N0mrLahzjjfrA6WSfExXGy
Q83MS5Vy/4lWf67zUtiBryIzMim4ix76GkeN3Z+LnyIiIh9STC/L2I/OIbtas5dmUQT1E4wvFII4
XyYxE/RNtznBmZQWT3kvgKuJP2LFdt0sEfg7abd20WoVRBKs1BZEvvtTwwT2PWeht0YdGE38ddqz
FelHLl3SsjZex+75Pcyo9pbWN8XtoNMpru/+zw6amIaTWM8Rlz1D/0uEKpqUqCXr7PXxMdgEi9PD
M7GBBYjmB+aRtD23Q0HwpjM+qbRGIJvJ0w6dvqaKQK6LkcJi4VQQ4ZnERaQsNA9FmnBP2FTWF1l8
nn/VWZl+i0FUiEz5TFAPVIhs8l4fuuu68Fi4WLAF4/MWYmMndmmIUYxWybTCqhgGTqPBx3RL5tZX
5Q4oDum4QvXC7WG30vIH0RAGxMuMA9CvHjcuusNx3ZjxCIeWX8QKGwZzARojOCc0tpT4y8GwTmKQ
o5v/S0YyP7msA6hkUKb1BJ78Fl17spIULhSxBywytpS/s8d6uzAXMEa2noMbgcOhLjy8jFDBevwC
PZoo6EneX9GbB/eyNItobarhU/0kcBJo3Kqn9qp2fZY2QKI3/YjloBE9d9a1zzabBpBUaDSs6p3q
FAaQnEI0MEMlub5Q0WAVSEIyz1J69GRK/QT9pTKzeR2F5zVpRwX9KpHFzJVFfpxEXGQeyPyzXqH7
cyxXfQx8Ukht+VHXKso76cHnLylN9Uz8hUMMae9USQXDCxs5UARMwY/EWTAl07+MKSiRugb11LbN
nu5DNTe82RFf5ljB6ITwCfHJ2RmpkueRARUQ6RL6DNCX9dXghtFuap4UblUxyfiNVHG04fal+1ZU
pCJWzqJ6bBe2kCq58PO3v/zelBU+TLw6lmAJVl6NZgspD6DjE24uJzFrL0dQi4a3S/bKvL3CO1pn
+lapZonBNmuHasIN0E/dr8VpGaQ0GDeFRYqeD4oLxlCrLH6aZ9a58HXmRKYr1bkl212JTltDJ/Q7
DaXnIX6rF+gl2jwlZe8G7r67dhHmhhL65nmm2pkeZ8CmN/uUPWnRkX94MyfaKshXUGlCvHYWV8VY
YqyzJztZ2RlQ15gKY1xthu7dv1JJf60+iSStxJAViTcTgomFIOqvO6YrMmgiRZG+zitnhAMjUsa6
Xm85OUBHbJYu1pigYm6AnpytfwLAyQJMdQNEDDDsX6AH6x00+UKJPXmBgaPpjd0LklCgykYrxS79
eOtUDmQp8YuDLFj+oL3thAg9vnFx0NyenrHCIk5t88g+P9r/6gah0pzr20k0avxnFu/X4BBkIlEY
EyuXxDG5c39U7sJg8zS35/27NueCAg0cBku+qa6xuzXHJNM0MmuvMomujs04R10UNpOyah0Uuz7h
XqN3uLhIyyfLvXq29yDMdd2ypqGoekWvbldu9Ws4IKcgLZkGUChGGwiOjVeAEb6mSh3XYVDYaE6S
KQ9DEFCJzG6vY/qB84obX5xTJLtELO0evhTkUQ+WJmv1MHcYlIyct72YPi5Mklvx7mbOlpfLveZl
hqWGTNwbonqlxv+BGzZFPsmg0e8lfxqOWqifHWOGfJVr4lgJtOyXJnwSHjVjUSp+JG7GIDvbCtsw
z2r2ZVxSjkGQZjaIZ+8mV6d26ngkRai8uVyI0Vfqj8wqun1NsP2+PbirFx3EO8QlO3t85uaq7Y53
cyzvR97uBXQpdD3Ijd0GrDO5WdCPDKmKf1QkKiYSOcCd+ikd7FX8RPxdB8xtOwI6sMQANEHhyq3d
4i2ny7pa4he48fRUUQ+h5nRxvoEED03PuaJ/vid3lOxWvw/QatD7ZLPytOfSW338hHyahFgIinqT
OJyvMf4C7sFK2MQPTzhsU4D/RdsFbDMaeZ2owKgN4H2AWqYaGM+YQwnE11J9/0TO/zgpBMOyAmCh
KGLZGY7F22xcVsJuyoylBLunWDDkn3m2ieVCIgnyyrxJpBh4QsugeGiYgp/P10xkydrKsUYyTRbS
1uOuIRaQiLWomEY1+LUQVlpu0A1zCs6gzKF5Qe+n+jSLZw3sUhB+lCo+raAtbsv4Rb3fP+0aH2td
SMGtaDz4P3DAxun6w/PMB6vabZODWHzvvegF+F4StH6RmomYRZZRks1u9umM4cKdF1ZGZQN2eHBO
w1wdSBqELNvlh8IUx5NnBUoTlpq27LQijH8NTVR6nS7RgDjW7SUw3/QGUZ0qVO/IHClKZhsit0UY
ePQdAtx6kU6k4l4tPZ7SEGO426mkwiU20+fxcr+cdDPzZ9pXgOD/TlsHBjbqHdk56/q1lAZzwT6q
y3XMrbkO+wg3LE+Kcp5tSxfEdGhCTFKar171ENZNLcRrL9JAQNJ7Bndw8nDh2trLH56Hv0DkQnmk
yodPjg2KRQ5XhGEaZWFpbD4LRHZ7dfOlTEJwgd6W+j7MnpxmZ7YZ94htMqHPm/UCGBUOaWgkTo/f
8KlUN7QWjJ/aQsva1CMFr8U1Y1Gn1tYhBl5M7kLSII2xE2EJRxITfQEr2r4NbQYlULeB+dndIXFD
zzG68wkdKJAx8Ei/fUD/UlW24G0CEb+juNsDVuTq7t3V1MGR5yTAGvXqAABCN45PS/kWcXt9Mkdy
gXi9kbOSXsMmtNgO8fTxVpWnd7HbBVDgjbFdP/p6g/UuZRsJ1XU5Jl+VTDgD9EOG7BB2dt4pkMFz
PmhUdXrnQJScOLFhtfSIOk/TFkyVY+SEsKBD0ZMKIKVZiTBzMI8hwSS80IXAJcTnJCVLrPrESYqe
jsJp5KueUWoO0hjT0gDvNmJyulOyXd+1bEIq+SBShRJlHnDyqERdPgW1utzVDUPYmqaixsrry9TL
zJWQINdEMASlSqyd4QIlpYtUS9Y8SJxTnECxiocDrJznuPoBg2w5Fh+wBo1a8d0GJrn2ZZgoHqc6
zYxy10KYXQI64+97TS86f3hOqBq6wqbLxi0fnAqNFNklm0r0NMKHPg6475YQSqjwV26jbcHQhRpw
+Sc2z//tP6VLZHsXGZpij2dmVtL2BA/pDiFBAZH8WRBHh6VHQxWUnPb2zgSKU7m0JZMsrtLMY1A4
kY5lIPF/ZfUjtI4pz1kzmXvADnYFdoOCUxxEK1y4uPf0mkfJVVTtNOPxhL3KrHq5jFzsQfv6C6kl
KEr04mFYPRIGL7LWa7pHei/QR+T9hMCvBl/XO6nwM2S4UHGqBvDp+WGKC1cmWphUWfTn2EUEgGfK
SpkJY2wwPZFsK200LGrWVJdunV+kc9Sogrv6Os9rneM119ChdtWMHxPGzOlg3nhA847c37GlBMb2
9MgIdcv3NLts3FpRbdGKAzoWKUao5UqlfTmzjS6TRwQgZyzF6R24MTbvDY/8dfBA8vxYYOOrVJj+
lggM2AVWt0jWsultXO3SWlPYADvhDkTql7X9PWYhWuzi4RXmotTzWkWNKiMk3d8IK95rLArYlVIL
h1K0hPq/ZIRXlfZSxFxMkM1aA6KyAmGDC3LQ95joG1lEOXzCr+0r+ME8l6FMoC9Db3AGPD015Wjd
WhQLS3k+xpGlLwcDdaKdh95elLHhxCd7+36yNbwK0sgmkLm2wj5DOPkPKN+cV4KbQGkLRsGdstmU
WYyDkH5lDY0deF7y2lWoI6NcUIPKu+Wp9fp0jXFOaS1i5ZYMQMUe9vcNNlvC7TWhGBLeP8H3W0pP
nY1SC7E/5jdtvIELR+yFsNr5/9PQie8vzuweMoGldEUh9VAeJE6PyjyVmBakhovx01yhI8yZeoRb
pRuLshWrBfPm67zc//oP4sbSMNA018WhvWw7WeUk+7j9Dt19FLdojxiBQdfdr7jPVUWcXPfqqFuK
u/HvCkhbinfKpTdv/01K4q5Yj7617TMz/yVi51qSSUtynyODRrAGlWpeJXX5y1gogE6zB4HL8t3w
+3/68gu8SK5MbHhl1x7MEiU7C0P64N6P92v1yRm6V6mKrlHw+gXnt0ZB0qXM51FgkZimmf666R9v
3Rd3qBJ12Bue3OWSvjs0KQo30s25l5QhGvOd9H/JqPkJ2gi/8NjMWJ91YyfAh0vu3es+qeQAHkhK
JeYCceew//AF/QJi5vuE7hHpYLqurXeAOS0MPbY0qVWwsECF/SeOA3LmlJECp+FEouF92xz7TZIW
xe6585QWzVg6wsyYFtJLmlWKklmOrVkgNDuUHRsywSpDo5rBxgbqIpZ0NxCSinCyZ6FW6n7mU712
2Y23TZJoqWww2nnDSQG0lcNje4FmFfTWRPqx1a9o7ryCC1yEEg+796rNp+RizH4jroa5fnLmNZRh
xZamhWkEuHCleTs96PGb3u1oT8NdjWUsRMfMBOgbKCj/XUnaCPelp6Y64ayR8tqx+iwJQsU+C5pK
ijxwDflUU8hZvm+gZj4m4DKzwWdcMNZK3lBBSaBgIHvG2z/8lbj3AgxPRvLpTV5E1vWLu3NpoYrw
FkvXJVJBmojOkrSkrrMc4B3A6dHEGuycDF0t0sa8oRJfugxD4et5/9ft+CEBlog5eQOrEA5ncLvP
hxwTD7OIlCgHGYbNa1rCVKUgMuH5oaYu0KygtaycDTT6h84xh+j+RFFb0vK9pkj7NgjCZkyktD+v
pKsyk8PAWHIiYp16b+utxr28tH11vrezd5qCkLXmfjzYp4LbN8VSSsJELTaUFu+NEL83uclFlujI
Lvmn4d62556FcLj92c+bbllYyty2BBUf+sLTbg+pzFIhzz18G3ihc8XdUyjjP92xrbatSzvvHseZ
/3W0X0hSXEUdegliBL54Pb6DJhKk0j5F3DBl2ZiqGEpDyUJAWpOTqvT+xOEEaUl+lNhih6/UMvKH
4Ca9229BkgfUQd4cRLguQY2ItUUEBkI5wlNKZ9FjGOaIP9bhGZguWDwpSIBDvwa9rzuP6qzfb02R
G6cGlsVEhAEtEdg8/IA45Hx93v3D/PamdQ3oAFtIt7PHkJNDn5tEieQ90tLztTpDUepsb3l7ts5C
dmqBIK5f3qs8NPYJSt3il42JMlV8hbG8eBoNOlEmn2pMernUVIo0BNJnsiFNHTWiSYauGZDkLKxq
s6DxI2u13IdJj+p8L3E/oJFwhXl1MdtFznBZLYdXrKte3eTWtVp5p31YrD+b07RuXdiHiKqByzsp
4yUl8Tau8l5zEG1ZYwow1qI5zTbiA2YjbPAoPEOS/ZId9QgjAwfaEnc86pBITKYGZ9CV4a97ggzp
SED2ZR7T+F75rLeSvs2EifWS411aOhNAA2af7wnnAFg+qLyb0kZyJwmKtLHXrulZgmDHeUZYEQvP
U6cUH864ASo4zKnInu/gUbNti4lcWPOkN2gXrt5RL5ztYM46oQD+TVw7EzZDbfmMcDShojsbIh/m
+HoAym3XCf8vo/T6fDIUPrwHtx0EbPqHhY9+56jZURJtHR3pCjatTETN+MZWoSM0zVMHDy/sRc4X
I40U98eZWABiD6ybS0ieSMj5/Q4pejiB9IusKtucTDszuf8ASV9nKGYGX9Dqw1BShxVgf3SegA/v
mchAPIHywoVUzLD1GYyrI2OE/wV1gCYTXNvqFTvwPt+PDa0+QAjfrgvGRxwTGkuM984JtLpjBhZR
c2dQI2zJLxbmNENZhAgI2HetaQI/gRud++Hws15TZl2XyPcZAsYPov9L8MtY90Fv+FMD8j8YwNIh
9Wcu2fUBSCnyFK1BT6DrQ40eASN3+PI5zutGHYSThBP2E46va7rsXig+ClN2WGm0EuT31KXSwGVD
Sy3Y4foRu/6Os0b0nyJnBWHZIxc4HqtpKYRc4uhOuRMmoszEF8yqRCL7+MR6lArRoNCPczAvkGpv
kr3AHoCNp7UozHHMnLGI39NmQvUbzpOZJK6bzN3SppIsPzsht/Jv2t39+oVP1GZDyX0JRQGWFim8
PqLuyiG/RYejbRG0KGuZ3GUGbkQorehwamqhOiE4sybejxvFUUz+zZ4rzMnEpxJTf/JoTQ0765DG
nQRMR2hI/TsGcU3oIVDKTj7zrP3O06lGZOgrPPK2XRiuLxPBKLSr3utmd2YaOZq98c8/MVuQkb5l
oBD3MZz6tXKKDmweVWVAf5ZeyBaWMQHTqiQeB8+8Qf6fut7WR2A5SzsjUtLVBEytp8UhRRPU2EEj
UnmUSbljIhGmLemx58y0qtJS/tB3Px6Lq/QbQ5eCBylIQU0NpcXzkF01VL6kzuVy9k87xAA7nYvO
S3J2sL9ldl69i3AkLhQZOLlszSCojLCcTwXTDP/YtaEYd0EnTVW+zqHC92K3ZPvAbefKrtjXx3yI
YVYOPkTkhxHY5S6TZ7Y13AMzZ9E7PzwTEiGv1kmsZ1HtTCZjiiwiwyDsiAasF85KBSaBGj6c8Xkp
zWaGD1fzvuJ8oGyrdwpHSel8qBsMSVk6OJQX5IV6nhIIIJeH8BzmJ4jaUStHFApkxJQHl5obX4vm
jMB+WgoVjikAM0PS6CuIpxciS7B8Uwc6UQotA7y9biAnkMY9he9G6BIevPtaiz92+Hp24fFh1hDj
63RFvWFUBUjBSGovElWwlVDY67DSmwlnAdojiybHgwxjtJKjqLN5lKPlyhG+U2oz1/NMmwjuWKf0
JLDmTwm+XFTWaAFe7XtLgnrYt2jI7bzLi17+kGtRxv6NxFp3n1xfPFcDDga/8IPEe430y1G5redv
Q5TGtFzijMwUb8OiZQaxNaKbZCnc61OhgXWp0fJCgwOQ5geKEDvEm8+mEWVRuUjREvmlZP52MVtB
PrRjG8ePHMKniWP92v6y/SVJBqeMUO6XY7xdN7V3DTqiI6rMokJ/UossfiRRkafBI+Vdtnq+IpYo
gngvci0It7bLvfvDdFpZq+kue0ba1jzbS5s4CA14xhW4CPhuXSPPax7QW1LTMMBRyx5VlATXfyxv
XuVKkKUw+xJ2jU5XIxM3HLt5qsHO+8vAsT5G4beU9t97AvAOEBKTyhuxII7qcU9aXCt3bLn0+HEP
bsPFiFznQzd9AYe3SDYPDviPOFdV9tuWGX7Fy1XjEpELt34UDXza4DUUQ0/XbqE3S1+yDQptOU6W
l48DJCNKKWPpMrGw8aqAWpHTSGUlYOPiRGVIkVyYfja7/CBFy/iSwnuI2EzNFUIeiWe230XvKB7+
uHLQjNSqheWgN+6RWAHBH7ppzFr5Wfz2yzIlly1CuZi0Zx7m/6b2K72LSclN6BXilsC+0Ymi66ah
RmjtIscacnSWfY1z1shXGdP9zTAdLVZ7NwepFRKNuETICZccbAJ5A7VMI8mz/zxZFVqxCrp+n4jw
hG7qIXkmKP8dk91gfbyoNDte0aSOW6D1ADkzPfIzOvYNNr6pAcPTJN1PpaFCc6IOEC0CPxrg0Rdp
Sduwoih66Fmayl6rMzPrYTOgnjOwDWRcR4JqLp4YIDrmxwPpxpMBPzBMdtITf9N5J0gbiH3hp8V1
b6WmKoDVnjoweA8TvomS3r/GqjWUois7jqrQ90QY5yGtH3ITk20VCB0j75oY35S0jtU3i6Guf4Xx
0sqoph24zdx51r5shTBYgByaI4qXIQP6LgCpD2TRQVxEtFTTZm9OvhABZPln1qJb1IXuZX5OSfgS
7Pgvvn0XBRTXTVWV1Lq60ErbvkTMAyGcpC+SyVeGqBRXnEW7jjr3SKYJYxUbDqeHER4OA+pHouWt
1vCtoY5x0w1qcC85LO+A4+yFPvkphffT2ZG2eJjODX5RQUxZPuCgInD7kky9bCH9JxVGQDSofK0t
kS2Lh9xtTJh823BZOukr/XBuBTp+srOvrmkak1+Re7E5cOTMXdhKWp7/TBCDCvy2f6s6iZ16u6Dw
S8fWt1Dg4GlV/+hDegscoZ+VfIC7PIADHgnzndTDX5VCJcgM/SXy/PFRr+jtjsN9gHOnYAxYdSVP
x+v4eWNLTz73s9ATB/06Dj2dzBlPLIMB5/9mJPRT85L57irsPdpeksKm/SP2KkCl759EpBtro8QO
s9MGisek3e71Q6Hmvb6/8zTMV2fWrMY/mmsCWQhEo0dgFff0m+zsOsXZ+QWmDA+arZEqLllyuaGc
gKsOMyCSS2mJWiPLYGjQa2cOabf+AG3TNDsuxl5UTczPbFfnkRnJ0ri+8sVoUlpb2M+NvT8HCGPH
jN/90nDpGxq+6t30rg2gQpVMxmXi23FnaFbL+o37TrN2dXk0ACiuzDO+MvmVr0Q1yAfkZChQ9uLm
cs9sf9KhLC37xUN+4a+sAomtkpTpTuygGJ+F7DqYRQ3y4kXv2N+Ftao5Hln8iZt4sxFl53s+MaGd
DwQSD3JtQX/1K8Upiai6GAmEI56hTVw5e/2z0xLTb6EV00BJdo8EkIvrfB7pDJKcm0KGvnptp2Jf
xDbQ7CA4hKMQvok4/SfMze/JF14N4koO/0PQzIOEfXsydFebAbG0epGGOI9ingceiM5nimDgLnrg
jfniRDHpV2hCQg9iWJU8hpALMPkyOsJtSQTbcFJ6n0LC2IoW/U0j5OtFblQ+asOA28m99rKXQmPu
l3W6bCoL4PzF/AXh2rBMizzV57sHHRR/6ZL5dC/cKoUpOoDLaK5W8ljKHlbVQoKAQI8+iMe3CD5f
yLSzWbanBSvK2S7rP070ibcPiMfU+FRout7qGgqA1wztl5Lub4n5LBp9e6feIgk6/POx7bXo/Obq
vk/5EOSM9He3UBH6UIGJpEfuTjq6ITyDvbWzhCagXGGJEwMnSwY0y+J4M0aP1AtMGB5HKNlMhhcO
y2AXXcUN8EUxg9MV/9zpTT09il6xvtFKcQF04rca7vkv2mKTt7tLXOgfanicCWE/6bOrR2/xPGVw
QN9NvO4FYyr3cRXTQ13/j3cxThjPDN01aJlfn1GtmwZme1T8dgrl8HSosI+MyHZ0/+5D3kxQpkJl
+C+tkJWylfNocG2+K/U8Qh6e2o2Ups2Td5+ewst+BZ7DsiLnc9b9n1RpaCN8ZpSMOQQQut7qhGdw
hmVbnahDH88fWxvlIvrPgqhMm4S3gcpK/2DmFxxQrPSVexGdZCsNKlUXt9pneUvdMbCT1mZXf93N
YX2hMRvsxPWDHziLJtIvsdWfdj5uFsDHb7HWe0auyC2GnEKMtQW+gKIrZtT9/G4IPDAt/35KQXL9
LzL3FtujHDMMlQRSZ9iIVpFitcSBAVhhSEPP1iNVX8dcQ1MbnO1f2/ctPB7P2By1GcwkMAPg90OU
+X+TCfcQuSVd+Fa+wimdyRMkoAyOi9fwu658r/EaxzX8A/9hsObKtTIzGo6UBf1hQOVoUoK8Aegp
SZCMzpA6KJiHyjz/VOXumoP/OTc8SexpOI2NbolxaT4f0vA8afbau9w7VqWRDFapyO7UdegEc7b6
FrFM29WSEtSiiZ3Srfcmgu0ynsDymfgcphiT26JLfi6wWWyEvvE9/IgXff95o7wWgUz1SatvRx44
IRI1ZwIDmC/ewj6aWWaNAVl3GWyT16HHcT8a+o/RbdP0o22Lvh+2X44bt3R5Rz04uhuXZe+fqpiI
8OzpG/GQejubDnwpk7j/ckfdkWekfH7NfF5Unen2M007nSLTx0F6aPcXAGfLBVrRB4Mj/eJ0VPGN
zbeowjU2m+PyzpOpOchzrHRn8G6dndQoRZS4jPouD4eGxVjRUg5I0TT+4OYuym+5mCutnMK4uAnR
pQSI9IZq+RtlvSIEPRzC2vf+chXDb+JqP+mzrStMrho75V3jzp2rKJkzRQUdGSS4yuEhQ+ZprnWg
Rf+CkrYMnEvxI7xcl20E/uz5W9ZiJhKA5EvSoNXpEzFpSAgNUQc6KQJy/ntrssJTC9Nxm+vETpsR
/28IxHqOzpw3zIecunlw+ohh0wjzqbz0haIvmbLgzSFJeJ3WnAJeRiZYX6VI55AIzGgEDAe1fcpK
vpGsjAJ96qPg6mk3GcEvF/RB2/n2AoqBGN7KCnBXXaBb5d5F5ilLsaPd7zGA0q2Ds3xH7pD5rIm4
aFxptpoo028BAphHU2+9mBJ3J9QEoC++PDcE096sKlVXUXlqZewy4udAEQQzTk31FX3D1weYv9Kl
RFCA24rE5qbmKD0We+qalBOJVn5lJY/OBhPLiBQFSbu+is2owo17ErDdX99Z6HSFerCCmSyrQxif
2Na018gQecg3AkssRqHeoBLbfrvw9PC6aECT2JJkljqr75xBZtJ5NOCVSM+/UgwIFTFTtcy2CiCN
e+cSORRpljw9JeC3THN5eIipNhVXpQLHhXfODtm9OaLN8A9PbewIno2jB2OvSWvr13IzzxFfIhjW
+BwdX2mHj8WN2eSvC2bKDHJ/B7xJHILYYeW+imN9rSsbJ08T/jcqhEHeO9r4G3IvbhvUA1/nWv7E
hBR2b8IExX3fgBARNkxC/6Ou3GpPbOMZsTM83Ov7PB0QI+fjQDKYXwgLS+cC/hiY/W48tpv2USjT
K3+b+pwCW4CacEGJctIGJAsL5VLnvSK++4FGzt9is0YGnXPdBLlirsbLuacJLwymeORraXMWyRvx
vPx+ioLSg5V30y/0deVibeqF+RpVHp5i1TenBkVSWgNpAwMHFmWtNEs2mEBp38R3Dxr4JYv0Rzoy
D4W6H5yGZXyTMaR0Ns2O3lPcOzcwY8bfbFHuCuy+M39xpDE4VKJ45CuFgMtSHiCYLAaYjkO4KrE6
MiUA+CIwxO4GyY1Jt2DP0ZYx28PWGUZMT9C74bKNZHpRSj8zy9a9BizazMxovz1o37bKqrqjnBhk
qeYaYLh9goMuAy4Dzj00GXRMkS5WqyWxwyz/19jkJ5PFG/VvIXzUvlRlFSUCu3My3DAD+JOw6cFr
2GvA70S9Qt6ApH/myW9EYlganIvGneXwUofu9aQqpp4Mejfg4R40J9QsyBtZUd9lQwztj8XLyrBz
D8uqgKTzxjTCLW9fd28rI1WiBicEi8E5TZcBY31/YC8O1ZZcEw9Qyd2TuLJmx19TjgN/b8m3odXY
fVDXMN4PEpkqHScuMyT7AU692e1lpe+QiRMIfzNwUwGvzN/htLW4qBtVY1PvZ+bnldNgIgNRaYh5
tnsuJdwNAsxlYD3Kp/bXAk25mU6X5JNH+f3FT1wyAdtnhLezfTulv2hLIBl/FG1wEMY6e5I3JYXT
m2biaMbXsLUyd2T4T2g/eqonhKJbjedkcxYAz7i+D+yjA9tJAtsRLmTUrFHDreS3TAJ8UY2tzWGL
yHqUevXxAYGQmPUcoSAO6Lgh4aQeNQlab+QcTOHBE/2BH918EufGjPsyuYP3cr7WHOsRXp64UtUd
47dd6ARIzWg7YmGX4fwkHJgroV1cszN29W++Bov92YHf9CnWzfxqptVFRA1XeL5a8AU26PH44For
Ikh7a3yS0h5la1ZntXdbYAfAOFEqAeUH/prfqFZSOY8dOGrpn0wQ/WHh0vTpgO23K7uYfDiiejsM
tDxbA19QayPGIajEA2+cmvJOL04KYe0zPhtJrKGxhV9oHC3u9GyLbTQ0xeond/E6cCMe0052xIwS
GfE8GQ10nhFtTczwJ+h+dQlCyGVftBsiaZslq/OpmweCKn29Zcg7JeuUdrUzX60ID2lDzwwOZTQ3
2KrUHpkisMikYPefplOt5C0n5pWHEpWMmcuD06AqlEk4e8Ui1ctHX5peXupwUX6T6886UJMjdRGa
QHD4fPhN+2Ep7pbk2PGQwBz+yD06HitWLo3eLaOZ3dIHkNIaQnqJyOScX3ZDsBDtcnjOj6ptOPe1
xP4xdUkNxleXU5R6At2sxQG8gdnaMN8/wX1ZJc5P0X2IQXWavqY+dctPswOZtQjF0ZBGLpFRjyfH
fQIhlg6A3qcIe27MDrdsYxRIg8gszMNW7rqbKjwR7qJ1pfzQze4xADTuaJkR5iwA5tNd8tKOasbc
gh0pJGe9OL46XWUkskdKn5uEnFOeAJGXdtR7nHppnphclnxMzYAp/KwltIaudUMbQCp6EQ/yO2Xr
KzPZNNbDQT5GIF9kD+3yiROtY2Q1OVl4U2Oq4FucsMvWO+w8whU+5x8O3nb0S5eBNkPpVe8ThcJe
jP5RxMmRWhDdGlu4KMbpmBEiI9eMbCvcaY6lazijkBOMhVccnjblXKjeyP3Ova5aqL/nkC3gl1N5
/7TBqZKBsdeabiRtH0SI2cmYv7IhfeKuDpQ07EHht8X++88BpLat1LQ1SGCNNhckkqqCBLC3a0Ry
xtLKmfGYz9J1F0nNdM9iVRhhZ2tn42Wpz459+jmTsoaeMp7uWvLi3YH2SooRqKEz5UDtHipNz785
QnSKwGrUSRNKpgMfnpGAEKPjlvyihXCv6nl0/uMy6R+M+lwU8/JGPDc8ySxti8usOp9ndOw5E/yQ
UTK3OwrbL0AVZ2pQMgThACOUxGnoCRGsw9CHe73LTdpc6WvNN2zOYnihhrzt7k2ue7SFIO8MwQWk
CDsLFpg3ZzRNvIAHBIeyLZYgJhW+lGItAy/8YWGlj3wZYE8rz8b9mOH/f34ESnH1nviLmZuBmKvc
xQAmAyJOvS/6JhFglpBS2UIyCSiniSXdem8/A46lq0P9MeL91qOpx2utfAVLBcZsHl1/WsCObB+R
8MpQk6oBZvT7tUUOXXZ124hMS0qksV2LjpZnLQZIllHlTzOjzENSHfgGRJSIum9uezi1BqKfrtBq
UgaFmW8ytsEodP7NGooL++e8Ir9/2F9TQ84gPQprBM1wCdk57kvQv7ud6xu4Wc/GD3d1bDX3XOOQ
Q0hEpNhSdiQ2jDUm0wPQBdpoAww585UlZl7ZIDs1oAZqC0Su4NGGmfDa3fPB1LwOQ+xS/fOWETG8
e4ZrFrNvVUnkxyeOc/jpCvLQGUcZp22oHTQiPCmda9VMGvWFNX9RvpJY3DbDz4tHvIXU7W0EwM4G
/EnZ/qnGfqFbVNHx9nPCZjeB+ccnUiWAVCVYTKMfEdE6uy3d0nKyo8gDfugifvcG5By3VPbrO35O
8DkLKqsqAKrde8bwMpTAIav5ES6AKDBRkcPiUTbSA8B2riuMPQmKbd6qih3EJ+Q5BQCbk7A2L+sD
3EF9dgrs4UG4RyaTmdRt1TCWeKp/rlznfaKcoehoDkkQv9KNUmXKiJU3Gc5PePpd1uwyVnUFass1
0MCTwqTyf91iLAzvWsRk80h9iUugv6xKpib5WKK4FWd/yInExNeG16BVtvfSQZQeBUeHZQ5sI5BI
oLB5EXENzE+cjR3W5ozYRghtI9/f8NgR2tf4ou8BcxdfWcYjA22qC6B8kIRWSN+uXCmaZhRak7sM
EqjVawJPYNyd8vmaLKRTAylw7CIbUSHMkDj2Yfo8jX9KT4sdhTDQR6iWTD33tkVD7rE8gF/9IM4Y
s+Q9rzULpVFfka53yEPuhkKsxxbLxXEe36bB84jC6d6mtXVC2qhurD5r0gbkqq/XRp3zqnvd30M0
TodDG6N/lcp89g8/05h3Zqe2+44Knnkr8jtIIYUDH+tqXo8ujt927gs50MBBBj02ojhz0HOpypmu
APFbOY6jhkRjyG6N5oRxfdyBLqeHHpcmDBZabop7/Ga19EtNhXGJQzfjAvhDpmkV5XitFTgNw38M
zKEUkmbFwtTB3Q1DaXnIpZdl1Z8R5smEUrhDy9hx+k5AkEXhm6ohylTrE852N3kwZjYVS2Kzbwkp
lvx1fVsUsobJqS4DpM4qWwD0EsZiphJMfDIeRjpd4FBSs6gGWgO6YnhX9ltrp593fn68FRgbTZjv
YchTVh/PRNVbUv3DG3TNMVqAKSW+LdmBsjGif2n5y6wVkG8TQOv6bxCi5Pd6v+8AcAn9USUueGjN
eskCtvzl1DdJV+crEgFVK9xRrX4YC8FNjDPKXWf0yAedd4f/WsUv9RkFPTl2bWaMUqedu7mkjitM
9Zi6SCs1rwwIylyMFgsP829FkfrC3Mtk+7CyTPwSsSZf+Rftu239jMhMGthQHi8oaUFCkfdaqeyn
IeILt28A6InS+K3YpU4nFyx4wIXhofKrBQSL0yK7HAItdSf28d/xT8GIXq1uEbnusxOQwFKb37Mj
b93m+62l2MlFTMmKOxFRut3MpBFWdfjzvqMJkZBRvhC9zDY3R0Go6GZAo0+xArBEkxrcWelyE4XT
yXeSIYPGKPn0awe3QLDF8mg2/E+cipMmxRwXe6hL/OlrilL6yA5+WBe6G1aUuPtJS4I7IfUIDFIN
3/sGaCobKeQUXukgMcLg1rbsFjRaRpMBoKUtGZqeILcHHxA+RnepxAwzpEIrSeleNiXP2wOFeBNw
y9RmgHmbSy9kB/sfZJfUfdXGp+uIzrJiqVVK/K9nJOYqZCdFeVjJnCWLJjhrb5q8cmAVqaFRuPy8
n6Ma+zqd/962TBJwqRjidUDRVPhJVpuge27C2HiAtj+Hq3NA0j6uRjO/jhXOkYiUsATBRWxpw6mV
4gWlhOW80sMjBUIGiCOORDIe8IXYxqRJZ0fYGIH+w/RmSzhY5tvHveuEBEZl6OOt9wy+9dweoX1m
EE8ensErxZ2tXgnujSY2wrlA6yRiaH0E5Bw6PYvRBWGQo/yVu/OGKMYi6cyugeBXvVWVF3tR4fPp
dZz8ugeF59hgdtP97gIkKXknvec+/cjtHC5IO8tCVbByBq/mg08kLos7m9N2o0UOyuMydu2DpjZA
sJYHd9QsPgydANPPsAvxA4OxLa6jDFUFlIs/1GhRvr2l4UcxuCay+Mm4IF5btNLcnq2+Hnrbtulc
UTwbUEEsZA21MMA4u6hKzO+DVB1Djy2ZDzsPh+Rcm+stKHpAF10KumKSsoc+Msk7RZpjFP5aCBFT
Y1Mq4X+kOWgVtUvnM7P8LB1FByH7dAXD6rhVCV8OC8D6LX13zUVgKER7kuzqX+oOVlg27vNyAcep
P2/AxjA/hIFCzzm3xGaoE9gh6LN1HHVb42/xBCx2oSA5KtcPWCiPrjoRZ785V7t7fbjh1TebCD+y
Jq6rWrSqoS+Mjy3U7xLbScMjGRROEpcx41O0c9xA6oUE/6yWopaesutjHw8vaa+iszPUrpYKolgF
q9EW2MZlLrkmWwoIQXBFtBeW3RrvpgWA5b8Ix6BHcCQJQe3o6MvsKymAwtjhrCqInjifvXVZAd6a
PsAAcDM2hsZKBDSe1uXJg0xjINDXKppMS8wfOXqjaq1gHNZjo4qdSPSvZueVxpH0pjext7D+7nE3
PqgNP5rod/SXN4zk1uhLUEHUlXH2NxI9/pgqHJgEgGzNCGiu5wtXcfJ9ZuJcl7J3qxI+6miW+9XW
YeYte8+VWtWVmB3oM8LboRYyk8U9fGCO/VJRssLzvbpZMDv54dBke5K0zrqDcJDtOxNuP9wAbltQ
XPMMwHVzBDwL3CnXbbez7kYqCrYeZFd3jztpUh7/O+EPSla0kRebi70kojVCwPHVF2iMwOTEYN20
A+bo1gQVB5ZyS30yMlKGNZ7H4b/r4YCgRIMkUOGnM2KCrKKQaeZNltppPAydb2r+AMMKj+NKyABR
JCBo1HVvwX8t8+adBbx9BPp1VskHVL3k0UkB1pGPNm6sEzH0gEnrYsxeefJCH//Z+/ExFFV/yt8O
iw5ELk1TQzX6nrWfNKReZ0Mb0Zehruy2vnb+xM6W+9Q01/6ufA7muOYfv7qVHHwgE4nUB5DSGHBr
gXqUkixRq83hC6ATUdR9kqeNMF40aoiJB/QrW+6Ct+XrvcmYyEufzszt7yeaTXFg0Qp9//4sit5W
ova77pLQvahU0njQOkzW0d45PJUfjDz3lBSGlseHnY8aF5zal3/ka0WI17MvI8PjxL7xu9SmFgfm
Wj2wKHjH2ubk+AnCcusAzfnJEK6NKX6/bvRadF9R9Y+AxGoCTiezxy0jHfWXXhbQKsRTnTV3XjfC
IwlYE3ZN7lkgDirdJ9E+p6T/fu0NZ0HrobiUWSiHAQDtnXrnJJLVhrkk35pElbJC9VBF5y23MgY0
psxy0QXsD6Z4aN/V0KrIhXgH7ZPgGvvH4G4NdXVMZmckfi/+01VEFwYMAoZYVEZjdIKHT9o2rOXD
ynqN/LSQYptdgzX5BvlPBf9DhCzqLdRhRSgei8Ni/AtQT1UVLqPi9Wr/IUG50goxAoZvHlDvW2Ng
YgHTELI+eZpMyYl3g6npQ8REvSt6OPcjoO9+XKZWHdbytxz70NQBsyAj7zSwrupMH0UktStgi9z4
XMechHc+NjjbShp0OPoNETtLW7/gFMrNfLSnMNny5TtyP8X3IFNUmY4yszAT2NcjTaayyqVGNoGJ
Ii62GD0OW+OGy9l8EL9qxhzlEXK3j06cTy5DBZXI/fVxmgdhsxb80OfGdEWMmTGZ3a8VKKeGh4Wy
bm881/r8U6zSFLP/PRiF3BkRinh2nAXhCsVm7+t+wiynY6o8bk9qiMW397C+HExtwbK8mDo8IXl2
JtZXpkvEViuV32AGTyvvag75UWyXkj5HQGiKOgLoW6z1IaGINNZAPi2ggbtcAjAbOKNStieDwG4q
KG3z/xdJUIYZ+66Vy7uwPBOC0DEK2yYnyaS0GJidR0C+n7xGJ71JZcw7rVtMhZ1j1cIVQB9ktmJD
mCtjohp60bSXxC+0zrdzZtTwMBIgIbTZFMlIrGRsg8lvJ/jXeB0HADO14pUXnUqz3ussG+h8Tn7W
mfrr+dSY0oFyDs1dByO0nFscDSPAOBCj+Av1kRu6oksoh8TMC2+mnqEuyYWqk6w8VTscp62Hug6R
1spmnofXlRq0acLrhMzY3Z9PcI/Mybg4KFSoPBgV38JfPz4NQAJlXboQOmvGQoP53retU8L1OKJB
WChL1Cmv0aRv5PWQFI1UM+CPNFGzCBekeE2HkxbXJph0YuzzJjPCAwzJ79frBegFuP+aZruK4G8l
MTb/deut2HLPq8lVzHajBVp1dKk0fXQL5W6wEz65P8iMRwSs3wFgDqTCU5JZiY3r7TRgJVHctN3P
eX5I6ozIbGj1q4P6M0rdNjw0UhFXmgEqk0Uwm85Q7jTNQ0SbEvTbGYHlsvzzg9wH/jPL3UvlqXf3
6PniRRqe59MoTzheSUm9GaQ30/bhKvdzwbvwLnGCYG+NE/Q41ghZekki6xP6fPY9h8OQQ1l+WeUR
iiDqVosXDu3IsryC363zbVMhzU7+/pjtCt0nHh4SxvWbl8FMi8yaCaLINtOit/HohioTkLQxE0Me
emkE1drC9ujumg8BoMB3HaS+tD7rWnqYf1KH35Nuf4I2tyCJbbFkEPMSlzc4SfICsnpMj2mo4OCN
AyJGD3R/m6eT0HPICBaFcVNlGDJNmy76DV+b11Mh4w5no4SRz5uRDfybU1leyN7CXKJg9TR4IYJO
yy5TRz2SJ8U0IYVnZTDVTUKZn+lMr0hKql/Yd5hyYKQJs+qz9z9Ffst+MpEMj0laVPaVHsg5fM04
FeIehf4VLOkEKIhFJHwbUWvbkhQMw+/9n01ZcZqhRM7Y8FNcPVgvKffONxNtlRMXf2J19AxVO+dR
4gwwd91p9+qvuusmnEr3nvyCqpOUTnBEztnt7EV1TaTB/4mPUiz5weQhAWElDf9z3fO+k9hCTFrw
xF+Re5w8C+GYo6nl+qVEeIoO0/mIA0vZ7FvNSeehaSCAbrXloNdv/Bg4mA/tv1fvTh2HwGjb3+/O
ARPDHeyTrRGcANBt/lVeFhb4fML2RAylnrwVYV24OSbBg5ybkdUsxbvlWP+0Vsch3+oIQbDvIm6r
zMt9bGrUk9pCn2d/wpmDykDx6/Keww6ESCgFZjXxhZVclNfzEqrYq26kuHDI8Y0n+vSMlM7Fe7E5
zcyfxwNOeuS90m2AYOH5SCVybUyAMLK1rYH5V+tv4b0zjOce9CgvLaEKbRwZlLh3m2Cuo8a9PmbC
xFPxMwnflH0VhLsjnWpiWyqRUg0eud4xCLQMfhFZZsFdcK0VdiijYqYhT595fyiuebltZ33zcOIy
fEj3tSbtDYGjuXtIpVQx3HcoXv5/JNSSCQ4wVLMNcRwxek2o/Lj3rHWzq2hMNZEZXfN3xGdfjN5J
PlNWfQyVHSGY2a/q6iiQuKvfuk16zIEc4BeUpqUw/p4etlwvRrk0I62fx1yLjWx5fNSWwkqhIedD
CjbJuuesLH6/uG3Np7OyznSB0QyaE5kljJ+bEY7Zz2liqJQT3P+vwOnTAjX3zp/9tWfF5uXWM/cp
LmZ3GxXPrNqFp2cqB0E2LWbQJshw+GUc9qWVcud4HqtuXdwnUQIL1/ZxzxGlmKYAPeXpGQ9Bo7Mb
tJzX4B4hk8o7JxeJV3vXvsWrpy9nWM5nl5utPmovz1T10c7VlvLO++Q2SS/QgOrvsNmlfXX83+sX
+b7LJXbDRagV3iJovKS7VE03yZJsLsgWXmVGT9dg2DW7NJdXDloKgjnSC9DcxyNghdqk72jfKZdl
GNN8EQS6bna5ymK+3MoFw/lzpp6fdEnXs9ZhfF4IPfYIJjQr14THwaO3ezqsGqMZIl9oc/CLvLUt
S/MyiR55HcGMuIxpqTFJWNZoz/nUA8FrUhq6XJrU5aDO1Q1mmlKgg1tkoHwdZnaWGXEtm2WyXQ11
ZQb+qyHoHUdymYTtMeFexbXk1lC/kzbYyyzfP5ZkBCObojGAZ8OlXyBGoqRSnazPL2nGp/OCW3c+
snAlBAGzCdU63VbkCHowi2bBI/0qMNZKW2GzWrCrP2k5fzVO7yjmzGxuM9/xpxkuRPEGfs8wdh6U
Zk1b3zs6yqFf52aeJlv3J1DmEwM3+wN/WKs8qmKZV3j2Fn5ZXLp6fTsELg+1UlAzEQRs1RFDQffe
q3KRJue0NEVQ5XLj+eN3UcMOBfk22OvvmQkz7Zu6Lk2bLvMRdGjiNVy0g/FDjkTFzo01eKk63eDI
rYAiSrUDgD4FTOFpnXrhus45Vxbw/WjOarJcsJWXmc5cLaWbwFblZlSjVJJuikfv22xkVSDekuPZ
jaySzycyJ9lSi6eVM2GCXPldtZ+bXGqhDQmRu0PYQYXP3ESdwjGXr3G+WKxPqrxia7BJbXpnROxP
ppXpXGRs/YVQpy58k6LKs3/6d7rAWzf+kQUQ8Mv0JflrYFo8TgaYhp3gDur8FlOASajN3Ms1CiBD
igCrUfyrXsbhv0YH1HocAXnHN9kob+3tTfBINyoHtqcZ8Xw4vQThND0qS0sooax0gXPBCpmRckVY
HrUAYQL+KlKXv6aDRTqK72nUp0LzQl7TB3zZOg9dSGtkHezMXxq5Ta7E4I8/DRDTpvqW4zjjc99N
/DtW4niUm3zTPDLhDsKbX+LOBP0r4UTENo2ZCgWX8zZnqLolVNdcwR2DOK+Ygj+RoiTVRg7wl01Q
w+dUq9mA95SzThyG+K2868hh7QX++yI6kBA1qg47ndkpBrSy4wBgCucPRjtpmmGYiI/pfsQvZcav
VLIrH4MpcUyhwV1GXSVa9WtNBiRORv76bnI6xVv3euLyI+5Ppdh6v8bVL9/U9CZ8XKn4D21zOZkh
q52CcGzDowsQNf3ByjPEW/TrNJxlpObPXmaCe7emx5rFg+dBDS7kRsMdzT1orP11IQUdBkmmb2/H
BS/PY7ZQjx6rNfEr+YqmaVbGRUUGT23+dcBmEMkMDjizRwYrzDwW+irTDmNjiCM7fBLPsNO51vMq
I9bBG66m98Svh5WRfgSxL8pICdqrJb1Hz0HrGLtUBSpMnpkHaAKAq8KXlTqQ6OaHivyY7UPOF5py
s78Ltc8bAG9/5ohZ/ctsWDVBmoSwhd22v5oe88SAtLV4dSPIZsQ7dS3PnvL8g1DFOofv+/xh4WpD
KM9gqRb4Kxe6HDykg+8seGGxCN95OOL4i6Oljj82vX2b0qKODVd3ShMaW81hThNcKzMKuq2N+eux
sOBZeluNxkm0yUWt/mDR44G+lVF9HSgPi30hQVD6oTujEkmh94sj1s8qJLUi3kUeehMaIsqQWhmG
7+IVDJknVElbQY6AJxr9k78qqGVEg8CMmDzqtXI7iN2vxROKk5kufUH8meHUQMsxEChuK5YtPsme
PaStYHjZnSVlmDeDEMvUGa4TZWhCRCuGwr6iUnoyPlbdoPP3l9THlSXiRE4yhsB4fpKGYI/YzZie
Vt5nyFN+3Ldnw+DWS/UzWnC11dojr/5ryP1Yrv+eNcgM7e8ImA/sI+PUHsXD1EPYcu5QxSHG3Po/
d8gApsbp3dqX2nbJB3KQJU0jPCoEA5DAwcCcUKt8ME78O6eNU7xprJtEPcZUEkrAUhJHeYrBWXjP
CGY9jeKJhh4u7at8iOTRxDjrvWofDvMjWwb2/ValpJOCT/zvboosMBmddO5oDCbsZaawZOmc4HFk
lEHFxnNOzehlKQGJOzUdbUwMh3K+0vOR6ZWpPEA9cJhIJyTl2E6TzCSjugYyxoTKCHZAkbl/nr5O
B2MdgD6FtyPmT9wMOko5ZqtbxuuiT5P6xYEUvIvp+spqC9JKpdtH8zgQotZXlafpY2a0ZcYaiA/H
YrCsti+mbJuPorYjZteObSQFstOJeHT3kzytN0EG/0gbc5c96dM7w6XpygV2I1iI88v0vF9LL/hr
Ykv+qtu2A2mSKBTdg45pi+9CluC5vsGO36873jO3dwotmWfT5/Z7bDop1F7kqClCzS0vGzG9r7Pd
D/3YPUjXisGJOH6oiL236KyF1QVTplheOGn73moGv8jLLuuHese5RHCOVIhdk/jYpeyHTrkwqMac
1W/fpKso2AZrPudz/utvq3fzG7BS9ir3urpEdOvGjlIX8mXNRCA5CHjxYQokqn4Ga4f450SAmfCI
6g01kRVXHTDacVL4+1vaKZrYUNW+HtiCpXknLZ27R0zRMyk3B/ekzerIj05pAvPRWAYbH7qxJet7
VwGKxgXVU1XdF9qoinPNHgI5N2BeyEQINRAbe5ZzcAOQFsBQObIvdtEfk75xMDgvy4n05oH5BU9y
XGgnNqIa3VWy0u/i8sT4JBN/H3y7PGlhq7/qrazTqqCzG82YWV7FpoC+1m0DxDwzY7OHcOZrbxKP
rvQq/D4iGeDgdSnvGOBr5N7T3Kv6oFAqW8QoFcZDInqvBim2EUv1NR0zhbF8LayceOOjXIXDshZ8
nq7Kd7HXpINzUI860JgS5tIFqzcavQPQVzOjQejQQriae/hk1WPZmvrUdP//cb7MMs65LvSUIHlc
pDLyXM+UH61pRCl12W5o+6dlYbowLBhwqRZ+oLU78w63GikBlHD5DrXY23t+F0MCPxWFPt3oHOcI
qFUZkOrG14MHZh9ate2YUPTvZAApCFKlBHrvR6khUcRvgv8wsLwkaYsomqnNSnHzIpHf3xQADV5t
b1wYyTAigamCb7DxcPBiq8WbYGQm6Rqh5/iYVyhvDxovIRDtEyQYTLHLqGM5PLZTzfux0KTj73V0
3IqXm4gE/xgiCbg1gcs1ZkxivvHHoipN8FlrV8dSm6rtqfwZ4Tb5aDisTzvzGH7mJOe7tkKsevwB
Gnz+/vuhbik+cDAxdwUGcgBdw9jMhn9MW4afUCEu+z0eyUNToxdjS5kktKEisj1dPFvLSMx/1IV/
UnS/yeCCBPsaYIm8qj3Zqm8sgN2k1MttBFzuEzP4RZyhz06zR9K7JCZIrxLJif6rOAl1dTBQAyry
Ga6XAtUwxzWURIUDpKcaRPpQaporS5BavBGYYpcfPn71kANqPt2QgxKZq/cyER9E1cV5gbkcp13w
sZc3YaXpvz16PuGlZpVkHgCUBEnIPLgxl85gF6CItJAQGp8xY4p0n9d70Gmmsxy3yrWI8uCCTX7S
It3Hk3Tzc8paMpjyUzT0Xgejiw3Y6tLJEJU+kq2HrywVP9peGZgoA9qlTQdoZzVp078rFdFuPfpu
U+yyNODvert2RknUGDDGwnKkjlSMpk2/d7405vZ/g5054z5AKMySQOBSq3E4BL7tXcbEUZnGse5l
+yDDBGESS3bQP69JWueCjmDEMJFMYz52vrEOCX44+J7LbolA0Zi0gmHOtcn50KBAHQdvBU5xCCIf
egSq8v1BVGx6RVHgMhJn92xXXgl4gDN6vax98CnBtl3i8vGBhYMJT0urv3drJkzTaBewbW/drt1l
2T3fefqBqBT7snObGzS8Targ4qLT1iJy/pZr/eDqmlIrKHJu9pOxUE9011H9GkHKzn4Qdff35S3Q
we42hRYfZr3N2RcWwb9HL/M98z3vA+xCmuvGl8+TYGwuOQkZEzaRGu5uOrSXsVUjssrdD/g/h4DK
WPqNewz1q9FM4grOzbMo5t/1WbrqAw6Nc41x3gFRs+snOTgwhSVIoBE0MwGder8NyHF3Jnu2UrAA
jeefeCfg7kqwKIqvc9ZLRPg5Whctm439TAnqRYkrOAepGj1R9hLG/1FlyJ//QeLxK/63O0nu3Sar
3orirRqbD4tS5rpBNHQTzUNbVTq/77ibpOFfG2s5PvPIGC8Dfs8lzsuQUdv5yMKOKBPLQcle9izJ
kqpZc3ITHkQbduMOh9JGMwTE9zCFgtEkR0soRYUSBvEYFFoq7KYFAAleNGM0UQmu5b3RPV0eV9BC
ksxctnYPTKJPfZqt5N5JiDX4QdvNiLk7idn7oSMYlVjS5W+FtYA5XvnW55dmDrmEDZILKpRe8tw/
UO1mxZISRE6+q1q/ACqLgYTjwkQQK/B2lnyBpTCcHUNA3TZiGsD9vyG/F2q6nXXICvfni4JRAJK4
cyqdVLcysSLzzvbFC4mpyQRqrl2ojdApYoNXgFBBnRh3aVFMyTTyUqSil/lHJVKY4sVcCWqhmMjT
K6a6KkwK/k2J30H2PdyMY1Yna0S/ReussIaSLfoPHkvTiyOe1hwiBYVnFndhta/tkm02siuIYH+X
lrHnkkVMEwkXPQyknBnxF35XbJWTLVJaWxsSWjAeyBryWnGxA6rhpfNWpokWeSbTY0OzjCe1oO0d
1kKbh6AE29NM4PZBQdBZMfTrps+cS6GCzbK+/uTH6/vxAJBYl2a52nV+4FOkjcvyd5d9ptKUrcqs
6a5XjUhngSyyG9EBUbyZCfkIzHs29pQxpi2FxgluOwYbT6PvYyYg0XCpon2Q8Cyyo9e8Ux6MDAaP
tOs5Brq1Ni2ss1s3UZx4e/WpNiWvrjlxq9foKzgAGXM5YA7uEwCmcW8Hs8KZVKX9pX98sVgNrjn3
l2M568hjLqg2W8naJw1e/xFUIykid6CDEPP4ICBJwW1d2w56O0J6/B6e9i6Z0KsXsQvXZxj7Yq4i
w09bJv8a949POsensfrni/jKatuWuPPZrYLQ1YjhsEJ9l1a641QzIlfsi3fo1/qdHnKXCOGWJihm
GxGwGyuwvP/84GvwuPQiKMAnT9DuoTkdjIFSj+D6XksWG9/Py/qZ1pFXAr9K/4JyduJQLadaP8Ub
xb4KmxVATPd209N+daBXxxs8iwnE2aZ6biBmGWOJkm32i1+ya8aR7FyypP6ojNSUnyWh7AmQubtS
Gh/48dQDOEuqr6t+rtzbht2BDOM6sGRHCUTAEFVxlIaCI6Zs8CbQsAvgRrLLYcJoSbQULTBlZmRW
oC+6XK0LClDeEp/7Yk43cTnBXhRhxcmt3f11bxD2a4LcLHHD4uEuXGWBht5+MQYXWcpDY7ffGTv2
77TkYeyOvE3w94iY03RvukBhtlFZAOcDH65rc39sCwKobifPK/1AkbxCrh4Y6I9/8J9xPSsMLYtr
LfWsGMc/G348P7eQ6y1btOx/R4rRK7e9sEVzIw8q/Z+Slgdke3U+WS7Dct1dmScPBJvMHuCdQoXC
o0UKQXZ+kJgnnBEYjwge9dywx8Y/4ewkOCzbaZc8mAEE7Ce7dHkfD7McphKQO9Og6XuVhVn79GD/
IUFXPoJyspk0jerpMEwqbEx4owvXfV4bu5fyoemgMX3WLFlATJ4x/lePa3eBJyPjBfKlIUqZq6cP
4f2g37E77oXF9US3JoSZvdi1223S3Yhp/LagrxvyegQofCzOQMbRxz0m7aZ6cxNFrSp4YgFpvVQ+
5yTLOqhA7fFqSIy4Vgu+kZVFYmhQljDYTfafAZJu9WWWyeYxsCWjGCdQbvbMiI+DsoWf9zet9YQ9
LfvAIjXzgYRlbm9vJi8O/dL3BRbbfsyfn/bUCMrhrlROkrzGSiIfFB8S/roVarsOL7lmJ+OrDv7L
ibXqs82KvXw0q9Lp6uUI68ZeNEcN9HsunoLVxVXxpBLn+T2shK4kDJXGSedMLqRKIevdfYht1GBG
6yQ9+MiQZjQ44jlBl3cwmQvuWVZr/kmuyUwOox7bFXg+MvhTV7p9OM8Qc/uAptxj9aB7NpKEWu03
fFVURoqjiDCj+8elhPpaV4IbqOosBU8T5PKbOSUjMhKu3BuzvT9lTQAsPV9pnlxuRUTjZpS/ETnQ
Um2qmVNNSUf0kQKGRrcrzVCt6yto5zPV5v+ZVuun/nEYVlWtldBF+drSzzy+QVHwQHiOFwlHDy7b
Skd5eKDqOr3yxRd42UwzcDsfsgb57MGK7gxDhPzp26FI4zQkE5HePBDR72WBuPkIGmxHfLvIpfRS
WWbf8CFAOLe8hIltM9z1qqOXoYglyWvHBY3R2KaMPxFQDVk+BMKKSllQyxCGuh/BoTBBh4RQOCO2
to95EE+tuiGB7G3ZkSpWqcSGtkR2eOZUEYjtxVUdM3u//wc6gwV0lA3LfVJLebA4S4TtV31J2wfA
cZgBO5xXs+W57f7r/ksEJXFWJ/D7H2Xh4lxE1ZJsOXhQAMIza9nrptg1DAKxQg0hb1VIiibhFAC9
4AqWADJfKjKagO1hU206OJUtnYx/TkNbJpsEaBmIcTthG/AYYdVqbJK26gRapy//BWrib2B65lOE
xI+HDgnO7Pf7TR6JCJo5HSmd4/aiTqwXjwSHeB1B9nzvPkS3r/0bMwF5ZcsMKaRS7rGM/qEd+jHc
QFt65OdEmsGRkaigJtjWFAyGaKilevZ0CwobnqtIPZLifFJL1M5SscIuIfMuZ9gmNH/9j4cfrR7J
caHHCWI4qenGVcRIe7MpJIjkZ4y/yFTd4rklQXnfrendX3SAUgRYGZpO0uDwYJCLcBrnTqRqfF8r
FWNI7sKPJEAU4pXY1BGA5x/LdtqI66NsBU/fzN2UaboifN7T24L4bPOpEOJwGPsjIJV33131pWc4
UGw3+BrVjIfkQjRHo65IkIEUVxWwQDs4WZqxBLSWvXBN6R1WLnsfZnIZn6lUIxR0vugd2oLmgwo0
sxkxSJ4GbToXQ9UmeofwE4dwTSDPakAI82Bt5MORtUoll6guwJ2tFvbsCGJnOywp2bIYrlbnHZFe
PgdzETZvb95tRNW+rmRIjN8R+Fld/tY0yNULl91WgSUyckv/BGlu1MRXJfdf8clXbKMRR/ngrh1p
3490X91GfKoDzuVvEWBv8nBOWCu13NvN2uUFO0+1IbZOM98trLIQGUDUyEQ5nvhg7VWv8o+Kn7Wo
RWQRVirT64YEsxT7z1Pp8SxIxLrXT59ciRV44Aq5S+918bsOJm2CG27dvjFDzG1XYp4yaVZQpF/q
wNkfO/TgUmCkaSp7wKOTGV4VMapvTvs+T3FA+gSDlIPeFpMUJ5NyjJtQlj+yTWxXSn5WdD4SAW52
i3hDzt0hxx+ziXtRgjb/oYTvHzHMxj13FKkAnlh96nP/YqgKMK2oAL0h2fzTTCXY5Xdrqx4OZCgm
lqBWZiqp/nRZDdEGluDyMz1Pf3YhegWGf8mEMNAo+Ar1fBF6u/tcRbQcRk64eN/TbAp+hssPtty+
npgf1RPYZnSseQaX9BNEffVzlBVMe9UUNXo1lVniVsW7xHPOEAVI+NwDp/HDFl/IXASiTbvFeKXU
e6UJV7ZdzxOoNgbUgQDQHc+YlSnBSYO5JyKVt98wu+E0M66xvKWjdw5rNEDFyRlymzUSer8s3pD7
z15CyS2ROFF3FWX57uFD7HzqrVz+l6BBKr4vGzseeXXFLpZZQW49UJryOIsehGHxxdfwNpVFwNGd
Jpv7HLys4zaL71zxe5eLdNn1+2rUby9Tr6JKfv318M2armDJ12Ki9whiqTmXqT3znLRqd7bpr618
Xc48cYFOzO/hwqIrfkuMV0pC8Iz7uPtzT4+EOE6qUHWm931YAQYzxbCGS9O8ENqSa/apU3xNn7IB
qMNS0MbM1EIEOWZQZcRcSeE1DqxetuAQqx0FoWO4bH778pWYvkywwCBIT0mwDokbtFMbROiHtB4x
GKTgIakfqKC2WyurFap3tPOYhkxmRlhkcATZ7x0utSuc4jZEjgT3T+3s0vZE89J/I3FDS3rN9TBm
0HP7yIvysfSuz7YjwyCqCOtWnNqV1m95nuk8NAiaxnXv+M9NiLxxcDuwm6EOR4HGRi0Q3ZjDP8vz
dQxXHGR+F9/Ec55NG3jIxffK+lsO48txxa14CFpIQ1TEx76q0dsk8GVlzo4/aQScnj8ApAMXMP9K
fKbcI7U683USoCKGioR+W1k1Zs6dWK26G0EoDt8EWkI47ZbO6rlSL76BJVs70awKVGaAMMn7AwTY
QDWbg6Pn8TmwpeShGf3G+ScEX4Gbt2wSRifef0iO6bHNYxSNp1hAztoM+cYB6kleeHvZKtMjEwO3
2gVW5b2K+3LPwZyYNWW5cT5bdKG2S/dDh+5CIJc7zwwm7YbQD4hShh0HqBkjYZfLuzFkl9c2fmex
CU5dOBkyOYQENkqptCKQsoZ2IajSsVnxQj07xeETBz/T4uvB2KlvmCXb1BV21cEviKZIWuTMEk/c
PwNAaXSV2eK9XZPBFL/C877LmHgjMVx7JQfF/T+XrcgHSUeN0XMtS+LlZSWpEROzLvaznrUCtytf
6T2DNYLLlURlLvd5e4I99WeCwW6VD20xb0v6OmKJYRehrEh593ERo3DoX0g77UY/GChxh3sn9uU0
XPz/S8NHAbo80Nc9fJ0kWS+EhpCQlT1PKrbNpA+NiaaZvo4z6SQeotKuaI00D/nJ61KpqCgr+pL6
Dudz25GJROxxf7NuyQD5DSYMLkrinUafCqhQ71vHL27XhrCnvykHW83DWuFwWa+9tvq9dacKsjhf
qmaHnht6dzTMVn5nYTHAqpo1x6lK38TZXgRnYSricPQgfucdpCQRI08U7Q4HtfBNNKht2v5mC0my
++sev1taYTm01JjMGF0GJB59UDJBqnYyKZd2zkb9u/CssE7sIEiwGFrbVoV9DCzlcym1HO0HaWe7
VGv3bksAgiIEkOYX7PiPINiOiWpfWz4XaLgRz6J8jdDteASjNCAPk8StLWn94f9uYc6oCPAvOR++
fc94cbWFEs/EFmQIf536RKpDHIyLToc4lLy86wm7LynefPq5xT32TLUJy6tlzE/UiiAkvqGuzv6u
QjJtsIK76wBFgWUHd89mwMU/VsKaFV5jRIVCg7d2p90VfypMVhdZOJiRlgXoJ8n4h0kyJF0gQBBn
KQ8QDz7OsIMVuHmK7ctZZgpizQoAR+llU7emKKF1EoSQXGO/G08S42iS6lrdQ3vzfaSi8lTobY5b
2EX1iHaaaD3rz4leErvaODZwe89ONPIoWa63jN5GGb6CWfWZ/TgKEX6IwjHyuzNFH1KAl+jpkXjk
pOsYbeKJhBbpav70eBMLSCCH3RoMvNoqHZQgLIHfV6d0l1NgW8UeMh1RWf1Gab+bv3zgDvwsega9
Q6bvqVtzGaeH/hmvr0hcSSZVNXl8B0+IAc1YROBKLpCQ7BxSetSVCJMS+Ltom46DRdCrG4BBmfa6
qC6Bsegn+3SLkKOdElsMvvwEJ5DI0GTanxDenSWbdbHZdJ/vJjDuYowOO+m6g0vt51psh4RPzRak
f3jmmQ7fa+Jt5fOZDdrqLzdZrAsfBxDVf+SDE8Z8/0cN/NQi5OZzcSZ0rn1oxM8vKq3UtzMQ84TP
A/EU6xSyi8/eDX6yHGLrDABz8oYVUux7fG4ESpTCpnS0oy073A4JQliJLmdJvORkrTc+TBNCJ8xe
/jNvFupM4fduX532BN6v+7yJXPh9VIcIK7rJd5sOgUQFcc2vndrLvz+dktcq8gPIYWcJyBN+Brlx
JC2OTJWDdG2MdCYeOK3GgNM9CPH9jXV/6O9/0WyyZDOU/PR1FpYSGLlBGDvPVegxtCWrTc/4ZyVM
0wG7FtdMPHsUcU29brZdDoUD+afjyOubdkPTqJS3+Xq8E5NtoLflIQFcYlZA/QgfqV202FnUW6ee
WZaIOpzPbO6dJF+HQ7ePtcG2oxySSFPwe8HVJgzqxc0IrFdNToSQ4K1l1Wz0s0hnaigw8L2HHfYr
j7T+mkaNWUkBh6J75+hqHoWAwBtkyx/+l8QzAs8Gljl9nk1coFWVjibJnW7jcnaXWE2LpgbV8svs
RwRrL6TOo5iY+kvCClIg/GUZ26ye4+Tn5BtqOwopXIjhbDSEp3H1U1n/stvC8FpVSJ6mpl2gvrBB
cKU2AFdZRK7XmGKDLDQ8l+Dzr3adeUNWSZt8tHikliJEUt15Sle9xH7sLqUZrfN7QYLvdl4du9JZ
o6foF7f3IEc5d8Ly+JC2dL95Dp7/7YWvPmVz6jMFMNB1MEMeEdkUG/ZyEPm6YYgzXtAt6jQzXCAh
ui9BQ0fwqbz60HFByWM6bQxq93MAlQrYGpC7v8bOss1YlUY4k5Dr1w+KBsK/EQBmTm3xqhrUkFwA
JOCm4nVR7dAGpKw8Sn3guIwmPVbfYS4ULJFhpxCwxhLwWy+Q5FSznPrtOCKe/m6nSID01bMllAfN
wvDd5qr8+HZbPp9WesLhf6ONVBMt6ZIUp4xB8U0Dqia7b50DuAZYWCBVQnZVbdTo/H3MCLnR5fn5
yegW/zhIpvF+HCA2gPQo0jhpoGHDFwZX+7RVcp4Zu9ws7NfuMHNERyc3iXHHDrsChoRnaeBPpGyQ
wNQ16WKYryZjsFmjHunLCmHxIj0Hdi+2W1hSy9CVqNxhhTt8qiOBOGIRLJ5QseAN+qiEZuzkOZwa
vQZc3esORkoxBhl4+w1WXyjYhOXKR+3wsYwzAHQPR2292q+ZhAsNTmACOr7wXKwYQhhYjGKWo/Dd
o8/Kg/7G+NjlegPlyDsu4ZrVPpTIjinQG3iHD7SrLZ9OZsfpc3WX4uDqTQd/cqzPBABFwJd1lpti
nNqJjgICrPm227bO5Eo4fEz7JYzbXr5iIk/XWilxK/HsnH042edAGEVuLOac8wH3re/MJHemNh/f
EYSV2MA8BX7VHfWiDdz4a+tTi1ERiNeHk1ZTnreoJx1YFf4pOiptBQWUDWkewdXbj1Xvk42RTAeO
ObGR11Y8VO6/XQuUlgFvjLJmvJixczYbsm30Wd4M2v3uKXFTngJfS298+bzs3Ca2rIZqiedkS0GC
Z1zeyQiotOKPIQJRCU3+6poh1eNAPbLSn5xOIj/O1EkJkhWY4UK3bkdjij8DUJKE6Xmxzj0g41jn
EJ5DXsXNSf9w6QU6u3dINO9gQI+XPPrF0ALHSPJ5a+ZEoDa1Us+aLfCey3DgMxfReswBMPbUVRxP
/K+9nu3xuguhdO5WJ0Iib1TIUjo2bhjL/H5Gs+w75yQgQZft6wkQumGKwzOprbrRgXQrAC8AHURG
eKvy388Cwc6blhDViB8Dht0QzR03C8Y9TWqBuYfSfQiJmXDBouhOAuzZwie5I/35vSwT+PTmRaMq
Z1y8q+57UkxIq0V918ifytrg5zyO1GAh2ZcuHAX6wsxkSwZMqzBvjPjOWE0HYYdsAOLU0Rop0wZ5
aqs1fd3ul61n7RW/92KY4sITikyng9lML4wBD0llcjkmjO1mY6/xPon8Qlqbu+SFvFbweXZCeEdm
1Ax/1D41jJ93LoVWjG71Qhn1WOraWQ/pYB6e8Jg3ARy2JCbcLIzzbLKmbxLOJ/WnU/kyFJ8n9HlX
RbN8RFZVt9JeUEUlS4jIJ4HGmheHbHFs8FGxtWUbPAbqM8+NtLpCg0IS2p+GdWFlTWUerg9fsWmV
WjfljRaWa8MlFhfWYqbIjWyP3OrSvBeaZnXWII9q95nAobclpTye0CCd8NBRJnI11C/Qsmqa76xU
XN4Dvz47Rg1fimumhq+9uy49t8PfLW7zv7stZ9Q+4XNX6XWSybTt06O7UGAfItD4cOxN/f2VG0gq
1djd+D36gYiuEaYponf+v4MYeGLjuiy2yrCc6HuXz2iTnC2mLptLRFZNHipsevYgmk7OHRvIeMl9
z0X9VZdZTarICaHtzyUJOmYeo7DoCe1GDGttisc4dAEXsW6aa847558bXsk/Xq0cjc9EQoWDJON/
Z8jkNK3elpTYjKPiJSOotKj0F/okkqaGDjOYHGo9sIWtibDrLkT8fmrAeHdjRT2bB1DSjaNYqEhK
i8j44t/rSycpmnazs3Ic4xNsNwqxtm73/4uU7aSKHevx6mP9CI4IPYnQWILZV4JaZOFeE8gHgoxJ
3oz9ZG/mVv1/L6bhylgd4wvXb6lbl+8G6t/5EDU8m0OZ7uYIRbtreywk4LngIulPm/gUucPVC/w/
vkMi4XFQTvM7A2blmBeeEMaTBDqS9MENZ/A4WhvXoRhc/Zq8cYEO4wnrJ1lqrgJ/25fySsFzZVlN
gu7JS65EZNocMFeynLNJrHPDDevE9Baet7JAsmgbSuXzX1zRHSy09cCK1bjJ9Tup5kKCsV55AXd+
WNd7u4E+8rwDZp5azNZ3ToZ3nj0JPYCvwxu3YrY/snPYA2nthIOpOhs5+Kc1tyLRnr7W0Szmyq73
slj/Ft5OPMZbAy638HmoV9/sjrcpOmwofFGzE+4eTgmITVmkKxGRqEgfcMB1n84rWf3tsOz268x8
EnSi37G5MZasJSO3ZlOAgrsqtZrwnwtBeqtvTX1Y8eBQE+2zERiLRx5UtVacd4dfcJyWMtBjmAHm
IhhK/HpG1m2OGkms9kr37l25WT9We1/09U2OtqM14HF6BppNl00FyBRPrx6EuRqWCoS9qsmZCTL0
OCPD8Ph7C5yAV+OAfeRSnRoL88mWxvqGXubKuZX8l/bnYpnFI6WZu4hKxjHPX/R3WV6RVRhpD9B/
T85TcNg7TaHLYDRsSyjHTU/rwERGsPoPTvFP8tytkAykWvUBEkTzmpJnPdYaCBAlFllWsioPAJFR
6E/fvYTVPxI3Ve5P9RD/Q9p8Y99Bviw9S8bIXjrmGxb42dpZe+QF/G/9mdprVr2s1aOtOhuRD+nt
Lc5iITv5mxVOssdgiXGHQ9Xzb0gDYSKc6TEX4MRqD4Y5gQh3Ql7oD5AYbCOuK9Fe7CooZdxqcP6B
O7CPeKGaxkFgPAji1nz6yMqZmGJC/7e24tuo3X8Z7NHFMvMmEyGc4j7LqvsVmDz3DUluWe4YFs/E
BgU044ZBOQ1D/GFocS0tyESaH+F7LbhSqdsJPqmeN0wVuYIIVc1FakKOPPDXHu5k+EX6wvCQdOWG
uizJNJVfR4koRFCLL29X1Y/vLridGip5atQNCR1uZGlDnHN2SH5eFRuQ+FK8SgpLcoeB+7PNNktD
Pj01IfQuFPfkExPRMg/7DFuh2N51Y8GIjfdmF1OE5TM29wgrngZjX+341zKymb71REX1q2OV/8e+
D5vtJiKqVC0oZMh2gi03Mq7ja282TplgeWL6eE65RhBrfIgGlxAH8WZhhALs74JawTmbfM8JxNyb
sVEeRU9jheXsc3IxJC9LvYyPyXRXa9+7x4d3UaF+pgk4v4JvPqZBROczFApyRtvEMuzc17Y4SsoF
A/xKSppJ+w2GQbX0XXHxeqpAaBIt+7swPv/tapz7On23AxGCu56wz5Oku0Nt6wSYWeOXJxMdC486
mzzEH4F5tV2qNkYIMmlDktL3nhaRiXxzG0ZioDSLxA7oEQQN6pQcZRs34j6mT2xfRcaVNrrj5F1G
KlnVYdrIV7KxK6zzXw8401cPsThaexfyANxlc6HL5Kgw13ovacOr1LxG1tQpUybibVNXDjv7OtYW
tvvJpuuznZoOZgyiS3TT3KvWqaC+EII3/A7fb8p1pq+AT6qxGFo8G/+7fGOzINE9UVaj4eMBnmu1
IHZpaFVY1CnDEkHMpxLCQVSjk7qsYpRJrusBQZkCQgYOV/MOGFmXWyA/kbSVzPdVvwcKWJuMa8oO
+UVox9NG8oF4XpfeoIsJvIID+PNzIrjmVPEsYDawt4fjd7qzeZoZFJjk4V4nJ+38QVKOcdBbAaOh
FBXb9KtS5rKhWPooGFxuzrxucrZ5Dl1qUretJSk6G4BkV6WHOAoyOCErKzuBKkiWow70DP6nc8AL
zslsnglj5QPXrVeImsdCjOdH65gR9PsT6NWcvePUoy+bHqbP8ORfEAKZQOuLpNul0YHSCuWBQ3rT
u9dpEz+qA2QXP2bimL6bhtweGoENuiTBSemas4H16NudZDBE5oAOzJHOOt298vkQ25La9c/KysqD
JLWrNyHHFfGwquwFzACAUf5YkwXdWE1f5TVirqYj82dJJS5pVsK5NA+HDGvc6apVocCMaX+6l+Ry
jCsnE82Nfr2Di6eVPxmZqC4RGXQ3vRM6dhUjhy+LqbRRjjcqIPX4zuzQRn3IIrtysAd59tZOXGwl
VrZ+PusSEuiCk7BEcrQMgbSBYu9F3kfw0Xfo3WApiRK0D5ryiNGvx4sh69xwi5myp8tRueckWlck
eeyRS1MMdIvBNPRK1suqFhvfbi5bDTBV7iQboLD7TjwGiBQ4ImaOv5feUlvVxtQZtye5WzPn6xy3
tf44bqHW9ufuY1qPRlapeeti+zLDltFHK8aa2dUTt7GTjZbyDJ58OSV8ZDPcwi7gLlVzrzBTS0ph
t9ZNgtBtcDkmqEKbyiIkoZWlnTuNw+Unvx3pbWBbKuUmm08YW3h2S/eB1hjFr6TbVo/x31c6hVY6
9QE0UEsZcmUjLiXXB0s1HI0kaCC9kgROa/UEK/8quUiV3Vx4mTpFdrXAIB0CPsLLbPAAfb4f0PRj
FXHEop3sODSAYpr4rx3l+rO7zpnn1nd0wUAshi1k9YoLNVUXOxbdEYhtPQnA5HfwKo4LeF+NgHs8
QBllyZAprFy5mKy5oSZq5lFEm0kuU3uyFoaTVV6x5ZJetnrt28SSzB6Z3pYt0sbRty/hkqAStGQB
1TGfkO9bnzg/yhxUMhn3Xmr9SBuYm0nRjoF3wHTddo4PwVBvqDT74not++LnySV0SFIZujqsUoxx
meV4rlmR0rK3NKsZRHnCLtQwX029mdY/8NXFelbzXs2fWO+5gjSJhDD3ZaEPxc4m7hADCT5zGVUR
LZHGcIH1WVUdtBWNsJKcehbLQ6tjG7RXUB7ospqUifBI29HrSiX3eGbkXOos/EL9cFAyxbqxYjhF
Y1PBTlmpXpJZChhdf38Cl0pwMY6oHU9oW2gWDMLwjRqPJnGyJzE3UC7KK099D1vTDRZaqHSLJCqB
fnsUa7kZ5/mLk52YP3eKEpTIDp5yuvrFrwKFGB6nUnN6xjkKbIGiyhaxR3cEgkfd2o0dXsZEt1oJ
Fsrl5NPjlyZYPbj5q+vLR3HSP6ltS+hJQnmwhizIqlea7P1MTPgV9Zpee/r08xXrmF45B/4KH6jU
+KkLR6+x+AEzzmPL4NTcaJDFiY8VS1HtiBCYMs9GF72+MUs3R7LHwwf1v8vMRGPdJbZnbHHWYL9r
kWlGxXROz1MNdUDLRyNNNqbtWWjhdR8gO/sAJ2fNfU1JAWI3vtyq0X9kaDpCMs9SYevJRDkge/bZ
vOJvR2oxQaxsmHiAeUbGpkpWs0pzJfzN01vXyuIquZUNb281+TfsBYTbFisimKpu6o/aSzPRgVnv
dPgQaa0j/+DkPRPvY7dzdx/lObdirc2jJls45dk+lnDMRvxu5GffQfpEnUcvW/147vtLM2M2g4Ac
u1Zwn+gWOADW2+41sm8/s0n+vwl+Ke+JdcFPkGlmf4wU+rhfxvmrX/n99I3vdq34dn6/3MQR9lk1
CFZhiTDstSepcbBOo7nnMoWdpFmfgwQaH8qx2RjwpsY9Qp/CbCr31TVSPO/IpcOdsZfUUR0ymGTr
1Jd+eK2NOl/H44I80wYsaehCfzwsk2KQ0krIJt/urAf5QSX1qd1++pBGaYAdUjwC51C5LEnideJn
2GByEGRUjb5rUhh4DVgXOAHYsPy1K9YFQgaqyeto0q96lPoNxrHt5cPRhAcSi/Kcy4uSRxWDEGSM
h42rkxWoHDb2fqCkSzRQ1+DJyfvj7NFwT2PYtXctHrIqMgyRdQavbCVAm7z29A7j1VZFsw/ayUmx
/ctBUW7xP3g5HqqPt4BuOKSgNBlfxV4P0RaFfW6TCjP/Q8DRh2ntEaVqHLKMlJr+sy3DI4t8xqI4
x771Or+egyNIQC4fnxA/xmwH8MirZS539HUOdl4ARXml0lrbmN3BsCG+0oTPKrbDo28zBw9GyS34
rgfSkH9122EZFKQ+0anq6Asqm83LBVua2HmYGpnpy0J6+Iek3FqXwKd9YPSBR5TyKDmnTBlw0orH
W17/3govhdAoCIxW/kFdj6UPhIC6Cs0clCbdb5FqmI88PMfYJuQ71uIMkgWk09+cvoJONh5/242c
F+24e5mufLAQN9rCltlri7f0F/OkJfr8eLJbdHXxkjeWHHzeBCRuZUiHESlxihXnzzQfXRZKRUrW
Ip6rA5i53/q8nL7QNrtmiv8hWbtcyeENcritMoq25fvS3FdPQsP41KiBeOFswrIwumYftIXpFoHH
aWs2/dIAELYDGvhNVpPZ+EOJCaxThwRTyjioX7M75EMQEZh+zJ+D19SDXYZi8YAAdm8MVChfh7JU
4viEczv9R72o6wPJjP9sZ3jx/HObYWGyOR2Iqau58vl3L+7RlypWqPprU3XoRWlrPDFp2bKmIdtx
U7x1+WvKpz2IhswHbjV+1yZsySdsR3GtPaW17PbrTZKwNN1HiimWcDSJMrJ05BzcTV5+/nK6heU7
OwjZlTefPfEUJ9rHh8iKJ2lN0bznSqIwEcYzKsRrUmgMTJCwLPxXheDkxHuiOpPWPUzRjA98t5QP
A0qlTAQTvpRBm77LRDgPV/9pjjlTO6Gqxk/CVMjC/rUWttDgHbsenMN73nXJIGswpwmaRx+mYSaO
G92YwBgv6hIwWT44Z5VwYCzqINGgiJ6j2F2PhO6E15cUK+QR2+HXVnOhbjP/i7FJgpNPZd0SeYvP
sfbI17HVNB541jwouCnA1T6CGLkmtJwxiKUNcRt2Qg9MkBeenwOEmsWmvT6WSssoHPQ/kN0utuAb
hTpZMmgaQXlWQ1LS8zKCfPgcB5EKopRtsm886k41BX59a4xRLWHiVdw/HhaMKUhhABrnLwB2SaMl
6i1eOpeSbla5WqIWIlTloIuVLFB3Qzaq+o67cCT5RTrfKMQhU2Z/uW1a6FNMBe8hXDJTv6OLEEpg
fs0OxtNqI4thduX/h2kFTLqTV6GvLpJ6dpV20QFrQzURes9ez6e95wa4W0d0KoAEEto1IWebg/ZM
mGq/2nv+1uMbc2KlCDSo4pCoPElrNuQ8N7QBw7mfqfMcO3/hFoU4bRBiFfyErQ92AEdks9QpHJr2
zY+aPmvEXaIiNoWrSVAdTS8wqD8ym4AX6R+j2M5KixqlXnHvm2CavTzX0PVQJjIGVJ+5mpYZholo
gsqyGukcXmQQSd1YqonAb9jEFM5j9p54ZV+0QVq4MEmHG6QREgGQiFI8aq8fo6tP5woY913MFFWG
YHCy9ijuANASKKTnr9zQrkMzGaG/NneN5tgmBhHQG3F7dwRI0/2GKMPeZHkl7NlXXz7cURUg4DnA
56W9ZFR0iRUo0SN4RwmnhwqcI+2bymmb6bic1pfRmIpssitUTBrWlHtlU3zdD00SxqWZ9dZaE14J
OyZDUd+M4V/mx36LmTTxC6gQfVEOIyOmRje5Fw/tEHSrBo55UHx5xROYTI2eaiN+eIJKzRIWOMtO
wOnyKZ8882ZHsBEeHoJDi0RNrtjKLBCtnQxdhiCLOfnQQz3dNq/6N0A9jqJ74PPopDmFI5wavYtQ
YtXoR3NBVOu3h2oVNr4j41Qu6ZEMsxi2lpTX4SCrXIIKrbxZnwjGkIJNWjX5Q5YT9eFSazTCafby
5AYLLnhehuyKQPtxdA2iXy+c3ee8QwPuNaeWFMf5gGIMkZNhkeCR3eJXU341n8VXJw3puXyrC8ja
a/k3LGDWVMyafMmZ7fbxWn5kFiQpDvIu2eOTJKdr4AUy6LitN0IWz0k51iyN5V57Mwb0aRRL/cwf
pl3xCB5FeTyXI0CpjnDr9it76Bp8EFLEgROkSWJqORniE3l+iaeBxZ7aAsQNjvaaALaXnuw+qsaP
B8deSNNJAykwyYT9dhHLeuGs791gvK/CLyzNMoNai1UEAOwmkBJWWTpj6SC4itDdCBvji3uCAcck
wQiZ8h6FWYfO9zJaa4cHMpR8pmYCisCrhOYXrXI0AEpsIrLu3TjUwinAFdjIDHpX4eMCMmuuMuEe
G1tI2rFVQaLMHg+L1/sYna9JTnCNxaF2sXSxKQh5FV4NBRrMAUS5NXIXlT69af3lZ7luzgShABE6
9b7gu3IIR+4DyZO5uSqBjazefnDgYtk2qZSn34wA54SytkzwVgD9BpvW6TZcCNynIXrB3pCIxs8R
LkNtl9ayaLLHM/MNAFg1h7fWzcRorsyWpdLSQ09NjDiToZSM7jwaUfF7LIWho9N3T7sQfkUMYM4y
ji8Ug/FE0Wt15gZ+up+IO5stZ8Uk8XsdzBImPcJcfRZLivvxYxkKLXH1htl6tATde4MuCN06GNTm
uC7vIRVvQMCQWCotGMWu/2hwlErY5kExPgsqjK7oNQr2eVJwOBYy2bLpzhzAlT7qOH0oMpr8PwOm
8d0LgZQ1kc2TTss6Pp5eyf+aTsYsYCZSt6F7kweFvCaRVq8CGTBJ9BlBGuBsnKZMtHsujzY8oCkY
Xc26Ez7RXSvLMfDkWPm+KQqWUaBmsqVsQYeg9UMC3g1bUz4zxK1LgoYlILJOPs1gjS0fchBsMjuh
8vlHtcRcPstYMQZLbiAOl2gQ36KV+7PkUdQ/8pKprjufrdZ6XRwRaINNDcCt+Qp5L3W5v+aYLhp0
/IHIzqCg3fJyq6JLVGv/ClUnsPYKptUclAesPZHOnNXkTSBD5mq2+ubZGF++3oIEAPtEdNiZwkbM
2kIdUSJ8Nw9SgiLGVS13bHlvX6k+ouiZvvUVM8KZwF5EjchaaQd+mXr9G2UouVdL4h0TZ7sJDxCm
9baXm48nT/TA0HVGML/aXAYKKwCNsmRcT82f2Iydk3WlmOIQWEcfkldJUKPvAsIQfzLIcGdLqrpd
l2bQNo0ZvazbhnvTqoIshHFiHxmQpHct1lvMcjPDtnDuL5gg1FddsayPaXz1mAjldTKpcqvD3XAm
7mphEELu7XkmClU7VCtQdLWGmwtssXW4VcSrwX4DZLI5/JYqshJqKIufH3gTyXOHcjybTiayuAaX
0u4IsxUgFEi8wmscWSZAJ1Fvp8frUDbokq/Sr1j7nkdzTrRot1iKELh2s6N9T5xYtfnUc/zYJlId
wFgdMxoLBpoa1T0HCXr63pMOaNmPdDdo0gHOUaschpD3t3QPWrqne6n7EWQbKfSaC09z+bLNpHyA
3CIpAT/o9pubJ+rDtbt7HTDCzqnpY5TgigkCKnrCYHwaIfq8q2CC3bg2su4jRMQwWtXkOdV9FO0v
/zDK6usnGO2W+Eus2CAFWO/7WEeN5eNG8zYtNAqJSu1BGszA/Oj0HBWqdXoX93XK8kE5hQP4J01V
uCqQ3TI/K4lIOpJDXTjqJF/ApL2NG1h5u7yvnF3JvjYJx6CzR/nm8nLVHvheFNm/FOb1H5ZHXWa0
nXIOmWFakqX7gRZtmhUqkdBtj1vYGQybWJQ6/DE60HKx22aPSjozWCYMDiRmkOSwMGF0C0YSTNHq
4U9zo1l99SMb0/WzlXkaePe7eZYDgOZUdN3T64twZ10dkb4my4jvFDnFHC5aN1cwlS/wIUAUtnpJ
eQVLVDgX2nEbbUmTTFBghHhvcoL5vTt2MOCZDKzPgFEVchIvtksEmQ8N3NvJLxy5Wznz1A7fsfRu
rl6jnuP0/19veJT0JW7AhFmENwYvHIu0qyvpOqtZrX7k6x5lTrsiMCtk7aaXaEN0zHx6AxXw/XFL
z5sAOyrKq387q6bC4+l100E6mmxvdX1ZGl+SYbweZzTDietPNU1U7pBV0f2je73mLHVXCG4398/J
n8Bz5FDK8VDgaTZWZtKdZb6PbVjq2pYz2mY5OaO4gQEk8dWpRL/UE/ZZCaWHFrJD3I4AEiYgy0Ng
I6/SDHMESgBvWUQtF6t2Q8jocdToBcOzKZFuLhzKYCncK8/lSQLvPhp7IKGOGNv3MEwnyp6BweA2
wZDec2L5avytfk4vOQfsfvns+WI4m1sc9nhauYH2dXLHWCoVjK1aU94ZRYV3i+MUCfP4pGNw6BVg
vHPlNuxmwmDJtOg2D4ZMbHWYVol4bAng8SOOs8K0Vsou6CNovIcDfSZwTtA3jg2ATddLczxC5Q2q
XjPMs9Ud1a18bwY94VEFTajMobwuki+ceFGZSqjN25zzhLS8l/9POG/UK7RbUS9LSnUq/iWe8mtI
A11Agju22J8cXw+6jta6HMuXWVns40HocQrYFXE8KsL7kJwknhA4bdpodBZJ2U7k0wI1Xq5wmS1v
tVTo1o/nL1OefFKA0AJ+LYnHWDBeul+wDMs3Q0flx8EmCWjDlhSqOdS7I63sRKE6tECtNz0l6gET
XH1GIjwj4guHxTvZ7+DZvHod7ICmIwiFVJH8lVZvVjLwba+f6MF9TXeq5pvKKglXoJdurxkFt7tf
T0IlkJ53QS4CkhRuq4ltsmil2dw9cSW7ikY+vCAZah/25xU3ePiplVDvj6LLnzIYoRdMyqMm6Q6C
1Jp0qli+ySZqJ7i22N/CLQkGkK8iYJBJV4RfX/ECP34AvngxMaONtrVgjnEC4ak6TSbKgaccMl/b
WQZq3VoR4GJ8x/jww3hJnDD6QHdP8cz/FmcZW82qbhuSYUQFbedgCs+yPTp4RDspHQTooXiYpMvl
et1T0NBg4zJCV5aM8ybzpIxmdS0sBcCeQP8VmfJeevJoLmpyvEhpNdwwbBsn4qbR+q+YPZMxTUjc
4yvmnsDhiEklzwm7XpMpHlfqIl+3WkelbrI9flcuhBJPa4/uQEuYZxxt5udbqw55vX3IEPbL40j3
6fhY+PFDayHDRI3x+UU7NB4BqObI/t32SYgFrwqGFsZsGd1vanc98Zjwu0WbuyVjGiSVrQaQhYJb
ygyYzzPSLwqFSrz3QnkQJjIqcwCYbP1W65GUYy7F8NNdbIizIrjtra2wRJE7HVJj7E3TCgLoFXrl
VjRXgrkj6/DjqkMBxiFaKZy/nq4FhZuNbJs67WrN43l1THqjZwuM9Unbe3GqFMUre2hGpMX08+4W
1QuGKf0WnPuXuoO6Mu9IVXuel7HOMPk24geX+rKW34LjyNCLL/zRp/sbCS9TtIK0yVeq31JMITri
0Fsh8aUlkMTy4aITP6ZdnqiLVEioX0XxuYPvVFB2Zr7oovoJnr0Bc9zhWjQzO8iMVAicibbdijsD
f5uUMj66KnYA1cxDOk5wzkGsALBdra4vno9laUu/pAG+nxD7jk5asT3t0zTjlkSRmoDACJXaVxwN
MAJyt1CWYRtEmxD8lP8ApOBt/Ya4Nx7bwwvKniHnO/vf4cioeGlqSLm68iZ9gTc0FuWcUPFjQhoa
nSY54SmTN1Qn0PUSlQu11++eonlhQIuZwfVLhp/qdOxgw+VahNzHS7XX40WbJdXEQEViYevhddqi
65E4PPl8uYrniH3KU1C5RadzTj8jyz2jOX/xTNr5mS5viTgwW9rtMqi1OBhwl7G1zljIiazxso+D
FIb9l5OBiDRv7Amt7JfPxUz9mnM5bOLahU6v+LN7PSdyP030IKmmTOSQH3NlSDXvSeAgHhChYO86
pWVFt56PN6+TdIsYlUOPrH/omAqHF2WOD1tS6NiJKhX3ljG0EhnzT8RumlX9GUXEpJQdDp/IJ35o
kNs3Ha/Ny6xQgfbnB1u5hreJUXTdm4dcPWtFsVN73LttdivqA6VwQxEolK6IzhAnVaknQI5aulSq
JrjspE0jp9h0zpFO3nKZnKekUKmeJAgKsfo+GfxQgplWf04f/gQ9d8zFC7ZSzyVFczV5c3sPYxI0
ddXetYK1EqOxh9OvfMS4+yV24u5ylr0SK9w90pWocgz6dkDonnTWHEVHjg/ORw6uztXfMbbqCtWe
q/M8kRHuBfmvGxn0BHlTbyiLPUWpDPuTw/SXiY3lEZDkEDPrETWMGIJ3E5Mc5hce9dbft07Sp0o8
2jQbew/HtOayxPBEP6GskBiSr3Jf5qzHw3k+WaDbF67v+vtTLJomL1GKNoSSEtSWjIJpKyhBAUur
1VHCuWb5ynkykKpsnHnsehpCHAfwTn93HjZ50fY2hxd+NfgAReda0d6aGU5jYz3PHqgYCg8yvi1Q
RUwQHvGi523H+Wkf09S1huzZ8GeRpdiCZvrq3QctLeOtJKL329pj2npvNKo8pQtVzFvcEJsSOC0J
E3ChG+WoZ6kxcWdwY0rLkSusugqfyycRei68Scs9+hj4GtZtMSiDx4IC7pcsF3erIvfefdlbp78u
HLi+TuNYpc/ihUhV3yhpIItJWq9hutAwduirZZkmw6G94LJRwtv4dj4SVwuKbFtpTaaqzFam02ME
FqN5W0e9CNXfm4S9f3inl5ar0TyTOlLc1oMGa7T4RgIWmMMohEUOxf8eNZOtQLFl6NLRiS8PQkMT
ClWzpIwWkL20LXYkqodEwA6hbMKvBGwc8bc6hjTJnCdZenoxoZJU384Or0K/7qZa99e1pqqDAzST
qv69AF3fmp7Mo7LCcTzNSfQcK3Q6CvcI5uzvMMTibz8pIF9vYGMy/Mv4hd8GnDv9zH1QSwYaOt9C
6axoyFYfcKGySNvG4jmTt47eIaSz2YyaHlYR95dOhZLGDJznSPhO3schrESfS6gU4NWh/gYvBfgs
a4UYmkPpZH760AzL++QDT57gZ9lZKy1mY4URdWf8JQ9CmlKsEHi5NJ8iKryJz0wkhpZtl419B/7K
WHAWoU+ZhaM8cLqhkS+GNJRTUEmeKqKM1vgLgQU7+c3yi0GSgpXEYNErUEohYYfYJ6zN6huWpshM
zqLbPsrC1hmRbUojkMmb3K3g91LYODYc96bQkv64tGxhjGGp7irJ5i3cu/83HdQ1ysY4RO7j0nPO
uQ3v7+U727bHz+L/8e2Uj7Uc8IVTHJn5wqNvg9GbQ4jdyTAcTk7uyn41vx78IA9LpTgHRIShXzXp
i6J5khyhiOkeGS1vXPRgvCCQpOZ7iodYKbci9wyNxgPVwOH7vKubC9hDFykH1FYuNxXEbwQVj2QG
KguJtsFpQkHo85pyILC5z0skniJ7sY82x0OfHk38baNHhsdpKBvo123fs/3EkaUliPs0MIf1bOfB
h359iJQmB3whBRX9gJ3Cj3lu5/S9s5oeStMHkMkylkMf3DsJnqRD1vNVsWsFIZ4mAl315uFvddnk
2Tr6KbjE6M08nEGby2if0TlHf+pkAojehArSj04qQfflygi8ilS/EO8+3eGQBY7br13JUDfNEW+h
ArgMTsolcBUFEmFKPx4Uvc6EDjsSri3COSEdc0UE5U6S3ryh7rHx55HppQdlltOecs1FXSeFG0q6
Pi1TZ9yLYSFDZy23LTMlGkW+lxx/uQhx1JUtrJLMMgHISwLrUgFmFIR5MaNJ6/qqfmPHvtvP9rjc
0FLAUiBgFQ3t+LUlWZuVgQ8y36WDQDOKB2JEEAc8goPveRfrhMgF4epQR2aHKWzRY5sGUJvJzprY
6bRNufPPVhNq+LgOjklLOaYoynXdh1wK8EncRkbVgbhAl81YlzpDlqOSMB55zX5u9fjnozfPzKGs
4P0X51bTRYlku1dA+1tJfuW0wl0o2bIDdjXM9QHsAa1MlYNCS65gvhZvantUHjvfI8052H0E/yu6
tlxKR0+m7ZwDbVCupev7o9apoQks8TopQBcL/5qYHgfSP0dkrs5KDKTKnW0/isench9OTqBHxWBS
KHMU2bIeZ1Qotb6h5jwhuN6NThr+FvwWs5NOy+VgsZA/C7l3M9z0s8evFStBPDSxoB5/cgFC3oWo
EWQb/HWEynzYEMKrez+x9vVDa46gDCgu00zvsqREszMf8oRmtq7a9VJciaILA9DgkOGYHC/lrD8L
QcmzIJeomPgYOYD8KxkSasaox9N6mpJG5rTfn+DsNNhHj56q++O8jvrewQMRPTu9ZYckp8wgj05X
FzduNBYsxBe3XRsDo0LtzQcbBnA4e9k9dafB0x567CTSIS3WKTvTPicAlhr/MUH//sFukJQmX39h
u0Pu07rJRZ00BUgRfrD9az8IdNEq4h/VA8gQVjjbFKt0tf1i6W7zm8q2/N0CQIGgvheLOH7E0cBY
5GjCC9IqBI1WhlpUAG6vyaYl96tMmnUgdXm3kkyVRdKrMLReyGXgUU7dX2e8VQPA6dY2pnok3E76
O2Ze7kBVuaMgVdwqg7p0PxW2VkESBmiqtA0X/iX+3yxbzjO61Lzbesfjv7UNdnUWYcm5B2C8ct1e
uOMGoawA+9691cUwbuyIPqoaWp3MGOpCEBX1+/gqAP6CwQ3lskSXwVPSCTiGIFZ6vsEX+s/+1M/W
kq1peKQ0YtrUuXiPBHnzT1A6pNifEyQbyPGrghc0Dh6S5qZSJpTwU5vaFL5RtAWaUPVgRop1S7/H
/9rgl7dOjWIBfNDgFMtKQfrev1L4uDcAFvymheodMcZvsF2O77bEouprqE4g0giFQ80g8+eHDuQg
MPHEI0dD7eHP217OZ1Xjqwl5r5qFNNVs5puoimTm22XH8qZGop0sTYwupolPNDZpMl/VP5nXzJR9
3nzsk08bbxqpziF/bneHQI09brENNdvfW9YrQm/VImNADRM27332AfD5WIqjJcnhBBTGISz/M8eB
SVs5X6gT3TgRXU2xRc76VhSKMvGFK5Ns6C9LtXltZF8AZyduCsRIKewrUqzPtIWGazMtdm2BEUq6
tF6NS3HagsYFQKl5nnJwNSShrrFVic5CuEAzKCAHOEPu5ypr0GAJ63LiTh14IO0nyvQFT6tDC05c
G5rPmvlHPiHAat0b+3ZvtIWlMrnAVgYmlPvVPJ8AHE4tYKAnLzTwXdPNJOAJ5pzR843tNBb8JMk2
CIxm6Ujsy4R9A3nhOn1RviIqTqzKB/tU9OYCxC/AOV/ftQ0400sY0rSQTJXR00zHdbFT14+f3I8n
0OcDTXmO6GUxp3BVoblAA5I4HNJtRCGKZ/joZpMCh5PpdkpBU64tvpq5UyVRHR/M1duJpB2LoyYd
PQTXrtHhlshPYp17FpXYTAPHj/TX+3XxvcGAlGJgqpYbHJkryXpl8RwmbfMjZy5uz63Q01RTGf/M
fZIvyTP/fBtBDJfO9irORwZ8EYmfNO5HvDObjEYGnfHjVTvKhLtaSmtra+thGmVnhUQwXoZalMqK
F+gJFxMjJL+hJzHOOeNMhN0A97EQz7nE+xBXa9/iZDI2pTaJ2vTWI1z81+9wouzEihJy/EEYGSVX
kySvcSP1ur2JHiXScbuZHVpKXO7BaKAbQHaeCNNLVlNMwGw8gd+yIxHPQE6jNTnQTgiS7+M0BPMo
C1WV0ZQGyabpC5Y4uxzkesD/Ti6dzFIaN7NUhuazDu6JdcJqx8ml+dNrdHyQdVbvHqE8mPyVZ+Ae
dff0aWAwz6CWNvXrKD6+86G/aWoKtI63hqdVfHytPAVMUlumKbyGkZUKkvKA4Kg91rWVig1/HXg5
oQd3ClRihzQbVm7RRgkuGi12mLuM7AKQnDZM1E0CkNvbdgKL17J9BqeUGs1WzmnZkefBHvwdASLh
i7MD4is9ZZWLFojJWNg6hRAB7vtYEoAAutEV2wZpc+m8GP/AGKYphqctCwPlq8OUefREZKQVuENV
B06w7HTZpfLWA0nAi7MQwuZEFe5XTwIW+WCu39A7BFm5PwQN5rdbNiWIW0A5MGsI88ZBlT/flw+i
lzJwpjxJA1jvKKv0AiBpx/sFRXHWDk1yhJ/BiIpnTuaMtMvDM2pHS2D/5JUsKsB57zhTopNgRnz0
SyXU+L3uCui0WYxvbqrUBjxPvRzzhpM70oY+Ici99F/UcCGJ2ve/RVh42c48ErqiKMOGmrGqUVVw
34GIGPUorBMa7RyOIcm+NpxB/m8ee0XmvfxVAopOOZrUfx1pjEOxA6rhIhttajwCEVhZeJ/W+7qC
ns8YtqdsNpMDxvpoFYF0BI88u5HMFHtmaFQd2tyCpHaMiBrDTKZ0SV4d5g8CG3DuAneCgfoh9IBb
aC65WtPxljeIuQTlZ2TQpk6so9vYGm7oz7eqVH8jz/c4GhKdhc24CVwiXeGG78sP0umibDfKev2Z
VsBb6carsIQb/qg16HmS8z3+oW0kDmLhEtFlo3G+8vBGUERn/rDB3CMSJ8HUoOJd7TWoj7u0/hVH
X2fb8k/HPtQh7YbZSswS1jTqgKD7ctOTucheyCA3fNj3U/lAdPAyNNLvQTI/CzDOwUbEuGl1+cYv
WBL3tUyuOEd7UuYnZn0D58RX7shYYQgqvupe0tWkqplFi1cARXiogOoc6v5T9xOwQgvA/lpyctcb
wMG3OJGvNXI+YLq85bOTjprXBVfZTVRJ3KzSmNdHq3FsUPTjBTNeSfqTtwufJJ5S6jEJxQU/LLLA
Ixxx96hMhm7iBvXSlTlVtOnwZYpu4jqYx4e9W8GaYKrA5vGfm34Zn1w8UjFAcQMZwemGjzEGZTlm
SKZzuD96mPY+iQugwVFaqBWT2daNBNNXAKazhoZDsqzAEmfPqxHFHRPK/fiHsYqW+7F6P6+DI3Wm
NLM2BjnLSAFxmcqPQKdQjP2DT4FucId9X4DdQ5fad+acZ8TGNkO3l0bufBz7xEfSSvW3T5GYdV25
yaYSgSJxJ2q0hnCTgR6NEvFmgPzCmohSGqPnFvfAfMyWNPQLqS1e5nPN6+XLr5JgqDqx53CTivPP
U6Ksc5xZHFKd0F20AKTRgZ29erwi2UGOeXn48yzt2sXlsuoy0g7ewM7SDzeouK07HUDoqZb0Dd6C
eYsw/ayNueiAx3ZIY7/wC1HJaFusZFViYkvd2TjF0Tyxgdd8pUJbWUGW3B32os4HEnLsMpPXlnJe
Zof0chTnqlwY2q8OUXzMlO9OduCDPl4qcjOtZPHO4G6LbCEVoC7uoKLlp1JGK02N+aLkNI0vY7Ec
A3l/xrpcLa61ElOrxY5VDvsassxDb9OyrQnYHjsztW9ys5yr2cc06TJGXzc15gqKX5vKgc7N60Nc
g+0lM1+BfuXEeByCNwb7Kyr2A9/vvf+9NgkgxzM7pv/zXB6OCxV929i5Tf8TtGyzKIZsCaQ4P98H
dD59RhguiaYasYhzd4pIhkt0XW3z2l18NxhCSxrhsf540KFuxMOYyyQZruLoLomRsh3WckNd/9+8
TsVrQZv0O2iVxH3jh0OejhjEO9G7rTsVbu1IXiqxHWotAWjTuuM+bjPFDmmCXnCuvrVFibtSiQcU
+1nuTpIs8wLbd1x2OsgKlUvYJLQM0NWHlXynasUiB0mnXpnXqHIdb6zYKUfigQmWz6tr6KqPwD2P
vJZYsL07z2lbmnzIw8E59kc3TFs0R9yx/x1fM+luSTOs9PJUWaWqOq4jnzjWQRCzKe/vnoAxjQ69
XxHb2YtjlFU1sFl3Qvg6xeTyVmio4o2fRpLFDXrBxG7V6Eje20f0bqdst1RjeBCpBTM0htZM7Uwh
GAA9Px0HT/DFaQVHPwhB16F1wfmShww2d9gqfVF2gaRBZb/nPia520LKf0S0W89oY6HtrE1gWGw5
TiVqjn/QYcDAAPGXSQkO7EBG3DqugjY8q1H439wfchSDAfWlyN/jemvQncHjn4fv0uIH0lITq/0C
e/vjgncRJ6+2mTVO8pj9y6VdAAFtVdDQdOZy79BK64b3mcTxJxwO8NNTMFNLJdUNtbSNY1IUib9+
R3z2sxCF/29QgTBCQvFcYQkN1fbPW45H0kDXRUU4AaZdHNFitatjJiuiAqG4E8RPR+yhX1OVz6Ax
zhRXRlBudVM/2LXo4Rw8NjRGZPbiPzln1B+MdMCZt1NS0MrBakj+G/FjPsoqDg7+I5FyUf+fPANd
L37sCr446ovlRfeeP3ovFKtJWvsNC+FAZpypHMxAQCN4budC4dNqdUn2TcCPXUT7tgi29qsApfkR
vOWLq/JML5P7Xcm40y5P0XD9gmoxmD5StwaGvjG+ZJ3WB+dJBJX/NVv1dFi8QGjcT2WVJvJhCxiw
eHETqUNFUxVbwV3cwI8Zce5VL2c+LA+iwF9Z/C4OxZUJhpsYkTPijpJnVic9N2/sUglaEbDu5Obe
uXEeqswT+Bw8+ydKwoGMmVmAlNRu/pzo+Qw4JUJybmACvXcTK0c3KT5WYZ3gfyncfRQXaYsllI/k
MpYtaiu2v9A7a+1jixnQI0FCmmpJquJW1p/Jv3prgxLTiOlxouUq4bSCGt/uzKmXVR98/Dh0rH7y
Iv7vylEHDhioYBeVvn29K6QjGmT+pwKVw/2V33DtjXBmFlyVqDLHxsxVS8GOpwmb5CFoDXV7DVKc
EY5r9WcJf9Ibk6sG6s0k/rXp3G6AKM3+X12kbVVRZm9n+id02/6YUj2yrx+xlS+alV0SaqRES71o
k5ud8R3JbQNJQ3pkg52nzg4yRPDXdlm1kidb2HiNxQcirJOYv7nu/CzD6Sq/JwSFiZErdvQZyWPG
lmMCkzWSMB3oHDLEub8WLJzoc4Ov8sfTCfTlWOxgucJtDlA2FmnZngIQvvs3+Gr6qkWW//Q6Wm91
J2qPGUYB5ugfdMTwQzkXriwo4vWkp10YDf6tQmyYj8QH0SESgEwkDL7meXbcKLC/HcBMgILw/UMo
AUSYB2t83fBTo+TwWYKQVGIkASBbPJCwXPjCk0ge56te3+RbXEpyAHJB/damSoOxFryPr5lCfHKT
kNGOkAM/1kUhvsxJ517jMUsio8r0y2JYB8H4te5GFQatFPemIdQuk7RoKo/VRxkQWPEyujIvsDaM
LtwwiQqL3qByJSN8m32o2E7AfCOF9T8E8GiwHz2B3meQYvU+LW/B0hSPi8/YYScdo95N7YqwuvHG
yT960jKYqrcg31u+a3PUfSqnrnmExUFw5iWxvLkq+NdHv5ve5e1AwaU1Fqt4KaaBd6Naa4X9GgxN
YM5nI16H0VwzNJ6tNMreoxXuqJVbWUWKXyzDrf09e6d6AfJbQkoxguR3kUqQ9C9Kl/Koaa6zAVKJ
rg2L6cQ6OHs+qNOSw9YtZY/sBX1XbOXKHAORMv5RyhcHop7hFNUNANa3y0huSDVEbr/dCa+M7aS+
W3eubFqjQVnAv8LfuwlqwstmjOuL0zAIMjRis4oxpysUNtmscaFv7vz0ETlux7PTIWFEhfHDcW/j
EadOYzAukFhUVma1ykaUcYYd1ZPV62BKC9Eeod0xzyrKTO9OeCy51HeoNgAH2+QMRkWIhw6CD7cy
+9hsyayHNGH3ViUR2SGmuG1T73PQwggHuxe7pHuzpygbEswfB9l63G+j1/ACgrIEwiVplZM69XGj
+XfZAspWKDgQPFZyVpgetjiPsWu/GPNz+lxC9GF9ybKx36jSeVAOOE2veF7So9rTSo6TBmra3ysj
VdkK3zYLMrcSoLcXst1WAhs4dwHjbcoFhlkRlU2cjXd4nL+qSPFEaK5VQVSMGZXkPaDi4w+aoIHe
bnEYeAnneVAsW4b/Wd0PrL6Sj5vrkSaJHPQLuOGaYU3WxIy5N7un/GaZpPzi57LekKyEOQFrdN1Q
oAYTHu9wdGlt3YxLPRUZh74F4ryhKXhxuXfxifuVLNkM2UQ4kPGhyYOcZXS983bnkcgquOpzF8aO
HFEIVdwJvei8Q0yC5Au/qGuNOqumR0iBfyh+HI+bVM8JvF0w+oEUl7tqSs8VgtfmPJ63p0VB0NDM
4JMrPwJ8kX/MQAi2H4Zrc7dlyNYT0QgyP/U3tT7w92p8GkNG1jdsXgB07YjWCA90RKhkjOOTusjQ
n6LkWzgbnkEuMUoUBA/dClWthfYA5QadvYvVIhHdAvvDKg5KSwUYhbnjp2Sg4aIan54Rkyf2UkLK
xMwKED5S4BIWZIZOorGeJMHqq3PA80oSaY7Bi4cRZD0Sq7JbRaa0aXjhkCLopzlRNamrTNAMR1HQ
X3RhewqLFl0OjU7jHnpMpd/MOOuzclVeFEEDUwoEx+mQXWVJyv5eskak9ovyCqBjzRfQptlLYuVi
Tyik5B8PTeUkVa1gVoCsWalTpZR+gCIfW9uB/nMbC52itUwuPvE/9wYSLQcytfanFeoTwz1HJe5Q
QeQ0IQxHhuyKBF9riAzOztgiMe2mW6a004Rd6VMfAYNerGrZO9bYO1Bjf9mL7jcaM2OIeHt6jm49
HGgat+9cKKg1kzyyWtf5CG+3UQzksFZSNvSoTNOfyAsXbk0odeg7Eh2tEAlufy+dfUl3K6++khWa
JGjND5Oi+994EXS7JL49ONd1qYio645dB67XHzGXpBbGbuuowEjLIla+SnadR9WK30VJVrDai+gV
86wCe1mpU/OXsStc2dJe26YauBTPeGrtDN2YWUxRnEkF2X3sQoXBdcINDHWmN4vxISSITophSvql
XI5SpWSU/SuRlUEJH7Oa7e+LLhyt5Olba9EDeQBB1AqP8IwGzshSX6KohPViHZNqJbs5wgtut2q+
8YJWtxjm07s2Jkh8cnUH++lWobxKtiUXcjQyKrOcGaFtGiRbqHhq/5Iu4PkYrEmirCMlwfJxv2yi
PmaLT+5GAC3SgU9lBi/29JwPT6MI7OYVhzWFdco1ZHFRMUrXq+EH8hEfV3Yp3WIrAwjY3J8J/mFg
+RxA0wIv18hT+L2+e/mBYRxlH43F+PzgY5IJFd6275zmUhYqsC6CFlZtwEqb2y32MaHeih408oFI
5oWYXq1dk4c3Kdiaux2DMXUiH2ZIoNP7bR3weBIsESi7tmrd5CRgdK9DKf48irFquLucwN9O0lK4
ciq1iBRIIW6+wxEzY5VjTxiEP6ZHblxrg9wRl/KzbStqEBlhOfw1egkDVbccnFgBBKyBkNl18Fe1
CvSz+p0HNjLhFaWekuVsyNqzGKB+oWhUviRBdM5F6OV6QT+AFjnk09VWo0LTqbqXCWJOD4tV3Wq8
TCBtGeQlP8VYR5Pj7aVR5S8sZUFXY1rPhcPH5yts/7MS7jlHIdv+uQKKWc0K9W10HoNhDseFHUP0
fMRScC0jssokgOfi1BJs/nMdcZwvCIvluwhns9hTgGbmbkd0z3RmQaa3VJIRDa/x9i/B+HSi7IJZ
LzNvCOkXlitWc6A3IkS3CT1bKMvqKklxc9Q0lfdQTSECz7zOfJFQi+2kl6dQv4Sl6c2DUt5kT6hV
yLy5jUQYCQo9M67+I8ETeM8QUiIzoBXvP6JyAiz1kfO2eXCL3uR6W+2L/24o5iDSdaOWlZPvwbND
Sc8yZVixvnm3PKNXWAZjNOgKt+16VgE9Lq+8x2Qn47cNjE93rIWlDbpt+Vdsz1bnC/GhzMYv2Cfc
62k+FPOlkV6LHGNZFT/vO2oCKnAoy7HzWc4aRPHlVYo0uFrwx3L5lwcm69jbAc29O00NIOugseKt
kihrx07FumPVMif0DVaJ3F1/fZtB17nwFtzwZ7BWabDsQ1QbFPlnmHlneTN/7cJASse8iDQFJH7v
ZytZ3/XPa/DVgNuDsE4hUFszlhNS3jz20YcTAOaTxm9mOYoTF1uX5gKsQNwFvFk5ktOubZC+LaM7
LgL3yScFDWuP1RhX5yrHHZlUK8XVnwhcRjoz5RjezwKtXG4h3ECmzuJiFbDZFP3Gyuh4KIKytuwz
eNDhy9ZvH298l5fLanvAR1h1jyI26inQkgHPEbcc2ObVB4EL0FU4F+8sj8YuQW7O2Q8GKwivURqD
TVZrx0ql8V6u4XFvjXdghNcOW6YUcszgUVwWfTJRADPXrMv1AVx1GiIoldhfifDSFXRfLOJNm0/N
kYiBvqGvmjTOku774Tz1eplEwxKORmumvR2gRI7Aug9tIKKBTOaAFvOzXGpXI9AiHP5iZBBu0Icv
oSZMIvkzEwEM1/oOPKOhfhU7s/SSK7imsQtovLgM2R13zhjIKHxa6N2wnAuh0dmzXuOZ3vH5oKCO
OKSlCvgMz7I98THRiO7Eyt98Ing0mfbXBUmTzKev335RMq69d8LDLLZTaqIMxHFSnjfOIcrH+AjP
nnSUgoGnC6WZ7ei4OYA+nAAlxU9EThRh+7TwWlGOAP/JkA2zHHMcoF7Bs4qzS2YkDILcUIV+lCwl
uyrTPYx0w1LbjyjLp4EfQtkgDX2sBj7G4cu0s47F8ux5/gJeXSBK6qMycUkzJt7YbY4YabIftNHi
uV8XIeXh+i6Hf4Dy+xUHGS2wTcruCXYWVIh9/jp0cx+ofPjqYSjQG16tWzogmuLFMChvm7v3KG6C
d4+a2G5bU+txIdOyYQ5Otyz0joq1Xq2+n86vtzsoe2wwz/fG5gmJ/FWUm/2WvkLPtzOuAq7cyK5J
R3IBNwm2OPKOrGw7dB2d4kSYloQ2KWKITXCo757AwJLkso4zKRAi1Ellg1exbAjKbPioDRbkjhmq
XsdV8rl+DuBNeuD9UQzxB5VVIXuD2LDE16XxNG0awD7abOiO6ZY/OpFMxFAp9ZmvTLvNQvloCtFe
CQWO8kMMezbJIt1B0wll6xFnzbeX2OSy13w+tcBadnhGu4L1n3eMBV9djzBUfrWAqBCC8w0ZeOA/
SXFvJPge5HjNQze/CyznU3weUweb2n7aHQgQ0PJxj1jfvRW7a/rxQ2eFXoNk9jk3MdofZ/0qCP4N
FI9DjnnMQCZSUwOzjlmUjVltoNPPqW5OrrcYrzVC7/3VrmLffHGkY/cE/465tjKwHG7jH9IEpiRU
EjMJaYihp2W1XSvL5JMqQA4Fx7jvnlnxB8tHc+5EwhXVtINoZeMXFCH1peB04sJhHmPNlVNcJMz6
H5F893swInnyf3F6B493dKJhocXM1B9fyx5VTIkLbgPtRdRyxtDw42MyJEIyMYjRWNohpqUazLC3
TiToMRaVdmOYNBdWJ/1TD2E2rXp9Z5JnY6Bp1AU6fTQLHQoGsUyZXspGJo/n1/JBh3FLOfr7AYBq
fVTJzvmNh3HDpuFTc9ZAi4RxqG36h6HXgXqYKxNROjZ14vw2fpjgThI0wAl2MFqa8gc7GJvU3vXL
Ks7Whg8HdsjD2vjG3ESKg/9aRy3OHCFU7BQqQT/7YxOJeeSwmnrU22h3UVevZ+MTgcSKhjhdt9jC
2kj490nKJFN4h8rIhsB17/9jblQsCQCZaDmX3HEGpAQSFvEzsZNriMkwHI4paGO40Z9tYgD/HnLK
OpZg2hEiDaQE3GXV14P0VUjPsxL0I/oKMBFLMvLaOG5EEILR6KxdgrW9k7ISFeEMbP0MGkwlF7F4
vzrmT0lon8GY+OCBMJnERlwlLiJ3QqFpYEBy9lw3wxukhLP6fW8J5a2cQmR6QJpczNZRCKfokFxk
LPkwdCX3CS57KOb5LUJgGly14pIwK3cJtwT+PvyaZNvWdHEeMpdn/qHva0RCN2LBcm5qednswKht
GyEBLim+B7NjPdBzwqaFBXPT4ShaG/us2pRjudHQELDZR8LLrJzZqanMZWYR4u5YTD4v16xm3wJt
OBQREB68EkwyySOGsr21XtsajVreJjFXahFek4Vb1TO1mirPbp04HN2BzqDI7fBEKs2nXre23gXR
ewDL4eydhIq+wIng8YFj6pMUdg/N/ihdK7bZXpZanrZbw8QWSFX8qGayZ7Ul9QBSml7QFTdfVdwa
4mtmqz7DsTMPpy/StDB5juLztSIo3c5rNgEmZCzpqos1hnO3ppeN1JiMVieP8c3gMTHABqwMLfeA
lmM0uDM9WEyAmzCZMQ24pMJO8J4r4WaKbxw/NALkBku2PW9yyMzhrjpE3AIaOU4CVnkajEHtOxd9
GMK9Wpjrf3BL8ORTB7oh449DIFf6keHluSm/NPlEUbAGBzLWS78aiFAkK6QwswmpjReoE3bSEAcq
dq55h64/pb5VXRUI4XmOt1jtZlPNTkPF/6a6wG3FZ0b02A9C83+tfGtSp8GsC0ZZp2JtDtf3tyv2
Qd/NT7QuI9gg4c7YGHJ9MNyyL676IxOvwxPsb/r9XWujcpJhSSt3nmWHGzKYx138OBWWTfPCS1pm
3tCd6Ul4piMHwbk8FtMJrDR9xi0T4XcE8xBQOcIxkFqbBS6tNoDA09MOArbMiZVhPgEl6i6tX0ec
yM7ZwEbsq57Nk/NcOwl1BlAPUbjwMs2o+/lh8SipE12+XwNQeLcmeXq7MD5mwRcZLd99ND6y6KMe
7330E0xT87v8telohhczENZxeR2P6mjkr9BQMKgFJcMomgNhZscaEnwkE1BMidYbOoI4tmbGzfhe
fGOZc6jZ+5XNIOQ5ImRfnlgny0yxynf7aeGYNjs6GWGqy6jwhnmoUoofpObNBSc/RYMdnDQzUqz2
M0gJ4y/6c5uBHTsgjrak8wtsYcyYcfjYI6fLMDbqjM8krGWTMvN96SXchQDaIYJ8GTdYOnVeVyB6
67tG+6OEAdhDUB6kn6wa7DpzmqBhjS+h4eItWRKnTgXnhhYMzSLRmw16o/qctRjtrCFfoZXuFBhq
U+4vW3TS4CKTtgh1T/gnoGuSjZUlJyFRnWMucdslEDgiBLWsGzXJeZ+c3H4RwcVjChtkZQVtPRWO
BVQcCKSn2ddqN31LYaZGtmWJJt63kwFRrVr4ZNjPm7rR5mqUVP2PZUBLEGJgs5EAexXjrHzCbpob
k7Udt+3WhHX0uVFM6eb3WT+tsx1N49Q/AqYEKHsua7mqVnwjc5rdHDDFwv7ys1qIVW14EW5zJR1q
LDqS2E2DIp92Czt12H/r97G1JQrxmNaKSPUZpNNrLIsZXb9PwLOM/LUJlOFpYobsnf28iO9P3Fon
4/dnz0O1vSb2g5cMa69tIRQsG5Sc4QOs61nDPHggEe51TRrUzqU+1u5cZsIyxsxVX9t4or6vQ94o
LmzwDM7ERaIjbSxrDMehJxLh1rscGh2isAx44bIzwfenKNuk6gQp/K4yJfA4QP3zk/2WpkaPss9W
zVEoWk7hUk16ns2TZ+MxGl1rtO13981vBDGpk43LyggBWT2aUxqcWJ1EXT4MT4ji5TGfDH9ID5Gg
FR6ccr8vGFv7mvooEGo9d3k23P4oMIAiplXSoKpEX8yxX5D+QpCcyr3Sh7SBxlukudqKDD0ti63J
WwNHIk11ro60IBll5Pbep4j9o4QflGZ37W4EmG3tpu+DGkcbedSkt9B+xJ43RkfwMxaApfDoFLDJ
VWxKAI8N9LoSR3ecT0iVStx3McI7d3mgzqkCyWCsUwQYxSfTCnQwDnXzTmLuIa4BGUz1AvXUGFcd
LvBs1CxjPha93cX2kCsq/PhX7QbNs2o++A/gQvRtT4+nlMWBfrwX1lsFq0NNswTp45yZRcGZM4bs
7y9El93Tmw78Re9kAKJB3FdZt+fEVI01IxlmamDDfl7tSeMsuswNUcfiyjB0Ym+QyabtZr5plDV4
t6W7K+ouetwjVHshLEvdo5fswrVBifIRDpVffb27jmPp6luBQw/3DKodGWXxJaq/lVnGLSKr6JVk
87EWPcktSqnH51YKhfCwlxR2keGXYhInmPMIfItff7z9MdfBHLAz1cyBk9AyTe2vCtupyCMiCyoY
KYEac+RluZpIWiSYd6dgOY1gELEZTO+ZtJkeWPVPCxNbLEIm7isfOzwI2Tdg0N1mNPSVt8o3lQMl
PS83NH1OxIxH6tGTlHA/vXj5oI2hm2F+1H6h/3CdfpuX5HQ2atk32y2baW7k5OXm/QKuXr/+8mGx
iPo6U/a768vnnhgPHv4EfCxMYLyB4/9h7F9YSdDxxpUFLkLV32+e/HAechDVNg6pRxonX1RZECOV
rmYHwex0jQI55dQtPE0IjyOvjG+I828i5zDRvtJXxcKhefwLwiU/YRQLB5EKNrZN7yyM1LYwlR/K
eJv3LoJewBsWMRxZDLufLOMnSGIEKU01Q8jELb/2hs01XctfehhGKjDvLx6vCHV4sRhnm8FNl7Wg
t6S0q2a+II5hFM+SeTsO7PCGc70amRWWyJnxvbUfXl4xN4GCbDRa+ua6Ns/bm00Sz3BpMTaYu8b+
GW0LFBpn0kZuR3cWKxDc49pi31g57J5c1gVFIyNTxSCw1h+z3tNwCzkob7NCcQRicyUiWppM9iZ8
qxFnJN1+rV/e22oDSkQ68IN1C3aMZRAs1UJjBrDEsi5eK4iab/OMRB8Fn1YT6PqyPtD+LbcqKIlo
l29i0BsMRQmOO4+BeCm0j9AH2yU66jBIl3LkY6KNsiPj0iabEjrsLaqfRfkb5TBQ5avpq4ZWC0Q1
aytzSELG6k0o9ouFTHxgtE84kNsWQcgMht+m+K9qf7bXqJWYkLSihxIkaQPQujCjFXekZy5ZLs3a
gBmeA+LFDEu6Najet/aqrd8xmcKH7kcOk/wQeYYhVbaRGAry0KAfNJqp7kOUE5qiZ7FcH+JQc8Bb
R++/ugPD3qeIIGlIgRxicIJFxGzbjjwt102ugOgKr7QZNO3Gi9mZtpFWV9/wWBaNiZ5PGYn4/WQx
BstNz9NBKx+QfbxYcp+6ykNhPuJaB6CeAfLi4di6ndG+OLukTVUtzlJREdrVpYIvuSG/7i5p2Iw+
MaHdBI9T5l10/v0esbRn9rDal2iM4Lnh7uffJ59Z0qBfZg0y93k25R6b5TRKDBJVMVEh3mb6IH4B
gs8hEYDoQE0IdCI/n/KpqnrwDcQwxHgpcUqVX6ai+dNTkUw2H7N0QxZ0KRLd1aSivhGNW/qyyKpZ
zYykn+5FbBTesdsdlvjJV1YcX9QhChPyestn6bc22iWLLJw82LjsvWgesO+nfMZCndcsP9Tgm3ES
wjFuWXlefDTui+2x8uKlUCkDK0AZkI8Qm6D2DtOpufXBKH6J5VlTYguvlbijY8rqdwlVMhiao3SJ
/dftGrLokXeLNW4HwqBdmVMn6qqiZMwM2Iqxb/ChVzdVmLBA8QQKYl8NeBlb6JhbldKUVG6q3Z/T
Y3IR87Gdpkhab23elpqnEx9A/oQpGa3FK6j8X+vo8ceGcPNAQTypSyNG48mu7dGId97jooWVpDNt
XO6FDFNpbCsiQW1hwazyS9hUum87KzRNGS0ZLbY1gO1c2fHJ78HmttrMf7R4ebGIg82aQclzKX90
HL2l1BLD1r+O0SKcfA8RUv2zwF0cVLO/Ir6N1bCwg6L00CpqaNjxqpbD/LRnTJrCmJx5DyVmvq0g
y87I01Ym7p6mQeWOcmf5CJ9j39wV0SXEhoNjh728diOstIfIvNnBXEszw4EJ44OTaACZuq6nwjdo
4bDYnNhk9SSE/fxsaZihetMa29U9o3WbdJp6QTOwgvDL0WhLgYaRFTDsiw+NV4pfML3Gwk9MisHQ
U7l7Jky9A1SdUVWmOt7Clx3Lp5VOAk7Pkkgg046g6uDI+1d+eKfffnfy8QxwPXjmYVz+tbhXY3Gp
LsFNP86EjiGdo+xpEulPpL1vV5cFrYuhjexxvutUbmnR73iJiTuI+mID6sNYpH2l3ZvWeQoyB+Ri
wuU92oUpFzFcy5+uK1QtejOs8qgtBtlwLHmBpcujQwGsrWZB1zug4b+DyE9IYeWsRHwS+VhKBp9e
xxVa0Sy2QVxZpj4MPNCF8oq1mb7XEP9qQl6ugsfMl+l2FhSp6LGCuBJ76tLoaOezgq3oayy3ORrn
jwshnN1kTxvMbcgQvFCgO3LLzVltjodZFkWl5YM4P6zmvJjexj4PP83POiW6SI7XqfckewiW/SoV
FqEyft9g2aSZ3/tVzK0xJjVWK+diPtUg3sYmd1CJnqjcCnvdmY1h7GAX+pKRBbYIgLN+qnNJUoFc
rk9RU215S4DjXYrZt+0kibhrrQo0yuuX3MbQiRW2uITiOucJtUoZZFc8Pb2pqT/ZWBl7eonPHpYP
OT1BHUBNQAy1Nu/I24XQJwlN+UYteCbie80Ahm75evc4fzJ6TmmJF98DBmLfuCKgoAu/QqJiM80F
/JL4c741E4PJ2XtnSkDB7W0kHASGUM5G3gkatoYFe8DFBuPk23A+DZ1sRytvSR8YYh2Fui7gWk/r
mPemPVT/8xByAx6ut2dmYkOiOCFcGn5SMJm2RBpsqg0B3YpI4cQ756wNyDNfXrlr/GJGMhk74HQv
ybT67y5UmkLkMy46ZoDptEwFsGLz8rOKp9g/Jh/nYY5/ADdP/yhf2iMSB/iXBxVsD37JvPBwIHH4
jQZ+MFoaQK6E2FP2Am9VSE83w7Amhs20T9EJGZbdJh+RXriBikiPAjJHUTYeSJviEdBR3jpyNo8Q
19PnIaKQBV2d7hFkhGxU33NxwteRM8FVdADaf2nQtXLbYkFeu4yx4VasVkHJ2sgQ4GmQguDuVYOH
QR8TIbu4rvrlB1wKL10kj+aER2XWxi3hlhKvR2v+CSxDj/+wvBLubzZfsGjT+HQcVfwr92zexLMm
U/qVFDB92G6MiTQasUMGf0kPEFrLYD/vsglEHHTeIfWpvUxTKfM6/hRRJsxum90vJqA/GvpQFZd5
i+9uNzEVPfY3JnO0tvIKS4obEV1QY3H5qIAaYsc1MBTJxaw+mVN0Z8A2SEhZszRjPli2AzrgZkIP
Fi3qo2u3ffNmgJKvvYA+LJEIQGHLeJoXCGDfeUefeVhUGmF39S4lTzkpUy+l6dZ52+j5/aGjABpK
fbRsp+sFmn/w79pCaOPule5+LHDpdtmSp9pHCUvGZIzlqsCa62dPUzb5ffBoBj0UZUauN2dLD9EA
6brcdZVy9syg8/wqZ/g/Sgn6WeL7WVJnqJfa4gHtOMlj53dm22liZ3BCdlc3ZHVCkguHMC+Lu4l9
d94wu1BCT+7U3jAoO05cJKmICT+f5PL4GvMGRjcnPtWGLkcytVeaUvGTsLkyOB67nPl9l91fpvIL
4g9Wu22TeFdsMjSjkm6T+AK7yUOyE4mW9wBX+kkzhjbN5d00iuG6TZwjJS0oSlN3td6xAm5j5MwU
rMtZYp1eUEI3NzpzHpE2w9AsVYY1J93m68savjJdjdLJkw+1eDSlIaOEgya7O2Hgjjx+wkL7JyTU
niUhkracLwdQVLUWwi5sT4aGjpxwtI+9CJNYkh9+Z02L2j+l6yK4b6VVL98Q6HN4kBx2pctIu07D
mWVxPmWF37kiH1tZtFRO5zbdGDv8tqpWikyPlauKPEJtFW+lTc85V8aziHzwwuW/vEWsIDyVrVTA
YW9hyGLi4YtOJBjdWIaIDlt1LdcynXnA86kn6vwcQZ71ZwXWYk2TbD14bVFC3fv2kdDZ7z4XAIcb
ng8lj7WyyeCJmza38PHQzmU1ZRekFuE1DZ/pwg0O71w/Sl8rvs5cV2Q/yWfg2Bb643unVJOCpfOU
e2NX9NWMSf8doTEF9LeBtjsTXj4/mpZAFz/FlitIsTyvvOqNEV/De3OcI/Toe/C3+go4iw0b+mD4
dvkABOxEfbXyNq1zrVPHYZ/nWtZ577AUdCPrSABCwzmXRYehQUuppef78pyLlA1JOnNTVRE2OdfX
OdHtUL4NgW+duF3v9tMQ6/nZJ4aXzANwkKOjzVxRP91Y6QJGmfNcIREUeWhmPfvmyAQmV08LoeMm
SZwQGW5m7Eh9wGDF9fV6qrc+lSCbVjiLi3TPc5JU8NholMWFuDMsjibGghBicIg5tE06hba1sUxM
VyNQs81rD85qG9rwSFJ/GkuWlfoGlkoiNJvluBg7TUXvL5M9Ioj3SvX6GY21yPsgN3uZUW4dNWij
/asah4MRG2HYovaAFQEkOAKgnmrNt9TioOjgyWPeTX+xORqmuBDqrk4hNRQViikANNjcDQFjrnmR
aFHeJUDXCWxPBOIiDLKRbx5BKYOLtIHSAMogQBspmwpm5eXsv3kUvufedyFdAHBpHyVFz9v1YuzI
C0vD3uUZE/QGfOFvtp8oq4z1bEivlBG6TlxOPpiaEFu6u3rPljJnAUZC1Ruj0UEDsrUi115ayequ
iSyAXmvBJiWKa9rL2Ro9I6+h4LyObJpe0sqcPbGDM+4VE7pgnu5Ils/jpWZQIbS4m2T4cjPRPom2
Y4kPdVib10baSdrlInsEAHvkASgpIZOeLBAScFU/pelJuQw1jJz4xN8RL94fRt0yYelp9L5TfJIR
1Ujv6MtMO+2KYsU/sj/MkZN/bRHDUZ3AGMZ1ns9PPV+2OIuboiu2IzTZGiFyBK8VY3Alm15gheSg
iZaxU8WzAPcsbKCEq03kqz97b/NkmNqQlz5Up9zIlawTmXr6tWyw/Z4Vzu8A5ORqbYAgoUmJrgWD
pr7E2bg/Bwz3qFAqBo4dbG6pTp6yW+Tkbbdgzq6CNsYWua9lT79086/SCpGrR9hf5N3E/Iw7YY1/
bw++VM5Ity7c5vxLBN5QVeIY871ATkLFdkg2t0+PTl8bkix2X/rrjEKqq01HXeENQNWvljucwxSd
r7/9207Eyllp3AKeOwHOYT8lWLhs0fo54qQLgRkndaeGUVYxLod5TW9M79GphwUOex9LGsLJvE4T
7DuOE8UnEu54wJ1LZZc6qgaxuk2nyJtxOznPDKNEAmk7hR8VB8vgT6dZ5DkPhyA1ZLyezNz6Gbi2
hUIHI50Q47m6sXkMFpw7oKGbmyhihIroB3DQhkdhSAWuW5oax9/yGMdnqJFegN+qm7NivjI/lWmP
YklIxlWO9oxRO6DfMtTGES/L1Tlj7Warzi6pklX4Zj1f8JEQu7dIebZsiEc1+Pr0mxuTgrZSvsv1
m5SiMWTVxASbH4alfTk0AOhuCx0iP21jJVpWDDibDqmobT+2Hj2ZoC+iPjRBvncbuIIoNsOzoQiN
io5vKKaLVIZ6EYXRAiEiw3xfbedzayO3h/sW8IK+Y+v0cO5HhHh8+nUEzAEguDJrOyf6iAOG97mm
lFZtR49k7yUvrLFLMLEStih3Dpb1n6ZQxjLqf9HwPfLWxEiFsnH0/bj1xfBwEvZ8III3ow6+auy0
xAPkio6260DwIoFKAcfWTTv6nvAwZadEGyzR2cUTt93MgIfCPruSVbeaQCu4egqB0wEtENx+JFT7
VM3M8uDdU4mxtWFGpEfb6DoDJj4kcfEABrIyHdzl9btf+7ZIxLRbE2/tOYpIDdQPKcv0HFJusp76
tUri7xTky7mJ8viV8kVsL+l/K7OOJYG7oh7/8jTV0oz7+fh8B2BGRIB1gtiRm2TeqE04Dg5WjION
qUSKMnBOF0xUvI28S2zRQ/R6saPEkVovayQLPKk3YPdxIQ2T+jhjq5XyziwW/5dTEUUHYwD08q6b
uae01VqDHDWJbenwi0UhSHOMBU+hP/cuCl5pp/SXk0baZw510jciPvZk1qZ3ac7Rb88ZERqunlpj
2xc2MW8zhARitT6oY+4lDMQK//7zozFqyBz4MC0K7VcQwA7U6opVJSdaxrxH3hjgH5MUT17ZHWlU
f+Ehcbn9c+plM7+HEfHJddtOFma/gxsvVBN/O3fMRMHH6Qn802VyhiA2yKw9GQF/ajGMKhMrcVce
OHtPkJha3Cw5emD9S6mKQeqC9bzbK3zJXDhH/jTK923Gxdwv+nlUEPSM+/5Xmyn52gCHHJ2akP8l
5LWJ8ZvwsclsbrSzCrq4JVtUcpfkqy18e3WgOo6YcEVsoLrUdJISGRIq6lWy4tz7AsjCJccohk4y
2JWfiuRl+ERd5/cHjyO6b4k/AsQvrQxmSNw9Yf9rZmTl0MCcAS4oxM+s2zqBz5hhWrdJToTyW2pw
wNst3pKz2nLvJn6u7Xvz0Zw3KwUsMe9oZmL+iikclUauPcwswcudUfMHm5u7/Jd+9OenAwOWbE+o
deWNoq2Mjh4d31ARHsEMJdx61YoVi+psUA8qiC/4dFKIJCJiFuhH6yxOY1BYp6rHAc7dYIgdfl8g
nkte6cVJMKWFNMpyldXPiD+T2tOMNqRb2tPWpBGTt/GdCrNqXHNf/IapotRGG/PMKMrT//VMKE7E
DlvfWqC60nkH4M6o8RvHLeruOL0WT5ez+VbCtRF/gOvV0IIYsuTppSeBfO0tXAz5FUyrxRHi5+wL
dF09MHTmDH0U4xzcucOinC7ettnyzWA2PFBy6teXlHmqwZVL48zx78fzYEF5nTYXGeqCjrMFCrpB
OAATJLPVEfXcwHGveYeZULV1CGDe2s6FF/croCoVK5graedvLfRlRBdpV2QArAs3L0Uv7dBSP6Wn
rAHT4IZqh07uTM52bU7uMtlg8MVr8O4g/sAxmGH82OW/xTiMinFm4EJZAUg4zdertNJhIO7rzl0C
IFpeRthOiwzrvJHxpa+O0O+mhtxftLp1LWOtd3XVaLlkecMb2pJbmerp8YeH/EbkSS8pjj57KGMf
tPxF14rFWcMqTCvA1BnKC5QUo2y90CiC7xGPqI55B3sJ2g8JxiviyHzGDTnmGRK194V6t0HeGRRn
PR59T5SQs4M1FLXV4sJfzg+a+gTLZ3Je1lPG1n9M5Po+ZO2Nb/hYf5i5r/dlREQOIMbxlGI7Dy2H
/uvCQSfUYYLRLanDLdgutV47CPl44WusBDctqRPJIpdcX465E1WyR8gVFWVXwKxrFrVxb/ef7n0K
cGmSRD7e+cSOM72h6OkXQoatUnMobLRIGD8IqkTqAceBahImQ2bgaOVF+Mb42AeyGvJNG8uwaUMK
sk901lL7HipKzwehY2AubdUF3JxL91GhjcMw2FL8yLyvWpfpNKQ7shGKq8tbYI9FatNpVP/pQO5J
VF+MAc7nQUhtjmpw3g3d8RJ99unljhGnJv9Q2CQIqiAwbQHxIw5k8QAPoRlBQQYQ+BYqBV4QFVEw
Yp0+X1PGP4ZgPt8TsngLP0tVrjsJHlOQCc82fMP1sKmmAE4AXeyB358jzMG50EhYJ1GSt9VHPcTI
tf4OfePvrcQbiomuFRm6psFtLYlC5uZowZZrkU4MI7qyGNqPjUq1Xxmw3INQJX5YrQnVA5oKBynB
gLVICgZxIGyGEfCs8vxC5KdipwXFWi39xsHP3J3nD/xG1AMdeHS4gDZWggbDaUPeLNLnf5FiBRHY
ADFwrEmcnPXpM/BfoBfDNRxTXU426P+lCJw5kT4yAwaPQ7g4Mx3J6pFpGTdQbKAc6/CiV4A9hB8k
K9Ft+vKcllsz/PD8gOCctlkz/2jAvR5oeB4N8iKdMhDjZNHCjpJ/qYov7jvLoO+S3owpJGvm2Obq
oSH7sN5vnKex7wogWsiAJkiH7bBhL0LRiSsEgeyv/HiVbeHs9X/zuNQBSeJozabWtzAnDx41LBpG
OlnS6N0moKc5Ywo10ATp8l8HcQCZbRWbC3Zly0S51j+6HEyBqnjdVpwROaybje59pjSod44rqaqR
ItcjhQr1fIVdEWBF7NvxuhEP8CsnDqc+91exgp7HVqcqD0IZfVjj0L2o3I/9xKmQsQAc4+/WhuEE
kyCXzmEzqpDoUQFDyQhLdZ/Gkm85oadA6f9+AuBLKxokSkkP9dm8+AYN4doy37pvy0Cqr+debGmH
VWrS3CVIVl4s+ecCrJysEY5BtP/Abh58O2Fqw1JHkrDtQIWaDRAjID7Tp/xPc4fJUOA11uVOsqdf
W7Sl9qqgBCfbxGlHrI+LH5b3fNOMNWqxaMyxlV513KWfnvarHoMdaQ0APouC6vVFs0hQgq6r0guL
dtjRe+rnzXKIGNE8ybPomfDSTRnyzcz4XfZSYSKxpQvWfC3qnUYCqOSsPpB5KOGTIAXblBXVbabj
/VyzPh0plfquc7gyymbeXMozr2zF6ZxRCbXVkRtoIHNUmmL86jfhN7glCCRAOZEZbdFqMwgNZrr6
4k/pJh2FJJnXsdVKizbg0eq2SC93GKURHEQX9m1Sj1BjmwMDDbS+vXQqAHvRfTDlWdAQ46ZXIlY2
RJuu/VVs2/bAzVzdNFKfVkdpFTUTFpFRxagkSKaxf3iaH65e5aW5YyjJuQHmjKw3MPSyvfKYeY/1
tjmiswOIqt+aS1JuQ1TzyAJZcXmq1+j1v0K8p7HNG99UUkc7a7wOkjvk/gTmoIePEfB3Rz2rtk3n
dK3rVsm/xPvdtGjJW7YvcqjCQvoTFVo7jUTDX3jl39aFsxDiGEzWoWaOxBPWqXvHo0LNLlmuvh0b
tNM1K3+LxUomU2CvRg/0HEmep/E72PFDLp0MYlliniCRk2uvRK+TY0Y2Uok2/o9iVATK9MJoatDX
HDftCc+23bXmPOGAkfyp30K1AnA9WZLHljqX/UQLEVvjIRBmIbeaffmjtR8OhsdOOMfpHBAyUdZ8
zSs+lBj3op4tJkiJ364U3ptgBucCXkWc/R3jkL3ZNl1vDvv6WZxpkQdBhykPJVGfMpHkODk0xxQX
HRVQG5MNFWLSNDW1E6FUNwde+p2ZKwZaY5IR+gvXjQix8jncgs+Aja1tb9Xa4c8ZgFLqhszv6mVK
iOksfjW1rAWgsUf6Y0LGlzG98gGSLXCk++TfOc4jsedNKfR9l3YxWQ/0pjDpn+3t0JF9xVwUKQmS
58Y82d0/50a8TNSWK/PYY7u83/qJgRho2lnMembNm6nQEnweL2GBeldxBvaw3/+4Jqf8DichqYcN
xUQFFNA7wq13doWPnMruWyEToH8H/o+msT4oMMiLtxqJ7ED06ls7omDp8enjJFwwBdMFRtZQx06K
Gby29VbQAx3CuMOhf68+iuWbxmw+1CgWxofoMTpI9xweIEbmy5E1ba4PT0KrlgGrw5I0b/LpMMWZ
sbXMGwKYLX3Z7UCBOB8qZbEGh4XC14U21hx+zOjOY7Xe78RY8JRaSn8L6m4pKWVkU//NkhxdQTj9
ocuTNTVecQRSdHnUY7d0GhE15S8aoew+Nr9IbKAl7/dXQ6vHSPtEWC652s81L2gHiaX1btvglNvr
QRHARudDcJ/rkC8J5CCV7bwl+UrlGlmaIdYpDad2BmH0rF1p8iRsUEbTRVHtAR/x/0/hXCbu+rWR
tVW/Wkoka+gr/nw9zPRKadBYc6tW80RRRD0cynIVKaEks1YRIhoXetScRRAkkNw2oBhTYeyCt0o+
XafxP0j3qAAK7PSXPQv43wB8CgE0N8icNAn/1ulGVjk2fGmWpvWvoweZGJH7/6v0INoYQgP0YRKN
smszJWv3Ulu4l2njNmOh6sfV0nnaR5z9RdKzG+FgKf/lYJ6XpOu2SaUybwM5Unn3Ts894uZeQp6A
bkl0lEla0XhQU7YKs4SWD6R/42h0D/20y0csrsND7WEE1fSQSuc0+6kSyJhcK26HHgLa4lJvpwqu
rPJCI5dtmNfVMzbL37qXiX9t8GgFz1+G6f08eUASeinnbzItq0PF629zZ0MQPJprvUjKvk95NEYH
t0JlfTGAWGpA5Ud6wcmdYDM9133D6+plm7SBjyMPANvzWg6agnuZUeJJKsQ5KrroCyuh00oRrP7I
HDdABTPrkUBBAlAT+0kLVXsws7ezB7ik1TUx4y+J0dbuUg9jX9lE1GT6xJ24GwC6mT8MC3qVEqX7
8+2taK78lcukC5BfMDh2EM67d5M50K0MVbcWdSl1K3kfzkNKY0ONKFraoEGR/2wjczWQzczhWvwL
D7BJOKzvmApoGTiIXyCKCSq4UonPqYzZorAAaW8z4DTeGXU6/EqvEAMSYe9XAT8d4gXax9WayzzZ
Sut/+iYgoOk2pQq8sNAncN/B/swsbVh8Lozchi5KZk4eKOpaIUlvs7a4sT7MBKf5vkt3PruruIgH
shVgBBlsh1b0VDIaiMeGHifnw5nIeMkVcNN8pFMITc7RwpjbXvnwMuK1Wc2ZyhAxIAcWzQSXr94O
byacUpgMp4Zx0uGMLxGSua1lgi+AuL+uCVb7T33AB/yDElxW8Zg0x9A9RA44x83fkMoGwc7f2hC4
F4uvm8msCOh20h5WIFDfeiQLY/n6g0S6+xha52KlBDA9lIvyYvtBQ+Ir99Kb630crFLPpsCU/bBQ
v9kjhc0onQJQ2XUupAwownT2WbdMBBLueRc0/2h/bI0IoNneIybiEZZHTnMTe98J108Sy+vsKEp9
5UdLMakKzv27UDkNvcAnLwcukiAKv4j8HWwlW+epkFgaoVu2ZO6QmZQiShV4LEzlWfLvl0tFy59C
SSdSLoG68CSBPFe+PcEfGVmkjZj66x+zaf+WWHl+BAH11IVZUKeHj5K6tqpUcjiGGyLhtGIdhgnE
Ed8iW7yHMFiNzt3yePBZzgpVdFY1PjiNnvLjQ9AB5ZuMAtQwJ/aPUHb2I5hBFBle7i7ychWFUPD1
eFuuinwHH1zeopSCb2v11K4w+Khmjf+A6qkf5fWTYWDqO1IZ23PZ/NlhUKyu6s+2FQQAhOSwt53j
ZxtMxaKIze7vrPIFWXrA2uThS1wHeSzWZM3cyKHuu1U5Fzt3tlNY3pAxoq6vM9DBEBEkTjEaZC3k
puyQnIRTwDyfHqk118ZsMQv5CaGxW6TTtFcsNh55oiTCl6ardM6H8SvqTrWCNQtpp7UaOJyISYpI
iznWWp/1A+jOAvSUEF6nR4l4NISLCT8yQA0wrpV2klHyFrY/mSYDzRi3CWtDVAGX9vQ1MECPb296
4KoQ+ntP3Jh3BdIhqRDp80mz5ZKtRpcrOf0y+w3XrRCHe+b0yCBrPBB8M6K6awi6Asyr7QqL2wz6
fgdH2WtQZF207IatRa3Q/jMimhUBlqxMvS8jNtbrXB7d+dYZbjk5ppXoliQOdgHWNyMEfRnhVGtq
h2gVS8ClT2mHGdeh9xUcVPkowdLKXRaadmcK3tJiXyVkh2k6XCWNhD+ZGlMpFGuqYn7v344Jn5Jm
HBB4LdsvDDcCaLaDiY1VjcAodrxCky83qULaJOH41Kkd9zNCcuuqcGprfxiMMMWKSZzYVDEle4Nc
kHIVS3jMeMTWzOlP7Yc3iSgLad/zJV3oq9ncNZ4s8d98sDLACjuoUsCBLFiAXa7Y+8Con+MklZ3O
SRvFKe48vBtvfQFP5ZSnuNnfTJSrL4sa4fbQkWWmnfJ0cK4lhUzv0i/G1z3U5qBjGc4lnS8WjArQ
EHGNx0c293KbSpLbnJ0WvF3PUCNV7Qp7ISemAY2sXAKbxx6kcjGg16dM3EUq3vaElD1nrH0mkV6r
2jlrjWcJZYioayU9dbuqTp3aFcBIESW6IPZN6rJb63UsvBg30DHqP6HHbj7WaC4jGJahiEda6aqM
2PElMTjmfdrAD5MZwmpuKHVb5paN2GdTaw+QYNYPrjiSM0GG8QYMTu+nYEh0Z5nEgZ3LhgPIR9Rw
xqpWvc8lx26nPxuveR+FgQpNOe1uyYhia3uyUZuUh20HyVnlFM/lP95lf5Z2iDDLixAJsP23Bb8Q
HCUS5tBEtlv/8yKebJ6R+/OvVAtVYWMgb4A6S/DGA5vGMl3Md1PyYKFxSg3ai1sk3fUhcpwflTRn
ngNGUi3CtdLeJZrRFnXKSqlYNsi0k8rD8L3wC50+meSzQMqxSvHSEA7KygqWVO2CCGM3NRlwwmXI
KglOJLjm+VkN3Quf0LosJdH9Y6fYTkyUibGTnAeOhyrlVPvLqBvRTly4ssbGb29JKreCmYquwmsc
E+dQWSw65wvr0+iDAkY2C/wjP8SXirdSDL8njZ7b3sWVAsY130hcly82X7AZGqobBP6/3QRJF1iu
STMyDp7xh8M7NCMlEE3W++l6rVlr172ysmrrK+TQzhGnG7sIz6+4LOQgEDYZuIcdUWPfe1MztZ5L
wqueD6y/X0Glfnz2KOL5+oTuKobmYKjD+Cvz8Oedwm8B4EL49EzKPX5r7sv/8yFLPgQZEt3xYnaD
WNZB+9d4RvHpz1RjnJHSorrYURbZ3VmEB7i+RZulo7Y1MfNMVsc4Lr3rxg/1clrKX1z+QiNtVkcw
qozcaf/9D9VB3AUfatIl9A5/otuzcaq9Zb5mzS3V2zUfbfXZC9/v61BluC59vt7KR+brj1EP1Wg8
Hb9rsJpK+2XBEmICdAFH8ilECYg1ifuF8rLRjMsq5Ru9xTwAxG4L2EX3k43NE9WwH6WQk5AXTW40
I+7PrIfg+wB+RUpCeBKdM052kV9OxsuAW3LQvX7ZKsMpBGEvrdAPBYQPA3YB/KB4h36GEWcsY7KM
stgTnsDVVHRYenlWDzCkpaX+SQ0GA+cd4wssSMVApK93y2nRtkJDSxG0Ssy87Tmw9RLrs0jehsGs
MLtiJJIJRk9L6XnYz03nO49V5H6zIUhRqKw9eYu+3LqM/ZdGUrWlToqKoi8oDz5bCtArrQmgTuqq
uA1IM5VT4CGgKjD4RwuR1lR/vXhBi4cbq2+7DveTOu1jqNwwPrH2OgPoPXn9lqsoHQUVMRw4t4F7
BEPWJ1PaswVcYSEBvPTNTnlFrFEdxdXo/kJKrVIPhK1N+DHrkA2qbqhYBcsQEf99hmtz48FTFMRo
w/r/TBt+kyaMG2vRUaA1AlIZtdMIHdxO6i15V6d8bA7ivwKas3ZitZkPV79ug7IeRLGid4lw1iGV
uUecjahjl1+H6FDlygmUWp+Ho4Q6OBILbG7OX9mWbYCvAHJjQ1M++qkHCvyyMb8zWFs6hpzeR/kt
b774rUEkU1tMBI5h6Q7ehmuvBqvi51IjY6cCHWNUeqkkKTb6TQdIZt7pwZwfRdvG26GQGXhH01ew
+cHeReNfkkr0a8g/E8PVGr5Z8++RBpxoMIFJXk3WHvH/Ozexi8bo30hxFG2oNNnMCeWq/n3/vmP3
B+9IaFH6carnXIbWjsJTsZu/ZgTK+wQVNcpac+BjEC4S/H5P4o5QWAiVqW5LqX8Rs0TGpcEjs/4Z
H1jMGRmLcNwBbPOBmClTjEKFBXPGW30j3DC4NkMIbdrcVqtCBPOW3To0nsLatTWnOQdq5B63tAco
Cv429ViWDKtfedgqhcdpvrX2/v+GqtIJUPjKsNaS0Ep4ZiPRFrxuCJjnIP70OoJnXQpKb/UId3lz
bFn1AHhClZ8TEMMLojeykpj8raOw273B/spjFn4DKJMIbW3CTbF5jO5NWCb6U93vTiGKDmmYcEq3
3xYH0gZumzYhLrhMx/LZWEYHQ/4EFNZ0JeWy5ualzpLNuHd/vRQBfsrwiSDrjuBV30YZUq1msseP
ca8KmgtWcFK63iiRkCbGLWLzXrTIPxlYyQbqnkDlhBh0XAe81O3Vg+j4iTHYYjbJd2zn2bSc8ft1
fLKdebjiagAUEXTOqxqaHPUXTjZmLTUwo0CBRyjJO+RJYgFnOBmA6BWQSXmtBPbJwjtBgyu+Sr8s
SS863ME0kPC2Z0kTGHrAEeBSYaTGfnkqTIcvOijsb5+v8G2w7p6ZZh1swI+ZudKRbACPNy8ivxf4
h8bFFj8dpMwCTM6/JwWD3afy/AT0puCKXrgzZ2Dc66uXPv2vQQ49rkbgvO3loxrnVP82S/R5QK9g
V03mLKPN0OYOeimVhOfZE/4uOH+saXMLLUd+7XHGySO2TWmbYHYwDJUtjviTLuO1MPYIdBTRQlFS
6C0bQloQDU4i56ZEZ5OdhH5qk7urrscsm+awgXsmlM5OT0yrXPku04a2mf89Kwncs56FEoIQOwLy
vv6Q6guRacHL3uoQahejOml5hSEJJwT22oKxjlPLojykWBI54AZGPXFKVkiAShPN7I7wyMlBO04M
96VojNrmrlCQ4BsIhHHuO6rC9TQJtfh51mCHMavTGTBf4n7bOC/5PEaUwgZZ7OHChdbspSj3Mwtl
/E3Zr1+3ns2m4ZcC+oLRQg/YrOTcY4IrpCCt36PME5tbmL5PYspppxCKKDlPh83KRZNx245i8HxV
Oemmi0oybfqVvpW+LVZOF4u5+oNf8yN0yLr9Wc1DqveOf0D4Kt3DmusXvZ9udG8qsJRFCm2kd2SK
QaYof6xdoWRAhauenbBNPNUF1ZrO4v/bCaBT8jq0Z8IwsYhHUwj+iWe/afm2oZf5NcePO7SctkRG
R54J8adP27ysN04jtfT4ZlFsoojXTnrz3EnQRt8+WMt48xNWZm5qHgKXcbqWCmagdCRMtecDpuhl
4XX7QXsLix/Ae5DyNcx31yaSE0xW7Y8nrfr0BMgPXyTme1FJqR/AdLWFVLEH+pfNx9BbsYO/fHMd
5zplNJeVZmnebhYB4seF7GqKbRfXi9xuxizYQuR25JMLZBls1H1naS278GFNXoGUnGnjQOdyn0sS
LuqNEBLWM1Px/GeMIe9jppZbsT5Vvh9MTQoZGk2bSwRtAwu04oRCyWOlVFz4RaBRsRBy86wnwZox
/3uMw1cd5a9JfsV5hHeyBKyH68Sp3yfAlBTw4FmEnNHAlgilHCpZwPq45kzu5kEvI3uRrWUiIDaA
0Lt1ioYRxoXyi/0XqOasp2oyXePA8ivASY8QogsHheEp3wfL5VGj09YB14s24sDA4XWmieK0wXq4
TDBoGDCeEFum37dhg45RnUoT4ckToffmDYHC9lpXmEjwZEEt5VCNc56f94DbUjVD2enFvC/P9kJQ
voxeL7bfcv9HvUYzpCuoXZHYEv+RIW4JVUVz1ij+B3lZ+8gM6VMgdtXjMK7QHJ4CfigssHlSEovs
cssDzuY7IXqmYePw39XSExJecoXJHOYDmbo3yIUCDfgDGk/gH1Z3uqdUYfCnEYd8zS56QxYj6qQy
Xi4fMcQbpGzLd30mksonW9BE4YkbdoWT/JkCMzocFxtzKyxRny3wJewkIvAAvB42PpGE7iDP8v7R
1CbE1kiwmj9nblq3s9oXspuQGGni5WFxsdIkYG7mGNRThWLiR3ip96rK8pH2IWCg9ih0S5RmRNHT
48X3C0SUDfytYBC56KJvq1x5t9oAUJ8lAKSwwVtyNrznXxEUgG2y9FsTPVuSBLC29emrhSr8FlMM
eAT6jgOxBBb9GOLWRvqxV+O4D7ZynNTMAuw6b4tcSI1HYtTXsUGNRkA7wYewIQk+cT+bbc3zT/Mt
U6gazxvDbUGxsYI98ea9qQxgFa/Z1FkfNLEsejw3LCJ+RMthF3J608rd8Dxn1Riw9K3ab1wwSKx1
Dejj3fKZNE+f4AUFVjsadv+Dr9Cw32n3cORkhEUkUOQ+HLKXudAi3XtllXQTAfPc//9Cbt5X8QXe
b9ODGw1dOSylsrg6JlFDKLNfX5ArfOV1eJqktmUwlLdmddrrxAz7t1Ol+jp+34lhNILVLfqCA9R/
vgWX/oflH2/sepNzZeeBZjCJ6jk6CdzHEkIQzUF3GW/wu2TecjO178fxWuF5Hh3zKl7osdCQ4+k+
EbCU5S9gLQiwj2URXsDh7IB5rTLtTkgHYrO9MON1y+uUv2ww2Q4PiQBurG16jLW18fPp5ZMhkPxD
+oIWFFfhb6cnWIkiYRVKwmj19q8UwOmd9xIgujkObbFZ6Z235pUYr6rCI9ADv6EudBlQhm5HCyhB
AE1oHgyOo7Ce4id4B3/v/3RGy11CvkyvkG/qtvOcDlxKaPcYVx1XeexjfUErYIC7ucm2kBYBStkM
EZoUY5z+vOqTfOXrnb8QQdhu2psdumFJsrkEZvIc5JviZO4FN1Nx+Mnmg5bltIY7MvD304Md+UHm
P8/cncJMKqCB0AjBdNbn3Gy7aixaW+9QDUqP7/K0P+8U3FeUlC3fsUUV/h2s7Qy7e50Y4RMgU8iU
xWzPEZYG/y2ePYguHGT53AREdAY2UKNGVBPUFThhAvePq+vHgx4AOt+TGdAGkaaSUN7KG9RhMDpE
OTB+4gifmFOK+v7NtsPQEG1nG33CgFfoY4MeDEqohp55vjkzH5xYtt0JE6U6iMWQPGrGxQ0kb9Hh
L62Kme5gvLrBjoTi2jDHVKQfP4MlO0953ATOh8MAgFc6RfiDsGoLvcQdNyqjYivGX7BmnMcIeGkg
AR+CVDuFjhDWlFD67PLNoppMMrRv8t/h14Brdrn7IAHYc/o5ByYy099OErlQOiI1ezCpQaVCsYDE
sun7Dahs7cmHP7zFxv+rGWVPO4wueyvyXgm3cIxzAaqOJZXAIsvBCwgfdUVoP+2Tw6O0nVw8IThc
BVIzg1LVs2oZfovYEkefCELP9/X2ZVpLMJ2MP876RbQkm514ODnq8GcjEhmSgcQHkai9kOidia5y
qK7cq89JDl8Sx4pGmi2R8c6JhUxa3txejQJIcQB192iXWVWsJtBKkSbos1AbhNk2gGv7C/l4QTn0
5z1PR3D+Kahdom25hzExXfXoizJ7XPZOLUS1kK+a3NSLXH7MyOJR/NxH3a60ZFss9xLOiHFJ5jaq
5wqpsJv/nMYkgMjo3Gcxl62dDEGd5ljYyDJ77r2jRjY/GsgqKLlfEnZ70CgkMaCwvBjqStp5N7Ra
l3l62VO20l/+UPPadWa2emLmDBMtFI25CxhIO4nGQSiL91yVhNrQGsSZeJYFGtz9VCfG9jjc25QG
f/A7BKgDtfQGKbi2Suws1K3+8QZlxqQqUOnRn6TEEfpzUv8BYz2FMIfJwStSz6HKbYRgo8KMPWfd
/x5YdEzDHkHxSOz1t5vpBcVZX6ISx6eD/izwmtb+pAS7t7CkRbGdQP/xKap0APYHRBZP35x+vW8r
YA3bR0U39jzIedeQ9Abr3niv2KgDRcprMkXsEPqH39q2RWDXi7KaryIDnK/IeAIThR+hUuGD5/Z7
X5MZOM2fyhlfVBhnFBPAZFV4+3NUsS4T8Ivr8OlTYKedVfBLhN22rsaa9Mjy/T1AZE4IJ9LW4TsH
1KWfaPEwZ4YNaFEfeWPRApIumDdRdIOGMf7ZOX7swmfPKaXDWlEL/RI/e4xl1qz8UEo9g/WroW4f
lIDlqi4WZsEF4hy6EO+PMO9zk5JEjiDCfcrDVXPWZHxXUOzYFT4FTCCpHIfknH/7YJKW7/L86+xf
KO4qm1vhgtCdO9JWFA5Cwmz2QRwJFOP9Cj7cvDPN+mQ66m4O6tVYWRHg+jDbD1uddipy9kRC7/xX
7zrtT0KmOS3Pnryj3xbVn41ruKNPSm5wAQNIYwIOKFaCw1oNdDwgqF6P+zijsT0uH6ma7VMLGRUA
pak7WPeDfUEJ4vttotFdNW6EYNXmMka2/LOFbCHc2KTEBoPtRQwRngU/GEKm/Zhlm0iJS0Vf8W2K
JFQoG2gUJIy0WH2Cs3WU7PVjzuBpJa/TJQXWDZIN6HOlCSrZFBU2+wZIweCLwI5FyVDc+1SqvK35
fpttrN3i7bd3iNAydglSdegaZ7TfvRvXQx7452V9WDjtQBCN46gJIwdpanpAZC/auGjxDFlnDr6B
D3RVF24ni26GUUhHI5xZBMUhz1YypAVimjFFV7RmI/I9Al29UwFGyBmEHhD1vXu99PznkU34Xsby
TW78xFqNO3TsI7jRq4vd+FTTyZuApPGbkXfNP4Ywbnolg7wMGOF015nkLxSh/vasYQbB52Auxm1o
gL4+fUHjvQYCxwO54xUEvgFcDnAPLF3aswdLQddEh8Qljilo3FLQV2KENCExe/XriabCTfpKtyj4
kqhko2jc2nXmOr6vX6Ri+bqHGvvKKdD+4hoTXJng6nGCrOFMTihJitNks0cJ2kEh3lt4tXkvOJt9
TW+BnYElRwaNNAz6UNMk65+2QShOAJaJz2TqGDGIWD8CKfOclkiKVx84KXhKbidiNuXn6AlsT1VM
p4OsqyC/o39OJy/5jgW9am44/zuZpbGea/+pyVcL63tNakvJkg7syQX9a2XJ3sxJiskfQYDGjDtO
09P5G0Rv/pu1lx2ZFyhwqtBs5vjgyuvQ9jTUC7ZaNU8yw70GgMiStwyzSAsn1rRDAddeeNaplR96
+yL3bTu5GnbZ/vyoleO7lkZY6Rvhg806OQ1hqxEXpE0DqIWCasoxS1fOpTAPnbJIY3KrDGw8D/CS
3QTkR0U0VGBcNdds+ZBVnUodpb64bYjNK8EmreE3Cm4xH55gcbjZmatWlTKTiRPRk44NqBjB7UQD
QzCEwgMU6Q3bhv8LvFcbmokib223GGycMtMgYvycBgq3A3KDdtl1ICslxbRGYVGi9PRb8ufhY7Cc
cojL+9qyK/Lxr07hklUf26AkZpdcPSxm+IsWi9MfvLtUQCfvGG3+nkYQlIhM6XMYJXlDJga0ms+g
Pnw6RUrzOOfeEPFuQPvur5RE7zKkt+QtgVTmY9NwEfMSQsK9cH9g3OTpMrgpez6vXJM15aW6XwWV
pG9NGpXL2jj8jXTWUb31LJJVJvZALdZiBM6UzrdCcLgmWPoWVF0OCCJJiLGG4zQxbrLpYCOGkdVd
O178ctPcVjxdMFanvh32WCmCeYGf0m4XUFLpyzdtf+FdRMSyIY1SW+SqZ4dwpy9vPxc1Z7N2MM7B
8WOt+J5nB1207DPcjv0GEyJQ1PDPiHGQ5+MmWMJ+baKYecyJGoXzokZMCvdSpE+0OTGsaWaUF+3U
/FA8kobckr8GxXiVpCC/hN9aR6Tvv04zn3WzYTWTKBOel/aQfpcUs3fL1739LnCYY8aqruubzCbc
OpczvKJMkA2T9D0WEFpOPuOM2MGuG6G1DrkhdGYTxqN6q0tdBnUmKyOTftCtraX8jxFCFlGqRaxa
CfPl6uXzJ52lUMsU6v7/VWNcygOoAY5A8sRrU2MPITpa9oulLEkIiYgmyoKj+eIDbg1S7u2ClQT3
loY2ptQw+GMCTRuJXTK+c8hKWEsL2IC97OIrPfn7sAkedxg1cdKQnOSkgD4fTnL0ZuIWtk4Pbrt/
g49rW8NdFoCkJgQ+MKe91e/DYJAWpaX7jqnnNtv0E7Tu4cfWYIabd1+7aGVKmsYDGfd0QI+Xz0kn
BUbYvlIRC3SZsNJpb2+TYYZtfCvCWbC8jYavuedlB0x7DUjFU8kXN4gUflFDWqindvJ+gWRDRFpr
EYtroXycpiKsV2/fsG6ZMHguqauQtGKrTlsxtLkfxNaW2qal/T2tQkYjMDxzpu7IFxBXyUOjL94N
Vl/Tzl1g7cZt+XY74h1J6DtMnJokZRobMIehkNSY4WF4n7BrVWPzdGPIcqsuBWOvTDNy48jslWBQ
uthpsjq9Maw2DBbh+x5oDW2T3rrUiDPY2nJyamnqfdKhxqdqiw/pxeBWviFv98sZ5eBaghZQ7ssq
hT+W+DNOCxSm2bLZv00+/0LA9Oc+5B2qkxfcUqi3ge+JtvcS6TthOLY87kP6NSahe1sx9ksfukHq
a7EOXbKNgGFTMstKDoEb6BkdqDn/q9pAJ+Fc6TUjpND8E7mqXEg03e/wg08dFuUGldVvwpq++ohH
Gm6BYZTv61U+pGXkpQkhoo9ayCpV2dH/gCDIomXk9wlIvgNQ4ArV0ujHBZIK1UV7ta88bKFqfC7F
Rm2SfbpY+lJs3efqqM2Ti59vaDqUHUJ1rDbGQYiM0NvQDc0FmVnlSik5WGApqILql5uF6a3QtsUT
LqCVdWgURK43zesuO3QDeWNUO4DwHbmw9CEGTPfZud6fJ6xBwsf+BRsdFmFFRQ+FqR7tuYH8D19d
iPTm6JG5HT7+w8fCK1E34PZQrgFC0eKS3SDhKCYCB0ZK+WiSVPlu6Lee8ZUdiyoUj9V8C//p7wUP
eS4vuuRaU864n4qsGao1NmIVIfqDxh+3dfPRiasxBUTCy6dlO7hII1HF5D+UfOzP7WG2JZn/dsJE
vEGapJ8BBs34l0GmNfDt9QEusS2ESNKRvXZ9eA6Wa5v+I2sZSrVlwuAQdrGAByIL1yozHdQItIpz
/OVvDrJhuNyQuKn3km0LZ7qQAIYQFnPRFmeQVlAuSbbu8emFbaPIsDaDAZwhWCCU/Gg04WXDrbnK
w3d6/E1ySW/JqXl5pAhhhOLs3giMAp8sItV/FpU7WTZwlr9vqCU1DJV3kqzbcgKCJHCYo+7CqSL6
yqDCJi/gKRmtvgiyMKunBQCuGAABw47sZJhe5MGKSULhlNu0W7ihSZb+rSML2iLLyMyjBUWr/Xmn
tHgQDh8+fv0NPThcOFwRrNieB45yOxF0z5JnwgsfUeBz9j2daixfA297z2NrPXuZ0wYYOSzRnkss
u5HKBz/i8fOJFxX8YY9x6+U8GFzH5ilgXVfMD8cv+f+hok9dZHn6bY+lDjhYPYMZtqYrE9aTAWVS
foZNCS3STQmQkcPEB59sMVf1UIx97AHK9X+vcY4Jzsl2s2CgUUwX01ZQinbWWrukCfRj8CKiEwcm
B7G/Gp9qGxd5Zo+nmxQIgAeF9m72c2eLqUdx5MWXqzmTEuFZNcvNuIZ/BMRcszbimSy8TTBQPIPF
69Kuo/FRUA3ltsW4K7rgw4A1dv6jBplHt3RUT9eKJAV36LonqrtE+2XBevo9qhDK2ifLCq5Bp+0j
KuIXWacuIdCEswDudim4iw/xHIb+oYGf64Hh8CTCSGUDpd0phLOxt0XelretbqiJWnyFV5wUzEFF
PN73UaEJ2F2h/YrKU/fmsVffKao/sZOtMuwHW2AKdqocsgTntchDm2pjBSZ8hYqlAAiJxYsrjb5u
UCclMfPQjIc5QqqWsghebLkDCdskLl+2OYSJGV7R9NgsxEO1Rhr302DM5YxCexcVOW/or6VPBMLS
2i8hbP0Mf/KIYzAH3srD3mVuhUQU1tkpMMMw+26zgX7sPER6vzZR0e6zfBodU4bKrwLvc2dUVvzz
13tZ9TUPt0u0uMDsbZFBhUKoHkOZ7scAoFAFE6DhB/zEZPuf/0eifVCrKq/9w0DnHwDAtzYfN3pq
9XGy7W+B4X+OU34y4etj6nrg5b2FVfSgz2MqgQoY6knEyhivFeZ6t1PZY/XzbFND/Y4RVtxELllI
dO2af9XnQCSL2Aeo+O1dQAvGyCDAcaXOefVCLTF5C2jBmSPZ89m7YsQuXAVrw7MPX25xsZ1x82U/
NCIWpwWPxY0ntdg89PLwvx1POdZe4MjPWEW8CV/AQyNhWH0LVxyRQr+ST5LSDgydDW0RysJ9oj06
zZxP/63DANkavL1bxGJtEpsyiLzI8o6LLA0rEg9cc2esr98pSaNMll59RQeLWPKjA8tNc7+gNP+t
sH7y9kobPiLPP2iARLOJ0yHbDtHmAjrbZiG5u6OQZgWlp6jb/xWlovASD33gV5ilt2PoTmwGEQ0J
2EzLz8W2nFNUqgwloyFRMm2oMMaapFYhYavmIYxMz1QLEUsX552wG1L5BoNNUtF6y12K0/WDwsuG
iIK8ffn9Oml85E4qCX1S+EVbEYPQlvD1PpkgL5uSVQJSVpX0ayM+GsJrsR5n/BVf6WnNhDPh4xQJ
rUrk/ONr9doZbJlGEaBUqG32pRRrV/xli83FovxtNw7lQXNWSiXak68FVEn4X++5xHOGUeWf6L0o
on7OYLgCXzlFuPZrC1FqDXOdQxWx8zAANCbbJW/XA2U9UKur3+LmGe5ST4BtDAADT23XKJSuiS8C
1IiIoyG9Crqrq8eiAwlAC80JMPmcEnjSJ+ku4rSPATV6PtZnQhviq1qdklk9csSp/CW3vMP4PrCi
NNSJ/5bmcXJSA/SX4AiZ3PNEFkvRlCKQk9J6KqOHA7pQslF7b9EgGftI4RIUEljs1ZfeOEj5wBym
Jug8UmFcJ4Hl1npdHDPVhVimnO3U6L04wNcCOS/FqlxKLMgaAvN1D0sT0eJmZkgXNgfUEJF9w9Fj
3WshfcSdcvflfsKPH6Wtl7fa+p1/Y3nYvDEl/Ap0e5LOk5UFVlocR+D1DUgS3auqewtEqzOh/zHI
u89AE4UVfq9uuK9aLTDpgVmfSKQZs+e2aZUEbOtEBmdVXxq9t2hfiWnDOePJR1WBZ6rwUCthyjbT
g3lAg+bcTp7hMLBdA4lt7po0EvWKqr0Gjw97Tc963NL3Cd49DM8wWkGoU3jQQULUIl2HMOJ08Qy5
EVyb8BbN4lNfc05a6mULS1qmhyNhmM4U7FphDg90gudrFuAHE5s8U5IpR0HbM7GJJyowUDZPLYur
yzfmhsJmzReJ2Mq9G+ErEX69+McW/iGB8k1+62EMpONlXaGnKJVdZ/VV9tALKFEHAF/DA80DdinH
cesr2mwUiaCqS3nRvxeVTJTU0fqqHdrKu2fy5x8IeF54ZGijAfbSbLfCpzhMAOg6yjFmb3ZLqyvF
ydMY9EI85Doea6MCzqGABidI8rnXCtxUo40WIUv3uoub94zKEtxVCW7ImmMcGMAa+XZE0rfIyJD/
hKWx6oIbx0UsMDEWKa5g6BLXCP5LLX19yi+vu/tM5d2Jho6hZXB183diuw3wuzTgTlsZbo6w+n5N
24Vzm78AW6p4NRpGRvuudUDCQRcM4FhJ4eTJsT17zCsgl+TiJqlRPIFbLdRKFB/VMctioDV3qvNs
ZiGaJzJ1++1AtpxwL2Jl1biDxccrF7BQPhXvM42egkE23n6SjS1m9zlOiGcR+5UtDQ2rSk8ZE1dy
lWcuoe0eddR8zVU/2TZudaUubdObtw/oBbB4kGvNwlM8N6QFEQuLv4ZvA5e5SuINANQkUXW0istt
mg1ZOQaSM/ZuxUcRxYxNjCLzKwhmowR4FDMnrM7BB/BPqMFoTxw9UTXsXLwd7wX0CuBKw5dGGs7R
GoPZJJTO2Nf5F7GRCkOFyQXFsa9oo3EhM0hd+nSPOVVH3CFjNq2IQvoKKp+bHy3+B/edaUUCQEQA
tTw1B7pCpzPTeyLud5I3JCOyU2/ZD7qlXRyvafvj5CRr5t+QNHAaVDHQIk6krfLLNjRtxEvAgpaz
hM/44jH8KOUEFMB6IJ9pHp1Vc/JqJHlCd32+i4hIvrw8reyRowVHdk6TvO5a9NHDxHyk6STZtGTQ
stFgFYEDA/Hwq8dsNmx/asK9dUdSf9j+hpboGm+GYbOhVcmoJFiynBJpsbqIg/cdHk/r5Odb1gFm
tV3xODJL79ITG1KG8SkURfcwP2FcdYkv5oiuwhGJYVH/DIwg/aHTfEsovAJ8GPIBPHTx3hCo/pAf
HagVCIykw6SCDMDxY5GYZKgW3fhbZsxIwpvY2HvWSMfgbXQi+sDeuAbRPAq8MQiZBVTZqK/hYx+V
N2Fxdl9QKAToQ+Ll7A9sPDxp3I9Gw9N6cH12KDWuzs3uX8K6JyRayUVahK5vPXuk5DN4VsjT9dG0
uh7qJJz/E6XuahOWp3DPDqpGki6H8D/7gZB51/E+0m83UW4IdwX/9moN15hd+emN+12EjpSvh3Hu
0bxEaLTzjTvM0gJYxYXjuE6AqYQVYkqYGZ8/KZFOKoXqCNOemSudjEI6a928WKNL2FWrPq/ONrKT
1ZszCkELxkL7ZqGZ2FhyvFMGeLZA3dUJ3vKSHPrtNoQv8Ax4VEiwSQzQAR1y8uw8SUSw6Gv/mfFu
V41whnp6WEkaDsn+JLT2mf081NJnJ4yKKl9HftY7InJ6HyWiC5uIqWAVWtpKujd0N1Eh6B5eGsYz
aWcoXpSB3sOOxQq7xcZO6rddbd8qdJ8phft87EO6A2Esj/5sNzitwbEVl7JD1oHDdPP9N2rv3BiL
QiW8OfIy2W/RLQyIZCQyVXSCBpeTSd2nX03ot3viSX7I9gC/sByMs4B7NZmBQ0sEnL60mA32xSlB
uc2j7Ce9TFW7rY6V9j04UR0k4pino5kxS9pAa21w3ApHo7C2pJZ9WLbfcrkpRqoKMA0m3iyU+zTw
FqUwjzcyJG8nbeNIN49zTb7yqjeU3H+LczkRbZDrYaVd8pPxVMS6TF+4v6PfdZB/e7Yg9x+1bXwM
uYqK/XLQNC7M9ppGkKybWWBkKvYBWRJmKkDXNkEQ6aiJSKUnc1SS9CKxwSchsLEU2tpCwFfGYBHU
vSIwsAPdPAvqqzlT0YMkuoSrI9UvfF4PjOFS3yoNPvYUe57qfTn0IAF3G2hWcLU1pQvTIE91fCqh
DTMThBii1pvQOwXJsmi6pmD6/DzQo2baYU7a31fyB25NjiJw6UG+S7WEfMi/v7zeEuhvpZhGOCtG
8W7qWo2ORng5hdSGDhFsOjUFjdUNkBFLpoXmbFoleJmE9iab1HrvWScdIoGzPVPKOOHRa/cuk5oJ
CYqAr0O1ud7ZvA00z8YSVhf8h/A1J4Q0FF7aGTrAKXtTlr4w0UDMP2A9eZORopGGDFQ+PHGKhAbs
Hek+IXx1SSSDKp+rHaVCHF3sxImUWIKfgM0vq4porkFv4PhGYGnvsoJ4B4jtAIFH8hW0w7V7thOf
h6p/61jakNDKKdS03pwElwvcQU2xBECzWAPTbKVCJlrV3qYDDQ+PGf5Hbsnw4epkXjl51m3R1urc
we6peoa2wMEPpcbaf64AtQPqvz3jY4vEqSm9BmLCscQcCuz9WkA0Y7euRYB1ebPU7vVKV0OLHy3D
EZWhmgXEadapi/etQlMMRoNqX7JQI3bo1QTcGbTuPflQe5S2v2zGe98m8rCON8boXM/eg/hlpq7R
1eLTuBZc9d6b0DLUhOcZvvwKmH2BMBDWl4MB6cnmuDjQi77Qe4Ct+ZwXb6nfDIz/+Vn+8U3I7dLO
j+0n1J1VUySd0HcSW0hScPqwrWN3HbtzWhjlBYE58ulnWmUXfOwL87lc+Ftg6OujWfs1lKeovLUX
KA+vTneQmYp+GlRwEVkrU1s8Q8jIiqFVdm0FFolFbLTh3QLZbxsDyoHIYDtVdIzEHX2pRYtksUn0
8xbC9fz8MH4/f1E1MCIsRmAf5SmCPyE0Ts4O4ixK4brBjkM8HvBFzVQLbAbOJXRYGESynWt/8/ZW
HO7Vr3uaRnbAt7/fcYZM6cCX1bdgKhnfHfMkal6oTC+iTnvOvQ7LPCXXzMaZtLyS9MtjzVtMdhyp
Y5RJSfawtLWhkAJEdFuqdqoJ1hcF8D3oZP1I5FssiDQqjcjt0Tt4+vZEMa1kj1zkVxV4aFEdDknW
kwoOkNLraDruI3WyokGBm79TnvPYMbSqC7rFGczQMq6cxsofckcKrRnihjGizREdiqFxOGAMDFgM
5iyfD6JBgzV8Ff+5Wn4FBjHZuUFgKEzOVhFme6tkepa7jbDv3x7b7/FA6O7MAnkvX9XaNNWF89wN
KRc1hwddJ6GOm8BVC+5+N1ect1YkqpzDCWSQJSmkgzugrS/yu9bx+oFNVcQfDQApxRxIVXSeY5s0
cpKW9yGPNhCoEdJf9wmCvGHIWRtqprKS9W0j/YzxAbxLJHCxXZDhsJvvaeWjXQf/VXoNCZ4kByxt
mnRquIxQfTKLuZEMRIkKOOFo/qNzxh1r601WuDJLptVdnIe2FveawSRNt2zf8cysNZ+hQiFLCZlO
a76LZbdBgqUc4gz2apRdHJE+fMIkOXdjeQ6iGPADRWLQwiINibAyPjvFTcm2026LJ7x/9tv0BqWe
nXf0ZKVrfUSMEQajaMzzjmPC6YAYZXLOE9KHP72RI80XIdhejERm7SdJLrSDvC7PMXDWt8bMHfZe
pEYXn/uAhsFnjBQFiiTD36TDxKpXmyN4sS9BqLjKcMV8rWDgHuId14t+X4WDXKsecpYkBXQbgIVD
M9llFn9rwuVfskCu9ur3kb9GqwTQ65Hb26cmPQydPQkJNkN3+mHnGoS2W1s7V66MgvYthgM+otlY
wQF86IB4qetiRHtC7IDcOzdogt8eFP9DqGPtZ5j/1SgzHEDls42n3NA2fprOHxI0a6gsPyXAmqem
/WhUqRCVq1/gRhNInr7HdePjdBc/KSE2D+TE2hJ38lfWo1/ytpHU60WMGQNWaZX5TLTlhYgVe/XF
HHH/AeoWw9MbYuW2OVha5TzRqoeHuUl0QpD4qDMHcsUjvzlc5aRzMDCqKe8Eg0fwp+jQd1GHPn3s
Oc6Bib5pLvwcJt1cDrjiGMmeWXuoGbt8gouxVYpLv/AETgN9vWcckvwMi3WRH24/hTpRWJ4CwYI1
1vta/XtsgQnoj9DQrVX4KNVUzDoZAGLcmbXQA8PYZns38wrggFNnvd94R2Kh5HPWsKIbS9rAzydO
0s2KdQbwE+My5GIvOPyl4+OBrmqbR3W3ck+1Gr/QtHi+fhyOi47FP8uQowvIOEZ1GpeWWbzIhu9L
oZfLnPfu+0hr+leGK4Sln+n7gkbczNVNLyIeSx/f5v5iz2PZC+6VL+pg2DAMTn1jjA/PHO8FkSb4
4nbXq7IphNSBZZdTpYIvjsI8Q8oi+M3e9wSnhE0neiOjJcIk+RNE/oMwdqSncdvmtYho/C8G0PjO
lcaUPTtZdPi59GRCdLqfEl5YKcbeeIcY31iwFUpeRYe9UEFVdGn2DR8aoDaLVmVNdH6PVbEJM1O6
O1EamSzavt1QopCAGEF1FPA42FW3qo++4dbBVsax+AnB6OjcFHHtr3HM29yb3EMTwmfXz/Ua2Cfb
XedQnAVqeuC+/KbZA+ufBCD3/ATjG0MdIjjIetH0Om1Kf3adhEW+zbWH6u5ZdyCj6KWy7Sag6b2Y
ZPHcvtliu1ON55nT+gckF/cwsHg71ZCzDzFva8+bErW+YQ58F3ho7CDnAxpuetyVxvMtVB0YqOcx
uK/ETIB0TTEXYLQZ9vKaUUXOYaVrf88Rlk9VGdtxPendJE7za/uY+sV9ZZqPTur5ejCj13tp7j28
jmJTegRoFHPfH+ebDHFEJ17uW9XEqwdUR0OH3hWJRC3l8W+atPPdN/ANfmYp2RqeQ5/H2GlScJHC
qAr/egTu2rtYo4bI+lUbHSeynSXDG0AhFseKMmFMmhSFh5ZiDLkSqR5s1gWmaevVorlaJhtQjFQ3
qbsgSi2aOmpsRq7x9qoCiwX+JOb1/ReXa6kXC6H9MCjiRFvP+PMD0DMXDJLScEe3yVg8NZmrUr7t
zNy3fVIVQwPvi46bWiVaS71ZLEL76nJAssU6NPClLlxjdW0o6y0N4n03cGZcwLcr+kjLr/HnyMLa
Aw667FoWLeAH2smjhdBQacZ+6iWGaOL5DdfgAHVeDi7qtuxgUaGMgwgetj68I0E48oVw2x2ABO48
8GKZMiOT1TBc3xpb3tDxZ1HoIJfEQQ9OedU76GAYr5x80Du+U/f01pMT0tmeW4s0jSLmWxXA/+l3
tPIcchW3bRNiguieNkTcibYzLY3icAMKiEfarMfFekmpKOyDziWVVhqAkDZxmcNpkCBixJZZwChL
XXom44DCxPY78c7OHnmWXBXCLFUFfKBIMYUiajH9+a6z4ShmZzgIm/4FPDO8Ouh3KndYod9fHX+r
RZCRJey4A91fe8Rzy1rLeI6JYluC+iMnXsqZ/yMd9GIo3Pc50+udS7XS8YV4SKMgPH3xEMk9uh6a
o1Dsuq43fbVF+fO0qU0HDVx2nxgUGhE46LnFrTGtyIkzLoVT5YF4Y0O7aTO1vPe3t62B1bApfhn+
C7325DGEebsSaTcJw085XN1bDNrBbcCLxA5tMcpBZcAy6FT7sr92usocTK3604P7xqCjm5PyYpJf
Iht6ihOc1HZTDdzyX3QN4k5g+Uw8fkfZlwJPtQOKaTPmg183qg0EPsl4nowYXJA+C2MfsV+/TI9C
kyby9PNWHzIp+6QbM5I02uZR2fAMu6z1gpf9G0AbQ9rICF0PjGFTwZfbAomWUK2DmLck6q8s0p9h
V0IzypUvVlkr2DGzWjGUnScRRc1yzuccwC0sYOtI8BVh0xKC9DYpap2no+tkdqgqimKOxSzJfybg
Y575Q6wyhoqWnb+MfO1QCxWLlN4Ul0T8DcjqBzeYEGyMfnafEosfnb6ip9NREbHGKmGzQOe3Dxuy
uO4OUi9knPgdT8tigL3nSwrikeogBM+mVlsxXBzcYj2sqHfUFWItRAsPDdlL0pNDSCJsYRL2l8tV
bYmtI91Z8pyFhveJjlk140DB9xXd40083p5r+FXghIuPsmL8u6zdbqLvcfKoFNmTFkQDespAbI+4
7HZDI70YI0n1Hl36NZpP5irQPnd16VBYyOFMaWONrVB18Yw6SBBrpsgbz3q0O1iwgzN+J6AM+pNS
xu3jFHTGElbvjnz0IcfvPDzU3mkbS+v3On1EBr3zp+j0oksxHO90p9ypUxeNQP3C2ah6y1179Pxk
wNr//7GwA1p4rVMNGhQj8THYaf+qKl+RbjJFgMuKFMBk3KqUklK0S2bbDwlK+4DUDXef13QTGeqY
IvOzVT53+eIXFA+DO8tDScKLb45YXnlEebpMgWXXdEfktdNDqjbGbc+ifXVpijJTeTmxdpkzq1OP
JSBt2dPPVgCGHSACimgaHpZ0bzIURBy2REzlUrwivuBhxQzyS9xiu0PurbugsIWGmtJGmv/LQnSF
ZY0y5IHDhWDawVsAtnpuFwpPj+T6jRJ6SAUm7vFm5rCE3PLCnBa8CZ0u18Ud81LMgvqOdjj5bJW9
UbCUjTcqzvYt9HUna6qAayefJR+VIFBFkJ1ilFrufYWL36f82l6V44rbMveDXfAI/aRsxbFB7Ksv
sjyIk0HfeeIZ+QvRk8UhObZUohdHe9w2s1U4hXxe6L6OE3GFIPSGAHPJbp0TMZgGSy/gvMR4pUXu
V7VGaX8t7pgChxzGVVlOF9jXJRkwDP/iofcQzbl4izvOldw6/VLoE4qmzOoPvOzimkFHahixS/1U
GM97heMo7PK2uub26YyDLi+s9QU1bSG5HxMOgMcgIqrRlp4KeAIVlumiIZtQ/Da2a3ArcJtkjfcC
rz/Sa3wpREZOJsY7Y02z+gy7Gp2gV9/UFaQ4RKV1aH8V557F4p61rRgkefDeXFsIxgzw8T1Jy5eb
gRvbeMB8UKF0+JpZgp0KcI7z6cvSoPgbP5R2YS3XiDmcO1a5DxBZXaX7mZE/2RL7BYH6p08gqNjR
sLhJP3twC7LmzSyh+x1H34sQpUnMvDYSP2wcz8Y6xFBdfQM8McsVO3Ysqy6z2NJFdF2rsi1qYxcn
j1Y4qGQ4Re6Bp7z89sH5uH2x6xAW7rdd0NXmsvgNHz6aA9pZ5EK2kDK3GwDm7QmJy40/fL3Ofyxm
Nh7H/qcdQwAw6PBYZ0GVEoFnISiL30Q4FlAvOYGC6C6qAGkGRflCtOi68mOxTicx+rzlAYGftrCR
lW9eArCYFmXxmNrOIVJiSmNbh1bhUUAWHB6I3zZdSvpkPI77/Dl97z/EEIRr8OoINLyeGm60UeWS
8nWofi64zPO0TfcSIyzPcDQmrpM+xwmLC1IN22LGxfFRm4mzIbc+XL+q212VB6JQzJfjRqliURxn
EeKwK2QnSZkZBMi5OHuO6YdNeDIrgfGCMkb+EPWVDXPOzyUImK3m/2lI3m1xdXCCVsZyxw2ukYlh
cIUK6TF7U+7rlw2V/EgyxIyCA09WgV7ErDEXViUunGq5n2HHK9xkplWIspf+8nSKtb9c9xNOuMf6
xE70RNxCTWm5EazfcjdKySRS1gYOYIEtBfFMj3+5GwaQuFRd16Wf7SqM0LyXeNYyIJVSfjAm9A9S
Otmo/z/CZw1bhsp32A4dhHsZCyD8VNvA4wPlwBcKdE5OvbIcoqh0GJIKdxCn2f0bclpR95VQ3BdU
/3Ku5aawjTfFbJnQ14Qib4xSpgJt1LGdkJjf4eumM7N9K5Ex2uL/XaPs0dYo5e7c2FpSFOT347Us
AGASblczJfoweIsYPkxKXXa2oGhZjqUMQDEoyj+bhB/ONggJfYR2jIqXdxLK5XHT6x70cBOP3pIj
/nguk8WEe9NDspYindTS9aAliM1lN4+n03qVBjdikVO8U57stBOCB3vWq9JtvAH4zToRGdzKINJb
meX3JvfYrDJh9Q9vRROtVdShHq5kkv0RosLmq1rzS4Q5RBgliRayGmrafBY6nuRAsHSZbV7A7qn6
kZSkEeWMCPQPbuIyrzvfkm0IUYNkGnt7RWTHQY07svnWGWKQ08q6TYaR0HVdm+PCi9dadGjIPvDu
6Af9jgCucQ2ZnXz7QSV50VVajJrrAeJaYW995rX7J9PG2Ptg3eHGQu5bE48yk4Zcbl44kGlNoXnr
uKY+oD4EZj3/or3ho5PNTGykFB8vc1PYngg7EPLFHdysObKFdC2qVD4qcG1MyoxgDiIie6MzZt9u
f/L6rGxuHmg0PnR/tmdlzgRV9P9pxaT/h5BSQw6x/FOZoHQos0b3ux2UgHH4ByTMBZkO7xN/+7mN
xuGLXMDEgzZTtoRCpmowSuF+wNZZ+rxx1EJ1ojELvIFkLfWiKZoVoeMz4FzLSzhBjAsnxpBqgYmk
sCM2BtDCMye5K/C4FkwAESyxgLp3rOWQr+B6unbuPdl2Uo8jxbP0FPxHpwDObxjHmvEuUtwvM/t6
KbcnT7Z2JJ8bFFvU0WX0RH6Q27EneTSVciTb77Nr6OXx5D/Avmc9lFfYBP0JXFOT+5lwHMp3wJUu
/g5q9VIvfC4O2xyqrqKAjTu+KfgwqT+GaRd1NMojwB9tzqYxzmspvyt5xSD5o6u9eMcXo1sqovFp
LS8x/uQmlgy4Mwjnutx2lMEaHWhvNUbpZInkLP6AUJx+lP0BM8uuU+nki40WkxhiJ+uXR5iQAUF/
Hzr7FxdlZJgX1kqXH4lbVDahP35wzW93xP4Pbj+ATB9D39O5Y1uOnXc2k6kR4Lzpnibhv46KLp18
+Yxt2Ck07XRKWXRZpg3h5olUZqcbmpntdopFUjE3/FXi3O4kA2r82siRXzgaaCc4NXMEicZ03kcR
J0l+TxlXmvVr68TjKc9DUGoT3/pe+WoZ98vj6t36o+FTv/hHk+hhxebtKOsfccZZADFt3D8iTtye
eeNU7HI0TXmASHtnitxBzClgCwWY6xO8vCUJBSQScZj68VbeJbEYuGZsH5BOtAhylWDDL9kHRfGn
jfHgRFB1FEXvUi9Pk98svuUBHw3+pxozPbScciNKPpxdlVUFkd0Ve0LvOyyZP7/s9aY4Oag4HOOE
TvAftv4NOIz6G6gaefgF5GwgafCbr76E9Qc9GJQSrpvJhQSiX2ylcYT2d8TTHwFKsCC3VnS9nnip
V8RZESVkvwmkH1OaHOeYdUTQKQnH+kcIyLM0TY8S+M422tLwN9jnaSJbO7Gs8TWjrJx41Lk3O2rM
lLUQZPYZBQmFtelDldkmFz+KZZKh3+bEQGY4PUvq4L+07U50/pygAwYrwN0Wv38ndxBqSsVq5I+x
h4y66ThQFwpd4onhb/ni49PjmoajDmv6iiwq0wh+VQefR18RaGuzk4EDvTOwz62ne1g/hcPlcx+9
gwRC9YqBkyCzUK/oSq6wbtBME0Z3+VmdE0OAqL51i20otZEqx6t1uMsOq090GQNaq+VRNvr8Y1OT
MvL2E754zKqoUQWV0doJaGQPrtQSJ3nxIzD1IkW2ZFwH6laKDSwB3F3j/4F11Hl5uK7WltQMJZl7
OJgx7vioXx8Is3M8unEBd/dHS3uvzBwluemoGV7moRktFghn8I4xl7E+8p1GpVGM3uw4MbUYAT4T
tP5YuAklCCdXPY4Z3RcihCYPrUQ6hq4T5az9kIbfCNtdHEwWITg0Lq6CY8wyktF9sIiubJIX1Kgl
EwxXJGPPN+mt4bRYaMyI65KSGUvh13p2OGd99nQ3etrUtuYHMJ3Zi+3PH9rYrbhq67UF15oNIM52
zVCh/lK6PCbo0WaxVUvmLkmIuGK2ui8XmXrigNNv/MJxEPFdSf3LK2+J+I+xDdEOqdzttkHAMpnH
ffLKD5hwfUxt5nU7b0UprhaChlZaT1oD7LA+XZ5AaluqD9RWVdPYlXpszdu54CJIUbKPGyDSr8pn
RXx68eCMxYSQQgSNq45+EaBvHzo6PiSSBFUbxcprVJhK5sjqkWNH8eQrEO/aalPinV3mWFc/57Fz
eCPoxe3wrDR2YgL6XilyMYQhhasa5BlQxMZYAlXEOCULONBJKqYyZyh60hXagdS4/kdBuIAUNAA0
k8oSu9VuyY4OjRM6KdZtl8dCi0OYDwiTNjmCLEMOLJ2E67MCJVXE/evcqISuVVtEq78SeiN7Bfvo
r19BHElyl4Kg7pXGF7ZVKYDNnroEAy4ZlAcVIzFCEImRN5k2MpgQgdGF2FuZshnymhJ/tzUYseKD
RnyCW0KCq8W0oVi1Sc1pkqaEf+DZEd3b8v++YXibOPlLm80oGxsS349roVlSzSiXVQmezPBAWa3h
QsSGrPpgTTBrcgtUWAeUxs7DwARVZ3415xy36Mus81v+U47oP4ktlkiLulEw2tjZrb+WclxG+gpu
YZpb50CPYDVKqJkwsM8a1ZpdxTwqF1wOcpFNGw+zYoE8lHouLuhspIC44lif11rs4F8KTOMDiKXE
odZD4N9V6kwxLXhgYiwGSOBMREcQGoX5C4f846epVFyVQsNoI61DMH+yvqYimPUK32M+Q4SfP6E3
m433KBlCpLhKYlE/i1eZ1hqeebgZMKN68WuvOsbZFUoLoxZrCVegDwffP4S8r/R/g7ul+/mNXNxn
CqDUEs0pTlcJEqjT6GTpkq3Z3AVi2rvLMMDg1hRqICm6khtzP6+6V+4LriHEX/9m2qNNp4N0g7np
YMao4rq7Gs58y+BLR8fRdhIgDZGfRSH70wvGfyq67MF5lapNOqRCWe1HQ2dQ3eFGjrNJC3zN9YVo
zojx1TwS5uFyaA//TXAoxUwCJYXS12I6rYsDnA0WicOsxwa7rypaKGg/78m4v8BqNOdXSh4XWagQ
c6nkh8NIBPl0Bbt5i3yqCKgKuggyMgotDtkNKA/kApfHj/T9f6x9Bunp5YUMl3OPPDRpb4htuIqF
z3Z86jlUkAs+Z+bcx5dyPljiYXHp+F3Q5HCVSzn6yAO2es0iJmijqp/+jy7SwLERC/X9RZFX2pZt
CYx22PPDwAEnb0hpHbhZi4E1UH+EyFlTG7lbcvV3IeQ9LoRoKzvWYD0Pa8f67uzxirQ4oAAEwwNT
Cz0APUAZLFCuzpPUgazrAY3qQ2/T6q/Hb7XZIJ9Dsk23ZeqiXq6rlkCtAisEhfFXzPYNaWfh98SN
P6h08sUTkiPF7zW9mKZAwIrPDGlCqGKtaI/zCF58jgDHPLnCIuh11SDdexjnhMFbN6U+R8XEub3B
wVqbbZ7agOYEAhwz+NhR5PUldQ2CH9JSOSpI8cnOA36myR5IlRAGNnN3sBf2Nd1qvWQ2wnc6+E41
2GNDqxiK+K+5JzZ8l5ELjKTHRrrPW1isaW+NOmfwiLaRE6N8L+s3625fMoi4c8thP1TUmHdnW1R2
R7D4N1cbfGpmGfMrtAXj5Lhbm7JRdqzSR6KR5jsVvwhF5F8jgsb/Hhk244sbzGExUE9q+XSmnELr
FD/y5jIW0d489AbkT/V6o19N66fvseOyJvbxLWv9JU8gXeCjjyviB5xXjOqwzIEgRFZBtN3npaZK
6SN1FVDXlr+Lw2O8ERCJ+NNjJojVVoYVY5EgbPadcQ2J1vKMDXFiqz3L7yj9cTaWrJ5JJLYFi8tH
xRZ5pBtDPzNbTRNQoNDvGnz8im0Kmg8OnLy6l0HT+0B7jm8oE1CsSOYGP9WW/5hHZdx8gew75Vv2
z8Mztrv7dZIagbWlld6p6/GKc1aTDCyDkI4oDsKmVhxICMgQQKdnK9i/7uTVAlewmnPWTLcAjnDu
deXmWOJtdPBe0rYYrE5cv8nd9RqPLdaOvYA4D1zAiWTVmwlW8J7oYQB0zbRfqwbgWPAAr5pIb3aj
xq3rS1UiyZg9d++s2CcBYEf/qaNgo0sAZzpWSQWeHjbjeaG/0mPggElOpjmD8uYqhI02WTDuaxDu
xv80e2RZooD5rLoZ4m5JtH0Vy0PtUACps/n5sDjlCq/0ODXVAdScjHbJIFfCK8qtR89+J76nhPgQ
qJF/mgFh5mKTvai6+WSDJ1gU7Z+RQnLEpR0vuebq//Jf1qTEQ51J0poq+ckKBgfRYgECcXZ+4zYs
y/vYzshj3+6Ez9Ss7cF1+UHpr9aBH4peKW5W0lS5hkQR9Xrl58sQ2QPdL96dHrPPeItukcRD94t8
HPzjpFOkML9XjOSy+wKZNda8vuwmm7PJAgd/ndbwq5Hi1mMzp0o8pdCjbIZ6GVsmxO2w+0Lq8BNX
5Qh8gs/40k2bsf6/Ruq6ocrZJqKPxn5w3MdLyB7jtKYP/Jh4F4EHfE8JlHyCDnW4ioJf+SkGKO88
10/7JFRaMBRCiEqMuUep1iSE+7KbVIUJ1WiXPFLGuKuCG3QgOAkZJGyah8j5NKza1LbgwcsX06Pm
weOERUsYSkLmZPQ9BUoT/pqOWd2izErkompHKomPWYvf4Cpu8m1ZfPxr059vnHBVcKuwrJzOiShY
+M2U2NcQPVXMZIQeDtQaIl5vkg+2+IHBJlLDGoqxP16Z4B4M2GegtI1oA7pBTFMb/16zW7ML67En
ODRD/NN5uzgf5Uk93qSe1N/9WOVWT6Z75lIytIlxXNB/WwTHySKm9K9lBVS/D1ROQbzSbkNTeMrX
RbATQzVMCIPEqRARRc4bfHVTagn87gYzWTrU5Fozs5Yg8BkZGgNFiZCL6qceXaPNvfU3ydvFziTb
wIitb+JSvnxoHkC8GjC6GJ1Z2QsqAKnGc5yCrPhuOONtGc/kG5ShF0lsLzO4EX2+MN6DPGbuu3Aw
e8b09GGEhFfuub5Sy+SOvjiVxRJWVA3VY0sYSTj0ilOPYGr6DwseKfIOnYre3M7d2vnCuvjFt8JP
/QDC4vUL5TJLyKDdfZflZCyWXFqFQKplrJRU8K2/aDiQlw2KW9Kzs+EGf0DjWQ/UPRASu7kCVpvd
LG2ipJ5mg9tbolIRX929HKwmt5UlvliaSATBfJ5kHGs042oJiFvgdLuL6zX0PskeQNMg8fobniKg
SpQFgb8vIoFmfv83RLs2kXmaEJ6qYGgoQrJui7Q0jB3gIKJBKnCushnbYP56oQazODKO/N2tTILD
dvA+/xISUIfynpf0wOSm5F6K1je6osZynKMKMDBcRwv9WilCQxllgN9f5PM3kGDcdbO8fmPvPELU
6WalSmuuTkwbksRt6OwoA4AYptNVsacVcA1WLq0wopGH/mBfUlrWrNrdeH+7OFcN83glrDdIpd1Z
ryeeIQ0TC4KKBj07E7T30X+JGLSx2gL/SwGGNxayoPtKN1CMhzY55qAkkZB3QjeQrAIc12U+pg5M
bJDeq5mDmyJEoq+IJTb4cdWHAsIyttUeVM1ESGDdAxjd2vbyjGDhDpGeLPE0RiL3k6BmXxvIzYTu
x95y6WspFbf6/72gYn2lKfGi0q8Ar7LFE5BSsb5r/9B8Cx5UXctJ/v12pdAS1B5CiCRHquAqDIUL
wNhVLR+ipHLlQs+A2Ne1e/lCESprTwLW5wk02PFybCxRVRFP9ohjjRlIJintvROZWNblGDmrNIhz
TqwV7uW6zMQ5yl6trbemB/5dYsyFMa0CUQHan2zY528lxcUZq4M8JTzyWSQ1iW91Gz6stjhpwtuS
VvwZ3+LGcj2RfJe4l1qulY3dHyIFdG+palNeP2e3/iTMvQT4EFOpdbUqDaI+rbEaVM8i7fFPmfBa
UbqrQFbAHyIjg7poFaoMyvttcwJinnrMTPDMO8ZEjQkk7rfIQw5jaWiEZeSxMpQu7F9YJKedkJP1
G6E4WEH5q0DETjWlobGFOMo5ciL9EUr/WoqAaqtoKM5CsK3qZXMxq8hlWT3EyLJjgU0P//dhFawU
kOWsLOavtRLEV4MkEuW5gH4Y5FeaIYfaqUHB64EtPJb3iaPvqzsFAkLFmZR2MdiN0FOgdaZ3CBAO
7OoS6aiPD0eLOJn6rE8BiWulb+xo4nxSu+4b7uuMfsLLLAwho2yABLoh/FtvBi0Ua65g7tS/X4CP
8Ylj6agIqT5Vvnk77FHeliz56atSQ6LDM/EhPzNN64IhOmVQednROpnrvStZvKlu083jFhxsS66X
AeY9XgjdFZnJaWXq/rJW4MfgKHekHdQxFeDdyEd6dgrC4xzPvxQJzbt7Ls31RI1rlVk8kLttwnDU
PWTmwlZho+1uZopoPjC+jmxzYFXH3Ffiy4RFAbX5heFxVIH5xhhjsxXaMKDYslv8kkR0sb0se4V2
xb3xNWdbNlMBPAk9C0AXbbTT/Zyw2uttHIFd7KQGN1ansHBBDnYdhWihPGmRWtSB/H8WJU8nTHJv
2KhN9hZ9yumhS9r2JFNLsdgv3o3EdgqkrlZ36jPLoXbfQSPxtjMLtKDZ0LCd3emLLlPcLcpuWD93
2ZGIg/0xfCkkx3Gjq1TF4FJROAOj2hSU2R6vLIUTx2OHlYYI1kaxZRoLPez1tiooxG6fc+aiBDQ1
RMZ0zm0iHpWcpRSBfNZyB5PZMN4SjDnnRd0ShK/lUahmmEOjvIL34D1Wj9utV+mJvENG3CK2nBpp
Lx69RVtGjIR8L3vC/El+iAJJzVfp6OceFV/pxZAFUNm7e5vlU8oSXpi2u/dsh/+VvDD4f5gX1CbL
GDypuFhpbc9VIh+6n8BTksXNdLnfV+p9Sx54RLdt8XQ6yzqex2241uJ9OhW7IT5j0r/meMeIW/6P
pbLXQZQIlJtkgEq3+LAoCetuGKmJ/7EEQOtye2A41chpzYH99SapGrNRAkf/vbKPX6lnBimIhoZt
nvJ9af3cGyq0nlb90PvsQqidytk92RrSM5YhKkRzmvfL9ns3n+GcfguLuuVK4gwtXFGduj5QmAQE
JG+VV9ADs9HE+k+hgOn5QYEFI1Tskeo0kPpcmkeZEVJX0TrTqdXrSNRArjG4sqBObHoX0vXARFrT
GaTm6MOBj9Om7Q433dghyOLM3uwoM3ZXqECG11G65CsB0Rdiszn2vWAhvqVbKJHS8lKKDPrSCBT+
f481CDh/QtvCyJu//AOv/PbCuBfnhEAe55J8NQea7+aYIaPO0TG9xZ7Cua8yU6MDGq3yi2gEmuB0
CyES8srpHmwiK3eN8XZk1wmNfoPphURg7MDN2FnPqCY+BOb9K9kyz3+6L9fHTMjGKSQKTNOhE+/k
B7rcoLaMvpkj9QcGTbXKvB25Qbg41wg4yi0TwixSU7mJGYm/6CdYOxVdnhpiiQ1JZxic6TesBal3
wLMMxOKubpQC7DN6qm5U3VyLcNvm0wmie4rsP31rvSVpEbhsJ1UXfn7GQx56i/IyqVVzfS/FTgfo
H6l1DHQZLhCBASHX54OtzY+lGaEo4BHQbIxFSZrHZCIEDgfb7DOElWBSzGeaaF8jaAOn94yIoOJS
fApOwGvDPh1vNKw5Sb1F4qE8smkuyuenMrDxM+tEnfZhBmoQROIJwolDq2FrJvvZFUJWuUIkmm7c
7XYFskE9O8E32JG2KhqAaXpCk9scdR4Uq80JPuPrsZ4J4XI9Q9wdRfa7Ft//BhZoiZScYodpOJHz
wLjWqeT++hMxMtB4jzopFaXtM3hIMGtvn02qdd8elOo59MQTlNDIqPOWuprcN6uvegV3FAnAWDRA
IowkqpUSEsy5g/jbRIa6tJtDpoy2GVP6bgn75dT/hMiynX9SJDGkTKdonzzcrmtFBIQjsRVap81I
ZMtZ9Anv358CEdlxt19v/u9QqY6w6rp8y36uHTLp2U3RYzywJZ0JepWTMv03KQsCupZ6NJTOR++I
5MRW/ur5vkWKBRCUojVTI12KsGcyACnNZs6DCv1BVgzmb2iPy6qdYhgoqIBbRmPbXLUnKRRIT5sU
fTYwOvlA/6L16ROL94GpGxWBLQqV5mC/kgamWJxvb2VR+1UckHfn340JXL5Fi2sxwAG2poN43S1I
5fONGD6b6gmwHsguIovQ7yY/kDF5kfwIdfwrcIjVuOWZsaDqUy8tB8HyIv5ol1Rhc0uHdMAS+mDU
1rlvqoDxnZw3lSVTEuWsGAIh4ouKCZBDk7SEEUvk0C1nXfWXSH5DlTAkwXK02Ckz6za74mcC0scC
KzXjef7+62Mm9voeq1tuKflyc0j41Y36+4ralOPXoRNcW5agKkSA7NtGy5Xr/yAJTmHDzLv1S2v3
JxS/d7Pt6KLYvR3BA8+kRWOcnyfxvmSSdZUEzQbDzW3LG24K6ZTI+AUY7rH5xXti9up3+ebPAssY
Uhw6pV+tPDCzbLJ81p7Sov8E0SN7UnXKpNW9uWx0O8o7VpG2LyaVdDBIpyp9puhfKX7WzlDoGst1
sCLBEqitQ0rCiMi7qlt05e89PnkXXlxIEGUamaE8L3w2JMKZ62qpWB9NjsnVAJIgAMZ/XSNNQeud
PJWWmaYl6qh4L0zx8rkkqoKk9Pnng+EmUI+92i0N9ttUehtlbWpRs3m8sW8Xu8xNXDcgBfmyQq0H
Ghv9CyaEoAvHxCPeWR+MsuH1LnM9MeDHjDJX9lswnfWcbVZJc5tWZxFdSlf7fWKonfOQTkWraLwu
Xi3wVXvA/YxM5KP3NNub0NHSFvEVE9ePdG/R2IuP77Bv4lkDf/NjKq1XuUdZkTdFJ8kSBQwdYrft
6x6QRVSdXnZbcKOwv+ck+qJmhQUPawIln68ePgadFNJ9iDPzxDmghMohS8BoBek5OawH4f393GSY
Oi0TEqoLzYSldmTaMCFFzlqEO7ApuumaK8VrFPnt1kHJh60XsjlVBe18WCF8iHcgNd3tohXGAdRf
qr+6PcHok/0DtLzCtiTdj8CHfqoNp/AsPiaPFzyw5AN9yzoR1z6rDTaT7mq3cHqeNG8BFh5EJExB
k96gTqssVIFJiSY8C/tWz2+L/YuNNIuXHqZWeZloF6BSkCs0nzDkha/IAn4oUB334vJCJxfJSXWm
+Ff3MVaAIw2zqIqfJiVZqq/2CmKjAVh+TO+nbltitLO/d64QNzIQ/zDsbbw7GHw2OnBjdp5uKgF/
KqyEkIIvNRdva5skbv1VPTUrYvCpWkpvZVwNUO7LfaffAaQBsktneiWBO0NuveKfOGbkNxlPdnvD
J4/pIW+WA+mf2fZTDQs6djELlFLGQk71JCG+Fout8kgBo1X3zbFpvmyvvuQoGNRbLo7czKfIV89o
CIpVgnDpHm6SIOFdAjlbXmu+DWjBIBpd9bgkSgYX2fPoZr4ZAZjHwlUuhKtdlbfe7HFhCy2lrZCk
xH6u3vpxfC0Rfv1k6QyZ9KoIggDb+6pvbpULxM+Qgi7OMV+tLtjBvhD/mK7z4U1qWREGV72ke89Z
U9fEzUyNHo2qjT8blirv+uTQ7k1Gv9RG3P+yeEMnYKq4RDK2OgT+83zHmHJ3uW7liJq3rEKfKYmC
Vzbk2LMwjXY0JQb+02+eYnl0Ga+IztQHjDrzJCfVNZt+Rutq7/Zq12tmtoupigLtDWiHaZ2Mg+bu
vZfALcvtFulw8CjzLyuMqqRMMcR3ro8wFi6SBfwJ7iW7VhYtx3Pw4i/ZtR33epwDOZsV6tXfWzoV
Ao9WYda1hQr7xgSIkqSBFHmI5oANXzbYxNT66FCzc6O/Y4nIOqIeCkW/GnsJoLEIirXXQRvAoN39
D80SXzgeTCJo3NhDE3fIJbJKmxPRHKB/uapgIbrRJcpJOx5CnNWEf3I67cA10zNk9/PVX3jS0t9+
cNBCNYVCZQ5sNTczib4izg+Ct17QUzX8C6beVkV34Av3J41usOLoFbBoVk8J6/Uj5HBG9hoIbL8Q
qOzUTbOkoSCbEsuoOeQX6qNDMMRIEe6JTORuo5j/gqLiunyOcMH1Xe0voaizozQIcmKZP5ztfoGu
qNhzIb2YO+PjNDGZ3x7Z/E81wyn3im9CZ3Py99+dV9E3sHG4QmeViErLr7qXq2608bK7oPpIgXXB
zjo2LRqW+livQn3TMI++9ms2dd0pgpUnioZDTNV9VNs36aSD42GQyP61SaKTfqzFXUJglMY6I2kK
oSDkcEChva1EU2CbeN/G8+8kFSXe3Tf8oBfCgBOneSdQRJL1WmOlq/Cyg2qpWxiWfRNQVWNafD6r
zdQZdn6p6yH5Gp+E89//kNodsmHdePre2L6tYP9UFEE1wP2ByYBer6VtvJARLYi8BrQ9XvTPmIye
C2j+npcGiyVGUNS3VmbpNPP3hnHqTG4loB7xH6MllVqOFgfn0pNUFjUsTnpH8esndv7jYeE7WL6X
EkIZupB+LzSiActdr4v+PWNrd6py5hed/IbRVU1M4HhE+fYX+VKMusLpMJRarEnkTLUvIIFnkHAD
aiHr74e2oGGPtrrw1/FcCkx83FEgzDN5Vonvp08BezATGkY6BQ0YGJnY/QkvGIbLqowgv7jWPS2i
vDLFgoB+SBVzDLc5//IZ4ZljSfvE80SyQtQfOUiKQci53N2un5JfBubGG1fRU6ElFGoXPM5p8I+I
N3otaOCvIj+a5wuJrJsdTfehD/6qxxF+ozWwhB4bPxE10lUD8MnQHuzNGe87vRkzrlGcvCthW/D2
L4O9RfnHgE0aeFiONDM/XNibBs5qIFGWlBQD4m0KMWR1iBPxR+mfbkkbUqSfLcZT/Ni/L8fb6a3U
amq+a3z6Hx7Qg+o4Q7GoFIuJUxMb7D3+3gmxCMu5nnGz5oxQkTJKI6e0Mp4sqfBBKBgV6IaKB+Ii
ir10qdaRQ/noYfvdTuA/g+TtWE/G4Qj8a8yuxplYPsnHc495eglK7VvoMayJjs6ytrjRFowfiJvR
EEhbVCRz5MEKzV10puSeOvvi7KJI9WEz+8UBS/BtxmWJg+fDiY8EragFFMzb0meYrqJ6rVVhyn5d
e7jAPBTeTMpP9q9WMQw6TEp3GIOo0UkVyHYMWYE0rbfIei+2QLnxTtAP/hmHwd5t/Xo/zt8Lo7Bk
0zY8dSdsC8SYYbLMjtzTxYHq/tmZjm9j44F8XRIiPhByiwjhTUv5f0EZa4Q93RJ0PKnQxBMgMvdM
dk1stGOuGarh9VLtCxSdnnUSouoHFVYZbpQZ0gSCUE1AtnfccXXH+2ybGJmkBoYnHKZQQkp9E4SV
MWJVVY985UG6ICqEqNAexNaakClprf9IUjKa8PEqr9BgxMVQKhSyPluK7FlqJSQa1ALN5gEZAkW2
Liiw3fxv8AqqDbM4MlJJ733+KaBCCJSjeJAPQrckvmCjnrya4mZIVmOfsCJ+Ia1yEffdinnFhU6D
xLeRcoG1kKh7L/pItuUEg2wNpbBqRy5tvfpE0DNK4pyR5XCkJ8muJAQ+QUhWPPz4zIIbIC8p7nTe
AKvJ9l5BXafM6A41kezN9JEvNN4o1GuFZF0Lc5dtvdt1gFeEcjWagtYbCQEH8xg1fik6LVOUWNoq
wnLoCyUs44PsrjThwYd8P8vuNN+jTBrVWk26nvbKtJSRDw5PmTSFEDh5pvpsE8gQuYpDJr5JVG8q
P5cOdozjqsCg1tlCT1YLUKJSwiWl/1esOwlQo5pz1O2TGtA1GpqszjLAkXwT5XxVuoxfNAZ+4FCc
M2vrNTFZz1Vc5Nj+8haw0OqDrIMn1RqL//UTfR2Jp44LVvtu6/aE41UPreDohZWIebA2syA6deB0
cQN5KC6V3rApgi5COoAP7N4RPgSxHIysx9FVfYdMde3uRBMf8Pr/w61GBCU9rq/TazwyU/BBpjxv
mw8jXXxOtRxk3H7XR3AIn0/LAWFXJyUUWX5mNMZ1JuEl6KyrH1Z5xW5yqY2sS16HdXZxswq1qQZy
JdFajLm/527MDySqDBymTuPINtF2tbaKZXh9dvvpP4uNh7uSyIxfWNgI1fxmNziYsC6WFBihHH+O
1g+vH+HjMrEqyx9nvHzG6RQW84CvWcQV+Ou54tBlZBUFP/F03yGre7vWsu3sp4T3ZdNZXK9QLsHY
F1MdOBxt0N47QJFZ22NECtRyhRo+waOSn7jDPPsbAphsHWGCpq8RXQNWMPNSAEQJuqHmQBn1VO+P
Arj+tgDL//RaO76XPXYcuR2o6QFF1K55FyW2vazX6J7TveaByNxWvU988fYdsHKsqUzWAxsnklmg
/ZSRwSpjqeR64UZ+xotKC4K9XkK9WYz0ba7gvnoRZssMc/Yl3vS7cw6YoLrLLzLR3z065Kyoa1f0
uhOa0rgqGGUSezwjYbmf4cJLWJdhBnLykeiCYoa4FR4hiAK+UaJbLyzLmq0X3yXAepTmaBhJogHd
8xLn+GOCbdqAksfYvSjj0ztKsml1o5vSRg5pF5Q9p4sLFye7QWeez+KEK9tYjr8fzZayh+ewmXK9
9KqNhnAxwtXwNQKpVyVSd0qWL1dHz7/Z4cCLIX91vc97bYLKcX3VPz2CJTpl4IhsCfh0JoJS6obX
xfoWHXkmWhXbQ52Vojs9Kn4rs3ICD5FCmIS6TcDwOfCcwGsuvRyA11LveYk99hzv/feRSnEWiKV4
htMaM4CU6xsvsBHPoj9sGKfSTI+9yC3aURRmypWChg8D056BAIYyu9ZoHwcLdgXOMZYJ7VIcNiIP
jq0h9J3oN8gUNdcnX9HzP1FeQIu/0evgEW49MSOdJ4be6cnmJpxFC93Vi1oKfHFBTWd1fEG29Kv6
fqMtOlnfOmrL+N5eu1Z0N0huBOIl99TG8wc+QRygLnwEgfJ75HX7G5p4GGB9DltS8FK6EGyUWgCS
FcPWZ1RxXB6A1BEOSxfa1x+mLYnEOu+u18jAQDXdqmlhyw4Wcvx1RWYUmcqvWA7JhLBWwlVI3OYU
MRwUGoH55UxGiqLLo9qX1Z7Q8fRBX8s8xRyYtuRYY/R2CjsxVyOO18WwP9JJ9U+YlsJX/h3akzG7
wWiEUiW/tgktwO39fcRXWkPhfZ2Ndls1LubC8kzkJshRa9Ae9ONRwfTZxmYdw8K1FpadFxUn/3Fr
6E5MKnORrxqZpjQvejN4BIwD8hA4YNZGMLLUItExEbaeJAyqEBSkdq5BqkJIcdCNjbOx4TdtloGv
2D5EIG1Oh5REenBp/nmxachaIklzOLsgTY62mMwkDpPp288F51M7+POm//F94mV4O04E0b0Sdz8d
kenXfFw+X1NQwJyvKTqY910I7HGyn7gXYZpPuWVTD04CM9oD8p3kd1IYKaRpdrcBN+xoPA2BmpDc
ni2S6YPk5zLrnxd/wbhKToh4obmbm+NBOiGsAaQBGgWKT2J/1eqCWt8Lh86E4q2EPe+aXOkZsCbt
zVVkQes0fJN2N6kL1vdcJlLmNjpHGyud5qUAuEgndz2kx7ItY0oNWlda55u4hr1eW1aKBOld+Hrd
fi3EAFj1tIq9z5LVDhb2UwKltPIEOg89/aFXqf4meS/Ent7AtjD7cCYzianj8Jq/VmE92Q+bsHD5
7EtzOACWVMegG693rx9ZJL2LsEUZ1oi2lzvrP6jRFKYveYxfnRfO9f94ahkVOVccD52FDIo6OhaE
wAcDGePJFwbm1XcN76veU0ecvBsqOt+N3L83ze/YU1IsfKnOm1aUjUs6cShDEdOUqQaGNsHTZd1C
QKSYcK3s7dKq4N2UpTExvyaxLtYXiew2ZAJPZkVQZ7DPNzTbJaWeLk1W1yAj0K4SZGAllkCv2Nqf
3HZrU3XB5htjpMKoIj9TgKMI0c/ipVJ7aBccsY3UXe7Rxpe0KGFQfTNMku2fDW1GVBW2Z++70OUe
33lQ1dSI3JtoUmKChUeK6u5t80FISw4YLDr0hVZnuFmyDj3hbM/CXdF5vfy+j3PuLaS8VIs5x+VD
v15K4Q/Aoc/OB1o8uWpH7gZLCKlzhmp+bMFBsBsUyJfM7i/WP39GYji5GJjXU3DcS5yF4HH3ecFv
3UyP8ZUBO6nokRTt93mXlAKa+vuwTw48yBU91t4fAuPsCuDzvcwJQviPMYJvln4vRN4jAIYOzEpI
QQAcFtOBMNfTi3Tm9KHZkVFDO92u3FpVrBBucfmPasODW1xWYd1YwD5AmXeChqZGkgLDLFhtVwp2
WYWKVg1u6aUVAdj/aNsmjxq7nUsGgj9yCNK7WpF9sn6xdcfFeSBZSEnJb+dlc7t5Qnn+2zLSMDl9
cQVOPZG3jcLZYKDYJAb6NVDJZigjTasGFjZZwmDYUl4M3kEO5Czdo4EqFnqZd/VH4sH4g6YlkoEw
jsWNUteujDlvdCAiYlC0RJLOAKsiDfXdW+3r82RE/vr2VX4tvXOsV16rAQB9XE+O/FGIa3UIwqmt
AMY2hb1OxHbQCT8B63GlCW9IRzhem199lXytaPdPCqhY5ygJdXtOlORILwXB8TMX+hVIjFFEhjfG
PzpzweMtYng+zpaCiiix+TdvCwro3npidJPalgTmH4GxUbd6WpEQh6GBSKmAhgpvWfC9nAaFnoLq
w6mtdJDFj8ZRiVvpSh9QppSYUW+ja7PwnEaapXaHjS4jDOvpoQ/LXrMPeTP51TUX4cN5259wJ91x
uunKP6M5jK/ULV8Re7MsADB4jKdhoV4hCZQ76wh2yfPCOXu+8OLwxm+Ro3yu+zd8OpQrAgHPVLK7
2Mytt6R55WMGJSWoP5ScGxPs9eT5JSqN4WRla5eMjo8GbZ2UkFsDagRweIGYNCKMaZK/mYL1m8K+
0aCHkgQcjYlcQXgOZJW2gzlEhkt0RcDE4X6VLi2vor7SR8h3VdDfAmLJp8ZTSrvxkoefgF6aJSc4
cBlrlpq1JZ3MgRRzpTTwUsjC6gpcZYJu8/ZN81IK1uH/ep2PumFl6TQCBDObwHkv1At15Po2VonW
PoVe+r+sVmLNvFxJ/b9sZZZXJ6CKz84C/ExXVY6r2v/AkaoRwE+VHGRQ8XXLQyOGcyJJANA9JLKJ
AJkMfUlA0stcPAFGccButQjz1K/21vOuGibtXnejrnOfjjzt+DV62bG2JmB1L5R5oPmiLYqbgCDt
cHd8Q0VDdHxqc7/Rr/MIuCRDB31sRShDfSe87qi0sJXWZZ3qTfiFGkAz6pBrP3n4xzGgs+Aaq5mD
TqFe7WMoRFcYWuok78DPTY4YIxv9vPPLrtL4cp+oYiliDkJ3hU72cmKSqjpnRek6SVg7X4asauSk
+PzJUrkZWth49xyIj5JksqdXlHaTLsLLnr+4o85eKunNGmnmPnCEG7PvlQLbq9/u7JGu6U2xmrpX
2Yc9sbQkwglGYX8WJmDVbyh0OqQK8amIhI5s7UoGSyQBVQ8FHRXYOOTBsE4VYloLXJ/ZZs6qQScf
MwJuFj7nyZh5NhjgU6HrUwxvt7aiNyLkOQV7CWCGnI/wKWW5gImTU+ipXTJe6jyCi7cWXscbEMXj
IiF8I/6T/nQKNECf3Vj8xZwUPyeTD3GI7fRrAYZ6kOK3U+28vSmuly2oHEqj6oTa/WvJtviYwv9B
wTPOBBSujrPTN2GZpvEXkNVMAgvjcx285TpINaBP+eY/T0CNBQkOU3qt3oHtrcbsO9uUEheeI9Jd
3A3oDVlnHmReIiZ6HoaYbTgSo5TKt1TgIxt0gymdyFD86GITYUPurklozwHtLRh74Hu252TfTPha
JM+B52ntDB9Bd9lDaLfeej4L/7Yyr43A3fu43wa4bOQzAY7DEZQIoN8rDGOh3Ko2hGln7XqGAg44
xjNbx4DJ46LIru3KOTxmSjTxCXnMDBd81FqA705DHOIlTW7xshjb2pqCrw5cuFtzeFrXdynAsYPY
Z76/L+mg2rA61UnmUWSqSKuWgaHunnN/lKzBC9k84IwDQ8k6ci/jSILS+sQBp1D+sRTnYv1abKYi
Qa50wo3esUIKErrTDSy7Mc6HuFFnkxRg6Z0kdV+PmB2CQ0H+G5CbGSKZb7ygc5AMBFmkvu/X1xw7
I8yU57s6+NlFwCr0Q/HVjHrt6Rgs5Hd2R4T1sG4LTXzKXJ70GJ/MKLVSLkNKO+KQPCklkZr87OBN
KTglImvO2WUMiieoeJgj0mMG6BOisyQ26IYqlBauwK/f1VSTej0onPxOybljJzE1eBDINntOC6MI
mg+UQPrFJhXeyAee9y/bSVL5QMsgYE30e615Nxxc+fj2eAAg9M4+T7z14IgA5lV6EB3SlEuvrFt9
aYtAYga2zU//nCDNDOP4BB4mT/lIBZ+0+raYaH+YXi8kFk232XTz7OzWUvD7Z0XwQW8faZ0Pdc3e
VlMivwcJQ/WVb4XoIBzttUoiAns6gwB9RvOypyQEU+m+6MDh3eYf3uxVSzSE9fmCKdy3Q6GGRINa
raK5yMWsUWR3NS2TuexMqPE4wX+kJlXFnl28HeLlY8/UOdFDyvMzo5xCBZ+B3zh3HNWO/WpdGs8k
3vNqz/OrPgATNx1Ewo+V/IdiIaOCCIhO7ppFVMGdM8d28FNqkha8Ojop4DzF8DdcE2mZE5N7ljkB
exwZxDZjpwTeoCT9CmrrXH1Acu4avjBCTfQmVNAR+oLT6l0UIxLqF09IeXmsDh51KdxCEopFc33n
GkeJdKxScGmlnnpaRQJUWBBsy8y/73mVfy1X/NxSc99j8wdu9O+Gq0Pw2nd4+1+ejuVTddFi917E
YqXSlzi0h1KSFiqSTdaoi7/jedeMOhpvwhljxgLXulURfZI8JJmoom0feqDUtn00HeA/LVyQ8cFe
kTv2xu3WNnv+2UYVfaEHkW2WKmE86BMdjwzgppiyw5nk1npRKuDad8kmAUQxKZd1iX7NZaKZygup
17vPefeXsY4xD6SKhipZZFzztvTPl4E0ZT7k2Wn1d1qvODUZaedUrZLFtIHIl2hYFyK47J5TqK2r
bQdmVZh4KxHB9dtJGZsvq7ZaRsARQwaz8wreUc5I4zJdza9wJlxXNOgDCgm82IqPGUEqwoya+OnS
3KP5SCHzx6hy0Vp4ijJRa7vh4Sm0GwiW3Ut6L55KiD3he7o/J3tkNcTe0rJhxC1e+RqS6dIYx2GT
RM6Lqg0tNAl1jqmh56xmgiUXkL6Hh/C+pwRPWlQ8Le6yirFJMu0rvG4GvMaar9x04ZaNdlIyRPWC
RSOna78xcU27nZrk/hivs/MezNAq3It1xElPUsvyaXzEmIt5Q9wDwnns3ngewKLHKzktXjz+ghV4
dL4PKW+vAHUYdHzcLZ1HJulsiEbg8GYuVELkzFwCKv8pdbCXcWIlOCvb/5OKDIZx8QOx7A3KFyXj
lLHw+jz/bHrProTIYh8NtAfBuIPDlP9aWX7gi9mjGBWfU5IK2KXBwvP7RPeIhIj60NjE1uEJ6Ct4
jjp/8b0y9JOb6u54j4TlHhu7N8iiU26uQ4kFuGgHqO24R0/vHNGcYXPEG9qUMg7cS4KyJ3SyGho2
fCVejZQ6wHJNfIamDjCwOzagVoCDVQkFtN7fZSNVHjAKebynGpPzRvCyOA2jnJKHQV5uc0pHuigt
S8taMg5gWcAa/7XLWJdZ7HeRJQOGc13rmpjdWB+iPCoDCzFFpd82PJqnJvk7FcR5D2oB+6+6CJ2w
ft9galYl0Qy8TpDPDXMjOS4WxZAd8mYZu6jO3WXwmIEMQ2Z+C8jiLgC7yGdYW4GJcQvp9E/e3AN6
EhvX2TqNlbY2YoUm27eWkzf9fOdFZamwrSQkrov1QB7DHKgoZpzPjlmPOSKCKabxUXO2WkHkGuYM
7To90EicORxSwwMACg5p1m+xHDOkRD5TZgeMvEE9P4oJ/3TRPSEGDF8692jPQC7DML8i6cf2D0Ar
2iVc1Ni9Gg3sFL+owOt4WTaJywzLjqNZzOSg3NhMFIcCZsdKG9h2SbTJnkmadUIwTULx2IIbgCUC
a381qF/ESUNc2y/tCkHOeN95/Ddq/tHWMPojYS8+6rPQnHZi7XpM9NDKvlC9nUIVKhltAGhomvS5
w0oisS5zTA3OX1qP1amfNtHDYl3Ettc6Zv7o29+YOfgEZfrgD0gk5LNNKN1X8YteufI6fmw+pfBg
kxjj7NwLMNamqh+WIqV0khJJTMHiZzXxtvyFJOiUF2Y4zRzTIpHBqHSF6WJPLqqYAqbFyGoMtKhK
LiCUXfnIbqR2Nk7CV2kBfbo7FreiihQHbhwYC5YOzNXoouIOtOz8ORPazMX6g7Jd5pFIiZtb1oof
G0JfHr72rX0iMT+Es5yTfp/JSYq2L1fFQpRhv7s3lry18eKd6KADYVuVSehWEdng1SPfvO3R9Ia3
ZXGZKmsFFgIAi8nTjdRq7kwNco2euOgOVUkmlRTbbhlsc9c27wFYTlAgGJuhyPxb9aNBtNpM5k1E
zb0zlUHDN+dhCbJ9WvFqvGvaVkBLJRTjeCR2+sC50gRI+THoI+G9Ovrcox47CTjHkBKjlJW+Logl
yXmYbMZ+8H+Scn3Nl5r+NkCkPr5sJcyKcKsIlNQ+4bdM5S1dwf3rZjWJ/9PkQPeL5sGdd5YrUldn
Uf14f+4L6Lqi7qExZbhkHZR9N0StwnODmaUtgJ80oj6irf/u6kFXjeUpoSlNrzV1gCXJqRP93MDF
AMvWhn+5axoGckbpEBf5J537eMoXzTGJ5qMbowABoD2aFO0920aJNkutiiynOo3OaLpZmeNhMboF
RY1rKxhOQ3iKX2B3l5IjNYgBV5GaPHxM3cWfUlujH0T8tyhOg+EVrtgfHujk9lz2sdzB4uyxJHkX
70nqsWUzMx7jFSznCZdmjUNJVziiG+ent5/sMmOdYDRyDT+AbjxfiANN6b1ndCivxUBukihxBfJt
NeBolpwOkT8Bn7D0ExuwRdQs/4sQk5PFSrkKQKUb1ArQuqqbm/Kao3OjVPJqxxpUdvY6lGiB22Bp
hQdi90jPACapr04Vg0oSxpDcr5Llpz6FZxgDV3YhRgdRs6dyeqXByKW1CZvzuAaHRY5JuMyWI1Hq
MkBBBkjpiAWGE/gk4JbxTDl2cWXRoRCn0GUtG5Ik9H7FbEtNcmMd9lZieqLMe4t4EzkYcJY4lhq7
6yoQpIBdaPCqJ2OXKf+UUKlc4XTGQ9MYD/b5Wx9xNJJ+n9NslDGeobfDk65Onumn3of9BTDpgpfK
U2hTawfp4g5syfrptkGFrY+c0Lx8lbut4jKzeqQtNbMCspNYAzKZJjMorPgwOwTbDI9L5fnpoDg/
mCcENs43OjTxytAyJrBueQq5m9lm526gj1PUhfCgDRqC2+ULzh/G8jGuL1IXtgm2PRCRAgWzHJz0
SBu6bQCRF7zStdIO9Dl9IeCwVs2DKwt59eIvvTGX3oDQ0Yt9tmIyxOuuPd2oVZcAmdZ3V2L8knqJ
ekcBwurvG6RRkklpDoCCvfgkg7evpDABxYe27qzgRQ+Ylr0NK20Bv8v+V0kraD+Ztl97/exIDZvM
zelpdzEtXXelEU8l7YLolYD+hsGYO+TsCFAR4p9zGFgziKE64u2PXTEQUtqaUFkYAXb3qm+wc8RJ
8z6Bp5A2t1ia6szpFO4Fm/dRwpnFV5aojqiA2FQYs6s29YBsXzEfFEcBlytWFrnbVVDdto8KXoEH
kx+M+J6xYXryRIGCSn7+0eMLB3WlBnJSajBTmQw3tAg58SP/HGs9f5Jacqxz+c4hPp3UYi2KfWxa
aZMXIru1gBfYsbK1Y4t2OOSRq0bmLU7Wd35sjk15KNOwp5bWxeT9l0QzHZMkI2m8D2QgyuZUlL4g
PIGSt3zcyUL3OkgY3CJEzEUL8AtY1Ixr7xBjA4uaQxJl9AJdKWthRY+hmyaDCjrh3xxmBt443d/d
VMcWpEbGrRJ6kKYScHzVDFHCz3d1j6lkNYHm4J1bIgkOei5AmdTtUBpo+ifpwmiokwGWmIOGFmOP
Icb2SvK3lP9RJ3Q8JnpwIwCV83A/hhY8Apd7VBdNVed1gP4xYNwWerfjjAMuqoNvTeZt8KvoZ+Ng
MmOvb6dBYrVcdXOcocZw3hD55amMox0o5+qPZSMCRKVAxg9XzacIC8Ho+nHHHOw2H9faoE+RqEhM
bcEs4sW0UnEVIEnUJo+5W+8fRwVQbLXYmuMGO3tnHHFwQoQ389xfMi+21k39KO46GoUywfPrL0oO
ByCP4xxmdxj6FYe8V3qZRhTxWyGPb8d6plf4dbSZH/Zf+ezbWE1VQJDuiav8m4YSLrJ51jimLUVJ
JVNd5ggxzZHQYhKXCdFW3dyw514UyV441p5n2HHYMxQ3lnwyrpebNNA3kHnAylUikYc651VQwlNg
nxKt0eHsy4/tl0tOq1EulO9gPIyagRW6XjK2pISDvQlcOfZmZhrbhLcAhcvtMovZ6sN6w2m4Nnu+
5KFkDl1caGCbseria3GX39Eoc9sKePMcyUqY/jnwINQecQ3kSl8zgPatScDS1JB/T8SsFn3Tum2y
hV+EmTmyaeBR/gJGWy6gB54Aw0RtYWDR2EGJFib7jW6D5+eXW6z40bRlH64XyRz2/j95wTRSlYJ0
RggjL+jeN9DZ+2DJrQQNIbI/piSi9hy8DUihby+luS8VqK2NCu0qI3jgQu1Mw4CeJAvegcgPL51L
ZB/x184NXgekMpABATcVWftY8b/ogf0bcGfm6kGzhe7Qa7cTXoWYyOw//XTH2jtsd6KGsrxiDD5J
Kbi+jAJx8cOUSsbsKwhOORL6W10DucWhvSsvQPOBEdnn+ZEhks4z4bxIut7pQWdvpcK4dEjFZeB3
rV4z/Bm31TZTS5LdRDPg/7lFyObyR1H/ZRkzgzjllm6w82Gvt/qIjSQ8dmAu7dCXqaIv7GIUrXFp
qw8B+NYPE02DifeD337Bso/CAtmlLzkcW+HWtmOazUdfYKh5/XTObjm2ls9Hg08l9UOhRk/Jtwut
UN1x+WZIh2fe9G3CtNhpiyy5H1Ie2PW9T6Y6vd6nTxjZ4zoIQWuBnJDJIKzj1kzEVsz2xIEpqz6N
D8s3AlNRzvOTRW3IYjKnh5jBdAqP3/zEhNtP5Cor1RPBCy67SL1FRkcD3IVGKVQfdGuOf03BVV89
/YaB6D8jAf0ba+a9P/f51firOrSlUm59Ht0LRQrM50B+uO/+j/AAA6cBb7Chn4DToui6dHIiVs7T
g+dYzB2hKHczCq880KbFcFIT0kwAnhCe+/JdGdtODEMA70/3irgwhj87wDYB3dFmr2CySZs0Y0HL
654dCA50EYOKZlPTikqexutDtJC4oWdNLT1dS24AuOqxJM0iZWtQie66jAvduS0WLwCg6YTlN8Og
M4KJTfWGVHrzZEbv3NYEz5TB62Ovc4cj6ShEe2p3O7qiALXjhHnMiJJMxrQEQoIjSqssE1ERp1JD
rSVF4I4ZnyKDJEPlAIPrcY8HI5pvdS3YdgAbg/U3bwvmvuaG3/sVUnSTbNIINH7r9+o+n51BR4K4
j8KFVKqgcNeh+FLd7l7gVvHbKW4dDNa0/71gxnDKdcEuzgDO89Uje5VWTh6ao239uZyhxpEHhUtC
caBhiC+AYWXVHcYwklVSEeGvWDJUFYJX3Px58lbIr7rSCjF4Am+mjk00lPwkVZ1muAxGxnjhuu8q
7XiZTKyWWw1pxFJJKASFFePrfPVHxM80KoRWD7j91psyK8By/VSxZJ7fNfTKzrMtrgWnv5TSUxgc
rNG6PPcpKCjb9arghEa5IpKLd+1JIQETCmNvT9eZg+r4VtvhfuGN8TwDZ++aeox3Z02p5xvC7ANc
opAlIeV7tbohZY1I1If1rErC86+wCwx0X3rAqCWiJBiSUzrETWLPmZWowHZBYeGPMFzGaSY4gBD7
GmQNgvLSxq6K19/YEqN9dQb4fX5exD3YNnA1XGZ4OKGe50+JX5LeDwu9Smq5x9fjAD/BcwWuK2oO
TfIgLR39GjccbeYpDRk9UM7ECiBXJLeFIdePz/kdJXB39l/SqRMLM1XGen/GnmFrFAQ7JH8P1fMo
S2c7UNqpI3qEctwhxP9+IUIKpoKClB7dgvngN4AUirL9s4I6NepT4B3my98ZtLsR7w9h1+aQhBsJ
jZatoSKSIA8i7ybXUEmOsM20sJHGkZJwBpB8j1iJoiDGu6uigbiUUOgoLu+o7mz8VFNlTLlLdA0w
cb2YI09xQ8Tglbv4xbR+kduz319JfbH1/O7Qm8pgT5GRLdxrAlkS2AgQhbi/qg2kwxHRh+h1ig3e
1V+GIG89QIL1YQJlckFwn23lH8v3tdDmefXek8E6QGmXiR+FtFSyceZ25kFjB50kdxcDGpJnLWHN
W3SjWgRRClkyW4fat1Kw5x+UHQqA8uhG9DPWX6aiH2kwmFG25Ky0SVmi05iivkphKLtVhjNmAnia
/TYm+CelAl2FBT2jONaUQQnsklbN8uVjpBe9eQar/GZ9cGJ0BtgiaXXlPCj081oRI7dQQE8HlyUi
vD2a7TSVyk55zt3TftNSHcV5XT1UsIoy7A4LNkevcbYrhVhrO8/smX7APRdA9zdrhN5LM2+eq00i
A3mayIpqeslWBW5ZKxPTAJpE2QAHjaACNRj610PAIBZBzWfCoWxS7Co35PMb7gOowxwxrN5bhPEl
em9DPAhGGLZu9FPoJzclDeJhLN1KUvQLcIuEcDjfjwfgdf6XJf9fvun6arPi1NA30vdXkQfCIAxQ
bBeRs5iUlcs3jeHRSOEJoYJj8XP/SWglc4fJ6ciZih0e/8/pRoEgo/nnkpLa6CkcEv6cYk6bhufH
AklgtoV802Stq0xUG73c6VW3vi2KOd7ay1zRknei4lqOa7FuI61HCPZnCGyt8IiTCWuDhRX1SkXH
N92yw0vp+CNVuy00yVVxvGGIih5h2jk35kU4qnFCmQscekWAxWi00/UBR2XhLs7b2dQNQqBlyrbQ
avzF42j77Rahx7D79Yn4roCxUvpuupHslN5JVejSgQYQS9Mv0TNxX2oKLj4iSrvJuA/cvSbzjEpP
9l5PHiDlPM29KsZn/oQW2Mcm0ohvoKe+aL9bexChTKvAydDka4ekTegVwGiDEnxRL8mSUzwWJQn2
1Ju1O/gdoJBAvduKSETG9uC6+imFoXmFt6PFisTum8rv3K7oTGeJUBaQOq7qsLSb/uUsRRivnJEU
Ijd765pvIAmNkncrgsHg7Ns7tp9cjqVIUpmzEqBQrZ0/MgVv+rQIrkWlDgfpyT68axi7ZnpIupdf
hi7H4ZguemX3dA2xWlSDpeb3ax4D3iRk4Nq9B6GcIGXsX5JzpvIBjhqTbU6rZEtLpjqb4QYHwYmV
ibZB+xex9iuIevlhCb7kLXOhNTJ3HnEpgy3vQdOvP9zFX4nzijqmJGzLjb8eI17Z1CK4/1us9Bdb
66CU7aRf+Btc7oXucPKjSxNx5g3V1JbjI+o8DsTdjNnYPYjc9P+eUSQZAqTA0MqUPGWvBq+SR08+
C4aqpabbxWJt8LoWJZfVWE4BMIl0aD8ZbsU8dMcH9oWBeNliBVPBPHEwx3HUThvR3MV9Uz+ak9RA
/uEL/mWyl9Xg11Zi2GhxLcYOw1CUK1/29inuD0A+eY9EI3GHgKFXfSVPdZ/rwp0rVZFELZT+wv4+
8oDetY6bc1rIZfPKmOzvTeBENXGyssG/fuXZ4Rd+Km29PZvWwf42qT85PqOcE0RYMzUETYS+wHUf
zTE6NDaRADDjaJ01Oe06LjaiLYCybbvopyTHznPeYcQH45HEgyfLqnZA8LnqtLAFXPloD689EoUQ
xM4f0xWufIE6XHs08fiQjSeaIlRJiJg3gxiChvXReqw5Xu4SJ23Yiw0ZD4jGD9/VruQTssOg+mj1
5uAfp0dyX4ftu/HKd3KBQqnkpBLBJZwncYl5fJkJCGDoytMTIc+3yujuaaky0+F7Fznr3kkB/P9a
QRe1rdzDvkRoDDPppHK0ubPG0Y0R+XAhD0rXTtnTpmrKNMfBB/K8VlF7wrpAy+ANSq7PSccVv3vt
xFMLq7Wfw3+REZmtBFImraOUt+pb+/HJxhl6fvB2IceoRm0LWuxq2uHOdLcXY0qORUt/wUPbedcd
Y3c2w2oVdS7QKEKzSqML6uDT18egx4d8Q/n8sJ3GLAFEsR5hzGRX2xyCJ9Sqy/UVMj08VNiTHKlO
oBpFjVTTHOLdb5Jgzx9X6D6EDuLvdOwBq2uH/Kp6/Oc0TFPRtwcewdS55p8ZXopEOxIRbCWckfuI
JQFFItdZMRR9pFgsyv+fD6UUN1sL1kfBFeZbaXDtBZ1a1JgLAvZWx8aeYujYrEj1zgpfhhdq5MAC
TbJIg/PGd3h6zmExJpUYJ5E/n/m68FMnpa+XWpg69IG3oOAJm+5h48J2QwIWVEh3+PhviZ/psClz
7BhRm98SqpArz3hXknaKgfl6dQaCHmNP/Ltb57ga+2boHrOvXMWwDj0Oxr2eK39VySYsePCa9PD3
hiOndZvjNXj+ZTsvUjx2g/Yvy7vqO3Zh8CSlXwYRVZew2RK9El86nn87NBGfbHzXB/poR2Ug9TEZ
OM2+pPKXLOwAEguG5T1lyxnZuGpnAVEOAS/ylnNGFbOBhkX6Zn/Y6ReBtOuUF7AL+kEsAMeDzS0P
jZpNOwIxSMIegMZH5ClFtzVqAuaqO9C9oHZifoNndkAaalgy2xNJ2/rx/OKfHUX+6mqvkKzX+gp+
olOpxZBPpRDNogwIH5u3nJ9H/TfPo98qMLQNaL68e8S61MC+LeStiURlOflrxQtzEKC8amncmGda
FldVk7oIxp6fjE2AAgMPHP9c144oh6CNNOhEn/QGgs2c4Im22m+CmBl+lJuPxVA0JiqCh3uCbEXT
twHdHoZJLIewYBjT5Quvte4JVHPUjkvfOG4nIHu5Faco1OXnrVXcYMtTo89WLTW7LlCUFRlMxfQd
onCLWOcqGFX5cZvyxFhstqPt7lo06loNPNQ/chR61tizlCbb7GFQ54LMavlCoiNo9HgLktmkX9zy
1UPz8IwRdqkMnoa7HaaQ7NEB+4p2DHGd5tldB/ljo9XrUxHIY3Mejzd+9QCPx8mTSr15kugUIv4Q
TopzfhOEf5NNQ3i1gh2ezmnFAV4V953a0kL9kOlGX4/9oM9m9vqPOaTELnpPbVHyHuJfCg2t3RNv
AlrtIYdrze4cMzvs4jvjnsZ5ducDxnsho/cHtLZ35Pg1ls409QIYsf9KhgHBro21HxZB1zP41Vy7
76vf20jmqY3WY7Cg/CtcPtRnU9e2ren7kPORKQcNEKfxaID3OYyxkS0XNvDzpCnJ8/V/emjvfrbR
CDT3rrXgAV39/lnlzKeRikRda4kgCYMztp9LsUBrdPU+9kb7sXxt8c7tTvUiEDEbIUVpwLCle2G2
yLc0Jj6xK2MXLvSpqz6ICzZO+F6m/AI9UXgU3Afg9NggYKqzj1dUrvYEOTBiJg9Myj5BtaYX1tqx
+JgiswbceCG9i+wC9+ftHJQrRpcjo/j4BFz7u9dbKGam35ytE5mFZ54tA9udsJ9UY5EXVu5tI16W
dAzSGbxnlZLD+6kFpYo599ksF8RMyWxqbDzDb2A8XyfDYIue0vbOpZY/F/iKfL29AMpdy+2f6kEr
rNg7KbGiba7X1LhREl2CcahbdvHdfaNAhMj3V7TGRh/MyDW9XO/dNDfOhfxe0Oky0xdpdDEOCHJ6
q/YV5aVo6TAP6UQGuVOliQih8Vf78NPG2WvcBRpzpKBeWa1jnlh5OtQZt6RKif3c1Y3x+9QGmRPE
bC1f9ldLGsRyoznM151Mkkj8idr8kM+D0TlP7m6k6yXMiL+QzJt6ozLiD6lFLmCzE3Sq5+blH3M8
kA9LCvyWn1yjOaKXQaCV1P+/mQ0IDOKguVjpgKFuup6e49Q5q7uVtSZlo3APw57ehdQTkzy5ghXw
68mEOk8lyGetp9wslwvH0ioJET5sP5dSHrqzAiUhraDrFojsstUmQ2Q12FKOILH1APp8ozvvwLSe
qyZ6PvsenKta4zBnriFu1oBPBlZ+Ftrf3sT/3gRmbWgRCWI/Nd6/1xyOMxz5zknUPeRSHQVFsj3N
zzfBvK+VC5C0YPLQBtb6GTlbjVgsgmX9XsbBSCJKE+N9C2Q38nS/5wJlou3dPO20ojknPn8IMXV2
QdHbcPuZLKopg65JMxvONY8bTowyJ2Gpug2XXFOA4KUZyDsbpe+5m8yOyNDRD1A6TmOzVx0jEeU4
Rbgk5n1FfYFyxd2zPC8ATzshvuQV1cEEeYqI5PKJ+kofv7cTc4J4R3OsQN9TDZJZVh8TrnojxKM/
OvQtFrwmkd8nlcvLZ2Q3+YT1WmMnmXdrsF3O+SxX15vA0kh5JyQh7obQNdAsEPAIljY1MwKB8fwX
kkyTkKMsfa2YmhXfxIkebtF1d6RG8v8+IR7wHSD3JKmfIF7wbGiHlfEWM6dzDvWNFYBgvkA/KL3q
xWC3hUL0p4IL1L7UIYVWAa0FryY06cIE+U0ZbubOMOeQdL0coZJfiVPPYvgzF9c3/fmo7WqBr5/m
mgdI7OV2jOQiQfpyMvLu5CtOW4fQAH8eX4MfmhLtMtTlv6tDzsXrVFmKkFpVHNgcsw7UVMUDdoCC
bGi/+FHaeWZsI7PDElOmpMrbvAk1iWlhpLNts14pzrQgdL89Wq7agd4oIhkv6VdHwCgwc2oGIXGT
Thu01CWjkFEjDOoakEXlL7TBqO2Bc6SYjxMOM8bj1bD4JhTDuboPq9t2/e/F96ySH6MFGOQ/Lq+x
KMNKacY6IdlolqWFC9Pd4ggX6xUaGFsgoOnmjw5HvIwaO3R3cnSWOVSV1OaXdsTJhGXx1x7203/+
b70WbmZBMH6R6mcpLuQ478smFDSP8xb8Njl0k1D3IZHbx57l+gHz+eu77dztG7NpTLHfNnPO2xHo
JdBCONsPRvePhNYNJPLsxF/UpVODiueVdfWkfIh+C2XUTAjaPa3Mwy9X2q4z7zClB2OBky+KG5mw
7xDUsiXt+w8a8MXYflAnx/IGdffpbG4TX/+PLeAJjflBHiaMiYnKzDJhqkYgB99XnY/A4032kUi3
W7g673vTRmyV3E89pE2xNplS7S9mF+JGgDv/jvAn22kRguXjNmeAo91RpYtNvOiwxP4s/Cgv9fDa
RuPRHBWGsDv648oln2uLh0PAEvMoFJmOovL97KJ1pVRis6mt6wYPBaUsuOx5LN4pXAZTYD49aEra
+bZ847Fr0qkYjgyNwYkSk59oGUzheWdg4x6M26oRzUzYOxgNZGoihNmdfTdJoBKlMdGgpfkHHwbf
DOWrdEaa6D2hwlGYnYSxgJfRB4NdpIGE/ppytvr3Rttc4vbMJKukCDQvm6JaD9tkjS4/x1VUu9ew
okqtvV3bOjHYHVFauUIqMk/bRHn5bV+XrXk+E6FFwdtAAWhc//+3FPrg6/EZAs4i1xHmWq2pjTth
mEo9n/tAueGRk4+nmMaBlUL/qRLVjuCKP6qevDERj/QldtXURxxEv33CCBFHcxNvlI6vzyw7AjTP
JUAfeKr+rC5ylzQKXC6frWCANTh3HKdrlh52u0wnslVGtzwXWZTChtfp0nOaD/kJLb4icPA6M7pl
CoruRYlD6FRXhsISaQljlKAP0bj7+HuLayQ3PiGyMsP18eV5DQ8Ta+tMi0tnmw9xG0Df23oZxLP7
wMadfkInTR95VlVA+8tmGWgRndWAcrPGst/j2ljMnvRXpUqxJCyemMqYzr1QnfPYxXrtHUsutZAd
za83MiB1kMMtkKAJczvv5mLQzRgR+aHB7ggmMGW3AEsTBdP9mTb5I0KuC1APhpJKWjsi4FsaKU8I
78gtZEC5UWls3VNFDKntchf8H0VtNlVWScIw1bcNyDiY1rEwxSi8EEYxLYtHLZOWA67zoK7oG7LR
HcEPKz/5GCGiPa+VAE3VvnUBnP2rducHgRDAA5IUtodNj52/wO4GeucoUjdTpheM73LjFLiLqyK2
EWuC7RPkjU3RiAyj1WtF3fscxtXTXLcGTdnbbF6XiGEQeI4pycZyZljwX38Qk34SRY/PqjkmCxqt
SLlTiEd2RIcb6FCQn96nwhMLQA7zeu5nt4n0rEC9VFOjOP8UKYclk4Gm3+JnJ5Di3DEWMvMFPNpn
Cdnb6GXL6XMzQByBzTrnnqjrairq8/F54ojO4k8tj10A/KQgRAfaNMpQm6UNqnE2jyB9pxjaQ8J2
DHIuZOr2OJo5AvzltmpdarZQJDb7CyJkMGdgteUxdnwi0fWUXaKqCO3/kPYnDatJjAnPBvpolgjp
p72+1EY3xf271CjPKZICzfOllsj6bSrpwZb3rOi/X1aPEOHq6Ss37F37n5ShdwnFhrXGbVw2WqkV
5NFqtS6qR5/KEcT8Gg7MX83hOcyVNHzL++Ywg0scqlAgF16PnPeHwFLicn+aEHVBBPyPcV2oO6U/
uAYOd9gKZ2JY+clbhsUQ9gimSmWUVUSkuleFALzCNGsw2Zy5IBQPy6cDU+EtUzHKWdCi1jtgTCU2
Z+bLc4wcz/15CjKv/39bidw8kIj7Z2nxhN4vI6B8T86iIAMvI+G46cuwuWYbbBXSYKl1ig6Xr8xq
9BZnapE6ALgtLx4SWqJEKT1gzQ4fJqYSCJ2QGDyVyNaz2cZ42t/921r3ddpEupv3ruRU478XZqGy
3frw14wwslvMaYgbj+9g52aCMaXJ1NTtadarJRMMpH85LS431YmZrBZQ1d41weqaEok1rq8MeABH
YCKbVouny4PAlp10tXrfRs0Pq2qO+CoGb4+1+2QseDlrb2EULpHazxtaeIhj2SlfTuHbZob19tEv
1QDgOjTFWsW8C843iVnFUXX6sIptD2fouEFo6sSbai8+H1WNmUlCilK4b/VFdEa2RDKRqViO4QP9
sK9Chwr9pVYpoLIOE/LedTrpnYwurH8D+QVSijXQ5WddB5fkjfghc3c8PMaIf9fQ9Wxj9y+sqdpz
UzHSbCi/8CP8/xZsnKngVmUzrSsv4GQ6rC9HCL0BU2JQsrZt6txNjMrj3TRPQBCEnm+WkNn6wmg0
aG1Qgd9VwdJUemBba7XuGEG63qqkLbRAjhrJ7ifeHWpei12fIVfgU1b8xyGh+gqOElJ17NoTYgrc
mV882z7knfZbGRnIJWXPOYyDVXZDxAMudyEobJ0n1Ypg7BZqWuGVC/BkKKvkdccEKdAhiTuC7Buo
RnXO+z22srNY9jKqEx24dvRUNsqimlMrAScAUmkjRfUDI7+v8WvX9Y3a1VAVR/bVI8RQqpliq3BU
QsxYqxTqbsBGfcjdbYn3Bz0sybFn08Y4TQedpTeB8yV53U/z1bQti8TMmh2E6nLTXeWAXfvn5DAn
LezY/FJ8GpwI+/LZbqQPdSaKJ8xXr3hCUJtU9U09GJNYy46UaSdufnrahVqVgoFCiLiHUfxRy6tL
5PHgrT3ZTWWcClt7vck6IZOe6loRBNJD4CXkS6VAkNU+G9Y6d27kkPwNeaQassRviHb7/XMANJu/
ihIzQIljF4woToAUZllXakl+1H/7/FBUrbOJwA+jEU+ps+gT7vc2vOOrVEFfSjtZRpaDiMYE7Y9O
zSO9ni5QPpsHDVA+DZdsn0YE0agouHBOYjHk6HWVJmH2IJ2zNjB2ewECp8lt20U/ftIFhopDS8H7
M69c4MzaAVi4lobNj6BPHtOAdxTqQmtfwVwIyQczIHFVWOl+n6YrJxriUDaWk9LsJzGJRe9RxS3N
Ii/myRxPKsOyaJri1rDsIXgkGj+Mem3VD6XhIOp6wQsAYtBCl1mkDPugArzNy4AMiCbJnqOthbB4
VHtIhcJ4HkSiTZES4Q5PGFG6ElmCdPZhNMWs2pDi+d4FAjajWmrXNG/GYNcBgrvJcnh1WuZvzEUp
qfZy9Lk///dDdw0yFccIbRRKHhmAd9bz/GhZ0XdHm+38VtFad+dwwBe71RYrqoUO3Tt/fQLyOnTM
0yCoGaZONE9uEEezN1/5XmtxX/j9kSNRnhBSVS9ksgNvGdYKDsVFUApTVAEnhTbBJv3gfUU52KT2
NkAkR8A1J7mGcIQy/6Todm0sb3v9uvgcdoFFK2d/HOZQXZXhaZ8myjLhxeS5Bzp9sUs94Gvde7JB
CkC9oZklxelkA4QpY3CkaS7hZZkFMOcWbMP4Z9qc4RsdIvS37SVZqwBVZP/DJj+vw/+fbNG7S4MH
8YuBWk9RESjEPDicF9//AfeKjZEyOG9hbnGbcBD2eY8kXIm0+s/NRZPauDKsP9m5GexU31WKHvjs
XTlneKp7u65G5WFruH7/We9rUk4bJBcF59gX0Qpx4HBTW3caxU7NbzsQqcvjV1Z2mJP80kDIQscJ
9dfa95JY0cWDHOiwtUHxPWYe3k9romCXrldbnl8G1DutBL69tlBJEPa+XpRd6wM0uV8UgDHLRHp3
KZ0acVjTzMn6OuZEZF9V89CHDwWrUCcV0+ORm9ax5ZORkf4Cxga6bYvxwF2XdF73jd25LRwj0c0Q
mnjN9PceYXzZ2HuhsZHSC42wpamN+HCjkagVv0tRSL36NjEvQsqDcfEBVQvKDyec5S6M6IwKILGk
ksaXfR4guJwFW32DRh+TxONIP8nPgUlhp03gPdktRf6oWpHF11Ybzvz55y3e610AkK9BE4wVL8LJ
eC4/VSpNuBVpAEHOVRQN32TX31QMtwZVgx4ZYB6cdPgpvvzdyuXUnk1j8FcSY6SyDT5XgyZ76P3F
hVf0Vu0DtEGJ0dqvB/DKG1PTrfqtBr8KBFJeVYtSUndvbL1xIi0AWu78YiWCFronYhr4p7suAXfZ
8f9lXnYVqvxHNcUuYjWvRq74OqELo7hkz/b2etsj5SpcvGkFgJHu1gTdsmMS9YY3QiKTAi/tt3AX
KEa1md40YwPb1z11EEaPRQ2oywheMzevz8Q3a40mzAhxZJl6PEghMmgnvsjQ1piPxgBwfjYv3mN3
9kt31llfbZ7BWX7pxJMG0alKUdU44t1b0VOCY36GML0dIbMxa/Z8p2mezhCpqWZLRFqVaPXac/gK
JyCvOMiU04nzHVZxvM+WwhpziHnLefhVYUyJV4KVFsxMyphNpOSeSO/9E5dmmUZrU71aGECWjPti
OxTSrF6FeUCGuLn0BdNWRgyoZXzKX/1tamP6BQGUp0ckZU0KrCq2Bqc2cUdNsvdKJ/DNcJTM8DBS
uesrzDGwRqvAYGj94ZbAeiLrRWjy16c7MrTDGGNnXOzyBDveuMfI9n7DdW08JMRaEqE7saO2P4H8
ZR3EPcD2OFmAVJ7oDzFhtPRoQBscBve2s8BDjlhDqXGu5Vt0DKjv+KzdqjbDgvfl39HNDw/TId/U
kUJV+SID5Nt9IrrUXuCZXc8SFxkHX7SB6Sr2yJn5IEoneCYRQWweYSLYWa9qkksGIHb4KPUuLKod
NhYzWhdN6HR5JAWlyZcl2UtKBWeAzN2HIwDgxuX+IzKhqDouZq63jBH4FVj+AL5lSuXcXNxAsi/c
QY/sp3CHysqiKmFjv3/OjuiTl3xeteOlnZrPsEeQCfyjKtd4VOxv5I14tWmoYY+6QcKhPlXVhOjc
SQqbgV2gptuaZnc0axE9g19w5k00E8fCBdLzX7VjRqmBnAbdzGEjD5EjUz9qDldF+J95d6rTNmiK
AyW9CRL1K99YzGDjA7QaLx09LAq8jptrEklEomB3pk+Iqqniab3pj9B46ZohuYkmCgYYG7jalZUS
wVlPUNeHdTq4nAdbOUvsqhSw0F4Kgfuu4fIG0UuLbnXHB2z/kWlFKBCcJCeAv1w//Ps+jX7U6qnG
bTGAIweb4ex1ZXcTAeh+pf8m5Kr2Zbraah81dP0h14l2NTHI1Bf6ULFszrAM0wJZdMD19FChK0Wo
Fy4aNd6QUKlLKTycJ2EVS0HvZxXGae0oZW7msg0ZiyCYM3nE6OEWN4MgLmwCREagJvoj23AziHxu
nmD7MDQIIAZgEdoemH8LSJbD5mtx40aw+j6AqfDiiFTp0LinwnhgQ0cgTfsCjPqe1qTsDWdIu0iv
J53jKMteYo5QpsdCNTvZrHHPPuSRgCNGcFsP3XID+SQJZc5NLvocjX9+4smnltZmEJVBdBJw22+k
2eqM+nFQnKTwRoncgqDAmV2sdcTIj4cfSS/VVt9+B15b93oyrEVyGYDpEhaT2NBR/fJD4KL7XFu9
ZffYN42OWU0jO7Vco4POfpSuKdH+iMONH4JzbefZ8eomDVLIbDjDU0/IJpmpUDRuIlSCdxWsOfy4
wKHo4UEGXoYp4FufC+fH39vJ/6S03zqqQFAMjjVIeroc0zXm1p+Uj0GOjs20Cj+4pc+jL8Alh85V
6iZ/a00nFzLVfurV8rPM4Q2QM2WsaOpfHRhf2cm4eQ/v856GwRdbvwxgvgJ31GgcI6UmbGiJUjwK
hF/fJG36kpBY0dsSNm4mP9VzTk4JjnelkTbOsYoFjCIH2oLlXRalNbFRba07VkH4/Rvw4a4ubUFm
gnjEttwY2eY8lYp7zK+u7P9kHN6FTFNgIRk1p0/W3tsdu87QLe2tPlz1VU/hx3Mkf057F+Ifh+XR
varoz5ZYXUYcYr3WlVMhgPo7Hhyo+WsJfUW1mMHHSQPfOIOCRhxf1rqE+zzPRjVEXAAk42O4LvMu
ZCNwtntHPXAMkDEdLmqOWuSglWG0A4W8ZCZ0DFLvGA5R6pyZyZL5T8i9HAkqK1Fygj4NglfBdmag
4dwbzOfuVMgf+62BUBYJKXzf0ZqDI2FhOnLb5musQES3kEtpvsxdXmPeB/8TA7RzgY4ce9AWYNDx
BSXRf8cfiLb3Zmsm6ERPurEmkRUj6Mu8cb5pqFlRsiII8JoamkLV127RxG+yWtvmDInL5DswT9VP
gktrWixUfEBHNB+mK9wGrA7kKsrVreX/8eZiio5g/ig6EUClSMqHkzTvz6Ili82vO2+yQuII09CO
M5geSsjQQo8FSIR7d+RyrkDgjAya2kgBjfA3URyzSmIXkhiOs87hB0oD8jtyZ2RFTyPGe79H3kLj
ANiTigPijNbiaKHon/LtHyL//1GJjA0z0L2KrgYiuXFtGM+X5UkK1bhR6X/VrJfmVMq3e4oKj4cD
9Z56DuMQ3u39pCcSvjC0Q0NqvLXFFIEK53qaFJzcXLLmaeFPeZ92D+jHL2g5PW55eXckEyXm+vy3
+toGh6JHrJqmeQDHyNf86KsFTjS1a2SAQjWlWYRx19S4JknNMBem3CoruTvmkATH8DWS5mj7ydKa
5fTV9exr2eF7O5WMxoJgDb4ttZtmycrK1Njhp6XzKvdVFf4O6h8r4mQHbNumUuhQRtk5vaDuW9Ar
LqcRhUlCq31em3Tp+5LK7rEhJYID70dtH54IRoeDVmqCrMTvys1HlgH3xuL3eSOSd8nv1OObFV7n
XJyW0ntwcDDYH1xgwg4K/aCEca9smGTKEWVOc4RAHe6LjO4bk2eAaEAWwNXlYYth0t6X3TkkcbCq
/imwUVR18q5Gg9DCDsc9ltMTMoRr2/BxQ+EF1dpozwFGz63Buk1RoLCLmFDdQZ5oJ4zIAuGruE9o
8Fa51llFuOjqJD5H7ljWOIjBydOxm0abt44g1P2RaSNHpEXb8qTPGSXUKjja1ZEB1m6Knvuk+Mib
uVASFXVlXJJzODzb6qiRa7oKkv/IfpoxWSx46yRWfH5C0JjT4Zr+5IWjuZlc0arXyNJdvaJGfDn6
y8XhLf9HZ6+VbacFDlVs0JgIu/zS7C2kd3Qvwk988vV53eobOmfL6U6Ax8odtuJflEcaGEUyXGOt
sG2EadnHZgQTmJcGV8z9iO0d9D7f+zZv8UWDjTh8Co5Et8KsSaN1bIFNT4rl0e9YjTjKWloYLC+b
yrtGtofp1ThMM+ALdb7JyZW8pkf2s/LXG/KdTBPiRjvgb9n8G8KtyVFme+lTHDGKzpZwwiGgcUwi
zJsx2CBb0Exl0Em+QKEauX/jKK+wk2//LQSjZt4/ctMINf0WVRud0GsLpxXcFXBQuEiz8MFpU2R1
fT8xMi0Kc5DHxlcXBnhyd/f/lgMlFyATksNG0dzoE4b4bJ5CtlCCIEfI53bGPWm+eLp+YqHm3f60
0qEjELDfYnWf8wI6uTW66JY5NXUAW6hapctYG1k6o3S05wqyQuGgn8QuK7h59PYKLy4s1DbPpXaz
OKTdXv9mF3s4xY2LxqUSoABWM4MiO/nMFb6viRT1UYV3B6TkMkblq6JGUfARLy0WRFbAWoWoSI1n
Y/m/kPVmRv5mJyaF9ivhl8RYMPf3KMaWixUTbDZOgqXENMb4COoXbIwAvkDZQChe1gARNcrkhqqH
T/gJqZgjJ29yhKgIu1VhfthwpCi9FYy4P+DSQKqN229oMf6Z8Y9f0z2KpqQmzr0PmVQ3kefpKhCd
Mg2z7SBaLqhriZ7bj957/2irsqYsACvOnvFPsA2d1ZYqxWyDcIp13YNZyI8zONhAWydllexEs8s6
r4zwkohI7xp/+nEklI3mWk3o4zraj0pZLy9WD7TOvHMi09CTTFExwtQHyVxnFNt4ggWG5ue69/lu
jhJ9hgcgNYK+eumwOPOJtWi0aOBEA3ehlN9tTVDVhN++W8NNFotswWzo/amkxI4pwtx9/Y6NPKD7
P1555vh0JVuYc8NcxlGgGdsHIfq/ll5wKIWVzGCiaoOjxXv45KLTNvIOHy7FZp2cZOYlMk0w/vu1
Eu3BK3LA8kAtcwzQl0I0xgkfludnp1QUPPWeyZefYBvzltBT5iEwQ43l/1KmEPbLHDmPK/ayZX5y
kiklfBj8yivvccFe9e3NXAil4RwP6VL7voFAcGndU/pn1wubcp4vR8VVZbyGDLJUPW8o6tuL4ELu
xpvk4kkITTdFfnmbN4auolzLI2zjChpWZwPVzZMbPGxm0hdGeGwQNlK+Dm2fHDR5RLf30BRyIRjk
qalgjes/0MLqHy7bak8dqyRKe71wamq4JGuvulw6j3E9K2J7jvgZcszpa8OPCQdkSUn9Rqvagv14
JnmMHwgZBG8xD406y54E/K2lFqpi4U3aJbJr5YYINJYhVTGCt5svd6ilna+/QRgoWV7VcBAo8ULI
PDDeNHAUIeA+DGf+7Eg1hFVoSiPV+E28DYUfa5o+NDB9wjiZNHNGqXAc/NmS9ANtP23V6SEVSLvg
hLWQVVv9wVs520k/Vo32860lyqv4w/CfIVji6eb1q4gSIDc3YwxESP4xGsyI/lyt2oQDQtjeHfGV
hzZttnUCNRGSCIGDx1/I/2I/nU6Oelm5EG8CRNV1qAFmp0baEklvbarE7v4nFe+/8zzYNCZZ2WUb
IkJQwCn6Yf6U61cGil7thrZ1pIl2ToqWxEXqkPyxUZ1r1pl7sHcUBhCGHuH/YDRV8FGnD3pMiuMi
ut96J9NGWU5j6j67FZncWolAnRwRZVGoCpdlz+nMRxRsTIB8+DPu2J/YeGVzchvQwQekMomEfaQy
dpAQS/faFeRcuk9KJ74F5Wk3XcsxmkIulmMJqo5+12t8WB9BEyjQmhnngzQR8YvvsdSieT2RuAFe
z0e/S8CrNUnx618GvPf5amTCrG6MtZBK2PBvr4DgDQC6bNkFRUCC8qvPl6H+12Pjghd4u1HP8lFy
K3JO6rkWy8bc16yy7dG4aTFIq015UddUmysco5AZAbdhMuKHmGW9N16ayB9u2VJMY8Gs1FOv+PTE
AqDBnH4sMg0v6GFoc+dQJHNd9WdzxwQHFUGEZgtIXFMJ69vid026aeU6GOqiApERFEuSlKM5xJDn
qJ0pd7vUkLDWhsD2Vlrkpc4pHpL6xgmWAIRrVOBZmWL4Ix5jhMJsKl5ri/5VqGJdLIc8XVpcDCCM
MzCvVM+Xi7rNvST46YS0xS38zBoFiJvt4X3NzUFu3CZao0XmrriRq9S/hBkWKPLcEQ9zds7ljx+6
0oI6seVL5C0CpD9rfsAwYSq7JBc/VY5huE867GblhdEtoNIOUXNZlpLm++6Sd6c5E9mtdVwUO6S/
ezfc+EQ3O0NHm7Idj+cjdyQlxsyYGjEOOlWNDIWZjK5mYLQ4GwATNHXG0OHiN5IhyrDEeKdxKKo6
OjWQyCSTFjSEQqWEIbLz2zQXS7KPXmlkDIuaH24qlwZM5hTzSaYzp7C6vYP5rVNA3538hyEeTotz
AX8zIAhMNn6WkRtmu9kbptTr17qEj8eYb+JlC77FxLnuTLBUzNv/xyMhDoDo2jVduLV1opFOUov0
4kz8f3mlZRDE2ctemikkI7tS1dNxaN5ra/BSfqKMSm6h/ivX7VQR8YmhGasH7nNOy92FrbQSw5q1
OxAoWvwhDpzC35KmORPgRnEWY3uFfjo1c5hjbC1Sfg9ONSKcMs+NAOoylhhEn28pvqgNk5zeXH03
Vj03v7JLuHaMAO5pmu+m43AzQyhuN9MQd/KOa52y9d1kXyNzN1x37ZQVPgKSTcnQGlykH9ke0b+u
sC+4C6aGMbShr9JRAdUvRUGtmZXtb3j0L2lmhUbvstAnlPZ8Gk8S7ujbgYhoP3yyGg++xOsC5x+o
rRK1yueaf2QkpvAALfjrzUbETzeZEhIdyQHm9Ob5uWd/PEdOyLJOK4kTGB0AmiyozAqO47A0ovPL
1tfa47LCYiHbKCpMi9mm3R2dNvrbc4Y7dkODjwYaaO0PNpreOu+ifTG9BeuEgCbD2uaXU5y2vDmn
yprDb8dyhl36gt3etGJ8IP2ph1M/PPp0eJOIpz23pCE9zWPE1Oxm72okUi0lMV+H/3cqJPPrYzl8
Elyn2USIF0sVySbJhXTsW3NaFIoz1D8gRplsRqGeOodZHKfrJW1r4Tmty0eAdgMPujcOYVCs3ra/
ZHGESdDliXJrJm3DxiDf5i9y96HhzXY3GXNMXcB909A4ZlDbB6bBMSAAYGL9k/FSs4vgbWMIHSQg
uQqzE6bR72E4+IkqMK/qvilWPHl64xURMI9uPclLqCllHBRtLBQbhNp11SxFmfe/MPFskWuZJkSN
Zy+4tUIkytcNMcdqAMaw4aG883wTGPctE+JcsrdJc2SCslNgb5kI8J/e0lqXHjLMWaLRRn3Jv1qk
xhFEJgDebx7XtZBNGtRQ2YPJkZlDVXCrQYJvvb1W6ZOkcZv3IEPYEdiSPKunfikxmer1CmjCAqkx
HjGasFOPnZw2gTGMZh+jz1OwYQBLS1UkikqKV6AvoChtWjCeAkCwBSLBzcXLNZpdbqD4/DO9EQFW
Mwg9E1z4iCti8i0/reMOgxuJIKl+KtvV7j3gun7+cZDkdhVvXgJGYgyI7NE5ZYSyGRdib2q5JUDy
WxhcYgq/ks4PK0CldhxnANJ+FVTRP8xbF/+gHOsEmpLB+5RODJGhdAiRfUEvGqV1eCxnw0wYRSxl
PtooGITOeI2mqWz6NcXDUd3jBjb8uu/TsqiyU3gQjl3JLa/eRTJu49LET1Z/ZBj0+bpLW0HRnIJZ
saNYMYWpRDyRFY16bV+51D0E/knalH1vTJY8Mq109IPujPsXwVZMvu91eLEjrPTDRFloscy4A7Oy
XSEjBYM2p3Dds/TOM8OMZxFa6iH9ZLQDnNqWvmmbnfVxBBzROMoy2FreMsaPmYrOw86ydJhvclSi
CGUdj7AdlBPlx5bI+DTNQYmibLNBXeFvXL9Hkdl9ReYLNvST2SUqhaNBu4OegIyLkE1R48pbtraH
h5X9UsUy4/zd7VtHVGsN8vjGiDkBCsDIneFTOLt+m6ojMhS35NBziRAF3W1K2F0QJOvyCJvl8Pqk
M71/JbfG9rSfhuENzRcphdMbaWbDJwuw0FgVwzjc+K+g7LK05GQ/dwt4IJX0Vm7q/a9zZGrQM4Bd
ZQBDqfyMr4hFkCaYXG62gbaf4Y6x6yvBoioZKk66rQq2Cq0l8YxG3J1TecTBjSy0muEHkYBaScoQ
yHT6QTCGd/9SYTL8wjI09H7IWIlKDe40jnx/uGX+Z1dcuFwe4fqGW/rCfwW5p8kJhAkR/l+/IkJx
XM4Yg+Iy3HRHoZ9m8r8xkHoPm7oIWusKzPZWCJ+LlNb2GlNFtW52SaCx7W8p+hqhWNdTkPaaQTBP
K5oQ3QZl1VWphKpRg7b6Iih1rTe2RJFXeMxlwAy5XWazaIcEm0WfSJC+bNPyDAI3y8iV0haWfAwQ
01bJyHAimP0SYpqDCWfvz5UuIdySRVU/Dokbsp8Zpi8G9/BecRZjqsUaISkA8htEeFw3ey1G5qh8
CWGA6/k7KV8fWyf+zD7Q8GC3x735rzaMVu0f9yKYoKYueUrWWVp1ntUQFI68U/N7SdTEv32ANOmi
SDggqd85qPqSTP5qpjV7WjJ1loU2jaY2LXqsUGzABCQcMM7e2V9XmzwH8WA+hcxTLBgI05QgW879
h4aGHzvu9XV8b8gZWSIN69XVpQb5kkZYpntR22u1tqbcI+X2qwY3fIF9HzWMKoJ+HmqN9j1AKsIV
CRQZX/AzPI5YSXfkjHx6Qu/B5VVSQtMTG1PVwQeBa9lEhArywYwBWlZjjBUHvM5u5vEJoK4D2pPe
cx3nbsRu1DBriAPc7R+W1GZIzl6PdUH6LEGVEH0TJehUPQilnUTCSMxBaR2jW2KXBYmGS968USpU
KQNzi2Hk9QSnUVqxoTdt9NUETIjpdQmiiqqYXVML1yzfrDmwPfXJLpZsTEFb3CXO+wyfkcyIOAHZ
8oJdsbDURQhviWN0oqXJJ7x+7IltWg4itJM84HXPGs6cWulv8c/7OrqqpSdFrtpMQI3PY6ubAdsP
jznRiOiYKRPDWL64qHdhNd37F4lQuVv2llHVR8B5U+NuGY1X3YgB1aTpsA6taZpALsTRwM/hq8Hv
hdlttovivrA13jdydaJkKlcL7cwz6NZDMHhk7WxqRXaI3vPOh8YnBiCJK77DtrZlZiK3HEkXTpiF
LI6btlR56heQ3ldvz3YxNoYh+hLtoHUN2vBkb5KEspxe2HlLZecbkPfbRSEJj8G6ZJbkvxJ9Jo0/
z/wRREECUsIwYi4r4f9my3H4ZrdeYNEykRmfFsEu/+hd/LJCjf1A/sYNiZHfxN4fQNJElcS5UA09
zm/517Ww4HK6nZ4O9jqTjol4GM7jmjOE7xakyzz5xg+Li2bYImcpDfHk3chMG9eAsEiTrPn82uYZ
pJQldpoRthNYsANaE3oNu7d9XTPJX36hoZcc5tYqWOE3zCYdLoEWAPGs1ng4Ws6ZPZvD9T+9tgv/
Z8oEEmcovUSdqQFQ0uEOVaiLQ6FCQLDzuf2cmkkYImUbOadrBu/Q4CT/ZUN059G/atQ1jpTsYBW2
wT0NF9JS5xZnTh2uuS7AlOfFl9r+H0CqJiqqPPwe2TCNrnnQkTh5vdP0461TIQepJWh76w/gbYv3
3qOy59W2BzjyAxlrLGYeiq4uGJvvpMeFjyTIpQ2H1mj17CFTdji+5DwDTA8zOS5ZZEY0klttw+Vq
DGqEkRtVYKlwuc6UUcX+quJZ6T6a4VhniF+VQFH0i4REbJma0aZnOcZeXTpzOKK+sqamSQ0FhNlY
0SsRehItQ1AuQ55s0SNV7Z12ZY3wTwGuZ9g05q6QkuQHhp29u++Bg6LK1ANnnkTfEXaMlWCFGhRq
manlOLT/nInhm67d/PvtAVFBJLDzD+89RMLD/+1winjJiXYQeY1aPQTr4dIo2aHJ58xut3ecch0K
vT1R2wGam2+T5E7UeSPXO03dJUDEMX/VpBuGBUM2RLbPSZjFbGCcXzHyKwf1TTqi9hRxrNP+Kyjb
R2YwgK64f0XDRWP2GwLXNDan2BTMN1a9ATjtAhbxXjxMfuF0orJZWTeBWca/JKmUOQS9HB7sEYLd
GXD6mgJBYct5owtaFCPPvftjQ48rk6trI4dGIPy9X+YQaQdXfUvqvFrfBZM2eNOiCL+P7Dgbpmbq
WvE8vKD1Bi+zS6YUN3r9X+ncsi1wp8gTUfqxmXNqaBe37i2ScP2EjtWtIHKyR1C4MNiCcZPtTzmw
ras3tgHg93l4sqW6qRhh2p60B5TVDMgJUZPxbglYbVpbwwnTY2LxeJVif2JV47+x0xxldOh4ZF62
Z9Zo3XboHwi6CO07mJ76IhkAVkjSAIITmRSKIVHMnRQQBdY3dG0ICx//DYA93Ro8AF3RYv/n+A4D
T1V9S2EPazPIzjBbACtt7VIV+VQ31RFfhvouKPND/1juvQ7xxjHeJSanpMjShOPPz9fUbWA0EDFn
mOt+ywUeoR/hThJRmbqXAr6JVWprb9WDHYUC4wYnVLJWAgoaUceSEArEmpUDVagIwz+aFW7nU9kG
/MOGlhxlvh1lqtK6unGQ3OjK5+9McMJ2XcbJLKqJ1GKexb38+tLmguSWCbKt5IBjP4YoO6F5hVnN
QsI3wn25s5hwOgq81tJx67MOoyvRdaITWWY/tQ+ZUBfwqkxxr/cRyhPMCg7R2JFysTus71TgWFUt
eLdRrfwW1gqLysRCAndWV4lbrrXYGTwhXM2I6kFLyifJnm3EDuhbck+ZdGDyApcFI2cC0Uy/tUwz
3QdxhD5YQY4F/yNdvxZx5ez7stvhpf0IyQuntuuTBfQbU4KRI3jGXfF0t6rvxlMk292k8MYoUzDi
np4CYSXOlx39REd4HjM7xq1NanzAbPsNUPIaXXkbOI3jLLXKP2Y6hmpKkkfd6tcr4BPlmH8wc90D
YMBysbKdAsalLFw2jlcMug3t9+XA7/HkV4JrXf6jM7ygjETOslAxYxNbE1fEiPEXmjB9+GgZ5TE9
oBgWT1DjhI4Kd7Ux3hSONnhT0CD/LYRqwqAKyovDL3EKQWg6xhZ958PoIUS24caVNIUzZ1YSp/7s
jGuCECLlQzLL9b2O/elbxDATJ22XWkrYVQpg9YT+hD5GOaqPBJkvz2PEyPcw3PlJXQqZVlFxnPHG
JrtTGdKTnNCzhNzXQlYFGbs96e+Zxkvrvan8Pbr6EMnU42xawTn9MXb+gB/82Fxddr01gv3AOgqP
md+r5ZPntJ3z/nNMcYxVlVejofICGXuHrIrrA0JZIIMnYoE855+t3MNGJDblu+ZO2Wt+qVnGZ0Vq
wa8TqY2toTM5wrTk+ARUp2FnxlK7JBlcYZc4sPE/qpD06pGVg7aiZORj4MRUCeCzAP0+dvlkZgMF
/glU3P6JV56weIZOnIuuAWZCShy6PeMYEq+W+VxqaC4fS1fk9EROOoDPFFTMpw6GBocVMpSdbDUz
L3vffeb3bWrRVyySNRkE1mOiAirRXJWbKrt6F2wkElIPGsXs5UCGyKVE8Qgf0ebBbKgT3rJfh7Nu
Yd9dGPqgo37EtFb2dGdeHHhIyTU0PgjxEPIPXrVGSSUz/oqoKHborgYYkTGDaJLXPGFBHLB+3e46
7KeGmo+XjcNDxg6BX8V72PSX8kcWGTcwKJhugTBka1uR2qiGMLuz9zFtj7CGQm6l78JJIpseJm3F
DVqR/j2yNQljDR8aaEPRgXjLAvunf3GD+HkZ9N0Z0pTi8xb6nvSh23VCyXajOFPJ8eDkt0V9g94c
h1EHtQHtJjr3rUsDi6CA55oVCyL869uEAyxqP9lAfeVnTOeVG32Yj8DmyItAyesDopIgm/s7fETn
6E4/Lf3k3boeHQSNV/YYDoR81UjVr31WUyyCi/jPPfYicOYhvC3bLAGOAmspPQnvKlisNmsCN5oD
1p6e/hEU+C52yWsKqdNCV9TU/K1/MoFQc4YDl349vWtTku/8G1wQCcy3w2m0+zL3/m3kuJE8aE6u
cY3nHVUd1Qeh0kEl2La5x4TGZQ0sboV7KPrWhoh8Ql7ObfXBMeWtaaOJETMYPNPUb60hTX8FcD/L
p4Noq24RHYhGM2bd4XqG6jJAtP+JH0slWTADaQhrm/LZ4UsvpIVIxbBQztsXQPhJ4MQWoO9ETBrW
D+BfLOn8TRdXYSni6p85xuL2G1gKY6WwahFT3mwyqSvcel3PChbK4ZuFmkmahcI4xyF4SGMSu5p8
zj7XW7JSgx2WgwLcNtjdFiJZB5rbKN+AleQeQE0BQz7KWa32i+VZhHr8eNrMo7uKE0cgUlTRclsY
KdKkePEF/3kipZqjKa3f7pRV/gbLpM28Q2yVV7FFWp967BYIub8GL9Xg5ikiO2NN2hOR1QO9z8OG
GDS9wiLGDH9P8btFyj1/cAh6NpNkH8Qh3vf0wq2Lezsy5xQ517OhbCLS1xaF0IP8zQupfWQhzteC
i5vwDj854bVsBHpWpLDJZ9hG1EY1VFcBZ4hjQn91X3Rkfd+95M9gJ4baA3QJOtNXt3YGn3B585wj
JzRRGjJacLKOCuiOeQuIBeaDHFJGexeYS7ZElIbIY4BQTDBBX656ezWaYFWpt6ctgXzqQwZHvfhF
OSOLiMNpFvSUL5mhqC0HpCJaBoko+zPTT60UfEeKDw6pCoLdeCCfMpStyzCh1wTkiuxyS6tXOL4l
sfB8ACj6dY/7EV69HBp4WFsPdALf2Ov3BiaZLEWrjuaqQGdwhWxNNUKDre6yv+P1E8hv7gdX2pYU
EmyPoirxpxvS/MK4Vox7eeTgz4AYYxHPk+S9VbiT1lTa3E/Ht2RmqaZWt56lsSgUhYrCYuW3UBVN
PT8djdYXRK3FiVHmd0jY1dsd+W3vqIRaWt9QuE31tzTTLLwX9/uxEaLDpnEYuaQ3pRP0Esx6XFo2
JyvAAxLised7waaxeCPgNC/jF563a0iGIpVesrAahyRZxKnbfrhYE7wYi+OydHUpR3GhUs3IZHFD
emYz1RofwOPLqOzRsuJwTqldTcGNlhb7YL1CJJRwLt7/5pkS5avUOBY0D43qKc6Aoj2uQQ41Tw2J
egQ+DtdZ4jEJy43BM4eoI4Fb1j7CyPJUMZj2ruiZtN0c+b+UgkyFE+Eu7VmBswADTvRxYJJIjj7P
p3Kg7qDEpY0GbX4uqo1EcGzKJNRlselC5KUwAeJiAPmzTj675zvGxBzULB+qxgPvjYCcS5D+I0AD
cfz+YQr1mevRNCRjloLW4o2CWR4rp1je/REi6/sUx7X8j7Kzgw7oST3rmNA5ZWjmLtqfqeYLR4QM
+dEbzkLh8HYxkWdx2HSyJKoU/qLjh6oETgmfCqIylBJFm7yHnxxTaWPwNp8KQW3Qzs5x4Q/Kd7zK
h5lCf7xpVbCSTqOp8xj3vXHO5tJaDaKOJOfdw17zjcnDXum42UqESRj6bRHwYAJZiZpvDZYw0WeB
nAC9zElTXpaHwxf8rSd/wOKSp6uvsy0h5D3XpQQUK7v0fR9hIxAcsXTyqI6yWQr4Z5KwTL1GrFeL
Gsr0gaoeu8AYHgLQqShBc5hceUDBOydteZuPUHJAxK5hrVjlZcQmbjmhUdobDauvH/8vB0wC4thp
3csLvN5D1F6m3QkBgGFAek3ax2tqqCXdlZA3K6R92YB6frTgrB1I7TFMPU49V0fbh2i4LxAyZ4vG
9v1pJrFodMxnaalMEXjNfGkfJsEGbN0t2XYDKuy6AFlXMqVaW0leixf43lx1/3C7BkJQlXcKN6yM
U9dTf4fa+xbJnggKHBANOHUaVYELxwE7yKb6HJwVpEjm0IFgT7ESrj41CNF52VnAfqNYxUNhqb/J
XXYcu6zQpWBbxGmJxF2xl3kKONzYNfJ0AGPqCUnBwR+ody9xpZ9s51G15WSxPzjh8AmmuQ16tKrT
u4MMR70toYYBTMx0s6vgUSahwPqizPm+aq3m5raYkv7EY8HY/1nrNEubBRWfzdlPv8hxijinLc6S
dLFe3jvIVvyi2Eta3y/ItLIg+1X5BmtSfx9nKdcUndu304HlfNcZTx7/U1+aTs32qlVnlh3fHL89
5heKBAiRw3Bwu6v1QLhmDkJCpDhtJhw4eXQ65+CXwx93NWCKDPSUDpD93tiS9gYP3aPLBpcDQ8rr
i0xGsCvaEzRsjSgYWxPZecLi5CBTx+iqkMaOB7Md7c1PPzRyeKO+a/VUJ4xsIK+CqVPEcRd1tIFm
JTA0wVqTC8VE8yGlub6X6w//q2HEIOPBKAVbejZi7gZ5zUyoWYnAG3dplwAVNAc0xRiulQwAagrp
/po3GtqeH0ddUC77+f2IT+j4xFx9GsLcDrnZQECWlZ0GqHjdQPO6y2H6HNqm8r07lG3V60ejllCc
zu7fdjVn+vkCRdDvZjuG0XaBvAMe6hy2wPwDjchmq4VpLKCzqGhiYxUone1vjjOsaja9/p0YfizY
U2VsDAhLi5Q7KOtiYYSlL/aSmYCh4EAhzzhXYkWzJ6t6+HpHe9M/XH7uqslcKF+rvuCcV6/o6osv
mnpT/RQJKFvhLatT5h712zj/Zy+lzb9sNiKeGpiJZmyof9idvAEonYvW3y+c86f7ol4nW2r7G+1M
L8BbDyQi7OPxAkzIOZJrv1Mmg0TK9p2bCPcr657xATd8mfIEF+ITKQAIIle/MMbwzLvLW53CkPpo
H6z2XbvhqlKaSHgDiKPkMwHDYJszcNh52UQ3uZ5losGUNTP+L+4KXVZCSQBwXIcOb3yP6wP4b4s7
Scx14bt/yohAuRvLLrMsrmPlepdlzmVAbmaoWvuDurXj2T+wXN1vg0Fy0ceV6USZvJmppfTkICVd
VhLi8E2mIbC+fEvhVWAo6DNxsww1QPmq+RkWSH7rVoC0cYB9hZ4M+bApsfwCx1AAMrycTLVAtiOL
fHaIhj550q6dOZRhdQqgvQ0PCW1qN9sUDFK7AC8qpDFf32fFqJrrav5CrXmYo+KTwUdX8SScV+Re
tri/15LZa3XPVQhzDVnPdV32R5QyUzaSc0ET3bOF1APaXpQr/pOi/ZqKEHybEj1W1+Oqs0Hw0GN+
WObS+XpCb/I9hDEywd58IYNKT12ZvFx2Bnt+yLZL1vI1U9rmEduWXFAC+rwKCSaypsHaKT15SVsv
u4V6zsBW8g0Ni+fxomSaeYJ0W44BVD8K4CnypCOLytUOPjkqiVXdVsQMyAlCK14Rvbu1Qdb1yX/+
j7jumtzTraVJMgQqDPFOtFNGk2EAf0nwoVvMzwNt6h2Od7irl8Ublp400PjKj4RNbWMzI/wX4W/6
pE+XZPMXmtQDheVhU1kauQ2+iBaVBmZe7CiaaI7Vfu7AtoLbWjSkqs5Aan0EvHvrlKof1zwL8jtW
Mi14UWxMtMMsJLuTH0VTBEA2nQjTwiFGSW71fKsa3rMVhCtZsbKSbcnlju4mmf7pKzWabJ09ht5i
4awYXFyAF3NTPhEJYyctJwM9G/C9GEuzzTLcz1TU7l7p5+Zm1hyVRHoGDWlrJfEeQmZfk3nXR08s
M7ymnn1avZ2+jMbyVK5IEU9VdJlq4IjfWei089bQWMyfTk9KPdag08oBNB/XqxdoIJHKRr3f9idV
nBpk2ciiO19MFsrn+WeFD2YezishomRIT/hMg1pDpdRtINogNIdrYyrxsM/GLIbXgGsq3Q8MjG2e
ZiXYwR03/eggI5kuYSM27AU23uwKiTj6q2ojXUsGpC1fTmUrt4yomEvtXGu3wwaD3bMKVVQn9TGK
xPBT6I6NloIyjZNEiymuRNtWI40GIBpE9KKTwydmwiDyEvj8ADciSng+6xzLuJvZFHNM0JwZn54M
LLRkffkp7zIHJdnVpVBVUMrSC+p9rOQlht2TlUivdoo97S+hQtTZs9pMwlmEBcS4WAWw9w0UjoZS
2PUmDRMP4olL8dwmeog8pAUVr3uXEJIMkJOExwqkEMHNrtJ4hBWNkoiW1W08hO9ZJmILdXiHTXk+
17BTJkAwGbunoWsiyjPmyLWwFzNPEVBHYHy9XKMcMbEt6l24EAHHiYNbT3B8COuUcXvuehDZf2or
usS3O30lja7SHUYQnUlRJSkQMDfaUdpfXqvOtmvO69cvtMaplXJVvSzI9SOQA/fY3fKHMON3/8Ia
zOBGwJ8uJzzj0LMoItxMoZeJaslcvEyWZKkd0FW4vI+oDNKfPaeTh2vfqlv4WgPEOhadFxhVt9hN
lR+LR+fkV0F4fk3Jw+D/Paj0bDGM4NJluw7q+UgHF/XNW9IPzOpV9Yd43klQ26itGjWS1JUW85IQ
BZvYLtcqDN0qEyPgeUXhpReYihJutS3BTs7vWsiK2pZsQ8ASeuj7L2osxttwArLwkC9Z59vjnB+/
YICKhFwFxPPSEIgPWcz/39qv7g7m8To+wr91W+qvH3dHzFTltcxyJcttpk4NG3DlaKb2DZWAtSoR
ogj82X9ikitF/oVYCKgxT76B0eGmrPj2fZuBc3/bcuvg8ObVzv9R8+PEsgHIhCDkcErJWbHcaQS4
IAnYDBccaofeyJV8JpOsmvQ8IsT5fbbiwS2zx48me9Z2h38xCZpGydFHLHan12UPbZybKOSXjtob
uF3rXi5XaEl7ydqX+TxTx+f37sCvRA3/JqKMlIK+bjrtihLqF7lMVS34Zc2hb6yDNJV2IatCMbt+
lGrW5VrQI4daqlA+Q1qsuhP+DA8AhyUzPfbh4z6OSA9xcE9q8vkfllgBWtOgLcu02dqCRwBuZEvt
A5rS/Ifbzw7s49k+fzxWK9S3sLkBUkjjv24FJgE1tTvfgwVj08hXJh1fTC10AcZCEsqNgWg7HQti
0PIUSgKIHaVt9XzrK4hxQTXGvqgtgwxZSOiCZzHPaDToUguJLrepPF5Lexn4AKB34GZHCOLL0QqD
wgQmaewqRlx4iAOcLyWEWGdalvC1oFn6IlQjQLNLR+ujZfoU/FSeiWkwVkGnfKbyTfOkyHr6ZZRJ
39+9jUQV14A5epv2+dSUZeUl4g+cNYblgQyDWcQkrSw+KbSQ73zkqaZgjvt44BACxNhCfoE3zjz3
582HRO8Mvs9aGK6RMSkVeh6eepTxrJrBaKuJMglTlTr6fH6KMAU+v4G0PywXoFF5E3lBd4W7olx7
5Ik01TuV3VWUVCSaiMY4/Qig2/hi4+0H7jyPNgC3o3szxonauU1aRiUaHCQmHZGqtX2y4Ie1q0HA
GqvVEBYxAjxCTkyBvI6aikCwkwTTmt8HG+NsP1fywr/CkiGOy71VnaD2wWVlEmNaPxI/lp38FcsQ
3NH+10xKQSCzKE+M7jTnuOOl8phcQx2KJ0CiARxAHiCnJAu6cC/0uLliEAhGJxgpUif35S0smyxo
WOweeq/sm76OoSi+ues4X8mGT/NoPyfP96Iho/yyYfcGILhC6gpBRuPqv8v7ZLE9DXBLSm30MfpT
j7lET6l9ufV+qgY2jnpQaZ07OmJXJ2u+Xlo0a1lxwbpefuQh2UHw/8o3bgRoxqUTzoh7m05qVQlJ
vaNRgaeTh25m5vAETIpjIHoF6kH8WfQLKtGP5J/MMUlz6+IWUiuqqrXV+KBwJm5+XLOjpHJUzMq2
Ioh50zmOs0ymjroZyvjilhTBhxlFoi2J8WojNJM4FiPZGpElq4hcsLYTIivpk/Pca6BbpcIbcQ04
7evb3Y3l0iCnkRO302GOWjqupmQoKgJf8tsHSOhGfEc0S9FlFNcB608c96Mx9UyPX47r+vWAxFUE
/N2gQ4Rs2lsDaSaQwXcsOu/YdfprRkjWsdN04yxHs1oqfN9JZGmLvTki1q5bS5M/eksWHH8LZRuv
zZTUHzZxdNh1eJu4dH2VBqquQylmyv6/nV9RM/WeY+2KQsGuFs1YBsgOjYRWBcpIQ4G5RU9xKQzf
w7WpX0SvjKEzqolCfqwFK7qRVojJCaTsLN/iElCyrL+4LqYp0+Sj4e9DCO6F1mKYayc6pxLn/rr0
6EBSS5PTK4kZyYt6jmC64LQMdG9n6WsA8H6VC95ROD4DAUSdJ8h48TVKh4oXYJHZeKrh7F0q2Rml
8i10YI1cbXIzcW684db4q9YaxngKubpht3k3YIvUnYz0tz540AHRsZqs7HY/PaKB2Fi10ThfujQq
ueV0gnmiStkG24b7t/RjmhJixSlhHJiEcWVJ/uxhzrQf8vRq+os/ATz1yTxzkwnTPpF//eh9gK7M
Wb8XMsCE/23FOoZoA1oov3LkGVzqH/B045OQJE6uWrny0NRxeI55IDUmljuQSSGtnVnCRl78WENI
eib+kD8h1lDLSmmnEUmBKOugTBmiPWwFZfc8fbUhRrTcrK2RpnXjXqvOPGAtb8zpOJ6BLsgN4cyd
c4VL6K9U7E/OQkwR4r4haUJTADOdzPfiQ/GKzS270QkIQzl+tkDiEm5Flo6+982EEZog+kL7nqTD
pWoKAOZOIq56/S8YE0cuGgapT9GQiw2ZENTZr7AN3GGVqKKJI+kEixAmggrflAwtI65RRsipJ2rS
tg+enPZ4pk+Oxk7Lxr11qC7pXNF7hDa7pNZvKktgq+pip9Y2P3IXTPuJ7c48pkAcYkBJ+oeXfeOS
6owu4TKUK0b6s5JOMyTQzFDfTh6zUMmaNwgaCUlZT6MbVgAe/gqEhfXDOrsGfcSrqltS2kVFXFWr
HcDtd99yqnr/Ur1zjph7G5PBUUrdV8mlJfa/DPgOZjCHNJKGLKeJOUvU8Far+XN/IUQaOyeRyaOX
4iFUomrBfTDPtklnwJciI128Id7Df3IupgOuOIvz5bIG12IcrjL4OJqG65BJcDDC4YuYFUSF1xm7
/+sLAE/hyk/220XhS5Y8cAPHNT2jzswAnysZEQ4/0ZhfDB3V8ez8AKULw9rfZNumX2tU9flCFHcS
1O4wY05THJqJnWzsZM4GkkuX6A+4H7mT8tdxa7xUmQ8V7pexBLBzNEJKxDiBPFcxXawX/xxwxAbt
HjPVrVCvpSs51d+oJaLZjHtMP2Pcz6+m7xUGCKdIjhIu3dCneAensdOI9tK5+5RsFAs9Qn6kzi8Q
dSiHSicou4znbazxTFIj071uXo7PG7clQZGsB5FWJwoBy856aqEvG1S+K9pF3KjzTwwo5qVOYmQF
BkQD7PMFPNvFeaQKhs0+D590ptH7AJmQsRk2XE2Z9b1GLaCzIKrwaVi0qhMcnqrq0XOroGufaR1f
bFseDhpB9g79Ud4iqC2raaikqfHy1BUaJuXN0ljKuA+U3X67TqkrFAy+a8gfqDUAM7u4IfX4lmvX
Z8RT9mzlXrbtuTPID7AXzviPEwa7sDA1uIN54dIDWIP1NKdlcPSQOYWWJGkqleVHBiFzpDJ39Ta8
nyZWlYyizConHw11ab+4CpFKR3MdgST16IevGS2f7fF+HDVkBbBCUsUFZDvvK0LMKqqL4dFswBJj
X9hOk81TaRRvc0ywglRLtuCJQKHaJOV1tdTsJu/nMGbCGhJ0IhH6PwLUCHUxigN4THRoPLWdUtLf
L4utBmbRQlHXYWSgbp7t/gshvjEgMJX79vYe49LUfxNDVJMgm8L0Pch99YHZmcqXtypT+sltJosI
X3dx86hnEn7IUGsblkH3byTTBkUrFGVMR6pfVHPjjgg2H5QJ4+xd97UZHwuGAkzQMfJUaDtBg2IP
zKSfsTMDK+tHg7dDeOAqR8QjGxOsk+8hCuq8LSuQeqAExX1tqsOtF4MHE7yGlJv9xpn0+PF2Siw6
M0gjAjM+7inTsS9TGKMoh9sFJl7MwWji15OtUjLZDlfgxAB7od2t5Jnplbuw+GRbuMHGqIJPPXtJ
ZuyVCTHL4XV2hnxhCUrUjBuL1InIJnr1+msAPIXujrUWY7mGeUdU45u1pGwp58Wm/UzxgwxeYToM
KrADkdlh/zYFzod/v5q/Qy/cszRFErVU9kTuUZHB+ISenASw3biYyiKcfxMpDllTiFDVI4fuoP+X
aYCzoNxlf09eusIn3dJkehzjob/U+m5Pr6M04t0rXSSI6wsCv+iIV8Ha+GyiOTnOnra8AN9dR/Zb
d5T5gEuX0up9RdLHW2E5Ypo/Z27tiPeeH8F82cLVd9mQStsVHK1XjxKCI03+MZl1w896oYpMvjVE
FrJCUf7R4DIgoUaqDrZPncVPIupRsDLR6+mU63wppRX3YcYQVKyeHN6BUpwFu1KrnvVzRxLodQfd
w8qXaj2JWYq8POb/YS+v2StD1NWknZdW6/Fozko/TKJUSj1AH8BF8UeZsTiSKMvyBSEBUBwOCQTf
3NTp4N2nYR12hDnVWyr7W010YdKchtjFnJ5K/Q7yjKk22aPShVE3gleD4fYlQ8fNgX/etgfrOVKh
IEqIpUOHeCePXNQiqYSDlFqhBqfMhvzEZBQX82V4nCYMR8ktGN4YoSFqGnKTRRtVWFBCI8TdcJtO
PBsEFFL2GEH1SPWwaSKDYpHoyr0gXA09EhNII4pm8hZI+Mi7Cj59TKxciPvtZcv9MYvznTqPWZFo
E28IYDmJe5apbno5UzeN9F4TWga9e7PAsLSIZ9j6qpcm+trGD7oxqnlojxCrG+Wj5MLzeOU9G23c
ycmIYsIUQy3qWaft7cqDCLE2wAmbW4ip9UysVOYAaS7UI+xvkhSu8G7JePqufG25rMbcne1/5wLV
UZlUG8OIM7qN2qKXhE0VenL/VT35mybDAA4rljp+l+DEfA0HYLRaXr5jSKW5a990tmozmI2Y+C0l
ERTatOFShu+uHt8x9nnK4cZwOCvvJXgKXaFQfLjnWuLUWTkx78CDYr8iUQlWX/CIxE7HgiyNx3xD
zU96a4AcLqMysJGXOjNSczL5LNgIjJp42xVQBE43d4JaiB+/7/28JYTMIHww4j3WX/MW2ecaJ/BG
mQxF1Mw2V728G9qy5RzpZhBGv4YQsZjNWH93rxslIh1+cULfdpFZgGDFpLIN80KkTC+bjKvgNpg/
whF54SwDwx/o3BBcZGHzRE61E+PT0j6q7/IAHKhZNOLWrroSb4J2UqFsTmgNAnMvlFIaDmpkr2+n
3Fer1leBc25h1NCY1gxklm79hUYdLefPPQH1b1zKy8v0ngwzgrFWlJX5yVr71dcEy+QFSO3sx1ot
CI4F8d2gS0Et82lCNYAEIUyX/wb8xJVPj547olHMyKa1OCk7oAzUWRAlds1etToV18r2L0eyM5ly
eL5PAmIPFK8ESWwcaPbaOAJD0w2aNQELDNkKUMJvPmT6usbUbtbn3JWZlIKKn6d/aA7+XsJGHVRo
IwYVr4QjFre7Tis4pQih909k0FONX19gpIRMXMIEdwkqLRAa06WQIg0vtimD5DkCwWuJthq0P/AM
QaQ+u+/dSYuvT7ItbehSRU7VAeUBlpYKBymYL2MhcGxlUsAFLHlcmBRtks8xjPuO3xbSuPmGKPXZ
Af7ZmJn3qUqu4te+Z5SZdPSXUJ53EdDW9PtsPo6HRSymUQ75XMMKFt8zxCY01IZVnMMY9BuxmLLS
IaL5HW2FU/WA3wiKJ+ldKlS1/kq9IZtlty1pgu1uKQ1fIYrvy9k/uTBQdbPTRubi1Rg4Rt/ouqkJ
zDwmJOftDdRDz/WJOtzIMow+Iyxu53p6zOtrx2euY88duZqC52Dl9o/DrQU6xncD0CaFkJ1RXV+6
A+jkDR1yk7GnuvfkMA/n636KLukhoijQT/OSTh2N7BRzd8POUuMTIWmEr+yp73qUVd8fyBq8D0mO
ntLiRnvDxPbRMo/p6UH0Y6YwFqbbpE43kOYmos/GeEseSp+T6MLq8uVrE0yCkNcgeGYFVP0M8Ze6
VlN9feVmFqbvK6j7XJCxJK40ugGmMf2wQgyQw4TNNdcjlqJcD82AV70kKn5+yRNanJinWdPpe05Q
3Lhk2Vj8rxt5inNvHzO6naULSqnVdvn6nXqNaD8r3Aai13riZKMgnH8ZOZ/Xxge1aDIfjf8IgFBf
QOym1g84qaWlD47oYOHf05Lxt0JxcawToL8/CqGfgHZenDKG+agq/1sBekGbjZ7GwcXZSri4YKhN
IDkaMzQuZE0ZJsvLUxhS4t9scAR9xLP5gT9p6R3VRfCgGNAmJxZ8cjG5yD9g6TRs07m4Eec7Lu74
i7cjECENz8c/OZduYMtduQQNe14hNClhNyjSiHjf7+EaLmHn9f7uLZClkVQgf1lkM7nOSrwLIQE6
gsiHEUMYnMNCg5k/Rz1muZBHr/W4uc7SjAd7kgM1m5kR4WL60FXVTXA/DsXMLCQKdfEE8k2uJBFb
RK9MYqLgDiIlUE5X1yQL1X9AsxZ4L6h7ROkfRALcqKpuSK2x6Vtem6iGA0OgjboC/mJp/eaayASF
asGP3NzJbMnbvjxis/iCTFN60l1UAptj6kTOIC994Rb95TVc66rXlA5uKr+TEL4Fg3HN9YT4cJPQ
c8pC4ng2bbl8NzfeXE0WwoBRirIwtRqydjmAho4XsHf8Suq/0v+SAhw+xSCWgvyoz6649Aze8MlO
79P6dGAN6Y8cQLtp93vOPsGHkEeS39HY/EltpUrQ4PjqTdN+QEAtJXSIJgmjlQ+D2mu45hNeyt95
KQ6H6+7vyam11ZwZ3zV3x2pnQMEVLCA8KwGJw6y71W/D1asJoNOZ/X+0Rola/KiSMOjUMDY1C/BG
TKHZkzN3bXoZAb9/PURXDXbDCbPyK5uRpo3FeVJIYg7vOxrm5TL2Rr2+5bkC8pshfglITMThvvE5
EgW3hPWaNEBNI+TrdLdTxATOvs1Jx/RleAWwBJq1ab2ahRMPOX29jYGxXQmbaK+8bReCyHewOHeZ
yJPw8xlf2CfyXZ8aeSae74eaKFiBaFYsev3HN+S6EJsgsKmmZ6191d9h8KFB6PPVa2zWYk6hbroU
DFYpqNKiiW77f9S7s1k4brzCZTjB61fdSRheD6yazOhARMPKCv3IOpv0pWkwfYA67xlQmWy5zGY6
iXBI6LajYBsoZKGQtxBM8/+kRrcucYtemHRAgZLY3OZyUnxKyn7zprsFeVbrpTrP9rbqcBOwmi2c
G0oubW1Dkm6Tcqh8TwCs+QyrDnZeoLggWKRPcU5TXJWRiuOhAFHoeGm1zRacsW1nIDoC2pTuhaz9
oR/RZ6jh4SUNzmEoHORCqm05ASX8mCE3UEt4IppuaoLuDx59PfXcCXpoXUJ8TzYflpCE0jttlczy
Cw3Z+lHFGbEkkLnVC8hIv9Q2FpnEEXZZvVVDX0+51IxXX9Qi0lE+8u3w1X3shdAiHpGVap/K7116
nVnHhEefCeSzJnZTQEuMC/46kwdFj5ryDMUXN5gBK42RhiRiwNnHZJgG2N3iUlmA70Ui1fLVV6aU
VZss3WH6X1eEKPSXaGo4lgqU9xk8H8FyNXXdFre8UwvVZUZHge74uDTTbeewLmWXUDjvEQRZH2+E
S9KGRC0lpiY05Jk13NJWrRAQbmVEcSdivUG/ySjpGavWELk2hQ3Z1mAG9fcwG4YuiB9CCyttIpAs
HmTZ5OnO4L1cNdG37qufjN46VJ7RSygUCe7KDIMhiAtj6OCy3PNib18E69KoZZIYvgMT6sY3i51t
iYx9AYsCZ9Q0AVVTGQsZbn1i9KJq9liXw2TEoUPJb/Uo4Vmk6aHXKi9AbaHl2XlbtTI+wwmR35Yy
ZHvprsuXzA0ySzBGqKNGrYc4ZPiXCWOR9arqKg2XdzP70RPoK7WDPPaZg32acw+/T/bP6tfmN3Wj
hNlGjKEpa/c0iYYaaUnp+73+x+o917jWB2M05waqYbjR16rHD9NzvaR+n0hIy5YU4j2L/yZ/LKDE
tvrLgZDNZZ0owWzoUnX7FL2cRf9BiRkOfhNK4cbDGdQBe8jnx9+PF1oHS2KuTBMj+TJDIKHsUAkc
OTy4kTrRXIDVF3IK/8tVjRfZ7nRYYBTl1FojYcgwlXIUTYWgrX4tbrnvHBQuhpdRri8nsTJqXN1P
xQzwxWB/VJbCQOIvbM3UgR+bRQu3v4h8Y7MwM/zooAEudSm80dDnXufgTidAqD5u+e18zroTq3jU
9lvrmJQHAqJYHgO+0G1CVcJ6lDqvzK90XU9+r3O9/7eZjnQkiOZM1bYaNaEKPuDU7Z34Kwr5/cwA
q50RQ/zIzC2tN0QKZ096xnurs1XqIEPa7gMLXMPy+9gNTlJptw4copmrlcPJFGPvbaLfdywA5pga
BrmUyJdzDZKD5HLFYRaovOG4AJszLkIN8506JJn24V/S9R1OUSmkZHBCDjsZkqM2p2kmF8UvgW3Z
fgfFCXiuhtWT8WEe/BudusDOKPCyz/t1ucJt5ADXN/eQZtZJfoMaaTpv6VRunyBTet+6v4/V2njy
ESEx0a0wcdDfgZwwazzntkIZURcLOaXjYsGKgGK2mcyRoCWk/rY9EtopRCgNLY98QyETp2PW69HC
jofT/ULV8qGM0qLcAsFMFnJ3NEnOc3XRzbH854+2mq7vWfTDh7cTjcKJIdybQQBSYhRfGVQhj9EO
SmkKXm8VY+FeFPGnThNxU6aPrJ2bZtnNd3XoO1zWeCmEx9LlMqqYvl0T0PQ0yhcoG8ZuD0aU0atE
JWF+Bof+JxsMlbfCGSeWeE4XTtJ5ZhqJjHQ1xamJWipoFZjogMFKaQQIlW6F04aFNQR6SMjU/2a/
HbaCGzFX59XVKJdZ85C33N/ZZPuMJDAHvICUKoObgdMNLyEUbyy0xDdP0k8STPtwnBIHMc6wgoYJ
y3eZr+vn/+Xta6wfo+YszhnGfA4iJpqd6zJmYTQAWl9hK1HZY1AtG+IY7Kxj4CakmmHKz1v4H0+7
4rQQUrJCCiTbjdRkytC+NkWAVhufM7LLz2BovOa/I0PIDZdlzJYUUgahf7NB4bX4RCg2kAtZtNr0
n9fgD9vEQUrUpsHn0LcNMH34OrJZbv72W9YubY2WUJUeDTUJRMh4Mb+BMGOjG2tpkWC5i9fHls2D
CJv4qZC8EL8Msgzs61OcqusgGBpk0fR9Aa5djp4uf8jjapfac8uksELc6Vr41SqN7SRNktDewzhK
Y4+HVUb1EX/APJrGa7KeDrvxwXAbcWQ8oD6ZVL6XsVTZvGY/+JCThmDvuM1sPUz2R/tG7rSAHmgF
9aq7MYmubjVQz+BV04Cfvk5Dp/PDdaXCkjUBD5CfnrQAYLiO6/aSjVcaoAuS+ZFaJuvbo3p9RymE
/J3j6WB/dEK1i/jJKvR9wOEw5ZOGfI2wowJNRfwZl2B0IzXRNgYAmU5voAQyfx7WB0GOat+YQJ7c
FKv8Ae/W5nWmWqeTFN0KpmhwtSRlOLrHOSL80XhrAebGe9SnDeBOKTsDCw2Ln8EPpSAbX/Ha3gT+
EkqVoVx8rJCrhmbcEkKjuOLjnuvwD0f6MM8Ljnu+z+7axugOEQlUQrs8k640cV6tcsg7iTlGMRFg
244MM3TvyWfcxgzvRN3ru9/Hv0CaLMaRWzYpoSlYarAs/UKtrRF6YBBAjnLDAw1q21riu5WsD6mT
la7loZJw/YBNE2MO5CEMOoH8ZO2r5efoTbmF36EV1gGPpOJQr+b0r466uEA52Jkr1hiQJIqGi+rF
5l+jebIJsaLw6AABpHN9ImcQoWxLF8xfUk4UAeFnPe0U89abnxYl54x0WxmLVsm1EIhI3YG9UsYh
XpJs+i7J/cndbw2DbNYAHD3lZQ6Z2BZHnsypj4BmtfCzF5utxULUjA0SYG1/FSc0XWP9pMZIPzbU
HEvBrRFzlo0M/XJsW9eoxRzzkIVGUhxXX/6l1DaC1NHfSTfNq6eKEn+aiRNFdu+4BAHxsCVNq/i6
cSVIzFglrzpxiH+v4Ut4vNJYL0XVJ8pZfnfdy22DrMBvvTsUbzlUCtnXebOAoyF/+S28mU4rmPDo
4S8WrJ86N0Yc57+52qwjGhLUBkJyTr4iuJ/nGtZD1lJu0Fe0wiTPV57LT6tWzj9JPFaPiGrDgj0S
TKmjFTHrIZN8tfgaEOYEmUCSCMDeeGytEb93BF21MVckJKXd5QRZVMOTXWjPo7EgCC8akCSj8dIS
zu6Vj/RT6WwjuhirgKrVjy0OVOXZpXJW/Qj1l00ea7MrUtwWo5KjiOXskaeY+EyC+nasCFtVF4RA
SygCJS9JSY1corl0IaUPVeSRlAXZA87nT4ZF4tKSWJELInLgpyeTw6mXIMjLAVU9ytOjMZJjD5sC
01kxPKEuFjBEJUXAgkJSqYPKOfuE68Xu+dMvQVk2PaJCinRP+T4RK9+qV1sBNNlbsbvdyXt/kecJ
PhDTcO6QXhTCJRsr5CFQPXeu3Om6uvgUJ/yC1Tp4OrHBYztd/5W/4rhA1a+ZFvQGVBchMrwnhxia
nhxZPEeX9uwGSUet0VDuCySeu5blS8fB4kqnQUJnDWh+xlANkfanL2uDAc6LkAzzHDKr1LamOoUJ
clehJAkoGbWxY+Ot6dDCKQFwk2Yknn9D1CfyTvcLcvJywUxaZuMvnsRmYYhnLRONO8B7S/WY8IR9
gVfzQlXRRI+w2JxY0rpR8n/AKihy9mZCKVMORaFvO1uXJSS1LSn0gHnD5yj7Ctv1rqfASSEoiYAw
oUNETCMhwQtYk8NpRegYrfqf2AhM/7Tdy+Qoc27jssXnTYHH87b5qKMRY/UMxZjhnxMuvpX0cPcs
gHuo2Pmim0P9DtpR8eerVjftJXZDQBvZ80IWDUSgwSkLNlu5Nxt5ys9hBXQVP3D6orqOmcYJeYcR
3m6zTQ/rjrbnK4q/+z8PrQ3XgkjoA80M/0IhBtIj48W0Dy3r+o416ZU7xBQVb0g97zdNAvHH8ZYn
n70LOqLHoWTXhqIGI0er2ruVA1qCV73W0qcUoCIu4WtcAUxu5+ABtRCQ61o0y7B55kb+A6ESlad2
boSa6qBqD5SzYzA61YfTWH0MdX8AGnLst0yfSRU2+CTNTrkH8Oef0TjhV4XnxUDCkGSDvu4Kcp8C
ScBcg271OxSAUG7VlaTJ1CAJt9M3xwbHcujIu98zKS/BTPlB52VQK955tPSladDOYWcF2YUOVgEF
VsJiG1chmPiqD3BtlcZEqp35/8uC5TrtRp6+74z/x3gAO9OhcRcskQh0F4lcBnRf2zHSAVbe0sfc
mcf0olv+4TRsmZCodSBmye3XJNa3gQ5vymQVT3iO/SwGkAW3xXtbMQU2/2qeI7hnx0ZLoioRYwED
ZyJHdbpQvD30s2ukHVlVFN0aM7x3ONNR9zlRraKbSA7TimkAeO3GwsAKtfeQXmFysoY3aVbIqC0u
tg2x0MvUmXrRfaq1qSUXuugu+AERP9LJRUK5NJ+5bOa9lsdQdm0e8LtqSrJduWV9eIrd1pjBcO8K
jp+nesSuHwbbCcCGpeFiQI/cWFfWi59eUdFyYBtyTC9VFaShscphVGSYJ0AAw8WtlxrM9QJvpDgM
c7kx9VWkC25ngmmoLV5HfcH0UaDwhB9ZaGI8p6z3gY9VAkPMDA71Es7EQClHvLc2EOm/+PCQBc4/
l2FFmT7LFDW8BWICzAy/X1bonNWF+gyxZO3tjm1AAFHpcaHzUcogE6r2UugRRPstKj5L3+ZG3VPg
E4XEoduelJPlLuHHxNRGpryzFlrodSMRh2a9NL1+tL+nlX46bMCbIefWBBa9sb69o2ODLSqfx5zu
6ECxnxm2O5WwcbGAIGFWyUESHpqNaqQD+XYuOkz5ZqbEE0LZ4JNb42thdEffYSmYa3j5n5f8jDOW
pEnHBa12gz1Pd+Jhedtv0WecBwxf5cU4DrIt/thQJ5V2fKqjF+SciSPmvFHIxv3vhsr7iS66AYmB
HgZWQs1GvCzlg+geR25aM3szm2YWqyqB8Bc2m4+B/6xFjve3mRarn/6x1orrrp5djySwUIIKHkf/
aUDQxC6gMDzioUSmhrmYBWROyjbzMZtyAZh9yjeBVIw4DpwgKY8ebKWwUwZTSIy5yAr0fHPcYRa2
9/Hgqk8UCia8F1sPXtTQTfgJNdai9wbby0mBmsKwU/WfQCvYWDuPGLcPpFUo2cRuqly9FMrhVVkZ
C1V8W6OVpp+ElSv7cLc3JTqXZlU2Hc9NE+3pbxtz4V8w8SLY+by78xbw4DkhBOyUpwgLCPDq5ZA+
ttyxjJKs3eXXA30keCUAdf+JpCZAP8ua7MQzEy7ngw9r9qaXLvzIQTNxHapK5tMi5BShHYwEfDXn
+2hI4F6RxE3+rdCqk74Dvv6qn5neip/egpNeGWxHzda0agaAtEwE1/lQP29Jkfu6eEzKvr1PGK/P
MNGtaQ3+ffJ+QP0PxY6wIcJ1Kp9zHH6MjPYKBr9i9P3I4SSH8gBprRNeVNTVqMHBrvkclUPxj13n
OTEThVTbl13x7lvAAWBgJG9xFZpNg7gQLQ3o0305AKv+fqAPVz6HJEScL1DjTE3TcMvQqc4lscvg
qXzDkn2ppT2zS7SUs60VtDIFs0e7010npUJIUPjMGYhjTQ+wKWoFGXY0aYCbdZbA32ZjY6s0AF0S
MZgxqzdT3Bk4qijijAmNHN9mjlNAF8+n1iOA2p46sABKArhKNtvCYvfi0waJMFQ56lvJ+7fuQBUJ
+TtdZFkPgfusHCVf1fcYd1BbtiJWuRXi92KhY2IoOt7k6vCBGuriQtQs5yC4F/QaYx+hHQ5GWzZC
NZF9QnBXlP/exmUC/2sxVElj1IUDa7ZPO7TuKlm0aHw///AE17xErDEGiL4CQvn25B+BaWTqcM62
NbVHZQ/raJ16V7/QQM18uhnryusBhwaPRzMAsZV/UJqHPq3taZcWfrRMqrLgUYxbFCEjilhhW4bf
6boAa/RTGwMrxjUvtIaIC85vl2HGYBWUumoyZy5Or9wdNqkgYbwgqqtXcEdqToVouJCHa1Vy1nTr
+xwECOdshTR26gFI6k4o4Fm7TGSaiKU7/9xL51i1OWsBE5LpzylG5F0kzgSIRgmB6HsVuQpv8UOs
Qo5Si3udVY1v5aqxKmLLzFjwZso5EK178Utbtq2//REkM3T/3iIKB78288+FO1sxktlAkgr9EToF
5VYdkerykyae3fXKNjuo6MYFGab9+EPqQPnN2ZfbbUfNEl+jtPEJdDX0/fEvqeJF5y8LTxaTpeyl
kfuigptFKpSyGoDldmQZHAKMcPWfoO6wWy/CPKgKg0wnnXCJBJIC/8Y/EDqg32stabaA/bFkW1+Q
0vi78U2JajtJJOwmRO3bmXx5d+bvpAgJp2Zeu88dcDZvZfrV3XOivg5gtiTTOfQTleDmGl8blWX0
nabXr474WPfwlv12LNkHjmxLarAQjc6+ArOLlEhanBIV5fEaogrHgSJ9Mw4sSodhd40NiSfSmJfD
EjKwrRPhoh0L/ZNU54WjH15xYkKS/WruTkSVGoXrqDTPmcHFEZFGSutr1CiFPFXiBZoUeEGgZBqO
ogtg8RDgg3ti90Ix8rgBKUR/xb9lYH9ylNJa0qszOtPInbgLsH2b1qexpEGLjFSsx3Z99w0y1XZ1
jPykIXliQCRfNKkkdCF9pZ63sUVj08B16p1XrbmEDS71eYcksPclSYIKeg3Uw3to7msIjaUi8iLa
onuPP50cjw0OxUdnF4x0z/XzfKKkkbNFyMDs3n6sv1tAWPtDMjxj+WD4nHYUkWftNTpjSI7ZvDTM
zNpJQvq9tJ9bPhaYrCzdMy4RZk4GJyOSHEkoMJmCzjfCwIm3p8OMDX9tiu+xysNzyls2z9Q70dVl
CIb9S+98PD/3s/KlZT7vuV7fBreoBXG19W+ytZ1v/3j5dQPQo7M/Zbmp5MNyHU/ApNlrZ7IOrHi8
xFzOoT9MzHYKZiBuy4TIlxIN+Vla4YLOdv6ZMZ63HIb20RZY5jeQeo0ti5PZR9HEY+kTr+hnT4m/
uguTc8UuPGxD1tUDxfv8d2YosX9cXVqdzHb719cCDk8Jw0kJHDB7d87DQMQozJbBhv3KwVUgn1ff
reRWfmKOsKBmGomLWvCTtnR6uIJo+a7oSVMioMh7YqZEqFdGCdcbtUGIwMUgPVGj9UmCIIE1o74S
ro6GzDPXAdtyFUk77FfG4BMm+qK8tEsYnM6RLiN2XSq/06sTxHC6zkf45ij8VF7XbjKS2HdJVS77
ojCX3ytwJ/elTLsymq+uHvclPzzy9lHguD/NikG+tXRU3UAcz2Q2vWz5nrEdeDZBBUCaSgqMfKH3
i96/4w3ZlOL3ah1QOxAbquEEHZQTvWRni5YneRz+u0RAjbPdlS4Cq2FNY0wvx6ccQKDcNs8eJLYw
aA9uTOEelazHLgKNqp3xMYL6zgRScYpGQvPfLYTsxPjVUDk2hwlhsYf+IKv/K3UqOOQ1V1z/zKzN
m4r6z3FtdefwT12SQxU8wCh5yBqkjKVI/K5GceWLi9EuWrlzIHfir9afKSwS67Bjmxx9YKRvSMQF
MiMFXsim8wUAZAfWY+z5U31AmBMqTe6XjLO5tgtPlsp83+qUZlp9k7vMEuL6SKAOB9zOKCrpMeWV
OLQu3hCAPLFaIpBYABjniwcgdJ/CXrPPgw8D3E8iQ9R06Ripie7mPDBSRLqYyLPkSc2leBZomsNT
X3KxkUtGdWF+HRiEKQpYVIexpu3gvQp7Sq2yuedyawfJzf4T0Ddi9iIbZG1odGBpPdhpOsFbVKnh
lf21XtgoGe6rMj1tOBC4GQ0tUCdK4SIjto1dO1O6BYAvQSOIk8HqZpdSpHu0hUg62FJ8lPIU6N3S
Q8QrC2U8qFmd4mpMiPYzQUONpT0bZmJhM6SwfGlT1xBmSZ7cLByLccWXyDloorBTRAlpVwgMlqqL
AS5ilx/WgDsNbjh4xXsiZyPoHdvFgSlpUKwL7fjLZujwn2/lxu6tPcZV23WFJMreuOLBymTelPi3
OTJYHMgEWBKnOAkz1D6f4+70V9Eqh4TTgTYbQNIMtq689zi12SFfnV+xgdP8breCut0NOwjUzKkM
AGUROA3GDXTcHsKVXcbBTXhDjdAvWz5/wBr74WmVgO/SBu3psrN4Au4J1Fx9sLyzUoJ1g0RQh/s0
u/kETO/s6UkRViQyrDkcVTYUX4c/anxgIKnRc7aEVh7BOuho5FdKgzG50HJNek2mJeQTtqiu5t47
cNj9gSADAv87arEye90fY9qPFuPM8kTuHc4kcmYyAV3a0YyoIxEFjQ6+d2cN5SfOfZ1vD7M6wHRR
iSN74jXZqb+V3jx01W4H0mkBesd6UeiHW3GXO8VVJJ6BCjTZBjv5kXC8v4IcOswalNt5LVk7H80A
V/Cs640LXhb8K88AZaosyJsUVs9UATCvjFyyVbiVn42YzAnwh+ZGJCg6bqrtl8PZa7Rp5WqyOJTO
CsX6GfzoA8l1DDIaKNrJcgiGNZQVb4lJF9Myk5/ybiT1btACZKBOfRlkIfOPuSajHo9Y5ktkG0pX
qxD18SRjOnA12r6RQwPnqPiFLyfxxiKmNAA25AA8/szI5PWJgbanLWW+cUt8yax+eno1NLcJRWYH
/9Opqom1j2i0dwatS5M8RTtMyNfdxsihIsR7YcIABMNUfOtR3FOWW5J+wte8//2EpLRfFykiWAvW
j1HSeqBnhVSLzufHg3mF7swlWyLyRHmvkZfxm/1U8Q+0SWJLdr9K1xaX6JGWK/ZZac5Ax7AAfCun
DIZU2is0gt+yvbAmChD1Uhyw74ZFlyOyKMVnhpcOz1ExtmsUqYsG44C2WlHdnOQYbSiUode1u4XD
SwfjeytvyCg2lgUIWqkZdoYpHk9ZYIu+afti0ASrLp4aK/SFQTERIZPgVTPZ4jRJ3s/J8xDfkgLH
8y8KRFeS5CvBARAYdk2GvZGIDGeOwr2ELWKq6Z5kocNg5w6AWGIOC7Z/7QCB8Z4XoI+6zgjWlg5E
+lFLpQuKKWSb/Yq/GtzawMELqxYg2eFiNFvt08Zuok8sxYkbwmEclivC0UzdXWeYEnHRvgT1xvQW
HXMJgETK6wqnyMA2cTB8OUqLiBBPwP9NNS5f+eNasOL3kPyhyZD7MjX81kq03jfLOUzXLnMqdkww
XZbduqKBMsjX2diuXaH+TPaBxGFltzxBqMoOrG8tlcXRgZLmCLSI3Dygx+/LVAg7koignXSqMJxR
RBC7xkLyj2uypcGW12ADBqrnS1luBhmNNLO5HwN87XHxyMcA/v06a7wVZDtJy302NqR2H4eeDGtq
bmaasgNl9MgR7rU4DFtPmBJhY5qO9gmBhQvYsXirtti0eWHaMahaoogeCt1Jp5KJd4Q0Alhi/Nkw
/yVgBCib869z+NUq+k+g3PVxaN0EWtSA4P5bJixC6720odBRdRzVpSrvRGI+7tOZbAlfd5jMxOwi
udROGc4D2sblBC0sPkxOabWHFXKXJx6jhS02ABA2Q3it/uUGV3/KyqUFSX7bQgYqjfDr0aLpo3B/
gCDPId3fAM8EUSD+Wd3HzHj5VJWebaJlRT+n7aQ6Y2ukvSa6kNa65641CGWYtqmRStI2epYOzyDU
9+P7Pm41PEkvnweDQFy5/09ta3tvI5XICDZbmIfpVg07Vk8vKvawRjgYLV0AsbtMNiwqXKnMVtk0
QQYK1q0+gwk2hA1znHRx3pxd+7vyVBYgIMJeNGRbq5ECV3HQV4ef+Egc4qRlDx23WkgGPLtyZTwr
VEwrqLv+R5kiUCo3YjSBVSBo6pl3Ql5VMYnO5ChcMXkYjDSAIeOxZYRUbB+CmwhmFYQt9uKrcxdS
itEJIloJSZdXJawjYo96lA99Qj3Da8HwRlADBloqTx8XpanAss8obpBKTtqo13LpDkgMhzyJKRkC
rz1RnVU1M0RvniC0aTPmHEEi3J6TfMvugzjh5PtvYHCTrCIW5oV9Vni7TZzMFuy6G6m3bWqzcyUL
43JrmmTMG7as64oApuF/1AJTFZxU/Van3ja27N6OiVzCkuuce9N4R+ehGqfG/Angz6Hp5060VWo2
Rhv/YkJj91dADPJ3b2GOo0nhF5uAVoU3xVOwHIXirgKWQ1DITzAoagLt4sEQQWQlzhBII2PQRYO5
xmFKvee9KXmYH03J4hINDCh/HLRB+knrmG3u9dXIdECFBRKfNcqs+5q75lrAQmrEDnBHEdq2+tby
Vhl4P2ekdvhcL/DRnTlFE626Ut0CPGjPkPlrpgcbSmejhF/9PBpbZaIyi2m5yZx5l3/jH77KjQ3M
ET7DwYh/JLZZljldi98bqfduOEfH58klrhji9HGbEfXpOG42U1NjCTczysd2wESliLTVuUVXE8rZ
5MW0bGkc73ZvWN1NnpdVix/zL9kJLdQwi79aQrrz+aYnYwnBjuuUd7NHJhle9Is29T8CdfVKncYJ
1RCo56qkv5j8lsSgredRdaSspGNh0ZBcl8wR9z0qLvNt92oF13tFPY63OP8KBYm75BIRmUITbziY
THoIV9jozL8IbEEk7HtUoz9ZqNZrE3s5qrDINWRliX+V7gZ7CfhVQCDgtiiiH+SPSr9oDHWvLGur
Watw3Du/p1tcL08JUR++AhN2gSbbYTQmqlW4ltQqaRmANmHCd00jnxikQjBsOwbwbSr60NLRv0PK
Q0lZP0GccygCnzXTnZ7xMjE+n2vI6KqKRODhD25t+0hjgkhWbqHkD7GwdXkEG0UyBD18YLrdY4SM
QPuGxZZtGX2/uRXwqG1SUON5vH4P6Y+HEBC5TnO3u0DXJkB8QfnSkHxrJMqOhy31R79JmfohcrSp
5ayQkqi7UrY7ozE7wYJPzg/z19/lvrMsWJQdQW4krb7OQQI90FkYEm8QjvpHJKt7z9Hq3iUzKV83
LaFZyhBkgaTuNpcll/csHgEyIyvX2zM6Ea9Le1tIbHZuu29CwyyXxw1txP5abTpkFJJ9WniCMCmx
NqeVQeU1j8iMocpSQDbKan26AMgVZYkkd3/ESZfbG7lnJAjD4hG7RCFmipT1g5vhU8SpUEXARLp5
Fv6/w0w9lV1E9NqCybbROHcg6RSEBebQoSr761UQOsM9JLTzYiF3FHz78PNAlsDDBsw8Ih3FfAsL
Vju4Iq4v2s7dsSssymwXp7r+7EGckh1Gzcho/vhkxWjtJUOhcqthsmPIW28q36wA58SMWqCrdU4E
fNg4KxawEcAwWFJGO/aDWf7mLOkE4suwGajRd5fxjQ/Eubw/SGDCf9Ho6Sjql4Xe0KAOvFoOWLht
OE6SNSg8bYfePUWpGf0YYBwaxifUOdNiHeM8VzjRCqAQfugdhVjTYm3xHOiJ4iL5AsGRNtM5OASk
mKNHixyuObrFgvYVrYi+93pGRDj1tV9jwmznhmQIgUolvnWagRcdgQUN9fEvBeVlm4YYwTB4+Vqg
h1Rq5zwAX5IMo5JB2Z2jOuE1PYSd3dlfcukC05EV3lRxEt5IbjM0Mz0iQNa8IWqJfvVUmP5N9D7X
PHPRiTVdk5bcao9LjSA6Iq+X7ga2PFO2a3BeZg4lqCIy7/Wu1sxF/5kMsgkQjB1iljJj2B3zrqkD
/yBeCN4ymz1sPSjU2Big94kQe/WucF6upfyTZzaMZKaaOACA/v0UHp7Mj6Dy8B4F24hxDCLy33iU
BOX8ASkvGt0OclrpC+fnT2XrKtJaUPH2ZayNHX55O+C1h1aAzPAk12P5HJXGtml0SoaQuyYaz9A9
9z90z8bRrw1Ouk4PbxxQfB38I1FOAFYJiImc+bYiuXvyeTEMm1M2PgYz0Cct9OOF/j2WGUudQmg6
9DRzttPRy1e85FtLgwuiavZAl62LqVBTXAkCMlfetWrXV3ojo9nA9bby4QkKAp38BT5cyBXftKoV
ZCwNjfDrwiT3B0sbk1revKNmdJgl5Fp2xqgJCMeoKws+9rH7bJ8JP+oWg03H8WO3nGoKnPRGK9SS
lavt5JV6Gh/1l50V/+rRjuIe7yJnG5JmtV38h+x8FsMSTSgM30r1nvAvubjyWS2jYEid785+FXny
n4dN+tqSqmgjPBwDuGtBmld44gJi4BZs9YakUFAwpwqQNeubkLcyY851AYkFSypDDyxav1ywKXLZ
y6FzbEA7Piqt988e0yS5rTxUxTQ8WEgOpbx5NbnuI+FAji9kcgWgrs9D7W+0Vg2SzGR4YNGmtFEg
Z9ih7y5I4hKpN2rIbkx0jbgmrFN1EDeOWfdc2PhTHND/rF6c9AoDLJqpI4T3IsLrFU9baUIdcYyl
4pAR9VCU1QXuI/ewdDbdV5zScOthhMKs6LGShQ434a9sZ4syX7g1lN2Qv8+0eATgHS1/ceHCmq9p
YdCIgZiEWhDrIBY3YTQaG37prCCSJSDT70pWfuwgHV9wYuL9TaetKtXPSepSeCgxMRMHic/eW6QQ
F1sD3RoUZwYD/5rzUiEE5g4oSQV8zIPh1BCPrArj/DQhOZrAvo+ATAzv3LJxXPR47fmce5rUbD2n
z4SNj+h9sIJtDzFv7T964OrDfWCMktqPEaPQJKWVtectCzwbTG3TsvMQ2bsH94dMtNT3pJVWjQDc
6hXTGkQ9R+xEFxB4qkaAyo77+OMNyIAYs+wcywDpARoBXNv1/M9LOwzPMGwf3v9KK4ohOptEJ9zx
GTCgcvIpGmXPCYSZpWEMx1UYNYGj6IS9jlOH+NWWRMtnl8BG/N+AVBqaAxr+tLhe03dFqCLHJAIp
d6qYLGeJThLGX/emF5aYl1wIF6Yqq7i4RZd7qFESumUMfoSCcR4g9FOuOV+llo9x4mHAWxIeHJ7i
EbW04t2JMxhbCK9Q0ISZhsreS0HtDs9GgtKk3fePrSvl9eQul+f57GyTzhoNh3ikUnrV1qiYx7GP
xEd/r/IjiFpWHTD81t85T1MEpnNX73GRGNIwyuIYinWGNYgx5zrSOvQEZEYinGvqzDq/jzS6HBu/
yGiGgH9bCEDkLTAEHiWk1HMfk/m2pH5HI13jpAAJtVaTdS7hP9RvGOoUmWk/JU6VR21lJOG4KMkI
qS9g7+luwFmkYDf0ah56IeALb79xv34zbAjHdbt3OMNzUnaK7yPSJdESjmwtm7CfatysKLGMF+i9
p4vOrNGpXSF1ze1mJlKkQxfkXePu7UgpG0QbIEfvn2gaef/EswQUsan1EaDSzvwGjTN8yEJZvx8f
xUiHYOfY0xJr1RJc5cJRxgi1hnk1Uhcru77N0EQa6k2fYO692DKobVISPDJkWbhcyPqqyJr6ZMhw
/i7P1ncSDor7vKbbgVLNMp2I8eQdh39ojXXWXok/zEX5vlPCazp9hJoiNJFqIJhlPFfbP2tLIJSB
+EURBfvo3lp4LfBN+hnWcbePxu0SHKEAFUWRTgKlOoYnMnU95j9pont0JVA2/Y2aeLbCMmdzOqXN
X7TfObDXbW4qJJb78CxXVCUHSSZJULnv40bhMpIlplFO69YeXLh8noAueFp5w3sEoZnH3rtQLAHy
t9ISjU7HaZSl0Ls68iS0f8gvzObVZ8Q2D2yEqYOZCAZSRqX9ZFf8LAS0F9Qu9WKBZxml1IWHBefO
RcfKmVp+sx4hxhEJqp2VwoJph2V/iZJtnL/wQ+uwuNuEU2j+yVGZHPipkfH2GIS+9XTZ7j2Y/ruN
MEj6apqqnQzjGSjumKtWfjFO8ILmtYMsUAJviPwEsVJUw4b78QfHQfB3PtANJ3M85XEbLBGN9MJc
Or1HvNxHMr2wKq/EDwNFzFUsowF1v3/w9Acj+oIJVcO8DXJNze6xXxFz9BF/pjqfnxQB4KDIvcej
Oi84QeCn2SXsa1zy0YqSYqHu0aNuG1Qo4FHVNSucnbvDz+1og+GoOPZvNt4j/V0RWm9/4ZsVLQU1
qHVivH6/N+ZgeEPoQhbk9mz5lP7J0DCBtchM41pf/sdcnVYUv53dtiVeNIhXye2LtncPKdw4/zDd
2l74V9A6oICCxKfepZHEca2z7d1r7eTF2/LqZgxDO2BJy8kjWiNRY3mBkcLK5QWq2AzlCVafVU2D
yLmVay5B5ZZau7gvPbbZlleZXZgRazmMd6SzFAoTBBq2pPGukLewYpFMZd5vyb/FiDl9Srjrc4Ac
qRauW9jv+YHuKvlVr0NZYx2AHmkczPmxztrKJ7PdJgW2bTqMudr7nPLyZqDLfeyF/GulFZuVXZlx
J6RXMr9ch8DzOg6nXaZWmq3IaDBtOG55F4o6+4OwXE1b766SburGv5lOxo58f063o2GoXcVooIcn
zhJRpD0G26XyaPoBP2M7yOoDtyUlysaNfNnBwgf6/SsPR7Qtpu/BpuNrZYHU9jbl8zn6w77p7jP0
GeO5FC3mtMTsurvpdfpJ9xWL8BPPlusvKUPZbzUrq6UWuRVZ3fksP2v+zVMAwNk8CYUu7429Dwbq
Iq3wcQOZtlnLNwQ7wCZK8EbuxsdvYKkm1fsNQdRxE3I0S3nBiEsbP8/reXS6Ciwa3cLpZ5l7xA4X
IiRvf1uuCceIP/PMunFW2XsDakkJSOpHdJDD+t1VlM8u14kv067flcgN/fPhjBZWlvyrFvWSOPTZ
LmT+WTSAgV2ioCokhNXPzoFlzYev8s7QtVNwA8OWYVS+KS7IzG1sNEMqaKdxBShVhcjfdg6itD3R
FmYye9PwTOSXOmXzE6CwgiNjYw9NgGEVCaSKWL7PR2f00pWMrHpieG1fMuyRpeW4Apzl7LEzMRVb
Dr+oB2/FwFEN8k280xYlc4hl/ztXrt904r6Fe0p8gYfmIPn+pGSaV6x2DTSdmctCf2smzlV2+HI/
yHb7/bofnFPCB/JVcVNptCzoEJrTR3ni/5HJZCmPFVPt/VWlizhnZqosuRa3Z86iHTyhjkeGWdgz
qe2/clHQWm/pMzXwny8TyP4HilUR/pQJpce6Qy+MzJWb3Cynh+/hKHztWy7lCFB2oS9Pwsbyk2rp
GqF+UbFfu3rP0+yaTMZUIAd0ukcyfyH8oJNotuRh1dKrYTbYip2otEelXYGZyPfWCXWSAK0t1gG7
iql0ifdiUXPUqfIzQ6DSyX7JNpAWCrs2XB19+ZBwXqr2bOjmrlvxW5q9MdqyvHB3T9mcshtCfX1o
dhW0WFdk4Bkbim5z5h7Wv95fogxK0IzFNLdxu24wn1+cr7gru5kp7AuYqeepVxuM6VEsbrJ2FLnX
ALL38GLniGmj0R0scqxwgQwmFl+Fc0Vul90z1K2Ri9DLqDH8XwPB7b7twwSF9Uu/NMVxLFkG3ZX7
bExVowHkh0IeWV9I+fWHoEuA8wr6OFTyTqo7U33un0l48VxLsmz7Cw09aMgwlGmSM8h+7GK4edd7
TwKeAGR0i0HDvp7BVoeZd/mE1keMTD8XEXpbx3NXJcpMY1KNUYN9/rtFBvh4W395sc21Ny3nSn62
585douRwBcyoHEpXWjuhcL7iOBfPC9RvkxJH5kF0wDdENMkmrQOTlx3NUNy3O5qvSn387YatSyh/
2swBN4+QM/yukja7RmNAhpV6x9vVc2vCgHXnm0GsejxtpsHn2fcFpwbBh4PLTU8cjs/eHFOVKsSN
MDHEwJ930PdPrMRtOks5sCIKmq1aUGqLowm5pDOQ5eqo2xC1Wr8bE+Zy52z4Ap1KGg3AqpmfJyuF
zPLPxCgri8DG6iPml5vdpVO111tVR8ta9Z1UBvPvCvtg+hY9YDwesV0PVIVwlm62ObOFN6y1adwu
nUtNvDKzeV/pdPb1WLt3LW2Cri3RZrJwHYyoaJkDkvrlThwGQQcXEyzLRBCfWYfCEyLCyTSeOPVd
CcqJEZ0/7hV72Ljr5rY8aaRcEzy9iroNFbE7mBScF0xW9BbdV42lRJfS62pHex58psBdHPva1Gjn
0bxOiy90cddKkDYo2PUGo/UyN+a07ER+bFmfdTn6EQbPx32bvNWMIs9mdoErxx/606kuQzobIYUx
I5nhIY1wseimzXPvUHlZGK5YGsPf9jz07ePUjyfwR0B4VSXPT2/XNGY8jlO4rHBcdC7m5eCv6KNB
+jNG6W1osQc3dBrqdxLiMvc3/QXAeiqekzxbgTmKON1pDRWma+08T55syy7wtuYYW0pSDic9Llbg
nmqL7mSOUOgCM/mYUQ3ojQZpuLQOTBcd1bxaBD71MA0Xbn7eykx5NiF6Uqpf0Kdy1L/PVkY5dBS0
iqC1ZkDYSebr6EYD3YK7Rf67emaRZWizbk/dmPW5K2x2UpozkEjmNxDHkbt9GxulcF0iBu4R4u5R
gdjP2xcQ+fR6qHt8l7ztimlgfVTuYomtQBmkMVntUvgf6D2xh1LbVZyWripM0nXeOyfYDaGC1K0V
oouQy+Mdz7kjyRKQnBk1eEecJgU3bZI5PKQHXDRfeWtsHEhrgrG5LArvpzNVSPOiFiz1zHRvL6+f
7Iyr6DJukHG9fmoWMzJTGkui/uS8+2mNgj9zSfrPf0LP5+EtuvDEUN678IV87n4TWBVN0TCy7gBB
OWYM+NKx9Go8ktSeK/O/UT1VT35gCOw6vf0RTAJDY5cLGJxyuoFa1u/RdJot6w51PvHhKHmZRehW
MXLH4tW3bsQb5ooq8bHaMNXbLDMq7a/HPVAfgaj9MIAnegze2qI4C1XCRqeXWBDhQoCMmZ81HsQ5
lfZiQj2/dd+D+FcmzrmHlLz61iNQAVLIQL0lp/W9sbG2XLihT5snbt3ZjYd4B9WH4Cqj/ufk1qdV
PA+dpiRtjcSDgpGjPsxodBMq2m6KAfsTDiEOEojlxx5IZjlfGkB6dlOJkDw2RwOH7NFzRJn/WDGr
GFMeYXDwATZmSsOIO8Cy6yTa8nPQaEAo6sW0GZjxxNZfCfZcB8uFhxoKFJwhK8PpkzIqhh+IG7+E
JemWCBNCCYP4Qg6Z0kQHAUgQPAc9smDek0YujI1p9kDwplHidff61qmjybPyYeycrhHd5+tfX9bJ
jkJA0j8YEJAxdGkVsqlnjLuf11+i5oqsXw1LSbikfNgpMY0JdyuNWuXQgYH4CsPjAR0INlfXX8zx
etdKRcXV+YDM+bF+2mW2cCVn9fD26BGbTsgrr5qnH6xmd2n6+hrmRqXZNBYj95Qc36Kt8SDdhHGg
zj5HdIwHrkX00q3LQq2YFj6wUuuq7Z676c48GiyeNQzxspNekEcWSGdUfGI3X/IS9W7X2jAfuD3H
dR352Da9F9wx0A1WKwhtpVxTFBQX8ynR0ZOlDdzWh+jokCtNxsgogRQxtyZdotlt9Ut4XTTjbEUT
XAYmU9HuBgtYH/JyYdFMqZEPnDyO4pVeNldPZwuOTjQIAFsZ9W4Gfw3+pM2U8egKRVFDAwEYxOdk
F3aYa/hRx/oQ2ghTREfHao5Qn2oHmf4CGtls63Z9uARGqO4WvS55HVRc7FrgXDerKtsVeMEjRI26
95vhKF36BWA8XphrJunAMThBwttQsfTurgFm1Se/4HoSmrR5HE7eNVN2IIaqHlGr5c/l+0o+3WI2
oZrcuIdWjz2qrnz6VXtUT44DFmMhedbfnrgtgnUJvZuPuMJv+yhc4E9MfEyBRR75SMd5qyIdfIFS
JE0ldaGJ8K3IypvmGS6J8whKy9AtWLuTpytfLh7ItzurBB529mENZjm1JiRvL66wbYZjHKtAf02g
Z2BsgZ6ljyMXU807EIWH+55g4/M2sw4xxYvG8BVPLXb7AkgyvtuGW/xH401EJYl5xZjWkDkLdQIV
fqWArZxoylUhjUR79pcVoiafIXdBIExbV8WltrWB3lxoALBXQTkK1YaSCAgrblN4PyZQaBRAPTTD
YDtM2IP0YAEF0Rd/3yCsD2BEPrVKVlxKYtUnPaF2beQQcoSNBnuMHXrUy11Qrx+dX4g3oqOcJCVE
txCcLPUraXXUEdRmwU3/GU562spL9Hhn48fQ9cXhycFmNIrnqgFrouOkSxCFVqNDwJz5jxDfbgkP
B4quehLxXSpFUf9OHPPiYxBsgiFLYd5OysR/IVInYw5RmK5UeuezVJ8Ujb54wqXE+QGTSEvh3O78
gxjM9O/m6mdMjVuKPcYeeE7p2KIOxVvlYilrHbDzhlWC/z+mi6Ok7UVrkiGh5TFd/KaU3htnMdLP
evu20CffXXZAbTpQ3gBWIsqXr9cmIPVb0v+F3p/ipbhQmjRpTznlPWiguLdx0qjx7jf/gYpaTi4n
PuABe7peVgonWheNsz2ZU5Cb1qQWCOQk3/OHVb472zdYXj7lxrQ0beM2oazYiQWTQNWYRtmx4AC8
PZ2DanDr1LozkjEARoRDku9x2pJlmS0/VK31QZH7NsiUkWsnTLIA+9Nd8xH0yOquFPhTMJn2nmIp
EywenYuYSF320sfPqedxoPS4vRSdpFwhK//EuXpv4S4ChXaRRSKcDnRYjYhqRwpnb2VOpbxgVZI5
mhYlUar81cgGeYFRNc56xHsJYwydnezD7jKcnizOPwIdZOYGV1vJcl55Ksx9RASuSfaiJsZnu9ca
IT7VRaZhnJnuzZSFW3F9/5z2LFFDObDRj13L8XqDU20LkvsCZdWKqbHAfRtO5ue61u8JPRZ2M3ao
lUfmrjOlWOl4zx0ttfaQJAgX2ke9bOXmg2JuGDzDoNu7g+NAwC1SEITfP7yE04m9tjlzYqYuASSE
YBOibEjNZk/F2bVFH+2KHv8ZaPAKdKTKNR0KXo7u/y1Gu174zxaY45fVdX5gSg5/fry+gy4UYIA3
DKot6h7wPlsJD3OeSI8BTls5L3c+oQsup5bIegSBZALlvsTbI3v2LgLgZulsuqoY2teXiOKIy3oq
FNsn4FjuU8nMRbVSqsElZ/T9V8hoSjgZ2s+muu/eTFvNKFQOO0PDOf7e6ocR995/8MWH1Xu3qgf8
QsMMwijKDzUAfm7em5Nv9z713X+T0Ru3iA74yVSZ2iEeygWqmFihs8najVqA4nbrACdhI+oeBdeT
rrjVOPi5TV0IbV2y7zu0tLcILrSTgTtdcD06upHXrvYHBj9oh65U7cY6gBXBhD6DQs1dW9B4Vox8
EsloQXAhRm5NPe1ScKKZqb2Fb018i6Bi38ADWvSLIznEbHnhxZyOgygq0Uzpa4RePWn8OSckv8yn
cNbc3/1zpXN7FqhmRLbyi017PmsAyGKIGuyYM+4qsFMznUUndYauCvd4YCdwL6Hg6x9Nc1pHSZF7
Du0b3qDOn8LLmCFLQOvLaXTWTM8XhC8+SPX7G2HN6NysWq7L1woYbdP3vYyQ7FW8MTMK628yOLFW
+07yF5FujQUVpAMjNhIUBgx75lWNjpBiCaWqyzqQCE9rZM8dTL2uEY+hLZiZvsWfamKp7eFqSqoz
sCUPcpKV56ioHSSH5a3Lr9PG8TQZXrfrjVz+/dM4NBVeFfkVsI55hJsDk89V6LU5nO+0ccVkE51N
7D7uoCxNd7GW/QM92FbIQmLcVG4mHHrQtf8wQYWv1QeZPfNleWlUuvEdQVmCoeCwi69RCby/0Se3
0YYWQdpwfHKaJBXvpgZh/UIC5JN+SS1dnHyJZzxdTfiWjMMUX0xkH7hNCR26Y7QxTgqKPJjtKOdN
IopPoS3HUh8/8XAFi1BOB2Yz2ZWxZxNNhdKMyUmmBlhc69a8Ao2qIoO1F4TmHFI4hmNvVq+FyuaU
cmmD+EXOma5q9Hmk9JPEdrdhQk2s5cYOnpeDON2t/I+SYry8iBVuWTm9JRh4KJcBTC+7k0GxJikx
xtn7UnavQ+o+qzdzmrnOCs5rV6x68PNFQ+X5OOqicMaS3ll1q/PTdmIqd9UETRyExRDKdFJd1pim
PcpyaaL+kkVi1sc1+5lUGdKiq1q4RlSkmAXS0YRlaaM4vtTfavxBb4BoCsjtDrGS6pxJiExwCG7u
J5wx8t4vw5G5cgWpq2TDGfKCQ8Z71+obc+ebkwbbnfMSz2f1bVbkFiRM16zUWf61rf6WOQ0fI/mX
v0gjjnfD6gG8l9QoQsOQZcTXPjmLz/XKrcCTTan4l6Zn8Jh2ZDuIRYux6nHklx/e2lc3fkCIarIM
c8JkSjPECcZC3ihwDREmba+C6S4Gv8hHN33ggrqsRwWU87QJu0sbQuhdwpnDOnIppDmXS4igMSXU
WY4pvuVa3OgbWsCBdqV92eUg1EWiNSO5C2zN97+bkrr7+miiuBzbNHh5dZvF5ogxH3znQuKx/ei0
/nQtiSaD+GjM1Stzquf1MXxFKldeHUEgu817kjiMadEmLO/73addwn5HtCLmmKIv45Fr55tWYbUF
BDh3MQ4pwsgAg6FK7U8YX6qHXGo/tlkRrVg0d0HMhb/o0+8c38CprMKgQi1K/nxoexHtg3B/ffUQ
5giX2uCcnwMsQBl561Lsgw+z9v1tuFbCNiSpTcmlvdYb58HNQw/UAIo5IoamhMDKwB3hKGhFYeKn
hohcnL/SuVeNt3JuBqOgl/k2JveUXW7Ij9ZJis5wn2cOLiONBDluYjXqxtmPWWy0qvJEw6Kqy2sf
P0igznm2PY8VyYpurnknipSf4ZGQLVV7PNbM0TQxGUmo4N37eGiAhjpsns9dSbyibhjeXHauH+Bt
F2w24H0LQ2S+qJwgBEb6J16PuiBIIqbJEOiAnhavStuakrbEkydttf1EJVNmc4N3jzgcW4jeiNp2
+vn7A0qqr1FEa5LWrguxT2fBraZq0VXU9bPMiQwxXXS/QSmKje2wxumnB2KiL69zw/T9R3kq+DG6
jWljIh/3VMPmFIB8KEgSk+4i8W0XPbrHT17Y+Wu2t7++I4tOBxjUeH681ipiNK4sqnSE5tBGxTtN
OwCR8LPDhs6U89S7QPsPt+/XE02rKCgtZxSqE7RUvvXJ7tX/U+Uw/ehu7pNgGEvUAAMpdMwh62nS
DnBDI1v+Jut1+IGWzmxFMUcXBycX/GZ3y7vPnltD7TA5HDn5/b6nwOvdV8/7JxWimUHMTfEdpwe5
Qo6y/5oZ4GVEt5gueXd3DMgBdAI1k2itaSQF8hPBP9ftZoTSmgLpJHJ89Gj4f4X+apiExX6SHLMB
H1R1UNWbqgmh6Z7dMp+HO9BiaaxE7CJLIQ0Hz7ZCIItybyD6IKS/2/uxQGzFTTRNrYr+a14yaWMG
a9NUCVPkM/3Hdc1Ory8LlaXID2zpNH8omWXr0CrSnDQYlNfKWxWHh4NFmoTMkXP9Am/Qsu6vHFLa
9jo9Mn1k0CALN7O6qvWs7yd1Vaya3mpx8Wl33YyZowDmG+qj1dS7BSb6GfLCwPAo6Q2ePz1Q8RVX
b6ADzWLuSOilB8DIMRFxlZETRM2zpd3T0Auv+UAL5pRxuRsZb4WYynlrE6DLUc8jc01VbNIYOIgC
EHcMMR3ispVKfl2ne7APKKnvA6lotWLOBLTij3UCk4waT+6NONaBfKVyR8eud0mVugjk3uZz3HHT
CtslNdcLXL7vZgHnuTc00bUZVT8iWNMlCeJxEHjuoSSDSihzgUln5FECXbDBp5uemo4S5/nv4f0t
lx5svp11fl36ddtW2oJ9+q3hYZ6UyEob3E4PcI7D/RtF+Zlylh8Gk/a4CFzILMnbzQrACV99YaAF
whUhbEpGKR0OPmki0ZzRqGSNFmDAKePv5WR3V0HqDieDGYWZ/lxV5qmdzhe4smEeFLlORBXVPHNb
lF30sHkcTBtP77l0+7+dQaEsiOAX9pZZoDKZF6mB56gnzSh7KRYaE2HqZkeczVK+00rY017M5PgU
eCjR0TPYJpasqjtXtNjBm5eW4mKAdAKo/FM8XbFGyLfKYeJBb6xLT6dDQaX2zlxmlx3SvTCFL7v/
zPu67G2JlKL5VXuCH0SMYhgXv+THPvbROJorYybJy/SPAd0Xh89WgotVc38jkCDGcA53j2dr8TdP
QHfnXlNlziz/p5KwoRG593JC7wmm4fVQLu8GMjhMF5B/HJGanPGNLpOBJ369TN7rz7Jjz4tL0UHA
yTZCrPJjYXEUHd+X7cVmZc3shwhL+YkZbOJ28jXRp1vBLIK/F49xd5dQEgZHPShKlcGG6hgIPi/E
VuM7g6dAO20yQ9pkQ7cNzZ3rhkI7y6Rk+i1JRj5/7j6Vdvq6lef8UKT1HgEM6NcyQFdZ1HKaro8B
sxzYDOx/qBZSK9arEU0a1vLYmcfHgTWtwvMlzF3quC5nFlkEGTIHyAh8xPm2fhtxgKm/qkdL2xO1
r778ZVtsxEfppQEonByoK5O3ThrqhUrHp2pBa7ON14gUQKAKajoRI1EX7H0h9ecMMbNbVnq6xT9l
QlxB7Vcu3oHk63pJlrYauVfGzisoYJf92w4mexa5TexETQc8ZCYVBtp00R+LXudLIk/HnzS23sep
ExJXXNK/wpaRHeWvugTdz7yV4/1puyd6XrrmCPIoE+Pn8/y3tJmvl7xfmVgHiR/682O/wc+ZASyX
djJOVWbyFZv3MGsCORteV0d4mydTFC2oJU2c6guBq0L4Hm+wqdMYYm42lmqMG8CSZNgd//R3JfB+
tU+Gv76BQzBVpusDdbL7AtbIGJmOt4IN9T9WZoK6cKgFTNJYpVvUndrZ7nTq41rT1RtvGLRQmwoO
RO2xDWw1a9Gt0aNUpQk40Jj0JrTajiAavCkhZJCF1NMH/9VHpDQ171xY/3/YnLi7a4Kb0/520x+s
0n3RkgojfsOwz3M5lBbOaCr2Y+8JziBG38Hr5sPhpAvp2N6y9487A814hFR6TkV/5TQ0BCVNA02S
w0sVYkd9LxoPxMwGz+hFcUy937N86g3gFv8p2FGVHb6BTfLy9eThJgehuxdqbAPWqDnw8og1DXpO
FKKnsWeKqD3zDgOhS9fcOqF6/KCOD7NsCejMclNHM9fCibDMKc7eVgxytHYitQmsSe9kueA/QYnN
Uuz8XUYDv4Nj50elEVZ50geEZthb88e1lUFoqqfFmv30W6D+RsuWNHqSXdHo15pqKAo4meRxe/k2
fP/q84ORQaZuWliPvOCgaXOzh0a034c3o1BLVXdCDHLDw69s3xmM2p/fwT0JpLQlMZQWkYEoafCZ
/V1Ltem39HNYbX73XPYFcmUeiww5rASyAsNDihNiP+T+dP1qOaugv6M8lkvxj16m0DQdwTm5hmI5
ITdROuQnkdCbljFUahg+RbcYq1Pc/0eMYHxSojsOYW7ZtBNy0L98WR0SWsXLrpduH9XLRlRM7DKw
NpvMbPHmkTixsrLAquxEJX0mIO+AHB5EkG7yZdRcZ5pjXQLrXO5nwXs+D9DtNvhfCJc84/XLKDqf
XJA5IX930vf5dduJx7wtQFCX3D9CQh+y98eS/wLGQiNLFtJKvoQ5+ZysSMHl6AxsPGYgbFxJGe0p
vxEiL2dywnoHVwFeh28fq1fsePngIsFc8M9WjWSChXy6ORg1iyD47EjlbYKF51aDt8esXLnLf81C
qxHnjVBwnhCHhRIJ7DF9cwYq3QwHwvq3A1CevRkcnP48rXGGJ7CoHR8bLe04gONalYK2QvZTKP7P
YCNqdyKEow+RG9Yy7rpi3MfmKqLC1u9KytmJ/KqUARP1fTH6xeQ8TZhLW8e6rV/CIfBBB8b/da3u
KL/U774830ivxMkoCnDjRX/ABJ9Zfnb/X3mmjE9xXPxtvfCgc33kP/h5U+dEtTxhwJkE9cDdWqs8
klQLhMQd572gX6T0ZU+iey1g/hIiGuy3VMbkOtC3t/a3KUFVyZtSy7BO0fxU21xTUMnN8AwjAMUh
Xj6KWI0ILe+4rJ8uMxfb1Ql4Je0YT8Z8U6amh6NtctmTsQlP2xI+zMRTnYKHJ9MLejV12DIGoKKW
yjHsZazQIo1bIRXl3NWSjqWwHFD498TfrAZHyMegoTD15Y3sYHQloBIdUbP3Fdt7kpvk3cqCOsXE
LsTBvA4IdWSxHaNGnRuL4NsBD5qWkWHbsS6nihPzO3KPqaxF8HdaxiTXN8ZTmfmJA+Q2sOFSGP21
P2O0NGI6z7In6EICVvmW5Y5uL4kYqr6lnIl4e+Y7GOcc803BrL9Q7Qbu0NLBnTpb50IAfsALsXWa
Q4nn8xfmgJdDn3mEH3RvPXm3aaZRMaK7O4XTn82fP2NJpdIJuJlWsuK8r0xdHvVNuEHZ2/czaH6A
gqnby18kvkISKJvOaQHSQqWliVuVsp2atDUuFG+EmE1lTslLg5WltSliE7dTvl1SGbiY+hBCQpN4
tJN505g+pqgM5vgKQ7Fir+yA93Ai5z5sAmnrWAAb1/jEnjn56GQ0dyutvqYb5B6ErHGsgK1/FCJz
Vdvb+nIDuqqWCM1uhfTaf9aKMP08EE3ITL41SSsVlYI6nxbA9ribNfSRxOx4xpRU7/NIY2ZQpYt6
F08WT0WIm9LYrVQ3jkLVNsAKsVy08KjUdUW9XzOIxBV6pj/3YUwsOcnBm7S8Rx7X4U7NP2U0Srmj
PRCqsBfbEiUogbjB7rMYExhJU6oITTjb1vp52t3v4tmyUK6wT11WXSUgO5pjPTDTcizW04+Q95Iz
7wgGlpFv9oH9C6clwz4+l2g9rRvMYhw0CIunCk8iLwrlz0oNCj49CZfZWkFKW1yc26dptPzQAWX1
X7aIGF3VsOIzbfiYh6rxWuTWGlyUfGLKoTa/a38EnpzqAH0FX7XcfbvBgdr11xJnGaJOQmCQ6Ejc
LLzBUjZcgfuFHaYFM+FBgb81gJZVZZ8qR/jQ7Lw8ExkXFTWruS660fMOPQ9+782iY4keMLXqS4/S
9dnKc/UP/tk/aoA1Ki6vEaMQGbowTi357hqbHZvtNvTVE/RlUnbcJQ651coAwd76lTrqKMook6NN
SxOEWUBckH9K8xRNj14FJG9TWqjfm4JKXNgAg7DqW/75eYUi8yKXPpzXMtWNRTE/UK3DEG/tdgao
n0XhrelAEmt1lbjTxFd6Y083ebxfKZj1Pl/hEMp7gdaESeyCArLkA4fjB3vp2Uk4gzNQ0AqwmWYR
FA49gxrgIKzk3NvPRRdSs44nZllXxEO18GHdbCycxbA/vbM5tGFI3YKAn91Nl8oXAhOuQcHVIt+U
CvRFmtG0ouv8O5LWR+37+pBcV2osBAqHTeou76dP+THuBLE8BrS7QSxzbmFtTDZjj1iEM6SMq5E7
rjlGKLo0e3qij2XGb63+W1kLKkC87BZjj582pJRVhBke9tZEQFjSq0i9l1650fgdhxbvSJIty1Rl
MpPpzMrVDdMB7X2hv4E6A5v4gOGRuuruv1ntDSWVHLkE1wZSkR2XXpIHFlubdYq/i+r1/NtBdtfS
Rrw7oWHaoAwi++uOvTpyDtH8UjtLLV0wIIkcG9HMEtwLLmCYkmMhn38ztHmlem+hcWqUW2IArXCE
3Q4CuWV0SenNfV+HkaWxcSjXiUltO31FXRL6OlgkoruqQDlbskgwrauMgWRdVmvcTtkDhMjwVYzh
PGdzQMQOPSF2GpLQyNuTINuJJHlXv9LLgjLLjjyP90hi6rzv5eJhDR3HXhUyMOvdvhOPf7YXRj4j
qf+slKuts4e6uOq6Lt6Lw6O036o00Pq8ZOVC+KBeJ/I+L/AT51hXZj93SomFgxsssxcwYC8ZaTL+
FpOs5ujKVMkxbyhaGOsUVTeWnOg7fIQGb/PmwdiJO5ls6dqQ/6uUm8cTJDS0uheRuNkSmk6rXyFK
pUYT6EV1ScRfXTjg9L3czBIFLzwJbvAgPPfBkJR0Fsd/y6nWaJbSquElNYRQnMxQJ+OTj/MnJKmN
UQL4TET6megM0QG124rfx1SXaittaSl71QyyvF7gzgVuI95a9iM49qGiqk4HAj12rjh7EjHj5ByW
LvU2nAlQi60x6/6MZ+h/KSWd1XxkQ9Sra94UfS9Yu2TUAaep6cXlrqQXIvCV1ptXdxOavDSnM4bO
vKZuUQRAbGbB3QgZd0PeIYLiRtPsI0a83ey/oGp4iiC9E/btWr7K4WVRmnR35gVjL7A+ox6gaXA0
YJiiAjqDHmX7CP6gJoRxWMf+AxPgimALI5+FpEw04GcJ4sOZH4cBb5HwOnTngFEeynEnwNvDQVeu
dn5xMhrH+dT8VtYISMaN1shydA40So9XPynNBEKlnL3nbDqpxyQtTzdAqWzki7WuWEO/ylwP/RYq
jjL6jiwzZoRYVh1AJsfKeDkO1or8xrERte1mOnAUf+XGDzGR0+BHxRlYYTuU+xsFvTwWfN1CJIxV
K2DkzI6gylSNh0jrboEfvr11d3AP1U7JMPT3+nwT9NiSZGeiF1G6+ouPnuYsb3DWrlQFuFdvE/P0
pFSlJmJ7XTpBP1lUVVTCW+3CLbt5MBN/kW9FaXcHnQpB3aIQ7pvz+cKoN9U9gGyazlb2AksbyZg5
MnA4mvDgTbonWzp5wWz09wXO5sUpWLD0AwZCCw1SgP2bXIPDTkfSkjrZYK2Jut5ahzEmVUiXQz0/
RCupeDxvDZ5SZxv5/CzsRCKx097VRb9yzwr+vmUANoW+w/Ffs3L9oEGOo/e2prkj62YNdE44bbbJ
9BkR+yZ7Pi5f8J3nP6bivrXdu3rT8kTCP76xLQ/yHlE6Le1+PpdWJaLdIjRxNx9B82CyMLb5wXpd
A0F40TzrM7ZcjfvytKyjWCwm7AJ617a8X7cHZexhCTGKS7iUuHqZLXb7zkOGMoOsiaGmU8WQpZxo
IkEhLW8Ci0erdG2cZScZeYzotuzPdP61YuJPXc6YB8TL5ku82ShrfdpY9BDsXcETsoQc8aqjbNz5
QYP/1/Ga9voRo16vlHZnfpKGUz1F7X0kypWjl8zR9Y+OP220PWSUznOlWYmc/LUI7gpaf1Rn1B3G
hImUD7NT7b8R6bII5x4Rdj/n5haDIr/Uo5leD4MOMKeqEXTHqPmiBl3HR/nA5R+cn+NXYmCZg6Kd
U5d/pgTkkKdjA0gzMZxcRiYrKvIkTsiFEhDtwx33X9DjHp+jMcsnv93tmkh4W10+mcWY7VEYZmAO
dxbPx5rx2IObAC6H24qy5kIGWO6FUrXdKYUKsaX+jTqQ3Piu5o/aAfXdchPQbmK51M/suPImmy86
sY3o5lEeXFTmLNgN4y6BFLR8EWPUL26C9wlqdRMq0HxSdjZeIgmHkK++9OgitT6gDqokpPDM9I1z
mitTlntDThOBWQGktyp37Bpv9XtPbeAa+YzBA5xTmXnMqH7g7JAnrBznsFPPmUxNM76KqtHmld8U
Qm6WYTeWLo37a/uVsgsLxrdAU9TabfWgaZTnDwfbN4CaQwwHheRxdoXkOD8JijKNByRySnQhjQYx
QwQfdc1p75qeWoQz0qu1PMZ2TXYHjCcdT3tsE9+Mh6lTvRtJ4rxeMUAr9NeAQFRNUuAY4YRkcrX7
oVtE7vzDeOHue4FzvYnFdjWji6IydrB6QLAB4revkqPl6rNRBm1/irAf+ALZBh6Nxq+I51lDujiE
iEFomjB8bJOTxhI2dZ90kxxKQN5XhPQR0oeZEyqT50SAx0DknijRbera23O0bqW9A26+UzjHIIqj
srAT05z/+cmo4cjriKQ+GgDIOmJL5cFI123JAqMTuj23aBK4YuR40a1THl6BpEZJPy2Y2Oq3KH3+
4GH9DXnZOpRC5gaW+lGzhV8It3FjnVsqxFv8t2VB9sGAhxno2ZCJ/PY5llCBxi09IazOwvdEhuwa
bj4pUZpjsMDreYmGyeXitM9VMw30WGh7AqKw35c82WRTibVF9VXyE/fAHVdiwRkMH83um00dAoxy
K6Q85pjP+vGHtu462kXaikWQrgCCQSClA/77f3v9VeUVu/XIH3OEYx4VpOW/kchys0QsqqW1HyM2
DtvqvYN/5OHSllgdO/SZkNZmWXkC/GgM7V2OwmcF2DkgTCcd1LMFv1ttZU0S2HDTT/mizLDkDkHx
cxBkVJow+h5YNMyqbyjBZDZWbhZRBfdkZGfjTFkJm9V8lLZx6UUMvrDJdtLFA8ixykD6yNH/8UGO
+oqpKf9qOZxmZhY22RWSv3mvnBc3/YnKMkZprxmVg+7Nw70PgS5NWHcPsTJLcZFTAr+aavGKHEqh
uFNm7nMBB6Fj1rW1QIM5o/mvmkJttn85OfC92H0+tU81Tbkc1XCMhiFyS2ryVyJX2dbCa2+muD5l
5ostD6XhAwq3ObCLMeJLsI0FdrEfkBLEZExaDV7JLzuZs2HlUMC5TPUxtZTQwgwKwk2u0C/Rvtg3
ryUaQrJnR05tnnjmYEoOE5yr8jHh9N+xDvCkOTNeAUlqmo8e30a+TLddhBeTV66FGY81g+ot2xyh
6+tcJnWoWO0bbQOkAXhP43hF7IebVWW+9NaGNL+oY3OBfKJQ47AXULh9zq0Rit1fcfS00V3bvfHL
OoJkk9I3ar6NCBHBkOLkYvNahavQxfM3588x6K4Q243Ni5mOREIbzMp1i/CxdaJ5SZMg6U/zCG6y
HG5+2RffagMzbnMv709ml5QKdcqDGdNSXYYoG6LcYdqWeMiLhWsJEdbtYZK6lx7wWXsvVcutZRdj
6WoozKXHbmxHH5IRL7i/lNApzMDjMin4BCluUXovoFdTZVCWIT26xg7qXn0oeCD1B7CN06nMYCS8
wT+0q5pbPqDvwW4UxA2Wjy2gkQChgtbyErSTDGQNIqwFOfNRbwo6Fr9wNX7jf40CuoPeBZT1M/Dn
1e8/X4VAiTwG9jKS705C5fS3dchTc2Z1w+tGYTuVVtFbpqtKPTxGBFR2qMCYfzWfl0KUqCZjyycr
nb9TV3W+uIMYW3hZvIlNxxCaZv2zdjDEvuO71DP0rEJ1kBW+hlpSq3Ge4c6eOtlJtgCQ0O2KXgGq
oF+MbD6hMl9426GDl1EMjKmGvrx2DV8xYz7+L7TTia8XvzgWt1ESjY3vJedEkj/b3JiGeTnKIigA
1L5nBVD7aDeJRbLVNwD8mPRwsursICImLNBTPUrHU53rEFFLz6gOGs4OcCcTbiaiefmXNnB951r+
7yyVl9F9/3mvaeTH3CtdCcVaqbJrkEXDbesOw4xMhVGAAWUeIuX22jcSj6pztq5xYUZ+x0L34apE
awGCx4MnsZ/sjYGb3FQTWI1YTGH5hdGxlkOT1OWpNsGfbsYFEwN8n3ayFOrS0BSCsdzeg2W7+vxl
vVxHok4v5R9fNTQ9r2tOAzElSQndT3Lrppun/xGaIDrduBvVMXMZjJyKZdWoBmXv2f+A+m5xZjnX
MMwVWbIuLmaqbHvKJ0yEZEUM5Ob/MM7HKRf4P/ZvbNaRqXQptLXkJdyUIlKQyG0qyRPsCoQoEPdn
YAhY+QseRihIlHX16EkPjFjqNl01DWaNQk3Wa5M1YX/7TDVTzl4PAFI7CAQMRt10RoyHGEGj0eK5
Q59qyax4jiPPxqihdmW5zBEJRfY24VFr/IoOM67ywn8HFeOjrYlExeJLh6K5jVOAb4D3PkfXWNbr
8OQck+z828FnPMZfvXoogXxghgwIBm9/lFwb0yre1xtuy6yskkXaePWAkVyQLGGuQTGNw96i4z9+
VtG00vfzP/fSIC4sZKU1pOYx8nJGqS2h/5uIZNmdMwFKvJy63TDAjocU5xoVbm6tf8nbGcI3hG1k
FV7Ab10xV9t7livq1J/0NtWns/RGuOAvdUVhaGqOvB1qYAgZR1nDLr8/3Qk5+Fmz5QUw7Zrd+/25
1EsEPXcXYjz04hKW1d4IrHCx90iX73o1b17p91IOY81/26go3X3VaC44ukw7D/ND+ybNBrDZepNa
v+tQiphEMd9Szn5D71RUQ5MQPcnlVxeWw+UXjAsjN656k9NqECwbIuh7oknl7JRkNNQUnk1z+o5q
+AND7Bf3lil7oOQPurA6rvvPchCHCnaCcCnIQagd4xpPx+Mb10pw65aYeK7KpnE7p8DapBnlnQZd
e8jF3H65oIkd4X+xvkVOvmi84o2kZk80OdzX5dhrmbUrVqlhasgvvOJsyvTlOExyAZ52SeWt7hXU
/EB5TVnlzJOqgcOyHYdw45fF2hPBSq8uTfx5qXCVfxBr0y+EbazxxeT2I3Kgf9y1MQ1DtAyuyQcj
S3ClOdm2W3e7xZbu4JJ2Qo8FQhm904uFvuJI7poh3z5gspoRJUkzf9bB6+hAu/65IFOV7pNPmSCO
nCMuI3z6cafMXmBQLhekaThkx/+D+Keq1SoDJQW0aL2l9FhE7UysvjbB0JpxP0s6GTKgm3iihN5F
dh6UnuwbrKmhHA+85/06Zd4uthaIxeL//He9Ki0a/TLy2OgRfzDVj+WfWwqCjug8bZLe313YsOZ7
RKm8FbXgSUYnQN3izj6c7rdpdQHVWH8yWM9Ff/smS63FEQnQAX9X7CBjsvN0GJt4t9nqt5UZIJ8W
TTd1shSMv5nHP9UuzDyoqx90YFSxggR10BCHc5B08YYy0d5uO8EMZB4n7loMz1wb18PqNho0RPGT
xStbItqhu/jEPvukVLnJVFRwbrXtPnudC1gG324KKhfEOCwTXvdy2acdh1ymIFATT1hWYZjnJEHj
/4cnAdnQdH8EQuk+Hz9wyOtYNZRNUISkl6ba1I/Bgv67GDfwPgV+32SQ8U17rYTH0X9WgxonmaJf
1ZFpz97LWYzhZcUC3/kT4FUOUXsyCgQlEe93FuVUVuV4nLoxuXNrAvG4PuQoM7hWzenS1EE6e5yJ
ZwpN/MnJomKb/6q0toPgHOKOQUOkX5sYjVP5/ZUw0GW982U7VcawyUQjLl32bt6CBYRydk61fUiX
qKXYrO0FqxjOiS7igLXl5ns7wPaVMasP7lz+WhjsRTK3DHAXoDG1EvhPp0YhMWXvk7FkbCj6GhAL
TKh8UCivOphULkB+jffWGDaxObS3d6dOsk4QMEpuN7Gj74F0tGpl82i5D+ZYwf3nwtLfdXm7Hrrh
I5YpyZTQ+QltJTKdu2ORsSSqP5yVFBRyTOqBV2DxUH5MAzUlZyXPDrbJFkWdnTpldQK9wfDDWb5H
YEXRY/ol3OA9VuuE1w8lv9NoKJ/75q+CLQlAFj+zcuUwG5z+71y7yB9+28/wBwKBYLRvIBQYg9+P
1RjnJdXMHaeZERUxGxHXv4x8aZA1HsIk0NzCA0y21cDB8Js+GyBGYmFX1cAC725la1hdR7eMnW/n
cZvcYNEm/ALp84bvkQblToNHGa8u5qfxKrPunwcKBDeX4cUp+N6L751NLJB0FHjplxyeVJSjG3s8
VgPCY1CtYU8OqAbghfgX0UrG5Q5wpZWj5kg5Lk3uY+M63hlrp8eR+qiqNhMReXu5V10XwQwCCHgx
5pTKElFJ/QFq3/7H1QJl112OJIGsY0xn7QqWnIJIqm5ZvuPGw9AT7mcBwST+RCAEMJhcCBvMqff2
66iIUUglQihJSiwDr4MT57yqxlVqIsIldrII9A6rVXtQmITjMxKvsN8amB6Y0aj2WLepwZKUkDmc
i7VeBkLb1cYlJX20k/SyxPyZK/jAIlwLWrUtzPm3XNxgcPhPlKLKpVlWDzDQfTrAMi5ABQIC08lm
CFTWXaMOX+iObaglE1ExxX5T1qhjrnhfKn9VhEVMG0o7ewXLp990f1Tx9HTHKl9mpH687eEvckiv
+SHLzdc4GsAkY5kB1tOKSM3DzGIbM/LbQLCwb/3XfmvTMw3SIBCWjb876VQ0t2ocyz0kbPi6x1q8
a3iz3thQ4k1HCsTV4+BQ4ZqCSZNJD6TUzO81YVS50fhVR1dKwde1UwW+5HabOhTjGL1JJg06/vvd
J50khTq6UCnPif0+h6bF4WHoCbZA7WR2ekelr3rUjTrpbzQHNn2QVYjIWC8BiJtk0+9T6r3xChjl
MTHihfIJV+czbJJOiSpWVQG78TogSv+K2zVDeTDuNK+kFyfINDwcBGVDHqwRm1G0jph+jE1AYlkJ
wFFGZ9q8mP4K+ymyNLi8UbCacCxmdbl9Uh4CUbpdSnyhEF/WfbpBky/KUy4Qg4udDTe8ft4ZwlYw
q3ivw7v7UcybARlHHW+9ypx9nyhOxBLhr5hF+BVsrcjwNCqu9lrpKqIOx4L7ieX0o/jOepjVPyAZ
cKv21jkWpFyHK48n7WTY7sFDhpJlF6WQ/EyJu2xQKe+jtMfQVnk7TX2eZ/8yNhHSoIY1sDofME8a
ZiDgyiYtmct8jjathM8FOvCDTvIEC9oEKxBw9zjqV/XMfvyr7sGYw7rvh8wOXFrM/k0aTkE4TtzX
V3G9QbGNxNwbLIBt8X6osumCbUN9od6ORj/62zHP8N8CU/MBjX+5EEsxOzgNZG8A3IyXtVVXSH/4
6hoJPMauEOI7lOSeZPcmeATcqofjvh8DxlII2ZCPXty9xNr7qoxOPM0pxqJEq/wn49Ir6njOGvA2
tXbM0IlBHojW6hAu0nzLl30kDoso65Lj+6GX5FnU8w6eLmAtARXly61Mg1bSHJLgkFb3WNopnviR
OfbUo3W9zYlrgR3UfsgefnEQ3Zg7D71uuSfFhShPwokbEtcFVfBbSnRFdmFX4kirWscMq7nW1kw4
RpiBtg7LEzDetO+aR31gqF0n+J8IsotJbVVXiEoSLruNGn4c/eyfogb4AN44LokjA2nP9F0UUSk7
bTR3qq6OkazRqn3wMX9XQKh43/T5Vct02otKFBRCM575kApQa28B8EGhVV1nGNr9aUHMM29XECJF
8SJoi3E0yxD75kPIbMyq4LiFIglXFyy2OOnFvkhqjxcSk3Ld/uQWNZ6rAY+fkou//4UjKtxtEUa0
pDRICqnpWNVeuOfuXKmrEWUfbBI5JUjvh+DQnaAxX812mn7sQEy2mFeCwJs/y6iZH9tqvYZdjiNk
rJ3/SLQPwNzT4WXi38NV/sh60F551hoeVEpf0gkyrGytY5qw9VAOCDWiQquS7NiblGBfaYg3AQ61
lm/a599rdk+YuYBx2gchi3xo4SpK0MuqDR1pDQp6WoivcEbH2nF45yb+htLw23vES5OImY1WIafn
i8zjjmiG6AxiBLcEQzn6ZPqfqZdzjI3akJ0Jo4eriILZP4u611OxeKVOweX5XEKjF8B+gCNfE8eW
68MFTRhqagw2fCPAb+GEOGX7G+PQ8J0ZRFrouZcAzjnDogpsaZV0c0iHP61cKciJIXHNuOMO6Txq
W2hEPpsIzd1/nzt3IjmPcZRKzZdIyoDcWdRZFC9EWy+5t/CYMmOikv4gQEXRt+80wHUg/IRRW6S+
aQ0AosB7QF3cjtBrcRknJb2r5AE+Jmh/foosgWEmXeUoL0TwhtWgRNuP3+yqJ3XU/7iKoF9AEt9v
TnVXFJ7IYT1xyR/ZCPRwklTcnpURoZjAlTGwzMy1o7xkcPwxGYyK+b+1NLj628CXRB0EKl9OIS65
eaPZPP9SCopbin5yTfU/FVhVfMmu2u0doZVp6WJgRNBYR7n20+KTFSih7p937srCketzmAzNGlch
rkscqMmNEJy5Cy0iAfdGwfQ2rEr/y9B6yIMgJU/CMp5iUeC3ASGDjgT+oYQ0kAjkv5i4wslHfGhh
Ua2Q2TXNrEgRA40wREBN8WCZRSDd0qaNZYtSnS9e2BDf2rY8noE7qXOG90Rrkb09SX7reZFtSFlm
qaPvDHZm8xmNVeJ2DyUtBxRjAO3OLrB1kjWU3/UU4KgK3pNQ+k/8B99mYCAzWr+tZVe1wD/X7aR4
XLQZabaEI6vIAEhzfAaaj6WZWXye0QPloGCZYz48RD+mPapCXPFPL81Yzatc+6cznk9VHZ9twxKQ
ZGEw+zzVZgZJX+qRHaEex98MGj5nFBfxpK+jg7J0bCBY6rjhpShbk3S2HH232TUD8hsPoW+Q3PKX
hpMnu5ZStJwlYI2DuJISeKNbCiEh3ULSGgb4jHL+iZmCjcgXoNgBPmM8EUV1rMMaXg1mY8df4grF
dd1grCN49FX7AfB08+0sPEN/7/+Xn2zcS59i6wm05XTFIIkAcHz3cwRTvKVlr69Y1wjPCYy4GYcT
3MZweXpcjw9LXdFU8wj7+aZfc275x8pcCiDbLBiCSenaYa9bNdUjRF8C4BI/WzMoQeWtLoVA0mb8
WCE0a7dPNddmmX1f/euqsVONGb9vEkOHvmlDiCgZMiL+dA3NB/K4j5e78WGCYb9d5AzqTu+fsXso
YFYHHPf4bkRrpgru58P38esozYNoxdMSLbsIeUsRQoREqajK+6ty/ufoDT2IzwT//y642F+eYDst
9rdAhE177zTX0jQCn+Ur5KMqCH5pc4/upkXyy6na7Dkhhle3O/Nh5y7Y88aIUFRhGXInCqfugwgt
YN4G5xE3ZgmBQ2YXwIWwuDmgYA4SJioTtmSCm4SBmXGkEKmHf298FtJCCrb//cCDl0Q9gm8Oifd1
ibLkvQYnuwxAZ3TaWumk/RVTRPkY8Es3fxYoQQjUkYkVNuKjaoeg6GgpUb5tkpdGyh0WOIrdRmoU
wxiDx1Q4YH2gFaqYTshAb5SM+rsCaLJd2fjljrmtOZAq11t3Fr1Rg2Wi/DrtgdhCxLZhOdubmtPH
XPSc4ZNrzUFScJrof63kXvqQ1p/PbFSFIJdPFQneur69xYFjDRaK2EL8U8LpWxsXZyFv23wunzMj
Xl266fbTqmcLVWCiXrMBFJwGy3dOm0W4MJizlF8W6oMU8aJoK1mc0IzqA3WZyAs5xxWQTLKWOr/b
US9MIZWWScEZ1JWi8tF2yrzjT4lExgJjFgitNgpVp7DlE1yfVhaGN/5Nm8tBjq5lIqVZLFfmWGTP
QBmaL9hB9WY0U3+tYyZRzJCa2rULCJpITxs0RZeE6IEtVfWum2oawZZW1Sd+M12ClAn1EzXkklDv
mnXhwlhGkHMqyD0rFAqdvoJVV0yDLZauA3SWlMR2m69xAiUWdGTMNXmbJYfjYk3WDyCNEvU7W3mG
S6dp3b5BYs8YxBoZnRUrDlNhuVcPrBitagXnPmExkaf/9Ndh6GthzMTuA94cROSC9ltcXaHjvA4g
CmSBnO3cUJjndld9SN6M8ly2MPS+eizHo94kizRPHm3+R+ZJoGDM8TuNw9eYSocb+9Y+23RCy81Z
k/oQVCu8aIgsj+5XYxpOwWJd0hTIP+Nb8MY6WkLelmAqrmou/mvw5eXAAbYGeTrPQHwuFoSuSPKS
5L7w72HFxjDwGMznDAJA0yOa0IL/ekmWP6s3LSaiw535qUWaHkTJuKek8vptdRyrP30A8bYSfw8B
x97m1Dp4NAxtWRqlfnprYChbNoxbnwHeraZOm1cl7gu1POrSHbTRWNIMPluMgyiUNKUjagehFO3j
yi+Uc+Y0yjwaIVvmgN74EvsbXP65kdfByuNtQS6JYlKy7XFp4ka6snmkcOapYf3SyOedt8+aNK0E
p0zXB7uuG3zJ1BBU4FEkdE/XFZ1zlk4F3OkH7A+kkepEg7R2TZ1M/oDHuGaAL6tmPwNR/rSV8OzC
CMuwouKX09WrYL3Qbj20RyPf7mcz8i7pP5j63RTmUOuQZ3yQY5sKwioc9dUpSRAIyhke5r0LkhmP
JwzPtPwnjMeeTW+54pQrYrsJ8rf6et8Tf3NHnxTJ1t+rev7PBUiki8+dND1VsoBqyvIpTEDJgrPF
CUiY0FLlol+BnENyK6QJx7CMZyW8jbSbaGiKCU+5ri8uos61LFeiZsSo22eQInWyvySUL3AQeCZr
SKdB56fGsCEX62sAM4HOvpOQrdc/YDZpharqQOddH5NsGv2p6QoCxfhezf06jdF/5t0Ow/GaaRlZ
sZbYUFuyQCq1+xgGsZ5Jq4HGdPu1JyvDfmsQR5tGTQElqfIW24A3Q5KeajVsa/sSVcDa2qZqA5e5
y+F/f3Hwjtt1mHELTheTPMsuSf2THJp1isanNz6Wchjyez5JsC6LgfXJcohXbwDX3m3PhEld+7Hh
dytPtMLSOWF6E/EYOuNQPuRkRGvg+N3uc5cJtaqRkU+QGV0F++4ICQ/EPsuQp4hm8oljpSCqGyjc
DKz2C+t8EujJQg34lWEMDIOtAfN9+eCpU8mrX0cP0inwzY+2HKltRfJ0V46qWrphNpwNzgkq8bVv
uDABh6p1ZEgmH0hzT/Vvye5b5AIm3jeSjkFpkYiQp62Vpqm2dsdwCUDR1L68KMBkJrEkh2WgqygA
rkLL7xPwB8wUTYUgSyUfNASfqUrx1MgW9eF8I5jJxgKumqzdzkSNONi5q7okbwQGiM+mIfhn4mtJ
JH4gHbSEvSM5qnVchzhFJWPf2+/6UfR6WYDMRz67QhUkqIDq2uV0ST0azB/e7q2OsqgaPSea+U7I
MTZHRCYLubeR93ycULiUf3BXxFfNEQiRqlgtkDslozksBGAIH3KkS/dWGKmusKIL5/rr2gDFiZLH
YsBGAetPwjBhq0BEsLloxbWiv4EgA8hBLPFubQnExbQ5MjRFkidPc8Tko5nmOZscYiVVD0lbCnmo
wR4ZArbquFgYjOWCi7la2+BNRggkhRNlbNCb/SpCiIv4MgcwF/igS1z3V7qY/jpOQkpXaVPZ1WXp
ZLEeT8btNLfnH0PEPNLq2jcLi0JSwebS06yMEVfOScD5SJp6h8yHWown2P0PUxZKtbu2xzyGFJLI
KmWxWrs5ZAyFHyD1F34EHnDMjKHwkgePYiUPFNmHnM974BU2h+u2BrJyLqxALCmzCPFjBJdpDGkH
0Ao8invLYSjOYZavb3/CVIsIWjtCONu11RRa9J7M9KIVN+1jWnU/GDTAFxDzogeKA7qW2w7EaOWv
NNmxg3yeBdf5tb13Eqm6e8B6tpvsH/qQosdjgWcxB54pTTMvkthTbrR4NK5ETT9I3rq99/TU1XXr
VvBsTu0i+AN6GOa/ST4hxvbCskVx1wQE9Qj/tSUIL+z4GwsHnB9jd192C/U4M+0y32ij20tS93KS
5SlqVs/m3tdrmM2oiE5joiRFLuV5EcdQcEJ7J62YN6bXR9wYTYONqM7B1JXAECNXu9mNbdI9O4ik
H3OiI7AnmOE83ZSH9LjOjaXB/5bifo7JBgCo8m9hsSuXU5HLwhIJ/s3JE3vz1VPZblGqYgfyYz9h
uLeEmETjZK6GrgfwfqzZ4Dhs65YVpgfDWWUZUrLeuPniXezHrROeLO1x3n6t21kcTOxl+iUPjmHe
iCSMY0Ve+JwzHuCkrR1PKS2bHb7GJ7chLxOzm/foEedjlTwIwol1VVNcA1rpna3jG0q2qljskFXK
2LPC4DIOypw1MeoQN791VBM7CND06rFo53bI6D8BlJc4pNF7Ha1p/CgSeLUzWxBE6ly1aq+QYl+h
17Gfhix8dnh2ztbD95+uJ5J3Bam2xpLCJWPjcj5ks+80/Om6KX+IjFzH1W/YhE5/tWkQcOXr0lFM
zDTBpgvysbgrjU1fEl/JTcDwndYzyR5LNwIai2bIyoQCqeQIGDsUu1u9odYtfsR3ARSlQnzKzliD
BujmsKjI4EfWsg5zAV/zwVpe1zp9wV0S9hFR1A8CgKzBLPneNVW0rRKNw7qc/Jw0W5DvSUwQ0lSp
gqCUlr0y+kXBWcONu6eu5g4ZuMkcskrjBiDeHaVD0cCEnLsZE9cJsi/LpsmfvVWi3giMKu5Nm8ck
YQ3HeHsIKKn0I1mAGHk+8PjxfnlT9HbMx7Iq616oSBkPcsy0thgfcA1/YenqIItIpy4sc/rSyx9H
f7V7etR0QSMq3IUtYOl5CqDv1AaAaHmOsGXjYzsCm8Y5e6w+QJs5nAtL1Abe4wTlv3lpT0D6zHiP
KCQbXcNgzTV29ljjQCKbxwhF2I809gKZs5hzFWEo3vS1K4UEauzOwG8i/bVBUUyD7HrwYUXfNPg0
Uc8+kklNX8F7VWGbErdqVT7e0olbxoGkmbzK//hFTCj5WPN42Kwcl3iLwreiNIBUijCbZzG023V5
6bY1NO9HuZRyrYkZhSgnWVyUZJCeB87vdIOfGR/4fqXeTnOczHR/rBhtT84YRGVAcIrQAJUEcYtM
VECtGilIU429d8BcqHLVc9+XtfqTlEZ185V0Z0YuX55HWMk6vZG1J6C9CkvQaaM0Y3pIRGtPZIXq
153BKf47/fJnuWTgv/d849fx3R2VEMM4Llbt1ZXEZfD4G2QTArsh6xqgZu+CdxfzUapk9mRfJCDq
cKFYBVwdR2A1A+dvyfl/Q+NLDMyb0FBR9HG1BehoXeujHmWlKOldhwCFtvIhAE/UFzZv8sfzv8KS
gVFS4jT8xvjCp6YOdnbGLmY5UdPIBLvzdfbVwBdau1pu5jA/6gKHStYrEdIWmjVKLidtDUE0x6fb
bZqmCVcJaMhsL/6G1saM+qfZYKS8yI0NO3fRoZNZhcb6V+JQyd/oG3C1Ap9RK8irny6dH/kXRJts
WXMGB39pp1KW4in7yaeNiXK//y7pUOZr3hVDF8H5B+dC+8V036GIZ0EITtp0i5ltyhCZlDPX3Xlh
Fgj0uBevEgw5epu7BGcjxMhVVgbJ2a5RZ8s0YFi68vFRJK4BaB1/zac4BIHKl+8EHaBITSuLBCiO
c/Yar4S3ZnxTpA4H8fep75jxpQZtSuk8u+w8eV/vxKiGBddrKjaVP2BIFe6/hY478wu5OPh0weFx
SPfTwjzFBVcDn3dgBAOAuA9utPuI0Bm7f4GhELejXOdaQavbN4aKfv9zOK1vYIIVUf3M5qgJeBHA
XC7vblS9ecy3xdlM0Z5KMvI/kZUYt7iJjxCPhYaaLyvISUYPZyiZ+2483mfkeiAOYZjFOYZo8Obl
VlwD0Qx/Rl4yhoxg8XTNUQ4zKTXoZ5dd4ZR4XTXaH/e39O+Y3EobevFD5+/4mj8GlqOu+9hkpvHv
Wm6YDWvfj4gXc+4IEe655/UWMWe8+5cB+pQk9rI1Cy2lLFW9X7nqr7kqrwsvs+ioIaFpLnFNs7l1
ILaHRyAsgqGYBhMTGl0V2evJTPSEbNYODvwcMtUjEuE0RZ0PbNTyRVvyx0Z7XTipVWgovJ8irA3+
w9C5s0d+ziwwwBLKQnp5DzEXaUXCfCdbpPfgnr0y/QDP952CsQmVG+z8kD+GORMsqPAeuc+RK3Xz
1lYcKg72BcKdbPcF+8uIO1eeeehDp6BfzOOh9nGpJmtDSo4zXufkK17p7juyLInvzgX6TjVQ3blK
kKSfOmSCHjLKJ9LTAlnT1ondvBdD7IgGD9HSRdWCaIIz0qn+NS2bHIuljfnhSJ4kvdRjTLlbIDO1
VT/LprgqEKxEweSecDP4wsYVM+MCSh//gi4HjybjPZjGlfaeyPT+UtACWkErVHKAPPcqNcnOA98+
u27TLHt9wSjCW6ZVPGO9gqFabEu0+MQxnOix6bi3XIP+SY5ZaDaVPjAwhb48v2WcON8N5tLF+Fhk
gm2zHlEpHhkonrg5XQvOze/hhiJWfVzgUWVEMOFcO7sN6pDbuehKYuABhr3AAtSX6ZAMDDrsdMWH
+yIZypnigMVak4KfuYW8yh24tFilRR/nnXqnOU+2sgQ08cfZT4aDMEmUT5tHVBgiBMTLSoJVAzmi
zOyWwnbSxVP3dldLslMe6rx/l1UEJk2JN2U+ephWNC32OPCId1IfBspxXGCdKITCq1xQrYDIu3gN
dHkPECZwWpsMoCKqKs8k7/YeLWxYyqKaojto1RuPg5GhT57YRu8DjwXGUWDwP3B9M9IB6eOCZnkh
YuvwOrwa8hRTmjDzO+eotUCU1cv5Ya4Awh8DcNIueRONrAJJXfdSd6YblRK1Ci/JijONunygQWJE
7VbswzXbWakQGk1Eg/Uy2BuAlCgpaS6V1Hpy+K0THtLQWNSbdXWXHtTZi1k26u0VS++kyCFmx52a
J+JVs2jzgZM7DtMV2eF9UTmY4cIV6GLburpo8byGbps3hRMtN1pBrmH8wGGI5SH19qePMEUEuKws
Ins1+ufDGpKT2VD1FW35W/9scxM7pVaKPMd/hwuXViewiGSGUSHZJpGYG5GZMVI9cZT/XxH0bSKv
9klibyBqF6ZCicz36YPxgoo2IL+ctctDCInXUUTMarlLbdLh06jt31i7wyatkSStJeqVpOOm/BUz
Osr4ouPHHk4y+02NmQ1T1iTi7yLa2tdCwKgxxwp6ztGWJQRSRCaVHVPMvkwRdINUPjO6W7OXtiAE
P86swtAVVL4rqZvPOipoIPVTzK1jXRjkzN/IjH+XVfsyWeSuzgUqo1qLRw4CQ+qNh3LjLKfQjh9E
HkzMl85PaNrAVtzgOYzvgGRy8Bmyns0Haa762IQS+j2M4Oq1W84SgGYyWNgymM0Poo3hXvZEVNXw
UhXlzolZtZ7nh/MNNPeolM9ZOH0NUznb+hcaJfiSg9shtcKgDviDlERFyWGW7oL4n3g8wOFqqbQR
hg2QHX2Az4Hhh1o9YpP0yC4A1jQb8W21Z3AIurrKBUjr/85LJMX6nIlxgsskBCPAQNW8QGuWKYy+
ykemVoV5GgU0KxGyntTrX/4jmUY0C+6uv7F6jEQCpI4katKCvqPxR5Oq9hBijpj4E6451igR49Io
VfFiztZZnrRaPUyWQRe6HSnrdlte1zK4VqdJx4unXYfIrEtHiZ/3l7NWlxMu5u787+1Pz8a02llW
Jcd9vjU538AvoIXTfkw2kYjQ8INtdj/vLC60cyWvV7JqvQvH6obxKmnlP1iEC2aCMlc8gPAI8aHy
jZ87SoBVFz+iqRWgBVfBa0ChXELapnH4udsZKIqpAgoAqgBfaLFp80nsa8cf37013JWSe0kpWLpI
pNuckz/7gExQtg/3sSRi/zRmdd0JrT4O1fXzzUnx9jHDy6RP66EFcIimvU0h+TQ/JGv7Lf8V9E6s
F/IK37ckK3ZxcVNxwJWbQGJ0G1Axj94VExp+htlFndH+iRR5nTMIOddKCP6MT/ws7RpniDUQ5xN4
tRny/sQWRYl9+YEFaINVjnYMmkzbUkDjXxPr+VJh6he+jAdnq2NnAHLxVLBT6zRtXw1j3QCuOVTV
GSUSP6vkxhdtShRiqiXsHjTaKAi37RyrHe+H4Axz0c2ud+8iuHEULM8fkDNwK1bEqD+ojH26wJ/S
fkulK3hZWrNg5wxd2BY53WrK0zmuQvdsAs0yOfH82zBMeM2o42HqKQQ5X2QOBVTEmd7NXairjCzl
TDsizyI6Jbq4yplgN64yXqyo+Wx+O5cRdJre8PZHVKYaHy0CnXD57Rc2s5F4Y6v8gObKoq9gsTtx
x8rXHkcWSLzAEfnRTtWJYpAge0aZ0PXbKbRH7qsuQ5wbATHWRBd/+HIjb7jl+K1jJ13lblp0ayHQ
MXirepo8vLIEKwWW3SGeHqFsJgzm2vGgvammMnIupcYGIoERmNnt0tWzshrfcqQBe+Y7HWiGqFDN
7Oax6Ul5s1ebALg6W1N793kfAL1/p/ZyUErkwyq2ZjfcrRyGrAFPiJMAUG30tab/T/ZXoNVKGvbR
HVOJwPpbB0dtzNC/HBdKpl2F68gU8dhU5iNcJA6Ks607mV+6JXqn+ZJMbYzuMa3jECfwFnl8TPoY
n1r9jVMFcI7qHCpHrYCIQrBwczMUg8wzn2a/U+t7kzoFEfmkkwiKHaU+SDBkzTJV4497F54HQSH3
F/5oTjJDfCjb72Nuz4rmguubfJPKwYeA7ra3gctXO2qNIzUNG8HcVimGzgy9p9dduox6x13qkOMr
5e+KXuO1Yt2hOBia0r1v9LT9RUHVbSYq0yR5/c9Vnq6rcnTgTicR2fZN5KormklOx711YWGmC83z
+X6Czzgy/KsmgyPRsPOcPjB4EE1t6VWg+8gIRPoRj2eMdwZKm6bezm986v+KiYdLJw998ScQVyoi
RXh6es6+vfL7NfYZcYT/otv5zbXuq5pInU9jn1kqLPk0JQZhIvLjsGLhAm3RavUO8n/NF2AIAyVE
9UjdUi11UWL0nqMiMyZLnuAraNzhbuO0Hrm8FinuvpMcQRJjPnT92QR/iKei8el2VpUz4XHDsWGx
PjfLhiWy/ISIyvYYsyx9amojxoQjmdCX48hvOevLqx2UO0qN9FJR7vf7SGEG9trwkX/3C2ztlbwr
LjCVsFSvD96zwKPREPXl9FWpurgr2OhcN3hdyM593a865GNQInA3ReYvp30tSsC3dtcOx2FB0Nnk
ddDtk7+ekVd3VgEbWwh8NdRy1Dkjw43a1KrWdSrWK4sP8rwcIIXVjgjcrIGFTPLpSUT0+MeQIlsb
5Ejmr1C2dIIfRZ9tGgzL6Y3d81aKnyaFkVOB6E7kaLKn2bwuVrN9Hz9530cYHFJWq6wJm7RmzPjL
hspdY55YhtvtqKTetDTIo2CqhT1P3yVxoQJy/EoCuETc1CiQiLRHlOdSji3b0s7KgVcA0v7dhQ/H
vrQtFDzN9tI2XEv8gUJCIw0V9chSpR8mzsDwXBAAXVP0WPeiRfdiZoYRu9jmKPGcHDjH5skkBuhB
mbXnBe1RT/bqdiQw/XfMOHyEEeC8cGwvJPWQXI6H2/vTrDG7PwlH4FNmC8mrAJzIZMJ72iKb70fs
Ch1tOU5MGjhISIp/N1CZiAleI8ro91OG9T2WUXbhAPRQg6KDgTkXCMEFNqr7FvAZLQGMZHmE3WTW
tLJtEfflRWwpiQ3ky9dJVElmfuA15x07lu6IsfjcX5aD+lz9bdoFdPVWq7+vNSiRMScLNpPNGTY7
6TLyyKJSZA2GRX6smrXU1Lzq1kGkDsNcbhs2y88lG1sCyft9jBKcj4H0tKY1kZ//Nnl91izClz4I
G5Ccu+kb4Sy+tcygLPgoNFQEkGtPkLgTQ6VDGix+S1vk2Du3fvFDvokHZIlbiw65esNF5phzGtya
JBtKRroX56aS7DlpdeRr8UXxT6/EC1W8AN/PBsRo9b4gRZ5b0ok4shV/jEOU6pdiWoky52dulwV7
txOg8Krd4c3hs5zmCPBqhbhO/EHclSZjwxjWBq6j53UEFQ82riQVbL4oFghoGSueUcxpQm1RfUjc
NBKXbjBONzSh5XM4ZIIx4iJwmkjPXKWVG8w0c++7EQsxiJbzFJckB7bX9Qh0wL281EgQku6I5/sF
OuLUcqSGFs3yFwkLbrYNS9VnOl3BpP/Ic/X3Zo0+kf1erkSr1BxKFnh5b81m9flIgRN943hbh5h7
rEjrISycLhxFWGVxz+AHAxdjM+v2Sb3CRJutbA+gOPYirQy/yVb1GtZuk7PT5gdwigaR0R0aERUC
jm5l4SUIo2i7JZAQlMcsdGTztGdpa13AHHoV0R3zJqZvO3ZXK5ewkxSpXv9DAlyksUD9PDFP8znl
uX4hFVdd4ViJuBzvaikJnD+WeyRDj5FNuqiv2yTdBQ7bbE5loX+dKs0bPHWMn2bUhfOkjBEKhnaJ
OsyvOzkDcwbZ/hcYTiBEmbBCG2ZPSTpnp7ssOaP1eh3qJt0iRFyqX71RKcRLmQQlyhX/1Ve0dQZi
GFnznsDZUFb/ciCf4RIUWPY2/V+YNCsNg2mgCa2Ej/BOKqEC1KZrZPLQxeR3QP8K9XLGBa4L+Efm
58ul9yXX9JRBInsZY/mt5yDbGirV94oyCRly4ui70bX7WrbVYqgz5NqYzeBLdQh98SNd4DadnpnG
GjSwRMq0fVR1mrJuGjOUuRJuty+2Un1zXBrvhbQPvG4KT9/XwAAzcodgyaj7KddLUf2zDvXiecCR
uN/x4Wujd9z1QYyFTdUIHthF7ITNIDhIDXbbHurIaEhVA3zOO5MBJsVAPjUkJkj9sRsoiUH/8JOb
bNM96T9EtS2WXwDGCJJ26HdOhiEzcSw62KYJ3VKFDrKzT05Poz+nOOn+fCN26ZhEd8RoGPLrqsJG
56sNXOgkgkOUtpcrgFjP7fDIvwNxp0ToW6UOwrjee2Yu6UaNTE4V4xHM77nNJCIsBWEU5wkO1WvC
KLXq9LF+hN07AC208KAEA+o9PztoayW16w0FRbA+OlrHMN1VdKmucL9hVtI3rwAvPGJ7Ro+Po+8e
mHmztXiNRhD15Pkb2pcyFd5iOQ08Aw1tW/X78mgOc73SWexEp2kD6tX2HSB9PFGix+meZgVcLsJx
fijgNQCfS3g0uIJOfOU+7eVYRHa5eZJDxAXiUehXx3r+z81FWvvQGcpIsFJTdnTxitr+CUiCCuUO
1IHK1m/f/TZVHugpGli0mFViSgPhgvgvZJhwdabxxGEX5MS2qtTtMLwFR1DpTovEdCVJiPfDMuv2
emMeKpLJDR/gQcU8xP5W9IaCcel0eoRzEPQIkEiqWBhZb07o53RApJLtSFMbkVTrwRGeGvca8gN2
iMjHhFNSoi+zTjv/XK+6RP7gJBisu6OC3+Mm4bX14uUZwvYV75V0wjjDf9wgRAQrr/uBwFyeGTzE
OfQcQXeERSr+UF4NmfdrA2sAWCXRC//cU07Pm7DLAFZubl/ueBsGEdLN/6SWiVOjWChVJk3PGWW/
nCrzuYNkU+RoJI1Q05EAIu7K7wphTUNTq3XvyzB35XYwBNkIdE2qWysrDf94RkBFkolo5DgvvH4o
O6N83H8ORFljldb4tcZdcwV3a3Qg8Y9lyxI5YzbfqM/uyyFalccCftWZiEXbkp+IhaTJHDyVq5S3
Z7V1QIA2HmqSUo9HnCwFMgiMwS3PAMjv//iy8Io7SH5iO7CsUa8l8/Z/jc7VS/kzHTQ1JlNJjqvJ
K6CRCF38ZR0TjkZd2NHgguohjyr7sfrC3G2T1eMYfbqY7M+EdbyBPm/1N8GhMamtYwnnZUqEaE/w
pMCjqlNO6lWqNYj8VzV0+moldxeHhi7qHcIFGn1ZvGxX9hab42dz/Dc7A/Qq7xmiom7nsCpSfLfX
U2TdURT0WbcEi/PEjxqWLYC0T8AIV1U9Fw9eb317Iq+WeqdVsWa/b5cQ9V1r04dEFmbvKUDaHczs
3xEIcLIGjd2bHhLUkWeJDd11NrsG3leMJP2edjSZIEbjstHiTQN5J6tdtLBm+YuSZEXja8Vimct3
X1JorEA4yYmqfA+I9h+jS8H/vube7bNlw9/cxS0rZtA/Is2scTp/PgJAd7mHm8og7routEU3D1Sp
U+rycK259hcuzuAVddhZ8S0/HtPU/K3MdhAsvLlOaAcjlMRr4EghbMDcmAF7PKP6+HfEGcVf2dIQ
NCtkMDn1CcxPsypHWuvhJ5VUhaH+c5hP7nYAzUVVNEEY3AwPuIr/Ll5Wze5gwTDu8rNT6K3S7gT5
h+v9Sh5Ljv32UYFp54vhXDuDiL0a8L931xbQk4Wy0Gimyn2sXvYgPt9kzpP9I/acRcLswPxxjcwj
h8OUyf8Q7z9e4JZb2v3XHd1ao2ItKe5zxaNfnYRpgKWFhqgKtiaZ/I+aPDERBLJMo5U5rgjNHQYV
ptIZLEC8xiGKp5GwWUOCgQvx3r2US8oYgqiHLvUm8Y7UbG/BXcI7Sz+KaXpkfv+TLk43XOZTo0Nz
0Y4G3ukkaUmnxTHfoIAiaiB3ZHWVgEKwbaHtQGr1Q3Ik7zPz3vKferLi8atrIFDKHfcsmk5qkjfa
PRspKFrAFUk53xqfSmLspwmI7L1N4HYMaApYI5HeNl9jPcQlHn1Igb67THS1dHL0EGkVy3MzecFP
WFKvyyJR1MI/jRNngMeRGlhz4tlyS5W0Zb/jdU6oEGE2Re0BmHuXw9Ux4VjCuGovRCTbKUJcdPAM
XkSrHA99NneEjlt/ZopYEuHN/TjR49XpWNtUS5vWUa3ASU2SfD++GorS+1APi61kyr3uoszV+48i
FW3o8muYXz8HEpqX7t3xN+eeXHP4eB3oPTmWQd+Yyta5YkX1JjA0AowQfobLb/UgX7X0CEBQsh0Y
aCRUwI1Xf7/ieWxKWldLBfis8VyCWsXSGBaFm4QneXDNVB30pZ0A2Jn2Xj9rc+liDSZcUZZNkUzz
cfMGQuQPqGUMjzkKg0VHuRKXt5vDJfJblDyKiVl1aHNbfLzkI82bGGNwU80cT7i36FcposOX3Saa
GHGlv5bh4unZkzHd8Sn2YUIdk8eDfnbxqcZztmcBUjFcab+wLMbkTnxy1nMocLhViFnBWueL+YAY
i7P7bB91xDUSv44eJeaAPaCs8259qh3/bl0myexJ52HsIEPm9u9PZZtaUF9ISQ/8Ga898wRatgBl
jcEdaahefg95Vvzuf4wIUNqCCp3RDeHxz0MGpKkaBNZKhPu0INptDgippuU/KJysZ8tZBL/Sf58C
jWSXGjmrUa2H3x8v4WH+r73gXYekPYalX7E71u2pv34W9mQyBE4hqZQH36aefI8+ySug77pDSQB7
jj1wvXAsGJzKMyi/zijASjr0L5lE8iGjFuER7/pUBzqlvDYjQVnCyJCK9mT6RJPBQkPkjLRXXGYY
Uq1qTI+JwLgc2ZHT8jOv57PaSRMeANIpIbmxQIDzDRFb92GSkCu7H8RGlPUT1in+f/A1lLICxPEN
bYYQJRkquOw0pkyI+/Sw6/F6cumWFbUUaFofhcm73I3pmTnVDbh+216zDR50I0As3AJp96fZdoc3
1rpuu8nlHA57BwJi65Oqt0kvMrZn+QT3EHZRj+/dr8jXFc3aFnTs6HeSLqRPYpxgbmWdTamcheQj
4Xyn+RQgNnyWETE8nS6BHeuFuLVSAwTkQ80dTbeCAhLiAqnd5SGnA+CMIGGm7Ivp0p2d24SC79C7
2yxMdN0/dduZ8GwvOibgaiG2Hr6+WPZu7XpVn8OnLDkxiafOy9ZL6en/MeZp3sCn3Lnv6TmPs0Op
5qzBdHOFgFYv08XbhbQ1xbNUO0WX8dpfssaaJatuW6CfeAMZOrETyui+KmqFNKUxDxfypV5x83bf
D97WEPw12P/4IiypafKoJpgqVf1bejo5qKXpSTwKVu7pi89M3tY2CwergQhmZxZH2qmCODZ5i5rr
RRwqDgwf3A0gMutdeyAxZPRS1c/r71MMcJ0uGXaQtIq0UiE3E4jIl1czO3LNyAPGmSnTYGfuD9qy
1E+joIcwjVVCDnvaY0afzwv0qPbqe9815YGEfz48xVrlyHx3R8rQ7viv2PldA7d0b44rRxmpzPXC
sIXN4FnRV6gpr9uLb3tSKwqCTmlRlt6mH9zN7LbxwtrcblqXtAmGFja2v017EglxXi4dnT8Jkluq
XXkE8IpqYJ/Gxa3xuG3x34E0hPTjP7ByRKHNhZg+M7dhXi05/ogfzE99iWB93c+yMo0jI0cvDOZD
fbVJvqE98f5qn2R/CH/Ka9QL42fvYPuqM7JMrLPlZ6C+13xu5Ca6iIL5EPP+1vbCpstwqDILrmeD
iBF89RW+sJJ8BvSxqcFXVR0IExjWQRbd4DRI4c0fWqOw1nH0Fp/99Uqv7p0G7nCLyZeXGTX5BbY4
YO64y5cRexr1g5SdMzW5y2dxDr9aw69WQXOh9+oIdTLKSXZL4Hw0T2L6PV6HZNyH7Qn9m7O3kZWo
7dyTMk974b47Om0xID053dfcu1BTQ7F3YhkT/KpibfGXI8gS0pwAGY0vtbS4+qD6yI3pOBgnGwY1
Fey9F/cPR/BRCt/vxdzkAfMD27PZr+w21CP6z0jyHRfwVHwlMOWS1gTmtvpiRL+hC+so0RVNvTZE
O/dtM1+qxU5Ydt8xu2Xomy7UBuk4STqhgWHBWtRX1Pe+a6OyGLQ6jNU4oQO4y26zDZGea9YAeIFW
d+sRUqkiDQpeggTsZv2hA5cIXIoAbWTz6dGXUQHO4SV8nrpQ+5+xX7OChwsoNmZQH971DiI35Pka
M+VBkKVkyX2/PI0GDfwgrkiMqYuJMmwDJ/A+oXfBZJ1bDytfUvCqpeS1D3piRq6ho8WRbrM412Kr
XDxWgZi5WjLi5+u07sMDq83YuZhvgiN/dU+xbesUXUcUA1ze3OJkH8NckRH0wBGrILDuYJxTmUss
JA2VZyUfZ7G4wfgmuxhuGoyG3raeoVx+IUQTT863FP1UBePlDfT2kho+9Vir/A4EeWh0w6y7n2D8
hb5vZUpH2FxZCG80KhfELquEq5s/ikt8w3i4bT94BffQGYYayH8djK3+vG9viiYix4DjEr2Rx4wt
QFLD4nt+90LE2JTyWCv9baKi96NNu8tTz8V2msuIWTAfG1kBGaVy2Aw7WOQvvMmS7xkuTyVcOmS3
A6GeZgW3SPbHDgTjw+SrXepmlAO4dGtqw5lJvU+xYk0i81oD66VSZ5gBBlMQe/ku99g7q4RFgN02
CtbDQPMD/sghfyFSidVTUfqxVFpfxNixNj0Bs04Jpjqq8D7PxSTxAXboO1wkmG3yf2gAT9ILPq1d
0j4dX3Txvq+MX4zMRgnkNHrAf8BdFodoMXxIa+RX3Me0TgfOEM52aFiBK8PZoc1M5W50t0e6Cq2U
6lFoiLzi2463iLS+OdiFplL2WYnPcr8fapR/35HURAQrITwfSu/FrM1B4U5tWnsTIPjEI42e9qVu
GfdRipfyyoZKSuAzR0dKdUYL8nem2wOeARiTZf5qsgUPPtFXtaDo4kzq7NzKvoJhrxRbnXkU2mnS
4OKb59G+wCzxWw/Ol+Htr0jSzShqR8fzfEdeOi3Ezim8i3ozV4gANc5+7kKb2pTJRjf+DRz6kYFN
49m06dvg9GUUBUqcpQz9S2OuvgGLhrzniUoxa1/Y8dQ6qRAnrQaNDFSQ1YEmRPJNJZaoyqY29Gse
PdoRTVPZ7kN6bMtDn5iYSI+X/YPcS2rbCUrhp6HBuivQRQNEtc4+UO5B4wE0fiRrlEtFzTP2ycUa
e9lbtM4lb+5qQpgd4BL2U8xIYH/2UqiFy4XfXnyreZRD1O/2MAUua4ouIqo50emBlDZWpiCW6SWe
CY8uOliGdUN4XLqAV7mdp5EHM2C4oACdixXZuWqQS0pbUwr6HNwM8wERmsvZ2GiJnPOoq21cLcOW
PR7zwwWtTER2rNDfdGcbSbrowBFyqWMX8UVR2zErRRkK45k4SdZHizzBBktIdXywFdTVBpcT788B
/a0i5mlpBCADDsCIVVM6sqBvgN/wYo39nMJpYZXsgmgSnvK1qtryVJ7wInvPKa/vCGot9LAe/B3P
HOQSQeSkaxBpzlukJ305n5mK11SbkBe8xGbKaKqTGGaAxjJlHtaFL28is9C5Ebc+mY2vQu3V7JG6
hpZri2V1qvOjCJ1Ahf2MtuSeYEAMArRriOrZoA4uthbj0WekX7H1KjjYvGxMsFQM9RIyolY+q11D
I1qSKqfnXQk4WPlEij9fhXs546KPPJrN0Y0FW4hu/KWi5f9j3JfJRydqOMVS6TdBLc+fkicKsPoR
D3646rzvdEyR28Z0n+w74TurtAqKL3pWDXiu6zogqM+mPP5ZApZxfAqesrqeJ44lGA293vjU5Cya
dAdvMMsXqawbIp7GvakRt9rLOSl4eu9iCERf/qG3YJlM+cj7mVOhA72MTRQahMSLy/8xpEaCAnDC
+lGjM9ku3uickGuUImVBwC1T0iBdUmi4opR7o86Dq1aC8NKUoNIgH9QYXQeg1pbhZJl1AWznFMPv
JmyStBmcpjwTZ/e/SPHHw23z7Q+sYG4LJ3GuaXGkh8/qWBAfoee0ljkrBK4l2zAvlYiCEWSm4JCJ
3VH2LexkJX+FQUMCUWZcAcSnefTVmHoEqiQdsBvh1acfpXjsDtdq8KDeEaYOHHX/h5K1jhEfabtO
GDRpQamR9Cto3wVCwLqVxMFd3M/80grfAtXFglHA8jejFhhByznm46skuehELZKCH/+AtKcUmJsz
xZa1T03qmCFh0fW10jgqoD9Y+n06Yda/3XObudeFogbVvkj41UC2iDqcl4c3QWo/FZEvzlLt4iEU
VKxJZpv1Je9hePE47Ggy6hf4Hdk830lNK/68JP6VOnsC/aEf04KcDCpg7TeDlP10Ql+YnZdsJ4G/
36HninD/xIFxE8suFVahxeGtWlxuakF0xvVVt+QpiE/Dq8Ez3I1lWzu9icZRX3y0Yk4wrjbiXUuz
MA4X/FOc5KBsGU6h764hOM5jdVrPt2phoWeirba8EUmU/atEFO2CWzYpLf2Jw5G6KN/e6gOXis8a
8F6IzLN7CCvPFVv0CXslWcJlCfuWzjN5D7Dq9Zxn7FDIYOi5wl8H+61crxDIudFW7UVWKEJORpMX
pNSmk0LyjN4ngMGI9+DtWLkQJcXCxtG+uOAAzdpUs8DXgUln7GdtlOspR5FSISsoU7lASOEOBzaC
LLm5brvVGflOLbNVy1rZVRGHOiSrYQWh1aN3cXWkVM0aZF2HsrAX7qNBHz3wSGsCgOdlVH6XD4xe
6wvPjUbsXSszPwbuEaNF633D6CkPHQFUIqT+zC7iHSedoXaxUiZVPYflPaYHCWbLzTPWch8lqmw/
lWb9p1VIEmlPkatH1/fdUl4oWwr+XeAEpbn5dcAGABxvtniKoqIjdzbMzTXyL62QbV+OpIGqDbn5
qrbjFY65oFH+/tWcqKVysb6xitwLwaWBiu9eOeY5Fi7xng8RVuSp2mkoV4sqq8cdXxQ9XcyoEcS5
Lipn8lLh4fv4gCp7uaEIwnoGDI8421UN+aMeSzOPoZpO1o2BlAwhSLoudixe6rWGgmoGn5Wue9UH
+T1//858gW3Uz72H2pDYGQI3jAokXIQGHIb2r2jkxJ4gyANd9+SNf3mLeZr2SfsT3FQs6Wymff7A
czCXCWoB1nXbwNcE4h820ZPquH2kzY73dYDZM0Bjxl1qCQ4dsNMfVxwCCmHOY1I3N8tFSCIpG7ZA
S7Tm/wDpL5GckJ9MVCW56n4tHpx6Q/0MjFx2vCTIbVPz20gsvYG07L/hMlzC4H1xakyUXNDBwe5M
asBUG2plltVUgPEqtbJvw6wm8Z4GYyJDDTmhOIZlJP/RHTWQmsOrKRWoiIcaTeUlscFUuZxy/8YU
6+SAvLZuISYpc54rqzFy+n8qanr0Q0g5JFJNvv9egHTT8CwnqQtlXdSzGAmbF6olvJ1Ec8ubOiyB
GlnIWyYb95fGkKz3WbqjqOCtrUe+xSulKcWeFNPpoIvI0mjexG3NCTUoWsjRpUUKgqD6rmXvJyft
1cT2cnXE6ys59NZrm/tDxHaHNdcOgLVwMHR6TDDIXM5PybbtrTi56sHqp08F6Kmus2jVyxHEMIRS
Oc089+Po2HkWtiMeI5xgB9COd4Sq9npJIB14Kw/l3SVBHTwnvJYXahKaVRJ5vTlX4rAgO5aznQ19
fOhP7oSEjVAv5ED4mbCf7JYFq/54ZNl5o/+w7ULBKfROOY2x6EeATLrCowsbbHT0T4ORf7nanTwg
hZnTMmJTM4GLlGFxHrzJYdybSAYJrGWWN7fxwG8XN+k07e3TtDUEthPoQYPTWfi+C71zFfDXl8Ub
Hu1XfHmo4EUxOlMzqDjO3hfEZjB8snMI+bsZN8Bpwmjrr8Yre6P3tQ3QWK7opBM0+8OZp2GhbDh8
EhaMBCkPT3dXP1ClWkFWuVncpCnGlEd3ohYnpRuuSNoHumHTa2K6Fkux3I+NLw3ETFWC3gScTSV6
vkKKfOSsTePjaZeihrRAcIDynoPHQsXZ/KoF8WPkHGsVOqfB1knE5TlnVT6RtOodb7cx/SC07TA0
GYR6gO3RSTqbeBDed1+EwANDtijDwWSNiBnxHC5VCFvpTW3oxZ+J9Snee5FMGr9sogRAumbwKWcS
r9NDZMjRmBQHAJ0y8L8eFkOUTDfuTi1m92rO474lc63MPeZ8ewtkO/Yc24vqn+INmzDz2XeaX6ZZ
L6gkyG/EAbiApkBMiTD77QyapK1XYF82vzz7t+cQuzgoJoCOHCUXkYgw6yqWquhcEM9cw9YOn20Q
LWh+69qW3yaeAfvr7cU9pJhQzU4o8wDSNo9A/h1p+5W8ECW+Lb5zBw8gSP++7Smp1K/QIpSgioi0
NOmRtRMhCRE2jO1lvibCQYUumfXl5/U0/CtPzvJFX77S2SHBGeE+qf5IYY34INu6D2q2lq6fppf0
qmW4lXSZPQ6Oo9yb6h1Wz4RuLf8PWlNxYpYX1f60XLn/BK4HvvNjDbdPsJoj43se5+lWAIG/v7R/
yj3Rjr9vmJTUP3zLMKI9jxGBBlzKCGHENs1QUWMwwVj4K/NYgDFgviIqA0YLczpfnPFUkJ/6cz2o
/BK5qKoAZMXYk0U+ZNpbVJRbTBSQo8gnaQsmryC05936M3WoSqqtvhGOgKvTRo5vihgu55wpTwBv
RpwPiS8eVx4qPCXPNyZ+PuOcUeBEaQJYUGSO6XMIl6MyxcUuU6RmYSiRquJYfTRVYaR/zhkzqKdS
r+nBAxJybefksyQHqraiuPMm4xjF4juHzOmZRRfKqqK3kfg4lbk7sTd2or7yhTryx+OOAacdC3st
kmdI6WTCbxnZS7COp4gju1yijB84jdAafLwMqrUpguXxSBqX5wbOfoLiGOeTeWlFNa9VLQfBVWpd
QK3kgeqNUR1DJIS0XWilkFtiUS9asuBHZ6qu3nfjyYs2E9SOGx8cx0/gl/bUBBYLGBkL1w8XCLdn
bTirIrd2FECtxRPN02pxd1ZQPqq2+eJb5maAqxFTc+8Ff3lmpq6Vf3U1/RECsspHy4LZtV38YCi7
xY1OpZc9ZmSPsj7bpRCMDwJHhTvU2Mh1ki8AFi4x71kZjAQchZRwuGhVPBbQm44DNO7FU8bffErA
kyNDqlAPCXTgqz16cDydbnZsENwAMTy3JEOTy0SvajemBrv0gG6KaalNse06LDZAcobTmmCTsV7C
CsPsaCAHN8wyJxexxmuN7geVYmy53kbbLWXdUur2kLbsDupNTMVOZw1pEJliTMtFMchiYRpXGHUA
etTSJTWxluyNwHJPzFAxWUlDSY2v70qYkWfuvG5wvd4zMDGDVIUlettLph2ySqqmD9dHYGfEYUDI
ukvBFaNVs5TWwlkpVRC7XzpK3eOrjTVQKE6Bp5TXfxdb0FkEs8EramBQDMxPzSfEr1G6reNZGxvn
lBYcLCwhBIwp8biE9ZDyd+AKy6noAca3VR8QPxh+QTP0N6xu4fy1OsxqU6bLLS1mSX27lbns649E
FwZGOHuXiCNNL6Xeufli5i+LsuWhQPUxSAfaIY/MYgFYCYjJgPwjwiXCClul8NzuBcsjl9H7EICC
DMu7qZ3r615ro+hqCDt3Lb/3v1UbPkNwbM3liosjDdxj63cVOI3jkAeHIg8n7IYaa2brGw6iGwss
JM4tP4THS36cVan13Aj607N6JI7PIlq5c5su3eKotAIaufQSeQ2BRM6Bd/jhRnQDtyD2yCrmxcyQ
wshTPy2+ZhBBlhy6u5mJMPnJd8JE7pM7Jqz0GLufZW+DhLnDTOfEqVTf4hpu2/LFj6NT+twrG3W9
dYQBR/BnLMADp7WtLMI2Lw8M0chw05LSpnqq62iVS77jKYlbAWsNSfnZgzsfGNHzYl/2gCX+21t/
EvmmWrJnOcaVGOOfbDI4nsdImcovvJOMXR5FG3CjfA3vgRhHjT21Lj8yC3SA8K/VeVnWAw8rxeJC
j2DgUkVbIihBpnUvsuRqYQ2KDBWy4VziNpPcpC4KnDnbvBaNTa3H6IIKYf3TUQ7kf2o4HPSVcWnW
+vQbp+pIhN7Iin8KoC9zVggTCp1udiPeg8blatStFvi8eRE2k+GuZ0cYGYUIz8OoyDt7sob/GKDI
YCsP5LwE3PjbZSzh5dHRfuN6YkqQ4D2a3hZzZtWPD5jTJZKKnDJBiqDX0EL7SrB3Pl7Yj2KcyIlR
EOYBhwN6+ATTCE/WPcbB9ER5MNfg2Exenfqn/ii0fmLao/FZr1batXiDSypojZQE1ppi5nV4jMHR
Usab2OCk+feVKuUnKkPsSI81c9BOnJzp3eAMnbE60kQMEDk041N/HClgkl9abOHBj6AkA4ac7bpb
4UwYiDvfj2SeJsPDPEUEhqHMdwCk12nBmqvR5yp6UQkauxLdwiXoOt6l5ER+m3z8q51omUQmKRGD
yGqhIji+tNkFKvQZjWmzm4/FAXheUcGzfNL9Gt7m/TNnxBXvtxBjNcyUDsH4T/Uc6C9OwIb3/vMW
VisyGq53otsM24EEuqnHL84lmhiHnqpLXbxHwPvLpHdereiZfLppqLpLv+zML08/T11s9m1SYqgy
8CMpjWhNXi1L333fbll6BwOcVEBi0S8VTN0EalN9ArVcVT045X20qGgoEr0FX++DtpRTHVQqhGOm
bmCoTQsrOfOEkQm4CAWxeI0sr4Is6fOqDWP+HF4sUES97sTRB++jgKcqevsDKCqD3J13gjFcds5k
nDDKoe0FDjJx8aHuhpyZpNfZlg812i6kHGVKoptUs3q/tPs8puC7yJwR3NmxakR8EOfO3fkfYd2x
nu8nGLYkcCI6mWM5VxjmKo9/yDSiG3bJ7fW3/xFdH5JSd3PKJqPXNf2wg4qvknGjT5grU6DTuho6
I77KkVnzX9Fo5u2Jz73MSgNpzMgy4KJC+V5cko5N53y/sjWpRiAxaqDc8Gd33QUtfvxTZKiBY0Mx
7O9/MkN17FcTG8uOpHvweqkxIAnrnmuABpaOB5ZiHQ6IjwUtQDMahLO+v0qt+XFqvQIl/kzsRfks
HQ9ugVYRrWFGKdt9zbxx+sK5WbMw9AyVK3JAieKQLA5HgIDMQrLpS334j3pejL0NPyYBpKiQNtSF
ioXFSFpGFqGtNP8V46s+ut9brfVK8Yq33FM4gF0wFC6/xw7IKHQ8UB8uRtYSyXIq2ZST9w/1gGLg
EEDBA3TPSs82xduvnHTqY+YcBM6yfuOF8GupuQfmzqFx4SHay4yd4v4zeGlizDKAPHFS4fvjKVnM
7uaw5QvSUQrsq1flu+Iht7f8qKQqvTOpeoqkoIWEfIAYKKHcogP1IgFVsGCiSJC6bSbGbCuPgMws
k72H+mUbmCNNARp7yMO2jmzeXMjB04xF3Sr8OJvYhHS01t6tLEbvWJXjyiDJrA3GiImjjUBcV1l+
0EejO7E2s0Cnnl4E9LEIYUu5EgOXCUYWxIrRIzoV4SizdX01sSGYlxmtRejfVprqMvDVuXkyRfkt
HU2X9GR35bhCZfCIEtaKKCvQQ2et4zQy/6ydfiJIcyVZu7Hnm5jt5AX2/cRUytosQAG3OG0IJBXZ
nF+i/A51wBdALwSTL0bGLKtV34BaEpS+0QRLP9R/yTocJIGI7pfBBzfqOmVy9IKiRbwEF6SoIFJg
08lUJpwdpU1nECFWubwk3QudDqL62VORIIfrvcdAGo+4PiwKbvc3+BxKNetNDKmCbYdm2LxfmXsN
TYZSWyGEcck4s6QVtWRpJdxSEdczEPlsbpD4g6l9BDleK6Lr1loYb+AH7sa9dYu+LMjCIwfbx7nM
3SPyDVbyjCGfmoNUsMFQibkEilPSLrSdsH8xVx43HApfcYNTadbiKOgGRZPab+K3Gk3fBoLTCSrb
BCT8qwDXsaFHxOboWZGH/tP2gviP15eCK9ya7hTKhbDA1R4ImZa7FynuZe151PPnb7wtey6RSO2T
RYz50Jmfv4T67XhjtylOmUTM7JM577hhMy69/5hi7obRwCy0Id3VFgH4tUUi8NlgTwtYBEpmX/1N
mW12TV/axuxwKdL3Olwu2Sr0BBgS8HF5aRGgD68iXogWD+TG10yJjaKSRaLlQY7bFISgJCyXsvqo
uIivOcxtF4OzRcNJbwW8Tg7nt/9mMlhsFkObWveAkGIH6oQIuffE352BBoh/ZzDvt0dJGhfa8pWL
nNNWUI5wzLuHLTUxGbnH6AVyfDahvQk5XBTz2Kgu45SRix501mB1pegJ6dTE/OVvFjlwyHpPEQpx
pIAbDYMS7UvrHyLWcaLpK1iJI0NvjWvS9T1mZAvIJQU+oTS6S4OIBQnhfUCllMkYzlo+eIiEyuCa
un0/WqqfUUpw3ocf0JpeKMi4ABp3ODK82nzlZ7KaH0vmIdM0nGZcecC+tTpJ0OfL9nJ4ieo8EfIL
CvYLxac9inaHxvfU9JeMNicxGFecQvqkkhQEq/LIyZjPchpbdKzDnN60VEohcK0ZL/70+0OJdYMB
itRJYUTWUbWH/8i+pE7MAmY5FPyDLW78rccYKZmaXJGOOCHbKPje3WdzShy6D7TveADa+GVhHlch
YE4+ei1rhp3nkQ7+CAElGtBQ1dyiSiRI+6nkE/mpWflrrefuuZ9mpE4SzdHINX1Rn4cEVR+YxwsX
TnK4NnbSfvNFRCXWdyT/s1VQ7nWRRo0Zmsa5Dv3QUeSJWQqmzbviK+DdiGDBddWzycbfVFSmDSiP
cOWNSwGyQjQlD2D49MWiKlkmgepIkYFHM4fLiZmStu0HGOWKlxl8a8mfrsCsjf8Zwq7G4q8MZZWr
ZYgU40FJP0bdY7SFZ4uBGxlTOTICPQi+5/nt/Xls3RGuBrJ1m/udUu2SxxSFivnrtWn9GsYGqs6U
4UU8IWo5dfDhloemCl4NPx6eQ+aQmYt0BD1BKA0BW7zNrlyjiN5phG3UdLwxXGx4piHuLsJ+NxP3
XWk48rOGSDlGy8WbST7rJSefLmLcYv+/2AnsVIcWTShF/19Xaq9jd4PAwZ3jUVT9GT2GRgkTpseQ
aNSlOq9Oy23coJMP0PnZLLZLMwWUFbWnuV5GeINS4JN3KEUCKoTGhqZO8mBAxH3RZh0RH8R+6mq3
dq61bsJmebldC+64LrgcdlXPYYaoZea0MfwGozgKgc9lMmDsPDzby0l0QpfDDZsO1DWHF6HsBzdP
2zZfBes0opxYmWNm2wZ/EfxGzhPDPA3FUnHsimd8nlShJR2bhd9Xawft/re635OO4YW0mEPYqM1K
YiWHQexFkb7RkFg+tuw9n/kj+3V9IVF7uc5sxG1QOAXP2IF0aMurHUhflsf59f/OijVJJ8bn7SsQ
g1MQXx0YdnkBfDD32UCHr1vZ1tqciM0044Ak8Sm2bC1TCENObEUsE22sVimBgOUun2X9nK9mDRC2
VmxI06b7l73qS0Q7j1hWPHqaokSFF4VJ5quhFuRxNq5BcJnEiwjRW43MkcC1lU6uoV1zIWij7QTp
762Ti9Er4Vq5fzOIvXSl5cHIjp7CvloWgUSJXtZ5BOZs//jU54RG4juSpneLmscQ9NUO7sPlqTqJ
NqWQpzHPBO6n3+S4gTPm2tk8yenH4uVv6GigEfJLlKsRyUgG0aLTT2afHbnmIdKnF9Cua9TiipNx
uJbYRP1h0lMihdHJnmowwrjir4gfwW4ZVqn/6kbrzqxMNsYykEnylvoK7rr5dcfpX7zTAGxmE0G5
tlb/xt3XP55kn1h5v4cUiCX3tzPlGC2jWpcaPbuNUYSOl/b7VuscZ1sWHXGS/uia8MnPdOFCY1te
8WdTd6kt2wOXNYFIc9wWXuFwYyoDKmKMYy19ruZb8QuLW+O/74ATqm5OX9buaYx2vrTZp+f48gON
X9xzLElxdBlLJBF8eM1E2jH6zCJsu12+xLKZr1efroKOem/NNmbveHIM94vUq6qZGhWwOuoHF71i
O8cBQ8Dqhh95LqvTw1SSGTA4hNsfG1YosJHSDEiIBda+abfbSByQGCtjLVzbuU2CdHlRqzo+uLLw
pKTQqXYMa881U9grrOHUIiCCr6IcWePz1nR/Ep4Nh76/fOn9fyvfsguT1zl8Te9fWXJDYH3icJ8l
U48RLkgHckwoEorjkLME/2C1nPslG04wYWu9Vv41mgla9bwesh6cstuITQwG5ulIwiIbH4I1SH9l
ebKMwP47RiTg+15UHNERYqwjbKGLNc2xhvVW/nesovyFXuv51mJ5Sxhg4Y5yK+vxkP4UlidJUgdQ
W2IwsHiu8XS0iknJGMm+n6rbdqxYLgU1mC+KKEZJTRdgkzaydzR9B2IPK5k5ngOe92ZYyHvFWWQa
2khYX/8hpNsygdzKjsiG2ov4HB/E8DjfAztYidAd0DNyke/ajozuj/iDfys1ovAa/nLcPNS6setL
WPajy/PYBEGkdTlCivcFCAD2up0uAVM5EkaBaHg5HotoqRV8RRY8DtEqLEraYy7GXgiDReer0lSZ
ZAja8QFfqlJV/AiFf3cob0fupLT1pf7HeBYKZnTSvqc7trFm3ugNtU2usUhxfLQT4aPMsDAWIKGp
uBxB/2u+wppP0L+PmQ2svVNBBTbwyxQx3tzjCbRarJ4u4U4uKH+s7Rq+FbX/JiMfd2F5++SupXI6
n+yWXTMcXKJtlK3VpvtKaRXisSFi+wipLKCkLDPjeKRWqQFEd9oqysBPIVbBCVdtVOQgdVhPN0fp
wZvR+itcLtTnyYB2ocf6cY/1+a+saQckDSL1YrDDxa4+WEzMCuxSbAQnZb6NlBQo8SmUsS2T+iDs
hSonSVJztZKQzRu5GGuX+NeMgBjp2ocDylCzVQFDRMYtjV58WWhjV4R598uZQgs38N/FiPsuSobK
tGQozKkFP3cioUOGXJByh+2qTON5XlKfMCPl2KTNV4D/x8buwtiQj+5t46OYI0MB4s7tiesUaw6A
SxDilgy2D6eK6lpAI+3m96ahNrYaZ13sx55efiW/ipZBGuuYG7JFV67BRFF90RUohjrAWB3maQHF
0Z7kTo7cq6vDeB43cncV1wZuNPXsh2PAmGiF6K+0k17RQJInuXE7FBe5TTBVl5oZ0MVThgcbGreI
GoUxQmBfJc9erw10jiIF5X7Ejz5gaZCLNhSrniF9+S0P/5TS+roVrXjkjZbHn1Ugrlvcbbz7v5bq
2m/kEXYO/NZAMkQ5GuggBiajvBCT5xzmoq8XAG+ba00chrm0GUtR2CS1wy3ioyShlJ5wZ9nrUt1C
L3TFgKcTwo17TPZameTK3W9Jnv1ZBr2UM5sJOlNmQFUEO2Blv0pdirjeIHTJNBpoW3C8cUJvaQdE
dT0uq/95w4LdhdZ94Xsma8YoKFdfdffsQgLKBElHEKytOX9azFYgvOZ2WcLVEizHjthS3QismneO
A6pNhGNCImXLxcjroQQB9iLo/8mu7BMHvDRCZAhMUDVwpB4vsv6MP5QJ3qX786HYt3frp45sHSPI
lwyzH0jllZJYv0srs/HBpc38kkIKcZ57Uyf++uhPG/ZQQsycl0FZAYZRrWvURt33xZcidZ4FZNp2
vAsoIIvwc4vM92FYszjec1GbbPnPGSwHD5Ww8nGrv+lopUq8uL+5ZDZz4bmjfVVGqddnK9JIG3y+
DYhU8l3YYyUrm/Ya7c2lBwzJR1q0lxtTWUeJgjCs2y/jRUIKwcCy+yOx2NG6gQU+q2AKMsoSk7fO
iZAgvuFSCoWfX5oZ/JzgI86Kr+gTTexMp7j1NYpzsbBKVVXv3s22n8CtF1RALwNOhC4srtdTHdVP
iMjoS+fjELSo56vih5be1VcjCi8olb6H2doga13Zsd6fe23oka80JoHxGmmE+tYkR5WCVpTs7FjZ
FEZLiAqES/TjbwlEbrbn+4YHGa9X3Z9x9ke/2Mij7QyppXXJQ3zbyq0QpefZxK7a+36DLQxMZLBS
EPmi6sR0JchKk7S3zraB1KvgddzXKalf0S95/NR/kEd15SNsQG0U6VTsH19ku7o34peu3/6rY1J5
f+HNnSF0noY7E/sDERkLJGwdO3DDJsIIC3hkm95EaewxjAKZC+O+FJodW8yo4bZ4jURiglAQDwMV
vSxFPy6gyWytmakBpDka1xQSBZ4E/U7vWsH+YYCM4bjIqn/Mtd7D7gJa14sYqaZJ586CSIlaEnX3
U/sYHAjGikV4+JkoqitsMLObDQP7HzIEIpHM6sI3yf7QAL77dE0g1ZqiJMWdvtC+VfurCw57qTJA
pN84/HZhK0IiyjvCkmyAkRgkIYYUD8GfQRDnCaHy+t4mNS1M0rUzRgykxx1bQLAlTh2/OPFCtNmV
JPaM0C6FiLNIyoa8n397IGnzoZ9JxGs1mjtvmV+gRhY/eHpphBFj8flIPrG+OgSstyh0wldkfIWj
COaLfwP9YXSJxKqsVWVaQkwhaXjAhel4XxFuxu7IitQcOkljS0UPw//FNxYJnKv4KSGgD3X+c8r0
OMz9ylBXPQWutu0GuL2fM85muQj75HMZnMAvchCjl7gz2BRlYO2aT5K8l3NWgTOaJjq67qcoX5rQ
Z6sDRxDA0+qLtPW33ev5JIS21+jaz0LMb3Jm5YUu3/JwgC8DmIGfXdM3dpceKtFv2KtcXWDUy7ZZ
cPS/k+7RMgXIO3p0FDE9Jpv9vcDlHPsJE6/8cdOUHc8HOoXduOFU456xIZfNOn2Rp1NnbNEnJ1mb
Z80Bt9bbpC+EMkkMPetR9/mXG9U6xxMFnmSplM0lPRhAGBSQQj4ebPbeyeqet/mvliQxXikl3kQz
SCBewMWqsAHEIB2joVSyaqZ5sNaTehkzs0OMbE7pG3A1/V3vyo38kqJWBjjpDRI8iYzKEbIatWfD
WA1PJQAZU2wnMiEO/w8WUqNKriEZ/c/AlTEFQ71hY1oOE3RItUeuD+OwsCx7oUcA27q6Y74c3ODG
MEa4Rt5MbJkKORn5iXMkFQUpa3r7uYLYGv/zIZ0WgKpjDbSxX+XnHgJqRZZEsYdvH5qGoRI3ygeZ
5bPxLwDYB4GtkscrKzk3dax806doNG9z0ClLxBADKhhZMDVLOr81eASmZLK2a1psNHjecD/M4szZ
9y1WXRyV4bMgUPdkwWPGM/Ikl5/7bD5f/MAJ6XWo+aZITlt54GuDHGxoGqSz010bJzjIT7LcLfBj
0OTlIKqP6zvfVSdirF75lQcz1q2pv0+gecmxxgNoVKfJFc5rqogXRgMFGzT7YWDrW8wnuw08QskW
jcOf3WkjVgu5iM4kxNnro8GKfdII6B4KvVbtx5+0MjQprm67PYFJ3TCHCHemejbFOBZwQp+ISZH3
xHK+LlgAPEkFtjLZ5+TRNNQvlLxWUKu1XKw7t0c9UzHPiDiuyP35t5EHpARE/ogSB4lhsLlub79Z
C+RL9kX70mBmD0v0iFS3wvQoKG6g1JHMvNkBsXAUhB7aWsKKGBY2fvI+xT2JbtOhDJEXqeHSSYVX
zYMm1Y4P6SidqsAxndBY/2AtP6yltB+jMzc7ijHd8ze3MnFki9spzJoZPv949O4An+IgS9J9HpJr
by6fuD/+oMyuF28HsaS404FTInIjInvnfc8JudMU2p8npxK7K4jvsKkSR+Tif1U1lAhEt/W+w2BI
lmG/bpF2I4qniyGYN+2MBnrkI4l1c6H4t9tPzdo+CaAyNM6HPEGfw0IPsHa4/qJH8Oxnj3hp8ML7
PBR9eiCC4Tf97Dky4gEL/VR6uiMI/68TFYNfBjrS8XAbZKONX4jTQbjGSfoGcyGgo5GIq3SuRSok
OPctrsNM+WC4ZbCV/yZa2Kok1v9PaKFQ1gl4JDdj65BGwt3mPT2QuPa5scNzOhfRMzDvz8AXihVf
OoAMsYn52UXJFuky6P3nkc+spW0NTswIvYZbEYLB/1WUjN+0+QtC7OKT/wLrGI9vAFhn/XFDD2LB
8objR5yT/PFDfcWAnCaknbNwfpwNCrDvlcgD7wS90/3QiF25oUFkzJr8geJxO3UhVYWoVgLBk8Gz
N4eOAhxgkKp0zj9cSKYqQPA/sLLgNwYlOgcQ3UTmxzo9SFJlkYi8pPwDGGaYi3UlTsxt5EIOL2Bg
OuIqohvpq6L5XHpGGTUT6Po4GiRa+U0prcke48LrrIJwZIumi4Tt1eWdNKlBYySfW2YhJ4/e5WkA
zxVF1U7zVXh/sCalkFwoPhYWSRjHuENRSyu4NHz4BZHgYqYy00HX6V8X66Dz76qMi3X08BB2pwrF
wu1gUq+e8A4tnuhefYC4Hk+arEzx5qMwmix0HjzGoa2KTU8H+RuCrTXr9WySUAJ+cRX05Vpu4Kc2
DQc/AjE5pw490rgH0RfcdlG+zUzUNqwUlTubhgsKxdajTw7NJp5Nls9DvYu36QxWOTnZsVYCSKgT
7INTLmsiZBL+JeVlyZ7h4xKttDNQBUecmIRACW+TKs1Ggn0tos92lb6LSN0MhXHGvlmLn1IRWIy8
TeISFhhIUV6hH2uU1YJvUM29bIVfjimPavPNV1MkF2uFyXoHPNYajDa4gCvoaMLrxgdmID3V6wVu
4od9AyKesiZr/7/trAJHzJgwrssi841ZliXAFsAd+2zIeA5b2nnaSQ0qjN3y8EgToauV4YDMvNm8
NcTaO6cErHaG3eUI+eE5vjJZsAJ16pzrlZ5tF/U4+5OpL5D+i2CbcBe3z9dnFresqW21PC5OytB3
HMjAMesTHAPLHFkEx/rTPGVG8hV5UYlSMph+Aanc+KdJnxyIo9fDasbaoNmYclM+fo9IkDM7P5KU
uZCSAQxtL6GALmt6feuKEScLTCfNhbhqcZbPX03gQ48cD9v7j5oqFWMsw+qb51NCRsa7/ZBMzFD/
mS4gIIL0PB/wE3zvtbWKV+OdOYv51WwMQKVBAMV1RBqVh8O1R9B/CehXuqnlJGgPrfA+Lwdtlxuq
w/NOKqnVVrjF1SII/214b04+6EkqroKCsqEOasqtSHbkpC1UpP331qTKjaPVtCnRUm5D4AXSFyv8
rouji72BnSpkIZpNzTNu4uCzGLKpHGzbnKeiFHYCINdyvUB59N8dS0PvefvoVKhZgY8CD2o6Zg/p
PLpRqjEqtzrbsjja7IcGnp5QDJ97zRFZPN/9KHzCIT0XEvCveFE0NNbBVCvf7Vd753p66EncdedQ
tWmEl/4Kme/rpWYbOo7ABJwfuCJ2RtqSxjD8ApOWrYsZuA861anXW/qCYO1JE+IvQNA3iJEnJPdC
ElbJva9fa/fBnokUNmKt8S6c5T0JdPbVrLupEXHTTlu/QFSg1C5bFoFL9HP+kxxnDUjOOI9sH7i+
24cyj2l60aKDbVp6f21CsnRTNU0VOwIxGV1VumSmWoIBZFb7oWX5ph+QWcJ5nEc2AFYUGp+/wigF
TNUBFQfVF9mUm9EpC00RTQs9pCk9SU4pPsL71c4eGjjUklgNzvOr2BnsuPNi27SBIOvuGNFisOMl
fCPQzC3Wi3IO4C/ksskfNRdwUdyoEOaHN/Ah9LjdXhhl+9+RSYCL8sgTGUty00Us7k8ZKBzX885U
uUgr0eENDLEf6CgzrrcabBZcku/g0ckpbObLRJCL4OP6iOtsKKPntfNspdOOcsLysxvMHtvoFAlw
v+70TzrRB00qZkfNNGOaHqym7Xue/qcOoT6TVa1dVrO4cuDXOkpXNQGMgYgDgCf7LMwRa/mFkKMg
j3q+9aoxAQPLatDhrs9dHdWy2E/1rsVKMHv9hD+LSkUhnWUnWDli2KKb7xZQ8Bpmx2ZrRd1QLY6H
CY0fr2/9LcZKlP2vGwwFudIjKdgk4GICTgb+QaauqL5yWIUBKHCAk/EEswSTllXp42T5SKdkYMlX
q8YapGjDhO52g1OlfIjQ7BTl5tX+HRdN7djkKEli2JqSSkqd34zYhdlByC4bdRaKfh3+3xvm+xf0
0/bXBLb0PQ1Uj+jUQpRCJA0rQHmO+UciIxmVb1VwMRQynolB2cTk9e9RCBud6cc0GqKEiPyRePW+
+y0dpq+kHVRE3qZQ2CiKFcRVajv1gfU3pKtWe5MypEwWlpVz2WmKxHqaianu4A9nJxuq+8/zycmB
qwPLAoUfzE0QqzgkN3ozxpifpMbLkccvmGzOZDTDhxROBfThBB46P6CpsHWefCJe1mhZDgYMRr2o
FoINa1aRMMdwHuLKMaHCfH96+R3/Rf9aWFuz4vPDh18wajUKW2FCasluWcdFQGGNPiylFPC/32u7
CILZ8wmreVzSdec9dqUsSu2xhkHlh3moJgpEnGtXAhTv1oXEbD9l0O19UFwiy2p1xHQuDq/3EUAx
SK4qnEXH8lWU3zLW0KIW5ME90C+xXE52PrtnQ51fM/d2O31Ii5CjFQhwhctQt05DRK7K0GRQeDQC
uEQEgebpEF8BFBsL3HQ+EivGrwQJu0THLTStOG6NQL1C7H0GeNdGbAXoww86rmZyCCZyqSybVocH
re3z0wWtzdhSt1iXwEbbUJmFq5dmY1AbX9FL22fUQMb/+rTF4hTlk/UfACRu55x8KONXGtm14pFA
mv7CJ3jbCPEzvTm/OBR0kCi8SFG5Jsgk4s5D3nBvtYE67VCrKXwkzMxhpvpXhWZlO6VLq6QwV99H
jzlB0n6HwuzSV6y4HwmZHmv65MB8fnh9dhJ2tXJRA+WqIPN72YJD0oN6Q1eTH3xys+gPVP1b3v2Q
TeE8wNRj0ZiPRYwqauE5ndp7jSqIptYK9+fxZQ5X+iKupkPQOjSBZ4X0eLptB9507QRj3PoV+8as
yCGUkZj7BwR5iXyZ7PS8SAdaRb4rV72Sh4jgIO9R8h8YmpceP+HokycAj3AnZm4ziPyuHJadRFLc
kuraOUv+Bj5f/st0yOCCbSqPecwe/XJQlt9jm3OAinUZqXttJto+679Qpx9HHq5ERLb6RgCi6Shg
UKSa2C8KgPlUC0Dg8ClDL+3Cb+FBXynMTspYxksrpGH4CTVqKCmx1swtzHzLYbudUL1qOVlotDkH
fhoiw9qT+LObOK7ZRRUEcvFGjLXJNERDpxjkyhixeq8iIfkFDXIjxthx61YtTBA39smpVCxWM2mq
Df/g+f/u40SjXUd8L1jbnTbS6EoczKM43PUZPoTTa6NjvIi1ZUiP3bamtOFMk+fXIHMG/Vm19uQ2
pCgOU4vl5jMi2Zh6k8rKIngS8CRhfVPp5L//0uPZjSoyG2frBqOFTqxKGO8G9aXvwPgfYcccpjoP
mHCbatLulbQ8nM0IRGw/b6Tdb5ykiLtEWdI+ZXx7K+w7vp31TJmIMlRw4OeI/QKLZRX9nZ734m1i
MiruENE2wcSLnzEDM9jzbqxZogl+rGBMv16E9z1FGpzf+l18mMF/7DlGnX7Cfu30XqocTg84pFad
CZmX4UkgdL7UtZ4P/4YncytNqQw6Dz20JoW3NuKANvA2EKlWPaG1Nrg2OKqEg9vAemJlGtqy09bT
EU1C7t749O3vW+yTLXzIPWBpilKAFtHd1QXh9MJbDhi8U4/TCMLGMJK0CsTpuzQKMArub7DX6phc
4cTkIhrAL6kx5z5Ono+k945cy4fQ3iVZY4+9GktSRvW1lCQ6GVDDHHtbCi3g1kDvL2jfopWYeucw
CosnDm36bCFoTuAHOMpT1/BJdZQSuiW/3thIx8S+MBnLE3XwJFir0UWXjFJI/FvjiVf57ClKjuZT
SLuQVxILOA13eqqISdA4htMxltRgl/qkKsolilSlNmv9j6N9KmAsNr3MY0yPwAanjp8v/XxaUisT
kQMOg7BF+OepCIV4L3D8n7c465iyc0ikK99Nh6cxLkMLeZhtl4fcBipGY36zasd7OWmdHXGLKZUD
rig8ggJ8SrTxSk+1MztJECkigWZkNo60BCrva4xQ0NaiW9jxIrFS8zFCfY58dy2ZDvelqeYVdc7t
itNlep+IMzTrdj5U079lbXVkr+r1XDHKDfYKAaNf6zAkC/hUgZOdzBJNC1XF/lDoQN8ltAfyqHYD
kvbMC7R8Z14knfVrZBbNZX2VPGmohg45MQ58yeJiia+SMg+0EB+TjSEOIXdyos992DGBgjdFzHed
j/4O77L60IKWl0IyJ+JhVKAoRBLpHh9Xs2Pj/wIg6KooIfUzEvXAwOBDqqu27aDSq/3kIH2+ZBBF
r1vqHKkM6x/S1dC5nVz6IScRDuIiJRzOAe0OUHMQpUd+DPLsNhuNd2rT2PK9h/nkrDWKN5Mi8HnG
wQ8c2gKmT/YTyoMI9PUN1sCbHBhQW/B6kk6mDOyEBjAu5bBD61WsqbgoX8B1mWCyJ9Spbcz4v/fd
7o2sV1ONjsJMxexmbcTG2XzWYf+goj6//skzMJzxN+hZVUsFbF9EWp2cpATwVNUq5ziM9MRUaR6D
PNKAlrQjyfdhHo+tu7vv5c0ydhVALPSAb5gIasIqgt378vSFh6ZViQyKX3K2k+vBaZ7G7bINSQpt
qllSxnH7A1pWiwrxpBI6p2mc90oNzs7EqaUfhAqsb1IZCRWi54xsFsiFJLhbCCalgdGjg/iWm4s/
0H1ZttTZJLWVs6boDI4ta8qZDb9yiscaQIxtcC1CL1pY2QKgKEB4GNDz6WnYFA3R4qSRnSK0DoY4
lNJnerNdlXjG7721Ke8slvaJnJSIJOgXdAJP7jJZpEjsz5tcGLyKWhrjOq+ulpxuP/Qbl7fYdkJB
eKseoISNKUPCNZvnBkuMeUw6rGhjwHc9o8rHkeunha6cWrj117URIV+2WlIat5+9Irt/nZzAaAEK
lUbIPcxOrjSPW2z1lj1EIITNSnj9FYrvjwniEQOtl/5Ka8bPy5Fj8scJVTpiLaiYAGhRp12hyP4g
QVJ+ABz4qCR4wvZCKWc0F/pC731etoN+u347IdP5tPf9faFH9PP3QP86aNsN8UD0fKD4vrlkkEub
2b8l1+bMn6QHU3T5KVn8TW3DTxbCtjUOMdTc9zNE9hTUNIiCWcWFUsrgfmIwZCGvTE4JFbvoyXhh
YPzcauspIxbfCvxDsjWtExLIEUaI8hsZwrzYjdt1EW1AIx5FaNUKHSVEGPd9MrCmENi2lhs3puKG
asMarSnnM3X/i+eEcEdyZTRbM+y8TAaJQE+2iilLy99wB+H/lJj7by7NEQKkA5w1D1mFfoOrdVlj
/BOe5Aa9ifsryWkxQwEMReuW1fZaSqbgtx26thWM2yBujdo/17ao73vWt6MfRpE6M2MULVaSqyA4
q2YgdI5+vvE5QVKXU8HJgIDv7zF2yBBAgWm4HFcihwG3TVepamHpSP5Q/nZnVa1x9Liqgbr0P+4/
XnQZ0GBYbodvfHtkAt9TNE8OLUnnlHBDNcghgMLF7+DapTl5XI/Hi3wZ7PJ4S/f1yMyRET6WHfu4
IirEjF1SPpDpit3TIiEDKPasA6i9rxbOhCRW2Env7zya5raZrAix7JPZvBDTshrti7PmhJiInORK
a+8dbxqMQdm3CXbFBhFVd9T2bGrKS6Amgj9AFNCPdWFpMZqTkdmKY8/ebFF995Xs1CDgdV5Ir7L/
J1sPG0UnZ45f0aYKVTfS8z9XWE8K0Q1hNDgpkz2ZwXPxbyJlYKHjnKpgKh8pr1TpkRSmeuTFXcGl
31W4V5Xu/CpfJS7/tlNBh2Ba1/tLhwxP/gDWi39mYSgk44l7vka0g/hznaBzNiHC+te4qZ4zml/S
Vf48lHjZY3Eew4p9Nv2H5S1BTEMoKXzIfJmuaS2MX3d8JHIQ3hoiHYcy71CnR2xljDWR3vQ5zp5h
cKUlq622rJbJOnM/V77RxsmVnoV4buK+OOk24TWwp8h8ZulEFskyP7iq66bi2uwzHwr3H/rSaFqh
lBSML9R7Ey3sBKTnFwa2Rr55we/s1yzjTGV5ocwjz3iJ/TqUmqqtp3Aaz7aVBHaHX0gJLy04KluK
tNuEtlAlXCeFvFlbhoyncfmqX+Y0Q4rPAOAa5gZJvxkfHsmr/oHkLz2B9ATnec0e3oEUawWl031F
soFjoBkQyW65SEzZh+YgHv0zL4HK9QNBD5PtclqMGqj2Vz7Hmnskd4RpHug2GKoFAPu29soQx+Dk
M6WRPuZnS2VWFtuQ1xvXm/eBOLMPS+3T0jyc8hXSxH+sTo2a0oyDREgXZDcBkDD0T+VyJZVj18pO
6O45Zgt1qlMhG1yOUb5NK/k29X9LeibnD9t2IoPAKxqvP1bdsTpsPLQPeN7qbpL2nGxTcKlLgmNM
dh8AExWSFgDVyLXBiWnlTj0LN4doKA3ap8ws5UTtjhWxukI59aCGgx41LericfV3yDtVlBn3LPDS
TjDT4uet07gztdUkrPMHmmhWCpYCy4EA8I5x7Ns1X7hYY1PTEPyvDSB9qyJueIQODjtRRln7Gqn8
KtkibgIFYXbLcKpxtN6DS6Fz5k8vmu6NBSmlgROiR1PF/ivttVw6geP+YxgPvZE1lvsxcoOtrCff
uEtQ7GUq5orI1Ovcs64YgNa9I74ef8FYHW3fFzq0OTzYIKiYHo7Db8r+fiuJ14PG5mzUHShrtbnh
eCgyKm0dWFraUl+SLyLN35gnC1Gn0xcuc9K51CEYcjcDIoDoJaKQN4foHlcnbwocyzeaXuo1bFsP
yq0hjpxGKQqEAgikFFb9pdyYCPUFP3Brcvr3Xcs6SZrIALtF8z1bORlBlhwLReJSALfWEu9ox66D
lKIQxhB9015mc37RgIzqEekhsifEyN4c760Xv+lopYkIitTo95uXracM+gMz3VA5CAaReoN51kfV
tazNqYqbUNQph0HH5Io0AWSnfKdOmCcP/lgV6gdqvypeSaGubARJchz36ohdqAuFALuolAUs137t
pPWZChaXSA7baDCzlsUgYmDAtDMpwsOHClv1lGHDzrJePjIhbpBsFW4b3XEehQKeMDo5FuhzWKGz
XyA3+PElmi5CdhJV+DI53N7XwllEBSJpWGADLDegNfdOx3OaNZ3v2C7UWzadNASbN9CeIpnih24O
1jxrtoAc7EitJKP5oBKdGLe6aPJJroKsWmj+bMSjkYJMB6plUzX2k1ZVw/hULiaxT87IzGcUXcxt
ef5M1geKXB5COaqi06yiNnXKxFuzyQ9bgtke+SDPiplHJIEHwAKQyO7rltg9OeO34T3/guswd8p4
/G1tvt/bgaf34/pp9v/AYPAIGzJdpKa/P8V6MJdESlEG2EFbyi0+9uf0h1636bSyoED8qdWJQU7e
sMITg0+lEjxytYDFhSy6Tkpu4UL2P3gQJtns3QqbBwlXgA8W74kRCnQRLcDSPOmLJ0G0y3S/nUzt
F/oqKFSm0cFM2IGrOgZkwbKaWFjQi83+dVyVe8yAFJRU7pGSCOHPQp46MZWef1C+Wyc5/AIoQjmH
S8sF2vSlpXelcdJ8SOjEMrKgfzS9qb2MyZ2Nh6fdQcTEQdOefFThqh7yzoNCPHeIvezwNXp4UZ/L
sqCs6uPSjSHafDN6igckMbdqnrWbKaGuY9BPHhJKFByhV6pKwDevcso9bqn6ZVBc1haPWxxB5t5s
O4G4xNJLV5rzO06BZ6kzhsQoEezF+WAJQt6eZ5Gw4G4QbDlbGmgjQNKMSakhfTl8Vqav15NvW0+h
V73E55ui7JuYXmOyGZoNpj9BfUSgvTEsQ/GySQGMFcSASYCy/4EnLnXY5UGvx6yL/Z1oicYB9F+r
KNK/QJUkx3Xr/XWAA3iNPX+CL3jhyS3zF6oZ86E5QQMmGBaWT+VblJ4zwAX0CqP9gX7gYM8XtXxj
wAfKK5x8xyGZyJDtkMyjhnLehuKH3DOfJqGznt1Pq1wsS1Xe7ks4CLSBDKrXFwF7RWkc66T8dKhY
+DykSnOtvf+IyIb/SZ2gGjhQFDZmt59OZo03HD8uB8imj27GgQItJUycRr/S8udGRVoDnXDrVLgr
exsPA1+Sz8NqcyclniiF1S+BxRdexVNG016Zfrn1omMUfX0hESUjoIRu7e7POEEyMGhfIRbV7QNo
0GbVd48P/bbU12KqjfcYWk1z+FmOHBO+5J4ZG2GYf7wrArXKXRRLHw3QeUI0R/HGZK7qaLpoOr3T
Z93xc9qyRQ8HT3QM4IIcYMFM1gCyUPTnBzPaiKKmqF7XTpRq+bLyOYWSichLkZwYF65y4C1MJd3C
M3dd9dkjuiO6HBy3FL5MeQNqbTijLhUZHx8+rx0+1ZKzel8sk1/6IPjnNi6p5DS3lSPfg9M1pEX4
lYYlyypsEcKI4MSedA2mRCAPb1GvsGshFrjYpCZ7KH89Yc5gfEdpcKgNgDbty6rCRNlSnYZp1Veo
0vwh7H0kPp1hLk4fNAJrKTa2I3C1in+bIeS+0ke/sl/vAqQJPFYgy4N+vWwNW1GdtlM1PsTTFvIi
OjA2hr3mXoFOVHeBUsHM1TBK1RpUXPWptylkpH3ncPdazjNVteOJqg5WpHrOUoo3+C6r9r4qXl9s
fxzGyeE8w44Baxx4oYlan6XKOxw4ITCuf9o03OLuM46IFtyYCHZTZpnTXNU1fFgE+bp0GfHQx3e1
K3eJ3FPvWQO8pg1D04IcbzN/Z4sJ7WTOltyMiP28ciTMZ8vhRfvPPzJ6kZlp/UsbeY1JJ1OyeL0w
iBnwf6zIwbm/VLOG2PEAdlJxMhpO60Exr+KANznRQjgn4dvuoFrxBuCnEHtKHGkPmQTbDPc4STnR
wOWFy/zvOIpFSlg/cAKoxVifI8I3Wtaxr/IcGmzV7YaPWZjQEEwJWB/IoK6uLIy2NKhncTF4Z8yV
47LA1xZv9DHNeT1bhAuFkYvMn3MYwJo95Azm50G/0d8IbDXDTuNQSyauqRjLARwsdlJt0XdhYL50
kj3PXTrdG1DHayu43wdMeZPW049OOzBgIY1ACp7y+h6OgedTVO8bSjvcbliVtvnWAgB7JvqSQS1F
PRBrxtxluZQR6Qu47e93dOSiSMzPX1Z8EhT4qBMRcrW+jYIBSUA8nWHYgKWVtlS0dsNftS5gHEzt
Lqf8EuvPc1iahfuzV4n5puKUV9ccUQNL4CdjcFon/ep7vYtJA+KmbKDPDjNrMhBKYbcwuC2pHPAs
tt5YoSkixvsMMCi/IgDJNoQp1EnliPJxiJ/6z/1W6LtG9NAitt9cV0YBZurNkl/fk6+lpDbcIVxy
uLm/s0OMCRiqXr7wLUrbsTnlLCc78HKfFlJ6WG7JDoezAxriahxBEPCH6U2JgsQf6crTjovSStHh
JB0oQqth5s10Z6Y8rdLkijEE3DwOxUKM3d6jezxzV06SRADw0KI1C+40a5UvLIhemsqRD2qRcVhW
Mg+0WsAYy/ZwGtp4Y9AY7jHfW6qJLKL7NTtPba6nviVhwCRG/T26IC0Z5GsrlKulo+HYGxoT2Ju3
MOmTBG5VoA9DjOTNSbBS6E1nh99Nj3zRpPRpVX9cQWv88GKIT3F+zKxLZNlBm7GurNC2+SYgUBYX
UW2pBxHFxJOa6ONZiHXOPDvaIOy2yfx8RC3T7iWngkOmkCjiSh7PLMvA0YO30jlBVNPA+61vAOZn
NSWzGuJA0UwpFC1p0O8CNlpmsURZ8KYWHe3H+k38DAIDrDS8rQRNCBm/N5MCrwNTu1o7BKAsEkFm
srV32vnPSQqJq1WGYucE0C22ePJ1cVNDnkDdBBj0W/PiFBa914dMQe+P+fNkA52Yc0CXpbx8bg7D
/zyJC874aqxaijgMkrE1FOU1Wr0r5dth2h6pauih8MDBUetadZ/12N5IHyKxdYu+NsoIZWQpSdes
mSgTng8AyTT1UHC1n+QvkPi5G9I1BtlWig7a7D3aM+QW/cDFQbRN7GQyVuh2Am9FLb+0YP9pLHSg
N100UmxrwYv125h0zf6P5bZWpgYeluiTrpCoB6jO5PoycvNpQH+2pbNUB+dodV1TlNrWb5vfT/Fr
TtN0Zv08ZaniMgASQXwaqKcKhnpprJ8JEFMJSSsbv47icfP7+6KPar7DiBr9RBu9P7Cenn6p/MJh
XI1j5iOLbcd39zUl+aS+7wxRjw2eG1H8kjdZ3et6l8FABfUe03pMNA644ye1PLNqxRoOH/XEzl95
KCjho9V5Qk0gblzk/m8eoI24d6GcuWwHJr80wpmxNQg02utY6zrY5RjFntPtQi428ZzoajJylOfA
7mpR+p+guCbXnOZ9F0UpM3Y16o6K4duam40TC+Muu3Qu7Ed3aZT88kGFuXmO2KY75lmDH4/ZItU7
/4rx2+6YfiRq1ftn4DeL9IkIGR7rDkWpflE/F5/qO4FnpLIVs3KjHLnetbKLc42m9/K/s8u9SE1k
LqupHwpoAYzZ7Cy6YJXuVExG1xG/iOB9rAZbVjurMAh/NHKenmevGJ9NAEKZ5U4tqKhNlYuv3esY
6pK9L8/+hAsHd9xMtLjeaGZAVyofwnptawPETBriCquutrjHaN5H+88Zca0Oe6FO5ontL0sVwYyS
kQbJY9fSgou43dQDn3r9DIZlIHfm82SFfx4lLWDiQsKzZFy1c8MHdlpJDzs8IAdQVSRCepVBitC2
14ilhMvC2riIT2huUR1RKkZz/MyCJPCj8ZuCtXlsmp3XTlkhLD8vFnUDzvXDKosc+piwv/5Wtu4F
3CvLA7gK/HoR4/GT70FBfokSY324dES2nq0XZkHok4l8WtRqNI9V/+VOLL/QZCBH9czj5AK7ON3R
n9hy+tGRGOSpuSfq1Zs613k5ZVXJjvtikPR/8KZIs2YYqjICJOrvX8F7uicdSEgXuqNYiDc9qy6c
qM9I33ogwr0Pe33+/ud/c4d8QHyZLVfeAimQKuxf74IQc+daQNwiEcX/d20PesEvIlUFLQtT5tw9
Vz/028BuVW+8ZtP5QKUxJX+7vyrbMIuAGLduAkNZ6Txmw85CbxuP32/j2AuEosXHyFmA1+OoMxk/
Q/MloJSJTH161ziH/zDBvlGC+NptvnDkKLxG3NKtmOlbbwhR9YvoJwJx8sotKaJiPAXbGUQ42GQp
digM53XBXbQ5YHHYk8SoMXEMCcTrtZ3EFxba1CjOjoE+tf3WIjWoII1xCavA8vtcTOdweJIc+ySp
FbNv22GaM54fSTCjdcJeYQ4RS54vSeP95OFAvleqcihQrnnd7hLe0z7EnWRYXBrX2HGD97S40/aK
Ah47UiRX3Hvs20NusADT6fGlJvWw2q0dL3B92hqW/5fEunxenVTnEwh4v+zWbVrb8BbyI2AR5vyW
edeHcTKqAk9QAyB/WoTSTTPTTDQAWlBpNu/BV+2781Q7u2mnOb3Q+vwa7thiGrUAqAoGpAFenLiG
ijnsoYyO1YlTvL8agTJx7EEbpx0sdG9SoixiADX44steDXiXH708z7yJk3Hl9FgPqxqdTplV3QfM
YIcVz0YJ90KeKdoIbXujltgfWB+HBqftbDho4ellDsz5+AoHgqGQrpdTe13KX4YGzGcA1F6mU907
rfYRXy3wX/XjNY62Lf/XMRfQDvQCHWuOnBKtSt5PJaS56wSI8LIluotXu3hFjiBl96PVlDOVm0R3
7F5esDF9qW62WXKJtYbDiPgmjfvdbUkvbmcHYTcyBSMIEJrys1wVqjqWxSkRb9caPg7tG6Wkvn8b
8snAdCkfDZAfmCEzukWJJkEprTvS58y3b55JKv0Bzor11MUHOJZS8SfWWzsxo5yshsQs4EQl0RpU
Ei+n4yhnuKrTp6UsUbWJER8f/RYYS644chi176qx4wLugRry+1Dl9QYwDh6xqWQUPQwOakQfZUUb
jeP78HgRHqIGQrrtu6Yexgo/DSiNjE+PtSnZ6UKV1+A/1NCWv2FuEHLi368a6Tgip7JjYA7daiix
Pepm/6dQDOTe5kb9HusC3KdhmT89BUS06J7QUcIp2r63fI6xmVWO3dckYzYG0GcunB+8bASP3C7A
Mw1HzBEdJxF+02I7zwj52fSg2DiRY94qDs5n03rm/vfUGWGAZrqoqdCuDgWKqHusKxtyO8SIMdrM
+QwjDOrOa2LZAq72UgG5mt9PpmyGPvMQmmMr9KsRWhczlw9FUBotsgixUbQD3JKohJcU+1pwkKpq
2EpYBUnYQS3b3rwdCKWSFiWrU5m0EVmLI+CTm0Q0RBbMlDI8rqKhUovrLO7BH7lVr4T4F3YNze7L
/HJHM3D0D6awaJGpkL9YaLrHAMXq34Qzq7eM+2UG1JpaNj6PJqeFqIsB8Yaa3xxpjFmalfn77Adg
Zzc7QiGnDWPWOk9kfN0FN9rHaCWeHkMa3sr+rL5xdV99Q0EJEx1t4OUOy8cZ8ccHCeKc9jQZauej
ggConhhs2C06MWtMuiMtmsmYfb1QLxd5aBqthkVrrWv23hd6YrNkh5rT3KDZIKKPSrUy+LLE3N8H
VeBAuFmuLRVxcYP15aAYTIPQTN031pe/PxgH5RnRHCVonsV12FP/zESn5IbCzGT40EvSIAujB5OQ
8Z48quJ167eScGgmhJYb9LBHIWzXM9CKfFyJ+Vq3nlwrWK9bf0ZglfRq5OJMEguM7gj28Fj5ZWoZ
zxO9H4s+1XChYQMOiFYn2GYrt/QdFHdCiDowsQ6lQfrxf0NGlhjDi02YuhdBQLdEhmJ2DJYdwNmT
9HMB9yIG9pEgutFxcIllANW0BnMxfFgy70dLlFa8kudERrgTrtrzh2l/FYTLfRPHP/74T619nAaN
O09Uo2vA3TSlsM7fT6ptQXXN7/RmQEuwYhhn1ATP6qTHA8gV3GMZiEHKXc6YskPPPmqGGXBql6Z2
vZguEKIYm089WDLUGVzvSrOoRTZtBcJbz/+kuMJoMXZCNb1sN8l6cDMUyDvdIlJOHSLj4/PNO3np
g4k3I7i+UBfsLGECj/vMXfytTTQn1nYuroMuUxcPMHbScclk5jO3lrJ/BiXX3H1I8QbfqRSPcBsM
0n/Y41fqW3HEYpzBstwHEzkE+2SnF7kWQpSL1ucouyhEcUy00IpfsdvHOeBrX/BDlKNpA/TMxpmV
UuYjYOIDxIoEoOVIPuPKqPnCeF4A8mdVbI0vdV+egVKFQhzn30k/5HfoHIpwkpMioAQxcRPoqxCF
yxucgyHv2Jri69QdeeyseZZW7p7VE8Q7XTu9nEcXbDRPw1h3U3pfdbTgge6zqar2hV3hWjy65g2g
O26edNmjnN/6jhADbdl2fIw/Nem6vqz0N8LPz705wQSu4+rbakfXcwTueEDd/9thCM+lOPa1brKw
Zm/SeYX8OlMe9y0BFDFFsKtc5awoUGumjqcIs/4TtFkQN0qxQAX3MgoS/+SH8ImV8tcGEaCDBNw0
FaOSK6OKYNIk2iVpecJ4cUKPYIpI7VOkh46mmQvUxrXVV1Em09VNWB41Q5Rim3147XUerkU0L4Az
aaCBLu+SEpOiD1IYGJHNir5rJwgMhYwpqu/fmELepVgFVLGHzwY7+twXLPk581HgMlb69DbpZM9z
dOyG6DFAXhcuioVHW6kKzotyabRvqL7N3f2GtPF82HutoP3Z2wjfRvYKVXD1ZO4DpUI6wI7+2DM2
li610aB7aWWkxmweDWC1KDSLnDlHMLNtn6DncSzQkUeJFnffddLFO0xxNOVTUUYA+56dUYkXaDTt
2sVuxSVUSx1Kre9b7pQTHl7eWQceCywjz2flFxHh3ebinQPfgoCKte08UCNGTnQXBN5IF9uZZ2yy
UcuxVEru057Cc0lnPendWLCi1PSWLuqVwa0FEsutjH3h2Q4R1aBFsqUlnJB0taCnKpJWkE8rqrL2
9jHeUI7Qi7uL7MIP9h8i4O9W42dD2cZuY+CEnf/k+mFcdGaNIMAg+iXPhdnaRlQT6xOZLuRu8mg4
CFNWTn/+ZryQry5IkOOcDqZzGnXjTryPKTK7Ac16Aa7KPfDFGefR69hNvXNnYLV+jSYOnTKv31Ry
vR8wwFzrzKUODx4GQJt8yADQXG0L6uPoxK/gKogxAOJMnrTvWMHuWHDea9XNldPEiGrwRlrqJmVk
WHmsbMWuKXLTprvxDOAY2sYpT6NVF1Gq80a3KDg5lrLKyJwjmAsPs4pRwOtEMveTj/WC7oePnnjI
Hry21v5XnI8AW0qLCvZ2UQG2o0xNO7VYjZFdjEkKc321agKOKHCt370vdoa0dmfmM55qCfV3rfN6
tRUiRVaYUiZRAlmEh+zwJVQruJZZFLZiASicf3o38IYj/EJmCjKingWJn28tDeL4V1KrhvoPW3p2
qCv9I3q4YDL15eoWMKm4pEj0YOciFsEMxp9PLMv5O9RizJzJFBv3/pCtr7KDlRUjKBUuWf99XY6z
36LadRUeWNv2KKG7uMcAjqvg268qBRFA+4Fl9PwXprwouWJum1oRuzI3aFH88DNHvhl5+UxoaWya
YppggrkeP9bmvK6unygKuRZ1B4lGpiGUU2lBJ60vn1lJYDmHNggrcglUSUXU+SiB4kYBPk9mUlpd
YyUJ/SZKjcS4Q7HyXizTYMpXAIK++rVnONBC5y3PN+5r+kXE0S0bPBu2mon1LA4pIpedoIotvTHJ
Fx0rsnFhZ35Ofbb8Qtx7pCJYtVqoGx4Q759hCpVnec9DcwbAId7XRV6c1/OJCvX/H6qilf+IrSD2
cHvZXdotlcpdrmElULiPanEDqQzw0WB7sOZT/wGe+vZ+cD5BEzNvtwsna3garDPduf7u5lUCvHc5
pUDSx2OEiH4z5hHquSE215Sx5yeYobMao+aUpINzRDuXwSHTD8SxEzUoYO+OiTEglj4pCPg2EOIT
41ZwcmvgdaBNJhT5MJp4TimVt3PGwjR4om9LLtSkzvP/WOedS7MfKMTcc8bNEy1Ir/csuO+rBh3h
OImIaJSVtjpnP27O+SaSzHVII4Y74t+3GUEUY3in9T/p75FlY7jvCRTFWjtgWeNrop2co0s3qeyH
jVDAxB88TVv06hKoklfKfl41SVqI+FgMz/0vWEUgfa8CMKXnJsGDb+DMUNWXCJMYzCHCGp3M76oZ
vP4ygIPtf6wMXXIEx7MH050GnfqkIAKdUsosrTfSae7x+PJ8qb6zV2cj3r2wbqInTE5NlyFei2vU
X3kMlIFTqjiN22S94wZ6Yu69k7xP7asZvKv5SSIyba5RthET4ODaMk/nyfaS5UXGoQ59ywHFxp2k
dt7hpFj2hQgK8xXIBlwtfW1XGmEkhTyckfQkA94AEp5nypN4MDLuhw3svK7GPzprhFcGTxjRnGSP
h2X3t0BOUKg78Mt/8xUKN7h/sdIdpP7HtBX0YV9cfagPjKkny4PEfDka5jW5YXcu0TyP1djahVUJ
TJPF9NsGkFj+RJ6ZgwuUXVoG42QZB54cpVG6wRsUnMVoh9zSzt4L9bYNrxV290gXsM02Mc8ldTzp
ycY4XfdiUtHaugTARL9VaZHGEaeH3RtQahyFc6M7sGA/iRCENlO7QWWXQU1jyMjmAjiEeOO7r4H+
nfD3w5CFY5lcvsQ4Z3vhZEyQA+yVeLqL4LYUG8+BneePJddZ7eg1j14+vJNR1zeo3fz9tguDujWb
D0lU/xxpfma4vswkP1z9UjjBQXNxpzN6+0XGy4mMYqXoszGSGdPxtV4NV3GR6nu2UUPPW3ogmhgy
GqMmw3iJNSeONMHXW+RtGG7suxvLiZfSMDXWLH2huPAB5DF8HEQhIqRvFMLXRpsKpF9AublQJIJ9
MXYzTfPeXjl1n4/kxd6xIeDpZ6ghuPapPm5DamhW+ngCbnFzsRGK2IlAgeQ4wwWNIfsyQ9/Zu27I
QrvlILMWtPSSk5SklGASX/puhPfJhGB/eP/8yNus6EwxSPZc25GudkbF4kt/IBzYu4bTSg3ET/tU
gzRY8sQH+B1IT6vJCUvtUFmeZ3ijhxS6mpZGRvK/BXbZlX7ITdY11LXu5R7Ps91sMCoUZW4ZC5MY
NW7LelApaA8LfbPTsk+5DYdwxa1t2Fu61647BzmoCWrCgLFRjXHC2OcsmgikumtNjeXLyEZq0nFO
Xb1u3Cq2CMOWaY2wXitJ3R2gDshgV5OgElgXLW9YI6/TbFIZ2qGwwiBwGn2lvRE3X+VTRNYxdf/V
Hu7aY8qJ8EjQ2vVUd90uJlAQ3pqGINspxnup64mtd9FVib89tWZY/PLatjlFkpHzjIvgqRs+vCcf
FPpAv3O3O8Y3JPLtHthwTL/9m2CyE7nKVmajaPSNPZaPN+EW2dwEGJaSTHD/eDOwVVkyeFCkNeez
cpHizxQ5uqcfPSxzMMuFYjQLZPEcaYv866ofYjlfqO7IE3Ueo/CzcyNHZOCX3MEEG05U3k1yiAom
WSKR6+vM3ei/GlXljtw3ZZG6xNDixVggUppF2//YcDPDADcbnGZrh6u3ZahlnLFMIBBHqetxoqJH
z4ae5lpdpXlx71Yban+KrV913GzsmtH8vUT+PU1EqsyYD7gvzAp4UsorhW08dFgl6sIjAE7a6t9a
uSisxPwO7hmxlfx8vTCicBLJpRqpxb6MQlTEIfH8OPlBsXMyWpFFJDC+6PoMto7td2gZuoDQs1aA
UXEjdUCQVe2mFPMINs3pNd1frtRiqkewNpYlkbMzwbz8h/ONPdK+ntH5QFDB2CXGx0IdMtLMP4hE
FaoUAuqF/B/IIFH1aIgw4AurCAojUaahISuNRvZBiBJfhKV8NNvPHnW48w/kXnVesJH1CH1B2Pgd
SM6GQyqSuS53EjUg3nS1BGzdgiljHQzH9LfZISxd+RjG9HnNZf1c7x3sqt+BHZt84p7fd524eeuW
cDKR2zimYge0H7UIx8jgy1aroq3WEIqkEk79y8rgkB9bbXUcoUqzxr4PCWxy1gm2jMG9eTCcokcP
iN2ULvwbyy294yTZkA3JMf9eNUFk43aFb6VLNNzfcLzkyKybHEyRaj/EQG41+3kcylZAn2QUp4v7
4Hf0iR7+RzcVzr1o/SqLjB5QiOW79wC7X8IH3bDJt2zUgSJ9caJwkEdGuM07DnZEgOt3FMtQhrqh
lQkpqYDBDXZAVoLQxSgIZSKocOR3u2fLfRTFxbU//YlXJVdnrrQmJm1bzDcX8pE/ccBNQThzUlFj
1NIc4+5ia53OHVpwomIJ5kQNysH+7I8NU3MNjXkzAqjl/ec232B6pqiZqno9moJgWKHCt5Hq66hl
9yI9D82RXUPcPeVsF4qABWUYncXl4Vg77a1qV/zrRUKbTBzesHhMhhLHqq4JXjJIqKvv5YQl+I+D
YcvUaYIyzel6ZKuEXZs6XebvQE9tLpW6Z64UZbPqXPhAxNSS7tBcXWotXxx7zecVBioudJLaVvNQ
PVHOYHK35Tc6jJlLRaB0Qm/1jn2niaQ9oep/cpAlsiEV0X2+nkVa2NkHENSL3PAXhkpwVdB5WoFe
9RVE4QuAvrCbUS0HrS8TlbrkBd7Ahki/FIiElQeZZdWKolVJn4V/l1Tg5c8r6qLkUxcb6WFNLa65
51RYj7uKXZbi4uII7XVrkQuieggmz5v78nAL+5hkIxlR8YHxBZUI05jjrMiUJd1DRT0NNPYCGXIa
acoE6ozvmbDivz4MU5CvEwo6INynKSz7q3A8TVVmoPnRlsOtbnxd0MJxlnEgmPFgkFdnaKvMTrj9
zDFoTfIkjRml8kXSA5hd/Y4hxj//zo7wJQ2ym96z0CjFieFC0TJeFwwuPEpFbiWudMBZcaHU6HFS
NGT82idP5xbg+7eHMAr7lkwhU3S0yLn2DfCb7UIwWCLAkhmCRAM9g8AAhQjsvSwi7UJeXrWCYD6l
hoOWYylLbdu6E35O/xcKm3PWb+iCowiOqciLfh5mpObjpZH5848+ATR5kg2Z3eEQJCxxca+GWfEe
N/KaB4DmlMxdbtSThMltJLvaCPEOF+CacRAYtKWOgUaCv0Vk8vD+S9iB53JYpLagg1y9oJhGrZ9F
uVRdMHvz0RYhp0NrluA6jXCkzG8PSAXvkMB+o53xY7h43l4eyOY41zZsieteCYjVU5QODeEADfKy
WRVLfHTmuw1xjtNF1vQngWV6WEZYZAHXHal/KCG1Ddw4nOJ9jxKSeGowkiBhPRf01RDplBEROp7W
JTFzxTk9H4RRBnRJS/RQ2Lj/XYldkcXHnybIQuA7k/VgJxIlhSPabPB5x9pYDSDaBJ2P+hK8ewAV
F4EUPLYSWk7zNdGWPHbJSD033XRKzFIA//Dw57RFE+9sIS8+T4T8lzrwL31kiI6yCPbWsZwSaOYf
PSopreF/6x6VBy6TjVrn8uEl9TL05sy9UXG2tldpIvj9joGZmpzPJ1HLqsjvRTmc5k1WZipt/s86
yyTrMu9bB2fozb9ugFcsF/wxhN9V0yTXFn9fm0jc/DWCtFJZ+xjzwtJkFtINQxZUGFLnMXlAPsh5
XBVcn5RwBSUIz8NWC7vKs5DdpnVMVoTI70vNZTQISrhp/8k1V+8CRPhOFyp05hCBQtd8jFKXUn4g
3nU3L634P9fyOpFQgYi4d8qOH/ajhqPqmaHKg1uoqbMxnPvokok2SyKPZ5rekPvs+pKZO0UcHuZR
J9oJxqp5uPOyM2rdHVX8DMCGOW/0siXewu4ZH94uYJBUc75Heh1NLhJA3akipR4/rrqNQZuwLfJd
a/fBCsgoMFG6MbZPjLUC2iDEph9QhoQtp0qe8OCYQKSm0zRdiKI4vdDYfg6rkBy99e4fzIdGDDNj
fhmcKc+OjuxjaUdlBu/ko5FiI1a+sk5/fgPpWJPlLY2KjGvG+rw+u9g1b5P4HaO4qTzuiKtDLAS4
E1OIqDehQZ6g1Sp1qyj3DYlh5uUcrb/6X71w16BK1FnRjjo/3stsz0hwKZ+81fU1qzqSVmFqYaCg
mP3VU+3X0QHN0GX9PXsH7oZlENwyL1KisDKu1SFVQLYa2zCI++uoybMlwNqZ004CpsdFfHiNI/O+
dYiHUiNKzWBzRfZxoTvAv4zQ1UadDwtye0WfwkRyqkf5Yqm4AbLLvXBZOXk6TtPyy7L/Enn0fE55
CYbPrgiypAFL984EhBA7IruaNnGmrFPtnvUT41XXw3dLpatn5TCrxlk+gjkV4yPdMCAHeLKTnefZ
5Sq2AVdsY24l491PKXYa6xX1q30cYMkl7E4oi+S0/uklIU3Jzjr8aLAyYykB2hUzhd2IZks4tiVk
bEplauhx4SrcBiQzKN68WgO1GUsYGqKWC9Fzkt26mAt9plPKNx+XulsL2XXNlMmVV0v8IlLwpQAd
ee0hSU1S/ZmN1aMOoMbPmPBRSvaP/nndgW7RXutPRaWnthqZcsK4u7HT/J8d/uMqNAa1jMrT/XlV
r3EK4nQIsI8EuCCcUdftqgshep5K35eKknJpdMqJ6rA8Nt3Ee8fLsWf7FrxqkUrEfSBSvijYCTY3
sXIOXLtZfOWNSpk60nLiCF3pm62XrHNBMPBu7u614Hey0r5r8dWtZkyqjpFS9xeO+2YTGrTSc9CH
U90QaxnUld+q9Ep+iy52N/z5RDA9IrhmmCDaDIpiPJiL1QtmOe2ZkMr3ybiZ2oVWHGjjE3Zal/rm
cUpyHYrzwf4U60EO3PEfLSfiIy3p4w3NFGnW2rMr0hGbSu3wSKA8rT2JqZoDEJdANapJz7PRMiJ9
I9z/vjbI71vZ5S4syaYQoHH0RDAE2irrrJOvcxeTd/fZvg9wZpM0cHfQGajxl3Gi+k2A3S9YNAVL
ST1mCKZY8lWxBxyeKNdySn4kOITYa2Hlk+G8uLoJFRYWS7YMF4qrsEs4VPQyn+puvsZu5jMx8n0H
13it71+GG3Fq0dc0DTyZECG44sQfC/bV2IALQnIcoYHBM6HW1N87gKfa0i5fW+OAfKJDcXn3Wkis
63FTgr8AxrQlx3ykQaihR+efLqer6Vmo3Owm3C5dykS6gjkkkVKurg8c5yJQkFuODrVnb32T9k3X
Zx0VRrC8iCBa5skW0Tb3kCUToHwqJt6vAn3KUNHD+4xeTUJYzGp29iiHx38dCXYlOawbnbIvQZxM
4QVO5/GcVeKjrcH61NfT3kdifVWUh+RP4zjA2emB5u3kODrABeQCWXwbmMH0oDxxhyez1JCQvF30
QPOyhuUAYN/kW/xsxJfQxt++9ChZ5xFxSTQQ4Rp3Jjm21nJItjWC5o8JJdlu9FRwp0TE70rgRPdE
yShGwLITeEiV1Iq1a1OQSEU57rymHfpIKvEXxq+MH9xq6SQRZrQrTdeV7ZYhuBYv/KUWDbXegufU
4/gDxInNuWkNGeXFQLtscMT7ESb/g8xO85kh2XdviZwrqZADYPwf0wy0qiDH6yXdpgqcsmwDZDVU
9a+thUzuiuJaPFXdyaj4W2RJdv1pPWZhQwtOUWdEQtwF6gXvbnLFFOSWNMjctwlL4Ooh9bXtnU6m
YdyExQ0vVzP/VOc0rlNWs16vLVWFSEWzJDSc475liGYEYcV3qxPPm5kuJcaKwmpzmsI4p6JGroNw
qUMtxazrQa/SzTdRUhDwQdxLxokuMkrSsE5hHw9TL5kXTnV9ocyUJKPiwgWeuTlzOxAJuj2l5nX8
yhvKG+ykaWetMrlNlmvXSibyfffNFD6OPUQK6b6EDkIqo3UNNwFhk4ZUrGpRlVbO+9oyW18t361x
tGp9SNxWU4XMQwl0OfbH4LXZ6QZr6NdpsIt2gAE0qiLdvj7mWL3qeFjgq2mGQ//JBFSUXjFsvUtQ
YfGmzCPMBgLbCERC0HHsOoC8lFQQTIcPEuyHPG3Shs7v5JGhi6t2Na2MdMFHkrrfjL0BV2IwfQXi
3sEz3DWvX0MuMHKOW3MHtUkJkyPAT+L7FhOOIhsmqRagAau7mtrdBJOdsM36k4Tk0LOeQN6T5xTG
p3pAMtafemdJHsq/TJT5mzpwBz9r5nIairWGWBmO/Sui3VMQdTO2hD0hyj/9O35Xsq0ECg0U1gtw
n1M0PGGAlOEw2wxYxUFbIG8abVYaiFRja96JiLGI2KlJV1DpxonXAYHlzHAqmplB6LYJubCQNrt7
/CfFpArYriUv7aJo/7LDa1R74Jnht3stLSdiMr+EIFkYoacJaLrxscf0JSSjD4Wt0yLxzqGFcL+I
n3S6mi61yw0C17XPNy3CxY+gojh4dsGm7oVvKyi3GCUKS2Z9bg9yBMazzLE7fpnu7W3OW6GQxoKI
rR9OSZ0lHw6hRts66fh0mGw2ABaorW7PKOvdgj6/kaQcdOfMQ9XNsOFKrlzJqPGzq4d2+fB+Je1h
+E/x5sBXvXpDzRi1PidD0L10X5ltjpHYmcIngDGoq6d+NJKY9WE7XZFbFkXxk0iLxABSTWYWYdm1
kUrjd93QTxwPyrtBRGg8JZ8zJ32cTTOl2qHPevdRiPH5+yZPTqjPC1Pj7Ly4ZvgW9VdrBbytt0bX
Ni1FBBxpOxFlWaVxpZLCOomk73zhDXBJdM7FgSy8EkDbIbvK05NRI+360qnbs+0MvxTtff8Vvyqb
ZDu656eoePAMDW/aQ7A/qOocHEaxRnaePb4jrp4Ms5cQ5RraIHeJv7yLtnPrhJf9ASmLdt6a5owj
P/maBkWqA9m0/Ic2BMyI+BdseynZBc5ag67jZYE0TKs2lezHqMOEW9FZYpVxJawZf+OqUSNN3Gyl
f1XUdywmvJYbyjPndUUjKiALuQgLx16LK03Kh/T8D8zEijQZm5u6YRvdx933MXt0amoxKBC7T7al
TsZorWMRR5b2Ra0IfnWRrVHe7UMDhIBWEe8e4tHchcd6CRgwWkhlH4HvkzIx6Ioj+8HtoZQKZ2rJ
cPb45zkT4hykCFMZhnEafUW0PFOctvo0zyyMWBUQrMN0tAEd1UYbx0K3lAlMIxsPMscZlsloYxb3
Vh5H8S8EHnrzzcSrmycrE/hxSlfEv539+g6vOVexMp7zTtabldMPxiqhxZQMJZwxnX1axhxFUwT9
q7yV6Gmnm4dpvL0cLH2D9CilInrJ2sETrio6r5k5PNMK+Tw16/QBMLsCXMC3jU+oVKwki6f7LkfX
Qpcr+DHNpyyzulB7rxsvxLjJ2ylMut0NlrDfNpSel6HejS0fh8GkLHu4BP4YlZPvBkJfySrTqtxS
1IsiWK3tfhF8bmQU8cEeHS7GAENRhrwv+UfawdkXsgXyUZjyOYGAxbGlZHJKBBePT5OoaUQUuztt
GbJGpEKL//HOqQ0foeKUqVFZ41GCBi0ro68plQEnBULt9RpnB/SYd/B4p9eY+Lyk1oeKnFF5i3Lq
CSAtNCCLzunO5jpEJB4yCGutREUe5ijE8OWCX6fL6Eywp4Cjzax0PQmHNSHi7mYK1Tz6AnYGymjl
oJt181UMTfRwlRajgNtH9lFWzoZa/JZbhnlNCS1huBZA2NXifbHqmid3k9Jue7rERgIAwrIFQwZQ
970B7k0HT4rOxttJOiVFFEo9ao3wzLQgYchvGA4/FJKzIS1APA+8X0II3jMGrYYwMV3xhyn2RIZX
SV0eUWoC0O+K3iwD7cUloa9THj1RU+BLNLa8qIfzOTXkCT40wUn6k3BgZxdKOLpNiwAVd1J54YZN
7PU/V6nUnu+k+O4HWEmBVnXXgekjnnS+9pBA3ZlUCjwTfWPRCBjoE7RMYA0wSKChPc6NyRYfxE83
FHGtd+pmVl1leQIcIL+d10es8m5TfG78Cl5LNFLhCnkAGuNkdtFLXv3pVMwDBcPNgYtrmU+CjLha
TvebfnSHS9dBwIKXz3GHXd1AVWRpVH/BDlxFNp3TpZN5LoMiPl/bVqcM/uRUGdYwsZQ3t6SItHiL
tRJRoiQaFdKv1yYxsj8b5P5XHkyiLE9pfLuTd1pC2lUU6wMkSqv9qH5/gbhnhrDxTfXPBWPttcW5
Q/0Fyt6A/6fIbEZ0pQ6A+NNL0988jg7Vg/gLtY+OXVDGYR+P71nihHOOfToSkqmSMWgttoQ1shdh
H19N74qM/iFDCSs10E2LZUCOFFMqJsjZIPyskC/8/8tTZz8LsDNtuXu45kG/2vcWObDSfShcXssQ
Y2HQZJ9lhk33gk0R+JkrlDPAgeFPi0iHaq5fD4CDHFD1mmQBA5FyeQmXbUS5yBKgfw8FPNCicac2
oyc2IU6A6JuKTa6Lxf1SG9r6FFIZc+guVwkgKdUH+/tXbkkDASByBPg3QDGaEmhQIMVDEw6ionQp
YmW4kGfokl5IJkTjDAwX/JQ5zhuAVlUam8siN9WBAtAKGxZZTCW4uyjRnvOraacUNOHSwNru5GJl
H8d2B3YgsZ3u/GN+hgqkwu7b5SPguCSH0CwfgnN4RwNPs46NVS4O/O488x8bWlaiv2imrnXjYua9
kRUkoSJU/rKgFNqS6rV7NBSDMezTAtEblotChLl7xZnD+BRlfatxajL+CeA0JX4qqtylya0JAPmY
JXnRMPVJtb8EXvdeKMq/ejX90n/J3E09BZrVl52wN67lzfG5RPrZe9IKxN/6RytVFwtPNIWb8nNP
0/L1JNyYpG8uRqsbCnsbagrGc9ZvXZIgUrrVR5JPJJPhYnKcI9t7lDJJ7hH9qpRI2+H73BlT7EvV
4m0wE+ixlO4wWNvkzIXXZMJya0dFbQHayexOdPxc9ksFmTT7TJab3LrDg3OCDLlB+dIr4AqQDqjU
VbfdNDOpBStzx+5GC4gbw6ZO2s+Hvggb8y5h2Wf7We2YDnJX+sI8TvLnhL/ziiSHDWm+ZA5F7+fg
LuWETnVN2yxsU9kywhubMMAXOl+0i0YCWUIweDlolU7PzkpZEujdzKfhyyow3xVV8W7JrQx3mujr
dlKxt2hKMNCjJKa1vz4ZC79T6IwyQm/+/DYGEv6Wehpz2ny1lY1bA1stIOr/LA+mCzQ7zAbJISpF
r2l7kvhJnTaYtBakEV5coEu7yetnx6YJWplAN3ayR4nbjmYvnR85DXEw7JaFPYFz+FOOOtqqsstN
FnfAP8kHu9qXNqyUlAU/g7K/+2aZlgimHOOYxqrUKZF6Te1t4YUhP64Mwgble62Wpr8yc1Cf2jR4
F4V7fCI1zM15Cu4IJLJ7h4kdD+LjowtfQ2WaXBzihY8p+twv4RykSvoxD5qI2imwzQtafYHl+pRn
Gi0fcDKi3Xpgw6CD1hx4ft17bnnWi/0bhTKSkkLRnNiR3fdwmUhJXPEqR5p78eJZfagG7GqVVhVF
Ai2vqHBn+E6lkcnWQx/9GhKXjRSXyt+oYTNAOxwJEkV7fjUgvBtOGHJx0fZDWjdHdkpJ/yZ6mHfo
/FEtNRTb8e4CrALDyLpGhZIUoQY2xMDP1V0RMTLQArgfzLtI56tn2BGZ3cun8I+tieazsbbQhHnq
FOPmCJpGBS/GbleeJw/SFpFBaPODHdAK7UF2nM2o4jIq3vZLoQ8/T8RaBwHGMUsdHY58dfTFJkcL
vnSQSxaDpxA1d/2cW1wURQ1qyS5zm6S4SePzaV+tod9WwGbeSWu2iY63sVqvo9Wcclj9dL+lmT9r
e0vk7BchPaxEtYqW/XDkc/KbTj1AKF4HGwpUzC9IrzyV+nbjzhpCbAxFSm8KXov8zYAAUwXNRtrt
dHJFx9vVfBriaU3wyEzAgs+i8ik9kXcxeLJOqiDMtYTunplYc7dTD9aRGghdvE4REjWQJbd5Vsm9
6RWztV1gIFfem/94YpRY3PnnXFnCUeTHPqHQjDE94+wDxwlbE3RV0NR8QMGcwBPZp+DWYX9TJlIp
nsts4/7y5zSShRpw8Cwy4tnMpp2wfxp787tuqowS7kCbsI/b60cjigOkHnI4QPXNxU00tlc00jsm
G2r6sfY6LHX+3J9HOKbHpGnJkrr61IzRK00yaIMtgp77g/muI5uOo98sFCUBNZxqtFI5zt8z9VIH
2UU71fwsyNnjPgiH5pwJ9CrNRZ73D63USR+C0ViY51axKWc2LKm1wMVJoJvjbgTxvaQTo/3tPOHB
FokoHb4NLSe3Hi+8kZKn7EH2NcEMecuKLHOW60tp0O+thwbL1pE34kk9Ze2rtI24NqcRxdMHHDtJ
QeSDeauH1LZL8S+0sMIUwTumWLegduXwpnebJdDjlntzsE0s6RRsIpxFO6DvbYSgt8K9WRoNDEJD
/bkeTqS+pBTl3Ibhavx33eMYLnRlxfDqgkdeNhLBOAXdlRC7aeszAtzWJrEmzLHMQ14+nJ7BE0gW
w69eSG7KughtLTLk6YoyUzJbf+P86GkAWFN6rYIdHsCkhSy7ZcAwexq8cl9bPjxoHtNpm/ipiTLl
orndK0qXSq/utp0vUaSAbrS4bugD7J166j7zWV/WVTPTCRIhiV9Wlw9ws0z5hwD7A5xtkma22/Q7
bZzH5PKB9H344hleeGnVjGKLJ6bRb16tzsBc1PJZzGJ2qmuEjkuc3C7hmrFjLic2TFeRRTjj7X1M
nW9sUuqOZyWaGD2u+Fn2UcAuTDuPJ19xiSfFvB0JSoEUVx0HQ9wQmPJxXaUwfXm2v3FFt+vEGxxT
UtfjZUKHPds2VwDI18mvhfaCax8xDJQqGBsbxsOScKU08/aST+V5x72RiklwlyyStIoD6d9TIpw6
FvwU4aN/I8Xl7oB9dHS4f5VUPbjm3xvAQv1UXn3hzg0QnFnED52Ver5F+GZ4YfPiCY5jLasF9XA+
OWoK3Cf5EoFlQl/cBgiQ//Va3ZekTnKdM4Zx2T4rzOtHkBD52g529IKDtHT4hWKAbrhx5G1bJ9Rs
gF5uIM5CwIkEE3HM5Erbv6DxONEDZm+icIU+aXpHOeKD2UxtqdKKxEePexJIzh+1NjIGv9+64uOP
g4AVCUyyv750enbKUkEY4fK4cCy/8rrGV+gYOzwhM2aHVNOdpcK11w2QTlKLc5zCGipR3y5A8f/g
SJZaY9/uKyBJkAl9P5B7nRp+vEot1OEJmirEUKw8gMtWqaHptSYXlkwJcjgEQCMLfKcBG2KO9KBq
/ZXWBeL6scqbvf6HqvoZBd81sELWf76zyDLms8td4Oz5wro2Qs6uCRnc0Xev1VE0OgbQ9m3s7cIw
HWBC2WD0Vw/BMJ0CS8UPwrx+HxroGpggyt5CWiTWHrqYtVV1AgtJHn/n+4cUAkr/MSpUZxfW26lN
uP2/XxjXZXCBUASrpLl3Xg41KZ8XmNTQU6YHRajjsfaUx2Fc5gsvyCiXCu/ktglooL1eUrYMuY73
EeNr4lF7D58MqjzuHVeokFNwJcIWZO50ciIufH3qxzq4882GdWKNAK7ZYKWdhaVvypdxFSGv6338
oWrc1qRBM6vdnjs/XCqb/dSFbBZjyRwPSez2Bluz97BlDwku/mwo2RAlA3h2b9po4/vJz4WX+Kj/
21hIVZtADjDxjKOgdgs8yffuSy8O27cXnRnnYNLcuZBgS/yK1pQFF85cM4tUAuxT/vdBv5Yb28er
hnFWHXCGrOU1D1CpmBqJ8ELc82ynoQcbE1BFAhbz5hTO7vSa9qwLPBCEZPP8Y9HNZ9JOkiAaEWd1
gajdvzQeFP7s2xhtZHNOGl+iRcdOQT73nDB57c+ujlaFR1XV/Qi/HDQ7GW5uxbt+0CJEBSTtNdBQ
NwMADq8p69MXeZjyXo0I8tcFPkeJy4ur/IumNX3l5xogcrJrhbFP/V2xQgxnOdElAJIvKlicjezu
6OYtQ3d9UEQXb4zXqCNsdmnX/540hYbLY9vNEAJAvPi2OvvSup0JjLik8l6Kms6zIQAIHfVCD70c
gG/AEugd5EE3FEO+8mfIY0XTriBZmLu+qzdUmexA8U/8NucJ7V/g4dPTv9SAeOdx12ladYwlszdu
uICMhFoPhA7OuuxBJb3Zs6iBD88SzqOq7+EP0pX7aJ4ASfE3n2MXnIkBkECmu+rb+NNTkquZ3pBm
PvNlEGZjyWtO5K8W0YYD3tQJnE0AhmANHPkQJEavqCoYkyJIWoagT/z4DC0A2CmTKRjnJAnoL9Mv
hXVXHVll8t0huJXKFkbHeRkRUHjvgq4Pq2hmDmrG5enid8ugPEiEu3ZzY4fXdeRpFR+549zPpEWV
tzuAOv8UL+b0q5cAQhsDlb//rcL0/3evc6xXQv72u2veUu4+wguYW2D7NJD4ywf+iv5j1e2snPy7
ftJuVMWwv/qgxRbtce+P95DBg+gMbGl0BhmwR42jkhi9WLBiBHSEkYlJeMMH1o7k5f3CuF8YoSg4
uU6gcgKLrA4IQ/qIjaKPSITat3G429PJOqytwtjNXPCMXBv9RnuCq5ebpBcgqicx2bFCipxyvntI
xOYk6vn5tAWs/9DhGGFJgKVAxh2/VGyFtI8ntjUkr9VcA3DxhHM9pJp5/F++4eXxsW2PRaYWinoC
i9wpw2hHlvlcxSbdYqroikIqkAqWKUFMwefL77q1nHvJ8iR19Qx53eqzI9HxOShg0t1Zjh4g6qUM
UGD/ysC7aQ+nvlpGTStE51++1iGyVGqV77e1sCsGLtirujkPoPGMF5KZdgyLu/dSK/UyA9VxSY4r
duorKGQVhYSko9jLtRcNC2bb8brOR1jyp5PKOs2DI2KYi7xU4quKHtNJHcue2OhcicjkQq3Zm6oh
RN7E1PMRekJWXbz4w6hrxu5+2w20cUHt7UFSPDXQ8AeKQ5f5f7y5wACimpzJtrSCxaiD5Z2UAilx
Qq1nv26a9xskNVB8kk7BoDvE/iNrdg2tXCO5hh4CRe0MjeVuxbMJtdkPxfdZW4Sj5WrcziH8eUXA
4R8ZE9g+tjebx7vdBaAIVw6TTT4450ssl/wsJnQrbU2YH7b4t0AccH90ASgHrOpCLfH5OcLqXvbP
InDS5KOomTmZD6aWka5g0tW+61LsnGYA4qk0/Mz7pi0MjcXmHxowSnhgxmQ/iIj0636ZWqJVjybu
NW2xfH7euPT2AUjNtuFdzhvV9pIK7dVbB5nFdMqFTjCcQUyouiwlO2RrDzcOlvELBdgp5NhqBmFV
wJMejbmNvTqNp03auh9Okh5C3x8jYRbnAp2Olsxn0HXjtob8FONgXVuWzyc/ll5mTW19r+l3zszJ
lIXrwTimEJPE/BQpwcTdxCqZJOKJ+vzZmsSxlhBcTLxdHIGOird7Z006NIFqFPchHiE70LXT03NA
xL43XTXjhEoNHV0yTtTr8dcDj9nQl5KNOX13s3vFBYuGIis6bgw0IJHJ/I0vZ0MVAu/5aTbXXgiq
K+y4dR60ClQpt5QmuvXQLkwZV++5cCKpH0p72Sf0FgTTvGDbBiEbHyxrVSmjmrmws595AfSc6CWM
gHSigXPMFdZjwhgh05ehcBI+f+og2G9y+zbhGZBbcgqvtj619LxWBC9/ZcRXzux9DhvJ5CIJtxqL
3ZNBTKTZ2E1wrDETGE88/tuspLrzCgw7sWTauFrLYMQUAuI8UHO0BPUaCEAdkJ125berDXA6JT+P
9THwHBzcfyMDd0DVpMzO+dTyBllF15HAtt1mCjZahG5k8AmtmBhqq0pZiTo8lHCT1fRQb7mhFOQx
AJZ+Wus39cCa8us/iAtbaob+v791MUMlZhNVbFxw7eNKIxVDCL3e/NzPWyCkdWOpVIs53W3z2NFA
DP2p5HVbKW7fy/GegpwDG0Cw3oBlfq4ghh+W5FPw9cD6+M8Uwe1/MO/LtqE+AsQmhmeZ7lCgcKnN
3rqwI7dgzvFP/zywXzIQG3P3D0jwcklHgPTJNDRBLST6LTXt5UNiQNPGOakOu7StDtu2tCCV+E1S
dVmPtGNZ9qxBegy2BPD9OtIkBbPIaAADHuP1gNRu0Lf+rBvUYtX1pS4iC9JCaKhmMUPG68ynZshj
KoYy3aaBurXq1Q/K+lXnaxHdNJX1wuXNKaRI+Wsba355SXGf/N9B+eFO/JBJo4XyExt6ektIMa8w
5h0I6Ov83/6iwUpHZkvJIkCl7Cv/VjJD+OBnCljVqSlRVFbqD9vOjxLz/y/CV7p7dfAfCBddLsq3
AYAbQF9zDu+nRRf0AxVq074OzFDdWNgKNv/V538kHm2ZAbvPiGTzpCtUmkkqRr27nsn97iG49Ra8
AVKX/Z/SpixjZZgj9UJwPruRIT9uiBms8K6fBeDEXbyqPA0JvY0uuhK+OKZ3m2sdDCGTRF5y70xI
3FaKG7E4VRBkZH+0f4p+n3mthfJXUnUkLeimmCP0b/Vn1Lx1iuySJn2S0INKFCrlKyj1OH04pWkm
4CL1mAAiL5jQllfyth0pklg0JtK1YCnIjLWgGPuCW6GyLYkVF0TDCMYtymBYLev6G8WnTzk0ZrVX
nqehje2Z4HopnjrWZTievjZyozRU7mSbJH6jwaW60vhL4r6h6FYAKcagdxQP9wDpbtFToBfO2D5I
TapJ4tjVH6Dhx/FhH22iTy5YnvXMVwDhRsl7AWiljr57asKyX0nMoY2Qd78sJo+s2jj2LZ8ZEnEz
2Q/GA7rQd5NvRjnu6VV2Nk50XsqSHaGsKGYYu8TwHH86IFlC+SQAGDiVe65D3uc+Dr0GhMrOuOil
OKNO8Hua4He++ybtTgrGaAGYVpYDIYTomMgPvN3oJ5Kw6ZG0wJ9AGR5pgI4oZbas4xfAcI0WRjGQ
HS2MuBkbe1Arf4QXva/j3fLxvKeg4Anwmmeual5V3a4y7D8utwSBK+e7TOFUuVjTX+PvIj/QO9Zh
tqYlotMefU+uYiM1EMY2qyEtAFzc6Iijoa6JUSgmyGBS04t49MZQsNOMcX6aJy17X8WVnlmw0o4I
zOyBmdAy1I/CluT5/P+POZvW3aFCaWsTHdlG20YCjJLoJK1Kn5/wyODVBnzzxnHJn3R1PmrXZ5uk
L/y1JxJwq93xyuDz2lcwYFZxOp+iWIflKGhiLzJs/5Odbm98VmKMxdHdpTgTJ9TOa+xABm0kmbAT
dezjt3q2wR0xJ5sXdYxC7Dop+6su+CF3/q2EqgCc1bY0l2yVMgYVh+JuKnpqw841C1H51uBGRduy
p0SzOx45W1plADpAnHkaYILug1R5jcX05ChqMYFZnimQN6MNTe7qElTV7phZVdsTjV+fkMKRjZ0a
Gl/sa9cZLzm/jSv1kKOPHrDZBBcG1u5hnKp9mqeN8WRcBsUm1Nukpl3ew2cMo7kEazqYHgVLhoNL
salmWQ3mHkmbmaym9bU/IV9Z3qo2SCEPyUew256ZyGd7vch47T6QhthrdXBXeOkXSn5VI9v356lQ
OKuWZWqpOTi8AUZ0EIMohTWfMffzkDUfQgpWu/vWJP2uFxiuj9ef0tinVmjSTRfXGCPGr+otowFW
oIfclLM2JtDpwYjlS5DksC/DGYbAV9govYui+tUTF57htRJnNfGMR+d3ZWb3IqSc4vWyzTzPaYKG
hVlbRY0PuenlKvuF3D+/ARqzlrlWusJYWzkFVNTUjse5U9Bo30pRYMFqYF2iIiu/0yZ3wnvq4Zsy
Jx+FwXtTxxO4M4+zM/T+t1tk0g01ozchv25omFcSuEZ6+09YR0j0sSj4MEBvsvkOkPRECQqh70KC
Az2pogmULPBOAT4b/O28kL4t2dchoxspeBnXggfkS87VmA3Xn5SXXdImJVvWkazh8MMh+l+J1VOD
v0gTL05q0iGYM9gSgPEz0ddU8OkwKqmTYt3B32N3f5Ij0HDeM9AFvXmq4yYVCRIlwzJQKuwTW0R9
rkSoJgLbXV7t196rj4SYUKCr/G3b9X2oDaGrIzdRVi+afXbjf1pH1dyG2NWZ/nG44ApStEtnnRvK
vCDmRlBbiNN9n4UjIyCpL3XDzSbs0pfRsx2bZvrdGC9PfvF0EEuvJXM9mMPcwX2toMMkTCws2xNI
lr2l+ZOiyAcU47NCOgGfwpS0UNcBb7B6qqxd6YlBRmqbK1pZhq+K/JVGIf90/uqHYfh12LA1xSo7
bXPOWw8BjpKeABj6wSrlZPFg7PGfbAaRyMH9QzVPqb/3sY01kz+m4NmRKrDiZqJJ7iqELisdlzHR
38mEdG4SfxU2sUn2CRBGfs3/X++oqOG76Bt5hI4WwbgSVIwzhdU8ZTDe03WkieLmJ3ESe1hioaOH
PPC/Vcct3pwE2PzSfdBEjWLYqTN8XTnMNe1H6D5Znkrub6TQK8DcNSOyMv6iShNvZi4rvMU/8VGT
Mj5nZDgKmQPgjzvc0kS3NBh+eOYn15pvlpyaagGpvvotZgqaAlOq0+7Hcy/rzfGVszcFoEeV4E6m
Iygf693w6N/rN+615C6UGBInW/cvRTt2HFnG4qjRPP4WdzfiGnPK2dnDuOMO/iSaLlHdhhFi60+8
PMTDkZfg6iTJzeH2nB6Zp2tWni4BIfHDjNa23IXf0Mtv6X2OmIA7RnRyRAblAhfYLIvAndDQ66sk
9FcikVb+6Or6E6WBA7eaRFmEALytLOatY+6Sakvv09c2Ck6YsR2XF+dLjnaUB9fhLJHL8jG2YYES
V8XfAX53PjjFGkls2tBp7r0cK9tCZZXSb1oasu+YQ4acNPoFwYu2XDLbROmfqzwyCwB4qm3ElhKr
ZCUFTrLUyNsWz/q7hnkBRgcHGj/MbFntw2TkrvIqcZUkRIC2rP1dBbST9eqyBz9b68oxL/HScH6J
+mgUFYo6apvISO6X3vDWMBR2evdltZTZnuf/r0t8xBkY0RlfRwoylXa10yFnOlxbUbHVLPwyPq0z
r/RttcAS1WW2A8MQT6xKKsEHAMkdS88cph3vh6uRk4w3BYC+8zxTug77bLKoBeppUaKrD7NtdX0q
puyCwhePVHTmbG/qXpAAEJoUV3jo/6VmcP3dp4zhdcw7a6thsdvDiIrxbdhGP3abTazfroZTm48u
mpuHjcV62WcwUolfk+KwEMvChtCWRmEDGBe+y4QFE5e2akqptVB5bqOBKb2V+XjUVYs+0hXfYiXq
DSxuynK3y8uVqeeonZQvWm/atv4aSDprmL8SUwA6M+c7zJzAePvhnRvZRM2BerfHz0fY6X7USTCw
Pa6jTi+7WMa5940B34tyBIGJGouvjYDPkEtl9z5SFHLDDHEHCCLx6EeZmX7C7y2K7qGZ/H6XmYPl
Sq0QArtIYNChIBduy+tdUHlzDrWvFG2f5qoghMRY70LsqC7zS1ohjGXCfMA2oP5hEsJ5PJg7otzc
ofTSIx8eFSoCs9np0sona0xiBzDa3MLnjtwcrlHclYKxqXmvaMV1D2wZAb7UCw+OoNtMnonW1Jvz
hzn3WqCE8NsMvkezSpyukHtx4+GncLruUbFL4mZSVdcG+6rUcswE8shVIbz7i4swl90kow4qgKwN
WBH8d8pzxy8GUOFKbqQNDRiP9BQA/fyiXblfiLpud7bEQQCREyWxNFotwd649KQUXcjfrajOKlYc
WVZG2MX/7y4vhY7OW+CgiPG0Sa2u/FUbFzX24eUuJAH9uRdjAmybTqIcDJJN1IKFyejT63iBGK4M
15/bm4H4PPon+qBA0CNC71+D2aEewsuOhPzYD3t6PgtZswuH00VWPrz0gyCSa2YxrFtbXI/Wovzj
qhwYUNHN16u9l/1X20l1YF8JDgKQVmvMotgiXca7ZMrLzTq4g6Rgq7e1PBBkJi59lUcIX6cA92B7
y/F78rd0wZUe9hdiP7FciPyx6F5gw8eWMmsUbCzOwoBeeoxfPU7efhkRBvkf2an4YaCO3EwLIZGH
dQ4F+HOwk1L1iGfEW7SQIOUAG1F71DvLA3SrRqFo6oVleO8gQqZjxIu3m6RFyOLm2krX6k3ouTWW
K3KELb+vODVu1TG19sJplUksIk/PA2V53EgxY6tNjJFd2OlAerNdRaRqB/tN3mMm0ckERnb5w3bD
zPF671rKjOYpmKYyzDe9IUOu/lHI6o8iNup79gLZX36wDNn89kPP2+T5cTSAG0lxKwP5d40oT65b
DHJ8lMS6FgAPoV3q4CiJv1P3DxhHDgHXii4uXEzY6ZGVoIdpFTcwKHT2kyKrNPhBDdYKpTSzGx65
KDQrXbqK2Ff9o2tO+KK6ifjZ6+95rzYmk3slMTQAMq86DzeeCGXhmqHE7wavj0mrLHsq5sjjyzE9
u/wCbR5gOoopW5r1GETISL9YeEk7xtVjMbAVz2G1vFqEEYPHKrKNRP2BpQAOf+w6OR2eTzMLx9vZ
4zgWIrArZ1truewK+SqhvHOHl8527WTka20tL5SL7wlv8vyzd65NLMxSfEdeH2yOfmriop+TaUbW
OhjM1vrLLKVgvYwKHYdrNpYN9lj+2nrg5Iq3jv55KCnVYEdpfz2svIMCOWPHaCh5mE5jlg0D4S3G
Oj92ldOyDcPmZ3TYXSAtqUDyU4sy5dlRHeD12HGYkfA8bWS1/Dr+1vrTW+lZJ1br9wJvkiDgpI+W
rlVF3zxpa0SVC2gZoHDOLn8pO2oxGJo2cZ6klNXtFCYM9AgvNW3XGRN0kAQizdCfnxaBqenqBFVv
Buz/jgdsOeEU/NLIRbhPqq0n1KKOPCE+MfozfC8sCzpJUOvC9XMqdm5ynucF01Sy2bV8bBWHB4yW
D22XMwO0Zi7i6ssUzZ5nzkC8ClGK0KUkF/d5JrTcx5R9zRvPuE8qYZ9dLe1Lkd7PxKQ3OJXZY3dB
6tVwkplyJPBi8SzbBO6GV1tdjtwu7625ihK3b2L/7T4s3JqzPkMIV4bJqaNLXr8HpsrmVPNCOxIY
T+7egOzAZB8ipIfwd+lKlSmpvD6RJjMCcLseDII9djAet/A2/AYIt3OCS2x1eRBW/iHxIY4bQiX3
CcEJC6uV0OrFvo4pnGtDdix5hifl20gc+T8OkY4hM/Z3XW0/OxdLaDPBAA4iKQTEUGAw/Sgkm7lH
JfQDkZmlJqne0YBIqHmJKoeGuGm5i/pMRfmYusdv/B/4PSHA7WlW07rJuCMTG4+wDso/+aeJlNOG
F0QeZSvK7+nNULVwP8ZA7vX9GuT0CGbSL41lsr6Ik+iJsEeD4sXR8MHFrqeqBl4XpR7QYim8ohsn
cbs/YHe4+WWoBMR8gPuyxKU6ujHSmxe7nR0zyKUtBSIomj0AiyIe2EH8RDcfNNQqdddn6nJAWNnO
++xSkMijrlLoeC9q0QqB9Pwn0Wb+pAzwQtRBSt8hs8vhiC6vDl9iCc/qrtiF4S91/Exvww7msA6M
PshLmgtZADncrNbxfe6WNRU9PbG+yoV+EIF7Tjqe0Oa/TSORSdN6uGgFT/rMuZtF5vaQqmV32qQ5
2grvaiNvOwHSlFomXgQ7GXhAT+PxCpPlUaC4UiEDIJx3WHwp9Zu29bmlo6XFf5va2yaXZzMAXrDI
1jLGMEQA/ChqGs6776tzuqnUwIcSO5VH2pTqhuNhcGDstHh+hImEVMro2wzzHYoEr/6Kug0tg0s1
aEqrmynrbyK7RibDfhHDundvfSkNpA6ZT8kCLD0Vt319GmRWjxFDZRwKtUP8IJndf9ZOJtnTa16k
QOcMg4tJAEZLCIy3e8pBbj/sekChKhfvG8CXx63oKk7/KNcHBrIl1cFukTXQ4QE4oCBU+1ELnZYc
1uf0SGWS4u4Q2OaUYcdFtXznCl/9YDmyZqOK80Yo2xtdBBngWe1PWs8LBHHTbNUJuFj8LJnaEg3+
EFqmA/ym743jQ1GxY2GgV5YXZKwnE6DoKI0ERg7jjEj2wz/J39vkar5cYm9MQKrzLu/no1A3zHkm
8Ae2O5tmW0Hgo4oBLVURVdlPU8hswT8Ad2sFmSp41nX3TKwSBpoNyS5pm6pGdcLecLAQHdOiGNSJ
J8ll6+qKrYPqq5lHhAbXP0dTHJKaLa0jYdirOSzyDxdi14CFrbKovF2T4qq0QT2jYtVV4Z8ZeIfz
jado6wR8+UaxaH2eeiMGkQSz7uer3TU8w++qw3d57AJ9zKfyvjnDJwL7vNL9XqHlS0O95PxANgen
qzJKxusWshgcdnyTiL+52CrIs9M8fu/oPhp/eBy+53jLHi6FIY5SCnXAEBa1y7vYjn1r0dhfeGc3
ukjtrArpfgF3s0mONl3ISLG07eurBW4y9wD7wUbpH9FYmgKNRjpfEpvOtAt9OW2OG9LzMFQ2semI
adjaVqQbi6XMQsLuHnc59aVkGqCF3yeM73eszofs0PoIBihBfViUrRdsxA3G3JnhPKKocKUQ2uxt
GV48LMsm62MYidfmk47o6ZhnpYfjz5hbWTnqwaiIeTKdXvoky6NulI91DDzLWPJuCyIytyscJKi1
uQk3oGp2xxD6jEZgcGwsCr6Uo+/p9gnzRHG7WXXEqNq1yj7/Ja0AcluGqK/DZ6hQLfsYIQLI+FPD
PChWyOCFTsnRnH5sS2EBu54ED1fO34Uaih4FFIP83BQaJTW2Hv+1omlH/rt7Jm+lGhIPkiU2hnVB
2oyOGdtHfrqT/mlErUcV+Dt6BnspLnKOqpPfMM+G9vS5ZmP+kX+0tZGYKPq2zcgiRlmlVzXg4ksp
9CDs2cEA7SuPeHLwAWhv9kYQDC9yTXKLW8L98NqaGzGBjME8xXOPJflwdY2IGDjeoB8tN6GfJU5F
w5b3Bbtku57xUOY0kPuz784jxGSE2u3vsTmdMRKCg3nIUJObK1oOqK1cNY9xr9pV2xzi+G/whDpe
iuNGisAyPtmukIxYPihhOE4xyrZUFPqkCVJAZa7vssxmx804NM0Ye1g0G1Y4AWI6JwPObNIgRtuX
RUteepxyUXzvCtjgtjQBBsBbbb6oxHXbiVyQ+oOisPbgfqhz5zZZN3rP6Cq0oEu3PVh6qE2lZCIb
vi3GD/2ZPOSOZ3vdBGHyTlkQi544NqN8o07+H3qPF/FVvVXKzdQmsHFaYqhR3aVADLSG3W11HiD5
5/aI3vGfYYyX853kSM+vNXESlpqz04DRPLuzsZ3KmjPc2Vz/HwflBWmrpRAPIfafpNt5bf6qP8t1
4FKDIECgeIAJOaV5C11/Y/jsdcFeHfIkRxDoje2vjuoaDO/xe9LO2iHLHpcmE5zkjQ3TwJe5844N
ClE2lCqHJr3PIrkWRC4cEaeHVTsYaGT25Hj6OCg2xg0KO1fqcpBJrQC9Ks65gUZ0KNfkmDLDujBF
WDVeG0YTi3na9MiSz2WzN89yfGZEEtc+KSoGzGNT1tiguWORNXzrOC0MN77p37GpETpom+MHQIgh
wc6l/Tfqn9NxY3q/wcpUGNNtq6mwzcSOQ+3HxgnvoyBhnwoO/qI9z8BMA6A8BQf87yM8VyNwxcrb
7RYwKXV+U++KF99wp0D3tFjGeai/UV3pxpq4nKmN6VfaJqK9FR7IvUfTgJAuZBljvnUFxp+TwbqP
ZzRUF7UuFP2GZ8l22EJ81OJyarPiiFXmgcuuC7htsFa3a1Skjj9mqwd4gVAiPm9z/FzMZZILmE7Y
Q5cxUq6h2iwlCRNzxM86/PbQImdZW34MaWmIKOoyS3G1vnKCncSylQvr+yH9k9hL7LvIn+V2JU/l
B6uRK3oprpSCXoiWzwHAh3Sw0fcR/OPQiZi+W0NKaUcGiTZEhhEyNEPgZtBfXmE+jARFk1tu3Pf3
gb9Ja0a6YZY/npUyWACTORUkcdMvl5TrB2u0QG1MDRjoIE9b3TN9IRc48yXm+h9myhANxpE5cRtt
g5swgr5e6+wWS56xQIqITyKMePlYfPsczp97nwWaE8bGoAg1MVuQWqGiBiuH/whmMprHnhG1CD2V
174hRCJpduutR+t8GiqY+oYAsfQTgoK6fSUQ1TULUgq4NL4UkyW/qxp063VIIFOyhyNYiSpzTOv9
GNOLNx67FjF37jVIAClVJsxCcpUBlTLinrNRo+doqlAp3ykdYYwDuGXXMTO7dyDHmoWvo/7dq2Lq
jXsaG3lNNAYswL1T3UVJdGOfrHPbJDYPlsF3Ox+sW765ZoT8633q7QmIaeIVS/uDl1hjaqjBxElr
0Ep1fFdSg0+CrsS5xnd7FG20ORJAQEPvmQVVt+P+jDD+8VxcfM5xmBBhzwr1RBivfgY9IdZem9if
cheZ2MbQ7RpdoW2Sfj0hVreSFV2MVP6iTqxsd9JrMYI7faMqMjjckjL6/jZqeh5NkYRIOggv/h4C
zlJHzsN6kRHb2mxCGppqtl3IYLpFgNkdRDgs0mCC9H/OZPuVTkzSVvaXpmjg+f0NxkmYcj22Exm4
12sitZcFwg2f+wvQ8cI8eEQ1f2LKFG7EPbU+dxbTC6WlPJXO4wfNfPlqNV3moswG2eto9XPJmqF4
ZamXVM2pERhTV4XOd/jAob1D80RLxjMLcPSMZtSD9Hrj1eVvRW+s9XavwZRVQ7xd+AkUmZwHTGGO
o9Gt1zLD9tSqRj5r6huMmpvLerGkZKm2HWKihVKKyD6l/ouNbmsXCiX9LhbWUyRQ4lQNagB2hLu/
6DMi/4TRuQUqfYsO/6uFueNwsHIVIaad6J6DyPvY5DBYITqqE3AXFr3ep2yWJJp3/eJzLpe0oqlX
dlAy9IMCZyVgNITNY0qwDjHd6TQMeGNpmBQp1Ax80hQTU3Vamwg7JVBUADsl1A/Fx2TWRSY+RDbC
7qv61evP/3jR6WdWeX3ZVv6A2AZfsD0ws/exwH2oPVbl8CtW/B9N8OqzxexzgNQveUO/bM9JARAf
h0Jo9C8iNRM6Ld4A4Pw+vEz4V6BsRGy30sj9Vm7U9LAmvtscRhVCmbV8knDwFOOEA4t2briOxVok
Bu/4bxANJtFr4tKbypZKk6DINUGYNdZK4zoDc8zVfP3Nip31h2Jj81uOV+kVbb+gcJln91dU9MHo
TmjnpmHGdn5POiVajXM7s8G1VK0+wANQnAtA11AQQFAQ32uh1muCL7GEJ7il4CHqas/8M3FLXc5U
d0CCUcOQKwTh+Z1ibbjzE4wY9U+Q6ZpHgUeaI1pAvzF/3MP4sv04dJ1iGjosKW0YYTZLIaTCDVXL
PSddaJDWsHhBz0YbIjb2H9GPN5Zqnk+hO3CK4urzXYBrbHyS4gneXw33sFyJQ8NY+NpBVhqI1xbZ
smtoQJOdRSsa2+uUgH1fIu+OiPBy88r0km17zkPSSod7efET2fgjAmefHODlZAkBI9GmNYx+A01+
aoxOd8MhvWOtZQ8IZVhufmTdXFEEzAOar6m+7JeUALBTGja3WZvaJ92y/exQyOcJCr+6wE1jAWjE
0AJZ8KEpXmWOiCzM1+nS8FKDWJMpIvJxVFhwFxFKFLSb0SbeaJYL+aSUCON2moLm7k9TJQNsmjVh
A+JSM315b5evR44JIUhvsJKyPxcjnk7R9NdTpw9tTBywb/5qGz/Dje/j4nDWPf4sV2r151H42a9p
BMaWB1Jy6VLQHkCP/lUe4BAMUbhjhC1SVezyJ843Tu0T65ZEKhy3W6PM4NqpXJfEmUJZIeuX8WMz
ixbZF3yu/q+t9p4/Hy8k3MPrUAw38MQEc20HeYpqToHxOeN03KzRd51D86AhfAAvD78e9gatX4KU
J0dMwbaiKa62jFu+IgIeaMVmYrvltd/fZxFQokLCR5+txtZPbfSbi/1X+ZZOmP4Shr4UycNkrWrY
2fzQXxvX6rRnkjUWTITk8F7hF7I7qc0ZXfU6B++14P0nV767NqO7/3+ylPeG9mN1j8EGvl/Ybau+
xmWf8H1yWvaQmlyV3yX/gnUvmEIJoxp0Ef3ORiF2S/jdV1xuPKawxMIQJOUP30HknZ9Wj67c1ouH
a6Nn61bOqnfvy1TCCsce2+85vGP70c6+PYDPUsJSnIbo0yjJj6T1Wzk1vb3xl/CRppz3dSeb1p99
r36SI2eDv4ofDmPZge6WxJT2SEPOF27+DA5pwIZgYdkvQZoierU9Zui1o62RnvmNIs5mY4qdOofV
sy+hCUYgYggZfnHzjByuTp1n4Z+rV1t4iNuEGATXnHNRK3crqphFe1KN18xq6gsHMQqCtAudLCHH
04ZpUl7AeXjtvR8nIYUMCEE+oh9O/uSkOEQKiJSStKHepzUN64IBZV1Bo03NEbYf6OPGmhHEWjZS
AlJ6GNT8asIkaqZSNLEP+Cp44LdBwuUTbCR+VnI5ZseHvHJBVFTOxFNlmwIGCROPB50NxRRbIaoW
NIw0R7bZMzNZznD+M3cJ3kqaLi5/vJTs3hgVPPVhN7TcTugVxZGv9flNUBIsTT+DO9w9O5ZUr3xA
YBJsNl8tj9GTQSE0qFC4AyBjI7NOiWhtVY3Qa7/6jSpuN+yBe9R8PATI9PC1s00mVEJ6GT2ZFwC3
NMj3lkK/S2r4dm1OhLgbQ1flRs3WIe/eE8zUYhDu6r22VTrgSlF28ennWVkSj43Tcm52iOH6gcFj
fgvtMHiGON600eOULUJ5yymjQ3oStGQsPADI9SJxPXiyrX2Asafk9aq7ZTK7vClRFX91Vo27TKFu
p8c3AltzBUfzRwvCiPVX1TM+Id5732LKhYE8bcuC427K/1oiVsLeQGkQNxogLFo3NAKMrHLqAlOF
JE4U+hax8R5Be8gte9GDsuWH+UTdYi5wYvq09/hYarOW1n9Pr74KwtomsRa8wWkZdnM5l/lPe+YB
8Gfca2DtmMAntpxxG2Jm8eAKHS9IaRh9kb8ufm48D0N8lXckyXRw7xVSFUbD6TuxC/g8VJtqMtv+
xz5MqNcYC4elk8+5g0GRDRhnI46YwsJHnAgXOpQQtt2eGxSBo2VsxVLgmUFs/phezeF3LANQYno3
JyrenCfS2rD1SfIBwn6wZgeZNOX1YricvrgveILN1QIRuYIEk1JO09/vAtykY7+PL9tKS0q3vwmk
clRwco174QAJPW/9ktpEM46gGGlznkI6+nIpY0AM/2oxtK7Q21y5XyNY5zOnt3ASJb0PbzYA3eIB
fB2adhJbWYsFuwSwJXoRkp2688Z/GgDmHvOqYiNb8eW9S6mZSAe2PbquDem5dT2CFE5pUeFYxZUM
8kloAOt2I6YPQy+ED8orNZMAg7RlmXIjtdRfi6Hl2QVcq8Tn2cD4QiR1CNwaSPWl9Pmi95Ao63qG
bObfw32BCnJQpsSJaYS7ETIhOm7e9jdE11AKhr//JKpfyceL9CxSdNsBfNsijQP78U9FlbgbIPPD
VmNO2WAAGgkYVzKyMHUhHYvGiRPGqEhRVl86vI8GNvmq3dBZTpxhuPmUIb4RhOLoRRIr4rfohMTU
3UWyWhQlzZa4ix23aqzfLs9sNmoDoaPyNpi54s0QEvvTaabDte1wMx3hgYX81fZA8zpo8CyKezIz
AWJfDQt0pdV8jn6hC7mQZDkdxWJUGpEqQtGfQwgGdi0aEXe1Q8c5poNnm44ktGgH5szMNRDw8mVx
yCuYmnjYm3VadnTaFsBsn3yK4QtXR3d58tEoCuLpJJb0rIURcv8qjw6rm4LuMq66noDTSnTezv0I
ioMwEMFnuOGp4DE11k+DmJIjc1nV5/8G427p6km277WiAED9vP0krxwcKQh4eGd70QpgGgRVdV/T
8KB56bhk+dDHhB4Z8Sf4Ge+CERBVOZb/G3id3MIlpuhbH9mGfjIuzv5Ur/ZfrgNNkvlp41xvMEDv
LtzzrAMlOD7XhWbro8RMkoTnq3zBNA4OetJmnnTS4ZlvGmgq5DNNhGnMce3++EiKy7QpsqUcmJPX
Hbo8s1FQNLeWixI/VGxjH2rf94ghCO1loicgiVQmY6cy+a9CpU8lZvKurYaujIhW9YnUEWwP6WBB
4KsZ19S4xGQE35AcUacOSY7YQ0QbFnIlZLJcdDhv0dIZPU+5m2QnJcx9gcwW7/UJQKqnmU9/pHix
SLy/b+IO/vdlrA7YRVsQMWdplkX92jyYF7eus0LXXWOFruophs++H79Ff5AVd2QDrbQEWYubd4kE
yYdID1PuyRDV9wwIZJtxv2syqf5QBcVOtewzB4tfmaV+mfTQ2fuCGA29Mg8iPIVen9gFlc1MTCk7
KB/1Vg4JD+g5zDhYNounz62Q0io99csvAMN1B3uEfAUqYJ6XI3sXSDm7UG8diheZluUTI07e89pZ
O2h21uY7+A8zyQkvUnt2L/w72rzNvh+zQpN3bxPan9FBjLnBWchnK+t7z6zlNB0NrTO8nsIaUOKt
o8qMZ8l3scDmmaedjMQ5o2RZ92xWOvdqP4embTilKLIgHLBF6LhsNXE3A5GkZBjZhCiMPeRBKfYc
DnNI+CnMi91pNY282Kn6qBUtME9zS5ec7q1jqrVAoeBpJRhF9l1A355DUQtPFxX1MY7q8lLSInDj
96DavA3UloRsbnDUIpRe/hXPX30A+H+2W/HmV4JeDCt48lBR6us8t+yQZJHgcR+27+3iaME9mvsg
mVPqirYSh21ib3yWGhnmhJfIz8raqVvLeo1ESIAByYfkT/aR9XR8KCgiOryd12td7BlHG7IzJYiH
ISn2yWLahaiNERVe2mhyfYTpoDlGZo5SbARcpksIWz20bnrwNOF9h2yPdCNviyU6+OVtln1hRP7d
dyEdghcsSkZDKx9wmWVuntOmKeZUrBaUwVmmrEizA2+ymyHTjhBrMyuoY3uaorRWRgDADVTREDEt
+d3DKN9znfF5GpydIHDfZ+N+kIQFMlqWCIzlsV5pBGHgH3e3OILFUUna+DmqnahuPHzpX6xlOp7T
aSpmUUn8GTLIzgHOWArcSY3f6hv8tK5YEXD7kXjzkd6boSvnx1z2N7j19+Am26LRRIsY279dMd0L
cOr3Ejs6eQuHNFaDey0H8Cz38rkWn6rP8XoKH0IE1EJjr54R2HDlz9WqscBeL66fMRwlDcQ2l8cJ
OewWk/BLziLY1OGKTw4hFYnFW4DvxnpHGwIVuj60hAAzpitDHIoFVUvIf3vmEQvjPnYEtDf00FIL
gkMbEETjS15glxCdbTQKwZDA0B3CFXFRFv7wGTV4Yq2hQ1qVjdOSi3+2/GrAvsTpyOzkUuSf9Q6A
7VojXaW1HXO9q5K8ns0KnVmxs7BflOlLPYbj0Rz+zCP/UiO0cDJgdtcXP+qiEzie9NdycU3s5k7d
SoGILnSSGONCqu5th3ikaw+iZqLkEdggI0g6TC9rCbSXsU0T8PbDYffMxzVCZta5Vv2Mg/3ag+XS
A7TfCM/Nx728W+NF39KXKUQkPxwVgWIht40rIJt/QGDsaVpPUMEqoynOBewiPxnYqAywq1F5CLuj
X8ZWFUx82KxA1JWuSeeLVZ0fVicRiOhnTS5kAApkfr3eCfhDUXaT1fSc+rEWkEbtaLru/XsrJyBI
ZBy3+FOVgb5jKyyLtanvRgF8flEODB6WcVMg1hJ6Wq89FqoTabNnRAR24IKuNzyr5Y69LcfcHmyH
xuRVtmIJvAHAucJHmBtyBp5bsKIZS8iQv1EB9U5+rp5pIvBmWyxg6+qFkNB4S5x6EIzqpT+KJWps
s67+IqYv6VZPpgR4UaUsckLL3DrWmvFUiTTmphXyCOWhQEsGWWWlvfKniOH+ujnlSnsgRWg2KvEH
6PrR/Umd3ta+0kVsQ20LHT4i4qmoQ904KBhpG7o7Cu53t6kbWoHD86Cjh3GMxm6dPHKkpED3sNk+
PZikrSP7VKTiDlQNdIvXPclJX7YVDGNjEB0/GpfF/e5VI8te/6W5Hj3UUnljg9cIwemve000Kung
TxdygeUtYEzcWcrUh4Kvb4Oa7xCQu2pzTcYqVn0qaTsdNw7C87rG6hSPEcEUpcz2PF+WZi+951GL
H++wE0yoFWhfy6jgyeH87Z3bZpgLHva+ZETpbmEcpJ5u3b/Ov3qjIot79JWfhCBSVveo71vTUCrG
0A93QHjYXTOG6k0s+CmQcKvIRvfaw7pj3kveUEQ848gJ95vkKQlYZusDjbNCYCS0/6pWDPArXtOV
0i+tg71JAiNr/ktGz5E5FNIc/10VxVrwGBZYt07IvCvRYyvK2uoIj0X8oMTW830wBKwFICglm586
YhrLP+Lngb3TeBQR4RjI4C8R/bJ2X6jRf7z21FHANg45Z81fD8zG1BJ0g3iOgRGfZjJiL/6M5zZg
ZJUs52ebm6Xyc6XTsxcGzpiAGSNrvqxSYVpt9wF1zLpuwt6xFFFiOfKA3tAhgfPjvuYVmf13zeGz
jsbSU0rk2SdmV3hRCBGwbTSl+Mi7haBQeqbHmljxsu4hCEzO7IF7Bq4a4XDmqTSPeXOdof8jkLOr
kyYtXUHct/Lp4BqQqXOZUfbt4YdRdQ8rgOVhipxTxUQh1t/7AYDRYvVsld65n8joxsQF+hat65jA
DvMug6JGqEObCfiHSQBc/WfW+/Lmv2cDt5kgfWqENsnB4FK2AEQogK8YgSIIYFX6bEWaoZKVjrwy
LH/+p+0QQCXTk2UfMtMTCuG+ZurBXWrck85qKJh44yHqPMLN+mEMlyS5LX3NWcwMWgp9WMsC68f1
R+GvopVN3FPcrs9Ywpea9vuxVJxQJVUdzj0xZxjHQf82sVJETl25goU+JpCohro8k+8im3cQGVsc
8vlDdukdQfwqJkNOxYlDH8CNjddHDLpEB1UJqUs2UjRJxVjfXpOwYdoDbytxmlDiELC3D9+ckNYe
8/4EZtyfrZTaUaMPqbvD08kWEyiePPrckf9dVIPAr9NqHDccJuGEPbRj6AQNAvO1Tb2pPlhox4dq
UVew1qYIOYjHZpw78LNKmxg6HTLt47AHs/6vKcWQIPe4wNCfJCR/sA3dfbrd0QSpf1LoEqQVY7KC
3aDyhLVd6kby5jQ0PUCWEYPenBZ0MQJUTWbCcyV40lMxv2ZoeGdNl6EA1g1jyaMQ/FP3g7ttMyUZ
Q/N+5DIuoGYGzISvKSuYxkJFHmblYtnxtDGrWCup+szQ4exgwNpEnRD3kUvy0zenQ9GWRNsg4kaY
lMZmHxiypFvmp8FraJJIMcF7s5KN0TGhKWg0d1ME2gTLBtB1mLKrFq4FWLiv+gnRK8/2lFqrRJ4G
Ck1c55HQ2A1Oukz5JHAnk8iN7ZfJjEJsXUFasMILOPzTSc7eMVYlmyBKA8A35W3vCYk4g3PVkyw/
nrfHi4KaKeBIW2CSfcBOotkovmYXgOGSc0ZdQvZ3YCx+pm+3a+nU66nJwlahsxCZrHND4OKj4t4i
Oyymb2nLMwH58h8kQKCAQtvAg68vX/LikbCkaU6GN22/eG8jYvmbqjFh0Qya7NH3OtK50TAC+Lvs
xSkc29ICW+FtgyV/eYT9pSyZGR2vqh9cQIfsk4voyGw3CmLfoTY1G+JkA9JW3y1NgI54E2ut2H+A
OGOc7Q8Yyv3LOQ5BtE9fLJczgrC953tFOSlqTJNrUuwy/nrbIjNL7bhfTf6S6n1ripkSLf3aTsur
ypmajbFhOeWEsBPalRmV4Rz/3lxmtldqwWjEcsXl8TUiuY48pi/z7xwrqSaoFPCfHqOnjVPPqjfC
s+D05uWQk3RzuXFU3/DrFZhzPgHYfQ/zqfp5tOIPLWpKyOw5RrGRU1rwZ1vJY3xQ7lVCtBwpJQJo
h8I08DW1wIKf/CpFikwow1/v4ZXloMPWn3YtbdpDrml9/fM5rlrqJ2I0/hZrJf2M6Isqq3fqSm/o
/8T5ffP2rx//AVfcSPtCxgUkYjsGSryLNs5reaac2LEM0cCxE4CWBcO1NH0scKjs/p4/p6DUhRXP
CuB7czw8loowo2mPsW/E4+jJpHnkHW6hAL4UkftNXSCmymHUgF0PpaeWP2gSwWI9VjnLCeOn+/y8
a2o+rffHvbF/Iqw6+beLK4ZqcPw7OMa+CW3rYfO7JL++nGkUujbO75ltPrvGhamKzyKHUDbY1XmQ
oFRjakdSO9pnS0DJQ3C2X5dLk8dV1G6rbbQ9BRq1+eL6PrFcEaf1QiMi6TEWVCogYZfov/FyVkhN
yOnTIku4oNzCexKwnrkipRJzptcIhoFxqQ3F3aJmX5I+XRzQokLGE1u9b7W+kIfcn7S+UrZohUmC
qkbwMWaFZiLMqhAapTDXX0J0XYR7J5ZuHipK82UICW3qXRxFSmYxrZ5tYCV3hHD8ieZyu8z97EXs
loqoUIVhqKbMRdZT6oX0nZNk1t3+DtPvOC1Xx+IEddQkfwBt/NdAHTO21wlkWQkNk6Ns0UsvwyNQ
+C9gGUlptcbAKF2DX+RSvBsWxQOYQtdPH/Qh99BxGwQLx9ivIGaLgreRdFbCQRqKfGAn+apcFJ7J
fEVxj34N+L2JiEm3768qJBn4A11ctd35p7r3sGIBivTTgHivRGSD71E9sF+tk6e1Sbt/igs1ofI1
xfYr1wKtofW30OtsYUgsq6BtQaV4mfjw45c2V4FuZ5lcTQvXlW7GypLVuxFPbz2Nl+dVB4qx8aqL
Dq3n6VaLZ55WEKtuG/yV1QWqNA2Mzd8mC0UHdscwNMIRzMYeGUzoff9F7xtpCQzC7Djth79MBVTS
9enj2aunoe2PO614eoGUPJ+5l4NgUGscYND/5kye28bbFB/5c3HSIiHu2UREF3gjgS/tXhsE3fmH
YQVLvx5QOZx94AOunpLJJkEf2T8iSZkn5FZXsaHny71NP0opSCDQwyvl4Dkf8T3jnCWvoDGCEg8c
0HORJRIggY5hNLVFxJObelmCZQkff5T/sXmxs4PtnFiC6WphWmCEvzm3qikcDKELMnZxn1JS1Jfg
KkIh0QlZIWAHlC5R3ULe4WYsjso06OsYU+T+xn9yh+nP9ahOZYUThJrGmHP1HEreZUxUyORnj6v+
ZM6o692kbKhXeNg7ShQYjHigDgh+YYhX8Pf6cjjU0Sby6fVK5XNJDi9ZAHIAaMWc0F8YOSjyhOOU
Shxr+nsbaUnpnmAe2UjjFEhA6jiCPVL1TwGqdWLe+7+yRcdKt/Fos/mHgjL2AZY9mBHxhWa3iA6u
qtN+HRYMNb9DqO+COsGlAZ8l0VelyMyYjuhr6CFKMVjxwhOJ0eTm9arGtWK23PdvDQwm40YMkjYE
YaEz0saT+4kDBGdVHw6e5Ay2bNoBLzLOsskaaiMZdrx0yXuU0OKzyImfjVMXYofUm0y8jYE1aUXN
Mo5vA61i/sk66ykglPykejN5UeliopAr3QYFFTrZ37aBqd+UsUC/nva+TQ1Uqeguh8v/mXhnMZMh
xgrcnxE9/6bz68JAibqoK95BOu1D8xFNWQzLygd70OpVJa8qz/UhFOuNe+hzsvdN0Ar+hJFAyTVp
1Bi0M6ouYasU9WAHRk8Savr4N0dmsVndxIFCLAEWQ2qsSCW+/yujtUcyIHd/cNthXlr6dwjl5DZv
2MXtzbn6F/bKnBOoTxmy/c/XRUqtXlwgwWzDr/p6jeshMNjpEs6K11xQXRDgUyxeuFXzSX3OYpfj
wOqKyGyuxNxaz0joP2Qtveie6MWlF2Er5dkTz8DGzzGyWyxnwrNyIsKzbRSWjVbVSxBpmXf6Q23S
M/yhoQR7bRJQ/Xw/ucTrVk0MdEha0wUO5isCNVLaPxKeUCMtynsOcPbZhXojzZnGj6SqFUJ5cEtl
xvFBN+z+2AT1GHXMS6DbGHzQiuPF3JvA3SDP3G8EHwScwzj3FHZMt8bdHSPmYL0UiqBH1KGsN2K+
5cXSuyiSyz4oJ4xQqlZzPMYSXXaTbR1AmwKqAyjTqD5fzkYtGQ8MNlxGcvyCqlGwykCDHZzJ40Ih
LHFinem9TAlXGgmZDuwCFbcaPKhELHcew8UoNEnnIMNrFp1jCYvNxTMq2JdoItCIJa5Aa2PhOZii
uwhOPgo7xlk/zvCM5p724SwzpqxWq5AkzP/P+wba2oz+SEe+m6TtPUqimYCsBdQdQqTWTdVoiH3u
yYttUqUb86TYXGYSau9HKUBkTQvIu7OtbgJqDNb7XerElNaJNp98pFKytZoRNEAUSTBiShA6I+cm
rf2qmZhic661ZWkgVb/QtosbVojQZ5ZTL6zlfbT4K1nGf3v2CMWUQiP5OpNjuiGd8Bh3Ans5+XLb
t/0t/a0/wYmmSQqNCnWiAJTM76TV7JflzREU1vRkazqJ73HK0zWhnhPpqfjmsa90OkagPkQWitAn
r3VDceLZcfqDHZyN5AW3FqYcCxLZkqPzulWCb/6Vp62uU0U3t1GcpKYQVpfEU7CTpm1Wji3PWRu5
d05JwqlPkoMIXKo9Xa1VR3MoS/DkqDJeFRwQdz+N7eFA9Y0eCnG7K9c6SgrM14SqAFd9Fm+i4NYr
c1TLaCcCqnjCftn/vd0ahCzV6gh0mVa3yqskcu99N33GCAFBNJnwS64Tu1Au6K00qLxV6qVHnhO6
u+BdsezjVXv41YT9w1B/38wUvVJLJJFyx1vNaK0ugpRrXjmFnA9F1hrOsIv5V9sutl0dp76rY+NX
O5r98Wb7be/sk2e/+2K7iSpoo4iMV98Q7LbF/rDyVFzZPSA8OCh9jNdhWoeOkub2W7YapObjXwXu
TJhV0GW7bbwVAeVPfqcCCxTJQ4JbEI1yXK2ltJKgIUgMXeCeNJuixuugFGzJHprMr7unoUavRdbP
9rbSxnw9h8dKerTTlS1wUbkwJ67asW9o7Hg2oCGPFy06/BggheZ4E3BMswbxiPfi+xJ+5phqTRHL
KSht2t/SU9jwk5OkmnFjFpjyElpLBwunKToYn34HKC002w7xJuJBrUW3YIN48nCL2Lgu/sSLUJik
gpDIBhaXPfoI6Ld8vT1j3dVfXFsLpPyxm+yqolEMPoSu0ispgBlwc8VoL2z58Vzx4umt5mN/Ygi+
jsRX0jlQMopnDXP6Vz71mv/Et4/+Y7zz7iHtbjhOxflwK6XC5LB1Uad89dc3V4NrxDeNNtd+cXpX
Okore+TDqpMBJbGvdFbHSGA03GFtea4kJ7Tnr+vYcUJKBVs7FGlu7tRDGXmh8kWifWBbK1MAi7ZA
eyT4qWNyjROe5YTqVnDinyWi0noVT9QvQcfvgV+q1gSQGh2RqESpm19bHETFZIDJneJ9pmdjw4gO
WgRC+8wMqq1/7/4SaI8FRpFRyrhoNSj62t+Om5f0m5RYERipetXHVDniAo6Rscsx17fS+irWiOAy
cxeAL1McIvjVRwPVjmZl5wMlUz09TgNxy1gB2f1a8h03hK9+Kw/5gyE+Qsywz8EduC66M6RxSe9Q
rYh1mTjB90rQgkVGzIT/PcAPEQin+NKmE8EfpUb9rDldSEoOe7YNU5b3t9lYTp9tfaSFdpRCLyIq
2gTeepdRpfzEJWw8sUOvv8ajaT9+4bicaLypdVrakrXbBbW0NFAsB1BRMhWlQWr2B+/6en6b58E/
LuhBC8cUCUIf1D28ZB9nodatgbGNR/F2zFHSPvlPCCp7C06KZSbfBoKKZDcZMLxsWKiePdOPQ4vW
oth7nAPsSL30Ke6t79xp1oMBkKaEpToxXhIk+O6cU8N+Xe14mlpCxd6oGVMULWXcF3Z+MVtj8fL+
FPJ75BCK8bEJAP6ZN+biC5rxNoRDkgKP/Z71abrzl7Z+RKcxAz+DbkeWUlySY7FqGQ4xqRMaxzYe
ocP95UYHIqPSw+8Mu2BPHzNeNnxCWfthsxO1T0OzDea3EFS+8mAJ1dKF0D5n4kGh07CLXtG2Wo8P
DgUcWJ1Tu86lgYJL7iytJSY4e30Sp4rA57yddRJgu94VmawsmU9Qi8pPVIdMfX6uumrrt6UKVnix
g03sQrECieGvyE7R6qOXcp9eQohyc2xhZCAfyH89P1u/6wc2RRlNy3ZeNSxQ53ehj8ppDIqZoCY+
DlZpDuDKA9w0ArtQC2cvR5LNP7t5i70yhxTQgazZqMnXtE6uP4FLhqUVP8N9MXPdAhqI/y3bndNK
wD4T8XxXGnecttAiyALI1TIqjpO4mPvjsq1ndmbi5F3w/063Jn8d0U7aibdGN0mEZXk4QkDTaaLg
RcJ6/3r/WrWEupslJwUrIGl/YNS8dtewhpfha1844JZlmjC2HpKQk2HNlvxH52FbGWcjUb0RQAp7
zZbBuRo3So5J/XgY+/VZ5teWin6doM6fSsQ7XTYm8Q2YtOtp6g2uWzwZRLGSgmKFHfz2Ube8D9lV
LE9u1G6mLIiZ3OQzsSwVel1qR8dZvQ/CEtXSlRVpo6w7VCHRX599c8mPLT/YEAUCcKbQi7axOdyX
ViDIXN3zSGR2qavTey045ONw/T2R+25Jhe5TetWv9gJUmmVjcpVsGOzd61gx55tz9DnNhmZwq6Wg
lWrbT+PC06ykCCCmkVG+GCWo54W3Vw+7WpfxCLwoYwYHXTxeYWgVmMCY8x9Pv7nW7SEQD2FX89v7
DpmnCmgeoT25E6rjtHkq2Ou5vXI7AHYY+OpGYp8lGWGRtAMQLecM4yFK3v11qi8aX0ebj2hK4NjH
UZLlwulZElMXLUnteUeTTL3FYnHJDcNej29hp2mzo6zmMtZJJJDdNDy5igl3Zo3yyOdgLeMBnmjZ
8Z4h13YfdgzAfKa4T8CDBOjzLyyVqCDgFZjpeUx9ttYkTyusWZKYL0mm3JPBiOqH3oSfAbFZjx4F
aQg5YDcGqrpi4Odlcvwr5+WSzOeXcyLwTrrCpIHZH8C7UQJx+Eno7XvLOhNBX1zNFxW7/KBJSkYq
qn4vkhMSNRkb6m+k6Fx24pXzMtze3mgXI6h2MWdEL0otO2bKO+xiS8enl7r239BmKrxLt+4u4t3h
C6IUdxutVZK+Lrdkdcn6UqiJEAIPRBtdIgfvJVLD6pt8GoVo/wxf3xjdRkbUNOabmUL0+lOTyPxB
IjGZ0C3RCWfuRM/wiVb0/MTBHZoHffoLEY9HydRelt9MFY4uRsFANIhTOxQCDn1Ia0Y165Ez2eBe
JFCAvpqG2r1ku8j46HLE1pXskH4jFc9r6KOEKqYwVYMpbwxjf4myykMA3MCjMo1rxvhyebJOTEs0
Exk9KyKN1NufB8Bvg7dH5I29xQD49fWOL4PCDpRlgTFBS2FutNPBwmreio8/C05KHJCwQiGVjGwK
lGH6NGyPyh7Qb2a6GBEnkfkHaTp2nezM4iGXREo1HOg9J9MtXPGwoAgZyWISwFvK/4/ncECwNN4r
H8/1AJYC3Tc4TBQILDrg7EQTJMszFwF4AuPnvrVYRRxIv+HFV51fq/W9N/j8cgt4Puwx3dfjeVzM
V9O9WfiyMSRsXJEh/sIyoTgxubC+396SsDJBTMwZjtB3jhYOAMAPPEwQxRuCjJnjYfOquEMkIlvh
hskQC8F7uHAqwU5maSGa/GnWmf5hhu4x8An2USwUxDbfXAYpZtotXslvHTYvaxixWE5N6clEd4OW
shjPFvuEV6ZCWKH/hqq2OVaxuEqq5OJTpIQwD6SvXWaPlnEWw9+3bUCTXduwRu3ugFQrY01UR2Zc
xY2I1sbLc+p+dzB8b/T+dJ6bs0R94fUSmBYM82xx0tPWnfzIjhwyb4qz1BSKFGIvbc27SQCaqEjs
lLSNeBghPHm4IqbFnat369jK1eJ7baVIoNQUYaIPPmYnu5jg/Ohes2yH2SPdBY7F+P25dwOD4S5F
cndeH0r8lVSxzDy5rjVlmyAHBC59RVLGgYFGqSCDJtY2Fol6sJjM4fOdheK/pgGhUvKz6dBPbWt9
2NJiRBKaWSoyo0Bdd3LoGM4/xbJIaJA0U9FPQEMc+eI7s1o0uIIl+Jh0nBJok0QVsdvbZRgNKG35
EWYvjpmE0AsHabOYe9a0Tj0FPfKyQrDWGJoIKS648VBnVyv0wGlxJ2ohRhqPWP4ySRjDNtL2UyBJ
y3fiVRhvmEmguwKS2Gonz17mpFEBIZ1/6JqUkRSShHhX946LLYWtKK/yrH5dVufq8ODPxE1lkLzV
hALvPxAPg6yKoeWaOO3EpvZLnzkw8wZFyQdtGxZpqiaKwsFQnN/FSQOOjHiMbQBBq1nkgs6cmohy
/NSaWpwdHiCkpIpp+3KWlbeWBb5DNP/yuO7yIiQ+t5gbX4tlL9DpP9FRdmL9++SV4+T5jiPWKB5R
EOqVV8Jy7Gm0qCBlJ4eYEgaFehpFGwRTKrg0ZDtsw6/jKzdwY4u6T6H9y7pTluxu+Kth9Wd/te6R
V8jTz76hEXMYWvoLH+H1ueAjCZLYqiBbfeDclBjUS+eJgzscvgrU69BA3wQeEehFIeaQZiUsFrCD
2CYNoEi0ZPxco2Jaj6kYP+s4JfNlivee6eB1DsbIeiYMikj43CoARikbuLYc8Weho1hcBlVl+HGx
Nrl77YmKT3MeSS4qoEqYm5FR9UEX7vI9Tf9Y2IUO62SPCD2YV6Z9gaIrWpvxue6loG2QcAYvrHxv
oHGOQu7XIKDVWfNOwT8ym9YdjJHm+HnviaBggCgCG/2ONt6+O+HaExw1EzKc++Oq+g6CbbzGHPlu
C1f9Nw2T3TTdboavBZ8mx1ILkFJOZQTT61Qh+TF0qiPqitSuQCvdMKeCitzoOhx5O0cPTmZTcXVx
QOHPwDqPJolyfVHgD0vM8JPEbMIxrs5D3wCkqobrHnfSnO4Nv1EOIvFcRyq6l6/cJbPKF0hPpwTQ
S54ngGLntxxFZ1FgURyOp55jOOa6Xj57Bt0UVGSEbSc5XZU40M3ITQmII6DvszHeanoOmKRIcZGE
r6FjFRSMqqIYoLrnRC2Q2gwIgzmIr3WvFaOTRwpBhDCKr2l90U5K6ZPLeLZI/P0hxd62jzg3azgs
d1Xm09XhUb07DDScEFU5X3Iid3yi5KGxDeQ/G8qwWIbY4zByKNuU/GixZUid7+H9Osfyc8fN5xQL
I/PJbhrLIj9OR8nWlKJU96PmCdsqhTkz0b0iyDoUWpoZMBhCKe9sfNWZ5C+1bpOuo7S/Zk7Uz8HL
k32e5gGhjQRIlHrZgXdWASpfgVjo9RybZvjsTXNmIN+LQnJTGraXpluaB0JIq4K8x5tw8e3sMiVw
0I4IDWwyU4msxymVfdm+73R26+Yb26DhuDumvjszR5Mu21uZuQMZpZzfoQq/yvDPzwH9a9NZ1Mnu
QDSYKwNlm+hUevEiFNzAAQCMtTUi7nv2gwFwllT1nXg9X8P3obupPVmqUJDYR5C1Fcm1tWw2BwBo
5CuyhmEye71UnipWUHXJfAhrxcFY5WY5LugAA8YKC6X82yVQ6NiYpUuZhXHnVQ+akvKfM2H4XpaZ
52YroPOTjnXOkeewLQPTKYNLOBU9bEpAbtZvrQqJuQuCjolAHCbGf9Ca1igq4obnKcRkfolLj3RO
N0clZI+CY3FLPsYlM7ghAV7rcRsRT1DDn2vaZq1hdYsHBimPW496+rbyWDeDUb3ZncLMUhV7+EBA
r1xthuOve2oOZyZBdgr+Yx7TEx96ETT/30Jpqd+J8QIqapA6Xdrq58ExcQkCGfTDmnAqN+yD3jGg
wFoYoaURdlURtJrwllLNED6vJh7Ets+irOx9tw3f4KzIM2JnT6evUNW7Kos5RC3LXBofJlFg4Sta
j1xiBAMjt2bY3WMwmqoRjit7AB9VLaXMSdR4FD01PfgEDkeyB7J82KS0L+XgumjiccL3NjfnWjwk
WLngGlgQFWOONwypttaWv26UVLqkARq+ijf7LQEEIeAVYahLhLkroZj8DTVprxSPOdyd9uGMyUWY
U1p0f/y0VcRJ3QET+mNIbb2PZGgqVECEWwTMRR1044bIAcIxawBpImdnXgSibRrz8c4Bh86VtOk7
SS1ZoL79JdnkM3h0mxlXdO5tgxa8TTqmWROJqXrs+9XfJ0pC5L7fjy/dR/qo/YgiEeq5YSkC8L7y
1w58KdPYaN1BWFhgf8QjkhtSWReXxrkWSmlBGcsvUhi7RBRhPrUFCc1GXUUD2POMvRR4FpOR4+gL
Nq3VCpUZTe7Ecf3esfpMMSaGyoewGbZHcjK3iPF9wdq3Q/Ii4rOH0NoSdVI+cM7S3zdvKhJqUgmz
jAA0/XAM2U4t6xIV+J/xb7BAe8KqM3qOa0HR0RoEv3khB1vjK0tjbgbRqckSSEof4Z8Anl80dx23
FIYHnFph4KOy2g/cJvJIPKO2aJ2DuntMhcv3uVvSMPYAUN0pBIUtgXeKgiznw2Qg68ItJOpVAak4
5xafxlAYSfLzxLKw38i4Ty8TRuWBCS0WEwOoKitztMy3ArbcOf7uhHfA/Q0eE58VK21URRkZr47V
HqZJI4Nam/O27p1BkSxVH1/EU/b1V/TtvZBchBI56qhsnD+rIzPwxus/me9qVn/VrGliaLDKj3R3
/qCHVkwCgrRMHli3iAygWOog7Oq/HIP1w/vRO22j0tuJZs+T7lcyiBncZcLxQ3cg38H/5Ftz0z68
6vNbM9cojAq37EcTXxMMEYRgr3rCwYzhwpiV+8LWBwSKBKDuxN8Flv3vt3B+KzimiHT6YQ1u2dy6
jfwrGqnO9pvezkMIEFuA2DbowvK9JmGwyslIPKOE/Akba3k+lOOLyhejgqo67/PyiEsjWhuhcyp9
QL8ff2wIN37NhIZ19kpy/VeDeDMgL7n72p0P8N6MhteIF6KlAYfCDlM4X8CiR9PI3NUev4upGrpg
nEkVK5f9fhSie/3BvvIAXHByVw2AP785lfiPDNOfAg3w662MK/mT01ND2xGIU3kupGGV4uxCChVb
2CdugjWN6euer4l6B1chBHVg/0wbE4ltkoAZXGBRJVFbqiStMJAAl9DQOC2Z9OQQeEIEwnLUhy/5
T8BMLZbgdxXNFvaWZFytFmQp/bqBd6pSnrUO6x/PC2K97qif8U1AEV/8H4s+wgPaYnHc5c5nS7Sj
r1UE5rikGBnY/5JCjgQuOFAsMfnl1CJSn9JTYtmNHm8W1QK84OvE4gyrhz9zuyQ6IzZGd0n6r9r8
iAcLqkgg9q3RF7Q5Wv5QWYPcyyMWQpX3TsBgUE27RnklDUcAiwic43BhGXBv06yn9hjt6iFdNAZY
GZcp8S74xbyTKB9tNuFLf7Wf7+05dm2CrzqSG8ChLo4jZOaJErsu2AMaR1r1gBdMY+ErFnvuQxdh
jXKsZHq9fzbGkkRH+ttEEfwcwyTyhVpR/nZQPxsCgWn8x8shZ6VeAQepvBcUxFt/3ai1KlwglqB2
CyCpllR0Ff1pS3w8PMBKs+rqgPHctaXf1t5ro1Pz1dSqLtrBCu8vd/4nPIzeU8SCkI+s2yDacc8J
kdlo+7Vow5GeWuI5wxR1C00b0Ye/4AZMObRXzD2v6R/6d0h5/KqnoHzn6wWs8um++Vxg7SO/nfjx
WydHxIE0pHMb5Bv6G4PG+cMAZTMB8MlAUo14jdUTwfdO2cLxt6G27JWNVGM/GJTiPfZ8RNxRojPG
7slVqT71BMvrS4sZe+KXxE4WpUD0j+261/pzz+dolmv2ujURUEcWCUq+vwNI8IgRxPmGnDuFtpak
YrM/DS40pDxWHQ6HJRqdM6XTIiUtltazUbVly9Zx2NQas6yp0QcPcS/+31IQvsWvR0kATjuWUZ2y
TxzgJVGu/lGSEobokiDZTH6znUwYt2Nd/xOqSBDL06bKpsSzpiBxz3ysr/W76USrMqqI48WaHqFc
138DAhYBJwWCkb29z/i41y6j0BhHNwAZZn8GRwVTyc9lSRMWzNshs0Vu3BUjgVETrauj370/2C3C
FstHADY3Lo7d4bdo9QTdTWWVoRy8GlqQ7vDMG1q6QshBJwt7ywwDXQIkXjZtqecYPYU+8S/pR+gc
gbHvHyQ6ePMS2zcrjuTjeXc54ua3Vu6W6SvSZHGLXq+23wHrJWfVzpbI+v5deDjeV1/0zi9GY5yy
K+93saM8VaBm/RjgmYUa2dcJmtNRcw9ijyIPXJlWmiFx13MCLVorlAY+CrCX4jXakM4/alDzesjU
uINWcqQQz1FGAoW+uAA/EvLe0ET4i2O6Xs/aH/JWzY2DLJL7izqRK0e7v5CMBQTypG+ZgR50yCaR
BVC0O/uB3o6aQU9VZkSnInHLg7ZIZFbPZEHvmOrQtZISk53dnVHkmCRCdKiUjd1ia/s5FxX3otGV
1NNOI/PHLImVP8Hd5BVQWmJi92khXBdKPB5zfW0CsCKWi+SUllb5b8nJaZsxMl93hhqisxeVq6DP
tSzylIJyGCIuQ9jo3zwfPo53SvbC0E3tj5FFvAkQp7EoaMJ79743EGkczxtPnzLWcHmlmagJhp3w
ymhQdwZsDEYHqGgD4N3sEb4HT55QrvxifxjmhCjEdpuVyqYRxH1XVbEYAm2eJ3E2kE73S5cOe0m+
HnWX0bU0a0FVy5qebH6vki0Qn4jnYZMfkOmL9HmKjXu1LE1ObyRomxFYETzBRXbOI0afwDh4yGLf
4eRpAvyt62bi5vVTQFqVwbDjFBVOwLx7QAYkZLknyf0oMyywsMFN1Te84UkYnjoB7oL5su0xjBhx
yRrp42i0Fw75XnqtwK9HbIVOpPcs/OKcTT90LqRFxYMwpu57oPqh+sDR0mwKWcwlF1pyoomhHXMU
hjMyL032BMJ74Sxs0X0z31sPrRClN0zKIXyME/y9mzWjRxtER6V1uSGXfyDdUn1imxJL+gO6Rc5J
8PfIC8kCRDFBFaCDpSKg6ojO0sQ2pxKC8jritvupJzj2hhS/Co9GM0OJbmnmD39KbWF5ObpaJWo3
tzYlzgeaqocjpkpEkdBxkycLmDKvqcDry5bc2WvaQfnt/5iQhxbwmHeheN52jwz7msrmAhkwfB++
s15/Jv94B/OC5oUusMdHDj6IkPFrkt2daKxgysh2dXaN9zWj85LKVaAuHpn+SO1WfRJg0Lq5/0CT
PIziZDIUbH1A0zc0oUi0MupYa36gO0vN14Lqr60JK9COQ4eumSeOfA1kStUkea0T+L54iO2ySx9H
wrktgQqQpPeINzknTfqwTN0JYPVFnBgt3/T4xLrlU80rWa3n6HhNG3e0zIfgMSoJenKeO6d8MmZJ
mu3qULma+hzKS2b8/MvpBSwuXIgEmCLPoSVxRCinNXatfkusF+N+FJElnCFUUjBnz869MBEVglDd
GXhwnQYFVPsBzf1qvezAirUd6+UZpQVPyH/uSyiR5Ahz1R8kDv3GR+/8Gm9OP38alRj92WLNueyU
K/JCK9RaJoTKI3nSGC69fMKwIF8YQlfTRE/3EcSse3MIDh6x04Mw0QQAqXpuJXklADfB4wuPsbmy
In3/vwRQEkO6wZNf+q2FW7B6MnA2iY/rtEc9emrtIq4GbmrDF6orpE/uTO0M9nHYRaU3T8lYFoEx
D5YL1yjgxE58GL7sViv+48UKtDS6dIukAhQLownBxjpPvnp1OnoeqkN9KXOfOFwDp7x5cA/Hi6Gf
kdL60sZz6uMXX/lyt6MKFCqYU3DKCT0JRZipXIX7uL8zib8CscszViOTsbK1GSou2og2PdfFJPKr
uzMCaIVtp0e2HGlVPUwMH6+UP+YH7NUzIaBo47ozMWBJrd8e+iL9fJgFCOFev9qZpnny9RBOAQ0w
sL7+JlfYR1D1ztL6E7EaAFcz3rQp5lrwysVpoFrNT3qthJWqSHHymYJU8S0NxPeVl+MQyd+5RXx1
oamDU7CMYbYpou7dbiBu7Rz/IqLZ1rrYC6N8d1EP02k4zC7P/4N82yUVQuU0KR8Ejp6Vd5BF8PhF
sus1DoJ+enJ5lK1pfezfFa/wgHhfOI0R/57WNeDcVpvUBgwytNv2Zst7QprKaN5xiJQ3V6LdrGK7
ExGl0OGdg5YE6vI0Icnfp+zxJXatcFcIofsXCGDGV9UHu0cYAVPIVlPUvaKuIG4x6pVQYASA6U2Q
eWMCH5A1/mZ9RuRLJYys0QtCc43tJjNl2ps1m4Uvj4z78yU/0BmIAWaUigwpFnXnaoDr2lNAL5np
0gGLQfrqxBCZbocSf1inUHEv+fXJqJToKxRlMLiVva/zwwBm2sXUoLNfpn3Mmp3YPDLs4SbIHuWM
QjPe090uZ3qNljVzKetUsyOJiH1XrGaSfYz6aXyvl5nYA8OSpjEBnDLznZQgdb3RtXcYwVe/vXEi
BUYP0UT5GA6QXLbsRWbj7iZhtZWAPK0O6QxLfmkvybe/N80Swl8OD/um8nSgRdfvBTlsQ7eI0uDk
g8LoS6qBa3HbQkTMG4wkz1QsZ7CwPDfrk06TvtWcHKWWYa0eEePsvxFZNPvWKrPPws73vRNGN2gV
/hRJkhLXyjfWvAua2hzNE4Xqqsn8aCxCzalzNoPpG2dM/PNOy9pQOis2E2QYIpnc5qg7nTjOVPVb
y3qbO3ggaKkziLL3drJOVyuHlqCMZKqR5AnIuj9j7aa6c10xrmJooJYTbgeFdQMCGiHhGn6xftfv
08ce6M/4mSmVJrmc9P2JcdPKaENXuhlN9fCx13N69NCRdCZcNHtuNLs3c4CpbkM6bnmbhLgbQ4QU
dSFPc9nJeRwxHzyxiNvX6al8UbKRm+m/nvBwHV/S7Vzbi47z5pXQrfJWX/MC1gjqhESxq1fdWTfK
zrPMZcAjJB6IC/uYuwG3/RsUOyzPmWICOYthce3kvNTG9yzFCEduy/yJ+lpWg546ALKYFvUu6sMI
aFAXEfSUxrNDj5wku1f1crv45wb98FeKVY1g04a99hUNS4ROWpNqHllWS5TdVJar8G9ckE1D/qMm
ANaTI9VhxsLjSKre42C6G8WkyEiJiQo4Ttd672nkBYYycvM3Oyj2DMdPN7h4GGIoJ+csCr+7Ga5/
eSypUUtr0XsQssoVXX1Fk3zbUc4lqSYF8zGk2uHRnwxuP1cWYpIZ6S8iOkVudEH1XP8Q6YRIzECa
Ehyh1O5Gc1MQjnKunvW8ekKhI6WQWrMv9pu6d2GuUacYjJdYfr1DFUhczeGDFfqqcr+I8SlkdJkS
DcDnSy+tin/Igbbo5+DrYTH+nFfFigCr1gcen05Wzb2INL7eXFOCAZiLFxrCZrQAf/B/iZTdf5xm
YyKVaP0aTiOXYTjYtFWHi0clduf3Q2sSsh/gT9rpXiW/YPvtG2EAC5iql+5JGeHTLdKyACJ25h54
ZUPhWGNacqB616sxBZoEM2+I0BoEWHYUR8tzsPlu7+4ZS8aShpwEptWQEVvhByMcqZHc7PNpigI9
X/ghkB8m9OqdrUwc1tZn0eQ2bCgJCovF7izMsa7rz6w+Jg7soxlwrxFP2sC+O9JarxS9fMPvjCaO
/93h9xC1roNoDOGZ2dDkDIrV4vv9WS4x8yEPiXcpAdpbwzyBFoFHfdfnZDV3N+OGF+aNo/1HLD7d
i3BzsCAnig7VPjXbiTWEOaWx2RGf7+O+UCzBzXYa+V+7o7b9N8HdwCwqiRMyVNx/eju6U+PiM/aR
ChU7aV5lV9fBsLS/qJX7VoDgdmfutSMZCx45p6XQW0EnF6uBAVooAk4ypqu0d2h1sP6WMQc1023N
VfRpVzAfBd5jh7a35KJ6QRWDQHFgmCzBUyyd1lbQNqrZv+2+5pDR3f6297C0D1itr8G+cDzFtbed
P5cquiqSnRI0IHH8saVKeAW6cyEqSF1WrrxvZm1tVy4nMynuwsZ6i6NZWo8qrFX5QdQFVbtdclXQ
sSexbbjQPsnNnEycQnZFZWhAEFpG9nSnAamPQZqgMwIZjxYDkvQoHUh0JGQer4QwZGvqWYajcOgj
93DqU5py4WeW+AJPFvvVEM7zPvOxjpT5EKuhnEqwyQJ5XKFactYb+qVbdd3iNMalUoj+AIWgsb3T
gOvuw930lZGNBq0FlI3ek79/8eHwHJ6USSxg9+27bne99iL6QJmY/0N5VFY3GSXoio4dfpBZy6Cq
ZWjkHpaZOgM1tw8UGBbBb9x8u3uGJ2ML3pg+hsXz9mhiX6YQfxDohuJ5w96WAKuh+I5LSF1YBSHo
XT0KFa+LKNlnNQqM2QjQLhpWJ0XRpcI876JffmDzwEtMpp2CTUwek0DTiNCTuK63Kr21SRD2x0Kb
svtXD/POcDrymNJEJc8Stda/Lpi5XKOueQ/k+thjqJOF25KSVLxLGboEjZ81MHZjVyyfaVCuLA3w
ZK+obTj22nBs225TKYpyTQvj9ElX3wmHaoY4lY1RuYHyS5m1K+0BPqgSwEK6786e+g3A0ivdr/ng
aRMiCy6QoiiETkhsH81vC8dPvYvzibM8CVdQ74R1wAQEOq1AvN4hKgIvHO86T+Cger2Zg6e1k0wV
Sjj2ztsKF/Ep52+dM0djQjHxpQnza4Q6dJuB9h1EDqRoGNhxv9KgEroOWAuMPghVqTD6Q4LroPNc
60stVbbQ475/SvEN1O0jeeWj1pa6nr3I3y3uBaAZ37Bw7pIAshWt8W3HIYt2xelpVXp7xBhFrV1R
eRaC95CD+fQnKWxNP747srhOwyz0WZuITTSqDl/C/x8eOr2aq8/CyplQa6iOsMAx5Wbxjzpn2tWm
CyHV/LfVmOvJzTkQxL1Ke34n7X02Vv6D0/zzu71XDejs/1RWWqb6t/76qp3AltiV2N016blUIlTB
mK+odHak29hJX8nOh7C7bwC3ZnOlwbV2BgRXI/ssEk4qPbQyA9WAZeFP/VLfeLer8jh1LFjQLNxe
LeWb58d7w76Z1nW7uI7bQ3alWw6jM7JtEM7bEJzn0mwrJQ6dChOuYiFACVX4w9F0fwO6Y+BzWK73
9mY09nj5vX2FSJKorWGndRhTgV/yXJVYl+cfJujPEw1eQMNy4j5BJFLgmlesuXrkq7N14lpEW354
UBPO4faBU50+/EH6mIm6AG2O+NSN8t0x8VDgw/BVRw8WdRLMPPToqMYRYfwABaKszaeslFI+2sNt
t7MLZn27GYoiY+FjDGwdoQWWTILPOnMo8eusHuiesjMIZ43q+Ypwb6wUTBa5G8FkzHJNpAtm0HXD
GFtwcNr+79GgSnPmIfc+ajMIE9vZLPZTQhSb/6IzOWqPW7lMStuqAiODn9Alr0Gb1bVIfrNAMCSv
pYdhgcD9mYhW28tXDCGEgYqsE3wpoe8RdNgIrSQ4x3IXvT77JiU+9gTlfDagrCRIYf2BOwjk8jwC
/7z90Bk4iuP1su62OY1+iIuU8lgmBrYRUFxRPEaOPvYhg6yAcV4ngFdrhv5rc8KIzVW1MBYySuax
ZpFF/TD4KOBWXA+R9xER/s/zIQta3SsHefFLuDqPluKIwZ0pXlpcbr0H8fAYbnyTl1qfpYujcB1R
tvtmtbzgezBjbwAivPB0yPav71N28gHLDRz4XKz3IhT9w3eykQSi1KlJTpFv0OkdMpFXmTtQbPms
pQLEJw/aVkh5un5mBjPkz5msp36+SY70xuSjqNKsfne9xbT1b5ktN8vFsOpaiQkeHE+gJQmyQxXU
HIQdKnuPAMg1Z/bF+mC7yP5Dllgw6syClaa0bV+DbUpMNe7g6sOdigMnm6GyNa8Re+Tg/AOuqni4
4Dmejmolg1rs3sOwRgTDWZu1AK1FSGVWss1tb7jUOtRaQc0FS5ohv1NSxMXx5pdNDE5SDZbivIDi
G8bR2pbX0f39n5H99K5EkO7hZURSFAgP6xZyiiozhwiPix6wnuXLkAIJpHHMy1BNfi/2T130pcEV
OQhY/Vr6Sfqkg5BTbvnv2IIBXGJ+RjObxSlzaEHgyVuMB36C9OEf+RD1sPC9hW12AFscvqkKcQOk
2gLiOPBUoRK5vssZC+Kj3gJ+AikiB3UjUHq4LrgOtRMFw+5rRXZfiJtWzPUI6zhzwtW4ZrJ2CSj/
oShIomTOkWp+7AGhRsjj+SWWTMXFm3otb+Sak2+mvg/unNqp1NxnZTP0kaSW8Z+NzUhaZsbEeHzl
fyzU+PgvWIIiyW5S9cER0mSSOwJXvTjSZLpKVeMgCE6T0eY9AQT0EbD8uOTU1NTIMjn+6zDwMuVf
XdX8rim5D7WnimTyXK23vTgSw3xVYFwi+ZIByBfCjGENYxEqYo8hKYL8k3qeYaDRBGBXPe0QXEP0
LpIuqc0TJjwb1G8yakY1m98TFartTMaxqsg19XAayYF6+ncQKGpHGwUE+28COGa39flKiFn8oU89
vmEUCiKLoKOKVAGPQEtUnr+hwSYUzGkZmsO2hoYbdbyuURIrSfPd/U0y6yQB1Jw6+K/MFGemON/5
HICkozc5jjxHjNRNLIDK9g7pX9TWI8nF8eoXRDf8MMF0q3CTyz8f2YIsZzvlY0uDSicjeE8+jj7U
ZVGKrL0elrP4wr51IGHMwFFgn8noJvruLSwxnW8KUeBb1yulDh4V7moslrvdl7RjmzaixbArg2In
lwVc+nZkj2ZwilqIvYVEZhBR6gKV/sqF6/zCwpgDrIHHURukR630a4buNlJPIY3nkX24E+sFdt5E
Vo9VZlJCXByGUJELFokPRi0lndjp/c0J+lRnJzSgwXDpvLpFxFyOOJMtdpbLvtAwQHdgqjHsOEoW
1jOwTxherqxBvZpAVq88dU4ZJamiO20kkZVUj4zW9kO/0iRxgeT3+VcFXBdgzj++GrNXYxIeyz/G
gkv8KrSUpYYX+rUQrcV6ibndfUXQx/aScH2gCYNIqQkr9T98F6wsuK7BFSlCP3Mn5NotVVYCs1AF
LplMFQY+DnPQ/DlYwVGYvjZwnly3Voa8Qe7I/W2XK0mlBBcCpoVI92g/Pm+JyUccO54UWJzlIE0M
naPdRirPgZ569i81/xwFuN9+NDz7JhEBeRNGY4UWbR0VXfIzyhdG3vfufb5N7OWBJxPjjdygEqeu
GSHRfmVbZqsxJ0P519YmPHXy7u+ht7QvHJOUpl2ShpLRA80pIuqzleGqSAYBeHC1oAhf34fMVgBR
b1ksL9PxsEBbxsrLHRNiI4sIuBUuowe5abtCGvn8aSEkqzoxGH+jloCNk9m04d6hNEv3JYxd7ElE
lf3hgS1+68x2ITAPUYvVwsMxFuG+H3wuUTT+IZhefArgnVR/BFOCF7ifrQMzOt+narvVwgMyVAG6
n60bvFdC78bH/l/A6ut2A3xzzsmwKuUFDWL42MmKCGUhz0IWp29AH4ANgVrFlU1iZRKMigXYQEya
AWwWYBaWasvnbnJtMlpAzXq7QvfTQuk4DK8rppvuwBsEJF8WvkBB862O1Bhfx5Nii0xw1AteExE+
s47Mwhk98f4GAI4kDu/Bk+ZgQVCI8+7PiI7oYWQ0NTqv/r53pvkrStd0SAkzbb66mBSqyI+ASMKX
jlERjmv4FS+NP66czZapcw4P4fAMbSK7yju1oRrS2dEf80Pd2SfZtGYV/OA8fakURdmndQKcg+lD
E4PpxD6P7syZbJw42YTBCjj9RcbeflE4FB2tMw7rDR60RZH/JVEdde7zBerWeNmrU0RHKbN3WbVA
mtmQgYWX7jj4c2Z2Ag4oKCGEVZ/7D1gbof7Ge1QZPN96f+rLnCRxloKpyolu/ESfxUHthL9sy7c3
Asg/3YklpLyorUfWJy6zvtKHFynOUc0MePj+tvFkQtvqZ9KgvYSVfOz++ZvvBd/USKkNaw54KaQF
LjvPZlEra7rPxf+IG7xlWsr/DfN28S1XEzRsiL47F/MGiVT+qOv+9FWQd0fMTgjEYkmqBgPh53Jm
MBZW90Cv14CODUW/2l6V8q2Y2rKymEpAdXvnfkmbjVNT9dZ2yWXfm/88o8QzlbD8ULhzokBJJ4vl
q49RfUOZMGcutBqVOT2N4/eTdE8eGU9BUZDew0Gckku85CW116vO6iq8qwQgmAWGVCO+zov1zWyJ
1U7x5IOnK7Y407/V6VfY9yhoQp/Az7XvX1mOrgF1IDA7H4ez09rvG6UHu5aZa4dLoWTlDYCHSWMr
vJlw8oOlzxpBCjAjM9kQZEFyxu5hF8apdxh3aXNyPXPllI+YiAC2+RbRH0izpGwstH5yb/PEcTXY
xY9pVlC4+HuYuKIijdfCZePPYhC3HOLHX+uU13jQxTyqB4roIzQNRc3qnLmoLy8SjqQgv8AjbsoG
1n/OTwnjGMerx/JFGnDP1goBPog5PsaPYwqOoNc+OB97XKR7z6cWqZaq8VBuJNoMIVxYWG+k7cpY
t5VGiApANO5/Rx95JPn9R1ikkDoifSSsLER7m9NIBRCXdAzcO2njTYBRGsu3WULsJI0GGvbWJgc7
1wzsXr+zUm/MjDEKDsbWKvOiiGD/IlE+lPO9oxmpbnt6ibXLnXVx6lZJbFrKWWChyAIZ7/pp8DMu
/Uc2DizX7sR7JbS3YEUDUrfoY6ePiWV0KUcuZVgaDoTr66o3Ifq3614AGAjDEEciDS7xgT1my+qq
xdsR0guU0jOwhdLNwoIzts/3OHutu42tMyecXM203AfaKlNhE88rI2reGcsDG5zAPP5VQRQ4oQzB
bCNgTU3F5AoVpcowRQLDhIkKvWc64/x+YejdyMyC+IeOJ4X20ay8VqF/kpKMafrp+SKbNQwaPpeT
vumyPLYIPmXcui3Ex2J4t49Cjb6w5zqL3aF5TRqcjI+R/8udacXJQAQMgvNlU6e8wvT+f3u+iffT
5VzLhd4Av/HLip7dB7YJvKvDu/T4Dfrk/ZcwTU0DDl0DUaEooqd2ttsrKlWOIm5/M7vSjOgx/OL7
072IJ1XLNmeiXKiXE1e9Cb8QNDEBE1wADlIPm+2WU+jIWwnKg+14WSJxV+C8H69Uk7iSlufCu084
RRtmeiknlikzMG4Cu2y5uZsPBTkaXPyRoh9UJrbLHeUWZS+y9qvQrKVXPMq/06V2yTJjS8PTSPm5
d4I/zy8csefMRt5XNNhnlNtCfzJcuGf5UT5OtNNgQnuLzogBGogglXV5nQRd5UE1ocI+mtB62CIi
4m9Fa+RpjksJRF0VMAuitX/OJqClErRBheKDdMDlYSbcwbNYlZs4DfcaLU8QzePHcRw157QStbBr
LncJJmBguzHtge2aVOgFGq+RlUIpvw23K0mcvnHFJAGlvlQkVOQ/28RkpeNUV9dXxE1G6itzsuFW
ozmvt2vV3rKRNaWM8t0LTdA12cbuc4oyF/tp5HbDki0pFR1ZHPlF5CLj95bKX09uUUw3UYmjVhIo
pmPt67pQoYmntg17SiQlvBPkJItJ/cTDJ7SxS1zAZeKkF+SI+wbEUycAUQEff8zwofchYBRtSY3u
40a3PzPwQk5Se5fuW/6peoVIqhXlCw8rkJV5WkWQIJ9IoCW1WPGU0/p+/szftyrRZvOWe2PTZEsd
eFbWH4vtxcHXzwZylsN5zgOm7K0kyCv9gQ6NLay1enzyFm706l7XWbGhCBC49QUGVaeFIZWrZ2ug
+A5Hdz1KCwZcZZn8XkRWJm1Vd+3cfNP4OdRy6PGTfy9I14F6udTN/CLLKGmwEn//9Tp/NRjAK+sg
xpwRNXkiVPurb989Z5QeUDifo4jN/0CrPWpEnvXczNk19mjn08O/9X5/HYBbAaUCgzOb7MvvSzVT
EvRGSIVg/wxU+awYeDEweUj1Rotldz0clAwJZwGhFzrG2NhPQDvL1tsTIKZBpNmsodmwCPSyxn8X
5z1hw96Vnk0MYW+IrpgmygwuSXH0P2PcXLp6x80FO3MnD0GiRb+7cVfkY9S9cHC+vKVmcUFgoPTd
UbdMNzAEi9tN2WGUjMG63Y6cnVnjURg15YQFmnIPPqUfvlQHxNSgdcc/ZQaj1wyG0aLfduEszq7v
j17O2SFSgXMCWkUVyuYVM4PHqUU0sIuKMDyPuK+BqmyhoAYhJZf+w1HwKJLUZYySgmZ5ku0pJEyr
fB3lQ9FzMaPFcoj/bUqwxgqk0kh5OiwyVEyeS5v35TkZbUqbnSMO4iNhILx6IlCQyQDBTI0Y7sB5
rsbWQGb/YjxAyl2Z8BblMl9j/nyVYzgm4tYX6CMOfCsEgggfZTgPa3NxExZodvNqJVsKMpP/UUnr
tqOexztDMrIE1uKu+ZRiGOqq4n7swKfJoibbwf14IY7ZdNl+x39tgui2hTaPBQSjOa6op+KKTa+A
U3LywNE51VCdQmc8mJQGe6tnUkTR+CQjd4nDO7kZc1WLW7tP8EvTNZLHp0cZv/VFbXgvU+fMQUGL
L0rYNqqvvK7fxY3nT4BYVR+vWTKwKOvgdDk6v4aJKa4dORlKgpLbQ3L8MWt9U1Wagf5Jjc7GXHtB
rB5/+OiknKZcV98E0Tb2MjVcdt2Vy6+ZO51VhN/QASZyTihHtewlhLj307kxfYAE0wD26uZt4Nw9
RIusPMW0ApSMGkawIH4Qrq+An80Sl7Vz55Kn57oNQpna7QEflxXG5b+xtVnrGuyxY1QfLqOu3yJw
066xeVFVphH98LjmMU+/1dBFB3eP1DAPH68UEmi8k7qoAe4lQTu9ytcop8SSlCkj3CGp1d3XvG0m
NGjt1bkUfeq+il37jqVxhCSgM/G2uh4fSSQnBZQe3FMmfh20rSuOdli6/iKrMiaQE9faRGKarzsx
PFGUvpNkBUSqCofnCsohyzUfGO+w72EMlL+lgfH8RYt5FhjYcDk8t6Ki2g2dBzNcHELxPt/DC/ac
b9P4L/Fl+S/Zg9EfzcitXUr2Gga7REj7CLSpbfIlvtp/CX1OPF4/T3OiEIA0r6x3PSTQvTG7pRND
MV7lDKAB6XJDbIZhitdZbkkGW7g5wIIZuNj3tKuKIL9n1qwFFRqe/z0XP9vxoqfxm40kqBOnk5IM
eJG9rX/21lyA+qzSP1utKOmQult5l58X/zCvvE1g3kuqwvV1Q3/VjogEMprtH0RH8LO1bkO95RDB
beqPNbs/H/H9xKXwn4gfLj2SgInum72ncfL8oMVmCKKX0eeZRL5M7OdclW5wCV5p99bciFZx0hZ4
MOlQtSYgPJ0SwgpmSY0c5YuYIshR47bTIha8SjDxWQJ7FygcnbyP3kzPXoyQ48U2FRVJ1hmcoouI
x6wbtsyI4NaeaRgQ4L7PwuEbMmyUfmZ8/d5EheGGNMrRvdXB4xktqEvB84ssLqtZUo5apLDYapox
EXsEsswmpIhSkpJOUWNav48avE7oK4slSUOkdvNqAW13+rAFUPhyCsvQ3xDLHjIf0pV/iUq/TGAL
2xL5jFggHLc6gveon/mwd8TSrlB5+3bAZ0tgXC4+B1+6AlFfn8ovhU09hb4WThQYSe0zWg6ymzCd
CKUFAeHr9gVQsT9mL/C3eUeOKBoBLFQvXEmH8iCXgh6AUPtp56l4Z6tI50DyW0dhk7TS27HljNOl
/wieAFGdyXAR2DPBT4/RVQXW8cHNkAZavqvgqQjm27joxveVYtWqbBUxPQ+qElfcaMOcK/+4PdpT
MfsAniDpK9q+6TamxAg1qXHuX7WtQQbzqW/4w31ecVFz5T+nXEbZlWcoICNdrx/15mSFyJnP22cp
1umLrb2xS40qurcAMrTMwJ28bP5Osob+K2vaRjCNt6OMbLgh8kuaYriEwOJjGgEJyADDeEEB1IuK
5nxi563tP6HICVOxUhKmHpFTW84wSYHhnd1nf9wAEbemfKjCeUC4Ol/Gm5G2HFhI1c7q//oQgwjE
I55vSGAFhDLmx/pwBBf3L5aiY513Kf7C6WidN8DKlmz9QUApopsLA5QegnY0Z5bMfOcuaDW7AePT
CjUxoYtKZhw3OqkFw7tXcr9GroUMOhvrzIwg/qHSnuZ4paTtRDhdIB8Ub3uD2hZgX0wviSLezFkl
MSmxzCoSvjZblNhV5SxYSjmHzfVcmI4/sddBLsj2c7egc1WOOccwfI9Y3RHokoqlYzYkAz7fACZm
71PQs+FEhiPeVBoDmUoBYXd+hQ8Ql08UbIgVf85V0HoGiaavGytZYbe2pJauXA68hJjRSVOATOpX
AKpLI/XZdlmO5CRUqgMqu6Wu+smyCIopllJk/2FvKUUN05KbYI+eX67BrLaST14rW4beGAfGeNYM
a7SP0tyCqpzf2fF4t7tJp0CSL7BSRw0UHTAUOLiyLOF6/e6zou/FKgigojGTg75Wg/6+ySk9VjjA
/yybVCcL5nAlImk8aXHrV1d+49u6i/xpN9Msm70gN0Ml/3X8jNJFRdquy3CSYe6JUhofJUvg/67D
SrQD9yeyhBKiixaTXGOPThM/GKTXfKzT4GlzF9ygkFhQeFjYDhXEE7TmlSwGyydA/opb1yAajW99
xFr0TIdW5Xkm4Lj30rmsPbYdMxHpxUvzstxyEaAdFTH12/0/Zy86B0zcudKn7wbrCyz7sMg01BHM
7yqCdp1gDsQCOaPDUiOT559jJ2eD39Ww5XmgdqwGy5V8ZM7gvfitPwTU39eygVCeEi4pEu/ii34O
mO0pnPL0U1WuH35ajFWTMJJ7mx/u1ybXbyX+zlLZLbJUl/I9vS9ydTaf/Nu3jGa5Fh9rTEYm3WVb
mNxvICDmjcM/PKkjMAcXarvJgNsQCzJR3EXiBEny4Joz7KpLFQE+yHRwYIDBNNYCPKePwjIQuaO+
wqWNZ8HpjqbAbFbSmYCgeccYiLiWsuhus8CuLyei38i04awDmfUPOxN4bi6GHKe71YwG3qjuNrlo
lrin0zd6FHi6QUuwHZlRQPHHBijj4tyRA+mr2US8QM7BY9FGJxyeGk5u3ljO4PGhCGkoO5aVDt6B
NkBb8lS2ryRnrsl6OVGKh8N5CEIFItJniuSejvPPa0C99+2GaE4fGquV7I4H/En06KJRJGI+MhZz
GVQhWyFNqYfzCvb/TfRL8jcLGqMeWi7fJ6xcmYf60mVbyRtpw3mWKwtcikH9i/bXIS7W555BbDiO
axN4qsiuoBEw4WMju8VWp6Jmy4bIicfN8MjEli+GWBnZKDF5HdmoAHDHVDi5+T4DGZs2I2qR4W5e
U/zZCyantY0fmMjH78MEc2hFqOqIgR+/xubZJgTDZoeZk5vWSCKfmZt6H9P7/vM5clc7JUXgT9uv
k+tsB3I8C8hqSilteOewv3aeU/iGDTIq43UrwHtKrX9A1RrFB3Z5k7mFfN96Es6HPs5u9wZYix4O
7iREiGgIVrg+rCsqv1Yw88uCoWmRdB+8hkyXO1/A5+cXqgjjACSThlBM3G6OCeS2uAKLnyToyAaP
Vsgd6i8BV+r2DgplS8FDrIHwv1zTb+etEBYSuUkn58t5/+Mj6FSZR9ciN/kPyu6jtBe6rMI/QdcF
zvvbbw+WVlkIRnlxq3Vt8pzE+BMml74JdnifaltQ5ybY6pr9BVb+cp7bhoD6i8HhoPPgAaS1J8hL
aPoKzl+xJqSA9rvoNESkHqaIPYB3JOIfgUFI9RDPoyLFRlXPx5hXbsQ8qMKtjmabnfDPV8FEzrWJ
hboC5ygTXv0LZY4VC+czOfC3hBSuJ8iycU61ZMYxGXnT6pq7EM9c7g79lIPNT9/e98IEUm9l7TLB
x31FHW9OHvR3Kly5FrlMlMUQFXn2qKdgfazKbEIbslFt2Dyckqci665ogPuC0UyZ8KkB/oN8TrlX
HPFi/VZyI1s469QZAfnTHpb63xdV4UiIBIBsxijPitT746fYPBKDO/SEsNTz0E4dx0caLc4WXjxq
/m9J8WVA55NtnNfeei3j/Z7xf6R7UmLaW017X9gKhWSh8cWxra+c+tDgTF5K1aoHds5rKRS6GDXd
cVqgCtz4frP6zJKUwF9NxTmIFW6YaG7EQRFXJDsgwxC0L5uqiOxGN/Gng2O63xxDYfF81SNPgg8A
EfrUgO/m5BYeGpHvmP54lpSBI8Nto9lerzJngKmETL6X1hED/Mn1wJO47nvDKZ4aufC43Z9bWnu7
ZikdAliOGekj5LbMBUe8XlNq1KTB2ufkM85I1tZLpCQk4nn/YCvkdlNP3ovZjRdwBCJjDGFU9mcu
QQpDqX7gsd6A6W2kiXR9zpYewFi9kxLwtGtb0Wxb4CJZ02sHQK2LsOm8iZeec3DsOSZHaTMc1L91
CsdfpIdZ20VJ/aDVPzRgDyJaYn57ov654UgYTgMflqXu3N0M0DnSkR+p6sb0huX4Mw/DT9Dgy8rP
hKqe0IBMSgaUM55/FPUq+TBjfXq3EHPXq6daubtTxYR4Wf3MMV6m3TwTfrxAjbEwIxoLJCZh2ETb
WVXXRRcjzRVxyfMjms+zBOYczww1v8ME2CJu8nwj70QUo+C+OdOij7dSMgSD7CkflgS7WyXQfP+c
CngI6+1W0QRmraDJWd39F+YWE3nHhb+i3aXR2+WFu0YxCqznHhcyc38FB+xuV+YJxBMgs9QI2VRl
zb/5UNwLeRTHaw6FODKkykJYgytURKEr+1T06U5WYBatkgm76hGbBpC01YqjKOXlosepFHtohtpy
eX6d8TOaPf4AlPbJ5mvZI8PuPT9+NHK+gx5JlH0A2TPfRvKeWU10Q62h9YULYY0rssxdVf3W0WFM
8jyMgRzWXZvt6LuyUYSW0zRdteDotP6SRqFaHrZfY0E0d0jE50WLyL7D/T9b4RWHKWl+FFOjlzsh
WsKiIW/yp1Qo/KuTstlrbslZGyzEaCFqpuMrt/odq9/DlyaR90iZgzouSvYz0k4ioG05oKnnFpI8
A34vZ8hCSsiH4FJOMKV7+6WzxAaj9Iz3GjUohLnkUm6CyyFrJbhsyZ++4yVdVoRttnHRQLcLfuJO
v6KuqWMHFJKZFjrgKSOoQQFo/b6WF1oYAD7MfepMpYt4W4QACjDa4DZtZC68qpVfmt0iG9bIrZY9
10iHEypzzeAlzljLRe5vaNKWmStyk6Hizb7/Yb8ehPTtljgjGg+kcFJ1vbqs5rJP5zVuFEL+0lkQ
h2tEw/1GjPC9qjV0sL1GB0oqBoMaM8DE1V6pArTp6VHmDU+Nd88hi69DuQd986AslfW1fZYdr7nZ
2IX0qopHbVldqgT2QODpCo3/j8fdKsxfj5gknafZXnzBD85JAWSMYEMHnk50+dAeYDzqpRvEWkAg
Dr5sb9WrVCMhJRKsabsY+IsOi5nnkYgz3Eylv7sRTVH6r+q/gHBjjnL8tdH/PfZrvasI4pXHodsU
2LEhMU74sE+a64sYtw55lWOAxgT4Gb3KrNVeWqfVQeNcQ0ycCRN8tTcmXIo2EnYLa+d8OFyIFYwe
A6clk+Tj3efoqhhQvCNBZlnXAmklVbw3K80njRL/+jHLXN100t79tL4hL5nlemrqcexzqshCdvTQ
ys0asVfAX+XksszI07f2jiXpDXwF3fNs3EGZ6azU0YiZyLjHmzmVxeXa6eYfwug0O7Tp3FSVBI5P
fwAG7btm12jMABW2Wwet8pUujWhb0e6kxtZ48mJEybTyvzPD0is4A6Qy7f8YOLjqBliK79jRu5C1
S41ZdhuKeSO+FzKI8+ToKmbTWJnRg0HsZc+Qom0MmqZsO9RFKO9wP9fpDdU892OKcIC+G3w0qxao
1VipGgBO0PpCRA2hOd6FsLLiXq3Y42WmBqP8sgJRfMJv1PYaRcGEwtyiP/oxeV+gmuL3Kc497q4X
/JEW/o1ZhofX/L0u/C5IIMKUrK3RvmRLKbglVNanHy/RztVDU2JFbBWoSNpYgB6Wvg0doiixnQXm
XiwDSZYrNlXgW6eoYd9Cp2+DPcKqQZgB0WKyB0r5AxPJxfxYxL0nPV0a1766cpSlDG4qH9B3vX6k
wQZEGaY55vi+CBkMYdPAlr1q8cvx0kwXrmICyVYbAgYdCJ20xgWpKsl3PvxVsFh5+liIF8y2pgS7
q+NjKswxzeVFbdZOjI5XUZ89a7uyNg/0QF4swesJgcBlC2bzyOZec6YAhgoTgMdE3xtRtST84LAx
V9pskI3tFQqKp+WNQMGnlqfhGZFnyioGb0vikT75cfUlBcXXE4XgWCOOGMejkss4LD3vyejTpbFG
t5rfqwL7u6FEKAY2BaP2CgWvwg24ktkeseqk1Ungz8AsyxqkCsHmmQBWVVhVUcDVCzjYZszdrCON
ysASf0I1GyiFhu5C7cIu9FJj0Crt9+zY5XBIrYQxwRnyIjVTBvghPL7PkLr/8ta5kTR4u0HKJmjV
ElIKayknNr5bntLe3abt+G8SkxL7RvqJN35mDwoaRFzg8kZCSQtlDkRb6uF0WKa9M5dA6fwtuJDR
Zgp921nbMpI/aX2Hd3jkCVxho1UwNkCt8xhR7z307eZ00ZeeJIYZpti8NSbrThFaKuTigO1tVeDW
sNizwJrnh78o+mx/fnSYbUw34rzhKFpFRaNEG91l3pYs1gPFQ8fbl1D6oo2oy4n58F8GyXD6azD9
TXOblVBVjI+NyNxsDcyTSpqOMg0JTDO/vuTdbN+ocnnBMpaxC9OP6XzTHq7BOPpNVza9iZIJHtSB
Fpq79C3k5pgWeFXsuEIGHIw1w9aPQIsnMNeajUrI8RaKLEDfCNZ9MNodEopVcISQF/HydBUhErSd
wlg830Nzsk50V9yLvwNyPMZDyVwTdnHh5TUIh1Siw0BipZZ/NStSy9rAWhyZwwiGm9nMuSfZSWt/
XASm43KrObhXybLV1tgNhqj/Zn+KIi37aHlXcN18WpZIrD5yFPHuMzR1Y/cDf8dSfOqmKyO5Wffj
PyWEggnZV+JAUNWzplL8m3qd7ajR/Kzomusfn9RP1T2wJoygNP74b/JIUg2P3pZVJx+epJklgYIe
4oo2icagc6VbOSU+aazW3SA/fRZrmCUYs/gm4malY4UHu2XrozYwCdN3uIaxzdvJ2b8FnHbE+y2I
HfM8LOIG7D1cfKl7cZgSCUneovDSF0kiqm9KmdRe8kqCdKZ/L+Rf5He6Yo9bV5MWpZuNqMC0ecmC
dnit5vTo4rWwswtDUX/GZavpGo7xATtMNnYzNvuQatnwRPAtxbSVPa5ArRZ3r2Fg4xJcRIj118Md
vc26W8P8RY054z5/CgSlURNpjnCOhLn6UnEuzZ+/VIoxOuwP8v3Eag4w1fx9KunlP8ypEJ4D6TOG
ZLXqI5wZcADO2BtTNFkTB8Bp4nEuJoEeUX3D2+f/OWQ7IALY+Jq3gff+q0Dj9DWm+RNSSiGnxOoR
fUFM0GsfXVIFDtYe+XuAyXiwt0z50jJrGW4ksorCPJoSwZZqZNy9nBMEDEuRLQluY8iHx6eR7Tj5
UVKt4vE1JLbZL7BwLOjI6kyk1qdYwzHGI7nD6DtEFSijeJuU2lcf+6cd+p1xHDatLOjnUIIE63gS
52DNP3WmCWedI7ceED8GG+43AWsN0tQ/LZ0Jhs1Kh2CI8iVv/HX6Cs+UT29qfsuhGAhmOtD58QNA
B33fpD+Ou1ufaBLn8uIPb9nC5XDJ3bolPNpNnakocEE8lnVhcm4m+N0Vz4YB5MqFz7VHzWU5Yln1
ojJjKO4wGzPz+HYy/1S+6uPqtSoY/0XPnN81FXj0ZvZXTHK8qmab79UH8njvbBHgfFp06QamNyo0
Usx+jx4TIhvTLZJ9a9wuymF+0qpMklIOjBIcgXGXcFVvl5FKRVxxBjyq5p2fhjTtAUVJcyCkqY+h
mo9fGkcE20PZLz5GKF5IpsD73TssHUyn/3Cuqp3YyYh0gR1FXqJF2c4jNa4Se0s70iYpg8VHMSXx
/g+1TEFDzFx6vM4b3AJSeY3FS6r3BmD0yZzMEEfGIMZzQFYmU+Otd8QwQj8cXWLdAEyiQnwzXjp0
LorRnfczq6x/Bmvo8XJ/5+C1T17LxTlPJi014BNA5OQuPApPBwRelMu96mPVRQsXNof5L/N2bRji
vsQfs9pJAkYLu8x1iv3GOhi2oyLEcUSVAmO5sI7BatodO8eSRbnexNBJUiPhy40SdTymfQnmRFqc
LMYQT1kp3RXD1BEpU4FqE+K6YfsrAWwbLIWa+m496vh0yinCyBceN79X5GT4RNYryZiQiK7D6cRO
GgWNg/+nzHoKqRm2EHK46HHq9wyRd5GSao4X1xw0GbRkWcJfI0Eh0VxKfMpVKHyv1Gec2P9kFy8I
6DxhATvMLlqfhdUjZ+3GQucOjHRkhd6ANhuLmK84/fJJxe5SZ05REoVa/PdGpYR45DAl2tyTEo9D
rQdCa4h5H4n8AZ6ZJsD2rXTpMbWYJYPh1HIrLIDBlaLsslShmz8Wa7MwR87a7+D7m7yOEChIHWKw
DOCZlsrlImsDTcG1voE7XtrjCiAGhzOU5X7/BOq6qiQfQea0erHI9FlAFEEzrh5697MiXAnoHzH5
UuSdR6cmxWSD3B1ul9Vj/opqfT57hOclfRppZhVaVvS6T8snWH0ddktNk/Dz2unVszbGyk4LaiAf
NfR/Tr8Bxe5IhjDTVo1cpksHrQQfz85yDoGM0n0FhVPzYoat6X/92uwZaoBYmHDBDO9AVXlo380G
+8ch+HeWXNc8BbYgBwPilfbN0+e2ha/h/IjuJFoPFehiRuIOQNCPnOB3kU/Qtz1jmoU1ZvGMW0qG
Re+UccTVxYkLC4kNnDif7xulbnUOKIojyGTkcqV6k0W+4YVDE7JW2IR7K4welraE9cpRVycvPeVU
0KPdh6hoB93xFWTyLghyg2bm2BQdw0SNDrdUOdYEVsrUKSgVvIesN1dfkTyrrhpIQ/WcbtlcW4Nc
m7lSEMZrvm2hIOypcDQYaJpG7FGl4+lHBrd0A2sw9o9iHUkhNDOH9/oS2qW2eg9gawtOADukhFnN
RwiXWklIF1Pxd5mGqVGSgecWpAhJLjmIc1XNRHqJcPJy7JV1NZAEADXTebl9yBGclveHdqvJ7HJT
uhvKik0QCTpiU6jYduZiwZGEZeDJqxhc/5sTz+pSqV2TwNASBH+//1rhvCd6Q84k5p9Em+xGNxy3
Dsd/V3ZgrPKQK9pErM05kNaBZqjgMlEGgm1tt++lItk8yFjqshaAIHMuENcN4SiB9WoizFKptLtr
OrEAY44uVv/u8okt4gdoiOkrF76SuJCVKXMtJd7IObH3HRhm3eq9mEGwk4yj+voBtkZZLgC1Kvke
8OnTRuh/eMwAJMRBudAB8AWvtQVVafDEeu5okGlACxRzi0cNma7VDe35JmPY+JtzQ06M2yr87TXa
ebXMVFy+iZwM9vw3tUzU7kl+98KTnDFGUFKgAHHvzt6ki8uUxZZciYLpf0tQoVMVPTXFkgaLvOxx
Tg9LYtWbgJ44uO2Hrf9L3q1oaM+qLKxHbzit+lhwIlyCeZdEgRhJWqUedThwqHQow7v7IRbbkhGZ
vYMEOV/vCofGZ/xH21CvEmS6BXf82N2Eo9HvmkQ0v6JNJ9cJ1ciCKs1a1XmEUkE2przrma6jG1EI
zdsj1AiYd+Tm0ZrI0EVmXWgI0YHqJBwQ58QQ3vH34njg6iIQaYsK8qm5W89bdx0vntO/Rk4ywEZm
5ELEi85/yAjc4RSC6LgFumM/5JMpYizlSfueda7cITfoVy47o5CxjbwyLCWXvf8ek+c1cJ0v0lR8
ELW4qvsg5KQAfarpYEUYUFErP0fMI3N/GYHOL3+8Inqwv8Vxxizp1ngSdKUgiq/Ss6xnjKV0s7Cy
UvvGOxHMAZcJl0uALc8zU1CDMrDUdsyvatJhcs7g9MZDxyLl+3mKEZz135EqSry8qtJ+FFZlKi9P
bWRga+2dw2YAwU749zP//LMqSkaXKNtluHcfYckGTS7y8isxJJOjC4PpskJAg6der5dgRF4YQ0hI
LTwDofnVVTtgw/5Gb4z+FoD8nyFEyqtJsWWLGpIIuqK6ZHXCSZ/QeRMLwMFV+a4I275ZtpUySIiv
OvVVPOqFb/eO7NbFhC2hhvAyeOn8fMbKhmQUCbhDzBWTZv/hi16/xU4zDyJuSzJXzUbYLZ9axtAy
Zm5tNS7zpF1X2WrJ3o0VuBJJIf/1YxjOIZp9SKIqf3zW5THNRd73i9CAZGilzTkVYzmk7fdJs4Kg
gdgLJjmnnbMXFNsUExWcSjnRuS74Lum4rsErKSXyDBb+YuGk/SRluxlV7MrUD/L9mGfP6aFe9zXH
nTZL+zIG4uK9yXkv6ya26l/hYT0yGE07/upTBv8H0IcEvzGpQqqV6TIhU7ukC31WJDv96MCAz4HX
BVSVUz0q0p375OzwFzqPN7EFUrKB96vlBK7yLjWrERoRRvRQzwxU7LjggipOiy5Wqh0L85gx2SXQ
D57XuqDm7c7u4tzjZT5HyuZ/bo7+cW+Awn3Rql6E9kWG8DTvKP+4o2dL4hcO+cPrcyD5XuihUrHq
rGY1VpzY7f5CmP6Iqu+vs4h/WcQgV3Tdzcfp6/FIBrWlmim5kCW0l4eAT0KnYVlwQrS4F6II4mjt
xz4UMu84CN404JexL++SpQ3VG4XKzewpQ4qyPHVHAH6TNM5c6vew5LBYgwIfDfzzhelolscVnukw
zasHUEaYxLOfmEXHdaObtUpPIEhLpLWbaiEytWf1o/pFlXrrbCwUdMIfUz0H3c5Wqg56fFM3cci0
j32h0jZWi0haIrpq6+Q8n4YoLNXmvRh88YPAilLZc7pPMLwT3mUF/IqrzZVW85FHgLTKpEZlEA8X
hQUyP1hRuN89KbPMkfBiIUpZ5I6ktiCUhNPAYzSrYv9H/6SlXOp+85soeNgmKYgm/xFSq7bHD6/5
JjBwSQBxJ14ourX/K9vfBIbmeeBpQz1rSJlNyllCx5OsA3AE8YooUBAThKwDlLWCkgIoTGZ+gyeR
8+ev1/C2qJOXnb36YGWVGXJ2zpd2TOB5GjjTlFY1Q4hn6DedA31f++YvZbkl5AHCCF0aKz6sKGQ6
rZaxGHF1QfFq/1UT1GdStFf+/nZiQiBS9ozjMcTwkZLuTWnkFA9k9j+hlwDzMoZNLLKrcMpSX4p3
O60uziBrLeq0gJ3QzbOH7dUHalIoH0fv9qbjsxyLxoo9NdwZD+caBNvW6cJhHJ1Gx/Vr2F3qsJFI
J7icMqF74k3NxSLATn1wKiJVsM373JuwOqMkidaL5uzSGriy7XwubeumC7v1JF28nf3S/5Bf4vIA
HArfNMW4jjfhPIaKeb6psa52SPdjhl2tITYI8PjX+1+sMIBh5q6PddBWevAPnPuOy/aq/hZkyZx1
R1PMxAq+xI8sG/yoNDK1tZv7RoTfVYC9YaQhRL2FT1uKGPg/UJHfu+ae/8d0rs+mauEHK8CqVcJw
mVRl/4TtDQ+oyCwftOcIrSnZao3k7+LZFbQD7Ddd3eQKxtvpHIzVok2sm+gUgWBrSXuaAYMbkq6i
hrGGbfe7gxBQltSYg0AxFmD/FvB1QbLvHgSJ2t2zGqHdhmCeSmnuMOdT1o2Ck+ZbWJkdtMD4p+dL
QMXDFJBxMITqZ132vjfpYE3ksLGzfPavYcpeLq4WEEL506q+DqsIEVVErlI3UA05MjR5Woo/NKlT
OAyuM3JYsMyXSFJ+b+0PI4XfnIS2OGY+1xLmuiaCfX7+/uhxZhHbV06m5z4O/8bHm/J/awKwndnh
+jgsMRqbh8wwkmFqF2f2CErMNn51iSX+nitxBMgzJi8+1524rOgbagD963GFr6fhGaqc8M/vpUfD
MIqVK+ZZm1oSs+cktTbv6W76PjPmiqIWgO/DobDxXDRuXtY8sczC4U1c5qB7m6JkvNxTtYHJhzQC
f19B4rqvP6mFUAN8CvXiHcT4hFrKE8uwLvnG5HgX3lYg6rLUZ+tF5/dEYjbi2JTg+ktXjeF/gCQE
z46oGY+FB77iMZB+2/9wvsMFm0pedJshxRopITC3JFo3e+NhM7BTcc9nzXI3hWuX+LPQLyUN6pVq
DRbep0zb60hQ81kvK5vpUyjvv9jmdRGyPAsSmV76CSqRpoWOKeU5Npc/5EGyCq+gyouuU4z1bcz5
mEuVGEEiwPMnSTgnbipbR1X2BPPTfFaYQ0tjxLK5e3fidDhpfWAy6ae5D1s0ES7Y8GpEpdb7j8FM
mTe6+oxrp6EPWgIpBRj6NsupRc+aZljXic6czMd7QtLBEwV9JvPXszzrw0XgZGkXQCQh/f39zUXR
9PIxv77YTIQctE+hbcKF7YqzrcggUvx1viKdzznl2rm1ENZRJ6EujoViIzTYKlJdbH0brcHhAn1P
smFzfT64T0S8mp1c/H6xzg+A6z8LUaD/QJncNfYbLWeBmCGTqoVZOZhdn2SCzz0jlqdJxwGsMtd6
oTLEWut0Sp6f/E30tSZrk9ykI+r4vMnL0/AMLM/FzlTEjykeVFN07GRV8zlmJGFmTexV0y2XlKIy
gf3OWKnF71F/dZcOCVMA0flpymHKYWpVCDS83kmQAD3SBEYpsWxBm+J4GtWW2bd48dtPP26d4L2F
aoOogblzspvpHqh60LYjto35Tchd7lFbh61frclLBcthCX20DU2zB/ZY1oFcjaJtkWpkly/da01q
QtjnF6GxnvdvfwfSkH3NXvqMKdSirtowb6Py2p32/3hGR3AKr3XUNtXhXTzh4IIofkxcvNEirT6G
d3E7hIOIaUjnJZipYfLuBgRWIEmU7TaZkhu+6oDjTwhXHtvIUoKnhqYNmVQbJwY1KL/dy6Ms7gKI
q2nHqksXlwyZdJJ+I/PYnAcgJf8kFr2E0YnyNPS/64p1KOdjnM1t/XvWi0tODoqAIOt9Vequ069P
91mOJWUXeP/+C29yhDFs/EA7IsmVcrPJ0QiDC7tsNbYQ8QBQzYqs/BJ14spl6ck/+/CX491bjpJi
p06NSDIgEQC/s428R3eSnrp5EOelf00CdvQAU8ilcjMORiUJSZsn+60R6URF/JzfRk6ybxj5NqsB
JTGaNsOMiTa/v2jzOCyCBVgyP7nNU7MCz7+Wssl3xQLMK7OyFErpGe8CMJLybwXdJQynjbP2SJgf
51SaL2HwUPpxYpJeTwEtH28Cj9+ZimQdpJSHXs2qoxevxywt/ma3lzpHlfVf/hJ8rm0eozuc6YTZ
xV5CzAtq8ofl9AwiTWpq6KEN/ZUebEeh1WpNopJiPvZSru0i5ZBSJVAfm03izXjGSSZ4Y+j4dRax
rLN7t+1VmYui39aXweWGR7z0yyEhW0aOxW/YU14vmTX3PF3DWWnKHhvG3wnNwAm2li33tVe6NIW1
Db2G2XKPgRlEGEH3BhYW/lA1hgApzxnUj6Il0aiDBAxL9oOBacG/QxUAVoQc8kePigok4g8umOCi
XRliiPPQIUU4y8CiqS/V0ejjBYvCaZEMTRR66XnGkogpes0b4q1qitrBD8Bu9NmxL3AbuFz9St5T
QCv2/CUWFZ3k2CAhfUTMPbnQfTjwWB19pNbhHJ2sTuMNPCeCm0PM7MU4/NUDwcuaL0zSL/5d1TmO
HNXRXrSantQA8GXEW8s8ublYPpI9RMDOybEmiQeL/NBr1RifOS12ib6L89jUhTYP9mVfGrL2fFxK
T2vx5nFtfQvF6H//7v876e+mgj/Gv4+OBmuhsLaShvoaiSOmIGNLJfxiZeiTP4q4u4DTuQoEUsLt
5P9sOJT7gZbQuYzGrIBEtT8hCxLKBAxlY+UKAiyLcdP9PVwvBPgWENSE9Uska6qezZ72bz/saUhK
vFCaq0329SyFaZmnwAXnEDPdqNwxOgrCUKL2zzKywSdHWH0s6UibsEY/+Wk1V/cSN2MNvK/Y5iEG
I75n9BbYPbtmlSBpqExAYu3F0FQsdUIpXg2/edmtDd5cxItvRLeU0TfHqiZzb/3aIYtbw83iF4vI
VdkVHrq9qH35GoEN2TGYN0QQ/IRB07qOAbSbRSjLUPP1TQYgBpTCmGfiAkLJmvH8NTusjaDzalJd
sNuHnOyzBIO9ydKa2jrTRMRCBKDT9/cuz644Xj4184hZjL4DnpPzzogVWyXS/4OeHoiJO9CelB+b
ty8gQdBhp4B3oQGqH52HUuClaDnAUZoFytJRZbjeOXtrKtkz8l+ObJPazIRS6ypSXWM5p0sziYSx
htFVhEuX4sqi2PNfpIFgY6lTlwlP38XzwsYJ1Y9vx71W1QmqZj/jLqn4e2PwaugvntpYyA358u5o
yEp7chDfK4c1Tbj39j0M129/m65nCgHtWhZ656Phugn60dpHo0jmAF5nRsUbszto9B31TvRSjxnC
MjuMPjLUImBUztZF2FKgx4t/uhe1oArXLIhHUMFOX9XRt4o9ZKiip+LyVzysG2WhOj+SLFdKf9Kv
M3t0Wb3pW9pS8QiVH+1j1NCQgaehVzc2u2ujI6yKvrtCIBgnOumOcsh0G9oHBeqk0pEJaaP5j2Nv
4SpLmD2DwrMgHFz0jaxeO8tiyufhSYFXQZvHwRjNEEVE/P5zdsedgoN5ZI4JhpBRDCHuan1QnyJP
ZthGYBtkLFkLCFtqGCdoHp7cejqJlrJqJiSzs1Eho/DcmZt0LdJCFG7gcCx/bs/znI3IiAT0IYrr
qoPyiLmS2Wj6W78MP/uw+82/NVt0plnoi9lmixeveAReiOmuKAapYuStopv1o4h+VIfa43t/LjWn
ba6vSN5olC1L2MzR8qmBtR4tPOATYhrC6yE3bg91B0q0d8AW24+UWM4QGxd7ry1aC+fc1onK5PQO
eBMPTX473c/sECJoyjpqJMKYJUlFZlfx6jjwTqRL1wpzuy3A3VmqGlx3WzvhA3h28bfPoLXVyY4/
gEDfDyJ/avRZWW9poPeQpwgYqFsBm2pqPsq4r/QtKTRtVq2E2AqerqLozGW7MfrnRaCHOk0WixTp
ZInUNqMxzxn9cBwGzdJAMArfePZFJg1xHH4bkRfcx1yzhQUrOszFpg9FSoyQ7xzlPfHphc9gaIkG
gOhSZ/CgfP+Sb1YCCGDxKm8sysgLYNt+JSpmbMZViuQ2M8xBxG+TEyNioOf44uz/OC8UzWP6LlMW
9gxtzjHsDO1AC9Lipo6B7xLLKSMu21LLNUWyWNmW9d+d4LXo6q0Zpd9VsdMSm2H0fGNyd/LpCsoc
ivlxudKDmDCGZuTnL7Hjixk9iZxcAzWNOvdrcYZSk5sFLYwb//Oetn1I6gIR5h/MM/Un2M0u1qq8
0TgiUeCdPENnnNTDCWlUqexSd9kFr0S6tENKropaQAXJ6X6QDX5cYXBy96aUfqj7fHvtQBFdFWV9
dcG4Fk3lfuqP1ksTY+0XtMv2dFZwUNxlOGV6yoY7egri3prWt00jaPiGkn4jh9quQxnugEm8TuYk
2TWPLde9vTAxORRI6RHtTyUjRvs/VwWkMYXrORSNlKCQgbz4GccaKlDLNsB9xb3hDv25L5jMyzMy
jA9JMtEvwjxcdB68yzdKnYT6ZVa618ZAiumWbmXZSGSYMBZJzSzsIAC/ESHsaBUcmPY18sGxDmC4
k/q5hLf817weO6m3FWGixj1MshhxYivJAvY75olVzfh5k4UQ/fS/RH7+V8x5XrVTHgOPeW9e74R+
vCI9nxEmYI6t4ChLfSg3d5EapmrwIkxOWJUZNwT6JZaMTue6o736HlNK3RwhtHVTPM+2d6p2+ZHw
SGoScSxQO6ErfE3t7WH1kvsYiljxzGFV05Z32BC89tLswF2cNzA62fxF9cPPGu1+bMye86UZkLJ3
IAhfUI3JssD4YtuPjWKDKslI3wZ69LE52uYJIxLNwXYY46vNcjvYZDTMhxErsOaC89gmGgo47lgw
ArPS80jf2ayztFVeAOwMKQIupEplHSRHZgElM38h5YBUOSEi/tgVRxzSpz9c2e263Qx9+nXMNvxK
tQsQis/or2AZ0ZL01ZuW2fxO3fBJ3ROo7C34rk3l9+gKQsZppHxrwwQ5d/voa6uG+TkYs6jiDyEP
15kX7qL8iZ3UUGUyh8q7fkxc4V2jByZamx3LpWCNafoiuia8xxvIkDA2ILgXRkfnWXwvsioqvuZ/
PEHMEqaxStFZ73OfsuRj1gm4RTs54FZRaU3Z9XQXkdWQ63oeIxUrEk9oKvRDXcf6Lpgm/dsfv/yL
ZaOvG0b0E7vEME5uzQhk8UBfM9WFWSBK6MOL+kBgtP0FhFSmDJAGOjkz7LDSlKmTAOt2/5mFzj58
0BJ2Xo8uZ2YERE6QPxQzkcL8D972Ueq3qv9X97xEe+s+PhyLJlLo1W6XLqXqHJOyDer+Xulx/aGM
CQXKSwsGeeFmIHbyilHIK4bAGDPg8PDLsw/FwkeFd7M21wmk6qUQt/GlJwkrSBxRm0FrJFCUOcQE
m7jyWfKZRJex9CESimR+0KqrrynZqRGLw+nmOUP3LRMfcGr41ofVc/tA2bz/bxU9Tz4ZYruajMhA
9ex9deoSUHMq10WNftH1aNeVqrW2UMC9qJRHwMXrnHFv5DoyzkBmVRlBrgX9Y2EcwtopVhaaoLMD
2VWRBAnhteaQghhc85+82NWODVUFOJqSwDghRZbEZNdn9kOy7XKmRTteDgy7aPC0Q0JP8WyjhYq3
dGOBBxMDgcHW5ha/6HIVM7YmlUG4aobtnUVloHGj+x9UyvSkYiyeeQSF5weYtZi44g9qu8zycUGl
av/1vNHQGTvJF73PuMZvYuSUhkI6dPMpQVpmY2i/sqHQ7n4cD9DxDYz8bUn068NNAYaWuldehtLK
u/yLj6mACGJCgolKq79KZYtirIa9nuFH9Xg8/2CfXwovXv6QOx1zZaBRB2RBj9/Sf7U9g3eum4qX
9Xc02OLOUXF3rZbhEdvU04IyEb7I3YJmh6LDwmczHDj7IkYw1u6m/V1OmnvoWIOT6yiCTE2483os
IqX/sEF67hyoi2jHHhlIouMTVMhxft50BXPwGdbJNT4Ef8Kj1o9jmaUoX0GDlDKkAG78WmBEHAwc
YqVGAUUZlg5yp8XRDtndSlT2l56phyG8Ozj/BvoyMFpZhoDjn7h8qm1rDHequDwIksfauJQR9Iau
f/mEv21k6hcIg4pwk3ORRo5o0mpuPtPlST+5WKg1u2I5/sK4bcVqIjoUzpl7Suuru7twH1K2eERH
4il3dgGKwuYgKnD2HH7EAssewG1uruSVISYFAjI7GpOmQ+rE/LkWFS1529ll0uGzPaZ9gl+ANSLw
DmjS2quRSb8PcoFzC/3KUvvx66wQ4Athmzaxa8kxtxd0puQ6WeM283pAlx8DgwbF8W3JZakKCtkQ
z4ynOrcL7o9qjp5Ns0Ztcd/KDF5kFoakODyFMkKHeijH3jaFquEvp5z78iBzLGLXzsE2shbor12Q
sc5V0Oj1qjGKnumA1zgk4KAoxb/8FpJO/Ad1mEj2AaezMx70J+ln7utLR5kESs18c3OzEtvW+fom
psjf4MG4S4pExvPeJkqTBnxtmSJygoULcCGianrHwON28X6wdwQMP+9U46phJCWQwNNwUX9I7/H1
p7DPgcM8GsQ186jUPv1Dat/PXKrt7HNqTmQ/Jws6ub7YzEz2ZTP1m87PMXdiQlzS5RA53IggfX/O
huprSQ+zA3mss+JtzcPV4o7+SJmSDjIuEZWNHN7F9BCjlyM4WPO9nwGId9ifRqRSuvPyNM26OL9O
kf/SpkeTrnfwIebwzHCiX7ZnR3K2CG4CSoGqn7f71KagoSpDadp5OocSaXZcnYoSSFPqVjTAJZxG
sAFdGKGxK8z94iCFyZ1gZD0bSEwlG6kyZJNuhLpzJyx643GujY+rgQ9NI9/0CJ+cbZspb2ciisZ4
1dJzHTYeKxa5eBvLP82wkkvim/oIFr0MaIzrDeO4bo7wNW3meyukP2CSvA4tNjGe7HkD1wqFM/g/
tlEHXD154ZemkRhh6vSEzSfAT3v4TKlsW4Lh4R6JN+3isV6qBCEwM0P3vRSTbUHvPDzQP1D1RzGF
sKlNr9vfw4sqipxM+7bnHuiwbWHnbAABTd9PW7aWlLj3A+wGphh2/Ds/R0VxSQlUJqLp2Wxs3uXM
HqfvXxRVX1sN+YMxiOF3IFrh096CU4qLzVRh6Bueqdrh5NvLZEvteGKAaQo6r+90LXAhQY/Ii9Fh
mpTFxhksq2ebmFf/kNHuHmo2/P14UV7AMC35oouGDWlvigkauWsBgyg4iUDwiQr7BIqXBi3MdnQk
Evo7V8nx1Q19ZxR+fHFMoneNc7XFe5h+0ynKQdcXRqiFl2ab9/ubHyrZ6I78d7VprURjpP2narD/
q8Q1+mcBNpSNIXGSEs0OtOXd3KhCOFKNJ+Vfv7jhPyvZ0aPq7k6gB8ocZ6bIJhRANRVN0J4sM8F2
J5FhcyKZGZGmbG2XpixLNvzKod22wloNNEDMb+C+uYuzZORPzl1tSlhzE7QIEzxxU8MAJpa3Z5zQ
MVTdK32Jyj0r1cBdvOSqsx4af2eyH8oz347xRrqH8hD4pCQo6K8ldDQJ5Z2SaLLnN6bfviI0jyEs
zPRtqoxyyL/XNwDulYHQIBLEJnj/cuE4nR6dmPwGVvJLhzgxgcSEDERPxkeNKPtCZERq4OZBc85V
JtVXlgOItB5pkYB19RStdrmuNBrCViH4/p2mFWQ9axuB0dIexL9FNtNRyPQTLumE6ICAcZjatefw
WdOvQVhbqlcE+C52C0elkQ5xGpRaip4eSTGE8V+OhJJkBs2gdkzadQVYSsSD+dw/SFK0JiT4lbnp
Kkt1XeR2lHO/nWsMBKunWppzDrgZSESo7IzlK8S805MQmEWgXCxc8s/PZok6Vi5RBv+XxmYfOf8v
5513tguQki01fzuPl6tN85UCpZ0rEne5O9+7Yb0XoX/cNUrX/92pJzIT+H+uJcRpxOP6mX4gr6tE
cRadLTbXUNrmV9j4hzRMXXjvvX+ffyjXObgGUsMG9E35gwx/zwj6r90KxbtzX4wx1if7s/k8a2zr
Gfoi9XQXNweGCAkyddrm0sVmql2SAB3lEoEBobMJEbZrTEPz50QeftMFDwZgf1AA2llUQdMKXV8e
jVhUFHWsYcYIsEZRRnD1WzT1WBUR5eXMTbCfLyB4HwSNWMYxhWiI9REyhEB7XlMSSyg7B+XaRRVU
pq7EuhhMb8KZd/4JQvGWMiuj/CBJuE61LXeK3OF4ljsW33VuaOpdX1hTxF/+NaHtRTfMgKsvKrQW
yUxZl56xwDs61yIUrgrOqi5+/iQcXDnzFOyX/w7zslM8agswrrsdHYABx6itt7kNP54gkKwHEKqG
pm2Krg6ZiXT2yYiYSrGjPIPfisa9c8BxCoXnyNVooQBGIrRCIBMuM0q0ycoxWSEWYeYoqeNByrPO
x53KutvyK82FEub4tY0llZ0LalAPZyvONSzRcG3V7L7CaD6v482oiaES41BRBd6dhawrsFvRNPfY
jnoko+gmflkWJkv6PbIDWcCNz04/0ZyOyw/xtZhGJnhw50cdclatv9Ptgzo234XeN8nbW4Opu0UW
JU2ria8gYS2RJpoJLUac/7KBlIFsU9C31yDtDMO39LnkHRt6PtT5w8rYqOOfGPqgFq+m6s6wHNTw
WMpNiUgWczxNSVbs10GWyN/rb/bm7DkpateYQIQDty0PLPIuI1Nd5NRocLHfQ2gGKHfJO6Aapuw8
AKvk8l0syQk/B3Qh3c9eRDxc5StvnAjRubwMZIvG6dYy+7Bo9reoaI5k3lXcjL4KZx+e88XMxpQ0
0oLbahijpmmG3a5hg4Nc1NH2utMbLSxJuwmUNQCLsK6qgN2dt5NqZqUTjhcbFTHlCN7b/WSEtzGj
h2FRkJezp4Jz2hGVQYnaKBYXIxJMSRdQi7lMSLc26vlD+O7zpF3xPPMZ2OrmTQgv30HTMl9BCqns
/OCeCd8BEx7o1bQ19qz6i44z1OwDClojRjYJSq8D3K0Lw8v5lyQO5yio4Ubc3KMEVjNyH9ZCoY+m
HQtQYJbzuDZRu0r9XWnWg8MhfK7WoDbvdtfBUbnJluEQQEAVL8Cpdia7pr6Crfh27K8sT8npKYce
M1T+gwp4eob7az7VirWqykOo8l3jPHkaDWF4kmrCRy1rEJPXGOKU6PbAlaWiT3trjryEPjVueXg+
oLnAOG4RHwOhOb77E2SyocogaXen9l/8qlLY6QSvwaHb38FSgjypqoUUklOkG69P3Vfezr/MfT2/
1xK7vFFf+os8bGMVrbNh+Ayvhaha2Dcb451t9S9bOtu4La2+OYlnsekBkc8wwGHukWzBWHp/ycBj
NpGtLh5v9Z5HpWzJ1frTKf16B8Ay+xC1NuPht1PQUwVN07XqgksA3x3ZZW4QwOiqXcP3uuPqyfxA
m3oeB2lwe6s5GVKqY1pa+7aD6+dwKvYD0wJuDeJFnypOLWCHNch5ild6hvv3j7Y+VNRGZhu/sCCh
hzlZFxkkCoeN0vcBi2JH713n9lGd8gfqwAAPZWE1DP7MFSNL1u4QZzEWoTUOK8k222lTngQfK1ky
/hCMa48GqRcLZrflI/t3h7E68bMZPFlHokx5cEL+DwZ56fyQ3eMQ5G04r0ZPA7N9GnNZV9NhpgSf
2qq+1v/upPYO1T6BRnzQveozq3dYTKPUZcevlL6q8C8d5S4wl7bEmPEevoFWzCSEk2S8klBMiQ1R
JzRSrKTKxPDBKqzNLJP+7/NE49cWHFncdbrnzhAbZH1njBQFobhQ5/ym/IaTivR8/g6EajD/oGBR
TmzLb0JgK3OpCfbcCfC5CKaKIH2KAImO4gz/tYZBxYUMxaQ9Sof1MxJyGiI0epkMCbLp2EMxZG9c
VVmiK69RVZVU7cLLg/tDBZ/hNPVhxe52jpdasMfpdkSrSsM4GegPZM5TsEvyfhMiUkY4QVDh1jYR
TmLaak9cT5YN0y/9ZCvNxJpVRnphuhTXPp4bOiM/LuifZWOpcV9QlkAM9FWkEIV+fMps7nJH5zjT
FzowC8UZPjWNzpg/fEise+pk6Cn6yo/RHjqU9u/Zwl7wTnrXeeofoEF4X9J5/36m2n3/a9yoAuf0
Ilnsd+zhtnZbByvOaiTah5LYHgDEYML9MKeRKVBsXl+JROA+pRtm8a3V/JhmHRUQ2C04ecM6rvV3
LRpaXI+MH7pF2FX8kwZPQ0gAC8NmVdYANEDZ+gEUM5BIBr65nhcbgOpDI/2Dojne2HxNLOd5x2GF
Bb6TkgaOZkrQt5okC21yAM6QBravZghVVx45R7pJvoJi1rqifgMFY3dfiDHcipNl+vxZnLWhEA8G
UkL2RWIV3SiCN3pb1IQ404z4zfQ34UCXaSmFdSShsSBJhXbh6BgtFgRGE7Rr7QIAlVuSgJRxUFqk
GjQ0ZpSf3Yht/kbgZPXOYF5cD/TycXnZu0CLUv9/4GS6iUvYnf2VoZTxXV4n6jQFWeTY/rZgRnVe
+ml//olHWxI9z73exoX9+beRn4q1HxevlEnXPwXQa0ge31pWVLOZo9QgszX9/a0pPmGUFmEpp2R2
5eRs8Gfz1HDY7tgmkhMPBJDi4EfQ2XC96BXah3LzI4X8iXvSWsxgyzttyzvHm1tFzLPKPQvNbvAR
VoFkC70iC4zCAhukHhRhIFw5yXZLqXbh6QIm2zSJyQgKVNSFw/5O9hyXH55DNG8kwmPB7V4quiwO
T9L22PTei9tWrTwY+uezex9yfs/kc5qrDOjlMRldg/7UIII68eUdLZ/Agj2UG8vJH/LpinJU++0k
1aDHx8QQQMc7Jr1nnAZ3SS7qfb5ui32f+mV4QE82R1D8Zg+1M9Ofx6KKvw66Ti1S55P+P/kffZ89
cVtOw49N9BbwCpABArssGb/0mBAteE9dEVuu8UQoQDdAgvi/aiat2Y8EY6yp9NIOn22kn/JeeeqH
mXZvhMUCKHHQb8ft/u/NyOOYTgIAh22mGmNX3IeHac1eBoBuOxNA+k3tY2Maox3Toj5U6O3GkLSa
Lyni4uLFW9vV1Bya1EtKKe3gNTmMRVi7/Ue3uxeSc+gUZC1vwnpkQjWR7Rc4rl8623DzCTqMLwoU
XCRD4zWhAHSk8KUqI30jpLhLpYoTtbRaOCgK6FPkzG8YFJRAV+3hxx04sA1t/XAa80cUtyQfi6MG
W/DwOWnOQMX+X/mBxp2355FW8i/Ji9rBUG0GRtFQiZYoTD2EEV3F6gvvX2R+RK2KpSi+5XLeBxen
Sykpex6l111S7SzbTKqwsZptr+eXnf2gWVaowcUuuxm22DtkBM66lTOIbZ0wYlILRgBx6I9jW1hQ
WSMV64IgnctB9S9EKvPHbYoM1ziqROn4jPoV5HxknjrvPdF55tvOLybltAdZqPTpVn3wmb2STUEO
NJgJScSUFncvi7KlkevMvzmiWniw46mMs1aA7zFSRaTL2qvg4nhOqdPFkqu0V7yQlu1lhk5j3RbI
axbpLzVoCzmoIgKMZHXKvWcJCuQmm/3IkGTgRP3AF1UYzFOjEkPs7HX5fyTuxVLCfjk1A7sYH320
rUN1O1QTEk3agL/q9ccOHmcFHpc6Og9wO79hc04hWyweg29eOExI8R7vnLXg9C6HG81i3HeqSTZv
gzl234R4VGkEPRi3i2rDHGUenV0ulzY+IF7bJfGmkWUMU9luqPSZbx/sO4dTjBrUSAUt5fjughmS
5hBqa6eR1CKnWexwFqPklNIsgWh4YudG3zaycM7w/3aMiaUNu3F9KFKjeEmjCYeFcNX27+zQSM6Y
//frgArv9n2KSmzQOqDr5fqTlfDlpoIYfYCnFr3SafBR0GJ6Gud6zL0t4n7YgpAnoKtTnKQbatTD
G0mL2zPBTu/DCl+Nt9bqdzHmLHwEvoHaxZonWpAgt6oehSwJfR6X2DgAOFZ38JtSAC9yEeGFzPA4
IIRJ86ID59zLY2wmyUB9L8gUhXOmpU3owAKwKWAfskPK5FHRop0ekjHvGpCpjBcMTP/XUMbJk03z
QoBEM/GX9CE2utNByhCwosAVtefwFcyQS075kSkivh6Uk/3brzH85UfC038ZmDtHrwnhU73Tbia5
9e2uaKTbeElDk7YEvVxRjbO8fbbKk/Ca03OF9oVCP/Abl9YHmyN/S754Ow5mepGDv8U/fAsGZNqH
+lR+vT93p95I8waDs2wyz7jv3HiOHczOxk1NxxkAuKl/jA8bmiCQnnjH5r0esljvPeP2j2d91irJ
J3v/nccS5lLZsBTLQATULqljNf25kB8mcyATLL1A3RrM7/Ue19qR4uI2VRvFnzEM/PO6RIlGTygH
Y61IinGqrfUWghfixuMpnbp8Kif4WMqV4tdvN9fNJbXtuWeNjofGQaXesnRsx3M62xHR0iVBbY0k
o4OYVlENcK7EodzQ91c+qIvFDEBh7FuUzovIukU+TBSyrGZgJExfA8zo1qqV2BKASAZIYLPtiZH5
BNdtUE2JV+oOCaDZxFE8Is+zgzCqldP+hsag4MQvQAxQ5sb5yvhZO9oWx7BZVzKEA1YZ84bSBHKC
Ms4RwLrU4Npe1xP+sBWT2ap9OzsNWFH0vl/SLusve6Ux3yC7UNjOEnsMxM60kiTwp+JlvTKGMmam
la0IWRYQ1zPHZ8bBfpxkpOQ60L5IgPPaemKAwFRviwMcp/Zxma55enM2Ii1fdE4wc4xk+HAQeL85
7rmDFoqUYQQTLy+/Gh47C1yIWThnT5l0eoYG5mMgXrDBVbhWHj4r5C1EjATLOV4VdSMC4MMGK8wV
ZhjWSZB7Nh4keaj8YtJXrTNEC6SUJbmBeTN57J/GscSKkIxT3ybOKw5hW30eOhD8SH+ZTjJyYI2p
o1UF9RuErmq6H66zgf2GgewKSeW40E3tstnLUke2o2FTAAEPVW7IQvUD/tukmgrLsGmwK759yGct
CA3wNNnEG5j+Bwd4o/Oi2tM2PLicAzVC3MwHBRfkB2lp2/Diev3go3iWaQCzJtcPtPMKmjdGiL1B
bxf5ssh0BpoczKPLCwRk0NSlGUgzvD+yrsTIeDZQTe6+UUN25O7vEK8Ymxn1f8ypliO+E/IQlbMr
/8vYsRCZrFht2ZNFpnPEy51QUANdeh2+sn+P68IBhGknRArxBjXN8d0zQ/8a+AN16+jlTpCzQUck
mTU1N8rGo3cGXwcf07OmKcG5CPMm8rErMVO6lEEfpuGNGgehi4802uGO9pkgvn9OOf4/GYvAuFia
g2Z/du85w8Wm0J2PlaS1jj2wiYylhx/tptz5rFE6kNpQikRQMQXZvUyfpoMBSPfW7IXxLDy9k8Gd
nDuuPylHZ+ld5fCbx6U9xExm6ATMCFUQY8YtNEwSqXN4ILCiW4cdPDdYDm3ldHXd0qYvdNLAq4WX
dPm3xRyvXP5SBKZv89Z8tJOHKPWaUfHwGgeS0I33w3Hit0z4dcKkCyscd/0bILt+KjCDBdViudMR
+TN5eYjkgShFZ3IIMUHLQtQtR6m+BhnviDbolzn9Ps/AlZCrJouFskGsO/+fPcwOmATTSHmE++/E
pVVSVJO7Df1TR88Ez+JHcJpVswiYTG7sXBFHZphA/h9SBAMKNtkBsYv3RlWYfuWjRrwdmA6HAjoc
30LwpLU53264SEPo6edt3pWl8bpxlM65EqMac5AD7mVJlGxfmdC9XxZhdhSxYLwkDup0bjek4NhD
ESzXyvKpVdevzoXyUaGs772qrP8vE7VCt/N1BHH3YQRaiToVVdOU2mcehDjGqR8x/MEXNWKPgr7i
07YuDz0OdWTu11URWumhIL5PbEdHIYygJdDTBKHsceEWXQQcCL+qTmgvYsipllPDT7C4DDmHt93a
FnsegHDsjnRE93QSmfHB/Z5axagHs+k+4F8nJqp8SRszTelUsTIALSrJT1r9ymdk25S5upmlrW1u
JBJ0iliGNl2PaGNz7uZzAfcUDvHIPrGwa9S0uYPdnGS18oLdbiBn41oS0Q29prGfOePBfMWV+4Sf
Xt4NoG/vkf3vMrD/P1R8yOlf8fUDNPoHQXaeDUTbFUr+ukAsAsiqDYnlDaJbQO65ts59eDSBFDNe
7E3TNdrq48IywnplaU3v0n6cH5J3W6o30YUguI0nS1KLNwpAgx414b8EihsvNqJi0AQajUsZqZMB
1C+8ImWl5XCVC9yxnY7rCpCEfHeNYYlC/nzAsIoiKRjfGHlhFXkRSQfX0sQJ0fdp0YECjfhFdjjB
9sk2tV2A743PJEnAP8mbkdc/0JpKPtsuoyBIrX7EMrYOL5QXw1JBldxKhpyBgDGUjvYzAv60zWf9
c9Pe0qUv/dLHd2wQiQf3iUwTV5sR0aHkJ/FmMTfEp3MtJvzyYhlo0HtZji03iMWR2mLV5kdHtG0Y
KgEFNM0JslgLCiJwKv6aY9rdDR32ydLAOsrynuXw1hwaYbf53Unoh3EYJqtYUoj2daxHyGpBWLTr
liN83tbDVF1q410IasvsPTmd86mDJUzkf74wn5lx+JkRoPmoWfMwZMBV7oCDl7qAmsKv43YnXRvh
cpnmfnYWAbQYehwVBSB/zYI1DqIDWeOC14hMLej8MdfSJSujEi+k/jtHWz4gAMiEczxmRE1gVDy9
RvtHEe5Pv1ED8ZPHiCViTxx85HX/4HWorZpX8aTnWYF8LhAlZ2CE0vO0aj6L4LYc0UFtfU59XNWY
cKd/ODuYz8ih0pcaRa1nJIIwhs6zOVAZMBpSOM1oDEVnSo51EXoxw6g37J89gXPd7RNPJABfLJzJ
2lRzuVPCD8sOnzQ3BZGbf7oa9N1KWyksgVcZtVlgCyCnYUekqFdpLme1sa36wf++LAZD7cWbngVM
hG6gY2D9EZubyMCYow1Max2BlCTbd/ZKczO76uBFSFaN1b4oR2cMAhfuj6BuRj69fGDxjsEBqgFJ
ignrDXWvoQ7H3AWAldAoxgY9LMiUX6zKSH2ICTT75tkYCXf63ZpaYIyEU3faFRzg17KTgKkqeDgO
OCB3SJpF8J6vBPp+RRt98ZfrDSEAIwh2vlbMQ2fHY9WnAFmNkPTvK1+lMHRyX6oa0cbUzDVQjKWP
vbx4qvVwRpTr0hGEtHpJJB07ld0RNZqEfHBn3c7Jio08QO1jPWu+2+srzrAgHJtsfvNzea/3It//
PvnqMohGXcOYgr1ZamnkmZ8aI3weqBdcbKShw+jUSkVVVeJyHKyNunIq2zuoHqmg8s6L6Hg9xG7l
zlEkzuD2dR4mcxtd+FxYQChNH+IOZYRi3HaYg7gFBsAeQ+oc6kEGxj6noXT1vR13rCctCDIBbqwB
wYxmxe4IQflTcFkYuSMkEKvZk9nXSuYVE9pJhtbZbeLgZtblxo95Jp7SGT1P8PYvm5Ybj3qwe/nh
0QrPQVqSU1gre6bwBffPfz0tv68Lbfnndzh3e/y3Iy3cvhZooVnAqITGCxQnvff//eVWOWD/hbnN
iRt0GRYhjp5+Pvw3Olj4hBFASzc5360614ToLIg27JpqisjqgdCw3g4F8PG6ijXd1f5tFMcoM/cm
e4uBrdbHVDCeZgacPwftCp66cFiwSV4Xaqrp272fDCaWQlZuIYgWQ0n+b7RYB64hTlYmXUNj8iX8
OqK/Q20Grx/zt93g67B+xIgJ5uGJdLCW7tBPCCaxQCeR/3ZrNS9JfNFbnZJ4X82yJ4v97v4yxF1y
iDQc08MiggvFRPox0G3bdF2IvUXtq2k5tJonFxYqtckvj7hZI1e79ZTZ46mKX2o7EF2ZujB1cbye
wTc1DKwLY8hnIY77G7z2pKLPme1uAJZZ1iwBKBsRUdXQvlR8jXM5jfC654W5z0iphTdeAot4xNI5
nIf0Y/6ebKQzKltJ3B3gzjGsnNiglG2faS/HenO3UTpMuWk4YZm5NV1eVwKU67fjR5Oo92OQi5qd
6ZgsUoEN0tDhA4LAQpTDVY/qlow4YPR6SvZwBWtyGju3E9f7d6i0ByBUYbO6dV8FDO3R78puWi79
3jCXpuR2FudoOKJ6KvGZAeTgDOaR/X5UZj+Jmny6TBdIwskOOGR1joI/yhAapnwxtjQL91RoQVg0
gHGkQtR/+exCTGqDB3GBDykzpNyivxFBk6KI5+Aw7ttMwYacImqsEeKJG3X/tR2IgRRb15Nb8lum
rZSFDxBFDGesllR2h/v9Du42wkEt0Ru9T3+or5UZYn4FbfQTZkdJ2VLBa/Elm8FCchSnKDylCnyt
kElb5uPOuNiGuAG9ynm0SQ6yrgFhYTw1Pc0o8oWq4NKZg7AsknJXiIfJxPX0s7M3dBP0H37Qa62Z
tNoKIBw0SkO0IWdRcvYM+s8KyKSVJ9yw0pRKux8GH8cf73/QAqdgw6I/Q6WXM45u5pSuidK766J8
wbzZr1/epA1jIz50xaOIiMiCRRPuTKacjqFtIa/zZrIj3/z8LoBBAZc1lhtgPgRkAJuP0eZ0DdqG
Fl2VEoze3Y0rSde6SCfjfzz+e/nHKDmIeCMYcW1G0K0JwmliOtEMJgLsRUA4GDnngbAdEJ/P7MSX
6FXSmXLvrPD5oIsdWanMV9OvKDgETRS8Qb+Y8K3bvRPNeo6o4ArD63eSYZ8pQvLATThgGM5wfR2M
A8H/FivjfV9MAvKsTmKVeZ7yjoO+BT0Nz1M/mouSiBHIWGeBfFMzzxvbHFuqT9C0I1kUftscDdJ4
BfWK9R7m/r6xQ6KmuSzcsLalITtsxeE7Imwmo3GahFntBfTOiXcMSRjMVYdMkqVg/e60b+hOOris
UqXtIEDg2pfoRXXh6TAIkvdxY8m+grcMcu4aUloF4H/9h6coWuAR7xflo7gm0M+9W7nwPrUPe5LA
eVCbjVNLTdTO8548sk+tKjThve+tPQBWJxkfNd5CQufXGJRowALifchsz7T24s7rB9DDRWG/weiy
LUqShtTwvZ2lmeXt0KmTvw6cuG9cpuiw2fgUxaYeJ6OaqSij89RCAq/z/zI+1kZsN6Xlbtp+kAC8
XFBlCas/XLy+W2eOwZNbbiPx/tD0jfEphPvoisOyK4zY1WhqNXcQG4aI9nW8BtY3WwdS/n9JDJ4T
vxmu7r+DM8g+aAr7gi2WS0BSGOuxgpdr6Vuyxz5FKxqHhqAbqkTKaa/Eco36plBpirBwyvXHoB53
Q0WYaNPkUrUSWiM9To4d6K3dEbx9y+S6QlNdb6uwWjFVJNuvRXv/dSAGBuabBDdkE1MAUBtWZYOH
o72Uwm6kQmYaPpjgMdIzHpXH8mfuQQgEra/eNP6gq+N7m0bzJ4vXUm0OqhiDjz5E8JazoIypoISX
wB7pTn/rmLsViqyVb9otH3r2AxXYP0xYr/tO9ci/jn/pp0iFbDeYFNCaJhJszEX1PYqtmcbT8khj
A9nIh61ezJ2SjSHkZST3THlNbDm2p8DCaD2ZoRcKS3uRmdDt2U/f/Ilk4v9c4h1sURbaUDxy3+Fy
Rj2PXUu5C2SgA3drL0Zco3/UQUe+rv5GvCWAJ5C7o1jWqb4Tbx8t7KcZXbmd2fRlX4RuEHaeoCVk
DXKY5riiGPGszYu14pxZmU8TEpvKq6229X16Bp8504oqsPyu3EzKcoHMJFRSi7RQQ5IZK9Ppl5x+
o4VSO3QhDB95p7tR/+/b/t+PLWBRw3In7g6BwNsY1rdXyXbgt1VHD6y6qrbwVnDjUm9DkeHRAqfE
C/1yUo5qWkvmQQHLg4rycLN1ESeieNnrjzFcC28n9b4DrSM1FDco4FRgZRSpH6zpnC4ryUoAOdiM
iudFOw/4MhV5968ps3CrpShp9fS8/8ASIvept1g7qJjh7OsgQo/sSCVEwf/o09a6jxXFfogWbLLo
sSE0JbVNeuy4FK3ljR0GWVsN3JEQRCNIddiphZCpklwgeJrDIxEPU/q8HLIjC7swNrJ5YFFNhWQq
BM4MxNwVyB7LQGbHlYM9U2n9UH48rrR5/U9audSs8VjtgFv/shGBhlgPhZl1g3KVK+drHxfPSvKp
pjB24b5Ob5Ug2bEAUv8CI/IDTXSvqsD481hizPiE62tT/ijdsy1f+2XNkuPFxYW6DZ9MCupBIH/a
3z5dkrDj4qmy804qTK+saMle7DLRI9FAKqgfYFBKAL4wQUcFi8WXVq0XKV5MZyXT2Qm8JjxcURk/
BOs/MP9qQyx4wu97V9GX8/pih8bVxX7z3odOQtx8z3aJ3vs1eO2CbBsal7DZ9BawVhsk/oP4jC34
dtBU2tW+ol/DZb+2A2cZ2M5qpQGQOuLXHIcXNtl6N/jjj2ye5YveJLs10ehIX70avgHr2W9eQddO
EQLQKIoTWu8UxlumsmEGSoNjDhnjqFU0M2+66hFCE/Q7FMFyXDXuf88LdOuWrLG87AKmyNyrLXgb
XAEfgoBfTDUNPe+4SobW9SBZnMWe4tmGAQspNVJPrPEx9jCShTM1HlnztGEqcKchPeOhEMCNvLpK
VJ5kb64uhzP5j12QWYi3XtYfmiUHMJE8W0o1I+Q6yY49GYY2X1kwX59JZaoaIJyXD5Ryri3OHDEc
1ZdVYeiSnbcMb1HO3Qcd8L1JXejGHcgURdBVKpLow4fCIWDl/95aXaskQAY2SED/KAA2Ujnk7RPh
wQxoUqtkaD3GNYDmCGO082xHB7UgvlCCq6k46Diz9S1JEaiD4ZY5h3Q9EgOwYd2wk6KeWvKaCXMm
I8pJBmDY2GTBDw/hqzlcMBjHO30tOrxRA85UMbdwV5QqV11uX+MMP15nOurS1PhtvuDZKtjd0n3y
K65RnmwrtCGmbUOm2rp6/tpFOrv4P8CDpYPO2JL9yWZHUPakuJbygyem06sRRM1qbMXPH++3tVQ+
3oHWC3MykpkcNanXmlHjJ73wGLdcU+FEpYucCyc+614KKYPve/DjKbgop3hKeIev2GH4cxzaiu5P
4X0r3rTTn5T4dh4ChMGlJRQrlJdqjxN8NFoPnKJz26OIuR201kLEAGe1zYQSqs6ssIxYtjsr/X0o
ApsfzRgkvI05ehRA563Ihnc8ZR9u2Bp/X6xfP0P4bJJ11mFnZsoaQ7N0S3f5JDlukJCQsy5YUhvB
XJkgsJAUVJhebMIDakf3GxZjG2c3HehLxRLN2b5fb9PwvfgxjcV1paYIsdHOIYUVYkKxrf85hvHz
LfZDEOd1BpvI0qjMoBEDHsPpD1ym44gOMPFS1LdUPjlFM8qG+gyaZRYsi2R3mNp3kl+GQSv00xaP
Z+eqN3wbWDXXiKn6faWesmGRgeswz2LPmEBY/R9HQBsNYMCzMV9qjfYHIQLZsWmd0HiVvUFRWh9Q
ExWEHbavyGJQH1JgQB9sT5gsYmde/cfJ6RiimwMdOGPpz4MCMsfySapN/W4MnlgS263NREJ4M6Bh
kBOlqwbrxFcbKz/abaHKTxBadkIYvh5r9x5G2a8QpnBTmx6/pzTeHBBbHjjoo0GHiFxbva7hse8l
gtnGNb9uNu8c8DmhfrIiX8l5bQXKpUIs4Mtlj4A7NumdiR9C8dXwjt41tDSzfYOR01LgdGUS/Doh
wSmCUGPoxJGOsywvVp734Z+ILxM+3mcDir8DOY9WqZQ0dowlgZeqxzLxU0RGn74HjVQIi4JRNQM4
2nKvo8j7PAy51yB0yF6bNuyoHdKb1/nxlNutKpJH08jTfEyBAyPJrPPDzMG+/DHXwG+by8r7scoe
QBzmwttmi0lq78/dr51iL22hQBe2t4H20dAa7YI5CmrP5Pf3zlFP83iDFbu9y/WrtBwJjkjAhW4b
kMWcxFKrDLlsDAwu0PyF8v1NJeY7iXe7x/F/scBccwwrNL05kOmi78i36kZTrqyomsNM7CZncoFZ
BvrxnQZqWXZLFkr1qFpK96/pUtRYR5DjK2qQYlgRK8aubeWqvtxWYMg44pTEq1CMVi3qyWJcKefD
e6JETRN6S8tHYAXbDzqpvQY+RtuUY/6PhE+KGzl0XaIWFXIH0yqoJhVQwa1wKvPyiEIiLdML4+A/
nRMToSQdGoHwzOz+CZLqGhg3b7ImHeIsxxElwQuz3buWc1Jbsddf848+0rXW+20GRqSdNQ4IYqJO
Kpa4r7aNFqxLlYSSiTR8unZMB+ietbNdviXLVFHlsDqORwgRBEFJs1HiVz8/9c7EkJrE/dA20pzk
IoBouSfz+N/XReIqXSszQCVcV6FQlyCWLLQGNRyXA34becC37SILWbjKfwh5lBrCEMZZyFxoXllB
o8PuJ85ZUfnmkwxUBU1l1U4Z7/h52J7o8nLI9jmM5ZvHETt1SERFs3Zlbvx33mijnfFAs6ji3oRV
IGLFlIGn6CNGNOE4xrvlM/0nPpzxXuf0bh86/BdMxJzRlLb2ONIxpMjVdFArQVk7B6i48P35jwCq
rCMd0P3DLwBuhPYBZ5DQMy7mb4eWWB8+9BJj4zJb4DHyET4IKEr1o0OGkXbitSZUME6ScrqrFHNV
8gkl3AOpLyTruRo8/Ocyn7oHLQxI/bjM6l+1myIog23XSBEVWxGHLLTdD/iFEzlsuQWpxSrmUdd5
GL5vPCXrHpfCmxIDEPqRRQULkTdOKYB+vdZBX+mA/2aDoOJMhhi1uoYz4Y6NDq4dlhqUltEABDU6
zRb17JRd69AvVldU8oDpacYChNuGb/f5EQl2qnVQ87ttR6uaI5JUF08bP0S7VBKfv5SKI8QJVm2G
CpLBKyqYbUqJgItGcQhaBoxZnaKCSa6VOwWxrynv0YU+SlVXv4JMGKS3kKs5tTwADEIPhjQJud9C
EJtEAXaswFjP8vzbPI9iO/IIgByv5kZfc2ac7vkEGWNLOwxNapkQUugIMMNr4NHWNGWU5GW++5rJ
GxRPjfhdMzbp7B2E/hW6yKA93HZiWwJZiSoOVdb9cThAAwTeY+u9MGqTURY7ZJkDh8ig9TRa/zIW
opLCmX6uK0xUJIe9ngY9Pn9Exw3QXXzai/kRTDGKvzSsXPYMXx0dnKjq1pj6STzJspo2ArZTfXps
VfazY7Pz8bWhNUNl0eFA1Ch1ljpRnWnBLasR/3Su/fNtXC8dFHXZRpOXHrg7Miadjdq8NV1UdIC+
AM/X+pIc6USrrfjpNErbr1sFiRAXQ6jvfmN+QpveT1YRQ9siiKHpZeWeky/ATb1s1wG//S1n9qhB
YghExfy7YxTsq8puZWHjtX5D5TXfziSGIoQSPr1F3c6K2X+q8beb2AY1yYysaX9Ivu0K623bxBAm
oKMPWkTJTG7bSjznBoER/S9vlGX09xzxLmGcg/XlvDWXgGg//gX/KwOUtiggiNqOA4npJNvrJUvO
jJFKulfSZOgOHuIb9BL/38nauQcywM8iwyBszSjonV0epN4oj8ouis8MZClBHknM6X1hy9F8vVlC
e7cqd/cVVW5fz3DAk5+S4ZIYC5mg+GUpNJF/0IVOdN62zfKlnoG/DQeArsoyGzQvQAtRt0YLyZ1l
lnRrBJk0PpbA6UQ6itawNs/0Bm6c79Zss+Mu5hno7JMmVNAP4zLNa59SPgLwCbU+tfwe5IVOn01j
ae7WdYdKxu2Y6hRZcndrrm1d8U7vpB2OdAYTGk/8Bs4U+Ydtju2hsFQuI0R3kLtt2CRYNFTyBLN0
GzSizG0RekfNTKGl5zLbk5Ql3xidMFlrbG5DqNiRqJjGO7KqCHQHEq4OBlcCmXr4LvD1k2avXBY8
rgAr6+UgR3ze4YwefoQ6qgrBei+h4PNfU35/UNacaTfbplmSmdMzbIcQsdmpzQCOi4LEbp9YipH1
sAxD1QYn8XDs9HYGcmtwC3BB8+hK+7vMzladpRO3o0tMlpPkZwahLxrp22fk41c1C1mW5VgwUFMK
EQ+CL+6YPxPvRU/1JByV66KjkFXwc1JLqWjmcHcoiVkdFgVeA8P5zlD/jQMg3k1igcxgg0+q18tu
tm29TsLVzzxwwNmnfI0fc1eYdjavNlZpj3pPDlzg5h+o9oiGpG9ATzy2O/iaA+OanUWYxVeLhOjc
gf1nfnP4y26lwKsQ5Kh7IpbQMzHdhz1Xr3LbZPJNpU21hK4Zkgnd8mw2HV3VMH0dmAZglwSaAGlL
vutIZl6/G/1oEdL8nI6W3dfVPDx7tZ+Sg7TI1npa6ZKBbzUBqPMfn6nwxX5mVnuq1xvNBcdEMMiw
vcs5fYh1bAIMVNaRrXUVIJboOElX9l/cgHR1Ng55wZCDBd8aA5uCB0I8dlVRnnOhMuDrpaVU0w4F
W2snj1MpA4bw0P3E1LRZ9idNPa+wlzS+VjDnj0FhrIQPjltVJhzH23C2j1NV05YqZUwiQfFhA8Hn
3X9H3IuFqswYJP139MtROruTsGCbQptkJxnSEfrNS3CUatOSWW3bYtmfUaefofxNODVuanEti22y
3CTB+sAWaseEBKy34C3xxfCQQKJWV0cbCJETKTadfXllgqIh7jMNDIyJSGwLTVGszYWeUwOEa0Fl
1keF44kdUGusiQ1wXQ8dkSvjZzrsD0noXO8r1vc0zWn4N5935ndUcxxzW++BY3x4ZTdH5ruE5ovW
EZCDUNihiIjQVDmYvZZCpHwU9ue9JbcUxauu3H8T5Cmn2RHDZt/f2/jMllvvo6dJMN+J3+z4T02q
nZrIuF+TD7Qc138gxGR/FzM5EeH6mdLOJrTwXPbuE80XvLKMnx5TIxNkJZJ3kz5+VoQn80WWa3/L
9dWDej/TyMvZxath1CA1utvv1bxCdqEIMTtGHobKk0Den51xQm6o3UvBQfRX0qC24xg0IHqigwHs
ItLJ3uEA9fcTe0HE6NTe0qwgrKUu7gR0FHIeBWJmOur7nGjsTNyaA1i9bRDZ09BQYnG9gZdosWWN
6CwcIvSmGdi9XrkHWASWIhaIiKVfzbYWLWURporzA2u593Ji4arciZhBN+cbTu9Lg8PQzyFnudLD
DA5/Pv3Bmo/Iiiv8LxHLAoFKSflml3kdZw90XTQUlgrupG4+2R+ZQudU4tbhmsUrFTimzj/Y2GE3
kg/IFABKb04bZWRo6wDh8Q2m1+N0f8mPNaLFJWyOWYi9sFzwj1rNjd7Mlemiw4SjoMdiLTvcN5vK
FSKDMj6HKwYEwl2elecseJOzcjbbnD7J9bjnVplaH2f9G0bFl5Es7XA5xNHDlWe+q6CYIlibjK0U
lC4HX9IAJnYZAezGOAD0VnK3H6+rQ7kU+nPFauFeqfDttgaKjfrb888uqE1wdR6FxXmpP8q0oogh
wWWQEVgZ83n8mYHQ4iHssWp9XGe7LXm19MLbdqjdWzA3bd5y3lM3021sMMigZYLZGeBlG2pt6y++
KV7W6F2pZhPUeBRbaTHEjAmtrGB5aOaJutyeGAVhjxDI5VUMrUGY6HBE4CgbknhFpzwRtpaAHYoI
HrS4Dl+bNwUzF29poIMmfWc6cYReCNxUC6rvxid2SfTAhCg4kYzbi8S9IyUu6zezBryCtPL3MvoE
4kryOgHCe0zXtUdo96+/gikEhBqZ6M/rAurgu18SsDFVeZUESh/a1TEqL0YGnTLmyjWFkUQc5mYP
B9YsYeTPzzseUD7UjY4oP6m49YJJGfPBD4HaQNypcb/CS3PLcJb6K4jDTkRLYIsmCMoip52k8ogo
CodGxTYJe9B7ytHCogZ0tWZbqpu7pzEtuzmaMvJ6OvR4GH/7tk7esjsyrwxfrxShGZWcgX6esQT3
ug29oeZwd6mCe4/GS/XYxt7bcZKVxnSgDGTo5mQPF6IXP8jNJ42R3CeyyY0v0N+AZE376YfU58rk
rCf8Jz8fT5+Z+Phe+ycSjUN+IPB3mfHXo+KNWtZeqKaP4eGvvi+OKnttnrz7tOOJVfy78yXD1U3M
DL0nQRLlmk9l4J8TP3rtFalEgerb24oaRFRj5DwJvB1jkUqwlptsiuCsKUNk7YWAisehbkL7OyJ2
BtViTP7xaSjSQHzkrc/8pKjJfi2V/KVaxLYZ2UYf4zkn4BIdDRTzgP7PfCvKXenIK/+S2WAkbhmM
vB4O6TFogNGOvqA1NpE7mVpwkKczJYoufk9bJeBmZ8kgMxAWtK71ryKmfR8VIowLEOhaqKU1T46M
Ofuo9G4wRgYp6neMzjc4CQDdqG+iA0IPXfUQrUk0e1yHWcS0O/Drr723pFgEw45nyioD2FGjQaCI
2/G0tfsPamTuU6Zq0hL3Cwu8wQRoghsJaKmvvK5N2Dm93heeEKsCe9NTtA23Njm6pPxA4wZKtPJU
NMIXuUIiOUxRGkWW4qUuEFGfkcjwqYfCT+RBeFj/isWnHcC6tVYdE/BWFmYsdz1i+v5OPWgKwO7S
JlFKbNrXCXBLzIpyxPrIC/jqQ42YYkFxIn+2cftr0+JTFmNnAAcwUOBLO4k3Tni1y1PNvEAlSzAx
eTJtva4lqGnsIrJozvxRcesypzkNZrvgZ217tUwUMTgjFUDeyltCyG98JQpXKoCdf/RvNVt1kOeq
w03C0QTftUfvVp8JfhUyirzSEaeVr+NC4sCgv14RRJwZl5tn4bgN038j0KqarRR5XhnKmJO38ytG
bopvEFhHC1OQ1GaPhqKhuczunNdmazB5UeC1pzBRvdnmvvwn1wseqOQF7iQqz25ujzQZXcYYXgji
FSA28juETsFyn/x+AI9Q3JtY7paiv3WB4nDBI7wW0WIYChN0o++zgShpMz7tTZ3dwDHqyvpfyeYL
ORnI0WfbiomDYfr4744heO88R+4mI5w5iBhzMl+pzm6TxxLsI1zwLcC9ORBhuKq9ohpkrjSXju/N
bqotsI8EauH2NuXdYiLCfiE/qa56grzip8BOxwP6s1USNihS0pb3T8wd2lYz1yZ+qFlWwBkTpA1M
wi9rBi7LscSYeX3hWZ85FgOjb6lKATvE9CXTYH4ijPZ+VJar+NS1kHHT3CdYFaLuJtP5hEJ8reXy
U0fM2Bk5SJBxYPy6P9ofomxIZpAk66pDLgnyFwO/Qqg4b+Bhe68apguMgneacoS80vQa6A8cPzGk
eSmHEwxxaZfEnPGyydapqtYY7j2DLUeCSiQ9633bQa4SirHKJtPvGcYUAE9zuRrvBY9twtlmOkUy
Un8mZs67jHxdK+OD/OOAVCOS77KCprWY3CZOoSMs249jdyPbWg7pAQ2jUuFmwHEIbuOXPf8LERhe
dpNXT9Civd9ZCaOwvWmpYM38GPOPfh8jfIqkiFSq2ys631uKnl5YfQgzYEh9BHI5/4QA0ziafqoT
cyfJgHVg+sD8zpZSSOOUOWL7Ip7jxzWIapWNwxCYuQhMN9saj5QM3HbgzxK5wYn6kX/fkBWepRmW
PI6hROrzbLGSVkUby5Gsy0ncm6l7dL/z6tPKQRCJIahrUbB0DYpOKBufNxRw70frcMauI/YJB5j/
hviSwzEHvGejptuck3HgG0DaHBndkVQ1YCnUfE6P4uDTeU36vmFgV1q6uicRgYlP1m2k/IKb3JI/
/zSPl8iCXBiBw163d4mcmShBUie9nmm4VnLQXwM6xyh7hyz6+BEbT6ja3W4WJ8cBNACQvZprR/AX
6o60DIkTc5bG/hF6bRN+GiiWBN4vtcUVX+9KPlvqMDV353cOOeK7xlMNQVf2r7dDXE8NSJ8UZ5r0
3UhDh7AU5CcH0xXV+FZNS7SXPK2F7YQfco6sR0/Qr1d6vIiN+HPEkELZyqEQSihfoBfWzgH/WvzJ
36A6jESbEnTw/wVF46T4IiAQienmCEARb+rgXW7jVlOAANvrOjyV/Vx03O1SeNFRPebGhvHW3Ul2
3+bys8K4zY0QKcr34q7iLDnvaxzpmkAUUAydLwozb7EZL2t5IjYQFLSTzD5/Y587rOQXVsBXQZuh
8FtgeftQTKTHHeefUx2UVXMB7aT8N09ZVRpwZL/th0MPLxSBWt6kzn3iFl+rLZSmYmro1+t+OLsg
D3PneOheMBwYycqLhKlcNv2Qxeosu+X79JyLHIdpIoU2J5cFjOCOcnIf1R7KtMseWUIqmwo3erW5
DCMqHmtUFCF7v3YIWoy0LieSW3wCm0TO91IyERnFsdkyUiM9VEQXcpE1tZ5wgaMpxe08eIZ64H7w
QdBM+hZ1WLkEqdhPc2QQoEhC99oassZweBg9sV0n91pvbaUnRFJS/fuayfBceijfYZpZgERgApN8
helfHWFQ0qZZ+gDOSoyXWhEqkSegONGwNDw5sJHEZbwD3rSIIvNZTcKSIKny9l3iAootgF23JcfG
m2QXwMBSsx1bX3yBFK1WGn1i0QEbBYwNZu9fXsFJeLl7L7HugnoTuDNqYRoPw6YdmtViZqkB4tDp
W/n69p7ybaQA/Jh/4qZQjju8zZwy7K3V4flDcTl8THclXH3HILvxv7bRB7qq5Uja8y2SUPila12x
9Sa4LedsowURyh7rI9HLfT4kjo0+ASkeaGz4OwZuTYC+G7lpJddhSveoW9WBgHZnN2ETSx3hLkCx
GLVNiTw4IGeB614353ZqMhn7jdolyjo4BwfJKSh73eYcSrxKNN7cpI0NHFkCgYehOyVLb5Bts5rc
OfpwsZPbEVeMtD6iQpTTCcibhlP5Z3Ozxv3QVr4zrUbiQvwsoNzT1U7MwhDzyKsLejBYoC1O7RDv
Gq4sA781uw/OLFeLCsKB3FmPLnuigrbr7Gc4qCB+jSqeDnsioQirK7/Tk74Jf0wXBs23VEPeK0Tu
rbgzw4OxzLONLLdNiEIX8PBG5Fzh61A4yV5XtG80emByqgmJE/UyERJ4YucqsOiRoPVM+2NhIVuI
iBjV86HdYEKDTwERitEK5no/+zJ35CpY9NQ0cTzkyPOuQg1pB6aj6+gZFu5mEfUFMhhFBvb75Z3C
yLS40swKZ/PJgIs7IqWPCc64FpAaPGgahc9nGRLu/+I6a+ATG831SYZJNRTllO1Wej+mzQvlvsTG
hE6LzoSKPe3HfTg5gJw2yOoA+gqBCp7jUz+I6RcyhHLMNGzfXJSvU8NUCJy23aXwwyVIn9qKJlWL
mXO1Eq2uFeyMc6ByVEvYsgDh0lLxONf5i0+r4Kr6E0VjkpbA5ai74IaqZefuN3GSZCbBR3RIipCv
tB+zp6Rwo6fdpYoE4YIW1zC+LnYlYqTtQJTBusDw1uRFKyp/uxeqhWGLSARaHWG73z+CS61sRYTd
tZTH3aI3ezdkfP3nznb5qm0QjBn2wwKJhsKRsSYPXNcPwI3jx4luQdPj0RP0oWD12rbfVM5B75iu
3pq4K+5A9g1YtcDvO/ar4gmgwo1CGNwfg6pElFefpz1oCSimiyHefJyzJ+3wJ17hOBI6k+SmBe8X
zFddEIpQBbxAdfsG1HCO9+WjJhZk52oI/6QHPwwFkAtR3Ja7XnLtfca54Cq8O3QiWCsYFg2du4AQ
v3kY3vbrZODROTsoAPVIhbOISc5ak3w11yqxcy1fPb899UTgrLALWHtAURzSKMJ62mJpSYYxzrS4
I0+4M2ycEopbjmGK9nVJX9/vD2AOY57yc4NnJxZAnRFtdv7hJjpx2TjruTe0vVibbjCc5CiAnXDl
1LTGni7Vc8GjzvlXmuKpMw4ASDoRel32UFJZ/aCu1lPO78iKRRWifTE4aZ3xCoaycwIgJ8kOU+/0
VzOQpUooF3AWIJgMCwvoHHRXYM61HTz0KJefFgghqJi7X9zPHF8Jk8/G+5NKv/lDt6nkx6EnRWMS
oA1guw9cK5Fbz1XtAx4KOMQAMLFRE1nI23VIv4iVmjR1P/1Y8Bx34eLTmmzW0PuFZi7JqRXe+oC7
K/OLttiB+OjvY6VWJknxJW6iKdo+zpAQBxPNexwqrbyu923azeVGs+FpGFvKpZN24ccOdagdaLuc
yryelgNAS7nAQ/zFo5vvZIP5sDdpRTSRvDSMcgoSlKbwEUf/ktE/zVbidRDvByXkMajHEzt/U1Bd
bAjS4CYBIVSSgGYYRzOMfG3zLra5Xirro40zZsClrvA3ROG8UKGqGUGxOZj0VNSKmDmxtSHGJpO+
w+JhQEvLDtaVxnhBb96HAbcqSpySoSc3tPVXTNU4IlDt1LXL2Hc+MuS+IAzgQW/102zHYuLPsAIs
giFzp8cj31T6O6vQ+aGESNZqNdexi7dFMQhQWSAb7VSAcC2JQrwZ9xh+PaCihbhvD6JGyxH+0IAs
63u8ma+rQl2zKNpW6kEnpG1O9pgP2FtD3dxQ4NeeiLvv/c0qfMoEqvOR+rdYream3vRMKfHFZojg
MZ4M2z+3lyp5be9a/nUfKFKJRJpGpNHHueNISvO8TlvaaKzH0xRslHsWvnPBr3hYRWBPT7k3SgsG
nZYYI4jyFESVpVM6vbK7Q/iXg0N9/pHS2nx2axb0lqqmth/2xb4S7fKjQlk9V9IamcYjrkUMMhwt
lASuQ4qZUYGHCedZb4hOlulIOr2h7U89FrUB+KmjRC8OH0k87N+EEmbNvHLwR7u7AAXcVt4FNFIZ
UjbUalkzN1veLc/+hkWlKJ1YJOj2DU1eoX1mH6MvObsKP/1rXhagpmlDukYcQcxHyffO0UxKjins
9/Pn/LTDYiE9aVQDaTh7wCRttIqb/HOn5tUgu/bc/xe9xZ17Nv0slLI50l4oDdXynhFhlvyAtcvp
i/CYdPLjZNTCUTgADum388R9n1o6IL0dywktFKpfLreXuIPcdBIOhavUFkaDTQ7atn2Kd7x5NqJk
Nj0G7pD5T11+2lDTZQbR598VnO+Rrktx7i9rfEIoosnz3oq4+n/LmJVZ4DN5K9PIPGzoStUbMhyT
F7eELdfnEcnmIh46mIc9+N6gZsVjKD/faEvgRA50vODjaMbCC9L/SIJwLXF1qpQXhvBjDMRrzlaR
TVPc7FRrIPeNdCus1exAGYnUqiOm+FbRnFDR+FiUBh8GivRjEUUwEuv3R3wL5CyS/CNecsES8g1J
dSNiZPqqCJg2AN0CGy4QQkc64RarxpZj2JMmJvZSRnF8fndhiTVZMGymuukyoa3yGQ3rJyqEmjms
7NyiQjy+aasc8zVD+Upc3eLKT3E5+h3R2mzIi8JthExZbFUt+0tCzeew2zzeE8oqnAgYNyhoOkRr
V03lOntTJZGm7pxEDE5Co0FoLuTluxFgSUncLzQK1lNKrlWHnrIWDUnl8GOWiOg9GfHiZ25a8PFl
9nbBkRnfvaQJywT08QyRSLM23CNqsCpKQhiX/NMP/+HJN90TQCNOf9TfcGl1g/F+n5n+p2UELkXQ
qhE78NjtHPIFuH0gwLeofgGYADgUYF9YAQ8dq/g/RwY+qAIbmTvUNKeNC1g6jBCT34nvNIrj0fTc
LSOn4tMpW3dakaXmh2xHjJn60ZMaX64rPgkZHieqBvq/wH+0f/Sim0V1rYNVlOZl9fPmAfGAH5FV
pPMPoJDNqjQWMbIpUJc06Ffc6ZNFCmoCJjuFP0E9RlEdcfmdJNm1VJ9Bg0j58gD96WsryGeDR1I+
jLjNJGeVwqH1bspV3wOeQzZiVBQqzXChs47C7bqfTKi0npoDHjUVI4ekgwi5z2R34pD2UWUN4ycz
fwubVl4kpQkYyVhZg9P/YrggKWtTUs69/FJw01Tad58NyOuOJ6h6cgsi0DCqdDeMKJ8LT2Hhz29B
xOc9RhdidAqlR/omSA+ORawgnaw73eJE6aL1fphTqTxuIjCJ3fQ7hIzTu18s/cb0KIx17X8YAdRP
ats+8Ye/U2JvZp6gaGA7Ju4H0Y9ELe9XXuYeq5bNyX6unZZUhLGTH+bryvaSsKrDm5VFfzTFbPX/
e/EBZdKSXXgHyjfbdxAWMOUfAOnxGrL+MBJvSG7uSZyVHmBJvrT+lNdXaqUjg0XhlH0xK9GUIec4
QJaeGo8vXlir39j6hF0muVfo6JEZDa9YHqZeCe0IorriwqzIt79oLgp5y2wFSMkA9agXoXcrg9oV
rlJReHqlXHllZZ+cnkEjiIN54o880E9B+md5rSfUYQe7aotoNcLzAX8wMmmk5ySQ6g8nysLeRFEe
9A+6kJM15U0TG6RAGP2VN2Qim+K0s3m6qt70be0n9JUwPI4zgaNk+oLssEJF4eqn7XESjh4jrzVs
zw/Ru4X9qxjDltUtQuCU9BDtrD/RaPEDawYAno0pC/Ff1vdjdFrTDpO6cbUBmdStA+Kk3OKl9Oiq
dRTfzUaeyNBfQpPfss7DNuhueu0SZdovEnv2JpFrHO+fjKgUVVMs4IaRlJDaGxtNuq0jRtTMtZz8
LXDTGV6qh5hHE5Iqsjsg/S5fepFHOCOuWVHfX4TXfHkFcVPfbBttR5Z75WlxxpTr6zKaVCw2o6Qb
d7oe99PJS4z6/Odhl2xkOCt3Lgb+hATG50Av93UECy8UM5fI+i91nzH6WhLTgoys2l/c9qbrWl+U
8MeWJ2z7v19qZPsmCrVCQedDEcC20mbr4oLBixq29Gblnr+bBA8Joi67q3lFAudu3hQgf/EKRifd
/sjig1Nrgi7VMJnLrsPgBPKyKyGqDo2qI+QT7cYy8gnuqzasy7uIT/2tvnupTjvRYBEX4b18ooU3
Q1E1pq3V0QsfwPQkmOpVIKfGqkgS/VMOqJoLCRxbDrldIdC0J582Zrk7UUZIv4B2kyv5XaLdoy+a
7ow1WpBBMS9TAML0dkiNZwGE0J1ajiTeBOHGRmVlhvRASsqRRZfp7FOGbFvGzQ0A3TDLwapSUDyF
6GGwPHSPzZvcqNwbSNiRZJROfABJcefJyRUCc0f/ZfRpBaNJgkUzTU7HfaHn8pRrqmLA/lBTOEqk
G+obtS7tT5UrhDjaxmOd4dzWGIyWXax5nJ7t8bfYUY6jowmYGPZMCrhejeIWo5JVxIzVtRzn3ShU
Gwa13DFJGNml/Fp1hVJHa0sUy1EEgamXPadjPImS3NwqEuKt6dkzB9g8bD1i86XLVT4o5+/QXOmS
dW/agNZTuN30IM+iaALxmsSBPV6YApDQktK79jaCp5Jb/PTrRT7n8i/t/dHDoTt6AdSJ1koiN/4b
NnOw8Z+td+P4yFynaYtAu1TERQoppPKadPyX5eKhVvokkcGplGAWYj5YEsBhptQgrULFgE9fMjV9
buazZN002n4457JGpU+HZC6uE9yFWpTfk9yRMg7PijlDyP3kTf8jmpX09OkBNwItudfJjscGRimL
9YnPQPyDlVnbfjmI/3Jgx4Vmrv0CIJDRV6SmTQ9UuehQKnWEzgvlBzBZvOIcdvhDuLQaNgMs4CYM
hBrKHbywZDNlw6piqBQt7b/6S4FOxPg2AmsxLe3SpcPA8IcXYccY4uS1Y6fP6ExcqFBTfkMD9wyX
+yZSF/nBNUDqimclkVIMqN392CfnGhHn4Z4KW9PhjoHO8tv+hFoWHG2MoPbTw7fPnd9qqrtEfHdi
VfN4ojUqIbxRynr8cq09ndE4aulDGIgUf96MQIKztm+lbeAuMzjnpRuq7xXs6CfXxpclnsZI7vgA
m2ezXWdEx6ukvJ9jVGe+FTxJ0OxCNsGQ5kvLeAFgrsBfbPZ+BYl/uBIt3haaOaKXzEcSvfGT1icU
ANjlX2rYtQ0meqtOnMjdeF2aMc3stlyTdyz2Ru0nlW8t9I2mzZq+JYOt+REU/p4KPKg2W7dXVeOy
jjZkwgwIbuRqVggD52n6IKJoBRqVpAXrQoSKzYFJtOG+tBXq+N1LlbEqkr3CmiO5DWUBUCT8uSLQ
vC5c8BGzC2YHq8ZofW+J3H76UPuPVcnCwZ6hIQfrH3s+vYUXrmR2opsEon7ZeWgz9yJmDYGxBlgv
I94y2pPfSrVYOuCreMywKIVjljmvWWD6Qbylx8dOXse/KmQwuXbCekhfHSPyQfi2NFwD8cNbY882
7Nj4W9yyQ8Vsfvvq4v573tdVx65Jl7GzfftLn06TXXpAVQP7jc3hWRbBQqYCHmFkxd2wcMBGVdL+
OVmMI3jO8SGg/00lgUG9NLAeDr2kP0dEWcCPQknIFlNtJyh1iy03mAXw6JDtIbXZL5ytF2tqJJl+
by9MbRi0z2fXzTizQSHRmVkydFWKcIEpPU3I9n3a59tCYd110TyZLmgrBMkHRgwMWqZehnMUH8oT
te5GPuT5PWv/BxNmB3P1sDBH5aan5BypILgkx3jBtCcaEWA0d4pQzftBcnKuBiAOv0GfEbUBygEv
oMT0rXex/MKDOzupynGdjfb27n2WcSRzi9kg/ZRROLN8caPZMD/XoDO3Gcwsw1Uok2QJLMiXUPXO
bloFAxltNpn09+P8mb1Vb2awNaxrAwdJ8RnOTiOrOHFayuIIKkkI6jrvOrft0j5RNNVTjq5gCgEu
3IIVjvdh6i0h9ysyjnUoVnSjDAT491i3pKVpYpYSojj0xsSrXA17NNRq6dB3zAJpmMhtNqpcaqru
WycgwFS3TpHJNz3w1+28wW1atBnp919AFflb5GrZYWaAQ5WpFXesR1cEbVZ0p2EehSY0TskZQl2Y
aSmkWxeazgWRrP5mYVHN6djCDGQjQjcfyc1qTKjB8KYLORmYXs4oAtTyqwsNQ0sam+ALLUZHhGwX
rzWs5xBFflb/UjCdLsIbCITC4izrOkZC6bzh7nGy+ZN3lmzkVQntR6vC1WZheuyxp33mGYCma67v
XX200Rgj9nsCV9ox6o4oHCt0+4JcvFRJ5+4O2KoGrDIPtpfB5AnQAhDS+PM3mXpPARfeH41kt5zA
msBlJuyt7LsLVT1c/CDxaYGowQw6Sad3m+zHwOXU0QJosjh5VGbPcua0OM6gq2NlXtXNAt4w9Pyw
ALP2z4oRMqmupj+mr9OtnC4jiNB0Iq2fTUd1PkgxMT/3uvTP+3I/P6f49icQCFaHvYnBp4QGUWBy
t+QmjWMg1ayVoiorWz6ReX9bLDAlwA2EfMoSIkuucqMadlnljRJS2bpQMKgz9mwrkeC5hoM9GAbl
Pp6YQsuzUOeXaVXovduyCcjfq344udbtdSwq/cjMDmJOh8YMy66OQfV0+Y+8JYO/KDX4JnDRDVzF
HpDpXtwp9LP8PrjWSeb8IEX6ZYDpGw0fssd5j61YMoPEH9zEcVcDugBDdU5cw18pS0dCbyRDyUow
C4GOr0FW/Nh5va9tYkZtBU20WkInmbkLSHi3Hwz0YbQZP91dTgLWKXXhDliFRZl54f4BV8qNGT59
mTlRkbmJyEsLR2MeCjBcYL6suDaxuEHe7BmgxcdygE8umOanxfXscZucPgJ4tpDeReClxHhsrzU9
BuoiLQYUjT6JMSzfI7Uvcwfkz/nR+AXa7LDGCOoJBT/4YtAZrwIGdl37df38B4NUpiSGpBowxV4P
JL/yrw+g9MqZSNiCLzV7rDN3q98OFC+POpJj9fiHB3tZmC+Uzg7PmabQS9f2clrrMgCK/EGvZGLX
Ilv0FbQ+HvFp1uKQgNUKjfPXVJJ76aIbAsm/4lmhnLs04gbbKMbQy2D0fFD2AKT8fdqkafmHjrg2
cdU3mP8yzbVW8qH3Xj05jakBUb4fq9H+CkVGdLdTSnv+MfeugOa8uCBdwJCQhIEdi3coPMKZO14D
BbpJLBlU1nqqrhOTdj3/IxX5MbES2UIX6F0I2UtBqMPR/zTsVfTCPsfTauDJ7igeDUoSQbPLCrVp
2LIfL/QtVDkAFL2o70myYVzCM1kQma8vLksbW+u1L4zpNp0Nc+Kj5q9v6hFUrPdHRUx2jd7XlP0o
H11xZoxMnolhB9rFSiibzrruA5TCEngBRIsRsGDef4u6OnaZzLHLCqttYXRBN3yj4XQl7bAl2te9
k7iFe5xmotfDVlxKJtFqjqxMg0CSOHBakXQ6lmOMyHsEbUelCwtQNPUr0dwUHJ+yox+NXaFqI5MW
JZGMZcZ64tfH4FgadzjOKCyCfUMPL449NsZSk+sePxRF2NY7LeaGOLnEOo+qQhqRdVR4TZtIKLuC
C93HpuLd+vhCIUjjJX+4aVAKW6z9nmwBDydpsS9n/AaVNsh7dRiYyibMBNmP4B5RC/pxzCjqk0pd
ascWMk+CYCGvs2dhihjOSvZXweAYuJdp/X1Voq1tXavYBPMHgzdSl+MH1fNRAQteRlUvzw+WZ4sM
qxq6A+1sYdqr5tsrIOqYNKJU1mKTQFssfc959rT4pkBsp9s+jeZy7xZq9uHs5j5OGcy1q6AqKVG/
31DkYD9y7dTjJG1cpkX2VPK8d+mYjYb8kqbvpL5oxYhvU/0IWTjGjV1RIX2pFNTIAcgE15ZvbL1H
Cl8i7sUbQdxNe3IYh9XYlBn1LpIPA72NUDRwUe8b7Lsb35xb899EfwtDz5Q+fscT9pkBVa11CR0e
adP1NsuNTGXYMy/y/IBfva+Wi6GXg/OX9st97aE07UxINtYSXnXHwt6ZTyFlRbZx/WK6ALdRUrnY
yI2K730FoL66WOmmMs/eb/h//tWNomkJ4wfnaaSjTKZBC6ZLuDA3ujLQX8ZjXVLjHLw1EUfEd35p
x81bCrv/R27EemW0L79+4HRajeexvPCrIqRMocgFL9UaU6J2+pv35g5k3gmJ8v/25w/pG/2ttDiG
I7qfvYtyL/D796oL3jL0k8iWYPlYecc3AboQ6rInsdImukWw3ST7t7P9QkCssoWIrzQlTetjTFPd
K4KpxwnZO2B5+1XdC0oUCYNDQCwL+eJKOwEl2VCXykY86jeDymaOr0mRnIn7/RYnG5HE0IyXocqL
r6HyFXBOznp+ILHtCRCDPm+WZhKqqbheZqVCIho4amVZpR3s0w9qqMLmu8xk9f33hrBWXPtV0+ng
iiqMdvIM88fHqohItRNSCkvcHAws1sapx3rB5fDxbE+pASJdmq4DpZ/cGj7PhlAH6DDLFuC2NLH2
LET6zf3UOVftgSJ5PFBkpg0L35PdcHoRQVCduJ8kKyI5CQK/UZEtd2l0WbuMEQoH/59HfDZaYqZG
1ryaaITK7HD4cW1RzLFAjbjysytRx86xAnpoauF3sRyzfoDE6VZ4aFSmWkKP0QXpKegGDDOTr08H
lbuUlfhn9QSsVTBwCRcu5rdiPxf3yE/YYFh1LYeMP8sb4NBcHMOS5TgfSLDTJO7nfuiS3F59rRSn
23vTa0WySxiWfcT6GLZhQGGD0JxQsTRFpSA1vmwPg1idkrhK1xBQ7QflRIx7eMxDBqOJPwO4qx8U
kzJeTBvYMqZoMX7ow3081KiILnT7Rq3qqLgG+x6R5C00ThxNN3nKoXr36Cm3b8EirxHpnFXAEAM6
H5pjcgz4SRmrtjLvIqTL5+LVt+crYApiQKyiSOk3RhUYNHMtXtCY+VgX1Fw14s34WA8CPIEkH96a
jzJp8UhqbkW3BQ+vUFBRzdA8z3HoWaIESZQ3M/OcpitJ6xe/+e+5xQrYcw1svpOjiINwXbQZZywd
3QQ4OCNga5QSCcz/Ni/XqqWN/JlYkqvjAnrL2XGuZ93UK2r1gyvqBeIxifnNlZ0Lx90aPhk9Qf/I
aWtJbEpO4sYbZVbetzb39SJ1mLSdGNvNqU5TmaOVLP92shyFIcrf51af7Pdo4xBXaBDHkI/wU2yk
64eco3BY1Wiz2fDwlSjo78Jf8Cmy5PZBUEWQT4roiXg98s6u9vlt/9/1UQIT5JeUXKdVwDGUs/4T
c+SpA6zH9yFaroKYwuDYS9KXFc0qLftvik9SJHXSPVvOzeIdUXdcnNUEPxnpiBkOnJxJXe5E97NZ
O8yhNtt9rDC6TPsv5RvUeuSW5iBRDNWtcHd4Bt0qm/lpXJbQK4pG/2YziC6D8ZSgp/qsWtrppb67
fAJt7BBSdeOORAfyGPVRQve4Ou90yTN32da+GJN7juj/ozms/uK2xOB3Rsc1NSqwGeH4M2/Mf+Se
nsKBozRk7hygeFEuY/l5XtCvRn/DxLJqTlrHuAEdCNXe4x0YdV/n3uzQmHEDH4gUCmjNgtZzWxvL
e02faoXiZ2Z5Qdw10apfaO92ZrTkjwQe0Fn25E6R1GN2TD4ulojW08FcLigWGzyWmZW9uZc2dj0I
3plMvRBA/tTGE7RaTloa00rK/UdbUUovZWkrowywbFFtUcXUGboeszXhN+5ULhI3ZuVLzQK4HYQz
AAPzxUvAoQMAU5baTdJVAJMJVRUdXrnE7QiRIIZFnC2UVGhFYCRdb8cQOLSnZAQvPLdPKc8QSgz2
GkgbLAwMQnWhP4T1G3cLaMTLsKXTU+tO2QZoM3gSE5f5Cf/VDATMM6BTlooqKOOvvcvGYJEU3mLb
9UupihAsv+UaejcetSVQiJi/l0ch+48bGBHEmjHGKrULSdzqRwOqrb1ySEwhZbGEyE01BbfZ4q7Q
3kTwje1zuOFCDRb0hqF/NYFin4criXkHXRr1vKPu5kvmfvPzgScF26wgDTDi3OCZWREHfszUnfqa
Dctn/P2lLL5ACQhzb2kcA8nruPABPsyiYgh9iq8d8lQBCYhDZdrDcmYPwbhUldE1/bHBTOzzV8zf
cXwzYvAB9b6IVCDOhyIkh11ZUXQ2tMIbx8g1kyGEkMXC2/PtwGWdx9PbwTTxUl3neZWyn2fBA2wp
MMGU2lkyF2+EIw7FFrOu1sPEziPk00IwhARwTbYdwASjvuFow43pMpqRNer1FP4Dk0mE1LWT5DjE
DodtZYty0z9Nr/C+Lul+LQfyNWypjuo1Hs+oncIBjSORKG4hsKK/0WGKoOqGDal61bLBj9prpLBJ
5P4lxuJmgIX7ZlmR0n8tpI9EdFg5bdnJRIR40rB3kpFeqQHCkZ7TWWHV2tOG903HZLa+6b2UfhZl
DrZ3zyT+Oi+UOkU8+3mkFuctNSIvUmtrKDZzDbS1NFLLQE40dh8GPr+payFywOfStjtdSZrUK5Cg
RGUODbnYD1MWFXtXDzxG8FpXPrgEjBkw8PpXOr+otBNPi4TKqAcm+cDb4Wql+hcxplikl8HxjPdF
P0ZxV54La+n/pA4CEU8AIJbTZOT7B/+h6Z85DHME8x0kXtAs7GCUZF4d+weY+yKh4PLg2eYXX64Q
+YOeHSoFNlJFCIu+zFgJdRxgdxrjQwtVXTP+wgExHhbUWLah/jIRk+2mbxz6+aD9SO5XTPffz8ci
2T2Ao3Ecnho2g5278X2++yysgV75rpMyoWQWDbI+Tq37rtG+0/v5TJXw9XkhxWDM3QO1piUwHi7i
2HBq3gqEXCMaydKzUFhI2gk7sPkVuV52sV4LJAN62L5L1ef68Jo9WN3m467XTQG7BfWfkpk8aUKC
umfD3GclJ/IC7c5yfCDjoMOmh68tyKk5EUizRZTN1FaKWjVt6w+t2TZxj4JIyBsDWmCWE5mUEXjS
lEoa32hS5fZrqUNb0ZmyaX0LJzsJ8QZ/IZeKI/FG/ndqo0YOAg/nkh5dRdDrea3Y/ukbx7Ufa+H/
LOEqdblqGWTmPTz3Qjj2xZfVzguHYpMPujbHQ6/RUmOa3Mcsf8Em5vBvdYugj4Ua3rOiNkBhUZ0t
P2zMQEqzrArJ5iif2AJTz7RPCULGRa70Y3JgdMIwEy3mbXw13kLzy9JCv6zDx/JpzgTeG9QY3yVL
mk0e6LX+99nFunIuoPf0nkt6VEXvdhKxXAMEE0WVHsm+FTM6lHQmtnJLy7nZ1bVe4LvgJIb98w4j
f327Q0xoeyb0SWCimMkxur7w12zC0XAslQQoCZbs4kcAQn91qsM9B7D1PrEDUhQIG5zApgoVfMUQ
9VTcMpjmSaEIzUvgWYy8u3igskG3YXHlwJsDG37b9xWQvNROo0/+1tWv3PVkUbhB0xLkAXJeoLdQ
7Jotd1zFlH5MlK4OYWzV60OyBVttUw295pX+xwsXy6b0JuOq2tdY45toeOgK/4Eet89sezkbsMu/
hCZ5Uz7aVN2aadHngHmu6itWlEQEqrpqCgyAjtB94iV18JOsFLl8jYYAzqPifuLTR+ojF26wfUn6
KxKFfNIKnh527W3geq5tOal31pZsaTkIJgKBCmhcRFT379diIYo+6XFOlM+d0e6DHy5svZsgL+Zj
Q/UycHESBGMRspq2fCkZM29TbJtR0Zqg5HPh7BFH2v/2iQjos2z1M7Rw/L8KnGGcovmE37OMfnDb
qn+Iuwkp+sChBisjUJvJSYK32+2OPyBjfAhSWyKPDj+bnYyq21Yi/Ao2hkNwhGMPervpOIMkP5o+
WHn5yBWxgEqPSXIaPgyUtI35sUPqfGm4Dl3EsBMD0OlWEJsS6p8gWTJfen4mbq2ZMiNJYw8wTsqv
e8saQcqYbql4qfoJZ2g2ZgBtOl9aL7aL4WXmiLKuoKL7JZ1tuaD7YXn7pX/61Dxk6AzQmMmnyU/c
MSjabFuHYFo1J31MTKJrboPHJ0vRyS6ncZuWYBuqD6ixI+nl3UPIjr87FR4dwY559ud4KId3WF9v
gGQSQ/0fPDAS/oiGC2zSK1ym1MQTslclD8S4A2xMakhs7fK1PV9ZnRSX8KCr92TCJ+Q1FD7QTwda
0+sNfOUK9UXiiDd9BK3jKOnw6h3Ak2oauUjIfqaS/VfDHprumMK6hS/K1X3BcArPoKEC2sAzW4zS
6qsLTu55Q7jraqkKYANr3ocmAQLEwyYySq1wionpQo8fxOZAki37EPNK7kQu4puDqupby7MokrQh
HedvAfAr5mHkTld2scspZNn1bjDroTnuYwMgVj52NyQRX35rm1HCpPRfBaEdhU+J4oZpPGEMC/Ez
32dxsKx9/iJcs/VdUELHK01fHBbo/cMdWrMa/u7y+CfuKqMOiVZqXrWkyqAY5WqqfNJl0DJ8Akil
BLpszGCsyODjZN4pAX1O2+THNu4IQ5p7i8LXzlKExkXwRk4Q/bpkVg4zjwiRGsdg5qlY4gmFNBO1
tIEO0rIbeSXfPRdErcn1ZWmxJ6bt31uSb/gMny+gothEt3FXsFnPqjZAFpVQs9IWUpa0Zh1RzvWg
qpq0AwVq6sQAb2tEkhj8CUIa8mf5vVAnLU06Y5zjjtF5au+iif3s5d0IaojtAZfzo1vZw/fSvqaj
vjVsEsx26/oGHnKvZO9wzCRNX3Gj/P53UE5TVaQrEXsWcvdaAzbfilFwyXhTKiOSAm0RKNsh4dlO
rBMv3eX9LmMeDDGUAA5cO6tLzuFBDBs11QRXeMShLnJYSiog5jRRHMcX1SDHPAEdeLud6Z5rAuR2
SsNhRrb3yXxW8NV/08zbcnHVlxAPDn/VfHV5/shqzcy1P0On1e610LvKgJvGCmc+qcY7kjeMraS9
DnPGozOQ5VhOhAWwz5hR/i+hreK8BEVmOU+8BJa9+V7OgFinRuYhp7W6/9HsXXUmU/WNajdXskCf
ibZwCiymDtXSCNH80d1muzVpAG7yn4XhM16nSJQURFktVtVIjzzU1vmxOeQOT9C/CnpkPrw+uO7F
fHKLd+Qr5Ck6ISURk4O226hZoUbpapyn8aDYKDjxUrz7xyXf8NZJbFyEV3JIiA4OEfOMmkz4oiV2
+UTr0VHBCUe+dkOdnscZmcTgIsyxGbl2K6ep2c8K85gEvcnIBvi29pRxJghd/Tx6ZR0RRD8ZNxMB
ROyjMy7ILwdyqrFCP7Y9S+kYw1a6ehgrgx3wJxDukb1BdCOM2r2OfJ/Xv7M8XXRaHMkr3G9rRypY
TnZwr5XOWayOnrC4iyHAHMt7aY8YdkkmEWPzYXT9B4/2HEZLlLbCchMtENa6NzUChSBiaeaPnEBB
2uqpxRJk//dgW81zBKk6fKgH8PobZh92O4f8WLYz29EApZlzzOjY3qRmkzIOcGjrcVD966lYKJiD
foZEWFUhyIaQLDX/V1KB8pC8IR3laVTGV9LegllUFoE2ybmJPMqN3qY7/igtxnzmUlZb11i4fS9+
PsjV+AEvDLu53zqhEfYsyGrsVMlFuP6gZ6e0tiMyWnlxaaiTR1e2mVxX1i1da1GUOoiPg+K3ZnvS
OX4L0BfOl1b57ijMobJCbJsSPgdQ4EURsbDYxdkvWTSENFwYbxEJl0EyUVSTnBTxwl4Sjl7EkI50
3LgKnhIewtCN5YnilfgtipLRhy/5SDGoAjlbzgIyRJz401pMLH5tkZHNUygirdhjstbuOKUyzz2w
gKee0daGh/8dvzYhd2r/ftcTHAOgbtyszhiQGoaxe0QjA6G+plaJrf85v2e6RTSwYCmaaEIeCsMj
XlIL9rQvI98uSrDnIyxqJ4/Age6reJZoogxeFez/+K7uWqva3veNMigqVl8x3TzDXc206glV22TR
zuO/+/H+9mMMtaZlhgvl5c6QKFgsV5Hjy++8LofPuvHuWUS1O65c3xZhVba9+eD6vKkfeUGfch4a
FIg4jePVuimIFG20R3V9ggemwc79rr8A1MsRmmQZ7xrW1hvKMYGwPsyAq4sF8TpTRNT2HgRrhNRh
ze8aaOQnf/Ebgldr75P1+XeVTcdX6de9mfzJuymt86QURedhQknwppvT7KfHpu9gA8VNbIFpxIm9
2XJdjqMQA1omktdeNwSxOrguzJJuU64PpQTZgqyhvvJaTJqY95xPkqx2lZX0dmIfdAyrnJM9Me6W
vpHFkMn4tf3cGxFrb4DggZKGaSuRPKalmKnuSZU3dCdoQ8PZq97vGOXJe9aiWqOZycEoErTtdpl+
LB5XlmoJA3OTWqgAqUawMBpJZ9JMLpV1Tmn/qGuL7PPGvrlpxm/4cw6gCs0yjluJZGKm+ZAbBdh4
WziJYSna/16GE6uvmdYVK5J0SIs5JAbH/H86RG1nm+dAwyVoVV04scgQd1FIFj3xkfI7oAzH485C
4h5e9Y+G8A+swIai/uHWd2BwCvz4p+Mc6fqBTqogHu6k+ADpDp82aQPc9vsQUrxlyuY5Xz+8ylL4
DsmDAIJ7MC6zXWcETRgEQPve9jBIAnGyrGelAyI26eacsV7oFR/QMs5IwOFkR8L4ZMLbf1cm+RbN
dxmsH7iajEKmoeTSbd3GRkncDO1mScZQB43H+OMzGIwizfe3qdqqNNXpGZw5Dh808DjpoRVJTKZQ
szipPguuf5c70Aln18AcBN/mry2YIwWT0olrmRiRfjyq9O0491x/Tm8h7CL00FMEolkXELz3xV/R
dUQYz/BEqOrLhAKyPDAjnzrTY383/nGAm3zNA8yzE/VddGnjiZvzpLo7yzdEgopDmthFNCwLW9b0
1DCDXhtBORyh916VGnbFuK8peOp7sq9gcFC2h8Z3zQUFVpbvNhSqowHTAWTjrTLy/Kw9oWa8kj4h
bitGG0jI85AUBGgcyUkcXF1vUymHaGltZJPNOqoUfYlQJiO4W/RNvuvSdSc/1wflVYTe4SMZ6v7s
iRZ6ymscqC/Px7mgui+syM5e1TlQ7uYjEbqQa6P/QQBVCElRt5aItuOuTSB66HwAj2xKTQ7punRU
iMQBwQ9sTNIcJVnWi1Zy7g16GPUiM+44obvQS4aCgkYVCqbBnYxctkEke2Iir1CNi3cA+KPKXju/
Yb3PbId8SCiqoQEEpy5/3rWI+npk9rq9id8b6VUilBPI/rydMjEljeNTL6kOJ70mXJYHh+kgiiF8
0W1r0gOC0lWkXl1EqcwOgWQrQ8mMqNAbZlzRF7i88Qi67KlrF3Rh8Rzb4NJOi0it2I8S6ATAmzu7
xDdqzz6zTUnHvNQRwHXsIXWWTtTn5gDtEZJX1yRkPbSWLGZqfUKH4VzO2Ir+npihNtznat5HCT8i
5CH9GgkM1Dm15ImYDaCULNM0wnWkbX4KmXU6kmG4pBWW0FHFybkwM4u9W8RHAv4gsknH0RE9qQYh
5TbJ6iRg9VnsFm3eix3Ro1T2f2FokqdpgEKGJm6m429MOPD11IY9ISHjL7qyk2we7K2aC3BrFLNA
S0EQZKaQVEnQ9iFc5tjrxqEfrCt9ulCIm0MwNpwoLWS2ZV37nK11AKA7AA0+dlgFrvkQbUR3jnKg
eBCzGYPoRVY/40mb117EYLY6dFzh3pgmcG/446O+uNwocE1Uafcoh/EGfl41EuFUm/Ldfk5BCvjr
j1bxcxaBjZrDeU86v+wroI/4YbRhroepdDj311ZUKfqUwrwSaVYXS0EXS+iPZTkIHf15ipgETnA1
NKki1KBvY5k+7cJSl+J9d1RvPhOjoZlSL3GhAxVwyTEVDbQfZkz35UuXrcUvAkkJhAryx4A8+cMT
kZA9hc90z9lNrfOKgxfNnZtENqr5o05eFs0H45Ol+BIpr9koXMpUQOJwex6X+Htv+E9fEAQIi0A0
ZUMnaS5tDaBNGZ4SmD9D6rOPOzHEbPqPxFEC3d1l9Zg8Jto8WT1aL0W4tiYpB27fRSljNLTq0oWJ
GNRdOeqApXlppLRC1iUFTxzXP+bJr5KzDIvyzuhGhLyhGsaOkNhBRH0yiltv9NrgYmyJG+RIS1WA
sIxX4PnflIx5A1xbNzAG5OxNsQRLTKTbWI52LU28xcVJVLiq1Q5ebrdU8E3nFiIlNPOrwd1R3UjQ
JsG9od1qDF8duNsbDdCPsmtbhKUsY5d7K0jPhr4X9/yvjR6rhy01/5RBKwflAKr0Cz6x6btO4i1B
41cIkoImorAhw8RI9t2IKohCTZYXvknWf7j/jqZTgtFPz5ga/ZA38Auv9zz8s1F+nAJi3J2Eq5Oy
pDUPbhgBR51lq/ZXarP+HCoRTsUyLWYcEpYeStUZ7yI4nkcLa5IfWy1DM0ev0J68iIT9j2cX46b6
diOD9eQGp4zmM2Ej5AVh500mUyj/KxbklSPEDp4ZfnSewVAu+S7uG7ZcGufaJZnPacxTOuAOA5Ur
yoCyE6O9/h6YUSd13NkPF7MYXAiNTu8A+LYVkJIgBp+a2zIjlUktRxvcKzQmmViB5royXEI8mVIJ
9kq+FjYGSCBf5XfrJc6Jd81BcuxdnPIG8W6P/9Slz/8X3QUy62UH9jwmXOu07yltOf15intYvFyx
3CYz40WcxCc55UzvqLYvdU8F2PejElGLPRM0PbGyp8PFlicujocVKqI/Vnus0VcKJVWVEVWnaFxi
wvrDd1/Y9W5D9oJuO+7LJPw77450I1p30DkmKgayULJOHASipreoCPhuwcS8jmAGezHFnzqC9eHk
zlRf1AvTZnteMjjFJZBQK8QXvTS+prP/yHmae+aEXoXY1dnUKxmp3jrjnJgRyX7Ljt/KS/RR7MMQ
AfcMlMBsCDlY56sppSYX09yIti3G9XxQ3Hi3fY7RdzbkyXNjrvD/MfJFQrCJ8Ja1ZUX/h3H6oG9x
NA+xBiH1ZJNEjGBCQ5j5QUoSCJnDyKPP3x8vf88COKFeudQX29aPTj1CPOJZXrauZ/xZz2dsTARM
1OLsdNszLQNUr8ubrh2EwfyFwr+9g4aHwuWA2iX+Opt/iEYdCh2A+/R7sWSZgjMrbDnfV/HsS8R4
nXj8hY65FWi9jSVkuuGIJEVaSydF1KQCEyuujtywcrPM3HJCBZQU6mCrX/cM1CCpHysX+XjNCU7T
VGHfY42mmbSXpHHMUcyOjkyZCzPxpHyuLEYD5qIjsA0eoQyb6d9+vMXBfl251iI7nLH+qa2w2j7y
qcpH5vcAx4xpkdSNG61OstxYpord767QyQ8oh7VsbXqV3F1TpIri1xAVE1Vzmk9qr/UhzNLhg9TK
BpPT10bSOS8Y25rUvxafrBT/1aR2pMgVpU5frNwG808Yx1yPPO3/T3TCGNnUaL19OEYLTV66Kjq8
54HKN5uF4NGAvwlSs+3nKHivnoPWu/r3Qzm07I/QKYFh2BYQutqxgbhfFwVX/qZD44BZTfJKEsRP
v5qq33axk5T2mRqTMaAbG56FYGsrtMizZnQ7QslRRdwzbTkWa8vIdkx4/ku7qOfLHDsEH/YhidrU
U60ODVuA0ZcT9BvWhYIYD6Qgf0jvwVWYIS8Kj8aUvVtiJHJ4HLu/Y7H9pPecBfEDrmJPHP7E9lM2
9Lyr3rqEXC77j4GOkP7jNyQqZO39VgDX91hQ1YUhM1pZtgS8f4xbufAC1ww0X4QDdEULk0GVF7wr
oExdSW6zbVZmOzMIPnKU2ZPrsytXx16S8Wefo2y5Xbkw3TIEUYFOibbi2w8tG7dBydlWWfgxtyhE
z1lyseAG1B9Rq34gT54+PXCvE8+k5w88lXAmfuS0MdLp4huax6oVqVcQO2s9Z9eyCpGFW3ndl27L
1fYcjzqG2R+6qLgmr2m+QoTjm1iNSZ4AjVvK/HrBB22OZo7Yhfh9Xr7wydByQd1avL8lL76DGLaQ
KwJYF9E2EH5PnlgTPLHRbOCfMg8ZdAd81SefmB3RF+lSw998FS/koZaPqh0Hsvp+VZJNzTBrdZgW
R9NLg9xFyDO0TBTRQMyJ6qlRnW8ZdRSqiUjnYdMnx7+qGqzBWEeOO2V6FXUZJw34OVDNqCKA1CkZ
9iyMT5N5hyjnSqz4knBw56FIkQw8lh+9aAK/wMucbIbkSongH0eZhu+QSYt4IC4aHQnw4Krqan9A
HsX3dujMcjoY1kDg70O6YOEIKA4sjS9FQ42akW+4nj5MbghFnEonxG4b4/du42f0eeUNdYDY7Bs/
3QkVZSwrd9JzLBJD1VJQy56xmNqGaxWDCuKTpn3QXVoiLidBi4PAqh0ctno4yPAvWQVxGLo2bIXk
Evx5pNQVe8p3ZhB6P0HRkMUmxC9HWzLD34ZVUeZa+Z8BZUuMFJCiqwOlrP0sykPH+6slnAEkVC3o
clm7nmc6+QPiXhrpYIqojczztm+3VuvFh5CXFCOX1ex2vMnJ9lODNwjz2luqV3yyvB2W31B0kvea
jBQAWkNTmz/GCg90IXhBkHKaiowZqMcQJTDAw4fHBPFwFRcH45Oq09xOfh9esMRSjPjia74jLtp0
gMk5dc+Sz7nmqJNwspZtrIKTTPuj+vAJErcGFZYYUUdYBdawDORh8bwbjCwG2yD0FH0AcDVQ4Kzi
aqKtpSY2wJM4+7jNeKEF4sQ1wZinBKeOg+YB/nOTvCvbpog+jd2dFtII55OAaKrhX/2dtoxkRgeK
xUAOiXB21s4IXG+ea90Dq5UzUXEMZlz9pmFAETtwlWvOXfEuP6Cn/bgafODvjMDuijPed9khAj9+
ZIAn/F4moHjvPBGSd1snbHa/aKsCgK9NkHR2pPiolYTQrIZ8OmNp7kBA8kplrpAaDAir2chLYAei
YG3Il9F2w6cKAj27KReqfEZqCpgHK+V1ZlGfQr8bFaJDeoFSYAgurHRnGgBuqq3lHpZpI4DQGN5g
QO6jKG5Hfs99zFiXsIlMxACAuM62VQsjPtvc2xzeevbZLkvdmv5rWTF8ZWyDDyfU6+OmzjjtyjXu
3lHkWSpcecs3u8TPyrqTZGF4yHFJtu5PIaBy9Axjb09+q40+OEFXAmOIz5UgmeRDhTdFkh3REuy0
pi71cypE6hqiFyIwVdJm7QkU55LIG9aZqNq02ZWlNCrHTl8i/bh+AR27NSzo0JNwdbetRlaKfrzq
2UGNfetZCfdRetz8HPn+ITn/0ylWDgvyrEp0qZ6uFc8F05pWVM119hjQ6nui/XVLh2q9Ypf64WZX
THC3nXyez83Nu9eeuJq/YZDHqtFMr4nMO/Inlq1olB4AA07HoEESyvUcXY+rs4CI6vIG8B0NCXrW
Mc66m8OmAKvRNv6cHE/SIBROncvGIpNuKuxsCkRlemQWAC5HPft/uM1agvpuH4E6XANbhdgA5Wh9
Hm7vSU05GThcGYcS8hExbTIpz9gDoDue1j7v/FHMEQkWqmxBBbl3VtM8VJiFfr09+xMhaacojfQE
LqdtlTDUzbbAe5FSy3sCUD/RJy5oLnKHEQJyoffgylqhVDi7CJny9lXGencJ4F7EXaWUXqKTt5S7
dYaWIX++UEAZnlE+4sAdtS/EM14VtJAM68gaJu1luGYIp3K62kdEJnr25nPf5KH5KMXTzlC7TRqX
VQoj+YfFu6rGbvAXQhbpcA4PPocAjIqJOi+1Ml0T+oRB/KVS0LBephLtxfNFd26KBHM2R0SGauUg
m7mt4Czouag+f1bWDMugk/4sR52LVUQn0lr0pBPW2aGcKLX4Y9z9bt92KbY3hg6/MVPQWocifd8d
DvHTtBu5Khmwrdx/0n0rNVnEJsBKpvKyYhEohfaPyb6W0KZTvmnN9UZa1wTnuLOyFcUzIAsexNIn
oxBB2iS8RhYf3rq1hB4xXhYqac3ll3nBp241N46jfGZbGTGapAuxAnVQMe3D1TOvvtmYNBWJNA8g
NZzJUcVGvJ1qzUbLwbYw/fnbqcceY23zCXKanKoXA11iGpUrb8j3hPpUVy8N22m5YIfKgmSKK6It
C2iuUY/X+59kwmjmpzelSHL0/BxbOKFPYXCcgRKuYjJdMAoW6g5eVzEfvVAH70CvSOEao9SmMQ9P
ULwttdCTrRxJ1Qe9EKXdkLN8V1pewlB+DnfMZWt+MUZNdByzhivoy9z1Uhd9f5oHiduT3H+f81Pw
OHI/BY1yKxFBRM2SgNfpiErnwBFU9Fhq2Tv2tBPnLuXwZZgjtsNcnBvC01FLwZi5UWLpEtlKKYKF
icaeSy54++FITfMF4u4Ypf4xT5p73oZevLDCiFnMS6WpbYUidTx0FubEBva3wA+Dmw1W6Ij5aTKR
Hw/fCaCHs3FHfnpYKFbXOPgIYYl43s4fICgxl/tEuCtKoN5rrIuUM22xNCgupKW/6DyH/HDHRP+Z
3XaNHEO856qZPzIT9QQsD06OaEHVrNi7xO3dnWy5REU/7bKeXYuVSwda172xqazuNfQLFK/ew8L0
BvveYkS0n4exsHCC9pj7OgEtjyZ8Qv4kBTh3Ae43PCZUsVRoWwQ9yD1BfJsPRtZcoqud2m+56Mh0
riV2MOKH1YOjsKo0BIZA4JrWv+sLz9clJB07U5MgbVuMsghXSh3OhD077uP2Oxxs8pRpzxAmGv6s
dcfwNwWNzbN4G+wA2fk0bLfAx3WNRdW7UnvfFQmxetwJy0H4GEBQXYGmUlbt2SPY7dcwpHL0bZ06
Gkc7tKNCKV2GWvJM5nTUIb9uGdCxuTG75i+lzznRzd9+Bu/BEUDpLfJC1OSMYYCKGofq+FVs6v0m
abZJo2KpLtQx1cdIckLqP08E9KyPozwKQmNzo9ZN7nCWyko4wxo2lDrMBsaGoSSxaVOu7DExkpsf
AanX+rtOlCFopNhXnCvThes/ZqTGJdcs1HsLK9MVStKuK70i31EggAeNdCrJtvdN7uyXeQRGH2Wg
0VyErX/dmqNFh5HjCV1cyUIEC+aehHqHafHluz558klmp3jXh3npwMItXOXRHKvPszPiLmcjACyO
Dbayr+ItDwnBanxiqnmlKemGFMDYnh16Xguw5I6QB2n5QpI253RWzaA939ktUSewu+m8xvaw4rYd
XpKvwSjEEPWiPJABVGcdunBhKLtnvuBjp519P9Lav2GnwMSCAl/ujQr0mNESlSYvpsttqlIQ48qq
ZTByOjfjttN2GiR7MB3D8bsSziFzy55mvK2B+83ZDN2+O1qp4c4zzb76ME6ETYzyfPfHvfZ3gsnY
22ckHodYVXvaXCK6qAJcbyfQv4DvDDIU7UxcVEmoHsqgc7afXIdX6iFr6P3/oB0iGHMqISgapJdm
tgnRiYytmsLdy1W4wI8b/mhnIM8G/mkBIYU7YB9WNnvJUXu1frkIrRj/RmAJK2Lv/VPEhaPWmdtZ
KkVriuzcLABTo/OEug9Uowg34HPAgOtsJTk/kaDcSvzRnVaC+sh0zjfgnSwNLhrPGW9LpAn4axbl
g+PHojenCHnv2Dna9ARvlcA8yCwEigZ4od4grJyrDpFCdgHiVFW4iy6ptbv21bBpBODFurSsBXzo
Fo+rj2q3B1jIp97+c1ZQW7snu67tRuN8dy8cAsrVUuJbxRGWOoJb6B9sg98iXazgvrTyf44wFdGe
0fEkAoyCcAEyOCW1kbGYZHZchDZA2nkp6eDX//GwExl9VaJccn3/T+6yWe1IqcbqRYZtTyCn0zR6
/PuLjPGGdKeKDY6fPr8rlufUz6Piid81Vk/tO+JZ1q91LKD/yncTipuYXaxGjXOcDNvF1RmNsMVp
7WCEfFxtDLGSLISsFUslNk/Y1hVn1sxDc32r6PWn1bhS6fUBYeX1rU8TlDeC/97f0b9STnys7kho
yM8y+HUfy3FsWCwwTwR1DuiEa1iTJQYoMRez+ZY+6m9VbXy1EwTxQUtNZDPJ1nw29XkH1yhNkLTJ
gMTZKosG87Zej+48VPdrtv3CmNSZZ+Uma4ExcaZm3aocqMsQ6u0Pcjb6nXjhLvitsdX1tcw+dwAT
E2h315d3peGl4eIz0KUnDbjkt2ELAXVMqwhTAGVq7fk8qrBe2lOh0au5jyzZVZ0eLZN3ZB20BQxT
/BC5GtentxKdFVLeIkJnaD8RfPutY1iGmhChZHY1QpODyCuiZE73VJIOP6YpByQtGaTTfI8xZzeN
JExLdCGF/lQgG9O/Y0/5EdyPIzsmCgXJo+tuIpgTIToGgQtjohzhkt+M4rsCf3VORrTFZKO9piMe
sc+d5eGk9DAOF1Mz3jHXx0LPQZs/8mvzmA9eW8+GWrOybAw7QlcLMOVI7wecGNwwNs3Tl07os7Ai
HaBbsqjFazmru1Sz8hCvf55u38+708jCDGJ9NGne23gV56fkaJbf7tJUdwn9fNlW5GfmcmLwC4TQ
f5FJvEikrlbTi8Ph+7MdgzRJ/QxQMpXZeHFRPCdIZopQN8nOlgPM3T/IFwO+9+YA2HQ79kepTrJg
kKHWQaHvB54wCKA3p+hrmGHR7Gavc5c46LKqCyqINrUL8/SZaUmbjOCBaRsaG7B59hkzf0UG12As
d+9v96S9YfMAPgfZDMfN7Pt/OWuVt7GS4nJHV5RIKBmxLIMuW1So6ijOx0deiyO7zm/oyuKG3cXO
of0fhbz3FUdL/akXHyCvns2prmRREE9kpqsYM3ISVTmQ6KX87KOeQ+qy0PS5riOJfiucXp2A+zjA
EQxdrZIcRqjU6w+OcUUmFEa+kAU9rLHSPty1DfbtWiaUHxN3RhVdTtU74NWAT7U6M5yuLkbu5TM7
UoiMQehItBO4EWyt8cAu5XaWJ57PeSIlPcZSAc9BXyZg9HkNjep5ixr5A27995XOhrO5aGkx06IZ
jiVQmzmFLakaFRjDiKkUSasaiZYnL30itpXnQ4EicHQWkfywsMcmOkW+m8KKOrbhR6+kFnklVr/w
4DYqAn5kPqeGD5reeCzvk4PPpM+kEob6qt0wEnh+T9hb9704OfXm8Jt4PRv0ePoRWCGAEW3mVdx1
UNWaFsMNY7HTRhtlPk3MFZpjQFLzicWz4g354raPCvFujhOSIbCSo5f+p5hv61sv6c+PYv3iSxDt
DEmglWFhq9khIh+WD3vCHUzjHcXeryv/tolUQxQGwG/9GkmQjg5Rn1B//KbJ2nXNuClhtn1s7+oJ
BFal+fCDrHpl5VexUZTW4PASOtdYfqUsHTgoAy9eFHMBZrZmfuwmzluqpBpvIjGIo8kP/8bGQBg+
eP/cFmyCppsTS6yFTqqQoJ4WGygahAS5t5XXf8uqMjJzgP6QFVXJz5+5LchZgT4/Fa45OOb2UIcE
pCP0jxRKDkBYrQj7yFYcTbr65uvV6vvXm/7rx/rxut5SXLXMlB9DqAJBMr7wzgVMttNePXOg2+bf
sSUJu7hQcEYmG7sdkXk1wf77dBuR++m5AiLnZ5qqomsKaJ8sx1jJ7zl8Ca6gy3udXaTuXl+MkoTq
qqxLFHBeNSqKJVTTksSXed8Ez+5ReNBDi+XsEtVV4mp450hF6Xg4w6Q4KWlrTkr273AwHXAngcvB
n607jJdZr5oUzkXi7BagvKHEIhtY5/aoRLP3F521cSZtvxTPCE6NXNetBg6Jj0STPFnLjjb1S9Pr
YHYhso3t1EPFf/0lEb+2TTlGw2EbZp8VvrjksOLSw/lHM9AWOU5pluuWZHCcROS+Jn3dE53eSooG
Ksipcx4eOHtAMoqzbRtN25LA5cMoFQ3s9ZObA0g6KXSbS1J7g/EO+ZvlkEXMIBQ9I3T4+Do0RvzR
jYhUA6OhAOB3lzdTvr6GsElu/Y2U5SMM9BdZ3X6kcZbKfLQ5p2MIUBM4UqIGrrgwnPVCSb/KtcW3
fi/ySfQ+q6iIChL/TURjljHC9DVJHxLJZtLnle/gIX5QlI8iWsbTRVI1ZQX+FbPrfMMuxMLhJHrk
FGBf0PZu948kp8HbP3uo+oe74ZE1ZEXiDxc22QX9TnavnbrGJRjPSlR00+gptbe6uZuO9KnfFuBY
yXfgPsUT9fENsffzCnlOuNu+gKm2Z7TM9UnQx1sHZLlsBC3a0UAV/lwXETih1PJy+ot/0z/+VVEm
z/zGWSIex4P79x6uttBBNq26uztca6/zqpevopecUI0N0hfF6ZZMGwREy+B7uuJWd/r2/qNWhGIT
1d9Fh1Z2/KsV5uOmGYVqw/wxHBv0naHJ6nlPA3WXCpSmvZOWmCTMM7ez3TeJ0EUrMGuk+38ncm5n
jEZ2WlxfWacjWgOOFsz2uh5bGdQ0trefxpitqhB69e/3BCYzvd86A3bS9ZtUbAcIvXHQIZWw4HP6
OgLgMgfH0uiI7T3E4bUkqV5ECKzSKzZdmDA25vQyJ15xRdLySxK2U3WaBQdIvmyWG3JbsoddnbIc
KaXrSnUBKrl9XziRIAHqF6XYvxotuBudcHXoYRCCSmDQqwgIuYmK8j39klqfPo/wDe4D3DVFAP9w
lMOUJZYmOZnbVw5L8NABGfgg8MKnnivNTwrQDlrlkkNTzmCEB/tjFxtpefro4WELTg/Iea4cl9TS
DG9qn58JVrhOWqERi+tC7bWM2fYzooaKwOJKt/r9BQnRvHUes13Oa9QkTnJz6RuyKcgTpSEyopW6
+orDJNuKftCHpZm+682JbW8js0ZNCXyiL+BpAZGQi5prH3yKfE5mwBYV+Lo1S/WDYIAxvuFzqgGi
9vratz7otuQRFUnrM2Rg4xFxyWSOf255nYzAvcWvb8NISVABgLe0kY8y1mappY8A5Zb0Xr/whETj
fzEsn74GGjjVldUnoTHerl/CKmdTQKQLVAF2piN0YmZZTMrPrEHi94YSD0QIIgFyW/78WCljCdB/
FEbPXwQrDnJCqbCSRCdK2n577tx1Tb6kszN0NWpIHmy955VUK4qKrV/AHGFgnaT7FFdNYc66sSV0
gDQaAc3ICx/i91iS29NkL5WnTDG7ooISCkdG+Me2uddtvxdFnYhqXTSfd6EkWqAPHcsEyGc3gFup
xUJZyP0ZzBn1SiuWapNEGeeWSgB60yM4bUMYq2hM30Hjxo8BsjDD5sih5Xxtk6fRTrA6cWj6Vxfl
tntmlRjytDxuEyXXDe2erDcyFI/UhQSs+3O6GbyxKRNEbawcPEeGqoSG9Aqj0RNtN0tZ92iqd8rk
rvMYuNDYQEZjsUhM/rgpSdOReQBGumwhrqJIoTv4Cok5rBlEFxGEEdQsGkIectU693djyNQgDeqm
uC+zRuYgFEjrSoj1yZ2GGfz2HUvve/N7JbiRlpMy5GM6YBS0zZDKE7ABxkKW52U01s88i1WyGb0h
bH56jnQJavLxSncP7dX15lbN0qCHZXXWRStXfc+9AiJ1d8mIIfoYjR/BiE08242a4LG/kbbgRXwy
Gd6rfJWLk5wZAIfuj+zKQW/0kBCnG4GhsY4NdQrNvL2BduJRnOoH2rUQvEwBdRlZPMIqEcwzUAtu
amLXP2gDYg5p488QAOA2fUAMY8QjRtkd6QWX/AW8hzht3bEMhAUhqzSIvASZ1ecZSJTHcZyTcUx3
D/BA4ze6Uyu9kPiAiZ5FjUAtteGKn3MG1ge7EmnyfIm4zCTscM2tngM1oPBkB1Agg8r6eMIJw+t6
HOrzlHoqRDpMI3GZD3Bh4B+pUjNh0MpB2b9eE8fvCFDJepqoA9fwR4WCIWbi+ADWSXb9xfxubgWj
HJMxkhDC/3dnAI0swqto7j3NQg1VfRSJgf4fYzaf0KE3MZq4jeBR1YVgjbD1ebI7YBHvzPfzdFaP
uf/O/+oSYn63+7Z6KcRKqHybFljsKbucWK7HNZpLP5OQFhRbyi/ZW8ZQ9LeG/iczVsKTkQdEuTy2
e8r4kpWy+y8spKHqj62nmL/Qh/K0mMCwYTZ8jMSDE+EzV+kLjyYb+bayBstkcabs8vy+XGpNmxgF
EjrHpnXZlCAHIko0GAygE2l6IbBrvSvcEw6XGTFE7V5Ey9Df5NHMEa2qVNxYClklQk2T+OLtJPVb
bDg84FVcASI1SKTVNDMpVAuhp+0KhYAEOfWSpsbzWM6NKUqAQrVsQgdFfDkjNASS42hfh60anU4o
4hQQ483siFDEXZNkOs91/XVW/FRdcUH/TyHyT7QSgNfi/XzUZQpnKMS+gBM9L3zFWuEeCPkQMUrY
mGS2jViM4y9PRXDZqXQZvHzojMeqZu0OZlIRMJO/OgrV++JYq15sXKsd7ebapt8LhBxd670X4t8H
JKwrnQ5F5MNj2FwamlKNKYJQEOwgNSzuJowW/eojcQu/9ej8wOQAhJszcbh3B6EwHUmcClJ5yraG
XY73SFAP16j+O5np+GYH9MV9udtzqd1HyjZz9QBpliPumEnJfJsyVtGZ85KHVzxGITRuERDvESNu
ZHKMVeDGhlyMUHbAVjUedDzFBSMTRXkWJOryqExFqPvFyEF9lLzdAn7vcLTU8DHAekokNr6CeCWn
B++JCN9jrvv8O/0+ctpbjSL2GykgiTlJDuAYGh7yqY2aZ5SBk0rH/KjT9kAIhszLjvZH0Fkvfkbv
GRrQtFf5vSCFTpcn6nxBD8o/kwLEN+GRxjMRiJTpqFgIzafTC2Gt/a+CpzQ2pPCxaou7FHY02e4b
Hawm5Kd+pXOCZG4bJ5Ms04xHS9UKwsyB1euAhNgpu3Dt5oQksNX++s47hJzrJ8qrcXQINspbD7v1
SEQgiart0yP0PgdRb5eSuSoLEH2J9oN80SNjMnLUHZj/Bb1qf75nGZkqxkfWwNRC1xeJjKQP/lNL
Tu8/oFSU4k+5AvozVGu5rTSCNVLuoQblrD7yI/eO9VYKRWIxQVoe/CF5mokX5L1apaCurxWsFm+d
m7TTsI2lX91n5BvKv0AvhCSOYgOCDie9fPTmOQPasdimWh4lZs8vcVPEDL5gh7yduBEd5Vq3V67h
EIR0wVtL+EKmXKYdbQXzXBoYsg5+T1ZyHI4GluTNFkN7c9eXU5FeAoPCV0dqvSkGbKALJNTunn9d
HPNffiXOQIMrak7qevfgV4Q+4IcqcLdLewK43RP/Q22RHqOA+4wHU9aP3ZJhAjjrcOa10VtCqWlq
xDAYZkfkCKXOVIIvQe7C9cMh1061H6c21VPINHlD5swVttOm+QepZLCvzNVfL9VUTInk961T/Uvc
GtJMBawXWNXDVkxldkZL1VLPQl5TJPEDMg9aUeIx4RSsPCag83oHew/E8xtXBwFx7RYFe66CEaeq
TlZUHoJPMvWVBYDsqkuk6vl9tY50vgzw6uJKuUplarEj7PUgBg2qMG2CkPi0XumI/hR5QcvbDng6
DQR3wCHFz7VA78ayG3aPQNNxG6PrBDNlUCStUpSBBgCfZpCwS122dGEoJpc2zHX5+kIZFa4NljZq
Lj3mYZzOQEAWK+6Bzy4WbSlTKz5ESYqrHRiC4/6tYRDe6S041k7NRUkDMr7GR/z/u6N0tdJFiTeU
DwzBcsmVKmSvDm3NHwkOt2II6YWmXfogL9Jm19EWRkT5D3Qz6lpte7ziDYzzzGTKHkdH1NaamtOp
RLtueyZH4oEH/aod1OGlp6tVmBBBXv58RWXw3ln0d8nWASg8WTdzhGMK3dJOAoWMMTp47gbgvAMG
1bhrN4FrkywHF7TI79PAdyJO/7OVmkJKdedmu3fpkz1d03KYZfT6F8Mc5O6xZ1c+Mee9IbpVk3WB
soLFAbsSHiROG078BDY1n0NI4DDhI7Egqhz8VQqZZaYEqjeeejbEX5Ahg9avJVrmmZ+xx80DkUkb
VqGReqMCTP1m3ClURfvB2yE7MSYHdoINWxksrDt7zYV+aMJF6B4ts61zMMg6aX2mXoA19EpAe5UJ
bsV54Qc3YWdFToetn6HxuKQ1TuRXW8JO0oarww8MXmX8sVItEQWX4NRnz2dxca6Xafz41ORz5bMU
oPk+TAk0DI1OrrrLJXgqHJbz3ryNHzlmSM2IZDoRfh46kCX3IIOao0EsflxNKM0Lxysd8N5Bm2cM
hJxY+qkR4RkOIp3k49pLcjWfCzY44BUpJEMjs2OWwTf6a+ppuBrdl7QvM6LZ73uf9DGWwklizOx+
l9nmmBBgqx00aYhbjuRh/y5oo3+WgyUQmJYAfqcEz8IBTKoro0IxIV8WrRod5owbqwzkjDIaD4/N
TH8VN6YdIYS5CVJ/GMLtsnrC+MW8gyIYG7Dit7AGzXdyiFFt3vvBl+P+Odr8k9PVIm6PBB0Nwq70
+VM+kNfHdKVy4fGgNdDvp9HnW9VDUG1raSPW76uDp0OOdyfxNnhw+ujZJoa6RgbXrBY+DzqRbOrW
CBYHlVq900+ncfmjVef5VUGJ9geqUO01XCOZAdzg70YbWKN6kQHgu1SlYcwdUxuSodUKhJ2SUWZ5
WEIAlHhyOfSXRtAtM4hkAd/5itG3at8gmDoyk+YmneP0i0kaPJ3WIWWCfZjoS8GBODS+RxvJ8bi+
D2gOf55UgkOBy0Mhb8+0p5HWwn2voz7V8OzS/XUhH7NUktPzbZ16cM6CAo1qSpKUo0RrY5WlO6YS
5wrk1SQhEBbxd5/P57VZpO8qIi++OyQ7BaXZwBXtdOu/A4BAsMfCvPivi218JfHwZaqE4acTfJXb
4UCDN+z7FAPISSrX/ynhGQ/cTdVwu8WWboYsUKcZ2Zq94onTx8p1YhX52VAHdb9B8DaNzQJFi0zV
ZRt0HtUXhhJt/eb/2FBU55cPeIT9wW3Dvd0ao6IQD5WNhL4H3sHUIC7wnPjmdTE+Wh+c+sbdf0am
YoPud/1iJDYnLBS72z1sut/NU+UNP1wMzvjyOW8Om6T8g0sm918sYpaSG5hRcZ97vP36iQdHZjUZ
BCeOqZhiqNV68S40dnP9QcWqsqEclcazJON5u7YkxDtxEQmtm4yW0/eVzoniDo2W3IZP3Cv8Knko
h5ofYQSLPKDl6rdLkmCIGIbCGrscs0hkRSLAHu0rPKx/V7XX/PgqxmZzfhLNU3ThuGi6t4e56+dG
T5GUBnV+F9VnZbFAp89LobdC7vNcsLHLDVwK9XxzT2cI9DJWDei1qoAbTuCWWbpWFaZ4jyJSv6Yv
8tTbyNfthASu1VQ2yIXTncf90fRX/UnmOMhbyc65iVIVJXbeUO6D6qVJFiawQ8cIyKaWWQ/sqRqL
Ha2OvG9RIgcYls/IILXSgtlnX6srjZ46j0Hv5mVFXSvf8jTzOxlhCM85a5voAZqK95mWNY9t86Y5
ODy/X2dae9zrw930C7onSEj/9PvBrqbwLJLkVJrPS6TUFULRk2WTtsBBuMhQgZcReOYjLvzt6/A1
EY1aNS0u83LE8gv3YNe6oAV7+8zxYaR73k/PkLWNqiPqqnL+WSMBvIP0FNMfZ217dAgArqMrl1OS
RwAirTVQ2Ia2AtURrDGrq012A869RPkasvfH+VMsaFQjvHQ8KzhB6/zbYo0NbjGgCvcILl2alVex
McFFBtfwnPfI8DvJS13KYxIH7axKa8d7sSlPj2KzH0hN6jrSdW9jsP5cVH/r8rzgJhGcQloSpLvJ
VziJjMBiUvfnStJq/YTtb+DIBlIQtcIKCvv1sgoYehX73U7dK5kJRYiApHqMgvU7I6asdiHoSmjk
eL5QMkeOdT0qR1z3sFVpVR14nLzYwi4XG9i6oHqP/8ALW7s96fw6VKFdB/9sY4xc6RhZJ7c7yoTl
4HZQfs54TGZ6o+uiKi3Qk11RGv9KkpL91iDC/wn/OYN4cbd/kA1jiDiTlpzyH+bFeDj1XDizqow1
VbZPSHKsz4o8WwnbxjaWH8hGlHq5UEZ4+K4f0uVlUQ9wadT1Gwbt4449LNu0l2OFmUbtq8fwM/jz
YpGXGkmXbML2gjVTWo3I4CC3AQY/5GrZFXUIHiNrmiaG1xiZgc0QUdgJ5+WEhkl3WaI1OXSWfiJt
SkRjYVBXF/bM0AIJz3P1f31I4J0FVBSWyvcBar0mYoGZJgMsHiNya5irgXEbg3z3WDkSLjQi8YDy
WCe2qjCfDIjYtQZGu184UrRhamhZ+uRHWZgKGsXKchyGY+dlmRApjV7rlWIMJv715chsc9WsgUNU
VXJKjCWheGtFrwSxjUenFWOr6uelgaMb0FLxegCsbTUWyUDCW1iL97mi3ROJIZfBxLJ8MyJgb/En
WaqBQagEF2BEn2s5oj98n+EtPg2qIQqickhUfzQszvp3Njy1HLI+llLKa4M1wwUdXz1y1E28ixFV
SGteI+k4xClo9F7/ET4YA+FZuVHMzWJDte+hlOGlWjLzhsz0Ib8Zz3TQWchPzbQQz3GLrISboMeE
NScuhWWgEfTNfVha1oSHY3fv4xbC2d4XUkWpnU0+in2yUxpRecAwjg5G6fmkdyKcAfGJxPbD8hwZ
mio5dcsAfnJXM+HIq1S+30mVlW3D5IRR1ksvHS6wYR+MI9PeC++w4ot9tid551Ya0rUMr00kYbsw
cJjeHEVp0stONYtOzXcWB3zDJ2zgawKzUDm0lnogRhw8vl8c//gaZGwxaJedihCwPQ65dMiFqQ9j
NJW8CLxRZMAmvvCegucFcdHb2sEbjzvG6/MDSsWzo8wCJwG/WA48HZc5cM56z6gpFIWnuQ3NLLvY
A+auUR1qMAp7a34/pOF4aAB5WhxKPLf14cY9R3VTleqT/TNnQJA6ClYdKDZ2VZrCyjcNLVbMgr1w
CQPbXMFXe9ZSxaA3BFgUMJj2BJr5bd5X2lyQrPYXMzK1zmcMAwC5PL4L3YqxYP2D/UYEwRZYHW7S
N4yg7vjFqFENupXzIulWEnVDiS8EinfykoIbosCiUU6a9wMiQAzKo9ZAYHXnoWJ0PS3AfFs+xKbL
/aIFCSaiV+yvgyp76h9TbN79PjA+jEoM1uSTgY4SnxmDONyDLVpXIe2f1Qs1pzn2mj9s+f1pDEhK
fLCfgDhPHKBmTEdFucTQyJt8JtJ+W4KuxPhPpUywcVjDesfWacjTkRYWUxynInZWmb8lCdT1frtL
moO6cnvIy8X0F9xC/j6q9ZSgY+xuvpMrz1LuwPKa1Q8PGU1/Lap1OEJtMjqEKF8A9z6Ye46J+nMe
0FxsbNtG/8OEuOiMiBuxJqtCKNdw3PTfhH3gPcxo4UiSUKNDvCCg2QLSP9UOTUTIyDBbgx0ht1eV
5Sv5xIEaT7LGijfOwwJlBqC0Bvbw3coh3dXZVhg7v5jKYjnvtD08TNSqwQ6X5tuRDjRsW798apCw
d3BLBBChV0YImsmBnl0PH+oKM0FVdn8VWauWBxep0NG+Ve5dyPY21o5Q6mos8ZuRS/4SaS4HTenu
G5I9OI6eSZWPEGHvyQxwFjzRTaGJLCp00sESwrBQaawzXlWlY9vMPghoZK0hpyl505BBnTcznHlA
72djvr1EJxJ9U7VpxvLAZK4Xm7vY9wfxp0QtEVxzRXBGbFgTXks5yhnGdezqPbVL+29VIb/6Hq7Z
N2sFN2zoHSyWIZeSK5iOCK7ZoJWBKxGftPh7JQnYyMQrfvCgSfokH3BtYyESFXUOJyq7ymhGEz5N
cCYhav0emssYoxuUAuS7UtGoDzwNq8Lxy9zUYxe2QhLgYW62nurJrHTOicHYcDG1R0bDcJMTPjg8
NA1D6c+TNA6nYxcfHdxU0JNY6Y/XU/PsnlPvSmZpwWtrPg4KneCs/Wnwk5lzoTxHBniMf98dUfrU
b303WFb/bSuQEpSnHAvXrt6vm8spdKszNy7SBQ6ifzYSbTkUaRieo9lTMRY+m+AEeVsd9kxOBnJP
IBiBhoRwCqityNDxKY7pKSGVmVk0JijkBlnEC1ENqQmCt4Ivv7aFkIHU+SHebl8CXOqHomGjUAOP
Wql14JPyjAJy1avon9gKnEJWrA9NC2wioSNnQQsNzTLesAG/rh4pHygSHolB/nk9ywMiJ82N4f/Y
YGBvgERK6PSKIYHSCBfRg3A/WB2GDOWXuIjQ8FpxJMsvvO2DGn2AW9MRFJe3txlWvrApLg7qSXGE
LL8nR06Sq5QwbQX4vOtbG7DJtTuxNxguduITD06cKkdiFMneZUj7D1morSR7Kopa1/n3yVF0ZsPe
1wQGTUHpGb2e6yjdvnBNECqgUWJ7kumHUCOn/DVg5pvXkXJWDuli/8ubPf/OH5D17S4c6PU79Yth
DqW2B0SD50dTKMRhhF8C8I+5E4evjGwxh8ijq0QDcmA/DMquti8NMsVUqlxwyigaMbZFIaZ89FAc
hscyynsf8aaPq2mgXACZGInhP0vZ66N8saiuZd7yQ5wvOcTwP5mS2KUGigae4ippf0vTOT9ziYxv
cod7NeH9yfQvUCrWo3aBBriRiZlygsMs8+hQ8VshqKiZblPdrkQsn0MaWOvoVSK7gYXWzXc8p8Jo
qr+XpBQFItmm4EbYqXnh+ZqCtlFIWfK1tPN32ONze3daLTjeNba0uyl2bCBXKvuvX5u0BsKPXXp0
jl/nA30oyd0p3rUHoH1DjrFiDDMRLC0gBcRHHKGJGntHbY2yYWPt+7WrqKog2EMcxDplke6pvGmx
zP9I9FzTTQ4eJk3ph1MRHeaNLiI8X6/fw5PiA3YwJ9rwab1aN6UOG7S6ScgK6hfQ/o0PjvZyAZtk
zA2KKeGevaCdNwFxZ/kpKqYYh9uaNXjtZG5iQohjUlH1o3ik9qu/FuTGApsbG4PnAPQDOXienNyK
5qwet5Nuyph13+qgzbfRGwOmsKsxUvD9pR4G3P5G6weNWTpfkSAzMT0UtNASscW4lUtW82w+8ZWT
sArqvjEzj1MHiLkTfKKLn+tAYb2zTh2yj37WGLb1JlYVH5T5Jv8nPJXWOum83zex6WGQmHFV6DXT
B1Sa63tewNrS+bxlO/JckfJoKIAP56rBX0yntOhNCsEuLIgSZ7XEFvPl2E4qvebwwY0J7yAOlpXS
CQWqoNvU+zXDJvPvz6DQPN1MKT9j8H47DBMMJqSEunbzslSOWEVbS9U8uXz7XYuQ1S1t8oed5jfC
R1pkALEjyBkNbM4/v319sNDdUX6HvUEoeIqI7KT2AnRwO8U2j+/dhu0xRf51G3X6hMxzCCK/k3BI
LBH5yKBqLUX2oDtF7oLapiaSNr4Psm1ZXRD8XHUAqOfcOjsgptCD0DVHxSDmPvdj+037Stzb/XPa
Z9wm02CBoK27tnUF8JGSQTBBTLAWq+bEn/KvOpRpQGZOfTtC2/iXVYWb1q7cstBz2ERpdXx1FcDw
9d3ijDewJr9gqvRwT1z7BriJFn0IMcg8WXxbSIY679wNbXZCIDgd4/+BsJDKDTjFejL0QwQ5WbH0
QDoFzp9GYwWknT0eyR0ArC1r5OmgzGUTkMtqz9QaKU7UMf+TQdyag6XRGrXQ6ucgzYTuSo0xS5DA
E+3+P2YkW4PJu47qF3PVe2BYdSrY1oTcexTcAQynjqOUooWrilBrG8/m+aoP9B3W7psy1dnz9xRv
crmBmgStnt21DsD/d29gKY3NnLF2QFxYAaUCeh5zZ5fvKjpVR3umcuAkHEgIh26rQHXjW1kegH1S
qiWXZQrFGBv0s6Wth0Iu5Q6QHyEf3nALSjBYya3yfkIwWGsTphXpGY7CILn+w2qGwYTUIy4BbolC
jKfMwTiVLUankEGskqf6JlZ8yJTTVJW+Pk+Z5/0ZnHKINFEmvjmfY3canmMQIToGupHCsq2U1LqN
wUlWhaG4mg46UdUE24/afwDJYtf+YHutd1RK9ALKYFz/rTvAS9g85TajYRPVM2prDbb8rjNbPIMm
yGAfIPBqTcIbfRFaiD+3gaR7Ch8n/VJidBhhU/CBJFL062xC8uzSTsSSRABbyhT5Lk0oAVV5g1YG
pyIF7yU4SkPOHLiA3XyY/9rzOd6caYo1dKWlI7YpUl1VCBG8d2ckNst1OLCriNFI5+4oH4kLrolC
RKj34TL08nGZEcpzCC1R5Tri0b/6SQ6U6EWWCozTfOeSD1kni7LOeE/+6g5NWXN2IWa+ge0Acitj
N2/bhSZWG53/BZawRWDPWE87Cx4X520PrWkpK7rex3bb0ZzQMmNGxB/hj1YF54w0KALZy0hwizhj
X+infUINpIhXXA9RjnwVQQYJFIiREoF+9GY4SwvBUhjQyN+mCOjPsMA5fuvs/u/3Ou4EIKoDvTgM
nmIqONx6PJiwgBNt3fxgT7DPoMJvjDcGLJIUcDhkI2jLUPX27z7jUZhUuZ/15adO0KB7Ua1sQiGN
QqcfMFDdVikEsm+kLSsGv34MMFPCjBUd+yRiXdGJLJGBp55qnkDKa9nGgTWfd9j9uXiovfgE11HG
Uyfrx/3DorhJQjBTplZiMRg9r05WOhJgW85d4uMYOp25am0oQTH8IZt0e63HArxp80d/Tl3SUjpS
Ij0Uw5IFpvxpmAuKz5093+ca3lEcl+G51pfO0MJsgNj+RfjDE83r+vO6yL5wcSlLGLVqP91ID8in
YoIt8ptwFom5sPVXbhoU+thMqRVJO6aIHpeHL5V+LpQBkBIHdEQPw8lGzOC1+86sUpFobJoqOE89
GgrwWPlLVraUFGZKBX7I2HF8dPM8iUqU/irEf1Ybf2XkB+jFH2HKxSWC9qC47buNQimSU0MG0b1f
jDpwq0TAoTXgK2THptDTYhftqVNRwLBtUZV8Q8hhbwrFjKsBnJeR9QNX7YtVppDrJT9wRv0CRu3b
+YIi+y1GLXlGcn+rdLZfZUBd5dalEBZLImYSyPWDyOozjbaOhRydk5yf85GqhpRP1/Q6kSD1cMCE
nPSDfy4Rrx/j4TxRoF1zEbzP4iN72zDfKIluSuxPdon6RVOScvtk1hMxSpgXX/Y/T6EuIzjNeaw9
UXuqT8PmZFmSbNUUMde3h+zzV6Uo/MTdMwf/XlPHNM43FwgiVKxn6qrEhAV3TmQYMjn915RQpEH0
LjHAaLkN1xT+v46b0o4Pwyfx4ZrIIXEOovRb0nbmgEWB55/QKTczz05nx+L6w3deAEFiTLJP69TT
MXtaY7WqDzZh8M4ZEFKZvySfD8410d/w30e+9OUXOhTkhmxYtoVNtawMxPbNWLed4aGUK0pj7iHH
wLyqtx//l/armo58dZX8Nl7IcqLUVehmOVlCL1pw1sPJD67VDnRMnd+ZBYxZ7KXSWh0TUB0jlTiQ
+QQgk5CH3VPE7lWGRlAsq7qMzObrQvk0fezd7FRTBF2NRu4XASKsGP+fBwRiGajEN6v5/hkO7dj5
DTcGChWfSPjskfJGjEwwo0WMYlBMRETPqq0jpItUeb+YZrNQt9BozspBH7FHn7I2FLD07X77frvJ
EdOP1jMqyclooO9otAX7by1d5gvnIUTjEbFNdjV+4zAN3s5rpJXfLNmzVIbGHz4Kyp4u54nW2MYq
yp8CnY4ZpIi3AhJx3jkuyPGcFvYZZttmCNY3H3DkeQgZsN80YwdIsrWCAtgg6JcQtIpYkSZQp5jd
MdvoXddX35ezpbIn8/r8bxAeRoF8ZecP5IkoKsaj/r4gBG9I61VfshAOVztZWJcRomrUlRzsG3T6
5OOdRFmctohG64aC14tM6KGpgrcGGEiLVbp6V0obGysSyp6uQEUzVqeJojHMytFVxIT0Ai0cTMP/
XcbUAaHw4hbc8T1F6yY0cM3QEL+PIFEMqC/9SyssRJvlPuIJ2eZKxjuknK3BlAsMK098R7q/ZVlR
N7R5wN1HXn3sTWRVg+DVkYkxr5h9CUT4QESCNxufV94djaCrXMLW04BArRGq9aPvLXMmZt/oYWWM
ufH/s4I1fw47IISHIBHn82A9KLSGtwjIUyJEnnq0A2/3xplSkKk/tqSjPMzhcFIt4H+uIhjel1K4
DI5cVPYnWXm6DbymUnwxsPO7Ou+hT45eeGfBVq3l+RPxSq8qVtYhb3xcD5k148Ssh2jFMVt8Nk/o
TYLMai0YqcfovcpStpS8/bBn/z70AosQHtVI0dArgrytxnOcc/NCDNvYCniI6Wd/RWTliE/h3bWQ
YweSHeaL3Frs+mhVIeVVhq3VV6DcWHhFz2Bw/U46U944qA32EVeYk/i/L1lVnixWsRUECoNNJ/0d
LpRhl3rXPyOdupK2gG2ZtIAFdGXcaL5SSfWqxcZVE6Y3itg5bsHPGGBQA6RZvPg28N1mDmwOBxid
2y7o4voBfDehGHTEQoI8T4FPMPdxgVWVIWYptT8Edha7QXgU5kTT+lUBroEtmAfUcf/X8tqAx0wQ
AYXr9ZRY+1qzIYAxcvWBAClle9f6GYE3UWE5wFJtrQJtKE/UdcLcFskQjRfDyGPVyMXOcizh6bRl
hP4VYtRbUWVfFcOLhrNPvhWMNokzInirEwe3graCCcwSfiKnVQm8AoOvMOhkU0Bt31JnSavE4x4s
nNvAcvbzMb+C6+xhMRZLu5lKvDuUPwpXHKT0KFCE7Keum9H8b81bJEPpaZ4/aaWTcaCQ+D4y8Rfx
K6vzmez6bV7sO8qiE9ZfArh3utlJzokNq1Q45MWwph4DUzvDfZdUdVXah1p3CLLcTU3KlDYRUKSO
pmL4Yd18AKJuS/0wu3xgdr6/hqkJwuekQf24X6fpHDo9/GXCBPpwmTIvJKhItt/Ul1gDem5MN+QZ
LChuvo8KMDOMvKnKR5mek3cH2grgPpnk2UH8I/9ecH/tKYQLNM7J12FAjFjtmV6j75x6Rrs7weOT
qMMPNyZFXnuaaWADi9zj4lFk6mRL6m9WfnZpeNHFK/qmG0YJovhy0jmsvGlkN5yTHh5e9D7BBEJS
W1+Rn4dF3Wt7xuc2oYxJNzwakE6tUmuWB0X8CfMxfYwdRqfuUBOnzS5YEg0WE4/gqesn9HnOnuT6
dhtgK6JKMgpz5sCK+CqiZtc/i4GM3uwoDL9RoAD9AUIxcGsXBxf0bFf8ZiGq4lkIfxYWwxmr6NXh
fHP/wbYvn5RV8mBWcqVMiUVy8TNZ0FsOEIYc4iNMYTy8CTlVzGFaPWNq108HM75mNf126w6MVpAW
6Ky1iKboC64q6qtYdxYjceoOY+Z7fHqIzeEdEb14IsAx/Msp0SeUkxIbfm65568JKv/hk5uhAZuT
wM5hTHXKSvHYaPeUl7SyUU7DWwcvmYPmmUUugkWaMn7HbFrPWV0+hUI/b6uVMH4Pbn8W5TMzzciq
NxbCW7F1YSTi7dKUN+5jnLRibm8OiCQ1IKNRuZSOdndu1p3A9HWN8b/zmR4dCWQ4H0OZHvjNDCB1
Ebio8O+FolB70NUUBbPO+MCiR+o+YyvMZLyvETTOwD+EWmT613F91pLPWbixT0WL7ergFp6CenlP
nRM3u5las7Jr+UOA3n0yPUuVal6HGiQfeeIgSXLR0Ll9PJFQt1m+Bljr+7cBB83Q/uFMWnH4MywY
6OZFjURgH9wgjBlajao/mD+50J9a0bDZDDSQZKVMfRTbDVphWFusFATCxH8Bkpo9yNsMVQQWs1qG
nig27qi6HJAUB9Pnl63G7ZnwjFmSIP5ymoI5IiPatM917lkzrTB9qWTU5ILM3+ST86kcepnkUwlr
iheXRVboN7lyrWriU1MKYnADPS9FrykAERnUxRydOFgVuaM0mGkNenuzpaOl4I3QymGBN0Xh5K2N
NEvvH1xqAGPAsJeDQNVpFgcOV2Yks+9gmoBzRKConj6QZgo1yblW/Bpaiv2zQBjN/4tRuCMl7yEg
sg64sfUCJZb67ssEA5+sq+BYfcpId/lZ5fvtE647Cl//2ovE2fpR0LmZaoR4qVRmsVYa1+A6+oWw
T3fOzVTZbbJ6XsuUS6+V4CjDhVUXR6z7HNlUa2DXU80hXNsx/ABpzgi5/mv/X9B0HcS1S/DHyElY
A4M9NAVyQYt5YTqNcfDxy/vZg69TuPfg+W7I4g6KboxxEAjx3G5VlYHKWZPk1k2DPv5iEgvVVJzf
SWIoRSTyrMo15m5VjPQQKi4wM1/zS4uff7I93I1qFgTA3QUomGFHMi6o3M8OzV9uXn3Tee9TVtAm
kKPSjSadubFJvtvAahyqjCLKSyaGU5jp+CyYNkR/tfBcrJ3ODVhuyCrXk91ANQ3tzhU2b+V5mg6R
h2GPNfdvHNaFTQNKJg998Um+piCHdtJXZfRmiSgm1IRHqONQXB1Ov5bkIunld/z4t9O6mn8nWz9/
YUdk/QeFdAkTUfp6muZi5oPnZ/nQJDP1ZLW1+/U7bEr76w+yFemUu8ivXXxd9XQ9kSvHPqoWv35T
G77EaFn9rAqez5c8OMRbT8yJMTUVwH4Vk/6ZyzxI+2wB/a3ZA61gPMKx7K8DWpGkBCvvwTz96NE1
xEL8/3I9aSUvzGT/wJqmVG7clTQKrNVyKr0y2ipZ4CmBQlq2rffiJSj1Y3lkzbVgx1t4dJwEFODK
WiLFubqHOHFu3CZSfFd1Q7Y2kbiyqAJzs914BL0221r2ucsVgOxjZLlal3Kzf3OfVcQi+dGzB8+Z
THN4zmaLTtAjStcvnvgvOH+ucB3cb+fOOOG5cD1l7FMOxYW56VhW7Z3SswgAZWBacDLYJzFIlfqp
Sb0jJ4t+8YCKz58bj0j8sBVIEVSw5U7sz13zLDINKcFK9TcwbjFrKPhtXrmNFxGfj5v5oAh7mBVU
CNNxOP4lLrh9az75X8u2AJ8QLk0eNIsN4H+yYaMA4gwOgSUTbW5DzkXcok41BYanyNWDycPPjuQB
C0z9o/O/LRoPf9HOpW15RGJk8YeYETBNmYWjjpE0ipI5xJ4URZ35ON/bJ8CVstMULdDQP7ObAyj8
HOMkO3rCpqUFUiJnsyOBYfGHvdap5Md3ZTocwf5xCc+QH1SHdADrdDBTq9JX2ExM240WvAzo7HCr
IjkO3XZbH4tDh27L+3hZXA0rMxOPVM8VSTsGFSdFrPnsd5+Ra4R8zsHDDsHesGxcQA6eQoz0fPIa
UPs8umWV40GwT4bzP/GJi8FMs89GzFHe9d9B641hOZE9XrGtilT7kJDAYcQWxJbHwuT5KqrGjByE
EK1vd3hLQmIkzdBuq5p8Sdth5giz4SzgaP4D1xjP+A8bEUPCJebB6z/7rdye2w5Lbc5XIUvK36Ba
urWqGpbGJvX9ptPZ4SGyfQA49wfuZmWsFIz0w/SQQmYNFPlFQ6BQfzU4bl08Jj8+JWZqhgVmfd7E
jCQWWovntCISaPsoOri8054rSwBe7tbcW6U1j93kHLsJ46fjElXZDAseR6po2toiyYi1odwo+03u
yr/wxzmWBzrjIfR827KHIxTmaRkxf/PKsoyOY6no7FZ5zoRSQ4sWD0JtxYa+WoIWy7Psfh2LgEMc
K/hBZ8+VRsOKvj/nYJkDnu0qOaxCY+isSYANxUyX/XbC3J6jFX98d1jQPNuVId4W3cxwp/mXeN+L
TKB8Ucjx2dz6nKv+JkdzIJceFZti1CTqD60FsBCJcl8+L1/N2JB1AQFe/R2FhwDZlg3U2KBPVKGU
YAtGd1yvx1kNqmK+pNno9t1PZxFj/us/bhQh1tNc/vOkUmLHe4zkNzGyXSuvPpiWn1dm2g2MU9MC
5HO1xL9Dg24K95Ronwv0v1viBMVJHlGklj1KZOT42X4lsbLPVZJY+UWlej1Kb9rSWlSLLxRkTG6M
2nOjkX9DKD6cjMIpUlSNmtI05IVTlv6Oeo9MwIY5ZekdCoDAktwiFIZSFW0qnp9C/CGnu26kuIPb
u3bUSeBfisO9zJOm1R/v9BRS6xevWgtCswUuD9Q2YECZaIFP9meLycDr9hXqsJ4ttZ1Mvan9CEPC
n9EKnfII+VUDTyx5ioNKuFbUq2i1/gMhDGK9+hZbaBx1tLAWM3jin3O+SH5+KOWQwBH0VSLwBiWG
Km9ejf80TZme8mflNI/fUHCjv3N0mjOdz7TvGOWDmm2BAO2UGtUNCUJR/OOEfqpnVmPbFBgH6x/Y
PhqhrAQNs4I2kbjvwq3NZXphqRy3fUmxJgbmKoVx2DzF5Iu42c/jxMMpEwI49KZD3LC8uXe4L8Fy
vIdxiNgGXStVqNkDGxk8YPadGjvherDIh8o8WATvx00SaUNYxVeX4GBOYNSMts3PyD2ihcY5ftkw
SUwpo4cPd1vtoM/LtrueQlUrliKEGJvhvo8a0jVT3WneTCCgwSMDtxAgvqoZEhOsl+JWouWeRgts
CAxOXhL0PQRj9RZ6JN9TLHC/mcO4AVnHpgNfJ98Swnv8tvu5Exi3AGngbnRuADzx5KjxbWrkrFAF
Qt1Gn/bQgxx/WpKUxNtFTLP3nVg6+b2AbsTaQqSrIwS3q/mxqgxIpr4x4uZKCrz1EbG7rGAchl7S
JeQQy1ddEmuO3tIsx5j5jiuHh+4mufUar6x2BdTOl1yYvPyOIweZ85RKgT9fj2HuFaU/JjnzkI8F
m/ErRX3r6aIxxxsq4zOmQTKcK5Uxar9Hd4frsWn7dvXgiQltT5anFUaS+PWP6xwMYvPHGzilTbMa
u8R8hCBOJXrN52F8v//odKHKuqJW4XmWfzmIuPrK+wSY6nweVRtCunHvKI6ffy/bsMBgKivGg6nr
iuuKQnrH279zBmeUv7POnNvyozLYTwlg4TrOy+OKrQPFk4Q4bm6daxLiQPUReM+ZmLsDJGOULRg+
lwpEduhZGSGf1IwR/lgqHeZHDbjKKmDkS9twnKXiM2AcPkdLzoiwaEzODSe6Twf/NZYaSlu0JNab
KPDMD951RHYASnRY1e8MMv/mFGb5H06Xl93xweC3ZykJerDEElbQ9SUNXEkazZ9b1S6RsjrwBG5m
Y5TniX0kUCmWkfsK37qe6vh6bSvNpuhcYkv4D47U4Rd7uc/KdGiE7UwmkguXt2esNN8tlNaw7Xrm
NO3B5ID+EbOk5G4rmSur1qi7qS8byUJiFgHNmfhPCo5LD6VXBPcIrP7pN9gnxv+9gdZN28uKE7T7
hfXgrD0XCy3Ck0fEqV3ZKr4FehtO/Q4uw8aooJUeR8J63W4tmMKpV5krVxJ/J1GFBdZn6pnLpsaj
GShbi/vFuwwRxY0PUmPlpoPFuu2kQYdbqM2erc4zwAAfCONkcOvFwHPcJzkiyU5qDQf9XLLmgxjX
uCezB7irmfgXrwwSNG2kqnDLfnpf7+wYD0ZjRt5FPRsH3Wv8sRXhb1WhajllSjXPLMBf+iB3TL3I
eyabDw8TUHem1BNnknnozMboNgvIGHX+n8py/QlhEQ2+2EDmbZtRGO8YMXxmC1U2DZW2YbLBHYk4
Ictuo9TXK+Ydfwhn2yL/KP+Im2ANHOgoTMkhc11RcBgyCBJj40Ja1SnWOppcC+GM+tCg7d+7tFo6
SLp+Enis+uvg3mlR7Uw/Pvw2xmgsAAbXmxp3pCc0ZhE93gFRiNZ3PAFeiisw7kG/aUgTMvIVX2w6
y0Ih/k76y1eRIPmnsTfj6QEQSxdnVo42ggtHBSVtrLRz02oEkndlFqr6i++doEl8fHsvl3ichuzN
TmKob2S2Qt6issKR830u0CrMYshKSEaZQOoO2Lc+/KzO9dK43rVR4gVAg8Vt6+VRhEbRO7mWpMnn
qMwFEuml+1RLQuZVkP2SVTzwEo5bnWMs4D1xIqXtz53d1oPah91KaOzjJiZk2CtvWRPTexUBylai
uG0PZMxz5rZiSJkCjBF87XxDYO3Z4JhDpn8NvGwwJgK5hJBoGLtZeggqjWGkhJYMLQXf2K/U4X9a
bC+RKXt8aF2WnnzWSnizRtlf3APelHbFp/9dIkc8lJ0QepZ2Ygp4MNWftChyikUXNiG2e3wqlEu9
k53gG5ouSV+M5L7z7UF0as5LSAmlon62gzSPT1H8U8LnXlRR2VctzCjVR9GNZDmg9P+u3kp8bK2u
aptXyoosUJc47yRr9L7N+H/ccfKdTGHBzn5YZblM76jeigFbyHTmIk/h/l9i7d0CFxMwXeGidsiv
FSePuTgcQ/FrhToRbG9wbwgcu6ql1fqLt0/NnNVhARC7wSSGSVJLuQ4FNcBdy/OKFlxCGlJQ/LI/
l9hh9fv0gnCYx4c8UIDfrHHfNgJ1yjzixSe43oGqYH4m8rkfkW9XLTlDe/op4Qq+zVlANa/xhn7b
VRcJMYvdRC6ndZai+8r5HeWJK/UKqfhbJG5WO+TT+f1gYnUl7Uc7nNs5+cXKy98UPfzL54wLdUH4
miA9lz7sJ2w81N7kqnt2SYgalT1mZYnVq7wN/zrLdgMuKbNGShpZj0lwxGxFJ7HL+bLx+KsYvNX4
uPtkCnJmm+1b4R4sU17LteFIMfsH1h2XZSFaFC4t/WR2cndXrniTsUbhaunFE4/MzBbpGwtVhWUQ
iLeMJ0gWmDlB54+zKbk3UgwN05bHeEHbg/Dvc3isBbxhVERiSBee51pCbPlnegvIb7dvJoYiXL64
IblkKdTBrhfd0KuorZk+ThF0JdDryp62r9zHEfwSFf8vXdaW/KtPnH+EVXH1corXe3FaL/4Cuy3f
VKMzRrvq9ey4i8OnkDZ4kAb4aUwQaUAaYiF/fnSNZ6ySIpB/BA+NXV1HCSqhbay4o+RVLCawvX7k
OUJfLoV51laiPVvXcZMP/ejNLmyCezsLv23wgP5hsGDidZP3RPPmEN1VSa4Q1NJCvL7IqxZyMwcB
NJ+uJmVt8PDuK1uaFl5DjirhcUpJWbm/CI4Phs8DZjOB5yohkIM1nBmmcBvV3cSt3eGy134xp2Qb
/04by7Cm+3jl9AqaUVH/Z1yppvarw16UKb2Y5qtXiHaPyU23KGoclIV7jd0c7cOMWsJEccEJgvDb
/kbv44c0jjrD7gUyJK7mA1esP5uxNXP2JfY960hdHRD/NyR4g1DznIy2pHRvjrI0Pn9+SRX1fj0/
1cGpNbqq19p8t+pe8myUC8jbRXVyewrgDdlcwcnk4us8VQpqt0nNkif3hd1u602KSpzsZ5QbLNo+
YO4iVrfhV9CMdbNqD1h9H3dZO6kjtzrWY5lrsQQY+n2VyPBlyFBXgDRbefOz8QoQimRTKNE0PAlQ
J0XQu6LzuQp1LJ3HkxEkk8hVv4DNFcww/11iycVTqyI2gm6JdL2gObtmOiFyG4llAiPGHyHUz22H
SXd3pzJXgahgdVmapHWzOtP8fXLmHH3sLwCz9hD33sSu4zHhdBQoU4UxWf2ZX+UIBxbXy/LFx1g6
ZUXFQ0HY/xL0pOwk4D4fYs7z/YAZcS7XhIeq+jAAuXphH8qtv3ut2E2YWWVLBuYjOu7V0h6udsIS
lbv1Iu019t47Mz69U1t3cgjYzYbSDs/k1uenPaAmRsTfx2qZQ1AIAICxms8fNYTU//aeqL8cR4P0
2lBsqvZkEnBsGCgUaN5KTyNOdhJYxuT54oGSU+3I5cm45weeolHiMM9Rf5GwuR++4P6DJST+U7ay
9Jkb1fZfWyi9cItrAokZ9sgGLFC9iFVJA77HyZ/o0sNYQ7wU9TY+35cCzUh4EefuHus32ap0GEHc
7XIO4NUL6sT3TJmiKMfT1zroXSKu0TkhcUzlE5H4Oj/nMCz6lDkclwWH7vlS0xP8vvJpR8TtJkNf
iFxr2Oz0c2f3C+0EZUK81qKwP46xOo8Jk7iTy9f7fj3IDhTwOcceASq3l88eRtBRP8xgjfC1m5OC
e3knz/57FQRDKWqaU43SDDVTU5ydAdsXWgQwro/5cseoT+kR4yNGo++LcBsHA5rzvlLGodNN5doQ
kNzzmnRoIDxPd3gfKM3x2cqcikFSizPasS7MyZbqw8bbBptTDrlFrXkvhh9xb9yqESKYMex9iiM/
Fd2uz6UeWPQHkR6dNuqYJ/+KQOVFcVThnG9Wjlpf3BV2kkk5bb5z073c+2Ec0KuGo0En4joayaYB
rApHbR+GfjH7Iv4hBjutQkJLnF0VDcL8jye5pU121SW1MKgW5+Yi6ppT/yhP6trxfB4IkIb11eik
WXNlhAbkitftkedK8vsm6flgVapjG2Nt1R3XpRjFpdWFa0EfAi7qm0Rp34WzuR+qN/J0oR5sYH/z
n3AfwiuPmhc0BzcnZ1SA0FuWwnx91VvJXTiCqi2cBjyd04F6vrAhdBGT4XWkjtPXnl+UFK52YOoQ
jgweQxZ6PnFUz0wpI4UqS/dpNiVw07dIevpLSds4b1oeGsrUD50pnZfsy1gUGpB49OlxD6wb6vXL
MxjPni0x6rDSnOZpXYgxgN7+gykCaXlRLNWywiQY1YcI+Qv7ojXoY2gXyPsbSac6XocCFB595Y3F
i5a0/XI8xkmX9F3McHewqy1XmdbAQotp6kkUrkYr9BjZQp/e9xWlF/da9qVZ/jGYJzNhmof7nAWe
l5PhZ7QWxT0XCA9r3fvRZXBO8i4sT+e1UIBgxAdYdNhxDf8/V/QXx4R4XDPpSIdeXEIIn5CfaOfQ
DxwHkrv9YNxF82qQYbzfOihOXn2t0mD5gnA1gRTtFthWdAnD+hl0vpVn9+IHZDSJCJtXqgilvpJP
MlVuMRLjqGpoZy/dDYouWV5/RBivzhO/9ZN5XrwqpEQU/DrCsqvSNSlyQ34kMcREqlF1cVR4xHKK
I/TRboyFtKtz+O9nmTzQRWdLjpDzep5Z8G+nz6oWeuExmfFEUtrkpq2XQXxYXFfHX6T0ve4GMreJ
m0AXN3FcEqcSTXqBy+NW+A9u7B5PVADL8LjAraWAizqp/bKTS5rnHA6cJURcA1khqTfaIRmOIBAz
TBqgb8tLZ4CFP45PskeasrQJ1PWPza/CCCoTaGxv0UfKQVt9mQH6ASxBNbFUPHqRmVjpzNIc7ySw
PT/qkzoUJIUiLOqpX2Yo9ug/k6/x6Vf7tuvc48+lKDVY5XRETLmFgnd5XKuz/XEIkjyM7vW7lDJ3
81Oz/pAuWxzFJiSoPTYogKdqubteOl/JBAnAFB1LpsaAlijEXCny03izZXrk3zqkjhs69q2vi2kE
dlOJyMV/jzeplZULk4CKLmwWXjHHY5Rf4AZ0/k3STee5FwScEGgAI+9YU1xbPa3/V7Tq/Sy/mK3I
pFo5NJ1rDUUYPBBqwBDzw8d5x+2TawHNeCPPUhxHbl7oMR6CS9dmdFgyd/JacL3B/cPun2yR9Upn
7C8NFFO08r/izYa0OXwvVB2aBqtMIQTxnEUNgkkk2+rsbhMh+UJ5X1t9CCWbUgWqqnG9QRc0jHnx
OQdU0F8Pr8v/jybKMoGH/OsYa+tfu4nq/cVQFM/E6X5tvfXvDPFVFOSszGjg9o/p0P87hFcXHet9
CZNEotM2gJuTeyIFN0QVvC572c0mGBGZ+z9FCUNWsEQxfraevbQ+2vgjaUtBvmHOGkYnOZpiQrsi
TeIOHTLpYNW7HtBWx1m6BVKFl91Ae96QJb4/WP2CVsfvnd8MihWu/Fp9RtJiSV9y1VaftIx6wVJd
7Jvt/sfe2EDi2dd0R9rd1FjjDIWOrjx6kwninWB2vD7bDQcu5JWgzh7gtemfSPjGkYb5rTHV60jO
VffZ83P0JkUfEOlU5q2WMLWiUM6cnGpSQcI16HSQm2GsNtKqNuIiZfXpxVNadyNlQe0Cn9uNXJFJ
7KTdLGWe4oiHWU/BYAi17Mc72Sb9KIQcx+s8Vk2drF95dw1uAcxUaouuHubHBkzuAnX+DTpry7T1
asIansvjRdF0JsXbVwV6WEw9vOlYYT9Z/E5ZWtMaCl9nAmp0p3hCWR6ypB9tLhh8t9tjZ/ctHSah
0eW4erLpjIQiil8dG0jDJEQAqziFpfFrvuA2kq8FQ9DIlEYgkp10g988TOVebXx8KMNmZ03Uklnm
Dj4BWvm6bsHrn3hHLHzfGFrqkNXIleU7K9toAvl5yMHQX/QhFs6qi/KsRswY0gFHhSFSrZNQ7QPI
p/clZ4lJUvBM1DmYNFbmot7yII3X5ov4gJyCAyepyk36FyEhxD1ujMVUfONVxhGGUzP6GjwTq4u7
XqvicjeKy05qcX5DmAZHcl0+eIeVhru4zOmBXyuoBMRTuyHmxEZnRrcIo3G4n4K0KSByWaBja6Lb
aWpdX4GLBs+E+9o7iVDHZ8imbFQ5CoQID8+ghUAzgRxq5U4GztngsYb5dH8qmj/ZqwYrTSxXLpMU
eNqTF46xjQYlKb84E3eiuLGZ63Zjl06WeTPRAWfBkBT7suXUoM/kxUz7APvXnHFn+Z7EJ9Q6DXSB
kzhFqYcUzaWLf/JYaJM47vAKFMdiew3QHgI2QVHIuHJKGUMeXU0q3w+b4OurSF3Nj7TSuztTu21N
R44yhMRFIB0ibxuqmXb9XpIbkqJsLXDiQKmV5iCNqB9ozyW8DNERCsdjLzDesSpPPRpRlGy6y6Rp
chhWTgawFUckTgMQiG4zU7jrGdYzBDegCzPP94etnlU1ScpK4LK/qzn+/myPbg1p0JnVMuu0idmW
jqdHxVwRf+hRUJ6EA9TVrC/T5kkdhF/7UM6Pwpt090Zvfq/XdlsX7hTZmoDUZrn4O5LHn9U5g93p
UohS4DXuNdntffoBzG4Dm+MUI2u4YeMfQyntnmxkjY323AsEwZbf3yEV1SB9j7qLPpDug3OtLuyN
3xSXAsBLFDPn6ebGk0GYZjrjZ6ZLc3xGbYZjViLKyObK2pc61vBIjE/G47NMXRIwd/FI2KiePQon
POleU9DDIlpJcqF4U0pQ7v0lPZwlM4wzezR9uGQXr7yMhTIUbRohjdW9d7Yg6U5P3nNuYk0pcJVS
jxsvcvNvsupp2WV593JycLeyI9G28m9Nunk4scG8LftgRSDmVhzGwH600QcUV9Fs4QIjuDc2BSk2
g4OiHTqvAIsTDgjXGl0C6bBiYSUpEZdk4gGinUHuQFqebiSEfgDPtD7tP/kOyKupvLo5MEYlGhbG
kqMM4B9CaDvDx3AmfzZNoLMHy6Nd3UjHvxQsRtl5gP+JSj+UvcL6SY7pT+8m6ZpEr2rbrAMbJCE9
O2bX7fkG0M+HXcUkl9NmU5vcuAxPVptPNcHv39M5XVZnkYOCnxg4LwdqPkvnBKevWrm7Z1FP4i/r
OkK7fAePLLpHsYZkEII1Vw0KdL1Ew0dz8QApLxiHp539haOqL1jjmv68falMstWyyavux5+np0gj
GY/3bLzzW5Tt4b2PRyD7ycGE+VVw2qhGsjULhXBa3FNSnt/bTLHqjC7oP29zqq2Ughxt6HgZbzNK
Quwg4FqOLeOsZ9MTedGV8HamfJ9fr0rYSyMCUGrbkYZYaO08NW/n4wTOyLAetvgtjocq/K6PfzpX
fzJSJ/Z5VK4KgSBBnrsCkEVUgQJrVXOEwibiIv9tEwwohP90jLKYZjnD2vnHuJ5ms6nwZlqjzlDS
HnaCjO7iyHY0zJ3eZIoZIMecXpaEIipBheFoYKYO2DyIOLFKrunAbZ4Y9llNmhi5S1kWR2KXIMG6
PwoUnXNY6K6APIa+qdeKU7opAXXifLREnV2XrIbFViPmOb0ESHgiiUBqDkMDunJhngRKcnXvvrzH
0gim9nwgX4OSYXXNk/QOV3tuFryc8l2NF6gt3ByRCM5ORWET9cvfWdHzI3Q0F4oL1tBHtFcXsrQU
8PQ+KHCBsndlcsS6Wum45K9e1Qt9GYA22avtvH4MwsYRendEhNHHH5HtpxDaKjmlFNPakotKn1wb
LRut61ECmwGcKMc4ALnnkSrvRLlBDgFAdHiIejE7aiRUIympEsp8AY5bF7asqLg2AJzGkYE5W23L
IvZeh/uigUalBEoNzBOHVTLPPLkAx9pbi/XfJaV6iPH3zyznl1s6iS0NDhLQPbfXatU4zBm2MR3O
siDIcNce73NDDVJ9qNd9U6WGfaZYhtQBUPAAeupjDYSP4KjTd+fazZhgaywp26QcZK0cXsr8iwLD
fhzBOKUlQriuY59ll8ws1BTalh6aE8+RswGCmVdIZxJuUimz5BBVaG6WawBmdrTrmYT3n2xvnnsT
mWomJtaKowdCWY7Z+3YsDKiT01L67JxqJaTyKlBzeSuPUzLPAPVuOiP5hrisjverzPjBG51o7v86
PFEpPd79WNBpXqKI2jaRiLwdasRTa9Wq3krEpedcc6+sK+seic771HDjaPj+/+aCVuKf7e+1NUvl
Yg/iXyUSl+ld0ezYQscDXuZsjmNryisq67FzQGehx2JMUywmo0mw6H/YLM4N54BOfhgugWOi9Ff1
wnkc16G+BgJ72FifmAGYDKJUFeCKSM7wEqUzU7UFgKB+v0IBb60UBYtduLrLrRys3jDiPsoWNs3L
gbgfzjn/YKFbd6UsmFW2CJCEDhKEmvQTGjuzWxseu0NGv+IiG0Sf4IPAO5bDcT9AqTAFDgY3B1Cz
IzufZhNhviDpKXwtywZrnMTkRIaZ1xXg1Bmo8QAsPt7q9kGGCjd1mIajL5J7g1etqgsDSeRd5xBZ
cH3rUmey+fmHgQCsznrhiTzCzijvAI93cHJ+X7Nw7/TreB+D3+fFcZXsSiR0G4mWaF9jN0ZXyo7R
nBy9adrIKxt6I/B1tyWVHJoYYAT+blC8wYaYKDQU7VrnQ1LxuIW05QcDTID6K4ec2520ZdT+KB9Z
9gbnoq3m7PSaCHzAu/n8Ch6buc5d7iAW+NNcq2WNNtK+W8rwryjF/PdL8n/WIuKwVKG98NWdbMja
SFT3Fp3J0iJRyzAFLVyg5S7RsWDsOJitO5IF/VTp8+ISawU/2mvjqTAYOx5UjlB6+pgIfVkKdZBw
h/umtg2YK+bi3b0m6oJPg87j6gTN9URJKJtmv/V9tuk3g9J9qgqNaqjwHUoQo4zqSkzHA5wKbIRM
cpkfSzdOXS6w/D+s/F2p/nJeJsfFAJVLt3QQe/UfZlNuy9lq65G7+Y2QPj+BM3pZm9+A3Mu8Km08
YrzyrWcVSh5rVfVMTuGtIuM8iV5XOu75arc9Gdy4CMTCk7MeLjft3yYr19UPW9o4bz69n4wAnUki
MFJBr/jOw/OM4bJ1TkBD4RCdPFG4IEH4QBKUcUSesvhvvfBsDDUIKlOaaBAKexfrriJB7wxSw3Gq
CuQqjozS0l3nW84hPJVEG24+/KvH+Ms9lfIGTSk1eL0ipHESUcocFJBenn8rgJDXUpxfnIssr6Y7
6JO+a68B4izD2lcqaIv+KXgOEjdNUzPX+qbBfESH6VM361jUZV/xtQrASHYWGxrPImBqiQDP+KuZ
QF0n0YvuNvwbOUxVAcWxQECq1fTm3+1vucbQZZFC8AiKIPwSIOR3DJv5knwE789pSnGxTsJDuAUy
dDXkrPA+tiivPInWoTfOSkcFGdKGOhna+Z2De95NheHTKqExXZ4C/1PJSWZA1ZHD4zAMsVgAQaRB
6o3bsTg6XozycKRbJY5hJ7D5Rs16f92OImYgNjKuzUMLc+X6qwcFr8RstbGnY08kklSgC4eDydbE
VyfC1HgrGtIwTlIoaUgfGM/+4N3et/l4ZWcmoQKHylr8uZeHCkJ4ZHOhgQWuEb2AJU+ItBygViMx
DMVYvj/kL59a/S27QWAyfZTgpbOA3Isefa/0tjICLS43DPXkRNtLi8ernYBJgSbTnBC6kyt6AUQk
+oOE1BUIFfpBV/f+WiSOkgCyqzAzm7+ZdXsoB8HiI2glDE8TVS2tAb04H4i+9EzxmzbV8ls/EjHW
vkfvFkdjIWHg9jWUFmYWtgOdhZ28jCDA74U8Qije2KBWu91AuVAyoqWEqRhl5huMWvJ6+mZ2sAVm
dCpdt9toGZX5QSSes8+opUMK6/sCNqjYXq6d2tccPBJB1ME3+1Ofh7wJ7tUIeOwyzXAjcDMQKdui
p9vf63UDdbdCRMuCoMWXrIxx178+HocbpH8XR+UaI9SxveX+/a0faegGFMqwN8kUKImK/zlYg7og
UQdd2thqm9uby5h+UoB1axUFDRaxH2EPoZ/oUFTfP43sg7slTbfE+eF00P10NhiWtHXNXOXAIPx7
t9agiW65sNNUD+yipyeRyRuyZFAID3cWVN/fc9scB+oTH2UDcz8UdrSqZKxD3ZejDCkyWZ1GR1qM
53c8XkTYV8+ntmuk1dqV7beCXHVTnSW8CFXZnmgm2XaOicW4/7nFwLHLftbD1BSxOGr1okYzb55N
NdFPN5CHQO+BKAF6iKTbeRef9APPA1cfjsAOzeShpCz/7NPwEBDAbP3ADgYJbpM6wwiAvUff4Nno
PNDHy4n4N6qE9UKDsdjPkbfmf4+euAVBdokWGiyxvo3cpyw1glqTaBatkjbr6SdAbLMgDkbEDL/r
jSkKTLj/rTe78sjz7neq/iC90DFlZK1Ia1ulLvKm4RSJSFvjyT5PLMizxQVMFfwzBVSkoznv2PiA
hPdEQzmLkXeOscPu7KF6KjY3fPzVO4nuQkYrbGhU+I0/Qmt7fTl0ezWvqOR7TqoCzegOzHxv5xV6
koWZ231SsczUdxXZdbCHGSiKnI5OHwtG8cUSuu9XwlUYCK/a1zSG32JS91HmvFOWXWMhuDpXX0uL
FzfYaZBRckC0XP2ilS2xBfs+TL0G9/vFAaWlYDUV9xyt3g6MHqD2pXOz8ymhK5mvuOIFDXpCPuzG
FKMr4GHXmwauDtpUOlsETdFuozQSHzPl8LG7w8Bo4pf4isfotuBhVo+R+qyHKvFb+9b6oumQsAYW
f5zgrDMujqGL9/czIfVt1oDDduvkA180/UYeG2hsK1GmIuAAtN/kyN65iporzFatsHzqUyNMBbta
3nyhuvLoJoI7axZAYW9vQYSvXyKhGTYw8jS3vU0mTwFg3vfIpM6RRhtPAIFHkRwqoe7wKCNpBtN4
9YxEikWFvrdqDcvY4b1Map+th2osf174Ry3/N6VJ3TnDm5dIb2YMjf5swV1Qtergg/LuIqPso8zY
Sbbw+B90I0mnVFKqMsvdIOnz1v45u9MFzV29Jn9rTatXRJNZyXND4AtP+P9bERnYDPhhMZXVipTU
v1zfrjBt6Cy9W+SO4/sS+b7iow18Mr4t8/yVErhQW2o6y8irf3k9lmDHpO5Jkr3QDU9ZzXPb4TCL
SL0gK4ZGfuu6iSVVkgcBHeWzMC4dtv/YztCF+kavnVuvRTTh5KQ7RyFwucYwKMPzOU9fErD4UN7D
471OLTnxzKN+Yi+GYaPY3CNl60125GKCiXUia5mMGiX5noYeZaLwq6RDROS4HqYtG5tXfvDNbHdx
ohLo/g/ikM9uI4SK4qSAOk3Pg3GQi/0qcvxzJSQAbH7DKmdhlR5fek2CfMGsC/M9WiFGwIjGw+Ao
Lxc9wUcrAqYav8x0eArvChXYoKGhl6j3sUPwTye1cTRMSy2Its+TBJG1S5tIvF+dG0Np6t8XpUzh
X0QZAgUOcffYyhLZ1q8JMDluI06tM3JV0F+lIuwMBB/GuC39KKk8Jhm98fp4/UvCfoqwOEHR9XfF
57MOARhTCdsMPcx9BvAL7/AKYPxsqO67frczG5GOQpJ2kfsetk0bK5UgNFmqIsYP5WYHgF0o/MZl
wop/staQUyllIPfljXIROLvOdL6TP155vAON9G/Q7Guw5sSMZVq7x8JZJzjdw2xxqyTwDAWyOsRt
ZapMC7n3phXOzagXVS4WDFv+X93t6pgmlDFsmHNF4RCJaTcoFJc7wd9TfAM24fcmYO4ev3EW54gY
gx8jHrWvZelGVV3rJf1iaKdoaVflc3An7pYQlUHQLtUOeyDH4DYGq5dZpKanLfORFeadiicbSqIA
F/x0eOrTKI6Kfu37jXdPVJ8XHdBXJmJCYn7g5d190xwt64CJPnIxtnWig9bU39QgoyoFUeCau5vd
GfC0X0Ow2JoUzO9KWB8yWfl6x/SxU7J5HLH00qs/orrMN9hVy51UHEUDO8Gh8uf7mVpzDTFOHkRC
1gOlLD098hF3XToH5iZRLRoVFp+dVxugNukZ3oMwtR+X/XhjCI7nqvRYk/PLq254xeHC1wiM24lO
OSJJ3LriECjbm17nXMDgBf5yZ1Tu1NVto06Nu8BkoQoTiU4Avxir9tWl5hbmyStvpUy8XppwprVF
x0vb5FGqlkS32UstVO6oxAtQCy/TaOo2DCmTOhXl9aMpxgCTHAaSo2+Fo38RAe7N5A+RzWhaYkyJ
qicrYAhIb4QzBjOPrVg54sZ8lXjhnkv3QgrBcd7nLuCy7oUPzwjtnT1H3tSeZnlTG+R7TV+s3Pr5
bUpmj4s9FN50GJNCgnnqwI55uezcIxcl9fCX8C00Z566MtHJVElQyiZOYMIwxcPren4XGMseb7+P
6kjku+25ZIfPUrncyxFbVTVogo3tedDxWwK9WqTE6NymUUeXamWUx/g7czALDafh9Y+roF7IWRfa
lPM5wNeWzc+Ag3trf9nmNuNkrLWSpcy8TCkHsNxmp4XtQ+uof7nKYxxrc0DMyPhlCgTnYsyGftHU
ISZio0+07ZuWNYmtOIJR5q2GTUby1rHb0zVnVASz/ahHsO4AjcKDPc5JPm/3MIRwQmyP1Bo9PL4J
m5WSAffxo+9Qz+y0KBBc4FITpko4lcR4XgRkf7H0DF0VpsIciRCttROcEKkZD/zTCVn2078Pre+5
Vsg0WSP4Bz1ARsAFgRy2g31ZrxX6x+VeZreCHgVns47UXa3H6R267oy5TUVYc1liNqtA1pcApX1g
uppN1VaeF31hhJ3q5RfkB9lTI/atGcCjq9LhjqR5pSiEOCVB3lKeaey+v/VlQAoB1gzU+gugmOBO
bHVK+qgpSJR/DN3eI2jDrX7Adh6FBu2ffsF7RVo0QeuRLm1Noc1vszhv1po4JPfbuUbQ59dQsr1D
a0jBziL8+fr9ipHU5LhOdB/VY2qU/A+LR0HfggqoHJxGOvCk4+CSXuoX6ewdV+fue9pGc7HI6IaM
2fn37oj8wEJKzdxABtsNOLeHIneusZbHdtaidFJLSqGB0FWYCfb+QdWE9ToYSY8uDgQOgCBTcEM/
1vpj4Wkxnon4cAbwPDZjQ7UkAvuYjcqkBv1k0BnG0zn3sZne5nHzb7GaIbPeHJzhUX6AX8kIUa+V
rfNdRToY7lNxkGgrVFCONl+ryY9CrLgjhaRfipxVsezf8imwNVmyt1gTzReFPtIE35BlDer3Kize
4y6FmJOLhDiUJsLb1RwOh/gFyLiiQvYSysY93X/ixWPrvCPIox13JUbUP4u6XARAWqs7KJS329Av
rdk314h4oJDg6M/RqH16G2PepY6BiLI9yygXS+wSQcyz18kpR2Aoa8sQt4SOWqb+8F709MfxvfLn
kaDgxJVJ+bR9/XLtfMkcU/yn9tyO+5fuVZlK/0Gz4wEc+AMnebiJiegbFLdl0/7sDpfn5DJT3pOq
eRJ4pI8e9klcBV8siA9wgoDTytR/gMkpUUlbM1Oi23qsp7tORRVJREPDLMQrkrUoTyj95pqEzyfw
LE06RniQypSYmpVC0O9Sfi0ZQfFJluWoZxPW78a5gLQ8xpXX7b1y0nHv4kQMZhIRc5SoeMCDUc8p
VcTKJc+fFYp9Rbp2AQm83CamZpSIGfzNDt4uZnXhWW3u2AGybOfwXkJSY3vNzhMG1uVwZlwGGGTA
FfnnVBFfEqI7b2/nJG4yyCE1JeC+fRYPK0G8U2PkSJ7uw3RB3oKU8l+qvMVxCtANg60gUQ/TFceM
ORAeMLT0HPL6Escd7Y8R4piQkktJVgFmKZRO2FuF9BVwSUZXHjukLX3kuDCQ2pwP7VG12/OqiJ0+
FDaMFcM6xNScXM4lVnKKZ6lJZn7pHrurJtMCrWgSNAz7DfbhU39lPC+jm21RyuaOFjz/NB/CLqkn
R/WDA6qHGzxOaeAzpmXLCZnb8gVjJBZq3BUYS6OafMDlTxNEseZ9/5BD64oh5mjawXni2ZQ82m6F
XM3Sd6+I4XtEPbv8xc9Rt8FRrgTZ1496XTKmQbRucpcCHnuRjsmDVt1YX+x5JX1vkqAc4xwT/huh
v+U9PYw+rk7v7v0vD+/QhwD+6kiVgccj/IMv0Cxfm62QB31pdDhU47xe7sI/xT5Q43x/r6D+Yli0
NSzqXI+paWhYrn/s0uJKHmk+SjkUb5ysj3QbNLsDTccPxEY2z6/JWivlZxS0tTrZuTLkAuOo4aXj
4TIuzUuMb6V3YibOjKZn3egICbkRElzod771Dgy0q/VZ8oDM7zmz/SFJg7diDCjwu7BD4UZ7umAq
netOOQ2rVzZQ+fqHs0D/0TgkGTEjqi8iXaVtiDI9oQFGNvhcSfbr12fTj1LUCrvsaNbzHQjbQcw+
yvyDtdpyiNF2gFca+7xRB4OapbZc0RubGL34bCsYDfOepdScNEw6R5u/uN+LvHuUy9Ujgu9sWZX6
vSOqixr20hrxu4OX/cT6M8XF9GJCREDdrEY7s4enHRq9BNR9vz+vByRvf3+lrqtZtav1oK2ulocr
7PHkgOKy78YUon5Q7zzsJ3CPhjlO9BmR74xIiiWOgykQ7cRqWUbGoFFt6Kay2kUhcanmPyGTO1dR
1s8VDo4KNw9Rm6gVeoiW5w+x5v/lG2NwsAI4EXqx+4Jpe4yPyjvKGRGMRwcxdKd3rdrUJGYvBNoW
fbW9u3+pcKD/pTCzMiaF+2+EcNuKVZBO3aARzQHOVpg1Bsgp4W5VTOHbY31XkRgWt2eioo5rEo7c
8zSpxsijW8nFgiuSaPiFV6w6xuyrWTQusz1JQMh2UEmN3cm5bJ3o/RWo98M/eioglzXSCkIw4T93
cQcRN3zWfxTo9gPk5KVMPUlKv9ieJj958sQ0JzEB5B+g6ZmNS3WlPFB6Rzv2mG6NYXCLPF/NXlo/
YrlpG2TAAJyzZd2egY0pVlEtrzzguTw+03+1A/dMV7DuwKvBa1A/qU/7fwEN7sIuXRkusANt28ux
eGxpMyHPYTTZ4wPGATO0II1PYrh8OKDGa3sE77sbhwPORcTvz/a04yVibhcL+dpjzAmaTJS27uI9
MF5O2nGi1X55z58BYtpuBK4jG7wxElu03lfHLgnJFI/7clCLwNn5jCT2n8ih9kR51szgUvglHLD1
IsIn0nsNdDxyF/oHjuQlhXIu4t2BVJ4z8mYxNnJ4TWNbRntZBBz6biZC39ihEPPAbEUejv5X5UMb
M94Rs7qEL/Rin32k4+x3QqTVObcQIw6lR1XiZIOZPjfn9RApkWWMAFFZ93M0ZzqgYvHQBNw8AK8Q
nV+wJAlQJ5eW9zMJb7IBdpTuCXK55+8rSt6vjTq3Cq/ukl8MKM0WXCgMuKQN0Csn5zeIPVufp249
GbHBGDiCtZwbaETHCd5T67+EhYWGKdszVq8c/sevhvaB8p+WuAq6z9MzlzIyFWol84olcNnDRWnR
TsA4lgvd5nkn3owCnvSIbuNSDpxiTNHu6M18cc5PXlkQUYOE1YqN48l7ycNUc6A1+bIlRZNOh0xU
6y8fkrUlzfajs6nuPEdEBNNHCpoUQlvpfsB0Y83JSB6dPzDp+6t1tQda9cg6bvHKRGV5MPAhNI++
Flg0fcKFCrc9WoBKnCEJEtE0/KpmIe3fGZr7OLYV4RHbxx/1Mw1WdWwfbKIp0YOe/8k/Vf4iD9eP
R4dFPLf02bwk3V1cGm42KO/j0AnKB/Dp+a8T11YM9fEu7hk1eUM48o8Z4jKYoojIaiqPxjoAjZYW
sn0eJS49ls4HdM0nkVkLcBMlQMOfCzjqnMfvuwqVWRA1OkOc0QXwQYDdzHjshbqu+wK8mgT1wKYZ
DUprTlihPHLQhlfzbCLO533QDJy2IOeGabRz2ppQegribdBFr3QoRTgkYBN2MNgG1hivQP8+f94i
Ia/kZWw1GW50KBM9L101klBFw/XMFsJ/Ex3hdGgW6FrbDalJfDoNYKn55RwCws8seNMV/2O82Dzk
e3o3gOZhcDob9KUq6aiBjpuO3nttyZsT/5r4JyjTfEqRoplXi2R5RkI2fXAlSiILOl2ndH1jC9C2
m2LgCWC5ZrZge8QcXlF3LZ5eeoPKOzyShYUY7aScNYxILJpAxss/N0Z4EcFxRVFqJOq6uEjbNhoA
ChrJpwVDupcC/S456e+aPJJk2ZQq/H5jh5CRj6CMpWKmKmqyhHDRsOlJlQh93q+xQC3bjNJ21lPd
f48C6rzpmFiIWCbhbC3LbnHMsUjWI0c3ZVGQyhwb5oq/+AJmzSA2s0sO8VZhdv6JaSaFG+Zv49ES
J+pWeBIOKH1+wLSciH3U8lMC51+e5CvxyKmMKWWdw7SJED0K4A4wLtJvz4E/wDJsB5jM/J8zc5EY
8QoU6wzCOel85dplBR0RB8H/2roVU0HJYPMz1ZUP0gk9YZnGwKhUlcMGkfWUgaNKlSCw+0qt3Vjt
u5azmmogjyVcBdQMfYWNZujoAwGjgEGk8eSCKkGlIdsNRxfSu1SzP3N+A6ZY89YFj+taNirq0N8E
cGklfd2Iu7P2EZQl6lzhiZYEHjtEwuaBXpz7ewfv3xsh84iRSWoMF9uUm1sJ+UjJjC7f5W+uDYVV
5eseGwVP6jtZpdRNhBNIPxmcNG3eonNJC0kB1bb6ZRJygKut3MVKDlhE6wzVM4ipXUPPs2+lyzTJ
hTANVzO0n5bbwI38cG8B3ZK16PqgNnH8Vzwvgj+IC+upNuOfK43mQflMWao1IKsYNYUKCwfmOYEp
3YT6+GGE1Eip/80gP/hKDQ6WpqPjKRFGz4nv6Bn4Vw9ZLYu0kx1hskIeZFxUxdJdyn4xvvj+fW3r
qBvC9TQkKaUbdmy8sWBs0xH7AG0hKSPdd2/z4bPXpICDeseV2hXHCjeZLwW9IZtXyDSiyS2yyvcX
L51WQiDRmhFzJ0ZVksnyfhWadJz5IcTOv7kfvZx2++OLrj2aNl8DmTuUSdbUkjvg16Cb0zcqAVeK
RBAwLjU8feAtMsiYHS8RYslX/Cnlj72gHXdKWAGhZiulvFyTT6IxqKEtqGYmjTH8zv8VLBd75OMd
6aCTurL7rsIwUYzleQD8SvL+ZTK1YKGdH9BYqtrpaBSTicIFLOb4UGYv7BJO4Ec1oF25MOkoByAP
BACtfcCtoDemXC2Cx2SawI44WE1sgNGtOQgV6ASwtJrlZ2T+aC6EWmEXFIOu/THXNFv1G+RU/Yt7
DpY1/CwapP9uHPfFARSds8nEH4++7uMep2+7N2q0hYZPACstAtpGRDsTfqOprSQNpnZmCVB19V13
ige9+7mT+nq7dyY3TIJjFj99pieQu2qrkhb+uODtiEgFtO/mmAc8is9q6RRbXu3z5yIm4eeoe9FA
CS+mTj9FdnR6QaMQN/RrtPcAsy6guNcPFB1PdrWHOncv/QEZB7TEompH0jn2Qy4GS8OZ8V3CujMa
tLc5DMtAu787gfP84qisNFwEqSyqyqiNZGvFLwUap6auOZJ66/lpMvDPw4fWgu894YBCB3Vl8+pW
U/goUEPxl4aYjEtov3mpoYtcxyhh+2iaYObugt7mXEYpSKswQDZPrwXjy2t4iW15mV6R9NV70DAY
oB2iib3jWv/SOqr0mv26OVLmSdrxIOnvXIEXMLzuM5cmh9enDJcu7oTtzJNr4j1jYCkaBIMFszX6
2aTNkdPERQ8BEmo23/HmYU8/5ciLVzi3zubmRddtB3DRSlcdj4kWBqlGT8jU8z0tCl1E42fdyHCX
fN8x+ng0aVEeAU9en1xkr6apDpijSg54jFROMu5lm7CvCYiJlGAB3us5MIMLstppVBDqdey8AfeN
JFYNQpEvFtiIn7GK1Ewb7c4I12yEVRgiME9k250rNkpKkxkxXUYC+QvKInhMLAUQ/SKeV5Ux6Ze8
iroEJLCzx9YYDNUVoThE3+kX2h/BAKXPAkiCwErfzzqOjYX2ShnEVFFbsPSjxRd0+Has1VZxJOyu
Rmpu+byh819Q1p0CgQV+wcjdnI3YsFa6nSaQCpqFOq4FnqXBVnSjymx+gFmm35gpZLXgXjjspHQq
I9G/je4ddQCDSg8817mKdwtMTv9tOJyobfDS4+A6mLaSt+MVFbvFtIIMF7+s0HihKmknUp8Sj58A
36EH9Te0W6tU+09CK/nV7duSX3oLyjhHz0SWDHx+Z7sdfJ5utmlO8gloisVd4yYRDLn0cKg8G3aH
ruIPzrwhX9wRDtxzrY3UxB0jU3B6K7s91rh3iSdos+vGHa8qNCptZowp6PL0A/V9Gpstc4Egk/WO
gR1wEQG+1HfsDlD2Q+XNb8w68uorpVPjLWEqFpdlVtt16dEk8mO+dwpELURb8VTNlKXPLG6b0SJy
C1LgSgACDnpzxoEi6PBi3HxGRQYpEhdzMldaC9HL1mhGluKW89HVPo2uBWgT8HSBKNzl1q146/ZZ
Fp8E4GUXRaedGyUuKZswW12BCAkgbJJmqBUUwQKq5rFGQ/XJE5qRWz1AjRciTeGE6AgTNBFPov2G
0TOpaxJ9zPmblWAO3FcHmKWc1k/kM0aucpJrMRQWjBXK5oNO+v8Ji7w8JSFQp0Cmy/TJHGacS3yv
36az6I2NvW3dxzZKUC+zqv8hhgYf+DqZCufrn/w9OUdoLQWo2ywOXOWNKOVn8SiIOnVNDV/04ygL
SaK2V5VET1qjrfhZSYfX0zvNc147euFoxEoC4PVZE2bYjfGCJ/1oYGpqvXxmJgz+bPIVb7VIUXOX
2AMzA/6CttigZS3pLe1a8RJWx8lBqnd5WVRP/npw7ErAnwapgEOS9N6HSAMHOCL+5IwHstkyBVxP
yI54s+KDN7SdsYTIWnM/H4KeOpejPsLawhHhyFjkVB7VWB8a8d7k4AjT8mHBli9I0RV7zfp3FNmb
vXXTtXVQmQGgbkPoQrgxEV8EFAq6NcxCEl9VgUkHVHQJe6mBrxS2uVw4+jqq49VtqWwaGfclnIf3
CjQj8NQaWjYSPgBOyele8PUzKE04eTFX2Gkefb/FyBQDh+J68knHEya/qo6f37b+aTJSG76VwRoz
kZJEHhzbtzV6KNie62nOqWYp6AXnHZKLVbb4XPmubg5FHlTIcBBdChmppInCri2cEai/a41HxThK
HYMqE2gWPHTGX+R7CbyFPXBmaqKbQtIV8U6uoKcvW2SeV284JHNASvrxNaoQR4OnPOehfNw3Y9Me
yWYK8nM9x6fLzs5RLzUh8rg8sp76zpHYnwX0J+zPR0PgUyg8B54tzswAVHZ/9glUlx5WAiY2yoVl
ThgQq7hSvPdgcil3EqF2SrxMp+L2P5Z3t0ddfvjYcDdbM45vav6O6IqTupy9bYsF/53okv4tuOXH
bmmgSZhZZ3XeDfPktO+gHN+2Fs9fcrO+4+WiWxZq2kOs1IlJ9fao1C60JqKBxQSKckqGxZVLcplf
G6nKeKJCOr7A6NxymW/lOk91/49lxdZ1R/4UxHLdgMdnGAWoOlBFbZxxssfCUOrN28eA0pC/mc85
t/QBA1FcOiSYmD3IWT/EGFQprnFUNQDjLTOltaYGS0QYi0SV2qsbLhIPCjWJMsw/tY3gqgm3KAp+
cAldfX3obNflg0tjSZ63KUCZg4wG2LDjkjLATgnvAOUh/eCVSP5yQwnqN43Hk/80WKYAPTSA8gD1
K3qIpSbkH2eQYE80CbzFq4dmJgfrS/j7res+uHODY6EsG/JjzeKcs62DBjVIl5F3AzNSOouvEnNH
TxiZ1hoAwQnPmcT2a5HrHGEVYPqewidmBqeIBP7VzitCGvPnB5cW2C1MpqXLJxejfTajDDeAIG/i
hXuvT3KbfQQofllZUVXH65dMtg1ou+RaOey6CORRFX1Xke3jLiarcrPSyf6ki60nAIi/UMV/YP5p
p8jpgQgBOlawgZzpfjWDJDPqfnDyj4vY5F051zqyDUkYc3+fitEzs/q2+arhZ8793u07oOIfSO9+
oUnpEcClvuXiXa3RUXl8a4VfBzF960we54ZsaPJNSm7O6slMo3qu0TRknilGc8wCkGM0ZHhy/d1e
pjXOrrKzDFwFj/TE39/0RkTN8plqjIdRCaJbqyegEOhR//3cmhjKQ2Psc5N+8e9lJT4EqELRFHLz
hJm2c+o5QnNJ38+tpjO3yrmvrr0DwHl50Sf8rYz//HkQuAIo0Eb5ZhkzNO+EcF7mevrGVwgBTYAB
XQDyjoMvfRgiVfWFKBxYnfW72JLOql3e34jhNk1yaFJhRmCLrjgWDZBiDZ/F1crv5riJ+o94T6CZ
iNjUqIt0eAA4pvgZ+600FAranX1TlauJJ1s4BvnhL55FQzAR/hXam1XR3EZgfKfdu2tZRd0m1Hao
LRttHYTmPihjn1jr9Zn/03udJRbQPw7Mzjs7JMDuAykI3FY3NgzyPGVuNDyIbaWZx5RHsJtOcozi
a0bXsE3Q6roXDW3K2oQHCbK02R1ilhljgzjZZOW511ef4Z4wpfCpsQcKuVYX/FsL7lCgVGPtebsS
YG448/9isDV2pz+u3QLJUNxZoeDRsZI45QUlcK/bhcYlk3XfvsG3QNStMcB7mx8HOh9cnFYkwRkT
pk9MX4FAElOcryYAQ5omb/xStQAXl1IRYDAmiqiCJV0IJIVw2zAeFl5sRdJcCOItv6vnYIPWP46N
MGkKxM70mOLqrTZKnsSSFLOZV30rKHhs8h8hyEjBHEp565D+RwLtEMgd8ZrfYsG0QxkEEovx9MrJ
EHEkkhwAMzfjCQkz7gkOnfSqT8Q+gzWL4d3M7Y0ECIoG575gsVeCDLSXX9vqskzHzI4QxfeeFgYK
yzxXtpq2o/mNWp3jM+/Fd3v8vXRRIlXnJNSD4jzAO0vS2omt+zVL3+D+Oyja877nSrnudKFjmiQ6
zPLaj0Cc1jrRVYCdE/9d12UK6G/faz4mdyJXR/2YB/jPNISPHWRmK7KRoGUC/2CutwTWxXDCCUyF
m14Zp/dgV1Xw+NGxwO+6UySqE7J0OwTQtzlv4KLIPTbzbcykamw2TbNDoIP2KDqW4XqOa97EEP5a
SVtxYiNfe7gkPhH8jkFXfV/nynI7+Zpr+IhJi01D56xfb0wj/ZYZNNzwKhOfO0op08YMbuwOTrMG
k+zUJItk7HJO5dkGS8J+8HzVQoHLx0j7hM0Q4rrcf6x5h2aU2ehUtccdAoV3ELLrQUGuUWozHS0f
4F3LcwZ0gGgtX5uXdIiuawtF56VLe8ReHKL3ZE/HJe8pAdfZAenCDlnvKTYZWfD6HumentQW0UwX
RBOVT7YBl7FtDa1g/wGC+NAJkF7RVQdDN3f7JX6cH1eQJCB10kpCww2TeBAXKewYa+8uwpHBalyr
mouad9pO0bFEEGw1e2/Ap5vmQVtGbHG7q8FwshOz47+tCx5qF9U9vIxifYh7vIBDB3iSVIPNsNxk
Fzgoz7VwJticaVTql8SMdxWPiP9C+P1zDih0aDcjmvijhAjbwU7cQaRfE+73bnQk0NRFykEz0wn7
zgedy/dU1trJ8f5OZdLEiSyuAFNpAjv4ceOrUOLNWIR4wN/N51Vg2uXUo7AK1tBINMjYkdJgJc2g
vYSTwccAnPoqMY1BrQmX4Y/LqBVT3BkDrqEvVGebzyNztOnDTxHrqLVMq/b5ROTImLMdijUWz7MR
Q43L5TIJUeYQo91tweB+mQLsvBAOLUD4X0HzgTYQjeFbsea2y+bhzn1q3RKDPmc9gzGADvGWX775
kEIKmb/QbdeymHHMoEgt9YF2HeRwN8i/LrUL2yDY8Mg1p1d4uHd0OgabDi5Jo3PxVkukKU0ggtd+
ED8zUgMHFaTffes/Zd9QaTgIEyVzKQW5d8dwPSR2BVuqSe0OOHKC1+N3S1nIyw4HHhV+aEGvWqyd
rRV/bYUEbH56i0e3DAV04CD5+FEZz5t0jbmWSDQfbt3NjA9G71/ekvGeJWruF8ZrxGiRD/TAT84P
uSCXgVuS0QeIREuZjCOkbQzJiX0p/9pMeXA9L53Fk4m10PR/pfncvG9mrat7HMLbyVvq/ja7m2Cs
PqtVWlBwjFgP5IbhEMfJuuas16UvoiofmutW+iBHAul6pdhIvtQG1cQ4VKIiz+B/oA3ovi2iHGmM
R80K0Ni4SSJXQ/jEV0xs126xZyZ8uvE8ERESkwASidg3Lkh80LYTcfXinUdxB9f6Pp3w9MNECYEc
RBObfhUY5O/zuy/YlDzfXSnfX0k6ZvV1iiUIyuT379nLlAQrhjBLEMcFU7ZNzzFnw5FutC4B6tYB
nzly4JrHRyT92RLR8vt5cnYL+oZaCAJO6YGGJ5PyKEFcdyXYwtOxxJFkfTrY1GaUJ42kkiy7zBWw
OnuL7C/zOCdFDRBgWE9Tag7i7uj2MY6M5xaF/HwIKMvKKW2sp9unWHTTOeaIUz7aKUAXSNawQyIh
vSf6qilhmS7gSs8JQfYaq3eQFnB/Jfz/tCreEi28J4Wh6ioIDrMNtHaXdixS0BSfDMo/sYquUU5F
N1lgig8OGwsFB0CqxNB8bXfxM7An9MEeLzCXjxyvdOrcma580wPUO57wB8nsjqhMaw6Yknkwsd2L
4sMs/ONi8/z2Gp+MVBS4TYJHXrCM022zQMNZX6scrcQRRfYo2vYnm+v/U/9lXoAG8HncE8n1PMdu
a0VgabuHDEP57TQ0ntj+Jtx8TkUWtbBgwlJC6p4J6cKTvTE8eeKK7SbYYyRwrqxltg3WuRKC4hVc
dcvrWAKhRIsObRlH8yzHaHyCaATgk8jEXFI6+tvc3A6N+FjrRg5NPnitsNfT68P72U8E7ABemM4Z
GaFuaLBXItj9uniPYQbOFj7wW/VqGRpKodnK9JKfDjPZxq7zW578ZbwY+GJ3lmVa7KUO8Sv8ETIx
X4sGgLgG3+GxCMQUNW3IJmmTxpqxdCMhZuI4IInhIzDIU1G4l+JYf1qfuPEAfHzTadqwSbSw66yf
LDIjhOO5V9rZ5esatqvMqIIIRZpRRKz8xoZTu6U6dKtM1n/6+YpUcZBS3W0+Mu+NEUx5XJbuky+K
rRrAHRMZlHIO2CyNaX9YM7Z+PCR4EUQb4OGvTJ/DIgsu6t1m/ddY3eZa46RvHF0KpDaWLFIt5WBk
rqqygB3TbjuWEHw7cGPBMEx7A98zSbbCnV2ipkGcQXYsFwWXe1mmQkjdz08QJ3hzLMTcIjXU5zoN
5JNYXZBBXFGVrpT9Z0CJyGZivQ0tsNtua6/YpriFE4RM3nYMNF3D+IjBzC3SRA/D5EtBeg8fZmHs
KcAhWRHcu5Un5tZ7P/b6bT+uJ+wT93LdkadlGDCqx73xY4zYcMyyVJ6SfIbyOoc2dwqn1bBNjHkq
/2Pe+dnNhoUnKmexGkk0gea+x99PavyIdxy7DCbcGD3n3U75PUFBY1qbdvdblekwrcThN0QApqkU
LYQKItY8XcN67T0cGi48I+Lqfk/cA7EfrmbJ7zjir7JkNUGUTtHc8+JhVtz7TD6BBBpaol21dhAh
HlflCJon0KTRyPdpDBuQZlqBiCCTdt+v/ONCLTZWujJrnHDOHajvOSse6uIUeIrYwvB/jJ9PA69k
gc3c45if1qxfwvr6jXu9nhd/cCUFOt5P1ve0+BBaju7idXx+96Ik7Ryro4KvTSlARfKoCx4+3XtB
7LTyeJULOMA6blq7hXRZ8HypUCd4hxpW6ABsi4qyUNL6I81GKDHkfuEc0a4AOaMMjaM+pg0HGdSo
qXlbTtLJSQjtEEjFpkLA3Iw+vXNc1sg7XXl6wWT8jJKHv+rwYvvbAzm7umaGJUb2aiPtFuoF/n0H
XxRuujFA8/sG5tP2sQ4KV4r0rIQWEvZE4m9y6vf6Jp8z5MIbC+l7b4t5jPEhl0MW/nHoGXUz8QRr
LOPUSnFCQD2KVLHYxxe5gRAZD/t47Q/AHSJHi2Jpmi4NDS26xTR75YyPC/Gl6Z6Vfa5xT9fS1Enw
hsqyzX8OkUO8flTsbD6w00T3oz2WRIrrByP9oa8FUYMe5ASkNIincwlJEao1iM8sr4mQX3c6Bkzq
i0BnqNkZetgA6Y4+1nroBLaU/uoBGYn6cJNt3RDXNE06P4DowAQfoYr1gsWYKOtU+KXSd3HZOBjl
EJRtze2i2WqPA36aJH365jlfpfSeoSKPM2Ut3mEBTrroc+OXOVMmynSEBQW0UXv1D6OBDJjnMcEK
pMWarzoqy1WgS5pm8e9XFcvMZLtZHmMvEJaZXdhgGvuwtQI6wffE0N3R2KtVPNlnYbG8q2sMgRHW
KaGEzrGnXBR2gRxFb6ReXX0tToxAbH6sYIqnqsOg5d6UxLnfCOZw+eNyFNXS0ij8ChqmPb71cEil
MCVerPxBDO/BzsTrpgCqghMdwc1N7bX0Ab5/Ft3teXr936Dhg0x+euXJg09+7qkbR49czIVMpRn2
UllsO1VAMgXPwkZ5qkrmkiwBnns+k1Am5HxOptIFArFWK2aWnRaUxSTeHv4awv4+lStSUK/lmST0
I/s2bL2fRxh2MZZ7GQvVtAcBDWKNAGhsXG0N/2kNbMcN5a+is4/Uimam80lAV9WrSnkVjvj2UOrc
zE5BTk09fb2jB40rN3IB59DM4nayzBFbPQl/TJaf73VYjNJSHCY67pqwU+5DMMtso4HRZk8BpVDh
xAVQqpfp7wM7M0nPxxVcXF/oSFXD6+Xz77KK0Ioyta2eH0g8+x377fVQZvSu7N5BRT99CKf6QL9k
7hkFZtubNgacrcz93YL3JdnhV2rXCH+srE2szvSnU/3orSB6L5ujZ/4xOfSiJWh7OCGKiFM13etP
ouHgLims3ZJCU+9JJ/XIJAqpn4+yOKiZ5MXi3jKE/EZzjdm7zqQlLI9nSZ+SU/nArwq4BM1QK+os
uSkq6+WGJ/vbI/mHU9pqlf5tCbh/JgXkDo5zI+ES7bX1AWsFuCxZ1OtUDTm5OlHrbBg/crl8y3nP
BAWvH91hi3Sd3bB3Xv64ZA/cWq6Wm37+iK9iymclUNKToA8hTRO9uyVxIVdrAPeLC3Lh1csRUEf4
3m0ngP4lLUnUeHTphIE4cxn1laKWDvXuQ5MHhVpNoz9AUaZJXWVyfFjqEJde774+lj2Voj0JBq0I
n40Kbr7ilplBsa/Fvgq9D2Fw7LmEyhMDH3xIMG+9Olkl4kx/3VaqS7xa1bz3WzAIeIcghWjlR7TU
Nz6nSMNJ4VlLfh/6tHwC0+q9kihkzR5FuWaPXhKaSizgss62ebiyKtJZCLxBjKjkAd6HJGXAhOPQ
Obf7JLtoYMg/9yZnA6VfD3xhVhVrFdS6GRmdgZuyj6vIdWT0+i8ZwUKaL6ZNdz58e5YId6b22Fwe
zs4hwDekhFL6oIF54Jy+ast0ziUdm03vOm7tXirYN2rDVVLWpbDEgSvKq7qZUtzw7FCCystvndUX
D9cx3bWrTKTVDwZO88+iB/jyODLIR2YKbG5HKxR7JIvyQYM2iLsMgcyellFeaOjzWEHXPabPnIuI
JJCLJTz/2WANHceWT/RNWQbJ119cobZC8Rs00tGvXKVxWUiuJ532yz3/7S6IjrmOKt2kpbMSHjrn
9l0O3Zj3QtnwRbtuirNN47OxePhE44Anp8zVvPE9rKzi3NZNJi7M7/I0R9LKCQqvajKH/ADGQCQx
hXYBd6+HisDk3OsB3oMCpmwuWlDSzcusHEfh6drFnRixS9IfYlIzqi3lR7vpvdraREkFbM6Oo4ib
Qgw9eC/gB7TvC+xIVVPHc1edn/h0HNqsJx+jCT59tuVVaN50sRX6PLBMZIzcBVXkuzkoHkw7f4Yt
V0lgkpzU0HJtpxB1kfjeoU6flxcAyAv/2Zv0Pw7qReXi9WbVpD4r5lluMnE3TsFMPUm1+AWzl+wz
r3+ozxruBdEn+14V3xj5AfRaD2UWhANKZraQ8DgpxQUy97MUdesJYqABuf4zfcejMKNfVZ44e42y
mTBEg1zpH2XY4gmh9pwvLuJtCGmtiUJYLtV+7tgqscpGt+uApQm31nU0Drm+c1mHWLfdnpNK/Cm+
/UfSy17EeIFdkVy4z06uMLFCy7aAuPIZKDtq+hyph9kNnYBrEy17yc2CsOFhKpCLOdMpaIPuUeAD
uzmUvaZuBBRUE2gOx4oFvVwi849/hy5DRiykIq0Oul9a34iEKMRFgnWYcaTSRqdBKTz9dhj7BhVR
4PeDrWD3tTUE+5ZAWBAiMwO04pvvfdSjC8nsF6HswQz18cKCEuL6ZjcXn2qg68Ym+8U2mwmRVVWy
ZlP3Oo31GtKSruBpF7n6hjriVU67a4IjXMihXsugK/X6VCpDN/4QjCxbwzBV1XRVKtzVE04xN3/+
C3H0qMvRzk05faAsGyC10OR0OCiDWdrfCJ7j6elmN5itA7V4COcMbaMNDx1X7RdC3//D8Y5HErpX
LM1fLs/nVQYOH1G2HHk/AdQ550b7LZ9+xCJ+qgETKoVnzVch1fcQggJxTDymQQFRmlFJEM7Nizkc
zWjpzzFb86CGNesve7FmfErz7QTz5ZoqYx+25zLf9c/QcYX9S/EqU5wpXEt7D/TEiBAb/Bvbi2Rf
PDTX8Z4jcWpuaRCpm4CBtzFWIbeyhdeO71+NFozVdg7DIo4Pcpol4GO57QvzLnSS5dE65hjX1a6N
xyNgjT7KAUC/g44BTFjqLFB/2RWqKueM2YJu13tYN5l+fOXKSayXrx3vAFrdQZ+RXrmH+2I3Ov2V
MWRbHXsKZMV0eMu+4z8EM377feqMFX57l0szZqknLEoQM5zcoc9zpDSP23DRFuxjkAD+ZT1Go3TI
ywi45OGMj61HQJ02+B3AIYWo0alaQQute3NlC8v2gfQ9SMEEKFzzj34ICOQc1qo67qbpwrDNgEqY
Gj0XD22G5AbhEQxF8OeK4kV0az3A6Ja7fYzX+wWmZGv/FilrsxN6xo0ePhNr28q4DDKtoscMa5Ur
ozPGq7rEze0M7owuFmuMNjk//EhZ1q2VBJMaE5mgZLbDWk36Y44bZekGfO4d9mBzHFUqDzEUT7zh
XtwfJRmUWLMrTnCvTJyOKWQsHPQwhGiyDMjGTxXJNHESIYZtZeJxYjXwZMzU9qiwmeX8m0Z7M259
o0/S6KUKzAU94sTsS7bumbOXFJtLuCp0tVDwqGvABcaNOn+VU4Zm5Lnnc/s9Yvljc/gUfQImhCY2
gBtHnx4t/Mu5hPzaQ8dG6xx2qNnteADAo9iLEhsBqWLUHdFlO7bGkawrueMHZAfKE/r6BqK0Pms0
Qha4hRLS5XDK68UX2zQNEkusZIvVGngGR2tWpuL5wa+G83NuFIz1KR5b8Bt3x5LfI8cjyc+KsXbA
dTQ844WWMWaORQEs4vTiIuZ4z9J9ejHp215rrXNV+5ZUoX9nQxPtgEb1rO2PUmGtHKk6EVeuOTc+
nLm6LgRBufD6irm3ZlZcf/YtDfoNp6vdBMe0gQ7MwcPE5HWNFjvH/yQSG0+nlHQnWy5A7IJ1QEr0
12doqlI6qrMm/ACBQ4yiEUox8oLupturNS11fxrzd99M8FCuVngSov38Fvn5rgot956VEwKfGdWc
1wEr0b7XTo9/WSKeO5LFhVtmRwyWeN6sDODLh0zwrLf4odmxGWmy6Uh7mp3o4GdQWK/EF16EBJOX
/zUvSXjvpw5q0In4HJXTW4A2C+cQj2EA59HGeqJVqvMX/bgHhs61idVAKSL8MH0mDIH6l9jb5wnc
ZmltSMRG8Alqu/VYI353L0dhtO6Irfom62mMik4Tvniw7Yr0a081iBa5/WT0ytdW1jSCfnZRMeUE
9T7b9NrCcna9dCahaYkKBDSh9ZAT8BqLWRnfQjlrkSCF5c3nlnf42a70WTTj8bfHsgCzL4A29LmW
NoOL6+Ficnwtj4Uv6YxhYe9McNextKCZo0km2dfU7XDcz+7P9G6qvNSu+fRQ3Q3RLl2I7679F3e/
A1EafPPFZQoDEPLIAwTN+sUQ4R4PDDXDiofFQsq5loWmZkMHf+YwZKWpHPF3JjtvIEFAl0LBITwz
XQfJRTVv8QZNZeIBBBahZ091pfwU9c5j6Kz52OjLWwNzhcQyJySp8i1njhu2XVmo4YAgvGuzERxp
9aogs911A9+e00roxRzDlrTy5bkPtRZPENq4pCIfs6QcYRYj4g+kpqRrez8OFGuOkCP2X6Y0yJtz
Nflr5DZi+6uObxcZjaDut2SrPzTad15+rlPYXePkqKbpiAngVYUa6Dd/CEzfuHrfdCpQGkt0NQhT
G/6L1QIH1LCGfAAIJoKc2zlzEAuWbV5s7QNbKdSqUQ9pAYT47xkOA3Nm+UTKNX5pOtj6SttNmVM0
AYXAo3flHBJWebmrGYGEseFh66QAKRvfyYkHRZ7YiRdmWo98htpw6z+od9A+XwYm0yEmTAQI/uHN
S5BJFSzRKOJCbiPwwJRik48NM6I3HJMLdIFr1RtLnn8uVxN61b+Eq9pTNzYhWye6+9RymbIwBFkM
Gzbtr757iYAAOIjNwAu22/FpoJMF5CbacSagfs8Qdj9xPOtgbflRHlu1DfchyCrs3P9IN9JQi34m
RCjm3LyvuXmk6KNo5428IE+fE+hvrNc2akg4w1uG5HjJ2cK4w3y7AaAZLu9knlSY1WBCrraLJuUp
qU2LDqVZpXdXQBPJwk9uVPtob34ItYAX2OVpQFPLFBxyhEeant+gXLgaqozEB2Lv+TDItWVkKAzP
bdHu31W42cxfgLgnU/qPpTTBLS+PlzR67ZDz1w7qrqvnrYa2vXEXp/TzXUr67dU3TBjHEtFg1+a3
xuGkDalrH0R7jPSlPqsGYuf7+N1vPvSCTJI9ymwMVddwlRcpkaxd/1aZuFdc7Nf3uAbtBu1GkHgV
Ve1BwFozh31h+2Qf7IO0d19b7NGN75rL5TduivkjwfQh/zBQKzZ3GvBM9AuxBgSMR/M6DbXbZUMG
xoT3BXswRMsYWwxYaHhqnPWfn+al2pkRAaAC8ET4N588G4c9ND86Cghi/j1eF3Kjpe7vnb86N2e6
owoU2AC9+PBSjs1gCMsDsGZBkmuOD4Xvk22Om0PYD7pXAzEFXNr6ztp4OgFVYdGlhEMSAodgWjoj
MgZ6rND5iAj+04sMhS9AT9WuIPqciIEFxU4P5yyUeKKyi07inA2UD5RT4wMYAfnkkXl5KLDMVF2I
PZ/IjTU/wii1e1JUAJWiILTdvQjlLq7goGxnFcSirh3tPqVvgBqhngjIPuCc9HJycRl6gsPIGWY2
zL0N2wNJy3t8w4Ia1CsSkcrUUZ9VccE2VfW32xtnDmLQzE6esqKuJXAbO4PIWszDmvW0NIwM4Uhj
baYMVOpBge1+00i2ew4OSOMFYOG/uhsQ4HUdXhbqseOCaJOME3nxbGMDmGPAw0PMP5gF0TOPBPG7
kTsECtE5XM5Ts/8xz+aPPWTotyW9SQbws/Pqa1VWcACoE+X0+ydEOoSa0a9NmVFvZGEjyZFV33oc
7B67IfzrugrAcVq67++bOon9HdhgWUZb60/0R5yM52lvx8e3vLy8zQotVZUkKP3heYpNGp4BL+Yv
8EB4c+b7B9yz/axa5CG7SdYzDBMLONeTTLLkilOKCiCrUe8Sgo9ApGaJzR6FsCa2IUe9Q74U8+Sf
9x1Us9Tn7egj2ITGt2GrtMH7hhmk/OODbGPUuhHJ3rmS/9bA3Ccd4Wgs+mBqt3RjnP6I4o/kIDcn
nA9DVZ57IMrUCb4wyUCxpHEPviXllHbSSLKaCjZfXfh0b44OM1rxNnqmDJ9V9DyluMvIsugC4bOw
M4zZMWorKV6w4EOnaA+JxXwgXVy6nJ9C7uSuwVnUTTuHoTt8qeFLMQg5rwjncNy1Oo9cOwdBr94i
L/aJfHldzl+ZtpuwH2bYjyuJ1zorFJ86uE/ubA0eWXo2wt+63XXChUB5brnaaMEI/Wk2RMbz2QFF
54cm8ytzPQswbBMKQmNRmC8DkCElLXukXsbxcJZrkgz2INL4SVht+53csyl7yceymLNf/fFsp5Uv
GeU/EjjuPO8U22Ul+TfAiOCA6NAlfcEU3zBTyeHeK8jDeRSIFmwcWDn1tIXxbCdAbXQTibI2m2l/
IpmRgO+N0mhvc0kPcjQyfPuRn/UBz/L29QhAXD5oIeI6wvXOysCpdxn2R/FfQniilkBa8EBjub2N
2sywaP6+jQUA9hWibgOW6aPjb7+6bjhzXVFhld8Vwbosdgh/fW/WhTnpvFShlY6QOggVvA/sRg+c
RcCES0kSn6DUHY37pCwwWeIUgEAxNK7/ZMYokErjTkbmgJGQo+xK13Yf4btEECLd3xojkAaPQ5Kj
S3O3Gx6jG8eYxX2Se8/UD8wYRdF+tAu0WkUErLlEAy1vBRF2kCmNemRIIIwCIKZdIMjWv+L56cgO
VvI68aa3Ivw94yDm0i3Y3T1fVQXqQOe1ehIFGxpApHLSwlPEOVBt2tFOfQ/cAxtJMbrvj8mCax9N
uM179tfrZ6R8S7t3DT+aarThKfo2hnCXaV4v8yzZu0tlBWs8bBvJEPd91kwqilnRicCdfDdhKoSV
0p9OCcA9DmohgNQjMbi5qcifFzUbhlPqzAkikwB8BNq4nvc07L5KC7jTd9PXc4Xrmd/3npkwqDTT
NGthakWZ7JqoM9AdoX73538Vn7bYegu3kItRTnusynC2NQeSStU2AKC2ILLfjGiSAq88W3Ds+onG
RShsiWxlMGRau4S0wnze3y1miacbqAP18T+kFWVK7Ewt6QdtfhheYGp2RrWt7Vqz0asvunwXvMzA
h+zuFb4sShiI2wU+jAM1mBRW52cumj8dVOEhq+CGCsbhcuyVw/JDq37YmMhXcFM5hmWm0FPEJqgd
mpzboWrbx3xaIMQhFnTXW0flCc5A9a+k679XEwEtEfkb70uDx8IAIpHcN3fn8iNy7hE9351Hyf/2
snN0UsdYQrRIIiIqSwx31togHgHkNSKvMb+7SZ8CJVZ8ksDe69oy6MUdUl+NqE7Ngpr66KlLq9/z
4U/DE/eKlg9Ym2C+Sy/uzZAt0BWWA638meBdrY8vgYyO/Ycne2LDZUBKrliaoJAa+30INSxssKg0
QaX3LAEX83sBtFHI++98ZU3Kw5uwTTZ8I6Rh4v2WhCaKhCnMNsVMEebg2LBvBWtDVl+mtUuMJspi
QTxc5WIvPaCvjqX4uFVpH3GSG0aegLcIYdQoNrKV1CpjhP5T8SXFL4bowRfwBACrMoSPREA0X06a
nmo/FMrTLJSl8OAsC1c3C31Srry4STQjDjQ9IqxCEb3HVC1XDT3pbezbTW2yjYzGA7okCZudi/nC
q/hAgbnCS3ZdaXW+KRwz0LppmwJH4f6T2JUSgFFoxHiCh6OYuZ8JSy7EKsSJ6O3uMCDlQAb7Y3+n
GmsppyIWb1LLa5WaBCAiY0o+m+u/E5wt3N1Vjg8Y8oKsC80UFdJ/gKaYmDhLy008Y5LpHzIzDVuI
JjQSuAKejYz5aQ52oXd6AeqhoVWrUpjdY+KljOxPf8q8QmpR848JoatYdznUsM/4PUzW+EQlFJcF
d7Z3Nds0ETaKr0hrzNeJ/UbbI3TamqVNqU6Ua1+whdYQuVChSJbtdWPo4QN963BbLybrvfMD836S
aianWoZ/cadJF+cvx9e16ZW23aLxI4w22a6gK/sUkIu4933+UTuLItxMt2JYNrCcWsgXj0k//Abr
Jx+Gpvzetm9GFXI0wf2ejDRbzxMct+YwG3NbjSGTA5Hue1EfNcjl+U+ZgDjJkQziHtarqXnsk9lR
eWylKU1wjIj6nUdjoonGnm/UtRMzYi5u0W7pvfs94wC4Qa61VWoBv9Ga4Gjnl2VHijZljD0WCy58
6ho4AnlnOb4fGKSU146N17bA77vW0LWj4lmtooNPcqQA+4cfI1Z9U+o+5sxghol77y13ZiqB439Y
j5CYPjMoifGv00SQaoL3zdlLmHUeA0yONnmBvPQ/E+eYTfYWPj1aQp2i44FaYcOr0dmO3lbdC4ei
524y10pvNAe2FSWC6sB+PeGbQEtOsFjJ5yiBA63r+yzuzuqOX11b5n3R+tp+l0QvlYIRhdXk2x2a
6VBNA06iX3gYHR7fcKwLMo7F9E6/g4wkS3yPKUw+2N/P2Tw9csjjr2xBMWSlmL7vUj1op+6MDZA8
nzdKj7/ZlQ0097HR6GE0V+sn+TPJCRcuX5JD3DDZbCtuleIDemKjxBcghzXcjhJRwAtzsZ8zOltt
VSfkdCfcy/pb2tb6yS7N0DyIjaFB6dAvcFrEGS/beXBa0US1ddnKdzn+R1jSvmcmCAio21CJ0xay
26Fi0fM0Q/6OYRwGKq0Tv2+BiMfqLAQrmMEvLqQuKt3C4KkyGNpLGnjEto48FqN85LrBhIwXNG1i
5KbRym376FP2XQCOvyFvfnconiW+JyPqjGV3G4DRt1jJN3As/uIKbTc4rGbenl4/ttcdLLt1wdcn
dYnF9HeUi4sGU0h3bCEjUm+TiiIy41AzGRWMONx6yd1UoIGejEpK23/ZQrwjuceGmQ3+bmf1ICnj
mHvRSp1l/7kk4w6Ox/BsINq3DDgxK701EFStTT5+MRvXi0PLPecR7+8EXAcW0re5wM1d63goXRNX
dfxl7Zt/gVBaB2fhiOE6jQPC6H49sCUcg9NSVf9dIdyrjNP0nWEZ7Ga2ik/zZ6S/y07INyUhpNX2
boXVEkm7dLpJoHgMbkuADo/fLqe6z98voykmgj6oKBFFWDQJVXGk5CGmp6NDilnbw5bwNWYYFhj9
lVvOMW0Kxh0tVI7IfwWfZHsFHS98aO6D9lYNJmcytad/yuBzTtjF38vOqs+snne6i5ZXBORXzolm
gvMpnNp3UzyrMKgolawIw7u7BX7Qm8gd9bvRo7c6pfXcw5tvpCfqxFCIm3rSX/K+KIdDQAm3+G9a
tFMqxYi/BhPYbg957vz1K8MPeZaprA9xWpWINeOlOvSG0XhVJBEeEnxQq3vRovNIVFh5dSd0dQ9j
xZFJkWX2sB8FGjuIBrn//xD0uhaNs2wbkxE3cvlcbOPv35xCoSerOAryfyKhTJdwClqtFT1srH6O
YzxI2mErkS1aUBXYQlb6U6vSduKpPrWNPI4SAhpXX2ZZSz6SYAHJPOwmUiGKLZQaCSuYS8gJ/G5M
x8NM+ju5gXJa+iBqBeWTlF2nLHOVxp0ioh90KIgzLcPuvWZLOYkHLiJGQfzQuWosnB1CNuzBdzTt
E2PRF16UPaQEPiz34T+PvJycYbGIs29StuLNn1YjMBXLreIGXjyhVLGpxnPuRZto113cMgKYtUZW
hnlRComuiwiDl0Q24FqdzuNMoKCLn0UxQfHzqtXvgXZa2Cz3M1L9UcxICi4BruShpknZ2dSHBX5p
4eaTrf6KwmHleXT4urjzfTAJwQEgB1RV3hOo5/KLbRJtrgz+tZxM6m87Uk7gMc2bLMJ2S/LedpVA
ne+EbiOIXHWjhTjzQMx7kdD8yj7ODI8WURV65CWjQ1G1bQax5FtgfBmCQJlxJLnFw8phlgX5f+3a
Ee+2dt/alWsnrxh93t473unLBzkWL9NQdOfS/PPpcDXIXmSrqXjNE/2ZzDrEPhigu97Kc+I+mjfj
G/pLZ+Nn/1uGEJhzppahHO+tC96novlc2Vk6FRXtyCsMxyun/ot1Oc+l3eQakxyKPJ7p+/Q9v6gW
Sn58yKLiG0gVwdDETqZpBNVu+lrc8sk+yFftda7/X3YrGSGJQk833tmePI0uEgsLYWGFbqe+a3IM
PrTzX+sEl+8eGUngMKQDF1ZomlPaikWWZhKwW9EQ9AR1qM2TWFO7fgEbTq4V7KkP8SbefS4D/5qC
M9LKqEhKtPp98s0mvb7zQXjtntfNG4Pw/EnvZNOdlApadqvFmx4oTwknnk6mvYfVq1gAhF4oG9eQ
zmAWvKAWNjqe5M6HugxzPHi12v+fDZxzgCUtzhwThrKqGFhyMOswni07LJzlrIO9kGkQcWQTnZHs
zq0ky2VBS0K7cSqTZDPbMKJNHpk4GNZ1spaUq/75uT3RRtBZ2P+3/WFh3JZ7dBh2i3MqCatJNme2
5bCrRLv27Y2Z1T/Ilwv2oXAAZSX8nLvWagCZtU7cPGpwunIlbgLMAuXlh8mfyAbRRZSACRERvVRe
1+BzajQE5XTHuiJSyHnewV79gvVo5qR0gB2AmVydoGFmPEKwV4Su+AI9i8Szr3ZOjeRjI/1ny7Oh
mtmHOlPT93dO1+mbM3cX/D45pnCKaEtOM3nSEXtywQ3WxqH9/9NS3ipOYkjOOfvLJ3skcXCJTyOw
qW8MXEMP+Px1JOpnNlLy8qKDlfqOy4x0gdM6PTZ8uf0po5N+Kfx+AyurUUYyNM7LbudW3o7Fi46X
X5bWd2pcybCSwVeKJ5t/z48HcM2zCXyjR7l1TI3g4EYLmSU3JAo2e7tti1pT9yIU0R8YR6+PKNaj
0WeXB+xFvW907blYmg47Q/9NrKjmVUBCM+wBt2deDINFPA9samDcA+Bg5FoHeTdRgcV8/XFPgd21
TzVtHwmhoFah3VkJXhGRuty5d21PhZpTVqHjhgK5rYGbXevOObvp2+TiGm00sQYVS1Oj3ukzCqiO
R07Q9WnfM4D47nwOLqcWD1s5iAIw/amFTZuucTarwPTOb8r26xFV53vGSoSh4VEyZWjffmzWm7DQ
1nWjGtzR0l2yJZH+fiAYzomQmIigPEbUYW29I65tyQ2aqS90HqqOSaun7E8EdOvOf47NPVrbHc/Z
7iddOlWRNwVmWdJZemGga7L/StQVuvnYVHQTNDFxSW7a3GK2HLPYkKtUZteG7z8WQUFXnT9Gxq3r
/KtEPDKnP9wlOqvlFwgxBe6NyNmGR8MKiNDUj36pdyCLRHAgawq9hrRyd/JqJdjK1YwDNu8GQAtt
HEEUxoJpbOVumtf8TEWBu1Hb0JV697/5Qn3gIJPZlUcIJcXcaFE+8dxYn+y2VGTa675KNzHdLxVm
t1BV4sN27HgejIH45/c6sUjioKIbS8HUl2NQPbDAhzoeHH7xV1usKspGB36K+hq0jsp/AHd/iqLz
N9bO9SY+69ZVfzamUyiE2ji8BtF0Xr1/TqsLaxV1MXu/l6yQZaz2gYRAJ8qP3Z3cv3QYAAY0gR3E
ECOz/8chwjhpr0cQTs8Z9npOIOQvBdNAnoW5IfBGhTgKlZSm4pfpij7bR6fNkE/XJ4DFyv2zja/x
YfLgsvG35aHrKWz6JMm6vLgasyHeQOVZh/JBBQ3NQQXncEFu4H6YjQjsVbZt+4uQc8fi9xIZvoyl
hp+o3VQkRBUGJtscKTmT35FrbR5rL8eo89GY8oY05gdu1yideQNshhsuGIzKzESWswYI/KDFx+TW
pLtYYd6miEEOQbxr/CAFz6aBlHNqZ4KZmmBKYyXEav3AuOvkk+DEINCtcah65WG7S2FJb1I4Eo/E
i5eCkd44t7qqE4XQreJx+e6g9HbdzyXqW+sF1N2MDESFwjF6dy8ULi/B15vZxTEWkDek2Uqnb7Ct
5z7iQjk6xR+ACZBzomTSbiWFyCQWKz0ldaAG6Bvym5i2wYG/WpDI7HAnCvy9vJcb04D24BsAajYt
kY8AGa2KALrY/X7rIqjqgtXExYUd2z8IPnceiyAURjjofjTJyiraKKfe8QzRSIJWkZK0bClU+Vdg
YdIK5KDpPvHzcUF8qIdtUTSCVWvLVtjUJDxsmJNn95ovaX7s8Yyp0kA2LBkjiSiVxcDnxkbZzRNO
KfabExk3vH6KKsittXgbuFqgJZZawcwYe1E3FvhDY4dqcSRyVzdZwNbJovZ7GY7Oa4JDKWHigiTh
n/HH3j70jbCekNiwV5jODPazMLNHZ+MNh8w4oR6md+NOuMrqxyC9eBDhpwMrhPcI30m+3hh/pMJJ
7NCcw+07eLD+sOmBsW7jLBbjAPXO1yYMPm0PSGAHJsz4CVo+CRRq9R95e3I9/7/TzFe1Iy9tLmaS
P4giZkbQO9hXVGPJlzyyvHCWTPRbN9RrnkqjkKBfb+ErcKXNyY0GI6t55XNpjmCj4qR77Pl4pwvh
oyQFQMXe3qLukKKj11OCYRP54MyAtTE/raBXnqNVn3sH+S+kfzIA8ZMB0v/xzx6PNtlj39rIt0JS
jl0nH25r4RwJkyq2dh1UDbdIYs+wy/e9ljv7icVtYobAljfNcrYF+ZboPVrbnDCJIAx5VPkQlKwt
q65kAryD3q9Lx9ieAFvpmlejLSf5355jexnN9YVDpHgXOI/w+ajO3+uzNn52N8/2C0b+qbtIiK4t
Luu9PRqcZQ/2qolTFZ8oUuZcwZcqQ9OmcvhRGpJ5atvwa8fSjpMI4dHFQsWrXe8IvskUU/qXl2gh
l8frK7A/tA17t2Qk3eLAO1w4/r99ZzI33rQw8h0vQRIvxo/R5DagDCv/e3tbqU2P6rXxz8wEsdTU
83I39C3UUmi9pX6nPyP0UYLO+LBPVOyrLQFewkdlmCYYOPMXqJIxcXBgEpvg7urWrocf9kBHu9lC
syrZexYFluhZYyTN52GIoCJlS5oPEb48NiVS165zK3zRz0Ejq91Gm6LEJdi0DDRxv770vohI9PQq
CmmV67aHUpeZeK5EJwQ4eSztz56JPWf4lH/0tpGVvVzwo2//LDYS71rfI64OiHbINhta02xjJVjg
effuwJBfdCCmy8t4OnshygsgJk6DiI5CmPYc1RSN+QKLIeNMECO5cMaMyjl7F+Uii+MVlGNQ2alN
ziH5IGkHr8Wv9Qk5KsglliQcfDqQ3dUqsL8SoYQNoBCBm3JZdBrlWIGgbMnW8z0WqSu/XZvtoCo2
W5xp4FFXB9sCCg24QrVnSpd7/nM4fERyU51MThcxUx1vyygO3dmzv1sA8yBb0RrXlhq3qULOnToK
ECtGSRqlA/9KCa6fEpmknlEG1ivoTtzC9+jtPNqODz0Q/cN7hJBUG5ma5U7luDnVU7eEzNKb9gK/
h5FkBjBkv3p26MFxCEy7q1qwNJJ9RAJy1SayppeVhNzXN8o4NmS9VW98OILG1SafirGzmKWsIdGu
bWV/cvVEipJPlSyOm50HUE4QYoj7mV3T9KbgnkjCgfFIUwLE5DRtcyhKv5ikTBzFwVCeZU0QZDFI
3JnrVxcnhfrItEaGap06qEQgutfm5u/nP2lBd/FqVCd3jD4YmcW26jqOIJeE8bADHgs8ziWPMjGd
LyxwCyVUwLaU8zksFynVTpusV41B0uf8UdebGpYRYYTeeR2YR76CRsZbWYR7Od0gxbZUzocEopHe
J9j8E+zbxg/7wFthKcPjMJFRQpwexGrCg5q44of5b3BxrnNDHE4wChZ3lGLj/Wv0KBVC/Hi3Mgg2
YYFXy12KPv4KwStq+wd4aoIA0pS8jKRAQR1BfPY+IQbgBweN6AHl3/8qVhLc+K8f0xTa9YK5O2tp
fcgRU/F+fr3e/dv3LX1DL15XfryLBnM9TNbMx7JSwzXVrIG/0M3K1c5IKj3+DuwvbQhw+HG0UbXV
fEJD/bJNDzJt47h3pRHK6t5LUTzBrS6mhf1oRX9SHvahxwGzHd/cnTg96yc4EA/F4/3YdjBS0cSa
3DPr5peJVHqpQXuOWtMZon8GQFDEn7zxHgjD2U5rsX0Z8pHn0WNElqQj8IyDXM/8ECM7ahSOMrf5
Ox4t9Y4AH+95R0gapOCoAqLvNXDxkFsserDqlud37MJ9xPv9ZENekuPDTB237yZDEp++kGsyDtUj
P15Efls1lJ/+gTpDUk0sYOMcdlBMsSI56BMD2LjvoJxtRwovgzsivKReVDn+C5uX/FaInmn9VmWv
DoufmrNeZdF5Q/DeRcT8o7S49DBOJMSoHfrZZCNtyrq8dC6SjbwgvBF0QI4h+GIkXmLJmeGRoq7J
VQ8x4DZIzVOHVxK0FRCt1lmtdb+CMQsN2HJg6ah2wUzYGlL3DOufpsaOWjJMd0888qCeJeDaxrp4
x0W+9Uot6J9lOzK5CCrTCHLovAFPjaWVYxm8LApCKVHSx3ia98JVLIDRBk8ozLAWQFF76DMqzoOZ
pWKgsreL2U8j0a1pVZpKlvZj6+YaI+qVX88YtQYNzy8lv5N5e1pyBmbFWOKAPa41vtko/emb5JM7
8bo4w1EcM7hig8+JBCXpEDYmGNBZAO3gMv4lnmYS6W7Hm4qn/PVBhmh4imVt+nXDN1ecrUQnvJKF
DC2NGaJOyZCYPfKH8mUQBTfBEeXAZgrqY5ISUVixy8yb/Zyq7UOdXxPvmy0pashmfHXjuU3Nrq3v
86QuWnKuFKEZmPpfwZysE/dfmD8/iDOgnypIpTZYWCNSJH4nNLmT+m3FV9tAMDG1F7m6bASMjrTV
gwHgyMZ8TpznpmABflcKhncN5gGevB9BDIpFeMGrM8XQhtxJe33G68T+ME6mTFPgkcNuhchG4Z+z
qZiN4IIVcZ630oBc+fGGmBh3hlF+HTwiDYfnt3ThnS7/XGZjTViSP7fzw/Ov1MHAygUvyvLSlcvo
QsoJvAXOjIdGn03HgLSY70u+53cfK/YkJ3dXnmZtAOr130R/5ajr9StlAdGZJujNRbHLRxe25ZhK
i6KdXcgvQn7IJihdN41U/D1U7tlsPWOS0U2cwVqDM0uS1lO7+YFSjodbyktbhzPWa4Ycpp84IGCB
EunY1ExEJVFAjLgoapRzgZAh5Tl4EZQRum2FruuTN8m8RgQ8Ne1XBUgf8mJ/nTpY3Exb2MwN6ZmV
4I9uyEuCPwy4yVx7vEFTP8kKbZPEr+/38/YIbWRUzfwc80+orRejY0Fqc2EqM6saJvDlfQRNrsd3
Q/gV7YmEJqRivDnE1Kobi5ZVO2SW70vikj93ZEZyr0QsGDat8NDXzNeCn3rXtAJoHrsdiV1A/sjz
cBZDkZqamxvZnnJYOz7OdAESejnpkJBnfZnN6rAius6SkdmClNuHR2K88tPvU1NM1u5vyiinrRqX
4DtSRaTyaaRBeXPhg8CA92QygP5LYaKfidpmrfCJkeSKXd1xU4Ia3IQZLKGQdrlwsSZqC9/diw4S
8IGsNRPkT9YHZFrlun1VYa+2QWTi8kCT3mK/glkrB5tspllhC97yDy0pEkXLFbB1dzdlGW5Sw14F
Up4TajxL2bM0EYeydlPNjFrWojzgP4UkJ9N+i+ST9NmtAJQHaLLTZ5I2gJvsosdQoJC4GQqqbxUK
RaE7tT/WAToNnoVEwk0YcTqIIWiHZlCkOVKA0X9dzgMKf+TiNHdiZH4rbM6wory5MN0wgrIRUkEw
oNYnWh97SaTGVtT10ID0vpkri0OmQ2APDbUF/zULN+gB2/4APvRMlONWUZpRs2qbdqPwIQoZ/vgz
+nMG1LGVOehueJ/lSVA9SmcrITwm395I7cGaIN7VlRm+aVsQ/pdjRhzReu5BIdh4J6F42oApGsvv
57WuEPQ1J5mxQRjxT4kdKm3mO0n3Z6AHlJP5pLBo+WJRszQYWAxsqyhI/XWcCNuhrALYerFOH65c
t8t3QUwdiXPvb37YaezMbQCh0z6RYqUqwTKAeYw/3VTOUWJ+qOvEgtEYYd8FG6zToLczWalZ2uW4
EJBkZ+5FCnaZuh8YJVqc3ciO94lDFy3FiBYXyeqLn+P/ESp2NPDP5fauoXuEbEc5T83M1FtNIese
CEYau6rVC1/KdkPHvQDkv//YCuyhLQlpWbDfmsylhyJXEXUwK1e9gyrh4CjatCfxJsUAJexTcsFF
M/GyOZWsZH7PNrfbscbn+qutwU+DcQ25MR0tq4paeSbT7Vbz/uHWT0KwIw1V2i/BeubyWMJHFTXF
kANScLndbFYTwugCtAb0ltEkIifgqxrvW78tpXi5eNe3OgmSUymjUb82p4az9cMek6KShrO+076B
grKqHPsbm+TM9L45ud9I9I+eBpGM0bwdd/2CpnErpIL1tx0T3ZyApZHbAIHqfCNLbKZhlOJQUI/S
fr02RY1a71uvgTgQlzyi7jsSohuJfNmRgIkdtnne5BXJABt9l1RVETUdCGEZhJo9LqGPQ9kqF2aB
8xU4zPj1VhhBsB27l0kbn9zEjOrXNu6W77qhUcVOqther4ipRELkewUw1jhJrf5lNCbikv+4UvSh
5jJJ4cCrFQQJ/Ku3idbWdQeTQ/uofCqjIMX5+UQSdi7Jtvocr8LkCInPLW+SQnR4qv3qx6xH6YEa
QuZaNDUSvjPWX+Z3majdISPu5Hl92i4KlibZjazObgnNHpE+Tg9MiXiXbBm4t50dxIpFDq/4cilC
h0h4tmWTL4s52Usfih2BuusKy1+MB1wrVlOF8X8sCK1aFaDwjUzSytHEknCbddyDlMS15utQvzcs
uT0W9ZBwYTq+K0E497CoaggYbuUzf6h/YBb/+PHOqFRPGXv5OYoeLZkAA7Rja9i75qDFfrFv293H
IBgVDlMTlbJkRke4MgJ8FAwOQppROcqEM8vvUbWnkElby+xm+gq1mb4Qphnz58eNS0X47QXoTs8t
xVJL5BvT8RZiKwAo98r/qYbOVzhuX+kK0KVKxIn3e44bdl/7H2FBHu36O2TmVcc1TyCrp7n0+IPi
xhPWIWc7PvMZLiabCXw0V8dunPzTjCZdRxDHpRDZXhb4g1f1YC8Ip+2VGDWfWaFlriFxIiQDgWtr
TvUDk05/aUyaU02Ll2qsJGOecjo1m1qFWssnxVtlcaSh7eQQa4Mis5PZJI+/VoY2pPvAhmfIaIUz
wjaE8S+CnRa0qdqvrovlL9HBI+X0wkm46RC7lATIF8ockbNLSRbDof34WjYffUtY2HeJaf68V+hi
Y8cqdI3QFA3Q2ErqTZhDhlFWgYflScC7KhIgNfq7qbU5tUkG7aV9IYGUFq4ooQKumIX/juYh4U7k
2lA7dNNXyS5GE8fNX2feFkYtVL2JHiLRVWHDAfLKBW/LXknK0BshiDpnksIeJ7IPAbSV0+xttAo+
CF8yGyDfZODRQdbxf5jW0yCGBNPhsUT8kHD3bUdiLnDtLNVvw9hgZoMjQ4yYBXgYuboxOSRE83vE
YZuuigq80Yug/KFyA2XY3EcgMDzytFAOM+5JWNsYHPcljZhacIKeKomcyPxRUWA2c3krcNSznvkE
/PQTBgjmxP9TEsHXIHrrKAMcnp4rvPkjf5UHS6TYLt1NttzRYDHKdgLqiuT2TDdwuHywpHBADylw
8elukSpMt7P6pLqi6YNcxU7U5eH1IygizsmzWDNptHeI0GdJdpXdgE9xnZstXbHDLKXAi5yTUb/R
h9vq/xK6Z9gA3x4Fq1YJlX5vlB9foc3An4fGGMF4cIm6xHMRbZrWyRJSeNrv9Y5naMfJk1ZljUVD
cCHjmLxO0kSQjr5XShQOIYqE86fOybKgvBR4y6LatZ6uzlEo/KXm+GZV3JicPi1XBxMJYBdhwacA
kO7iSi1c1w8iGpmTxeJ5jyEJCAbiWFXZX/fMs92FWSalHka7E1OTA3acXu0cRW13EHaSanxdjDWd
hR3Wn22R1oPdP0HDTRfUzZ7Q6GXeK2CoqnupbWbB4jCiFDhFmxb3LiqbUkARf1J/YfFcPfZ81EMT
Tppe7UjBSb58QjVZb1wmJHtDJ00PtQFXQXvxO7KwcdhzWbmViDau339z0BYuyxYmt+C/dIBVuZyD
XEvJwc7C/MMtR8H1aMlKLGGhC8txL0nkG4oWd9vyI2bAaFA5Os8n3HsuqtZ+29gHfPt/HiPN2BT5
PEfhJgSsfk9ByDBgt41Xug26Pfq4koD9uCVOxvpHDv0zP2x1NKxsp+4amuQVYRFT35gx4APVwKKd
0NZ5aakODzQ6x06oBbRvo5yHjPkdvTp5iJuw+62OqZDA81LJjrlrdO/ECT9D7JDVXAA4KOPy/GsR
kmS0Cmt61DQTAeB+d4fK37JQ1tTFv3kSLZ5fn8WhZrDwTIee0h8O3yBdqDLurWaVQzR+wX4NAOHC
vjwS4cADEhn8wBQaLneOWxQCXCgNmwYvNuyMskaXIg9s18cbMcOgmA7fD+swSttMq0wFUhyo72nX
psuKb+kHw8RMWtFb0eCdvmB+jAMfRx3l53gGSkSQHaO74+9aEz6DNEEgeAsvaS8l38DoCHPoWjIx
mfJFkDCEfIJP2kuc6std8qmYRGBZ7y8mqbTeyNl8PVqr1n3ZJ4jtR3vk5fB1BHSFzG9SGOm/KzB4
dMaavsTslvVFHT/QXKMt7d6sSVAe1vYCYT9rLCpZ6u2xWwP3iuwD2iwx6s06Rbd73TE2TvKLQMME
3MJF2THsN/FYcteGcDwUJ6E38mSDzB1Ddmhg4E8mScWX5LIbbR6hU/YgUEq4gJQDnWmtgpeEB4Ob
icMrPE0NAi4ZwJCXDT8N3Fdh0l44xpKUf9zzTcePDR30wBiX+vl9E89y8ILWHtfMnefjFbKJ5ksg
t7SogQOvzXfSLoaqw7w+e1PoxEJ/hqL0W8qMsa61hrpaq5D2EOs6IEsIInZuk6JQWQltSOZlF3+I
n65PG/H61ILwngQDDnyJzfVdX2iUEIIo9bUQn+48ayD3hr/0gOluod6GU7gHO6MUzwNX7lg+ryIb
uKFc4FjKr8u6l7te7lihns2R6Dkggw81GJ0xCkxsivh0LQ3VkJM9qgsHZNS+3mamYmeQdpNm5l+V
rLTVCkPs/wMrV9+SKS2HjttVeL/jUJP2BBgp4ZgpyxgGBowfakMVFEXB0YU/tCIwL5UDE80dd56s
ro+6H88tv9wjfRHTbcZnJpNPltb63woN6i4fsODHxsE8YB1xSoXAmk9USAJOLsIzWTPn2WXfTX8M
nk+ExObOi9/2QJk+4IHOSMD5A84mEWe2P7HF0qPuWotAt2lum766wvautAw5pWTKMsz5B/4kHZRI
rAT6p9alhc0grxzurKi9oujqmF35aXKlPFX6CW6h73bev8YMD0GsBrpkIDGTfk8Qm8BpZMiMELxr
0wS3IlN/923PUfquw74Wh9cyXyVyNmg7ryWVqK2JZngtedxhk3d8sbLwIuB6C+Pf+6xoQMKN3ru7
Sr0QLcQVwk02+kTQ3wLQIsasq+nrO8SinRbEpY0XyI1r5dNNQwZ2WWPr773dOJO4so5mheOv6JU0
jEupHge9LZ+Qv7t5c3tRq3RXJY+/tl3HDQDYf5M/bzDkgUR/S/Z+VwisQ/TgxkxsuPcWNoH7oUGM
Ht/sEtDUcvCQRCjogE1T49blQJlWiimzIZ9Fh7BNkNrDO1LMQBXKwd8WBFD+nout/RPJV2vldjpN
WRlvk6vx18DGq57RIesfQ1BuCRjK9bUdSxAI8pQrDHmJXDyOY1IJO5ZWrqtgURih9fx4itnCuEVB
TfWdoDzg2VkR0HSaMu9HOrJc3PDkFBJzO6biezB+zlwKX0L9DbL86871+TsMH8706anm6gOSBDl3
psJjRoXlOtVPBSwuezlnkOLEahaEXHORCdPXXfiaoQZJ5Wd824Tce0DnfhQijcpk2e9ERkW29ke2
VAFIPJAgKF9qpsH1YNbsuTUH58ORt9NiSEVVoFnFCZ/mLch8QV1jbpgvZoG1oLtCXKR5t3ZstduH
zNyOZV5tNYGDsJUPA14Z1DEz6yOpoN3KLky/a6B/b4aBHnnAEZkPP7Cu5tTqSSQjrL/IxtsCn0CP
fbB8+s5gJXhtVG7JJ9yUZm0lKa8z5oLJecOYRSMM7H8YpYNvwyJ5irxIdPSbBXwEEvYf7v9mo9GJ
ZkJQI2wwJoOVxE8AeZPZwFgVAV+tjIfWn3j70yTfjjNhrlBdQvGNfGlZXFOPqoEmPheioecCUWFS
cMeR2mvoHRB8dYbShyLl3zH7MugJEQ8YanwixrYo+f+SvQNeV3jbvpt8CgGljP8liNuIih57zAsE
rAmhChgxE5sBdZdE9GaqYnvZD8UajlmkLr98w7wJr9RO7IhF+g3EuCBn8cmMwOOJPJde245bhz8+
dZyAJg5Ij4QFzgWiIl6VVOQ6z734XpbJbkWKkhGJqyTmNdzTLnHppx3r4DX0/y7YUmTde3P5Jw3i
fN9xkfiS1g5O1mkEn0QMOOBGtCPll37odn4ATEyglPFkOmitaaJkwIyVHTqrultF5kOM7cMhnmft
mQLJ2a9fHP4c1RSwFti4DWT4O7rbNfW+HO14DIHa1fgA7zvKV2KxXupTZfej8n01DyH1nvrf4WRq
LZtY7djgec95J9EyH+LP0NJDzFBkAyQIW4lNWQu4yISMTbrR1snwxVwP6kSDy2LOE5U9uD520spn
ZoPaWa7ET7shNFKYjZ0yhdv+7EqNFN54qmgoOf9zWh3gwO7khtLJRJY37iTMAgK4PQB1Mz3dZwB7
Y5XJ64BzBdGHvRP7psviUNvoMn2Hi9uhH5zaX+0eC4nYbc2enRL4AoLiAB/KioY/PYQybGAMMVVj
K8vnORC9bfIdWPvGxkIlAXsTohKTTfZZifCN/QpjFulSyCpTJmpoOOdARJgMY9ZwsPjGOot3iqSQ
mNiWQ/MBfQ/eFpCBJZ6EkKQGX+Iv4T9s3XmEI41cPrsjHK9zOqYbGEYbP2BbwjTXqBSaO66DdHqV
KSQ6+cL+KzRH+cV7eNR29EI0NmObSCufNRikFCakA7GXEJKz4oUNnBx2VSTwg+kTDjqj7PoHbqFw
dDhknkIFAeG15sSHlLJ4KOGOcfPCTJpm4YGjZpRdVAovpH7E/E8LCVvNVkumfUJmdy4+uK4pSda7
D7JvB55wJfwTg3U/i2gKAvC08JZS9bJlExjhyWViGW8RFdKmNfH6W447nlfsB70dNARAi1W9FKrG
LWLJA2n5M1j6HqZC1c56NAcM5oYwkQz3/bj+CN89sn2gzPBVFzIwgr8Ckg9BrLtLtfoev+V0kfjI
mrns+lOkuMNCx2nLwkHwQrBfDGKwE0YlbQuJkbNF2V/91xjnI5GNQD+BIYebLDgo9s5+hDFhttkw
/1NLy9xEe8aBklKpCIC+QyCb/2p1QEPHWRwYmkL13dfzBJdcBXF3hn0oA1osU+CUTWefy6k47NEh
zUCfyPipNLfhqYm8jc37T1ZLxBp3e927sO6dM79srOURNQ9yy8lH+uZKTTJC8Nm9mIqbGoYydrWz
apW356mFU6zYxkCvlbgL1ZvRBwRgbT87GUHvsSFkI9TTlDTOE8GdV4RXCvIETRd5lmkPjzuDePrh
UKt7nx16g76wxfpsCZCvwuCslz5z3jFDDAWKAjid0E95ysB88HYp0WZJw5wwDCNtQ0gQMSeCPIPX
/wOCvy2mM3pAuGhCSA9YiPjCOsFEJX5hnvb0WXIwB5M3HLWHs2Gs44AKlyYddB7Zg7EVJmO1rWGb
aJuMKbq9JRt+Au6Oucl9GJ1QeEYSaODMUWHguVKRq63sXsb2SPyJgqTuElvajOWjCWAxJP2GIFF9
5aPAeNFKHyN5RRGRL0JxVjdbTpMAdJsvIl8HbsGQ9Vlg1MJ+6Tjy7Y10wt/KfUuWwKT0yYKZqgNc
OhDTfNihXAU3daaoXpYnx9qBWDBIqh46kcmDMlJCYJ5BqBQEgV5Tv0OPomOHg7RXdII3S/skvkTc
gB32mnTPlzelzaVBwQDZ7x8101UzFq9vg7zB0AUS2Nvx2tvMqph2e8fqgYKwx3IRge5Pl3eCLFWR
79+CoWKFOuKjCsr3ctOeFtITMdctgjxmaAKEeU7y+tFqjVuLokdb3kGf0i5LmLfbv5EX62gRMKg7
6lU+3nkRxxGit0y8af+c69PrMhJKH8A3B7eNrYp3MLWlinlQHUryFgje5hVsmukZsbZGjEKYKyJL
pRgH2Matocn/O38mWBd5zgTZFcV1yyRL8/0zXiC4peH9C7kAjjb4aGEf/o+0gGVMovZxHjYkNbi8
1YHNGABi6GOgcwnNz90uXtlCKIxtzZfuD9AfYDhqayqXhO/X07J5I62RoETgxjdYs23fxXFkBOP7
5xwp2wxLBFVJVd96He6ySXCyb5Sg8qPMO1BDy3dpfoIbi/Yl7/lCw+7wwp2fof2Uspws45rAlZXG
hWjbIr6D2UWlsQq68Uw2VC+ZnyLpZOnAfyygG3lqy1fWJ2kksDWyzqxEiP4L7ycouUw+2g37GRIQ
cqTU6rgTnYPHRFrrSuyi2kliaOwZ2105VB5oo/HHaT9L1kTQ/N6shN3ejzu83BAG0xZqDah9jLQI
duGrJaTFWH741U/ZwBaJQMuUYBPIdGBUFHXUbgegedeo86L0aPkcCNESpItiE6lpYKNud2zQ3ma3
tonR5dDdwrm0ZDroDEgzN9IXV6geyAkWLjXrQBW94yBZFOYOV+AacuoC+b69l8WlF1qXu7BGZp5J
Ye89aY0NZsIQzFFVoTA7+tQqLBZxfONZEx3OsphnB1bjlEgIZI3whJYMD68JC5gNW8+pac/ahcME
NWxwRH4A4syO5yre0p0mInAkCTj4FX9Y6kgDhYF7xtKUlCPFs8Gxbp+Nh2rykyT/SF1RWU4GXFPq
MUoGCcvQquOQFitwqWzw31jd3/EY6qzpGn30sm7nKYRGJBwx2eBkHhy/0itjG5N8rJaBX9R3qC2m
HWq2Tu4vUK7hr8ExnPTy/AXkIGYZipVqLrYqWhc0o0LMrlVnr4aazb6w5LiNuxqelzTrkk3r2uY8
ExjkN2BS4Zc5m0BodHIYhYWG5c7QgXB/teRfuqACf/BsAQ/baI4xp3LSFWDS7Hl7YY4IgwuHbanv
5uckH8euh5srSsH8FDmZq5+Iroq4imFV0074daHDVmYVJLFG+M++P5RRGDpST8c0tuaU1aD+lWFX
JPwVERuHd450S9rHlYxQ8Mf9Gc1NAmEEi8sGDIo5JSCphUr0zkBlQwn0wDw67ZH9aJxj9XYg+YeQ
FbwWO0DsaNxqKTC7OGANkDX+6cH7F+8Dr/D17I2qe1yNjYU4nj7LxtJl1ntmQoWDD0VXvEMp6K8B
r5kj/lhkYPND15sUNDTwdb86ORkOWM31izC3FvAJNLNefiwKGB6wcfd1tvz1oY0AMeMnrfanhKud
xKDMbUV66tqeaKMoHTPN0jaMEwGGrlHMJvMjKf+9Zjufh6v405QjSUNxcaD2GOq5OiMXeaM0uVHV
1dvDKANEkGE5JEkTKM66oj1DMvcB57WbSal5riwhJ8lArWpQ0pjeQEXtBTEZ04U+Gk7EIw2fW3CQ
sPsrc4Qm0VY2GcbCNLd3OGpRRIDMJq6oSFQgsgqXJyNPI2BdX3GOy6gcyLTFPn8p1NoUqvzhMszT
c62r0527Q3QJxBCitlYi3p9BQntGp3hdVzgqaaNio2fhwcoJKd5CZCyvyyMj7+1S9nn8W8QEK4tI
Zb5QVwhtd2kGXkEaemJoFcBKyuUAsprbosEyUVIysGW5qSC8dMLbObf0Ynfd+gMqhn2DfrORhvoC
BPEzERwUWPt6TEGgkBZHwLKrj7hDI5VNJqDbGez+DQHU2H5KQgMk+b5SzgxDmj4WLxQHenXkjEpC
WRIU+kV2pVPlY1Sl/s1SZYDvddr9Np/Nq7+CM0dodprfS2L8yCV5Y4SWZVEn6UDFMmDCn1JrO7HN
ET8HPzCeS/iU/ijVGXf8Vvz+9E0fbkqvSPmMINC3kmOG8s14Fj1lBaYC1Wthggmy4mnIyLzuWBSX
n0CrR22qvWTEPKMhJZSGAEPrLaJ6pPti2dYXE5oRN3+nUkhgIIIebI1OsJtW4mjRqxAE1mAs969n
AvbMvtsW5gy7JzxCQqb9IkPuk+XLvNtXtONjT9SHDe6dk9ZrD5FxUg0GX/SFh5l8GHaLfgNVMVb/
LNwuMBFK77GNw8ZH732G7OmZMGqcozmcuCBYhdWXiVUs94AwcS8GbHl2Np0egwylzksdZ+diac1G
/81qiHKcFtT0GALUE4VflvFGK3yl/6i1drmaQWzZkUjb1zfBGR4PhEcNZtypHtCzOevNbzXqmtsY
ynd5BI6evzMtIfR6y614HrJ2fPJN5kUN6D7JIsU15Gw4POXQIoCQKzM7nuoUNA98Sk+IPABQT1Hs
tjpjhDkUYh9UjKF40bpCNaG+Ge4g3urn0JTKjWRKn/qALEBU9EXoOv53Xunmu9pn9otE80QHTu27
v2pBP6I4bjNFYRD2LFcKDsNVzQWrHh2PPcdBHbdP9N9Ae+Gx8LwV34NEqRv5Qd/EnBDu8glbCj4O
fEPWkvaU8UVz6Sy5xdCxBkpx+sQtEWKwHntcjTIJRx3k8pY9Vgt/AqQjvVxP50MkxAOnP9h8f8ne
xnFQp/AZdIAcDT+eMFkapdAdZcz07QGMdLNtCbtQOFkJgSuUvINWaqQtgNv5qElncznW+x+Q5583
Ur2safwwOPfcgwZyVTOHT3ox9fy7zHTwqTz/IcpWliuL57n6Gb/2MRnOigXC1jV6Gl5pqPKYBma3
ja/Gb6luLp+F9WlZxkX7a76SWbdoDJ9n87L8iOqUUsDTm0vuL7msINqoKc3UTfKljXMfhy/i0hv7
8edlh01iZdfIfc4WDg9qTvkGF2TPlUwUXAp7rriSKxXqGGRLfokMketPWmZFa45t9jXaxQtLGWOS
U4erHaD9phrvMQCuOsPyIRl20MJ2bTZLEzkldEDyNfdeLUkTkGIlRqR667+yGolKimka0mjUTlKq
PuEeVwoUrIZmACH3ogRCmpfBgDcjnRbioBehwxqESONfa6AusDQGylbEU3iCkiferuRqG6BDVIa3
cdSgjlvmGbF+AYgUQICRidknYnBH3iojdwkrYMpnieZZefeK2UrwobJ8iiTj4KqMim4qleTSSAwh
bQW2PCDbaZW1LCThI3tDfZEyUd0F+bsV6qaMtVhVC9aoSeAUHqjum7GKqoq345UvDe+LJBvkOcyJ
LxnARuZXPFkSM4qwiWAqHmLid4U09+JVSuloy1sw2vZZxAP+7ZavrHO7/VQxWEDUdfRH1I0nNXWk
M74azILzxt40YuWW2+XFTpq5zlwb7d7Usbj+6gnDcmdVBGMTdS4WCD9wFZKniPdHjGzJbnV+RYGC
MS29aifbAym3q+y4qbW/8qhnWqtKElUlU+8rzwXPmk26TyzINCaRTIpw46p7NzpAk4zFX7oqbLez
Pmn1kekUp+l/GtQ8N6DfWBOdrpSSiz0dEwXOzSzam029UN+7NDjF1t2F5iyL+kZRyopI3sEj/iPE
iFanGr92yQbIc9OYp/K8wuNMiHp+M3Q2mJHjjXqsNm/nla8Ls4+Z/6g1nd6RkmfEMQWaEGSotFDE
O7MiDZg9DOjnSsOUM59cD6Y+Ty1mocvMZHp7f1v7TUE9eoT9cYCoafK2MWXtM92+3guag9IW2N5F
xMjodnrwsA7gc8nip5e3agwkOdf7AHe8nqtlJo2f6Zd7uXwlF/2pj5u+Q/h1IhBcDZU0VkJ7KZYx
Apzq9oxV2j3QpJo2ydPnFebGi1+lUXMoYYaS/LW5S7ejJIMiRHCvnK/oS3Ril3zC3uBaFK+lWpzU
o7KeEP/QcU6Y0QL9GY6Ef4oOzbBBwOAaTyXA+IQoc2JnwaEg7zVLdv2xDbtiDM1+gBxoZj2ly7Pm
BohUz9DoUfHWU2fqQ9ZO4bBa9uN7zICOTVbpxb12+CMliTgJ538y4Be9rnXcIQUA5LH0+GskILVG
bvBhWpJqdiFo9IHposWEB1v7g06ArFKQtd6e+2wY+/iVvi0AqvvLJoG9N0TMBWu2CiEDgsW3kw9l
R0+jYXhfSw/FUvP1lGflRAI2tAtHeBDsDA5dSkitla40wELk4BYd0Zr2LY4WtmqNAuuX+0vZfNYB
G2LQBp4LyqwLrT2f3SwEQJtWEmiVUIpXXX12rG1f80uluOaSI3ITADnwlR4jfMZ5KkO7/MRiIfL/
9cvzmWYnhlj4Pv7l6zS/KZ/fPBpnbNVa9ZgKFpQ9sfz5gGG4iB2owtFyzX7HDTOFUBvdtDgWSKr+
yzRpWVceC3zVYlYYq3A/XkgiROyZRec738+YS1+KjUHYjFOzWc48/USj7mtCi5BXAwcX/O2fKfPI
Fj9KBalDEI3OXCXGc4sK6BBWveyOAkJQUrHBqohX14RzUSZCbNZHUnvdqh2dbSnlNRO2euJqXYaY
w4DApoqd/v8v+QoD0r7hlHnfLfu3lVwT0KXhNAJwm7v71kcFXDsvqNtmiUThuOjsxxcKXu+9oVjK
T2cLXaOsOGuQqO71G6XTYX03ddCT6fvQsdP/Y3+0T++46kuhcn3lM8eL2M1QDLjjIsYADpyKMuNv
tVla0vU6E8fP5FvQzHxqQs0/SPWbg9847LYjU7GfRLWb08K+/EV9waxv/b+o+qvcrJ/jbFZUx9+V
tMQL1fE0d6JWqIQY3wHkT77gCCg0W0lSES2hjeW/GWW16DUOkkW8eVdAW/38XGiojfYjcPafARSv
pQG0CFILbsHWeXdlT/F+O1Ofg81yFTjEkvBJ8rbRhom3j68rp6TGc1ovzYc8SU/DRnpLP8jxjavj
0PVB+wGWDQAM88k2mtEDH2I86N7VsGCV/YLzOZhXaAsadUbhZ3+0JIwabF2mT23FsoY4mx0gYaZS
S9gOWpR/mErBvHb0uIXe+2ZliALYGCIEv7iVT68zlgsmuRmOehOur3okiOMRMrM9pVp3AT0HRjLb
SFEk7uoiL7BYas0BGp0MfgwChxRub+zF8IPWVO4f1bWqNTYYwBQcKx7XZAHkwgAarqYiKA1BuI4O
ymLr/ApsytGmSmq8+tEFpxxfU2HmZsSjEtDJEgt+jC4kaATbMaI2hHLyKKPM6dgWFs9wiNAOLBsX
ok6mqW1b6vUQq5qmg36mFl2E0P+yAscNC5bUma4iNaAqO9bSoE3nEm8lByZjns0tkbhCbl+t/6A8
13Kve/45pPvgrtWVhb7xMcIO/vUMalk5a0WfjrVhSgPaAoomubS48JnTmc21f9bDCrIykgc1b970
eZfGIYVntoUKDdup49cbcg/Rk0JqICtYZcmWQxV7a1an4dQnfpQBJrlUZRqOALF+E6w/vjaD1bwu
KJZR+QJ0MX1uiWszqnr+KiO/akTt5zv82EuaYAwkJLUiNkdAnfuKTTAqOKumW0K7NzQ60M2MSuNA
lRSZjXkxKQxs1DvPXxKjNhP/haxRl9VLPa1V9+HVo2ocng/bTYkeGKZEz4KrElYusZUU/hDRSQFq
79o1v5gMd/ZsPv6orvj9nn3WwJb3yk3Hj7ghwqxyqTchzmEaw3WyiJ7mtsZJ8o2DqpQQE9ZQGFKG
atK7p1rs3fj7i0PVjfyvLVoVoYeW4UTdNOrkPjHAOdrpRMn+jjq6vGNmLcoJSRZ6VNVm0DCLvWcF
lJF0iVcPGteOnDjAhQUdVHc/vvHHbcXjilU3dla72Dh4WmvV0fstEqomsKpdQgwXgG6QyfWqqrwd
mbtHHBgcPsEBX0rHj1sn15rS4f83S/JpxQIKYzZUJgb9+2XclNHSlUIqBVIeXJU6XCg2+XpGVy5D
/SoE5CsUNHomNRCXH675JEQJsgd7RFchEHYoSC/f05oZYsKRZPmQf+fd2E0PWEwcvJ9y123+f4Fe
kPb4lTcPya3BkQomU4Hqc3ywMxqSqS48MTdGlD3/RZMNfu2ENKRgzd0J/IYx8PqUcDKpVVsbzKlX
Vqe6MgqXTHwoccNwXR5SA6P6smQdhX7F7k9/YyvqnRHKFcxIlVgap9bk7A9qnFpuCLlYLRpRGeS4
vNJphfvvfKP2AW0wscWl2tPdRp5h5gix5ugB64Jcmyk06b8EsE5J6aNDXFNBJ1QhzGZR5v637WKQ
Owjws73phEOl7fIqs3xqrxYydxQPAg+bq3ooSgR+6XEkrctGWFRqpd9Zwk0hd1oTGKQhpvNUyBJs
LwKk00ZagMfbhyAlN9BqtSkuWFw67M6vo7rJq7Vci+krKznVgchh1+IzNT0bIY5dmAxqPN0XzkvS
otaIQmpSgzPq273k2rMfWLVshFVbkBX6hsASLc9WFVnTMQAPPnnRYyEcufJF+AHmiE4VkjPVnHfH
wIWNX3RNXTyR/qG28gi4IhxmVzY5B/I31Ct1sEQyd0ukFzfRKE2kgirX6Sh/JV8Wj9maaS5zYZj7
QtN5hrfL3yPa+3KtVr6Zw/faB8EKhv0rttZhlEdgqloma6CLQGPjcBaBOBBYDZMMOmxX7vbTbAXC
nb28m+jinqxDLxe0KwbLnwJnMMYhiE9kXxSgtML+K/gB+dsOCaqEdvev/yZY+XlC10u3854w55Oj
NeC3pWXeB7L8AyaAG8x95HgRCuPmKTC3LzpF4e7cRSIgFjnIMy8tIyCz20/T4OcCeXXA4JMfscvc
DrME13r0eIje3EAY71Ixp40GdrAEXb4zww1w5OwVNwlzMLNPWqcLsL4rg91owdZ2mUpYoSfDz3Mu
wMMn3KVnTIsz8LyrkmqH0gB+YF+u5lWAgaqlpJAYQcWIgDmBpO7QnyYButfGZnWvNPERlmjjzApu
5PLWUbtR7+RyTPVUZJKoGm3UxdfAVTHYRy9b4NQ+VzkXUldcKYNID6eI/FCtCth33nGmKI4j2qIa
GnRM1JoMb6Tu6Co7W1qN/ScwnGTxog1njHtuicR2tO6/Al/aoJCQuFtQrwkHLpX40H7996mK/GTL
KMRtL+5wN4+Y+pZ9S49qo4JXtwjZTLDMMBQ4tyDBUu8kXJwOKTyWRQo9wIaG8KL7Wt5VD/W1pIGv
osnXbKTK4If84Nm1UkSJIdebru7+ROk4BmcF7CC7yLjQ2LSz8O43l8zDJRo/ydXu1zTmBCOjcPD9
FgRvpwBcxdx/VH6sQtotrGzf9eb7NpWyyldsq6t5uk1PsInnWPjaYBI9K1Lri9FaXY6/W+TffBfx
Z9r6NCOanXE5EmfauSegN+6kF+iGd9WAOViGqlxqOmijKhuz6+C4ZqKGx9P6q1jpm+3LUMfaXEVw
/QQJzIVFbW5MAt3shhdcelyWOQ14olKnO4Ka5PvCOZDI360C/NP+kdi5s9GYY5BLVMAD13wIHecT
8n7sMEAmdw133irh+q2YA9iHvfk6XkBTpd0HDGYWF1Yv659eEeJttaF1RSVBC4bO4yU2X6yfoPlW
11J+Wih53TLcD9DmkxkX9/Ib8grjaj4msJEZDqXyn7FlVQgXqK8kpcxkaYmQPRyCgajpHVv1iRQa
4mAO0pvGkJnt8rO3pa2ozkT6o7kXeigczyVpU7fKMolnkBYNQ86hZ849e124MRJ0pdFE5Tn8c3gH
NjBAreAxsWJE9MAAkqSgfffhALMXssgfGz0GBB/CWyADsuVK4zlEGuF9GlMyybXbtK8SWRH/f37M
8YhRKCrd5v9tD12xvzHJ3eEa+WNk68NBT08yGaauEF6h/bYXYaRBV4WOH0fynUzATHygvLBOfOIY
aQTSQ1KFpZLLKOqDjyBuqA56qMIMnZ/nko1kEbwoEdIB4gbXxoZbSjdeQDpqjXOzO8knsWKUEgNO
m3TuSgYrE1+5lk0fyeHcqaawiK8SUpLnG22xDvpL1BiJd/irWjUHO5RAoE2e8x2TOQYTThz18xXt
osidG/ATAO85L4TSoWllI8R6ef3a8YP5/gyaXe9OR5Ff/BzQXULNpaFJjCnyKKCguRXAxNePjJV/
BpRvOpciY+9LpXEOFB0ugoXMRnld82mqZ1Pcqr1PBg2n792GKWRHXDg0reAS3M+hY5N9tA7eVS39
Gk/4YxP6xCzncfkhEqeK451E/iVk/mkExi21FEXmRQNQZ5/j7ZOACqas4V2NakAgVHsUbKBJEbOn
nPJeMEC9fSKJYbmcr9h9Nvgg26IWA1Qh8Ch5rAPaEQ33LKT3njLJTC/RHtPlxbR4PbnnTTYzJVRa
saEuOLOzr5UkRMmBQ5VTSRg/9bTIKK8BWJ4ahZke/d1hcsmr464V9YdafkEkr3zZARb3yRg1H7TG
zNoexjoZR7cGoFRHGdA81n3vHaQkKOh+abdOrtCAB9ELcHqtJevgNwtEw5ufR/RzOUtSNFVk9NpS
5dcUnFUuO1bibnaw2WpwlkxHYZm179CIxkpuOuioBn1xMIWdVAVEfNI5Zxc5cb31xZlOKDuY2WzT
2lQagk7W/0zoc4AY8LIsDrBw/vo+CuszPIi9fxDHGWkTdWKA8uSf0f4rbeMWRMNJbnBhfVu+9Vy/
tchBwz/gtPSMFNdnssdBkUy3S6OKuoKysQTosAJla+66QH0WGp22LBQdd1gLWWXZ6t304ICvwq4V
URmeVssRu4s2IMwurAMDkC+47SR05V7w8KaGONpaCoU7OgP0Xu1hKXMS10Y37A0j9JFZZXIc/vkb
39PlKZI68f41p8s/xvUWdWVyq6gf6usOGKslYYoV5FlgfQq2BW+ScVtnjVDm7dBRJH7BHMMZqCWF
IDMq+hW1+Zn6SVrHQMuB0y3cb+/Nxy++XPT4wssyV82cr4GYmyMumNxqxY8kG1TZKC7sFBfe6M4g
EIDeDGyRWqLxx/YOYJeMxViWIyBiQX22uhZlZ/sQeDOhCOFf+ULZUGMk4YGGV44KvZhVVYp4UKBY
Yd6hp5nRVXxQNcBV9pT9/MQsg/2F+WTXFSFubqrNl9dsrPkTcew/PY0TL+bcPKs84vOrSXGBHFt8
+cMu0MUqYZ3hisuqrcrZ1jAgfV83D/0KxFE3NgS5004Vjah7n+og7V6ADKAv9oscu1RZQhWUmtyy
sr7P6E8PVnGRHmIfab0Njowi1zrpVZ6NUJsu2uWM1o1x0tp+qDZhZTNoOfXTYGFcmOOrmjC1HGXZ
Se54wU94iwGrU04dfrajxPwbCK0/AnwW8PPbokeuHDyjoBCR6M2086JQpL1gdRsVEUQdl8k2upJD
bjIB+6kQcpVjh5uZ1k+W12Z6lmG6XhmvU6VrjwHZLFmYk513crIr2J0HlYCKcieuWDubQ90CKR3t
NIxPOYEXJfpw3USKLoJJmjXjxYJqC46SEwvRZSmECH9uInBYICDvNHkvjgGxsYaJn/og1e+c15ZN
WJkcWn5/12aFAV8GFuo5Cue8JNM/Hscw/Dj2WE7rf1JrK0Bmc2P9VwCGX3h0zv+x5qqzwJYodruX
zxA7tQ9PhITKMQwl2iW2L7XnspEp7B9mFkNfPF2jjjBzoQIR0DxAks9Rt2VqwAL9crHZE598iVS7
XWVZ8GF/dnRZ9AlXlh/kKDkOCox2AY11g8ItAQm9IwKsli/XvVJAD3YeWbsgFVvJ4MF6tc8Pifqb
LPNNdVHAN8Bk6nEaUJyirYawBjt8YKakZaKyNUN/Nig+rVU9zwzDK/45FNOPTi2hOkJRmGe8NiSL
q95zjpy1Q855TFe0W6EaHFHtQ1y9dduqfFlDxrkWmGicQehSXemaVyn1bKU/7vBeyAqyp/FAnsbk
r2syAA4ivokpF6HwKwjsh44kes1+PeOQQ/r5p/QhY9fO86bF+fG8sKby3ktgExuPbqGx7C/nUGXB
8mC3gj4tV3mcKC7E/gXJ5xnAZbuJpycUUkEH+i6H8LYmmwJ+rozedjpvgd7MHcrQC2qdpAg7R9o5
y36mf+eTveTrsaYnb/gLnovAh/7S4TR+oDttgDeusRKKDGhF4zvslmfmHSNQm0LZ9PguPg6iXr0y
/3q5bLDdkci2bIXQeNO+bedBJI4wAC0d6z+AoMKnGdsNHa4ZRt967HKstrTda0A2gJrwS8PC2UEA
SgdFlmlB1eiBf0IXxGUYjGQI/YQTBpF8Id0f5Qd0D4N+xXjx4rpkv/dI2r8gG9dLD36ZUAgDbjxU
DdOW+v2REE76T9qcqyI7CR+3+h3o9dQkXwpurha8nJtyODxp8jtksVPQ/choNQ7aKJAFI+ypTsTY
cqKcL+1tzkC5Mm0XLnCZLhjQoCrJ3E5HUfRKKdyXH1Ptm+VsYAemOKFvOUD5vJSWUoh56XwzruLo
MXWj3q78W0G9a1+NqZkkToA/1KJ0PrgQ8V50i4A5xu1J/zy7g+QCJhD5RvSL5zzmmOfvkC/3tzER
bFhGlVZzFXDjLh15B2tpxOYdgIsSSzq7SflksTTxmLuCTtu+f2G5V77Pd8SkFMa5nK4j35uxgdkO
Lsly3mum2ETk1xZdxKUOhEp1wkJf0LH7n5SJa6Lk39LjM+rTyM5/QqKbpI9HPGRWzzvlG2uVZPAI
z5g2JPSzRaI4fA+X2x3ZNqwwE1xJeSkYCyiOLDJtgZ+ahJclQFlbbGomDQ3Mt1P1Fhc0hhh6/6rx
a9v0jfx9HKoazGbAeRNqdwE/gx2DVdEOd1t2inJdqrUUVcAq+oRNtZIK1YpYMZ6qbRb1HBYuAurl
WfF0pg/EuRwX3xguzcd0UvnTGWkbHF3zRaNandF5JaLBl9qm2pZYpMte+62LvY4EcYLHJr3KDAUI
QPmYrkC0i8QHSQ80rWJIjN2ML6Z+E63lHgVdBYBhhkabVqzgg/LQSxJIv8s1cRIpLNoBKupt+3J9
3myUFPAbjCiPpF8SgTZDaPSOIDJGb8TePhXw3xxIfXyxzvQX/EgPw69Qjlk3x5rdDaIfo6jhiVlj
rSgjPtC6fJZ82msry6VtQS67oa/NucEhZtkkiVruoDZLkEY0XV9dTge4+6azROrxhlZGz5icju4x
HRuRbTjcnz9oKHX3+LbaO/CFlnsHsftr54OTVmacM7A+q9Y9t2qiMRkr8EQtIUrG5X+ESL8rM1uu
xWVZ2x2OYX5jO7/M7hw9EjaTN/+gxlu4aPXivpXuuGcIJnxsKPDCrLBNNSp36Cw3QTkwNjx4oaEK
3cJWp561Bbg84oQVgVntDgCj5dcR0laRGCgbSmg5m467HqJtfs5NMcXHtjiId9uIXysDhUm0373d
VAm22utw3KjuzlMsGc1B0BwNrKAT33kv8/jZSELKAYA4uAsHYWCkACaALV90eIedT4bG9Owb772U
n9SbrX4BKZJGXwapj9+v7NFLaNl6eqTrSad/ztDU4y5GCiqT7rF00aUFwcjkqNY4kspjYccK6rUW
1IA1MWYJVfOAJq88Q5Dt9NPFw0uNAVnKgJf8DrUwH39Xi30riqilsjJMIy1H72C4d3CptBlIVyFd
76fMXSggADroD7lIxGf9/Jf0e80WgLmeaDncRfdZa2BpxJkyQhtLXjbymDj+tw3lWFaFYvYgE1tM
lAMcBlAir2r7a7huamX2nTTtz/CHEaiWSwRncGQ7POaxKcQ7DUAO+ZffEQyrkBemPWnzLj8IskAe
PJ97uWqg8zBinmoT8xdkIRiFpwo3WEWRjJafuoYydhw8ik5jCywwXYs8S243h9Ggj6cXpIwDqUhN
iiRRFo8H2uajn+hoXQ3wa5D4EDIFnf5Siu2MnMES3lbJJSYKAwqLIvppZgCJNx379YjFa4qMjtJH
800sEKnERmMYStd6tk2KngebD7uWYqQTaBjneXmDi2CA6zulgrXWvDqfXwwraIHvYaQ5bfvIWVgh
GchdjdqJdazRiMs3VEA6ojeZjlN/sDfyWcHqK3bZjV4nTcE6iItbZ6fYwYlQvHXyVXbbL/zZj+bW
7ELMova44DSXDlfstA0eyOr8PXXuohMyAmpiv6Lpc7FhxYKLQ0GT+rrbNIWtGiS0M+F576TLU2Hw
McjXrHJoS1jMF4ujALcNvHTJjjrK8UXyz2KxDsEc0gZ8HyVLZOaFJicN09eTu0hXzmxTGkDHqfAL
TjFDdlaSPwnjNi/JrzetOCTwG4Fg9tS74r/EWnMod0gJUD5Mm/lezuxDwWfhlR+GbNbBbBRaLEA3
rTn9HthNjqrTKqh8Ot6pMCkI8DQPQNzaOoPxz0nqxAG217kp/eEzoRbrXYaOTQnfTdZag+sybDbU
GNxyvHqtSUuS5xFQ/rZY+o2+yzyVDHyUIVSqUxIydfZDAJZ5+ITkHlduTsAL0UX8xXPsEwm7VtqG
PFXhn18VCF1GF2LJ/EpRNcjKa63XfDbjVxiC2XzJdmeuuItM9vSa3+5lyJ51siG0e7HoCJn4IQOg
+wnoLMecHg+m7AmY6yRpcPp3FSasW383KUou9eZuJjMHbSeAZxX6BCOE/bmLVjaXYLT5XyeLHINm
+LmIBxpl8U35i6yUlORo57XGDRKpVKn18NTXxy5JeGiEGc/wuZGQ0z5DqRj62qGFsEyQ0lkzb86l
jPM6vSOHkC0MBouzYGQwozoIwn1xdDK+AVLI8sAkoEYHDnS9RygNaKbmPCTEQy56hc5pBQouijF2
jpNYCi0Dkm3XEtc5TOMby6TmuYF1itOIC0BOLCjKeEmavo22l7o1jYXXkQCY3y+iKw9b69SL7BIh
OgIaD0yGNf/WZKCLfvDuBeZLvYORBN1wdzpvNBTw2Pxv5wiHU0aeZgAitpFfCmcnN933Or8Qd+eB
KHdYMLUe7p27Uutin3rLQXUKkRZdWIJR+GinLp7LAO6ItzzvFyZSxUhcqunAl+dA0hopZ5Tr+641
fvo/oF3Uaa9rcuP5xNlCfFnlUyZ3vhfwr5DDWIA5gB3BvBcdzRItXB7KQqEnzDsBzrS+ZQscQpAF
AVviSpsWpU4Nw9T11Fq4l2r4MME8FaWHhiLMlHQ3fqfm6y6AyLYN7KlPuZyrGJvUV8ZAE763OJOV
NxpAQZh+bTkkiOyyUWjy5kr2fY7MF1u8vRsYq2WkMQ2VYXWNnopR0te6W1uqdyj32o7NhDplTUJX
ILrKoT2jrTtsUWO7ip+TgIx4VfyHYZgHZ27Wn0dV92RUqDF6boTCsbQD4ZRJJp4KdtWmd8cWX5VS
HieOViv80YgpBBjWHpHBCibNX8Tpcx6XKC9ieT2TGSqJElrlI09UktHJH8d693JCgLrdLb+X/A/3
5lrdPtmZ2V3dKmuJo3fx5oqI70Oh2sRRJl5PEkSsnrpEjcSvfuydlt5Hgd/ftPHN6iYme71M2HzC
YLio3F1d5A4k7yzhFGDjrR6lrZxjcbspgr70Nw478bR2JtDEHEIpx/ySZegSAmz6SEcS4f9DGRBx
OyEle9blMx9tkm2vmDli4mbn+Maknct3G03boxm40FYsukC1uJmj92pFDA+keSou8OOAOu9wbU3H
rOytZSgoi/gpc4OVwadOB/EEBla+Xtm7r0ADoct1xe96CXfl0bCYtWF1D5+xPqZwKLeZ62xNeRwI
n2r4bsEcyi84stfQELLknhMgPDM0p3WgjnXGtlsoHeqMQmHpTiwjtEGEppMgRzx702ma0IMWjFQz
TfHe/a2ciIeWGXoRzszPW7V/46bdnQ5cY4zOLRbVgMTuotGXm8n8JT9TAQURPGj2E3V+N8RHm1SW
crPs0ll77YrhtOrqTDNUt0FJTNCeSH1a/bQmyvehPeKQpwk9cncAdQIBhOEwaKvnGG5O44nOR5lS
5jqI7S9drGwia6iuPl4bRp+p8H74msy52PVdeLZ0pO6bgQaW/pWGI3gsjVzTu0e5DkasX54q7J3m
An65eCLIuOgkoqISqwB+VtT3xoK6Xwm1um1bvukxw+zwdSn1G5HOCGXVRIXiL0vfUEB8Qaq6lwpf
VEDWaw9lwfYLeKQjbFEDAbs4xG+1XGpQvM2v6ro7D48FiV3QcK4o91yNcUG+Nf8jhWb67xYej6Eg
Uw9zfDK0jsOKccZRXZx0TdB0rhQMzYg7m0I0Jezh1SD2o0HVgjD5M8o/YjMBYHB2CRBgQX++6Nmo
n/vWcbCE49DNea6HAoRUPnO+/8rbwxWUOUfa/uEtw7jbob/Fjz+WX6tIAoSf3Ha3ZWbOWVi8nlcw
DEAeI8zs562WONgkqI7hDWtp4+y3oItMsz6wE/DUvaW+UaILsGIiWWzypLh1VE9sGwXukpOX/GrU
ioAipwI3wyWuS8h7gaOVJCeLb8QuYUpGxJZsSLyAuJMtnMFZLEukhACClBZ6k5Wxewn+EJRuc7Ez
fAoB52kUU+Z1dhN1BynF0fLO2anyMpeFGeFCMsOgRzKx2yGT6uENcBHDNeNfIuZVLHFiV5lh4qDf
iv0TyAN91gelDnF7suKgfYMce//u2ezKOUmcQAWXoGMoJfUXXAyGj/DTj9xtVmEpUyc+mZsU0AtO
SpCR+B0E7TlzARsV+FtYwTnyPBC4mxqi1LaDnWQP2RCRk4q3yz5KNX4o8ZenqCeEs97c9O0HMEs+
CyY8GPRNMzJ6CSrKx3LPGP3XBaB5ONqR+bb4KydgKd+7hHojBC8y78KodaURDZuw33/9hWtvOXzf
1HceTA1w9yokqh6SjeymfZ/XU+qqY+HOLKKu14eojVXgaQiVEbfVz+MEd0dQjbfiud7NgiQZxBMz
RaqvDaF8lrdyqK+fjU8sefYx6znObilyeZXmTv3TwMGKpWPaKVqucnMGelcLYNEk2RP9dcyPgFjl
7xgDcGbPqWRPTyBWAycO4YMbhn0U9xn/j6WRGC4JAi3nrnK7A8knJhqb5VNXSoPMkv9lFMXr0Xyy
5jC6Uru0LKNFp3bNffn1tiNB1ftBiJOHewd54ngOn+bw+DaWsyfHPmMnH3iDQU7Aaa4GMe50qXMp
HQGaLZ5Z87gE9uOsg40BMX109ecHRaUTUlRmnoFCXu34ZgP1x8AG/RmhUuwD/kjmv26A43TsWhNd
gqxuTay2thtPQ99f24weehfhFJ55vl1Bn00dxWoWs8yKb6ZOTfRNp3ownWuUxtsuOzFsVHJUAK9w
yHspU9dKWWc1a/o+65nW4jsjSPzkdAItjizVX1ouNCghh0SGcEKVI1t9tzHDxm7eJfjrLZefrncI
5kJsH0Z8sPLmWl2gwkRLGf9N+aYrObkKsMiWWFqeQ/GMbW3j8nMjCA+S43/i+8b9jAjA6XrZxJj7
G1Ps17S8Bp3fnc9NOBDFUPQUDwv0KXbNPfaclHLcpoa7cPN1y+FY0cZYoSqGS6o2lj0CF3Kmwlo9
yo8h0zTVeoKslni+zOiYBh2rUrmF75TGEVr3G0xOLAzKkI9FV0DFOJZdw7IPMZZZVo6GUHixF9eS
PVB1lIOTNNCy9gGWmhWi9P6iHPQdYLNRfpeXz1ysc+E9tOPBZ3zWFYnodOE7LVFPXxpbQTRs9riv
qnG/7lzqEHBJpAFqpHDvkxnB4ykF8Pz4P5YqvmDUqu4f7EjBLwewaDMLyqzxdVcK1UwmEo8OwPfY
uMlVXJkC6bsFtkvgttxyEttp/DTng3aqmnxljoUebypVov0qtXRaPFIAehxQg7VsGGQFy/VmAAJF
24aYZ51splRafVcmQTgFDsIl3Vhsl6/etJnvZ6ax4aVumNtD5UYCb+5jEsCfc9wwsTrwyTZB2kj7
Py7uERRPPttNCf0wALTmpipNfTvzQI017ugmEw5K+vA8voMmFXpLT/C+USuMLoA7bXxvwJVT9qf+
7wQusfzYcKpiGPkUg6Yc1RaSHxkMbyE90o+hBlFh5m0llq8A9e8+gmNEy9XvsSP5WrUmv5Uy7okB
RLbKCpvprn1uMOa3KXD2MiaLd0+d7v4/mVJ46e50nOzPlYyojvtset++mOpw/awVdoVWSF1YC75Y
jHadALMbnxdkY7JlTJVTUHVnf4LU5lp4MK49YjpKbVV3T/GhalP5yJDqVIzBdKaOHgbT3CZg9qzl
4p46wwBHMHYJJkPZ26ifk42Ci0baW+yHn79s+SSyurcQLgVp8hBkm9VzAlT2HMce1sXQaZP9aKR3
Pcbby4AMsqGC7X105VVHzIOrkGZWkRoRI9SqFnUiUi+f8ApJjx/eH6/qFq85eXw3la/nQtwC6gta
RLdVKj+jquMD4y9kSe+eTlYREt4f/tSzE5V11hX9N8IlFesCoVUq9MedTJPpKtr/+dlKrZNd3RkV
Qd/whNUXDxNZYL00sDDvhApmaqye/yRLC9lnHkFZMVaJIkadF1C6kV58ds6Ii8hsbp8LG6z+ux0d
Gk9XAzkqTynyH87EDaJOwBiSiA8xnbjlSnW2RKp4vLNNbqvAYlNCmY7oFR5fsqTPK+2Z+Ta9jCjV
q7COuW0JoW8paPK95uO4jw+c/4GagExuDtN8DPlGzGk162Mp/V/+Bt7WYThNHLwUI2v72hNGzaW1
p0kKQbilaL6hxslmMwmxUwEGhdiDbf3CRyXMjesjazp3RUkQI2zVCjZDZJ0dKJhIRVKoNxANw4lt
xbL4CtFzVviCEqNweNeWIGOWr/fLIIitD2i+RabLlSY90kbqmu3jS9tm4izuvvQ2keoqGfza6CVg
QKKDVUvBOZi1/ROAnzaS5rjESTwX2CE9Z00k2+yladXlwfDvWEJVdh/okYRFaOAsTKj6WiKjfEbL
yGGLMyc1c7bR3hItHPKXUMQdJpqll+kxOOMnwhFxUsnDuQ+k+u21ieQStWlIMrkjMl0oHbGYOqv7
M0seuGcABkWQbSBpukAUjJYVBL21etHvYQU18gmK8FufovaYLBD6YbXa6gx/QjWgX6LcOQ/+2Vaf
j7QuJ8TchxVaPWAM325qv3EgOscamgRbGTGzRBGapl6m/ceprcXXRQNwde75Ol2TiBDWo8X0Uwb3
04Zl3KY1rNLOjchviImGEGkSYE8c2VohlxB/CnqIi1y30GWeKs45NpOcLVDMrQVIq4luKoglPYKg
4GISTIaweg4BTu5L6EdopQ4xfcQHrvsssw+hMWMwxLN0cqdvhP54OfHQKwRg3+GHulWIfAEXwimJ
JaewJENdhVVM7T6u/fIFSxK/iJkzqSRKkgQRO7T81vWJGvOkc2U8ohclQFrg26FA+ANalidL+yod
LgnkK2fBGsPdR46xKeNVhbS4etWsRBLuv784W5xqFiATt/u9fnShx50GVRRvMY/qazxtjDcsvHi9
VXikfm3yQmj4WIezY5jts1k0aIWlluAbQYpEX7GzxliKT/Ajod8l8R8uZoyjABqAqtmL2r7DPSoh
axaYJ3BVWq+4rMasW74VMbd9dywc6GFKEsTmWftVorIsuMu8O1f41fixgo6Ws+rE5AT024huXbh2
i1wADVQLFBe7fbWKi0cXIIa32CWQNZe0DaoXlaNSQm33nsFKYi3YsU8RJbTSe67XoyskZAXINNDa
uWBoJOc6QvKaGpg1n9+cSlyfFeCI4gRTH9i+oC4O/7tTRIKIG6pnilla5T3XAEPx7sGc0MBdIxVr
k/k96mMcZqp+EgCUFVTpdCnhIpMvBCt0Smj2fCC9p3P/3+3XzWiMPEG7b3501Oe1KblbzkFSQ5/9
e2OKQOyTg9D89iRsXkxF9zPy8Uq5nOXYjtjxVuQ4sS3fus2qNSilqP8WNsOqd9VQjFYhcZ3pZxPn
RL0oZpLW+AgnyZLYtjcphFRfBvZFczQk2wDet3Peb91qDYnsejvZWWjRmtgkH6XYPO8PUm8KA/Yj
erc6HxaTB8YBbNaBX521H7O9Kq+CXhSnGus/CZGxa7uS8WX3P9BoG5wugAuOuMqHenLSrIqFXSxd
2UgARisrJRZyYrB+p6u9fzSm3itjA3LU0ZFBg0HW0efsgDeyVhtyOzpBC5PDV+mHjbjWirT+ZvJo
9crSFZcIkKoFI/dIA9iEt7zCjmNNl0hybwwziHwv5nzzHbJi4CpKC1Hg76TvnlRocKv3w+xvotKv
BfYeuHhS/2b+6G71H76AqqxgsEg//P3EBC02FnkSv5S+ghH0QWEAlRLVZNNwu+RDagosA7b9A4j5
vEHU7iLsIouEAs9mFWtpO3JkVKtpBsEG64e+5HgmeQhaC8fXD2NqFJhtF0SaGsJL2rSGXgSScuB4
NX4qHONg3IGUZqn6rNW7fhHte8meB2pbwRNEMOAYBY9H2ANihNssRZCKaUxbsqOym1o5q9jLoeLN
kNLsxCOm6h77cRI88YKrFPl0gXPkWPmDseq5zMJixFxeD+CbhZzdGKPzed9FiRlSHQWCmxPFDqAA
Bcl6ceT9Zan1TkfrwMRpA8i14cQ06Tk+PO0IMdWUG0WeO+S0pmT9Txo94uz1sRSErWWYuLqM8r4o
oWtwhsvglJJ/qgcixbiHchgDS4gxdI0slr/hEZ26vSKazmSuN+K6XUgOuyTGSmR+X4dVB0fj4Ejw
SsDk2NsBQ/+TbOxpTGBc50t/SkYOXW2W87aL50gy/6AZ0P384lRW53oNysO0ejL1vFgxhkcbyb+g
RZ3s5ZgaW+u3TiOXtK9Vhp5PykMf6+6BIie9dfR+5Up39+FhUCIJJ1BQqfD9Zq8XB4y4LrpRXOGR
umbxnG9O1H+sZyY/2h6cCRTHtK4wLv0YmgQt+1cDc9vIcJf8Gjl26kVrFEKgGBllXDZNqKkX7dvE
9XMP45dfU9BjC8G9wyFzONGsYaDiEbn1CB8YInbs20384cbWmLExRz40oJ69kXVIQQ3X1WPCbcO6
6RPLNY48b3A0M1ZV2vLgv8mQ5w0iwuX0t3UjGHGfh/jfbBzc4rEOWdHf3pMvKnWvOnsi9x9Kwrdi
Mf5OqmaaBBD8FHdc6BeqD5AyJM9UKSeBe98qzCsARspTghBkv5Kap2huyYgOkIZvnx5jovyL5S8S
X2GApnE3FK9mkzMj59hOOmK0/1lq4Nk/didmCx2QKAhWrL5B2pjuV3DFFUPnQUcx8O7L/0KClbOb
RZfcflc6FhVZp4j8fvalY+BreaOF5a0ANajKW6CJSObqXVmppY07Lf6NFj3e8fa1F94VU3q88W3/
4gNqOpdizSNZVWtbZiy42xhR1jtC97VooXVKoOs1CP7XnVBSAQVXeD06uvS7SqS6RwtzTfnrgJr+
mPJya3+nKhWCkI690q2MwB9RiZM/DE1py4RgLRTaEP6Ibl9ocvgaA6xRjykX2xqsRdX0yD1exrlB
vuZtVsLYvjcd05XuaMk2sUtyPTWK/tNd/fXjR3ke4/S6t3f99rhOSkkTNLB1vau1Wq5eMyLbEhAD
ETRFrUlsf8ynsLJxt3tXyLGU/iDiGb88qHrXiqpV6W8WdKpC0N8VXAw0JVFxQ5sc3FzGJ/o1LsHP
Kz4j7d8e1YQh8yVU6ZQVhLhDWRWrpR94/d4D0Jxu52vwvYU84RZ8eSiWNKGpeyC+D8wi/pzAXPTG
w4wOeGq5IHtbCPHQ3AUtDm9q+bfF88pjzR4TYUHYud0FICG6KsWRky5ipJF3Bow2j8ICVsIO1vMz
sXfcezTZhRIpeEKq26rckqmnCwzRD0/Vo/+n9GCWBQE0bwiNzlgSTcpFstvFBOS7nIqbqNRGGSqN
WoY9gNsZXU03sRcQ7/B42w75lQ82hndKer467lViNjTDjBwZDlgBNvVBcJHfVhsxv9wLwRmnJL8i
6wz/aihhEIokII99/zq+fGS3URCD7SaUacvkxCbIdAuPb1t00RI99M9r78CqHZSF0pVx+L9yPvvQ
fsHgdTlazq2R8pIxf0HWR4UDkrMXW7q1ZIiCQIPznf24n+t6tCvckYScTYL3vWDiJq3uONGuBWCS
3LXTj4t6KnTpKSC16Zo3/HjvnFXsjdqVWV2OeBzg4Tm0P6Y3b5+eI3bwduHIjg4WXyM3hncyA3vw
ckxRyMAYyAMclkfNzR6icXFheIWnqyJrzFgBEZNIKE3KhAkdQPgCA1NHeFTDdbeAJj9s1hfwCHpq
Ec0FVlmqiF5jB6D2/0t8q7VYhsObEHpS2crRxfklzSzsj2JNIVE5h1I4Mv9o/Q8tBem7IfCd2ZLD
gO9RPApxl3btmPi9SuJ366hhqBCRodTnTyMtPp5iDbgs5pxQcbkjA7apP4VlxmBAQ9geHEZo2MNE
nHQue/iBDweV3LzNg6nrUZyOaQrd4svLQUGjyChaLuL32o8ae2MEJp20//B62iqOTWlo8p7HXCrp
6JLdVFVr4b3AQQ7nCgIAHkGe5E/lX6YkLNWfkw2drhgWzZxZnFaB6IA651C1ChXFbYASapQGypel
hR02lWHCLkncVEh8HocB3K9N2p/Na+d6VW1XA2rf5wt2kuf0cI6sIvqDHltUSd+m0ud/Vlkt14pu
CBhjWiCEaOhtkNLLmRnPyI4Su4eilxfK/uqYEuketLn7HuUv5E8TIo1775kLXkiB4mWfmRNX8a05
Q98zfKUvX9QsiVIXxNX0saxpG+E/+QaVZPOI3g82ayErl6veM9iHN4fQmeeyNgzafhvAxeapYw4n
GSWCi3QAbndCyWH2Rf2h+0hUINQs9d01/Z1t0FAJmPHq0b0+JBvnB+RnDzSQvKWhxn97X1Eupf+V
u29NW0NfZ/uPOWoVqSpA+3YKLTo/2ghw2VCagQmNnlkIGKdhPdfTe0aj45fnlJpwzMu9e/TQMgy3
7rg6iTBYBORyqBcKHb99H3Ire/lcFYi1z543IL8YKo9vUrrk8R68qtFZWSu6YsLZ7XDeVPcB2QE/
iiUljxzQJb8zlk2PVezgIfpFKCXJEQwSqIBYBbrJTFKPQYU4tvg9lsTl0yTwaWXTH1s0l66q2g4n
RPgPRi4pwTJOTdhqeOXuhCXB3iQPBzudvHH/eQf3khHSDAn1q0ZQdbnsZ1wFpEpJWl7c35pGmxjY
3P61shpqUHcc9pXEQhZ5nUnP9OYUJzszuLLCf03ZN3aehuXqIE21BUyCjSIJuEgPMxa7O/YjFiOL
yzmEwUZ1hQqT21lcDdpH/9i/Jte9bH1zUqBSEBI0XBeDclLCstK3y6ErCzoUaem+0NTs5oI1Osf7
P6GRNs67ovSZa5MrIiSAMZ9HYhkkBcJtBPQhOh33mRJ7bp5mVD6Ja4yGWAC9hNB4h5De9tHOVhcn
aDFy2ez8EahfPNGUjHAN31FIX6OxTdOW0FF6K36H5uLTwBO4WU5AHxMeH5XRtLH6Tosn5fqD6DUh
dUsGdKJHR4c1UzV0DVLbwag1VuUNMU0IVmgZptUe7C41FVHzMx/FeHnSAfho4Fnnd3aHwq7pl8Ve
K2rTbnCm1q8epcQ42YsBDjX603sgVbyeRklp/D2lROCsTWzj3oyd+keXpZCxAaYrq/8XX1a00mze
kaPcQYk6RXRmLc/CS7IxcpAwq/+6uK8P5r3fuLlsoP37DiPSrniZ/lOE/G4otNsx9pUh1qHbAEI3
tXmg4ZNMGeW6NIKUjltDAdkfD/ibCHFRoXDISvyUORxMC4PVCK2Betf1sJLGX3J9IfJlin3aJ7pX
/7MyA6FgVx1ZTDchrwwDVQ0xti3jW1xCVCZKDzaYA4Awnuz+eqd/8WSqIr7h8CZpS6XZlJ6UObOD
5zs5FSHZN3genutk8+44n+OBQtTeCHOXv0tjmaa+WVXLEV/1uH7UFzC38OjtIYaUAK7OXf56Xhp4
JWLB/sJHq0pzENXZmJwPTKGF8ypHZodq2Uod8QQHzs1tf+DOnBqBd0Etu6zTupuUxUueu/o4fYpk
EQvtrecyIyQ7Ji7PNVgyn7uUsj0Io7AyDhGjhdNZSbwAZu9UmRwWr6N90n2VENigwxrA3l+09RCg
DYlBwbLVw5hP/QDyTxDNaq/DaDIsfeMJ5xpMUdDSBoS1jM6q9yT8dmvq8kV22AiKgbi3nloUgRr1
hGMvUcsGmX3wqLIUOdNfsVuyatcjfgJeIdoNC/6IkMq4prY0CHdVYEB0TeTQVjxOEsYpewBYsDHa
DSBlnZ48onO3z7Wipy023tFIEheQvqXsCkSRuP+jB6TU7gw52zHLOSFqEljgeW3KPc2+pmsJYC+S
iF6CizOV4lK9pFZ7aL11pIRFXGGh57D24NpK9XFHsx8BPjnTYZqk1hxoejFGOPtzl26XEe5XH9PG
doMyAWYEiqSXqBzdwWMAMBzRlkKXpgx3oU6bTW4L+wLhsAA4PxUDRJhglRgN3Nbp1md1dyQst8Fc
l3Eq1PQC7xIJtgw945ZPVXUkwOz16jl/jR9tvZGMsuB2Ts6s7YCk2np8TRh51gzkxwTC7fwPuNx0
Oi+J8rh4BXW6VY+Axl6moZx81vyy58SWW/5t2Hjl4ZhSdDXD+hrzWxNjMWK6SE3mZ5tTvKFyJ2Yi
GAX1icKDaUk8sFBGJByccidZnXVRWi7l5HC8Z99iY/JbbiWoaOde2UNJBuxCl6uHOljP7lXl3Ppx
GVQb0MvzBhUCd0pmoAlARKkoqpb9sXj4Ju7lAYCb3vkA32X8MDM4DhIbphAaYTlyktacWYV3SEH5
rTVr9RhXcuxkU9YHRCQVQ5CzTDHpKIQBF+ez5tp9da4MEo5/NNgrB8N5ogutcz6y2kiqoYDJiPxZ
Mad/Im3I4slWdh9TIWclb7Gw/ZrM8UrY0V51mlycwVLUGS2AsTsCF4/de1F5M+aOY1vQhy9+6iR/
gvxFXuleDqk92LWvZcJjwApDVdRBD5HgwgxIVu9la4q3j0ZfXRFVuypQ02+1Vz3jvr2QBIFbpCKr
ZzcqViiVuWaYEkYYvyxYgNfz7Kp4e8IQ76VNe3f4eI4Flk1XeQtbPcoiGv5eJwhmb1QZs2Cabe05
MwbqpwU4Uogn8aT2jrxRRAIKS5b2dE9irVwjTBmX3XLo1QJFnEmlNmKpU1ZW6n1zv4HXYAWllJ3Z
PuX78ov+nVasIW9KO+glAVtrAblZwmCQr1yQ5LQJ0jQvoKz/JWV6N9Pme5uCKBLLrW9SaRYNWC1B
P4evyerWwV56HxxWoHyWUjxVpVznBR5+OtMm1BMCfkvYWy4xWlSSAYDWxP9y2IhYuTMVT5AsjU3G
xEP1G9B59aP4TzeqvIdRjyq1Kh3rZMo50TsvS3fkAirvZQEaRc8GHoCV1xcntWqGF58tUZbAU27Y
wYkQf4CnoBmlkOAZP7wGuMX+WvwoUDJd4ohCPaGa/8jBPzMx8fUeKHLWzFxDOfMdIZ294XAbgZgD
blUu3VvjhD8dDiBml9ODSH1EE9v5RrXq4DiCAhvYNisz9njq/f+XpAAYpPHD/o+bdtBFfaJNOV/y
HA0aQcPJr/AQjjngQ9zIjbAjeQ7byz9OK/vQlPleh706ly58dCLH5+mzegUyTCF0USBG5/FfvVYH
PqTtUevppxcOIjwOosnTuu6HIzMvWjgERHzbsUd7cZvtLdg04XyKIbx6D1b5WD3807xYE2w/fAqW
BarQkjuoyxl4Eu3txS/khAL2r3v2kmz8OFyspEZurPjyjNTdA4tR7zUWZbpnpFKMU99PA4xKR+Q8
xHwVYjLlReaoOhuKigyf36o0RXkpqLR6BC5hDEpOKMxvJeFMw5JeiryjqoWnYHADb+zSy1xZcHVG
MJOsmT9a+9ceu1DJ9cLVZObxEhYCndxfUiaX1DVebytmSM8sPck4qtBT/2PJCKOsE6HUCRGgKTlT
CdNgZRTyUYkEW10EOSCd/EfTWJ0XZswREVtHsATxCd3whWYLmoBJcvedpVI1a1QOcD+Npc8ghi+4
BCAAmbcAMORA3QE9+8dI1UHiB0Aoe8tE0ZlCEJi4vRv1J80RUatbAFtgUyeebZHqXtT3e6d9ZfGv
nt/GoQuYvI4rAh+9t73OlPWcB6QYA7Yf7Wz/O2fpGVqQoRg2VF1plwtnw6qPbRbaFVuphHIcObSA
kXY2f7kew0OyTmTEpvbjfwHtBR305X8w+BRUlPb3r/9B4c7Fp5i5NPJcHn4/zj5MO7K/DSHHhEK1
fiWEMF1nmRD0YveUeSuVQbr7I3I6SwRV7OwlCBbFM0ZICEMn38cTnqkdpkS5ezN0vYww+xNmN2jW
ChxEqN/IqmF4S/SWI9E/IM/M+QAO1vEcT4wSabVaryJEIUmRboXBMd2TTHlBZyuEVluFjCkikNdA
DiC03ABd2WUzIbrgtcxNnLHAiSXCTfaviVDo7QP+RCQoWVuy1dBwB+ERFlRhy7jga9gGieyouSGA
o8tBj2dZ52gOL65yFi1uN+LN9td53IqycWKQSDNEZ/DR+yzBCd0+GTZHbvw/nTMbtW+0/xiRoeZq
fTRbOx1LOn00rJxdJz4fAWC12Ww9EWHSd3gEkQs8iRvpFRuZ0ifqlAXhQDjzogP2gQdCMgk+LuZ0
mUUObdmqVGR2LD7Pk/eUDXYSWWxNH2TZD16bFjA5cW03ZlZvFhC0ABDsz5iidOXSxArPBUQRk0z2
EZdGL0/irYkG8foZp2wt+Hl7M4z4rUUGk9iC8dfdLt6b5jbqzyWyrbHnIczslhGgXVY5w76vyjl+
El4m55dMuFiH5SRg+b8ZOlERkmKO63q3r5CZK0JqWNFxE9KQVbssxrqTMi3uWHpqRMpD4Vkmw9A7
5JfOxCpxyTp6uwAVgzfZVGjvTizsMabgjrIccEIz3myVe2LYgNHCoWOu0iQxz0//2bmmIOfp8VaB
Lk2hI7rB7NNIh7QfjSx03mJK57wNGsfWPUsqABV6umLKzmI+A/3NcT+eDA9NAXhcW2FNe3TBVwgL
58jye8iQvqM2vveuRazwf5uM5JcsesTjl9DOxUEid6lkbQVt2y5T85liPyimVEf/8JmPX8T2a9SE
uMvSkYx0T4Nvdv7rc4B+A4RCFQ4StFzX9xfwv8+mykiIJHv1/TMI+16AgvbAUjJSpdiByjSH9U0S
TIsKiJvm8sFeaoKBnB8G+aYbtIXD81bYjq7ek2azmXysY3a2aLdUBcfzn3+l7dXo3agUML83yGYW
t5SEDluEGYwtwvOSZaTTji4ciV5mblF0aNUiWCeVrSCJDQ7Bup+ARaXvzBcn6oew0fBbgp0fkFHs
7mRjXcy107lCHo0YMo6L4Z7hwkRF6BVE7jVs/tNrDgeSqBfppMvX6KwhVyS4F5Umz+uR9fYlwcsI
NjU4aGCCoJpobeW4T7cEZX9tiWIUWrqbO0HlnLb5YKSFvs78wtUNzNmswr4piC5Q2pLVjSdY3hzw
oKQcjflOWXEWrTombhsU8FD4ucDrsir0t8w8J9jTzBREFUucOGqwknKsx8Tjb2vjLsXRsNptMIaJ
Qo85iq0QWxh0A658z7c7KrKZOPpbmjiGyZDYNAUavvmgEbLP6XGovZFmLGMR4ggHsJLs50MDDCjD
KyNwntltlkdGWML223t8AMYP8kx9sRWN6/78+khJoK11K5Bv/kyTpw6SeekKN4Kv0lUIJTzWD+ZT
MzMAx1nw+RXDaTYjZBsiozKuBIZLpCjBu1aJY1NKfXBpNHTOeIggzYzSJA9HyQ86/6ZPF8LxzL6F
C5r+9kfpj1p+vX4t/AgJHFwM+7CVbtfsOUTYFEbg4IhtJmLflZVn4uo6Kfdq9JIAZkXHKgi3Vzec
RcnXcXOezKBZGPNtuI+kKbUgkyRazObFD1EknAN0A2El05K4mVoylM+W2txbAwpgFkDVDME+nrRg
nNN/n8qZZkltdGV/VYzwSK+Jd5wCC2sIw7Cm0Aj1DirQ6YY1hyIbh0N5L+VkmZrAuxAIBKNDIygc
NBWkd8xepDpGXaXPtfaEPgxJbukmHNLbysFAIMPOVFW3c6WZMpcbaZ9K5K5dpjcqiS4ro88hVCUq
UVmAmUPSRuzHRkY4rvghC7WJQdpDoGx22NoD4PMAJkyD+Lmq/I+XdIjp+0Bsftx2teuBA1P82nkb
+V8UeZMzkLoqV/E83Z4FKH7EPwZE6Pq4I+d3+6AIXSm5n/o0+aJJ2lwKBICUeEGRVTY+6RB05RLw
vd5cJN2x5i6/qe3uFyVbBiq67E7bOhrr+8VTEyvNVVOu91LiGgNz+ALp9n7Bbfr77jHTS3AaVwGx
alAzyWzqRvh8cAJUPH8c9u7M30w6qIrf7AoPQzcyuyq65BuNRhGLzZyHebfMUQQLCNnw6DhUp/cx
vGXbwv2ssfyXDIBdwFxSwQB+59dURybLEpIPCTJC3crPe8rsf2ApRGXm13QVLKeRtj1Rrt32aHUO
F66aWTHlP6zGtxMq1l9xMNHv20pxKJUaEKgLiCU4BFAC5dm+x3O9aO+X95v/jZ638zRtPxZILwnm
CCWcewUjvmzlay/S5KsC/bVCQ55FGxwc3NcI/zWhW36daOgo4TQLvBOcpUvufEcu0PACqpPfz+/T
mttK9m7i0kO4oAQnvbOPPbw45VzAh/8ha+MWD+d2CvmzLNmu7zPKONsI6X8T5CbcEgAnRZk4aK63
PrBlQvFWWKJyBPrLkB0kW+MLRS8Q4wskhq5DQ0aQTDJpgHob5Z/I6SwgFWIAUpGfIiO6/xv++NyP
n67zc/ehMVjgIZxp4PCMZGKV10tuzPKoaH2UDK5f82Lu1Axh4LYLHlAilN843SQEyOnXBbuIR8Vw
RR7qgSJGvcsdzlxzxHGGSJATPphKRhSH+BWOmHxfS9irRrQnkABTZ57RQs1tsQeActLv2phIFXoH
R255EmAKygDu6K1xwyBdjoK6PI2RQDIAlLBv2FoC7blQ77jFAHJeq9vMCNWDVV2UERc2KzB41S/g
GByiM1FoigbCsWFeqXqvTxGrTwX4oSYwklZqb22SB1gEqHeAH7AZ3nO42RXz0u4Ex4YSIboOys4I
SrLz87EG1HWbtKeAvfdyJSV6JC6Hbr7kh69BAKqtHiwVHt98M2ap6JDSNL5o6wqJzzxjM6lIZWQJ
isXu8Udh1bMlfWQHCWCrVRZq6hy0PFOawNrRmGsOP5C40wt358MiF7F199JjoZSdvEUnu+fHifBw
BIyd06HL9HHpVfQ+nqM61ler+kGZ0sR/1D/9ljGDUOK9nC+pXRd/bgCKOXzinEt1Kg4YnZHkO3NO
Uc/lT3IK80G5OMlM73KnU/3VRwBxTGz+InnabZ1c4ewbbjv2lYeaO7+o2xgDQ1VUoZJQg8vTntdC
m/OJ2ZQrWszxSiUnTVAZVeq/cAL00vfsyPP3w34ORaa2S70d/PXJsGy+1qCdoSYReN+BxohXbves
UwgwswQGFGP8ubNAy9dgpRuUu3p/ltEI6rTkEtEdGR/V46wVeElHy+eIg6JrymKayEqPm5hX8F+E
TsCgFPkUY+wpBG2WSm/u5zgmHoahYrpoNxqjOhQOJiCuDEbT6ZT6yg12DPdWZnqcSVizl4kpyFnA
mVz6e3rNhpYYeXN7SmEXoYDaC+1XWl/+QjCJKoMq3rfOjHd6KsjczjWixelQzmD7netCcmyIech0
u+f0Ex3Cx5e4bBQGYCVMMY3c5dgeEjlX3Ae91Dp0URhnl7DMeZ8wYdAI7hThX/GSKvkYufwBYyZJ
4nE8Q4Z+1uGCTUU//MmzDLhszc/ZNbtU9/CADrvZU0vB5Z3i+rv8a3CV5MnMqrgUJ//3xsJud04M
OsjUI7dXx15raRQfz8+qEk9Zey21qKkULHbFdQnFFi93c6kl1oLaL0RpRP8sGiHNi2+jaJygvv4M
26Gy5iO09rTeWTPjyjCkoW3dMTaD6/rYi+k/TsUlYC9OsbCcv3XZWctsiJwQycKrGoWF37T+Kp+D
rDxk0hq/oOkqqIcfhxdyrWPuMj4xmNPZQcIzzODCqdOAukWX7IoY5LCwpjhj83Zkf8PEi5igI1RY
Y9YJsWNRQ9O6MllH+HyMKg1YSH//DWXblZPMfi8YS1yWbPX1zwt0YFFv46cSn3Jche3+uyBs7qO2
BS0+uAnkOP8s+q2thK52b/SL14Q98DWRLfzL2xPS7klHv0KUPGJBULDtnQdFpTc5aEtSjqdY8U9U
GR5HUbUg39tFYbYBlii7Nh7ZAHwVPz+vpHTfKtwq1EGA3eC/vOCBpiDL6fPmnOzYgDtpt2PGK+Gz
ksnwLwzsbIkCDVq7s8k7ZlUmg0gB3/FX7H3YjKK/gbK+XLvMsFseayIdr9XVfwObniqPHv4/eODO
UbTDYgMsUeEEBl88q2GYLyU5w3oxJ2m1ZY3p2FuzebP5NN3WZVzs0UbfOtFqdlZ5E5L78bANd7Ou
J5H32bcnzn0f36gnHvakTfxlf8PAO1KsVkLWvgHdrDaTsv6WDjtaxYUUB6zoRXQZX7maAtdmK6J3
RLL3xjWyaW3m8Qm8q9DiIEPtC+7PJ1pAowkBfI4W0rfc7Iakl604kweyjEjO6OAz1DdRHqLn2Ke8
grDrIJjl8lru698O9WOEFEHI2wLHJ7rE3a5ee3vZfG5vCy0bzq8hfyejJiHR0di63nk4Q6WjR+Kj
jyC7rV7SE02JXTsA1KpKckAiFnRxcSLZ23VpMNNswoRIciDjx0yonNsTJbirxBXMco/Ek7VMtkgh
RPWBm9mm3eQGL42vivxxcF0gLudYo9ptYhlEdboIJ1vJjmxsdyOQ4FTaMdGIFwLVjFzCCeXyYFkK
GlqM0DI02n2/1cotTV0Qn8XbySDHJBh42upfJS1wyXxJg7QuUH0Bby72A3xg2V4NaQ7i/J6hCbqb
sK6lVQ1sUjZp+2OBljECuAl+juTPIW8T9bWfCUyS9tVZjFexiVRQrNzD/ySuyaCAyIQYFoEpy5oc
cnP/7KObBSwmTIY+BHlSHe08rqLKf0mYjDQh3eR5Q21qyT1zT+qxglCwbYPN6IQf1p88yAikQwPl
CrrJY9qO38hfFCNTFmM87SYloBkgHltf83dqAvb42QyrbdJoxzlLAGmh0yaoDb3JA+CQtcoyn5+/
jFVO8JKdjRMAX1qTimyhfqVYj+TVnsl3eEZfsaNgUTHomvVVdvCMDEbpE73LNAjo1JhMhIyhHLr1
42O4s46SjupKbbb+Yf0WR4iUT/BgKP5zwL/fp6CN6lQZVIhGBCQNN4RbBp1hcqpxXa3p27MuZv8Y
ePj+erFJWbaoRaoBPksgeTeK7Ivy9AfSs4Epn3TSADR1B7RkPz1bLnOqsD84Ef/NJbIzx/nlxts9
LW4yqW/oRKGDh3DKQ3iHvYjjJ0Py9glikS3bMxIKByadp/kTwml1Xiv6nAwhL+kzVbnfXqyDMfdP
7Kr0VksNKcflN+4Iol3STfoZcCqtJW1isIoNC9sdLx2fHQu2tr4CnvTpVWtyebWK1IUYvImvjuPU
HKWhHXQOlZTLuXH1B9DKsWLnu1poCXtrKLsp5cm5bOGJwiz4/MzsFz2Jaajod4E01/1JhgFk+YxJ
7AicfuRikKglM2/PTtmizbr9KrFkn7ThSI/koJSsu/ZEt0r0qIdTq+vV8BJUtABwzN9pjVYqRNGt
goP+bKL/13wgPvR4o6DfMljgquBTZ5ZUT3HfXP/SzslNL6fyeS8cMgDCOn92HeK/1A7a43em4asP
Ljq/WkGFmBzf+5Ge9a4Jq9dSqhJGtgfe8KjhcIHzRR1XSDzVSJ6xX3G8fZNGkLo8QFPaYNarmqbM
YkQH11BK8f8KBrcLmwu5MMYiOoVzD3R62rb64aCUI9bcLYSkK/w3IK7E5u1aJEIzIHYFc3oCHeqr
8+Ph1r8FceBnNOjS28rZJGCyn7mBwiuaQw3t3dZ/QXhdwGzELHULUb1SgDLehHBl/R8j8+iFOmIc
5rQnCutAhLXh77Z1caoEXqLKklfKiSqpZQWaHEHO4vPNQaoVE/4ILxMIcGHcBLLqihKMpG4+0/gn
Uoj98GEXVL+sk7Rf1TfC3SrktoYuMoxLOYYNUs3qw9R4ERppNHBgjkd27htIOhgtYs1B+Wuud1fQ
6MCGREwsx8WDq1U5EJ+M0CEHX8r2FfS6FAKInpOrDpjq3fHVyZ1P/hE8KNZZs5xYsXs2brfx29gR
G9vBUeWbyeviGX8FePT+RI2c/4WH7Zc8E8oNAmBNbCfRxBHJ5rW5+VUIHb+F0K81q9bOn7ZwdytD
BPpc4uGT1M58LDYxbgKo4v9hprnYRzT7TgtJX89ChVOekmo9BqvN7DqvZbW/56k8vDQRTVE4cupB
EPkaBBbUGpp0X1/BexMk6sTjUba9PeFl+J9Zb1ljiG5aIpCJoob6F8g2Ybl809Gn96VWaPLonl0N
9ZGmSAayeoD+mLW6kaB85S2YHYSKIB/nk6vtxrhFKSoa80PfPSNugWIVukCxZbxUEWnPWhY8vnnM
krB0bhgQtW0WTswxrpWYoB+rlz/x64TgB9PIz0VBdfy6pBfuj7A2MqZCKIPnPQGvZOI/3mfuxMO/
PgUuvN2VyFWNJTrtcf7zne809kWWhUJUnZ+rXyJGcGw/op0ECcgxBZvX6kCFsxZ5/BZUAAEWi3Mu
7pypgwEItROaicARh8VY3eOE59vByKD/4v4NTsWoKutfrmUzRduA45T0uP/mad7ZVd4h9O7KExST
FrOj2mqil00cXpElkETcz/8cJyMt2v32R6Xf3PIUF/XayVM0fsmnI6aKXF+tN1ruu0y4sbun5Rxy
+TgJ4/bO5ADbiGnx3AiNtRU/IAevl3R4PXLzjmLyb3FDRP62YXVzWUTbkzMSS/ZfvVW8giOKK9dn
bJ842935FFb6ofuhNNMFUUXMw/JJPvRmok4KPWHvPu64YZGOH0ul7dFK5Ly/1wJomvMtbQsOxMBo
CfM8V0dFY1QCtO54dqWa+2x3xmoirTQ4XTZqsAqv5ilJavb5SYC65m+/Avli35leOozL8tjkBGTw
QZYAqJ1YAmTBnSCejufrc/Apy7cmPCP0BKaPkc0BalVpNEaPrPsW/2zyV0/gHr/ffSaTDaxHadNr
OrUkkkECNdKUxUjEjPEYIqQquObQTx9ekKA1PbdSapVJRwMshplcf8eqSlOLyKobth9ln6sMCIYV
uW5uDsPMsi7QqlYXaR98t6WpqDy0Aw7Yl6scQJ7uaGoqnQOVcKyYtRBI1koDfpwKKnEWkpBDAG2S
EpOS/FeZaBx1MGov4dhhvOhehjdcCRtTM+/V2DVk29Yye+KoiBQzYV8bhHjP0eYbqmzLKZIyqgXV
W2GSO8kw3xgbtBP+lZpQA74+PZfj+MpKvRpDKS/X5n6iJP5SAhmCR/52i30r7f4dpLby1BC/yi13
VScHoq6xpZXQUylzr9qG9tRcr+KNWkJZ4r+2MXfBfhw6DZ5XuH2ya+YEMicje7XuvmeF43YIxDU2
zwUJz4WXMz4Ir+4VLytSJgjpvz6guXwLTaOw0igFTN/O9JYWV2aZkFsL2TJZzVl61V4SKFrqvEz0
36V4MCtLyqfcMJ2Y+iuFPZZBOYVoYwbII8KGTZ1qLkVyiuOQHVDKWSzYP69tJMzzUlPRHLd2FOBD
U+GYNL1tebC2chW8A95iHxpLAs1d7RH0I09Q/I40GX2UeJbctPbTuPhgLFWDLdGiPJ9I/L0NCjHq
KgxYqK8szgwA6KUUYyZUPaUa9tMGIyM1+0nnNBDpQRFUlrEF7BGJKodXOjoUsthWfcVPF/d5pAtE
MpH3CpCSkmqjtEN/xYRTVRNLiURiSNk9BpqMnpDb2VkOJtg2Ir4u+gaMaF9vLXb/ybp7jFmkVTNz
B7JZSjNqgWr9N3ktZTfgisvqmMrSSF/EEbTWxs5V2SqUpCiSTDEjDzFrjONZ81TUCebuInj5DeUE
bEpV1ONWL+dvolVsJz+xYvZStRe0FOKBaCWaH+4w/GWSbUOQ6F+tCNdfNSZPTSVnyWB1DUqQ50Br
Wc+YqW/EephdhrsRuwbWsk0rOhZRyLKM3VPwY/CteTp29AjGNOkIXTh7Br6UdKMuySC34mNq/6Xw
HsX/aTto4jbH3dc+K6qeLLcsyIOmiVYwAT+IxEpaaqPUWzqA/m+yUkeUHatFYhtAk9oA52LBRE8W
hrw30drtN+nDAtAnkXmomnxE2srFV6uvYkEh+9dUPYThFWN4Q+t5MdK7fo6NDKJ5Nlvb8j2ke82t
iNDULYn5qa3hQODKHvL+axkbKOnSS/qLQauw7jOSlbTLl6m52JbmU9c09kN8B6vK4I8UVvFLBtwl
8h+gj4AZ7VhHbDZ8T8u3tsiJ1DH75hGChSNvuTRsqoojyVjoH0zoK8gSR7HAG7sK1sIUm+Dlqt6j
f4QrNjdGSMQ/wdpDqY9ku3VmFIriJzNoeu/sx/hrNuSMbMwaTAZ/Sm5XEFQF7it3JtYr1+sb68Io
okLzzzZomqEa5Z/hrSLuahD5ihSX65vI8YhSlcHGixO0gzmY2YRgVx5gmkR4ocNZrptFNrGxy4Jk
5v0KajflupaQCcVGh3dOdi6cFvJAfNLDLGLCOS8KS59kXwTPHaBX6pDZxPtTBommvXv46Aw2MVXY
Us9QDbzXzg44EOmEtg3A/KTI0qVggIiOPoxBM70MPgUE928Siyfdf0SeeMO+Al/L/wyZpO2kU3R4
ko2sy297eLrXqATgAkaTEVirVw2XrGrLjI2XAFLLkD+i9V2A+AqosO1q1wYr38rZK08+MgDERY3n
ZHRi71kkXSMqRKtuxk+7DIQFGJYeSNgJ4tDBrYXo5J5MCyKSVc9PMiZqWVYD8Xx/hHR7rIVPwLL5
hDub3h3aRldMr2qTktFEfoSwzPKfDum7XAUrI2ZL/Uhp2FprL4QomPR+s9Xm/9GKjMclJkG3dLDS
zxgk5y+T6I7UKepcBK1Ylnf05MYAUmqnl1SdTkvPgZcBGyIhZsYAabDF+jeXNixiI/Q0VzXGPQBo
JjCbzfXJZchu8eINfYCvLDnoN5B7UNHEscFE5ziU3c07hH15lQ/G5TuTHWRr/uFvz0xgPg1XRBjQ
6gTe4IXgn+TbeQE/93inUxHelE0sP2Y1oyWdkFqfSPh9NJvvqCPDLcCw+pwQwPVT9ANneX61IZvW
A3YVINY0kZ4iAZzTHjIwd4g4MM2Mu5vQ+Qi2BAcXHNaVXnk3+aBi8i63UIrlsBbtWB5V0ZB6VDEV
FcEBew5REtfhO3Zu34yUDscIm5be1IMkN96pNHCpm5R9r6L6tDpTgu0FOi46gu7b4xP2aecBe9wU
vFbv7tkRvSQ0aI/8I+o45cHO50YmwS9R/wC/8sCLn32wanRtyAymtFWfnrTwB+1u1tlpgaAoTYRl
LCJQVQw7w/ovXCKHE488ErTMfSAtZyhRMr46Wd32L+/1imWVbXZvP+w5m0umf0zpwp2uweyv2heO
5jqAs0uaE/2q3WXfm+hjq9EX2Oxgu7wPebQJj3Pla7t8Oim4ltjh7yC21rRICw3FTiermXvEaBJK
wk/Dw05YbR4rL3BU9z794XwtciGhKBi0EuIObjn8WQc1DJhUkrDILJgmmRgcevwss1zCoUl+JR2C
pH4BOdJ2kmzz6HlEmN+liVFzjU/9P0gNJZ1Q+qFw2aYBpd5F9f41ym/6d0bb7A50d3ajjB3Draml
6x2iPKyfVNUtvoSepL8nbybOpxPugRnZlzmvSydzAqUeHECyYBH17AqkqUbxZWijvaYbEBpK/ev9
V+tcNgYRtmIRpiyIa2t7RPcN87/XRXwqR8yr75QXRy1pcoXJKg3bHe/1rTetuyKXk4Yhshgisunu
71hEsB5EIX6iQsba7lRnL0FarwtLhhnLakEsmAGIZi5+wreTSysFsV8QJpP3b6gTpyU7LSpt7N5s
ZtKQ+nkdUVjp7VWXciyBwfqtR4hKKF24diwMzPnewcgIvOrHBPA9nwyyePVRvGerCwFozJAtHaPR
rSxiHqRDXIwhsXEDUP6BhntUrqpHczMV50/q+RCdVJtLE3neaPlWEOINYPrq3XN1AhVBLVba/Nmn
5jvUwQJqQCkFzwKfdggM0FiTxNfDxp3h3gevxiKN4rsj7pl3/gWL4jNlUArEzoQFjPjyvBEaEZQY
gAikIqX99qb5IX/L/qNGEx/2FQKPG90bItQz/xneR/zkBtX3ZxqYast/YVMH1yE5oe0qj/IF2kF3
Cgvuhrt8iRU2PJg+UMqs3br55d87RAJelvSmk2GXirpDF33FLh6MYeC3kZHtScRfiwFJPunLG2aD
C64SGAekD3bR2YO7jl1PNU/szFIRqnRGMtdACIhtoGKcO8MErIvSRDZ4R4yRj0t+8ug/iZHLs8tQ
9SuP2l43G/9H7gPfpbMqz5oHRMRV1Fp1GhBl9kYAbgaFsPip9T+ho9obw5Q5cRUhgmYTincVF7op
5VrSr5AW2pT8yoZVTjdtrvmN/mH7yNjxGvkW5tBToMntHPgu3OC2VxRrUFGLydeF0QCmGZ6rggty
N5PDJZfj+h4bo/vZyK3nvwFjEy3dVfKyEtF8RCIRoZJrSyItHbZHyFVz+piIOHOAkL/FU+ypd9P1
syvvwCmYh7OWM2g8r6cjZsZhBzCJ9FNO1uO6IVwUUW0jbfXWw44gwFPCMnkm9x+rQmBsZr5ApIYX
3Mz61EPIZuL/MsxeK1uHiNy+djquGRhIsCUT7bszr+PFYaZpIUHjcItfOYdxHpWDb0oqG9NahHjZ
4QqiFWhoMVMC7w3koo9ByyywC7qutQ3+ZEWr/Xnc3Q8wuNcFXkXoHOSIFBRGMV6bTSt6MBq1jwAb
/+jr8a5y/NvwwnC0mj/u/vgQVJzuTNjbguHu8cq/Nq2i1gXcM5Yvq25sAIu7NtPDkrr8ia+SDIP+
Rwuk900Apbgt/+qLP6WKOW8ngQRW46DW6lmuoU+1YSl/hJPGOXm8ZNLlmPglcTTz4Ub65DNRwfhW
GmfV0o0j4u1rkPZrXqNFn36VsCaISvBe7waqq9fMFX5srxdtJsLw/nKBN0RcjWT/1RXIwxpMVsXu
BpUk8Gp624vO8Srp3GEBRQFlnX6TOMw+mivzRK0XkqMr8qAf0fjZ/Rv5hcKmw1Uyb5FyhstCyLBm
2l4sqaZRR87IHKKP7SQXEL8413mWH3zMCfeIbTboIxRxtQh+IyC328xcwQkJV/VzcLwJiBFGV7O+
+LdYAgOql0YTLtigUOta5Malp2l+0jwuWq5XjSNiVES23wzLSlgqQu4Fj9IVeEVOKFK+2KACuK00
QB97nE/rdoX3e0Jyy+fZ2EKErqNui9B6maHhQ4pr8+XadHILNxfzx39lY897wSI8F1Z1BZw5DniP
cKYJHW8nydU7fhlWpmlm73uGcL0ImMYw1vvD5XuHIT+4pBbFCI9u8cXsKyDTmS7QEdm8bH6Id6ZD
Xg/VRcOhjdSFulEk45eagnI6PYtzHJVhW/uopBpHeNG6k3NaXYKigvUUSgq/OGmlsap41s8QWV0W
kfY/Z+2ZCv7/wCnpAd4ItfiAxUoWU922hWvgQK2REEaLO6fHInXg6WtMCp8QKTJG0H7Upz9giT9s
2NVV4GVdr3EOwnmvBSk8S2Dz3qJjT9X1DJP4CS852BYuKQvi+W0n1S5VSjSbSi71srkuPzUC20/2
8x+3It7og3LDdYn4X97WZBu6QCV4emAJ8MYNBDXw74X8chVTeeIaTk51RBD7tvfwiuOpsVTA462K
AxW4ZLABVUBKkZaFq53AomBGqCyXiQQj5VGsqBaHKVM6WqIaXRjttRpM1GwKvF/yVmizb6lvf0nD
ydboCq1FXaXTCBflfEOcfnxy/oRlSTxZQIKVq7F+uOLJDhvHOuhY6i4G49oOsD/SLgRNGfPt5M1m
ZcOZJf5GXaH1074qTp/td4/fs4iFkSZLYfrj9z+4JyE8xpokUsNxpSkVH9FnaMhMgg2SeU/T/Dae
dOOkr5M8VtTtS5N1OzTMkDHHl3OeCx8TGLNliLclzgBKDakqEMtUHLx+mdRMGvtDl9kwzATdEr2Z
PcnP5XOxKhKYQ3wN4XX3wwOMS4WnncIYODnzTJsbKU2ViROTrqABsW7cTely32cgax4u2IUiD/gQ
HhUBtati4FZ/laOu6los9yXtGmRdtn9FtR3sX9Qe7qKc7r7djj+jaK5g0UNg/deZS65Of0dz4EDW
Wb/cLT+BkAJHSw7H9WoJb3iF0OyNshvlndSsaZfGCn/YRlxSH+9uUygO5jubUIBwAiOLO/SQmg1+
qmUzMExYJDQjWeaXKOl3/KO+lNnRkmF1Y1Ub6vStGRotIPKr3CEMfdotT+HhMnMwIHZFyuGE/wci
yFPuaMosbBzQ9qdwgb4382kmtWrtKi2gChGtgaks6XhT30Zc1W7G0UPvKIHv6uxOE3eaZDnCWz8j
V5C5VTbDDsJfaJbiX/ACW/kuKvbQIw1N7bpmdZoxp4sq7IqKAwgV7PSPkTK11itM0q2NQT7/GNnG
hQMuC96uTl2RvEDqU5uJ9Wy3gx2aVFGq172ZV4IEdj5bXNh1teypP+EykjtfEKoUVEpDI+BNMjoh
ZCe+vaox4hnYk0tX8i4YU9UIyn67aKyKykNRx/EGfaan495lDSZEBp1tBIWFd0aCz7OC2EtwgWX4
kY8F0yh3lQYVQwdMrhPDsSnpKYgNU8CNX3g6gwY9+/0+ZsvrB2S+2R8u8fm5Z6bzwhWlJ9ASIzRv
KIK4tdDzVVkVb1dbziuWj0+J9eOsO7z2BEMA95UKpVu6Jy9XPD/O+k8ILF4FSm+EcstJLduO5Tuq
gG1FAKLbJPDzcrn4euPf9ENekJ4+EobfacWJMFCpfdzNrMd0ZvLb3qRFvOrMxHxHtcQeFSQ4lZKg
y1R7fOqczy+9+Cwiexevv8DDx9e9S0C8qBQ9KFUQSWP+uLVgopSK68Pl+RL6zFAoh3RS/7KTs6SO
jYB8dwpTidLlePankuzJk4EJmvht4JsPDyYcGPSk9IV1OTvTCRZn7qJAJogdafxJsbk66GCyMK1R
2gBBfCyzHPzQ2poVGjrTjV7C5bPUzur5wVVeoZUA/ijHwkUBl3CYekUjYHUoQzrf6w+/LssgQZE2
8RR65bBLK7vGNDGik1uloN6c4rHvITdbcriI3h7Y9NYtzyefvgOuG1KtTjC3ZEoqZ+9g7h6dLspL
yJuZjDJBUdOagmpmR2NyynVBrNY0v/pgjNqTvJ/CCVtksO1VS4hJDYgAvv7DVzGR5mffkDReTwak
1YUHXlcSaEvcylUAIwKLQ/+dWaqxmuS+PxjcJu+5E+cm6Jw7OM7ZYn6VB+6sPkekGu1PUmKAXqYT
HvR0/mAZbrQy8LVmJgosyC7v+8TWkONMtbyMLJLFUPr6TA7ez6bS4Oi+kR/a0uopE5wcmyL6o2AA
bdaQP8bS/tBBD0p+g+yhyf96bm3EG4dKk1RyAynG6z2wRZhlWOrReSzbE8mNTAnnuZFKTjZNXf12
UC1C9tEiH7wGaWd1aEtvN0O/3gSaLlyMBu83tDrJftlmBe8C4Rk8Ugyl6AFoEnP6WRiV4b7M1pNl
q9KIWkHCQLe3qpLIMmCt0hPBe6KYVHRQglTUv07NrVg6F8XH8vxgv1vaHHgfOqvVYo0mqX6X2u+d
DFmTqVQk2uI3VYdR6QRZ13D97XOXiHt0EUL/GhWmK7PNozzFDqrGH8UYioZOlooWZIsrH++742cu
xQVwvPBKzZQPGDnv1ajq0xnWDMFrVdIAE4lr2lWP2Hptvn5hWOKVQGvRAouPJJlMTxqk4F80YpK6
rsihNUQ92E22IW2ZK48R3o6nMkn9wW6kCo4KDdrZu79c6cVfBYpWivTjKweT1bSQFlBpb+7dPfnR
hJ0NmFqEhKqcCWF1vgmpZjrAYWS5aBJKwM/DVRm3X2kPORz134ATId3iwXXAmzypM0Y1DZXRyMON
O5rC4a6p30D7kkopD8AQhH5ReQUa3Un6+cDqQ8OD6X3EdQ8MxV589/Kmh9j8t9/Uo2ptd/CCrcIP
AMsnrJqzV+jZeVDDYG0jat+e0q1IHg5DpXDFbLdsJzhzy5+DuZEXR/FXMQH8jjX1I1wwYUwc0DUj
cBz9Au/hN+qt86z/J8rtyhJp7JZq3MH43CJTMJO855dariWFG5nrNKYywLJF1U4D2CTE1Kt2mAF1
0dV8/OUbSKUAn72Y1S2CYeNPG0oDp7m1keIqmAtCRux0bwcj5XKbbn86LUYzrjG1q3hp6v1gnhY9
4nquHtwcoWGK1V/eQmaK2en/0Gse9WOsakCcBd0TJiPcURpfEw1qcYycP6TMgBxXwgF/mAaof23C
xuzAGqLh8UY/2DqNndcXitaz1gE3rU1RcnnyKvwMOXXvDbQ1eL7W3sQ0ZL/ZfVLSFshIhkO/psoE
5ldXSzX08zc5dDnaeFTrt+Zo5ldTsJm0jafARYno0SG8mSe40JsypQT7BTjQP8OzHSM6LpVbp+y3
WLKY8lT//4nWoyHn9j/WfmGnzBb6vyqLTHO8MB4Vnpb+NJMCuK3ZSrXrT/VKoT8fXKKjaEQQQUV8
YFtsHPxvRFOeEchrmkBxNPgGjNMvA2CYsgkpmC//lZkuZVrMOsc+FRYk259iBQHTbDp5kQ/9kHpU
lTWXV/GEamxYUOwwDItWy3IEDGi+yRKcGTZY/Z+fl0BagdaZopHQhdxyzYYXLKQ3bVqc9Wv66naj
+tU1kmnTvSwk3ZC7GJdukU/kYXamf1/oV+LP+SEa2JCoT4431pwEcq2KjgDqNT+tjYKrj6PksL+t
n/Z1Bi4JYTu3AnhK1AS/Lr043gMow34i4yOCZIyDMh4QPsGqZ3xvdqlcl/oqXeq5TB+Gm+Y31bQ9
SYpgmTj55vEDbhHiGGy+oBga0G7m8XZWlKXqRCRO0TrBXMyiunI8rACrIVe6Zg6th7z+wCHZNMQi
M18zHbaNH8Bo6KLpSeEEA5OXDe3BWWstxon7PUbE1/92oM8qO7DD0tJq4RftLBIfWtzItPk+CvBV
I4dPntGqSnws2OTwuU9Na10H/yph7BNZ9MG6m1Z6W8C8u30uaB+C0yHYvWHmidGOsI5CzJa7rSnG
Krx76Wsx+l4qnmL50KVxIom4JH8jzfLVOvDBw6yErCdY+/unod78GwoogEnqR/6gl+E/oMJJEX8I
7O7o5jkvnW6Z9S5MwN/26zLn54tGTB9mlu6Rujin4ThyxLVKJVf+fRY0qIWiXLPpI3iMPvI1lEU0
ENYhxzFfUq++cJJHibYR/bEB+BD2dA3pszQ1ZeiIFVwhRrB0JgXq6kA6T64x8sWtT4vt9hQjhqtX
xvPphuvkwXsHvZ6w6IZzr+fKZ3TQbBkn3bntDzxosko7atatUlzrA7WH8U3/7MJ0VgtrGh4mu5Fk
FmRWyxxvAgmr+uRDGIB7rxWaY9vpNDKf9DuRdYUvI/RTagVyc6qEwjA2BI+fSx8J+hPmtCDNIRDs
NVwVO/OvGJOE9Aem5stLMdrZLHnxUp6/ANL0tf2VqXFJT3UhpKV7rGnfpXSlf/ijemDDpPXHJ2JL
vy5sLo284ZXI2X4ms6JWo+D4/QQwsVv2cJ4Mf6MhHSWXPkEg9kftg+1RDLZ7WyuTJ5A/frgCA0KC
aZqf48OLl/S4yVhHPjJ/jjVScfOv4V5HwrRp/eOatIWT9yGkgzTQ6Au3rdKG8HmogPd25+TlpxyZ
OFb6pih2fnIh5LAp4Aiotm9sKzFDujE9sZ9m46h+1NsUrJI6W1XD1S2gkH29+DmqvO0mXGIG+lJQ
c9e6Vq5Vc1kpIjPFd1XTuK7pteh5sdS7qAXzNl3j8YYyYpV6QDVpCOA0hcbIvBBUPmMB8Kx/yZpA
LxUBSgPu+Xif9NTeYKjp6duaQyXQS/qo7ur9cHY5wsykG0QBpZMV25tS8Wg20up/OPswjXN/NOo+
ho8+gRVruwHJbPUFcJ13kz+EU8ISmkxiFB/oSuVzP1BWCoochAQYnp6pzBU01Yf+xdQV8ZtEnZWR
V3mYqT3LlbVw7eXingXi/Jp3HO381PPh2/7QZwyLKIx7xBCzO851vbgOdboeHUfI8mvcxCfTRj/N
9cl/qL9EJxyaG7JCbChjlIMEP+5zkgsam3x81fWmE9LpxQA1kliw0a3736AHyYn+NTVp+mUizAp7
9kb/p3NkWZqLQA6KjaG/rs3GT6NWbN0dj4WvlGTU6fR/VppzWj3jerDQsdpsvlD7gHnFk1UhNdIV
zwAuMMqQIIm6vjeorRh24lS4nK/wlmB3WEKcQE5quY0Qt02M5paWcAdbGLwmbQuANtpcS4Y+rCQC
BLvijqGpqByv6rDN4ktNmfClVzoMZfASTmaP9at9BgolwxcCrAswNqOgSNOgi9J0sOLy4W29H+Dy
Vcb0KABFCLw0K3YIq3RI+eruhLwYIBWGPeP2qWu8yxihbjQmzImgit1uXQ5U2JK1QKBXSaueK0G3
X2bIHpmHLkkvUgvzqTlcy00aMkqKmt3TbhLkueOpS1kUv++9AkDlrL9AjLhhRqnajV+UCrgMTFVd
KsgDG+Saulw3RIVnb1X0LTuWeaVUM4+c3c+T/N5cXkljc36+Xcq3q7kdxZ/o9cZVXAOHOZ0hm8qW
hjiqEa9eRzCzGHsf8Ei7EJJgPeLyXzB/tfIfIlDoeWtev03A+FUJahYqcE2+ybrPiVIlohxoyj7W
dj+xXQJyJHOOjz6sxohVX7ccCRHGJSXsG0nfq4N/iYNPW/Tppo4gVe1jCQOX74bvUZORx/ZwNyuU
zthi2nwGMiI4SEdxeZx5f4HxtUNdkgUgGEwYfofXWWS3/MgJ079BCvkL9PTD42BWFr2/dvDFb8tT
Cmgqy3ipTgq8PJq1abujl37Pvruiyj3hai1nLOt1wpueylEMriE9ipoK7usPrUhL6KBXYFebVoTr
uu4od/20/wdit04H35PGxIccmwX8lcoa1ngILnyqjY8YbxZRNVbmt8dzhQjsUlE4EA3X36QalA5o
VE1AHyK/Nasq8zXMo+/3RZ2TgN9E/+PknkqjUQNJCrEpCZHTJrX+fIOF306roIE7ceMU/HyXSWxT
GZHCkJZJ5XNpnlpYbfUbPTdKaMNLVmb2utnMtn3GccYs5KNeydvokZmVRESX/eQvksnH5pyETdlb
gEtgJJ5tNKeG4c3yLsCrfS47vy0m2YcjKm0c7fbLpEdvutUkljSxpTc9n8ss7RE31Gtc1DLGseAu
XJu+W2oxApnHGw9BJD6L0uT2hZvj9ANl4q8Q1g1QPFcY8QJIRfaIdekFYV6AL2cV32RYTWHgj7N9
f8dFbs1jYSIa5bZiFiax3jgQcLxD+9QNvCFIxth/HXakNnIO1Pq1M0Q7SYjps2ErjjRMVyEKMjww
Io2jOUt9j94KR7oBtYxjEtKQ8PqH7aRaEUHLPswumVjq0JnucysB0IxSoUG4ZgVk+ItmKXISNaq2
/xuZjO/eNov0ZvxxI8CZzrzICKtmLLTRodXoavnLO+YBaosQvLMeRyFzYS9iIec3JpmlMz12taoW
OYeOJ+TNSZbLPvrAVwK/YPKlJPN1lO3h4jj99vy27E/uHrZPtl2Q03x3YExUoVjgAZWmBCZc5g3q
s1aDzlLDHj5H3SYxnuU2BadfJijnfplkkvj4J8eG+FIyE+apMxg5Ryzd6+1sjNqVUdY/2BxItoy5
vSJkycqH+M8Z75QCKWbjWf5VC0UCKN/18tqX1GARXTU/ujM6CWFRCruNFQyNykSIojNGKIB/DrOC
kxpz/Rgx8ScwNi1Crp0THQI7j4gTVOdzxLp+pDQtuv/wVA8whdFLeiJMQIwMnJq3HXqcArTEJsjr
9y5o+wHN4UX+MUvid+k7Ow4Y2QzmDenBfh8ODvoYKoIQgsMTNyMyxZioEn9Hh/0J3dcynqv85BKS
l1ClkDaUgZcaTAQNcbdvaUCpqKuv5s7O4H9n52pfsrNjp6eflL2bi6MjDM0st+VG9ec4iWOaU5Cx
Pa/qJX1egFTKI3WsSMp0OIVCqdLfDhQEHxMQ1uMByzZBZ//KCeWtIhqfTekok8QLNL6VoQKuKCco
R5+y+4rSoMgEFADInKplzUsSU1sWetkWG9JGUkj6WMlvT2KuOZX66w/UHXm8AOGt7AoJrAkb2U7n
vdhej2rQnlR3yygrZgVze3EI2YpkC//iuMr/5oRmpaElw5SqneHfy0RcUoEdsrugRf6EgwIe+FYK
N0n4/28IgtNI1Ulb0OyvOqWuYZeSSPOx2EJTqXKdzmOKvwvT29UvQW8NWanc/WMyGiPJIH6MfqDp
ruiVOaPdmM9lsO7819IQWdKNDidKMpGubS6ChPU31NIzra17xCKe27mYl3cvI2x7pWWymxZAtaQi
GBHeGgEcQ/0tbxWEVwz7/RA4CYIhNzKgyKr1XuNBlF2hb1OqwsIL5tu7EMajiwL8RgRUSHLrJ0pk
RWilUy7S8ebStErq75x/c9WvccJQ5v4sdWFktwHiU9OQbXAlnGn3wD2pQzseRLigqRdof4pta0GM
cyH+1sgKCHLVykQXTCbt6di6oezLyfdChDxAfkHIkXW8ZfAcNdXFVAS20rFsshO/JMvQDjIX58Qd
gfU/esZS/xEE4J0fafYU+fyA+0e4Zx5/BssrzXwHV/4ISkFNJw0ipFAt6ziN7P19Psu/0QAPOfa6
n9iUk1SvNsqfGtuc6WZoKfl7qsNbP8JanS9D0rFcKNeBf1I9jJBLvIuQOc8RTmEPgSyntC8RUfP4
037WKf3gRzzrN/6p4JlojINBq+qEJDmHj4UU4XvI2l7MF8b8jkcPmpOhDZ7zWyIBbM0RX+vD3Ren
YDoXiOjD3mrSwAtWnOKR/HeTNqv2oRQJRimynp/nC2jgrxyW+ZmiAaj3dN/pHvlnZDqYgtIunhvv
R0QK0n7kMc9P6IXoCLk2iK96Lo8h/dGgutxv9ypWYt6eEvBfGAgAcgMMzu7xiFxldYDHcYjemXta
YK1Sy0NKR11C5RWL9UXTa6kZmKJy4dBYkkiKwPCncgLc7elLyEmA9/tMBXmUnhaqJ8KzBgL9jW+J
0lgIQE6TgaZCVgSpeHMcpBGyU5TORYAWSS1JZ4NJRp5DDAg81VvGdYuhleCD0ApQJWIUt+Pv+fdZ
ANrHQOUwycPfk2V51xarzsh4K2nuomBDUcsDtpfJRYsKQwuGvbkfAeI4s8UVkWNrEdXuotsd48i9
3nReyrjYYzcaQ+Yo7axWhO7/zSjjbxqundxFbl2GhDYIMpOtL9l9wXZWp1yjPdHvH2+aaig1dDNP
99YhnwSJa9lmLfLuA/Zhy+mludOi2rUD+hgDPSPBOr1MDkwnepCB+nRIP77hbqJg/mJ1JLCqpMuY
STSM0eRTkrZQ4S/SjbAG3HAp1BpmbnCBv5wupzmWVBuIf9+aTXZrI3e8g7ZjsNjJ7PUZp9Ko3mEZ
lXwBuIlQN57dE3AZwxk9BGhnv80VUwbylUJZnoqbHxW0YTXDUH/KehccdcRYewF1WMc6v5/JcSQ8
1b8iXkIf0OhWMw7ubsYK0SAWdxs02IKKyv0M2r4QjWFzc4ed3E1WePO2rIipDL87bKiSRvosjMLj
PngM3j6FF0FV0lktclXjVXy0YYbO692D6+o3QWwJLAT92ZBy5udo+hcM/yanCas8YhnI1Tj6lz0N
zLAftJt2KDQDKL+BSOsMbQrE93uFzCpQ1UXEp9E9gnA1UsZBYb4DqHc7Y8Af05fH0hdc78rrYYWX
mqD6SlePUViWmglDxHtDFeY6j8CCAm9QbE5Jy1WvzsjBiBddH9VsDLTq0v7UUTu6DWYkz2sh6xIu
qICIZ70/kLWMFyMsX1OqtZhSKmRqA3dMbJRVcqEmlb445KAVKfhmZIpBWlx/4kwiPpoQ/zhu3JxO
SOAo6DwE2NF/MRyIJ/wm0x2XGcZQcvOFgICVeDT+bZ8CGGhdK4iJ0sdZ86LA0PeQxCl3FkWxjcvi
aPOhaW89KgZj0IFGz5w7+fwxK/XwXzU/C0tPlc4DRveH7pwQ5f8/rE8wExV5qL45m18R3YClgSJR
E+vW3AYvFOY+IoMA/y6hmhs6oIqzMfzqCoIIYagHVtlIfBbzc4Xdtt97Vt2r7Qc/d4IOEL4wwYe7
a857euoOlFhiAbYMdRhRMxIvRitQ353iSV9bFO1fJ0l+N20N71xSnO/P1tpZsUUfrZp9NaNfysU5
b3YWS3kKWCemJseDAezNJzqMKuF+E8E5ztI4+EKXKgJGaUdx6nSruDkY0lAS/ZLSLzDMcV2M/iZA
8563A83TR63TOGvyxU1nq6/i2Ep+cBR8M+foq16Rv6TOIqtEmhmVcQeGH1NlI2g2Ynh8vOVNo1nW
e6h7JmRkFrV+jh0TB+BdGI9j0KYpJnvXTemcPKhgL1kcPP8fdi0euTTYv88OOKUAnxVigEcex6LD
ST2t95bbsrXdOKoVz5sU1n46ArnCuUe8GI9f/7iKHeLHWzGasDGUK6IH5S94SU0l6gR+OkGr7ibH
pSJ4c+nVIeu/elNOX6B/flDyY2hcqYbrBVT4+dws52segcepXMHs59bJ9RobRdcvf/dXL+LUAOFl
Z3ht419FfxQPPJHjFzjiGXdaeh7NxgYGJICx6YA99SLvniCFlD5AjT5VuZ+KN544AXUrUND2+J7Q
0hDPYCAF2QL1fFeezXaeaTbROB+fBvWk8G08N5JI4hjNHO8l4cjSGawypaGwI91xqMnu/9/QWBVQ
YjCTQpjd2vxJYOiwhBvqxX6m7kD7D+2pqIYOPj84xERMHk1XV8jOD/LSczleyi7GISAORJsZ1PsZ
lNonNQAi+I62hu1d6QTFC+h5mWzI4h0QoxXHjf5ZoYShQRXT2JXvCcVkL2TJA9zVTSFrKfgsnfuu
B28JcBB30QlexCw0YqNROKctX0Snk9HStiN9mAbCVeBc1tFApSkWImK0FCZFNHsA2yAfyZRyZjQo
5EStFi/6rE+0KHWMjUZgVAMYwlksmgF/q51FO3eICZeNHzvj3Cv3XLwqFImqWJU5vUp/79lEY6kv
yOzLaoMXb/X0esZCuKFQNk9FH/O/Hq0e+2zysINvVerLu9Edkq5ghpnJA8utOg9MgWOoqNO52A5s
EUqG0vY8qMF3+nu1pc7uFEu0Mzt4aKaRi38rWt7ix+vIX8sk2WE3It3w6aIAd/qRIlCSo6cBMrpB
1Sp9FQeSqfpLpp73xE2HAXkxarUa/ICISzrKxi0D27yhHAnsmnkzdh3VEB94LaJsZP8dsxWZz37e
NXfp/CpUA8LFQQMCKQSfeHtmY6IgkLcSqqTMoFzx1/toMrg1neE9UOZMtZIkZUDvPP7JqlIgiciV
YLKxcZ+s2K9bV4wpsCahYDXrNStUZcr1bJ7epKCACk0rS3ZX0mkwKSaiB/aM6GaB+Qv52tFUnPqU
V6TAX7HvafvXL37cY6PGlILdv35FzvYxyzIvnZZFYSAnDdgH3z4B6KOGM4xn7ksq7QxlLB+lQVlF
TJpx1LSOpCt5VChe+WpK1oXeLEkw41/Dk5kkSKV77xyXWby1C6B65clhCj6V5HxUAFUQ2GHmFs6e
TCg7C2tqQDJuKdgKdWjE808bfEImgsCe+U8C2xO0Lz1aZuEgOZOEcoIAZtL52gdVzsRIL/3+r0Ae
J25r6gRBe7C2wBWWMznyVrXbghU/izGrsBB1XDk35PBfyg8bEg2DY7kb0OCDYlXpvLy/hSQe4bDw
uJGxeTHFok1XdwFEP8fyF0uG1/igVRMN5XKuq1jEADCnh3f5qQ5Lnt4Sn9LIzKha8oATm3dzKGDy
M+e81CUj2DgBaQY3hY2VNd6zbvhVNsssOELsOEAZCTqfvhHysWBYkOSsa1CFxvJCAs7W0Sn339+X
5B63SZ95fkIhkGKyQzYXyDKuTD71WLHVEw9It+MBoA+2Lq+XFUmDsiayglru2F5xJnlSlcDYPQm8
+7Qr1gxWAYfpxgnrM4HA7O3BvjE1WK0JUqv9fY8OCJE5HuAmnMxpubj3hr26PH7jVZpDO4bGTdbs
7T2hpWR/qooyX7yhgtgyqFfHD903EwED8PAqPGdL7qd6013Nt7B4otsMap3Or+0uo/5sF8e/d68M
HoIM8CP1nTTxJwIlW/NIYWTR4XiAQvJkzoPd3g2raNLYxNE2X9DiswcBbPY0rc3mSe/b9HrfUTn8
DTGRc1LSBaXH6sRTzfe+2Ywo95RUkAHDyEk7gylvjdS3HrpwHeWHXpDfZKZXMiLGTCOcTFASGwWV
k1V0IIR+T0uXg2mC/fa7ytHqGwkhAvlVHFb4Gt1l9LKRrAUY/i9y797+J2y++4dyXGM9dr/DXeH4
83H5kX1lr2+cejiklVGv5qzMXUrcvQjZfm+9lhJHJEo8aoKxGLa6KpL0kzfqN/P7Dj7dzOmuFCLQ
iNS3aRnYOQyWNKJFmzv5xa/xi7b+wSB/UxfLwdRg3zLL3cVMO7aEK782XZBnWI6R910ptvQdrhi5
LBfxmKxTlFHoc9TKR6VmKvhp+EjcEn8ER/X1yo03EXoRFY/4HplhK0W732jvrn4Vkmwy7XJ3FMke
38XDCU7dnxqN7VQEIJ3VAnKWKSpj5AiIwQCLb1z81iXqgKwjeui4O7Od/4mj1YSxyTsIOiX839Fx
m0AHv9zjg/y5ZJBQuEdzc4LWhYg+rooI1UatGGzo2xAIDx4OougKn3kNOwcNQGu7KQIcTjfZ5vD0
eDvpy94Iu/thUcQjQzPkiGFYPXRySTbGEj6owY1Awmm1/+rPXB6lJnwnSNJm5HpPd6QT3T9R7gLr
khD64H1TPbHan459A8F8HCaoPDoySzoZYmdO9V9w7pfUaS0mhrpiCJkdW+sG0kx2DhGYGrn4Cex/
bR1y/9lJQ295aQRceoX4cSEoczYrhMictMK6flvOoO+fuaLYgy99NlZHD89JpjZ5MlqUkwZYQxIG
9Yrj2yiTVJDGx8Ue1O/nBZnrPqRdCNcjoA42PmKUxSl9CJwcoWUel5kPEuIEs4Pih8+mcwgbBrW2
qt6wxEPljKk9DNJrSfBD6f0VUmZkf5R+qdN+3X2ZqlEPTmAwTyCa239IiXGZBGngbrgyEPRd5JaT
mZEIxqA87HsFj873olQ+2YOs/JYV7lprSWkaAz+R0IepeIAGNT4mXqGAUWkYicPqlvWTmWviYhcH
xZoU7ckOdFr94bLEOAMMg4T27WiXdneqAs9p5D//xdAJwgfpSGfg09aX60NlNhYaQTEu8P+uB0GA
bzLO7XK8Z6u9niOgdDOKPWnP/+mWfzuO89ZZoIibYdoTZ2BG8xhhuhKVjSTKXkXDXTufNu7jfv9m
rpzESBD8DI91i2uaEHc6ExZX/DwXQM8zE4J2zbDPDF6OBE5ej952MZbitj+QYZJBhXmIBXYkeGGZ
W5P4nKrYSqaFR3QeIu2P4jfIChmJnfuBuPojpjdBIk3/J3hO58h7kdm9H/rU7fFOMVnamvpxcXfq
GJZPgkCqBCdx2ectesV5/+KFy3f8BYFgi4jHwGR7VQIOkkG8HxWmak/8Ng9OSALi9XvBnTUAWcNn
xzNo2GtKPOUmXHmPRoxBdpZQxI1D+fx04urmAomsZE6GK2UxhIuSK/BKrUxP11rxVJ658KtPNs2L
p88D768BcGQG9Llu3AIU6FmsmIoT9lQ27Mc9SvjDNUclrpHEwNq7cp2UJXrHHnsca+Gu0b0oFkBH
qjW2epiUhAlyI38o4LPqjSmIMEnHEBjczwErlniWaEXN2mipY+oJ5qgvttZz6I+9ZVxtmpHmLtIF
o3/aC898Xguaqk/xiC2V2mgjNekLr7/53ve4agDQPJYShpL7Zsg8DqaK6cb8N9gZufyTJBbHqDyk
QUcIcT5CYM3hQ9jfE0Q2bI+kL8hg7SRSvQJP6FWHx2SJE8ByDeggDMGTDu1U3SWc8Sda/kV9MfCG
AieJi7+KdbXVkBiIXcttskcvscJBYRec5q8KnyQ/sPm6fY7pA6Td2hkveZnHiOnJrT0Ufze0QuMf
NV/K1VW9gBivrlZy4HCnLfFTp3bndAQtkmrFzaG2ZAkyKo6UMAYaCNP1bfMaceJUwRxeN5V54hH6
ccq8mbSL7/g7jthmicS59xHxaDUPzeIZSL9ra24/5IALvDgNT4+gbFOiyVxcOuJ/GF3Apq0INrj3
MBE9lyo7JPjrRzTPFdE6cASjV0TBlL2kmWs6KETr3H55iRTeJ7lup0+WEGyw73kDWR1Kjy+sVrSR
CBlG/eD1xOKhdGyvNwuUhxhxQ+rcEN1XHHNGr1Kof0c0AA9uimF54y3/k/ruRKWRATPfPqdTikut
vqrlNvNnTW06tKktIsQ9Ni6oSFjOACsg02o3LJNi0aSIcxqB9ffeTJCfxQRJwLV3jRrWlDWpNfbj
6ZV1f0+78uwXQJJavUFqoruJUFs+GujGQ+n7QQGIjyxLRSAERSdSxHkU4w0+d+hbSepp7sBNnrAz
VgetG+ExuttMhLP9C9LhkJql0n3HoyV0iSHVWQWKs+ElYfoKhYyJ+9mqXFuG8k3Es2jxiPdoJCQA
z3wDjE9S+W9QsOoqyvTpGZTnYALjt4Xpxt6zW+/aI8EOURPSaKkfmZC7JQ8hpxeCoDvPAwV/qlI3
kOUk3sVLS6zP3sjrl1eTrxmqnvajwvkxi5uRetdd5ABoMpTQVA6N3g4aj73KzIkxeaz+O8ldQ5Gp
TkaC9g0hfIWn8SJJZKX8propy/P7BcW4Kscwbe96wKGkfTHhwnK3DFRypQuwlxEVi8haBJIBJoKb
aoHs7GZpLjDf+q+qTapbp3sHgeL4lpWbawOJOrAPj3EHx5fdQabtKZNFO+IWv6m1EOMhWdskdeKP
HacjW0CyFxE3GnRTA7XFcZIOBk56eBrn0xA3CVsw2N4D1Kw1EsZ1EYHNLYIrjf6It3nrjsloroBV
me8xYnlklLozxkbRb2wRSvDMeRQU773s3WqPHECCtT08OwzZIGnoUu/FrBg+IGZHp/lD4c/M8VxA
2HNQTGGC1QYLk/WlpedCGtGzSxa4AnUAMrk0kLXmaK9ji1ErXKmonihpisuFz9kJra8G3m8C3/pe
R7U9bDmpYqqnzJ/5jsRoHcDEnyB2VcRDCBKv9Qxt7O88g28Jd+QBMOlMgf+houmbrpKsmWZTzgh4
503S0Da75NHL/N/C6ZLOaTbBcbbD0sQx+TQ1tTPpB+inopFVc6uCHZqOIi5zqtyVS/GSi3DRpa1m
e0T523Hz7xQxx7Oxp1zyilO+oPWH7+7mgW5FEXzBpnOcxZOdMTOuPa6gimZIJAxu37DQ8j3XCNYJ
iRAR3V/J0g7yrA5dppTizZGWOBq+HwyZXcWVGYDpTB7B1Ofz3g23KxynzjWp3Fc7D6EBhV4W7A95
Kapc5Kbe7VaQhq43cFrEr5HYlB5goNBah67LfWZs/37rwvgKkkKC3Np7Hw3fZ7RTXnMsVD5cF8mQ
ea1mNR94HJv9P6ieDwM6ZUOK82HTDdRuGo30kbEU4eFLiPoqulBSrxit22430wxwut62KPC0tPX6
+dL36IIn4gi5/LefaMTX5IO+KPCWkaJCKjoDX4AaUlweRBe64jmiL+OrXMdOVumiQ2+nciORYMAV
Wo7yX7C9Bz8t/75xbtBiIaPlBnL4bnFDCKxZHSDqOe9PrPjx0t0eF1WQsHl/Nn+3YCgiv9U2mG5R
U4OXZoagfcoEnRo9nBU5R79Qe87J6fEmD247N8Bc8pptUnOWOeS9xE6AIjdI8tDo1N9GEazkhlw6
MwrGsq0tz8uVTmopgxkx6V1NN+7pj+tzJUZwhdaIWgXAm++aTPgpEwMeiR12fEzcHKs3jLJwqRc7
+zVgCqXly6kGGiHKF6nI8t2R+Qqobj0Sb+oDb8Oj/msKFx2m7Mzhac8SeSStIk81ZODs54GVHXDa
uEdGOLXpQNmGH+hsxS8/KMa0O1PMjhVbVX/02+Ufm/mou75eu32UvGyJQXzfe/B7XWJPA8Vsx4qZ
L2jN7wZGpYDdXdeD4HBOU7Vi4voezonOy2s/Sh8lt63zFiTirRwvRTHiq2OApeJE0VD8YGtjw6y4
WzhCvL4wAZP890tiDWTiIU6h47aSjEPGKq/e20HMNrE5QXn9tFstIO+38xE9Z/MRhXJRRdSJIB3Z
qek3aTEX/mCptjwQwTy9M3l1fEBGfV4qG7zLp9yAIA3mwEMw56AN3QfpqB7vYhAgi6YL2KRRc2nN
uGxLsaVxLplfQRlRRM+2P4JdP87vd2aCHWMLIgn9GhcNqgN+yPgLgJjVdsgGstplZOn/fbdGIMGp
73bgAFUdRHt+RxbakbNqbPNrAa8Os6SBNtuF1tbrXzeTGtRieKVL/Hc4GYzP46EwPQc/Hi2WeBIe
J+wSZn/+PcbZQKuDTaDQJoGtoyRZXAUl4RacNq1Bs/g4ze44qL00l+xScWCHWZ56QvRejuhfeAMJ
7reT485xWy4/7kWw3LvWTkZPP7slr1KMPeBG82fAt+f4EcdqHGMqyH+X1mRzXRRI6Rbqeh8f6NOH
PAT8rHHUFLSHJzg7uTcR7qXtv62LZ2jTHZt5PH35udoVRILH6LO/acn0LkBhFaSz3NyNPYIXzEza
sXFmxXw/UgAY9tTXnK49RtEaUS9dcKCcxMiFAf/qgtugikgbRkzeow/RArIrNCONf8fMzToPYaIG
cIYJRBb+WcVwTtAqVwWlqrRr+xACGvxWlOjDCbQyforqHlNc1GyMn5wlIUkjT2na/dHel/9nxgWP
1dlOT8pf5yHgkG7uX5O5KArDjla0uMf3cYireEDjIGSJOgA2Ywq/Z6tDpH+2/QuGiCvY+WwY8Bxg
ft9U7vFq79KPCEAwWD7tJx34WlaFarzF85Od56HJkPRuZF6snWIxAzEfkkOJo7rbAG0cWkex1dlM
39y+ldrYG4o+Yzedaqr2XWmYAQ+GhxIr1fmuJo0DDwzwZGDYMmJvVZitPu+EaVUppEnwmPGe+FES
eA4frLs9o/yuJqJe+PVRwqSkIZiAZcmS/u/Wz/xMbGy6sGd497i2QCDnG9oyrUwLedpaq/hOkPnf
sUDAwxxnHQv36pG27E4xw3V8/J0dDVcZ2mNo3KVbQJmkC+AdQVBNLoYlbNEsTvJ1te8BPR37PANH
JLmltXgpyQFtITp8EsI8v1ZPuEnU4kU+idLQBHCP/v+GCNxTFV7Z71W6QTt1wAYhfEXw6TY2g6TG
7YdL0vq3eKj36ZpeZQLgh2WMRiPSfFrYnNzHCwHaciP79/NF4G7X/KA4TcHTrDpzcUGLZi76iZaI
8rdNFMd/rB+0qAFJ8HsAm0VtfEKvyeYOsxIr2hZRDCveqn/x34/sEnQwK0JJAXYOtdgxnhuiKGx6
xOcKrrZziw5sjfAjV74inUGTapoeITyj0F9hDFGNw5kvFgKwa2KNkIm07vYEmLoVeHhly1KymxXf
pXXwvTB426eVh4hsLVv48z+20UDi2nPll+XsxZbyFiiV8vIWkLO+VriU0swmW7MIjnAAeH/5Y7p5
olf6hyNFBT/JCgqP5BC6amNsx5c4I4spaSb2di2/qJ4C4eS+1Dwxv7gBRQyRbG1y0/j0ySngXg/N
xklIOK8FhFA1Noxw53oT9XaMgA6HhtcJfzHIz4B/7nb4/raEAUjJPa1neuxs94DBvlr0REtzEG3k
SN80hUOgl9iWB0Kh4v6qBNk5G/c6COuK3r2cGsXA0G8X3nItetmnulKkHt1EUYq/2ODPFhofJPA+
YNPil5mB8RLcvT2aTsxygmBmYEA+T0qY6rMXolQcveRXA1c7ARV3NWDkwsBU7xIN/qSf2bdv1cJK
a396lbhR5cv92T0t9i0QlNzBQ9ywvCHd/z86kb4tp4DiBUmlzVj1ETWmZC7pefbM26Rk/OOXPYO1
xlxUQPdhBohcRX3/fVogms6WEKTkVa71fCJMk2wJsyiO7BuSI3WN9zq9a9jgRtns/eUxMjdjUAfx
tUhF/bc2z+SiIbKsDwC1fdGHFedqlHsaVBwXBPS8dF8h1G3fzGrASBHd6lntkl2ASdCuJ/twnoxc
dAaqgUl0hkKmaUXEw3+iLNdA/rKa7a/JnkmGCHx55trAfEtQossWyknDrf8qTqHfe4lw/XSDl4iL
RxjDeb5fuvkkoj7L6wI8YkJIn6dXBdjI+I2ricpt6FwNA4FuHZz5f94I1XMfONYPXlC+xpOxqQJO
UH6kswhn+YJAr43lR8Zj0ov8ZhoeaJ4cBn1HjE4xSJkclWA2STEO7OtWXKVR2M8mwxc3tf4R4fGh
IC38Tig9i3WrCv/2ymUvt1mVMev5bQjSKQADcORxNjfL/hCFz2tuXJ+oDtBF9GmcUBezYjqXi255
5HHmipNC1x2cl91GcfuVkxLp6e6+KadVaGpR0hDnmzfaKX60uiAffRZGzQVK2cctwYC4x30oDQi2
+u61PoADQlUjmGiQNjnI4Oie1hIC16UeLopZBDer1aLqwRqG5vVGdvPxvcjUNC7ziAOtzf9jfDtN
scEiqFGJBXqG0ZOR5cugXVoVTw1GVleeozBqp0Fs2sed52pelv4HWqHGuPeUfohEVQcAPW/kvSFl
sS2tpOOC1b3veDdrjxqkI5Wr4Y8+Vb6/6hjbNtyNNzaAMiB0PsC9OAGMR5XdafNMt2LHwbWlF29b
J8D4jpqf/tlCaCLYIijRP2f+pAxisjeX2vLvp47FT0t5hh+XOG+Hb1IeARh/TafkvkukMZkC6ai7
VLPPKGZWbwSTwNPgyBprMbHWG0XXLl3etebBTcZb6RRbF2M0F0O++E5BEgyemfYo58j9gKFr5mVS
XgmluvxmIPpMCOoSRM6WTFgu9pNfwnQUMEVm9vg8O94RdSL8fPL2pHdo6TFSwQEH5IO4nDT2Gsz0
H+ZLeWOOREq18lm+EN1jCPRUi1Rc+B5T2bLmSJAyXhjGX32ST84iNZnJL480bGiwYIygAJMp0UCu
fkWKzw/1rQAFLNNE9Dk9g5vrLiQrEJqtEvt124txWafHaqNBRPUkOd32SWh3Pv8x2cY6PiLOJVPh
Jp5BCtRGP7hDuQ5f79AKukCrKZ+Zol0lwV98y4WdXB7uoqaw04Er9uFXTXPdP/As/KQFfiz57pdZ
MGCVSxg3ZwWuyGs2VW13Oc+SRnZwTCTpLsgwYol6UXxbpUyARlu1Whj5aat0Id8WbZX7+lekdEIK
AhLX+jhLWm++3CSzeuvZ42i5SogBZ1C1zqj3QKpFgldpFrX5raiZyMYDOlxigiPNiAGsIYrNKYjI
xMikSFmYSTHxUs4SQSZ2/82d+ah/YvIDkZnEjjN5H7kWnmpe1+y5w8A0J20G5wFSMgUzZlpfbHta
zDl7Mhc0A4qTNWhJtNUWiVEygXhwKxWe4TuhJhiQEwmAdco8Ywv1qyopOqidu2rbE9xAEdWKDkZh
WGj5emcHzvSpBk1/9OHp473Pm5/2dVWqjbAuF02AQ/wJ/pRZrwTTcAsFn3RewLCMQFTIE4yWpUDD
lEPdQ4xabuZpFZtYPjzonHvtQ82Y89LKtIgoSD97yWFOLLB4KDWyjWkcPhvuVGzNKreJcmrntdU8
/EYk8X21JE4LwLMNXrbtVf6T2FEHyuROGg5lrsX40u+ja3V0avrbVUy83cSEXn2ZY4+k30f6BZFJ
p2d0Te+m2I+2ZheoreyL2wXxsWtsk2aOwgCL4t00V64WxItkRlN4c3OEcKuDUzyRvueyxdBiBz94
2zMm1cAbXsgyjkWvWHQrroFJsU2fmJDgKvk5SqB0skxwPxj2bmgVb5DPFbXcQVH8p0+1o4bNVXuI
2ppLEmSsUpmAmgZeefuWX33H1L5tGhgOlWaco/GJv6Rfg+vLA+hUsjbH3ZslsA1ZEcfD4a+BwWMI
Z0T02p/rQ9aU1b10JJCeDOJvcyzsfEXPBy/vnE1sq5/3Ar2qWv1Kaoka1MmpVF37DGWjBYByr358
mQgaxGY7VcfiYdtGafDfltj7E6zk/d6U6tUyRPm7WxbHy3yRaifuPvgeAuU6TRog7Ag5SGzOTmn2
dh4ZQubqmxr8bmh11JJGVrDf3EMEJwxJpVKhOFzrfUd34Z0UzQBZK2qq4Ll211oUtEYMmtk25Go4
Fg+UCp8QvITjxF7/0vgp7I12H1xdp7nlqgVV05Za+wmYEJyTIKLXDuoWbHnk9/j++IaX7oLsdSlc
Y3HLxpb5qmzOO+PEApH1jLHkaOMFA9B2mg5tSuYoUt9BcuuSVj59CwVQ9pMgFJT3p0I3KBDj8Xo7
bcFoh4d8FvdrPFRXMQfOCvqtxUJ9gbqLEYmu1K4na5NLhzssVB7bH4/ZPSbqb3YHmqoiKSaBGtfM
bdZ7gMEp1iSoEP67g7c1EFYTVKEyzie5umP0wIyjJcVFfkBOSoWmywg/vwbxy6UfIBVnI+WddM2Q
vzx0rrGlTscT0YdkfehIpNohlF1JvvzK3AnTroCfORTNu5tdeX2k3LNgpk2V1HJHlBjnhkC6XphP
rZ0zRVsyK+kA2wglyNEBhIysc584658hKLBm5dO2omIMuT67hzlNinfNTJ6v9hdKsODLZIG5YatV
b1B25SWDwvDd0XEFlL0K2FMi20WIOm6HHRQLrL6R8cPSPLce7/lCrYcD/sd9TPEoGJcLH/MLy4FZ
XYlN/45VNecOdwPC5fQ/s8rQbYlja1HOvquM0JwiJFWw9qocKsNeakn0zznnjGT0jyvZlsHeVk9H
ECugNzSYdppIbz+zWXOp47cg6fy3CVb2E/tbEeeU9Lkg7+QzjYK943J0R/Ex3JUUTNkTzCB8tIDG
L9G5Kkkz/LgCclM3iXmcVk/Ayn7svMJgfMr6Kkcc/zt4/2iPr3TnGGAvgSLpypI7z+VawmPcxjEJ
bHfKiAx/xOXa1QGg3gRyr0L7SegOi4cmsda5w+Vd/3MnWqtBoEoAzzYCcrm+ZQkHkdNZXnrodKFl
kQ2v7UJwHAN3lmtOZYDHfVgoKcc9zSb60QlnQZfRFZ6eN8xpAXLvWZI5q8xxPvH1MENooyzSn4QJ
6IiL2ep+EpQ+aBfR9ZfxpL+5lZVCTlKgsLMBod+VOehXRkYz5WoduMQLrEIMYWZWbGS3NNj86OGc
QR/yy2q+JmN/e667HlmXHPKdy6I/q5yq4WqwpRhFX0j7fWkluiEdYbeznhNqHUg805mL6SDQ0fkp
LfjsgYGYj36IaUI+v8/3W+EwS2AvKKkoPS6zi2f+zOBH5fxfeXaaLlxXD75g0qW3sltZacneeQNe
i8uNIHs+/DzAfc64HA1m7KWD/C513oxnIUl/zV/5jvCtBKZB6Fx8x9Hu4+d3is2GCyksKjqOC3rB
HIUlDPhdk+YFh2FtgxxUktm3rPLSh4dAdxSLOjmFhGz5gJPF3oEAKXEQ+0FLTl4BAN9h2KmNKPAE
PqkD0bNtQKjfF8PcXcZY1iXeIVQxdlcmW4wT+h7KacyLezUP1RQLjdRQ69p6GJgwy4C9imOrBSxO
XYXiBLuk/VVrTcccgTzHahOrwl+DQzUkS3O2dVQ5Bx150Kc/k+wG3OCSlO2QkvkbKxo/slX+NvnH
F+B0m4Gr8mN9QzvVJLe2NKGeXk9Ov+bW39po/o6YQKtDl/KEzwJrVWJFjJcDNLT06bzc+AtwZSe5
YKGSXSe8EKYEWk06uOIHa376ZFWJPDrD0JKdT/Ab7/xqxcfX4oU+Z2lrbRSN99I78iVrulSe1hN+
KXJ5sHUhYy9s0JvWQLqaEu1SztL9T0D2y3oIu1tYVfYFgDYS+j5se4peYrxXT+mPmA8txqrk5Vm0
iF4gyxW2mP5NjvMRSYFXwO6w4OXr7FBUaCMOJLMbh17Nt+VqTG+tCrtASH02M2UXY77SucFRCMtq
K3wzbT89CG0C0tx1ymrPeTOvVNCrqIR/ZG5iZlelHl/WkyjcQl6JFX3gjFkWv5/dLoVBHVBDqxMy
xwk69VueiOAKqEy9nXqZ9rjg2GFFlXCHphDZBRhGad2xVQ0vDQbRXGY7fPj6jO6S2PA427uFqaoO
XxzddWiWboD8WojeGkI8lh6BGhRSc3PlyXO42RN6SGyrjlibKT6AwgB0+KoV1H207irzpDylTFFg
sY3KkkrgrJ2haqQlM1INXlVZZSrDqSknEYWwg05KhgxdjDkEgUM2pIIebUzNVBFA+frYb8WE6Mxa
wP29dOe+GrR6jxY94Kk0iG5HHNlwjrY5goOTlo4Qd8goxP0F+MiRKa4JSbM7SJvWrQIRYx71Qj3c
nuLBvgC0Q36cXsV0L5LHPPRExDIuW+v4ifV5JHi8jZ9g2GCG6665JKzCUdvAcseoAnzrEzJKKLpS
HDwN4d4nQP6oW7RzNpU02GzUGW7kI5pxMZOIeTTTEsSFUczJJS2znVO7S+yZPHcNqV6HVk+Ir/YO
xAg3y5Hogk3jSoH3ygwwnNoJBHb3068e341FBUDaF1bDmied4BBJq+uNBxrhvK2AyihC9/ZyUo5f
XS3ynmvnh//aY0gI09MUNa58AEown+ltTjD27ZjaZSWmhYhtUGw1xdcj7hQBO5DwjV/INMci7NPF
GLtfXrWj028io4XSQQkZsl1CjAHEdJKwqEIC/NiSyuSXXIbUjLxJCBCRRwXtu1eQqn4GcAWU54dH
XsG8dTYTZQEk3qRPzJwOhnUIyKxXoM3gqnn8K+OzoDRdFR2Hsg/oLjTU3dqDmteZzgwB6HKyxRd0
KbnNKV8UwMINbhUp3jAp6lXAjzGoifrfqfsZRi+70xl3N0jFwCYNtOBPimc1Zuir+74ACU4MtfIi
4qi3FLUWXqtKHfiqggL0ZCwj+mmbZ43jO27tm/OtplOF1YERAO2txLnF9aY3yZSdY+tAc2Ckbvae
uTBDcGfy5ae47mWgM1mxf3DeZWFPCkS/vn5ZkLJjpeYg3ZkckVXeAAtiCCUZD3eEgLkfWnz9bPlF
xD7K7a8v2gSmdOEgOBGAQlI3TNr/WS7K48qDR8vb1MSMqoZVQ/7+Za+dpCPM2ASbAILMnqEYz5ui
2BAmWk8Of7sceDve/wHAC4RTC4YGVAGxBb8EYts1GgsgyxHpuM4XDthl1+Rk/nAflHfGtmndf3Xe
0dun2jLLDhs4xUr19KlDMm9rf+rE1IMSLvCiv9H7WayFuFzZUYjN2aE/YSPXkvtte+4i9Mtf4/cc
w5qb9XkPXSURan8BGATolUCWaDJKXF9bink+1ePTggxM8BKJfHtgrhiphp3clWOIKpSS/fE0QZ0f
fP3jtIv9RdKd/am/1WLDeR044ZXBudd+MwVn1J2EozZyaiB0ujAsqs8nlPsX5MtoJ4F2oAUrdGEG
Oo2WnrMdxavY7dPjBFLABTpade81IlHo/I/rhcvzlyO1pWomLc26I+j5+8+YosqggkuR4OkCPxQf
CRIUcyfGybICcA2mUZLNxg8MhM1Pl6ZhtlqQ9snFTeOpzP3bPm0VVq2NU5NvqwJoSxwbuY6G/vEO
K9f4jCoqnrDN2QkZ9ccTa4fFd5K3fUomO8rz6+mr0WIaY8n/dvz0O7z9fZAOjSFTwSIBkwY6ULju
QfAp62PRXg7IalKebNH494qbbzmf1FSbEP0VX5ptxhGjY5C5T76nxkB7cU1IjukSjbF1c009S8ig
yA67ACaHcyXpRFdSfFalsOX2j4S4WrJDOIun3A7a20OiQkJJc/olJqcJj13M4X5D43gFAuv7M8Fy
8nOdh/CBJ6oSNSU+xVr4OuDFD6lnbWu517AOQqhkd6bqJBjFDvL0m1Rt1qNFhOkTq8FcS0uIejjb
A8zasJkBThTlfn3qKy5krm1PTQ12bVK0CaSOeVKb6aCeEe7eikPzgRi/PgDO6HoxNO5yi3eTtZP7
Xv4bQBCAmIPNFJHEASi1rtaphCOz1CRJgZ180AVSF6CMWHPUPmCutS9jM8584y8EkY67+azyjqL0
uw6KNjSbZ54afPInr4WO/GOHHAPnEwwCdzrFGZmihBHTT0lwFn7NMLT819OU93k/Y4cZKvkeWdWE
VefNzE/uA74wyf76iDBSpfQH1S30yhyG4UnTeIJuuN/kGHAq1NRdcTeXpIwnD20UIok21jMXLrYn
8V8LfLY2XKAtZ7t/irehTszhLyWRWkSFOshbkH/8I5A6hVm99zHTd9ejUivk4HvbrZZwpjPnLFfM
SKoUkh0Y4PyIZSysuo/3PYkG7A564kbw0q+8qEkXVbYbwRSPSwhonEp9vXsKPdFK6W0VyDm3zXAg
l60REJBkqOkRVTjdE2Y+2LTkPefbjp0kYM816IeoJ4Yg76Arst4j6fkccGrbhrKKioB+xEj8b8nw
LXpxDCepvsznoHNFRprJfzLetaK8m1S78pFLNHdol6Z4BQuVXzfG4k+PQ7Ne6R05eW7EMDFqQtPe
CMtymjkRi4PSz/2d+2m26fBDHrZoBFiZV9WJe78HGd/C1vL8WUfn+Rm45YBPvlqKu1uy/mNl6UdW
ngpwMVUACZPhXBOP0yWC7bK5Hty/EAkk2K70/ddM/WMdpDrudFsFf5JsIAXQyQF2Y2pmzPvJrZar
gPcRrsj5aawpNSo4Ja9Luz/OoX3alVDx16yz8Snfoxwq84XsbMuNGoVwJiL7CEUh4HuXLChNQoN6
LO8QX/5Tl2CyLmSvKoC/YMP860D+A9kPF9eIq+7SFjOiomufhvh5Nc4GaevcIA+cpcOPNh60sOi2
cO5TIKS6JOfTFDZHLiz1qvu/txMTiVV8K0myiUjx4TDramKz2irkY32Ee63sG50ccs00njF3y7Ub
wQuwVkpiv/aDvEMKWMIfwXjhBZrdQC9EYa6F/Zi5crBzc+xv8Jy+DTu6hbTtCjPCbvBgSs2I3nOs
n1UnkAOaRXp+ZDQiAVAnPimIpbt3DDjPA9WMx0M5+JJT5zPC+KtAK6E57pM1i/zh46PZa+o7lGJo
2VWNVrQrBO/gdJpvA1Mpplw5B87xxvcOxbnsP84Fc8HKpI6zSsVItRM1VCDnC+RpwhfwRk3ZTbV8
f9Q/NnN63pTICGxY7X5jidQhJFclQKVv75dGIPhamw2NPFkV0nn1W/VfvP+LXSvKBWce0OOkoZIi
KXsWOsbCjSXaOQfKGLH2KYWgyTfXCBu6xzLtZrYkB0QAsKgQbIpS1NejgS1KnY7vdKRt9KMdRoXG
LeXCUhG8Af5Z6imMXgYZU8P9RLx/TEG1raG/uDkcEG8beoR/pn53JQ6ZRu31XkMKR6UbaubuhYWO
0LapsHEpTAa9YCoIzvDcDrezVjM471AjzEPNY2P/Oo+fHE3Sl/CYiHxmw+19hVGwONA2i0LXPWDQ
hL0YMAeO2neW4SiUV4GVCVlOSo4eB5xqTF/3hzrdR0Ho5ffpN1zvZEmPNZ66Iyhca5U1FB1nBQFp
YgeZtzcEd9T3QPADKKMrJyGJwDATybgB8TRLm5qLtuglygMLmKvfB+cvboOO/lSY9ZfJ/gn/objU
56cTY/irHhgDDW10JM0e7uyDXw4HemoYO54l8KIoU+WJ3v7u6NUg7XMHaZhXny7N3Fo16bSSNq/U
w1NyZpRnP4ZmMGm0AzIo1d8jQ4hb5X9j0bYDHTuqe+0CWsW6K13RAQAfJ6Yxh+sudjq30f6CstW6
5rE7jxsZ4dDI2opunQC0UkfVBQ/9AQcLeUMW8ZNe0WGc7wExI+Qq0soMexZp7cGEoighzTwP0cuu
LWF8RLMyH66QDzkO2RAlv+TJLChUYNOUJN5+8rU/fL3ULePqi+vM4tWshW1k85WK8yajCQlWkcis
tHdlMKzPjfSNcWyDA4+UeFMc9YspY0uMqES+G2EsagPc/W5NyMpxWEEwvjEVsXAoVKocP+PMft2A
QjV93nsyA7HNmoVRc6Fu/H1NEPnrRRFUvmEL84jcw9YXz2tVjQ/QcKjanwjHDtPNkS8C8SdI/dC9
eyY8mODvYHiYtvO1FsspgwKvel+RUFgg0Tna00jZnWKXXnUiHFYuBME/J3itQSDkopuufIiBdhjc
B4kIxK51tfb3n1Wjg7jyF1FcVzmLymDJg1CJCuToNXBIKaKbA9eLYR6UijRIFcazlx2n6Svdvyrp
A8hZZQ8GhArVfMWB23AbZ/BNxD0NmbEmJDODWJHD3G3c35D2+sVOJmkyIkSJHq3oTrahdA9Y2ps7
YxLyNdx8TPm4t79j+ipdMtrK5PuIQqY64hxrnj7bGygXIZQ0Fy34/Qd04uoAiK04NpsboA68Gb56
n5dtYXqWGtCG7ABi5+MeWwsCc4zM7unoizgYSk+nWopx5CxviSSPeF07+4pkvDYwFj4s7JxBq+ur
iMrtEKVUZtj2Xur8UgbpJ5HP109UD8GZ5xij5wqnvrduDpVYoVXen+XHgso470v+XAX0infHJNqN
NWoTrKd1Qz8B1jLuaJ2fXj+MoDL8nuB8LLP3Nvjfk7vjkcTqlukxirfbki/4ovIF+UGKjfMHfZSn
IiC2IhK0VGVhYWEUPEp4qoPI85y9DjYUu2E0F7Lojp0x1d2I6J9UQ4DY2qMa+76VWnWukea0KlSr
mdF/lTklJvj9ZSzhFLeuWIX9EWqyLMxkVwWzoGkT1jqzBT7AM5H5GcIveBtNqVVqbZ0NGHsFSIIs
c1cPjgkyXSuI3OysmNP3yB1hi87EEOgA/eluqddpVW+sjoU1O7v/5uizavNF9xJpZ8SUFaY8H00k
iUGe+33Rmqb9A4L4Cio+yi5Cbqej5/7N32XZkULNwkjVVexbSwoPDhVTkZkPSY8t9KI5YC5T4RpG
8npVgETs7Z3wUYmU9M4SFzoesBs/R4Oh2faYN1n9basPzt10UNAdMH3l6b8pfA6ty9Iji5vKBlbK
G0YoY5/lFwu34Q+yj1epVLJ4h9+jpagFYUckEJIvbZk2R0fJnJZGzU4+0svOAMWhk/5WelgqNSox
DidV6Js2NhC6x8WwigYb8qmS3TQIRXmub5V4d0xDASwhbbqe47zcvUPMM/vdHwNciuIlAQ6qcV/a
hz8ck6TVgOxyL2vFdcgre0kVV4c2QnwH7WZ+AY2U+5fLVfAfSdPvgW/tzX8IFB0te8rFXdlIZ1n7
A/chvbPkpWdgUWAzEVkLj2+ADFots9aZs14nR6lNcHhA24Yuo0ILcNXfK4yQy3IAvVuy8pv8eQHW
e/uP5WYUFs9MWqaACjQjU24Y13IU8ShXHfpS7htmIr54AjoX4h7uPe6uTp/AOF4FoqPGFB5kh5e7
m1U3PFGTaFzdD2dHZnwJARoJ9e4NIRboeevfSSSkjLujRZH0ODTvGxLZWjPF5yY9rw9M67fPPgvf
TUjBTbclqfhddb/1JLsJ6bg5kd09YbTumgnVCVksMfFe8XqYHhQFsATYY4uLVqpuWDph50uOavqU
/hUNPnIirtcBPtzM9auXlaJi1ekFCwS22UMExOUnulYuNtxVJ6hu4OCYIQVlH2ewnGjfyB8m9flg
vkJdwPXHR3DXvK9dJcQK984vWCZrWZ/Opawy1kTf2nGcsrXCr9OjDsKaQKbKDNczdcJFCzu+JIah
daBqlag/dbVrRxeojdxWvRHe8FzV2gtK9/3s2nRKq+/8AL+k3csTnKKkrt952sQRCnvlfl9t1Hye
g6ljM++VJmqSjpeKdQtiELrOtgCT0q0nN7IrYIHFv1XaScZjGeNPhWTFTvq83sRexpPUPS2umYk4
VYBjtGKYO0whm9oEMDo5n5deOCwl23RlA9ITZ5BksE8uoV2/fV9Gij2W8OvU9a/iEt4un7olRodQ
9phFjGU/Lmk/qu5lGeR1PuHIbu9zDeM8moZxTfRc72H2WRvZSsDxGrlmEdwO0SA547WgMjp/YsdZ
Ispx9pM8viisfJWbAFvbf2G18wvwjAA3KbxN0a0r+QMx7gWkJvSHrro7zyVYCyPMzQupOlNzdMyO
5FJqm6voXDPd0Dyd+53bxwjT5h5jGBEXCJ2qdLeiniccQUQIqqarb7STpl6oipWA0Gaamxyn0QqR
r+mm/fVXAZtOg9vRQuhmDKyF3NsbPpIEKZtt/v0c5xfSfFj/r0ZAHFOHAouRtxboMaSr2JLU0Wx4
ZGd+rR6C6GL4Sowt/DXO8g2XPHT52kdCozTBE29vVyyYycUCQpjHfnabkeRgQa2Bec1igJAOHuxM
Fr8PRpO0eU8xJk6tXRUoPnF0RWuhE/8y/hEALDf1Z0aVLfJOJENj3iX7ghFPECMo8Dg70jiqXTsx
dvCQoNBnG22rUe8IfMsmgTnw5hsdeM2luhUtPeQpw9/xleKeipnrxAmG/CKWEmwHQ9wlc/V1jZi1
DRglplOICnNuEog36pFKJnMxiLt9qDEYHBzqjs1zPW6kR7XCrziWh1ZyzlnpZ+MODxpUwGSGzRmj
a4/JFXjkfy4lput2qHfQSBgywz21hEoIXRjF9dbp1OkD2yGRZbsAEr42jcxGdC/cucYedVk3GNM2
cTrA0danjwEhQIZ6uFwk4SFhHRrTw6vB7RpmI+kKNEvTWSL+4elno/E9sawR1ZLsx02rUCJR5l7B
XZya55MNFoKBV7SzSbArhMsx9UT9d8nvzkm++k/hAAL3KF5TId00bBw7QthTAZAz0aPu0l0WV7LN
3uCZQy86aZKsoxNHEtvniWMJ/YeEDa648fCf9mtM5jDcPxDURCMxVrJyFJ1R6kMmq8eFIHmjqJu/
1bumh1T8mD7jnmE7a+WRCrltjdz9xz7T1Ttx+CgE852KBGpqU9gVvh/Kk1oklpkhisTgKllGCAqL
A+j63Rf9q9HaghhgwYOFxby+Ei3KZn5uIDMDXSbTQqltAm3ruqQz7+h84ba6+wIskG0A/hKbion3
I/acFFELa1CfiMXlZ7Lj/Z64F2z0aiPyQ2IG+8uG2eTGQM8HEmbqShkQtcSjhPDllmHyjrAOcDyR
su8eSoCXL5rnN0qBdl2kwGqsuewlwcW9WeyRvH53l20zhgA8XM4M+rVVx+kgTC6KKbyS/KYup9jW
HTUUeiocEHClDe6DpOBEjrQKw6CyAR//Ay4NPXAZp4EIDhBVIEfWbvAki0QzlD6mYenY9kq+5oTy
wx//2Xm7EchScpCF62q/HbfJmFFf4AqnidLGhTsMveQfs3HNdZlNDCjc/5BlFx8oL4Wsy4jK1Ibz
2TKIFlNHW5+ZL3VOKKh7VVhLQnAN7w7YxUthQZHIhg3Rjh8QE35bXVnS3kNM9AsgVbwJGo1GSnyz
O/paaESm6MJ1/nLrWVwCcsnX9XJ38SWXJfMh37Jb4fVqRBawcXjbCs+zLqETmBM54gTrq/ogshfr
laV9d3YwhKvDfmPIUVqvz1quNt6ciB5QCKpHl8/lT9yHvrLWp7qdV7KYoz2Kst/nb9P/tywAWWht
u0ggc1t0tuX792mtdVKXNPT7Wa28hYT4MC1u/U9JspTys/wxqgNvJaYug6z6N0gI8ztxXYUCvDAd
cSvT8qodR0u6LZLAy97mHkWNwz+BftF8j0e4bj/Bd+BV/pgcxsgfLDTrdfXjpKpsWfmut79NSIHb
p4pWdkIA5x3C1GFlQNqba1o41dvxMhyljNIoOvsuI9Wokkb/4TnFZgsuPQPFjMaARd9nkKtJSRD/
eO3Gj0l4uPWLEm716rmGf6hiPtJ+lbBLYgHzyM2U6CCarvHCCmlM82Jb6J486TlT9s28chwqRgO5
9hbMPZe+GqSU4ny3mZIi7dUqpoqIGP+q5zJVaGposecFdRV2WSz43CTKNPSSvqNfIWcCFh5N2PwW
ECGDlNJf8yCy+Gc8cWu+wHK6JEtOXq5FU5/k3fy60SuSUm0424efdS0f9YQBBux9c8kuJH+7DjOh
BYmcBvvQPjJHmpne8Rbe4rCU7mNAg2cXPs7B9MC8aTjudqZ+vzllfGVKEUz8FZkKbI/5FYlgfLxK
bR0efRq451ck6CBM3gmUS6xU3PTODEeyyMS/G9a8kEubm8ikrzgZ2bf2yKZkGY74mkqHKtzVRe3q
Y8u7CmbiaZZETNX2zj2OvPeMh2beQwIzrJySAdR5BSlyBkoHjjJXVlVTEQyqek3BQtwt3HFeLNmE
JTXU175/JbMoPGFdXfsU3EiG3CTuMQaktmYUJPDjKPVA5PjexGcd6lJgBWZjAfcWDNpHGh4TibKL
8br/FCuRKlSkgHpmmFNNtHiwci4HYJ8gDkyYYqXrMIL13k+l5apx+bCm5y5H9iSx9AaFVawOidW/
69gi3aAx0JFSA6LYcBgpKQMRoiTvX3X2ph3O3qTtkqOdwh0nT2/ayucNPmccTHZB/wphnfHVqgjv
JpZM3tk5lgUpgoLA/v8uO5oaeeV2SySgDmDvhHMLP+vW0TMO6/GrTzU5bWX/FiT+Xe6rwxwaOgIL
qmDPg/uVy/JbQLD4nSNehdTTXYjASoQJF9/kYeDXFPxcDUksktZiQpndBt2WHNcW2fR8QuO0cjx1
x2ScjEogGKtnylIcCEM+k/MRzNwzTCGce+tajHSFgDaEgM1GvAHWP8i9KLjgkPSc4FMVQN9dyIQq
vmgUqNCqcc/tT+1umHOcOExT776t+XikjjmXXDVfZkRWSevzCqH2UKi84fwArjFkCsskCd1QZ3ny
qxqmVsBDyv+7BOwnavw6NzkPRsyU27HTDV5LYH02EpQax7udVvSTZnS0nI/JRtgd9GU9tliFCZ65
aHta+45SNJP84jZ0iC2/tH6LGOao+lXRC1mbbjaRvMlL0y+8Fm6nLzn0+4Mw2oUSOmLFphQgE3HF
Kbs/0m5g7rsUCsgSdCmhyeW39otbFxIdS5Nq3P4oNtdG/aj8xlNnsF/W7sqM38dtY5I0pNuisnca
HsgQn5iv96YZCch+vKPQD2yyrCG8/kn1zQV8eveVcH1+nGm0Cf+vVN9UITAltFtU+68pT20gHE7h
JZwTwIXmBo79XEovpYvmzckV/hNXzNTYCRrI6UDeWDjHKp6hUtRAzZt4vSs1O67kZz8QI12D6lAg
ZqP3qfQe/HV8FGFMrgP2dID6TA55LSM1whR0wJ/6+iXwzL6PZ8c9C7fgJ2WuoJUR4ecvnqM5DoRz
kcClE7DkCiN5Hel6UuTtySLljgazMzf7ZlcgdynvxUBJU++sQQKrRqxLhD0OWjWolxHFX8kKKs3E
V0diYMn6u3nRF4K/899B59rXsdAa4ldDL4TfWLC65GcUbBU+iZDHK394hSGQ1vz0pLdRFqEoN6p0
S7W2NOd991BZXCRIwSzoVbmXiCZDJVKXLqYGKQnCdpXupQmIA7irFaYx//a8ckK+z9cpnXA+R5/r
LV+ptHtpFXTDAqaro0ZufUhLZBTLJnYXlWkzN6KJctbAAdU3NT9dLn76wxfdkV+RW5ol4o2T1lgP
v9WE1A9pxUe9LrbF3dHQfhrzYv9cE7CesOnTMQ4MyUNgicnZ9kYxp0xfdr1Om+SrvVO90YquuKJN
S+kugT5+dhmjypZ+sAKVIup9MWB7lpiPO3ZY/9qShkS7mIZe68XZ+DEM/V2eL+MDcYAolKuWnT02
T/MoY0YkQiXBoojZXOZSXiv01UpHfe2hKnNcn9rYFqawSKYweHCfjl+MvghAmXDEE/eJhLOllqkk
Ej79pJTnZ/rQVYDTycYf/473yDk7LR1rGKDeS+aSnDKToIRWUoewsyGqgHrJfOTIhuFXLHMP4rHz
9tNmcbiNUWKPvhrF7GOlK9TwJSculpMjEKBKnGKdT72cMsm6NI6mFW9VudFocqXmarICDIYkDMDv
LyomP1sfGQ51gZ4dssjSOs4PP7N9R/+KwyO9/mLjSjorAfM9AdWstiE+nVcZjnb9ZH4RNSfKwi2t
yg/nAsp3fPw9RF5xHTRJEDlaK9Nc2Ti84aa8xbKKWXQPnfZbiO6eeDqW8+batrTUC5HN7kuoi3P4
+lBnrMUCn5ulMmYk/5N4fbhmsAp3q5geng45sr9AFNx6NlVHIRfnFv7fiWuWn+QJHlXv1lT6Wl4w
WY3aySlRR2Wseq5zniZklIXytEPgN64BkJHz4M5uR49BCgmhmXrxjnT/rdFm6dAKpdvuIlwlac7u
w+I78s5297Yg79GKgXZc66BMf7SltZL0rLBZooT7GMi4DZnzg/hyhcViOOi2cZXQFTdZJEyzHzyi
4c12BJqkHW/19SbE/x3G5IKFLwRzLoIq7qJJZBB4p/bAjVF+et2RAo2ZJz5o/4VtY1LF6zbX9a2J
/j7iX8m395fSC+4CgD9GvFe9lEuWub1D+gaU/7th8kauLyBauLea21Gnb3HUqeu7musVAdFIJMWJ
cbeNannR1E6Mps+IC+xCNSr2riYsafvAD9Kc7U42tzY6X8z0XSlJjdRB2Sxp0h+lV1uybJLzuA73
m8zFj5pdEFKL14Oyq4gNX9yDryYzORIqbl8mNe7KxRG89CszHZic7Qwh43bf+BJEcwlNz74F0kwc
rO0lzMzSsCq3rZy8XZSvI8TVmzyxO23PpU+MO+Op994QliFIcETLmtfKVwuREtMOJn00C7S00ny3
mulIN8DDd1mwMep2AqmIzKbXQ42gh79tn8e67rwidVVKsDTzMMkHOqg66VC4qle+8llWCFy8M+55
g95xJjHoiH294fDLFRGM4P2LEwVUPAWa1N9z+ZN8/QL/YDkK5sJJ0tjGQ4LsOrTgfDeyDqIuwewd
a+GM4oLN+uPrGMPMV+3QNQzDJxQxpLAxPMRPpDcpjcxzHIcFNiIK05UdNNBm/BBKw0X+0brwUIi0
tUUCGZUph1tMPREy6jGCdW3oIu09u0wPkGjoPpaIplYuOKq3R5KwX4o/GzcKKNhIuCOPq2ba11G4
TJa5eazr2QQ9up7hcU+0U+MfbG9Z3EdtHjLdje+qWu3YQeJBaoNjZQ3W/e1oGpuV07CIswKgvUOL
VFYkDrY8OoeQHOJ09FeQGpaDoW5v+GVmPoEXQwn7Mv/pRMhYJPAYPxe3Wmt01Z9EYFiBhw2L6W4e
8M6wYL/sTll8uv2tzrVF97Mc8Io06aQS33rkP/EjPmBHXqTIGGRKeS0t2zxgIu8WgouUCVgE15bw
KA4Aarw5vG/+rsiliShe+TYWpZvO6W7sc5Z8AdBWgOjNVupctG/QT7Qy2Lr/0ykbGQciLWf7jsiP
5zay3xzYastA+J29oP35IhGvDGJsS5OQcqKkAfLmY4pyHwHqwY/uatsaxDgfkV3WHreOI+DG1aNJ
hRruM1RsDlJQILDI2j5lFWm09ekOw8ZsRTF7th8VWE9AKfirRP0gkn4l5wl9nQy+qZ6vi1da2/+e
YnDoQQV1NzjFwXi0WW8fkcQM4n/n96hm29Vqm3cURctXUFv/UdtJKfOhbGAg6UGqfq+CJBFE9bJN
MV0A2rl+v7SF8zblZi9tHvFo5UNa5+Oz/2RBdn7KpQFBJ8ath1S479TD0cBBgnDd8eKewA5oKMPb
cYkFMLX+h39oLEl+BFfqtCFiTKv9DRxnGginrfADnaHteVxeOtrhu9Qw6oHgApgHI2T1wdO5/enK
ixPzNjTNYoR0Pacc6T8JFvB9/TWdd7ZehbRZocI6VWO+j7qL++NCV1ZayQIjqLA5U555p3p3M8Tn
aDfMuj1hVIROSX/pF/gjuVvVu0WBzOgyjuVWNRplzVy8MEG6vZX5VRXRJAGamIvdwQyf30Lx0tj5
+w+IOOHk9yeljASYxZ3CaJ/JusQNWj0i6q4bxR8UztpgDRQfnxgYInghO1JWxpyqSBOpb+USn35U
SQ793sjuvxO30NqJ42LLAQmauFSAWxbdwGsW0/tM6mo1S5Q8M/o4+hpsP68qj8rA/wy+gSuogjFU
w4aMk2VeQ64DbVyRJ6aaGCplx2rPlQnwoyWhbei6z77J8I8bGZv1Puccnp+//WeTlBY/Gj2ml9ht
x6y0RY4y+n/nOXLBitMuWqsYvL+7iyGxNOItPCbQvcMt6kKRF9scvGPRvJ17EdDSaaohSXlmum4U
pO4kCKyWr7KFsJga+q4YKBS206SL3cVSxffHrfU9nPD50Tr92rIPzRj7zNfDlp1MruXlepcd50fc
dWD2m6IJfKAc+abNu/hxWJbnb+h5v7RMxsjecpWkeYW1G/uuHUYOGvYOxP3/UyXznukzGo+QS8b9
0HI3wTkpD9OmwgN7EWq1dLCToNqkSiLz7NFH6z/sHitof6gu350BHGuyGAIXRxSprADZoH7lvt6d
YsDGDdPgawa/+EERk7TZzfFPD9gt5tW1UGkiKnVhkma5Y547BRigCsK8rrMlLNVg6+BSA3oscRvG
Z7YbmEvU2zBJY+JKvPN1bT7CVlL+SoSKB8P365EXbn8Fp5jWmBJIYWLgX0K/cAYkkeORvw/LNgia
lBG9Q16KNrC+sp9vuRrwg83n7uAgcp6NNBTcL3m5jIdaJNG2nFOXTxh4f96qu0o87b0Bg7amvqn3
vhf8EBXfpAieY3+sHKP5jubiaCddzD86nR1DBlzGbJvW9Vr0t8u+m9atjDDkqfku+G7q5Q5QH6un
BMmEfjl/IWQtWRvuqOtKGeThmunJIBcM2k+4tsWFsAC1K6YpQ6EiAWHLFQvtuhiT6ExdmNMD1C/s
WAyJ8czWMZtais1ePT7yJ/HrTMWbBluhcSvltnc09SVoGIEV3vqWNTS0aAa+/arFVZrSWM6Jj6Nb
M6GFjQmQhlQOys2zoBqVqT8MLEeFgH+d4f0uND8Y8/tRpGC5AfF8IRLb9HUfaFCPRbWBWVRC72JB
2/Y2+tZGy1YIEREsU+wN1k+a0x/1RSrem1HXYZv7dvutF2yZ4Npm8shnTzvyFxOzo03hKSUim8dM
0jJSa6RbIr/EvUwt7lPPvTj9uV9iokSmbpfRBmoZdqO0u7WNmEOVqK2CUDSbHlqn5E5pIIHCfDWq
PAZ+OG0EYB3UNgHIh0J06dGpFkStIS20vnYK1/hSptozQ3KWiUXMZ8Hc7pq6/gtMnc48hn9+1QHr
mPlR6VLwi4gc/O3LxblgUgbKjlD6079ueXeMVNPbP9Ii3UmGsUaK5oJqlStvfMiheAU0CgHXGWKU
s6YZCw5ni0PYdryKtsWmo5RF/hW8NWYVTeD4sokpAjrm6NmBfOL8pj6VXaA/iGEpdE/gVqgP0n1B
wPlf3cJodPIeaFZpVIRGEaIrzNdW4VHiM0EE9rSZq20n/v5utWkACDjunsS21o6dXDEWGLhUzgSv
S1Lx3tOmQ3NKhCo5nEEkb1RNAipWPjoH/OM4Re6kxqanexIcE43V06HslOMHHmuj9FKM8bLvGoxb
fxqZaw90GjHlt/4fd20eg7m99HhZh1RrPg9545k+GN9RlOjIugWuVVG/qXXeJ8QQv3McnJUWmFuD
B7m5JQ3c2lJ8Z1k4z/vvQ5z7I34lSNqCOWmPBo6YQQ+i/FNO1FtnOHhJr7/gjBmmiR+DRrVpT+EE
XSgXmjkiedp5iGkX8kBlIwRzExOCK0e/jpHU2FG9PFFPbs4myUpAh+YnX7tA5AKl6iqoASuZXx6D
YcYNN9dR9i+0VFxF+5D8ibQxhK6ezpsJBZBDY+xASGTWMqskvKSr8TVrmE6St4b6xj0QdeiuHH/9
OeUlJWOky8yYbfIc+wEKlpGpKpJAYpsUIeKqYgbE+0rCKj0PYkDkxYw2bXHngO16rlvFNrOTyu6X
crIUJYE5cwWmWqT8KtQMVFDMcjQ38U7W3I1wGXlsowjVW/DN7KTcjDDn+izeAEMvXNXmE4YXXf9F
E9ZPWw4S/VVKtO3xFdFlfMeGyZ7lYw78XSgT5Gn1Y0v+DLHUguAgMhhDtd7rDYdDPnj0Teraj8zU
R85nIyjaOVvd/keJpfDLhBA9B++U3B9aNVYWENnee90+iI54WfGBuLQUOnOyUQGzwj+1+2XLaeH8
O9AD/zxNfrsjn+lJZwa8NgPVVRSxDJ4TQAWW8nhwXjUloT/bbwsvrK7R0dnpg8Xpq/pNIbXJq1nh
3IUrhcCRvKygGiMVWTD1mOuNvPxwqBEu28BPQiYmcj9nadPYzuuI+TCoTN5thjCGq7eNWY/EqFmL
VKKKpoXatJ5Zn7CA/RxCQKJXjasixm9ri5qinxgBwALfs3EjpFQ3f3gXKTcadXvd03moRPzbM100
IHsqTa+kRw9e8UiqKFIU3y1QA0aFhaxgt8NmPB5DXlIPh4qTFxH7ouy90CiLL7dITCHjjavrd59g
/8uf9TUlwdstnauWrM17RUtQyBiAgCwRi81k3Vqftl80x7cOsTM0YDAQE+uP3k3DANHqsuwkbeaj
GjZ2VgY3jpCVLFvBTmPwjZ328XXxwk8E9aiDHaIAe4A5pZ2ddUuUrR8ZCjtPrbGDb6CzwYpAyYUp
xz852wTZ5/sWWqsDhL6dQwNkFp8e0k3bfIN61/Zsttk6k9U8/1BDg4lmq1QIbmy4Yqvm90yyKgRD
ti+c4CB1KkKJUKqmu2QmZf1Dr0TeusbdR3Eg3f8Od3sM7jVmdW6ICVQVMSIpuAd3GeRt0c3MBqHf
yXc0mwdpWS/62L9EsI7pxZf/R9NQ4MZJtXokyAyeQ99PYqxP12TqMqPX6/vUmMaTejS+1cgD2t4R
HIbIgmKb7CBh2QNlcPR1eJJwxWtL3E8f2rmyReXoLYrLAWZX2gddJPs+I7369wC7z4ZjipKo0feM
hhnQhcXVEw7hNO076Zmmp+S5y9/VaMDO1iIH/ekmpKP/Q2SofOUVYODiDZBETsV2NsMUEPA6PD9s
/eceQnJQnL4c2kUhMtKYT/hZo/gWw6krk58sdTsUgDjYVUOx7yeDc21YWyY2SfanFOVQmDKARbZO
YCmjTmN6d4Cyu1i/boTTZeMmbyJkEFNg1/hKZGg3Q8pNMA9CUPJew2KZJyNWjLI4hjEDO7LqAsLq
ttFDRmlP3elETJNHAhslB9ttnI8tKhMFJvgg+BDrIXNvtxnaa14gLNy1UbeucZHDjoJ6HZWKrGS4
aLZ/eGzJkhiWSkYBVrEferXccSe9QaaCsWn88mLHSB/mHDsQVStw8EUUKZgaujTxJK8400c1dv7t
kuSdctd+ir2VyYq6IlStsV3le1unsZUY1kucoQzy7uT4EG+v6DDotwG9lXHe5C5FpuytBFS4oz4h
DWeazNI8kKUmA6dZfhiSf0vqFl1TjDNnUqkH4mguF+2Xbh7Df92nlfe48rnJ/T5ZrQuZNyWMIjwv
tSOedLZvJrMOs0N2MajWPJzwR/NodYsnU1sypXuQaNy81inrksNUi6HalMsjBVDKlZRXrupNPLrA
ipTbWInNaYJ/1T4xq8AFTijVWhxk9k8mbtblUPCZRknPixd8ECoWL/WqYyTnPA9FnVFl+o/oQ8FL
SWYEJAwNeokRgWfRpsrJECsVd3RT9clC1sj/IFZyELrOV0NsxZ5p4ExHLA5T2I0Y7PyeQz3BTx6V
uaoPyB0ZeZybQHQJp/Plf0NcWvl0EltL5gXzsuLr6cZzJ6tZaJVIMWQ+7GKZSe/6daMsc7saC5RT
kM7SHfpgOqZj0ZVTz7KHdW7wchZQaZqerDOO8C2fgHim89OjV5ldPmwQSCrp1HAZrySQlPddhqaD
53vnEJRu5YsLD6eUI1POV+8Pq3E9kmR1VKzLRPz7tbK6cnZLXFwyB2AnWOBv6QGUcMQijJwogkaq
vb5kbv2sMFtUqHuc3OQ936CzaiSS1AkPQsQSR1MbWqRRk+3Wid5z9oHt8Qen7w88UkxLzHmXrgYU
W07hPnNpG0ZjZ8F6zvwZz41Qk+aV7hAMLyjDpHZZer9KoS3sLEFt+RcCvtJD0BpT87rL5X95GmnC
LNKO88YkcyqE39pwuaW+5+yT+IYaEEMZYQY1YZ2nUJ1XAxYLVvD0BfGMte6EfuiCL9f6MN7lJw2N
qcRkwdJY0efttpS9uPxBG/NGm16gIkE5I0tIrPFUmdadDf6DtRHUS8WyPVK/jZs5nQxKBSQHrFiw
u2zvtDFPKmeFAaAtfvs2m0Lcd0C+mQSOXgTNfnURWuMfB3SkWyNwQsSAGZbPjlt4/qTbFrCnbLBQ
zOrgoVBBKwH7A1RVOYd8pX3qLkYxkfYtRZdq+tw7ondin2QK/VLTz3nLC4a1eul3AHUWjMaqIuFw
5kKEYRTcB5K+dGAZ4iGRe6EuezV2KKErdR0mVG1kzd0FJXqsrKTe81eci9UvjcadiYcTKtF/PcJ1
oob5H8N5rXJ+JVOFMsKU+feqLUAcDMzdJdjHEm9HBft/aOri/RTQ/xziSIQgpTCm9jB4euJEYRuC
/NuredmpGyUQjBinINrNwWklVpn0QLAPFyDReiiMeIWlgzYjVqT2T3gNI9Qb96amvrhufOklzIL0
42m3HOMudIxUJ7ZrQjAhpOjA7N8Kjzy94vh3qRSqdSsoTMFQ9XezMCF9DmSb4hCPk+EsWOHDS2ru
rdWBEe20aqwrzRVnVyiFrbQCmAioS1GyiEoHbZHCRGGTQeCVwfpL7HyxZAFBYkLTKTAuPV1L4nKP
4eIQ60eYra50jsRIT/dWoECI4vHY1iCWi8irDyz/eqI+ZMMOgeWWh2ER+ho5FA0u6j96+iYeqLXo
osUd3ZGm+RbmWxkfLDTHiAwJ2/HuX20cYG2gfnhgY1Vu2ww+1BYhq1yzVvUNuli994XfyquD8brV
cL4EfrDtPGBxzusF/QasNOVlrFvUSRQhgqr2SZ1TRGN/lMzjZevpBGsvp4wbwe10DVT37/MbxGRN
4catIguuK/K6iXNfgWJmp6yyxTstd7USoLsIMsNWYZVTBHIBy+R5te6YHrmZuJxg1/7h7/wZIjxT
Xc3L6T6mzD0RA5x4L7JjivQ6wWHDBY0owD+LXHhD4KA+izp+buBpt6vQwJoK5ZVECxACckAp+cpD
iFPJymq7IXZoAh7WeektiEIIe/3myc7aXmvu8QPuyBWq9r9OycmZOnNJIZ8iI81wQ92THBKY3rFS
2YXgW2ywtAVZZYkttTB5U/ZAI9J7wvFCOH+1ZFLCw8d93hlBzeg8G/izE2+39w5oJwi3qOiWQg39
zlNAWR+lf/eN1C4GdqEGzvZPgvMcIk5DjNwnptq3utyFCpwztx3M8qePNirMNVfO9UV0oLZ4n9TX
mQ5RjUQJod+oGw9eEVXnss+WrCuxGNi/y2V0BsYwwsOzenqkTGybp3QaHkdGK/A5X069jsNRWB6F
FCdIuhPK5gspCQ6B0JQyibm4T3mv1B6BxO67HCBfX7PsR0+YuEljEtnHflpcc1Y5A+k3mup/iq1u
+M2Xd6k0vKYI0fGNQPq4txh8oPDEUoIkPnwp3/VX8p1QsO8Wh1Bt6iykG6tssXlLxWH4HF2MBCWe
YSEOpSD42bg6KBDliW6fD35FtIVW2yhqAwQ2ADEWyZJZ4NbFkiBDRGWD6oua5igVYIoBo7leMuHU
4wfVsmv66tl/R0yLPechveVzbqhQVlbmYl5YjqOFeS5n6XfSOj9kaTF6PUHJifLdHKFBJGJkL9+9
B3ZmBn3uk2xwKc+fgmm6pSdRBj6fPaIAr7aSl+C9lQYuO4Bci7xEgU33eERKTeLSPWI+zmCSMdBp
TIgGBHWQrJkQ5gFx55tTvS9Uf2nOOkTqJmCc1wa+4Tx8uFXmvn8SH6JaMfr75LFC9XW0FV1LQOPo
Mi4ggsamhySBv04R2F2N7Gazemudqi/qk5YZqk3i+NDrNirDJErQYIhGHwsArZ3MDC1oLE5j7m8J
EQgKilo2uGg27+nA2UAHlw7lbsbGsctrTHszfGHnT+vCJ3cx6K8k6s3HXTtsVVhvgfXqyqQ1zb0E
EHt6VV51psVTiyUHnV8am4yENHa09xgy+FqmW9A6F1qsWGi61RCvEHl3uyF2daJxBPXGQLdUWVSE
wbGHPL2OzS5zszZyYjfJTxeTDi9ZFqBaLGTnEGVwrI7XKL5pxsgBv2NHnWQkXnAYH71oTYHZZWxy
U6yZOmc7XTnD+CDBnsszGtEc++FTfuyYxHtGJZKuul2aKmj1CzeO1/frc/O0XGgOysg8vVNoB33R
YoxvIuCwT97XOPY1/1M4ZnriWG/a1+m5v9EaIFbmoWgDF9j+3yqxgk8mjUosHS8uR++6mhSejv7P
uDS8d3Ev+Dzwze6hArumQHekBkMZhXq9VPaanvS1lqGbJmFSiNcavGWurbMZtDrgKTdzOYSdc50g
nclU/4JP4q/GFYo+sy8EcXC8p12ixcgYOTnmT6GmKTTXdpZc5InmLDrOsRKcnZQT1uQsLGgX1+g+
2/l6YkJfIVznzTD+t/D1pi8iPgEmYmJRG1NgMRrqhkS4XV51Jryh/kDw8WZfB7kJr5IerQmcJNyp
nXn+xtp6U0falXbEoCZKB9pnSKb1vMjjf82PaCbIS+u8+Ao8jlM8WJjzJxkFiyRVFVFOV0yvIyJL
YYGRu5UMx3VJCovQvbkd5nNHlQNpv7y7Sws5viKfWIEnqcKd0Z0dsoCVDpk5y7jaG1hc7GEW+fjr
l1kiYnJi1Y+3jBnSSM2OvIPmFbAMsDtsG0kPVIw5VW10mZ78KqPg7WKf4lFN9vrtzT7mtRQ4GrWC
vssWzTVPV1NbLNh054Qi3PztPl3nLlf+rdVyQo08XPECDY3zIjokJDyv45vaRYpdJYjWA+r56Bd0
rWTXxmLspqHtfcafgvaAejXUTBk+eEnK+ZNwfSpPSYlpQcMXr9nzUZpEetvC8fwn/GoZvTxa+PLG
A0RvX114dALvsy9HwS0fVM9szn/SKNtskn5dPWyun5MoEcPxXmW6VtaYsV4YVM4mWqKClQliicKN
xdTGhvtoBOhamzDOGBFu9uklIiXqmA+wed5rvuhifQ8eNReedH3dfvAcY9Q4u9IbOKjxQsu/0mKq
S03kDdoS8d4V5y8iQ52RJ8CdxLmp30ErDa+EdQp6FzPDQfpqd1GZTM3dwIJ2ou60oZ4lBmpRJrDn
bcXKT6mOv+RJ7gc4cGwCq+RdAI1YkgXCAapNNlxF52FIRcWJKK4Ho2JPUBEmPz08yCB8OsscFnij
Nd6Eq7Qb/WMpy8vGvG69mXVEP72dWsRzX/fyM9tHyLqcWiZfF+n2fnzB66YQsO40iOnvaq+r9NgE
34XR5wqNC6uglHw1EUIHR+oXn+9WA+NUPX7c8mGw2EQHao0QUo6fCQY4MQ5381Srwx3jkNKqvVu/
I1UmH5PmwGOo65+ShtjGY1N1pWOj/AsavRV9lb5mk1JWe9kMLQnD4XKsxGPdWsX6SOuuvd41fcoF
4vSbJCGULYFGaj8nIVIS/ygXFhmzX8E+7pGIiODpOaLePcGQgRY4Zd2PQPaqloyV8HTEVzHNucDJ
fY3Jum8kRnD4mRaK85zwjRVYGbvjwx7v4dbRlA2n7Xvfr1CXO9Sj1DbjQHkBQjzQcm0/skhOZs4m
mhgVoOmrfU6pGlW6gWbtuAFKqkYlj9TjakCsYdSipTmaqVE2/zOuZvQsXxs/b61awSHoir/6J55V
lZ6wEseESPh0KYl4hvbCDjGUtYnx+MBK8ClszxlJLj5UWmYd49/7lxjz99m1o9uJFXc7NHXBAqUw
prbBmrvqV/fDjikeD7rc+6GUi4vzbINgaSEK4duAGwT16AsvaZKEwbBsBOfZYOqrFHcpz1S2+Ms0
jJdTi+VmsR7Fb7H4TPM7FCUs0xIqVvPBDAnyv7ybegrS+VITPl/0nChOK3Ad5WKH90deRmWzWICL
tprwSygxSHqdfxkjw3u2Org7JS2XwKhqQB1XrqWtBs+8m8IS2sgHclMg9U68PAfeGeNryA7/O7bz
C6jsVrtr+qeH1Y4SnCoV6YqOIz2x9GdnvTcCX2JViA6931c//R7sAmgVd9RohMYghC8V6OF1wWK8
44vNM/r1uhBKIVJSYKkAK1Erd5WDOb1c2HUA4TxsgJvAMtVhAt69EhFEYe1IgI6JjYIgCoQ7aYff
FntzCpN8YYLs1KlXRMrWuqohdIuZ8BMOBCrMt/JWSkHtdDq7C+Yeltrv/uTYTP8hEHcS5uyjmYgI
sKqx6jhwjz08VaKNNQfVptPA8TLBQcGVnu+aYrAF9A6lx2zumwx/QopfSSjFepCdnuj1+DYzJEZD
7fwmH42IejjpLSETteX7J7GO9rxWCKVUREMOKrGgwfI1tIPbyWKMosJFjkCNBlzu2clCoRlresRX
1lDlM0BWbtv+oFc7XsYNgvqfG/y3FmONg1NbYWAYScfLH1OrN11Pr3e/1p6bVA1ONdDf0MugYeii
vSnOve4XWV9Wsfez2U92qFIrij24Wi3+kz7A+Z/mUmc5hO8JHPYocbk1dp6gzb+u6BOZEI1XkUiS
GRNe2Vaqlu2m7gAtVqqLcTTgPoCn0M/g9+jcoVyVZvr7pJeXeEprfanXfgzrt8NcKyUZgaRBH8H/
VM3CuK0gkVoWwP5nYS83IZkZniBQl6xzyTbD4MxCfChWrNmFokg0GM0ZqR6HmCYSsX5wzM7Fr4vq
MgFHaVY8Z6QilDiEW6QU5yYZ2PtAOa5kGb5r3ldIvNbXyPJmayAw4jA8REQcUk+m7mkDZzZ5rwDG
RIuKpIuP5ObPu/+dkWjdMAmIwPA0WlQXzw+RFekwmVioQZUd/HdN/kA/DnUJhwRNTPgWLMuIjdAi
VrIn8wfPQWBzUXIB1U24gXMvWdLqFcgCG/xhw12apaxAMSnBfyw7hgc3YGs8KWH518HvYdtWw3xT
tpafqGjyS+y3i8v2vFLHSr81IbwFWzEP13g6ecDhWn9REI/y0KQb/eMqrITj2I4YZt7XpvT9UjKh
XcVQsW+yfG3CzRLuLjE1rO2Ip4EqNknNq8/3Q6jOANWSXUTl8HD9EX09fJkUYz46SlePktFBDcX+
d8fh1ZyFJ55X5p21f+0YcPprTwo8zeKDGqQ2k20kEyEQ89MyXW/yYlFJsQ6wXtEn2VES/2zajQPE
MW49pP99GHq3mD2mMSKBXPBueCvhoYL17CwyxTFpzNVMyI0fik993nl3fZ9fUGucZkQ+EjI6hblo
TF1cmmLoyl3ehpxus2CpAuhIjOn7wZqNTUAD+5pW8bDNktObuokDK3DdabQpQpjwWRWo5f8NranP
Omgbou6OFj5r23pHg730HOE3W8dJZCUKdyW252PV+fQ3jKi5tuBAiV1TQBg/vV+UCAW7W+GteXnu
OraSdbDke54l2WqqUqwP2Achp93An6BXLnfrH2ku4oKRu9cgmqLkPXiVs4F0ZMvYXYHSecQGgw83
lX1abX5t0ZRz5navmGvWAXLdOgbUxSUCkdDNazc4LZYkqsTUKCpCkU7gJYdmN+wq8W4s0ZxsV/tE
1k1bZLRb1ObMzSEXYjRKYH56Hnai9zYTmyUKlPmhxe8+wda5pcBnMjbfSvACD8iI6BrzkhpXCGt8
ePejD9aqZHbQxF5yGXUpOP6+TGLx+NTjQBYBJCitttnaB2/hHWfNo0SkCqZzUCdsATrzJfVEQD0s
HoYRyqsBAv40D3/53kQ38FFt08xbw0tSlH87lvZVymTdrQOwIeVYmO3kugCVECVIuk9Ly4pNtuJL
I99nroQAC6H8Fmf1N4d1K7bVNVsE7OXHvr6yU1BC2t2wgOvGcfBhTCPPTrGa2uygJScW45SeKDWs
GA1M0b6lXvLEGNb0LaL4guU3AM+dNv1pHW+rCOQjGpCqWfuHlc3/sxLgQt29hJMZ9r6Ka6PNDS9M
KvjzC24/paNymOKResS4p/ge20QIpd77jdtQci8KgmmxPlQ0zT15GaUbO59Tor5E3GUIZcB8c/wA
NFEYYWyiL1QHaF4mt78tImgNWs7X37wP2TOKCptFMP2N7ft/RXl7TNhRkzejt5VJqNFJqVGXXll5
w6u6/L+cbNds5P2PPIgF3eRDn2mJ49CoJiAF+jrhoHtOo2yR08khVhtXkOndR/UcwmsNVRnrmqZG
PfDR4PDA7EYv1Ne79Mcj4c9H4C+KR9UZoGL/3RgpF2XkhIiJBXSh4dFeLfp6eLTZM9VbXscA2ap+
GyILolV/urqqDgk2/7tEsIRhRcqSavA4skOhGBsOV307lREkgLOMTcO8WIFdfcFeu1aZG4DJ2mPS
O1jrQKIgquPGJz8LFKB4eM99DFfWQ0H7f4RupcTj4G0HdlwTSP4v/GZpqHdy6pCqgEtMrMKf8h8W
7FoyloeQh4T+/umd7pcIl8DXAjmkuKn843m2D5Uc7sbWsz9rRyBgIOKRD3uP0yiUQ25FbBX+C0AJ
LR1lXzmFLkE1ByVgpv583rr0v2ENVwyRhFj1MA8ivh+UnWr7b7YP8yKFY3VRmC17IRNrGMLOcr8z
AAzCOBqrXYJrNgUSETduU2FxHZZjuWZItUV7B4FVlhaFP8FaeLE6bAcdPW+B15+6jK9MRHQ4Ayjy
PJVGr7MHxujC5p+RAosBrpo0JpTDFcqlb6k/oYUSA2ZtJIJP8Wh217Xzwd6sq6pFabmh49YYRw0r
1Tf4Ez7k1yugmUY/VBCtfJ5tshW1O2AIivp35ihEWJAylNcg9h5UcS+7hvrr6Sw1GMR3b4mm8+sh
k4UZinXkE4QL2x850oNyV2gl1K76SOs91Ra1n+CQu14hp5kylJB11qxgDmt9aGvW/48XMTf3KEAS
dJo/V/tz1DnWdpit74I4/Ld0c3U1U4VKT8Ug7SNcpVoDhVutfim4F37nmulfdrX86xUcuclZvO1N
p2Vucz0A1C/6POfrj5XXUUN6+4c49B1MWHakj23FyuNYN3tG+k3KDGC3I98dxejxONhojMPKdtcE
ExpnHFabNDkOm4+LbOsTbq/3dIIyfdplhtwBweK8ClxN5xqX7oMCZ4HxlVne6z5dWxOO/76AN/Kd
FkrmbSInj9gZs0Cc55IOAgWP1bEL8T7O58dtoM0o3Ti00I4TEpuZTbk6/1Onc6O5qkm7c6rNZj/B
3hyQkj7FmCqlR4FxBMI2edHaIJl0zyy8GXZQ00y3ngujnLz56wRg0c0mpZiVTz9/tQSbFe+u8G8f
9yKFQLTwRWCcmj/WchaZAHVmSkQwFw3u31f7InRgbtFbYdcnXnMwQJ7zBN72WCeW5f4fI9GImLH9
A3akbVo2W2CTWeZBr1yu77syiDPlhWD4VERV8g41ko5XYE3wMufChC8duwXoIAZv7l3tQRkyEAAW
4U3k2U/LD1PPY7YMZV4IRN4r4OCwB0vd1GkDdGcraxk0MToQNTNkZ/BehXxeJIKP43PGvJVBlzaX
RqByfyQbaaFEL8NphO+0Uf27a6h7lyG+AW/G64o84NiRTROng7qsBBqkxE07645AOSAaryWfjs9Z
ya1QO0u1uPsKC5olKKZM22cOYDBTWhEVj213n7lZx/YoBEoqRAOyqZkUur3/TjM5O4p97wRINtv8
JTDBR0xarPeDxT9jVXc0bbAWXU8ed9pJAP4FenXrRIxRann4f2f14aXfQM1xtXt5wTh32ZdvCuD/
yE33tPeYV+BFuLJ9BPFyYqRAGrD6rrdSQ/PCm4H4yDvPWsNEdfl3cff2OGqVQ+EOJpH7gBRMFSP/
70Sk38hndg0A3CfQuS2xxZipo8rwKT8fL2sX7kNJaIC2Oe7hXReSIyQiqQMA5xjJRk4RT6Aqe+Bz
s4w6WwOqjfzC+3v2Lg5N4u7ehGcWldXQBIPgCqSPAzB4MYNUz2Puuinb73G5m9z07mzwkTBJoQHo
9JwXn2vvTYmajes2GFZHxcL0qNWPtnId9iJ/EfX9s/nhAGyvXNWzRJJf9991ro0ca3lE7bpaki0f
anZ5e8g/Z8KwnFY7yzbC6GUHUqSWYCkFfs4kD0bWdmnVxcpKuo6jnKpdtvoMnMPO8qVnvSxA9pBV
uQH1OcOSlXUFVVntUJA65GiYxf+uizTLoUwqI9Ax4XDpeXrhbGxFey7G0QXVIZJfh81Obu6hQd2N
1JPpgFmUm/rsvyJlJdJQ1EfzcmwX5SIVMCOyFqPNaq7mTHtwbbmqq5gig3bPesRPsCvrI9XzNAkf
4S9OToJgP0kFGYroCD52lf/JtYeQXQ9IBIXYc0k2zF/eZAsBev8MEb3frJeDc8vcBLYXI2mTPaqz
iIh83AtbmspYA0wmu04zMT9HV0rJE5LYrLy26o0H6twlUgWXmeJXGo5LwSSw0gDfKBzPVc712CiT
Egl1cbFbpuxIFbPvovU3v56vnaaGXmWro8k+3gGobrpfP6FarkJalXUvUB0LOGErFjJx4rpOv+To
/dE4810AlRt9Gc7QZYx/WL3grA5JFq7DQgzNj6Ux6Q6WE102z1ewSQALzT01A+/8/ePcGp1EMhSV
Ch2E0ETThkMkNWQR+tJp6nWJPNUr1Vnsy0vV46gT+M2jIyNddFYoB8s9KOpmhK41a4gCVY076v4P
trPfGgV8k1rq+1ipSaiv7HyZHGvMWRwhqKavCviS1an19WKWz9FSZaW+Kwv+d/zuGKh1IQkWQdyV
Nd+E0MiJisrhVd+P1vtZcPRu05rp8fXRVD9wESQ8en+RQNYz/IimqoFmEQ5g468Z0C1DMggoTXh/
y4trfId5XfIPf6HkFJFXfN6C2OMC6ypeQcpK25+4kUvGpidercDivEVe9pikZKqbLyC17kTjwYz+
FLHGv3b6a/CzyapmHgqz857SkxcrFQoKtBXpUzi2MfpauJma/vyNzTw4I0AzUgAvM2J8yQ2uWHTC
2VLzwTzfO075R838L75It2v6/ecqC8YCOYNy8KH160bSpOC0sZaOh0KqBCk78nXE7T8tyYRflrbN
elVVBhAr7YLbW0HxPbm2JgorZmmG1QvE0+dVqN7plud9aMLaBCjxKl9K8vKo9sPswnuCq7W5s/HS
v3v5TVVgYXu5a1g8p0+VPlghQvuzN3ujjmT8sDxtyFDaK/CSxxqISGGwA6iadDzRyzNCmbCz9BrR
aaOUNMVBz82uhU3nL/rlMyx+Q1wgttUbYW/7kDASRj9+3Rfd5uNCkuu48FBzWQ+CjAJarKH33nup
ipgav5Mh8RKo3gF8B8VmhGVQimOKeqdCbYDTj08yERU8OUPtu5hIgHbm8lPQ+S3DraontvhF9ZS+
RKGB134i7+jfVDDeibNVoqPOGHkcLEeofNGzcrGijQHHzdFxScQC8VqR8gtAQgMaUHAkEtYtppNZ
L2COC6CJVRydZG4IjLYLHwoABDoO8FjcByizf3z2DzDZidoqq1i+LkaC7/3typozL0akCXc3lfp1
BW8C+jSPNhQ5YTkWCvlF0YXcJLUaIsqZzherTLykM9kC8+Xu2E7us7p502DZhgcEDoeacxbZ4b/A
F08lOLSQJMnViPKgxeus5gglRemwh3UXUqvv5g5vWGIyo7WrkEDo7aZ7tQ+xs7Dglxg+QtfeIwzJ
V1nQ/KURVyOwIWKkjlWCC6Yb3SY/CH7+a8b+g2S7eMUNWeTZfZzqCFrfFaP5lxfgU0bnb7AU5xZK
y86xpO5yn8ivfgFUQ5wT8QEHSUlEJnKqfxmoJGy4/R7Kiv7pA/6R3WiDjoL+vGAyqckpWthmrTo+
hE7SBoThwOnZrNCHDnYStwg3hx/Myq/fYSWVNDIhXb4xaduLeRdaNbJJHL4zpak8etaBqehQusuq
Cm65XIRA4G2m+XUR0BEPqvvjwkv9MRvvbCi++Kth2jNt3H3KE/s9Ix7F8gF55hR5ApmHmnlMW7bA
/Onp+6mSPMrBWI7xfgTft/bl9ryxLGRclQpqKaZm3PBnxc2BRMOFzmZZPKQusu3suVRqv9SavDpr
XLyaQSE6nbySdKP3evLkPJ9BeIjJXgQSejfzVs6bE5O0lbCbWK/jjRlb3fLG4l2ZGmMeZ9BqHbav
gZyq8MS59gV5cOf2RGYkvqFq2WdFMEZhD+HfbSi4gsqmgrQHVQLf/DsJCig60Vv+dd0637LhA3hq
Tv43lfOy7kZagf35t0435DRy/lh10uX7IzMCKPpPRzOherh97COu77kaYIdK6dc2qgbp7nJd3cEC
9CMLuC5XSKPPPH035unznCCAXJzgeXbpkr+mxel5CFT/94+jvvIWp0fUIauYC5w9H3N92wbi60BB
Bdvrh822B47RDeu+k4rboZk/4NOd+ra3Y30eYbpCvO4U1RzMKSoIVzafTdPy8Y+6q4+vE6JCDMaS
WvDntm49BYYhjBsmNzEDf6L9TM5vfvA1vqv1PmFH0YGP21Ut29EUrBPdBtV0lVDQgNXlL4RXPVIw
5D96VKKGE6FQZTb+Q9YlyT1bPS3XJwO+/JtbS7l1jF8DkIDUh3Plr9M+rRj1zQ31gpouAjSmO2wB
9YucMDyQxrFmoXG61Rs+vVgMGEvsWqKeEZ6khgtMpFsqgKfpTL0ozWn0mkh/ccEB1ddN4hSibra+
0zlVWwpsSeUpDSKTsw+MpQMKwl+1AZVbliTzNpzCRE5ixyQZUeh9rqPnt0M4aJsg4C4LbmNcneJQ
5AKNw0zlLeRmv5twSxv47Q+SMSBoI96KEBrUz63wW41xRc9x8laR5ve/i8xGfM16V6nTOkBq0Ty+
9z3IgtPRsfmu2CN1EalQKgX3KKcpFRzszsmf49mjJTKPdI2dveqb7/9BokZzTONY/QN/ErR8Aoh0
Da/zHDIHVyz34SylaZkubo57r7SkVI3LViO1+kEtbwvq1CHKxo8fH1b9MuSosb4Ma9SAjIOhEFPO
nyfwqFEIiO9DU9mfwAXJWCSmdQHKKQjMC41p+xXOzi54FfcXZG6S2gaK9/rG0ob6CHIcAt7Dtx3L
rfez/nNPnhqSH8DDf/wmzLAd/gBBxquJNB0WNShqNaUbKRqQafAFsVMHFjAAV/tFQp26vf7okwj3
IFyqJStZCmHafcPblRW8sO+vVPAOFl0zUqlytnEqViKxphaWU4E8mjJw22tli4cYSZqL2W6l2GYC
HfZevPd85rE3Ey0Ac2XJ8P0GbTW0hLLmhO/MWTEPMYP/zD5Glr5PQcjJiKJKla/xHHDEqnyGE2Oq
1fR/FYScPvJNoMlExwlUgm/l5JaDrJRaGVJMgflX+J4P7FnKewioHO52BEZxXekJ4w9Cf7ktdjiO
7D2W+NDRTUV2Fr8ilYHUjX4mHmA7RigmbBCb2j8Q/x+PzMQosZG9/h1LdHL6d2aDA1znG71ArmO1
DFXfRbOPVGtPx5dh94Rx18xe2hDD0VNScGSZKt57iORZ1F/WZhVLCtMYo8oG/UQIaTp3PgwOU6Sr
gkDV2eBFLCBMI1009+6jYt3wuBTLZJkMRENE/tY4lNqMrzsrCnppUuCpNb8+w2rjcui1LdhAynlw
QXdMCk17z2wZ8nsZu+MMFcgYCTvCPGgIlQXHOrdMBXOC2nP9sqJgDiomh+Cg+S8/WUX5sE3ZSOsm
0zsHerxVNGG5U9uH6HFuyBvk8NmIcaGXX/BKViwuFHLYhwHZwFXBkQdNN0kOsiazF8AkBT12i8B/
FNTHLRa1wX/J7JHp1NUePK6VhMC0iJIq13/dBkHGE/ptE9DlK/xbzW/RdmJFFi9APL/sTveWzqUB
ghxF8+RrY/i4j3F3Lk65cXQla5J5BH6Xk8PHq9X7Kxyoh2vxHSoD3qtqkRssqZO8asegi5AXmJdJ
tPoRJepIfSr9ISGGp/7tzCHFbtz5ZIVRZLexVj5b24le/qnK0uCSh37jx0yYtVGfokyciEuGGAK0
dcS32BFgHSQ52mJtZ4KqavBkgU3JTGghzi4Bfq3HzepA7jmjZwi1Vfkxziuo0jkevkW1ziXcUWHI
yuJlTSule5QP3Gkwdwb/H7ns79xxKXfwrEcSCLoihOCWL9qlZ5+kTXIBmdBRNoemmycgirI7loZv
ocm0XYjxT92xqbMvQl2vfbop0Tea/Chnm3hsKLBinbPr6k2c8Xw70seynMtG67eMSahf0N4Js/Cy
vXknpeMGYgv8rM3gZooMiStEBejjouVtXU6MEiFwndUtZUjMCrYpj8495zWYyrE0jSuQxxtFgTKk
PDlH8vQQrnrHKH3UsgEFdlRF8jRUR24i8ODEbXN79KdSGsL/V21q5SfDzPRGRwbtMSmarZ3f/eRu
auhdfJhWVmzbeGbTTA9SYXRJq9+mn+E6FCA706KNuELur26bIvYEXK4uTpg22a+OVY7qLpX6SMod
aJ+cqfr5W7IPs9bIDjsh/k5BAPsZV/tKBZvnuVfUzZYADuQbF1ae3hTetB+92R16VX/P/80UKMCg
CpxecOXjBQaGyFEQ+JkIa+hX/Gkzq604qoQYi24EJJRtZYlY/E4mBZ/wOrQyqc43TsSo5fmuaNd5
0oc0i3p1OZvfEilEhwjVGiUMjvCUIZSClxjgwrnQfybJLiOSWua++a2f3TaNYzhvkUfJbtHg5IDg
/LPuc4Qel93j0tRnxFTb9Keu0PdXQpBMwu1T1ljlyfbGnTv+G9noI81Yx/781T3ID80a3GJaSYjE
Hy1H7Axy1wxLe2P5ftXFf2wNisB51tHCEQtd5fjtfTrJZsnZzgyJxn0oopYTs13NMLTLs6mHB18C
OiUX62OEgTQGHQtNvirZ4zvcmtAE+XsNzukRfeSKdu3sIwfOiUsL3BRrM4lW8T+DF5QknQBDdJG7
lBe2isGoFNfa2DG/U0kpqXq6KDv0zgwZNS8EGFW1KS0rb3mdO56bzDRWLHwBCyCfkivi1pg0SVsM
BYRs2BI5N0p9mgcHfuNovwlfA91YnzopAGXszpwJogOmZECAhdDdFMdQooD+d3M7NcfnZM1z8sm7
SjS3yFWx8F63+GVoJSHCbxWCT0VrpTGyCpujIz6x9XVl/zFsllQ+n6M0o4hb/YOcNcRsG3yVmEHn
VdcwSe1zUlMEmzkocvwA0U0xssU8rq/K5CMQs2cBA1YBGNs27tSC862kQK0auz0rHiNApyl7a/5G
PjpB4Rta7rcxTKG48k+SoRQYRDXbjcYyeZC2CJ/psp9EZgWe9nHK6tSLHkOjHa1a6lSrrFCAuB+4
JcHDkG8QNmkAZXx22V7rc2FSYlrbAh21bCNOvdj66jCDudrUJXN2VMxK0oYEj5+UEakBCMvB1KDa
vWrE6uv6KIGHAuN7iynSDIpXZl72SoB/TdJa3MQKBMgGcTCap8n17+pQYxtKmP2DwiJlSRGPSekK
FVt0viJoO6hlLW/Yyf4IP6rvTa52UoD4dOlFgA7tdtdj5nhB2Cjq6jNPt+4JQLtW4gUSWTr0lO0E
l9/FIvxNKRm3vE6+fg+mVEr3Pb6NfQ9c++oJ1/eUgMhxzkAI8jeWpccUqKcm55RJ2w6/WdXme1FC
5yZAQy8++9S3+9VwBziwlmPeWOJB8KaM24LvKugLXFPUiJZwaHNsXPG/ynX+BtCUJoFkNAsRKa4u
8DfvnJPyZbP7yREa4BLW8gQ5kbUZNt7Ex8M4hYUoK8OdvD6yEcOEINvfFFNYE/lVvxyr/KVP6Ifa
b9zH2Bo0A1PUFBUMOXawSynboQDKGccJYPvJCT3eFlwS4lfuKQO9fVqBhCR4dyTHaWdwkKFSv6Db
pIymCZ7rZrsWec/I+/CLYYGvZbgZCRqcVPlE37iFRXOZQzU9GIxcWBoeSem81yaPLXK9vWcdUfI+
QAFg6q2+agaVtnmhQH1FuMH1kwOXzMRhn+tPBzqoMoAGDN71m+oM4h9+I6/Wf+NXs/+M0Y375leC
z9clNVdw4Oo9+g/oKJurzy8cEkRKTqoHX+vratg1rmub/teJuLifXB+dAvxONpreoQbKk7vOOYOq
UFBLj/kuc2zyf2UCt9QmjWkI5Ygg+TaTlv88wpWdzDTczQqSXCGFL5xm3c1gj4Az4J5IkTDef7lk
Xkkcw5NcoWHwhN8qZh5fpKI9XXHLxDWjjQYDPgl0Jp9ZvkWgY6joK7sHhUBf1OL6kuHSRL+jOJ2a
1MMl3cuR2oPgtmgEDUbe7HT0yZxwLHOXAKETeJkifGNt0i1Ctxl/9LhSoa4istisc+yWFahZ+Uvq
cAgVMk+vNLDYbAeepBRpq0Of6StRl2L/mGSKc6aBNjfYRQmqrsaI/8P3xZdEjptiU96UzndVKxWI
woA9hhkvbZG8RajJAZUZvNTTd0y49LJ4sP5kX1rppTDmAfbnhbX0ZNmMTY4MsU8eR0bSpQxladYp
sj+K8byu/wEeScnvs3tAyNvTJVBLkaeoUTriq1rFKvcSbvuO7k8EQmOOioq0tcpnTRBrTkHJ9smN
33Bj9WFrhNC5tybj9SwOStB58N0P2XmYWoEdUqj26fMRughiHq7caL2X37cfyW8I/VA1zODw7FTs
32qM3n1q+exd0odmgi5pLRxkG4plzORtloJSDu42saGZKOxOBZG2oZi12yfhkg55Y5mZqlGbsSax
kuXmCuFSDuDcO6GODfnD7BnKTkvcFBcOD8oTCks00vNmEBoUulVbul/XF/IN/JIqk2mwz6A69txe
zOvl/hCtHnC+5ewEzvT6Ipu71uWaficVI1mCj1sb6vyUFyT8IKI0V2L8OffYcfg8yuXj53PmTqwg
Z0sOuFcdA7HaZAotklPP32yC2DwIibV5BvNtgr1KonSnl2pCaTnHbtGmtA2NHfKirW3VsSNKObgB
71pJzymWOZ47H8Nhghfz7yNBT2nWudek9YfcUiW5XnvtWn39660rzs9t0Wkt1zLFpd4BB9t9o2QY
tY+wo13Ct87T2sGkhIOpNDCoviY24Blc6fAcqqL0dwr4Ai8v24kw8mLOVUVd2iCiBCL9MEVghMX5
6T3gDnHIoLXyDPruRU8gzUZSMNCGTcxpJUGwimwcTs4IJ5zdXf64xYbew0jYwsXeYL2A6fiMfayH
3QYSo5+cWtyT89epEWAMH74vY3Ys4fKoIb/9o4hMYtjBKpsWWMgolG6F+gii0RcFxrifHPF/TiA/
+05clYqydYGi/MitGnu8v5397AWrCCC9p13iyEn6uo2hgCXsTHI6yl5owUctZzAdtr6z6gAmZ1sC
0+mKSJwW/Qbypik76Zu09L7Iwl+xjuqwnn1Nbb/1W6GzvXOgFkXmQZBn9NeXN2BRk6bLLhDekBBP
zvc/5iysVxJGcA7gxIbwXjErQjRUXHX7gky998VbgTTaWqy0SGZW++0spfvUEOxPgK/3E5KT/oLG
CecLa1vNm4+cWCe4QjwXm0mFg0S6GYqEk/IHeD7DMFXNofbm8kx9/202n8oaSW+SG2At5np17r2l
3MJtgYxgNj+yv8OJ9+Rq7517lK0yuyTd6cltbphwDAVQvKFnEc/hWWwnN0QEiaIXhKe0ukw4mVMN
OmEmJr9uOEeb2s6QP0TVBcesTBO1NUR5QfRWietwuY0T0njxQPS1WzwUt9dUJme91NTLdMV/t4Vd
Ph0wAXtBhyvZOEfSsm0tHNbQt8tsQm/XEXBXwB8A0IEE1wdspHGdLxcRGhoCCUSEczbMiWQljkz7
nakjVORGBsxYeVT5NvgoTqLL5sj4D7he9slAwTNBd160pZMT+3H3AF5NQ9A14cdRGynzr0hy5L1l
0kQO+COcOyoo35ZsSRRgAlFNwn/mSFym/VAEH6UH+R37cs1WFvvEwFRQ9fYXWPCuJuGrQXiOf+ve
pBiSxJM0PUTbZT5Bj6g1YfGKsin58kDwnEBXMeiUyJB3BKsre2fZGFbfkgZf0mRD44P38mqZNx85
6KmM1Grfns8gzjYJwH3ZgihtuvsnHrpKKeohXhqvk5NT6LS/3nTUZ2yN3QfXc0HEZUPKCyu5O4JS
pfw4gTjMG9gdzsBLc0pkN9K9Q00dJxrH2nThxsvtRtOBHhhGDNK7Eq4C1k/LWDLH+TGwoKcrff21
tikXFfaHsHv5/qCTE+sK18Sd7JRZlFWpY94IJ8pTOeTIIvt2lxyCadJ4kLVmpO2m1We076BnLjov
YZwTUnWmO5N++WzVhGqMqXaxJF5oqcXYyxOaHGfO97nNVLyjxdz5v3Md5ZikulgO0Da+5k7LSOI/
lKLPbqoy5twfDueXQHD1jyMEbMG735DAVRo7pdp08OYBoNsqA54RJAt/yVOZafkO2CwiMfzyOVaR
5IEjZ7n0cseyGXrIy/LmazAUUXluEkIVEaB4DfRmcVjd6yBNdkPVkFUQJbTbDr442Ad/BK92vtEL
DQmN9uK4xDVX16EvUfTcJRj91fOqurhx6lAiDVRj7SRQ8jO8wxnywGQQhJuT3i1ELRRs3Y4pPEcm
72MxEKSTA7N3ZemkJ3CGkViZFoTo9eWtM3wcNokqf8Z8LYSvrJ0CTWED3vkAoXBx4V2fuuWdUtQ4
RbcLMO9z2n5l37VWnsExL0OG+YwdK0kmvkwkZydXtoP6722KJjG4o1qA/0yUqujeHglWu4hRCXFn
BcxtHLpWdJ53YI1NyfcigPuSqD4Ho+vHH7MXmUsUr+RZjhFnAa8mKJgMN/Pl2LLGDrzixr0ruiK6
nVd5yAGZD1msgwDCZwD6+7rbOnJLNQkwtutFFTon5xrMT2516EfxJKPRNlmnjXBnhkmGS6Q3veK5
fQze4ymJbtTuFh5EeqTZ6p6V6Pdc/cV/Li7L6yfCRx9J0fTovSTF0oLdzhUmAcej73ZDxL3jRxfJ
Bs3vM7pkCOLCzJZCEoAzkjl4xWUnXpc4mwkviuOom//zyxsMmNQxVRwvy47dq+6liLacwc9AGMvu
wb+CAw5hI2Q9FV8Smv01q4LDFOquTt495SKcr5lxSVyi2pRiWWebH/zYzBQEORVTrRPHV+rNPC2s
EKH4kQue9AShSW73s5TBzIqtfvzRwF7f0HfwltIF1hsndwjf7v5uPeLZzAfIXbn0WamjpOQimx+k
kshQ4f49tprtYEAPkGvNUMwABpNzIlIvbRuUiRHzyKRU4fuFAyaNJeThVNDgVAtg7RYlD6zsA1ZV
PTW6/JZEx3fn1go+e7uy0egCOMFABN2pA3EJM6VsX8gBf7RcHEkUHtV1qP0fzD42/HvHsJF4Zt2B
k5HfeLxrbjEUVITVKnMuBWdWcFuTirQM4Yenmr013jLhVk/BhVDCvFtS8R+zrdOoIgBH9n+cyg5Q
Czi4Pwuewb4B7gBoGoEVsNdGXL2KqDQzYQS5HPuMLFHhZqFsEOM1q/Yr34fqC8yrUh4ooYnBfv2+
10QMKgI2RKpvPYj7sL4hXGbGvdyQ3c9bl5k/M+jAk6le7XDOOcO/nNpW4CJOwfwR+0udKIjC+nuF
o9DlH1bNXFskDxnzE8XsRaN9/fCTVn2PY9JAGfXukdrziyYO7161ZFaFVv75Or/UXb8DXcWzfhWd
nfILwZ4i2FAetLmua/jiu7gVvPI4WF6Gv+swQA1E+3DFORoidlnZsVyhsomxsd69kV81yDjLEMev
ksRdgnK7DON1cquB3A7nbJO5m3IsvlVuErQt0Otxus3VgxBi2FJc32ltG2n8sxLQ6OIlKKriUlnU
diDqjfyzhjTdCnriZNSADHUN0W+DtCMbL6FNRmaX+f6nKcywqa8qFwalN2xUdD8eEh1WBh9Zximg
x9NmTF2w6zOBaGdG7Qn4JSRYXmvkqylHF0xoC3SwOu6ol6mKkgFgC46d0A7QOmIQ/NdAv5jMLf1n
t1bKlh9i+8bNnyjifRXtJ2mrZKVSUyWK+rQYK1Uj2I+g6CSEDlIWhQiVGUb4SgKCozA6WhKH5hcK
30zCFTdqCTvh8y9SoNVfTHafpAG6qncUH8U78Ms99aWeDKDPuwC/JCwowdm/yPRXmULeHg7tIvQ2
++yIEtjgXTM8BbqQKUIFxxoR6ttoMCjrW8UpqG0rX8vjRq3NcbOY7hDQSg6oxaUe4XtCdqvjid5V
bidTpMVZ9IzTnXIAjVYgP7car/l/g84HUe+t7ZkuzcMop80fB1MCIsm3EnrBTmXT7QP5RHRllUQm
oJEZhAVi/zNiNt+mYnlJePtgq4ZqOMrkX/r8qzC9LSPVkYwX26adX4ksV/qNxl7O2mRemMErPExf
iweA3Gz9gzAmzXKR5tnkczmhcvlNO8AsuYEBBG6EAus+OwqiY6BLshBhVQD1+dhNFM26c8oT/lCI
aSdZpYEvR+1A8ShoffIKbGdHx1Go4eu57iF164cSLj5hABV5UsopPt5gfWKo3Zw6CJlb0/anNpaj
+ksF4Sbwi342bO88L5TI4CHG50+xrTLoPKSJBocgzOCd0QDSIFf7/S1EAaFSOwMVVY7Izle4uQPA
mqXRHG/9lL90ZBfkrbeQKbomS6XfXPD18/175bQpCzI20op/KUnx+P+HgNnTMMWGZphS3sXlLmHU
tMfTHdYA/ROVeP06FEqCYo4lrq7T9aGFwpt44cK6Xq1aUUerOg3jWzFA0HpK/ipL7guVHiGpLzg3
VB+lF+rMGBPldrf1009SKVZilml8S3smDKRinnn1tksbXeGrsuFfjbajYiLzPwwejQp2kJ2SdxI7
WlYPVHW3N1vfdKxJFg97Uq6wsRqAl2KwwNWRy5ODIZ0iCWswiFJz91GjxykXEI/Pz1rHcSkO9K6y
qobgq70u4z6t8WLqRKXC9yTMVN5yYoDAD6ODbrMc5iN8fMfioPFfH9bKicHKH3Ks8gdCgMp8nT6k
1wMH8j73rwoo4eQVPgap4Cf6Fa41FvYY5+KscOtBYj1pZ+jAmiRkSPR3KgkA5aca/h1sf/SRDbZi
Slhb3mWU3/Suiivg10+7WhqeIdmIcqoba93pINHQxQcnH9XLUqRGGstAJscvhOZIuY7I2kjdIWap
QKDxdalD2kfuoM+y/fapYgkd34jjqkgDGxVKQU9ob3iGq/Cr+iOdcQID4r3TTouoEE+xn1VreRsW
LUnUtRiDIGTrfrph56iR5YSFfRj98t94A/VPlfyQdLy9XDreXlrrGXdKdJ2KfTv+uMmog8G0JTai
Tqplsishrup3NvSPhSiTdi6LPuIAc+PpKm/8XllFuEMXq1xQSzKM8fFZIjktjJOiwGMEPqecnDJh
1M2fRD6g7XrdL/SbNLBOrKkYU9jziyoK27PWTbVyx5uN0wyPlKzSc1HmKGFQrYCv8HIN/++9s0c9
7odEVljs0DMj5PpAC06J+8ChIdhqYKSgfaBThZUC0ScH4M+7A9yAgjzQiG1+fN0YUXcL3RpRicik
d7cwQN/7pfv7ysbczFzBlmUp9fIPOTB97akoI/1ysaqeOuEvGa5VPORui4Xtq1P1Tpi4X8AGZNTd
10Pr7d1SwaH8mOUsCMXQQbSJxA7wbLM/LTAhdfqufg/2MdS4crWiHC/HT2MFwyZG4z2qa2RgFhyK
116jXsztxe7aafjlBgJDoK2L84daNPhCooCIROcu7cU5iTg3PVDyJnUk661/A9cMeVquVt75ad0/
nCoCGI7Nid6nPVRelVj8Yipno2Go9ujZu3OVjiu8DTIsOmAITou8Clu6LPqR+kIHDhfV5qPMO1H/
DKqxeyMQXJZSV9Rsa+6rCYa46uDIKnQOdRgrqwtG9CrY2j3fzClk9Od+VSmCjnytRWIKMOOPJcHv
uA/kHeAsJOroFIT9m0GxaBNWmGJIQ0YsD4XcNCQ5/xnkbjsic0rn359XHHjhN4KpGxaJHJb0+nW0
QwcjuVnz7jYeIJO7YYPdSvReUYSdwo4Jp+UNS5M4fg5mPwCaHxMh8xW+TJmE9AHvZBKGlB//M8XA
fnsY8Dv7RuoPXcNZZG4bQ6hUZSg2LIlMX44eGr3RerLtXfcpAzIjHw/ArJ8ZKE11a07sIEjWf9ME
59O9WFU3mRtyLfPKRhBusmLAFJPIdw8CKlmVK9o8kUDhB+LdCCLGcZkEUkX4ZjAtX178MxzsEiL8
IGGSHvcUgdmJowmOPoo/kbFsLx4rIrepC8T241gJzUyVkouR1nPDqeyaZ/QEhm9iFY33bcy8Hw3M
JeiQ4g5RdgKhOEIJNj+h3jJgNgbi/t0NxReigv7gefzr5d/vFXLOHID/eXPa0ASx38tZ6YTqXsQI
XmzcHYXHRGUuuG0vChG8dcMHBLy4k/pSAQR9yuq2C5IZ/0y090vWqG5ZdXgRb/czGAkiYUh30mR1
TMrcuMIbB4K4iwPXWHtr42PT6pojsiEk86nAd7k0Og4fwcHgZvb3nbk9dmDPlc3uKBAZ+CHMak2o
EE/xHdyxjBAhQJMNvwsgqZdbh8J2bu0VMANxUfRrAY+RFSTyjEi85K8+BCUUjJbgn9RfchIuv/3h
kp6WFxEchyauza2muL26u9yEU6WwBqr5fiojzqeEZyBrFzPncW5RgmzN7yvYwMA1qgQV4fu050Df
nft6wZoE2UYrY112dIW1h1GwgPRtpN72wtkXqp75GEUOc3drVznPDSHu6QaRznOVW+lQRsiH34ep
Q+5gqtbh5YCMQtAWVIjNKvCxNyMikr/Oj5OKtx1QbMJGTnhuZxVRIektoCrPGNBFswBHUn604BzX
LybILTGzTbOqydhxiPAd4EVHYA6I2iXGu5jgMAyFldYjbJlH8pC/oEqMO9/HyQ4U+zPv7TQZxyr1
BiGUVnuHe0Aj6qvWJJX5jyKTS8IFBJ/QMEC11Kb5qdA2j6r6gH9cZnJ5e7wraNvmRWAldK1zQS2N
IHwnAft/NdAY0LUPsmZYaH3h8lhiKM3zmQNLnny8NwFub+gpCcdKkjzgr/B0aTQfH4+6qVZq/HQK
FQ0XE8GvMLYrbs2xMgtuE2mEJrxb1AIvakwZWqckZ7VX+BRIkAyHtkhYwsk9FV4+NmgbTeLtVxQd
DrAy2/4TEfPBI8BQmoh5vTVXKS/ZMiQUM75NRKkm8oDr4xgnuG/5GiAGGmVc9Mn6kLOBLq+V51JG
SjpR8aczv/88P1aPnCLdBqVGLwkzqzEgiAN4Y7nvlT9GItp09zTs1D8pfVKvdwYQ9izuLQtYwh02
37yk72vgKw0A6a5bZPo+TsuivNmpu+pH/6Y86rMVu+KO/QOGVs8yA7KmxBIK//P0lseT2J7GJChA
Eh7e1CL4Iim8/MWrl8imwhyj6sDIhlb23+SILWqNymYKo5ikh1k0TNSKLs38Yg+IHwYakaufROiN
8rPN2Jhr/SfuX0nqGXS+ApZXvKeFAbps2BKAKKfXqelxTxxNXAtLXwZ3Ir+7qhyV43iuNuddj3ut
xg9BagRpk3YanY3Q3uteXw44AU8skk19wHC1hN8jqDCCo0ipwigEnsegIIRpspS7H79+ZudDGNuQ
a8dJ9avEGxyVPdjLqtSxmaBFf3PKtrE4re3R7/2GXkSz8U+BYUBme2rXRgmdYdW1lxPLwhOoV50Q
oDFfOxZXBWnj1YijiVPFarNchrVIAffQN0t7Ies86dGhM9ZKrQnKypzzdpPJF/0uE3/JX0WLhJGo
w+LsYdfpOAjTOaHopPBAYVJTGXU+ihcvV3n8ZhZKmkl3kN3r5FUl2T2YILWoE7DfQ2xbVnchwgif
5JS3gd9TArrR9fRJ8pxLobuDXmsyL0Y59kdXKdGCKKfhxKIKvUlaSuApu4OkHcq6pVrKUCojXQFh
mRMTwuOwfiv9Zqcr22txPRdozZXxmEjyUEFO7k7T09MXKLupTY1GtqEi5xxFO6x3vSqUzM8igysg
x8yNcD82AQFxX+/To8j8xRLabxrKnxjKs50YN9hc4xToWwYqbzqmECpjfC+GJuOppEFdoWdD/Y0J
ZY0gxbb5uiJ2cDuf8BIBxAubXqRc9b8nyHQnPIt3KDccwBH5pg6S8QcgJg89flT4JiDbAXC7OQHj
5PuJ5+VHTpS1o33whA5bIwKcjf/WW9s06rJb6/CtgOQk/4SDGtrJkrJX8VzTLeE275RiYrcNTEU+
tqIa3qjZ/cCzyRkRHZdH8qHzf6Ji8RLqpVLdBfntqnWrR63biQDSHJFxDg1X8zjkcKv4voTrNNpk
8gKOG5Xq8+iBBo2VAk253nSh3e7bZb5gpoOJa5+hSPt/vIl/lOYe/SbBmfT5G7iREhmczu0iQrg7
Vb50rX5o6YXGeePJ7Tq4stA6N0bPnFCSeVy7Qo8hLun9SmYhKVdV8BmwB901+91aXoCKLnYoLEdZ
2JQIPrmdlVXebUhHUkHwBe5fne4YG5Mrx0i2Jis99wipWlRL0YreccIBPQDsTRX3l7wYif0mNJTt
H+Shss0AMHRSX7ZomHfu0ySkyb46hfEBNzIUc/sRabm+ddx2rhmGDDgPTtlUGhKYlMglX5CtWfkI
KKXNkfdJF/fnWiE099rkBigtxbFc6tf1mVLoQab32A358ZILGBLggebHcUKJUiBCUTcFMb5PYgLB
68rpO1EEGRth5QyIcodxvFA0h7wC8K4RrkLHduVEVnwouPh9PYaJXuXlwBphgYk0XhDPUw07p9Dl
cB38oOCGD3CKa9KWS96xjdkwy1/EPxkzrXl4WHixbQOrWo7Rxe9eZpxHUFCToNVyW/0sofIXTbGF
nemgota21s7uQ9TCrBbL24rBgYNVnFCZWi6rsnKbsARCOq7sqY8z6l3/91FSc3rP/6iBlCRv9r8C
2OJ8JXFsTcmoe2m5STqv0ngnyfYiFytzRuEQVd3KxnKr5vor6d9J4tF2t+BekAqmjsxUDP/2s6NF
Bwjn5jx36qczpNfUhkehdiPc1d+kQ3/CV/HxviW0JitUSZoDYZ65qezNz9Q/6ZsdimBRELlUVncO
CdlfU6u0eePbYCIl2BYpNN8+8qn1jZMMgaCQhupxoLk8czlzaRLlhj9xuTrV+jPiIw1HjD2XqeIk
PosvboE/xSruiuEwC1QkpKpmrXboLEZHQn4RG18xJ6PZTnSc5NlsItPLoxj7iKmqEefRWlg6Ag3f
8d41ZZffXRwUmYabFcAPEVmFo8MjT2lxVm4hsENY20Yo10NlqKDwKhQ//z8u6mJXN2xd6UEjWu4l
tWyiTaxwx0gS+2vgTfwc2mpncwp1RriV7FGYIkNZI2mnItqXnFQU1TObjuMQXz3deDzyLxqRFHso
ez8XEkx/s+ynFKCRhUvq2kGiafj5Ilh07CH81hknu164iqPYs7ON1AbpGovf0sVQhs0BwURS9AlB
vqsy2qVbWmOP7bIkti8pVu6QZO6m7oe5riw6zimy2jVCddiwl0WYL7vHYQD2CTLOVPZ4EVdLpD0U
QKDBON6bYvEqdrD/AaGyjSzPK13KsiPQpAiX/UhQXJYrGxjOggT9GXfqactEPqCb5OIyvsblSrTo
IM6BcjBBqhT7dG4x0TxbwaJFX/ETSmwfcqi0o85mxpzaRV/ckljvUEAXXB8DSXFtie8xs54uzPX/
awlJr7vLOsPgWkyudc3GV35INty9d6VH59owp+IuZ3zYHT8f4RKzU0/WzWCAXtdYd4RqzLUEzfsw
o/heisxPCrLElRvY+dHsw/9k/ag9iMEILOe8qJHCb34MocXGt4yguCC7X3AUKTA9qs1np2cG4aiW
BIIUbKer9cHpMbbDCBgbTRg/6igkvNaUuQjw20OfR6EpDxTHdrtw8fUk/9QUd0q9OvnWq7AqRp0R
EYiZVL9DDi4oZItLNBWp7a+dA+vlvp2Mh1GUmutJdNCO0g39Edeybabr3FzIUlfS7/mJOqIV52LD
dX2Kp3V84/0z62O44sOFGAXjbk7rK4f4RgPgUcTJFNPWGzpyeUixx8SfpA8GzK1nX1CanMmigZQv
bAVj8oBC32KpSvP6nkjBLhkOr3B+3wGGkblGjwYlfU4t6Q5MmgDPM+dF14ZEpLcaRRpL4X4My48P
cwlLskikSJGpJPKF04aggno5BNfOMYaUiryKcJoM7A/GI27/0h4WRHDtbrQqD0K9mZixfXe0pOz3
Rc5mYEi1YyLZnYY1SjQKKg6f6nwzTfy9vnvpWATW7MPO2svbOfe+5PVS2Uj1sKk/Dw8UTdXzuhZ/
JLrGJ6ISIGWlgkIQ/XcxnECisRKt73qQ8nTPK7YTVxnvOs4Wxf/M/L5/PyqtqLHQggCQ4nGuxzVL
kSkJQcvxnmMXJzWumydQ0BtvEDezX/s4AdDTvJ96SQszjk0GTfa7MTJOVIKM63QEzWJdxDTHANky
3G7rXc/kOlFyAi0OPqWsdNy1gN6fkBCpM64ewBTLJBZQdkQSV5UEPnbgwVXjM/sy4QN7wYdefCwa
aGy4w+DKBQd+PBSeBi2yZ9dtx9EcqeDz0wjUG0C1+Pk0t/plTlpBYotE3c5ieDLUlTzTjyQ8cy7o
gJf4A1TAYXUhG9wLgm6LM7dgaFTFhc8/Li2CRcBTMiyubeJNoNUP9lO7Ds62UDzyH2zUBzHI4gkR
yMTgDv+t7cQ8q0hpWGC/PSA54LERetmohQkStPzCAQpa1gSuofF5d0QONc1SGG63ce0VK32Vzt6P
hlOBO/rMP50THMXztMt28EiwEgH7peqAaHHdnIjQrx3mdnzKjdUz8klh04Z6G5cJ/LXOkb1T5jfO
8cx4qda9E+l+tYXvXhIzhXjdPqx5qFNgQBS5m3I5Ns8TtPiHrVVJEqcUEK9pB/uB1P8QVJG+h7Iv
8Q/H+SGm7ZwLQ51jaoMN9MwjPtutM4cDKFsClUKCp5aY3ofgNu43mYfL7kChF83v+zIiWfWX+8Yb
fGRVh01hyAGKHS/BbkbZS6vZdiI4d1GZcxxGxcGM/r8IFcHqcfpw4cqTJk7OIdXUbxW6JjARKRQJ
8LWv8GxslZeICw4kbCxWql6oX0YcgPWITnsr/kvxkDWX+YE6PNPinvBcqvpV6ty+cgYtFVGYNNts
0coAgSD/DKQLXnaq7uc4tYgySvk5tm5bZmLqCp4q/XoRmbcI7RsdXaABZ0yGbuyo1Dp8Iq7aMJZs
4IMkywrtJJ20wbKtJ2iyy5vcwoyOuls7QCZEC8M5l2jXTI/h2AsrMopAaaXMt9lvsi+PH7KDWgFK
TGrpPgoDTPjXEYX7Aorxxhe5jTW+ExZPlWEB87OXehqm113bQyQ1O5rYzOhvyQSAfUqM/simbKV8
M4fXbSV9eKcg/t+vWXMAG3qokI9KQmeVghWatNCprxEG1gW4mtJzDKs+PxImlEI4bGPznIBsbYxg
5am5M5Xfn8WBFPpXstUPi/dcBjg23S07wIvUOAtoPAUTyhoVduuR0jffBSemyORTykTT6vOWf8mG
q4LFnTJkJLJZddRVxxrIEq3TxDROesy35jeEvqRFloF40kNdGlXqxWoCwM3Fc/gKXGWf2eLb2wJ8
5lFeWSjRJtWMoNyYX+GJ5m2hnpZ7/55jZm0XTHQcTfWecWjnpy7jJeupJQb5ulnHRTWezYXyuqBR
+7gPD9f9jNz0zlg89j17A+L+5kpicL5M2cJJBv9w6Ezbc/Y8q7u6tbVOJoBxuv6azB6PjHaWpBTX
6g1zoMdKy8mj2QQ53F7nAAGM1hRnmwHdM/IVVwbezwR5RlSeiZUyupBACZgtpMt0vgwnRgAFCskK
cIddxovxA7zqliUuKboM5ijir8gKTSGq0A24/dtAb2sDidIwSOsNYytFXN9jdbxT4FEVhOoP/7Or
RGuK4wo746hNk3dV4b5GPW4FZ9Bylki/B/7k2/Mx9zCc8XJuVPFixfoF8iM5L3vZK1gGUy70rp7c
mQN+x5XFgpHbrQdzJqaW/A84joMbu9juBVjmiukCSIOn2a+vEkjkTCqSmqEgT7RPR02KKW+3/UmT
/LTS3ivq5eo0ZBL4WecWucEVUiiqnGW0JhHQDoL4QfGgWPvKKttL5CsE4qYV6hELthHUpmKT4t6X
szdgj0wrMTnZbhowNTSy90vgLVg3/4Yu4Xzso9C9wMKRcvLpr8MI22HTFpWoqA9fKJtBRLZADSrA
EyvQy9edLTK8zEBAUUe0Vy10pLDwZUBk+JIsTy3Rtv+xYSBVILOI+FQFKSGS0PXw9usf4YOAjimJ
e3rJwEqiKKIhJk+g3sEJODXtoDzdNfa04bYzRxATdsGZQsU9CYg8GQ9h1qdgngEyNMK9aHE+9jxm
vNFXVaFHW5AeecPZPXJDJf3WJEXd+bHlieQC0CeLIWSOZ1DsXoExSQWU2poELI2+pPIXn8ptQvlT
2DpbPejtBZa0gXc0aVDBhlUbo9B8wQ5JCh3EG4G9IFBrT97PD++vAp9vYXbBWu5sRB01kcoCbJnG
onM/fDgzeI6UhCZ11iyOZ71CFlEnuCJ5deT1dlNWZ9ry7fSNQ8hyrkt8kXMx8UtwU8h49WQfSKzG
f5ZzIhKdwGPm8XwHZEqveazQjIC1a5KCLQY3bB6CcbxQN1z2r/khTAZ4n4/7CLqxHxzflvFRi7bt
znARKVMeseJlFQEambYuKi1eUc7JluvN9PFj5xlJMWw40dsMNtCdrMt4P6v9YFHHV2uaQKcXIER3
EprS6ue6nztr3d2pEruQ7eX3nr+yRxMZiVTZHRPUcWLXN2Ay+/GTDBjJ7PPGtyLg+6RtvKe+u10k
cLLtqrdq9CRf5hzsC7R6ZIakSpALlh8/k9YwqfnWh1OmAeN491FBFG5k8sabBpGJ47E+tpk4B98h
mb5Y4+xO5tGnadRMfYkzDZHoBZE2Nej6SRN0dZ9jtv10t9IQHa37KauGfIaepNgVqvzy7Tej4yZ+
5boQz4r7HheQBqNV6bdWxeu9vbMeWWdpwOOIIdK+3JO1ksd60ybwDTFs0oIVxZmqRSLO401+sSVU
UANHgwQHGdPjshG2jOz1tzuHz6rssdP9tG3FaG7H+C5XbxZjvFMM8EC1ZFIyj0gK03rw/4rdak6J
XMMT7jlUhJjvSedmUYyg9FCAJ7scXtqiWBbAhN1vrRb6I4VscOucmS9WGeh9pjISYJlX4+5JqjC9
molNdBKhruP7TWw3BpFbYISQgMFH2r0d1GgI9eRbIbNA+PM1wPNdTNG13WcCgSRz9EWaXrJUbfoI
H4180g2TTgJIBZYpeqN6ADPRLzA668KPtQWMSVB4e42a3GLxEN+weL0lcLjFuYahqKbwGB2I/zVm
rjyqxSR06tK2n/Z3SSCTuGHqotZ3E0LqGCXiqf366a52l2S4cNdc9pLV8ga+u0ARu8yBRhLDflNG
iz+MlgYHi4XqKOq7GLQD43D6Eia+FaNEsFSvjycqDCGvMSJX5tTSCt/WjJ+kd015qz1sP4E6sGDb
SjVgx0/gTFaGiqrsqQ4aVYE7R1axRR3emi29hQWAWNJSZrT1Iz4EFPqBm6W0x2XZUJP2kvHAQJXo
p5MOA3nCTndNj3Fj4SAPu8Yus3Ei8jprJN3XRYtr1hwg/DRv8MHpxRFy4oXO3qPQqf20pNqS6+bY
r2Jge7HjCi2TeejwQ17TTzzCMhFPuxxhTIB0us1lSjo1B3tVMOHXNMhn+bCk56ww/0pYBWA6JhJO
q3f9vypBOnJFAusJ+LWu/osE3nFEsby5NWCuqMuhWdM4wesaGBJN5AaGVWB+cLJqKdruORxF2uGP
xV1Y0shG0yZVo5NG8mJDPdW71sWgRXmgJAPyOeyZOnGkeDXdQ6mZU7wSXl7X7b3Fb1e0gAm9oLa6
VP9vTRWhiGbllFacOYWF0mKeXRrafouLqPt3m1dXSWY/vPlDuFeOoCTlz1NvkG+Q2TuyztwUVera
OZVNxZZ13p+ZMdDMj+5eHI1HusRVCvkwn+v9Vp7MNRotKDaut0jjyehChZkxqzq2m0UyqvKBtoCv
H2/LCojTv6cZ5TzQc7J9NBOnjDKifub/7s++AROH/m4Pm8OsVmoD1GHbuhocb1Ak89dlS+kruhCK
cNYKFLh/ZVUsvfVM9Vl7jaWPnaEHpiHJSvGyKROxzpqPPBFXdluPDgqfBH8q8+GjWhT4wSf4CtEe
4vyrDSrHeXK5Dxg/JDCfgwKNmuZ+GVWwwOdZfGJlEA+EQrY5fW0oU90omNkRHYnMm5qYs/vrrAOZ
PqZ469Dz/k6yX2Llc3my48KZbMLTeKoPbJ7yZJSjU+OBOPGfL7mSOe893CJoKEd00eavWSUiZiuu
MKXE0noKjT40huGIji5HGKHrJ1HXfRk+Hrb7TtWE8KXbCxdGV0wb2z+KE5UaPSIvr2zfWr5S3b/B
7Y9H4f8A8cvLydq7/3DOeW0WnVokKAgVamHfz8419bu3cKKEHX+hufRGvOPJ5kFkLqEJj0NPhM+L
5lViYluiCO2EiK6FhjIkR7gD0F6fu5cVeqngcZwVWVH16m9kjyujgxbsxhjotxEij3EkbeL24arj
hfN/nF6k6JqnViHGgFVtkSUnU2cuZI2AeJADNyi8HvwNkbIvF4NCMplkN8v2zpepZ8e8QjNUcoN9
4ZF1qwQOdenWgBCG5FnKte2tIbQEaQGpvoaBXgJ40GA/2OicDtMjssu1tT1qtoQreevepforfHXG
vML5O/KoaFCKSYObZpXgIVecutlnOeGcvDAINchsDFNmfztFnIWDSnwOZ5NGCOX0nZUv3uY1+Ra9
FitWTgaD9GofeI6kg/hbVtuEOtrot93uPN37S1iWjBEbDlcwYTHa7uVw0MgS+zsjzuhLNa3JIYn9
wviVCX/wFXrf2iu2kYOv0tIgPC40bKDBFkQz2PKmNVYy+gHzAKt42Zpa2FepulySMUmAmiBcjaPg
B3mweFWbZNFQpjDdTzn0+D7jkIrKWLVrFvgyXOpjEvhoErkCmaWH5Jx+dG1B40PVKftt77tG5lTn
XSmSpSUslv3f2Ct3YfvkMKsHM5MqZEPLyA0E+U+ycTFY7FklIhHFx0nkpySaRMm1mXrG001au4Aj
ANYe6o2s/Fphyfyd41YwcP72MO3jEz93n6AMr7tFEVWZghvbtPoCHqCEhyFjtanIYQXmAQ4aJ+By
fbubNfhjfFNk+4DsgFtBA7/J4vBzJ02HeULvosWK9Zu+tOFb8QY+wd30ZRnN0KVFLncNXHTDm9bv
3rq/MYF/aiXNbiEvINvuFOjWCqBGtFqVk+QeJBhEaDijJFmvBe5UWNXItwaxibTtiHDl8Bk9Rh5T
5qyBV0fL+o0cisDh0OrMipQ9vbdcGQTYryffMcMsGBtDdYQaXqLtTl/aSRbeAMOmR7Wy/IT3/81u
3g9fMS4d66/3qDoOwbuTre35AFrI9RHcTHSqCK782pIQ/dlLKAQQ0m55qhCUQB32TnZNg5WvH4VZ
1bczsTUP6iso7BtRFlcMK7u2hEFc6Ouo87o7MoZYh8QznCkTRQBni9th/1odU69H/xQFxuxZ2z4Q
+cNUfBl4C4kJ69FTR26BVveGRwDNf1qDp297uxwTO71lTUgA4cR5YvJ4sbTw++HYX5AOhx2zXsgW
JSFBA2e2bga8hIWbUWQ1nJF3FB1S60Emw1p365rd+efCZvy30T0eL4OpdnOTIHocr7QM/tObNQud
yXlaAnFgBZSw58Aml2N3LfMrAvETu+pZ7oeLsH+7WbFcfYtQ3J9Vcl8vJq5xiRkd8jTgXMmpVzk2
EWp3NfwJ85i1W0pPxQjrXvK1OdmkyyIyvf2SIRbuOgmESAX8vH/5bW6itM0YvC8NiGm3ArqEhgu3
8Jr4dyAYcKQXt2vwI44YiD8+3uQvC+rWK9gCUgUXDP2D52372mEmvwpD4PwZNzy+ARQq1ZYUNeJE
GRp+EFlT+snVO7AuOVixGvYQRerKfvC5FnNdZi7jq7py0anc3jim7rZC1sKeG/S0di8eRbYzgfL1
PDGUjOQclf6ggakLjIT1ZL52pXsI0nFJPTmLCBIkE0M/K7n++PcNvOPyHoCxkO631IvHPzVOjql4
lT/ht+tZNbzqlbHuA0KtzlRM5YU+MOtbG388Jlj5kca8IwQJ/pnbUmO648Gam/eTWDrPXYkH9TXH
UKSCSgxpq11iKaIEKuZrrHGOph+3+89jt8MtlS2hc4OLNbH4g74WesCzzWMwwez7D3g5zJ1vkzgz
BMsazUEu8Z2Bx1pDntTmnNyGgfl1PqDk5o7yt+N9PonPdmHrW+S/3Auc6LsI9d0rJQSu5mAAF584
I+OMwnd4N3FF8DvMYxtjCGuZmvhw37IubeFu/VCrnitLqAr3STvrduosbcJVG4Q+0x+Ch0eEilV0
3mtcrsruHXhyumBd3yNOizyggmLOOJRgXZ3O1ABwDQLlPSGcjSekKOhInK/bx8Ixe2HTahqsxFpm
D3XmiLVb62MlyJ4N30WVMrV+qS7VWJQ8hekVs6866a6mHRyaMPTa6HG33ThlvCh8ZIO3OhiHBFuZ
Byo1gq2AJWScLjAfrwIcpVL2z4YIRef4+MUPopu44Hc/FbZfTv6yeY9K0wA8YlCGef+hAsVDcxCb
WXuGomqV1bLMAey89y/RwNbV3D9fXaGwiU4n8Ia4n+EZc4dkfe3YUEFG5A1NIwA49j+SHmwr0E+1
GgtNdQpTEO2CqgNyD0YYyrAndjNEFqhvJToVw9ac/YCVyTIitZS/ee2pSW+lVIyW6xxOAzjGY6mq
mDKh+IcJe6XXA51TuMtDH8sUU6OzZyia0SPw/dr4PND9Y8jXhvEwZCh60CLZMxEd+pkQeehhN9Ga
wBrPPSshsOnnK9P2Wm6dIOSnu3YHfaDloqtVUG4dpRlq/C2OZkgHFHTdlWKuuUG+RohPcDD4C57W
mB/dWyo7fFeGDoebQrQc9hijH96399T7SN3SZnRC9Lqu5F0eFGaWOqaWVUVEWDxoA+r8VnVv2ePE
fSAuyfmX9xb1pO4L8umBv71Z1l8gtLZa5gfj1Y9hPSe68gkXltKP0mdnQEUWx2IFDtXSQ5jKIKWV
2B4YHSQFuIzLbaZUydVO0d+V6DM2NlPGJrPTZRLrjZyJI8XOUtUb+bXTP8f1i0klD71kl54v/PoY
uRUOhMJl2yWBpY34RYOFLPLI/pm7rBl4vToTqScWGmLyu4vnV0jf9ZNgeCaXZ9ckDLy2eOqaTIWA
pvlXSdAPhrSCXucFLksRTbcWhOPodZ7lMI/3LLNhWLju6frfL3XM2fhCoJhwfaz2XoueIp9oWFdX
1DE45fXOhs1Nz5mTgsK0sl80lWwf6/hc5oYa+5PB2NfUN38SbMrO9EUzAZHVuorlUuoNuBlMiyQd
J/jzTU/jUEMcAcaVOyawbLpntOj765a5AehxjxbMqJlUaNTsu2dx9jr4IetlmvN3avnAeefGY0kH
/ddLIib4Wr0sNh7FXpikLTHLcSzY1v37LENgGqoXfva34r/g4Z+lOqkBGdS/deuhwhIPRtKJK0et
4FUsS4zn/nmd/7UUZw6Ix74m5Q8oPOYoYk+C4BwtMDOFfzQQTJio1EnO3mUyNJb8aUrEl8qwIAUa
GalCL8iuamBJD5z57G0ODDZ+CHfovv9z0xtmnASvpY+naUEfahMvYJndUQ656eptCFq374Q/vHTj
/W0o57YkBYYm6X7OAyYK17gvx8XqY8/JJWMtVEpIeFWJTthdY0GzUPCYHa8Yx9IxqrIOAdkcBMtB
FDZWrhEAY23SlwJ1MJVGA6yEL56nfkO6gNyVSehQtoYpoQzarY5G/XVO8F2GHQDFDrKH9VWRADmJ
a85hTbvWl9EoEHdDIVwPiTgpJEKskZRVfAKevA/ZXhrv3FkJf8/tjIqiAdA8zygfj0reQsQ55haw
2he0y1mSqGs2ixtxVX/SNCbMeCk24aSdW1hhrEbG3sTgxU3ap5b/NfJtqDyVlgojcr7OU1bu02Y7
rgqk/qZL/DJKMiM0+kAF+fpC4aDJNOjH+yZMGoqOdRkd2wSVYkZgYHuQsiIhf4ayUFZekH8hVJeX
WZaWIEX5QVXI8R+aAG+u82I6tz2omTMYhb0NHCxW3LnJXBrHiCJe7OWLM+UxC7V2IpY71ekrlH7R
kRv1XJ44zpYRyRSXnXtqjYTEeDUlQrv3+QTQzlUPgdCVjJwyRmyUjgicXQZJXtfZpfH8SHtevmNs
PvIwqu5/PR7Mcj6V+yBF83tF9b0Jv3IVJ9oWOYHba1fQCqy11G4hHh+h2rN+NL/nFm6nS0ZzuEdT
cV7XT6acc92ScB2yia5RFyioXht0XA1t8FYF/LLuW2IVtKjmEdJWGeOMmyy/CbzuXhdaXAy8p/Xv
jboOr7wPSS6ixCqp0wU7z7xhNufbueD1J8W+gXSUZuPp+2pIIiSOI06nwQzvxBqm9zwsgRRiz2QN
LsC4pG9JNSd/Gu+4u4Om2mhDcKqaO/uF0Uas36MUITURhZJVNnVvkqVJVmGHNe6f7eUJo6W3Ib6l
h6vpe4iiuJpNQ+jiIrhdaMzDwo8994eg4OtIU6GJ0VRSrRcPiKStiphBOb9wNv28ctCzLSYi76mb
uz5rZT1S6uacmlismth6+93u+ryskf+qKn5EsJZOwvgU8wCbCyLE1E3MeewNfeGK7wObgGmc0lo6
APoEsmN4LB1adhV+L+1s6hTIxXWZHhVDdAEAoROsLsUQY+Ui7wqLxrjz1o5Uoih0JYZi+MiQNEOO
zEbL3mqEbKMU6Oh8ioj6BOUXQaSNm2fO++juMPTuegPSmzvAX7yynKk66crxc3YMkP8gWnP3LODA
2LxNyFuHYrAsMWzWSw+SDB0ZZ13ce3sYRDP1VBzvxFHaIAe1CT1Xd8afXdeFz/b0DzO1RaMjHZiv
qXwtcz0d2/98rhHKVMDCVpQX8xvkVGUYhljHSVuGB5Iz6C14B6So3wcXn4L/x8RRPhjkpAMNiMZu
jTKsRgmopVHeqUNsqR4uC3KLIMb2A+0W4j1tWDJX35hserSWCS5rq8OTobbOnMntzhUIWcNvXTQ8
yrAHYKN68waAlOfgMhjhBWBrOnHbNTQq5GQPDB8amjueJV9u+ORqpfOsQOUck0xCg/ZdimJw6XFJ
FTGlj1g0sQ+U5IkZl2oLzmeADHYNc31V1VhTF3nlPb1ed+mJeQA4B4KK7wKCedZoUN05juvMzKOE
lI2HHPqDH6O4u4wU2GlYC6WG/mFQobP8CQUR0GndXrqJhxK9ofljq43lOb4SLJxc7nt+X8wZ+lt7
UssesplsdFZlc7VSqsv038RTMfIFV4ojg5ERtGU+3DhkSY6RUu7isSwsIgjB5WWou/UpnAboPAF9
ASq1PHHhGpDzM8XsGj2sFZVt7EMkysg0dbxqyeGplTKdGkLZZExI1irVklPiO+cX4LY+nQEn6Rjk
FAtwChiiy1KGWoKk3kzGWuFRQANrpLXkMriaeHNRqotdFS3MQfDeDoSY8JCm5nIC4Om5jh71Mdsx
27erA5xD0eRD5R0Dizd+pWZFTlBZW+aVGVQMyYRKvmez1eN2mrZMC1z7Et96A5fcT8sMdQXxQA2H
yicJ9Z8gREjhwbklNLoCoL4xwyIMqZv5HZ1oCt+5tE+/ovYHv2DvLt4IEMAHte9dmoAL0vtks/Nq
EHGSwRzOO0JNmeCA7QIoDal5gs2TgFPd5zDMjN006VWrTPxNCCzO08z5bIPBZuD8xrGnj2ugMk0A
NZVpjI00ysD6W5u0aK58Yf/bm0X7RgiM60fUGRxJheoZjc7rwXkPdDGjlU0ooeJncuA7E+/0bfXd
oNox3SgyJ9vxr4obFiO1iV+meKb8iC/pHlV4pVDWPV2YJ9asCDVYRc53PFPn5lcsykBxAcxR/46b
qx+SyEwYWe5M+GIA/ZVYyJvU/nWB7jG3iv7Ie+N13tiPz0nyGFishJIbCyTZyuSGqZM3dWYGdW4p
WI2i8SWGLxIsdMDEgSe7hyfgFCw+wBISoobnjoQ1WJmCqDgaXW5nJW+n9IdlT8MvOvloqMkT1rPJ
23tDbmYhSDjZJ1T2SRdDlcS4Mszwu+c8QA+dJXF2j9Fw0phcMeusZIGCLLmw++vCEFJcmlbl1BML
WR9UzaadSGbDM3P9Ro2MMis5AI0whw2y1oWET4oep8zfRqWnoSvwvlLeYplfSYRenykdI72TxDOL
Fg38nI/WUnNKxvxHBm0Elp9AS26ErvWbMpSpaCO3euBzVhWSiuVPh9xa8a5f3xdQzo/qvlCLXfmE
InNi7RiuueR+cUrxCq9S7UFMALl4fIcBdrnAzRulek1YEBsFObTJHThsrWts7vEPwxqdBSYJuTHf
Tp72oTeZZlYfAhZe1MaZFj8vJHGXHP2vu2BcnzIUFTw0xnxEoPcqvEvV0HPLadsAOgInuqzCs3Gi
F2R6dJlAzJTyFGBMP6FL6VWj0ggjoR5/q2oVuo+uTayq2aiVsYrdQMN+mDDZid96VBP0ZIgjhwWm
LAcb/6044RD+zljWCsOAp4kRxXlk073z+/fwliMpJaqfDAhsS16YhwEiBC9+eWu8kHZ0W+klJrl0
0en++h8GduQCXE85Vz7qCZLN+kmSj4M0qetAEDx5WiytoPuJfvpyFtX/fj6Ps/TLfOcCU/8qIfpp
B1rqN+V7f+YUcNJGRlLdlmC8ks0QyV1Pe74eptjK1FdUkVmn9G5lzvRGMSQEpHkrw9KGiFP6q0wk
Lf7YHl/Z8AvR2vrt1xBKn3+P8hNOiIaAu2ATgv81S5Su+kSlaPBcWsndiUrQjiFIFrN6OVfbRP3O
/zLlI7kqZlHxpUp15zt5eR0qXecFIq5PkBHHTlVPaGEeQFYdetq+NLFKGEZBcUKTYdegp+cfv/xm
smzaGeE2lSgt955Yk73JAVx2C1E4LuHZHG2QDTHBRtK7L6UNmr0bYSBqiv9wbBFyMdzxb4QpUd+k
wfWMBnLQ7mD9UhI1S1T+QJe7vVJ6OVUOA+ZktGX8CLeNMWP/IWWhd/56OeN3StPv8A80P4YS5YrY
1OWDn4w0Pgi7hqgpvRYALwRwF01IZmACw7v7LqTPmom+u0oYZnmCxjvxFN7BV6b/xA9MV+Sg5AyX
EOylt7TTF0Vq2uECVp2LfkOJuCzp8GSl0F9IHVhVagsPcYpHWUMkNdR4OwEBwkIYiTW2BnspACOp
4etmP0eS+SxLRdrVxyKl9JdGadO2CH/3EhubK9y3cf3aiDtEV3Yfyq+BVGpy/jKXce/rR9xkiXXU
wI0x3MMnidumaReU4XGkjY5oWazb0hD9JoiONTsmx7mie3VRq/i/dUlsV+DhblSIuOwReqYP6uOx
uQci+tMHsW+v5y7FV/zta1ZJAi2HR3tmMnBvBB8VymVDRlUW0MVUiphWSYktGZwYswR2vQ+AFhe7
4MXlwKzgAcaIkmzi7jZWOvF1gvTKFqUhqKDI1f/roSjWDN6lzyYlOjKTKekRgdoXSb2quVWznHXe
bWeNH21MV1Bs9P5HHbyRbhexykCuA7tEi4dc9y68O+QwJIKP6EmgZxQUEUS8fhgXyPBy1cIzI1R4
RzFskbRpZNhL/L+faEQKH3zMZIhVv7hysy6xH/6XaxaIE9dbmDNdksU0K7kd0HwJKDUbepPtY7UD
meiRWR74fyso1s28r80jycjC9xU5ndQi/E/qFNraOs9EgH7HF42VjehyBhKyj7OY2pWwJGirUBTe
/N5pKXni/e+Fy8IFjdayaQCt/xUvKohMIrHZTXl7AEgwGW8ZRPLRroX5xHlYoi3pL6FBYWopxeBp
angZN+ZpKY4bB4I9dz8J6FZTlEvwNMKwGk1nz3rlMtqX1KJt8/N2MuE6P2CSIw+WjBVsIx0g82z7
VEl58Ko9a8lV2vmjjUIoOP3A55N+Pd64cUw1/7PHOexqaapUGRQ5xiq5hRSIz/VNqCdCczIEh6uf
PPjRf58EKCuc0V1c7cYoph3ce1zuT26k045LOVr/VjOSzw+7GQ9Y8/KOcMAjLUw2S8x2OvctZOGD
gaeKeMV0Y53X8wiyNFX4QCxmHSrYTvUoIZLZLjtyrMv+VmQRwGyYowqFKeV/23yaxcsWFKIMoOjP
5khD5LX10RgSrVHK0lqm1SPufwoMsRYEygEYrNhow4JhrvkO6DL1IrdrZliID5yhaJIoYi8ulqDo
NT3y4VbpgYeooyg2YiwFCFpEltR7dKpRhZ5uA01QBFuJ9ILp14eH4SvjQOwOSzmQInBpaWoo4e0M
QWjLJRGVJTeexqifMPGVeexMEYgrOLb07pk2pMdjV1Yfaq0aCiwBiNt2UPhssRrBM87w33Y2pZFc
seIVNshdCrxfQ9tZA4jdoWtePlmMAgP5XmRzosoxmBSvo4yD+iLXpP+QSz6vmU/y5+cHoNqWu+Hj
6LOBQxmlOc89xUvWBXd4141bu9/adz3Yvd+XI4Ei9T2gMZKQS2TWDcqAZcfVxZVXh7W5SRXDMkkg
13lDMZwIT8kROuEi7X+xtS+O6Xv80vwaSlMqJvLNxTX2f2+sysJyXrgUPotMVxcg/mgEbbssv7a1
ySmZl6nIq1waT/g9zKO/Dvo/kZMT/RSG0RdYlviNlfD3Whn18CUK7k1xxgglmkOTOWMFd+1BxRht
FbBBSsEIeEUA8C8XjfZBOTGNhcQzJ//j46TBEVL/DyZqSNBZ50OAVdfYYd6YO9CgFmlVIIE3433A
H/OgpJA0DcUcnFgZ60QZZP+qa50tQtUWw2Na22utgTcSWHTV/C4jzaYd4M58wFflXHA9oIU6NXIv
klNcqjzjT+Whgd3JLdh1/i4s9P0RW3ETuBbjBtwVzJO3svgONT7fC884X8LUoinX827v6dmIvwBo
z/ZyYaOV0gC65duddIwpRTFEkZ0ObOY/M8H0HPHfS0mkY/p47uuJpHOM4ilkM4Xp7I3gxUgJ2JaI
tEnwh/HwX0kzkyhpM/DN4heCYeKDSbbaRwnF0wbguDfsuzAhkuREr3g9rtivTturgGNbIgbO7q8Z
9zhh6QWhNHgMMOFafxrQ/aB1Vv+Kire/4mieDkvexK0Osqq1mK/LBR9C5e4DaIiFIxKNuyIDKdnG
BikS7KFUWNLPyY/lHcDXRLkaf5unN7gONJbvECaZA7BH/D5J+IqzXt0uik0ih37bVprKU0LhLSBV
IzD0ket3WzYJzOgmJpNgAzoCAZIgPIIqtXKBNTIsOgi6AYyfHv/8vTE7KLzG/EWZTb4u/jITw0IQ
7cphU7Vj0BLEq/p2XiWUJlkWvIthLtM7HentEy395RGfId7zdGc8ePtMXlVSSNtvw+1RB/+14ani
P6WBr1lUzIgk5L2PZsrhVmg2e8rLg9EZIKRoLPvYNWklZaOZl/qfDy34hG7YtNsc1Cg9y0wWdKn8
AfFTNuUuTOCO1QDEUCXM+WyzSg/kO8KCQOB4HpTcoK5wVOK5r/gTbwu7sVCqZJvs4SYXvRZRBdiV
Xj2oFdom62yRNRnC+tCIbf2VZDnqDDPyvxufD5bOYkjCv4rRKqVJL2jZ2RrQRV96i2+WuPG7ffyq
6FmdYiUZ+56BkRIQeiqXElgtzTLi+ldQO7roSPufLEaQN9oOYc3NG6KwwdiCp+wSOzTRTYVc48XG
odVp2oQPftn97ZKwMi6B4ltFWq1jme9FdT3+KVSqSG+rrxX0Xp2gHmVssSfKT5mucf/kkinSiGdz
+tM4sO065y6OyDyIFwSL95zwDO2TcqCGQ5ed5ziqltUPkAEUqFs7JLYg75Eq5uUgLOvahE/iQ5j/
yPWLB52/5IMfUAo6eYThSA+uO/spOW9zKecBiJXeNcjEj1BzYiz4NMvJsyK/DWyU6pJ+ybuvBG0Y
vOPSsyRPy73+j/wSWX0jhPtfezNnCzdaqXjR/0PqNT1ZIUhaplOmF+aLgqf/v96oUP3Y2dp8Q0Gv
t3gvgbbNPK5XblQDEaRFbTg5DfTOPnG+9s85DPito0l2hwlLsE7Mqkpc141XGGwJBNGEJ0JJqqMQ
rToyT1fhnfFd23B6itSLr8b4s+OsHXO3HACl1htOwx7wQC0aLBcD92gBvynTr8hAvQeoOgkMoDn5
ZDvzL0771hlReKbaKFJEjDIDYFtD41WVj4rEBwhVIZ0gRAat9b2ubEyx7Wq0FxcstVEahcKfVsK6
6C8xemkUNqV5L/DXWAsKDz1tXGApJdF63xZvmz92lXclUrI0WpqKK07pqzoIuBbYYHtgpdVWLB5V
QFMwlXyjIe0a/UyjTM/KKuAGfycbSZp0jFuXgljXiNo6yClGNr+HauEr2cvVumhOu3m/utFpntov
YrckNS2inNPsNIj9HpWohKMLRSrLFJwuUqPHOFROGyECw2ErJYgWPK8sf+7Y5EaCmoWKurpOpsSl
DlROKA3KbGjrUWVSjPysxisSaGDmP3McfLGoX7HydKHFk7qHKlkUNgqPoRZxSU1m52Y9Bg8XQOOj
RK9jvspZ0rVlDvxPLm8dtosgBEaUqRjoPHhMcIT/BsS+dheYA0GRsXaSubPTvN92w2OxF260VUlM
3khK9rIPe96Ns/Fu3A0QRBGDSAxfEB2VwMGxY/JzSxF8w5KFchE2OU7l9xgIYlgWwy4UOHigEQU/
jVJXeQ+aKx6UM/D9Bo1qhKWa4QEnDyFQBOM28/h0IIVUTZ9Qow4LMuuGmcwfcpe/nXDEcGgnHXw2
rU4VHWVy19hceEzBlkz9Tt08LiguCCnEDLxLDzoLADt/Omwv9rOmyFLUWUEnvXvBkH22lNDyoTqj
v+ONDFQnl08CQOI6I2QtlGUNj9iyQsdOjXLu4Kt4TlUBYc30LJXDItGlwiVcCQZ23b3Ki51QYMQz
ZfVST57dOaCyfZA9IuqF6NCX5TT8YQZexaZMfeTq+rEUXLs8Xutm/a3dxYqIbH/R/7FuTGy+4YMU
dBXQRV76+o0epQKR/JLuEmggfmzNewGpEVWo3mD0QNgI0qh8ZwSQSplQfxo1RoFCSvnYMqwtHOMI
ZaKEQkkcQQlUMkWRdZeMglOLpTnWbtKFSX+W6WHWmayIfw70SIwmE0UYOYvI7QZBwQ9aJUsuakW4
BhxDm0Kt7ljPUy7pAvBX/axjjld6l6LteHkWa3wDq8vXT7syrj8NdukhTBsIBJNAttLrSpPHhvbi
bk6Z65QHM4QuD8NBQTeFSuE6wR/dn1NE+KMFnCJh1AyxaFVRvIB/TAFg+3JFVVZBID1alNqb6W0G
QVlFCXCt8RoUonqRzzK9yCiMXREfAJmB86+icpNn6HoA3Ild1c0JC30l5yxxJ0SUTDEk5CHi9U8U
/NIw+ftO0pX8FDFtsP85qH9I9AGI/g21cOna5gs2xlbz50nGeQKk+xt8I2739b9XcOPSTeo6kZ0t
z6cMyCbHblo6T7S633bveQ3WVDIay6MJxX0X4ZONoAO6dJUxxnp25fbPJFuT29GeQooNxz+414M1
PH4lvx7CT3EgLHBwCo7lyShgFkhTX1uQkKFK15Iq57PQTWConP84gTfI06gKuWFZyp5vVGU5rXte
q1OmDxOSJSJn5x8xS7DecoaQgcc3oAT8+Fd3hkGRLd9/droVwhxuJm4FievxqujMlLU8vu268nrf
+vfCZ698lz+os0sm4mSywo4INnLJfYTXoz1lUKERXqjVF581kKFaWm2jDXE3/CZoOj3QSUCzYyvI
Zv81T45YaR+RtM1EGcrVZdQ46ZcGqi4vhC1lKhr/31DByQSY+OUxTlR4dmJzfz0W/JG9wX8RR0Tx
Tuf0O8YTsYb9LBwObJFAinhWMrFmk2qP18/AO/mmKaVa96nNdinFfSKG9bPlelmbtWI9QfzXjzIe
9JRZ4Ra9S6+AlmFLN6ouTjFUGc9IVE3a4MoWpBuO9RgFr1rMwogU8uPFe8pKPgQa1Y8MYK2b4Aof
GH174dVefA7qSsX3XW+9sGlbzHPAL975oGWRH6tx6HyRtQKLDCSwuNuzzSKzB96kgqvpDVFy5IvA
Uun7zJ+vcSxf+b93kuCeXu+AEob/00LchK9TV03o/HMJfaLQFBEzsClFuoMP72F+A5NbCizGIF6s
DizP7u3r9RXjxyHMwj/vv2uDh+/FvqUYJQEabT1Z2/68CcomUclt6PMJX88Kc90PrTOR4FcM6P8f
Ui9Ww7HYLQpV4XVYN90wtpM0rX0/BUYLaCDifYUFhe7IQPGglMnu+3wAEB4JUQkxgAD9io0TB4/C
i0JBL0ObQyTCwGPLsYsYfgZnK8D+1yPlwH0OaV3ZFV5F4CLHJToIAN0xfOmANbhbc4fD1Dj242Eb
Q62AgkDN9XgpAgZkn2HewK9lCFp8bXUwaUqE66yXz5C1dn/R7vLrG4juB3Q3gnP+cJNUpshhNPTH
4oVHDnmfYGMqK7zD2vcL6K/cVug2EiP/wuo9ogSshL5SrI1kqGM3MhDblL/4dMWO4S01BobHlb+l
vNleUP/yuYwDycAW/JcqfwaBZ8q7xfWkavnTsSzxdQRWu+mGPIqGBtodL6/mqqsAzCBuVpdSYi6X
e0ptCvuFYGxqB+S4W0vq46efNnZN+IkvSF16yYKJxi35IbDh4vd/mDoBkBpZj7BsUkyWpb3mR2+x
FwTPvsmrHuu75ebsxjYLhBIDMgQATDzx8cUqJnGqKtK6Q+VXcYLZ/4mC6qG2J4Vuv/HuTYGhEK+a
L7GD2NWjuwqJ44wCJIRoHLKpNUeKs3tqyEnk2iC8Llg78Q4rHxDF0pnlgp8lI5ZkuaZ3srWt5beo
HxyVo6RfKdZXVSarBkZGRYpUiOG4+rxQQU83xnCaszOLXUJBK2vCdslddud/VC4Bk16YTR9Ez7MD
1f/2CIjM1wqbZ097IsfSjSzlVziqEY9NaPLWAUGnY9OT5ZxCl4hEC6hnttoVu4o2fJstgSRfp0Ss
ZvazOU01AgsgdQuNY40Wy7YbxlusCuqFvjAvGsd6G8nM6aS2wH8OUToi1ul4xuC6rr/JyN2fZpQ1
aYx52wAEN3v+x0pia8k5CXA1iHtCZ4uZubIiijwjJqqz52RTOBL3EXsNE6MCkkT7Dx9piM7oEi26
onL1RMomCHh5HHWQ/HFZ5qEUzXjyMSZdlOZqK50rKfeepKDNAKV8Mzwx77KMSC+taHhPUM0VBhh/
Z+OEc629oxMjThBaO4doonvCOOLAptbGWjjpAUpD7kPtSUXXQaYX5iqTNvXO5NVdsuMnu8jvPCZn
kzk8iSVUcGz8YJyjx4ch2HK9QWCMAD2sPno7ZXIU2wsZ2BnNSX9nRfXSSeQ1LGriAj6+AAReEXaK
P3lfktrC4cAOpEdB28JJEs51yF4gOdrxdzW6MjiZmojDvP9Inmkc9BsnDTVomYEtJVcB6P4Q2GA6
SnALSGYqtwTst967gxqVdtjCog5FZp3ilXWIHpMFNWnXfM3fi4iIh5tsldWgEuoo3F7d/c1VRIVP
ib6jxSvGIZt/BJY+7I14kCr7n/Z9QTBOhKkQ4LbXj6LTKPet4VqX8qCxUEUfYZHscURnQ88cQZfa
vbELlHi/ASzz18SVBV2c3oYoWJs2F3vENQkwFoayWvr7ItgRAFLjfo/a4LDZBEkeLzsMzxiaOKMg
umNlDoETkE/TMfUfnEOHhcWzjKH49Bd0M+N9N0hUwvFnOlK3S4YKC6xfMQyrvg/N1r5I/+E8ETm2
Am8ktW6ZdYVyQc3gk/HWINKkaLIt7reFukIKOwWyJ+FKNJX0AxGOhkKZkU6QnVv1AQVHXDB7jHx8
vMFc9UGUIDYgEHssXayMCrIyfuWkb6T+PK80iOP4YRwlpm6PStzAYYPxA9tbMpmaVs3vCevNTSuO
G3hLmiBVDKEqlvuVL0KUQ9qmZm6wMMoykjjfuwF11HMwivDCnWSAdDTqEBaFmzhN/VIz2HiPiyjV
oYCUQfocHCsuOkeFErhqafwEqrVD1cCzN7VZHcGkj0OgH1CBQR6iSz0+jwVdTovFYqzhEXMWY7xp
GByfGcZaMPUPm1Mb9kx9j3J8i54V/EZRAjGjn2TjnF8YxZ8d+dDFtILD8iu90x2KFTOfwPita6lS
Xqao62mnzWXqPfY7JTqzLfunCx75WAdMvKFdLuG06ss+aFjg3m8SFWmpCEhLC4FBvMi75OhDRg32
tNstivjTUWoWuiubusmPcETKQo5V8PkGKR1+e7zc29DDJHCTNKiojjy9Qy/6KD90znmoOzcKjuyl
SiIg2d6MIAE86WSrX7n+SDiUvhGgtpqwOK9GmXaz2GGVnxHJNhpZYE2V6rVDmPxxIdKdUcOkGQ5h
XHp4z8GBlNO9pLm5taGUK43lS1ttJ0wQ21Xu2Z9nHZQfbP2QvwAA175QbbyMutCBleg6wmlEOpBm
oCKFtR0znIPlMd7CBRoeCp26ta1eXiGxzAGZs6FCBe1ZVi+D1MdM9rJ45JMBmCt8VtlXkLl8D3yK
Yfh7jy3qmIiMGWU3By7OJ+efIS+V7qGRpuOTHqUVNA+3WYyG4irqH2ya7CEe+nZe4JaCRkT8EAjl
V97vIEVTfFqGoseNZXIByjGXMU1AqHLz+7I/bLl+HrtAA1FhW+JkwCZ2ckEQlCDw/HE7bJOxlIzw
1u39SC6fdEjiT2yJuTUgntqkDRiu93d4gwwcUJqO50CjPu9X5ZR+kFQWmupLMiB9o4CpE2ztySx5
cCWVNCJHLocdhg0lFPnhcziFRimGaQeHrHduZzQ2aK/qzyPDIfiD/eWu43AukQRL24wSMv2pQRS+
V1zQ2V9pDfr2KRro8LA1SgiliLc4QR8ZAV0/1l/LDZZXQ7DLAhhKfHmcJw6ep9/B3fVfmRg2BGEn
hyxo2wiSAAwiwip3XliYLkEGukbRjxpMCPkVIwLANnAkk9P+X+wRtHFdIF0OHkLuZmC4voqwI2PW
dLceNaWb2fI5D0CKRNGajdH7GIXP76j694DY475w/sUaT7cKd3rsmH+qhM8G/gPv6ECK7rSTslra
+TvhrhNIQ98dS+yU4vL89HF6wnUdL8EKc8no/9KkCAyVMwYYIo7muYMkvMV41l6DOWPGO+4UPnle
P45T956kF6UFqcSSt6jniJV1zzqatE4ZU8oR0uTatU9isMhW88WbGFCW8nAKyTOx6R7R0qVVF9ga
/aG0zTJsu6tt6I2OsxMkP3s0Fi4op2k87ZKyngpxE3rveEmaNfuRuNqccRcUytzVUBrcp8lRO61U
37xepcSdYxxIzpc55R0SPnuKb2dCmf2BVJ3zQivimdj9LS1236LlsdBIPW4BGI9cU35pyFaNc5Ze
tMNTq//YUyP7emYGHVQbmM4VTYrGBN8LpeTeCTxppB01CPrDmNaxvBlsZJPHa5rAF0iH+kkOJc1F
RTwM/gNpjWj7nvBAFXrfGLPV1tok0xJCEvR68RWc9Aly4G0PU1Q5vSYP04j1T3izDrphWdvXjcSk
NeDY6KZCV+weN8jqkkdX1x8iU9zUnmE8E+GTulTumUSs00F2a0J0/8uTLd8lutNr+R5JkRirjho5
tx0d2RGka0cQNt7hpDdMVKSO/xFHNZw7N42j2wG1PLdDoBQJPK2O09JcvcEvCE6YFyRPUY24D79Q
Sqn5QswmWyPsKLlsZag17HraU5JqmtJKZR/PlV89Oqm1yZA4Kz74Bbaynmi4NOtwfosPnXrvAtee
vYG9WigRYGLAUMgQ+rZqpcqLErD22j0JLBluL7Lmxy7oeDPdoBQeJef0SwTee+nzcnsHn38VdzDh
u5mJpmY9vORLib1N5p7LCBW/UWgoktY8Hnr54xQeNguYnYBZQy8aCGHNb/NgByb4mwcvUpPaO45p
67iTvAc3cgvuuVLr+KDC1XrjtEBzpgu/EzHapi3Oo7wKkTZnIjZc5M8yKSlaJuqh5RM5DYShipqU
ta09ELbO1kcRK9lnqxXk/5ZGNrDV9VUa3hFscl7KOW5LKQ6opt3+m56/Fh1t9ckN6vFNcTQv8emV
0hgxkXf3XQuxCFhy2bj2ojpFfdRUToySK4PTUoakS43OoCRqMbnfuQP3Ol08vf2+d6U0IZfgMpVo
0ClRjy3ysCwinJeq7ddvk4bibgE8frxfP68xlXCCTifId9sxmyXuOdXF+EUco3NF232s69+rnyg6
YKbUI2X3bMOGqcTumRW2uYDT1QdogOq92T9pGr56O0qUXbjESqwlRnhJFmxlYvlvC86A+6BwF3Xx
gnZiHpazYDzoDi+9gnbQxxEcC/b8VIGyazDQXovfzE6vdBZtNb0SVG4blaN2pc/zvK2bMHw0TWSQ
JgkDymDt8x6FcsMYWJaacXsd0OIKZpLnAVy58J0hdssTOOKHKch+EacB4oQSmcFu0zjlduMV36XG
zTamR/Ea3+o37w+IKinbrSfD6xlQvKFxIeJbK2CAqX3U1l2sw/jIXDci/pMcsuM+a0VUHt9+m9Y/
h05ofQCG7hOVFP2M8MaZrtxhuiwkQTqjRWxSccwR62zR7E0JfN0i3qDTwXn3gnVC9ZISBICz8h9R
wGwkXb2azwvl86KGHfpJOpFz7mDKhAx7kbOFEbTVt8r2t73ygkA0LTXRewBSR8vPLhpsYCP5T5kK
BiyaXc/4ToeaU4uHpLm/H5B/OY6wIU6/k8TIaV5TFbpIXVm4XlVNvKitqKs4gu3OGp5QxgKtHQj1
JbSQQK1O9Kbt0rWBfnHVAIAWuqLa7dJJud75JFKkl+/paAErdxwXtrcQGYQeI1lfWUI0YdvXBX2D
xr3i2TbowOXH3K/fBH5zGJhUU4sASz0voj1p6kIITpTyLz0IriGlWWog8CTEdPQNMG7IqzEJKJy/
WUQPEMNudyCTHzPzXasZqqGF5xaGZZKATVcj7th8TOVUbuIdG2lDMhk04YQvz+QM7/dtyEwt59VD
TnjZoPYCBruC+VQ6P28H4W4dZAafFlM/7yNzVNjvGGgBnt3QNFlQqjmFQ4d/fZryg3Jwe+ScmKQ8
sAmGFh1uOtuFc0feB/0SOQ7UwjuyWlC224t/HyDMYJq+9pFaabOR5sASFN5TdoBm/vGzgY192mwZ
kHg1LP7U8yP7LWc1oRnq5m36NNLkS57Lzl28nkZICX/IaREe9MBbRQZ95jwV7XaUUbms+HZhzsq5
ZBG5jtNhqJdXQOJxXBvouVR9VPFbXt5FtyPBwsJDQqVN+3LxrE692ttcJLyuWiSKj5mzf2kHGoTh
GNUlLPHvIWLfVGqymaCPyNrmDYP/YGsZ/6vLAeDDFgOwZjIi0RWPBy4zydwifYmbZUWy0v8IJ5uh
BxGHX1KC5Lv1IJshQISIY7orGe7uoGpz4RexYdhiaqU+9xCPFyjau2ecvCeyf6IoVx9XKJWclRBo
6+R5qY6ZZNmsUf/KpvoPpBzGzLE85YpM1VcobtEflo3BpuvCoTwZYkL3sDEiZZeoHG5YsoaGtu33
nNBZS+5QIWL9Ee8Mi1Zhz14/sMvLfiE5yHikZjcAHpzlyIcsijE2aWUAjx56SrkPy4pFI8JxpVXg
8RQaSH3Nis+X+F7gt685B6pZspF95SOYWdta64vkLJAPCYODMsPKeUWXmQoSvxVPh2Os+Og5UBe7
teZUBOK8IehmI3Bm8np1pQ4UpeqEB0yzG8cWXLc7Zc57+vWNgXiCKVCpohCQCNix/9U5PH8xB4iD
B9xWx7RU6LmqxrJKrpP7NuagVZk4mNsdd10CusCCC+KWnbGo/OXuMnqaPevvlFur4XZjFyi5+gDt
DMEI8iv55PQA9hDjNMZKwtp5E6U0t25GKhY7bWcYY3cI+ZPpMh8jVZswyhSlwdofc7FTFPsNDXfs
YfJSHYaZUXHGEQEE2Xxyu3oySq7x84Vt1TE87Vj/52EiNWs1Ul+904kAVvkse0hfmmz48xH5+jPY
+PWVJfTgaEqh2eKqvaMfUT8zhALB+gFXLpjjmoyz7rGXImI34LgnGoLxiVfHcqLLUpZsZB58ZxGa
ZUG/0Wu8iOmT0AOr1RuV/AH8uluhNDxhk5CuhAL/BsJ3tZq+uvvgMwV7cCx1ybAf5ea2DOaZhx17
pa7oeGg+Xx6HOMUqmwuL4GhlivgA2+9hnXHNMQisR4sPAyHEs0BzRbkNmL4Uh2YyCufvyFMehD6A
+fviIy6KhDaokTiAt/HUSJRhEWxx6zYal5efbB2+kReKeV0uUcWwHvmmcvNPCVXJCbIZhyDQ/b4h
b2PJ+ESA+MMjR1mWAdTTs52RZwJgR4it/nGlwhNvpkclSISx0POFJIJbGa6s+lRU1uE/eBnkn4jk
vPyKHy3G+VyXng8vGr18H6cH77kx3FRANiCbIhq8khMBnk0oTvHD60boZSh+ynMiNaIfsHXvxQtk
cuq180rVV7b7dnLPJg7ERKdGsyZtpptT7vWDQSMGXBSYy2hdnhjRq/7X8AEBZaJ5g/61JFznO5Fg
8smSsmUvsijUiKnux2Bsb3aaigEqKkb1xmp0WoJ/70r6uItuc2ae2fTqJAuvqCq1z8gZU1/tTHE9
gxOPScg2e8pFruqTPGfvsqbTnnqQl4PeDs+G476AHrqhCW+FxBAc9gljFiFczISOTF/oVBUgfkSq
AI2QAIJgfBqSFWV6NziPQXKGoXT3X5fM0nSESeq99DurA7V3O40OHBOHquIGqFwWmzI21wZeM28A
mlXteVhSN81YaNuxNygVkRNLl1ev8N4mN4xH6/No3Mhxk673rzWuxooowpxjHpT5RFOdYo4v2Xal
7MlfXxe9TM/VBC8KnnAFKsLv8Oa7WayyCspf3cKuXmYAL0LNnOFHWIe8LumZiaDX7W4J0VC5m1yl
nwcUU9jEp7XSPDaPG/LYTvYb6ylCuEwsClPqKa4q/gvpDmrePB/2WZCxhCMd7WFqB1ajSpXBmUWO
HVq8qLMbyS+Q8nuNz3z7DFlEpgn0iE5SZkXbNPu0VuH1GNq+EV4wZsoO6RyHtd1T/VG0hDHH31fC
CnXxzeHHEq6lu/QAq9ngP6l94VD36hhscFsKXPQn8yXUz7BEkmFEtNxXmhBwG44dKA4GFjSWlqhi
Q4nDg7U02phWjZhTM323sIfw4RXVEdZQE149SwwZHpLduQyvHMgG3VfvRfY/SOH7bYJz8TTHSoLa
sISryFJuFRBOcApHigp8jFbiXjvMn+pXHF3ZNLXYrji1nVqYHSCemM8HThKF3YgOOE3WpsXWw9e+
DYhP6qsnyCNMnUXI4CBlEKSlGkBIt0h06XqOsO1Q+rEUhtBPOGI0QuTJ2s/vnvTHvE9yvmW74jlx
8Ycerzd4BDWfP9sc9iJLFTyYbmto6M3BYhKSLS5Z4YMLfP7pHzIwjpAnvWuhs9ZqJZ/VGMdHOmn2
c25+WkBHVmfKv5B8yXodielMfkc7IagdceA4yfdrFgEPOTFlAjnEXxEEa1ho19pd2MsFgvKyePh3
obWZ1UrThhqR9gU9xAysCCZYHA8Gug/fyhcQp96yUNt+IpkEMrQlrToZkcDIrT8xWgmY6zQOuHvW
Efq/NZlHYXTThr6HdCdKSy36/W35wW8A7YPWRVchiXyJywkeJqZLzQlyNLle0kA8dIuOhGPW6Ztj
sD5YwLyvu2bRoqViuXeQetFttES8ONNYQ4lWxjn8oserBaqkztdtMTUYgbktMDERys/KbydA8lUA
VGsMGJyK70/VZsLmx4aMWslj7MIReENHbnsm6Mfk3BvObPUMEiiqwvyWbpFeVeiT90wFy3fW0sYx
B9OQsbWnnRp1DVwbO/6qn1QDebKx31bRw+/QkQj15fUKqwrGCulF1iCg6zRHtbWyIkp+jDyIMX1t
2G+qcXTkD+HriXoZc41ufS44I9Gnmqtt9bdecaSbucladgKYuzqjCuEHEzGHAKxTFBNVQdGJQ6bo
SU34277Tyh2ECUNAPHIQANTl+F1mwC/VsHJvmmvMgZ7d//2xKNpsmP99Zygj+h8ex87o6deOSaiL
9ZCmyPL0LRpSQ491Q4Nt10WHIr+Wuo6yiNPsNYfWsfBb0L9llgArkoajC9OVpVTNf6wQ7A81kRoh
mVZexW8LD0cBF5wkj3UQAEfDenyPwpUZ/7J81bG476nk0GXYmM9HStBYkVE3HI+JJgDu98KW1bwr
4tWV7Ru0GjueFKYsF/UQj6bO6fYunfHu8aj+AeWbHUphe2pyxck+AfHEnfWsO0sKfsA78qfxsBHr
d19XKDh7xBSZNYTAKCtCa2AqFfk6j/LKwuot1Bnwe+Ese/XF8hNzDNUGx6t7wfk7xeg4CdXccTX0
SOOtLB7gf+HZQCjziSBP0+4FITyyBx1i+l5O15WMQI0q27QSa80n/WY7qgLVX0LOP5nMmCf4Erb+
J7C9KrV128MaiLGzqFshUIhTgBvYlwXTIMEC6DfMz+JdxTbc7kZWELJkR49sDBTNOVJWqkBdstuU
mOJ7qrQtZqoUvITO7pFhVc4Xv8roKTqUxLGjlVLvVcmihPzyUjA+y49Oj/0tr0u3HN5lCuwkxsX9
yce3ThVM20QgqRzlEtcdV/mDVk/mmM0R7rsTSFmYZNw8HhgUM8kdVMSe+wLQ+nJLsIjzvWu3JcrU
qnoQYT9QNEVgSoY4bPNp0Bd+MHGQjpR2W1diLuxfDHlI5PkphlH8YTNk7dIYQ+uFVnduFrnhFlNd
IpaEO5xjBmsMtHdE31T8AaZd7GqLSMDGt7SqEzvdjSMBG4yJwytku/O20Hgitzuc4FF0/AfErkrg
4oQjfo9FDm7B4T1Kj8B54odrwAweUkYt8OeWvF0cb4UCumIOuZemB+NlzCWpUMRwPvJIhuuR71B3
e8MbIyD0NLu2qTDk7ZpsyX73URG+9krgq7x0B7h/XmNt1cUKPvaFH3t/pjQ53UkuCrkAdMzRmcRM
BnOXcTLQrTBi+32t4ahm8msjg8Jzgi0Ab6Ko90bpNSQUudqNCOLE42I/5c/R4Gd8JM5WKBvcvxym
XF+Hbver1PqMnrkHHOaXALN01r/eh2vIjtnLMphIZFZ+O0waEdnmNNTUH6aOkbaMrHwyhirv8SfS
exT4Ocfm8M/aawc7ru6EpCSHIMwHvR1B2LYiF+AWN+pckZScVjVL2loMiBrRGgzuKhNnGoHakU9O
WFTqtqnlt5FKftc2d4B+cyjZ+lQk5sYpAByq9PpGjqjnmWaxedqpeRHqrEcfoh+eJGTjUYSo46MJ
Drkam+VYXQVMV0IyRDlPyP8G5gwvgciqtmUBwifx/hGIXJznmKyLXgIc5xCPktEqHQWPGlNbE1cB
+4iNhse3ZqnxcAG2XLkvfUNoISOofl1IQyLJoMBpBCYGTcZw/Kk7uo6aTf2nPdbwNlz+rsBKfvuU
2U9RLZUYCLZfOe+VYFx/+YA8uU0qaQhVmCcpXp/4bEHv1id+jePMtqfNHuj/A9CdHaN07io+VFEZ
Zim6lFqVFAt3kdpOl+aCGCcJq6vQft2EVqESCQrwGZeyjytE5BBzFvv9C40DVW21mVRBI89hSVST
CGQPzV8GGTQDQjkRTzAyy394QAH9lN30cfgyb2BQzK1+ZgXlpt3IFQru2ePaOWBbLFN8CfVPlsJL
maLNzzqRAXRx3GSOEyobUeTlupW8H/8Hh6Hl79dAcqw/0W/LZh2SGPs+OqZVOSDwcA1mHhAH2ay+
5l/N+bh9dKe0eWynksBWIvs8cACE4N4mhvEVdfylkGrl8u126mAm0IDuB4IUN8A7MDktCSCcA94o
Es/F4IhgLEkx16lg8gVBnJtQTGqpK3686XcgYgmrgMBkt+ahIkbyc3zAjF03EhGqYk6/9bm51MIn
102MkH5yq8mWwrSr2TcWVx49gc0T07BbczBQs2SmLwj74aTctX4wqNQT+aF14MWXbVrWyjYLk/fQ
98+tPRYix9/PFp9sPl+HZ/tMc0/AI6szqmAy2k25c260+hFiqJh9Le0V3G9bSO4qzlSx9op6KMxn
rHFbNcohQyzfsz+1wYDHeiP08CG21FJ7zNlfQ/PJuQZB/qcCiLkI/fYUqk70oILu+3BZik++WAk0
gtxPd3s4VKI4Ble2AlbdPKMT1NA205wstoliRlZ8SB14fNFQnd/ItD15LX1ennyBiX4asR9/K+hN
ew2N3H4cppSMYllv25KdNHH90YZ2XnB/VKrYQcx7iTjMkTQ24pPdMISkdaVEE1JYTeBe1ewPOUz3
lom492wIsqzmaYadGj2rrEwYerESehmvrYuoQa0BNr96VPXvu94w93E2MywX5wfe42wVyDxbfQLM
H48h1/V3DXNsuBrYpj1gAuAdjr+PiGskoBEHBARyCszGCsezg0Se2aIo5c01vaex7hvkSwuU3InD
9YpJYVcybB5Rk/Jj3R5lkgak5o/CDeGMuM0z5PgFYVgIAJWU+G9mOUwWDSW3e4chPmhqb7pQ2OD9
8rQfVqlaqhgOe8U21VjdjODZaE6loq7VTc/GN08hkFXmHIXzR5OxC+1auphdAm0O2NQSeWmOy2a1
PyGHRC2yMxvIRXFjp51frITjMecAa7Z5eg1TAjnM7lecRrCEBFe30hgYH2RO68HCmA+IyCcO4T3R
xF+veJusYkOR1eVgXU9NroxTnTsrKwSyZ65KA9a/lnfjSLiqh/zw0ZKHQvI+PiYbo3wHtm/HJqyJ
bSWAKv6jAxV4z66S2unRjiMOeuxkZIg6Vyw1cQVkRi5YQ0pyPTFO+0jYeSxSKyby9pS7X81pK4zt
xisu0douk4mkjMldz11aDucWuFsPl8wvgFVrN6fCxs/dSDRQ9cqUNSXcYce90qQwSDdCrPJhAY6g
rVMk4TYFud3JbyVCaGQHQHarSFDPWJAX0GwLW0ccT0E6qJnUocfdWqw6/AV9rvACxpbS57AvwO1o
AZoGzxqkSB2G+/8tTY9nORzu8M9WPovOjAWqQKYo5Qn0RIearfKT78DPe9704ZjAv8Kb/GDsELSS
ppFAxbG4qbL4oSUFEKmugjpTv00m5l9VzBT/afIoTmM+qRZGmbpP5xt6CqFqReBK0nlQqCgr/EX5
Ty5hlSZ8YkyQaTCH4iXOzM3+TuRUoYliiU5BCrOscMKA9JXCzDzOzAMvMMKWhgM5npF/KxoYeEm4
qCotFI+kCVO6u6EsMadoiXzASdVAv16ft5NNgAktYiw3JlEPplw37FM1paJqOBICidt8UyRq2OM5
CjOMHUuGW+wMLbvmg872/X7sSlBATYidrupkz2dTjEq+yyDcHGnMrd9tMZum8p98U89n5FLlZVvg
37xieFnOHEvqFQeaTMdpxn0e0FasdbSeSyV/5GEPPqfL1f4jHP4paITGWEjV3ED0VQOXZhsP1knI
ISGVs/ePyMZJD3E7Rqzp3HM0oeH9cyUbHPicoxu2hGnLCmA7mZOKJV63h09J/aUXcP+7JdZzBiAO
G14uQVIIvqEFdnFKRgTrdMOVMezIvLzMXoXlxBrg6R5IVmYatgeEdqO0zx3A7xGycQyQukIE85s5
0PNzZ7u/fJ28js7CssOY34wfAm0UNrZcnMDGD0KVoi5xztXyTgkVGyhkVl1z1BcHlTJFrmMUkWHx
utyvuleZdOc20+0cY+CQmKptv8ZYdP7z8PKHbr/H9UcPHTTAeWuN5cRukO2KK1rdj1cs2hUJKYRY
WCrTND2n7ecgplDxYGIVM2xbx7+J8szqxov1w+P8jmF4egRCkV7bSLwVPpbPubyI3Yfx5ScbFE+O
nSsjtp9OgKTJ1Xjon1Aen0jrBZJHmzbLok4N1kEEr4BFekOMzqb4bYboi/63e6FHj1cTEQAv/fqa
zxBvzZRoYU2IuKQpJ8zeyWLm4ulGTBDGAAnyRdnowiyXQQh57Vvm/e6g2mcHFDlOS2lAFuBPHlTV
TUFMnaDofxJi3BOTIZVr8QH9N58Vd2kEh+wD/Z3w8Wy4hJpYcndjd7OihJhB/kNtsDEXQrVZqbL7
DrQUMuGPwpvp61qSHZxWvaM1MG3apFSUt/9YIkHQDAqld/tk3hTE6KQvabmVZfE+Vnag4F3nw7wF
EwYqvL7yA/L8tWHyHKe6k7eN6H954266GQmv4gAtjXH/Dmrn4HsgbMucSPHyL1DTo68xTpcZKKkc
HDFAoqem0+0bsNc6L9btyvLCHH66x+7oer8yHHVE54qNMdBDNVD48GDwcsiReimXDg4gQg5ZM2UG
mB6nRU7db6M4Brs90TmkBAgIftryDBjnRFXJaT2wLmQbXtOYQRUA4iVt9BxIMl8YldDQn/S1vB3G
nkElIyQANwr0rdlqgVTHjJmD4dVoDLJE3nUj0G4fVEVf7UOvnSSg20PWn07BI/faZU+p6v8ab3Ta
630DRuZIHP4iC8pGAQFtvkKVjPLDUO68G9wl+aHmEgjUQR0c3zuagIcsfzoM09hSRResyE9uh8Kq
AmV/XrMB6RagUV56DyEjffEh4HwMUum9lIbkV7uYySakOlhvNmTsRyZcNZHjwhkEa0/kbbHtI13c
r0xrYAW9CfAUSLF7to1vrKssREUS7hySwcPcgIR8ZY5HolMujjAMFLd1It5akNJ5maleilHJf7G8
AQdg5xnPD+eHGmsprZ7Nf5KwLk9GlN/oT444u2hrkaIAa+7Za3wjvihuYob4JDzmIaui/d+x5M41
+EzRdMkr+2vSXVOqUhXZOGWYo7aTCnuh+/r8WLlOjxp6Eab7m9Zyzm7WCHqDQgjkD/LY0m1tF+sW
UmECQ7k5CtIajkcVDBYwOejKk1PSVQxQYDZR2egnpnmlXD62bLtAEE9T7ZMuZxVKLRAhY3dusMmE
M/u0kIZNNlEJTK4nQZS8LhQz50G/omDO6uvl4CUXX7RtU9aNUl8ttYYZv0UEbA8OEhFkzztjdOap
WnSFQ3pLpbzRIFlXaFQ6cC79+LvJr8Ipfdym6DcOf/yI2f/zf7AnVIxTITuhbIdU8yo5IuFhhiJ4
Zv8SC7umLD6Lb7fSE0mV2FiSTLdqREU99cPTcaLaIlnnvXuff4A1yaN2zfmtXzFLMNgHQvtqf2Lz
A6FYrWxjX/ydpg2vuAeOaFqNdnzBSmEpj3yx2c2XL6KAM1MkvhtMmg94cIkW/D4WzS5aN8z8heTM
KN6fHpJ4Fi6O5iGab8QHO6tiEP206zA0Ov9GEcnrinPWpfyUpfDXRW8Hum1i2cQtRFy8O6zGq7mk
4Pj3zPu7yb1TKeH+O9lhOm5NV47Lc/ywjZjqryp2x6Gx7BW2xdxRmUhbpKKtoTGxmzn1nB/1kiZt
5DgUsBheOxa0ovu7y6iVgbh4NNp5WAsN9N2siqqqCUkc2EH2ja8vScoB+wzCGdsynQLFsoYf0S3O
5+NkLvfQKvcqw+aQJ/8LMGPzBroH6BRc/I4Tz/rW63n9xXHk/rlExM56fm8BQA3OXl3j/N//MviA
Y6SoW8JOSXCdC3+d1ZnUAmMYVtaCLPw4OREaGGNueC2CLIaeRmFvNe1MA6uGBkd0tX0R7oaYTt0g
F09Rbtdk851PHy1qakmvGT8L+cSb6jU2Aj14ZOMtfQFALTkd4LIwPTEGhhzvrpyvH8WNDVGP5MqG
qUgttKZxImLXCPdNK3Wg/Qj7f9RhHKyq5PkrAi5DcKLY5kbp57gFxngA9gfNpRWYz8UiyzwLJqZ7
Xn/5Dfn74ZrKjvSIFdfwboI0sB1dAs4WaSaLdYmH3/xsYuZQg5h8yiYngm5LHID6SfwVxQaAUumw
YpJ8O4Vja9HcNfvBN9ppelcblLWroSVKpygMNuUnu0RBE8ZnzkFwItG8id9EPDlX+OOUzvybNarg
uZvcfNymtwWV136aUsrwpRbJyPK/x78hIFOiDZ0slqGvLHuLgj9aywghu0l7h7juIO8RnwoFmsar
KufELQtrqOOzhzoBvviItQVrxurHiLCiIJdOd8uqvlJlyZ2HAgyyMbTpB/PewMV16yY3B+9EkjsZ
rCA6SM9Te7BEJf70i6BvKbRfqTy/Qy3rphbtkvkf7vN9EuFR1F+/qvu0GSQPPCT5z50QrYnWmb59
kIjBZouhm0lv/UJ5VjlxPSqpiEiJRTYElO3yc8QUmUYkRXV3W1Ha4kYAxdhjMgWHjqUnIU36e35T
1vlYTU4lVGFDgXi4tbfJcuGoz6GM+7DxWlhVUV9x8uTJAZi2YkNOV4RFtrSAcx1xa8ugIKoCYe2h
ZzhExY3ktaMgOHYKqOZdOZV4FVGVKe3NBtIk78ZIiefCBLxFI4RluM5O1FUjZMOZ4v/Dy6wUVDOk
bbXc0RHNJ4RI35LkkYM2p7mhVKOzNu+bVTVBOAg7scR8rnUY6He6gO1kVy9JKBve3cd8XEJCEHMb
8JlAc1RBoz/MNVPDs9rxzUbTmDLKW1TfYj0fgJ2XUh4LCIwzuyVTw2lpI6z/NSAwIovvEnQqvsfv
LzrtGJ+A3LY1fvj2o2yFp4A0InUQzJ5dIzHWU8kQO9VlJ82F49GZ98MCBgRNkSy3QelvwU+Wr4rx
NxuHcepje10su7eHHW2puoRp4HKq7D4R1HJbmjSMSJfy9OK4L+Tt/My8Rnx8V/2NtBBg0ZY4kfhD
alHGn1fglYbRyXnD45B7p/UL1jyKlmDNfjV2SY/Sffh9j5FuIfuV6zG47pkD/aphAyrp2B/XR7iH
/7XXFig+UNSPDP/WWmsqNXl1YqycQtJw2E3/L07NinbIkwS8l4ffchU32mdPwbvXeFXw/lFYH0dC
GkE1soks4eKM1PHzxv4LYT7X+JD/XccS05BaAYzNtqgDIjr7M0rUNWXodhAq3hnm06Fk3XZk780W
AduFp3hM94a30ifNeTKWScEC6CyvBNFTWPHMfymmd5pEl4HtjScsK+DD6dVqfdzat4B9DXncZUqM
7lbaqrw832Kru+hXoFMnkHWi6esDU0a/+JMf4FbwdA0zhQo3Z5H7S3Ex55MZ8CHFPhwc1Sm1PDiA
AuyYy6tR3fbQDs9BS+ZyReUFKRvVp6SMGNfon4WPGCqmOsY8VivxU2QqxSOk851Cj3qyAzsu8jN+
WHmi+WnD1/s3epS9jjWK9IoXAjXbvi0lyon2cnAFqpFCKSgDSzGvYPoVXH8vcJUR1Va4qBKfbmOR
q5th+0Cknob9KVIGMzArDtdyIrNKwMyqLzXyadahQEZfA5uhFL3WKw99DcFzhTh91a4sXRXsVeiw
6feKRWgyxfW3Ds3xtmT+/lVuA9/38uu+QKoTbdTwyxHXxusSH2Gq+QjIdL2vqvfoDMiwgD/LsKtk
g9x6JH8Nq3aD3ya2RXH0rT+Rnrb4nfi9oCiRlHGGa+NkiEd6lrtbf/17q8nZOs+NOpVRNNBaCQN2
sc+TT86exZEcdyj9tcYmAEFNH59qrmd+GaxxQHCb0qd5bKBtd8yTNwjbDIIpnHCTleU7Dgt2dgX+
OqK+6K2BGm+CVtAOhBk0u9koUUMgoF7nrA8ALy+ABrLKhoYGWq6Po3dV2IJqI9mfoFmUnXBgFqWw
6FalvrhwW7pQZtzFuMiOwvsEHuf7vM6nWPT82ns5144sZ851wOMIqR1mOREgwniYbPBmJwa9cTLJ
khfrKW1Lgwo8IFBkhxD6OEKo+7f3LtJhGwO6KT59xGA32gW+arFqV1SLUGSyNAb/cOr5gfvUb3fB
YbFy17Ad/gezMiwTtjPKSQC022fN8nrHfVCHAY8EyblqyQl4//j3eJIevvy9/jA3A8SDR2T8R+e8
5lwIK5t7jSjLPKsbro58mKLOSs3r6AFKa1j9XQ6xee04cWXTAMBbGmKIftdb4uhUWsAVSuVLXKhO
F0hwc15svYd1PMCWbXIzKQafzxBJtu/Xf/GO8YGk+hcLYDim6p8l4pY8O37vmmqrYvB0Xyh6kg1g
THoJlj4CH03HP7duRUzhuXMzEerYb622wbO+kGTQjilYm8PHajF4paJ+PnHiHW7X436aYk3s3C2d
hhi0c0Rg2jadC+ZdWc0Ke7QxCZkSMRj2QEgo9DGJVRzoPrntQG8a6dWPz10S3ndPWWQyMknEa5E1
o9v22KQGJKmv5VWI94R0s/CXa6grLrVvYJs8+cJJK+3doaRe0sfROBhp+Xbq/4TPNJzbf2SHYDqq
4CUSJp+K12sxWVwMBZhrk8Y3dMpmRiypbzPw//xKFzsJHYkAjJFPQ7PWudRCRv89rPKgX5EXXiLe
blgkivOBVVBOCuyCt+zurUuUslPGv17g2ofoBHi6bXjqPO4G1cAueb7lhh6oK3D5Q3WrbfY4NDAN
mGvJD6Cg57H+/HCkCBGP+ztKDrfQ6tyYfRpn3gP+NMLccqsLCvNand2lz436Z62lts7rjRmlXdjf
U5xwsLakk0lN81TN9IXIi/jDgEbppTwI1to/FCoOsxI6HEpkk7YP621W6+VUQO1SmgvpElM4+KI0
tb6BW5LfK3bc217WmmV3D72VTetbftVCuvgjh+nXJdEwV7LUh2YCx2lTUIB11l9/ytviJvgzzbDA
kBhGcR7pf1DegN6PspAx70K2xebpFP/s9418vYJIgE904NolUIzXbE1b6Evq0khnJyZ9SQsukRYW
66oyc9CSKLb+Z/doVKHqw1/pAutv0FT8qWEdprP8buE3ebcoclNOiiXGh1hFaEn95c7S+JVnR46f
tQ22DegbjZF0RbaXaaSvq/EKdsU4iKTnUE2anPaCd8J18GhFhBaeTj/37ha8/ew1/wVnZEoKRiM+
YCTC8eG/oXWaueUnJBiZzwNoN5GVQ94aga5qx18XjSMsqYlWjwTS5NqxShltmdz9Bhqg4shryfyd
zAiCplT6e4Rm9qSeBjWuWCX5mLDwGcn3wBuW4/g3IMXtA2TOcnI5vJjLOeVAlYoQKmkexoZNldfR
PDDCnJEnhHfKhkvf9yfGCkCjoX9fCD9p8+747D/G/uTgPITU7HbAObJpbRXBtsGpeCyYSCIOnYLu
cl7bMla2lTFO1EycpStuAa0hr9H7A+BOJy6d6esgjZ5+Be1ALj1j+hAQ9hqT4YjqbmFMATcE0Sq0
RZBuCXwArf6E+IjMn9yi0lggFUfdL2D/YO2SzkrApa89YfaYARgUlSGktxF6QZF4GyKx7juLTxbk
CFu2FeH1SQkmUAspMwdTCALPJkuBMuhudScR6V9NT15kD0MEaISkVV0pnjBTY4Clb03X7Q1StDWH
d/ZeZmq5nmrCEXoTP295CW3/6P0hXl79wAI8l1UYO9dYVs3XlX18XxkZadC0ntmBxvb/DImqyXWK
yaS1TudzeAjXVkg6UhaSxYkLe87OEkBy/G+I7P7WxWGP4JVnqiut//XlnEkpdrO8j97EWyCb5Wh3
XN030PSHaCVyhzVnxojlXaqZHtPknJtkJfCDJFUtVk6j+jxmcUZwNolL3LqbB5d5oNXcE6FXJTnW
5tThZ2BbYsGgJn7KNKroq+zCQxTPV6quMsmk2KY7hxqOoCyT7NTWU4yMQ+xNmHzNBX73kkVXeH39
BXoJ+x6oUHo82LafED77unboSM9saDGUmAX02tkvQylHfUYLmZFi2lxxS0DORPpCDFVem2TfcWsB
ve8BP85SVg68mjgmAvUnpliliS9G9qcm1X7ud6zme4BFpjniZQtyYIFtjiAkh8wBUkD5Wf2dX8zv
a8jZZlXyXjAwPuUwDtAADZhAy+5ft32J/PnKRF1Vv413CPoKprXZhPrxBiGa/TlaKQfHDZRANkYi
u6lCsQhk6em8Ea7hGvOmRj/6n1cCZdLx4I/W/vSZOc1ADqwWAFwRUay62FtAext7tIMSg83x1WQL
dA+RhZLXnAAP1pxWlmNQ+czQEbU660JeSTaCdvh0UvObZSl9af0uh4YVK33xek/VhgescblcqCGT
c8B+UPcJdGylsVDVFB1zDVDf8QMc2aUU+LJVI0QKBLOeakj7yMdOwOb/DgAZ3Sm/5Kp9qz8rDqMO
8CxIP0GvtRZWm+inbRXUAm3Mo3qpVvSOOQEwgl0wu7p6rcrAT+yJuSvOl+fyEMrlG0Mm54AcCHHZ
G+SAt7Dgv4WriWCt5eAv1ESStOVJoqhKONgk1bres0GVA7U6NCm2hdsU7sOfi4G0/09J35Qa4Z1G
XWMuxqxICjiNNQjJECjCWAWvVTi0Bs9SiTmZVHMmBvY4v/l00ixXgAndz79edqrQBK6wcWB1VV2h
YgiWiL0DZ9vWXAZMq9pIVnx4F7l67L+U31G2zoY0qknh2b9+TxrDwVzvKLvAuH7mp9M3lS20t7qI
Y47NQ9UJ4nlFVV4Ex0UuekVGB0Tmeoko8oOil5PHRll99BmY+W3KIVBMDRviGpVkBLuePmpYm/TI
Lu3IyajilhuwSzLwJB4DvgHYRtqqZ/3kPTiHpNXMqmeKEx40TQRY9i8/J+AeP0XMGSEjW08fvTKR
/3jQ7n2jHl7i2JYuweaYtPfVDH1goON/HsHxDNpYqJ2XDJTEcCdGT/bKkAibVU/kb7RdPYbsZOqU
YhQZNxHrdFXj8bhGd9LYUXfoa73r+UObvT63ClAm/A5PbkGkExhI0vc6tlNK0ziZig5XAVHoGXPS
qTBEm23TYqemtW1GFASFKSPsfCo+kOsShBrieTh7+Numdmuuxy30nDxxXogks7Xr8h1vsWEL18us
eVVI76k+tYJ0XcekHAT9lATs3PimNqq6I8efQNmdV4i9tqGXgJuRC7WSSxTEDdspTaHiMF7bPhXd
3RnQbnOai33lkV5yZGK16j6Rl/Jk+4FsWhgS9Tdaa9p/yJvT4+lqcG7s7oATdFgc7QCGd44ZNbif
AZ9Su5lKYDFBtul3Mdckl97R95JtPyUvcU3eZ3JyjhVfiTuVFcLwq4wtDYSiDVrm4rvgbuERw/3U
7EwMKqUYnisAx9sZsysQS2CAP2aTKbP+q+s56NufWIr4KL0c2WJVSTmrMQJXm36cJqAhkrsUw27A
7t3Ra/SgIRHMugn+agybHDBI+1xx/1z16kzpjwHUc5dbVOUqUrvfp/uhqhJXDPwwS1TyLWTJhI9j
vJH99gYLHGfvgkSuG1pYRxibVcOoNHGvpnTvk9cuBoKMjTJOC80YQOIacHn+w8w1Dq+3dlJb2IjC
3+PdqTNJ7aUbiY7x1IfExR43TypdIYdiGDW3Xmq70xAwZmCZdRaj1+y3C+I2j58KUZ9t6vjXNvqZ
/nklKfsJ3H9tKMXjoSdTjmCJL6GxQ5Yg8Au0jGTqSLgdm4Bktm3dJqVUNalcUVxFlcZCn6dxPbA8
TpSCYCrnMt4Y2E3/Z+DrdjyIzMKsC9Itm/nXHnscy6F+BR95nLmN+tB/0oHyYtn8nu4YIHEWxZGr
8pY9iDwfx4dakIKJjtI7pPv6W2Gz9W9gSn0IwnPb254oGa+OZ93Q0WBnAu6/ObFJorzPLaKKyZK+
bZKkGPefYgytIkaRI8th/9CJHSxw2Non1KPqccAwI0QbdyqjQVLsIOLdE5NiOQq4TACdWMLrp0yf
h5AYxQ58aL2cgDYqf3ZT9cVvD0bE9NmBEe4aVL/JZFOLssY+4BXqR/4V5n8Uo40rtV4HGClrE9r8
qBlVjaoL0DEre8+Fec76jsFXu4EreC/a86/uoopq21oCWSi2ny28bjE50vFBNgmPYS1KShIihUfV
MnF/kWA9u98JI/RrBf8Y4SH2vwsR2QSv9oKIBb2OoS+ZQ0+z9Dx90eDcIGQHCwxc3wkEJy1zUAKF
Ecuhm4HXPmJOMwkSnCFzOw2ltG1/wIYP2D72Gf904nmw1l5HHq7J+bXjgv71+BF+sKzYtxyNZfRm
LmxYp9YjUwosvFEXgKeizAv2zri/v0iua7PQ4iqrduy7YwLsBCPfvaj/h0Qfv5eEn3SB/uGIx5WU
xKGm9RGazvDDUhTofA47lV+KZxnANA98f8TjLXGROzDOmt0SBAAoQRn5A7bMn3wZs556ReMhK4o5
tFEjpc+3QhrTkMgDAY8YwgqKdrxF/IwPt5Z4WRYcJ4oHu3eKKwLqk+KsfmewwDQzIRSH2aO9jaEc
9jalcihx3xM6Z3AiiRp51ejG3e/Lo52bbB+aFhhPJP8Bsl8oRP1M0dAKmpFoe3IeWL9yrdAGLYHf
b7v3HvD6oMhoUJtz7u0y+zpvW5TLcySE8OuWmKGNqRcBuDz490a6v/KeTnzPZsEK7HEe5o0o5Bj+
wKLh3sYmv4t5mXzTllQRGb8H3v+sy5G7rtksze+rukZkfHale6j66cKHteNaC/7CiRxoffVkuk9n
l6r1Jk4zDUgz6Qcey3Ttn4kMQ+9lpuIn7NUF83m0foAysdAxDNsZ7p9tIQO0/cW4n34B/IMOAbor
QmMCX1my6IuUZWHY9yGShiyNmr5orAfemL9X3RQMoYDFUPLsarN5YxaKm9poHihsbn9eIjsKwSr5
DvWVYa4D7kSzwZgkYcTalQCnzvP4TiJQtG49v+Sl5CbwXIzvdUW60aHHYd/xuHZe1pcxX+VRgGLZ
wdo2ilF/ZI54ZmOR7CraFxM1JBhAlHketDUTTYhDV2bzC0fpaLG5ygDJlHRBaCpJ+Fd4B9WQNTaR
tBgg9exz6mlUURyKd+0V3S2cwLNpyeMyoDb8R4Zw819cSgqusuDTqwKfOXGcb0gq5T+3GoF3o2bf
gc1t/Oz50/iPUrtWvNz8b77u75uGfJsH2oMCM+P9mvT53PDb6sRmmRV5eVM+2seM2aAtrm/Rr1do
jHyB7q7jxzMysbd7sq7ppfMy4Dk5lRXrbhhfKMaDRt8RcSrXsKApQF/qjrRjetUOqEjXmy20O1YP
Rj5UQvhOOmCeZSALqrnn5OzpPoWVh4LgyW6PFtQ1zzCiiy+KoY0Fo/0TkyzVGTPIS47stwuO8/22
XkJZDsCSTzOfyAxl2ap1r6rZsMnbrAZ/2jQpvr66xPPlt5GuFsvg84cELeWMHVZyNW6oJvoTovVi
Fcuxn8UxRfvD5Vw97tlVA1wkLEA+7+Q8Z3+irj2R3y7U/DrSmHRBO5zxiohYoqEb1x6trzjdaUiS
OBsbVgp588z/tNjS7fAif8snav76BsZ70NQPrubBofgg/wCWyu6I0s763WWT0t8oM09Uczugja5U
xmZGxUPbcESQpbGwSJaZ2ndw7kbLRfLV1Lzo8IqP+KRd4kDidHIfjD83TfoRYNWev5zoQuzDUYDg
L2EOKfT2lxJOQH0OB4cYs9/ZftvWtpfmpLMDO36QatAQB9Rm57wyjgr/qfLNWEQ3WDE21kt9/Pw1
pFsTdyRV7GftyH07L26JgUDvJdMxKxd6/i6I8/FmdDhmIsTDVUalaRVOVpKUsGqHsjWBqZ0t3oYl
fKRCkbVpEFiNEje8s70qEMy+nDshSzNoz8wH9SQeNZwhh1NCJCrFqr4oF/ZZPMD3v6CO2840MmLo
714qj6351IsigUvvr818Qk3mfQimjusSN/PBwojje8xhocq/QIj4MOEJjH0pTgLsmc54gCVT/e6f
ALZ+mPSv+/JMGKmd9zuIIJeQUzL3gDOjX8fqTZokwew7LtelufmuyuVkk0RZnHGBcmp6v+tVVjGT
ulPN0Y2VG6DqTb6OMebac2kgx2kJxltQURg886cS7nEG36tneJvaIoFyzZxULYLMaY7NJrxVfV0/
aVj7+HvGoyPF5XOTbee4wYcLQrQeInWygaLUHQqGjQmdrCfDYznRv+xUIAiuA/lI/oAWEjAh+QfE
SSQERmJ5OwQmNmWru6s0rwCE602yRSlRuVkxUCQHEWIod/vfjxL8ElXYA+kwafHD37dVf4MY52CY
wJrUj7LcPIwnPEfjV+bPQUp0JNMopibeY///HviZVLuzJLkVMsCXMLJZwa7KYRjfdmicTOs/bgP5
sWbrrijVcpQbSlNw2sO8UIik3KqcWpczTvAamUVlUD9DJOPisRfH7t/AbaUWnvBlvI+uPDe7MsCv
uaTral9+jytoelp6haYhhA0VvDMSjOuDLj0auvCU/V3avfKQSbwktsinl7BlJ+Vf6Crv+BgsvR7I
Q1X4yP7VxmoYxsM8v69waAMHIWiQ5QmMwB0H6hNJWvPM9Us/K0n4FYxop/kZmafPumHN5AVbylk0
q6IX4jcjX9Cs/eCePK1aMU0eWOBsk2ZQYsIKXUz0lIpO/4or01+RBumlg9ZHbpHspDKyoHNHW2K8
F/JpeiiprVJ97KYVR9u5XUFVRXXDOvsFs3V3wAosUQYg457GWhXdFKAkvEabRVrsiDekaJYcG0hh
8oqt9jpzyGGXT+J8S1t1Ii72zLPpdw9LPHBgwzeJaWyRZcH92RUNEt8k7y0vmwKVqp8QRpfbTiv6
qvapyHISiIhhl8Dp/Sh/uYt66l2iGoZJqb3Xho2spTalADnydwJ8lUFNOELwMtOkP5cMKa+Bki05
qTNDDPcbGAIQhK/m2BTvDXVfMXtUQLzYRbofJ7S6PSsEkFE9S8WUPcBjE6UHaE00lNRBxNHXJSAQ
6W2L4HsyiBMKUiG7NUge09oxWUmnysWTkt8XA2iA6lQyaR1VthNGYy6IgHFaPshpw4AeDn2ICjsB
69ipLJ9lcd9LXw3f6Y7a0cmJSoEgOnkK2tkLY3BEihvXKAaneIrxdYKdMDdAflSSQt8Ld3vqY5dY
nF+3qi4PFEVVAr3ZaJYveK3z2dE6f+3Mnj2KdMS9nok2dHV5qSY2jb/7PeXMnYXBN9pCU208hxd5
YOdcySM8t/15CCkZ1EQWbuzRkxkn4USPy6lT1PlFckOSKxosigOMRFUuh8EGNYnHzFSYwiEWgJtr
/WcJ6RGQqQyPL7DhObumQRn23NaRJbZUpa0HaowfMp41h5P/8i6cox2xH2ATU9SfcLXHozp6UF/N
CJ9CrVpB2C0YTYiOYHuuq5MTJVmYCaz59+z70GSWZgTkJdsWdOvkPIRPBJo7MOIxMoWhRpyPzZ0H
ID82B7ZHt4Gw//DuG/3PR2FjYGbSDKfJlrAldr3cqerEsvMfyyVKyFyActC/kN3xUvZyyipkvtNN
sSm2VBHF3asvUzDFZ38e5M7J8Y6x6ckkf97zllyUTGKX43EWmTCpdXHaK/8CzRPN6qI1Kes1CvQO
F+kwY9/rjLILaV3vAoTOOPOo2inqwSMgmrdgDdHKeV/MGjSDg1u9U7HZ91Eq7dcFhXPeTm9To2Qh
HpkMYL26KSEE+GiiKRf4qRo4W3M82SYk8SRuzPZdC0AvyQ131/eGLOsIklvgYLtVXGoaTWvGkPdX
2oAhinkYzGOfj8fkqS+rRes0+hELZjA/gKDFIOJld3n+wU4AVuT6Aq6evs4AZbyYhDexIuo+93Aa
vzD3kPVeAsUEZlXzhODrkseMrr2BtP1jNoHFEbxD8PXBoUWTKLzdfeQgsC1s2wH5+9tEi0KzGo2V
1Yf30QBekoVkxdKqIscUmb898yXfXZ/OOB4mzC1r5YkDFIf7GveG/RJB6dsm24Q6i8fiBOJS8Ssm
e0Ja2nxpn39DVDOtVOYvZs0bIpbVtR2rXAo0H7cNyPPueBgZA858slderO/+8POYuEEEQxLAs1m9
6iFZHHOUywYh0npbJeIJMMMSakeSxHzEERQ6Tzjl4aTO2Ds5BI6MVXrHR09GptMRlp4uTcr82XP/
WcELIN6vuqsaoGAxwCxV01erHWenNkneZ2dfCBp/4GFAXuupsTj1OrBJAdDEBb7jfuHVl9kku3FK
BiUxKxGa4MUzDNeOGXh8Anvl5ciMghRz06ff2jTm8i9kcnckvjALjI/z3f4x9cylKYU3w6XUkKeO
VslT/UI7SlDotm9iN73X5UkEi6edm0C2ZWZTbwujVRZNYowZir61d4W3UDV7VsTS00fiI/1V8l4j
qCpg+cc72qjgnOmzSHdK2oL47XwYsAqh+Dqsu3o7Q9Za6rxnKyV9bRERPFga/llDPjVOUOkpJIka
W/qLwC+LfIetA4Q6V2u+c0doAYUqOVWBOgZxs2wH1wCmpfpnW8iXeTKNfwO0z01taYK5/I2ZTb9+
ckZBETiCmMqsJBzNLCvw8KpNA1O1ilGTiBDFN4T0namKyUVAvAHz0HL1dTvjlL/CR0Vh78y2U8IR
h8J4ab/OgPuLDXdCSXBkhRWI1yUtHsFtQRPDxr7neT5LT1RlSUJMvmseEGhnOrerEnWs/kvKa1dr
irjExRgIMNwql/XZLO5asokfTBOOyBFpnYuxmTIY+ADJ95TUWLjLW8F90smDjIBvAm7qrkxzat6E
ZeF6Ac/Knl9xPAeuc7dHWD2b6wIM8AfWdFQfkuYErbfNeHUhYAcKa9TSQy+bSMAxej4mOBKfF0uN
FYfmcrc/k9Uix3amtCVm2sPhSbIUQvu3rLTIWRskB45his2eLidc4Fm51UnYDyqbi4FvXZN8z/kf
9qlBZcgR7OWpA99NeJKzEziiAXuEJhFBJUZtR6pU9jk2sjQX50C/kj6UiBEAq1/ktv5nYxmS2PAF
Wj/ErUF016HcBAOXmy17GiCQ3ZwoLMds+YTNxl92rdOhae3rQEvsdSa4wYUZ/6s7nhOqWJUevQgo
PFlW4b9IUMtAU5S9JZH/MpiUYSTLuJry4O46HozzW5c4JEXO7RgbxVl2GarC7FBD4DYuC5ISVgaS
9oT5SNYXlGVtqB5+h8vA3olEzp+nXS35TftF4Xf7FBMNuDwBE/NXThr4Ciuv/Fk5B6KBENgaf5ix
s2gcvYa8u1Aq1id0522lLZMTGafpUgI06JVgUjlYC8N5R1K6AM4WvugGpNXnCChc4ieuwhqL53WF
LEZqUb591UWH78iJ9be7X0Uzscjwv286XHtE1EuIu1YoK/cogRnxhf+F79thEVc8gTp8L28jdlQJ
4euHzABX1yUrCJj/UwsObIZ9qxPkzXigqaLPpn9zuLgLRGHCi5otuqfki+NBzL8DG9NY/rjD2KtA
0OUr+oCTakGr5zWbuSDNViJMabDkDF8XZNkV6ox3WgX0AcTfUgGfz6yCp1hAR0Uqxhzr2uoIdv1e
KhG+nv//dcHggZqj155/RETC58M18fzbtmuZ40R9e1HO64EuznR2EL9MX5sBNYEx/AQREdPiKMMp
83BustRXZiBvIMWflZoJCy+kA8m48zKuqoleqTRzPPb7F6uf/Arqcb3RyMrXfOhiIW3A5hOC6al8
Kj77GkmLXH5Wtl0or7f10f6Tjpbv9geh37X8Mo+AMFHhKZ7dFs+KjVSHZRTKK4P0KWo0fhp9TYQz
26fLFKQI7W+eJtoCDuUxZWWePb02QS/Inlo47fuzAOrykDpI4hEE0hY7NruONzWLsyau6dzMP30H
YfQ9Zl8YneqDSY7Oy/2r0SacoSrvFZFaUMZ1sDpO0y6mullrNWbApaGIt4NM1S9eGT/89A52Vlx9
xNctnkQXitcbGb43ETSrPlOuMagQfxPB7g0EfBe3xnnVpO/x5iUrXEBiLBqUJiJBO3hKX84LD/Fg
0JdHLoteRw2ornu2voOQ8pm/HlToE5jnebzkvnFg+Xes553dOBAzVjpzwqGNBH1s5Y1B9ssY32Js
mqdlUP9WjSh7QLfs5t0xK5tUfN4uKjVlDp4UnyNlGZRyeQQMqJSCZdi1CGUY81TZsvfvktA9i0HC
9PbNdg0/dE837pNUkep90cVqgVRSCvYKuTQioGvhE0IsFMU9uhyD7v9sm4HpOxvO05UqRLWRAsy0
71inWBO9blBxplMYAr5WY3mHav4pHwmxeOaLsZwQRI8gjWG0UAh2M40/Wd0J+538z1sCxZhgDkWf
A/vatqWBZym0dXi45nIMZE+kY8KxAX+UOrroZFUi9xj05nLcpZhbPe6dcXwoaBJTt0FSlWjwBnb9
mFm9lsAW3meEkrmVjt+R/3i4P8OjZuCIBKTfT41We3F3Dii70G/MSTT2nvcNby1/24kV6oDtHl4m
dezlVzKSZeXV1QCHXpW8fkz16VD/L5KkJTL69u1kP79x5dMJ+49u0vTvTgop5Op6VlPSky5wTcbQ
lx+UJQp/q+GqW7UYavuCYQEmFrl7LOVkC+CILjd/g72Ukg3xJKgtcWhGhnthjdohc8G4Lq+FFG9W
5ZquWWBlOVJdqBi6rOvPjZGQ0OnFVoLZJbNtHcU58A+GEWPYAlXLqaT9JQo7rxtdGo3fuVYm+NQn
Jtd3LYdT4YBtaXcaYLeFedS9ZA+znD0JywCjiZZEdiyy0zIRWv8BWO+VqfYia7BrfGbL5J6Spkir
jyMI1VxZr9TrpJIN7BpsDX3XldiLzAQiUi2Hsn/sWDT1prVvqifTza20dtX+FQJS8ekaGM5p2168
peMlWGAMJgNCbAX7vdkJ/0ln8fsWJAV8W/iUKv68zhhCtdkAwnMLDYsgkJ0uULF9Y3WVWHQu7M4h
j0qyLSGp1QKkFpqAOvDbvnG9zFIM0Od32vJjgULeJF0b+gkiUqqHAQ0ceh2+xujH4NFguaYcU6PW
9E1d5FR4cWr6IjBKsj1W+KEkuFhQT6JdsbBB5DBTe5RKlGlPGNzutaSKhNyjVoW2d97uYHdpKoZy
v/sHfx7xh34tBEl8Mg3untL+JimixQZOZdYCxRpwOCII03odlKfdBqQiLOKyxHfQ/OZIk4k2DAbz
K3QgFVkxr3CuFZCVZoKyqkfEioj234qn3oOVH0Mli8dyY24+f2GO7nEy1WcGIVbI6oVEdN5wmksp
52OoXcz/IigbL6Cl59pck1MUCPSUjU2gA422IeKI0jOEsJKJk2yZPWPc1cFwQUptsP2iEMmsysEG
Yu6fBaqI9ruKv1dd26Q1TisaS5vojabHVYWTo2Kt9/u/gnRrTqrKSEIXYD6DOWSoxq002SSDkJps
eBG5T/dJe6FVfJm/jEwGszG4hfji3TrJrLTFkYYD1On6q7x9K3D0glrtxUra1QMwJ64ltlunvfq+
4YuwzLXaXSPXS5VWfTN0gg3ueCp80k6/tKsR7GGJH1vdh61AOjO8Y8WXYoRNfrV9N5jqy1tFBpC6
NXLznNa09C5lsitJAQsZZfpGlFdD2iqwyq0ShfPkRE4erJzaLnzr8fq4MiPpRBBEHa29oEfa333O
ucO2SWrxqDbnFILaQ8wdzvRqVyvOETDCyNTB9aIiMtVRbiofajGT3T0GrUfNYqR5ySU3J4WRdUoF
lRR7RyOHdqEnocLG3lF/3dzpmTtvVNPZy62vKKZ1r27c+LyW5vt7cGb2X88Ek4yQ6uXuPyn/8TJo
iIiKw7GOw9p3AGuqqvoilpqx+65I0S1ulcqT9ysmUTSuyLsQ9tYKHL+UZN/9Uh2iPX7dDZS+9s0C
IIjlkBh7/MC1Sd2JivazJa7LLC+i/dyzL3ogc8KXsEHkWXw7IuqABPvaRi3vqzc9LcE75zSODwjp
UIX/7QE8K88DtygxFhy+rbvLZ9iHaUtPkpq6p+eKtzDbwnHKGxS8GnCs6mCq/nh7857ttLcvO4Pd
7hO/pYxpg3EKqDcmXq25Uw+6N/F1nZH+EJYEosDTn7fyBBH8j2YvPJlOEwn0TU+13XHbwUSPmrIQ
gvQuNTA4N2rkls/wRa9QzIxho3bD5QxL6/VzLBwWrVhISUiHd2LCHrYbSSNRxkx++b+Xna4Lq2io
l7WK/TAWSCBdPnQGqlbQX7bZRfxPI6AtIVmH+/OoWhONPy8q7to8lGRyVuaTJVLwtuxyclpZoaEV
shwy9v7bae+GpQmUpQzXzb3AIsrD7htI2hfbNGA0i0h7U2r78VPpmmG+iWJGOaMC2LabvtCcpVeg
xhOIe1sUThXzrbkzME14VxMzd5u2hyd9Zpg1F48l37Seu9koE7XOG34if1sFOsl0szvAQ5ske1tk
H5RWfAUwHJSEJ1OyeiSdDbZmm4A8U7ex2WValz/Q7Avghe2TNZwuPD8y0227T5XBPWYkxEgAXS7u
JNrGgliryRP48opTx37dMrlgRnGvmsFtmWmuWFvg9ITXw50bxi28JBsotXNezi0nnsUH4lquQETe
RJ7kvjnrR6YKqfoVbyTr9RyeXupWUHR7nIwk7SukQS8beB3go1wIWddEEe7QRGPEqR0OutALjpEL
aryifkqYHZS1EDWRdETrWTchPwVjrK9Lq2ukJPkX1UGRSp51KWGl/rgFs+ASt7kH5orRw4zkBO83
akm9+fNir4y65xoavyK4nxbk7T1oA9iX+G7QHmvVW//Fze3QrqfBLSSWpBjGhh25mL3AzWxdLhP8
GBeqhbtgBchLeTE5Xipgoe8cIRp6PxeUHa1Qr/9TA3mExRgEvR0IjK+3/zJI8heH1mY8Iiaz/SuM
sDsFzPflAmxtmheopreNZVS/HJ2lqHc3Rrd9vAy/ImyHMCqQHvl+yfbnmQyhlsno9wJQ09iGZAYw
ntfF7gYw4rSlqN/4snL5rwvfwhfVHDZXLgocAQKrTqwC0rvPdBvh1y4/qNz2dvjT5JV/mKlMGLzL
vmqg+x8bLKky9520MNJLnis/MjfNdQDhkNaAWq7mf26AkEg+NqLmOxZZtSKZQ0yPRrXxUgdo+hrg
wyuD0sDjTm7MkHYkRCQxhdtfakoJ5H15tgyTUqDklg+2yomSdaBl+GNePfJwD67j1OI4BqW2N78f
D1HMj1ckkdy6zgpe/9q/a+8YSFMWhOnKZzO75sqqZjjkeB99n8J0SWSZl7IVhmsecUuiquwhP+PN
IDNBLknYfphXcbA3CV5Pn98M4ld5jvLMklwP5NeczFES9irYaDcGbKaIqHDOxzyY+ZtO9KnAUIbQ
qA+GiL1jgQDk7xYimZK+PN0NtF1RKMocmcT1KiGNkc2JuX6Qd5h5bIfu3wMXxU2KYd16R2iyVD8S
K3OIHp+zKszd9GO/Z63g+xk7QzHY+kYHsMxCPmk8eo5FMgI0qif3XR3+70OXSjWiXAQki0O3oQBM
OADo8FiGCmSrDCBQqqe8dChYGLVikhXxvDA1DeiUV9R/Qf96oHOTyynzsB/ROWhL1/+zG1kiuZPI
mAqVvCL+X8DaFt4+EBJA85mgG6nMw4THBP/mQE9BLh0Bqjx598thrXROtzrTaBWD3oqlS8eQbnaQ
v+rMSW6H/1YAl8OWSDMvTPbSiRLE/iiMJXEQCk+ISjRbjXfiyfQdHGwCVo725b//PxIauAiNtZBr
OQd1XgzN/xwBPtv6wwDsX7px/JAjby51Iv7OB2zt9G7a60YuyCsDQUrxjJqwqIYNioe76NAHiVzz
TDO0CLXK4rhCCAPjYjLQdvhYMsUJp+FUwLaUQo/XWXlP1P0NsKs+cPYi2CkVX16H5k6voACIkpfT
Ub5qmDWTVbrYwygJwniL6RNs3LtKOI1LCmYbPcICSh6i47guTmXVbtkon55Q5f03ZHk9VvYjfP19
tsvn3fpxhw2JTxTLWgCmc5kTXN7gVvhBBlKCYxJQAp7nEGy1AmVrzWuoxFlPtmJTkwWNAwjKMGDg
w9W1AV82rEp5ejWmI53m9tOpl09eGOzMeDghRO6cDbMmMD+xFQ5CeDRRTpVZXV8rbtPe65Rhr/8s
Tf/1rpHSgaE4vSWOY0Gw4eMWcmSpX+GIAccPtbLP+2aY8hJdXa3ZtTqsR9E9Stzf6khFsE0ZkI1m
FPetJGX88Zdj8/+FMYulTSOTXPbl7xiLTD+c2YFTyfvCTcdl1Zwrg45ISWFQkAIwhqcChPOpSZMy
DzJjMulXkRizDSgEtW5L6Fd5mxz4yAhxuyy1ghg6b3FZVou3JaZqzNub8ZWFGtb9pZ/cblJOG2wX
eizzPBiKBFJa+I7eYH28mAZjmfzw7GwzleXOgA2vR6ON5l0JjFFhTmJX5ZEtddzpBymCoyENUWCt
HItzoUgmP6zEbg5tGvdtrUsuFQLQliQ5U7uJX9Th88OH1kEmNZlSe1aLVEhd5Gsjt/oV/I9jzayP
vBzljMhby39bF330F+0lunPd68vam87RW1PBe2bh7P6nn7SfF+pNdWf5PjWYfPCC9Dpc7NCinkkb
SdJGEjV8Ivag47yKeBapOzvKilIaxvGFbSkHNuEkDybJ98e9YmO3VWc98AH9idiFSRInuRINUMuh
2EY7nV4UEK+fyx8rrglpmE0wigYUtmBsGninRFSbOXF6sfwaFRx0jzFoISOn3ROwGI9z4sXT9ffb
4vDDVLiFGGnUkJYqsed0ts820G7yE8QPYavSnneUFpZBAa7NJaqa61ghIHnRJICtxaGLgBxXsGL/
llIFFljV1zbk8kz1oO0yyJ4lz5txuFmF8VvBaPZBsHt9rRMjIhuPQRO3fV/E/0hQg0dCIHyLl6Mj
OzyHoB3JiPeutfq5yyIxK9wCV2FcnFRzQB5iaWdc92KUGGa+e2HE8TkHaWlXIhvR8syMd/9AzQ+L
YV60ZLOeFyft5OZQFJBn8itPBGoTmsIRSr2CPJVq6n1bDP0CR2OLon4SUJk4we7VNLgJNiQlPM/p
3oGUai48wpG779jEUt9/0afJCxVhx8dQvj6SMiKC5EtwUyRC4sJ9PWm8NmVKWZ3cFPoY9SfjIfvh
zmpSzDtl/xc7K4iXdXzfYl27HlOkcVWarHW42fPalFqzIz84QzVJfddwNqnq3rZ5dHgtn1Swsk6L
+zobGxX/UnJ/X15SaTvb4G/1lgsSVA2ibRBQUoMZARMv39OKxiZ3GD++QKjeg87RPkJbWMywH11Q
AhkMyriXLt4MtK4l/lwZZA7+K6gd3qAw9pA9Gz83M/+zSUrbUWRAWiWu4XaX7zrb88AbtTcoQVkO
KqG9Tg87iJb+oHgUCyO33EOs//Xi2fRd+7l2EHCFJXoflCwrIOc7g8AfwRdua11eYEFemG5iuKqI
Lrb9lzeThqKwUk487IQ8kqwSJxOTePaF4AlRdMpjxsBkXjEZfb1mYCvI/2IQmRLVdwtBq06TXa8P
tYhMjsekgln5KS3y2fkehi0y09ZVYcV2Y0h9PPj6Jq0LzUkRTzaveFnD4BQ1EHMxdk1gHCa+4KGD
AUT22sEZTEI9ns3oiVn8KnYhnJH0ngP7oxduyVrlNhVAZ9bLLIkbbJqA93AdkOi/eU9OpN78cuW+
TBBMIMUd3KFQfhmzpM9YDerC8l5GdAE3/QNR4gJ7n9zm4kBrPbUWoSkqZKOUfT2adfm2vYe9gCmR
ktt6I9oweDnu7tOJHI+2mL6l76zZp8zUO/hf3AWisxSWh2ioIreN+ispOqYB+nRW6AJ+Qc+EdE+p
tKuxqrF7CrcE80XDlITK/KjmL19O2sKhKTHXC+FVu0Y+tvcB8lWqy+mk0GgwmtsL163EVG6cfASp
FCsSoaE9lAEdjtnA1qMH7Z/AYn+r+fedqm7qg61CQuLfsBjTI293J1qeRsW+zHMMa/1s4MY+N6cQ
ChoDWRXDG9PWqNElUpXUaVMOz/VBsGoF1XvviSmVetCCtLsYjL+A4icdfT8x8tTBtOMhMVnnx4Y2
sj4F+cK9C3HgE61NUCHvZ5qLM1WtuvX+CC8rbPQwGoRyEJsXx7QexC7KSiES3228bqbccWeFP+0u
H5DlTlyuoMWYvYVBj47Fg1o8/eGU/qP70mziwrf2JAVseu1IMYdR1yX4G32jha7Li2qg1+pqBvAY
S3CAoVR6gJSRt/6J653Ub8bRlgTwfKz7KnK/QyfE2WufZ6ciFTzO4Xskt0yD4D6CEHlr6y9dB5Ij
fHK9HQJyAj+eDV0MT+y8inTG60jdIOzTug/fEQeqj1Fn0FH68QdDnvWb/mD1wtRe/oO+wYWcSGmO
9d1k8Dp6g+pAxLxqht+cJ0P0938k93iaFv9rmvDVy/CYcWoZw1POCKietl0ZuzS7aRQbMQGFs5Gn
luAdCFNBtF0KEjpKv4WaF53PtkiYCH98UXhkMpboQemwCg6AnXJRS71hbszVU+2B4y0lQBObi6me
aI5IlpH5z0xtdzTZ24BNpzhYHqIo7froLHacmVIE0Q2dEVEdznkA/WFS85+9zDEy3EYhXcV78zAD
nvuTWvlE1/+UjpPVgg9Ueh1e6IQsmoz+4tDQ1jk3oD4WUHpkiExd6Eq9rt+1WulWf4EHB6tG0W4v
fQ82wvDB4B48zjsrCaXYLuxDDUYNRTLpVgTvyCqQ2DGSG2Ok1DrNctTRF49yMO1a6PjWSk1kUvwX
kfj5i+yjh7vp/8uobkr+wtji0g4bvY4lNe0/58AYsiK/Fn4X7vVzGS0sRTXlChU9JSQ1Sc/QejGq
cHGOwz55s33sw1eS5i59MF33RmDDhpS8IvdArncYAlfrEwDRdaQYHNJvHEpmyHZqJDoU0BysuKhw
rqPzInTN1EgF0YQCeTN+qcQAnAhVMFkND9+dgExUxWCA7mxp2gKUTcl993TZa1CfYcYxvvQbp2ci
vgWGZw0Ak5rz5YEswqNfqMIPMLl/Y7I/uXN9mFp5O02r+l2afGMN33xgKH0VtKR39fN5UBhkTHbF
GbFMJgGJmxW2HBwIgJPwWTaCAtqTmLvbe3ypmiXyHZ2HCZGJlIuw4oiCAP3nSK+N5N4xearPrwn0
XayfhMS7JzpRmv8gd9VVhaQnwUQSfl/YVHNhIaRYKau2UKs3gND/A0yUVCCI6SVN9092RNgTIWtm
ckjxL047miL/pc1oOq99TDDs9TQP1YecfSQ2AbzU1im0maxfg6fB0pLTanS4PP1Jv8GaLp2zJj66
MWTuepplLz6r+aWWA6yFXmLNB2uiZVvTpg4oGbLZUo4UtRLqLMvebung9sBQOQJrzs7r6KqmKt/g
rAxjL7agyaJ5CIgRSQeqkoxrUtUjDsFTa/wdSq4U5Sm5lCzn5SGbMUWF18lDB6KhUeQG2MXVu0Xn
I1aFKMkoqnTcU7Mlj2jKqEH5kqrvh+rXp/bxVgQg//ymLUCmGoPUYQ2wh4p1VtfjOlCcIvpxUqgZ
phDRvhXd6q/quc2DA9x2ZJgb4cDoecAQdx9jBDT1uPTRaUK+LI5T+K8DIaxDXhd3bcCYTxcvnuvd
FGML6e8AFpG87k6RaV+Sjtxa/tuWsHgLu8N7EyaCNzi1LdmKG3GR08FBys+JaQsS0afnW51ZW0fo
MLwY7R7kqs1XPgZQgAY8RWP6o3G9F3c8LFVAl2g2LgmqVoAptOf3EWQZvq/x/+YpDhjmT8oGjAxY
vwHQf4CAHqAlwIZEZl8/A8V6FZwxCgLN1LT3MzxGhC3kLPkyHLoijsAbCUaMsHvvffWpBcWOuIOT
xX+lQwymuuWFyGaJS8vquUSHdOaA81MrUOVoZPK029rzL8Q34ocf4juHG+R2sL+2FWMt6aabXiAx
vFbgBPJFO+ENM/cKlS9cuRFFQc/mgg+X8NstVKdyNchFEXqU426kjIQVEniTj/BnJzk6dZ5gRQ3X
/fogaceJWxhkrM3VdCELA6l5G5JJCEsbin6xkxNrccoI8MYgJMOpphkkF1JJ5HlsK338puukDcsD
bX45HiLf07VHcRhy9Rhe8FSpGw9smQd/LwNL6l0mKhBPt6TZhsIapYqdZuIzlsLo53e8DFju5p5J
/vANmGytVksPmWSsvgQnUmo+74zFyT8PprjZVxNJzfolcq+5qBYzB5ZjuAmAvGlqlaJNj/gKr7KZ
JKGwCket642Bu7924G3+RvDlGEVcyKBB1RIKvVEhYU0ZbsofkI7XAtRLTDi/2Kzni6miUsCSDSSe
f6RMypFRrJswKz0PB3iQG5so7kd5nuhXmgMh42z2pLtbnWXpCRV+rhJJpvevsJpEQoDmpvgIhVsf
1oymY7bjxwLXVozDJ8RhElX15YHVhbTbrXRMeY/pGCv4o+8sWCYEjPBiASEQEdG0Ld+nmvMsvLWp
KahBHkW4ObMSNFsaNf6HreM618SpXALuTFT36T3AuXMqMAIWnpSq8d323Sbrlksi7jPqhtfkG9e5
E4V9LUDAdj2uBNBbhE30PU8JLa9/U7g7moFjJ9rfeZQV/yV0ZTfpGtgyQj1wLTypjeDJMKCyxjPe
sDI/x0AGKlr5enSlKUMTONG7Q1rYM4LK0YwYwJJIa1E8o7XpZ/oHUM24IiqhNf+zkm2o0jV143bp
J7X6x9pG2m+spL7c5Wl5fjLpD8OQIhPUVkJeDqfbsQzvyDuUGgmRD3+5/8grmLCClxf0UHqpMYMG
w6b6bGwHV+wqRkoZRL0kvYGS4z6HR+kw76feD7Nv5LX/Q8wfavS8QeieasU0LNcGraMKE5il31ML
prTTWvl2FOGIpsOuxbgS+PhiqEqIrHRVabSxClRp4lab+0NKUEgS1XeA580V2QTIRbsM9txhQm7z
7UPnJMcO8uyD10JdqU5jljjWv2CXRWy46xPXnmTA2C275+/Ji51ZAZPA6vCBCrongNioaO2kyD11
jAmVd7Q4YkWaKrw4rlomqTw6hUGAC/a0tvrDI/XprDP9Q+eeOJXWq4UaT/Nqp2trN6kdTkFy2svh
tXgdnWARQ1Ba6ayqVpR46wqlpMOdo3RM8Iu5NEBizUGWGLxwIrSqlVmG5rTUJlBdU7IF98daCYwN
DhVDzBS259shrPt15WTf+CvKq8+yeXMdYnEnwZlOdlOb5luPVhU9meifV0R2gvYRD9h/KkGScSgq
PuiN+0EHgFP1w6xPuOk8NRpeCzFIOD7m7RnxXgdUGYDsB9OK92368/VFNN5y0DWPuaamrrrAGoX7
njTKNLRutSmOs6Iej95dVZ6ejByK5COcNKXD/6eZFasbNiguve0ZWjkcmARWH6xOn0L2HK9hozLS
TAFE3cBto3GxBnLbohgN8EOFLQ0+ye73alaBZqUyBHUBkMDjAZH+XT2by5C/rAHMd9C0YRzwa6j7
N9vweUh5iIUGlTXW7cQmUAZpqWrtyRG5AAFNtDQC/pwtjJdSZ7YzDWBDGnwYAvwtO6ATDCv5yrKb
3R6MCvXLoRrXb+U4X1qdn1pyM4PNWcq0VSR4yCB3YaF0VxUvjvhG2/S3uOx7VBcCmH29dhvgxUyo
3Ig/J/S5yE9uhGFtIH/Lm+989TFkieThf5mTikDRH7cyH9ihIDq24M515b/Ogd9V7asOC/TpvjQP
bV8mClE/6whcvqq3OTEafDjmm0AlbXh/Q/oOreWJ2fg/0R+aJ9WjVxxoZyBI1H+UmtK9/iIJDomQ
VFXlNQ6Q18ibCNPdFXqJ5xrkQ76Tx3wfaz0biFSRZKIhlL5J40biMjExYABdlpP4TJ4MU6aCkcsl
3HKp6Tq7Oe0xKoN/XwXk5xGkRMzW/KR0JzonPhPk3/1HMFZ9rjtUReZQ/MQbmfOlP/JIdapjJ/zB
fdbTmjAu92xGbwg1QH0TkS4YArTH2IYweEoze0cjtlKNwaJjvx6xlR5CtMfbZMa0jWnq6rRrfjYJ
KdJsb2K2/hkD1DEJzQCLZ7if5iKNr0O/Vqi+p7q+o/FOeVqTnSukIMW4HdeMEleNZWJqQkSQbunQ
x2W5Mc5gVaXA2ZogL/hAwZtHSLNbKrY0m2uT/+9Du7yFr/poezoR/HE+Qznp1bOWkgfA7KVmvVtA
RSkJS2pTXysNFWuX723pC6YnMCLkaBVZH3OdXZsU2CLvEsjMHC5HTGd06gFT3/DbqR/M0RiPs8b9
liYlpfZU6iWgKXoD7KmTojuK5imNwfx0goHUXqfPZ/UrjVheCUfapyneO6v6inrm+uLdRmiAhiGR
m7JQzzhYV8sOolrGCMB+7+O0RfJxy7RKUUji5h5qetzVYANzvjDhCLaSK/FRpVQyFG923ZL5Zutr
nj4odGhtYMiGYvKUK/82GAPjj+oVmx81O/3slSHBhCerxCWxaMndZ1zt09I8i3hSmAs2tA6obIsi
74oEgMWGu+0kD3RSGZVPInOMDB87BXo5oqJmZOq7p7gkJ0ScUyvoHnXineWbMz1hLcMZt/H5FFW6
Fb7vmNUZisTxeEwtB+8U/sVmP7+UO6OsP1brhX+aqNp2J/RSL4gQiHmnDKn+JV2pF7c0QhUg8YWp
4BE9GC5LAVClAMlHoFOPC3TeVugSudtEn8KXDxzq96FgHEzhgka44fmTgZ1zAVIy8M16qu6495s8
8HYDet/b1hpbcjG7xzUYLxB24mWRmqdv8k2zTl4U9IUr98Q2W6EG3shugZhAPjoAt659VpSvIAN0
AHcRIhIhR/qTtKy+HSr3ZZ9BT8LBhKKIdyQ0tN2ejzgHJaR8Kfjt6zHenRF4iuM4+LBTaLj7XuoJ
21Yy4jigrQlUsZL3R+VmnZF7CO/en6iWhPIj3waISHc32jw2GmDDJFc6HzZp7w6XSMv9hZwmEQ5r
RJy/a6VtcaNkRdBkYh0ng0fVxbU2df2WKNNKQXKNXFyszGkkhkldLeGis5RGfzTl7IZmqxbBg07p
x3J6A4bMoQeZlEUgsJWR85vS6JYRFvYH7BgUu0bgUlict88STwfhQsCuqQc2NJjoxm0no4KmpMsA
rC6gT4cuhx8tobrKL3T+0GdSY9OsnrY0P1OAoRX0hMhn5EI7rJXGlVrPGrABQStBl9kUfhkeJbzk
lRPbtDZ+xYea6DT9FyRxFYSrbnk1U47XBFdbO4ANdy4zYEXCV6CMvRcUN71HOanH2XdoU/FH71Ar
80laFQYY6R4YObVis8kYGShuMRt+zmAixbVHRMdxq/zppsPA7iB8mOrCL+lVxs3fYoAmjxtSTnE7
/kuEJDPfOMy5eQO+ihxVfX7DZ6EibmRAUSCNO349rjwq3nCdloMIFNv2EXV4s26i1BtQBhcdT9fX
xQoWXAx2Bk/HgQ5HxSwuD5CboScxIS7MfTanVib9gL6PUOjS5fnCduuyyZxE/t5vMjfyHDe0/13Q
G4kJMMGDC++aRGDbmrR5fZ1Hc/7NAtlDT2RQR87fV88oPL+zKyv9BqOAUKrcFSgZ8L6DTysqgnE1
TcgLiLfTuoJl5XKknTF3duQfL4xRzZGWpetyoI6dFVns6xGv1Dgy2svfIa5Hb1JHMIIJsQCQbkW2
/KuLXreYYBaWQLK7UZD+WA4jY1qGZgqIYPw0Y5fSF8BLJC5ZghV5AAkzPDvvZByjZZIt79t48rIx
c3ZFeBgDFABBwSy/JW/5w7ht50/YvMu46270/YynX3rKx45RCPDFwaDXVrka8dxROibAaZqi40K8
/HyVsmTYproi+vnVsg7wpw1m5adZiHribhNPC6tQs8+fewv19NNmqJILprd1Kvy9TU77bUhUxEF8
oMj6z0qW9WLKNeIXrSxSKkXyHaE5hOX9mdq+/rVf5gvdMxwhwr4A21aeBNoA6xVgtPG1IA4QB9gG
kYNXj6Avsi2LoDnDQ5uwUTCIMqhK8pDbsNvA860S2ssRBYadnl0jxh2k2OCXOfT39E6+RmPfEieG
V2/uaCtfy0fF9msDtgE2r61kXLq2VF2P2mZ1dCwBnBb6U9up5K1VHO2cgxguK5nI2brqsKmOpCRK
lsTr3k/ZjpP6OFhteQu+TAq8GpUuY9DfKcEE9rPiWiQi3OgiI7mbUMJJ3Se4it0zYEvQx9whb9E1
U7uqS4XQihzqeTq6LdJkeBPXXuxF2jEav24henZ4XJTHVI++mFEwDFU0DUk6bhMXOB+vS9cxWLv9
/E+/rpNenqZRdYR6ltWicplpflICqy+huOzXDa3o7GHnZzaKRRst+qXiMxCNuzw3jmaulli/scZo
dOhtJDpsU1eNBuw1fzZKhqV24fkY3tgV3x9x/8tq8mDvLndNWCpOLz1iENrAO3uiWrTGLqKWNpR+
NT6luxaGuQLxd1H2bo4yyZqWTXAj5hqAtFNauf74VfDzoP83TFPRRjkMEjB/lCXLMRgsYow2DPQh
DWePy0gMjQYcHUeKIV0k9XZtJVcxvnAx6olJjJ/3uQS8/qp10/LIYEAWO0UMlo65XQQUKdEYngsw
RPF/frF0oUm9EVADph7S7A0mBQlyAGEb/xmQ3nSa4MX3LiDYnn7l+xlvANjU8mCHVMA8qcruT80x
4k8GBa1+yRn0VW7b8uRTMm/ExBu35ZEE7VR00aIcmzGQN2pTzgBGfHsdVSLKg+uqaKylJO3PuXgy
Z5DR4z45SnVrRMs3e6SIevyGiTToFM7kaG2KEyuE3N7xJSBAufEdluwv26SgS1MdFMpPmdwsRxpT
FwN1yphTJVuugKS8LLY6dXwSQE47W/qxIIQGVAA7P/sr4+TnG00u5qU/CllKXxAjlmKowGJTg1wu
g2haGn9ge3bwTbiXW/GkFkClKQsc4ppcT76+U2PFeRNU0u3BQwmnfIw0N/iRlO3/8Vu0zoorhjkT
vf3I2WBsn9hbZ4PgFcaCM4Xg23lvOEPyffojoGylyTpSW2COIhLLQlX4f8aclM4pmVk2JPsKBCRx
9KN4MlbG29Wh24LeAkn4tqNyO0zva7FYsCnGhW76+jKFTqGnBjzNwR9l8yKdVKb6mMot+n+y+GHq
UwnWaBg3myvRWb0uA/YZOWtmGIirEHgeRvrG35TFAzeXUXQoVsWqmdB3b8cZxm4OmPIgecguxPOK
4z8aqknbf2i5b0mShJGVCbVPiCQ3WJ1CmvwEL0tIwGz6/+AFOuLjbVlq7HoXoYbz/2p06ceF+MHd
vLZnU02WrRtSkexjspAE7C4En7hLd2tizA9YTZd+kkYImnefJCPTqZ9MtX6pZ85Y7oGNuMKVKUg+
PONkH+oIyKQ9Zk4DAfSuQsvlkEuP4tw9BWJF03l70LS65+7adZ8r2aNOSbILGJ7t43vXdZD6DcIE
G2kl/LOEgpL6CNhL9MQFMYYp0PB560eC73ttTRbR52bbo8HiN5d1ZcJedPxi/WJK6sIavGUyEIPe
Uh+hA9GbaNOCEviTm8tCTc5bERMixasm02m5YVmEGFFk4CcIGTyZQR0ZKryovFbL/hykybs7DtmT
JHCDpaCGkFN4kydWnIvhD4B+y/eDE4WzdoESitZ666B0GdRep/ztL0AnNSWwY4vCUtXpksNygV9T
8uObmY93CCuG3lTfkz+gdh1ks1Cw533PTFnkEYwQ5iSy03PM4e5OlbdN43qQmzATtz92aj4FdLAT
u0YBl6xVGU73PqRuWDKXE8ehsPmLCexg+CoFG+Ycyri6S62SXCtYbSnsvBLHVEw2n3HzCbSRM8Ts
Ofi6SYXLSfDYyiBATJmDQ5WRDV023afdhaBOwwJh54o0HdKWg06E/sgJdllvbO/vETs+iCWqjbVg
P44sIPvmAmp7EmLOp5w4VaBCsqVz9Mp8kHrGWrys4pYSm7ChN39fBYQhYZ0NpLKh986hfrV89Ws6
wSHtb2hqeA3eLZ24/+qvMfuRq8FeGvKlbPtqlOMUgzq4C7tUFYouLfRzeVeKc+yHrGD875MXnYXa
t7p7qKD7KNJj39MH9b7CcCwLICXfBD1b4b4k0ThFh10MSdLBJZHeWEAJ16SnHiI36lcPt0lYd2iP
skn0CshMna2HbEm7Wh4gmJmiKgUMgAM9fE++P0lB3HERgWu+jIkWRReI/GXwbqi7KcDJZ/fXvflm
CcyvdIwXGo5nXzEq/qcjpR7we6/lD6M0Wg8VlTAjB1wPMc5KUHrh/rYJ58Eb24EtaLTAu1kBiywJ
rGE1xYeoLjji9JUbnhwowMTAli7UjIkwJ6ftKSGj6t4qhD3bFTmkx1zAnPOSYoc5oXqURKgOctzw
L29BKq/hfE9gCZsJ6G4xY0mWeOflbhmuMwsPv635405uOZ4HJosQ8eYrmoVyPbhxXj9NwyItbTtm
Ujb2qPt3Zm8zWCI2npuhKx9apcL1vmQlINRWd+S8WWZFVg4zG+YwlmKLRnXHf4roLgLVOnvWX6lt
WcOt9bGeBLUzcMX8GrXwt4wu4ROhq6/Jr1yd0rnMkPisQvaGU7wWqW/WLWmPL4m+0Q9Lksm7UzIu
ImontrAZ7JBZbwMj77zz2kYTlujA0Tqnn0qgAE7R4foIO4zhdSmSHj5S4cfXjMvQx0WVVX4gx4YY
UEmOwPbMNg0w+vLybM+aZ2wfYZeaDAFfen1dHf6oZzheLVxaKJzLdgXRWCsnm+f+wNlLzKxVuIv4
LM/11myuF7oxLfgiR1nKBmQ3GmmYCtRlVDPq9nwSo4XaGUmRPu7HU+bfp556YYa0IYRuNbJBSAiG
SJoYBj68amX3EvPx3EBmzbKihZQ8OeteuGe/3QAPMC9o5k2D8y0oXQ1Wa7JzTsmD5yDz+p8Jurr4
TRXkZNovzhweQh0klgQGmzk3TSosL+KCvgk3aNdZ+X4x3PXsU1+Hj0mbjhedGqSZSKV10r9Gmrcu
zqrhDrOIWisimk4cZ8DJZgsKUz+yyzUkgXM4VuqHDGcFC979B9jHTqND7W7AtuehBYzRH5w9LK3f
7vOaadDUFeSc26SY2wh8alIrPauf6QM9b8CF1j2jAlifSmxj2xAUPxex0yuxvJ8/WP9zvymdPFgI
qWlk32bZwJ5QkrUqSOouGyFF1eSNc3WwPcHGLu4f2SWWR6bb1Nt8wA44gJaq2HTOX8bo0kcn4sm7
OuwDNgJdeuYnkSqDNA7IZvcD642jKuiLh5w65QhaAnCSgzsU8hIZnDt7ocFs4qiNmB93TPG0d1v2
ltXCRUtllU8PzSl10n9K9M5jyXtT3PIJsIz9P4dPwbkVsNRm7nlGF6hzPGdp34YDWCYbxM+dhW/I
tbQknz9fHJM4ZsOQQa5Kpt3Jto6dKRJ40/4OVG5aJOjA/KSzrNx+1ZhazoS5KOA1mGtsN3/5ZzgB
mdwdbXNvyo66uklJZrBF0JiUSS5Dqf7F5eRMVD+Rnz2N7zTgtMQLCY3dT9xcwpj3d3AAToCCJ7A+
K8W9hdyYc0pBi4SUzZbO+Roeurl0Qrc+IQ9Faa8elU5vSqcKBBAb80cYViKO1fI1GrOWsEjLBwDO
Nw6GX4gd1ziU/96GvqM3uE7T3e6tqJQF3j3Q/VdMw6+QQ+jnGZw1ObrnTAkqVFkF8Eu9i3eSHupX
98fSeCkNTIfPmc7exHCLLDA8KTDkFqIhnJcWdd3EwGdOHKC1xDUw0pSXFZq/YSBRUn9X7OBzhVR0
YiVROA0M4nOPsUsJQK7F0h/eNpFp65wsiKRLpCwT9FP75V+Zde0HUPMxC0m9KJE4UGkZW63JhvPO
3UMiwUKdGQt9qxroHqz6mTF10HKsq1a2zpgG4gEPIS9DT2ZWTavRMaEIuyepK4edjyebWowalnVS
FgZLB7dGfRCRrL4sN5inzXZkW5Wqen7VjLMha1KuWLeXF+5n4IAt4Oai2a/C1fOH1cHdwOeseEb+
aayeJkUZnXuEFegmvm0EWkgjcKT/Vxbn+8h+xngxkqu3idd44+xEKEQoER2ICvAV6wAS/BphJ4FQ
eSNjpXpcw+d0FXVZR0YHHZMQGXB6JlxhNkweebWWDwaEbM6mtutcTsJx81swkUnR1TrhjJvn8Gaa
WVj/ISRk3RHSd76ZghZUnTlS6L2QfPbRGxqNWdQ6wMELCokCD2jv5lA8BElkz9AshzvCAj2/dPCg
0NwcFKaY1o8mDjF9lK2olHksoh9q4KKPpCytlXRfKhP10mGA2kpky5H1MaSonxEnf+bMWpxh5gp0
VgLxRh0HWlC+ksqSEv1hWwS9WKuc8R4c4ZWywASmaDgi5Jwxd1eNPXdldZxEvVHQo+1oMSR/gSJY
4m6SHqZMolo4N0A8Hcsb2sB0ycKpwJTwtKY4o+q3sQwPPJdi/NuT7EoCULl/FTDke4V0Z5F/PJ0O
E43Ek7IbWg5HpcwnSTIyLTJGMj5mqzMEC/+0Ei7pKIhrS3OhK7Hb0eaTlKjoy7Uic6+zug/Ra3MD
1RwDGCZ6yv5XueuYx4VJk9yRq2RJaMbAve2eQGGPuoKJJdTmmTN3EbTUAB6VBXo8p14wXjRlIxk7
uFTpbYPK+8q90PD+kX+4Fa1LYns7rhk+4l0FXvBaslMPLrL7kjersYvMERC2tnivV21QhL2eH0FB
QEJHpeeiinLyNA4X1XwzaJ8koeebrrSPxdL/74WxfysBQ7wflb17aGAblqfK3rnzyHWFBOUZppiY
lMNE9dvaAD65Bl5q7FW7bwiVk5SlMpfhFRxVjztxxjNozuB+Gxmk/T0AEuYudWEdgYFzfcez+Mqq
4SMtAjZ4fmJc2hgqmNXTEvUYa02Mz0Ee0/kBgcV/J61ZtgNilqqWGsWF8OiUvP8GY8upYU+8dkyS
vU0q/AinHKtK52U/FAtijL15TXVpy7iQdVSnQJ2wCcAM6scGFMuk+7TYHwAmjTH99EAonzojks10
QDLulEQhnPBgbJOw9MyOSMxg8+8bEuuV8V5okViwJ+7OwRiqVLLtU8m/jcCdfbRePXsfj+7qHoqj
m+/xzWf+1c2ZmeB9YT8FaYiNOOCtcBsriVlqIMCrHGJQ4PSDgHGzg3+WrQ0rHkYXb8jB7vP72VK1
JHi6QnijK5+13APDRmVwicOMEyl79qEfqcqhTU3XfOSRqM8FadIsUbiahVg3NuSEhcQ/Llb5C4k9
uTuXi06sxpLgPhj7cHHpy59iUbRY4740Dd9Vzu5bNbRg4ZWyjmBLRbqh2p0meW1Y9x0hWzDH7b6J
aNm/nmEn2UGoLQt9mGdKPZ2v2wOZi+ySgiPUmGclLO0Twp8o2Q2goXwkohJ7Hy/hUB6GOWFYNSxS
fKMHJqII2dDAOKSuH1DmI8nOIjuzZ7WxQNfLWkBBorGxTBYjXgavGg9RI1cBcZqR+Xpael2/VOSi
qF8yknOQD5+XL2vBMBiaQZRnb6gmwWjbhQW9ASAZBWcYA3QwrNF/hmE7IPlnmCxIxkOthx2e4pKm
GwwK6XWRevrnCKi2+RwRVIFqeAglXQckt1fp/q8h9Jrlqq6eO1sODbI3sUuDui2KKrQsncpT0a7R
+Nk8kKvznllx2ebbNiCChPWq7Vqgx962cxMp6R0Jf0RS4Npbf2TKfQuHneAZmC3eSh7KjSp+oLnz
xbP+kLtKCCTiw5M2X2uVq1eZTyPmJ/DggijfxE2PMZr8aphiGICq5p1f5auDiNZHl+vO/r1aKMrn
H5xvILHUN8LeVmbUXRxuTYtViWrHu8CXbczGkL7De7zWD9vSpJBXtMRbG3olNNoRdjxfZv6WxdBJ
Nob+Uu88f922nJGZMnk/gmTW7DrxTItaQi2TN4ddNp+Tk8zykv9jC/YnmZtXj0PMT+7eGT0Fco4p
qsB2dJYSVitqczyPKH3voa5lEbwVaDIp4qQijJtRy/4VR+3FLcuf3Qx9QIVj5ujTYlTjGalaYhHd
LxiPVtUk9f/oAWHP2qN0CwaNW46qmKqUbYbbPvZbw4lQjEeXlLhLhwiSRiPuzI4z9tLeFLZTKFUP
eCNQBr5bobedLs40ReQJQLJyTO6VJYdojYPw/RhUKdRp2xloBeGP0P/rrUvAYOcW32Ok5K3HnEgC
iGVHnucih6qK/ZCin/ZMvn9X59RBgGNPOcIWtQGgkC++vOJDQL5T+PVyskNDRV02dZZMoFE3OX0A
nSS2fhApEnVCTgIDAsUJBF1J/YfN0yYZXZM5+XN6Vufv2bzRbDzGBw9PiR+chDJMBpa8aWPIUxT6
hRajN5IbJT41SiEF1nYf4Xty70NiUY9dsLAbOds1+KhWN+/AFlWbn3DvvndR+Em3I+OWHFZ67Z2E
xss2Sd9Vf+4Fa1bQWHbUX4b56Msq4p8t84ZG4RUh3n2kHzIvybM8JgeXSxgWcPJt8ahYMPJOucoT
PVf2xaRNq3xrAgePRkcphC6R8vcRRvlPUYJfzrVGn7CG0TFLjdooLeIsE9QzX5udCg6yIRIgljmK
CS4w+panmqE1vWclpvJb/uJ2zmjqNp/XMFVFFekKJvjMaSYZv9CFN6SdyeMBwcr2Bk52EMG741pX
jHrOhxD66yAKjdSOIlP0L5sXvUoIbWxzhO8tUGcEIRc+ZUNFiKkjvPQEz7jQ79M8+z+5ypjVoZsw
MA+aVhzg39M5mY6maOl11Y+8uc1XfDn/MPa8wR9qsLjG8rTNKZUiVeLSev3uida9dVZQ30p7/IZy
vd4p3Hvo5V0k9P5Wj8P5ZhzWThXAPl/oAPXNInrWVNTtHdGGf3cIe1Xcx3IWpO9/0y1w9/9nbF3A
bWXvuu36J7EPWmUmBK7QsWCD6g/6+pkb67UiIUEIqAFFgg+TVN+0lS0QnB/voyk21qZE/ZvHvuZa
UEW1Fb8UyVI27BeD02wVb2FaKzeHggug9qjPKFwTitjHEMDJhDrDIe6RS3ysNNM3eeyLiQKGM5Jv
C0aR8O5PA5yi2HqFZ3T1rqsxTg8gXHPhjKRKi9a1LY0RuqgqWccJNEkxHLPScOk84lFOPSd++mcG
R08KStG2BwYYwxojJo40IvEXK0sa3mvihYkGSxaurrUhVHkBR6q8Tde/pqtnie+cavc1dzCatAcj
+lXZ0t0PEzhdLZRwGwZlCxLQJqVymUm8DcEWTURR7PRYRiKdXECQJo1/lho+aPTodcz3WESY3aFN
MO/GQRbcQ61exKynLQIjQs37iMMvnBAuyPsy5OaUFK/LmlFurC+S9hcFmdkUHUWZ0AnjeD7kPK6u
B4vkaMm2sqh0GbovzCrTU9ppmvGikGEMRVLSx+6qPzTn7BOIQTZCVMQ+mK8S5A6XK/TCgq3VzRmn
NaONA/7pQRbGUvK5/dFUs3b6OwfGqLGa3nLdE9JQvv6lOPj8pCDF+iZnIcNBQov/xAyJ5OaADHyA
VTll3XSujyKXfKq9kTSPzW7nMHlBwOmyZ62+mpaRodvXCV1mnX9QUd3quSWYOqf7HIgGK/NV6mk+
7JqpsetbB84aAL4WEDH9zEpybuKxJj3AzwbT7XlZNhVdI61tFFr2fk1PTxxikvgW+XmwFNQ5sLii
PCq+enMOavlgA/hAbkuMOOqt1Hz83VPeaIgSk0QuECwWx3AT8l+Fp8ENbSUepb4ul1p18xvoJrvD
vkggIOzRYdZswrpJklMtuZs4AwoCvk4veghpQep6Df6jqrJuMHiiKLNsHcVxqNJpx07OHi8Fc+lr
ZpYMGOj3trpnrjaO2Htpb8buWyfKBDBv5AIgnCez5tqpl+ND/E8h0OjFlELv93GsRcznXj6Lyg86
q/eYDZp9EAvDa2bagXngwgQ9tznfIf8nuBz10+4m2uMbGhMKLcfMcl5U2xMLFgb8+8UenH4foq46
g82PYNDN/tApRFFydIBvD0T8h0vCdTkrP0SwWqhhkWMKJ3SdNMU05TQrxgn5SK6eAl8VvEvrLon0
Q0Kc3hPdF5uOo3QIEOH4qmzijQqwKCERf5rGjLook0RXpiFy0fhct9Gfdq9taeOlVW2wJMvtF+Sx
Vq+YE4CNco46FaX4j4eWkGeJBGBdpqFyjSsd5Va/vT0pCo10ey6egqVlnJmLN0VVr+Vygq/DV6wv
xzYYB+wLb8lP1JAMAlUK1T/TaAfewbnzoa3iAljkOdG0g8KIH9ulR/CGQB1Uvccc3rcIPlG+88hD
ucOAZQu1GTYx05PLnItggSJ3Qr8UqUoj5OtciX6C1i1lnMvkRyqoBO8STWpyhQEo8S8vR2DkmE6u
ANM2k7g4rc+hgZamchoAA+tdPT8612GehXH0rkdUwcRvZlidXMkUDilZbD6/+fA3IvOz36wuxZdk
Ksm8Gca51AhISddsS0EnKOBWWlfG7UzqA6foBpFcoUl9NCwe02vNloeZFX652l4a3oGa8A0hbCbH
gJ0/qabT5LshjbYeuMOt1CJyXjC34kv1bSmN5Rc9p0e7RGNTJC7Ht035zxx1+FM6NZpDA9L2dF++
YgvffVkKYM1wVLRx2qcXso9llSqQIBp8h+KCFBGp4R4KXvOtprqvYp70gMgvsNgf+bRzTUQpOfC+
+Tk1pp6tvD6RoOGp8xSblDVO/qCvbzIrN9Pdo3zklBHynudIG7gVQVQmS/usjHcKy7YJ465FQred
StfZVdNvwkjEaiANc5z5wWXom8ze94QXl4qr1JQrNGeKXcnLeuAfpYS6nlVMXGRoOclpuGyT910a
ZYNlzkMEWaCBJGe6p6W+Svksuq31D9+himbBh6ePBJvMf/URJN0ZRW++spWqKbZ1Yebw9MX4G1Tt
KvizFPxg9USR8m1U0IeJG8rp4H5gJqUxPj7CP/P+fhjhpDruIc2X34SVOXYPUKmAQohGFqGQ9PCO
qNbwKyeaLx7+6xrQT+3pwd5QrjpWa87BJ3fJYD0aeD82YIQCf2mQRxbG1uI9x4qLA9uISTfDyAWi
kJMzK32uBHXPhUN8DRNw1snX7mSaf/qpSduwB4oGnw5UarZB6EBrRCvx+YyO89O1o16vSZ23LkjC
161iOHh2vhOVSjaUBBk4WTpdPaq1n6oxSxs8jtrjy0O1ifxr2g4JQJnhlXOAXvYw/eeAcAFESGKm
UGxpGQ1Z955xxh0I1Q3PyhiRaVDandRY+G2RkgY9Ae7jowVo/6uHnnDM2hazxXE1nVZPpEMGs8P/
FqNZU4E4tAJxfulAqH0r7c3eu/3T5Wgrk2e5DT0fQ5w76XW20huOSkBbwofhjgA7+KRnc6hBv4gv
/g3crEWtkQ0YUantlyZTQgemF7sGO8xPhs8huDZQgFvW23+1hIXhtvwLWbKIRXA3xvFMhzq/gLYG
l4fUVCngW6DRzml2sf+dWcP6DQ26On/YtRfTCJpgc1RZ/MBr3D7BVRuisMfu+qgBQsSx1BeBhU2r
ONbMqLElDopdKaVOhSAFsBRCVZ0ldEvuBptRYtRQdq1lGmwC17NVbO/oo121FxMB3R0IJ8SySPHH
YKXzJ3FhpSO/pL9/aHwGHhve3yz6qiz5FXRoo7xNaMVJlydK7U5AphsUVCWZLrhyEFjkCnXeCDA8
4If3gkfR0rFrdtlRr8Z/u9PKKenJuWsieA/8ewd4dd8M6DeXRO+BgWUdbQdWncuWBOXWPbWe022R
8IbAPP5AWVjNbD6G9i+vRHI7S0eQh7vfaDjUFT+dGOxVlZ0rqJSIG2afm2yB/ncz6Vc9s+YCZSas
i9GYqnSJW8appz9u+FTehzTAlgiDn1h1StUgTgHhOeGpMkY7kmTRTaOuqVYMM4A8w0YIoU6VVeQ2
E07K1k/9xWUad2MGhS6WFUcXvRV5mPhQcPHG/qJKZnxpOgq6LPonERLep84UzUEQgnpGQO4uzNYW
vgCZ2WYpuGd66vRWmdDeGDW61B5TxDiFVJ7kQFO5THea/W/5JZoTFYqe5R/eRnwR0n3Ec4UO4tHs
AXyWpB5BNtT+yey/tSDPMVjS5WcqUFDqW16U6TsAMNhJNZT8ZdnVKNPnFbD/bno9bgPggl3rh+ln
M4wSklFcyC5VetyPZD9sfZpV81aSwIwIuP3WdmrQllYUk6DUE4IVDF/DkChxXOfQmiaSltdDmVxI
QCrqbvsqAwijP2YO6x09TV5EQNDAVOqy9KcK1HR8+0R7txRgnrmOdvHYpesjZD0cmTkdyO1o7tZJ
CJtsVL+fWijcs9k/DME2uYFa0cH/63CkGfQpGEdgn2fBNahGagGO2PRGoGpsuna0+n8YxUgkwTUJ
S66NX3E6wlw0b9dWb4fGlwh5sIN0bGp21JdvevjbRrko4Zl+G2ncyjl/QYaazz8vNEgmPgDvXP/n
Z/70K6rKwGoW7yj0/dcn79YfAQWrh2Q/u5dc7K7HpZDqRjZ9dDR3x5MVX1Ilid2jJzaY3t9li5qm
tXfuL3eZ5tgBw3dFr/enzXoOZ90KSO1DuCvVa/Pljw+j9ZPsxlbWzuXG4hewbu483RO9MPaMLXuF
h+qDNDg64dAmsSvjlE6sZYyqPdaW2S06sBgi7NtuK12j7uhWwbNgIKmfKFKEWbyzzdO+ISnAkuig
cKL7bvwOmI4m5Fxy5gdvyXTo2DaKpDmMSqwGJbfcHpWPj9KyDmeIjCV5ExyZrIv2rIhF3HYpAcKH
hpwSQETVeUPOVbzqRUCotLc7nmjBJKfYOO+0BRO/hsVhCwnV5cYIrto96zd5YTJB+4oM9pQCODRD
bM5MEj8lX4fHcuQUiPJcWYx/nn+6ODe4tx9GICZp51AkW7UHnPcxK1ADK17FZxv3jcDJvXQrDJwV
a0MEqi1pbEnYLt9G/PGs4RrDtqxcBapTxS+OATWtx8cQXIZhx4ZPND2/XYliWw1ob8NNF2QOeiyd
x67Cf8+qQVDP8NPDqNufbOFowNRW4xw3yb8zg9+gUwPFAvCXtveK2Ci6gKmoNMSXDnlaQTnKrrIA
DgjaU8AyEMXIgUZN4IPte8iSyiM+KELebux9wDHfYo2aL6GscJt9uDb3J1sGjmfNeOynolnggFSu
5pvW4FA8Xs9LjZwEUZk9mcFN3Tr3XXFbktM/E/jTu6oOuuJOUwaMDS5vaNzWu9KUT30bp3qzL3i6
OzXOYT9tXXMeH55K0oc2OuKuyLrUJIIaWWPfxL4i+nKO3X+AMLTFZi0SKwEIDNlfVBJ+n67YEEv/
MTN7HlQEDbyewGTouBI1dd6inOIiLSqqDy80BghG+7W8prwG1PLd2Cttt9MPbnMtjspW525HOim3
P2ZWYu8A1HxKFW+UtqnsUWcdma1DaGS3MF9GNwT6wwHWJqgPMmE3fz/d4DRZJDluh8LlskAKcvEk
z+2cqQFejiCvxQXxmfWyRB8ysVi+IU+CZX7ZLfpgf4/pvYV3VEpCLGn7DblBEtKSN7GSu+C4Muu9
O7cSPZ7RW07n3TShJ2zl7QJXvSo0PDomTVfW2WH/+dOqJ2wIyMGLCcVq9fLhpMI7edDuyxYJeR4K
XZw+nagr9YP3B8at3aS2gmRzk31eRo7SiEAVf7cw7hEDeT/B78Dga6H/Lpp0WCAxP27D+hvs8M+V
KztoD5xPqyg76wTEMlGKxi1nbSOydgWp93zBpNDhFdNeqin/7T5SECijkjzQU7Dr8eMQY1akdsz/
m6fC8+dMwT5fdNLrZwWmlfB2ku3pXM/Nfm32friDTLzouv59JOiKIZoHXJYfDJmOuth3CGzupyLb
gfnbo0gVpKnMjd1AFntRoJfk3NouEqeHCSc36HrktMAnvIOcGR3ZffwUNyUQ+UrBj1viBC2d6IYI
Q3OjTKVcEYgwieMylcPW8G9n+yg7zq2tLz5vgQ5wRD15gLj6RxQF2VbI+cBHZ5WvgjOx0PwlLwMG
p/hNVsIGRrgDDhsjiygWRIJD2HzX+1IH14+j00vBnOADOX8IolGSkrCwJ5UOr45LSh0DHAI9Wgn6
qaD/TViGFlKbkUSh1zUIkwSX8JSaG9G51aTtUwBxMRtuQBN3iDrlWZ5y5v28gPVOWTsK+HrMzLeX
jA1UVN/pB5Fb9jf6xfsH7VCO6iSf698p71MyBhmYgRFUX98HPyyWCdmDuD0cC/G/txNNGUjro0DC
V3yHHmufRnQLqmCHIujiwZ3ItsDhV1Pk2CbLttJlfEHhcQo6vOTQLORcG77Xj3DgCzvkh8pMH30b
AsuYxO991YnX4RkFZ8hquiyg9P64gEG1vLZ9JdPDAbTdhhxO/8VUo4Xt7TTaPt7daZ5X/wgEA2kT
ntkRR0tSQ+aVeEeG1JpR0V3zpMDjCOyVpPjo4TTW8jm7HdELnLUu+kt2eyUKlUQy8lyWh/MTXigW
ERkncjkIAK3s69mgbjKt4dUbhxD7lHznUwTUkeencwX1DLtboMxUZg0kcHChhDbXMcyWY4xnQ6rz
8hvBKPGpHsaUFkv+4glY4rgdbCrI9h20dHQQ/DAmSscyePfne47wql2yGm4jjmWfdnp4NsteDIbw
W9uX4roFXXtN42qKhCleIQs0boiQJ/Qws6welCtK3LZ8vn0rb117tnK8eq10oaFHXHa2RpLBbiNa
3x8TNQaBrsbzXLr0NHKdt/DJnI3UwmOq6Wv2wEe7UOJLND/sH9zAbX7xc5jLmdgPFXhsztRRQzFW
Up8pvOq1R6wEclIsFZS85TFYOqKbSCqw/z3sNewIfP8a29PPVyK3Cyp89JjtkWU52ZGy0ghKTwAa
NLRSCzoSnrH7v/sldHgTRRebXJBo7XB3dqojJX8qjh+ajbofsr5qcoI8evUOLiF2hR0NwWejMzIp
XnKbBHVoEdA8HTJq/zx71Vd6qypksdfoRFdm2+5G82UgjHyZAQGyX9cwyKF90gSM/hDGgJrYdTyZ
VWsyF0WbtTJPSYYSDbkTnHWpbC4ftlk1jw6WPeAM73AmpkrREiTvseeSccZ+6aLC6+2VNSSIwoJa
xYYiISaEY7Ki/tRtlU1A65jq7yIVrZoxPBF0QLZ09vxcCJQ5XkWNVCPK43xL5td4pdexJrLKGcRK
4lSgYD/icr/Sx3xvbuwmgORsCMGBVjOqt1fjh9KM6aaQ9dDuP+SLJXn3cxt+e4n/czwv5Uj+j3Gq
IRo4uJAM61hB1oiOiYlOciVyd+etZaeubbEnflmZ6aP2S1ucQv1O0oLrkDfYxEyBV4MsaWqwDSz6
yAoMUYjbnG+Tf2kryK4sKr7tRmp983bPtnsH7BsnahPS52YVtTxE7416BA+mvbPn0lFqle8xOf9B
LT0aXo+7LoYYDQGW+1dtC5R572GvC3npZUkfd7j/nSL20DHCwx5zsu4aNojGQ6Qdx4oQEd7Zngm6
GHdOut1A7nnmjXOubdE9xx43TKjWSnbjqnsxApkQXfDNOG9UlB6TOMIUL21ktwrHQ0BhiRzR0VFL
THmfVQkzfl9iGy8ixBjw/P4uQ+3vhSJn/stoA2FVweTcd9pTCQaHn+s8pNCW63m9JKz81vV8yPTZ
Ux6moh52ugusW/v/urKwDXSyPnvawE0NpVpPKZH2slgX5LCuwwH3qv5jq+JpO4bEW0aviUj2X///
o/IsfCABepd+Qjip+zTJGsieGlpZskgvStJylFbsRGP6eyi2kVZksH5MiFSw7+1lFNdTXYgy9APs
vYHmlxCXNgMYadVu+Sh1hvvcpiXseePirNmhpYo6yFgqJi/Tw7UnLtLU5rcFYvtZE7CS+bSSNy3V
eiL0b2hHBkXRNlSvmwAZUfx1VxY0SxkfxHwFDH/5HA9olZt8ocjNQJ747pr+jJOMrC2dE/HRJ8Ok
H1KQhgO3wyTk5zJVwa6wOwmZUhY20wA2ZCiM7EaVKyQxFdi61o7PY6mrO+AKPDzJPwiSujKQwU9e
gpLbd2k7qlgfst3vNxw9Sor+VTG5T+BELgSaPg1XGMLlnkJ9+Xok56aNjIpVMCWHxBBddpwLvtAS
JXlmFRbY9rAjUgzuG7W/l1V+hLZ+X0Zj6qgEHwQBvWqIc1tnjM371ixfbf6IgAQzHg0VylpnVJal
FE4p3bjLR+6p49wb6/VML8120F2ua5s3CgDp7Ph3ooU5WBmjKKM5CSGr/0pfkjmefzZ7O/ADo9CH
ysMKFryzCD6k5CToKMX9gdD6BbkTP/rFOFOAk85vGXoP9HuFx3N7G3SK6UqvuqbSasTSAdR+tzND
Mr5mNFOvqDAXmTWw8KLUU1tbLvNC4wz9EZcc72O5BLopVKgFqyJBsWKGYygkJ/Pj5ShAZnIhUUsS
9Mbj2MXrFRqer5Rv3H0qtos7RWSD/toViukTFyFUS4Jv1rtQPRZXn0/qnfj4aqGUlLegLAUx9eDX
YFiyuWYPjkx2AKmUHZvQqfuE8XB3e1Ypd0idt31AnP5O1Qy3NpOUjcs9HgE/2eyfMTmBCqlDiwQb
PaQM85kDm+N7FYLaE0tFFLx5+o04EfIzjcqwuItYFJglNs1S9nfD0FhZwrUv6y23I14b72P9nG/M
xhmA4ELz4f1vVlGY8jeWRzqf5IHY1H2r5TnfiMgzTMoOYSj+SAVniQTF7G/+TvSQLBFbCzTA2GYI
T1vhJFApo7PYziGg8oUyEu5PYhsel3FyyUILumiBQNnneSXifyw6sfLkAxIhL+Qn6QYfG+YOWDOW
2VuEJjw5N0TZiGfowvOZ466bNXDvqa2qELVu6cIX6XGnzJeIx9humwJoSacXJcghfVNsTtLxTsyn
ieU59aU8eiT2NNzij7d4K7ZGP3mHRdOh/8ZxBZJ0Su+KqV+hFlhztvJUQUb35t0c94Ma7BmpVibm
lqfScyMBztEWuIR59cREz08ZEiP2dCkpEj6Cor8RsOHtRY32Rx7tD9p0npQNyZoWAmnF7VaPjytg
9USzf4yYWSDM7Ms7+5BvcazvlZdhfoVh2UIqX5pPH9j1swOBK8b8qdW1OXyr+ZXGpe4G1OuIPmS/
ZcLQkHmaR1AmLi+SA97CX1/kA7T1B8QKSN6DujornHe6v5jH17EXBiEUIbhWotXq/+9ELa4E28mS
4aOXh2p1NBqkHIFDZa7mW6I56SUPatX04cIl7s1bY6kzcm8pjNe+fdVUgAWHSyMxYuVAdsNhNdeI
2mucj+tpwvk9f9RAzLD8ViRpDWAtzCAuRIXTb7+ofHOieqoqCbVjgOBHqdL4ATH7ODxJIPKn33eM
5JweRMwzITThzEC/B++awGiQFpzUIKmQFF7C7YPnRE3aLH+RRzbGETKFM6WvB4CvNmwvRQcN13oM
T17IP5dzS4UpEbA8QRBEGAIKcMUaECVJ0u46ao57RTKxjstBvX04274nHrZP8/BSgq8EA3L2KU3+
pUZ6KIr7ggWbuKzTUlgQ1kZEA7uW2UFLguengkMj8kI/rggY2ZJH5NbVjcYbmVFOtHU2eiqsB8iA
h03hRbxDwQ0r+s4v/EaEOpukzmdxf2zbRPj6hEuBIxshJBfRV9yJrZsPhI7bBt88KPeRR1yBFcnh
VCwr2546HBFpT6WPp0HVYoWdlh09/WI9eeB7fKdtVR2utlGTKayP36EQLo9rlqOeeNrbikxucDmj
WrdFMW2Wi7ksbMXAfEoIhGavW0G7C3FTqymiuhGIrB1b7USLxL1mZHACoX0VdGX/IKH7Nxs3TSBc
rbFS/ZDaX4BFvKLSFkb2ccwS6ewsmehWcY779z2Oy7rbffhDwrt8q/2FPPWr5P0QO1hONheN4/gK
XYuMrjrvXuNoYy3m4Jb+dvfaABFi0vMFbR2MJ8KGgVK0tqKRhJZE2QjLiK846njxsQ7yKoZ/ShjF
tk+3oh3rYcW+nHvPfWskFeks4UQ2h58Uk1sxXTTJXa4JGKptUcRWzpMBb4G6qflvwCQiEsYLoJ7r
1IZJB+qFeqGU1VJKjv4+IflfYNlmzNgGMWB6E1E/tdkjoCH6C3AndynbWpft/nsmIWQbXT3j3pNx
aSocFWTx7BF7Qm2K3LOFDLWgBNHFaF3dPSVPeXJJpY/xzZ8TsQS3R3WwFFc1sW9ZN8T/bwMmgamN
ZzMOH4VRHiPsir3d65e1E5VqGo8RUZUX5Y85RTIH0uxEV6Jo+l0n76c8DCgqoZRnp7nA1RfccQde
kAjxXTllymJgeIfSBueCxOgA9k1najN21q9LphuDodV/20h9sRS5g7UIcPBijHvikDwQHftmuRwz
8l8yYrxmk/hoGhlgIVNE91iGMQrVeK44+imGWKnRbcrzVSLH6ZbfXC4SUSOuYcnZ71S6tJSJM2ey
SktjjugdsmQ7xXUjC/8iV28ZRfUXjRViw5AnKAfrlg82j0LWcNA2Ta8898+pklOLohoD50gp31v/
dUYdfaBrh3nyDCfzbfnfVYe2nj6gDtyP4xGyGrWuW4sa+7F3CJCiDyDAjKWuOAPGTQL+qIY4aoAQ
kCGgw2Y0ottA+o6W2ZDV6OjeR7OcyEwZiZEI2LKnUKRlk4YCi7Q9lhAI3k0LyJjA0qBEN82p6K1t
PEZaNGKqKdFPVo/Scf/k/rHM13p82iCG1vhuYcr2l7AWMCLYySpFw6ENee5q8WFADKnx/+HH82fD
/KqAsMt2wk4Gx3/EqxibejN8Km7LkNkr9ZMBPqMLoGXCK77O+XL5U3VS9HpvByzkotGjUa9caSiB
XdLfneURhNcVO6fbkyZG1wB75vsqpZf1MlTrlLs+uyDZQdyIwNsIcGwloFmvsy4f4UqlDoGoIgg2
9jws/AhQypyF5qKTX8nxPaUeAOqZhXkBssdrOOL1gVQJKdnt96ZKvzboqe0gI6rUUmt7Qk5odrrI
08GtEKwowJjQYxuGkgql8v9DHC0Rmu/FLoZA5L4qbDTOspyVL+mUNRiccsAmlWJMlrNpwOup0IK+
X3YbzAOTAfGNG5Hx6vkSaJT40zZH0almi2dZMsZaFjokJ3Yq6X2URxS079+Q8aqx4BQjonYA8J1i
mn+VUdxDHx3tcOBYwGI35CCe3IQN/3HACNcDeAgLz5xqUVHnjIx7S+EFH39LJRIPaYAma0X1sF4U
zBUXjS3hW9u6toxq+baiU032oDqxkvADjFZUxmZS4M1mXRLrHI5OA4bL3SdgfuZuW0RTvxIaYWjT
rqqAhBqcPoi2/kk+hj6irpJXnG5ELZX6OVA+v/Ctja7cu1RoA8mbvgrpj5UdbaFDrne2On5EMraA
JTqIhIYjeDABQA3Gl3lJFZK26hRK82iugVbFXJi+KzerYE3WTHfa4UHeNLHkVdzd/smSWpo7OSH0
BLvDf+tYy5k0yNVOBKEyjjtLb75lX9RNBYW4ADor3qIWDbjaTqohYzFVzkHx+/8DFJT6zmkBLq3T
iRJ5hoTew4Z1WrAdkfaUM1GSm0/upisI1IdbWm7fbjC+uAQ0o/1HSkOcy2fNPK+qHnaew0ZM9VHM
+d+b+zdeGolXqkOG83spgNSYEUdPmux/BI/QpwyHk1rHWfcXQ+QFqe+EiB2kfHZgN7cgZyRyjmCc
NiKIn4gs9g2s5LOtE5J6tvErU7VXulxUHjnH9pg1keFk17qy05wy4IhYue8zmrkRMUSgKaqILHp0
FyeJTuNNpKxOtSWupTMxjoS8WP2Dh7ZP0NZOIQhAUK6KWV2teM0zY6vSJtp/olz58qXvresECRMO
InQja8TSZN3gxCOYC9rcHFlka0KA93B574WkZ6MgJXrEBxlocIXM5vO0TTW1xSWr0Mj+DRo0TVYt
+H+BLkIyc8aUvecSEHSya5zJamxeOfupJ78YZ4sB6OAHuCZ2Nw4dTzp1bV8iU9+w3vpC17088gl7
7UPFygK+qgBcP+IdEgHiOM3qG7kbTtmToCcmS3diZr3FLYEP5GO+2NzBWRwQXSYyL1sOg2xof7OW
HEFvDXmNGHS6fshdF+eC2GBri9eMlNDsiM856qkmg6/+EWX7SPt2DVphXqIFnKbScEbl0pJ1koMG
SgUBZnquaegsI39+hxL4ROfwoq9tkfb9f2lakk3gJhJjFWwHyEQU6rZblfEq4L6suSsQ2d5+zPEF
C1Dfdo3PpieDWGw/kRXwC63yT9/jRf/m93kjgYjEhSXy3+70aCg0cgitNn0korDxOUaSxDQVKYmJ
xKksknmcSQh6wqajNlOWXhwu/EcP1eFpm4rHyOHex+hMRODPTHr9s3H7qrVZ2J+gt/7dE60Vqb/f
Y8Gia4iuqlhl1LKw0t8US359egBrDjBI5vZ2UZ95QBWkXK0LTb1NbLBl9yoYt2HZCxOxr0ynRctQ
bjtVj87OB2sa1DWrnnqgJ1OPGtmSLRAPJPm/KQPQZFufcVyDw34fzv6QYHh327B/mJjUDrz217e5
FmQYiFv643dDJPHjiUTSDw50ZWyxdys/zVIyv6sBbubWm1Q4MIcv1DHrDrMH88O6C8ZHkx47Uq8z
ZuuTn5gWRnvNApN1BAg/PxCFOcN9oYev4oyfcBPyci+fcXJj0etl3mbDXBYujPUaFZtSN2jwj2/J
vLhEdYUE6kQVo+6QUhOrvZ3IDlzSgph8x6e6CMtDF5R1L04dMu2nz6fU3UJc0TMjMxwuEQ5Lp/Rh
/u8Jz0X7wUtzyahzuSDeffKjvc6JS6T5Q1he1xz3tKtmvq06+3enqn6is6Cd3unLBjw5yq5sad11
GiMSKXjdnGGNN3+xkCL1BOgVEmtS3xoJJ0kdybJKYWDyIGjeaosLRDv/7DlloidmMLQEGB8Gh4lZ
O/UIQHCidopwApcIFpPPrfOphglLw9BfK/uoQKFb3nnFUqG9REKsl8gDFhwd2C4pW7DcmIGFgPa4
/+pCk6RDHWMnX+Mjw0YiU0LCag726RFBkYdcMaqwKvL011S5g9r2NoTicPa7lr+F+Rw2VzDpctM/
qczw6J5HpKJKraACZiuqnvglMIqhZPMAnnqHgN5QRzSCh+Lk1KmQNkeI4cyFqAvdxpdOeQNp3+6t
KKPAvjerh19ytYiT0t63a24F/FPS3wva2TCmOIs/+/2voEHTv0ZUMJ8RrciesMn4LqBUO9p97+QU
xRTgWOJMRzRVV2Gb13F/XbMOEn5+Y1mJfBxFpUug/jC4Mu4IpJ4QVer8q8Tt951HolBth1XgMUl9
OfPU0saISFlV//IHUpclzcqu5Fez3jUFMbe/Nz5X6RBvksEVs/fnnEQrpJLrXXUHIrEk+rkD3MyH
RKInsMtTxxUscNHpnQPTzc54qbLELBrndJHYSMdE/QHRzpNze360FMmxhgHPym6ugMPP8Ml1FH9w
RYtt4rdPO84SZjmxrXQ+lfIm4d1Zyof41SAzNLf0yfu2R03baVRdGZzt1JbNG+z0Bap2ZEz7iWY6
vU29i3JvHkNeD3F9+9a6hE7Kryy6KkIyjJBpNYyQghzxbEkgKURWGFJ4pOCkPZ1FBEfOUnv+DBQE
Sr9+eoVe5a6slHs5z+9EX+ecVLJcPoLl3UPm+D+StYv3T/q39dr6RolWPYxgCBbI/CLEfUamJa64
SA134E6K/9rWldgDTP2uRGxtMCnYGt6P9HHX4WHRZxA8FZHlLQWHzQ7PgNpxhxoTjbON+OSegJT3
QRV5vl4/9F2/lFxEZujwRQdRoUVPdYZgSu89tFyU0n7aEOBBSd8S2UOahTZmK077CP4s7hWIBgdv
7LkVyEWThV9Sidad71CrkZvdAzbchQ2IJQE/LOh4qigVtNasc/EFLWiLl0xH+XEn9ep9e6lBcY4n
KBNgyQcUDoVftEYs2abbgvEZQZFOaflOlDzqZ0d1fhvvHOgn3kM3TT+Mp0y07lu6PpKP1CX/N2dJ
j1PHUFImIu+ppc9db15nNdK++8gVPaT/PdBH3ugOUFjZZf3uaUAsZe86vUk1EOsCeNZlQv0gt3kf
aCRVT+rbwV6EK/DKYvEgzh8XYLxDW/qM4y9gwjmv+i575lhVmOTjUXJt5jyMv7+PQRmPy4ngu5H/
m/Ayxz3Vui7lsbI9LMiDHXf/tZM1uyFUg+AXjm3Gfv7BVIq1KwMVElPCSqB+8fsARx8kDZFDt5X/
cqhSLj5xXdUqwQYReMMC4BdtrJshIkjZ9x3WrA6txbV8eZu+0BisZTdEnQue+jY9faeVD3fmaovh
X2e18yaOezHHY2IUJpyiagHP91MKqaA3SqBf0z+dWIscKvq7Cc/oaxbIpPYAOnLlK35JlubVnEDJ
hGPwbAcIlQQzA64Sit8YZDdnVPnNEvHhhci4CerpLTyNZ+uWNHG1DpAEjR7kHKdHLoEQ8nbFGdIP
p2SFz88lbUxMtXE6qxQX+zkgvJVMQmxKXZamBlJh6APyv+QC4a8FgiXG8d13TlKFcLINHsyEfhM9
gmPIqn+74fSFX7pq/cvZltY2s73pkVDlNl/obGhNaOZiEwhzOaUa2fxUTw+NLERLpVzFg9s1aJQu
qYghO3w6eBcFmfJht06WtVEvEY3M/ItSzksKPXXGrCe9XA/GUEbghsttt75zayJSnFJURHGx8v0W
W0etXtL9HXdK+h+d0n2s7nS92Tc6HjypI09T+kxDASBWw+EDlFcZuLTngtNQRgUEZ59q2ZBMKTSy
2KTMaMN+77zXOkruTn/KkzqnUYZ3ckBel8j9taixbGbJLNYvvPouatCmVU8WtRedAfJiEnBQQL0Y
X3H8LhuAiz0ykvKHbuiBoVUW19emduZxpTaPjkBA53jCYVHEfBHUs47jvCSq+bv/QEmNZ8yy4Y5L
zNSCLdvbuGld619yG7jUAiWv2zdNCaSzDIZ/XNsEO3WO0pEez8HQrcpTSOQ9Luh/ED3nsiQDLieV
mQLodDmAqW7iKlsE0YnuCUqejxeYsVc+/HCXk7Q+dSzPmtyy4AWMBbj4/Zhj3ZblIbZHX/KQiQse
j+5yGiiskqvNcPzY3titjueuUaIfWIhinSZj5m5Z0FOJn3kkXLqkifqJYTfDrLwR/Kl1xnT7qBG3
IIHbLdtCT/cRFLJ1bfZqyFh1tIP/bTtTrPcxW2g5K7QrLpK5debFobliNh1smESyk96TBVngVORj
SI7nNslzgmexQf6owB6XWtlC28T2AZEN2LVVT/SfUznGifKTjk1FqH5pBJ4xuKGht9RayiChW/ND
xWylFsRzbTQ5cA6dLCo7mYK1sDqP0A14IyIQZ7rLmH6a84Dj9v7QPyrey9ZO/e0v8iclbwxVXAku
+7yhb9opL7Fqwe4KiWDV0vzAvVmzmeEFi37pcxEmCSL2hsf+Kgz/EPqXthRh7W+GRhuhye6MNBL0
LMYGouNcJTPJKNcf4kjs5gc0gAdMuCijkikqsptQllj56Ed2e87u/ieWmUvixP5SO0sMjHBYTvXS
D5FNjFgELAVZe6WCVlBQ861ey3A07AO2KjsfS3wl8gU6V2f+n7/aKiUOffXHAbdenMrblq+nE9Ug
VUX+egZ7V84bi2Z8+5kV3bCsYrCmT8a8ehAYsQ9zOANHryEmVjUAidMbGUO4Hj4wc3+c5s+rFx2v
hFSzSiTKhPeS1ejAMoMM1TXcmmLEpIxFoczu+OqeF8PAAZuppM7YTWQXLsZH76n3Qkg+iZEpgUC9
f0SKC1QFOzH57e+I5JO8nNeytvkYbC9cweoKvrTuTjo6KZIaxONrrSDOZv7wFwoIxSSl0px1MBRf
p7PtnQNLmSQk03T5cGajAqF6JBZgfssgN6isZUbdtIxS0MJdopMLqKbNQWVoBsldUOMhMLwIiq9N
xyZnlKTdHqO2X/fuZ3V6HrM/7NPCIov2Knql02nk6EntHHvqwUuTr6ITTx0JNsiCh+EF3V0mgy9t
1qKIXoBWj26hnJfkHYJwUEc8nwImjrE8N9hcP8IPPGSRHaA887ExqctybZz+ixlehDNyJglR+EES
teCwYMHmO99+wUqu6Hhbc0MwagUCkVyPxwhVhFukRyIpzNLIZFOLVJRU6wNxLMcNK8/AX2D3rL7t
vY2nfcwsJJgtqn8bTpSFT0Do2Li9og28Z/hYq70LxqR43IYmQ3qDJrOHri0/jFZKvLI8pDsWsraj
2Th/HhIwgJjcjdyIr90O7N3ci/Dzl2gQ5bwsl8QF7rYT7yogSf3WLTs8LpoIsa5Ztj6rmrsCB8XR
iLwZBZYwYY/ZHXhHWL0jcSL9TmOCmrtmgk82LSSM0wA26nbIrSjV9/tWyEDOqi+q6Zn8HDptbdnj
JDIZKI3LXaNGBR4K5nBe3h2+LGE6kEh5uxVgI4Y+gT8u1AGTw7TfSkplBbagN/e1Z8lb7441CMTC
n/UYqd8n/sZlqF+NJ5WQn9ikOsVrzFNk1j12rjiFKPJ/TGbc7ItqTVwpVfTx5LQjN888ooeAbkNU
d/R+OhnWZUa1ijb4uLVNh0ZGceadfzAezW598iOgj+jNY6imwwCpwGfcq7JpIWyNbozMIifBzeT3
by8GWw00L0FIFoHXaQ2f5bNovTkFkV5M/cYXBlt/hASv1u/c4F7J10E9h5v+21+t9OTTxEXnBEI2
bVK1gMhwkftwn6A53bMtEqjp6FLASMxy8lfokTokdQ9GknChaWSGpoaWtk4Rv/P1E/M6ai/WmWdQ
6JMwdf86GabUP2H8skVooWbNR9Zks9t129PPEHHabP21eGr7DSuxbmsEBpuDWwaSfoz966sw3zS6
7nZC9GcTH+AkLvM0fzlGhV5tLsqSw0t0UqXVIHz1tKVTviaArnyPqt463aeISyD5CRKT2CTN6FBb
z8SZzjc9s+gQSVT/k5ckhWExRi7Je4rpE0zuvd3L2V6KTNcBRDfu1HZZ4GMdvlAAlOBqpDsoMWEg
UJ8T9qmFU6+HO2izk9v5+W18BwS+0UI4VbNtPYLGmbaOQdbfeNXCS8QlIa+VuwLwfmhYmyqQ/Bs9
D3bWAvBiy71XE2N4mJn03vdOhUB/PeHVNfo+eF4Wgqbp6ou9DCgkAsIclTuHuvXN9zy/hHkZe951
WC4KUfVbzSvZJFGpc4ISJ5ftZ17ahLAmf+C/ORj+LyZUBeX6iLVudGehdpkWTd7WMgov4uNxC2xD
AMxVOdaB55oRRrAqK3qSZXJTHp07hKgOTVu3xS23oK+sIjhkvjuretdCMboRnajqq605sDEsVGDt
bTpwF+ucbF4O0mJdDtajitBxsT8Aap5amVjaYqq9cixCkCtnRVItj3d807fP/dHViKjEjmfaewuY
lR2Uxi8dJ9eCWH9yBnVHMIGKIvLUBPWIR8eoUdgfVZIPIl4Xt/szABdTjkWMHytlGUXF6broa4W9
PHkL56xvjzQd+QkPSOUkGIkegVDh0sBWx1Oag4Mb8A0ypgnytIIM7FYCoCDL23yxaqGaYC4V76uh
ZBUXCMavWAb5wn5EObKiLWaq8g4iFHma/b3W7+fsZhSykWz5hFf4+o2edwhJj86QLaBOCdu8irLB
FMyzrbcFPcy+K9xdFXOWk15JMRXkyU6mElzoVpS7VynWf/Gk44umFBJXNgEsAjXIk1dP62S+uw1g
BFfZ7dyAwwaelyGAZqyO3pUGwN3H1answDyj4VVvMg0lwHA6iMgug56JBUfRFBYwVpsB21rB0+CY
RgIP9YVP36kLAoQf1BpEblEP+P4ZF7R3qObuCqh+1V5Eju41MOGidp79S0R5G/wCFVam45vji05m
hj2DOnpmBXu+Asx8GdTXpl4H0/sTw0x+4XR73JXMRi77/Gw0spHVORNWNIsbU+czx7sljp4bvBgD
2iVSs+Pin8YFALH/8ZB7umem+/t4eGoh2lz7VFy2wfXwZdouAnIO1JdYaD0QJ1uWJ9nCz8xIKHX+
/YS4D2vbXejbnQqvGJRMFxDOfMIby5TGsuzuLQFy8N5e/lyVTbSclv14I/ho9c02aEii4c+qo/jE
LFnDfb453ArT9V8FggHNe3OksxamrzatG72ZXHqhZ1oWcMMaBUXFoYLgZZ6TpZszLyZG7sRWjRU5
nNyBHFJNnvxZcdvlhniADIckZPkKLa3ZyvShYj/8Bq1Tlu9uy1EWBMvqZN7J9PQpCVLTJbEXdBgw
fppSNAdgKl94v2iSpGrDF3CCp+VoCK2drSp8Pb5mj6Gy4y/fRBkMOGOPLT3TCRQSrayuXvBKNHN3
10yvYxza0DxBFrNENF53fDBy8xC78VNwi0Kx1uck4Oo7iSUkjmANRUHLQxYZ2IqWIw1Fja50sa4F
8iTiOD/WoEjn3UMBcSNH12b5Z0zIlGPhdNDH5u06L0cnHop6FaNIA0wcTrFKDZ7nEpM4ZEat3wCQ
u0JMUKd417DVBERslD1v+KuluIrSh4MRi/z8x0nZ3DutO3roZa88FHRO6LGhLQAQI/+cGF3gghbd
s+ZufoI0pEYUM/BI5uJNpVtcLQCOg3p4skgS0/higTkSboUk4IWYswFnjracPxYPF2M8sVR0POWr
9/9yAROIdTHKup0996qSUDfMGkpL/TfYQEiLC5zLwqZbm3ouWIgigrygVPy9JlTEb2kqEqIyJ96E
UGj7xrOG7VrRVyhzdnDj2aSSKCBrmEK61usBWuuSHiYck+17bpBRokDOpFHqQrHg+9cxUG5k0xi4
2QbL+Zg79Fbql/FyxPTiW63x2f4Gyf36srcFQRDLb220p77T8trVTmK0HPoD8eIjd8pqJZu62Qo1
paCT2+KBaW561h5SIIGNEDTz3IvM9BYGonh+oaaTTdvF8AiXyqXLD3pWfsOckT8WK8D3geDosgFf
9pLZuftT9xmbRRx10EBSrH7a3sovppx8SmRxvY6QXTtgaOXaQ7iJ/zJ/PL05AgT5ct2omXAapcvT
ZdQ1gyKRNuJkCGZDb1eOBsLt5nq63e+vC/JJhUMbVRyzKvk8sQCsdG9rBnKPl91Lqe1W81Oc7Dey
4ihnS56XqkwtDT0it27YnhOhzfUB/8ykbhsoK+Bm4hOIqkcG6z0ER/Xe/b021ObKq35kYaNAkZCC
Zzgx8SpP0MjP4Mp17o/F3IBxOnTyniFym8f/ZzN3WOGg/Xf30YRsFm+/80olHFH/EfwWom4O1F8H
f+Tjoz8E41oTeRWiMz0AuXgdxG3txRXhzwEopyyGkGDjlkdSZ0KbgiBLZZEft+mvaXb5DdI8QABl
GF4914/zXYXEA/OlYDjLySabmvh7ZYgDW73Ff/SlzPgSJGNGTWGTg5Yf3mJH8uahymg1RCea6jiF
Gn9Gql+Gv+/OcQzxLB+lNZ6LxacfMGLwwE/d6eCj+ugiXQgTB1DB+nxsS3T0RFvy8QNf3uLM0Nc/
dSLjQ1F1TgqAO4MKgaothgGiwOAzGlrWzsr2QK/Sgk0gCzrH/aJbJyc53mdfqLIqGOAx7aI4Bqz5
efg4sHPUlGKCiFGidGdNctuDLp+aG4NNGn41exwLttmA//9IUtPk3JJ5ejvJwY4Hm6xD/8xltpgK
NquIRYcx6QMi7k6L3rVdGr/C3K/qCsTz0CjG7a+N0XZBNnlxoy2CvHPwTamF9eIae3o3jJZEXfxm
W/jTidNDwgoto3gfPVutFlD+GwheCI2Hn2m0oSpKPPm1aBX7kEw6y6/xUoIV8kf9ktKatc9PvHC6
/rJcIn/A1PTHacH4QMKE8j+Ss/YBzOKGNkIg/V9XtHMoiumQb18BGMSVE060Hsh8+NmkpgtMLqKN
5y8AX6FYwHnDvZvZHv/r7NgxIqjNmz/imZmmzLI6oDxi0KAoeScA6jm1c6zDmlSn4HC/T1tTy8Vt
w9nMtPzitXk2IG6Id4E0GPD3jmOJMYXqXRFAfxngiNWutGkvwDq884NjxxhTRfNS6p63OPuYuSJ3
MaE73bivhcPZ/7Dk55ooLWvHLx6f5Fg583SfiHqfc1vbE5u+Vh/8SUAP0nxRG+v0pk29AWgOjkPU
IKFsG9zmQLhOYLdIMUXjsPjKs/pkg/1f459JQUHM6/rzvVRa+31zcqi9L6UHqNb8fF2yenyNPjjF
D8ShCuDecpPl1txFlT4b+sQ+Z8BH8HUIBJEHcFMeImIEUbibUAozlslQ8Zq0fj6vjX19mOUMv4qu
m91G+OJl74vD5xsrhhWH06b02NZZ/BfEfbdasEeTmwjG+ziGkrRoklx7x9AbJ56xzpkYEplmDoJG
9XWhkrdwQLVehvcqR0HXMyuHPovZD0SHTMfaFd3IIvGtBqIT04QiM7wEThrwxXEJa6QHcuM2MHPE
kV1CTKWCLB79CanJmg41KDo4DIsGPRmelwSBCadDv3IXhi6brmsAjW4zuKXi6vPKjdE93QgYxYwl
GEcCU3rHjfbLBHq0zGfD+itCf53mbbhYxt8N/DQ876/CTtpq+u0EOgjiJP0G9C9X/nScHwWlYCXB
D8RzCwrvFvY23mS59C/sg0l9fNWZsLpxv9BNoosz7AqUr7Mmo4ep4nsn9U/563IpmX02I2Q03rHs
qdPHZ+g3gvCjIMrh+2Fwh4q2xvrFQTlIMH438ZbYevSGie1lZ/6xqo06x8qK6IZfYRGYeGWUV0NW
6jcqHTb6iHJzrm0E3rfYgYN+cOAJGANejKA1BMxyhC9mgDIHhEr67asa7lEvOAVT159Mktb0vDDs
BtXUEaR2ov9C9hHr5POIesq1UGgmYu+hBWnWXBu5KSzU/vZ02dy+U8LFQcZhe+7uGBZtLuGzSZNC
sqpLDORVlejCPnsuwHgNhfOzVocwbrF2RHI7iwY2KRZ4x+fXFo16II5u0rokwBOqBQ3fSL+Il4hG
wh3Tqv3r38+nfLuoHJmOgBlFioN6zGKzmNVOchYPMkrPCxdsIp0imM/gEJp8eEz58IeLy20HBomH
NBxzmbURsx1a1AyhGqTSJwf5rbQpFPZs5qQtFTdp2wEJ0WXh2N7Gr15eSRMSyxwJS5K/5e2oXH0Z
2boQujqXDk7S7pBWseWYNNUYbWuvDC+4du45SSJG/jA8Eujy10VgMBIXCW7aT2HPCWp5NzWYHnqF
BQRT1ubA+n7txSyOHsx5c5scgqcTA1HHmfC1O1PPn9htjtnyAQ8D0IjzbxUPtgsfia9YIevRIAsR
7C1v39H3+02kGU2ohjUgrOCcKll8DoINdr/L/ORWm/5jKjDSf0ZPtR6JHy16rvFtqP0vEPe99G5g
8W9vWh4Xvot9d5xhvxUtEBOmuSnfhqu6f/PL4BfgCdInhUvdTN3VwW9bvDDEsZoahgWAIqNt0EYL
5j1oz46wTL3yXe1w3PfuPqzPnEMgZFSbKlRR14FVgyw2wz7nalnWFxMER1ih2FzaIYLV5yFQGMkJ
AIP/UyffMqOJ4RAQ5FaDfbQFyXLpEkBZDSF+CoqQQvHWDJl4MeVfG8RYmFRNQPVUu6AEpNqaBvvT
yaDqIWgL/jLz/Py997mLTWo9sRE9wCuurYBz15VcVoTcErgsQUD9waEqkh47PXknLGoy1uXt69F1
VMOPbKavKxoRch3qyWcy+UeFo6zIB4C4JE/r3UNVUgms87CdhlFUsR6ZW03DukNRNkhMKY38bMYr
N4cJMQokNGR6CLgIJ12ELMno3QVeIMk7XvYKIl8K+5SM/rIVH21JQ81UNtwunLMX0RzW1rs+oC8L
DVl5uiJm8ystF74YknGruVAvnB27SYAdqItgLR63mtlkBkeWsX9/s6XIxutet6mwa6BCos8+0Hby
seihF4TxnL7cBVa0DAS22KhGCi9w9aIvl7gtrIDlOkmQsPYVlCM8HbwiAnoAIfpgRG0Uqgaoha4Z
jpV203yZhBYdUI1h0uXgplyQ0d3WLCuS80HIdBBFeR6XR0x+uWV7a4ADSEar8suWz5I8RFiYLmAS
wmd6g01IehEZRr+FXsdomV0ZVksl3LgOYdmyBNcrYCEczXDuFx02oz1YF50OhdVqvgaJqfJ/KV7z
XnwfOSZS+jP9pP+D8lt7RgypayHpznw8r1HQKQlhaai9KRPhDpvJapZeoITgZzper+tWLYokKtaQ
ibeF6mvlFveEyX22cV8Up+w5XWDN72xSGxOVLSK2YYpniNBMH2pP31z5q0Vd4czyxEUCSt4H7XJi
BIG2Mywr72Zu8CrnIh4O+/0f5EcNpqjUPTwEVBqsjHfE7Meo5qCEJ6juIjLFjo0AsenIAtc//JjK
H6dw6mQ8yTq8wdNHL2eJlRJcrWnmK1Giy4rox8nUVnvKX/YmPAAU0RmqyJk8ZWbbW4FogfaSxjcW
v2j1t2vWY+ysi9ULr6BawuyZWG4ncxe3FVVLoTbQFb/OLAbZTbHvkDCA4kQo+brYYUZULIwiumZc
qj3W4BLyQ2iz0a0C/ArRHu7Ta7t7Z+RlLy9YrS5uNizDDjhubLg4Q1dPuC8Bwi4a4hDn4ClsvQY9
udLyXq58/1MsL+dPRs/sYiBLSUe5XTzZh0fMEdpAp2uKV7CohHPMPGWRpc5sJDO9muZsUescdNCU
qV3tgffEcvhMbkHXCr3TyNvTitYTGvmcohU08UeDV/rcQHUpUsglLX5rMRpGQRDlbre+nN5gkw44
12OAcrhdyjj1eXF1YdChOYixu3vxKs/fmpVQAk+B2gzX82onH/5juFysP4/0ZsNLBNvXeZdgayY4
He3HiqEhYPFLgeZm3beDXFXppewbTDpexuzfZAxhVZyi5UbqDpv+IiqUyNbbXLcwedWbiJ+0aB8v
BeJtZkT00BKFzHpd60GflNLNzv38Y95wp8YCpdAoJmY6AzIsUJUQZrBVUyLKfMc7zSQVUYD2bex4
FyoViOMv3LgkHxwVx3Rrkw99dQaZag3JMoklmXq415Efg7PVQI9u2Im2qfjCI8gPqVnpgKvm7UtI
WrMNFEyF4+nDAYugSntpTympv0k0taLl2cKf+IKgtTayD0EA5atpAXqL51NnxQEbHEntjONLSdDz
bu/13q/6N73TA2+qfspISl83+ws3dTo7g7yPtgmTSX6TEvWTWXiMwsNgHGwlw+aVg4FYYDtGY+dw
1Vf+u5n6tLvRbDK7xGu4IsRsOuiolTfEjLjVvgwA/8VAi5iGLkCF0aAmDzZV2RDp8WclNsdBxZkJ
XgmXCXIIOD0TwPrpy+k97m5EgODKHxKActSdeMmfm3+F8XnQQ2vULkEmXKa16zZLB9zNLv/S4BxP
fQP27+jSsR7/x1bFmsI/oB+hLqWXZLDskEPrT4XS86hVCMWoqzXnQcG4489hVL+bcYoPwlhfiwcC
xC+MP6fr0WQysGZK4tJXZQxRkR4Es4NkImCicomj8cCowtg8z99reHalRvPSOHRh41JdvhLgucqz
VbEuFYGIhhEH/6EqcCmOIFsASfg95eZmeHxvAjZo/R+nkDloa+tAzFM4ecK/RRfUPE1/DgFqX69h
jH2LCWCm8P+c8+6A5sDmq6iiaR7/5VygXk+jkn0G/v8v9gveNQjGM2+6ysf4neo03UBQu9n+npDg
FTm2FtLAqiaSfm5PWKbAPQ0y16twq5ct8XvUf8Shxs8BtgbIJHJSg/EYT23SRLUFS1P61Q4CO+kg
NSBkCWQ4Gn9bG2OajAYGcAjHWK5WyW6ICCb9BMM4rHVkNTbel2TNpuEqlsyLb+hyC/erEMU5RI7t
ZkAhRO9kW4xwi1g1uuEuCnrpa/VJGqAbB4t4pQ4g+yFzlCR5vNvzl8dzFns1xow/4q2hZvB5gBMK
tw0DgcUMDbNQ91V0TX+HZCka5fg/PCAlgxFTo9GIiTgrRGm1B9ansNIUoOuI/0i5rVRWxKI60GfR
tT1E+cD01Rf0VlakgDnEUjtL6TkUu9iwyQWgDArmevMNiHvN0vcb4fI5RL5MSGjhdvw/Fyq8N15o
Za7mix31nqIkIH0uJnTlJ3HtTkMyDm2UHpByvumeYcH2eB7azhsWtq+ESAKvlinA5f77Ru/KE4iV
nnVSVM1E6KjpC3xFojNrTF9XKq8AARDD2+xVkEvZhfz0aXA4baohqywAdxYju50T777bzZM8r7Lz
Si6N4iHbygm+hoEwHOu9zD5jfJmIvD1ZEMRXqr7I0ChYfDlJKWBnBPkKjDvWpnaZkB72flXfQik9
3nZPh7qsgEGIFiySJCnX5DHRUqG30MbQIdSH0raZeC81EMi5jWqnoNPSOd76p/jnADc+2YgJui9z
ZrWeLt9ZjIp8W4B5gOs/aYpPgIQl8Xjpg15QKkwqKyneGp8P2AvD01C6DZ72ufUayvqIBZ/XMdgl
Lb7W353rAUte+FozaOxkEpCCPlBQi/e9gMcL4B8QrJrisjY9fnsfulyKb1aPCGNYIUVlxZS/+quU
NzZGv0NeBixpIXD7Oh4Uxbl1KUzrR+jOWKsgOHMEq5WRz+HkT3YEd46qHN2XK8seGK9icETn/lC7
kDKWTDDvibkkYqHAp5PLDuGZh1zWsgf7E/lfQasWVd6yCQWfLSpS7ADfPVp9GbSA1Ox8IGu5r9uJ
zwl8OFfaRQJ6BP9FrteaF0bBG50WJVe0nvehF9HHaI2FR3xAs8GxcmrI4kjnYTU5czo3/S9ivKk5
QA0m9zvTDYDmgpnemmQNmeqGfw8Nspj6E2BJEE/C0nrSVwOFPHCYTSZr8sx2bDHp4IOO34tAaJ+9
uEqb7I2xEutIQR+iUF4WHk8bMi4vWzQjcYnVMlUZhGIol/t7bbSRXb2JPrUYkw6WmMjOJzg7oMtN
WtbblbBiZQavLqiNYRWBvPXzCcHLhEJ1S7c74H8fZIV270fgp+8ij8pGC0//NE5qyqe9hAAVHSg0
NohjrNoe6LMnBEuGpYD4OhQ6yetSMnoo7ZH3E08HqsYCbm4fFVCfRH4R7P/U6QluErauHVDaWOYz
ltkGscI7nIbJ7DjlYCAqtb4SB6hEOku1p5IjzoPxUEPUAWpJedWrQmRow4GE82ZrTkppzt4nHd7G
NXNKdyTpYKpDikNaGwe50VkL+s/oqk4HYV+x3JfZ3u0yWSvD0FFBZ3idXt/cPtRq/MjCW1AJPHNU
ZQNu4bh2PXJGYDx5yPEzGYHoKswYHQIsKOdH79gYdma5FPAfZB/G6kmtXqOAfg/zqVURCH+pXK+i
UF9utYxH/0UY6lvPv3U3kV+VPTpkeoiXka0VBvW0ZoF7qV3b5agAd3tWukXSrIBeHfasLqdt0sJD
m57DdsZDhZYXAyZAz5LMuM9KoGJRU5Kwx1Gl1mVtupwZfCZwA8Fiy81OJ/u22y/xg1xYNaPB+qt9
rJLKnBOhmaiuw5iZmjmYrrEqO/+vSgKvMHevG1Wyi/WWQ3DFOj/EcrMAyZhjzTHAD19ByD5rgzPI
ejrJFm/Ozpnpt/1xayYreP38o4ah5/j7E/hUA5v4vXhvqkc8x56Y1oqp98LGTCWKyQCCAF50NA6B
4FzGqEyyVOEdL5PDDx0nF3A0FY183O7VZG1qS1S1EbrJ7W7Oy+omI7hcMDjVgxWS+UpydILw91fH
GomWHM6FtjybehClZlDTy9opykYAoA8o11cEgr8ldq2ZgoUx/N+k5ig6ErobMsORB4QQ6lj3CIbb
zIY1GlHM1jWx5nQQpsYZaNQd+oe5wRxRT826Xqdi3Cg0D88ufkbansOfnEOA1B0+XwP4xZ2AGacF
wk8F+fiUkBNPFZfraQs8Y+UCEMAI6F4JY6B1RWwPul+pHyeQj0NTTWuONP+2+zPnAdB9Wsy8pRgW
p2NP3+3G2vMxHiBepYCb6VLSom8DJFBTLCPKD1q85ArynTc2Ac7o4kWxl6BwtGFs6p2le9cRWAhC
KNNJ259eIyo//A1Pdhq116d0cfXTfTZbbw8+geLKd9/1mBaB1wEYou8zJ4OlgQwrDoc5o8V3VoVm
ZFT8rAZrPanTh6p0ifBmyDWtJ6vS4buyyh3fbEF6DwVhL5vvwYrVeGa6kUdxnu5p2b8dmCcvlZHA
DbY0DZZYA39yfq9vdYpdSt90lHye21U2r+iaBcc+uZ8q5JdCq/TQC4e9AvqwfxD/ITdSaRvDJXle
kz3vIHnqpUFMvNcMf2bK+dKUAbuvrjJh+r0w80CycTM7QqmkFOHq0LtCjIRlbCwblrktruPILkQr
TGbFc6DM2n8CQjd12ok5tjMTJAQa+NSo5MQkiTUc5KX9rmANbuNElBwnNLV5wZr099GtTm0wonIY
x6l/udQJnlVtyauDVmIVe0V3cVq3+Nl43QqIxRtvXTrGRftPhhpiL2Pz0wBBRBRrpExLpa0ZYoP0
bVv6ImNORlARrKXJz18juGYb3K+xR5rXOoRQyZHCBj69LPYkmJt35losmPhEuLSCRRLMSGordWda
QtpcJBLKL3WTtgA8g04ugdApkiz+pFBt2PCOt1TxR++vEB042nQiIh9wU7CF2ljv5l4Emy5WYN6Y
2jRe9I+2ef8uG8BjwpqzRquxm/+jplND1st/kXHntpYQbT4UNWUexDZNdFUQDFMTzmJeDlFDISGl
KaxxJ76/eZ2A5cCLripAQNcC2kC7ioODtQLTbAItBMATstaYkl1MRhEKuKOUtBMUsNfsdnExQq9p
Px8KiLheNzu5JFc48+iOyX2ghxWS6X9CttJzno8i1s2DEPHpyF+rkpr++VeQbCk9Zc2wWVRG931r
6HBJBlCoetPO0IlX6XQlnYhMA3WzpuOWj3mfFPnBqSVK2v3U+hDHFmi7B66jJ12cLl0qIrZ88kqo
3v+g3li7ubaWah+pPsydiOI1NQLBhUqI/imWSM2KrEEG3rY3hJl6hLWc6gGAJqJ3SwFhCivobX7E
mx5w/WYxv+Hz/OVIlOAkMnzX9+ROYHjLgKDgbKw4inhyHQKgAVaY5JaeRxhadjlfX1tXh7lcJ22B
wnj2AGPgH1byl5RQsHsbKnorUMoaW5xyATjA3VElcjBaTJ0Q/btzwHJxPEGygK6QhvVJHDDlmASF
zhwMpOO0e5Gq1aAYJgqQiNMI6KPuFjFVqp4OJVNWULvum84A+jTx6DS8LaSxmpWAZh+UgiL5YeLE
sVsCabEuc0RCfL7yRxJn6M1KXUXdVqazXO+a6AeTNoUpwaFf5HHSAxVTNrMI/IQ1OsRSlVxaxhnd
JBOXdJc26R/yM88CD9jKvXAAzUfjxkCy+3tvhsmVlDifkSbijMPlSGzoZhMZWa1Xyy8L3mj6KPHb
kP0oD8yXmsfmvtYCW9KFCc7PrJlBMErA4q+Jb3dbdYZLHnZY0mY4Z4g09oycKOrQ5/B6b8smgz1S
UEIsh3BUE9RItTYpj134Blu6tOZaE/oz91TpdvyxRYkCw9+56zlZcm5myNz9Oo/k+C/W4RB1d5qa
Oj7fLFOni621XpMmps80tRNXE/YeNsaK9dPwHwuCQlMqEHR65LrmUd3rwmQtWXsFccShWz5ZINDc
MpiBFpYIQ80HH0gwYsH8nHkNnAZj9ZADYPI0B6cTiaQ+yki/HO0to9IAeHJdqTVX/0iwP+rDd0jk
Hm5vw05c3oRMjiBMF/CqiyRxbJRzemV2/F3O6xWj8ToJW8pYOh6IJP4x42l/72BG3er6V611bo1p
ezEe80dTrR5uXUMurGV7iVEu0cemM4B0s5Iv4R+rvtuAhAc6R7P4AnZDqrp93kZxt3ewVi1cHn2H
iY0xgdxc34txq6yqWGCjPQMzO+d5hxgfEmqhvErESkFNjwBXpi5mwMd2aLSj3GmOnsCdanzavWP6
1hEgp2ruPvImfmmTCOBxVJxedHu01MU1g/Y2mlucTnj5MACESiKz/Bl2+sNxA2TsUxdZ9/x5r3qM
mfOlBZKneA2wG674czwpTRg9R7YCgMDNVliyjIeuRfFCF69FZIXji+freGRzLN2IUcz9Fw71WCD7
22r5DH2QJgExi0BHW+6lwRgwvZtCOPunvuvhalX32uswJS0qbYbYJk+CDE/jm+X+k+CYfb4luglF
OSYl/gVqdvgXM59oY62THu+bNLyVN3QGnuzihgCmhXbOX0pHDwiJibbUEFnZzxhvz5BNx9acHEju
LQ9OpQLvB1S9QrElYkc9IIw0n2o707TaXs4BBv4+MSpqSyJJRcZxJAxwk1uWE52529zuPIgYMhYH
OwITyHGrUNbuPBz6EBed3WJm2htWAVJjS4Wf+xfUO5skfBv3iO9NqY9F3lixcEl2hO9yjUuvASTW
fdvlKMuFMgPaxd9/tQYOfhySA/SjwnXG7pXdkG6wamZTN+Qehd9F0MtjJK3gctsTwEMrti6QlBx1
mSpgVMUQoDYG1yl7YMNrAB50hnye2M369ZYK9lwxmSHVrx3hutgLHHkbQJSXxDLcqPMCWMgOZR3h
RNWjJOLkNYMu6COnysphA4JT9NBQzYmwTnYwpa6iVsHW+HfdBJpRb9ZOOZQxVtFEOVWb02YYmJIb
pOJTuADTqksbznqhAX1IPi0za77rfwhHjLhGptq7Up+Z8vnsF3GX3Dy8GHVF2ABntX5dXc2QCsnP
3/5qy7aZ0nFr9+pQ2jL9jDO+DU0UxpluC0AH9mS6esPARVKuwCfuvURGrhck/LDxvTtFhhUDZ45B
pdx1OWWviSC4ZnC6J0zE7yRpHvx14f07T6qTiE680cV5tTiwQGq4Sbf+cfc5ywPq3dAT48z5Bto6
mCJyL9mSlNjSTEq7ChPVr6CnD0LHdhGYa9bwIdH2FyagZEYs3ib0/V8SUEjjYb3qGJp67HhlPR/S
6yctmMCjqRwBwycQUGFGzfH7tIWU9NfAM76f3ySlgpwzo/sIkHD5NArNb8x4yhq8kD9HOcRhWziQ
l/e9dJBTqpj1LpVGepw1+vKtW/j6UKwrNT60fZh3fq6ezlsM7BR06vxQX0Z9tve9HDUlOv/A8QDW
Ovi9NNW7ICdpVQiA406drEBYTOgxZKrC5KxbfKMGvluzbOG8y95sHWzbtyn5LP4pbRs0711kJ3/5
2nNkFR88hnFahpyhhqklSknPgdB/uhJU3y+1ny25AZRttxqrdUbktoS9VF20SWoEDzWYpHJGOvVa
fTc6AC4P6DUReRfOGWvBoYikM6hKA+GJNH7AYgM6SaVJASd7YcTSt+JjqMLYYysbpHkZE+kXsbPU
7hi+sFjNTM3ZPBJklBLeWew18xrNDFD+o53RJQ5N/yYGGwziw1Ju9qO/NWcMywv74nrbXrIOWWi1
bkCsf7GzfY/XS812SmL39cOKR+xXnDTGvKkJL/H105Qk7sNtODGznnD9Pzp8v2IzSCAJ73ODv2PF
W9+3pe/W9ZnuJM72m8PrmqzfFzoDYy1DQ+bl953CznP5abgcspcEo0zIwRalUXPgYPQ+GE/O0IYI
fq8cYj/gaEMJGkzQ+IeG+cxshdQrclvWYwuxJzQ+g+UKDeQYNRLCzg9kpxgc6ujzQf+ZOZ5VN79h
RG+CJ/5LtEDKMDuFFwVtoaxMcW6sWWqLoslaf6CxbXpWRQjECZP7/cLTRGshxGZccyht6AABTRHz
NZ9YqlUaKwjUUDODKrllatJ8YeTybbU7X2rP9pSKMzvqt1ge+Al8+0VnviaQhOeUZEI1tSiwjsp6
1+KFTLgKgaFPlRZuvQS8gUQ73BdEIKwAzs2B0ANE0MZ2QywcPeLySs030ObN8xmUlaaFo6JjswgX
7rWIvn3fFGjUCwcNfhL3QGaZ99IwYUdeqEmUHqsJxWqWJ6lqe6kVf4o2QG2apPx2SA/o/1KLOsHG
LcSBhijQInK1HJBX7DXuw+wDPVAiKB9lsg6hPPBUTH9wLxhiUSFjvTy5H72CF3qzVcXH+wVD2vwf
FjU9Ki2En6o93l34h52c3TH51a4/lePzyYTiNo1akCmYjjngM3vydJ1ZkZa5TzlF4zksRHsZTy8r
FcxicvH7lUoTbDG1uLWsYwG7YiN5rsaKNp21YO0UemKpfymmvrL4tKGnYYJ2uzh1ToJEA8wiQgfP
9m8NNYpt/fN8KnAvwOdIYHdkxFW6FpX/KXaZ3dxKH6BQoZLpIDXFt5oInYByFHbUO0GMbgtn22Ed
52AF2HdCeujYD27axg5El5/3SNJaFDbin7HjPXmKri77gKyEs1NkeAbXusEjoqjEk1ZLwntYzeo1
TZlpj2qKysfcEI0b0OoVWuqbVaozKAHPT/sUQdmvzbvi7H/F8eVkm66hY38sUq9dpInRm/rFADXt
8O1ysHm8pHv9TYtkI/QtHcF767bW+VgjSlG/JwtYbOP51bWZeaRR3kAZFCJTBEn/V0JeVXFmX+/R
NMO3gdN7WtFd5xVjZkqp/A/MmWtW2rEMU5JTxiqHfvPOJ8MrY54e80WjJRsSXFui7T9mFVigLTbQ
OaZG5+9QF69CMTya2Cn25X/TAoqFjnf8UMq5qEOCPsPQyzOe3QrCxOank69dASP/vKf9PcP2eXW+
Vnl5KeVwIqbjwvY02W69VqaU+N47W/KwxahG1xWlERPGoDKgQRbFlh5EYPRfyyqINrYnh18XoSYi
xdF8G524DX+5CPfWp7R28zhQyzMfP+YiXyE9T5DlYizQktiTpjb1ZKjOSyRQReMaPIdI6asEaY8m
oaIPU7kgkGlLjf5Chi8a+JOqNcQkWjihC24hzCt0csAy01UCLp6UEWxpJcJQo9+KvVxe8tSvDup3
QUH8azKsi8e3riaeM6AyUZh0o2JFblJXTnzMrWyiZ9wF6EoGgjmQRVcjDIaot1JC50wsifJd3WFO
06VgzqfyREnM3BVTULdSJho9l7F7gbroRWUulCkFs5afNWN7ackpLtoQcBHcZ0ID2aCCfQQb7UKd
5L+MdTecilb4xc3jUjxe4bYPhvA8j5SqChGexTptFjktnrBoTZxZLkc0sye005BDogxuQvOcGMzU
RqSJ1iCci4VcHW/Re6NwbVaz8j08Wzr0HPfFeFxTwsrwsbOo5XsDpssZXHLHKubeMK2qNeLx23qg
Z7brkLG6DgRaRfqPFn+XB772w+hC+5jHSSxJ6np3ATCkr9Flwyd2X3FkTdp7nLUMkJOP4i+9e6+A
Y73xSWm1N33lZNiR/Xqj79HpGi2UcpFay3TNjUkJ2USyda8OSqSPw+fmKm92fiQw/Wv3Z64NZdA6
t0lKniQK+vfnT83wbhDOAbofKKCyVh+7ltw6Y9pzs83m+Z6uoIEAeIgir0E5XC95QRfshSiTuLCD
9kvsrra3AOl6FJNBwvVO5rVjHe9XDqOycMa1OfoY5Fl4Wu3rsCpVBQoARlpayCZkZJCqnWlTalr7
A2orF9xsTUybP8EYjF0hZEWnjKcRNf73g/af3p/owvpyrlas7xh+RDltYWPBgPQHFoi6NKfwvPIn
yj9Z24WJ7Waf2yR3wWF7tKkUqksEMsjizk3wsRGW0EKdOSlOJYW8FZZEyZrmGlkCXID4f6u0N2bT
a21L93sML3i+148WeL6nBm8fsbxlWi0ggyoOfsaBhA6YAFGS3Nwg4hZ5E24IEsEejS5dHOA39B/Z
UpUSEQGxo+n6AOc9HbQ9X8ykKmEFMlQv5Ji1G6j5UTawZQKdMHCve6f2eocmR9LeMCADwQpQLNJV
6coCP/VOlpoPRqtOJW3V8FlNNg/6e/fxA91s2bXGsvJ0d+YFwHFYmvs29O6Qkc6colVe8Wba0NY0
cigAoSkUdl7Ph7oFzoQy9S577GcGNEVCWWhLmxW0+IOXiKa3+4Nh6X/3n7rIMHhrDop99x+pCdBP
A1pPvJIzRLi04/tcOkbAAD9kFnikzdQ0vI0v6EwIV7ZKtdesnASK+C905d2OUv8NiiRR2++Rwjq+
ivQxbbOJ2p71hKrptpb7y7l/wD0nf8eMloOqWJlBp3p9rm003m6xShCbtkXuA78DKUMVAPihCS+P
xEW4ygiyniTjNOMxtJMj7R+LyPn3UznGeh8+JEkpu1onLEPbluFBxlyuEowWrnWzE5n7gFfvSSLs
n5pFbzS8FICBGhDukytuB4NpXTRo1AdhCv6JOKCwsvRLmw82N0ddZN/90I3SvVFSue53znXr1x1U
AqiwHehPlNaTgBmnmIW7ak6uywXdkmTdMky03AFnuWHop5j6d9cHfWZBsrrQPPBMksxS+mpgSO9W
qaOizDqOM/vlmEAqo4vktM1FyXS0VHeCeXiOUwdas51tVL20QGUS9YuxQ/y6pjtpV4OOMhChXKgm
6bHEe8RvV5QbIJLJ9hnCMJjOeLMpNcfT8YpzsNtXdnQ+xUV0gAUGF+6YholSUWyDhDvfSvfeKH8O
i+gHY5sx6vsxLwNLRMWY3gN0Ic4YzbR7j7tnYbZEwXz4a1dNxPxXUO8LP5bbUbq0oSfWDd74AKHP
XfTyJsJHLn2i8bS72Yf5wXO1el9biLVgQBNiWx8DyRJUz1tv/es+f+mtsndr4gRYrMtZF6TtgOsA
T8TZ5VTGmbUWDNJLlU9TEA7Kp4eZPpI0Nu6uvzj+CUrMFT+TpbTmdLDcVQ/S9f35OKnNKKAROCqE
c/WFxuXJSWTp/c8LbVuuVu14v02UdT9guDCqVryu16FkfAMRnIhr1GWJuDGp0MzgZgT/YK711uC4
vlsgCJ+QkiTPHAMYO17R+aPTG7EcYAvCg751JhnBQH9ywJtVjxihsxQERImckVu7y0QWffbOLxQv
3pABU2suP4JXeZih+94dL4dumqRbG7Iz/hQ74VMaaMm2w/nwP57Mx8B6LwiFNSwN9U8HfqNIhgOG
pmyay0VCfnHBV8JqvbyCJrWesj7SyH9Z9/5W+lyBogMIZgd6BiD7+0X3tvPyDVXMOCScQyFi12nQ
OAuMhyusbxlM/cjxzpkwfOBZ/JWeZXOPWS7KHDj+0bwQnkrCQlzixolM4JabEBi/Hz9bHVd+YLB8
3J1y5ZEb1ujrjHZiWDG/HihLVifeOJ0FUomXP4OQx80f6zkabgSKNwc2zpALTve/tw5go08kegfM
llyDygSir+5g8U2VLPOZHm0cWA+P3hn2FVTxM5LfQR6VhSdBckYaPShoPwuCNkr5RjRpfqmqLsCj
dCZBNFiFnyV0nnDjT9Rs1nUj50ooKiPsmaQfnQHenjBlddfMTm+7B+my/LN9xzzxX/sNrXZi/CbE
4/s2cVcE+ZczgYGkl/IgximBe42Siul2fxqm+cF/D7GalKQezsSgW2w3oHLILbbVjY2NDQHjcSAX
8lPcGcjUrp8FTf2ax1W3xqHROw+KyTSM3/Q8vEWo67cT2tjlo1zcnpGTTZN7LGABAsIF3lbFxQII
+zEwenkAzagSkKSBmkNA/W3l7R7VSO5fT7J3EPcSrKypdu7QudUphLQvxmDzH/RajhYi5qCQa6rp
066Q83r8XEpSVvucd8mQicSe9f4MJuZ+4716/OjpUnFfKwD5BeYl6xJhJcB5GFSiNQzIL3v0P6z1
4wyMVsv8cKMbuQ5IGyfxoIlF9BdW6qPfiPE7NhrzuyGoLrBqaHTXDy3mL91SDHxOrhOwCdQZAX21
ruS7v/PWqxjRpXgbZy4lyjEucIGgHry8C8e5LSlqNo1K4PG4CKQBQ5OYrig5peyQxmyuHXm3k6G2
vhapXFrl1L78i41apsaLTvjXjRInUXgu7zarPxW4VuCSQMylo0vHexfjjjA+TqUWt8AJ8gs1jRH0
q4oEYShHJZ39idFwpPIClyee+I/+YwLPbtuhOoK1X4LNrTm7mUAb1DQlX8sIESaU9Cs7iYICmCbh
cKaIUiqA9QdqHGbQv1Z8pP29qER2fBvXZy5USBqqRxxp2G+7WL0+mrdmiDU55ZPDcWHAQczJcmgL
6aE+YSNheRoiUG+Frsx3HNfCN58N706JtAWkNbozFYceM4rYbULmnb1JnTICpzQqUMOO3xJW3ako
DiigHx8q5nEXHj8XZEvn4A0x02llV+bG01Bf5JKkqx2gA/EBlzF786/KS9vRdWweHc5fIXaJwSI/
7BSiSXMvX/UjqSd7mQOGluBIfVG+sP1qHrz04ySefvae7pji+LMf8fN5kgi+tIxAXZDxgyGu6PaH
SP4FRJ2KFkpR33VmgEmvQIAvuFTMtiCgGT2km/I+tlGVwxpWaW7bkNiZug30Yd6vjM5u5QGleNlu
IsBed6xOu3FWcYuB4Rpxf7zSk74iaChUcxSSh+vjY6778l05eZU2J4FsnpP6a9PTQAb0QIK19HIy
JrJvpNfpGMUO6Mah3p7x2GAIpolXaUqGTp0qUe1k7Ue6IBltBCNKbeu1sv1sTJblNXV7dFFe+t/+
85d5YULz3WlaybL0dBWCESecxfetwltx+KMk2D5teStuPH7HFLIAuVFMTewVwFfkKm8gaEsBpWA1
HQIjKQBD8Q6QIjGFzKGqdXBSNamtPLCVXIt7J2JRLPNCDF3e7aeiGOBKN2bgtaQJ2wma5HtsL96Z
9oiEUvGKoudRwrz3v3oftzjczYY3p+3UquyiD8UBTOn6WxTHVJHfPXcbPrJ2wBrjFt0DLL3ldncK
CMMl9jtDlZCVsUuFF8JXFP41IJg/XeI88EnKligLKCIDvDufSVqKHv6rsVYJc/wNoqY9/JcGFIkw
DDdcBPcDunZrBymdjYhoMTHGDrA6IJOZjKzUKnun+7mEx3VqfwxB64nP+Y8zqm5l+RyEEOF8AFpL
b+9qoH7+WWSjJBR3CtintTvEJzSY5MHKMx4PDyYhFhYwbyKX+9NMEAJkTBkwCIOC6xz/XZnS0QO9
qAyceGTp66vsZyFkKAXKKmbFsHlQGQnSbszOELnNwvvG7ihHdQbqTCRttrYyFDH+oDZKmUzHjWkg
NZzX5R1G9+Ckb4w8x/kze8CsffOiojZDCBaUX8luAYGHYw81x6FJmV1OpNg2YGmqNp76ce/sMXVg
//vkq7Eig2hKPFtkE24phIlmNWsvKYUcOEgBG/LVQDBg5e8/jOY6U5HitP3w0cwqnU/Js2QVOmUt
0QpOq0iNf8q3RjONsdb7/z+1MqjZVcWJYf/kpjZvuxK6pjLlDBmEOb3Yw1EnzMpAwZ/qJg23g5U+
A0ukq0MBR9XdFYju/YvBoRSUgcWtoW1yqF5LlIcgYOnZJMoqqni65Nbn+FUSeWBt+R9yfDeYLAWD
QLN/WG5/vFdp/JUEDN3mCdzKEh+WYyHJ6FEHRSldEURMuHe+3JZ8DU2bEDHTKUzI3/R+yycCzNno
l1yx/gtFWr5rOCCBb9Jc+UiSSOdULJUYtL66QHpEC6SdaTv0iro8i9sWYN7/6rja4vik+2hP64dW
9IOkHZQloRbHnp+fL2sfVx87gMF3II4Pcl0iOoz7KcVFYAV9hqVEkEb7E345o7uAqHREuF2IyTYW
/s2PTNcLNbcHnqlkHapoYzcda4ch0QKzmCJMFju7oA5BDxjSxVaYBtRD0WXgK3YGzaYW5Xf3p8SJ
nAkLnS0kglOM9hb+AJvRrtVJLdJSnAvY7lD6n1QTvqTO76CVbnpynXLCyUjhIV6alPN8jWykeUto
h/ElKzBoa0BlBcFTuivFKeXNEvz/3bB+H95Ra1pQr1j/k19QVJ+t5UTgqVoLMF6OzMIHkRKEWrGO
648nxttFXiq3UhGeB+1MV8lq0CkAyaMR9wkXCd+HiWHddvDzK/I3Z287HjQHW87LOTNS6ciEeA1/
8H5f7fVt8+XrpsnH+WIeJOebu5CtdUvnTcKsIDl7GtwjEWcrdSEy0QqPMb8OUu8lxPgueqHpqUpX
78U5j67J5AoNuRB/lg1TVOfLZwnFIIJrhRbA8wNhnCi+gNGGLipPLm0o+SAwktGaioGl2Qcz3Ay9
bqcmPqNQ5gUr2wjWd0WjHwAjXXtA2RlyZakCrtKp3KqIf9ARdyyEoJ5GgUz6AIAC1bz0M3mfZh9z
Phaf26SCyDFoeYtFCrtDhUX0muA4nUGHjVgMoxqmZ2JMBxXSbzzAd4fe8udUfUWS5aw572chtTWN
Hxv9ENl0Alw142bJzBdqdTITBUYp/PCuloIYyN29Iin2q1A1HFhRysdG0dLdTi+NZemyLBBkGt0F
NpPdjcYULAfoFcyo2kxqwRvDgg8Q794j82l0JD5JCGhTpDSN5GPVejhXUrjhNeVIHfzpDas+74TN
z0zFOtfl7iRjUUyKTzW7/aD2uc59FrilgOnGmXDAEVigpJK1G12xplvUp4hvUru7AbwAkNCA0ia/
AXnW/JMJiH0Yon31wBukJ1D9SZX9Jv/yAR/ZUcRBeul/9JCcXkEJa1YSWwHYSjrvaxl+EOnYNcDK
ftRMhJZ5uLU62DlWnkO8ZvdQESbnFfjZ+ybqVmIr0DR0Z4lHNGyIqnwpuV/I43aLgm2XYJIa6llB
8mqtxH4BvMEQJX5cQ1fEJqxtrW86FbAJQazwPBSLBlyFTpZUxM3kzCAzomDmuw6IJouXgkDP0pps
UJMb+SFRm+jQ8jgTsPDgID8XTvomhhaHCNzICkgPOCGifIkGPAbUwHwig+y1GMkFqj20nkE3l2IB
0Ft+lr1Kv31zJ0tvYWQoBxUsHQzG4+jWhnQcx9hjk73G6SaZ/tAaPOp6sCfA9NTsNA+LU8BfNtNQ
LDbZkNHj7NX7BswFEywuPvionGAxzyod4UJ3/rhF5US9x6CzJsHEE+B8jXWhBKvIGs31ml+OLDHx
IYJkxfcXhcRCDiLV8IAYAVCzD3u78VcRnA/B0yOOON+cC6yqzpl4QPSzkKT7PxU6taHe558t/my+
+K7EV8xLFI65KD2f9iWTzCGge5W9IVZkDSOJ37QUymMc66CkMeaIUxEGv58ljSkak54xpvpNDmvk
Pk5AUCJIDTHx+EQp9vYFw9Ncsk86f49bug9SX7dBRC02N9nZ5Em2b0BdRXuMd64oPww54LQn2VQz
adJBJvE9UNzvU0U4kVAl1641NdVAE94RMEXJ0c3A880mnCFKIsWHFgNclFzzukTx7nX5GAmxM8XG
iiZiHS2D7DhZ//jNJj+84AA8RHF5p8WGn3yVmSfMLQegLOrh5SD2yK8l9Ng8lZ1BczLQQs1wk2J9
8kNCbpnK8PuCNAsWmy05b7TOlY0X/25WoWOs9BwhAUSo6EnalwAFptnWTqQD43VfvKfgEfxjmrHv
NSx6toCkoQBq4w80WJ5/4d2Qpw9kkL1WZDGaPmbdTAjoqr07vX8h0zStFI0NzbYn6GSTWJM2b+ms
Rpt9h4FRVVPevlJel9lV5399nVs3uvlT3rwNHIh5HOhs9526490a/UPtXzOs4Unlmb5WkWtgnyYS
BrwoziUZ95IePhLsEputOfRNkz7/eC7OOjpRNPqMtIWl4yM02BEI3JE1NExzG7dAa8bxgkRBL06m
Lx39fX1tK2Bj5mVpbM5p24gSb9YRh08jmq4AzYncHZErEdb6DJbQUVM/wOXGvhVjx5wlSqk2kPNh
zzdXe4VUUnxnAUYQysdi9MhKxUXZXfv1wDyFd3cp/AD80D3LFmn8HwUzQS4+mITRfoeGGF092kiI
01Vb8C4Vi+qJWO5fUuL1Cd+UpmrzHTBXqkI9fKtv/AFIUhqDQntIHpaSK1hqKkVh4W7WrPTbFJq9
aQl1MfY4pGX+E+7HuHs9lE9jDVFOmoTJl6R4aO9hU/hbaI2PGgGDT2dzOoJXIW5eCjLd3svYobB1
TgcZAFHcFSdO9MJfmAqq6vEzFqdZuWVudjFl/FnGBVVYJnOhZDJZKl+MtMFQ87vXt4l20oKkfNUH
NfB/UjmGqGE/rgo+QLtp9Ei47/VEch5wK1v2sjvhflkPyVjmpm9XPzOteRSgT0dqd/xdXNpM4ogF
6dxUwJhAvyBxa0JWQ1uq7nyH98n3bWXEY9FQz8OEnY01i6wIFx8NH7olwI3X6G8wO8HUoNIvAoQe
ff7k5/j/xnZTLF/YpO3FL2/yEJZGruxuC5m+AtTU/XbccM1mL8dKwjCN+cpFe4FAV6HAPaErMtOM
HNJD20EGB+uUVCC1xJc/f6gotzPcZ+GkfrotV3xSe3vFm1aG+l9d5DQ/Y8YwXDU9jHnbr7L1io3t
YDELUMlDtxpGdO2yHi4FSi5utcgTyqPz4beosvAgkrptrrCXxiQGnTV3EPSFAYnfW7tlmw4nigBU
+5HVteKLc4Rrb+6h6HCbkZlj9wh38A63cg6jygBKS0nXK3EJQv9Qmv9I+6Dknm5N+qWTPT8+ii+a
pnK42sLg/6b37Qc1GaupFq6mgVATER793wZSISfNxz/vaERW9usSk7cS2SlUh+phKP7d18XuI5qn
zjWnUmSz9wzMAEZstvgxNwNDiJSsrYOYmNTg/3cCewlD+waOnTUWpkqtvxI6MQWXECnxNGmkEAZD
+dX02ijlnDaT1Yi1KgyM+7ze1jxPgV1mui9mk5Gq+U2lqDIhJJpt+RwNO7VL4EBCu5OhGneVg4Dg
JSTsfJChtD2V3VPGcqv5oV+8KfEPRoFthZewTIAIs1RvEJxDhaRkZG0+P8eaLbh5EF+WrxmoiEzd
AJkgxyBpJgsfKAbB+NsdIO1Gj4D2XiKQDoPpkJwBCV+5whH2r73QbMd0MtHKV22Iy37Nc4zEFx8j
vk10EGgZMkYZ3Q2VHAIzU0pNVQEGsSg7MoOiORvvgAaVHIiHqIx8a1lidjNPyDFWes0EPeqJtoWu
igYiYu9vK6dEQxNVzqVHTYSMr8g83UTtgX0od5aAvkMOCybnCWGHGIO2C98trFfoPN+xJTW8S3WS
PL15IVf/6JeZEzzfXV19viDGvV/fsoeJk5cTc1NLYO9Y3z5mVF/Ju+6wjVdhKEd5nlovqzSiTPJ3
1LaIh2oF3TDnFp5fA41PvUpWZqpiDaXKXzlxd6YEZ51StQYPGXTfzJbRwzoWC9ZvruZvZPzyNOxF
SJlsmNrMJgQed6LnYln7bwc1/7H/zo3T1RufFpPtpQIfqT8EL42UHStA8/GoyVWgkcgZJqZDZeYw
dEKeiz3l3MhIovijTUtvw65em0XmzdymvudHZaD3QZSKdtkHTQjOqq8YV1o0s63ezR6bubdV0y+C
n7XvvbBw/0c/RG2ii2rooX7gVn0W/+h/XHw95701L5uM9hAps8/B73gw/XwY7ZV8htNcrxmgf/40
UNjgWhgxRS3dzA+8e6UhPgAmXpqcV/fqIOLBioBcarj2wKxjRHiVEH91PiZZQ6V42TMsbzCD9NWY
lqYpumE+qZV5TaE4dpm0vEt+0OYpZrBkbf0/qYZc5Cs5GBDR+lVBaAMlWA2JWAeBFKuB8nw3DJ8u
9+npNBpdMyhgYOsK2LVg/Dgyi0BPSpkSCN9xXteMsFvuEz1PBofBVjpeso2s/lJto17k+eKeVlsx
Tt+wGDXciBIhs8viYC1Akb2Ni92Namit7TVR2va7vmL68VlMwy9enQB469TpFavA3cBuWBpXAYz1
VQEHZVJGDN2u3NJFxWRuq/oaN2bhKiuaNk23v0Cofdn6mmwV8E5uaH/+871HaAjFGuCeHacGDXXw
d5hTaXhK3/pUiIwx1nGeIdfs70KW29u5jrntqsp0pNmqF74lqSlqf9TPaftj7e1Lypg4zx7fTfW7
r20I3KLIegcrPO0tnb57hHmBy62akgNijKpd7J7m5wwT3nvDVMfsB0FfID5rLAlRKit2F3IE4+5s
l2bL67ycNQN3mqY+KzwqbQ+f/LPmZzzWcMDv+OpZe7LQt0VTXJsQ29EQQ7zt3jRc62rM4vAEKuRs
DzTnzFxeSFLyXfKqthbzCP2HDX4dLTeiGV4f1gq7UErqUqRv9uBwUhqTMUUcAp18wIDjcYV9uvjg
v7KAWxFJCbxTQLcePUwc4C8wketp6530POU0L/C2jzXLag06IC+2VSowA5JAxRmhjKMuPjXqoGep
3sni1fS/ZxuFVEdRCyNYlrDiDbrPQAEEhFmBo9mPMEQp4ELC8YMnwhxkMAwOgsI/+deo4nmYHanO
2mts6F+vruMZCu3JYORlB7vltDUT7K3F/+n0HknBkoJ8KGmm5eYOxQvtxlsE7G1sHfOjjjpBjlWj
oTdRhFf7XCUWD4JErrV05FFxLmq5hMjk0VYulbiAmW8x1AoXiPjanmrlaswCKXEvsALOuziGbBTq
1mBav+18gjd1Ix8YX3lxFzyNWaO/JcVUAM4p4bALh0ymnl3KrsG+WgscnkYWle4cxsWRGRX41M8D
fSe15SQ2oHAIKpJpdPhmjnNXB/Q6NwDFfKBd6v8mIGmA4tXBJ4nG5/Fh4isYwql70WXuvG0KnZWx
WwAuyYFvD7t1z4tvZx9cB2/aAZwSlQG/RL0dnjEYkl6ZQ0FzTG3tv+GvbT0IJJjORB4GseZYIu75
ZQgwFGQ5y7KT6wpwAl+OocsTZtTPRFO10BGfREvk4EhuWXcg97+eBdiwVca2Hi50CqQaIiTkOVdW
KyL3Am4qpzYOtsY14IVbfrbPkPzntg4qtTcDEEaMdtS/lKO0siE4ZcZc+5trx/xGW6svIauQ294n
ULnxEL0nX7pPJC78DZUHq7r7fK2u6OuWeLsmdifi0q8+aiHrKn12ehaifADEHOTneXzNAbsoz/yG
yhfLDjtqeLyDS/Anmw7L7c7zGt6gDDxKR4+8MwudAk7X74Z5jnrW37Ai/TExF8Df/wjfpWbZRJgv
giWgWkckXB8VTn+2TaCP/XqTVAeSW5q4IBAoIYbLV9hN7QKOhUSLVCcxCvk2oVeWFePkrPf/otGv
0scupvfT3HRyTBVmT0PFww7iLi9hMvx4JMoPkH0cgeG4BOvaRX9BzyIlF3FS4yHKQLuNrsM6oAsw
XDItV/PuxXpnUWxziGNxkeukhatUjvhFsHjbVEkm0taXLU4/IOOAan73nMxB1SxPf6h9g6b/4R6S
fuLU956GqFhRG8y2jYmF40IBXo0HP74EiD4QorlPySHw6LBdoBv7WyKkAW3poAJUxYV/MUouEx22
I99sSqj5HCGzCc1JZQFFi4vGnWm3QprVztb4pTN5EaMuvMMwv+qDx141NB7Oz8DZpCp/J+Jhkv8v
80xdJ42V/hLIAGFxwzNYmhyBeTqzH1ewL11swquFlBXdQ0EdBFn01om+eUjTsA9MgPMeNou1QEfy
/kQv9ijF5PKPRfe4Uuik6SUMoy5W4tQtsLaKP7HzWm7ASSgtF7OHWbuCmnYNJ/EWxrg6EynXcDBa
+Ej1gH8SVQbyT/uqhhUkpIF87MkFa2shvw+UcBcjn6LktIjzZ3tSJy/Jg2H04gnffE/GNcnWMCwZ
8LgECmDod7GN7dUa1tCm8MXdI13FsyAT/gRrUYAMDknToaJYZKKsNtPZdy5KUCwPt6pIhGuyEpJR
r99WusSYd7yCLvPWm9Lf76Fc436y/a4x7OoAPF5Ml3jL+ai/1nGnmMug+TKR3wkdr73cOIwTpbP5
XgwijRa22jhTX48TBkWw0c3ZobtT7rN1hbwmx5VJHCXwUdUJ61+43+i4AaupYYoACeNufZJ0U/WC
IYn+cl6hl0UqEu+x9y3H8lcvx9McbPeN1cy0jOZ62Z65IUoqoA5qR3h5iF5oxwXgrncJiZmf9Uzy
uimmqpyzzRrwuD9h6xrFznVfLTqhg8CLyfdMX2g0sv4iSBmT7HC/fUnmYwdMPU+ZhN0vEDA2sWgm
bI5WEoL/QMaqTlt2W1IK5EbTVsmzKDI2UATzyorD5og6jrYNFoHNlHMJubPSCZOqXcZ6M3pDr5b9
4oR1CumUN73U331r3sVkjSn6B5uNJcHp5JYrc37QNjHP1ezS5/yqQ289HFhmHoI0JBDv3pIgOQRf
kogK3k0+l4kAtq5qGQdcwh5+jo3UoI1R0GF6PbvwvUQF1rAjTQw2MxZHhjlJI3Op8Xc2JvOkxI2i
ZsuIphzb3Rbp4jV6b8piau4dDkjxSnotF4GGE4XDVxQGTtOO85gb9sFxlTPx8tycaC4fBg5z9Qs8
QLtBMZMYewPjFG71EmonvFUd77iU8Jy8NLjw7mAiY6JQ76FJfQx4PoueAne+f02VZYUSfP8grQ/l
H1RzuKI1ZQfR7Ioe4HIjhnwLF0kuJTAQDbcP5qHSKeysO/pBy53ol3+etXFVK+QiQ39hZ1XCSpPw
FGbSHRK1Yqc/S+Uo7Lb4E5fUscQFWkSXy7aImulaUcXT/yQDy9lnZkZWAH3Agny2NXkgqc/cirmD
yfXmLUQi1nX4SOKpW5LJQYOInjTeYl2DjOoPAMGtBg03c7+bM08NTEzrAot27LxyVMZaZg+/sieP
A5p3PTTpq+8iZ7UGKB5+UI437zJvdiJzc/nSDG0u5yR6WjQQ2PCq6TrrI2sZ9QyHxuIlkvYq7+Nx
w1nMkelNaUd8fLXl7dB58hJY5vFWX70XPuv2QijksW9+QIzz8jAbZa4eEocWozL1ew5Ld9UyaN5z
BLFKCA7wkSWJJBO42KkwDDmMMxkmfRl1CT986e1+ESw3ZBtqIoXe4aHLI2A+ssFlcfMTrLozES4J
VYV/i88h9eRc20pdrKjjFu9lT1LHQHJZN7bNQOt/i5AhuF37Mk9vg9DlkNzv1dzjGHBC9T+NORYO
Tf6MfS9Hiq9odSNr+y8k1PycoiUIExI4aLMvm9Hb9BHFfZcyBelmapjvzQ1zbCNxqT35Ugd9nDek
x1uCZTWmkZCaNYkfHe0XqEkCvlGM3EWm8XhKhDopXDbX1EeOe4oQNyxjy/p5j0PEuMJfNNeVM/3D
vGl359yZFnxZSNn5Q9Wo3HkXyQ+RnEa9s9TaKNYcXa7ct+v82XlYhTZs+cXvLcHeO1zMVjaQH6c1
8w/+oEfyQC7J0243YPN9I25ASGrMl9+t1pnEqXwR79wGZfiMz0QHUH6lCGUL6VsZ3uLEo8nF6n6d
4OwXJogvVnUxfybgRsOCsKllqQ9C2F8rBZQYlVdoPs6gZmwL3BXdapnlZTIDk73AeLGsNfzcoSSS
ELuNSjPkc2DeUVP8VxO7OULBLl1CFc8dOAPE2EiaKphyLBDpBLaYskUb/6/kT9Pp3jDv92NtMLtK
zzmEOZ5ePLAXYEVcNdwk2r/CswSd0G4ggOnG6oekRsVVII5bSXrTGhbM4W6v0Z3+GSQ/Ll0TKILI
r56BfRDhiZLPg5Y7U9W3xfR2ZMv4i57bw12S6d3yqeMvbJA3p0q8CNOr2XIq4NvHKPpNNAmXNYx1
Sc8PGzi+NIU6PN75+fxaV5wq/6Q3gh5mjkV0Shm/6d4fw/oiTtGUsXAMb5TiqvVQjcbpbwODgfLX
HAcRCcGAIV157hbC8LXs1hg/mvq3FeNMk/6Qov5C2xSFZGtZw0KVhDZACsjtKlv/27RMnyYH6jnk
kfwNBKfUAP3XgwUNx72dOODyElp40pM8ix0LNBSu6t+2wwr11Cth1IwZKHrRCZ9dVyMFUUGnYFgY
p6evfcEY+wEj8Cq9NuOCpE4T1aFtTE2lp6qnHTPjwZ2AEa7DuFqx/IQimN1E9KN49m5jJYY3w+PB
nShPeOUbd6eX/tJHBEc+0NRbCFBL6b7QpiuPnoUx9rGk8WiaUitwirxTRYm5ohbPfh5z0XIQfF31
DFFrHei5a/fyFWGUHDQ7vAa9t3fm6Ip5bBnvWScypv3yDUo6ZzzRQ8lXBUXsSEE9J+4Ch9qTdGCZ
87FTAoHJCjeXHhrRIvG7NY2168RuuVxwIMW6qjLzv/FKArUkFB90A5F6zc0OjzExWxXfOp51sYSB
zi2HAxVOolZE3iHrbLOqws/XKUT0iDXsjU/CsVpkFW6BCOVjoSrOHh7QXYN42uVNM3qAEwCBgokz
B4GSmDt2WPUk/KdAEVIG8D49vuGthydvparfWTJGnDcll97NsXzQgDFDDbscsmJrX3Yw+Qa1Qq/u
5xVbgje52eU6zgZ2w9W+WkktXZI7xu31L9nS0lCMQcKrnbmdZE4HRO78dO37qReEoUjzL/x30ZEU
MG89lf85aw1msy98/kEkjzEuayDuEQ3FMR2VM0LH+ytwGBhwOvVWUDEZn6S++IpflvRI+LYRwuB5
LXKxrjYycbCZAYN4aZGjU+ikgAZc+VDCg+zH16S/dmn0y1rITxBv6cywrwhRv169w81xxovv4MUq
VIKuoyChRJwuhjsE7WnpNt27/NkmpwJixw6VnLcL3pZGyizlfYXxnAVrJMv0OzwPoFKusJmIWDOb
goS9qRRfAH5DJG4iP7z9m6MZPmcCA3V6BQEVfhrnPPcAycM8AJcq7B8fy+9ujHiW5ne560Gv7PaG
g6G3+nLXaq7JyfkjJIRYx7pT4jXgsz4EIY8Uv/i2qTDN/0UAmhvNbaplrdPZ8ncX3ufuWc4X88Pa
l1S2AltaqPMmdQLg13KYKesQfsP3GPTHczOBHe+8BPuqauOS9mprjt0JR2Nv9WYB721XY5zGIlUw
bHInw3yDMvVxMxxGfvS7+tv8eoDO/MTHUZsc6XETVilpXLsY/yUQoypFi1IzsZx8TZH0St34VYjp
z3Sne9u9Bg3BG6AXJUL5VwdSWDcA2/yYVE8cSLk5+MEuvLSWXKfKbGiT9/t6i4L8gI3ZzsPRdRdi
oB6KmHp2bkcjCuPHaIb5K2Vjd9tkuX0y516bf82zPNvIztV87GsCsKcYsONfA3lveafq9wEzzRPK
LzZwBK29AS7PZhaPf7D7VenRiBFnziYddYyIK4E3zNSZN9s1ZNyQXuIkFWvAftvsjgnGdg6ozPwv
1goXbt3dSJfsUwO74ID2Ig2HpZYks2W7/gguFVJP/3DX8wu127u0LEton+gcMFJCjRoutlWTq2F2
vQXQHFap3WeB+AM1z3BMJQoROzvWn/ovn1hHary2N9/ViUaxS8nd6HIvHc3A70dOXeB1owpXjyQV
lfhBVYwtcHbnRgPTUu1EljXGzH+NRgr8Wo7xHdIK5CrYvLWmDuEzeXkVXb7WuhnpEfNUVRHn9IOE
4pQnKBei1rApOOcPv/LGcMVHYUvOo8RWT4uuxOMnm8LtQvhWBuYNQot/pGvvoyaGv2Wn0UwG77F3
lox/Snv3z6cBDhB3NwFidD6xOESURD2NqcBUr9U1yFV0oi/lCJB4CYg3mZy2f1F2rI+WPOVm8wEX
CA48bA/tyMJ70reQqRlTM34HptXL3FazYrVS+uI0MkSmbkvoeqjq8GgSOTRHoK+fRsn4NOzR9ing
nHEh5XmEcyPk/B5Cl+VJn2N5L5E7uACXHgYnFY0ZX+yJKBQe5LtVZXsIz4g3crbCktlU7yeH2imK
qy2r+eKakyVAm0hNZ9+U6mjL5b4S52YFXTfeDGsY/RXk9Bt2pBOJhUwwfw5nDDJV2zw4PZWYCcaA
0Uet/PF1b5xBJxyfDIwgjjlKgphHQ9kcMr2QZJtiVKrKr1GNKI1wmLcb4k4mPPb00iZolAP3BcIa
LCbdtIto2qiyYRELnk57pYZ62VBl9u9AU3Lz01kS0SCghZ7FDVXfxCM7aFoDzL2fl0TlE88De+LJ
dKJEYm+cNMj+lbzbccMdOMh0+wP/6nG7QAYYRYWSlkqjCXqojNpiPL/hq9WQ3icJpV2amyQDXutO
uZQCWj67WpSCcr+dHBviTSjb94kcUpGpn8USEAz9AtW039n/Mgt6e4eMb+lkMxB5BFZt04yZp1M8
aouY90WSo5xI12N8ZBPHMK20XA5E0koKq5Dy0oAhoSjc/AQpifzBItFl/XgChCXVuHZUhZoeFWTU
HKod2J3acEFzEXCzNl27E/ceX6utYPfm7g44a3aYDJjP+xolPwmrg2dh5QZp5EyZym/G9LDnxGm3
KjF1dQgWclxRG9W8Xu0Mo2KZghRu0fqkL3p1gAfUo8cvyN3+f3znpH4xLXywe7gVyXkrimcRNxUS
/n4wJMHVWVcADyYMj3WMd8tZPcgLVfXwYTPLiUocaUrTQvqjfiuZMo+4873rZxUsifDWQ1Lq45b1
2QnP90Ph0NNRuSE8mc/TdcdaLFbsN+eJO2QGh/81gM4ra9IJBCIpDGf/n5JzlB4UFu1B+QYRdbvT
UGPinUPNJliEE4oCds7Hkw6BfeKZR4DLsvWDVY6YSBTqDFOjqFgbI5K5SrIE6zyL/LKQLCl+s1vN
4I0WhXzE7SKUCKcjBri/f7s1hFqlPDT56WLUt6ucJFjEIsGcqSruAqvdWM0cXd4130LYIs27gQHu
Wj+yZUOh35yq42s+X+Mj1B1ZyF8ySMqBTZPs+uc0Uc6Yx33HWSBFFCW2zpABf4KZFkSE5Kgx54NI
iFY4LBWaa6N4L57VtrKmNLzJYeA+Ui2z09eQNhvtabZoGdg0GS1Az+XnHEl3dyz+xLcVOWVuNX17
+mvsXCfn/vSxEbN9ugS5HuQoAoRuMlTKm2lsyQMDSwGREP4ugOVCREN+SpqeWvlZ4t/rS0umjwU4
33R0agRL8rxrTfcztxbzfU5O9y27sBVxlnvY8nSQTLjDiDrtg4RNpB2bK+COHWLZRXzj7AQUDdcZ
6Qo2O6e1EMpp3Pf1H6ZDlpu/DHyrIe8Ip7+D3FrIImTNit0G/3svmhTO07sFde9T1Q74r+8uLCNC
/w2HmxkIUjybNU9o31IAyIW9O1AgYtlFoO0RG52EV0rmricKlSGhQDT1bwx+Uc7blzBGl/bX3H5O
6UM26KmOinSfBCaIpg4V+KWGtdRx8GIx7WpkfQOC1kMYUt8KJ5gTzDVtV++Bn2PZzfhTbKERcSmx
QAe8kCmFKa9sfGeP3NiI2J0pdF+rauNEA+DOEpFBZuQy2rNEgOIFaqYTnwCe+/eHqCRncI1hxPd2
ogPh1XPvP/k1vimat/kyF3ghS3LPuNNUa0NKB9erxpSkA4mP/JGgGYD7MR1yYmW3JQiPkPPI9usY
UOfbI7BjVt2hYnkgQTAcHu/YNjGfLv0VAQxx9USUeMkEpmSa00eNO9L9WS6u79Ad8IUGfj4K1IcV
3DYHxrzCZhB6PWXence9kqTsTFA5Icdih4cJfs3RgM5l8QIRTKILOigeYN3WWG6ioGVIQerBKsdS
C5Vtzt8Fkr4etvShsLYNRKPejYvJ3lDt4CbRSRB7wp5kXznl5acBr5q7Tlg4CsUUBCij1j2Q/SaQ
5E7POCMpRoE+/06YhTKrSC2c4DFnl40ybVC+pr0udiJIC3jGdBvDpNkjQEIendvJ7k+X4IyS0yQP
pd5amkT0qr2hTczpxi/8DNW4P2gYlKj0UbCXnf9UyPa2i4EJnqZ7V/6yE0s73F/KqKZjZyadWr4O
kBnUd8Dil4IjNvO20doXisidc7Xe5VApjMIdzGvpYMTcCMwr8Lsly4gRcGPc5YscDvImfoZgJnsF
Z8N32d4lOani2XO0YRX+cFyoWrnsmbqIIKbPYdtEr/HvFW7uRoyyqORc7K+KQgZd9yCc+J2QA6VH
kO02jTMD30Cc+WUIel0fxGTyFGDty6t/OoeaEAftQHx5gkMmMMEc7OIUJnkowQxUbUCTymiIzgWV
2553QOwmZqnB7DyCJzWCI8/0EGxS79CiOqrInYt0MffJ1GJZivVjBFG7BqzZq+qr/Ok+4nP3vgJj
KyZpIMZwnrXdKTcCPcAmC0Xaj05NGAjZ9Xr6iH1UOPDf1XQLl8xK0/F/SbDXlh24P3m6gTv0Pkur
6fuFu9t0zbTk4nYkEOohh50JVgx+B6nU8mzWelc6YykiVGm273VxCnbfVM4knDaEDuCIcpq+ibjl
DNWvNXCSzZPxyZxkMqP/bFL46zRk8LCUq7zsmPbZd8hyjGRn43HNxvG4rCct3uT05EVX3e32+wdZ
AJhdmWUbjlBVK/RG0HcfqCg5DWyEr4vCW3eNIQPcxEVI9k7O8oW2iyepYovsZWKKXdm2Q+zZyuR9
f0Wua97pQCcc4nWA+sDhEoz9dUEHiBL3WV/qx6QhLlVrSwVSupBT/1dmfmsaD+pnT1D89RYfVU64
10G1+rkl9Qsk+QYyLTQC2vaA2uOSQOMsRONK+YMCzBCjm/z6KOTPQf8SlKbnQLiJilXSra7ZBixF
cvAI2eNle+q0ogzM50JjSAq3yi2WDeWUG+MUvjj6RbOD4uNOxTUtbvQnW/9RRjAcl6j6aK3bFiGg
sQl9+e2yWd7AwvI6hF+UPOUf6wfqWWOy8g402dyLxiBzQY2iWpQIAnmYuNU7PdBpN3R6Ef1oJyFO
h9NMHttKTj+AIwtPUz5PMJeoOJsAYQNPd1jVTWYOCgMUjPKxy1+uweX01c+CSSq/g6tF9kciJjVQ
GHV86jQZWIljAGeMYndeQDKCdpk7rTTJlB4HxJ5JfjwCLCQ3cnTXGqTzfP0ogP0IT4H0jz6l24jM
WOxng1gwi5tW19uuHeAdxccuxgjd9ekO+0JYOAzDdkaLMkBsvLIhd7HVIPQBdlACrRR0nf5kho4f
9I/S2glbyRNB5KuQLBBOLDuasOmqbB7bBubrOoO5N6tNBTCqUiGd76tebTBVYtByz11vqtuFakAz
mtd+iT6B/8kFeXSwpsjJZXoWTTcolpj9N0hB0+ik0cp7yN47uzqDQgJBsJ/gUe9OGaYyPNEuTKgb
WM01IPb9tpmsQsw9Pm2gghGhPZiwkyBqKhpl8hOnlf9AgZgpunkPNJfJ53+IQhSDhLVgU5pjS+FR
2JtuhnTnADYO8ssHVxI7Uzx62zZXw8IIg5LkZM65N+nU5arQoGq7pJQLf20q0hwyMKilhBm/aUXe
E+znQfUIjqW2PjX3rqrj00uOEGlx7NR7z68Udu/LYLBNvzfzVUHAqAvrNKMBJX+5B5eWrYesrGy7
jmzy/yCgkA3vH5CZxWjCJFsytsS7+8DuoKs7KEy/sNc6KlOROOLheSshLyMeEmYyUpoPPc2y7L3q
m6/NE3pOf8wycZQrMTrX+hBxJ5T72qB4RkxJDiNmbb8oOgrSE++Iv6n7VUA3Q0fqzDUqP131Y63Y
ji8X3/uo9+6WiKbX772vGn/lw8889dHe88FWpEhNnUdR39v5Zlozi/2n32RAVaxByQmLcU3YvRGQ
XQR3OWYmCXHLa8SbvC55NToWqPEtOmudFwX1WWCZEhG5QUz7MdkdZfHBDk3EiHiXi2vN8e+cAO/z
eGZBMuZl1Cwj58lcC1aokLosZvXb+QWhjs+OL355drCCERyvw6DH5Qv+XouTtIrzcwJNZOcXJduI
y2LZZBpLlf/Tp/Ew67RBW5ZqWo8tgpNEhMYoUb13X3RUMIBD+kxHXglLrdCZkrfxBuC+bGlaoBZ3
VDP7yDd+4s7uWjl9USZueJJNozFWzDhprm+zFh6imerfz9tEVyeuRes9jIwsq/zwFgIH199tE9bf
9j+Q/OOLD+9hSrvOvHpU0ehJBkBQuMwj1WCUur+xm8plCIGlextKmPirhbpmxA6kRBbsNv8o2IbX
g/Y7j3L2VkaWFMabUh3VVNYv8pHz7Bc1+2W2zPirOQmLpy5GfB04xI/tiV4mIibnp68AjNxKOZaI
7Ks0tH8tNALYYyasa7YO8w2JGCRlCXImgjHGyVFvJAwDa+NzGx7q5Vnj2rBn1G2woxC+Ea63XgHA
NVFU9HE7xWHBbg9EaObcKq0vcg4/tsGPQaL1LDnQTUg/rT0X3ET2AUbE0PRKqW3VNGR2Iow3V5zU
OAXaRTq5jDqS6oxMXafdyazBeyqr2oNQJeNn10xEX7AK5X8QWMNQvhzDf3tPmGi4+X5OY46qVn+/
VqQo/enkkUF30ogeYE2DwQmnelH7T5ElJjU6dfF3SPAXF0/VYAEOpz67BZ9Qw5HG7dfUJaBs4QfB
c1FBSvfMkjg2Sg0v6It54DWq7IL0pXQHGa8LluXUyYml7nBvdVQbs1fMliXoqprqldZ+hi4ALk2+
o5sYmZAk6k3IJXUiow7E7FU4e5AJzVbOHWPI6FjsIJMsz9K3ZX8XfRQ1SkQ3QpwUAmvcI8AfErOt
x2vuFi+nUk2LZoB/vVWUGuHJBdIMCge+6Rjf6ak/KyCOdvMukd8VvR+MbHsgERWbOQauItNqZ3Si
Tg3vvJuWfv+odGyTzrGxSEipajRRAsHCtilACvD5T1G8PmwaZDPacir6B7MTfeRwfbowOPwEAIxW
PURVRLnAMQY/Fo4oUi6XB9Rdyn91/JEgBdg4U51K5YTPtNZdCvMd3tuZpPYGIBlTMbmrVsdV7+k6
spM+olfQgFRUrJwtJajt05FBR9IoUC+AUUWjw/VziW5UCPL5NTH4FaxkvNpfl+AkLUGujZLMjPVi
cK221hobsoUFRc1q9yr4x9lsUiOct+Y4int+caY27M8EYeNwdQHonLa2rGpqy84owziMizomxHpU
hlxtJ8MqAUN3aYsv5n3y6CdodceKJNRx+I+RyII06hkjxXge9uSBVYIo4j2qe3Ez++0Z2tLZOv2z
YOsWsRNa59Z8FfXmTfi2EsZmfTiuwT7YK0c+Ig8p7CpjAnWZASyXl+8mZ1SQOSY0dP3iAe+IQNNA
tDDCHkOtzJeduPK9nQodjf9IeLihfiQZOUPn8r1SZBNl0jWQy3BVcwufQ1YYXq7BuBNzgeRmBrEb
Vop9AhVNEPfdO9UNqlnWAE6wo6vcaGPI7PTYBrehMNxxzV/4kwJuR3CfCVUfmolDBAsIg8Hs4iHE
aDFTJ9V8X7RYNkcM5e/Gzc1xCORF+HjUv3BFoJW17mc0CkUBXdtlUTM5ZrfI5TkoGYaHuGWl0Xto
ramYjrhfiZMFgvqTUJwALa9p1Jrp2erWEqmI8R3PaYih56/HQSiLkJ8pk5FKA5BdwqCW5fGUB0s/
OY8+Hi9JI5Y+TZDzdDx2tpBpW6459H/DfNu8FgAmhpW9i6380fr3WvP4F2sXlsSRAi81GeZFmVIR
Ykbszxow4HcEgaihYhPfqNHBdjGWjesYplSH11J8QO56PMOwYRAKZyVfXPgSTxRk22xq3FC1ElsJ
/MCTq48tN1m4tNmqus8RehrsJ215aADIHMTcX6kvf2y0G+LAW4mDqdSu2rNN9hYNiA5AOAFeYw03
pzTEFb4Kpbg14HMNQaDuDZpuK3V39NXj/vSBGX7S6a4Niy/+2hYBRPLGT00+fkUa7qEMeqyxWTfj
9u0tE6L8gSXKpqXnBrP7VRjte1jHJh9EamVahuwb1wJexqQ46tTO5TwCgHi+ZnHx/ymFbpAV4bMo
WzyzbeXqyVRHL2Zur2P0LGpvXE5zbCQcntVFvaxCGKZoETbiJQ29D9+dTyCk/mlTPCJrYrSiajHy
j8+nHmXn61foBnx2yTW+xKURY70tpDOGN4c57nQFaTDHimtWlsKWVMxHoTOkYVUsg0/PtIDoRxXI
983AGlv8DvL0nwYX+rvDJopr8JkTKxIP2XYUQsLuW9hv+TaGp7FNtXg9bQSv8VTCg2rp1tYIRn3B
FqrhUXIGesjFniPVWUjUTHe/aORBDrujGDb7LXiTM8o5dsxQcExFWYy/4MKmUXfukBLHhsCM7No/
sQUWWsYf3jbquyYtvnGZs0srIrzeBwn6z2vKyRsR7WZ9UfWglnX0qsAbXaqCzqnF7nQkI4PWoOmJ
SemEomXw7ATZmhNo9DBEBHxMd19RLx3XDbxmLJ61oObpFjBslDqBd1O2PY7J9N2u2i9jgGfPgbZI
OFEL36/jR/McLCpaStotDMbkxJcTUoKWhcSt0MLoiBMCTqkcBvoVkqVI65cO+fTBYpONq5OnvGW+
soH0FCJEBGfJTSovMPRwBn+ApF1AYdbXpmgMvznp+nhC53plMUKanQre8WnfdxVLaXJ8JMn5T/r9
VRaXYJlBKLIaRg8ew6cV6Fisg66smZvYx2Se32equ92gnF5hX0e7jUJufjuNV02YnFpsNi53a9A5
eUN6NkIGY+KPFW5k6ODAcsJuDx2IOnqzoAfQ0on/AW3FiOFN5YYNXOFARx9sHiZ8AyNoUbzc+tv/
ZB+f2n1OHNLYZ7JLVdrnzF6uRDOYyhqkHe5v+7H1eE58z28YetFlb6n5XgRr5P4zDJb8zGKILwOZ
s4zYAz7576lvRqEnkk2JW+YjDdi9FUM6qglSI14dXZVipKBqeiUnnejvWDW91C6vc+U6KO0mRvgl
+0SLYpb18hZR5jtwV1E4QLFlVSooiwZdr8A98ftQ2ZSCIAeO1dAa51wIbLnl436p5XqevCgU76yO
MILeA2L5PeOC+N2r1PuP/hDIFV/0lFFu+ESalWlHGUDfudKwF7YBnwntrK4qFdEwHuQq64/VpvD3
jbyaUTZhHfjN+AyNVVLvPeZuuxd9mbN3ixJq8EG2EIrJXdUMBYxGcGgUnAaf3isut2g8AEztGT9v
uhxKIMRM6wghrRvzpSlHdichL4ZkEos76te2Zfq667NnHHbqUOQo11p3g9or4iB3IcyXwaqn13JX
E2dz0staFC2b0vHUBH/Yajv9B2FjwwaLx8Fx+YeDKP75YAc3TH3X2cbbY4j2t5BSQYguBTkrhWpL
MM9Hdci9vpqYnmgxADo9b2IjGWFaUP7vGBowJca/5B/1zcfPRhm4Nmh712Mym8Kw+l6VBv1h9UK0
4bO7LwdcPoSH82ozp7kAsiZY5cxh59gzwl/o0/0T0vNlGnr36HYxP4MKMUSUS+n+mxQltspR2fFz
6pGWsDFvVppsCZk/dZW5RaFTEeN6SvXz4w9w5DYZB1qVTYQHRtU2HzRBIHiW2MDQXbN54OSQl8nN
7n4vl5hyXuvtl1Th+X2IJUfG2bY2ykkVzEX39JREZDN6YdixEK2l2aBNrCEshGMXfqVTfMLS0VUV
+28LZb2EBQcy25Njtf5k29ft06CL3g2V9+N7L2vwHD+EuFcPgwG4l2Q2VJ8SYRINuYqLKHbg5DS1
uLb4xcCjT+uXMHYAs1P8UAYAMRgk/iszZLnUiRnnRSUs7yokwiRkdzSoCL+e5BqW/S9Bw79uIWsd
WkKSyVzfYeMiV3+UylQcYeV4j9+OHKg1PU+aHBBaQFdldfThEtjNg3a31tbhVgMSZMY6QMdp5rYD
f3jQz2VVpLfMzL9CrvOE2NR7KrcxifXoxL61uSDCb8GpA9bALBguOxxISRkn+RCpbvTAOS9Z9EoZ
E5jUZbYAnlZQiKufNzp6rh03za6l7r/C7L9vMEwoYOv2kj+5eWTspxp5A8udpH4vQkGmOx7nnMAf
bMN3g/SAsZZJRASdJhBJyk1/+I8o6PdOwenDrK0fkF4igcnMNZS0oZXawBVS09G9ASCBZpthG+xO
ckJNgFfErTM3OUwlabuc9APVG4j8H+xrclQi569to7cIHU30FvbKk92vAaF+9lvr1Ss0JpaxDFgj
qWqTPoA2lz7Mr+EsEJNK0oq46JvwZqcv6s/Y1wHW2HMBmlEEnFASNJUicTmeRfOFSO/aOcH2A6Na
VRGac8v2+acmOR/H7Hwy5NPNB2aEsSxTbkR/gQ/50vKsAT63va1RLQZIv6TIFU4JEA3VAU64ahS6
aulZxvk+pz+43zAGpngB56o/Cm20nPICalyEQ0X5FtHRw8nHhxMdhQXxnGr37ddUZhAczMaIvuP3
OV3vMY1Ict35f5F/hnSy8o/vGF/7xRHa9HgSWbqbYmTVI3tJOA1InCQgxzUTWyn3Wx5oU3eEGXiE
WSnX7NCvNtJYFLkOqcC8/7jMnzWm3RPn79Lf0jb2eQUZ17So51gqkgn1AcfnG+7SBtkI7YZ9425Y
ULlfu+Bojr2TAdPJn7Tw3QICE1Mld8OYcI6maeh0PGyo5pFtO8ntOx5YYDPxTfAJ6lzGnUylw3UB
RDiIElqerYrIkruQg1GT8EueKmwE34zB789DbSUW4UFzyDo1h2Z/Myi6F0WyKqbuuD8u63iMEbTs
aJYyDroJQYCeOOZN63fFcentbmaiWNctDsYFujjkoJb2DwIvYHb8Xg8Jj+T2k3IYySxE/uUbYlQM
ZgTUCIerLJssnG3Ggw/cxXP8EXMuFvGcWrbCvkvlZxJsUwp+vMcsRHLFTj5ahIUUxX3GzsvLbx+X
22u6u6q7eI+bt5ZovW+xbRY9S20cnlx+NdRe37ZnaH0S1KX6rS47OYyYMvw9go0+ztmHipflLAur
5pdmgWYiePBghhlIwS6YFPE7gXVtj1xg3kLzop3jSkUrlntWOPi5CxvTXwo9ikx1bN7lICR+vTXM
nwFoTS+viY5vPLw9gWpcORV49vVG5YzI+RAsNVxDgv1LyTXl8Z3BynG8FGMs0LihExzVrxe+VaM5
ZBc/RvIBio0ChC6q8HmFCU5jGooMfBF/JHwmZE6UFEDHwQIMK6DDWkcZ/R5Y79oN2He5Y4yrYSqx
ZmUignPSCz493uahM2pbiJ5T0CaFD9zQy563TQfdefRhjCDmHg0D//qaSYj0ywwoAY38ySyDGb1u
+fWdTbdFJ0T3OPbdr7GiWuZNg2HbMdtvRKky/vNw+4MvDi8JuVcNjwhqQ5f6fG8NPbLV/r/wXr3C
We5eS4+CgrcQ79MZPk73fU6JDn5ArfmUXvitJWQ2bKDMT5RRUGOLdta4L13/6hvQk2qiqxW8OaR5
Mt7U29YTCkSSFhXpeV0Ozj0qAa21UT28DsHprABk6/KS7bBuTRkU0XZNozjD7U6JDMW98Y/Ig8gc
PQqhsb1kkMoCiuZS5fV+gTZgFTLPY2NQJnkZaBRsuJ6yBvms/+qWm8TxDOMBuW5AR9LCb9u0FGvm
X3yJLkUv9ctuBP9CyDaSA2HSaMqwLxsqrXSn6aRTeEUo5ddCI7AR+GNkqLIOqNcwWFPUqoIZ3/cg
uHAu3+xD8LV41rIQPLpDpzra3gXajY5AO8lJVBdDTJ3qCg20uBd3sn3sxqw20EQKu5kffTuJ3QCP
5oW72VmM6XNKzZmzSJtoZmTGf/yuauJS03L6Ok4t0C7bEUWhwafFS+EClxDi0oYy7L9v+2d0W5X3
0exyffJ4FU2XzNczIcEkR0uOaAPPlaQlR0IIRxDGKakk+H/rPmVv7U13SBhwoX9HSeTP2NuZOeqY
EwBZNzgZo7a9SyjOxsUXhgOa8LXXWmAu0SchSEIQdwWE6+Fv4qpLA21DL4ZVirfsOM/4mIRC/pnv
hzONcPftG80LGyJ8x2vsjMTE/XiokxFSQgRPjCZGB2zNKX34/LZGN+aVooZjZZc00Mg+6wo5o1rb
MoRusf4VRC52SlVZnFqwyot4qaRAPTj572liKHwcbD9vaAkGGoBGHgu6mvkCAvHzCtovG4mxb1Jl
Gz7ItbdTt0ZOFUhtqLMQRGEZEp/8KCEAMJ03qXKuUtSlNPn5JXrvR+iyqtpFSy3IVzb2/XeU8lYX
OncN9HIAbHXaboZYpy+5hoBJlhcBHlcYhDHgqMcQORcUYNxoOfnu00LEXhvb38j/c+kdMfhh0My9
7CY6B747CMF2H+wU3g2FWGB5j5LweGeQWE9G8NfI9C+8utB1Y9BTeLm4QdXvPVjspLQqY63O+GPE
tHgN2X5H1zdWLC6qWcCy6k6bgCIheIWMQz+ePQ80+bV9B0zmPJ+2ANFEhQk+3BtHQYlIZ/nKOAfE
WWYVeHNp4zo4Ja4U5w89/FtcgCD80FTS6o/WPBBtSilxx9cZuT1hUgGsJrdMNUctV7wi0KNlq+XN
FIgmsHUpOPADd98KXRghdLhVcZ7gCo46bjLDhAV1W7PLCSlbJJzdRB2DxjycRdZPQXZ7aA8GqTf0
YZZEnz4XZkGs2YIEXPzkT6OVWcmGetaD65Jd42vU2I8fV0J1AID6wpeI0jO71gFykPEoPHSrMbtT
zH+kcGPyyQQmGAi0Pjg/PMZfjqtpTcaHOBUNNfu/hKGnkg7D3Pc5uVRLZYBo4gm9kmdCQRS7946m
SpQWVWOmW2mximWW3MeFL2ctZSwqRhl2gtQiGBk795bS2Ypmk6/YVu8IwIj4TqVWDe4lyxSnwS2j
XS5Ld66enDr8YPxNPMYMKDasYuDDXfSBRgUepmf18dxaibw6tG1Fx6GYx7jVhZNXGRyoLsE680Mc
dWyT7FFoZGhBw+6emRACHe4Y+NV1SKf5TyEOFsZJU6reuSBQPm9mnXzO/4/Z3xRFGZni7FtoPYrj
eogILJxoGqbkRE2emq55Mjn1nGIK8E/O5/Equda+RISshPc+nvzBFgOggcYZCFvYYL+8ERekPg28
Nb7nGPZdpb/3RWZUNOgALio+xNu7oCHdRkd0Vy0FjTSULjkodqFWmtWr5jrPR3zXdsHzXkhBT80u
jWe3cDCjexU5EYeaqpCRSe7bXIwRXa+b9/Bet8swX8KTAu/TMSHCgOLXYZpcJxJzvLhxza6DKzA3
TQJ5mQx3iDRSlLmxD+xeo6m6nUZBDvNisPrThigavufPFAhBpHsjVW25uZGhfTB7xdLDrYGIbwfW
LwxUYq6SSVVlAHkTry+HexfTX/tG44c331X0vc9zhvo6YhvgNhLRfTpRmlQmzfKuWCYXwvnj6lZl
NnJSHfmSAMloW5C5AZKiTjfoulbUXo7bIld7VF0DCLR/Ml3s2ntOef440NBed6yLQYO3WZ9UHWlq
kWXVWurKOBCWaWxh1640hXpsspNFgmM3TuHMyt0dVDbxGJIuGg7SS8bHTKerc4v/PZT+xqVb9jWu
r/uJUq4bZVxRKHE/nsKNAl3VPyrOYs1DmwF7FrUqt9PR+BsNR0pt0S7392yyZdJaQVus2preO9fh
FuL9RbSQ62j2tOtyg7SsJf8BfBnIcJEHZhToWMLiSOjqyq0cua1/0FQwun3U4Uy3aPGxiwyfLw0F
1l/xjOrCzsWBud7iAIpsKM3hoIeX+LqDh3HKApcWQdrcJ/eETkNdlavxGvTS7rS8r2flqreSnU7h
jX1LeC88NC9h9t2fotBgB8kizxfhGViX4DUsUhAMJzoGddczpodmba6BOt8gBT8hLNCbnFcCJibB
q8GuBVkUGabWd5QHf/w7OptIt2FkdDvghx3AvZ7tNQEyQcz/g2GYKMLnYZ00kVnb54jnv5dtsTsU
gvqgWhVkfh1QoJCLwIz89YHzA+5gEphCrCIdkNsstA7WLNy5zgo2LqCoetZRePVnX5mVW30FSc5J
TNxTNPk1uhlenw4iHtlBEwPzMfarDgJ6QtwPe2L9NC5fc3ej5hXdD/xSPC+/kLZ9dNYvx6uDIef2
sDZGuC+9PJCinXw3EBpaR4YFXjgRqopCoWCyv+eBikeUozFjZy6qB/NlU82U/ru8MtDOrIVY7Hw/
pMP1sFqlzW2OSD6efarEnM0CjmHSITdMScmnPDfH8X87dKys40ZUW4xp5v3JhGbK8cFnlzocSJ6c
nOZkHZtI+Xzzy0XiOuoq6l451RUinWt8HY1P/jmfrrU+kX8NZM9poKaUKiMVWH0rOr6eYBAfpncD
bebbkovtfIiwzJuKCrT+q/PNRj4nyuhyLSvwn+ccMkjF4fS9mFNp917kjXBIHZcCaqm6kM+5QEM4
zNgMew4RkpkCVyOqiaTRCBhASckD0i91AkMt8iJ9dINWcOI+VXtRgsvdvx0e24VmNtyHiQkJehzg
QzjFZtDcDZ5I4lYNpVI+Tkati+B7vpk0sKtjpmBe8lL+GmtjyRg4tU0rKZYeXnFe/9Lac26uIWnU
8YyApQbDW9n+SrANLAZOBEzt5HSVaezHJoBSRcO09b1oTS6CX7CLHISJmKDlawpLpLDgYQTbisae
9f+Q2qW8RPhD5ZEJL5IfLyVnteNqoyGspegnEO/EvEYGggXzMMoorDDRyYqe5s0MZadI8xBkXrz2
xRUwppDceC0oizlMpku97W16SrpP+/cxIR9084XG0qK9Xt1jSXDtGzTvg+Btc45wTb7wgXsjqdpL
sRa6eH2uG5uXbSKpGFYzqLI51DGlEog4ykWTjPWPnSYEgbrba72A9EETiE1AXDZ7b17mSEYQC49Y
XVohHKgEcxNWKifDGk9QMHJFNtTL+iZZ1KqigDGzy0x1eBfCRR3630iZrukrW9fyNAqlcRJ35D8U
NQkZjqCwe35XzkWJy3ezd7/0/nsEfmAJ1ARuEbrNjCJn0TXYoHHUx9y38+x5W8AMEONvHebWmAij
U+nw1iLpYY7F+b4aBHQRHEmWmn/Etvqvcf8lWojedjYvB9DrEQeZVHWrq7kl+RDQvYDfNqKp2D5E
dwmXc7N0aK29ytGiX97atOCcH6XGXicbu+5upoz/5EztfaJzBCk/WrbF1uI3gmar3SEtDVXhp0+i
CgR1w11ysnBP5nN1L5QQz+s4/b14/3Bo9XhcVKLvDXJaAnPKbnrGobDeyMId2OfBngGlfzR2XePy
MrrEBo/anoganNZcBRI0H3XlSLS5OJhw1eeG9TdgWZgzH/bBD9/+zRNfCKcL/vCsKULc63IC2qvz
keAioWJAaQl8GElyyR9PZaBWvul0enEk/kNkw3KlsSAQ6B+N+6M4+NJ1803OF1iYwvoODOabL9QY
jETsjv34U3Zg4ylkoWpN3glJcVbEn0erSepSg3VuGjmpSdjFyicYIH8ajfDD6aEklZNn7zH1j70d
qu3KMzm+Gux5oNQHcz6CSRY5cCWMsCezI8Lk+8cqYUTgiet8WLihudmHmBncmT1eBq6fWJJ2hKKI
nlA/ZTAs0e3ngtMUHn3mLPOawHSsuoBx61UJQtJC/nCwuCx+6k/ur+ipA1ExJ1NV2lITht42TVnp
a/nXiLd8w0PD+r2+63+3CeAWiC7WMAk6aurpb3bFlj+VRYuAzN/KbqrowN7LROMi6nphOE4U1JOs
J0xDnPT3E2yHtxct+qomlex/fAD3TFpsZuCKYie0gwt+vtodpEp+niKmtrXc0ZvlXJWVewAs0SVA
SMkMH6RKm/X/oasPkSPmERJQwqdujMEYtuXkGiqDNb2ndBWNvZ+bqsqkhk9VWXER7GLMidbIzku0
bZBD3heRF5zGNHZn2CL1OM5qTy1Y/FepIr1Ya3va/HgBYRuuv3lKRQMMovE1caG7Ryj/wMBc51k2
dh2v0V2KKQ8J8IJ8jUYo8wtCfhWu+XouqlT37+JohTagoHKKzV83vfjpvNxPpe7YcimI6Dx61Oa3
YfFRbQKKuu02UPy2lfXF1dKoB+xGjT3ez4klCtSV2ce/wBFEX4d34j7WoXmWD6mhcf0U93B8yS7b
9wnHk3nZOTnsWM2tyuqsJq6Qlrd505Xqcn/jLCTMGgFd3h6kXyEZ8bU0Tm95sbKosZ+8gS6iPetB
V6ILjPxnnav1efDWMLFcuDOBs6dZd9lTiXm/llV6ICi9wJoqizJHVQ4ONtJaO2+6Ozsy/Cl/ACe+
JOeUW9ExdrW9htO1jJu/7wK1etP+5qhBvce5TbjYcGeAYZK9bO2sMCY7V804hT762DEfwhTdptcM
A7IJqAu4qpLEMWjMdUCoE6yo08G7DoxBKVXM3V7yh4KAgJKsYLBYv/F3cWKJIPOsBWdbgRafjq3X
zL/CZKe95uJUF7ALMudLOg0J8H8JwvBAboXxyZIEBYH/dNkyw6tJxi+QYhp9RzuSC8+MQiN6hDsz
AqFAVqxf/FEiBCLwenOBqzEWyQyGXaW0GNNkO5PmPY1hxr5G2Pl5RHDbFuJ1YmRhb8TSdfbTVvlt
k9+WK9V+p3qASPz7LNPzg0C86AKSenyaCFPcmQL2iQ0P0Y8wEau8mbnSoh4Z6frRAOaUDPjpW9Uu
GF9e01rLyVMOin76+PaciXU0mJNvwwDYzgjhfG7CyTKE1NWnMUlUUIxKj5yWApXF76LYkyBPBKRt
NhgbUBlyRjkoEW3C8KXSHht9EWy9dhOzoRCh/fn8KDmK8PjJFMyMXcRp/WlqDc77CpSf1LSJdWYw
Tp6QOzUpk0WODS1rsu/LdUrYKcC9AuYUfJEW2P2CxwGgnYX4zxQvytxvWnWdNy0hg0DprtWCrOQJ
jA47nGVXw8rbRe8P4xIDhB0ZKrjmua+8qZClAQc4tWonCDvX6VrYQyqxvIahK0VKDt+UUfhlQs7y
N10hQAGsRdXyYEOzpoT2wRj8RhC82H4NaviE0rAIV7RTj/V6a/TI0PsN9/apV6w+pO3VaQuraPsv
kwAcxamYsSyetYyfop5px1wtW64yChmEaC/PTS2g7ca60zQQp+9pq6IkYTvt3mO9rU9OxXr+D4n+
7b6oQFkkIBYOBoMp0rHqAB4Z0E6jd2bnakjZ+27jmLiQM0eaWT4utePrtRaWWZW217OC0+M0Gwqi
B0JSHU+WCOA1mHK7Sr1aJvsE2/GA1Ibsm7V602hzGR3ZWJPwCAiBb4lEt+OAVlKpGGlxMr8fm9E4
yRXTfaxXghhlQ1HQYxmmkOsaCGwuabUbVDhgnrmKu8pn7cXX5/M2ZRt/PgQExZX4SniNyn76zxRi
17c/naYmIL/9giSclBhoH6/Kyq8guldd5sG/6ikwfBsOAFr6NxAJDYQOeOp4gdQhry6GPLnSiVaD
WVqM10Iss9jgbNxfWIEZpb479dvRmPgcc0O0JPajABndm97T+T3zNVejVRgQp6PGyCQrVJceXzcT
4O/oCL/MgGb8YCPxzYN2lSEoTc7aBS79QeGo8siY0Sk/V6PPOBWAG55l2iaXKBB4JYv8AUkJ1urT
7f1WLJUQs3tT71r79lBmdHemEWguB1CXHSfrq+79/uI/MRgGEV2wnDCTi7rxy6++TsMXiabQDLc2
KSaJJ9Raa2aGR2ZQy81VUbBweOVap0V3Jj/5eQ2rogdfejACJye/PTy41nxhcDueikABLi/91TjG
czDnStE8OH2E8HD3yvBmPnVNMk09CNAwPMI9nb450I3KJXHEW6KbS94Sp2rdmLPmr9j6sT+pI4OF
0a52JQdyxoDHXMCq2w9ZYi0pCKQOnpPoSm5pKfQ7eLuUqwIADt+XVlsUkeQgB9+SjwRigyoriJsN
5I9YDCrwGeELalgyvVRgEcgS9Joh7xJL6XexYT56ov80m5rJqc75NcFMf0wwIm3fEW8qvV/1aORJ
bs36n0BmZIq3nNUS+GAx4GJ6/OgPfnUIj13bXnRhZ95nQdsU47/77kTLW9qIxNqMbiMFhLNbO5wJ
RCCKChVCjDCdzU/JcbomKuzA3Eid/VggrOaW+deqeC64OHoayUs4YYcljYErIfDn0b8Ma97Liyeo
kM/3oD1ToLDWa2FG+OwWt9PWXF4was/oVOYg/s+fxNwf5zZAmFSHfMEXdFHS6u0YTsxPSX85hBw/
SNo9G2jJJ/J+Xf0FCjUaJGky/JlAdk/Vd5hDq7VNXG4sHtlOVZgCkWmC4aO9elrg6JRsoh1t7qNN
4Cb7zP42LyTrpElEwtIJdWXgClQzjuEcaPLwu1ts825SyGLpqoWzkOlZrUcbqAz2CF072Ek5+ijA
yfLU9ntBb25FvL9y2ozF7xBAAATDM1AI4M19rACEUrrNvTD3ry8f8NFDhjobCnlPXfU4hMe+Bh+g
+A0/cSK+KthoMM4dV4stvMoXm4oEr7vmBM0MIk21r0xKfyIOkG78iiwMqiwfG8aS8r4032h8XNYM
qiG3wIW82/dgfxmlDpGYZv6q3qHcWZSWyYQ+3amAm/ht388TrL4YmB57qUMbk6ItIUHwSYvo6RwF
GZbMtgKeCmPtcMGzoJWI46XxjCGA/+SIPWeJSsykaSZzkO+1rU/WE12P4TIkl6nck23SGqbMV6vi
VItyWzke8tO2OfVnl2RLz5Lr2tpz+eIcChHnzjsHMo/JGa3+mr5JjT7XnB1+rs4c+X+rmH8INOWP
4rRqvLxVenjZTwoe/uQxOUC/oPFqyP6FCeoyqJy3FH0ErDTdydvprkech+wTihrGRGG8nyUCm+EW
wNE7ws+DNQql/P0jRNY5mnf9mQeSct7gNeDJTB1/B5RAg6CWXbJpCoMcCqHCmkZLjEp+UVCJut4X
cwBcIfsEbrDwuTXKKuamPtUP27L8X2OlKrxj8Am/IJ1fSOfbrn5OkdxVTlP1LjH6tfMsy11zmyoA
R51iLzC34LfREI2AqFypaJCBkIgUrJJVtDy3Wrs96ED8cwhxQ5z73jsEtQcNDlSLYixARaN7FLBT
1I5VLvDrS5Bt7OBFC+Ll5K01wCNe/uviNHgWGpnvGiOnHbKceyV7P8g768EtJZ99wfXdjsRdYnQ3
4dXw04fNepP9qnIGob1kS8h8BZbyYCjT9pvZeLAysjocXDXnLm/jHaRIrJRgVdScTqX3xuhsV0h3
rNs7nkGqt/uy/ZIZ7IXPK/Sdegs13u7YSjqukltU1g9OKuVag7YiNIhjZG+e1Q7ntEdx20jU+8xp
CgMnWWmod3/QEWj/8d5fuBQXcvMf2wzJjAI/uY1OaxR0gWaffHkK9Z3xpbFxv+oJEhHqVgBlH/Rl
ozR8EM/DvrFbMwppyqKyfSjApiCGYwwyc5pOQh3THuoY8by3OVFvLe74/TzLtWkefKuLjKRX4FMS
K1gJQIm5fXdpA0KdpQDD3OWlsb7Cf8e4ndKVCm39/y12J6zoXePyyLjA8kZImKwi3RMcwSeBhHD5
sP8EvSgnUOqm0k3QCGm4S1LP7REQXaPiiENa4dmSMbvC8glQs19+xFVKYYeLKRaW837LMTXIx89l
5YQX9UoCVmabT49UAhc4aBJGRY+TB4B/ZnKAzK5t3ni+SGnno9xlxcWFshiv5m5cZcBuTeCQbbRF
lIn4yAVbxxoWi/TpHuD8fAGcXlyskLgZHqIq/ou+sLRIYwX9ujjFpo3cuQYXwfSXGwKOOaREI5lt
E87M3CoKGBKhN6WriRywODvO1sOxaXqh2weL2BnlLWFpWE/jfwaP5s+Q7COAJoWryKbtWV2Y7nQi
efykBZYpDfmbY1cxWVbT3b/jNDt/Vql9fL4WRAo21Dba1gxM81wHX9mzqgBjRA3TB3yk41/Dz8iU
OYBtB5hB3dOLs7cR3ZkfDvfmC+BtcSBZxo8W0lhfXTu1ob0r7u0JoOyioAp4fh1QyAdeR33YLoyB
qdpbCc+UOUpymsk4JT91Fa4mBvJJEL0ih1JYDPrZCsGWWNJg3SpZKoK9UeoqNPqibs2rbtKBkD6W
ucJZn/w2ziYuIAJJeGZMp9SQa5RhrIP4HsyJdFSdR6XiuNVci/KpWRCotWX8YeJAYL3MRtEHK6Jd
Ped63fEVaCPEU4lCv7/vkpTcMoLBHRnSfCEPKkhwxulsxUo3mbidzIpqaqzkkJoGGWQoQaklXr2u
3hS+WGEY1dv+fFukaXKw1XvD1h1hm4yxu0DebC4SVJ0KYibrBOMsY6lTLSy7u+QKJ0HiJWN5pCee
VL713z/c3c6dphqL8j8eOGI1J0V5VpdQMj1BD/Cga1YxbfeaO4OKENQbX9vPzIiZScVP/drNH82/
7gcw5FLlMX2iG31dL3BXBCPMtRxv4dRNbbO7JqTBGrnjO7qUTUlq+vZXiKcYCO+Ci9HWD22JdwYV
kfg2L8xyCXdpumWKB0ltwOj69VQkUlnndiXpnE4Aqtez6MyMNiqqT2yrlfkK4JlD1Xre1ZSBOTcc
YxyHhETNuFOpZFmYVLfqjxM+SE+fXL5eLWaIdnw4sTvVjAXPlsIops48w+xws7GfamXDTTw6qHjG
1CBsW3uzob5bEwLmSdoLNLkqKfhBbahRXvrQFE9OemIrmxTscu2SOq6zYNKMo8lDI8dyf2h4l3FX
to33H5dn7DPFUH6cpW7Dywlvfov+iWo2Wsu8NM9++tCKcRAFYnRMJSswqUDwh9Q/wImPtX6GSVv5
7E7OKdUzP9nWef/Nc7xjYelTGJ7+/2r5+eff0UzKB2kfkuYC4n6uu3uG3cCfqFbMoL3S3iTy4W1a
wyOXWquZAU0b4g5GD4gMhJ5+qNtnj/jdigwSN5d0mm7Se57nChJR1HyCwXzr7HQbVjjZUwJCJoz8
EzO2zkPcIraVBIoZP0LhBQuC2yNUn7uQBMPWkIZSfxFPzYC6b0r1vBbjMVTxuj0Ja6K+vaFiTpWY
VXwy0Zp6ef71emzbX70zTq99F+dmmCEmIP5C7hEtZ0hDb7WvHDtZzM4HpVDhqUNsk35zpJ+y5Sl9
p1537bGq8i7P0w6Y0CVtqf45yJ9soi+LUf3x2oxDzCDlnf3IPLba1A5SItNO4nYonq07+qSl4hIG
piL7D16KmCqpipTikN+JJKiG80rO51a4sAExorMQPH7lfBmxEi1U0BQV/CEpWhz0+KdJjq7QndgU
19yIq9hQNCrxsSvDLrE9s36xUP0Uo+JwjzmkVy3Sokofsp54jtFFtl9mCZdXoR8Fa5H7Mq9b7C1M
WDTrYz9F5Had0ap+98KOYwluzWHxn3K5SR72597Xt0vqjsU/vSW1jqve3V6BV6AX09NGMCdfhRi3
+AyNpVGvGQbm60H7Yfc67VvOWWY7p+SLPluvln01HLYBJgIjWuDAHxsY9qiXB2Ohnhf0JaJL5W/N
T35ah0hOwMyZy8GiRNXp3MtyiWX0aD+X1+5r9YBJDiyOH12SUwjYrqOiax0JVxh+0jVSZa1p83E5
6lrExOis64xqkASLUo1T4hamERp+3dMDYBrovF2UQXdSvyr8LDgZkGRLcrfdOwZGhHumpl1m3++b
O9WlR9waYD93St+9mIVKM1InuoXmmDb+zau/EJwyqRyXKzvloy58UFtxdddyn5CscdeeXg9Cu/Q9
JOIerYeJG18wKKVo3k0X13U/6W5h+pLdL0TM0tgLnNJwArvNZ7AQa8RR8Mc2DTeR1Flkf976Cxm1
03j8Mi6iFpM411H7bOPzsCs3Iqrw6MNWiPIbYEZEc9oq7q7aE6cyLdwWL9kOWztwzDBLK9OH6lkb
wCqcGy4g6f/wQTGdYLHxZmiQbWYFiWDLwVxf1NmZfweH3YDEa11p/ZpO2Uv+t4t5EKOhh381Yw8J
5aSqw+Bfr5pei1ATQzYyMc94770fv2hyq0jQBblLk52HdxSeTqqIGVr3giXj1XF0+Ope1NcR8Ngd
37KNIZkl4P975ZPEzXVKadrT7v4NtQzxZN7N4UHuGz7mJz+OFucM4iu5Q32Ji6dqmknhppYcuiLZ
oXH66yULieNH+HYlbQGTQ5fo7RJ7o74NEhxS6eyMeZEBZ/+d6UgXP3CMhziG7MNpHr8vWrM/zfDL
yu5MX7gwiNlekbonyOZ0lV8pGUsMN+qjwuGQTUyM4x/z9KUydRpFbxnan2iCktRzc3H0ZRU/W6vg
gkymStUJQaw/b21ZL0NaiAVXAc+FgnGPnv9IAnyInDBvbpdor2ab3kMXEhxvb2ZsN3TJw7d9RLoE
2v8ekWMMK5pkedH/QGQSa3nHcAXl1/JxEZCSTy2TCN5ViHu/XSi7Ha8OaJ2RzD+aVZe04PiFQP7F
se2tJfM6i81NtkqfvVf4RHmxrObkxWfAAeoTn8WMre3sakt91BDym8JY3PGWGuIBvOBUzUKVfDO5
FU/M27eQ8hhb3IDTGMhf2rk2Gxm+pTMBg6GPkJ4Xs9Gv+6Ifu8jC1yImGHwwIB5746Lt9THw7E2G
CWnp1svCf7SOFgit3wQNIOmmh+DKRpB6pEM8iSjFQorIuyhS19ZGsIKTMltvmHzgJyUSJdZFqTU9
B6ala7MxRhTHna6/t2NzkLr2P9nfphY2qcnAmdKCEiRgrsLwG5LQgWJLyJQagTigFuPO2StCDbGF
EqdjDSLv++CgSf4wyk1aaxfHyxWQ/kM+b+EoG1iQZXQvnNwtgcPXyQUR8A5tmuYazEVeV+uOL2tt
SlVejv3a4DXBdzMXR2BtHyVXfY8Eamlxk2jJYH+VUela6iWH+KgpRYgXEkLTyYw4X22DxLMdy1CR
/uCq6k3gTnHZNBcW3bx+FY+c9rcrO/jyaKSDZiVub97Q4SrTzvb5vvTLM4RuF73cu3R+NW7bfchq
b2eXfJQd3DcJTMX6v+/bBXWbua3mtD1tQBP89xiucGoUW9BF8ylzsUGnsIRnf0RIX9afG0xuFKB/
kp2SSNL8VRo0GpeNAkPSRTaDiZ9I/GzwNu1oH5FqM4JSMKyJ3RG79VlKrlRnGcj9HAIA44ufhzWu
0vk01PsUzIIrrsY3dWY7ZEK/DkyHhUcmsaYGdMv0Ndy0p7+/uGvHM56L2+2DUkh2ooMF1hw2MURd
GeJBc3ZJwCHxnJQoJLuh7boDPZc13S3K1pvm9BJq5MnmzQp1Eeqca9rQlHMYuiFYAMsTIG2PFuEr
gtj4by7Wlp+xSHk2sryn12qLfV3fhlnRJh0br93rTx/+3vmbaj0rSWdHL7PWM/M6WL22D4I+blIc
LBdDEEwqg7/1F6kQjx7KjEtp5mLrMA/bRIK2kDGZDqyk//cVUL8MWPxz/EQO/r1ejdlYpQxxiMBS
Tev2cR4go3+/YsNHSAMOlX461sXpvH1mIYdfTiD3PFGwTb4FrARxxmCSpA1EwqtJ20/Xw0oulXLv
n2sT0KopxzN59WNJI/NxzUWq/k4CQZvaUlNdCkosmezk5brZMRKOiXozA78JTclhAakhrTc7+8cL
19YZChaLF1PhqMgtxd/tImF/CrJiMALbil/FypnJvn+fFafdY2S7evT0irTOGtoz+2CGDfPHSHp/
NxBjFM+jiY9FeVDcNdxekcglPJfoxVskPO7jFJdMHnz9qP4lmpcI6qbswCavb+GJW3VX10Fdk2s9
bsoxR4rvC+MYhD7qt8uFabWt/f3OFVvpMa4Vo1hFmCbr2AfwWYKTvQn7qR3p7q6fgFWnQvmp1Kua
DZyO4rtRU1kYOwLg4ERb0DEMCiw47vxDbwXe5V8u9b/24ruAq8npyqLR9JjhcTKvY4OEAOkLL4x5
rj8ytWPzofGuGr3la/v7oYgZuAjGilaCM9r+V9wIqzJhqtA4aysgfZAowefXXvUneNFqSeUhXaMf
4KCq7CxEdcqNuUHlWsYBDKi3yAo0VS4L5yeiUcXnJbMMFPrAy0qZGCAhz3fSamjOqLi1uITTBfv/
fD2xqHZ5a6ok1/3GBaM2gdPs196AQiBHgD39iqn6TVm8TAAh+Xdhmy0Nzd5bYEUzlAtShNblPgEa
bOepNPsaGPmrb1GgykB4cjcOOi45oqBirk6AIvsfbb3sGCGxztQoTV7XTW1kOIoV0/V3dXvTW35C
ILUmNFSOrTVMKD5knEk0H0lF64JzMsFVyT52FUy0M6tGH9TScW/1OdpYAinqTQQesSJNh3opXJv1
9l88dwONm3T5jAuba5uUY1fIrg6uVfIpCptn3YmYFZf523WBoOoQxpckaK9AWbnWZ9YC4QCekDFG
uqttcM8jgqBVEHgcy9sP96Q9a7PgT2P/1R9Xns+Cg0WQ3Bk6uFycEPcfYXfgcalgm/1/50icCqZC
xMlfjIJrS9bxYXdp3kx2yqu/ms75KmB3AS7YlF9Kze14k8kN0nPCt8A+3fNPVVpyURB/P0OQyttb
GLhTBB8kMclxSBdACsVHzVbJA2lglZoI/fDhnoPRCIQbh9x4RihMbpqCRW7oMnZfx3tTLRR8QM1A
BnIuvA67+Ic2BqePWmtgLp8gwwyFPZISWMOi6BVzKGmwuRlon8HM3QhPSzxzHdpV1+zTiAI8fQrC
KfLuToxz/KMUYTnwmJe620C56Ju0MWmJhjQulPNBArq41qNlcNgtMc1UfNoNBu3jUtrV88yqRhIS
qeHKxdcx2b7GvMcy9DpRcifn07+85ilsO1H2OF8EMQTBTzya4H+u2IOxqtDnKyMx77+EdFg1i8bj
rrqkwWEOlr9JlghJIBi/jZqKaNUlrB9P2GBgVLUO3TSOIH6FxS7gj/85jtI7hOI1NdaBq5QgfDh4
SIMgaIDd+wiTl/uyAhYqfUsGmNx4rtetHNwfc99+2fmbtko9JzBVibUQ5Fb4DtA2Z9ZpCJLCExfn
EIuuITjpjYOq4MrLCAcVvS2YhyRm2ZT5WStblQAVfzg02SIChkNw+2zZIQ5xL9JQc9r9YobNUjKM
XoaLQNlrqfimx0LifOXjDCpmYHb3lP+HqY5Xk/6P0lm4wm/IjdAUKrGx3JbKahuc+EqTMj7tkVLX
KxNZL57ITW6db+ekQfTzpgvkolgSWwZTsW0XFLzBmF/gF5MGRdaOYtfDHuOyzuucOxfah+cuZZh1
dJsqreCx2qpAmoEThkRsfJu7mO25/Xpj2ZvAT5+TLq/MruC4uzIS1OzB87AoL91Yt5y5hYpTkhJM
65aG/w5zQsJXMIPbgh83pIRNifOtSZ+ozRUNGRwFNgWWq3Uzlhgd/PWg5GPspA9Ch4imFhJn7LIS
NZNgb9EY+gdxoJ+TMZ0kQzvWu3KKbyyedqkwm/j02j4jGCQrLlu7bDOdsJg7aVur44xu8S7lVxuw
vMf0FfkVTuCpvIstJSqDMsMJBMb/Kp6+bzBu6uQGhARO/yqoZIbbvETBa8btZ5/R2RG2GHMMZh49
B1cczHxvgpa907NgdgUoAGwOUohSJPPtevxEk3gj8supa6Q0Xt4vHIvL9jbvGw2NWSwBD4aC2Cn/
P99fBJr0kJyeRqc7PMFmLGgpRnRgDaNeABzgC1vGppQCvhiE3Pwi5pOjbGhsAuIjqGfqVgjBNTkA
YNlRMt1VRVlwQoycctvR0nbqFsrvtv/kn+vDlAAdy8IW06AE9AX+n3No0GPHM2rHaTopNIwJqk3P
qp0oYeg04KnW5kbVMpUY/6rOZYqlFjej6exW4RBwsszhkhDh1218db/D2q5KlFVI+UE0h8BkFdrQ
vprUq4v3GNqJ3u3DtNhJeqVCuKasOgSd3UZHYeDN5DRwdUy5ovGKtkWEHk2TJ8pyrmASRsraHWP9
Zl7wvG66nqQw11F3wS2m0oLy39R+QLSiCj5RlVjyqsknDy32kSKuzADVPeMdD2JnxclEJbD+L+tp
2zuRBR11omp3cOQeuCzYF1wVBeds9J0Wwb3TjkvE/r4UkbHjpYjBRDTZdufisVNs1Xl2q6szg9bG
HhvwbfIFk2ojui504vClckCzx0mB3tfFqlndZrY93850hsvF3k3xqJ4UiFh4sh58F/3Bs5yws0jm
gEObNjRyeMjhjGCDJRHK/wKa8tfatkdCrGK2pm0ZSi4Klc46Uf/RalSz575vDDq64Vzy7n26Ez5y
czcW4I1lzzn6+PtAYz301frpW9XaJkflJ8l3NB4ktLKLnVu1FTB4YAxq0yGVWyyk94nxRPMfo0yG
WJWfxps0Je0Fx429S+CGvMX+kAjgZUrpgfwEc5zSW/XSccqzQuiQHrHSkyV1l9Jt6/2EiFRsN6a7
l2chun+dF06nY5UfXFwZbANE6sLTe/TcSxPDWdZeE5AItd2JAYOjjiGJmHOldeWQ+iEZ8YGXILLs
3jTno+REnoXP8Ru5CRSf7TrSfy4hcRoJfEGNDbDFFF0vRIGM0Az/V34+LYCrzjGiHr8Y9lCXWOr6
ZnIJ/xheEGbQNWN2hbsD5eaOp1e0zl2LFJq7csmPQD8I21oaVIKNEueHpOvaDhYS/q07W7rcb/H4
MRtWpQoIwYGLv7AAtS47j4Um5eDC8F3xUtbq8pBV3mljoKhZNdpiFNDNsJipALnZUARtaQ4GFgY0
x7bzw4W1EjmZfAtKg5S3YSPYzlfWIiO+Aq6ujlaDOgsrlBap/1/LueI1lL6l7akW5O+cXC9hUxrn
Ad3FTo5Sp5qRHuXConkixqS9HI8ZFH03j2Ze1xBc72A7nuSjiDpQUwF5OiHz+2UCZt2RDVyzkW7T
oBWw/TWzAgqTsdoeFm66QyW3dQOuIwSl4Dv0jycKzt4CPg3kStDyC68bRRsuDhGFdSSfrnagciW7
qsbxNFQ/QEDbgmp4Sebb8N88SNmsXmMCZ7GuYSI7A+15NzrJM8tg55DAnEv+9fZkMhE9SzE+K47X
ddBCfu8CjjBwQUoiwvzSV2orjhzK7YcV8AwQtxn0VTCp1mw7RNxio/NHhpcYJOfX7Z3OXtle/bDz
x/OhZodX2sj4jvs2B+v7jXiyWnM2MqPkNM+DBCwAYm2p7F9EwykEzwhnDvRfstLtfwN38GfEe8+a
YoxMp3LWYI42upeoqItGaCcvTA4A/KU34kr4tU6WWSPQeHT0X88/vBvCviIrkoZDT9j4rxVQ0i1/
kw0gOz/J8vM6hWiyeUqniqg+4Auku1+sXgMn0UW15xtTWTigJ3PghJOWhekttdigDHtomnUHuwnL
9jSYrTu4z8KwMJ/FMDGA+x2H1V1VIpTM+wzaW3YPjziblF+EUEeHudTOqfsaGHqZZ8J1boEIT54W
vhAJqJBmDX0a3khg0fq2KGy2cjamrZTss70GdR0xjWNGlUrvEa1QVsqJVXE5cnvnkWOhaXmFiymN
lSNY/BC84btdYiwKAefjfC1xykpn1M2/dW9PcuAKM+kNy7nsU0518j+JhSfCfp2Fe+K2Edldjmm+
RO9mPuoMNbeWMIW6MeEVYxTuGJoEuhxt+Stt3ejELRagxVUiuSFpnHKhJHze5sd0yQONu/CvXXT2
JMkFEdtVHGPMqMNO0136mEyN87ucMhig8G3RLsMZaKZ9pYap4aQ5eDs2BuWDlbagk+NM+oPAQ9tQ
M0B3buxJxKfFcaLEwmqNh25wEdfAda23+r2cK+xtvFA0EX6iHLra80h0ZuYkeJkJTbrXx3uZURXY
JZvtaukS8zSesfdkUuHwmkehGPLyI0nW4G/YxO5/u+FlfRtd5EhFrdJeh8olm1D3qKylrhhagdl4
kkUinNTgMF5mQdLPnsfcA8JHkZ8jTGTFiG8oraXtPAQMvZVVUMQbTquBCTwUzzwmjBGkQmIs9rkk
Qb+DUHbVObF8WLX6eNO93k2SlgS1DBkG2utdY53Ki8TTk5XpGnsKS9LA6Y8MJ7cHZRR9C89q9Ypo
/XPAT7Zrzdf6GpnoV807qi0s/qgGJxkftLuaqM/CS6DmtGjCUFnGfZLYa1rFPfiNJPP3Q3ZSFqwU
jPOF0OLmh92Q3rdmyXLwo+GGljI/XDhRAEYQ8S5+C0R9DOXNIO1HHiMTuZS/1hepUFIAsymCWXuH
e3yNn9NcFXGgfK4aJlMuZInuIOgsxcDqUAYFSwKs7rE/3aCk6LstXt6hGl7LaZO1DAPcwXQ4wPR5
rKEq44xoiT++fG1rksxz0Ox9UgC1HwLekwDfxyzC6D8z7OVM1aPZG/ryGTn88AvDliDxWiYme/aK
1yU5srEEabYrNTFHd9E5Z52zfbwAAvnbhcLSGmiBYoqscfvb4Ty3UBNOKFewq5M+CtWgm2Q+Af2l
WkS4Z+us5tBaME6Phox+wCTK+joBmrxFHNy+uikpDN/ouPEZbSPlLZDQpdk2mPJ+V7JdmcRVay3a
jojBPjWQykeCvKc03puWaMBhzcnFVg61XChO84ak3xxQkGJMbh8QmUGUwUBNd7nhsy/HSJEwc2Bl
CNU1te9yqXHODdORbJ8KT1ns8UQs4EgLpB1cwVeHz0agTXADkaI4Im8a0SkG3RymxVlgg2dOviB7
bC3RM9ox6peKDUJCpvWsNTaeZy0hDC4bJ11xkyO2wUpNYYnH1jfkqkU1knj2WUqNAtHyx1bg6/G1
DJcURykcSWDd+hSVw3cklE6jvgwuHsJvZgwuoIUdN3rGV3amLV/AQ/u6+spkyWIEz74nxBskSq0+
yIhGD3CvAxtVXKweScoAtDo5RUhjyoDsDr4U5f0smG9yygF6IXx1ezU489o8CsNiBY+QIYKxhwsq
j7C1EKSdZmDsvQs2/0+g8X34+clEWOyo4MTqjl0rr1Gk7hcUDyDdS3lbBhaT7TNuymi1bSK1nTZi
BeDkd9CaRphwlVEWG5UezYB0YuCpJcboYBdSSNhKLCKnF8DTOI7YtdOTIzjFVzunA2DBz+ZZ2TUx
qrNra99LXJX9DGQI1SYNOiHhzZDTIZuOqMIe/GyHtaO47OBIoVtaqPY4GRb3Dbqirzk1/9eFlaaK
6MirXXhqzcMNv5cAEDhwK0ZrozBbTG2hDuJZthiMa05OG+1aMyewycbQiLuZqArl0hjFgxKqzdvL
RRukpGr+4u86zGQLg6tQfRhBrgfYMXj3qTOnjYf9WkD94ZH+puRL1awMoDGHP/FiQOAt2KogUsP0
fb7AkSO4mWSRjIBwBIb6vJETkxgvYj8+35hjTTPMZhV8+2TOxElHXTTcu4/pVFeY1HLyo3ze3DQ2
bAbX846c9G+eiGJsTVF6jQI125K/bL91RABtCpF0Z5sfZqleSL8unDZmOeolRBJFCs+u7JT4orBP
Ti2rULVwcK15qtqDppnfa6qYFjEg2Jh6mPfGG4V2+FpH0S0aRjt8kQHYXIGNBVasG64+6xUE91On
W8iuEliBJxLmsQXBOFs5wo3nT5ia6WVjaHkmlo3G9fOlc65gEHzXXp8hQJQ2T+4v/R6diUXdAYjP
7JCAkM1dMOQKzBhnA2BastIFF3CeOHdkJqeFrC9gdbrsLDoNpQ/J8okfzwwSuhIRhkIxKwOMbFIJ
Md9mKHVmNsPbeN9evpcm8M5XBEQwCRgz216ydLdh8PFrQuxsxS4nA3Vi6GdTP/4ito40C7Hml2n0
gUU85yJqyDUw2lO87uUBpFScAaT4+ej+yUY98i1/Th+6XNnPxKt/BTmwAvcVmSfa0EfVNKNIguc2
P9yqFJiXltr7V88EUdGACLeu8pPJXL5lk23Hl3YNT138dJpAZ2e3Q+pXmp8gUyojftNYiiKhanyo
SP/nM3/PIJneRNkiWm42euAhVr2pPEhXTxG47S3EQQS6PixFPMMZI7ghWYp2JJOUkoH/nCr9L4oh
curw3q39LuGO3Gp3j/047NFPQ5MIi3Pue6Pn/hIGqcdqHNpTi3QEZOnxUFl71eFmqygerKSP6sOL
qrvocdbqRyyfOEQqTzmFuxjwbnXkaPngdN8cq1aOtCIdF6DkTBD/+xBMMAbtt/86oI1BjdNIzC9C
uti3qDEuQvgYu2OZI6DFV47aTo7HFEEJhFM+LMkfaHJl49zgv1fVElBGXjOYpxQYJpOV+nV1EZM5
FlXkseVBez2FyrYkpwolp6aowQdICEdzJEJ6EU82aJELWuRh2mlB4+GliiKS80alsBETNutVFI3R
qqFxG7CpwPcDe3tgHcV7ak1y7itmFZKwwX5+H58Ba+m9A4pl0oqW4GaaQ8LvI9/OUwFqIQjD+pOu
b8D7NaDR4bmy0FcsLJ82c5OxEJpExOm/fu3tg5lYBJQ8qxWeS/T0KnMuM17PzP7Row2I9xF3/Vsh
TO3TzpkGpPEPsv+j1cquismcfBRLy+8R1dzRXmb9MiZjdmrtBdHu1gHuSrlMZJ0av9ZFp+M/CUCz
HVbYEoEX9zvwCcyKuVpecDc2VCD4Fy9Ry5yeC78KTfvl249tKb5BdcNmhzbE8v68n+Vw1vOQrkBX
biyVu6jiBUgQ1y06ke6qFmJmPggTQP2hBferrW4Sc+DROLVJ7egwtdXSqGqxY20qYE7pqPAnTTvx
J3JNf3jrKCR0EiVL7EVqyTgZN3RCGbVmUyBLY02po2Vq3l2pAk0nXGEYiPTCL8AbICore2GCYADs
r3KKmn4+kdLtXWSXT79bjnwWRvFA5pGGxxUAtXYIhT/p96v1lLfEiNxsoZDOZNN2nyXox0E4qGIX
SbpuK26T8wIsUWZRPf3cLGy5Dx5KUTmLqwuf8QIrvempZBIOAPHe8GJPBPXeXLWirarcJlZOtgeV
XS3y6yoBBaEuRGSjz9FdHA0q3wadDBAkXpwxOsGbxCIvahw77t0I9+XNFKoT859F+UOSXuS4T625
jgE4LQ7QYbdVUf+Q74rNLY7xhFAb9nFmybhkGeQKn8SKSib6W4nmc6s/i+s0HNjXJeo2yvTdEUjI
LVEsLGx4NdJsM+hEMitR7z08jo0P5YAbhG/bXZE9RT+kG0gzo+TYYXJuPQqdGjg8wh83YjXIwBqu
Cve2ZI9YcX6DkoxzyY50WDLiloq1/vpI8gX8AKEVKk1Ft7GyP8ifKfx2JDnvBfqeef4BsroOpp+4
YfaWz0FR7OFDv++NhTtoncDWZ4EEigBj8oOI4sEyF79noYMunt8SIuUfs5UtwWhZz+G6YJluUx2v
yIiMzi7IuCZvNqoXLHWh55sUqEXYzaw3LuYiSlgnZhEp/u4dcmoObnq+6X6gDAwCbvfk0/fvEKus
op23VGEj1auKMzzOUAlzPVlo4Lqzkui/GMoEmBn6ggLVblBI1ApzB372atZ5qBSweB/rYMVJ+lcj
mMgGuY8WTShetGcLcoNbbXpT3sdbqJHET+tFQsXeN+W8d+KR2wyG1awI01y8EFm0boj7sO8aHr42
otL3F1tzN+hqMfk0a9Trej7IU9X0ZDJcmkUiDVCAhsa1KcaA7pC5/duv5Y1+DjBnQ/sD3gwxlTLG
qM1nltfXjWoNY59ga7vNFQmCLo8kn3UQOrcfK6Qz8N1ze12t2rHC7i1Jt+qEMwjsN0AfvbPhc/Sb
QC6MgP78gJlwS7IGryzKUOdi8seHUinq2e252HllL9zeCEPuu8rlRt1GIjLEHSHxZl69K7CDEHDy
1gT8bc5ltbDphLBu5tWHNmV07KDBng2+1xyT1FlFnGF+KMlv0xK+i11sqVOmNHP6R2SioTJMRuj4
7vHHhyMODr1xpVJYpM61LXTh817KHuQ9oV3OkXaYKw+z7GwjNZPT7hV53rg5WiYCTfDxsgnycYUm
AilXyRuEBoVPwiXnwW8W+i/piCeU3HE4b2XE/jNnr/G69siQZpbnWnVCFpkPhokFTngZG/jK6/IX
s3TOlHHFljlwsdGnucRyKfIKPTf83cgiexK9jGccf6MDz+85MDYymZnsMvIPoccSJeSkHMGpEXKr
zF6vH7kpK4BXCsBKJ6HMsmJRDic0KwzXE3vwaLTegp2WdBFWiYfZVeFm2oV4G5+HyrvTi8/gg1kL
I0fLMsvREi3OFk8Wf07EAwNePHVmBtDmoFLWz39Q0TpLbWgBRVY/Xz3ixZPmDbZZOSA0gWT1Czri
QfFuGUegmiGWvCr9P/xHw8WyN/3ysfVf7Dcq5rtWIayJWKyVlYLIL4QTnNEGBBfgLX5/q+Ux7t4M
xjd35FYqteUMD6M5WnxMUQoSCVrrpFbUe2dte1cIPTaJKc3L+Mp0OAOPyM3pS4U5WtFWwk8F0ry0
DVRaHwRYeh62cxUXhKgK8dBZ6I0CTwGFftfR2VbUSX4Ao2sBjhQz6w725m4Kb24zhi4Ys4qnZcYO
8tIHEK9PSZDLeNOVhn3dQAp0FXURG5EGuSywvexxoUTDYQU6/u7eUOH5zqHv5N293ejpxheJoi9s
gy/uS08Am98i6eZsnShBLvIt2DdfTQyK4UE1VpUEixs6TXbkzsP3cA78PEPxVyHILmZIQO/5ufJq
1/aaq5YL7Ip2TAfv1fsSVb3Er6IdmAOlJHtr0KJsDQ9/tPjd8RPrWFpmmKvK+OFgI59AWvovqY7n
60jmtWht8brfN87U0U7b2pxcf88Zp4rCbHcPTxzF7MSA9QAU8sZlGjmJp9rLhDpNgwqPaYeqnLGZ
m5HF+IEGNgKazkHb1MROLFpzGEyPP+xe6+xW9XdcNiu4+6jq2rhb8ncNd1uP2q4Qc3VCZbItSjT4
h7D0KiS+BGJAy0CkQz0rBsyJzMrSHEqRU+wBQk4rdiqykWPG4XiMO4OBQd55HVE4mwOxTuQK4zyz
klJnp324nAxdE5WyIiXhm5PXgaO/0z2vEijQDsgPUzCJfKkkBS+vzA4o/9jlxsYyp2GI6i/bTrLW
YaPNNM41Qad6IqPB8dByyqKPn2qM6oy6eiiFmFUbyefSEW7Qd36GSuVtc/+y4xECLsPbGPMHmfGs
r8CyZQSu1Izx8Xuw2yveOu5RZB/VWID0pw2CSM+Onu7QImSngGFKs1+7tJ9oLL17NpHqTVL7KNQn
A28JO3yZFxJhp+8rABBh63YRjM4qveCSHlwRLCt7i8MHv66jwnOmIcpF+Pw3QfMREG9dlOR0Qt0z
mLgNaKHUkSt/qKfHXirxi1t2NL9DnIRgZbP8G3Rl16GpEYGE5xLhKIFBvZgSd8tSasEaNYo69iub
qJ3JDH9oxye4Jf+VvjaNsNhbM17NPvOGKicyOIPslzzOiVQwwIWA8h6YEqMlQt4R3TcjKZHzIo2C
5PbR/SHFpK53BJ+SpYXN/WjcouAW2n0aHv0rwYdsWkNIZMEwKrq5c6bFvzEZEAMAisdz16l/mHfP
l1BXqGbnzAbCmcw/RMdXWyOAqgAmZByU0cVLcedosE5yuD0YZ59KKFzQfLR/MUXVHfYm7rvkAaf+
05lqtxsbuv5+KoOLAkek2UXhVfVdCCoyg5t8BUXNMkagZSUwsPdZ1rDAOY322/vmzXrhQLOyV8Jc
FHtb1eiALY0bIXMl3aqHXUtbtWcake8Mk3us+wCn9GjAqyfv+fuHJyVzGRo/NnozLYroXoes/0Qr
GHpTWXBxVJlBKPLBVq4MQmwR1LlfjVWDau82R2xeOkMgQrS+2hz8MUyP2vr3aD5lg8hqVlCKv7Gh
nBiXFL4ZwudJUdmX0AbXtogLqqmnJce5ffRv5kbUMT9GrbImsJ8OOj7JTA1bQBXiamdO4CKuVBAI
w2HvUcFxjzQkmHbBe9ySXFcjr74s7JlaaBFCYnXHXuHVWZ8Rhq3U+CtmKAYctmugLYx+in4wRhc7
VS/tQmisGtB7dW80UyuXV6rKbc1z5jRtrlUWNIQqc/BS4ntXzb5CFjqMfNa/ts5iItRFokcHOiOf
S+yUBvHS3Ffom74SbWpo/h8mUBgJpiYKvh0AsV3DzqMnS8RWldH2zAujIleJECyLhykepD3aiF//
rVTdamC4igRVqviaWi7rxcMSywz1Vy9U6RUqANPdFN3QU3pYpQFWB/dzwWKOUMwt+YhdYkimhRFy
E65PJdDdx1Ct+LAIJLrYg72uP09h5mFMIqBL/a/XZHlUppED0h3IGApqjM2BU0QQKhFKo0olWyxZ
oJvR5Ifinfstzvp/7GoWmZ8KLWpOrtrS0Sb1avViR4vm/tVN/uuBARZoiT5i5k/2mixhYe0kghOh
ttQQxSnAZ9gZg2Ks3XL7oYQsve5oW/Lb3z/9kbQUyb42i5vACBJbaE6eAZWTrFDfTdeia8e5mizz
0qES9iylfcB5VR9eUvj/LWEZBSSXOuERkDPlebMNpdAnyNh0YdT1FTGthRmntxC81oHvIlHQZ7L1
vgu5IwKbAkII4d6KskDgyLo5icnfJfhrkxSZyQyL0ASL5CMhDuj2Rfp9z7v6teE1RtW8ys/CjBFN
kiLbvwxItrhwE/1iY1nO0LZhz/cHxowjbgSX3s1MjGBhQWcV+fYoIgPTpzg81ll1jnDu1qrFxfDe
onUBJHncghVwKb4WdHd6WuVGk00B/6LA7O3JjRRVZrUjcnyReP/5q386d6tr6+5ssKm5LjNM+l7G
mSjoYmvXxaz6hNkgRPE3CN6X9t4I/KBTULre1QT+mHInnazSStkHD6rNLxX0ZM5g+K4pBqg9YVGE
OJdixqOnADYfaq2tQWT/u7IhX608rXk1EwgV9ByY329i8D9obVqM1EBnk6SeX0oHH5//smNZQmLs
BdG23MrIcPxJizjLs7raxXrxolNcbf8i7d2SveB+pyKn3qLUJxSHgefzW5FEId6bt8MVLfLcpY0R
VwLOsXDBQ9ktMphBBJRP4x+BYs7KRKGkcX0opNl/qI8fmxIoTG0GbyGHWRI5N0d/y00yT8Vr5hei
hvF6thHzkAxvxfcjVnUSPXs49ypf1UV/EmxI6AFmLM10tFidrS4Ja4obRVZg64gTtMSS/HimTqnG
WC89vLg2jgQCqkS7xLDQJI55TMkLHuTJQ+t14/YxDoL94TiEHQ/DZRBPydYxzlTiMWLz7WsIu7rB
/jzKyqAbmZCCwAY/SfWlDNbk9gCKbAjUzTpPdYH04xng/7M2OT4oHcxxIVEUGelh/3qupnkff5Am
sD6lqKsJEOThUefLlVwOB6P72iU6PF8JGvktUS4piAxhxxpw7GuT4setOZSA4n8apBP1ZNLOI4Mj
wyUY8xSpBlcQKbnnfx6XEpbcVJ9cmL2sS9WVuBSaOr/12jJikriCv1+k4btcXbbnSMBiP78sN0qB
tu7gdwu5XhsxoiwfwHY4C8GrAMfopytrN7Hk8w53FpeJZuAp2w5zr5rZqY+gALA1gwO7rTXIydek
iAOfKaOW7IKkldGb4+5dvDsj5wb8lbPGmGPL4arn+lFQMsO9dTyHX+WB+ZN145kvYECbtuE/EzJ7
PzMfz433iSSSrxwBzuNVgBsCzVztNY5QrypUfVCwVMFc0XcBUIr9H8zZQC6vJaYTg/uKRZG7oy9U
RhPpUBJ22SoG4ETziMH34mn1txKg9hLZq4IY5cFIKjLRpAy3dyupwAKwdLjNhI4SbQCjVarfzU1K
zqc/rBqv+3BuOK5XSxzjUrwiuU8WU2zYOup8N4rxCTKACMWUfCN9R2lIvDoR1q2OxTIkfILYCE9u
ATQWO0fbNzVE4lQvI7+CjMCZfdZIeoNnNJGKr5/GGzy/BdG/Smz53kPP7sXH42OoyO5ceO8zIB8w
9PiylYCzRI2/2eiwcX3xQnri3rMUx45URhTOZm/wQpjz20LkAZ8uHJGgJ1K+Qz3CrZ0QYPpYuAad
9hiCGEmKYzwM3Aw+k7nuWQWbv7gefPsY+tOZRZZqRvapKO3hs9TIJi+uxXWjWsuAVom3ez+VWalW
KFHHgThlXoogRt5QF73KqeAgXLyidD+76416Jxj2PvTgsjeGy3KGkxHcjMRN7QSeIbR9smH1c+Sz
xdq8ekHJqYwDVpceptUfNqkNF2+JEhUMJpnyLWvJfAYq/S0P2gZKJ2R0Uu6nz5yAB5dQlBTeEUfT
da7i2rqCYfLHa0dMSeBCbkrM0GReF8lcqU+321kgP1PsZk6eg5BuonxjGzGhm0zWEocq9Bn348O4
2ODrlc4T4pp5eNQ517+ydtyB/V9ElpCqYc9LMC2kYY/2GMOHJnd7etlIBhkNYQYPkzTTu1lsJNnb
B72seCo8WefYnP6l7pJqYlKsJRqaekXNotPKkJokVetCfshn2UuYk309jQJ9kAKMyJ0n4eaAUUMi
KhWTFN+SN8+qiHAqfThW3UyenAsO7NDrVxVtFG61axI9opx34BroNL+lCxC9oFAMdSFRBrBLjnNt
0kuog68D3l+QBHMyQ621DdwVwPwFWFj8o6fDTSIgVooUZyMn0eXSWxwjX9wCNzY0magbVRGd/uED
y1aUbY9MvJUYgSYV6aKLKFqlhmdeppZHep6JzIuu4wAVVsFeAev+LOyEGdP1yAtJtjAx2zcZTmAj
ZHpaqapT734emPKOKl930vEOWMNEhHOiP7jhwiCGuKHpY4RFvY+mlZi59p13VeIElXfhVQ5Bd7gr
I39QelKNBekRFeDHrRyzgGLnzLSfU3Nx3cN3LWlFvVFEsQLGE2baAxrAKshM2J5XN82RX9b9qtF3
MvW6eh8BcBD1R/PNgzSJD+d0wzPy7n1gKHIz1oXN7P6j33vd92EjvFGM2ivDM9JyTgN9qWJAkmRn
MZv1EPRURhQlrCPJhj9EfbDTqdFNeSS/Sox0BTjHvA4KZBCD0N5aduz+MaC/TufgaEfpVQ5lIBue
xZlNym1DCgzftAXe6Kk1URqvspET1F6FdDGPbS3Ozg8LOPFqE5JPt+MhF8rRJczardCJzJ9K8SxA
AmmuUFLnbqq55hBTR6JBBTKlOptjx73S8l5tesym8nYsaHuo9rRHE0dsEP22VHScz+U7eL0cxwVw
hEMjDH7PmH7uCXlED/6SJsz9Zpq81iJYpy38pFEvZjL+aG8rUV41KWjpcgn71xjbEzU2GIaSbTAC
C3aFkV89tHK1N2CVGhcvBRpb1xPA6XkjKQ6QX/K8ZSyNvtfpi2hbTjwO6R7IG9vWY1Z5awW39/S9
kg1VG+4B3b1/HbUgNZ7aKTsFr9y5qek6FsfArv0xNNe/KKaPRjZbkkeqD5lVCS3ST2vDdcgcIPgU
cBflxKaSguj3GRK2UpciK+Xa6phsfzOdKstY2gzklhVZi0dEa6wbhhJN+mMMtVruJH7LPHNMHp2j
k34vJld7WXlbQfANpv1AtUMrJq6NbhtBnOWPPFY1Q2ojKM+/yeE1Z3W6B35k8SD8W7AlKaYTbEDn
k7EYlFbNeB6GKGdlf7l1ig4CIREOnoYWQYPNwLLnRdQM6r1H9nRe9iT1KlcPvKQ2Sr1yYpiZLsM5
AZKPidUVwiKuxtB5/wh4pEbVjFpNkqxgqHR3A8KIiuox9Q9E6SVZ3oMZbTMya2b4dsxJGp7ji28W
jPqYF1+DoQBSqmL2w6r8BC9xV9nqBstGm1baapQpwjjChX/DUTfg1Z7dv7KKRv59jw04GMhhg8RF
1Mb65gA3SOB/U34JgkJJLo0FmI51nIPcGDtH2vpf2UkVbqsPkBN8dENzJhRoXXZ37n9QFWkW9auG
XAmmb409oamP9lf/5wSLEZDTzMBAtA8W8tiB7ADwIRvka6jeGaZ5/o/aM7imwxF8u8kaNNE3rCq/
+z3OdrxgUMMUSlYfkawSMakLg2+FGTXVIP4SP8a36E96R0oDW3skL8WSqhVnT9Sd2TuwkRNMUkDg
nt4CGtAm8JLGLVGA0GujxrOuTLiZWkcyOvw2vV3os11RhWRzwlCwPAMf+bkIP+Le5qov8bmAXYHT
1uxBwKNAznf4BhRaZS3r1vARmFRzO/AsssebBICCDBiEvdNA9sAI4rZgdqnUBRBa5lMJ7vb3ILP9
yGUq9RIB5FdCPb5xijWSIi2BmsCaDyNiypUjQCTnO9Kx6rDAypHSjN9CHacqy3wFJxTvymUF3Uid
5yi14WqcsirrWQ2LxDa/SMY19FCzobTUPUdH1C4ZXAy0AeWosneNiNv2cB9PfjbW3RIbocO9sf2B
3oet6RBewinOkY50qAoC3JMVxxS32UjslCEqVAf4LupkHmHUIH7/ENvP2Mf/sXcZKWWZ6mKNoOzL
gjlMq7OPqE7ZHb74Hh9ImGms1uyk9eBF3ZkRm/XCUXvJIeAOTws3YSQy6QQdeRCNCLbb9/Xp/Lmi
6gLApy9AElJRSPMdQEu+fU38nUdnKSfjPb6Xbgg2eAuZs7mvtAyQNRsR2YrMORhzfD8TnwIyiXer
bBLWKNae5rKyiigdTYZF57h3oWzMn4iJ3TDjJSON3IrNrRgYxRjnEVsgmXgvCUnwPn8J5pefdjQz
Rr4pgEMlq+0QdPGY4foF4i8JZaOrwK4TJwd07EosZ+Bd3V1ruQHKlbPz/d12GIT1uKOlkaWmfWM9
0prIoFF3emIj+IL4PbZmCGr4QyiJLCi3HVPXEbYMPP1njKcfPKHs2fXGoS3X1K/Ibc51wMhNLRWr
9cMWIibaV1n6kLRjwGrygzwaovynxtTSIsML0WqkAsqdT6dxQtB7Yso1id/MfVLIy5MIeQM0H4MM
bTlS2JWewvyeuIv+Htc0F5fErFapBIyrjo9atqzQmQJ4K8KlTsXlV3v3U6xsXJG+P6neRVl/X/jA
d1bbCI5FCARhGOPvgD+ogD785mQYKX6ecY8v9vBoiH41/ijaXLnXIx/nR6kfQuVN9gT/ttHJ++2f
tBxwk1u2GWCoiSvtjdTrhiXqRvDIxlESxQAdKnKNiF77dZYKS72rV7WHFIsYPTtTFzC8MJVGDVwU
eQSdPbymoKVLtaXHLlrePzAPLQyNa8laCKWDbfo6/vt++Aapo89G+kboSM32iUbO7An5DNezDYJV
FCHWJMhgYFmrLDqb6tB9Mf8bA7reqA66r+Nk28ABRiZ/7YEARsrmM6R10p2j8C+cHIqAjAZxoezC
aFOBeU6sN84UIoa7j+2IsA4dny0UeRH6F/2NuJySLspKQ07eCeShnZArTOQ9M22097edhxvCMy+5
oeH0kLhwFaLp7xY9jwAKU82fDE9ftvMBREqy/ngMA6q7NGBWzho5CFzr3M59B5wp6PdCHUurzj4e
BmgmZT1tc7WBu4JinQSnjawYbCc3kycxPur9RY7LRbGpaIW6l6/KMFy1GYkMb2pslQ8g6j1pK9zz
Z4opAoPKrOjK6gUiLWoVGa6SQl2yNbGGGn6u5+mB8m4TIySEtuq3FeCH08RdjU7EQSfK5yyUbirn
WjXVA+dp2iWqmhwGviH51L8QheSuC1VPGZwtuLVAacFSk4zLVJ6JGhRo58DxhsmFm3CjYAWkcMF1
WvoUu46DxUF5eedzsrbzcHtDO4vxVj//OB/shUscsxPSw/vV5TFDa6KIZi0rJJiRkvqoWJNg/bN7
FA/ZN8XcOzn2ysbMEuy/E62lqoniFQa73OWTJBHoFBa4RHXY3v1YmiDxjaYb5unaSKCPtW5FUMeW
gLseyi/pDs3yHsh7DNpWdNcJ5dAF5bByuAKz9ym9F3JHeHcFjAkixiIC5v0QYSvgeEnKQHjhMoBY
qVpr7oQCCdTBVq0iZPx79GB3mPZaLwvY+BiCSMYlQgmrAoJ+hIgf22OcYvuXvTdhKF64lcoMtl/Y
F//1oy+GSZSxm2SBNai3eJyABd2wIUtga0rXA+i4HymAgypeLRkCBqigWVJLpDnMttsfwOxtkRp8
C2/ixcCm/9vpypya8dTGOcSK81nizWnBBR/tLRBpOkd5L2XanpHDcV6YCJzsbK/wVd54wwHjywzt
IFCYgScDk7CpFIO87gpvHQRfY+WNZsYZwQQhYPT11qZiukTqpJfFY5uRCRQkASuuc6RxUKT9Sa1K
qPvSC1mZgQDoJ9C7MDp5Mcu85FsghK6xij7D6bHlln3gy2Rr8kwO2DI0svYiu+24ZyX6avvKLcjz
upnF+E4pXDoJPCvMnfBmmjgBEFU9ius8/3tEFJBr5HXVclA0VyKBMqhf0NpXArrR4rhbx26tK70/
93i/iAcvO14a/ZJuTkcGyJvJAXpQjvXcePyqQnuF0htTybu+NDzsICGGbpAMKx2EEp/hB3aQfF8X
f4Sk1iFqq6ZehOSXmSHBsbqdgTHaJKrGLFc3e4aiA31BYqQNiUA6VpFlQNVlcNkT9QapGP84jM61
4FoSM367TQqR+LG0YFePKD33KzQIIDMFSu5iByBQFDu9athjlXOsWDWh8/0AgZKm2OL6jUE1VO+8
M0wQ+jaD+AwP0JDeCUbq5Fl8nAhbYAIKQBBUlJL3r5JPaPaq7HavMbE4YBYPQgJXbBJf/h8k8Tnr
Uxgbxk4Vcy6F0TeIGPPDcfUGR34Pifp/NfjUvmtUTKDWkOV449k+QDqII0K8VGC/JDPugGU7KTPh
kQnyOasOqPuG31/lra1KPCo9FcwuWHfa8RWPvigIwCXZLNu8kHTREizBlWKtgWJtFCTXRgA527UU
RQxiGmR3uET4y52RrCRLXmLJBPWr3+NtpnhBGrwcIf0Y6AIr5JjnvuAvTVBVorON0hdOUysuhpj1
lQeoAwY/USTrg8zErOyJVu3P4WJZAP+VYBGgeF1Oh+lNISaPrJCaPofHC7G3vHDSC4183HxWiTSu
jqjBETSG7TPKdTsBcPW7F6ieYj1Ufd9DwI61RuMhNeAduh6TKFdr3n2S/bxhyPsvFoM3Z3Mdmab4
3Q67Ig8iCg3C0pKEoU7LYihTYzLu/Xf63LLu1QYLWvokXZfOlTOHz7cEQ6F8gxQihZ0bm7Rogadt
r2iOeASUCk9wDrbozzCbUE95RpApdRU6JD7ktFfM4Y+TtlwpYxofJAvjqSpPuSKCmOqtszxQEbWa
Qa3Gqmh5NaSuPzpyS+dQwEjpuxaO4KnUDvx9yi8Ce6LFQFrkirQXcaDzxWTyc7MeQ6EvBdv0IqpR
H3twf8ucl52ghJdnqeuMLcseZo93C54uCz9fhSY/FQ0g6meYYYneXo1guWTQSv5vEeqImFKORDzs
DEFGPMZtrEsNQhwCfIgrX9lPIZdkrCl9yWVPsdoswidfRGvZS+Se1AybeUiRreFVxZGrxa1lthnV
ii8kl6SsKmhCAOhohU0EaFzvCyTL8MFbPyogPVel5iz+7uWF15iGgwee2QqSbHUywQy7fe05zbpJ
G7D7p6VkApX5e6H4IF9fDYug8fqumBo2bkK2li+p8JOAe3tGDvShBeYGU7MMHovIq5bG0AH0muqB
tCMTgFQ3+wAruWj8U2PBnoyqt9HiknOLIx1HRne0PqlMLSv+Xpk6XqWnCAzE8E91u9ypR9axOF4O
2yVLRLFiPeDpfgyqbhwH2ebE8ujU5kV2TEIOxG1c3Xr1qkdtLxuM0suChZeRW/mslSLmQga6lTTY
n+160ZoK39spOFfUYwCojgP9OvOwbYSNd+iUcrOWRFlYVONh6m5md1WdGNxfZpy6LRa9P8RNvca1
TNwRrEZKYeROF8P2lJ9erzGz2byXaBKgUBOGU4gF43+7mYWNP0dGvcipLHn793x9gXdiAxrY8aTQ
YAhMY8gFCeFbS0t1sZ5q1DaExwISVf6iThBSjUdWIXYvMZYk+ZgFyYrNO1qkE1fOl9x5gNTRaTE1
eXUgZJdL2mr2N/zdVfVaIXN1FJ8KnBIX8/OVzP0vpSDRtZah9nAIvPUACAPvlI6t9yG74Kmfahqq
dPq1jXzwT41eYlcVVMqmlLkrtka2HPNTYgHGwww4p3Hnef2ZyMy6/XHC55wbAfJZuEYfzYAScPkP
v2hwwuD4VuFNSzEo6NbH4vu6AnZDkVkF4Z+3/Vi91umt8XqLR0IETZhg0XVXICdX+JEOrn5Dgxl8
pmq8NRM+ILAtgClxo9QVe/fmhIu/q68+NajPiu3njAAnMzUI0SwYNhFYaHmxgqdfyeM3Wj4/cjOM
qvQ5NxafDcABK+gMAIKwX2LrR1nAY808AgojBsScu5FdF5FiihqLdzb/XzUaylXO9H8hT+68ZzOw
l0JvLsNyaePyyNi8fXmGEIxmYIr8jxp2j/Bzk+mmvSd6sGhSOYG9SKDDkepCKWuKfoaQUd54GjN8
UY2j7fSo0ed0hgfqlHNgLHivZpq9W4s3/+bJkjVTDVLj62eXMpmUlZnPn3KlCdxKtwi8AVdz6IEK
YVj2BhU+roHZV5oQkkLoCMXpFSqnM4WED9gWpLgBxDtbXUEJYtll4eNiVhXy+mHLUWg5ga3ecDXg
jqiCuZmoOsQeRoqdOkX0aIjGsABb+7Vqfy8f9jMmvej1erW0TAL+LoQ++jyitlw0dvhbhdfaNvkl
CvWr87vtBgp9iikPSAfhR8J0WIlcImo9YHCzu9gZSYPK7bIyTsYV89xhpyDXM5FLNBbBuFzBJm5E
TCt+LEK/gtAnbne5MO7IaU4mDVq+sd74vbF7pfUOqd6wyZPFRcFBMmKkMkTHuzIRb3KU3POaNRc/
UL1RyigGybEGQPHRK01ksjPOx6zoLMPfKvgq1KGzPS9ypFrf2iMSVBgtaT1K6ckGtI89vz0YckGI
zG3lp7hJU5doIFzfJ67dVsCRJg62+D0XL3eoZl7LcBYeSqWdWTR0+EaF8xXyj+iMj89ddCWhCpg3
uDtEm4FEEmxWd1WS1MjsRvK8FYEmbpJJWdJSjZblHsftqLhHkn8Z2vfBodwhtC+mQd467o4ItowR
F/iPi7RvNILA8WrXWNR+GrYLDWbRHTjpLEgwg+POXeT/U9x17uSPcxO5Ev6JwM2sceUMvLS7bCvy
LI0hhIefDTf4qwdvxDiSldCpm8H5ZN+Auk4SMlDFY5bSPBnEMQu4tst8wd7geZIJP5NJ7wlIiFXa
+ULn4urCQKHx6Uvu4IpFIhrXCxJ1RV6nwCJv8p9VjkZScUDfzevdprcnudKx+0Z5ORF31CzjU5gs
dvcv9WJEGUEJWe4uJFQNar4DclFGCBLBv472FJFXPaIc9R9kgp1DG8stUIjk+WbUS0G95EV46WYr
OP2PFMXz6FfbR/0Fhe6OkHM8Jn1xzgQ9FHRgiAthLMGYsQfM2GOi7YNKMM2z48E0ujqzaY0codSj
M/HsMiPxMqdwqSSmzK4lgzRabA17XefSSsXsw0Y+Znsxt8BRBK/HMviK6SicAQ+y9BIj/EeHEdK7
UYN0eew8LsGJwDkAeEU3ey0oThi+9OGAfE1T5SZqSXK49f3zIALfan+lI0TajahmBdnpKepeOOO2
l7uC2vc8io0BdI849Lk57NfxgvHorty5+0DkmnQ0k1383wKLdRq9klQMgQaJG/KUAP1jAIS7Jgtx
FLVS7s1ZhJtvvkEr/aIdeFRd8TEvf8b42urnH7o6+iJx5JonWjFbeHGJjOXLnGDbEeu3B9BW1WGj
e1TTu3ZN50ylt205o5YWYlu2e7OICJHbb7uqc8K/Wnhp5L3BoAJpGglBIn0Pi98b5muZ6lD03FtH
bz8DZRwWBSsiCxnS/MQqYrQkt/RVEyXWSynnxpY5ntZu/RnR2zsBQKxe2k+JwHEfoCawrzB/bfS3
0bRbkS6j9dd8kVdaoq2uruz5HuUUkqFxhXofS1DXRxAamrs5oXiY53S0OYuC6MbL/AmB0Z5BeLxG
auBfkqRfGA4rsUYS7r0++eUfiaAZPwZQcMtu9u/ha+1EdwQNUHn+IkcNu/UPi1Ta/zsMmuiUHMYz
ON9COtaQw8j9XEV58D50v4T9tq1a1P0bKkAtbVizpOhthp0x+VEhFycY4CEkvJxTDlllmKBodUTv
LLiDGfS5NHjCqxB/5fb6mjycqPmLOBr+Q1PgWm0pfUt/dQ16RSz/cF0/XC8iQJX8avh7yJdQenpQ
8Qx4Z/C9ZYn6yBNSsmWhNkNQGxE90Tu+7EmuoSA0IHgWbSOAekjTOgAyUnyS4yTTyq4U16DZPZwg
y36YdY9asgL0XJ3mYE1R8UWl2m0qBRmWeFh0vOfIaw8SQRJCGbbW7XGY/p2h7KeGhRR4vwSGFsbt
u1jMTXcKso9G+iYfKyVctmmUygoN//fsmo35yW8ljK4DsQQlpEu4xNZUHAlhwXhl86pfNpPkbsSW
f5ETzphS2fZgmyWqFpfNb+jxw5VI54S+Zu0um6XTPq7MmPLlllGWtPjSQMbLFg+ViCN17I7ks+nm
1xrWHKJmgj5eWBVCMawY19cOCdrZRXYVmu8VpEvQVe954+rLZ0plUpvt9GEa1/eAvbMKb5UBdJgg
qRXJNw8sd+BMDszrGX7D4x6CwwJ2JODgG3RnQ07DMf9GtEJYNZtlSCE/i8azQ3z29tIqoFiGOhYE
qZxmuAuCJ0ByM8lkkNJfPCelptxGU5ByG3JH2H7UtFWMqbLsbD7zfQUsTf0/WsZeO85mtpao3CBR
uHzOFIXQkbaCK/8Xvysg/kocsShumLqw/0j4o1zUQfa/ZQZ77gYI8cVAKWjWynPZAf4PPoVk9Sr8
p9xhs7XkWhJnfeNIDAD0Gi5/3aY2gVGuCf9q7yhSyBWN2Q9mN7VA4o1qVc5XuKvbrQwwfhHOpSTT
8pMIfrCLb9xEry0Ozi9xI2u9ezLiVsX/sJRy4EBi0wpXM5XSBkEMWByhnEJ4KqQxh7nPkdqYUKlb
jGFxR2f7+EzwhHoF8qnRG1KMusPVknj03wapEOTVYoozYl2XFOwOVUa33aXyUZQA+FAnnSYB5V9p
TJJ3ubNZ7yr02yt/Ug4eyTZ9HuS7N2EuyjbYStU/DidB1uPSCeo8amAGbcjk7vwFmg4lGrtk7311
isTwT51oWuXdnRo8x7bvs9UHpNtVVsvTCuPGWmHcOZJjNMRApGg00tccUE2Y6RU2u2CgOLzH1qZj
9r38k3uD4tWPPM6G4z2lKS5R8O7nEx/QWqTGjDvS/oqdEJOkv4CsSIJfA5hsSDiCAQ8z9TUVo+W+
LIsqrNbqI/Gi+a7qE7CfHf+1fxYVzX9Fv5cRufh374WI6bN5fyvKSSY5OdCf3UJJaqakK5lOQmxn
csh1jl945sJ5jrIIfPdp2U8aUQbe5HKdLBf1Q5VXQAAE0uOObnv7FMaOJVr95+iQp0vDJ3Dj3f0b
XdikGNZyAfKqjNCUKpkKqTG/0AcxlwC33GlE8T//pcfcl2ovv15rbXi1kEgfit+rpV7ZCvKZjQ5H
iLwbAqNwHLxftYOAx0pDAePNXv2hmNpYZZnDqesoYHv3GPxi0qMTEra30wXU7ohiD1wU+kmNTu+3
JPKVqE4VGHIn1vEVY6E6iOwuL72GahmzmVMgQ1aQHkUB+VEfnPTcAjrCh9K/OHaX8vKIYolmghaH
PP1A+N+GsK8KsIKGtHt28Zu5/aLyLd2W8WLIxe9yLzXSU0omuV1FF2fMqChaL6E5lnnn767g2Bpe
ZWhPyir22TO/BPtHQFkMZTOm1pADfc29RY7sOh+y6coQRgSG/IWWNZ8u7NOquOoj4QCAYizESSbq
BVByev4QKDu4u9R4cghaoMNN44foS+ReEZkS44fHXTvevqx4sVxF/lmWfp4GLXGCIaaGru5sN+CM
jPgADqikv28NA0hymxMeXtXSxpr+IL+5ozkllSo6yThj6+jBXih1dwUKp6WWLPgTygt2Iqz2q6I8
17PSI9BKDv/RUHZLPrPdZ4ZPgyk5qa0nlDM4DtL3k+xNq+HXUlwkhCQE3yGLQQP9vN/gmI5gRz8H
weYfPzS6yxUU2R3EtDdzhaiQzxTcK1eOsOHw9UTZjqlLJLzAWjt4J+NiVfZNn1fctSa1tCH303+r
YVmZndUb+/r6iuwxMGtiNxxbdUYk712NpZfq/QGRvFwJWJ0nbTs/jGwdX3eAbozuXA6+JUCRiF1A
BDu41nriYG7mswT6szOnEmneJ+GPBmrakgpWCL/qKU/C6ilPGiirlGez9AJmxZeJmzhoYNsNlLko
7skW+vgVCv5GTKYLIAdMUONLl0F18Yfl/3mCu5VQDRUqYEjtXh97VKtCTHg4BgEd84nKgSH2EWQS
8T/lFW27yNV2JK6E9yFf8nP13SqFqTtSSfio/8nDD3t7L6q0Gz9d/L7+Nn7w4uVXUHVnt93zNtsX
lLN43/TW2JsF5NI2mbTdg/Z/Tz5S7KpTC8dhLfDequ2/f16zWE47KIMNK55DepfjTPm9SxD6OgAd
QzdQsLYBlzxDLJjKh5bvfJv+e9UYPq3tTLJrUIp8VzrxKWzTBb5UAIgUbA+Bu5IekCVwXTcBGT+p
l3nM4gF4gSlENYMA8sblX/ShXSCtHnKGIfXpWKQDdSzdoDxhwuoATT00kEwZcLRbga1ylJlZUol8
dIdArQnOhCbAxgGOHemY7U/w/lX1LawqmGt9phS7ErtH+hlLcdAhJzAX0q+aXr2psDVkh6LU3GhQ
gjKKS5/Y33LzY1Io0iVxdzg8Jro0n6oCrNt+mX5Na1lVctF/xd2hoNaM2n2OqH6Ed52K2XjlrVqV
TIz0hHZfjabk6WUIR/dhV8jEi6vAzhw1UBVz8QZ9uyhzasRTOrJ9NPdVH1xLr/Y5FZYeE9TINmU/
JRzkcf84qaaqT+dpcSkeB4cwHNd763o3gr9L4ubTTvukTpqjp+ya41MQuIK9aAORglVbG3Z1rg8t
1ZobtukETKNiTrft73mmtS9Mue8D0QsLm1JcvnSDnBUN82oHByFYH5J8HPgQpI0QdFx3GCaF2kxE
CiV2vx48C2G5bYgIKKPOffniTTqazR4R+Og7OS/mW7gJ15/3hvl7fu1/gpWjr+Gm3z+qgrdbPMLj
85Rwd//VdPu+LaujAzSKTd9kE7XBOSgDAdgIeic7d+dl/YlhGSUMMrGXiBeg6U0vwcsYuEfbK5lC
qFpsUjqyjCsDlI2QbiKpDFYGbTL9uhUNQU5YkSEEbermySaI6rApaLK5Xhc2cwu8U65R85UbQTrH
LAl80ZRcqJeqrCXIqNGWztmQnCFy8Q68EVvLNLTVJEFNJgOMEIv3An+GalQQiDCGNAfxGCvzjqgv
GdKnBvAJF5fqr89JFM691QBwF3LP6t4CjNS8c3KBgID3VYKCBNI6fxeFgYzIER2yE/A8VqLfvQob
zrpkSMhXxsZ5f717xBwF9ZgzcE9JB4HYCashRgzAqptK2qu/dqTA13NHq/KAYbv+Zq5p07iSJBiw
fvA2HcemCjCZtoufR6Cm+oM/wIAvGB/7vtWX9XzG+JP9B+EL7XITjJE8NEoCPxJRw2bEuNuQKB7j
cw19PnOTVey9MEK3bU+Zfe+i1MgYcRXApD/+RcJZiynJvZvGK5BVdg+8hNZA7tbj2RPND2N1oVvU
eMDzNByT036KlkpdfQxsERCUun6q7kig7UQjENIfk4AB4GXpXq81r8h2SIWLenthPLlvWxjcRA15
/voYH9yQqZW8ASUUxhEhqZuEsCKLl0y53wVEG9tGb8dicbSJyQtJBCjE5GL3cf734B4vJd31g6/T
zL0Hh621FoJIJf3kvmJgF/zJFDJ6FHjTXmGMvYB1OtkyMC9ZBOEvA/AkONWolFvCV7Ng2T1LL7bd
vCxGE4pPXNyoqwub+eT8JuYop9K6e9QHvLwKNCNxr5iLnuns9DGdcJm/bpt/fjsOoI8ZNCrA0sMv
mcCyrbfcpm/MjbG60nljEuV5/jXWrcWlLN4Fs6IY2gUssxdBR1TgJMUR02L+964Y8apNHCKMASy7
BkQuhA6uzoJITt5HFsh5t9W8cgR1DOCCR+DK625OQMYqL6bKfWfB1sX61RiVYtJ3nnF5FllSb3iE
jNeWvw0vp3wBb2Vxj2kx4jeTmVzkNgvdYZmfFyh9+7NrI1LVlBEC/kljp0HERnSVJ+3NUQaYqr4t
Suj1x+8VZqMQC7qAhe/LhxMmCa0qscdsRhKy72/3hIM8i3iDy/IrOeVPbWKzf5lAxY6Qnj/z2yfA
OWTMa4CJWPpa713QyWdPkXI69+R6gVfB67ZI/6iegzDlrdfJKgi6UDKBpHR7vW7OJc3Tt3CFgPE6
rK8EiA3N0TVoqHgOKfVblvGbn5nsCab0y8asecmyOC1sadYC0b0wsidaSt5o0JO60tZKX/9nGYZf
cvi8RdmSKJ5HK2qH4OORelt51PwdTnhVBFnqXWTSFy0La9r+1Jh9LpvOKC2iQEmuw2UXI+uZytpI
lLQ0oY/TCgWuVQQB1HcA4Ca5IXF15x0QZTVIjSrWDNpNs627SmSTripOwiagAcO/yQI2PQ+308+t
u46tkQhUb1vihJDoni6qwl8+FVb9PO51cKIERwsvLaBxOYwuJKNOnAJhhhh6ItLhHsg47yWYoZBL
k6cUPqGrWs6+kOQX9ZHiq4zqJhZfd6CVCPj+hOFzr6d6PEWJy5XsCGupbHbu3iDwbL9gJnS5KxNu
7+br4i244cbXsa9/VgnHTBRd2ImeoGH0m0pd5tYu487hBAPYKFGd0Md9+KsyxWkQewqcoOMA+P1p
Cy/QrAcbbQNyNVpiGPrA2YOhVNUgA9AQjW1jBeFfygm9rILTFACSFWpWR7HLrwOc3KVcQWQ8X+Mh
OY+T7gd2O7eHWuJj8YQFCPuK0zmon4a7+rRo2sAJpU45VQE5fTRkh1VvTmynkVjEj/yR3lWXRbYl
j9cCzo0pIeosRp//hPMvlSQnRJDGOxUs10AdyhsrmKIOcagXrmHM02B0+Lo02uX4LyYp7dL2K8fv
feqcvCFJ/HQ32/TW4/hJwIbIw/5rRzajO52NrM/ZH8EtRzqtMQuLbMI084+SRTVqkqHrWdCiMpBc
HuF/SEt52IcwNE/SdIn6cz0PRvekBp6WgD93ohhtnEk3dmnoMGmYV7Bb0VjJiJK849F8A2EDrWAz
OzI/qMXCWi5pRElTB86/+zo+UVTDGjIGT07imC82vPeRb/nnjgnqeeoPYhuMc2wJmlGiTwQyfXrx
isiyxIo9im/y7NF4F+I/pBtXp55Inhq7j6QNRsySdy3IE+FSGZosF+Diuoy8tEI/l5oKuaT6HC32
UiiWgDwZsOM/I5Ptwzk+GoV2fIsAaR7Dmw42hDAMngfFOYZYzAJcvH1WYwDv45B8p/kGkEiZrU42
ZPKmQsOxX2JXPUSwJJROx57RGmwc8sLhuRlQUpUclnfASi9ipEEyX9grj+iw7KuHKTvlkCn1IICD
Usd4DkXKmj4EsDzQs5gXlBxnPCjQsy2nv5xNSdUh5yLIbCZUEyDbbcfVn84LmOe4xoAHy8w42kxe
35XXu8aqx5aX3UNIhu6BcmOMZKyer07VZq274CSJ0Ij6bLZ7a10Pm52AuC9KooVEpgRSTenhTIQv
QDY94KlfV4xtD24e7NymGnmGa8HSeQzOaCuepd4i6wmdTdUyiEc0GZhGonKep58JgsqRfzGlc3ct
LCl5DttrwLpuLs3Dh+sqosWtxPtbtkXqqlSr51M3dBMR9XpNdwlk/vE04JGYMcyxCE6ggZEC4NDn
VHK26emmsxxeoLuPc1eq3zNDSEEwd9ppS4GCT6agzBhvjfVgJMXyFAEQFna2R5cVifvR7rqlHLov
4S+hyW0qWSDA4f5UWr97uIGxGqIvvIJobg8ItWUAqSKYto/WhAudXDJKqX4kA2b16RcUtwLj3iM0
8AjvmsZtid67F7TdtmRqX1+0Lc7YuFQmoVbaEQ+KOaHKFQUDmHeWnTj3ImeX/os4cO1KyLmndcrB
xJ+naT5z+gRk1Suu/kPwolrsmkZJKtVvo9Ynn35RVxf+y8JobkJocECwMWgvO1TCmKnPWxMjNjwp
LAs1pi+m8PD7EnFmdzGvO0o+jn5F7bskF/pqXH+dOqGRIrq8CYouVDaJxkAbxDiOAzrthwnQY9TH
7781ernc0FZrSZGoWvllMxIWhvwUnQZlVnWvXE8rlzLY8DU3GF0JCsNhvUyXsoMRgCNwQPrv9w3v
UwuF7CvqzP8d+ro4YYnoHdE/HfsVFtCsO8SQ4t8rVPijq9ss9xXXVqXbQF/T2E9vpHHA2Q8TEKg0
zhCY/7xCj6kY3+Potpy95Zf1Nzv0vUUZT+ewkkT85rcwfKIc22I8JFMhd9/lbcRviHF4K94sG7Fp
B8WOUiA9BpCrzxKmikGODGBrA6F9dBKV6pFawUUFeCI7rw1ZCbVbSlOcKmbqeeuSsAL4jNPevXQw
la9w305EcGKS3gpJo/m/1P8RZ7ic4vTy925RFyLjhBGtKVFiHSifplbfNyMWP4x+Azhdcmx/VPnZ
23sEIL8M+LBhxPpJBwXxdsiUbGgnJvE2GvW4eNvYIqMKdzNP3YZpwdxqUYZyN4saj8LpBBlyvS6H
lVLblDiHM0zitKfJpLe2tcM4xujOxw9O7VanrUOHYTumGVf8ZsbGyToraeV3iR55DKem9eo26Gb2
MiR01m5AxCPaHDiwe9vUNRYmIZg1vL0jlRopyKRlAYvBFpYqCRyDFh76h1HvYgzbOPdEemyIr0rj
IqreYJRW9i+3BVATJ+gonMjQMkSGgUNi77Go1NeQIfOgmvnrYV0QILB3dZilWiDQATozcJlQENfi
+QnIUUVCQjJBAFT1UCIWQryf9BetLe+TgKygsbvx3x9IIDoPHDMPuZJMnsh2EgpJFuOjHqAGWX0k
YK8aCJTHeRxAjb0vw0ZMiHkDmvXC929/IuvQCWg3Fcbo0vfNe6p4ivwTAqT0i1epmRZN5Ne0LRkv
I8nqQhRLGcHggTvzUjCxQkYkQAXrgrG3bQQnQzViWWGSDMXvz5IjyvuEfF6XINUGmySfTtykwV9a
yZEWEquxmhKr61+0DRbr8Pry8wf/SwH2OTecL7KnTGYhafS8NpWX2LuiWnEECHuaeek6nD+uooR9
fgWcpTbtr52OOiOfuSSo4Iw1JXI6dE0lWFdKW4VFFOcV1R6Mj0rV8Drwx4VIyNvQ+sqY8GGCOGcZ
I+2pna4ta6eh+J4QCuu6nNAR2Lq+LaoJLcGLZS9AJ5qkCsPXM03YMWCZiMzCnYMjnOktuiBkJGlH
tNEoXGX0m7N3rD+48T/oa869IbhKHMNXrO1RRi3imEzheHF5lTEhKXg3pNsySR99LBOuTN50vKBf
pyDLDgQxfEsntaQcfGlV5BCrc+AJ44D7Oni8TxVabQGpEkFbx3by6XAJALOjKx/eOrDHZnMBwdsC
lztmVwWUL2g5RTg4kcPi13SOgjdjgEUBZ1c6toBSIjJlrMON34UnL+3oIbsFcEGV3/mZUS+1h3CQ
Yj4bw3Kz4vKhhcNFqGTwIeRl07W2eiYjh0GMiOlOEwHJ8bwUmWBHIWuNL5Ftxf0Pab2AIOtWOoD5
hL9EgrOKKGWpur0V8mwq6EwtZDHdNnc0zozZ0SyYYi/lClg+NrblaOKnAkyw1IdDGMUHxeV6EVdu
J0k1ukylJvafYjich+suJAzYwC9EF+O1pqGgWsmzMfCJdu295FvTsdw2YQxzCM8kq0BDKYu6mB1k
y2r+rB7PgWbr4YF82Reh38JtkF6AWxoeTYwZO9QIcK8UfC4zd2LCHRc74N8UkCV3nGcj8vYb+OQ7
2bI/W+Sjli1rcMkftc2XXmMDr0MnB3DXQFgA+Gm7UQIRgex1X/9liS9CaOy0a2KsV1yAGdkMuYg7
ve60XGyty6ueyGg3qh/kUiyGS635yPGk1+poIskjeZDzho8HI5TccVLg8+gf7fwnAmY6MW1HmWAl
pue90raNev4ehdn/e6lpFeK+7w8UsIXRZTiijcALcT8T28LFYaY3Xl5aN9ZwRku5DHuLLHmerUmZ
s7Gox3jAxJpdd2u79wpa1Q0aAoc+usR8ZvWtvB6jv7KGyM4ERbTTc9OhOfZezHNGZdYeZst3+Y+J
zB+Oy5R1RWQaliRv4n7XX/NvkjxPRgA/9F96df+CbnFW6UjUF1SaKHOSQrJ6dqoHkea4EnSnlD/M
7ZC4LLyoyRRcM8eh0MdJtmizGBCFultgJMGhfWDz4/WVHyEIU33gzHMB6MNvMkX2m/fgCUPCmo7w
AXTZZ1VCGcA+jRC/Xoj7NdVRDemMHSw4f/9k41tZx5Y0DfFuG+HWQdi58hVQVJ4GjjJHofUqMGJA
RYO4ttzEY74vIESzYcJaqYG0BXmiaqbn4SeY1Fto2ypQTMM4cxKiXnv68d/jI+ddybS00RXIyWQc
RN7rQ8ib340er3KiZt4DKHcMYmlu96k7L0iqwwDuHX5o3PqAvbJT5r/c3BdCDdOywpVKcqba8ZB+
9wWpiCrcm+ulx/njKm1qVeSgTXdizbaOPmSVhz/kqm+E/zpV+4OQSCsYUMeBJdVm3kwjnDXpwtRI
fxQKTxRFN3z1a5E5CfHoa128UvsO+HdTlPmeI3u0cjSRJTGMI4z42jZljcGxZyqH9vaCwAw7ukGF
QwayShxYTAoIEcZIwBf5N3ys+tjm/EYg+PgHoPQir5QPcti45l6a0sf9/JkpIEQq082ConHwe6KC
HCEfz4S0FfpDycG44+5LMbqELDh3bNw8OwDLGyaF2tIc0jdi3jRHNpmsZwpKC6W596kkBmBTlFHq
UG5RFEIUftwlnRh2cQn+iqgZ62Ir+LxkRayPi1yPvzIX1+Pv4x3ef9uY28icMZgDh7BZPhV4QOyn
n1kvbkK2qLAu03bejYLGcsP69N9Mno+ZfDYxQQPNJoIYy06F/a/bUch0PpeY+0H1+QnT7MiPPFsY
0TduFc0+yKnv47TIcPw+DeTA+C1DMoapPmiKTDMRM2TdCha10pnKpcaYLrpXas9coZQNBF6ggygE
kfpYJN+ehwrejw4sPvDIPYIOdReu4/oJ4TvazK43qeu58mKrBG48g3yrjCk377yuB5CR11VtgO5m
tkqyHiS6P57805SERQwKrJsfzN2HFjH+oCdLzBsyWXl7Y8dVVPS9nIBEG4go9F1XG3TLGaHun91e
EO7MbiKeKf1CaOAzoeGLgvEoAYvDVHPm/1z2LvHMlKdlWxvEnZsPi0d9Vv+4OcEsXAEl5kcTsZ9K
jiMtEHk9trtsj35b3QJ89+965MlE7WySR16HnR1OPwkINaijPYlpjkOU3x+iRisvy5pE3L1s07s6
QZF5ufA4m0+dpTzv7raZiwHVBvrYX8Z7NIQBrtufM8/M03BRzsTgaXudakk4Ig8h1Yss7QJDpv2/
4oXI98HDCVs0EdmnnkRcp0AQFn9SW/LSz3C8C+dCHuiHrDGJ4aGlu19sof4TpU+/4oqQlYJXEOyp
Kv525cB0ymk5njg7lcQ0W1CjQplKP6Gqpp4ZrMpfjnMT0QEFpwblrb30ljHnoU2teaG+4QbYE5J9
gdh3r9vyJ0ETwoBrBR7treQl+fSPGnTsOM7JjjrgKUr+yWQtuVVuz3w04pmzYMHmkRzkJwkLAXKX
gTUmbze1Vy0JV11q96PRcb+pfzhc9D9eZUj7sRdcuyMUTQU7ovrjNDjZqW3WWDH7e+MeeHhetVsK
hl5cVwPLNUAyc8yDN4gv8gMYnGpNGdd9gEe/OggKw4zpu5ehMTx9p/myHxGTc1kYWZPnU3Zqbfxk
cGFQY8kO4owPl4LwOd8mcOWoxWvaRJa0gbEndeHgBxwyTINf2aghzvRT6akVqpsygnco+0LmtkQG
l8YNEAQtArAj5lFbB4fkdSLtB6bLMcC87L8Lk2u+gQOGxeeAq1vLHSbk17wxOO8O3zBrSE3b42ts
PnyqqRaFcl4nmZBHPNCZ+2ahg3GbPjfsI1jjodG9UjwtzA1fYxm832AHN+iakA1s9q1nxDwK/NC8
9ruxvt5q222M8mRSxFqjCLemjEDCqOS1p6mt5aUd9wKx9MJVANRIFiaAm2P1R5IvYEaMbfpgsbZb
EHCFbCJjkFFtJjZIzVh2YIThWB8xDVNYd8rHRdYde6WalYKpRHzQ6rPlbZzUgZv98ERcEeijVEyF
4H0eMLSZYW6nzLLdYnBWIQZp9hjA/mkV8R+deyFcSDTk0DCp8j8e0cZ9VW7LN9CmtgiUPcKFtlly
868a/uF0kg6VVbrpUxPAIdwLXlJiGUs4wN4CWg5oa82is073zxvB4WsxFk1d2n5k3WOof5UuEDaL
PQ/uW6bFfdKeQ3hfwTOOumDMoHQosoHmLk7GJnZL80tNbYhV6SCEpzL8wxH/1lohea+0s8JoY9kN
PecfM9GlUsmc5Vbk9xtGWVSB4CoKKxAePZZgPq7AAlHqFTmS5bfHP696tqMbhFksPH9AFqFxA/02
NYR4y7xbZ6FzzsbxvQ5N+zGibm0Pl+f6XCB4xTKGj9M+nBhwY4ed6uAf1UW/0+CM6/QiZz2CVpl2
a/icdsiinmQeoiD/lTqnYcXzQzlXf7qakZpe3fOzjK7bRLtVyk/1PmWg5/hiyATHiLIvBArifn5Q
AjC5qgYWxMD+/KRZ9GZ7MIiBOMv1FEf/Ipi8ymV7viywNAklAuu6UwZBCGMAdACVbjtdHAiLZSYj
BXCMWZqToOZj2LMTNxY/dYi+zwXibuqwvRcYX3ttvaBC5b0WM6+l1zpWHQkDARwLgUgfZqLLdfYJ
QLyi8gnZ8BBKgHIlOHPGlqaWdRrHneddJDQi1isomzXrinEo0TGIlF4a8l+AaZAoAjnXn9R96+Vs
01/HrsEuRCm6IJhrXkDjG0SlwtB/AdzpKBgyfareOBgqLge/BTgCm4j3/bTVNnsuizlqZgEHV8X4
uYAD1th7n5MCkOESICu4XIRDRGHGm+JmSYmvKAE5J0X02ETqcLTLXfk6VhEwFYF04SpInmaKeQ7u
coYX0A0+oXjzPr/dbR2hDFK3GYj5W8FTKQ8mSB8xQ04Ld5cxYLxssyp1cYXHMQihRjeuVZR1b+eg
qghXDH5mazKkKEYvgFZhYjlaYD8Y+NthQVi6+UjImooFaV+DbVdZ6D56r9xX8h6tGYwGovM42cK5
JWLNwaa43unMH8LEooMT4qy1s1FDr7O//wcvE+FjlGGyEMtN9wFr5c3XZbfuczfilpUInrKVVdby
g+1WLFfxgDeGRd2iyBroP53Czi2qVLo0cy6l44DkJ5/Efmf3VV5kN/PQj691lPGqz1jYxRcm+Qst
DrToTHLfstpPTCqzVmNmLjQKrXTquNwSBIfL0+ebxqps4NWee2b0UXONLJ3H1pOZrjRY4pSPEljx
zToFtxoRKBU9F172mWU9TjtMHbm7Ax2r5XMrueF1pn1Cic4V0mdmu01dAVLBTTOksGodsR8FraZW
rBN0M80aJiys99Ogum7zuzfatRUVfOqJhYqcLF/qPs9WeT8xo36emOcUiJqgvMh4hNT8Uj7YoK3q
HE/xo+7eA/hPA1HxUAKkRoPR2DgK51o6bMkRNY8sS6G0KeV2Og+MTNx75m0zdJcTM2SRClTh0ivR
GqMXIK7uICujwGebCHlCQpBiU8sh0/jwSW5UQQORfoJaCCEHDI4Q8lpBtGZIifRmRuKG0tXRl8rq
C3Ktg/RyjUpec6bLrq/nn/3oWClWCUWYmXWFSZ+aNeoIDDLxp51NULu2futtNCis8fxKrpjSGXH4
dnKNxCIsqGllmHgzx3/WBe85zeP04vek8uwKHf1ad4BLrLlW8BcneRQ1a1E4CuKzi8mJVF6glLsX
jBXBHaLDJXusDxc2R8kiL4K+jlFcRelmaUnTBp4Zj0tTJbT56Xv2j5/tQi0+5NHEI3GNFncMdVo4
Gi3a76eIfj8JO+EOt/KUogVguOx+Y4BJK7Q9w4dUVEwzc0Dqr5WcVzAo0EVy+clknyoiY0lecIg9
Wt6Y+madblCzgWQhyxOlDHBKdFBqc0V1UI17+a2Ux4cR+i1yM6++HWTTvlVIjE3gopai6NvPuGqz
WZiYTeQf2mPud7UTyN//pnpdxkGs6Tt8i0l8BHU4rdVCtD7ihx9N0tnz/WrnPgaAsaDZcnjvJFyy
QQmEFXuVrPCluPpEEl7/zTAIU2K5ByMh8TUv714hRdQuBjpJPFgT/vM+3xK58HOjz/759GH9wBSd
DYr5zJpxi97rpqVIXcd0rD8P+IeSGTGDNO65TGyxCr6fgm5lPgciCDZYtMZTuuqbmhpR4vycMCOg
nIhXP/gk/pt2Qbj6EBmCZPqbd3xvn+1FKGjKeCCMlNzPO1e9UFF/QE068X/9MYrPaJ4bRpeSEiBb
2yv4qzCKndHJFMB8TwXjNL684gS2AKwgPaTraGYlzwvUP7eHR50BvpmnfSiIsxG3LMfCRkuDZpjJ
kKzy9+nWB6KbHknGJFB5EltCu5VCOL+MPKySNaU1jI5sH3l4iFdVNCmigvk3Y2Yj8bo8+R7mrRZv
sqxyzFzoLlZNs388pZgMu4J0h7ggijvbtPGnq5/IkpC77EQ7DkO4wuCKyAIBzx/WivzeOQiSbH80
o06jdD2/jAo+hRmsG5groy8f0YWHzWzKhsMnwYrnsLJdqygwPNbrW8U+Z2Ug7cRW2AGkIIaoXd/6
zl6/cCRuffdBpfTw1JZKjdfhxZdMA2Cnpw5iYaxG8Qltl889a7Bf5nVTWvhXXTgaJ4nIHLZgPxD4
61rfTEiZQIasOfLohbhBuH+ep/X5MdcfztjHxMdq4tIVLsDmlWkJB6lpaA8LNOn8KFHufEXy6neL
Kzu63R0koxxR0BUAYMWyus7FTYrRWZ4RNjcIEBuPtfvropAbpPJt95+4UsjcYNTO9V2nExXhuLSB
H/O1BSQwEEPb9xkP/mCDmy/vf01jkuDd0k72LAav+cDjTtpaLyp/Ob4+KvFZQvMzwR7zoJzq0AFe
7q9ca+5iVZIUaDWzhU1WaOsCMXEhRFrNIrFseJdWQ0KdfI8OkMpolgKReZlCjoJNuxBTmlVJH7qw
qy7bI1TLLG3Ht0Nd9IVJ36b1e9WDZTfPgP0hMttQ8XXy1cttLJtmwvmZmtwXMKZsT5bF/uMQfan9
tk5y4zGSzNLhOm4csxIqLyRaFz+WupO0E8rbCSoLFWTMVDOAvYV3U977WTFh78dtH7C0DOMLD10B
jdY2gs6oK6rQ4hhimY4JC1PiB/+8x+huEM12HY9zz3Xt+BaNpgzRbju4IsuF0aLgLv24qw5QbMuy
tiIxvJA8R57NbUJO1nH8rgoagYg4kqHs73wfe2nnT/GZoetSihZuWzWB2PLdfmRujHHV+PnEmiOM
MhRw/CH0UgzCPw/m/A694pxCzDmwp0w9QDovDkGxFJLRzJ4Ve5UDIO9fdUhmsgivZ/c8v0ja7zrj
A0s7xp2gNPYwQAoMI0QxdhGQa5fYlG5zqPfFWLGOLXwlA++oAktK1y1qh17369oDUyacGoeOzeUt
xvPsF4hLkDYvFY2rjKHESpLEiAdS983Hkb8MheYVUxkfDiUTPAU0BkfAkQrkr//jiCdgzsYS75G6
sqE/Yh0+4aBUbF8FMqhKolWfrKb3C/WBgd6wLa7uplR9Z5plMd6cD4LcLCrBmRKr0VFmyVikyq10
Bzav8i0jKPvRnDW/md346Dn27psaIsiVrpsYYf2y0jCeRFZW355wl3bpgt/Z3S9MVJnDqXd4nEXP
Ru8p2pcrjOkHlw+iAk/g5u/adX4Mkg9jkCfaOqi7lqsAbRyKKSrjtTPPmWE3MY2DirdHSAF/R8+G
VgVTYTu3Y+mk7hXj06kLgxummKmPD0mdWBwAt0Xnb7qFI23C2Azk8dAsOJZmTEb1O+QNCj1Tiv6b
oZB3R/SCj8BHrGliBeOAsJ68rJwA+ATImF8rswVcU6o4SG3lnOJgeqrTrt/qmR0YUTey/Ltm4Ea9
vA3ZMaHAJ0JVG8zPa8yVJxfz9TYZ7dKxTTqMDukREZ3cIwSdwG8nOfc55DO8oDcJO11vWCc4KT3P
tR6UY09Qnm3MYQeIRGUWu9Ehjrm0Vzwh3wwcW7YPZ0k12zcmLPCrOF42mZJI6oPvBCGtyJFXAo59
Pf9+9DrKCyxZt7mGU/VG9orNHETLrlmaRwxNMkYdDX4GxrG0pmfn6UzmHGDLCqku44XBLDkO4B74
jlVf1yAhVVgyAdZfzaqFO4Oa9d1d9WFC02wI9BWWK/rTkIERXDCDlB/koDKQMRoGXvx03iiyP5cc
zpC0LnvV5WI15b2X7j9vZLvBi43ecleW+XwOP8DUozNYwgTb2A1Gdt/2iy8APytW6T2MEn2lQ33K
TDBsGczXTB99ITsnYcmm0PLJMNlj3xAGkohxNmzY42yAFTKr0251NAtBawrQ+FfeiPexk1a8tcSo
UHD/67ix7a9PnQtPRD5BTlKxPRofCYXGYZpXsiH7reBM6xTMkXDOdy3482R4DPxPbL+9Z7LtpxgG
avf52wqPeLRXzJ/ZYYrFmlShtMq1gHOwThdq8BKql+rIB2W1bzpNG+KIdZZkFJExb6Io47sKJKGQ
WI9AnQNaO2SkR/kC7MR/WW1fNs4I9L3jhP7/TLAO+8ZBoypAyk067Hvx9012boQNtJ4+RtESLws/
eq4MPT/LOYKLoEY1xrSzBguIlsbUIYRvIeY4QYMAl0dKUkos1KLR/Ytqzxqua8YjAvJvhXTdnkz1
1JRMWVnyUgWlEFP5wAst7yndPiQ0jWVhrK8PwfBTzLT0TCzv4xUhvBi1Z/+9EePVTr2slJECoY0P
McIihTOR0cHEq9qrB7lL+DAOiIJp1OxGxw0FOb8ef1swdjpLpZ6T4tsQWUE2QUF1vy1roRC2VyoH
y13mEqd6kYprYasZeITGyTlm3Da9lp34SNhHeOOdFMwHFQXdshMrs739NNLUbcXmGIfDzpZADXoj
QKNNsOpnTAO07Hbuzpx+c6WlRAqPuIKykm/ta56Z3PyqUMSD40yBqPSqOEImOemHgw8aidfnqc/Y
hbfwqacHqwCcpOBQlMCgucJ0FRYB29GB9Goe4JJcpzKFfn1ULdhUcuSTkX3TKisz6oO8keQ0DN9X
Sr50/gq5UAzKL6KMrnGacIMLDhiFzQgqCxKC75S9nOyPoGWd8DOBmViowyM6rA5ZzCNEg0l1jNd1
dubrp39liJU8bWZ0C6y2yINNs/eIemhxdIi+SSp6Q6KsPPcCzbRGngQYQQ073BCKQcxp8o6HLSF0
dJwEG9FlpztT35/E8MPbT/oBdCq3CX8YmbFiSXWsYfcYYHDpimqlwwmKJj3L778T8E5A4sOtgpLk
u3xK9DUl8GtO93VvR4nWnV1tfc4fTqXBZ+tYjyDVq9oIh1wczWkC5sH2xmEhNVU7BQZSveYdsIju
/85FVqkWbakrlbNKcbhLCViXbLzNSOTC1dfLDVnL1xEC6h7AuowajHVXm3BiqlInr0e1as2bYWAl
0K8EHJj+FsJRJ2FwNG7gWYlOdg4/81jfI1XNBoZZPXDCAYrL3kYBWnc8VV1/Ye/GEQyC4cdZNmp9
acIMv3xLAmbjnlTzKJKZxy70LNG0vJjdtfou7IZwL7/kLGtgGoQApNxTGdJTKity2R4QoI4NCC9N
ul4yxQT2Srlj7J37BBidVgeN3/fow40DHGx3eXfxbBNjHDH75H89itvlyhhpwiVehT85zKQsx6fM
2Oyom52cMjpQH9ICTKrIrGSljye+b6Boak9OkcMi4j+cvyM0p0poFYBQMzqeqQ5/lvBLPWQIkf24
5aY8rL80e6Bx3kP15F2gJXDTAwwzcgJYG9ALIS3VbsHWerANzGKIGf1BMT8pVtEXjL/rvAcF2yo1
TfIdPxMoqH/in8QlWIx25GLcItcEB3bRAVY7eTO4ppt2YrpN6uF2TRIo6lTG3RN0iV7SsI5Yxrg6
UliPelqsIRCi0VY0jMpqeJMHTaqE7ih7cOLpKYHDhiLj5j2DUpxGsUHglH/v4Sfq7hP9eF7KGaW1
t5ZO/ezDS5U9cJx/3SYfGZr7xKQALZViQrkQhJQYu0/WTiN+bsmUkRpHN2n6tPHFtW/EatBpYle7
EMOqouhkFRAvbSi9Gw7DvDn7qTt8juiWuW1bPiHV/HsGXo+mpkCygnY2cVqxXZrjar0yTisZ80Vh
lXKwuQi1ixHK4+sfFAyHHDWIbeQZAHC14aaViX+cK0sN8afu7vLcc0cXhCvojml2k67u1j3TMIRM
dK0azKF5ur90GY4raKz75YzVxFVmuHVyE2zgNKFNgdH0Vu8lvRm/YOUAwfFuOKcVR4P5Mx6LTU3X
Sr61PUVEdX/jDT/c/WfdsZXIQYqeI0CxqQHdmKHwL5VDskOfwuauBLIcaC58TlKAWVaNmjRDQLkf
Qn9Rl++XBc/YucsrqeZ/OsPRx17zZvXplCHcyeK+1Y7/6BlRD7gm6EDWhe3ERPFJOpLieKOYFgQs
uCRR34q7wQZAdf/nPubrBP61ot3nNh5WgoyYZimtJIiqgB6Ds37DlJ1Kb+EmYuKUaVLNRsIhzwPX
Xb1KWmC/Ch0g01nbBVLjOCdTb3e9PwKGSgKOjCNlq/I9k4ekDjdzvnLFBvuprzt5iyJMdR/PUlwG
OVdc/9Gf5lGHTtzvVA1pVRSNc/bnW/mq81E2GiMuQdqRMGP48n3N9hWVMkfbdD/QUdqcU31sGUhx
LCa04LTEordo3l7t72+0B2ELqKv61mGJiEKMtvH7bpYoNEx9SBPjcFjIFb/xJ475OJD1Fv2JJ9DY
txY6ZjjTJx5bUULjykH+chx7yBJgKlchRjQQ11TvWLFcfnw77gVpemN3tGx2L9tk5ZqsJ7AHdU3u
kiqPpzj8ZD0syJrt2Zeg3Kj4Jc2hfOdenPHIitCHfYxlKmrv2/WGmIQi/3Be7fmrXlWRPvik5MaE
mYMHX+h88oEBuPA8Ike+m2ecpoL6xxl16zig/EOOaOLRss/MvENIKzdBzkODklOH3UEvw/MgBONh
tkl8RaRSGtqCQLMPSGk4Jh2VlguN1GM9ZhWbBglQdW3xl2fMRaGY6Co066yrOGXEzlBzbzl6FAgB
2o6fzhTR6faofsuI1q+sSDax4XZmYmi2KRTns+r4SQ+/PtVY339Kbr/nWqPemQ4tGLgpPYkUFpJp
g4IS/kjudNewNuSFo9K07OvJOeREIunZec0TP5hnj+2Y38Z3QLmgF0iDqux+pEjNtT4HJ/z97IDj
4xDDvQTanu62kvAc2PF1My8LZu0ioOWsLBxTaXb2x91dfyR77+uWPqLLw/uq9HsFjORh9SQP28QM
zdtJgsajuNV53aZIM3hPP6p3lQzY2zmN7QSYm/xOZZm+hChja+xM4plIncbmvyJJPwvrRCsm1Ig+
fFBoouFjTtqCbZTMfCR5Z3Wsi9jcxxm4kOlNynqf+EywkWPmK3wsjGsH/iqHP4ys+gi6w8Ksi2W0
cMv9caByzZpLRc5sNR83JgzXXp65ficRYHsB6xSWCMjmlxAyM2f+Qp827yGOY1Kcn2zAAEJrfuXV
8r51SybiQQRyUppHiP6oYZp7dpDW8t3aqVpbxGIiOs5TYVViDrarpZhybTyTnH3VxLgfQGN5URDp
raP0veYOCE5+7wRjV4QRrZXb7ZP5pEXvp8xz29JvZIcyzHmvBGcpiThv9Nd/nKV2b/8VM+DlW5kJ
KGAMlTijvJCW/7IBudrxuFZjkhRw9AG4HuuMpfywKZt5YOjDcPiW1aZSZNcHAIY6TV8mJ4WxaAMg
ah77Lycsp193kb98DHCqXjXP/vBvXnaLU8MaUtRdheJ4QtM8qvW4eE84Qj718gqMvjEoHf7ksZOM
nFJei4pOlgl2w96jL92EkT31dlu+vQTXRpPA1i4VVAKuniMVZhK7N7huceNKACUeHeFE4J34i0rF
/FWjrdanYVXfdnFLL2et8SLIV/iXT86/KcgB743chsS5Qhn76lAGsIfmyftgCvtmnJGfRafZFnYC
cxy0BV3i6bhin2yQUvNnB26B4A0lCPGgaaaFnmJljxpUg6c6+4gPZSFNeNrgDEl3JrA72S5/Uihz
CRuwaC14IcKGEvYmwYhWyOeftP+jsXuzFcw3+IhDLe//HrKDXfQiSrvh95rIg7TTGMOj3sCmImD9
dykir9LRJI3oNMgEC61hy6DylREpLlV2ChEQW8BVKvfv6+PNY9w2PKcfAMi+o223QTT6ul90huK4
2kMkWfrph6Va3zfqn+Jm1s+bUqwd21xXXzSxDrso0RZ/m9StyKR+WvRO8fLoyYj1A2jSHQG1RoPN
Rt9oQxyGBTqrJ78v0xYcFtVqp+bYL77REnwnCj3s5m4iLgohGRIESkv3KCRgILlNyrxcLMZsbNZd
dvoA6oqX3ZSoeHu5dFfnRE6SPfKdGB5vy0dwBnlsuphzTz2FEPIzR/VK3C18RrJ7zBUiezvdbbwt
/e1F4Nx1pAkVVLwUYJsQBXTQVJz/ErUtzXduY/gCBi5YD8eKCy/J8OG9GY1sk/3NicQwHG4AkMd4
RrCD4nSBuBTflhzfZLToELVLoFLB8/wShCYToFTBdRhI+mDaFYU1N8Ea/Y4bFJTNatK0Zhc/7Gqy
IOTX6JJwHWnLLIJKGmjre934p2rfkqgZlBJ1pBJ0jRapIRfNwl2TjSZVXdxgAW6ww3GJpRo8M2Ff
GuSjuoy7PPykFFKMBBfXMMwEzypxNFK2RIRp5XV4iLVp8dn7WiVPATMqw0ACO5Td/vCtS+4k/A+4
ziZ706B+k1hPnBz5XaQUFQf+A+/nIXp0c3ozSEZrhXEZh8sltD8JDnLPZfJ8yR1M/U/uWjd3+yjH
rrnfc9VREXDpiC3XVqo854HgDK1KHiZa8Sgf6h85MkvActmN3bgYUe87dyu8L7uhQhF+EGOf0xMj
qrO1nMcpmnwUJX5xioGZ3I/o7u2I/Moi5vkEJ2PS0llc2sHcwiQUFl0VqF6xnoPkWgC+Zjnvl3Dc
f1mpao+i+vddWpKQpy30csaYCUejHoLXSu7rBXwmAj+HNl8TpCQKeQWD3K6GnqrYYV1hneygTYrc
FptXamly69lo3MZL9OEcJq1Xv8TvAK6Hp9SXMJwU/T98vcJ7HD3nJ4zObkL8/mBqwAICg63/SEVS
wYjjZEIyAdrMnVjBoivcsGjgxvNv2EsjfYEO61ljp3h/PHK/wcn+0mTbgaTn9BsAMU5ua0gxg0AN
toTCXzGLCXhwNC37UVaVj12dr7G18gDWzEGafhFdoYEVYP2Di3pHQypSzcKCgjnBawIt0JbwKtNL
1/WaaTpSLYe4jC3KSHQCfKpAg8LMp4kEdnh9RbUGYJKdsvKxYq2D9WxbSv5iWsSf0cdts6MDvyG8
FMOMzWt3V8VB6JKOBjC4ET2Hm25QEpFdtI2CNYGI5SuUkZdcVXOzkI/1oKT9f2bhxdYlmSUiPCnC
v8rA0pOYWXEtNmEW+64081NQCrBKxp8KiVrcm7Z9fbABSJ1tdndDSdMEjDgoRZD1z07PulnZ0Qmz
9sqf/umkl9n52Ko/fiq9kpRHtZPm74VDmwX+/nPYYG/qemVqVOvlDpVlvk5hoLUD3PM/+lzzhntR
pyxg0pDlMJGaOsZPr5ef9cz+tMQVowf2xq++tt/Vws1lI1f0+4I3i7RcDB4P1Gw+D+ZKdCcjjx9T
CQnrUT+SQqRQvhvoonm/GMN++uwhVY6EKbbfPJHJUu2xfY+uT0n/lWalgPquHngyxYGqzgAMTrbT
N1iJpE2Xb7iRM6LoR5mZ3uX0DKrmqjFlbVgH8JSKuJORzQl/BtHus1HlldYwXbEWp+e+RMb8hWe1
tUDqDelmXKYwruAItP1e903z+h2etm6J2uGO3ePx5IYphhFbFlpz3YMgCFt0GVlOyqmm0qUon8kM
6EFqF1X5vSk0Zts8NnPCqAZ6rN42u6ZIWGTyxeycUGbGVm6GtUKlEI7eHIyPnbQoWHkjtkh3X1hh
Fnepsyx+L944YHlY7/yntulfzv6FKpZhRtSDdEWMne1hAM1rW5AnrvNagRkB6DRmTzuwQgEVd/wo
RYmqSwCpkIJDdsOO+xTCTONEHPNxnZvRJeVPEUk+znRdSK5LBrj8zR94zv8UbWXRU5+2V87TdBvf
R3WRz1diis+uLFOMW9qUBiHMLj2CZwFhiTvqrxQ43Dp8P66o1eBuKRYnCsaeQYGclnRZ21/kw266
5QD0UAZN8SMuBQkvYghXt9fQ3DEwFJy4k8/nEKfZu/5+SAMmQGBeWmfpDN0X7z5M+snhHMaq5ar9
i/l0Sqvu0VJHW537Fv21Zf2zr9iAmAQMnvaWkEM4NAoZS5pSbb8qlSS77912ZUrILjXaPeMwfHfc
TxGV8t2sCU1wmrHXYhkiuYY+aFzcPNue0a3oO3jntoCp75t80HMkIo00MND3KV0NBNDjWfLT2tnU
XJI8JAsl1HCvBFvSSDf5K4jFKLcixI1L1cr/cq9cIhfztArWItyKn5+7kDNrYsIhOcaAIO1EGepA
02SvuL6BP9G6v8O/qsMThj7hDwfOi4nBhtd9Bm3K/gDI16GMWSb64g77mPAmuKKK+QjZe+UxHnHU
myYjqzSrIW38jbJQaQR+8xM0zfq2whhkjQgE3Ph2e3TfbgYnx9QfI8EEhtiEoV586VTEG6qUSaRR
KZPIKuBAn5w2Ku3HWYp+c3YrUc1R+qBxBLzIFofnsTveVUXhFlSCI6d6FucioIBgi2Xb7oNBwkNC
94K52qWOpEzOJ2ZMcjD+iRPWjp3/UdJHRzfRsWIAdKOqkDmddgd01PlO8AzN8rdarNyy7uNzKtWz
oWnF1vRGmvIh7DrbJ7ETYROed6Qce4cLs4z/ZJcy0rVAcNMbDQ7RaZDxjJiXDSl2xrYohXyD8NVd
zlLUudkj60lWnRBYGKNYPcPAbnCZkO7/tKAKyBosn2iQF+TuqPjxiyS8BgYusfzbhYTYO34vhdke
VLsJWMNqG+3jS3D4yMd2iLqmig/ly59o9HYCLgUU7KslfdUH9b3JPCJVYPde502ZBPuOnYUx2kLj
aCfia0o6FO/fsRyjI7NHINnK3PnhzN2uYNCeGnlbBtAmza5uTuEsrrGZR+L/kTZAp20o4qiBOPkx
Zc1BlhviTbdTkRBNCYP8zD8ZBuiWtlKdLtI6rpFiHAHl0GF0kpebxBotz01UhtmWqfJDlVKJbJg9
iOqOnGzlZHKnIPIGDVNwtyXOJZGsVaDUz3FxbTfY33q3lsn0wRChulhFbb1lhHZ6+Wp/Bx0bn1zp
fq/OHWurptcKaQcitLXaJgD557rhyeHaSR75k80Ro+DugOoI5jw0W+zZIr6aHpDvWGwSWnrRbm83
mvTf/sFvCCXVkQ7WAZrAim4pv0yNFqZgidxnvHCre9qMbjqDUHgv5VqNL0NoYaR1HA9iK3IH/lON
EuMsHihD6KJmR+ofDsSZ5RO5lTeC+5hrODXUFAzGWO7KdIj58xirsK3wJ/Oxk+wkLXbrcCFYoVZp
dCQirtp9GGi9K+DUlkY+Qk3oJBfUpTPbPpMuN/WrWeEZmYR0ws74SUJ8fyuGDQpdugs9s4N0N6aW
++z0hBs3lYoBD1Bh25yr4tzvCN15CfOoSLMNWst+Myedqb5fSZrN6rgN+T7UhrG1fN8FyLvCQ+d9
ImSv1Hx3gmcRhAa4xb6XMuSmdWZDqOYAVfVRkZUobQGKVDBxJaJw3y3FSfR34N4JMnoZ7UzFh02z
FAELZYf4OpZ+KgfrZubKmOmNsLGUby1t6Mwfg/qWQ4P+lnIZ5mKBbYqLWhH0UdEtuW1RgPFI4KUH
9EOsgfMd7odcSJRfgotjlNwoc7zmUL1W1I1rGrFqD/Rv/haXiprzUmdaJel6FVFraaiS5utP3TKB
DjQb1mZTovYOKbK7pTvh3q3y+A7eADSxvX+v3v/Jmw9lrWHiBxhWJ6zOQDVx0ORCgrsdL+Wdlb8n
BiWGORLbJ4VH7uHrNUZCVTnJWpTFWS+GprZOKMjNmqe5GCGamJs/15wR5rKrtE0B+k6rWyVMx0eN
nIsqPt0gwi7HnJeMMw6pCdNl+11RAxEIw3s2a4FZwYehEfHC5CwkdQXIf39QNpkOlfUY2DMJ0vlW
vVO0obuGPYwx+jab3jDJu3PbmNSLKznoDxdXPfASBsmq8oDr+qMwvxngdQnxFcGgWEat4CxjeFb4
7CRclZpGDH3N/7cBtVb4EoHOfnMBjqCE9OZfF8G5bil4FbQ2bwokm4V2MTE4UEFsalXKK9D7An7v
O9lKsq9rlLI8CeQY6EVXNYgDD8eDpLifhuF2fy09xgglucrQBM2oewfIbTulmGvCrLr4fnOiEOLj
bsUjjq20lozeucT8GKrMxLcsEYwcqYzbmQlMwxk6Vg3OwVTHHts4PuuyWhtlcm8GSdqWxNe56cXh
jY76cqkLtVnwQ/p7t4q3kX7s2jt7pPjqFB8t+kaQ2zIcGL8Y77oT8IhDZl0140Bf/wH9fFw8LxOo
GBA8JeD4bcJZEQw0huYDq47sA/3emK7wG+Bz+lSKzXW6EPsCIoaohKLwaON8ayL3ZsukQFOPNG8b
Ez7kFMoDeVsfoNlGSjjt2yovmB0gXOz3MePwrGy0lkaFvMXlijJx3p1p5tfu8B7sAxQNJpX7NHRS
NSc+6+0fWyZmQrn4QeSmPp3jJX5QJJo53ODHIUhVI8/Qy775Cib6lO31gThx08p/5iN8jzq8zSr4
owM8EKEuvMuDkddu0fLTB25EpZSN3TU7zbSZEaNMJKxAIF9ygG7SjkX5llVKsJ9go+VnZWnBMEuz
zD8lIdK9gpo0VXp+6hczeGx8M6RCof91/o7etEWlqb4mu3BdgV2e9OiwWweOXDflbkGJJAFKGBPO
5ilLvI7ct0Qdc2tkTup0HHoWFgXF3yDlqIxY+XZCJnUgNIs1rPexY2qocFbOqM7bIhP3TA88vzXg
CPMT2fr12Jqdy3U7+O4Z7BSclkBXAK9+9Y7sMqNfluOTqe1TdQVKJ0VaPlIWXSPG3H6MWJhKs+fd
S2q/1863gEu3Upvq5oHBi4HcidkCEgf5mHrDuXFFumS4j0VYYLrYFNJQf6gXnkM70QRL7muRMXlQ
0Mq4sh814DdXb+OM7OVltW92btGByJyhEu2PVqff3slb5B5GxZkKLQwd92UGOyBp3ksVwPX9Z+Ft
abr9pJe1kZFTrc/XApy9B7iCYPq4bDGdHhcxbF2waNUEMBHA8djl/UduKyJhOA9F036cF/aWmz6o
h7L6WNDJ7sLNoSE70to9hExr1zDz6DToBcfL9w+3Jn1xhM6YlU6PNtdVpkll2bUXGuw5vsBj+Kxv
biwhBLTvq6/UF5hfjj3kTUWqEp7TLcac+JIosBeU4dM/oYr+dS84fN5V6gwbhfA6zvuNjE7EpCks
gOnMJwPQcRf6eQiFGLlSWc861GtNRVggfaOxWb8ID2XW86ukrMWky7rBjQOT5NK4r1kA/xFikBzz
W4Tvjh+5cQfGushcWlZnxqT6XR0Ct2zpE2rsrZ9ZyHhC5mgnVIO9mrlGw/hSzGk2JE1Ogokwcvx+
QNB9EtHdlZLgRFR9Co7LxpOJ17eGuGpzkYww7inj17KZnfg3ods/H72FTWvO24wrxBmaDJLbsQoR
NEeTFBg5nSkd6AF0GVf86RmeotigIXRSdXRLLvCKw5FpsOe7FZa86GwKlEjnRfDgWiUGK87sHEJL
6o5HFzoSaWGMDkx7KDGGUIfBTERWzAxcBMXaA82D36U6xowvO6siq7BOvP+kK/hPMKVa0qq35Frx
ssYMOOxJYVZ5KT1V3uBpTBd6tbD/D5GNV9VTNjuzPlKb0SdKZQf0G4xz85ztcFRtvm5TcUfgIpHs
raMIaGDKvrpBSmDtO4AdHldadVtfiQ+5k8WzPqctieG8dA6/7QLcQujp7hDF/u5fkRPs088cw9ll
UmCDZnUFBfo5ebOXe12xT8cynZqNyVcT+KQXEM+hScX7/NYWyl+UwR7kbtaL5oYQtBx3BCiC5fNz
OT6C0o3+wrdFkT9qOLrZufka8kmE4Fxpi8wmUDdQPBfTXXbai7Kooq/EgAeVv0XvDl0NBInQjox9
DFLZd4/PJj7RlkUvXduRepwPVUcMZPaYM2WOmbnrbP+jqC51TZhY4iDvJas9t3mTiuZ8WBOaMY3S
D3b55a9RWgEcxVtRlZUsgEhbyrabZloL1//sb0zmSLbL4oSSnM1JyoMYSvwTUDuTDZ8X56cm49Pu
pH8aLkwUDbpk4A6L8BYRPY9jGpLzWvMY2I/Zd6EPDFn0vFPTOrQeJ0QZZhnfN75fQppJZjXRWPd1
gXBDybABlvicVEIBiEYRBlm87oea3RzplJI1n07q3nMcMIWdGRhh5YixkkkowVImyy7r6yEQCyfY
3qsJM/H9yPt5pGUXQGAqEIht8KfKdCyhJ61gMH1ZWDxwCS1ioOFnPSuX1z1aDn+X1swnsyGxoGZ6
5ou90ZOnG3w6Zwy51/OnPEwyYztsKu4MmEP77D47zkFXTvgW1GT2WUqr0bgZkCL/jgeRIcswps84
s0+B/8wehE7BV5Ih6iQnhJGcWE9VrEMTzHjdAd1sSTWSes8NVj0Ai868nt/ktnWrHfpHpnIkY79E
iTqA9rFFqOhExunvebF4uhVJSBZNbwEMss0Hf/iEqUmBoG9WarbevLszv1h95mFKsk3bS9Z5ky4N
tYC2ZK6DZc+huRbPBr5on9/whyt6omu2+h5BVGBO+hPJ9JeIPdEXBnzi1F0YSuosGlKSdYRz+Lq7
AJZaf13q22xxsvLoyzMfbrN1RxlYsg3nVCCTlNmxKThc54TW+/nbTZaCRnlaciilKOJWxE42lG0D
YKBJ1sPXqdbDneCSQ6JI6pMbkWzI1eXstjGABvA7sdzB0yt+cXYe97Dh3SSSUFsh71sa37vd1s6v
vYRiNMId5zwipYkNSZIVHazs2CjZGVhrqVyGBB7MKIXQGP3ROswQmIw1P8bQ/iib5REvHV99rsJG
83MBqOHVrid2sobfzeu20EOj7p2wzvwkyVt+donRETg985FhXsCgpXw/hmVHGYY5IvVjS2Z7FSHR
yvdx+5EjiMnjyqI7yrZdqlv78bMFNag5AuAzFxEBGjftR3y0xftjMrD0ULWMtkYroNmd77UFFXej
TWp0JBOCt3bRXmA3Vn3bhDhSjZD4JI59sBzjWE8M5EbI34Sx+2lylxWyWPHEl6qr024eHqt+gjhe
WLwiXF+sYsjSOPGw1T7KxpBi9toXisNgeJenzLqgkO8J721Os56Ot6iNIl2aAZ/fidwh8s2Wqrbo
XJYS6qwqFq9Gfgkpl4ktOjToBYIK098L3v62WL4WCniMf8LVYdd3NWgUkR5CtZimxxBOl721Zbcr
PzZQ9QrtOPkwKnuNGh8KufqwwIM8rWAGD1NY9PQri9s3tTp1X8xysyp5Q/o1hSQTSV72CjseWsin
56NpeFtt304gOmWd/1TjYTvXqBYqQaJy5LyNycnqKXSaGQaDYu3yXgkxy5EvULK2EbdfkQrIe7Na
krsvGwEjA5paLHyuUaDlg56E4fQlZSn3o1nXZUJuiZX3C2hH3ZSi91na2sA8A/cc6nHgX5/Fh52K
iW9vFTsqjBCwFLAgVqBFNIfdVTzuKLMxCufTU3WgPjoHED4Uj3JdSAT+QW+zKIgkhNL/yF2rHMVG
aZ7VAWixrhSfwoQkVPES0lUMmVIFPGFAVFv1AHGdLxEofzfWtsFhMoeQEUsS94CaaGqCFVmUmSGP
oQgkUZWCK1ehdUkxDh87Hj9lGZmTE0oxbd7/qFEhi81DzkcingoRYN6DDCZ2lb1ohV1q5fGI4GM8
DpuoJSg29u4yN8dGVI2MZZipulKZpoWl6HFu3786Yh1R+SCGybS+1eebdlK0jMO89kjKeJngLFZo
TRfBpSYXGn7vXAeztdIZoh3D0WzvYuOoFoXhgHB6CoaC+vp/ulTejcYbblO8VrEgYbBY7TOr+hqH
17fEZXvl7mdR0TaPWuWZOHjQ1a65dwzMSgXXoTwwqD6xDhVwtVwpK+xh/vVfLsajHJJ5bfrTBf1G
NAuNGAVxqQiLWyx15vWbft6w34SZ4ZHRZzwW3Zd3RGtZ/RIFvXf06lU5aE7buW6ZIm285fNyVUPN
8dIcD2WN9fdfZ09Br9OfK5Ecs1Oqu/4Zl5KrtOxh99gDhFFSviTu26rGPLfYYy0Pef+QD19IIJdf
5G/Y2qrFePTSUqKTAoBpjul2csmxfTHtZHu6BSddbaT3nZqj6FUE6PU/yZaytuZWmvmxz14aGfV8
oiD+DCNgmtT58l4CwnQ6t+awSwmtqnhnoY1gXaosrahXu5B3fxcFaW/3cQkQXASuzEnjfhqlNlrY
hBmnpz66Hpg3favdewyaOpVhr9DtYUBcbf9cS7kCwN0exAx0clstnR9/i90oL9FoUDZrXE2bpH9x
gn/ufF4OZi3GszUXhmEZePKk3xl61zoNVYdHlYPf4IpAVe9kei9J+m1WIOl2Gps0haj2VfqtA2jI
N0q052V7Sv88wum8MnYLWzehBycX/Yx6ZoUJsbED21++pz/qd2SXX77YHJXA9SROzX8V8Dg5ncjx
nQV9h4wcuVc/LfGn6epgkkmIEiVLd2HrKxMH391vwEdLrkgDncUd6dPdqCt0FzPu1riM4JPMU2yn
NucaFpjLRXo1u60GlSbb4ALujfmFPTtuQ5lej2LZrV5G+8APaJIT91m4u8PoOBWOYekBm2HZiOYr
m01P9Q0vy6K3+pFJ4N71UIWQmDEfIgis/FkGYXaj7hDwU9zYcRDuZIekE3y9RLLcE8P2VCZWAB6p
GI39a9kYofpstWW/PYlrbUi0cLNuXmCL28Jsc+4+fmIvhy8kdLCTLkBP6xQTC4bVbHigAjG2+lu0
GvqGi/EVOI9fjNuFoy5l2K4MfTTTpDohDT7igfaxEbiS9L/p4XfZ0Vf3zZ8TMcZmztKUYT9+Rpsn
vCNkHEaMRk7VVsRmxwpXY8txAc5Y67CUtudgdSwvDCFlJYGacLQM/uCtIFfqYbK4kkCcZIv0U9UM
B2EDYpQl4EQ6L4wSynCY3eb0XWMBP27Xvo4UMqbcKhD/WW1ezlMc5EGtpSa8lXwHC0hPg0l76r32
rlk5/OXoZNWB18QmLnp/pyhRQNO93j7N3chzozwQulauOlfpds70zfFJTnu+PmxO1R3KrzwIl8lH
0JFtXselODvYCfgWlS2FsUSs+CNpolNWTxKOrEQ3KKJvWBLiPVXYqbLn7BcJaHh6aW1eunohHIck
IykRmcIY3yh59kfizM4WdvLeH4zQ98b3bcMVcn4SWMPdwxCPKDGn0NFI1XrGCOm4A7WhRYzY/VX6
lL+LJ6bgopQffMBeMruDdoB5jl4inIStkPgG73xlboAhN8i3/P0K4FcfxS49Fq8ysGsI74mBKdwK
xmg9IJpntQPzWC/EQTCUg8WQZ1P9NhLkxrSVmo6uWv7CPkopNBGfvKw2xOiAIzU6iDJTxur7Vlhi
mRBqxww0jWe8kTzDik5ZeP7nfJ/XQkfyz9ZzDkrfxnRtFi1pGHpoOLEIMdTMTdBEdp62ZNwn5fTF
V8un3ZN4o3GyRlPAwmXzZ1CQfzYPbbUsJmEY6BNcytThCAiu3VdYLbmWdJej/Mmpzj7E66UGIizy
NXA41sw5uoXUeZsr4GY06OMJ30FZxZ/OErOHt90TWW7Wa19jGtDxGJHwrUV7xzukvbjusAYVg+cq
enHadrIOygyphvx0XscZ71TREVbKT3E4jqKvWkfifmRkn/0byjDt+ZiE2BAfs1Mr6nPK3W3zJNab
aUFoNT3dYhd2sKsMR5FTkQuzw+qpPw7nqMIvCYvvyKgii97c8ggsgOCL1rFKQHX2Jrc13Uxbap/e
7/DDOzEjaSAEGhh8Jk+cn3x145mILuOiAnd6I75Pm3BjpygbLZXlivXd29h5QcFhEK8I5fF19RIE
5Rc3HOz+OISbLFRnxws9qupCiFfQeHCgLwGT1VLwPr1mQEnY5si3REXtVj5LEyXXf8+rw+JY2jGj
yuSccckeN18lkbhhiwW1ImmasJDWEnjBoLkCyGhPRd5dySweatCojz+GJMXzhOwPQYtqHWF4jHUV
eOiAq3bluBLKdXbmSP+VW3Gt0tJLS28iKJfl+QaknTVqo7KCtyjTVVopC6EYuibcyHNdL70TRA4w
+c3DFwlQ54YQg3yTiN516XkqtcwxSJaRwAyGvUW/wCou+ztjQ/Ye++qSZP48Fwa3HBtsKpcOflm2
8hjTHIIJLipBdu0miDQJop8Rgum+PeXNiFKqfqRE/yJ9hie4Kn7I0O61SW6YUS/8mPDinpcQ6Zc4
7xH0WI1rp2aznmEK+aqciozsEFFYx/cfRgwjCpXwuzQs+C97GCVVpYeStlqb7zY2Ne4qUiO8vHUQ
cRR/s5lw53oaZ6aiL03Ai/ylxB2U9MSwghAF38nX8XErSuS7GQcy/x8NN3Qk7KJVf4cgWwpRIUbo
Gdqqm+QX3Ku35b58J5NFZBru7a2vtEmqUGqGARByjpnlPoPT274+WJq96xtvBKFP+fV+Ue4n8Hak
3w65eKrGDrIq17nl0M50Thp0n8Ie+7XLYKuOkyMTtY/bl0dxSJ87Bcy8M2AK7ZOQm00dNNFqfZDK
OzBy6F2T+LwraaxiW38VbAeAORmFJGV6/Zt4Lm3dvqdrraaphiNLhNplen/oio+rjQQhqZKkI3G3
YKplRFHiTEXEmHCjJ/73zGWzyLzFsHpkFNBuDV6xP/Tcr76Mlswx4QgkkjFfyetrRNvi+ViV/iR/
UOObg+lhed8xm9KJbNFK6JMwAnuvseei9/AZxy1VY8KqxYWj8KJN9/Z/XHwfyL2g9ocH6i4ZoF/P
CGEPopqFt/sdZCic32+dhf9AcONyP4JR9ViWuUdvv0y60Q7E0nx5F5Soox/An/ymPXXMJBFPLAwR
f82gyqOAh++sKCTeFX0IRXTKmgOJ4bgxyGKMITjZ3E4BgXQhlqR2ejuOjhGezdCVOSD1wvoh5yhw
zGDiVqM2YkzvMbm1TWZ1mwQoZorZLjY7FEwkQU6oyq45F1bqpABuQ18flH5RWBJMQ+ejMTa0lrLP
XyhLa1itpPxF/8csFKqSMkiVhNBFfhoJGd/fjVNTkvI8ntfRZ5Up6bbHwNiShaok1xAIVEyGrcdl
7MkcNl920Kmr1BkKOiTsS22KIVZM+vTJ7Zh+li6u8bd+xMrzus2NaS3PXVlbcPFwdCHKjitTbl9o
5vki+GZZMGKJ69VndEhQrL1rQNtg9KLoHy/yQ67TFs4LjUQpB5QWt4qTleKY404UtL/26nx9xwEj
23omsh3WYWgbNJhpfAeBKoOsaCTJgXBlxasgLR4xze0FUoVV3Y4Ebjfk2Y6AGEWlM3BxaXZQ9wLw
KyJxwWxpoNqBDyPSdAoAs4puOlT1xG9Ad73OcCmDII5D6PmHt8ZS3AW1rkOnQM9DAf1y4XoINh2H
sjUPI981UAK8v1rGAmM30YJ/ygmjuUm8qvqNPN7imlXmnuLglGsYgVqcESpGIQ4E0zs6VrDNql6e
EwfZkI6MIT22fCXeXi7hCPIOVRDSB3tfy0frZvbSGsxYcsQzwvTxZpfi290uwdQPFlWCGtqZQfZx
NdDaaiSHrXRUoj04Eir6LmSseZVUL/C/3YEo/iwiRLYes6CnkVC4jbXlm5L1+JnUM1sPu+0Kqscd
wOiZV0O0MzMeOET/cgFEO7hGD/0ZXH7JusMttT2XYpHTPYwbZXZXY8zceBuTRj44+eiMXh+ZmIdN
h16fXqDic7I/+VU9wgHG+UXtflYPaiFyGSkIo0ATFeYIYyiL+kJro0wLyraP3RE9A/bHyrjfFRe0
9KSFsZuzQZ8c17VDxWffpRfNQKg0hgKCkoZww/VqvX/3PBABKtU4wpu/ZzovByu7k4NJmcY/WVDL
/9UH9wcxdjteq3Csw5xZrx+6CAbjkYWAdyerwSrH1kjbm2wmg3Z3r73kEWs4VM2k3lajw9WmiK/z
6CB0Qfs2IhmHBJLXGy3MXYsnjNV6dsLkxXZUpl3nflyI71tRaLPDMWqQc/ghKUTBI3zhzdDY1ELC
EssyAo2EQNj+QN3rS1NACdFVC1iao3Y3/Xbl+0pfjXOrT/+sPCSaowoMp/9XM5m98iBF3ZdM57Kr
i2RrhpgZQMao4qq3Aw6zLmUdo+iskgp/W1gL4DkXstRMUOuZwnzzTMyr/G6Erbrh/80M6LZxZobq
rh+ONFJFy/CsvoizT0SZHaauFeuz2tC/Sr2lgshe3noaSSZYw0/P0KWutv/B3oGkeNB4Tq8cBzOR
BKIlkdRVzPp4uHazXcHJ/kove6W0rBaCbgm9MD6i65Q+FjATlwkRp2KU6Y1KboMAh1D65YXgug8L
ZEijNLBDQ09m3EgHcgYl9TdyP7vVFzz2FtmmB6mwSnyI4ulTM+ubTRNe59LBUP7vi3gYxrSo/dyq
o/luLrarx46I0pDFux6xBuf+Wl7/PUbOefWEMguao7vWa0WW5aqQCEyh0Jr4Ql84TEfd23uWxMZb
wM0fCWsfHcfeLGV/AZPhqlUjFNVxBdIHc5JM8d1MPYcrk1e4WzDgDI7K3lhov++6gFYUnijTZ+ng
lCfF1pAJDUprKc80piQ/rjdNstky/HZNea2du7OvRLfTxj20SxGyU/9hknbniprKKk+onGK8MG9j
OmzADQW30EyS7Dnaf2mx+c0z9xSJg1umeFUEyXaxGmDcqTOrXaNawzQlySIaZiJkoDwbUTm9DcsU
Y/ohmUUy7+KM6Ckw1iu9yWlzK7ScsRsUe2S3WBSnEP9Kk4KkwJPYtTUj9skDCP9Wlg0QZ/JEseOt
F2KIze9KotxI95SZ+8JNwMcT2W8psQjI6XjWwyBy7V7qi6CyRlfwzpYV1W5mX3hp6Cybhteqas+P
/Mr9Pt/pb+9EEpk2u6muWajhYpjMIcW0FGOrjX0JA06AIRb7yAZ+sArUkzfejFmxtOe6xFVtBXOW
o7AShU3rPxyQOVQ/qYr1SzcJd2I4dXhL9jxzXyQLIbE6r4C5VOpLCRmowWMzlzBfEIYLElfar8na
PxttJTZf86rfDaORtHbTxZIDh4glmoIPEDmexbNd7MOSN5JEoDjgMQo1nsmbBP2WBHwi86rvLcEv
dNliQBfYomZA7hPljwtg6kKu9LEDrMgjWziK/lJVV+s/yVPxOoFodOP085UKMq4htCtrFOLw1WBI
3SxpdCVMQVAUqFFCc859/lTcW3Pp3tDT4scElODdLOimCCcYJkLesdkGIKTi8ee3CPItANtbdz8u
k7jiGjyW2U8cwVi6VW0fOgTNOt9yBxcfMPh326y8kEpE3j6u2e9n3cjqHv0PtN4HGZQn6tYkcMw+
K9QmAkWweFaRXUaj6VseHepc6CuZ/bZFCY7p3SXFZwwgFNxZXs2Z8uPvJNaMb86GUdbhMunK/Tnq
E/jt7lQZm8EKzedALblL3rN3xe0GK7ZzPgNRWLaaH25k8R8vTtzDAXX2UJXUUk1buwD/nbC5NfSv
l7aMxC4bv2vbJixNdI1Jri+WhbKIcvefZjyhgCbRD11p24v72m1XKm+wPm5fJ8oEBRPawieeCkdn
1GtsSRHy/lYX7u3J5M8hVuZQWHKHwk7Vvn+QqP5jJSJE5DBT+84BqwtYPvzHconn9a6ZBEqUaA/S
+tYG+tmlZBwzqhgdpvRqVFgYCcpIdBjHtk5CJ5R0TH8gmuHiR4Q/OnGY+VSXZIGJedyp9m3fOJMv
HnzxmLa/hYC/mUUT/V/3qRAXx03jXZl367DpVEayVgcFBnBSZ31/lRMJgy7YVCDJaWqD8NTeYB7d
tTHO38UtpzhcvDMHEcYJJcROS+3fGCkLPZvBPPCPegBOAUVDZYFofBds4P7RTtKS3Yl+fe6bCp7S
khlAafQP3i/LQG4JSQOS9Lmy7p1R+ORWZJ1NzWlCKtGqK0MuMqPt7JiyoTOK2hghwe2bgo6wtLgW
ubZzoa6w5Y8LRMpCxxryuh28KzO8VNrMFSAXCPJL5LxEKyA8NsCSkzAvha5YnH+Hkt/CQAP4kJOd
3c8ri36r5izJiEW2Co77PIBuQMQlJlhnhrYF7NqwkW53DcnnR/O5BWfJVY7sZuAt8QLxUnxcw74n
IS0r0NiYjhks2QQ/F5zg3Smjv7UKM+6mLS7l4bzRaOFy7ZdITB0Wuq8IG89K+/+nW7Th/QSFBEHv
mVElTwRdMdxJijT7D14z5A7oTf9kK3Yr/Pm8Ai7PFXtWgRNWkKexnIOG32bZnrixmzWKY8MCyi2R
c/XnNxAvl44jnb07zWirf0Q2m5TflCHepL3Kcs8C49/4G+QZoCPWPZhJNHL8aQtuNIleVp1axkbM
WOLCPkiXT6aREEwbLfR329ohhfdpE+ky09KKh36dzB4ZkekyRYXlyXr3XApsCYwrBaYUUVHJWJvK
RH0ZjA/RSdYCZcvEXLSRrCzA8LpcEq347+3q6KdAXpUbJXBFYXuvjgCJHXlHmHBEmVzoqM7IgBD9
vMk0gagnMznryF8y77FE5jnWp95McbdkLPilmsaKkf9YokKMO69dW2EJR5XiG+9R3Fm6hng7LVA4
ZdN2zbCEGj9ZjD1Og03UvLEyRBqef7cdM9KRFkV2QZ/CYpMmiuYDuT/brAoRk7mxwp+g/xG7Eg4u
wKhT1PpiqXjasYg3IEZBfj5Ntz61SvYaeCG+7ve0+zHr0Ea+nPat8e1FWrpeeBnRea1jpXFo5tbe
JZNumKm2FG57X3rKrQSfDxrbivJV1qFhN+pQSLlRL3bGK2JYm/SyaHaGmHa7e8kAdURr0dXoXLIG
l0AkrEN86FjFSLqkMlNwjb65y2DaWk4y6/WvphmPRnR4EIjGiy+ckUTj9CGMI6u5iwsHC7XUhil3
kIdinQSoglUAEKqhd6PB5Rzs7UwO+pD/Fu/o5MM5IoHEg8QdXhs1i8KbWc28EmfkyN9CTRa7iFJD
pZZl0CpHUW7jTuwZFrSbT7QcH+sbt3UdgGHnYu1IbTtmLaBh9hzFpbdpc4+JAYav70wu8OAU8A0d
fNkQ/NWTC+iFEMIOHr1mRgKpDAjJRkWGtfGJgJzktCUNha/Vg11pOffbheePCIn0ByQW7AFty9KQ
tSF2YlMOqiUH6hWm3S7Vn2ZxiKzS/Op3j5gCuD/5rykPOQedytY/4Z0kMEIncI3hnwFi2ROpQWlr
18vG5dlekrdrAxXa0LGxliPXO/8GDRwYIPa6zMl+NlARLhaXTh4v8NqhCg8UEhrQiS6wV4d+Q29l
u/RQE+zIixAu6tjq7SQNfiqYqT7Gqcl42n44jzYnCxI3/AdlcP6eiaeZq8RojS0Ir2YH0YmoNRGE
MKkdsPKHXs5xdMVZ+Q7ataIxWozfY0swdN5D7Xcc9ARtBdCXvWxOR2CEG9IbuuF0d4s9x4POW6kq
QP4Pjw4sCTavAAeCWq9le+wmZH7DtHPEGqrmZZQi3xnH2q9hBp9JG1+0kctCWuDPcAazyeoaTT3q
AtAQqWOSOrEHEdPvKbhpo2OlcUtP/oRFBFxDZS3OilG/ic4iFUN75MwVsYhD4+JXJLDviXSixwon
Q+BAi3ylTnzHmL0ztsqnP/K/6umoeRvATl0L86ndQccQ/BkLIGI8I9Ks5R6jU9fhG7AGZ9Eje+mJ
uY8w1TmCVhrklBT1PMac97OEN8G28iF4T504oUcbCVJ7mp7zkD5LbW8n2ccAja3zfy5V9Hi847UF
/tTaD/8svPbqs2l+6W/d4/tU9QMI2/3u+tUWz6dA1iNb+AZBA+p56pZW7KlmC3IxiV1mBKL2tfD7
M2WNYiN+4QRYdP6YIMVhTTwMdmmo4oT9U9009DSJpu2PDs20VNScEaG0bIZ/WLp8BTrkI/sBhvIk
IgTXtb3n+YMpWQPkpdmJSg85jTwderYcaJaIaX/hEYlKRjGFbzYI1usRUCxcRIOpcTUKTmQ+X5Xc
fvMk/j0nOoJr5VdIkWiq1gUFM1q+H4O2QSsszzs8pdw3SMNSfS7osgXff+cO4f3P2ZC0hZs7kgtz
zJILQVTktjoy0nTXdCQm1KF/hH8mJ8IVM2BPnhlwOcaqkZjChZBd52TgKbiVZreocHUtcncR9Qm0
6cwYNJmDCAuwpsxP05S3BYVlHSK/Ej8vYV15d9NjvpZrKuKQ590rI21nvV6qDGSMySUkzD9O23z4
ueABZsHq+2OWAjPBhjwdYIymG+fN8nZix/2HIJ4+02J6YnIvVtYf8tiedjUm8ReEAocPWDL+2SvJ
TvzMMVHJ4iha7yN/a8PkYIzVk0zWYjhFr3XHdRrDKsTOnKc31ZDAoWq3KtaE1kjkqCY0cB/ZtBRt
91X7sYQYPYmu9qm396af4ZhIOWhHmWDpOLGpWVF9hJOotL5Ti0dqUWYDed0CZdQZrSTIFPkHkJoR
Mot+bLyNztPv6cKpni0ZaHvH/nZ158SdTtnmmpAsb3ewnGWBcujYw9Ew6Y7739P3EAIhKxgpEQ7i
+CSPUW1EbVtvtn8dnb+bNUNGvX2OBYLIJbbGOnUDi/ARFfL2nu5pU6ZOyfTctjfc5Mpyni53yHhR
vCpq6/xzRkLms+1SdpQao5K67+7GF6tjRyi5elqsFd9BtNTZLWofpDOPdDys8HyLzoxqilsikJcf
jrwTQP3iu4LmhBzueMeWV0vqXJxrzu1+hY/2DoxuV921MpEYfCi5++8GKfpdeE8JLHfojmcv5HvG
SV8L6IUs5glWK/LeSn4tXJMx3GUUNQ8IAS+lJ0ziyxxCAf7yS9P2E9KJ/kYqpHe8YWUdmdHeSTNT
OZeiZxqhhLKsxTWYXDdI/ve2ZoYJANy3rnkLob9Z7d6vcOmAj0/0y22kURy2BCq0uv0Sa2rr4yR4
2aVqTKfL+UJvMAxvQP6CZGnEBBwOelOpLYhRaXhAWYO+d5UQLaruFGc7hfpOHvDHoAY5gRFxD0dM
4e2RjZwu6WpHbel6H7BGailZO7tC0dipWoJSG+WQXdroakOvflB3ASdkQVkufHswKPrmsxI6s4p/
yMn095DJYDZDLnOTiE2WpiuQKGBhfOUsi5axYtNwKy9+GTmkiCRuHeM9DIbUlJO5b02xK8g3xuwT
Q2uHYt0d6UZ6VENK7Qb3JHJ4vne3QhdpwHfoJjyrYXZUuNe1JSTNP1J+xNU5yAxKhngPVT4JMu5W
xQGx60Whq6TToWuCDACbvsLrBK95jIXsT2/SruNaF86E+9KKN4J6ssGeZGYhUtH1EduQneDP0fC2
ZiPDWHuF0U4UKABki7WKDQhfF1LmkXpZwAVKrZULrr6q1wrIP98NtXYAdFRnafCoQisDmdpNqxQM
ioHiQT5HKxoLoLTcZcgHZLYscERTLRIy2EAq2hu8zZJv2+/iyhY6lYZ2lRFaXF0KKJspTHWsu3OH
fpljijuspSR33TRqoLrWF16Ik5PIBaTA3ew/gkeTnn34ORbuboIYwwE/3nx7bSM+Qg7o33QBpfL4
qklm6KU6aI5DiQ4vVkArosMgapXj3btombhgTF64sKkx5yFl7wFo/1tp8yDEJNATfJcWLlTtOCNn
A5dukMIS+St2PPkrffWZ/+7Z3V9Aah4E06oHuiNbxmflHPuq0Kcmzx/wX/2m/ENtr3VMIwkkCaDO
24l8GCZwSqTRYIWGv5OiBq7dHDuDkiZTX6vX/xjn2UHxiJTqumWV2wk0nTtvD63iqGR8aie0FzmP
TzO9Ns1uAA9l9W/W0isiOnAZolF4OACP4IS3ovdwW28mu9xFs6eQJVFSNd8scSz28jwE1FNb0UvA
N85rgXKDrPU1kOICvRi52lK8vZSig6pCA2EZmaPB89n0hrB8J8VZRjvUoY6+Lo5AOmghjs/n2vxa
1nUMXHLL2H5zVHdPOZkfvDjdys27McT9l+DdXSPFqII5aFKexfN+jxWjpZroD8ic93WFyw+K3IsR
AUM6r3loUurXxTXmITWppN+dTr1ZyjRSiZrh1lNmUY1+SWuh7cMBAlYNQxRsYhm85EKLTd15o6bt
Gf2J1RNE1GlRDZKfqPWFlR2NuYu9+TDlbrhIGenTgSpcbfGQMZE2TAEsZ4ptqnrlC1di8QRWi9Pz
mKvviSzAkAfcSIPFy7UnqDHsWcULqJCXW+eHqp+Gb5pW5u6LzoOABjoY1La7Wuk4Nw+qh151n6eq
QN6h5+PEc113591En/NfHs64zUtf2Hv4C6oLKobgGb6/FwyaV8higdXGLYcL5WDk1/VgDcz8zQdZ
C0GvFzcxHYfaAzz8fK4Eog1e+9akufT5HlUM5hjzKLy1byLGQjpCIBUg7xZoaVLLcb7ORazpJtJ3
z0kQ9ZG5gWkSAgVmAvJMf/EUl2h2ZMVxutgDH+/0L6rw7K4q9j0p/dL1yeb9OaXhFjT6cBDQkodj
5YB9pe6W2GzK02Osax9dUr/GK4y5p/SrmQCU5zXNJrQ3zLKIZ/PWOZy0XTigUKPhocJCctkw2bTI
5y3J6D140Pd5s1AU4cy1JI1KMNR7bqh4bR0HkvZ1ngFpXUXgB6w4DxQpmMwyVQta29ahaCZeFy2N
4/hbVPYHs9aVfEQ20+yrlM99LhhUxpMoK3fToB1fR+URhgNhrriyKO9lmWWDsKJML+x/dKtBDfq7
96I6AREoDGlb1w4xb3wVz+IPnFw6/Xq/VfkTYry19KZ8HrtTeRkJ2WPBtGJNPseBJShuDB7tC6hR
HbudqMNPWcqfzmeoXSxIoIfk0mtuZk96v5vU/X1EcoTrJGd+iFc4RZ2Ir0rUFjM8eDdcVlvT2ZUZ
HLK4HlNlMEfTR+MBpJAPsAbFuuBi0gUiyBfL3sVDOQ6Xz5jzLFfBeHSLYY07gY8wuJ8QDLgz9Pob
H/n7KzzVK4xRxarnmihW0eSAVqrgy3msnps8hFcoTO8vI94o+wpeqwo9UyTYIdjAFQszc7ShJr4r
aE3qGMHEbTPr/w9eNr34uUl9JtpViUZfHhdxamXHbkjy20fokmBWcXCVWTVdO9gG4uNWulZx6HkD
eQvtX7FoLaNe40OsvK5qKaNW6KbN3C1UYRQeVHG9l7byffrs+pjtixOVIwmrasMT+RsleaHadU+u
xqvQBg8JexDx+KUBlLwtwP7qKDfufXvvOBk3cYaumnqDrnBq/+qhXJmelJMRqzKVQlDL87xABN3E
btXSTEP4EMW6AftaVXW7f8YcesmK9lHQ94Zuy+8Nvg6j5FgRlADEmNnE+Lf3dHFk912E5RbmfbiX
Mrci+u9eF9nOdTvqijOWVNmuW7uPCO8ODP90eoZwABEbH7LLJAPr9qTrLzVWAlrjScaE6Mh2WSXQ
zAFqTdBLM+UCrS5qfDNoa9Jm2rhsD8/18Myr9uAdNgSiQVmjKur6DxaDUCJKbM3/4J40P5YBuLAk
a/KUu3L7kqaA1Ra12vDdTACDCECCTjr0LPqXSLnbhZnTiHGZjyoAo18lSljMQayaQ+h8KUQsLJA1
ZgvZZKaOEqJiMqVyC/EFVvlWY8F9Q293zaBj6DBy7zUSK2LQKbPTeIvRyV24Txs3dxpLbRWQSWxg
fh5cgqwGTaXrYJ3/heHK9fNrhWrkWjzFc998pWIUQ7Ux/kLVWFBlFlWWqX0q1fqZB6DQnNLlkiGh
vrP6hKVPN23VyLxmjzHL7WAoFEqox1Zfk7VR2bLXA4gHgYCkZItSNKktELtyTlu1rBe5l6id/dbr
DyOjDKrI0XlHISrzG7V7oDBjdYFEeWrE7eKtGjgguC6Go2cg3S9fqqpBO1xP3gUVqh/LDy/3klyZ
LMmeytlpnafczD/gcPiwPfCGPtZL1aVHqgmIJEOmRM7zSCtCCtn1vlVJa59hK/GLVqVyLggu4oUd
oQvi1p8MITuHl47sH4VsMEkTFMgPJfGVWz9uevVdwA92Yv7eOpKwJJT0rbDFsRQytn/lE7EFGxfa
suY349pfaDv/Qkl2sZlZa6ypuwAlqiVEjzrCt7mK/P9GjCAlHHJC01S6C61p6JPeHWIExxg+shwG
xGtW412tkCCQCq+rtVRKArzuJGwnNbnLUI+HI9jCuQpQDKmELZoY22lzjz3aLcF4hBGHApo6ObkP
x2C0KJpMNXnzi7qkCtuvets28DSGt7BibjCFSOBqfn3VAjmZ3jL6Y//zAI/XhuXzWqaYWiHMQu+c
BEjZj7B4HYPabFqgEO4P8n6vVjozDKd4B0OfJnXZQhQ4TkFt1cWd0eGG5PCkvebyhVWDgn3yZkq6
Ky2rDkncquq/1qLSAAMCr7cNjBr/4vaNUukt0Y2ZqUmaCcU6DXp/fho6EGvuzDAkum4pgtkOshyJ
iCwZKMOj9zlhyIRegdjOJOV4fcAGHsxeKqFiMekbxrz6mEa1OqhEz6G2sNbj1LeCwP1HAboF0IQA
58n15Abw6GJP6wAiRKIz/2RUcHoFIaVH1+PZv+f2CT5GRtZ7gPwP0pSWrhjTtA0smGtnXrGbBh3w
pRFtPvRYpzL4nkqLGls3uVWcaWIOWv0sapXRRFREhC60gIQJxqgwY5qy1T+Do9NYru5qmm3Ow8wo
5POhmIX3IIBmcydTju7F527BQPAf7kddJBGHj6fRuHv8KUdrsCLpB3T7gu+LoueBRRkTB/RMzJ/t
b4CHQgS489qoXzUIif/qpRIOJKqsIXkOKW3DpD5PmwF7Yx7Et/By591l5UFvGztnrbbMXucLD6lp
RKcfyxEqBRJTZPoxQpoj9HWxOtuMv0jVH/EzTVU47H3iUmbxRKtZPJOpRsZ0EtFo9ZgJKC015Tdo
mU5exQHBnVJFoD1qmyXGC+gskyX/SXMhZhYyGRW2R9YwPjdY7np2GoU1/7nJP8HnO8QbRqToofT7
W/eRwHlze2J51sfNpeU3rV27EBi5ubWzaudEvHndPkng4dVu5phcqW7jFbnCBoEYPvXRfz1SlIhv
Jh/aGy0Bw7fFrAPiTtPp2FfkyIH8sN8csFiGe/y84p3L9FvXlU2QwymGAFwURr+Gkr4/3ZkspQ87
Wp2QkrLBLGV+UPwlQNRAhPa1+gp3SfJiF+6SK8U7+JeYheJXYkakWNM/1gHuAOoQFw9OTIJ6uhDl
ta6/eEf00CHigkH6pjBVHGKXBDRJkC1ZnE46W7apdnRWIU7DqWiQotKORr3mcLfJw3KyIR+CGao9
eUWPU66qofFZnz8ouP0XJxl8YTTucpEgQH5+MCX6HWO0sLl4JV0xYg04fKc+Hi1kK2nmqDVU+bOB
HadTtm1j70So9is/8RwoyUvT2Ibzg6qdbHw1o+iNdu/5W4taczxwUPWtW9RjjntqXyTrd0xsDim0
WzfXseZJ3SkIDpv7TzNzaPH9aqdeEYmsBIasBEs0s7vHx4WU6M4DUWoq/1w7ZCKZ+WB8m5tDhDks
9yZHnZd2cojBRKzV0tIAnrIg2LHKFKDd6kTo2lTi55LOARKi/CXlpegYgB1jGNKUSaiiF+4xHVPb
RD9qUwpuLQczp3lrqD2SYmAVE39rHrnEIrnKAihUWKgDsBJ3mrH3RJfExp3GgY7UcZBCfE5qGzhn
GXPZe7TrgVuJ6Oo5Gu4yklWnIZ+CtJkDC+Dg4RVWQMKB8XSoDVhzcWgINZCrq+7mQcRxmY6/xnA4
UFL9U/8vJouCA3pnOY1BoSGI66NnzywPxh/YPXz/GdeMfqv4dz+tNii+iiYvgDx/YgSwfz4waaHt
visE2cRzoKkquRcUbQnRhSDyskeUNCwTdE93/W8P+z6nD0ogKPrn255uaY7HICPGTqovrdavG6sz
GBK1dsivAiCP8A65ijOWhXNf31cQK9P0VHHVtJHhoRwav/v/Qg9kriUL/BhQkuhM15+DIsyGb7Qf
X0VC7immSEC2ZKTKAALKncjWqy4pd6cc0tLcerbTIGBSD4B7V81xH+5gSwoizL5lOya0DzGF8R0G
Z0CjkNl9FsSzfDxspsMpN0azrq7Iz/Lu5FIhNicc9kzjL3opKyQAW+hgHPwO170sVIjZcQpdKDNW
V0UQPGGgrh6Vy3445AhcE3UK3MpbyrriuiMb5dL+SlNxiLAhC8yM0hYhZz9A7kRW4IT09mqUItCI
1u2O+NoJ/b1FKjX1gESvtPHzycxx7ZduKQD2/Lho+b6EtJV74uT5Auytns7qINAWDZcyx+D2uGE9
RVUgBaJL0l+Wm8d/2UUJpsDwa3sgR6jOoPzHQKJNzvd94caj9XVUOXwAcrC9t/rQ/h+2qYDifpCB
PA7MZ0EY+ge71+G/5sh8dI/aasmqNS0+joyb1IOKi2KA4frcUYDZaWnq6YaSjda0T5vW5T3B18bV
3UndW9UOEAELSQIqFv1Um+4aZEtTtKSqPlKqIaFY6oo8xWeXy5TGKQeTgd8LJdlvIJhr+Vi+WWdj
Soxtj/nEVFbwbqgGGAzN6HUvz3VDQTlgTKHz6G0wofHvVMAq5YC+CnrglCx3WOOzMPgDDBgBxqxm
j5kbq8inA+m6Y1HQ3reRE7Ie9i5yAfsnDUWyS2ixWzSNoRPVAmrpFWHHjofWt2yhZF4n0i8EbIYv
EcHfd+T/HQu8dKOs1DWp3M4BvVtaiNsQNGGZeeECHdD23lapgvT3xZ0kgT3+8JOHKKH7bgqBqa4E
CtYb5RyHT9PuVWkKMiKrledOeaBrFMq2NJXQ1IcZ3J/VPreQ3JMDKIOnmKvIRzqwmK8erowPRIDb
tUr83BgnUwW5+KBaFmdP8i3tBbIeg1tsiDwRz9HmpUzaAkLuH8DnDi2SYC8O5YY21nW6RGrRxajn
GfudIvZkdpcGdi+gr4MZNApYmBtGqnIQaukw+yHOlrGRhO1RSiUoFRpkNN7Ms7UEW6ot5DtMagaB
2W44j3NBKKMCadCYc+dDQ2AuG//qwWaZ3hpjqkoT6TvmedGe/El0QyiOeCz87Hboj1RVe9BxScd6
cZ6E89gpAuQ4rHa3qcsvafW8mHf9ilC2JatPh0kPYhQjFHrwrewuWfSdexfveni/gOJz6kPvy+sx
HfFydYwX/q6eGiNnOpmgzzK8eyovK46Xhj/cqrImYtj1gwjtiVW8viGrDZuDdLBbxjSEhWkVrPtD
FnpIfIOllqPEOmPjb8uUY5MaCJWOUAr2Kvu0xhYTHOmkejDnHQs5Do+cUgxTTD9GPHftObmMx2Hk
rO6xOXqsIRaEnujzX/JXNm7sQUFKMlATv8jah1e34mp+9IOoIsmUAURjbVkYM8Wi2kpihDvwGM0o
VxGZOnSMZQKCnfbiGM2SJBqCupQ7BUMeCqK1NGHbPjA8M+WTZ5OdQJdrHOADb9LfAn2J9+dnuTmh
PBFW63M3+E+RJGBa+5+NoKh2ea+ImnGC0tWt02S460HSJ1U2d1Wzgw8v7eWbiobpkTsflrUoxWoH
l/VQrZQONqqO7WrK79nrse0WPpbEsaTTYaHMj8xxtAsM+7qkkgRO6EyHScs8wZKp5LRR23hgqrSY
eSUDKSwfwfJDIYO8sO3y3SarhpZv95vimNjI09n7fUNqUJJXcSK4zUjv3jlTqbRjeY37AAYX8Xc1
dFpTpvR6eMf41Z+r2ZinsA2fv9tgHCJw4+DmQtc1vRkEzOIUSaE6xRDsQTAAdtR+hGaFuXrri9Sb
tFqIESS+9pdRX3a7kUQ7M3VXMnjGRPgEmuXKbeA93n/MhFR5PV52CDAj/a9bL6N/sUoycwzD+x7+
MXmx4GnKbqVh3aW+0FaaCT7e5ccwk1JO1CE9WHUG1ql3SCy41mS0wun3jZGyQG9QJhTqjui2i36P
iffrE0401n9EXb87HLG+FRD5lKvi2EsXl/Mycaef1D34Ve08VOcMMvJ2UfE++xCBfQnxj+/YUX84
nZ4PMJutQPPIZ3Sg2NWw5b2aq2+HeljfrlSlNokQhDuu1YaEN2Ky3LMSPj4HjitLls/BNVw80mAl
vVcIGmCuR2s+YhXYD5GDlrTHOOa9D5kMmbNqeCFOeNPheU9rwVrYzSE9AGMZbYrU2xdWj1BF9gNI
vQYLOZ2qkS3+aT7lBGStMMgNTeSdl2a1Ulc6RYn8S9hIet1rHKplE4AIr2Na5jA0lPuUlYhYZPtD
fTxgSBnPHWTZP6W9RA5XOjig4Kyfhr0qU8+Npm3ww4fwYyNEyULr4VeHAMVJj78HqF3o0avlREg/
NKKr81klEOTybUoiKyYpwiRpp5ZTAkwYdOmhJIRD9vHgOas6rK1WnvBDiL+1zA9OpwtXP04SxDEM
3ThQpx5bOhfy8epJn2IoQRwB7syvbAtrFO0wiGvNFu/pyHBo8T1wMkikOILvGG57eBVMD1o1DLeZ
BgHiPEJSSVY+oOHr2h2YLDQd5N3LkQHfI1VdI5NBFYfX6SPXMHssnIfhoBRr1GYtMFb6f2GlVkiP
qqUT4sR6hkvc5Vv6WOOf4ykZFc1zhfSkYXFxRGdV8Qm/2IlMouLgKAGm9sJvrEDsSeIwViX3qW/X
hDByDpVcPmSzOaJmXcYjQ/e0zUOxlVL9fNyHrijcHEmuYgrPXwqFewUzX+1X5LMsbhERMwJCvHPn
iAs4Bx9D+/fjZyFHi+W0n22bFOSoIRK2h7Bl90Y3nIKFsnbrSANIFpZRhVUOl+GJtHBi7aUmXndn
vmStpKS4+8SxgnANo3z9rS1md3qtOYEgKYyGNEDNVyPHZRS4fgxglEl43EecrmYtQ7WRyw8p5d2R
FG/ve07RrlLRpxhVRDX0hnIX3TXcPXYkVaAqAAuYIjZ0hFt5Znq8KgbhJ03MiBAGRpX0o/5B+k3b
5lqFUcnYR1cLdYwrr1hUG/t9AYn9Ucq2vxP3GQEgFBhYE2ltg1luh2SzVQDE1uaHhTxbpNebxLTV
Rx3FXnNsW2ACHZi3+fY9mHJvhXwYMK1dcz1OyFD8jWCVWJ2ELWU3cKcc+tZf0iTv5Kwiu1ZigvfY
8uKjVY3P9ionjoheUxLigdVBZa02XlQ2W5XKN2bC6HT7yGkvlz4tMXCzb0iKy4JHYcpdIcaMG81P
AjoZntGcsdivK/GD0xXn+1A/EnCnH3ZR6eeVBllRBzRkE51FUDQN+zWQNbj6gEJ79Dh/HWZOP3Wx
YudfxdHrmJGZmJHaQODZBsGmCqCthqoG8y44PsbvznyxW2+thzvgixHNa4e/tmvLIM43aoO1ZeYy
H+9YXcge30Cj7aGgfdQm7aacs7Is9E2NDId1HzhD1bdaHMz0W/OjScqLgGWtx6wwXxt2hHXjAuQ/
cHdTCcmaDC5rXQOQDz5/VHiqkqkbLYYDIKQjkFt44fzL20RFYjTboMTYGEx1nunS+QLyIr1RSd3y
YmfCkwR7Eh67uFglTZM8Qmby1ogApeOn/KlaBO7j9xr+IozFlVz1bS39GpdkJLxdtRXZbAK2sWxp
fBdnzG9xAzCsd/2t3PzaELP8FvTvZBjzBtSXNFR6xGq7nlkeAZMbXpkT4B+apaL92ogNZSr9aFTS
zIMEVwav4DWgMzXQix3gvsnN0zrxMKMIgvKBDyfZn8jKeMh6lxgCAy1VcrN41ABJ+6ae3w55LBr8
28hSgPTM5zB1VRXdmFAe0eEGR5+w91WVJNjLHmEEfsi6jrLWSqHBVM42lc/zIM4EQnTeDPwyDrFM
pwjdKnZIn7KUQovucHswRlAD4xgHFwq7FloDN8wSEgssj5irsnaTG1Np6AhveP4A/lVmM/FIDrZa
k3gq1w3gcg8Xpe6PSN+ZNv3/oloMGuN8BYknhdDNPdKkxZodzIEwsIfwOiSHsj7Fi4b2/wa0E7uC
VtElroAfvv1MUvGesXBFJ9qmT3PdAbhtGy2exEoqMspFhS43zjGTJW4xONRLv+N0Vf0vnK1aQEG6
VivRUtmtg9lCv2+f42xDeh6p6TZop1iNU8UDEj8+3PQUeIV6b9naepX83Esi8EZguLeAs/SGaiUt
txt0pO7cSSRSkTXj6s6vQ5CM5JrAf9u/oH0Bnoazbb6xhaIY1iLAI0gbLueJMQoXJCzyzI9qgtiE
4Ko79g5LfTUX+x2ljEvgswqy1BbUfKufhAjgUCAvXLQgFHiN8y5Rt+uSSBNORa4C9UL6etTEG9vR
1cahTJX9e3PnThq3Bt6EcoDIwTVCJZ2NQnm2UfO2LJBNw7q2uwxV56gRZ1mGzSaw8bhZzYbL8yon
PcJDv+d6UdQWIcBCnY8ni+EYZW/DEEjMp0MbEC9J1fsv88nHEkemlrIv3A9zlkjBxWV+GE1Pw+l6
RtL9B/NxIeo6MceLV0NavLnNHFKBu8H2yrU4TqthGhqf+wTKe1FcoMCW85xg3xO1H88EL9aYq/4T
0/QiDxllAZBacS7t8rGxbSDG5DoXDs3Mu4s9ZBQYLCrB4gWyMIP0UHyBYu5VDdSZVErfpX4S0Qfd
SoZNZuh+97Z46xXcO01k/aPoalIKVJRXTgzC2HtKY+wBFJJdGcgDw2Hx00Ddjqf+DCfiM1DvSCQW
ed7HMgFcttqF32JwttzxxESfPpvxdwXJlRfQ3o1zAhilQEv1s3tPk7K1pn8W3Fc4zXHUfPrLbQYo
kdkIzujbCWSiRRKIuS5WgGZj37XNIVdOjbjCseXNYcBhOtGQUH9I5Ahtzf3r8EDYkiG5lWv6x+mq
446Kslsh+96wZcYIsAUFixxdap6WkdNCfduwtqaBK3bSUdalczsjXxTanCcWNQKY58yOVeKBo7Ec
cG41iWp0aW3OWZ0SUOfn0rkuTJ+CUNjkfRdxdFuBTAY1vltepjkXijRNsZZiJl67CFuYkTwEAwGA
6gon/wv5e5VSq4Plu7zAns7BpcmFYaEhRG92j3C+0dFgKdF4U2fklasjhA5yOGo64BCA3nCwa4xE
8seiU1AdqN+FXb6FFUsRutBrZSsAgp/7N2lqJzGXsHDrN0dcJiH2x8Hmku6KLunwxgPg9wFV29H0
V5oBrSGaxmcrJt2MfgxVAxk4GqPZMkaEaCSXWgMRtM8EYHUUFnYBxweQTBHOmk5b4kp/NUkgZ3tV
Jeagvm6D4pWe3Vh3u1AN7xpQGDbDIwBZZC6lhCsxFIZEeX3mZIgX8HE2ajwPS7Lx8NZmBtHUnA1I
feygIDyA0/jA2NVZOo3WbzBq9z9QnV2TEmApT4OXiTnSXPrgzO4Y93aBz8YZdLZ174eTuVS6ovnD
jx4YgXrhvDPJcLbndAJtxMn0slkylz/AcLjJKb0rAlt7EIWpHeoo5ieAcznrtrq8iBIaqqymLkly
F73bKFzw7EJFoSI3lMbb4YOby3xeyPEAXcxdEb/uIjDxuxuEhBAEAlFYCn+wXsMmMuOThz+aonX2
/Wzhz+aCxd/p1RBBdAv64+OCzc02EmKlmalM2MUrzQuWO/Hp++FqMYBnQvYDwb/CuaxxgR7n6pDR
nEJ39USudlsDyYhpaZfigdiv1RIeOAv3rUmvW4PkUo5MhVzkkppWQds3ACaG/0iJUuH7r1ycYhU/
IAo3jnwqJ9Kofi2JKNhtsPhfWz3OocCpMnO3YpAozNnvrIl2tTVS3uZYqQlPjtGy5Qk6Twt5SG/M
kLauN60jGPLAt5iWg7Dq62B06/s0do9rD0VhFq4zncE+5TWqnUDf2kxZmCi/mXhCva7l3LWv6mMK
Oe4HDG3byxwzOt/J/LEyxJDi93u9SDNCvlO6HETIgONCQCkYQVBjnP2QW+ivFxm8snyv3rkfoEM+
+VLIj3oiz+89NpA4aJfrJexLqXL42JKZcbJlWe/da8HddlXT75K6Z9UxfID9utSHLc7RxSKixDis
ImvQCbVzj3NzzvlOikdGLVSid004nd3bepjh3pli2GpnSUh7jYj6g5Rew1IAczBT9yeHd6QFREfJ
6yQY/ov6amZsWK9VTnvSILRWgPITdmGG6r/Z/T7W8/G+92SfnIxPN0CiWczcWO2q39CgnWgOSGsi
Iohrr8yDyyfldJmcstA5FJAhaIDQxe4H6ce0Q81Ipz3yPtku+tSBC4SHN6/H9ox53lo0LJt8f5eP
6Oc8IpNHF1IlomFaQvdcTPokc0/5TTepRJQkLEmNev7WvZrxN866wO35Op5RR9CReAfwqRZYQ/k2
IW+HZMNy11k3OMaZoAjjY/rvSl6XZepGzB9uWgPf6aKSQDCMHE+NUhzJ4tbhypItSCej0TwsnFj9
oIJAB3VvfCXA8CQS5e7wj+laAF5w1h7eeaab849Pd5q0YayZLbdQs3B4nedIIAjBznjHFustJVBF
dIdfxagd2+FHuXZrCj3TIyaFXwr4gOCwOZxp6huobi0bEX+fVucjDzveCZ82H3oYRlM1FekpmuDE
xglW6q0FWJcCw+MfFLX5KIGptw7LoB1mkCrViq+uHRATAV4ytCbb26LILMP4xjiqgREh6L0xN6M3
1ZHCG+Q3ewHi4Q4ASqBokeKVPx4jPGqPfEi5W4O6nYQhYE3sq5NtsFCA5no/yuIPV9trMaSQvIGn
XaIk1WzrmcDCvwd4lKNIj3BHq9vmu7YLDlwXvKZ8Zs3idw5hkga70irMS4Y5U8rsqIDUSD1bImDz
5JCmmSrMPbU/kEpWnG2jQ5+zkfTGF5EyfMaq3tuSYaH8DsL16Q8QV7v0LXnJkoXAN7ZLUbeUH6mz
0/I04N8zUgu0L/6Z7kA4/Jbk1sUryj6jZnEYBkXDXbrD41mpxpbziSbOPft4Qpr0kWsnCNYxIgoi
21lsU+u6GUTA1TvdkKabJdkU4Hi9dXkctRHYLP2UVF7bmGsWjllJPQsQGr1oMELpm+THJ0jAjlM4
ohfnhOqZNcrcKffMR8eN6Pdkm6ne2tCm3jBan13fxvKufhstxBTfCpYm/YEZj0ph8X5IDbk3Nyrj
3CRyQBbALFANsvgywCDuFhGidpphXzhle+xjK6I0sUtuj3QEejEtBnyMAdZiSodh3ryJX2vC3zpd
WZjvx2cBzT2jCY3xrsMN/QpNMId6WJmA2remhIAruY02QiHwCj/bID2q6NTrHl8su+rMoY8snR0+
MCCPPt1Fk58jrMgIKM5rTOQO0JRaPC4NXF2CPoNNOShOH2v+rHIiWyaNY5As40MmJ5ZrhFYgUVJo
eS40Hwhp4PbwuhQOS2L28Y9TGZx6lpQPcin2ORVlr1YUEd50O4UoIPwemJChRSTO9NKGrbyGqCKa
KkoyPFDhzA+RxW5IxbtDbXJkvnYCy/q6x/8K5TWLoXj6eyB19aGLqPGKG6VZjs/6qtV0NYM5kjZt
ZddZlgzBFObWSiXphO60EyPxvvJzN4P46IymN5c3IvPQpBrcxYj3SbwSzpSx74jSiR/MNTXphfoA
/cG889ZknP1g+uxnttCaTwXK33btavUkcq5kfuHt8mWph+HsqbIl4xArRBncvFJDVe282qfuUW3Z
OA5jyTGCMVBqPoG1J/X9xAUz8Tq54cXH3bb+QlEcPWxdLy/JNJ/VEeJnmvsqCHpgZ9uKNIHGj4+X
m09SBi2smXiTOgodI0LkckpQCUbijuxxPE0BbXB03lu75yT+OjLTPFtRKveRfcZ3XA/TQVxatNsU
wrN0AJV2hDKesPE72X52Nux5KgEIPnGtI4maS2iEDpg/Kdc1xvRLYK1/4AuFJxktcXWKFXearTDd
I7stX48tbaFmWHRpMrAC3E7br4Nt4hFMi0jePbmbLKCOLYb83Q5Ueh0MeFE0G9TN8sjUyjZhq32n
ZAl65ZS+sMnAIb0AZZmvMTA9wfJ0k+79XySuzV8Pk9yYvkppdzhyQUdS+uNyA5LoG/GDR7wssk2d
dGxifHYeR59FFQUtG2qSjPGnC3gdY4vUZKqphMK84TZgbbgrs0VOOb6RJpz0hX+7EAVeULmGEMoP
DgKZicboxG+fwQsPiRUnMI6phcDl0/9ld3z6rBKWe/8292njWIhTxSMCZCwaSVATWZMt+QTDc73u
PZmkoR1R/cR3g3fJBT8pyLcAhmDvJocFOAWISMegM24z4LNbLucEoFO02oUHjkqS1pWXKWm/NMyn
WRBhZc10T3pL/y+GHNYNHPFhKHjyHHWFmofrep0lM5PdMFRZqFDlLcv08mxaoKWWzhftj2IQio61
80RpD/yBNg7jDXMt9r7c2chyWW98e1n8K5azLcAr6uZAf7UUSdeSoNJzw73RLSFSN3J7kdVUszaG
5uX3e+XHPPw70pbwOKaNgTaFCOcbIgBxsAPP0uSQcvQKtGHhjIZt18MrzkRmYczuuFufcwYBjIVK
5KN+J8HrBMqfxHjWu9K9vfHhWkWSHV1MHfBP4WUmy0kDHGvY5rphcnoW9yOZIgix+tk3qzoBJcdK
ZtPRU3ku7B4CEWzl/pKjjMEO6lYQbGKt14ffFUdATOnTt00iKwNt2X4lNaCANsaivP2KCSWAUc5l
ncQ0Ut+J2k4QR0PFyKLOgYO78bpIjBzn85R9T0n9zvGtAD5Mki/lZXqlJBkg9n//H4E+eSYG3L9x
VLXwVfn5rPm2mYlDvIvGTsRVy/KRhMmGMC7bQ3KQ5t9OajEoml6w3x4UVZTvFP2F5+sH/MDxYO/X
9NV2RDFhtC+plEe17t6pTR3aW7X3/ab9X7sT11oztMVjU3tkqdKMzgDbNPFdbSbzUGT1VZ+vnp49
5rCsiy4g8YsdMKLhAqm9p2C6HuLOAJc+Ab9/PYUjxleJCOooaznZNxfZ6zJHvQ38W2lAp95v8icv
QIWDa9lGu667Fh4W/RBGhoYXurEElKQ9nUdQPNlYy7IQOtOr2Mj9PI3dt+ZSzhScKDkX/VuEEPyX
UTWtClm+A8BP2+SjGl2bWwpo2BFMOY3gx40qo1MJ+U6xo/JZp1RcUIZARV/Mt/vjOReviif6jaHE
mvlkBVXt4egOP1RDSqO/rOlVoxpBz4mkx7w8lr05nhcZZIPA/ZDSQq/xHeJ+hBAiQ9EC2eDhKfyW
RVuqBMdrKg4fU+xjTG6wVY7Kb4HB0/abx/yY7CA0NdPyuCZNN78Ji+DqfMdx5+ybycQ5q7YJ42Pd
H7DONV74vJnPllgvUtX/1WNJ1nCWVZwIRwGY0dDW6ZM1zwSqKl5ehPKkpgUTq7iLExBDrseYs+K2
+sAgfXvfbqMNmWWcFNJXDtlZYlHyW8unkm61NK9YCH1yX7zpiTV79AFLk354RRl5/9P594ixRrxJ
cL0Ov/LLvCQZjNQ+hI/KRZpB3barjKy8WyEDebP1cu+haTM4OxBHAtOpRl1lLUYjqSPZd3Sptd+9
0zKIiJHkvQesTsEOUFPK+3+a1axg4BkmotYgmu8AjFqsq1UYQOo1IdAbZ0kPd8GtqqyQLgjjz7eB
C58mlI0zxtLQIksEIqP+Lzcq2UCCu8PWCgiLQHd3onzJPrxBrG2dcfPEvkTxUWbLfKcWnq9/19m9
0qqId0ZsdEcEMlJGxDnwyBZN5UiHkh4PQtVm/6urkC/5jPInZE0iPrI5rJ/Wwo3mDxSpZiZsqtUs
P1kfPSbBIziypbRxH4AMzkdp4c4i9TnQdddizews+8QA1d+ILhQOIXFT4g0XutNcwdlLBLujxnvT
emvfnGq3/hj7S47ke5AePepDEvKLxRND6CNAM7LYrDEqkZ9p08+LmVdmsbUhyGa9Ozvlkz+PlwF3
fLLFxMs/VbD+Obx80RcSfBACtKSDzxqMoAlhWqyY3e3uS9t0vf/DXBRtpcp8Pn9bzSEeQLUumhp3
vSgbi4/QZJf0hfpaIGKTfw2Fx6s579ospD3O/N1iuU7wgKi7SCNFgvW7C73136Vbo58gkAdngYku
qvbWvXLkyMbC7SeaoYm4iDZDWEwtW0ivoKVRYwSec2lDb5h5ad1Z6GvJvVAvZjIO2gNRVEMcPtpg
5O3ZunGzUl1Rz7EkxEuJODR+Ojm8EVnKuGFqcaIY01qqhwW4WqYjFq28l5GkyVr4HiEtYxAfQAMa
Z/SRkW8p0iAytVfKBDMMVOfwSKLeOxHTwgjsw7iIy+r3M0vrl7iZ8f5zz/Q1DYxKXc8NGdL75Go0
a0IYyutJMwvUJhN7aGKUkW2gssR4nbnPlk6zCzkZQH78pRrwNhjY20SqaMsdhbFV22ahfiJdhVsN
d0I/tCpK2AasmABK86sjDeqo96RvKWLMavcBgSUHZ7wngOaNk47MHkDAfdqA7B3P/UYgJAKx00ld
lck4K7/WXSDTjJQwQgjvWKRZL8j6Y3V8SSJ/lCMBN9By1TRhMXtYuCn70hc5aIeIYRM+7O/oo8QF
loVXoPvVxBFo3bgA+pi5LH2E4AFI0tmzYkmknIrtL2+arvVyMNJVf3OFYsM8+VT9DYY9GzE4lxMV
GOrSnAbF+qX/1387eJCEkXJSKTOq62KqTggR/LCd3Dugj99fmBlH4YwD9D14nSdQlk+4fKRirsCO
anBkmY0xXDQed8wQ9TYvk1to7Gcc6VXxDvNS4zDwxTjnL3JpAVe23+OiMV13JS3Kue/rhIVYWQvN
vtMe7WuIPr1fWnCIF/du6XvQeFD9wosLU2+3cNwYe3kiGp1I319O8oAZuFZwRLSez651OCXmYgXR
JxmvYsReoIfaYK/nWjonGo5A+fUz5kHLhm4yvLFY2S9UzD9zTa41ZiQs+PVfkPL4XC8HGVF5IvcJ
SUV026ArbLGE/gnIydhRWtLT5bwn3RWRQmQZ49uDOFdflqUtsl1oAed2J0Tmpe4FVYcxvmd8M/cI
8ENMesluFJWCtwot1TED0AWEr/Y/Nra/lP/bz1BoVOPL6xkGHTdECYJ9Rfzc5USQ2R1nXFjGvQlP
HARCeIRfHqiMDABLLVwOSMsZhAnDP9Myicjoz0SCk9cQ5FKRs/8mdXdr2aDgv9aqbOeYSSlx6O0F
R2rzvtEFAcCwLjTjFXdUiRz6n0baNTCQs+b9bXMn+xhavZ9hDLdSQ5nJIHzMfWF1sfAemizXquYs
QavUe9z1o++8UDQ5gt0hlfrmPK2u6msXs3Rwg0yJczQh4Wa8j5hWxv7E1Hp4JRJkG3WmS3P7nEP3
sfigrwBkQ8jq3nLvsPKUqYfDnecYR98u9jnyUcofIoCTv92DutIZEysAl2Wehq/kkudiEvsBJ4RR
xSdQiNd31zA+aLcQXTkAYheFtjOENwMRDQuwvgYefziMZdbTUraiWoGajPVRdHhU6NCje1XtXslO
Z91NbZJ1y44qZd756t3mfZp/pVPJlgyAwg9TLPyShq/Q5/HGhBZ6pxL6JX/n33hbweZj9NdG9w8l
ZH1b39IaxU9NyTf9RarPP5vIfVkXMBEj7ugg4+TcEriK6Yq811o708js3H23PckOpSwglVURNnTi
zfV22nP7kzbuovSrz/EpJ0PUjDB7wnY/38lDAF7Yg4w/Axusq77cQDscnTVfzgkCumK53YOI74ZM
rIpHVmpSYi+PzCUwVuk9H4X6M19z/Qv4lNF3bTS+eJL7tBXS4Z4R/LTgt77k31tE597rq2IRXWjA
Zxgc2SLWw54Y5btgChdFm/OWU89rqZwC/O7pCxiG/Fzjbl76fRI5GhtqZAsxOtBbV2IamURbnmkw
ZaLK3RKe2Xg+TNhm9YklxF4X61c/cMXMYwlcO3e7QzpziVt8ZxPtSiWK6yWmWmZbiom2YAhxFhVj
hwi+Al+tSSE6Cax2ZsUmzEi2013awocLrOk6wZljj/u0gRlYWLJWXj7y597mHpFYnMG4g/CrGD60
eal0wP+2vPc0FkD6J+cZ4bhb+QZh8MxB8SM2iaFZu6fmxYwa6Qzc8uf9uMGGrCYJSPk5NMFKl4HW
Jmvhmi2F2X+pv1JrCWpv3hDB2yE6XQuVjV30uBJEpujsp+gGoZxPFlXOUPXS0HlvRzBkZ2WwebiU
OpeYtmhnEHQiSYPpU6EF1FhxbyH9YZQ9fdH/8MhdwxXjqzTKJdldspl58ExgBFLN+sDAYw3WsgdS
GUosjhxyOyNBOBIDIOA1Ij6afAccTsl39vrUHWZ0qW7CmqxlmhQYs/X1LK16Yk1+EamGQsVzkFe3
UME7lOWi8KQtVApBXVvZfOvAqBTzMGhlUkafxZZqOw/z4UYgu5Ehv/CQx0/72GGN7vhuYi1LPpse
AKpXfJc0T/IN9Kiw+blWSTe8WdFPoKk5XFrJ6LQusvzg4VyqgbBBBgWsXFaBQyMPmPLvXDI1d+KK
M658tMA3ESj3qCabhmcqiNfZlaIuv1gUXUb65LSLIGNDLLwLfFlKKOpQpMzIA8S77G7q+sbs/Ad+
M9z/Mn/lDyQF51msgeMF1H/sdMU/V29M2JR0LRndgYU1fITdfeD8l4Fx8cfHhjcWtLKcy7JwOiz+
SWbXX5ye4POEA9l72FOpWQktBdugOZaOaOC6r5R6DBGI0uCXZeQZfvMpOdBiaFwsuMVhfdYBhYvS
HDjY8NSORCx2z8mCqIHFBZYOzIURbSETs8u+CEBFdRY4strirvwUkwX1pW5mUCohjIL52lm0dDgr
FrcYih9C1xtmqsFRU5HSG8i88XQixktcU1AsyuHOWocP6S/20GW58w6NEpil5jokIWYjRVNC6E1b
2wuifQwPHUOzh4OOdu4PyrjqGBhpDRV59mBsBwNA8Uydj4u0pEwSoJvdxFBKsD4+CviQVEzlfpBQ
GUnom0CBgDXAmlro8WAPuozwDNH43+iG9nUQaQibzmc6dMNnN033C29n0TxNI8wsoAXw8F5uHbp+
wOAv2lwndder9khh4RdODBIl3ruVSq7TWXhhnT7pB0recRO4acddoliszpo2BojtsZYuPOVyeoi9
bsqXGGgamYygaYGwWdmcA7/zgSP6E/Cf/+XhGFa6gFQXft/CuDghaaXei4PQf/t4oO/+haIhA9Ml
a79dHRir3zQZ3DtSll6CMZFcDgfTWV6mT0qlUHYHd7fSE5roLcINKH27hHTjpwGEzr63WTgqwbKi
99dj0U25dXAPenuKWXdSSEv284FQ4bA9OVtnW/ydn1yBmpkloV1HKqtk9GfvsgAhxVpMwbgmQwz/
kHefaa46jTcjrjnTg28+h722rLdmfHhfKs3MtBaMSXXpemY/6jBeh+oxoN2i2ku+hEyor4SfixP6
NsV3O39NjuYnulBX15WqAm8FIxua7YIdaQRycJPGqRJ5v1hT2JK2JmyBIOXrWVDGOVmAiaK6Vuvs
9MA8rpGYKKMNV3LLvsFrl1kf8MlW4OELfv87nBlvgABkMYobkwfPfY7UqRateKnpfiHT+ftXcicX
jTM2MnioBb1JhwmLYZUyoFOs2UDlK4OegErOF4BZwRy8R13IQ3EsIOizxcejR0aql0bkdbfdjOdD
8yNXda0mI4kV+Lx8D0+WDRllL8W6AsOdlSUm4vp7h8Hd007u8CClUHVMrhh7HdUEO8V12Q3IY0MO
GLhosowfR6Z26B181RQmTWRALuSEo/LtQVMV1fXEf5FyNM//HywOReMD+ADDUW0T9/IMTLC8rDFM
D/tYx217xdsUFXV29bUcTggTfcGkaFlsP5rRn2XtTO7L4NeHQ1n38UBmUEBHfiupyRkLbMJoqopV
573Fwjt/7iE93IS5oxtgXrGhPE/mZuj5DrYuVx5nOoNJknRbThiU6QVQvArwAxPjg5P91IFD4PDv
T6M5WqlBIkcOD11Ua9801Gi77kJB2Bg9wP+ZuyUjdL65nUvUObO6Aq9p+kOszw5cArpYvRS7NneR
t0xOIeOgdpnlvoY71tv4kSUyd/REvHPLrtQDYOBgEugVnnYozGJxdUJWV7omJtqxn7NXKLg9UtFC
DaTJl4G0hPjNn5wkmHe7ZY/cGASkigDbod8KaPsSLJM2ZBYHyMFPjMMTlYwrJAuml3LuzTnSqH3U
kFvmWRgCiSlAwKd7binNDciI1b0vCu+kLX1OXD1vuCNCom4cJQrmBbc4QY80n7Rs/V2LaYKfsIJk
FiYe6qNMFGoxNy210UtKC6APH6f1SXvk43Z0iqb1eJvZRZOzI8R4axYTWD/CQ8QIBFUXRgWXjcdQ
c6lDNxEhOZxVAn92MrN/XlZ76d5Gxiuchs+s/cTgRRM2Brz3RSYdhSjThTY3uHqP7Eoe+e5FynSs
kHSToPrzFoqUjGDBU+FoAH30z/Vab+C+d+eFbN2vYcGBIXkFg1zq/YXfbncxSIFN5S3H4ijSDWAY
OTgKMyM8cdbZ9YX1CQhsa+zqTHcINiepy2PSDRgtZTTcQI2CJ9+aNdcz3OQNoLRlci3D35f27O9g
7LFSrO15c38/Hb9TwUu3DSZAumXfxcPsTYPbuMETJmz89wKE7bS45guGnba9BNfmHd6ZYM1WBTKm
OODb65569x80DUHXR8YdPN1O+a3TYYH2ZfAkf1WkEpSFF2AH33pet2gSCEjjsItbc9AJiahHDXab
ybJ2e/hL+FnwQCno4LoUK/VlL25yF/TrIfEtfv+1zH93zCzLu2Bb/Ss6JhykDtsC/Q3DK1Baxv9p
BW+1QJvsaU3dBN4yhdUmWtHucNbuA5JBIvPra9AJqAriIDWbGrIErGp3cQtKdPzD4FyJ+VzE0YIJ
fbOzQAecQLx+TZ83YXCawMqbHIIc783qL9/uyYrKws0dVCSxkwDE2DrWDwX+Be6ZxDuKcLaklOkb
W4OA1178aWkX4f3YGgEshYkwJLqrjSwwkKXi4bVcLJQtsevHTQaqwYLe2cUczVREnuYCh3KxmuAE
0NThZIpeslmlZrMhhZy4Y3UzBhH+27z6WdNgOvtorbTkgxISYV3cA2nh91BuY+XlbuS35Q+yLbxs
lSwPZmc5yJa6tKJr9uyWliej6WgDEGyEWlmegHGHhW4cve1/EVt2sGem2sJgYhH3Q6nCT0Ocqa7r
klVzb4AJd6HeKJ5JKhn0twismR/myPxGuMSqX6ZKhOBvo29ShNwz2fdjrnLHBOP9ij1E4rT9lnG7
VsAiKCX378hsZ9ceCgb47UANZ32znrfLvdQkrndzPsupbcbVkw+l68NO8CHdE9y8romewWKnMovR
xdyumxGDa47E7O1SajxNnt6giKR7iFSC02Sabhm7UZExG4s0Fp16iE7z2t9mOX65duyp3Ku+90NE
W2KXOPHOl4liqvIIFXAdE++6yXwQv8HI7Z53j+kHQVHMUkXR74roGYUJuWidRWisw0ShvOLep4AG
VlXyvHLiji7ulw9eNyXPPLRUShz/PPtCYob9hO3f5+PL/1vYZj11+ck9xN/V4qQC8ERQ/PU8doac
n2BJEdi7UoNWHJitGBYyE7PpQrQ8h7xDxaNFwssKp1UhBCRQQ5q69f+wcYg+pNPOhjUOF9Blx6eQ
WlHGKT+XKVUbyxrv4xSjPsDMavrn2kXPtGfUQ/jUlg6gvIqe8vL4CADqSFHlqmRnGRJ7t22tiA7/
e3XeRR+7BNgYKL9anV+nt2DMjDFf1NwzM0BLXJ2Egw4X2LppapKBCDdE4kPFPwAvMNsYfS2YE0B/
Bme+YUskS3o+VKO6BfPq1cpOz+mochjsVPA5dgwNaEKO9jsRJ/Noz/zMNST/3IwjdsUKA6dS1Ko/
N6j/2WikJF7t78k56Orzeq1V4wPQbCI8p8gSFRCwlrdPiF97r8e+vMqjTa6ZaPxNSmnnX6iPCwld
lJpZMqWnaHBsEGxW7QgzzMpIrY3imbYXlJijEjUPSSQXmU72fbf/ucD0mG/KhW90wDZdUeHosfry
F0FbDXWFUqi+7x3lIYhxoxCwu0V5cMdRl7rQRqcgWSjDDf2yhu18p9ZMpzlo+ZRhi3Kmf1xBf1/D
KUVgpJrIrX1dDIos0UE2//EiklTSeXKBPmu73dpkj9r9phpJG05QFo+4LzOlFCwiT4BmgBQpuk//
swxqQzFYh8y0d/kIP3b7USRnLX+0DQQkew/FFbv9U6Tbd1R14MbBSCj6ppwmE+u57gL5C+6aznqm
Giv/nBVdttjyYioEdhxkcYY9tuIu3HlTwurmIe8AMi3t/JxXV7UUER9Trzx4U2+v3I1r6fFhQVG+
83NUtme6pqDa6QLay+W2JHRBp7D4Bbg1i5cOrQmtgBm/3BWKXDkh5RXt1b1jaRHRs4X3C8UjBXxg
Nuz5ktwQaF7Gszr4M/9KVALoEOpCu3+rq+2yxLAZ9Ew/mWt+10kv9TpnpBphYo0xMTbugf9nSC/S
mCyen2ikn3f+XiixW3O5nQN18g4PIRZhb+EjfEkKbXDeEYrq8MUK6dCOQDog7mbWgWk4fNSBRvaQ
SSNtIumHv1b+BHZoXts9Azo1p9iV3jogvr+XHWoM9+V4jnOXEamYWrqSMxmdpTPmKUlqjer6p1ug
t85BraHJG5sYrmnKzQRBZEc4d2jh13hXRmLkkcXOCzd8pjdhoaAIeUcEU3EsxkOFsSihDdLonuH+
SGugKZxWLcF525TyctUBmuTOwWRa99vOg543FChag3OjC5+Q8zosXNfzWgh5QRB07NYWSsemsqWz
aBC3oKajab+lbuargL06JvNCNlQMBylN5y6jDQnDP8zwV9B9Laa+v6OerN8vjHq4zgxMnCKjfX7S
7fuhAT6zEFfdp1tS43zQsMGiKpJULnC28XEapRxub5hx91HOAGV0/fOSpF9Ogg20dccP+9G2fiwc
L77Fq4rzTefTjUsDUVsUAY/uxLWmUhdYfmpb8OVYTEPAw/QUGYRmTr47bhdUNSOkiWvMPTUlzQbI
u+1M8q0+JzYxGsIoihrALJ2R9f+EclSu3VsBNOllfvur8HWQTcQJqMTl1n5P+mRZ3/tq2F0Ref7D
QRq3MRi8lmPow2/ndzZeWdCsH//pV9r70A0FGDGLJR3sjXGMtGZ909Vrz1+isp5MmZR1UKTx8Jrs
OHFbzl3y7ZqupyLf7ou1MG+NCsj20e3lyc3O3wQXs38XzOlFZ3ywgztZQ61KFHzQ7OsHKQx3Ru7F
GoN5YsHyGhuknuVmxFlH/uvPuz6Igom9uamSXt54jOyBiN15AekE+j6pCp5xacYdx5RSCxKg8/rJ
VBLwwuWYX3Z5D23asYHTmOQOOtiNUnEjCQqTfAZpRgGagPR60qhAdNnvpwn8/gAe80r6uc+cKjWO
cMmG9GGaWZR7IMym5wczSayJkyjqLQdQiJVnN35AT8+UNEGH2SJ3blT6rFcpT+gD5liEiKiQAsEa
AKl5XQq6h2S2XqnBN4m8vyvKZeJamYTZEnXah9B+jA9a1pcZQkyfJmkPvPmyHivQKSbbJNT4uJsP
jckcrPt0Pwki1TZBOPbvMyfLuekHqfpctt0gM3tO0/UdnjGF2zRyKg3w+XVZ5GOb2ecuVVhD+cKK
qctN6E7/AD9SJbWYGmOseD3BilEni/jInsHnfYJYEmDHVPouAgH7/ET+AWoHb5/nlzbIte7unFWs
F1XqgBlzHDETazP5cBT6nwDu9P5LKzBGKegoe4SLT8PYam7BTFtNna1EAlsKr00CQfhvGtyFoIC5
kskzKuVyhWzITTVyEKUie0+ibD3rZhmawP1hQeiA2ty3EPrv5Ja/HII8SosWwppup97ZpNRAShgR
PGlkX4etOT40jLu7zerRLRGF6/8/BiUQanzVuky163RNJr+7J6jr+MZ0DC9ebSnaJFa7Ik4egzhf
q0UDaQktRUyUr6+U7hEv/k3WHRO8qGqk7lUA5jMfom23Sb44pO5f1FaCh3U3fLr3V/XT6WlElpVg
hZWi3oR/qLIx0MGnb03Kbb4IpshWu9+hkL6w5M/9MxUXJ+c7WCGzeDgRpTKN+1GFdvbWGRqvvEJN
V4nyCJSGQ45H5yCKsHTv1Bx+4lVlxvwayY23z9C/2FAc942eVWQVvvpPZJG2o9HipRq1ifNr9kDa
d+0EIERW2Y8a76N49JQqrRnCB+GxxGtD1S69YRYy1qagGhk7trzVznQA5oKPllYJftTJzFFUcPyI
O/44KSSCSPUqLA+bQS+deUC25QSUqGxAg/L+jPdFeEGIG/0F9NcFVsf9K3ZpOEZk7lKfMYOkcwt1
AKDMqOJ72u878SAJgQMECfmBWFMibZ+JpqwIsmFrGJHSffQZ53IyN5H4wovYqPtEFGfqfdfONIhg
fEC8+o1fzxUVhir3Vb77gCowEiohhqD9OBQh1Z/97gUVHQVeNa2iI4v3+sFHzJlCpAoSPox/qFNU
YbSPYCezTVamxUyL97FINEFFI0xUwUexhcylw7Eba0GcTP7sHtGpFhC9qYK7ePa0DaidVLLgX2/+
K/29inNPuyq9IlufQU0jGb1tg1tQIdKXTmLmAl67gSW6EU/8yX0a8ivS+aeTYqziZtch9aklRrYm
T5B8+FykdHd+vmD9pXFemXt/DYhe77OyUiLncZK6MubeQAFHZoqmCsj7DfMqs+XbMDs0QUHQkoZZ
10OrlYH0xicxL5ijp7593Ijlvidf8mRfoWVCB09yDYtPjo47MWN9SCIZkUc5NBIVTo7ABhnsj8v+
LvMZ/8qvc2f5Cd4uhX75zPs/fT5ytm6Pg5bLRo04XX/bDibbkuJW6Q6TJyyDkoEPGINw2Wx0hrQ/
L0PYXv1eE8mESWBdxw2ZIQNR+WH3HpjcgjvwFsOptFVSMLcdFf6lednhwNwTQOlHDDtO4UFl/Ydu
zApMmcDIWSPU1K9MfxtkZjZfcCbKMto558Rqqdjly++6OPUgOaVlMYO5vnQ3BynmhrFfgR+AtgQo
vys7jTuqDhFifw0cUR46Sz66EYg3yCuyWNdyOyEOGjDY9oEPgBtC7YMiCYqcZAeY1Yu+8IrqZvd3
vdYOWVVo84pL4mwYskFVHIPlCnoXYr1ZrWQXeJkViO8dwUrnWOW3YPrB+6KIkM9sg+u3oGGOFg0U
lc8/e8k86O4LwZo47wXhXKTXcVgJrJaUAcpMwQqg4QywTnf/DB21BfKlFew2LtE2x2aWmpQn/Hzj
Vqck8pVhr/Y9NQox9Ln+DyyiatilunintHOu9P7+3jWeGbnw3Z6K5Uu1hbKmHivGDiwN5ueaL9qA
W24/pUCcxJCPEJFMyHfDNsGWOntGEt91Hyw7NMeJlz6oa8X2Oqn/oM6IyVjJV9ayRGsC/ZloDPVs
cU2kMYQtERBGfVj4cX1TGOYJdgPYUxOD/XQppMUVtoW92UIZ3b8CD1qKDsxdujNka+sdz/Q8YiwG
ZwoNp8K9hVSvIqP7sFW7VP+l6ZFhuMP7V6gSRBkcsCsgzLcMcpD0D3fTola+ChWQD3oxKQBYlFFj
R4xjPSh/8fh7vluS6yTqWjBijZu1F3bQRkbZYVLEiu4dx50m3eS+6aVNjX7X0cF20YND7oNZRinP
UO9VdlrDBbVGab2EuaP99XhcOl6KIhor8/Vp8WK9zJnqF9sMhCaoMhrGTs97rOGIOVE2FeeveViI
110A2/oVWwnpZ+235EULSsu370q1pbQLZBpKTuqJUawWf6jw5wbTgn/B+xtvi21uVfu+cOrMoQWH
3IEXmLS2THo0PihF8C26mKcVsbMsd1meBIo0UsEdASidlccZdnJHmwiVOFfH2srtsZX6YkuODxsz
6yhr4r5l4EskM/ZuX78Da+iRdXoSKhTOcju5F8trtHDVx6LMeouV4Mo0RcHtoTDYCdfQSai3p1bg
uRVMF23MX+stt0gBV2VGMx6qO9eJ/6Ol1yxrv0y8sHeYmOUT7wGBHyyRQc7vxHGHRWaLMsI6LKhh
IXCM4sOD1BlQKukMpgrHgZjQ93f7NvrVtxdhw14qTHuvwW6cagAYcqGbRVRGFruGzUno+VtWBl4k
dySr0Ec8RcQ0epJJX/2ApyXyKLxnYHhlbQ6ZbbfdBvxkks7RNBAJgOOOmZNIfvYDW0lGAigZCnC+
wPnRJLAvV59XlctE+jhFqkwNV7fqJpeXCMQhteTq/a2V6N/eAxus3mx7TGdGc7KdT0AqQ7edYoeG
S5+LX9kU0RhYjUlcFCm0KXcBZ2zeiWsRSAcizuDGCr6xVx3LB8/CSEMem7A8fZyCPbAa/+ANuSw6
shcdvpqQ7RBXpH8FZyYMsK9Nz7k3DE48+UmrENfqjmhhU0cvt/im2I2tjJ/j2J/LJyZWzdpu/+Mz
iFU6nrPQhcFAjyzdwOiUAw39KarjmMvmzRd3HNSgaY3kWbBOXa8/5/VDGQc1XoweY6RDFe8k05t3
Zt029724Eann/0WYZjsc0c/VGA79qYnJrczQIlMRi0nHv3d5sBH48QGcB8Ta3fyNToG7HvEYAHxL
B9o2kJxYUdtE0ymmjJ5BnjTem25GLBQyE5Xf8pGT7fJxjxSQms9OULrBo9+aZIPtYpVU9QFXF0/K
UD4VV+9mWZkb0SyTF3/xb7DY36mTVJrVdHwBblrgh3F6Xh7FrtNrQrtzBhKaU4jwkVEzmodNgCsz
YUbuqB/VVQwUCBtNa7JwbeuEXXJKMS4lckDIUFfiGpZ82H+C/XgpWW4As/s1SM9VGqCdPafFHHLx
ogFPUzEfDmnJQwH9CT1junyj/Ag/ZNyFkvRgJj0s5jKrngRX5KP4vjSxCiEg/hwJXhRzA462+SBX
MDzfDjqdHHwXNMM/NSdHZRKAToXStgoJ0ZtBIblLML+z8lzyGs0BDZHOC+ZcndyybNntzpyHDQ4P
i8FYLiFQ/wvfBHdwdk2WGHumVV+gS0s5FpMCS72XcGL75bymwFwEgrXBwvJH41RfDgQcrRlLs4e9
kki3fo01aplHp2QQfFSiRgi4GixlvI0bz9g/kCa6QOTEXL5WAlvCkzdXF1eP9EjBUjXb+M3T7umj
sq1binXgZnTVFvwDw3YyRC27Njd9r8qkujeL2hy6clGOjxgUsCRsVZBK9UKUWpxfza3a+fOpcdVy
kDDdbZ4ej6lgROfBip29f03Rkl0tsz1dKMjr24vGEykkAEJDxfQ0KBOboixa2+fGetsMXtrH/AtF
x/4+aL1Z3bpAMW5jBbo54g9HKKeBQFOWK7AsiH18ZiulggTAURGiutaiq3sfadrEQHIrQ/EfZbmi
OOaoyjIRUIRl6kqKQoQF9fU2o7tfMokMBvEhZp2VrLc6SMFTOtX7G31S20eYdVdFtj7cYyTP79By
OQwlvLDzjy8XPawcWLUfUsEtF4MV/WI2J2IsTClvwh18lZeJwiNMm5BinmNtqmp8cVpcFDLh7exC
97xHMtBaswjMqUH5EyCpcbRJiVE1JwjJ8J1ek76ddUOhPntc7khb+zZjNi0BOgt41p3ryYjTNuPQ
N2uvfTrCx9cZxcaiP/peySKDzJLUsbRPqoQ1MZp/0FaXfZ9QMPH0MdMnB/8LO6MKAjj6piDhvAIt
5YWWkMfIqfW/9dyRPq1JJ/RowYvXvlfJxlXpXZ0z9zFt9bKHLCWWjFdxZfnnh5xn5UDsZ/Qrfutw
eji0wtg0oP4YjsI2kXtVstSqwQ8hDZBECQGc0Cdz3CZ8nQglodx0RjfuWkCRuzng2a2lFOZ3ojWj
PlgXeccpFHfEOQmdJ9FRE3SvXTvCX1uFX/8Yoy9Nx8yGl/b/eb+TrxCpF36Rmcc1pLvCKToOA3zS
QJjnLmt1xb+p+cTUcIoj/rtWkalW1qi//TTUFiYULgXsmIgLfm6aKs+ucKAzRzEWS8v5JZfZ/58b
JjC88U8RD7l6g3wqGY0nPrjodrKj/u55NW/D2f5pBEorvDPf+CXXp7oUJGBUhXT24QD/ffGXhfHg
6A4+wjeVIl0rl+yA127hfbhkAKeTkPKPFuEvZje1uRW7aPhpem90Ff+3gcXXrfXnJQGVI3mZR7gM
HrAojEE7HUuClxsUyGROMGfZTgVvtaNhyYB+AZpfIVJN9X0tMP7PH+unELFznfLqb6C+IsID9snh
yclReUI8ZVI6Exfi9THlEdzMkbh5jcXkb/gOW2/ohh+Fi9MTMKJWVcTEaoOk8UOuwrRVtH7ISa4L
DaaoO7N6OLedSq5bNI6WMUWoArMWbA3esgeny0qZYG0H/Jhnmn04fCRuEd5IKafikJ2n+YGC5KVp
Ae91nZ07ag/asL387NWewAOaJfgU2S53JdCU3YDUG3HS7cNk7gekpomudfvSL6gm5cx0Slk1bpq3
LV5ZL1sRaOsVoJt+D9lqynI2VmAzqD1gG7JdsadaoC0LFx9AR5kJPWFOmnf+4pErpqKkXuwdneaI
Me4dapKKen4zOA+k2PP6at1c4m9hII8jM7t32fO7ZIozig+GVLJNA0BWbexqqLhHu2MmpiZhgUHK
UfAnAhj5qWg58My/uUdTzW0ZAqFFEtnyQFVeZ9uy2YEsu2pBCUXd4eyhylPAzPGklMT5Q3bileef
/hzFcaqBVBpeGufPJBIGqNB23lGsCE/FBPDwXz1aJVef1eU8l5XAIpQrr4gWF4pqWUFQllhHQ5A6
rALge1fhlMchIgQlFquovXhHPSJ9s9H37JLoIcLRDIX40kXnc8gd/acYXzK5JWkRKaRRQzlIwNsc
bdRD4UeBB2wcSqGUn7r1+g9PjscFI31V6Ar8oE0PJn2yQYEnPite5DqW5ZwOAkQAtNa5O4R/WMWN
uXeSqiSvRiSj6TAuTVZrRjsPPWtZ91qatsuywuBYJpRoUmsj83n+4B7+WPbefe9rGKMkpdA73Hqu
K/rFURzMm69gmK+M2OIhKibShm+MknnzeATKqlLXPPhxHqGPb9Dve9GqiFgoWQB7E/kk/NVNSREy
fSmCqMouCEVRQTEkwWp31qTobpqdc1C6rZGmElx9A+PhN0QfuTTC2bfMbZbp6ilT2w9bD1RmCnf1
8W6NvRBalgy9JzsuzGdEChCPePx/gZybn0itH8r3EMBKCupKGIlkttHH9NtWi4kPaZaVid53uLYr
3/XanISFbbYttIO3eR02WOkXO+FMDqkwxJVkRxBLrmWOj0ACflqh04SN5xEzsHKqestB8adr5yfL
KWH1azqtxOsWjxB/I0g4Ba/HZwFWkIG3Lz3eVOAwmmgsXxM2M5ONvNNi6LFYrBRKuVjyPziAch16
61RYNlhADKBPjqVdarDs8IcCcF1pJY2XP4eTl3MxnDqetPOGQrjHGb4yxBDepRXYlqB55FG0j5Hs
a358Oqa4n/152VgLOJMPCfRcGkwGX/8zbBrB25wV3iDZfPa8edME50onzpBNd91shybpAbxW3B+h
4Tzd5GCUcFN2NC02Usopi21zD1VXb56WpyXZagnLcRBvAHzPDyZ1R3qWUZFuBj5nfVhH0tQHq7rp
F1SDj2PulsuHegAbZSGAgv0Gudl6XN0foZJ5Yp2Xo/iSE/6J7zwXIm80v+i/uAfXBS8GmNLNT8ln
3yALX1x95F3Skzb1SA27esD9xZKVbz+YOoGP6ZadJh/jm/hRsmUFfjw8B6nxlIyFOak1JdVErz3m
59QL8/i0KZeh9DPLTscqVp303CZi7/2OUQCVwZFqy7liO1sbHFh9BBZm+Dy81PxZU5voY7Ep2YOW
xJMkUAakEsZ4KueakU/j/Sgg1fFDwxVntcQuj2uSVmRirPKB4eSV+xCaLXdwqV2zIzgE5xmXOLVy
BGb+ATKAOwZeUh/kqSapHeLQ4TJoVlGcOHQSB+D4+Sk9NfZoUflsQkU/xVa6VN4BhNoMxw3ZdMPH
ypnmqUzHPP0piusD8SFGFcnMUxJLjDI5UiQG8zCjA5iv+VGpI2majysh8mNOwpHYeVY8lw9ldFf0
lMmDbCF9QbNAUShiGfnjyDZBvxCU/6kNEvqFWD9vChtyHhy8fKphu6SMugvuIGoJusth72GQDf9U
zk+VyKeKtdlmIeIMpqxwbmP97nUYmoLAB/FGwxYVO7SfHnWuaqlV74KHCXaOcZTKDSmWnNvNaMru
QRgO+a6fGN1p9MHuibmbcXsi9Ub+9qgpektei1wdBANEBxDqOJ3mnY9HIB5q48IOHsNubU4+rH5z
/E7jW5kXyS2IMQwDcDiK+WXC//R+1awX9zlk1qMjBVbaZCviEZuuXf/UgWLnEomFTOLi8wWJ+ron
mVq2Yr9s/ur8AOE+sT3IvF9/BFRnV8+WrkwcISiZRG2Z5q7Tda6FSHEgz2VbrTgRDIy2B1CDgKWJ
Wtvm8YtiCKRVTJDLhtMSQoX5yjeJQ8rczk4Zx6yxgZIf1Nf+ATiHngP8kKJiWFPEJgoDAK+YmFZB
xmLZmQFUwiNS0wE0wo+tmONx2azNKQQ7B2algLCEw+BEEHHaHNBBl1cUrbXMp6lPN+1yCPgDTHdv
rnRTui5mKdUGQvBZmAZuhEWVtxT4du3v5zQcuM5U+sR6k1naCatZhrPyULNQZxTdVUxKEt272Deq
7ryRGYubg2nuQyLch0zYTJlpVxO77WvnkEqSTZKCz0DYHK0Nwbu1NAjY0QpUzwbfY72Rc9pWD0rQ
d5Y55zbp3Q9P02VL6cllNkmIfse1vRSZ9xuD7m1qQrIpnacsw06WDhoqj1XPateop8jxQP2R7adC
ejZQqyPW5mIo91rNTr6+ML6vE6wn11znbuIPlWjA0ItnxS/Gvvlny8KSBss4gnUQfGCG+gL+FDSr
I9rOsXvNV/qOgZP4vNT5+yZpAlamHP7aLFv5i6FJXElVOkmShdMfQ3bs36/n7oTARntyBesRMPfn
ORphqa1dtyvjN085OhsSU4lYui84feAIn9sqE5u1nIetDg7IuEz03ur+t3DoXWcDmDfdq9aFEsIC
SVdekoBfSRip5/Gi3lABdaVvm58QB7q75XSfMIEgtjsmTMMcfesccdhM21C26sxJ84Ay9eCA/hsr
fXS733tRTRyWyeiMRyovBug3DMwYS6l5ABPM1YnPALVQt76c1WGxAMoDxsW9iufqG6ARYT6PKr7j
TQNwRyj1nP3kWVDXJdU7L5yQuxcQ5pg34JnZNpjnAayMXV2SPsuPUjYYfs73MT/33n93J/UF84I4
C2VC5O9CaTW8VK+jce8BOhpE9KJFO0KNxULiWSE04mrE1jUMkZhU4elpg0nfHEq7Z6oz0S6J3B5P
O0XH1Z10zhwaEOzzloRj4XCeZGv7F2+g1i1LwVnffsPsR0Cy2GBvd8O6TpblGl93Ldvv3EsHX0n6
0XpGc6ryer6d+nnjZES9Zs0/KB8t0YLDkU94xqAstBqkqxh+0UfiL8FjxpAVpbqUM10oiStCn1eE
b605Z/O4McTGLSPFMOTbm2nBTy0U0HLL7ICwm/Q4uC97rUOfi9sdFJl42ApBrNlOP6bHasZcAKoR
cnG7wwprtmrHxlJAh85RpTtmPHygqq4ZwMnTMPj3rgXxtJHT2tSpIN1pX4BKKXmerTyAnM/zYSyL
EWgIr0P+tCNaaRP2fpF2ZY3rt+ZfgY3RpTm7u5ZL3m5i5BOXCFP+NGu92/zI9jzCHig8q6j9Gm9+
u4Hdf1/rrsUxjjWse5Nkq4jzABeWoNpwJI3wFrfpX6rKgnDuAW4ynFpWmI3t2ky6QoE0NsBu6dcr
rU0pps13BEdssck4WA08A7WbwQkisMO0PDtctV246pwsdjmIo1Vv2qSQngynSJj6dIL/IaAoRCJh
zy3SqvMjI+U7xaIloGbyGRi/R7p63mJ7q+UciwUNapQpKmraXG1Y/qljeOFRm6sFdHq0PalyiLyn
x1UsAOpo/9zEeYEOGfl+RzGwdP5QjWloAAKfSVvaKpmKWOP4j50giaJz/Ona/kWYzZqcpLJv2GkT
yeY3+AcGlIP3LUCDWLXfqKyarbsV+Nlc40BZzxCnCU/B6OZ8qUQsc0pufLdgL6461cAi6cHZx5Ht
PEqy44xMTSFK/pi+GKQD0pKC6DWaHHWgBND3jCxAGLGHbcVZPHG0YFKNa03zuD3uviHno1zs0ws/
F0forLP0nPhtWUmrQyen7IP8klrch2O3gbZFh+KUZ5Q4QxniueyDg7KFs7E4b+n8RYisCIj+xwU0
C4wT1X0w09tCHvdLiaht9EBuCzS5TN30xiF0tV3/1NZXI27YlrCiGVmO7NOwVzLqgpZQBQqEKEPU
8QA1L3tbzVOki/pANRvqckH6yJgGQOywFHDqLyUF3szTchyNBZ87eMtzZKinwtZFVKfHd4MvrJq2
XM4Dzxc51ZRq6VI0g2KgM7/SvWoPejBaoGYuI3Mgbbz+U6wazFhMCv0ZXhE/qHC6gMGHrna9Jr2f
AasLPeXVajIo+mPV13Sfh/lrnNfElT85kXbdJVevRA1SXj8DVmXlHYeSGjA9P1NAs2tOiPSoahS7
MA/x3mIGYSTdHYF1KUIfPO0VmspbuuJdTdgrsF0kB1lqlRjIIMoBQ3Q/w0P93oIiyGd7XXgO9Du/
hvDMM5ZRl4AsAuRlZ+cwhUe3JrIfqLB3zmuIyCn+3YGvnJgaQ8qHPn2Jo0D12riPlqzegF1qxs4X
CQMGdGXXeEm82uLlhd2iPmAG+RB3PpVSVxPEaM6V8xYTRp/0bNRPNDgtsFAlo+f4uJ3XRKXROk4p
SBdJ85i6u9/r6ElnqUs+apHOUi/AL05oLxSDuL2fv5/q5P6edPnk6K0cvwwiuI0zusiHttwguIkP
zUDinlXDByIZtF323nKe9x/mSxx+LUvKL/8fis+vYyC1YzSuFDQVgCKWBnV+BGG0YQupXaH7IpYZ
VRPdcbnCF4NAS6ETQSv5axjfshzxZWcw0U5qpLg79fB41sRQiYfVyn1BXPR2C2fOqDKec7bsJ3Wt
TEtCTTo6cgFmh7bOty9CwsOf5RWmvW51K2xRv1ypR5MYG41QQ1QMRyvOmgsoFxNV4xo/PsZ7sPtq
ZVf62c+7dhXGS+zK+SaKQOWe10FUA8mwXP6VDBdquWgVHrMeeMotgncE0cfTkxlavqXYpGEoPk5u
oZQoNhaG9sYoZLchKgVfbGsz3zHQjOa/EJ9NBG5XKp/mEFm5GPAsfsfgsGo4FoyK+Pgc/vnnhUhk
xwU70izUCCRLLp7eVil9sMrICp+Cx0hNb3Dy/5zkAIzAH+6TENIhS5crmGGiR3MljhIBQi5eVaTD
a8Pu+XRWCnWn4aEC4HGOPouOjxRNFJLrkP39DS+RoVQufjOsn9Brbd6rp7z6Fj48KK8mNAK6wt7j
qG1IJnQ0OGCa0XLhJO5imkmyezqjcQKAq0GcRcuJstROtQhwHZH95+dwAEbEthFm3LZ3qe1+Wp/Y
WZXE9s867xQ59Oa4ptXGvTPFwwElUKEOp2M0DJ1gb20nLqm6Gyy5mWrSc4cyaqRsajuye4ra/+JL
xKmDbdaF2XNW2PBw6VsXtBsivy1gn9RQ7NQxGyTI9V+Ee+AN3j+oanFrN8nmJsHnGoOY7GteZP5q
h+1tXhLlyzKGebJVmXSMlwQSL9gPs1MUhMq/CQKpnwIbdVteUfJ4kb6QuRXmgS7KOCyPNw+ORL2N
SVU4c7grE2HsyOSPM1hKW0kle9NzEM0smblWTZEAE1Lm6CutEmbo+zYXuCIetX5QzYSNYTqxHHwV
kf+blbiXfkoOdSQ7MIm9wr1ak1pBKh/g8SPTph+67F9mIHl6Kyki+KvE2mi0u76Wc83jV1zeFjhl
2B3MBWw2YwDm5nZAA2qnJKagUlcoctBcyjekpYvajeUrxbU7UeWbp8ASsbUvetBhW1pSFuOdgtQY
T9Q0sknYQ4+VmrUWk4UQgajHR3laxygB7iMs7Z18phakVLLWcSkzNnh0xWC7VQeHOHBo+sln2NM2
OHbeowi+8EgEzCKdVIyEg+NaU3heJtXYVchqKtFOOFUP4AFCpyGwAyYyguPJag+JrqNiCqB8uJAx
U3VDunQoOJwIq6JnGJ8XsdK6RQRr/tvI0vLKlLOarm6pOA4ATTvU9XiACEWf093BpURopMqnjba3
SPhB5Bg9rLc5bF71eDy529ugA7jGhoSNifDmFDgrPGZIGSgzTmyq7a8nLsJfAgT66MFnXkXNq7eB
bLUrjej3nedS8VIKwdB2fIPF3qQkG1IYQOcm1yvtR3rDlO4DNOlHs1/l+iddGJDV2jBbwJnjDPxu
NUrx7rzPriPiNyAVSchs+Fhc25fFTkGzg3rpBerB1n424C6AZu9pIG3ws/9u42zKDBu7vJmVyxUA
3BYxMVRTnYn2gy1kITYb1w1CfMjnKyPupglfYm/2suyUC+8Uij1B6N4GHYkUzO1lzlDty0P4WvZA
3Nkbuwo3cDUAtWu7STXJi9HgIJEIFiVDewZRHSOeG4il6J/uWAKsTHxlskmyMGr9Z+r3RRwxtlmo
1DefcFYZ01Y/fV5C67UAiW9c3TIb6h6dWjKjyB5GVGpd3wKiDdXoWrn/G5/f1ZLUOyI76Cavua1V
o64ItuSkZC/0wZG73SQWWWEEOJdvCEItIkwE9Z6MKSbfJ0817dkCrTHW4lw+ZFsT0sV9Fl+BLLQ2
rWEuEKfJ9rVxTbvHznq/yPiVnqGtfidnlF9dLcbJF6Ab8hzHyTwTVsu1WfG7N9Qek+fSu//Q1LZq
cFEH3ao0HavhEgs1v0CSSEdzc6wt28mu98QPFJSGdssrDuqoaC29DsYcfNNiFlVTkiQofDrW6A5O
Hr3R8JakYNTgfbNbWqh4gUPPGNh9doaeXepK+LeCpTPxxJ/Aau/UK6y7wUaK3QHLS4eI1ARqs3p9
0DD+0Ciz7IlUETBUINNKANG2C12w01TPzE8L1cLWBPyFT6DoswsyPrjVPlYmD7LTQR2Y1LDQ+Gk7
v+ZBozP3fLe48zNlhD+H+1xvHP2SHDoCBAN+PT+NvQEy8hqDPv/ymzx6B7JmRJ2WAnn0c6JoeeMv
QDfWI5TukblsmhQOTuOZ01Lwabpa/9GG91lcn6zBZCBQPneQCsKrDSaw+MU97MkFYy+LLsQ5eY0t
GVsbRwnOqTnjylxyAkaLWsnckSPCbB5fhiQvhfUWA0fbV/wVkIt8M52S98CsoOrudFxsyIZp0VzQ
Xp1MXNDNXGo/k4Eu4DnBWS+TnPXOgu5vL7GtMdHRdMd6pvBsL8vfj/6hl0qjG9CLohr3QBz4MkvA
cmvuUSyrUc7ab8l9sd2CfRRz2mQHTVTHrU4W3fb59bUcWCU2OpY53nKsywhk8z4/Sp9PJL1vs07W
4/ccgoJapkMacnbxwOYY5r+FrvU4OgZ1748lUm90f/koFbps1ZDan5dudGcRTh7gseq8gUqMLaSS
EGFETafmuL0MUlzCAxR1Iac/3+4UcFecHPc2aBJZHOI/OLxb1lEAuBTUYJhsINluXgHAi/2ObTNQ
u97a/jkr3pqhBOQepE2PRprwuSLB6Ux7RyvGD/vSy1akRCrDZMT068lkXCtx4hzy8IdwsPXv28u8
0mEEyC8VSncRgmdA+O0KvEvo3zdtkwXCUSMtOwoXcou2vhZXraOjEgYAjibVrpj1iuCKZrnn9r2t
jKZzmdLQu/VHmpqeVRhMBtc0NYLDF03qXUdkYGCTEyt1IAbZQdl9LOlEHcvH/Iq3oV7PYqV1O2Tn
vvuwhkJP1I6DX442YANZvA92zlT/aYQcyF9N+U7FB3Bli58KdhDSe32SpAB/OtMzKVDF4mgvVnQB
UQuD9LXSoZXNQ6I4y2MkI1HI1Yj3bsDKzmtjxTtfpIl0sjmLS4afMZa+c3ERiLEHe+eXPk7nV6Ih
HlfMYXbAy2JDzX/Tj6Cc0rHXqNsx1NsbGiU/+8kjbtdQ50G7CXMn1QHBC3/KfH3c24oTzSL2JmxN
+g8/rMuxa4VmM5iqOtcYqg6nYvfae0jiXM8PaVKDhGTzLZQEBSSRy0xaJkPtSI7KU8VYSG4xu+Ns
jpUwRrOZ8WAPy1LYT/IaL8eLxKdHvUszyDqiQeNlhDcY7/R7hcOCK7IYa+BT7fF7k+JAmmsOhcBF
IkfmnHFahyR+GsJHZOd4I4lkwMBKUsj5GedBStgeNMPPAUZjIi5DvCWt3vBcnl/4bt1c6Bbe4vQx
fxj3urGGfEhRjl0exSTEWD868gUr84cXvKzLsVo7ccllf//WxV2wlRItZa91RjqQwy7dHVdnJngP
ftueNw8hwBKptMdvkZr9Se3Oyguo3PslEoWEuTq5yzKsa9qqigQ9D4qeWSxcd7D7KDYD9ms5U+aE
PkCQKfTGjD97lAwYLhgCoiSaqwqQRJq4emQTWxEvsfSB5q9R0s5mz7eyN3aDX7xhTpusuunnu8Ma
KF+1KVkt27LPBY/jGz8dk+PI/IpxVjKbNF8baaXNCP7O6oYmEijJ3g3Lo2sJPIJ71yU6vug0kWLU
i48WEcTjGUK944jPBp7Q+gIZz+RDeoCHagE2cET3iFk6/534JdJ/AP1IavpXpL6Aja9FfmZTe1ok
rAw/lofpWTr2QhOTt5243HHLuidodq9Nc0Mav262XbvIgHIwJ8285oYnhwj7IPl2RZ1DKfsGSQk2
d9Tq9u1fs4SP2Nwl7zrrxOSmjiDOkGbiz4kyIPHEYOfk2gGnRRtZSQT1uSP5LAZlwdooAyhLY5GN
ogxCA9NDGS25oMxtkWoFToejNGG/aHjkwMEMQUthIAbj0ETfk0RdLLaz4MYSOSSW5U2aKZOHDAiM
uEUfA0W1uiOcTjjXm++mHhPS5qul26bU0zCehxEbMAbOms1k+yn0HhtEy7X/kbhDD2VX9MsoiY4L
FKY0KAyr0naCXSDlO+9TXjdXn1a/Za8t5yAAK7QjWnUiaACmODRL8vVBRILT657lG5d6pPLCbkNh
/tDoIMb4mat+JhdZaf8c/VZUpFHKcr6GdotI+8hfPK3RoMIhwwWKgTJbFlLwQnlYtQIBKA12bVSd
s58kSkD7Wmz/viU2cn1EjBHLPSW/F3iE3z1YXn3G5C/okvhabRE7EjvmDdsVxyjXM0pHHXpfLApG
VDntSM/O6eMkGQZ4KCrRl2Wr9oraM37kIA7FFl1WmqOOrSkMaLV/zRWhvyqpZx7eyurVBYGd7w0B
al/GRDsQgVQwhggWr5Cnzpeg3NHZeLjzePBYZElZme0V9JGUcA2tTmHeF5H77++G1Tat+oKDAgXf
NqZLGkbDAM5KdNBbCKiJ0hbTSayWdVrNOtb2A96Z43SYQJVhFHgPlh0UPWwn2Asetz1HOl8sYA2P
swYujtogaYrWhIJjiO1o6py7SMjP3CyqVsPkiZJMJrUr57m/6UPvQYfKY3mf1GQt070dCP6T9ZQK
8uwUv9ZUmYKZWnvxuKs+6zzHICykmVIgpAy6HOrFfqb9wfH8ubIGRohhUTCi85noXCmaTgjQKIzz
Ql26TEkkcvNZF3y/rVp4Dk8FWRvD4IxtBJwqyL5Up1vOxj5D0V9SWyHI+2QMJGsU+jxkFiKPk1kC
3+RaBS2bvJ3QJrb4RiMMoO32a3Z8vh0kne/nf1XwvLPwqmuRt2A2GcEwCD7YjZpZ4YVM2137DaEP
dkZ0uorfVNI2zAUI84lM2LK9rBX1gnKfAXZrEhBWXXT5OaA8+Shs59wieFLu4/Rzr8dB+GyjH14p
Tg2Y+LJLb4j612E2fo/+l/+WSEHzoyWsBRdDHhxtjQ4YUQZcwpbUsX68qQbYycjyjVMtQ3SHt4dU
OywuX2Y7Za1zT1Xp/UVW9sECVu/n2gcbtzifk1Q4VhFA0T0jN/LhN6ak64NCP9pokqMh3MW/IAdC
4zCtaA+jUbSAQ4WZd5cqmRKkZ2t7JZcT9IDgM551X48fieOa+uugKZNrXYf372757CXPM3reuLNJ
CPo4mHTjsxU+Fwn6HiQfzTIMHOYQkj+vrzGM36uBYVK291hyBW8UztiU1Cr1RVkO7nMv20IlrhGl
poWwmSoYOC7irYFNvckRg7OjntjQYZ9q15z7L4cVLfdh7gPSajcl8CMDJMTiAqQRY5E4rtaxzaxe
qWVslz5ANni99yXnSEQhpWEm/fcZl/TXshtW0YUlg4M6H1sNEg+wHIOJauh7vLrX004gLsf/rq+l
wZFjOsVTAhgPYNDnMPGueLDACWjl/FGCiFSNrS5+D7/MS239vpZIM+8I90y6XUyJ9MWKydBW6S8Z
K/gVSYr6m0inLrEQIBwh9y1DWSP5d9P8RG1SSLoDeHkMQq5wRZVZFE3lrRNjmMqD+Riffsc4QFyZ
jwBFbE2EM7/v3pwISaVC0zhI5gbfeOPqom0JpjBsoq2A5AnNDcjKFc64rJQPFQ3znljHKYkdnU0b
xL1AY/49wGraO/UeZYk9n8Xa1BKXJHgfreXwvSoIrd29ZYvWYkdlieaN+/pKGgWlAywFmhGoDrtS
pmyKKqOcz/THS5GYuYsHBq/d0cs6x6w8LuKbuAUTVK9PY6Je5rzlhf1bWIop/fb8AVuQn/poTD7s
Uy3zeY5JM7UHMdpeGrdQSl+f1/4G0h8YJo8WmtVNeu0johQHifeLYIiyEOzvU8wXoZu/fcGknETp
gEQEO+HPMqe6rSXzg6f/siyxpdcjC70/Cz8Aa+5xv5DcV5a80VcicWSLBIAz+lpiHaNsSpvMer5k
pAn3n0dJJJiMX3jHKCSDVgyAS3MwyWFr2zsBLjxzr0uXnEX4hXSU2ntuWjQEkh9l7/OkCk5/kPq/
USqWKDLlKjKXX9ZKSnyMWTxef4aT5QoDx3bFH8VypGId4fjSUgICgiC9CyaV6NOeVtCanDXtZtQd
mVG6aul8nwvMD1IlLzw8w3ntyz3W4+vtdiUawlGBSDuNsz8zb8eJNcsTsbtRTNs+N+h0LLt/7mCB
v4OAbJpQcynC6APjSePaMpPI/tuVR8syG9H8FQHl0fQyC1nmeGaUGlkf2QKIi+OIjlpiOmWV3bs2
wTddHXomQFQc/XYvbpEGvFIr7tGnbPL5qO+bDWZXJ0yMcMImcBNVkE4ASOmaFgHAnEPwzTFJgu3N
jHq5R4RujSo27ppTniXvyKwDNgbVsKP6Yh1tGxNJ0CFgSCWgRSqK1L1u0l5cKDvdGNZrviadKB9c
extNL0ste80TB0QHbtkx6EtkYyHAkLI4tQA1FuiGndNDHA2QowunTeljO2/ZeUqWUg/9V93JscG7
0JFJMgtVNPrPPtZaun4Q5SnfjDG0HQZFJTJk8zsY/CPduzBp3YWSWSgu80RCaCtTILdSv4g1qOrL
e9diSeQ8y3PQzwJI9TXnJLL/FLROdBGvxFm6WWQtGr4uOA1ojID/NHpJzKnAlrcgrWByKpKdNkN4
jVXtrn3enNnStrDgVEOUdb9a5CrXpCz0hoSb/vY9jw+uVcbfL4Gtx7vPMS+bbidOKvJbqwPC4CAh
q5aqTUe70ARSmOobNLyhFNJChev7EdxApyC7m+jOCHdJftjMGl8AnyMgGAOH7EaVemoPcGQl00U8
WmqCn6XDdjo1Ipebk8mWpUgf8KA8W1W62sIDExUoBUj/EByDBztokh0egPXKOHpgth7jpzMQMqMJ
1aIMQoh40uhQxmN83zZpooiBftnEEfQUGuVon0L6Y+/LrnC+IN17ZYB2mN7Q+D/hP6HZ3Pq3MR7X
LneYLbBa19YRymbgfF9ZUUwi/244cU3qK5bjGc/KwD4GtfIHziPhuBvtACgg0JqejIgEDzqqCmuk
zo4JJJTtdISy6yL3kJcFxXcHEtQZ4dfwG1XmXadWiyNAKWFEaMO3n7d2qBsQVwaYU2aaanmdPuCJ
EoPqCqt/StCmcVeOccqTYvPjE5do9/cIuN+PnWC6+fLsElgg0X4ly7FGaD0c8Q8D6kR8jwIMd/Za
tN8sEq8Rh22Zb7Qrp1+FoUqsuCtzqRLnKZNTCC4q+oYzZVSmBULg7hMXUlL+PtONk8BNVoqEvoUK
Df39UusSoOfswzW8/QeiD4I/uW5amV5JqjdEZ4m1YbVhlyueOzQztuLN/jQYwqzVEVvQn71xcs4+
Ft4lyoHl3E3Ee7fcI5dalX2aOuyL3apxFur0MZk6Ox8r2hLVR/63PIk14qGwyvaqZyN7zL+XenXB
feQCS1If9abnHEWWMhezZqxv758RteehGv3N2x+x57chzG2d4/v5PotI6qqNACeh673xeEw1EoPA
e6VMmvZZBS0XCS5wthn4uFh36bhbVOVn6HvgaSb6zl/zN/kPmr9Vb2mZFlplXuHAev76zNSJ/FVy
GcujwEuTyZ5pduGso108RCBINPz1T4N0ktk+myYEIBMmNSCuxPIZLZMtOGYu9JV7wJe/z1IoVNlU
81r5hJHnHRc8wzASNy8qAqWXU6bVHLOD6eX+TOUTJm8r5QkhI3xKcA6usKzjJub0PuVV49ZxRsNm
r4jwUwlWZ8K51ivdS1UwqG/aeihphh3UMZA41GS2UR4WiN/4m02J1nLVkTBncsAEOn8GExIGc2qd
vwKqNxKik5yQQUX7UwLzq9gA3VTwHrf4ky98K4bdsGwfWUWwhQmrB3o+nCdi6q3yf0ddDSB6sJob
/xGXvOX2Vy6FYoUDTIGUu8uoP9JDkzKCKVT643M10IIdhSzdOiXzN01kF0SNPSs+YbO0w+xzwiTA
h/a1lDkCOud3VpbiWntnWWyHHiTfYqeWLvqrKv9SNb/3s4QH/w01+8k0PxLfYOx9Ep/vXzfVwI/p
BiEfQ8bo3HYqyDMIu1KnmNx47y4pRNUJmzotWZC9IFWD0oaN3zWXmD7V7SWdU1ppiwKedu1Qx82T
wv6tlm1XyvcLA9+bN+rBAAmBo1LM09gynseb3iBXUVU52dnfO48Qgkj7oZ38negPPMELBNRLZfHQ
TUm3S2tNrhlEkL7nVIwhM6QBm68OZzg7VcJvSKXhN98qMzFbtT5+c7RLJksFjFeoUrnctjAr7rqX
KJG9pm/0RRQsQoF8LRxIGvSfvXLQnIo0TUUtA7+RP8Nk8qQbRDJtdxQvGkdjpLPLlbEWFua8xCrV
qBvLZ5F6qnjr4Yt7LA3OSU+bpiUjJcsZrAsa6WdaurGFyhapKMM9yDX28OL0/PLPgCeeKw4D6Q1j
jEnMnIq1pGJve8b33xi0lbQvAe6VgFkvJYSWgHsmS6Qyyn13/xa0y+PuIQOezshaWgHwhO15dIVV
PAOxbSBXr/2ilMBIKMFCl+jcrHxnpzpQs0HZfJRxXyzqmGsZKo6fn258xFZCLa2EVwg+RJdWv5FG
EnoPsQ4uZEj1f6FRbGCPsTEb4XNgEJaXonzFJMBXRCVEpAV4grbPdqBcImHNmhWoJunE/gii1xJw
rfT5NIf0p9rqmdBoX3n2+3YihjnkCnlmPfCdeDSOQGumz1l1RuZ44CBQNhyI2S9PwipQ+rYpBKZ5
hxohCzhh+1NYuA82/OKJHI4AXdY89H1S1RdouBMiRRZ8V4064h+Q3XiquWVjTgyGoZiDqoJdRkb2
zoVxBhGTEgqCZG/DaQNkZmcVrVo5s/mPZWTYXf0540N3XcL62G3CZDt6eZusjWYlJjk5l0OJv05A
0uFPv2opmXCpDfXfDwFBD8Uw5gzrx9qkjSbv4L3EOdW8h6KTgWmCA3EnNNtuWc+dc18Dirw9SaeI
wN/jfEGZAW47TKJkpLFl+lF9WbaTGTkf3JJql4EImxxqFOc+nWrPg3VkhpoirUSNKSNuPehVPc+0
F7qkoxuWxwDo5l0cHLNEwc9pbzjHJh4pYu7wARpqaIwuhRxope1G+O3tbXBNxXtEHAnXfjOUfL3U
/+FQ+z6M8aaXt2HXuFvihGIQcdMi1BBrSnwYUlljg7sbRw3x73ehKATE+Ir30EDyZK08Ne7OXv+x
sU0XVZup2D+bciKFG1xnQV837zl8iV9GLTZSG7n846cv0Wa68SzvRroJhYHYokgphqJfezbeVORG
vTHIKLgvYHSxnuKns5PmoTtV21DPVcHz4of1nnIpXk1k4hc2mkWbCLsvKyAzEF8e+8vDa2iZjOWE
Q8LhOwRXEbfwxT+wkjhbBHsQiMWY1NGcU5n8FPz9Wiy9igoZ42yANNZcceDULStOdkkYWS+NPBpY
LcijwFvwWiqFUuZK5025ah75lLa7eg85gGi8fRGokA5DDayyjQAzcF8WKVuiRfqlwQH9eKjF8cho
xgrKMFbNAhmDC/CILV90QV5qfC63XpUbKAHHTaFwHP5PytXNhPXxs6frQPzeX36HDaKswPoeBWOI
ZfphdcXurVu6GNFv1JSrIioKyv7+Oh3z/T1oJEFdalyMC9+Nz/vgZlmndn3Beq0hmvb+U7qIVr1g
7vy0NaNcHcNjR3rdfnh3hDkHycuj6Mi5ttLbFmYYwxf+RFM5I6X6Vr6cmBko/FjtouN45WC7rb00
OaY6dA9R+Crj+Gj6w72CfVNs4zZHlQiLfRgv9oI951PkICJ32kYWZQjp9RTTldzjPpkD/s+uDq1J
tuimijad4ibsdOROoJ65O0y5Og9Nmq9AID0mLqkY8NEKMqtNVOndEjYQ1HSSWPuIkf3XdVmqyJTK
kVbm4Zhvpfn1gJpwqN1ITPLkR8DRQ6IgMETcsIAoE2FFZSQbKWE/VegozWQ2XlAOyL2M9R8RWLAY
byVwQTh3Qs/n37K0xmkW2E2/jGyi6NQxGouIdcAeAmZvPRBLhWO6lbrM+V8CmJn55lCSAEj6wD1Z
mY9b78TQTSwwLbzuwzAdeO2NLRS5Nu1+hEUfsqOFvACqaZmjTMSQ7iakr+yKxNJPiFRA7v0XbN2l
BZczRUbozjq7EwxESH7ICPMRehnPVFHsSopagMdFYjal9QaUY4bBH95seFFTtJ4liEkZj5LyWb4J
I+eAo0WSN1GeHRDTu9m7I7ilRHt+UnSn35jvZf+gktOy6BRFy/aPi/Alm32+Lge9UCO4LFYBwsFH
e0p8Us3coTC1zw8tbdnT4CqGbRJ76zqezF0MNFmu5aqC1rU9IOVsWcpu0yVNsiVtugY/1Nrl4vsb
YJ6C8MygUyfpkQMtgF9UHxUZI20wn9+x0L4z6Q81ykEa8e5FHqA2/xBQYx+UIF2wHU+unGFmj+5O
GCXeRQ1R0xXWcQLgmGtSMhEexjOzaPWyBRNYqBPHvZtEalTMESGxfj5gTGqUgZGY2pTEpxjcnSMQ
xrEYjWizXFk4ccGeJ1hy5gMmeZp+Lh1C2CVj19kxpsZmhSRSc+gwe5iw1crtpcxmKc5mdO+mjrac
/AIxbAY+fR0c30dSYmFW3GOfol/Wo24RPLhhsHTWnp5q1B2NXjFV3mTqkeuUXDzo09My1pT4Vd4g
4l5W0O/I8YRh2dAqS9BXoyLZZLeMumLq2KBnuxrtN7i0ZbQuLhZtTpaX/qMk0FB0E8/ANWcAUJ1q
/hUI3jyHPwr+BTP5KTBqNxMdT1+IA5rNAqFvQB2nPtVuqluVjduHiZWH+26aNQ/cFmLMgMBhidOW
8Q9kciI5bLMSoC2Z1zs091ApYtkmg/J13PzTTmVwxzI+0hBg6xZWNTCDjeRUGixXP+v2mftIAT10
K/av8FQptZchV0RrswmfqBsKQycyhm2jPQERUvuvnOT0J8TMTDBc08lhpGvT6VtmeChT92S0PpYB
9EZ7GXJrAKDAk/f18tngFpPZpgwVK1W4rkhJI91ZySilDY8zf8NXUyLq6YhsN/IDQxFaeV7++dcL
WXkUhuNaK738Fk8sXl0oKpCAiZBwhZQ3ubm82YuWprnKGuK4yHbC1tORmsSDalxRnslLpJYjlvJO
CS1filSVVIQbsJJ5XUkU5dcBSo4Bent609ZoXhrr6GkWK059cCquYwBMEbkvObe/06eDAazJoA46
lQgOpFx8NyFv6PSNeAR8NWRkxoC+4ZCihF3D64crdrpnaLn43kSN384M5T1NkWsfvoHiqWvYag3d
LzgnUJRFmh0/FTThKXRFfRaCvlqauRlG+sPPRiZUnl7K6RnubTVuEXFkWW+itNFeiotWbqlKq9Bl
VfxQ/2PWYSXBQmYLjZ2y6/a8xY/46SUyyuVO3LhFQ/kuqmEIwjr/InZfGPr919+nCH5Qx2pWXMA6
a1khD2R59YpSwU8KSHf1esi5EZg2/ERU8UcS5w0gsStUb/ErwVnkQsT6txM8zSYTCOPP2S/6Qvgp
eWBKXqJOFfpTJrpqmbAbtCUmOlbA8eo2Gia+G/N+Xybeb+ZpsWCYMUqJF+KLkZYyfVhBGdd23jo4
NZPu+JKttHf4UuCrajZTyiyKJ+t9GBheL4LRZMEt9HoisghiB1AB5T9XLLECNYxVYMWapL8p98Cp
Upww7MgUtpq5uupeVK43pryv9+Q372JOqsfkCLgqKcwAMiN9816OKZxsKuIjgFeULyVDTMJD7tf8
XLiJ+yRDXm+SzMpul+xrEnOD+heRkuQGw0IYsSxkZex/cmnYURWmHKYKe9JCNZOF+Rsr/zB1ecOp
INPjp65cunte2Yi4DCrO3eoWbDhhb/EsRoDtKHLsHx2bzLdMFu+9hWjM0p8zJuQyM/H4JJ47j0OY
Im6Ibdn/IYnu5f3Up6HdLp+2wBXdfSSxV468vUMiTVIZzbRkrJIUAdu1MiX6WqJuE3wFPew3WUs0
kXLEpFTqqU+NbNEQkVKue2VQ4b5A5S9GPKYorWPJGOE1/HEM4fchl8UGBj/PasF7iWsTCjszqek5
SQSPqaSAAoVpl5EW8UQzPJABBxNWB4PRwFqurn+AmAfk0TTHNKsf75l+7WZDcdVGPB0LuIMBPFUJ
CK45DOuixpuxxltY2yNg9M4K/FBeJucIB9lbEf7hOgV+DIXPfrejJ8glh60/cZoe66nuTm3GnG0I
TclWTT9XQzdQ3ASeKmZqD6kZRmMtCAjGVS2rlLiz9cb0UCBwzroA0b1akMr4elPIICFJ8qmmRURd
DYJINzgmjTibvYaRDqEGo44GD3Ym0vYU9FyRGOJRJuDYAx9Iesde6x/zrIMMn9FOelfsn44raRFl
+B3O7QDwWttT5mwQA0ceaTJoSmEDn1WyVvVINF51wr0hjKDkMco/rSnuAo4P0+6vZN3sab0SkNyS
JHnuHgLroDs1u6XU3EMWDeb+xx58CC7nNFoMt2PIVZiMYXja5vvsUVzWUkFwYZN2oerLGE/W4wyc
TbjnoeT5b9qAIJkXTN2ZaMMqYnfegbay0Lgr6yleA4wXVkW390enjcmNryP7MtHAXrYxM9Dz0gkO
F6+EedSetHxRWG8AOxgNEXMKiaKrRNEqspAOqIM5eJnghq2C9Ise8OEDaxjnCOZiQKcKwEsvKCYH
t0+BTvl3+qlJyjf8mRBgBCqTjy4WkXVlmaH8HZbBQj+8h10DnduTHEngig5UavQqmatAi5ODXwv9
bNB0SqVA9wrmwxQXpZKzwgMq9wGAG5JSp37HtMcx2QHzexsBGpBtiL/4nEZo6dQkA36zNKD9QiCW
j1cKS3ErZr3/42JANyOTSRNPMW8flZtVeTcK9WO1n0CLqCktg5ZRmVyQOlRRPztT3QJvZ+5g0yJA
o6ORNy9/Er0XDLB39L/2kDV3RXjcRo0raQ/vuncWENzdTdPOW9qCmXqEcjbj7sufyFQ4KAxFgVlU
HeaSo+scUzf+V4Jrh3z/e2Edk14qEXwe/upj74yT5x4Sn1G6JAw18/ASjc32OhA/WjZhHrMLbJt+
9OaAxHmvJxmQpb8SGvzdSYwDQEdA0etKT1QgQ3G6rQ1jmdnx4j5bYCMDBBtjd9TftawCN+P0oEPi
E5x9HkXa4MCtft7ojsiS9eYNGkd1YEAGoLByMdWC1NSKpEcCznd+yHOX+YrfnhNYGNImjj5mBtrh
/1QG65WAwUgGRiQiMzL4knUXzOaaPySanSw9GQTYu/imKYmQhpfERM6c+oifkYtfECL9uLhd7msy
V/t+9lebkcDp+7rDVKk08s95T+MVPMGSuZoFeBeHMtz3mWi+9PWOD7wxX0ycd9lhsf6rj0YD7qdm
nXsKKUuqYwqWqZqLYZ79KZrUqQpA2WA7a5nABUGRAwdx5HxhGZEmn7q0jhbEScKGjvvEBkXkoRwL
FSmkU7zQkBe/x8/22OrH9V37dUugSUwkiNi+z66BBkPfPgDXO3VcXqiv0gnJGWbf24dl54k81HWI
tPuiLotbr5fqVIy5dH62D25TfnR/1WZ36YShSXLc0B+yz04Uru4dzGP6tULoQ/8iXjlIGjycCQ1W
kUOpLeCEdtoIEjD/dKWGzw1lG1+hi5G9dh75LW1eNmK+O5ADYEGU2lgoVz0RiNZPREunp7MMdKRi
Ah36jlTe/TgmPo35bFeZDsQzwFWMYg3B2q3bUI6SfhljTFr0ctkn0e9QGMe1Jfcc7/st7lVLAoW3
D7LmuMqbgDec2hVKxeq9OUw1hSXR3oz6JS2vvC7XjQUtDKYZjPKnkjilw/YE1iGy1PJLpqkdZ4Lp
C3ABCah+rhsPBZITLHjjrZQ/cSrGTz3cvtoJilX/9GkCUUGU0QQmg98LOnM1JfFiMawC914Dnasj
C6tXI3Gk5ayz3CQzdimLIGUVnI6LTP3YGeRYaPshQlsxT61JvAfDWHm0byIqj6uiOSgmE3eMcYz0
OEL8b5kKm50mzQ+tFkz/X8gVa+Xn2eQWuxxjhjqyYzCTx/Jri77CLp7HgmejHnjrMl7fjjrWSgoG
90Xrlly+gYDOKPKJWaH1jX3oAjN4vTLrKnR05PIC6HqEiI1B2YwlZjvjAzGrnttDnX3YDRDoFK90
+TbXvq3r/m/dhppGS06BTeeaJY7s0xABTBmoV9IdAKU3RmvgOU4R4gpEN9jxhONq80jPyp7XXYuy
WJ9rLhQDctt+12Z9ccCDHYzZn+AW+F9zA03KDrohicG/cJ/R5EpdViXOwmRLuxBMkc9RGZ5IHNZx
Z5I/mTF0Ky4N9sET6s4Q8iVI8z89b073mws7qRag1O2TZxOm20jh2H05e7TuzE2lcjOV6BMMg1aF
Z9AKEPYpeHIBN5xRhyZ2iO43DfiuDB8UZK66MiVFFnm2dMRQS9a2AKaMngYNk7wrLP53T2SiyuuE
/9uH7pxPBWlBGu7hqyvkBnjIeHjszWMeegUdxDdiWr/YpSszLs5kbXT6xTF+iWRfSEwN4kbcJ2jH
LDuwCs7NeyJCPWis2lzYhmdziJZHh0nQ2A7g4eULctyrlgfJN2Nfm/keCB2lqwgfiYKxegh4uFd7
9PgjRCXsM3jWg5F6lhSwlq66ZncpgG0QMU/5MSR0XZ+g2oibbLv3559CiIHnvqoGAROykABu278N
VnnGG8z1fDgne7LsmJfE85V25Q1hG42nyz7tUEssTn0lAbuiGvfezVj17Mvcy1T8QecXTR5YtUW+
p36WmFJlWyK/gyQ6ECVuXjrhR9YpQ2u4cWTAMV2cjiiMzSuG1dB5aC4HWbjchyDEf0Ly8P9O4fcM
grjdrk4npqdJ1RZECRGcKqnKyJG6RsrooxByb4COovITycpjstshKeO9LQciuvRzSnFB9yWMuWMf
K0FP8jy4DWZGqtifyYszVMW8ERIqFKms9pnU6mKBm8c/EHEuxivLBS6wnvF7rv3+wE+vzd7ySoH0
3bYvTGqgYBFOdbVcvW6pt/uM2NZce0j7ce5xH5jDmoDl2rp+CUjD/ctzt8DyzYUtEXowK94eWR3F
p+b1q4Y7kCc6K5qQxbhgPwtRBjep5tZn3lFz7As8nVfsLaFQ0rJx2rnbqP8R/iVj6kyIaR73vhot
mj8G+GfOa6OtzV6U0bGvl9iHmzan07aFCnXG6uR/fiovFeWB2oy8dsDgyeSCItdg+hSInUXKHxB/
eytYRQbF8d3LSYCD+uWVcSq5xoCGrxYmZFHD9TpqHNiptcVlZB4qlpb4uKMk2tTI71S9/u9JlnnN
2/r01xD34U5ERByP5omgBbOEeN6XYehmLWbEcJmYHt5oBScF3Yga+z1w/C7zlzeNMu+4jWaOS9Tl
LM0z8MNkGhFPuTnhKYa3bXRTp7cr99+SUrVDX2gGMXCTbVaJHsJCmqzutn5M200LAYIAL4rCY91m
2M9FbBAh4fCvLuLhJKpHOdKsMrRW9ap19bYvefU2e/S6Sx+OokcuKzDaB7cKabAL2vZyoKpfhCUt
04q51ApVqua1gXX0ef5fTgZR+j8YnHw8OjxmGELGK/xwcP6WUvkniSE43ju0Vicwaqda5+lbmA9t
dAd1akjno8/M4si56sBZLKNQ3Lbp8RHm55VzhxA+1eC43ZkSScNErwiRRrsGoACaADRY+y+CqxRj
Hfmo3BZgUGgCE0lgqVwy0vrHQyQy4Vo/imw57vX2DRdy//+H4DBOTrID+0jq+nDDbOhyGXvjKI+W
gG/uI8XFsbqiptNEV2Gr8vchgqXvfB4BtX+L166kt1m9Zeodf/jCIDnRnQMakTM84FWfAy8lpAge
XUjyzyCU20YZ+VsJXdZrc4IWxq1QGDBsq/mo1nE4KnujfnDyB94r1OP+UNiU6v+jQV3rs5al3hR+
ATus64sD2gZHIBjLUPpBNOXewbMrHcerxEAyWygSHxXonvMIRklgiiXz0KcUf7a0R8IGOdK/F/Os
KPXWJB7nB0F90bnHZ+kd9mEvInt1qVm4xSSb4iEU4b2S6Cigy1GQT+gPP0IN5pMYUAMcVyajxEKf
1H286WdCPtFSpnOBrkClxhQOb+orvYd1fvaPsrCdCq5bmlnks1j4Ud3h1GnvmrCV6T/CmlQMJDS3
HwU+YrBgu2t69bDPNqlGaN5zAhoLiX6890izvg8Yv+2yF5aOeu4XgyC63xv2a3PwPHOnEedRBZYw
GwI1qzLnCdaTGo66TanMNtQw8X07dpUBH1Las7urMrSkWwq4h+VP8F/4IHBLOi78ebvgk3NZTiSi
osTOzlkv+zy0pZS/zXgubR1z8vGKAIczh6zlIbwnUH8xJPoRvGRfJsFz4lBnSUdxTUNhgB0vbCPs
+h81WdVh/6IWLRVpG3WMnMAb2gw2RZm4WtfGbe+NFeqlAiT0ZHWirrHVLgAX59W5W/OoRlwEza0e
jgAoUvB+STbRCc5LrnJTB+e+O8Esufga8zhypkfLEw+HWVIEQ9yZaocvFq8Zx8lz+Q+raJF3pdwI
YJ6cMcjJFYnc512fFaQA3r7h3PRvIdr6AWvUfem2S8kcEvx5cNbvD/fT5JLMavOCM7nlNhanPTpY
d5FFrYf5mIf2nNzed0Qzqq9zc66Wwr9G0pmrC90YKbkr4R8ETgHOav9i8480/rK/7vdhucD5f1E8
CInXGBJzocStc/axzQnVcUtkEifsYT6u8ZtnpUhuZeAoqo52WkgoBWm7u4G23iOaVdDuSnhZ7fA5
o/UtvHqWYHZ2MijOOAnqGoEW9ImTnAVOeZX59BamZBRC0Thch7JGR1tXvtcYtobQSby1YkV4KcQo
0GI2hNXEubUwvEYswY17NE/X3LLbteQ39HCTc2m7vzTVsfaKQNhfASOQ9AA+IgRbuGRnf0pL+Y5V
vsITWrmH3saJZ40v7rOVi4OTnVdW3F8x3NMCPE1l35rZc7XKBnF0Q24WwdY3Nijcv/N/+HYDKjHg
6HBu053LgO/0pULSoDokXrnhJd3FDVdBFH9GSfNa4sL1IqTXYlQ1QaPGIuo1lF17oyAtgfR5pYFV
cPgXUS+1rly9dCKc2TYoUSnfeUveXOv5CjwB2U2ANApx0MN6BTnIrCPuUR1IOf4meLuJ95k7QZIZ
1TaDbkXPm0u5UlH3piQG/mktUmFgDydo+ZF3GgqP6UVHGyyLCfOEgQW5T//8r+d76TV5xGTOt6Dg
AGtiwH+q+7cetOLp/3jGEa5K3ASXBiPSVQOOf8FyAD4tvJlLv558rCMpv8tOy3Vzv7F6/TbrnEbd
bCcQezoQM/m/7QFmQFluodlcrU9S0FZSU3iq/ajXcy3aUbuT/+6cl1DPWGxj2HrzmBMMjn407CIc
KUow8049aofyoYawBzE/Pn2WIStoULSwZDWVHN2KKpHzgn4GACXuTkfSFS3QWj4wekFXugHMiT/o
ygCx1TDAP6cjfyqafyVizMuuU6ZWi7MTPEWCFCbScGWdEXnvpi7VMveV2VIroUmn1kuYmEJ9T3Gi
pa6feQcuFeLM4ngPSpszyeLIXECl/mltG2PuF9879/QtBXC3OtU87eYEf1rZBEwSLLHFeVD2sM5s
dq9q2svqqdBDYFuvSWkIovWoEmBpXOpCY/HFAWKQMtf6tZnjcWFVg1sqxjfMLJeLht91xxKSxuHq
HMWHtcJ1jG/tA2U2EzsuOXQHo1HVyAS2DTJfoPRyXrwsOTGjrf22JTe1zOSVqXG5aUIcatMLViBu
YGFQv50e0ndv5emG3Mrid0sttoZKAUppZoedulQa6u56uSCO1xnZPa0e09oMswBh1sC4UIVFQpg6
nX2jPOcpdtDlRBVfzoBsyNuVsfroISoXxIHohOwyzlKNFwNKBMMSPvxcyNyu8xXZA/cpqh0f/EJH
ZgsI98GPd/yiyPjvCQIrA4Q1CU4tZMkmrJctOxlriwiU/WtnbziMJPIj13lktiIgy1Az2ZJyGW8K
CdRIry8R3pLC6j7A1dPBaf8RQwkKnjwDbdovAAAttIx4i7c1YCzyP3lT83lgPorPdlyVZS3xLv/E
hDuvMqL/8CwmF9bCk27dIqZU10goEMMFgr+DetER67u/oUXrRYUxU4Du9ofjjY5gkOpzM5pOw1x7
s5uT7cCUM1wXJ2G0o4LIki347tlq1dKhosFZ7wpGxAa/vwDPlU/FzA0Gnrio+UckjMq6VcDJGgoE
GTOrYoEZIkeQVsb0z7SDhSjbJy8Bw7fk4V4T6//A+O38GuLzI13rd0bmBVkIrJDR4mnJ6abudDGk
7YLpWHSvRJYKDFtI7/SmJBu3Dr/hTKcXuR425j7H16emRxFf3wVe8s0dFJPGaFFNmFyxGirQKkJ0
dbD73UuqNlwBxZQdaufAZZf/AVnzFAevrVmBel1NKVq99vu3CzwcQ/VJg4AUglXkE9NLVOPLPAAz
1JQqgLTw4RE9V7Ht1Gy7K8zM9Y1m20VzDTqRrcsmGZPZjEeTXEn00fNrgfx/kI43s4IVuGym4aWl
KPsh/dMk5eFzmsqR9bizuZwgBzUkysQRO+gcRi9xNGlM+SgX4mJ7YLLnArscTCqWGdHJKJtv6KVn
vdygu16ZYRtMgxQp5iPFrlyA7YqPtB47AXZy3u1ZHLJyUfqne10npCJcYezWPULETQBveEGIAxZ3
Gu95E2iNNhv7+tKs6dnuvdPQe+nQA9qcmFQGJc9zJ1XJqRZuDZlWzZRklkJYfD0hhcIGJZ6qsPnh
yuO38YREvMlTNOHnNlY9iyU5aoP8aifWqpisKJ5c1oKju31SscmZHgRobPiEVZBpVuXMCRBAlm2H
uvPp8Zzre1Qpq+PrfGymLugTb+McgeH/wGjX9tXtxd1G+6ok2bXS4gBD7sztnoi3UIDj0uViyg6/
OhgRY9qjhCAxMsghj9aHOYB2IDMhkZXbMx4cncUsrqtn5eSh4k3CPc38OvNrg1Ly/KI9Q18zqhKe
agyBhTM6maz/w6+grzJHEhATJNm86JvIYB08Fee/efarzxVvX/g2YTZY07jsk2jqAqoVCBw3JD2O
7iNGjhELYlkG2S5p+yX7l36KoEFmx6n8o3j4/5WfbeT7DCGpG44dQ7uUTFGA3fyG638hCgUDL5C3
L2Nq69/gETT2Ntw5X209+prbY6UsW4bZ04DYUSRvbjVQEgclPTjRFLUIkEWPtwsqsUW5m52pCpwH
5zQmxl2ZbFdRVsy9v8DF3hnPDCtmVBPbMxs/EIgsVDdpo4SPsg6IBMAMrFP0VnFE4ia0m9metiZZ
8dVWtioKVVHSwtcraswa2d1biZ7oRylTMWkp7otPhFb7vbEDiADPcwjxVD4CErz2+aIq/cKo/ooQ
9JI0zHaV9xi9GHcWaCq7ODMsugfXmCjuwIpHr6YLLX+ZQL7bRpNlW9xT5H0WvngRSni0Tbzh0xE3
q+ziofX+bXJ1ZYHGYDJmdRIZRv54xv/ndZCpDER1p8/Mdh0XHDjZx0RiTDg1lU/2NxiRiXABoxaK
wZBi3iWlDlL/9TEBASmI1EKWm/39JO4fFddQpfBhmk0If1/ZA/btUeuEh7gO2nUKm+jNHLMXpVKf
xBYzuqIBCqXOCPF8LTYlGxkb48VcCdszvcFPrbqdnqBZfectKyg2uLJIulYiy4vz9Xzy0TIBAg5S
9NLlK/EiEibQNnmA4EpQDZskDwbokr8VY/7ZHfPiotisiMZzu3l7+u7ZIm+xlca1tJh5J3YOIkgK
e9d4RcK7Zs52td+u8VkhRC+673GYRYNObtv56nPmVm9gURNwSYyRzdxpmCFjT1vlNc5nBqOe7WYb
7nE+c5Ih8dyZgThunr8IajrNbu5oXyz0Fv8P4+xEVVZfrdkQJrrDeZ1ZZ+5ETPhNUDUMjBiC31Wa
HXYOeGcnMj2m8jb0C8rKBcXFSTCOS/dqnoGaF6ZUsNoO/Eo1/5Cz2n1yrxj0grFTqmHJLSiy1Jw4
qYGwPRdFcIMO7Sotd2aVKluS6usjQXJl5kkJRzy1wXr/C2IVzWz9yZKLsdMgms1bsi5L0BxXfuE5
PGLR2g5QydqplAkNiaum+fpo1BYVi1kFdiUb+5IkH5I/IeIgB/A1Nb9yyCtWTsAMgZ0FTn15UMCe
uKUFep7zNishJaJr8c1nueIrXQxdbUF34ljKLD2aqxa3UiPOmtS2esXbrbOAekbpY9SmH/9A0g+s
Hf0hknitX5qtFEcAal8Nk+K0R4s9sO1p/bcMb4eAaA3iJo+XuVEnyrWdg1/7PvsWTMTGp/IG441m
lYbJdytIHyOS3fNA5SsgV3LTeuk+QJOqOtRTiq6d15pdNaBZCMgsdnSVgZJojrNBglRdrW4Q9xlj
gMz4Hmthtr8SE34AknSjcnXmpMqPKzQv7u2WXkEhGsOk8RvkGdCnL0Ym40H1dZsNCkB18PEsBWyN
ydKIN4wLlLuhUiDSYXBK7pbKgZvq41dfYLKc2w7P+Db1/4U5YDh9myQc/6NyTA1UDODBbWD6R64k
RpjH9tuVtrJTCYWs/sQylApmPR0LQDRbMdcJ0PVnMOv905uWodXdZZrzwG+PHXGC77inSA+Apc8T
r9Nt7jSC7FHHM+KVEQE+ILrLs5tGCzwSo9isYLW72tPnGY5LhXrCfZ773+a5eoW20iqTB2p5Faj0
2Vqj8+Cre0mO7BAEbQMICHAvft5kO4ye9rEuSKxgx/VG9Qala5PnRU1PlEP3BGQ9fkbbbNp6F4jv
cBFyRt991qd3jII4x+OBnnPjYJ8SY7IRYVs1+eaQ6zVOsBVIs7gUGRqoVvTz/wIBcY74FU22mQFV
t1zMY4SwfvPAPJ5P6Di1ukm9FR2LxGeg7tJhVGWfqKnrAqKE+bUuva11fzlCknYe3RLpHvgltH+V
dADwA3WpO21aJY5UufCdIx7givezILgAYm5EGUSPBAuV8UrMOtQBY64CC+oPmlVlfd9yUY8PiGyl
QuhfqBmrNvT2kxRIXHMscYeP8r5fT7FLnRusP93ECC6MKTrczRFo9+0zcOKy89kWj+djTTmVAP5m
kHcCTL5/XswBIq8lyghswPOPiGnGNuk0QAIOiFdOBJGczWE6I0xjEm0UqJWY60gZvB+4NFsBR+HI
xjdHCYOXmnyQ+2XBuRPMpylOZaZW1uNZdwmVx2R3sMKkoj0fYVp7bzGvhitxiQ4mWrQqh9Cxw/sU
LMCPojC8JiXMBjfP+oZa2vw05jwy+WS/v59dvBXJcdua8mXAa/5PJVf360C9reMlgWXeZV1z20Nb
/91LN+3meBa4QmUOk3wBrSF61iW5dPFFBPPxjvDsCj4amO+eP2FugdR/qi7G21Oc5J+MhNC+cqwF
OIt4c93UHklPHTdqsTqTuHH4A9uwfTFOSq7JW7uyXUAFHJz5+R1dsnqfj1my7Z8FcobcRKZxbdUs
BGo45F85M/Jx8i0SP8pKR9pmBC3TtoNb8ChB8nLQgHucmAdWoxl66ygSNA/0CrZzyL4vR/23NF/1
2P1ip7U9/rV3pWdzpd1nSGE11V4kQ3Wvu2nDz4td9l012lHgXamnr2W5JnPxZMz+rom3B9+Khpbu
8QSF1F0F9+Gm0XmDYqmJFRLCv5NIaywZDuO9jBP3Hh1XqOxZ9qV7LfyWgYb3LGatKEKk2X/Eqa/C
tyZrpTXvgoxYqcwI0vRmsn6ysR3KpZSQhZVx2CrIF645yusdJ2ay0ARDkZxnQuzlL4BuQCR08G7T
AYOt40Nbs+H6NtuPtXsQ4EV+wrkoP8vjotfTn/jh6smgRvmZd5XII5X4XvpVQQhSIDwMPsIc+vtK
WMrn4hYUtNuCvrpsHYdSPCYpV1QOcZEBBi8QJ5zoG8rq9YQaNJ/7dkoWjphqDN+yIVaDw7m8DpRZ
ZFF3aQaLMVsgHjLXPgpY78BJ+CZtJeKTZgVSOcHq6XCC4I66PuoDae1nAjfgx7hl/aa/5x59AhCA
jkIaoro4AQv2KZJgO+OxOZV217627nv8eLx8V9+gb0Z0wLTHsjFGZsQ8zjOw9N3PYGt3D5hlbqTc
F+J1uq1II6d5M21tUr2tmeqH8VURBM5wXMUVjXzNap8Z1xxekF5VBivJGVfpmOlM25tj5Y8N4ZLV
z7B8ugtB8YxBbmhrxwLM4OZYsx5bplCbdXo0mlOoP/21LPqIqk3wk64TT17Jgf6C24o+I0A12nRT
Be4h7autrzJVVxF4RQHGLkJIVH4iB+4rQRuaLfr5yEN7jMKQCkVrRl2nXT6ADFO+G3xnITYhwThB
jxIrTcImmX1iJ1W09Cw5OCFz7BKTYq62AbPsU6AAwukQFdph1M6GGgnDpM/zwJ4PXWh3jMKmFQfN
M129LDMiE2CjTMvmx49STRtrZSA4jDb9ANOQUWtF1Nxyz2XdUINISnZstWsE0ffyBYri26kOIJEv
Q3AlenDuxvYkwKTNVA2GmT5BToiQtZLJYdk1xNOhmB9w4twWUa3+OLnV1eQtcHYEIi7pan2fRb7G
2llo+6vJea71ek3CN1/RfWqcC+BslfJAwiWeKvYBYtRs8PvT2BC8zKLid79jOl2wopJcEmJaF4l1
vEj2jx7H6v2L9Ggfr4NNa/aNiKUWoH/ZvuMpHvCEfNr99FdXESlwkRxKgrTY2Yd4auSQVQDsl6TP
IPBxCiap4WmBBvry+UoCm8M/vIez487S2e2Y+psWhsFQ5iDMLRdYANuR3WbSgDtxA6WbbFSlOqE6
zsV1gDr29d6/pC+vMN1F6fv8XIx9J/05FsYkEA0kT4nYcwuRNpKnjlVw4TJBHRaJQd5u08PnHXH/
prAt+5b91uMd2b/tS9U6+inlHOsz03Q0JfR+A8PSY4Pnb13EHRWBxXVVKqI82U34tawIXBgMNbQh
HCUZ8T264fIsHfoD9Hy2hIwgcEy82Qc1wot8b4ms6w1GIjzdwak5g0I7HQPYJEBLTPcvb4Q37JeZ
eU39g3nsDdX5dN8+MFz/SlH3AMhAYpicDYPYQuiP9rIAUN91pBpFiHmqOXZJj0Ldz9n0v9aYe0uh
nhiLA1AJtHG4J2Sw1VZHWLO6YrwC86zJlcn30VvQib07beDFtmjr070GvY5IeQG1y+9rLBh5RELM
UmWFBQQZTEF8h+3vjioGe0jwFVrTCDeafklKGiOzhVf1whLTscfL8IetimxCB9DQoZ2NP3Wr2uQj
UqCB+YnwkVVebWeqTNGTYIQWgYcr2NuAi8VmDkthrhy40Ng2Y8FN2hYjj6v0CfPPh6CKYcXu2Wwv
me9CvnugDOHaU0a3obcVa4Ld8b5DyJkVI+xHtRmYTOY9cQCkwScZ78eR9srdTLvW2RP4dhb5CGy0
hJV+fdxTVtt07jW/eGkBL+wyiBjiRMtGGytYh9Z4PgontVGdye4eCUJELesmH+iWd6ZXqDav2IN3
qNRMIDkyqoU7RtANyOeKmdc0l2l6XcVeYwa1IXnrgJXLsbfzakuCTG3DoQDT6EhdHaDP04A3sj1B
3zMOOvzSGsQqMR8OUSeT9fc/WaRpYF7zxTAUH+lWUZZZo4UGOHk2Houv+rx0wUg5utWIBsc+4JIl
suV5Z58E730U90euReOu+i4myX5V/SBRCoJL8aXD7SZEEmnnjDHgQN2RrbwmPD4/32HUG6u/PHxR
szUJ7H05TZLhFVIxr6TdxPd7rrrR+Y5NlyNR4TdgG+iDpItgPBMMCefheDmecfHfvnZ9x/QkDs/J
GB6jSOSxNu8GpcBRi2sdxcQ6fvGhKmC3b+L03rGVX0+7/rZJDiIgVB0eRcPuKL70slOTID2R1JE4
Td7g9u5V9RfgRe4ZP31eb13n3HScrcV3zAqz0dn7KlIfabhfW7lwEyPeggAfANsmQB7lmAWnKcYY
R4UjqdUoGcFcCE44SP9s1gB+wa0Rg14IIOsUYMUQgN13RnUR2b0mb5Ay1NDSfU1/xmzaD6miCg5B
vyCQSSTzLdRLtji89ksDffgDQQbDTWaMJtcF8zdRmVzqTlaHJ9rcJ/3NTUb13av5uS+OE5cRNj/B
fipzh8mo2gPpvU2v2uQMYIRn/6bRtZQoCUput0NHEC1E39brl6xYk64auRQR+JepFZQThidGTN6+
kKqNaXDJym2/G+dSyo1oK0BOt3RcEOkYTs3oH61qKyDLrn9Kcc07PSKNDJXtfFI/IUbHfdX/Cw7c
YDNahSZ8vSu6zQNFZ77BprARGGWdEFgS9B9k8xgS8J+WTwmLbYPB5IBx+erQlK2eOHeeJy4EWzA2
EUedmygHMC9NXRlNFKMsfUuXTApVnXEM8vaxP8WyZXsz2s4reniBy+airOM6EZOJMMIor8J62x0L
KIwlLp4A6qZ6+wGDzsZ4V66d53ukmjy6tsvZenk+0A1QaUkb0KIP6gTvrbK0AC2XLKoQjHM/Cm60
xH0OuXH+uVJjjo1MlEab5EStvgBWgFw6thmbzTj2nJtv1rYLIakhusF96lb4FB+m6o1bDeJd3zSo
O79WfOVy73+nFSp+TiyEl2TarXcw9vvVYANFauAvwQuAWVjGzKAvHzLdkKBKvi/L7QtMlAozRRq+
6ijrKyRpk0iughD3qgrW8YEIJ7A9EOkLX3AmItk3KrEyMPc4ztOFWQn8eXjvOr+X1IDKmS+WPElA
InZT20u90MNXq0v6hUbYn0LIYw/H5PfRQJjxeaQC/aBVUrmtnsjv+oeG0fWo7LVEvtevTaUV4CBd
awkSLClkFFIGb2MqPqnvprrcPagYpELgr3ocroplVWjKg5GPiF0qqLnWC5WOUTRNSBn6XW5lRqSq
Zd9IgT/ETASOczRgROGAMseKtwYGn3bRu79rUd3Zk0nkskFpXjsZb3YqAVHOCnjboGECjECZ/gWm
d9oUY+bzzYB3OYlRE7251XR0Geclp55QKerHwk4+Gh4bkbOdSDmTvVwu+aL3QC8U2QR+T+IE3B0d
TdBRu4cvGgxjH5IGauty9FnSU8TMpAreoMhZsxpX3N1UIUm21bW11N7X0Q1d4E3z8qTDwnL9pN3n
gmxl88qG4TQ7WyUToB/TTh6a0+QwVM3YoLLyUlhTvHZSh6xM7hctwyENmgLnYWLL7D9WoSfIT4an
prTB/FqE+EC3mhM63Lxh6HxPGy/tjzhNyVKQ/vgyjDoOb2szrlZmSensMiorukif7x7qZ2+5mFas
Igz8jLabdahyrYoWzsSPaWnReBrkgMspz1HvBzEZkUSX3Kg6Xf+HA37YbogxFiXQYJTeeMDRoX0U
l//bqgnlcyUU+gKc9TiScc2e6J6z4DOfOdr1Qw5Ymtxni1WoDA0DomSvGmd19Zl3cCz6J3LDWvY1
BR/goXmssFnqanTyxDY+AEYMlbcJn7I/KJFSUAEhscP+zX7/BzWuG0lv4/zHdpyPtRl9X3RWYxtu
1BTLPgspQ/aHKI/x7cD8hjeG81N/xczaT4JTjvNnOJW9a/7QUeKBppOgZpOqfsMZ6pyhRP0ifvui
j2NPxCoV3scQ6s/eOC/CYDYKSS/Cs+g8FWTh57+YOzJukyw3px8rhKeCF4lRYqzrBpwnlUlLmqM+
9EoFJpgUfeg6sGxZmf4vDagg1zWU1GOkj51Bth+eW054aWh7prxcSSJMwa+rsnRf3ILW/yOCPZ0p
50vO8gaZCwnQ+YUEQ4JlJRh5GB4kooE4K1wNK6UoXcRHgRp3rE/EST78Y3nd3qMBwGT42s7z4Zg3
duKU7gGgaaAG0hhdSDEORA6SvmXgeAsj8OjBVDd5yIdAZfZrkdMe5LpeQUqUXt7kXRek7yzxcESh
5yauKNAvoupDJYPC4wHGYN/G6PYpD9/dol0PeZKi+U0JBQABG+5HoYa2mXA0IG5UslCQSLswvvuf
/BP8X6U9mJsN9iZInhhy53TNi5+ppxGiMs5lFVE8y3DPSERauBBWzFw+AZnWEwwSp23ihZmlxMsj
uknLfPV3lQngJuyqpFmOYPC0Q5cikHHzvKTiisa37pZ0Do01S9m1rxT4t6RXAXkkI+/QM698maMk
GuHsJjP3oJhD3GRmrxu3ErnV6r3ArVzQfAYTUlFWCT5wwLECJlTaeyJTZ9GLT6k5tony5z72gmum
DfB4bnDHFKM27ui9hpeNOnL27YfPlkiUmTmH/3ovwnx3RGLfIJeFaxtrG13zfLCDhLTKzXKfdbQY
r2GXvAvxD/kiX4AchcnA6S1qgiJHRWYctJOR9Rvs6bQn2iuW4yw39TAkpfJg5fmIOsteFc8aUQyj
mv3tCVIFMnF9oJmGWlTAQtmfmmf8qX8oNAox3f27x4qlgq//5CR4l1yk+NI1tHYBZzmmeZssuVb8
ASpsV3rPdqUQ22AHv9j7q7pIJwpNVvRIusik7E8ldxOrBGlg+MMWcxTfD99V8xNu3qvwote+NQYc
K5whPisoQbL2gZxYNkpnYGhYzusFF2NmUG4VUFfP03JW9MUks5Hl+14stYR4IaD0psXCPwCkbNDm
KlldoZl+FrcQZ7N4LLSUfUgr6U0XJ4CL8fVyni5AcFVhuC58yj81KZU8ZqpsrkwZyAQksLYs31ef
ApM/WESx2o7xJF04O/u+4WIpGzS8Sd+bQcZxpgvqCnWaTMiZqc3hb8B+plEnxrGQRquQezDCMAXv
w/ey0CQZTa7Mq9GWknn1sCpLpbyMZGKlVxq9ZF78ZGoE11bl/APUTk79HFp5P2xdx/sEXOKIuhya
8LgG1Fi80Pv/zkCRESfmkiDwew8UhR4Gd3L0VGd1E20kZlBo2Z9EXDdxn7xaDext0mp2xFsBE0Ww
nwck73/EWWwjzjBTys/J3ukDoX5egYTPZoD0y5EIz8F5pWfkNWBLPr4bQOpJo7yIKlRmNfkYwaet
mFvDgdrxckIg6GfYxW409Nz8ym0wzz1kaF8TiCD4tevRA/JARXfcExScnoIrz4EO5cV9yLtArMBm
QVtV1iAYdzuJL6vZ1dLFjWEyXt9cUozVXabC5/IaIHKQqyxz3tk+C3u3+UgoHsq7qmm+9r7Ti060
eYTzsoiHBUon7TMj+erNRkOBwVnw5EUvBR7/eyTPn4P0w91uK9FgklNwSQx2JOYip/jVRTxG1e1M
fZLjZb0ld1E3Pp8/qzIupW/1adfBT6qNEdNRAZwh8HrO2SNu708tD7QqBp3t38tCJHZC2znLJPBb
oSxyHG/5LnoCA4yhjqOGirCz9iCMpme9Ld7z4vuA8Kq3BQ75gZLPJS4f4xk6z39VUFPXYSX1AYtY
IkNDctJcr4VeG4WUPdUzt9ynfWLIEQ3LnjphDxcTRtkbO1M93k2xe92fNDJ6AAVi8pwQhz+HcXZH
pYO0IqdYAggkQqtBydGmNHEDYG5YHyQRK2cM0pxqaAx4R8X0kuy/9QwR4Yt4FvLinrsxP5H79/rr
A/FIgmma7/Yp9Iz+YfAWfs9Tai5o9fA1JsQcmUhj5We3tkgBsRFWgIWu78wopjNcFB7nRtNzTDeU
CwLnNAxt/o6qm1rCF4lxnEQRppawuv9PCZceB2zk9OjoqKsJZkd+VWNaCRptm5Rpx0fwLd/dYc1S
LhbO+gm/vITr7mRU86lLd0rtZbXarsJKd+dj7zb0Rm+2HgPbqR4hQqhPP9UHBfnFINok159j0aZG
f9qxKrkWErLaO3FRFlXwrmdECRBhHjVbpMcUss1hx6PgGNRpRMUIscwoj2hR/6PstQ7GLfXMUfQy
LTO/mWwZOdYxk4+9QsJrReuv7/n6ntlsqm8FHBa0AuKo7zzieOHjLrVBTNotfQGtGHtKF4YaTOP9
AObAErOF6LAPKbqO558wouKoCWHxSM3ugFM3E9GwwgTKtfdIG1ZjErzjE0Qg/0tVmVHoSJBJQSQz
ElRqRIBXmAsIL61VdxjDgoccRAj4GJJWfwbnJHPRSc0HKJcDvrkH8Kb1L/qKaP8bZ2ihJoV1W9v9
trH5XePGExduxla4l3wgsvhNbnHMNko6+6h3WxM6TVXCCr/VVWGc0mfk20728hsYBgthPpGwSLYk
USpWD7AsvSNErZGEgWAVppfqnERKLVOpFZXChFQak8Iaeqyx7EWJxfRvntRlRSMB0mHsh4Nk7hAd
PrcvEmXrKVfWl9pGD1uIaxjg8LBu/WUFbOGreIZo7srpLru803iWEAtuqtCKOdQdEhowzYx6YVZ5
uflbLBr0auTQ4JM2+pDVL0TduYwX5Lj6FPR9Y3Vkf34iOluAmD85S62Qibi5hVWgxYz5ZorXqjkO
ioS4D7h+sPkrwGcruue3IBikcvEhf4Kgh6RaYDmeG++iuTITtvFibN5JIgN/dUJxcm1AFhhPYEt5
ElZRL8DeSYGUZBOKQD9ZG+NgPqmXg2SDh3IxjBWEs2QfVuKHv6Cx72lTg/a8ANuBqxdrVFOQjVlt
e02MPfO9i7zEuAA6Lkbh0IE5tZRexQ5cUcwwDmKrFHy1HwUGZcCT3G841CmNw1AGZisC6OVMK00u
IlCEqKzUR8BGF4Kvj0CSF5lvaEB7sFRjSOuOq5Hbi6PRDuUzA14aW+m8uGOAIdt0V5umNC7rGWf+
ay8prFQFscMdURYfxmdWXRpvCkEZrxSVy8Cfxd3M45pzeZ4vgPA448qeqtuMN1m12Vr/qKr6Ns4z
flNrzzHmsyf3B61uWpZl9HOJU+ySSnTYtusVQA4p55DyheOhIYXgTZkkMvPfkBogogoY0d7gmlzF
fGBcvGW+j+Fav373ZbFw17meUxerddFATW5Zu8HNEbMU5Yz4LAeCLdQOqhdwDGH54gg4QauhUc4Y
/sVJQnVuudjzcYQ2RU/XNaWJdZmuP9Di7z59xwgzHMrH1QxLwU1QXfPXlFWB2h99BGT2hmghUnGi
I7paBUanx/qwgHL+UYRq7GfCWutZVJx7mpOg8CuFaDQ45PsXTnx7uio2rHiKCW4To7CWTHYR5plG
wAarAEbKaUB8VN+dXehuiHokTuYCrCzDidomou4lsipPLt6zPYzgMo0tmmEmHORMWo0DfwJCiUSk
A7oDoOX6sTjigPOmZxFMzaCpjK6kyTrS7redbgPYj/edH+CKSZPNGN+6y9cBs+hdpssOkK7OwRq9
wp47lAd2QiyxsU40/jjqptiHUR1Xtw/arp6bW8ObrJngF44C0wnGXFf16tKwOQioXfT6EaEcJ5kM
TYVUy/r0LDdYkVbmMmzryoeLUiD5KQDChxcW409ZILkoKu4JUPakOEAE2Hsv+PUL73YWAORCTEW1
NHTJQD8F3Pav6Ut4+N3AIy4CL5D4K36FHfte36JMRtbSydM5Vy7NeerCq9LtrDrWRPq9MTuQjEi1
0hyvUEWxAKurdtbbUzmbkS1t/tqX2qW6sKFcYwrUJ5eKK8Fp10sIB5tgfKQ6v133s22QkZljpMC/
blg80g+NYQ0wzGQdYHzjmU6NnueNAa21AbXHhD9lHpU5u/hU3S+tMuH+6oapvYXOoc1XDNnVqFmy
Bn+phbzi+pDCFIJjczR9RmHz7Or3Pw1qX1GCrhSozUzlzZ+jUWT5IAfsF6nqCQfXzq1v6IIqyZLW
xutCgrms7mBPGeSkvdaakSUwp688UyY4SEG7Tyy7J2J4MpDIHIxZajspAaVR+nNQsLX8bzbkFpVB
GiCSuvjyq2Yz/fO/NwO7y6mzlfX2GGroaNy+W0am+1M1hqtoQDR0M5eKg8jxZMrsBiofZeVotau7
4E6UgKVKprUCHG1/Tz9tmkydQ6G04JzWnWWWSY6jFHje9penwtOOFICTt/mkzVP4fIfHsLKSMesr
3IZtclzXlh6i3NHzJMohdrXafL1DPoWP+jEMcjn1WPE9WZF3EW/bWo48IKn8tcIbE9WDeCUAZTDY
HOsVkbk90A9FMfaPjD/8zkxeS6P8xqNZsDVpMQPix8BFOuuhjrI6CQeVAYgeTCwUejXD8fpGeycY
chxfBD0Rjt3618xzLlqdm3mpbENYKMvifhnKgnGk0YEryKmV+/yAWITqAJtluQdeA+gK7wA0MEr6
ub0vzVnVsIzaFJSdgRmk43IeY28u5/1k2PJHTSWJJ9Jl4gWpP07kAEucFLder1T6LHqtErgLjzMn
N5e/zCAcjeUiN1cC3k/Z9L8iMicwEixqteutDpyZE1u2NMRgtyqHq/h8i1FaKYpIf/bg64v/oUdQ
QtYyiL8VV+TTzCYXa81rYJFBq3KyyYLxFMiNxkKRIaAskavbEFCQl2kwTtQr5oA+WyO+T/TXvXVb
y4/6jIJxq/srmvBK147PWc2QwvSyFjImOvF4H92SAinDvBdyTGxPGOgL4I9+rV11DxxaqF6X+i/M
7JUuQPGb5y0awe8nJL5CbNcVWiNJKrRp9b2XxH/mZhzJCrHIfeLZN+LBGa7952IqYn8387nveYYJ
Knm7S5XcYiJwwVi363sijOl1V2/ohTJUh+PRRi0DMj9VTwfZocSxuUeaJVekWA4U5FJn3v8FFaJG
SuL73aruDaqRCeIl51UwHFV7xU4hPaAmTP5O6N0fsWSsyrfBe83FyZc4y5TtWUDoFxH6ifBHg/yf
ly1Dwg7I2IlIz3gAX9j2IZG86flQCjts9P44taD9eSZjaTWe80UMbPggbSWW1iSKvGOvtKNPIxkH
ezXxLfiPxPX8ankzMDJVYV90bTrdcM7l0X6vIqI76J1Sb56LtKjh7eKGFghoRdTBUpT80FPFOEVy
voBlL9Qkhk4D2D+di5iHXRQ5ceeHgYerfhLA/OE85B3NYAHxjc6VDeWyjAfBqIEuhzzpGJGDbQe2
4WegtkP/wUYOQliXcKpQ8z5NoadLF39xbX66lYkLxnboV/l1cVWN89N//CyBDiAfNDE21TrcbHSJ
SaAScnTfnbfz79ZrgL1bzmGp3RdUDBONkLB20LOdp+kj7tYSjvklEPlJ7FagaYsawlDSoAQOnWNl
+IV/7uKoDoIAHN9rukHjnS2/JXRCkLt2dyId9NZpur/0eQhXu2HnQqONEIn3cbL3bneFyjQQnEiK
PU7745HQuzRCwyuIpZkSH3J4Gaq4TeAK2B3zN+22MgQF4dw34IeeNNYTsqWuT550gIUt3Vfjq2Pq
80GDl8nDRWNXSTnidMmSgu+bey/SQzpC8JSspH5lrrv8f4NTe7sm4yMnEGbYy++0HIjMBlCGpq78
z/wT9bp7txwGdg09uEWRZ19z9dg1u6dCRikA6Vu5aMTdAeE/dA/eOD3ANEqAGvW9UlmK/ncq3rly
FfgokKPdv8c11gzaIc+tVbiaHl5dU9OvF0D6jG9TCZzqeXyF4FaDXd55RM2vkj1XTUb1UnqDEYIV
wMeJzXyqgOM4zhLWGSHuO5NhJEz1K7NUayTj/XQNX5OSaeFNnc6vo0NxiC4sOEok5dVbKZoczLEy
ACt3bJ0smmSkrFG/WLG251DIQ1v0RBl4VDHyRI0V0OzIOTwGQQ5F6zEfJjS41+vVDrOhZ+UAfJcw
Y7+o+nyuubhdgDrzQNCrcaQzStVrYqRzH0xkZ4L53dnYhs66uROrhlYYys73uoJECHJklJcy3YRz
LbbUbrgdyJaPSPs4Uoh6fyiPYrt1YoW9w+PJXjJi0beoZu1nKZd4G7RzyR/mecMRwpjRYuIq/xRC
YpU0w8tuZtyYdsV7KUJQ8Ng4MFJeA2FGmerUPgBmiC96yyM4eMHw6RFf3r1IL55/AUmGw6ITJjfb
v5El9fPJm+KnB9XkSUH3gzaKV4gGasiHI7UO6Hc4TN1+zy3kXtw6hpVnK4+IEpi5iWoj8pTqCaun
dr3MBJIQmMsbXicvj8jrNjbRu3hwze8kyJwlpCSU+FH7SEEyz8c2mcDncx+ckenBwlXEwZLbucKF
zPP6o4/oce2rfhQ2vDGTcm5atRIKGGj4DFtQ/yAV7rjFq8OE1c2cd/Cog7Z1mPrpIBvOd114M0UI
TLo542AuJ51A4lMBhTO/NM/ttteDqvo/uUKSzBMVrNQgP/ibXlcUBdXR69ub9uKeOcIpaHB9vZz7
O88g6oQn+s+Km6w+OCKilIjFe1G1ogSypQDUz4flSy1/UtTc6qJ0fSeVtyja7uNiHcGTfS+/J//p
IAxUTxY7HAbiPQD1kEnSX4eUDRFRKJxlxuy4/OWv1+vUGeHLFKIMbRAqCxNFxKBV8ZGhUw1+Sliq
y0LEWmc5BOjwX/pO+bszCnApED4A1oVJtW4kD8KFOJr4eBCWTaBNPEVXCS0IXLw0htwuvp2t+C8z
kGx9SnAKBh5XozvpBJWlivmH6KGfATi59abp4Z2ZcaR8fzhZvZ0jPoMCR1ulDGglbd4q2OsFD/xo
DmkjgXSrdO7SWzLVE6bWRtXJScfs359y/KnIWz/wDvIJf9RuWru+08Cv2X+A2SDBT1sG3+bsmPyb
qe3fkFOLaa+mvhqNPFlx7U2UvujcajcxtX2Ov/ciKqs5n3rVgu4HtVnzRwSUjNx/uV8DWntDcYpQ
DU8bFadf5SrfRPjjTnqvpQ3koMNY7XvD3UXlQYoPuQlC64VokFw3WBBA9A2DvSQdVszQIzMjj+06
mcxyWGKDNd1ahlJiCz4YezU1Iyvxa26nPLHY/isumZJABb6z5ijwIN1uXgxfIrG/joRcMMYFWPaH
G2r15V1zA4dB0bYCyZHLRTFi7939opfXuUXk1PT4N6VPDosUVAIXe9ETsiZa7tzEeRv2Sc8Liw1d
SOJx2PilXe+hsPQcwWR/XEzCKTDoLbdy0DLb6H0RoEAIdGeCtqA5vSCkYAwRH+9//IIvG0Tn0825
fGeJ5XW75me6WQ1w++AVm38cVmqPIAcDsfvwLHMJ7z3dPHj1VI6fVJj5eNkUWneQBswWxLqrCanu
0CyuEcY56i0zvDOcFO1m819YJiugZ3Q7ZUcmjLGlgq3QMfeOHSCfBqYX5d8TC3eos1pnOu5RS+qt
m76b5Me1OmvXRf9hsywiZ5ZhzVEaWQOERbFcKo4X5gzjxrmNafwFOGTjcU+gsGSSLtgCH4ljlA+q
HGH/Y+lTEERDwmSO7UeULkaJQ2Z/eP2ygJe203DXiVIGQaJy9zvqgZMttyoWYHh826Mr3mF8Up5+
L3WEk3d38Oo4oVuqevqgHlFx6fCWfMijw013cr++RBqiSChqy1h7Dfz6e+tAZ84q1YP0/8ZouifX
q+ZPjCOnYx4+FFn5KRLlbGQ00FodpWPWvHBkql95znOJ3l+SVsvL1FJCmqGFqN9s/l0U2kNW2e2X
hwZyTmap7Enb808IeBogd7023CUu2pv1/MuMAszwITXYPzKnsCc6u4V4vhYn/PEZ2sZpW1nGEBmM
n8QrZ4SRwWwWJbN+CAlCmylwuuZ0WXwyvCN41PZ1bIr24ld4mfP2GDH23ftNJKsRSgnZXDq6tJE6
32cyQYObOwgZ3p/17zYj1tXOcoABRIn5jM/M4CCvK3Rza0wGF3Y2IZ+QXBW0Ph9nC70KplRxJ7OW
F3RvPFn9NMEe6rumgy5ExAtlNDRP+NNcYUP8jBLrE+K22vYkC8CbEhCUqbHZnns75VpdsBtHyGNd
i/8fDSM06mmUJsTgF0YMi+FmYm0zRqsToUmrm2IkbIxe1zthq5zioojBwCXdMCRBfa8Ghm23k/wH
WQmuIGnmZiCjQjfWodFjxxyDxlPlnYnejroHCSXENav5BP5FQRHJHjKkOU0ffc/ZURlWryZIFCrx
ekvGmSnYc5wtIvGSMSBlU4GuzKrsTm1UBJ8FQWU5bxVU/pQCKQYM1awPEMe1rA+VutdlxylNsr6k
dbb+4ZBM9dccBehj550GRmlflOsSxAxlYTEVxwvsyXF0TE3AfT9n1kbXLV9BwJ0S8qKuxsYLwvuZ
BVtJj00BSenfKq8pdH1D/OrTUB+E+RoMFvEdZaSWzxKBg2ip0lxQHJwNVP+vLveRBM/jCpp7Eepn
EoECscwSSdZCORIOX6CmefynL09qBdT0Fleu5ueu3vh+Haa+kcoVx3I0G0FfjPEYjTjQqlqA968G
5f8cadhxbdl/DaqCoXso++ax6Y3C9E06HQ1jn2n9RKB9n1fxQzpoV3sV7QDIznk4Fq8CqbNhQ5/f
ptqYuv8G9TMI3gP8rWtQfQNHC+pDs7SG4Gf3T+gtKEaHLr8hST8tYO5WNJm0JpjceV3iZdOLGYxu
Tcmmh85mo3I+wUXEnhgs0fzP5jLyB9wvuWsbaSKUXG6fPS2bP9mfsEPOC0B+PF+FBRCCxO4SEnOZ
FSurq7u95GiP5QbPlFCTtb8synMKHLW8UEnNXAeOe3Zduiri2uk4fUYiF/9ShmEK4NAdcpWwQaMd
Ux0bqifs5MoN70bB4e5a5+Co8KHfEvUNOBMAhHSOxj2SvBEnNI/T9JEwivcqXrwDXZcu5UqH7GjL
RuXJmkPN7nCiIKGz2dblkmmihCdU8xYZxKxwXALvYvCD0SQYcvKKlUZraq3cXEdtF+3RbJZJHwpp
9GtLXeBRGUaY1MI+1aADRgL2sg8E1mSEbrJlnw0wZkuQuQ7WUTQOgbam6b0a+DCWcGhJ15f9o0jp
/hEat0M2XGzcicoY16fuv1JacWel0HOElq4PSbjCrWTOfuN2sGpOnlNZ71PTu/4We7aEHhjYvyrr
5jFcrJ3KQv/bzSZ0cXR6Uqokk6gqdlHS3UoyfMV6RvgqlV0NSdpN50UmSThGi2YP+KvSLP08CP16
oIyJHy2ok5cbHEVqd9faAFebS3CIUyMfNGjwDwMyMx4zVXbxczHWlekce/iFjmjslwK8bUMawjDx
OyikrXEDPT1oqp5zwjJ2RTSnP3VP+9pmScIAx9h6jKJhO0rd8Lzuehv1+EVUtStMUGQIlArjbWjK
plaeK6AQIvlmKD4py/zAEj0ovmOLPd52YrkqyyEXb+A1wRB8nXn6uZAtSG4M6pUZT6qIsoAFRLTU
HkIwjor2rmekQ6RbmhSL5vexzIKvPQe5m4Ve0MdjsolWLUiXuGDab/JZKPXEaj4D3mNMBeboGfG1
8iNumNoJPlbGJyxZtModHEys2A3d63JfNYl3pBODG4QJnTOTmy8QIoQiKbo6ZzYJGiKOkauUn8sf
qJ3s77qLyGoVoz7/ND4BAkZjt43b0RgtLgX7INJG8Dq8OcZasdWDUUOfMWxncj1tPRgHwb3WUWLc
maY4ohaC/Wj8PRWvs9Ka5pkpcs9ZSOhrX4WD/FISyOF0F8F9lPx03L4DgXkZp2dKjor6NZGxKtQq
ESEJFyXK+64n5vbuK7ewa9OvdfFGhxiDwQwIMOFgT2OSq8vWiuv8pLEVuiCs4wO782fZfsGzwuEF
1K+VGNRO7qzsWTFaB8j8c9IfdNMAlbJxzWE793HvVbzwxP6t/lAhwC26ico7RdpmJ3Tu0rhMF7qK
6COuQJC+YdjRLfG66R40SlpiQZspGXzl0ei0Nf4GB2jK3MqtNRRSZvZyevNEbXijF7OdWTjK8H+h
OuyWeEm+LT8DBnUX4UPctjKAYRtPJjQTG7ayGIgvc9J8ZMX9Pel7mM1t3cvyKiFsb40gjGQxdx8H
BJkAvIqbtnEwajY41Gr86zETX7yEm5c2ixSS6ls3TNxiCufTdbpOWohHgLqdH2LUXX+PUugtObUt
EEdv0COBKKWkid9LSD85+8kEZ0ZPwe7ToJ5fm9Uz6CUMxqMW2BxJ5XHHvvLa/+GTMtBQHRRQwGTz
56iVpGnr11v2A7nrQH6cZQRq5lrXuTojDZn7XsdHwklyR9PDrVr1eV4pQ8WcH7IIDiGTCE8sKTjR
lSvtBS9bVO1N5+8XQhnaxrjzMGMyvgvdh1nFamr989Ihdd17i9DrvBumh7vHkA4eYr/q2OO+xUMh
KVzZycJGzammCnAMWXWhf8kvJWl4GmtK0k8oQ9xgoUqaSVtDV5RTdfapRRk/JgGHyr/YX6Fgzjst
JqU2PnLtFmeNr4mMW0sp6gIG1NNsohrJCgJ3xixRTTPiMBwqcsaHKypAclq+wvpgvYut6z39COj1
5CdkSe7c4xAHxc+GRGVGVp2FoHEevL92Nn1ui4bX16MUC5iXv3aO+57xPWaNpzOAWZiZmccjunsd
vPgeSGVT6Di+uv5SlfiYWADbP6KcoSFqkVHNmdOLWhxGMcWfuzudB6kJ+goa/8vpimIPx1uOMe9w
cvKv5HN8/SgW4j++atkl7TORvm+lorgvuwzCeng6BLlgeMwi76l0ZxCt46OBVKZ49/lKJHOZvJCr
I5kvlLpwyyt54JlcwdnYCLZAIY5VYa8ExGO+kZlOx16paw/Wh3uxnmz/H5Rvuv9+kieMEY7vtS8h
cSQbJCzd5Q3zLcjCb4xowxECYPnVLAndJMQCowNfZHSms83LrORRrgJMaIwHh2+lKUmGc17F6FOl
ghqT0t5HccLw1MsoLXcZJtd83wU+nTB/mS9m+2RYYnYC+9AF+QCuvB3lJ5UcOZKYDBPY0lMDYgD1
eOPZktzz6M4SiiBKhMOhP0FLpH0G+vBc7ZVbVNZsWgDBkQO57tbyIWLDYz4/PzbGXjzq5s9MKd/8
5NK9ZYo6rqoovak0hm80bkTptFOFjcvGxZc5+Bv3Uk5aTRju9msqZ/MbSkm6/lGpYLkIPgsyF9ru
GAIxBuDvu+pN/PTdLzn+v59E4OazwAIrLvldu+b3I662D0XTqthNkQ9ysQVAEv8wpDb1kcHvEGK1
EA8qn7gDY2gUdnulcCnPUiuXA5A9CCw35B9UWI7DmFlsDMeTmg5CJHQxIty5QZpUGEu0HHD05jMu
sCQg1nqlcxbRQb7AF08ETbsGxY9zl6EnXkYYn2doWfns4lzjpIeJenE5da+5MpJoPz/G8J7FNuiu
Mrkj2Lm0Qkcx5Rvuig9FHiC3HzVTpTK1DQ78fxDP7AAp4ClBF7CzEC23JVfO+q4S244ibNBC1SaD
aLi5voJalE9aEZW7C6MtqEmwU1SutkrDiPQScCLY5L8FKk06k1qMd0+drcIoTHFfo5EPt3fIcL+g
JG9xO6pAkiL5927EQHFNdpXN+VBYbMU7eryq8KKPT+EI8nUHC8QjNkkqUh65lZX0+DHv0pCms+Cc
HkjxcQRPazXNkHWqQNJRNuTVZa2jLDlTUkf6GbxZ2dx7i9cjB2yhqwlHG4jgs/hlywj2mxfdEgcu
QJlGLpMGlCCBcNwjRYLQGAiqnS/lnu5/lUhlxYEslOY2Qgmrj3+jKRZZmbLCGYExIwdzR8ko/vif
/0DkbKAsA6lNg7JAmSauS6tv+gGPpqqYwgDXYvHWDM1ABuanotct5M0Q/zLYUiGWmQWQ46rP2k2w
cczFQx7MFh+mpNRofTLit4vxch2Cs0hC3yY9r00E20zW/KBPXWNnzTxmm8CzeNcaMAgIwnPE3DZd
9CC4Poo8Sa2MEZ9eUfMNYBlLEQf1Ezx3tQdrug0WGvB73ig1HWXMYUdOkhnWY7ZOPJmgbiKt2XPo
q8EE04FIMUqvgPSbPKobtgKK54ocsztKbnmSgr++c4zkw8ipzdC3fETqgawku2TIjsLjoznYIszl
cSSGWZdCijKzCiIEy6bydtWutph6Pe9Ql8BGC0VCKwhKlOmNnVcLouxLC2SbGZOOt+P7nOQwZtPS
ceCGZ2r7lgYqfmatsru+oub4HAHeKiYkhAqMAhe3NZ5RMQ+Cu9AwoOHimHAgm8f00b78t80buaaO
hDk6ljVW/zeSBsBaOvusFJpd9cwpTpJMhlqBSNMh6mNno/qz/kaGgKgPL8OW1G8tvQtsM1P1Zg5a
DtTNrtoD1ThcLW9UwGbxlJIoM431zGAcBtVOrwL3siJO8EUQq7JpQSGfEfepbF5QpvDKnTyKGWr7
QAvG2WyScJX+BOhhmwKxYCjWRyd8YdoD7RCKaAuUtuh13q83fOJu7G209Q5kohGy6HKzTAj36u9U
Hq0VscuYIzQ9e2zA+8+oB5J45k1DhoOn6zEwKRcn/kgUd6KuqB5JW+47WpANUmUIeVtiuMCQb6Sq
IgAJ4u5uTmI0zpCSM/S7fmpMnxET6w4S5EOQpFfdkpgEmwBvuyZvRuEBatBQRkl0+W8x6c39UQqq
fmEiBf2sFdkPaEQ4203GrFJVr92mAfrwpkoq9v8AZBJ2acP+Tft1S7n7PGM/WjgGl8MwWGo+WshN
xW09yYreaGQvJVFJOyDtXnnqJWstzTKWIBevTTcZ7y/hgAMR74REQAx7tYjqZPKEAyZWRBvS4Bd8
2jBBW7zZJEpYieJ0xS5HjNyo5cPhvBNlSNG92hG/upUCBqdPOBtS7+IAhLGjJQklRIoR53yV3ALR
o+eckakf+XMZ9jPeXX/1IJJJYSYw6snLzCkrZ2jg+k9ZcdWyE9+ArhJ4OBKKlrALSHCLzEBxEc3R
3Cb+u5qEeFWbbAZk6dLfe5Kl1UevyTYhKhNNN9YRKqeqlN5pBjUNhieA4pOtk+3ZTzr0PvLLizKS
I27LdWLq+tWD/m7nIOH7Z3IzSFSnBgXONGTEJNjFzcdZrF42tMUox+c8j4eASeWFblKSinJmfehy
cTESgCeo5RVeCl5U4Un4sv9OBnZ/TpE1caJdh6WiZE6y4GRMY5p9CZNNlZLC7KxyLpPNm5aeggk4
+NL0qkUyWv4/GG7jNm8zwwQN1RR/VlZKv9VlOaJ2lKawFj3LMRIlZeJBBeMClYwNxrMPoC0N5Orz
/6Qmk9fMzB7LKkNyg+PDueObRYx9nVJ5Yu9C/FWaKY859W2fvV0OeImWny9mtg9NvCJBRMdoSAhj
d/lVgupjXMXwHYzvYSdBKwSP5yXXxQtvcj62V9V313oHeG3C+VQV5cGDDzkNo0vJ7277TpgLWR++
i7Us9WX+reLN7lAjQPFtMSZNZEDa5VgDxareV4wrTDAmXBZGkHMcDeT3xDma00+mOYym/38qC8If
LTEKjLAngR9wiAqZn4zenr2McFYGtxNSSvrm+s3vaFdNV2RQuwM4UmVUtQg4xIj+6gzyvrxt1hBg
7AIuehO/i89XQW9GMGDOLfB6CA+5oGOFh/SlmEysYTfijM6QbZKYNHpjBQ5WP1kUOu5N44xNFZWN
fvbcVE+zHr9cwJEruden8MA49tHM8bYu41LKx+PCEB12oKR/LkkPv4/bEgmA/czJ5han4ExQiRUQ
aqeliR6GLA7gtX3duRR0NaeCHjkGQjdVcSVqy+u5mpTryWMGBcwLjRuKlwt7PoGdCjGNOiiDycrb
oP0GuQEh+4kBOwvYZr/gc6a7jNbT2aeyNWjvlevG+KJNI4dLA6jN2M3VsWInprd3tvfg5MWcRZX5
Or+kSQulco+DLPSd8G3jb0cKK78klCHUlYWJDxuMzxgfTteiu1VHXeNwsejSUX1ryYVWIqDd9nJe
8ZR/yPMg8IMBvw76FCZqxjzLvcFL5Bj1EkkpfyxgwvjpZeXAk3m5t/4DrqliUkENYa8zgkhplxCi
inuNVP+N3CHC+pm794ieUJLLh8Hy33gQdmijCnL1aTD4cIRtj4ZzdAX5aZsEoXqXgTTc8qCSdX4O
fPXpJVQdAQJU0s+c7laULqIYcf+GBSswdW+5JD7IpBzoBNapZSqluYJpw/9fKxDtYO0xKpL3jBiV
+lCtcnEEVdtcKAqIMVEcZTd5/xFcE0XRiOghZ/Weg86UF7mK5aL3djjG0I/83DgjHDtNo+JzCyT5
gJ1hNEVERs6emmwUP9zNPSrz18ya3UYC4QhviUjQUcgXJ/9j8SbdpfIIBXH0Z04EPkm9wBGeB2ON
W4BPTVoq3E8cPUA+Et1shAIL6p03lvKaQSQruTvuAs6xuiwZ8IYYU4wl6DPFlV4ryOvgamTP1HoP
kXi+A6aJGFuXzNqVvMXutqP6atfM0hL+wsTg1e1kcppgV+illCCLTToc0qYu1jGWbuKjDU/fDcdY
A9yucsx+WzZK9WeQSXdNPclgA1faW8WgDDxNEpky+U/X/aoKSPN6b9zWsPR9MY32m7YYSSJT1bRS
3MIA7kLWiBox1NLesYzSlUCwc5r8G6H1DHodrOxOcaMoxBhCGWkEG2xaTC1DMIXvchFZGuNzpcMT
i81IYfB2nKC0X5YTUa678Q4RWiDs0iLsmoynO3jNy9iGGe53RLlrEAVL88mVEahoX0wH9UIgcOxM
62DBQFIwlQxv3y6G5Kr/QGU87TDSwJ67lwgMW2k3FXy5VyqISFjvUDH4KxjCmTYzrd3Mp/vuNYCu
m1BBfyfpIU6HWGQlYLBimoXOtdRoeUTDj3uiTU9mc9D9yRek4Dcjsi/dMa0S1depb5Zpovp6x9wm
l9mThMkvEB8LRld5QO0uIBdkmgzWuWzwdNVUREA5BdtGmaSoKYJ1yhZLVPxIRaijljQuWoDQbQ7J
/t06omkmwwjk4c08mODpX/gjc53jRikZWXviYwRJIyXeT1ibLZfhw9PWQLVHnUkRkx4wtxKvWtGx
FqkhA/wm2xm8P0QkqE+C6bauXq5EhKqAffEmBTFC9XG8Bbt2BC0CDzeJMoHBe1lHagVgji4OXMXb
xd7l/yxE2apTrwM39PjIo+QU+BBG5jPe7FiXxHXQeRiNn4BC1ut5CLGoLprdxq7HRXbqDAOJaZYz
Fut+X/TAWNX4Mp+ZNfe+NWFfoNEN3kGrWoDhM3dGSgvffW7ae5/GX6xuVtJ8TxTUfumFdma3FVGW
/GTCCOzv7zvV+bRdHfosFEHIGu7TErcPXeUJ54BMzucqxcf0XTwpSh8LtbDCe1IiCYzI/ZyIYNWa
E8PqcENOcqMsHIluo52OwTe/LsDPqUSVivDZTsSS6g6YgvOlfDcn1SWttd9CWrSPcIoF5pD3kJ6c
lrV6j0t+RGdCWpeQN77t+lSR8YsKlLZGqKyLFi+M7GwQqiT5KV9WSEAAm7FYdgdPwM8lXYiuXOGT
XJUiTIExTRUJgvUFB9Bo+wlKyWASepCPoRkvsi8nbVXOajkhE5yIhgYa/IS8es/5wRF1hLRbZxlj
Z4jkD42WYTvq+4cQ3ae7Nl+36HAeNDtzy0ddej35r0iIgtXHqeEYrqZQ8UQtOyxq34biSgcbRVky
NGW+q86i9JVZBK8KtgBjoh2C8UKODIQMysx69GeAi+IJsacTcCAiR9GHykKvffCzQD6D0I9hR/VS
q5nmWT4/89u+a56iAf7yZ2g6bpD9yL43L1YF0xr3j5An5x2kNaMj0rXx7vJ2aVMFM2Cm+d8+H5/l
Cu14IxNoLTx0rmF1HKPg8GDpMy+445pA0iVHCDAuc+TsQek0yi9hNwUUdf+3yOFYfbdecLytji0y
gKOpUahxsTmeIuMH7rPYjiG32qmb3VKjH5jSw9yiRk8jv283S1wcoUU7qC3j7B+Ox/NiutGL5Mlh
zE1h6aDQfCziHQB8IV1x64pj+GLULzgY5p+uvjsPvFx0N1rf1y/ITrdp0ucTSrZeKwiAKOGWTV7s
z8AA+Ep6LBEnEwZ75KwODTms5lbIJT1g5L5cwZmQIi2xz6ZjKU5jB7FLzz6eFTWqXL7M7Ec7uIgb
bKFZIGNTCSchMVcwj2Clhz5665KXx+0MrMehuBFEH2nxeCS7d/ZFxXNo+C5Flfdq7rRil0/W6LxH
YUqNhyNHzDGVr6lkU+0XmbuEKJcUBdzBN5aTTfNx/8qdxZgMEFad/rhAzurQQYH2vNcV6mDCRR5c
kc8K30NXEX5Ib6H9BhU7SRUrF8feaidfhfar65XTkJTEBKAnrE2iGbLsCaS7WXsWpRLC6k17xrpb
K4fU6VWhkuaGRnjmU2Gf2k6io8A20QWghkfZsLh/tVtlnsG3AMfZOztHQ4YBZCVvSeYLmdSqdbej
w+4NzP7C/i3cvwgeKq4U/hQNjBC7I+Ip1E4aQDbKCDCZmDfvBf8yuwg4uuxCUOqTD1lsq+o83Vfy
D4oVnNlSmrRdh9QF+re7GOU7go54rE45cUBU4V1LMMIKoePkk7EhGZLqqoszccaHyaKac0DsVEw5
lT+/RiLAc19E7gMSynyR6LkffQNci/28gH8FiFbNg1bILrQV2ob3rvWs67fxjCQWl6tTxXlRWb++
v9V/anlpvmwCH17oL9cJZyQ25iQZwq0YXFMpA52Kg5CYm+Kn+w+YUrUkbfw9xNlrGRJZSrdpSg5/
pjVW1s0F2c+QcegQ+GdUJToE6q5X0d9/uB+UU96SHhJ/fnmwRia4d7sufJ4Y1flnRatw/Oo5s8cr
TiyRCPxsXwn/roB/0d4d2ywk6LW41cnj/ygW2sAYLUbUa7YT+zruaUk+OPtMRHJCkq6C6jPGGzvR
4P3ZjK9Ou4JTBIz4yXyzv6GkGSV6ucu/lccw0DtLi5BUaR999O6gK0BO+MPWSaPKJ+qHYHqEr2Vf
S3fldCy/28nBSC8EA7gz4cbdDutWJzHzODJfCBLa4ZelIskYxyWBQpnGH6OUwZC45f1qj/vGOg7Z
sGIFWnCDl56z6FpYiZDv8/9I1jF29Vw22njAwRiGIqYH5FClIe42UJohnB+F1E2zvisg1fxzzW/M
MCi0X5gGHcr2RyR7eGZKjk4V7dSJJEG/E6ZAhqP34DKgAMaHHT4pRVCTG1aJtyJh69AdYExr9oB8
c8FL0OtkuqXtdylKY1gehNXm1asYevYHovIJ5MaiSNniBig+LoB9pKLVfeNlWW1gOElRb8p6//xY
WQ6E8qCL9/F7bSNCxVXdxlneE+a8NPUWMpdXM08GiLX4bk0JM6RUrcMZGZXw442sJ3w9DWffm8ku
ijTC/HaLgN5inwRMFwbkKKpIaTnx34gh6ghr9G7EPEvAaM9f8lKD4HE72NdF7KL7uZ95toZzoyyp
bUPGkKmrJxO/da7pAjhi3cQ7dFEp8pecvkOGuOlidjgafFpck9Pc5gTOzpZyFZb3syAseQ7KZNuI
0l/Q+kfuHPyFtOzVJwAX7YV8wG4FaV//ROGjyxktP88cxcLId3XrSt+vZDZNEHBMtBJq3ZKTL13G
BGSr4FzVW0X2kS+esfUKscxs7FKe43J+Kgb3vdlCRXba873zUYZJlCjKTXNqTrIl2JiAXC375Uet
lMAHwK8OPn6eVYyD2fxhlRpg9JqSCxmOXQmbP+t82MntWN3YHUE0ag6/Oel8viLHU0cRns3LUAu1
2YJE1p9BDY5Hpx2RqRzg1OIBXYbbWe7K76Qd8+6DKSrJKotm9oGjCn4ZbJl6ld3iVfXRwShNdSKT
JrHmEetk7CZLMCgQETf5t3axDWVm3BJe43BoXSm+FeYlBRylIR3bdie1IPxQXsK+BWAH01o+j5QU
ZDIzNbcUxKpb5ZLv23nEAg1LcZgkeI1kDO0+YchSTIjSUwBOeBHZahLq0n/fYPT8FSJ0HFW1P4kJ
4EcMto6/j9V3i3o5icOgHNIF3DA4TfoaHV5eN32COtXA97glhJ6tHGFNvqhh+0cRD85N9zEdxjI9
64LDW74bIRh6IM+CuyhaEL0bbwlRrS0RpBG5wNZWs82gK+n7JWsNilJEb/M/WL1BH3jGWRN9R5ZG
a+NE3mAPsRAGCQxU+OxAPbqAduFyCvMs8N4HgtU5yCRuFpAbi47PO37hgeutZ+AJpDDRIkFv9naS
U2JbIys7LMnWktzHbGtKt/8m7svpfUIDWH1BF7knn2Si3r3GHLc/K9Pp2cd/fwnTVh6mW25rGgFs
0Ii5jF2+jSqNTyf5gguLyjp7RwsZOpD0PMscQg5bI82q1xc1iZ5tY6qxgtKkjbv8r3DXmnYa1VyL
NM+ZNOTErVyi++G2HoZEnaNjlWFSKDFDuaVfcyf7JO/+0GFdBZ7+ZNDL8zRR6mIv9KA5OW1K9Nxq
jDxJDMAJKXsHCTIY8lCNAkdPC65ld6XvqlHpfxq8Rj97UbSQn9aXlmShq0VdeXgcsQF7JTO3qW+y
sf0gjEF799L3dsdcMjAPykHzxEfZxPvvnrj7GrpRmy7cPoY9RUSuhUdgEwCCo2WM5bmNAA+hlvGi
4Vf4zqvoN157krvQIKXSN91SQmfh6gUkIlRRDnIIV/iwq5oXbFAocSId1Awx3UnHKwDnnvOCTrMr
tV8lJoFQ3OosCTraDHYUwCXRuoJ/Kf/I7Z+FplVp6x7uAku16MxgejUhsc4Yh7uxnoKm/s/uMMaa
Jy2N3JVVXKpw8JLdE4GKnIaX24iey1vnLKygcKSQ5laIAbMkBphsC2adqNX9PlEAQ9fWUcguga8T
Q8rDh1Rnp8pxFB9+eC3OO0p5tOYN9R8PhC+TxtPDXuh/gi/tmxvJ44jyReVCD7L3Dh6c264ee3Ui
XDR4GjHKFxgYBTqqV79CmmkRKay8V8Sxw3a/GGHBp1161TppTSER657fWxJJoLg/2NaAFdVIWque
y+QFcKaj2eguyFQ9kG64GxUNKw2hy+6p7zM9ffNhvejxwwqg9CcD4dMm9HvFOI+xlCxgrepccprX
XS5FNZ+tI5XiZzehiausY23oZ9HBT6YZkpNxoGDYvdFOCXN6Vy/uDkPCr8IMQRS8+s711uWZdLYB
9Sf3mAtkhhl3upzz01AhigGHSvDxtX8V8QgGc6UeVX+vkutmNDB1EdKPSJ0153YLQZFaU5PJcCHP
uOty3PG4AfAJked2WP+6Hytd0VtN/xXJ2Nq+wgYmx47WJEVgAWpUZrwXZ4+ZRW6DPOwpfc4KrlUU
lksTPMQrKwAfsc20/etAFoMtd+GD0oITvGTOjd+Uhqaw3vx/TZCdbVt3Z9Xb0E2OZJXzo/O5NGMw
0sXmMwFuqmeDt2+L7J0971Gu2bdNS5RSI4P/mYU9eKxAQuUagwnhlYfsfkNM1ULfP1QNQSLyT2RM
KTKAteRxqTsU9gawnQfLl/baDDCzzbet9n4393rfCXl5Qxp7qzgbTsCCxISKOnzqpv1hcQINbIbQ
q1m8S+znrh2xfLT1CqWtQPnpuDS/hhdKIb/ogjTGms+uJaTRz/bL0yjiaBbk0N0mc2e1f/KxzRMR
S9vE1MeJzGQKRQxyMM0+U4FqrUY9823ojBBo7TZo7kkL4EEWawhNTfqcov0A1NfGe77S744+g1Jl
RVxtXsqm17Q9agbU6l32NYoN3yyQREYcMM4q3ZzWJyFz7hcnboxiJEVmiuTMK9solXQs5dGa4jpg
k5djvTo8rOKnHHCSwsnihMIUe6IL4uYvnKXqpH7K13z9lSFJcZ5jT+wEke0klAV/lm1h9liRENV9
zCV6bJ6Vy82TAZIP/KFykWSaMFqUDVFce6o8cJPvgy2TdCQ1VA8BN4JNap54xMZoPCBay3+/5rP/
wcnNyYZhuBS0S6Omwa5t1P13roZhkk9K+vYw45Rf1hcPM/L8QlIsFQh7k8prQxEQoInk/Ghk14Nd
VVdz4OGa0q2hyMMLE1zBGLKADORRpLKtzDwR7wPyIp3Ebwvbierfxm8i7ouK8OVJ7gUSOvzFyMhG
X5IKrSonzqwrNXYj8IdIyrSK450A4rnR+5AeQDBdErOTgbRsm7JucnjrzpfH8WTt7VUTI4irb/K5
HvRlmWGNYAM6rAef1VtMJYp4xYlz8nVK5AD4kj/jvDmJIfLfURLWoFI0+nXhap/pZ+bZiY6UrmHu
su8LIHJ7u+J4hTjRbzR2uf8hOVerlLaN3hgrrEO4aTsDp0oi5PV8S6BfyWk37KWwlN8mWMF+9dPC
YVxiF6yOvKGFAEMNy3KFii1+OhY/GZAN7EvfzHcn7Bky8Djdd2ISVpmUK49WgoiiF8pfXer2rf5j
H5aiLjVMhr1xSLBapkOy4xs8nyfaNME3fgXnyiC2CYqfzZG9sX1AzHNQybagimqRGZ67B+A/5o3L
HgN2EDkU/xyoirt/nermACRKSmoh6BqcRg8PJYBXPAo9DoWbLNkeuVLS5oo72EcWu/xSuS2OERYT
lCGuyBVjFGO+iVQ++ilm7dDlTGC2WXopLAsj6mzEFACZwUhaGDRy2Dsvi9+EFXRfGpVxRd+FDnsl
bne10ZEPbm0Jl8tj1L3TNGownacSOOmyHtORf0iMI6GDv89yeo4Xae/6163LTlitFjpASJcTaltH
qtjSgUBpf0iJmnXPJxTW5KyWrV6Sbw6Bc6MWJy5kh+38EArKMmzgt/FY6+Xs3y/TecYTPwBQTQ3O
hlImcBmHbWsp3rxbmc8V77a8kuOWEwmIAHQZreBfmNjp88zri+BmhjlCgCs0+YIgP4Q0m3cHXnld
fvmlk/noGaVmNUNXk9v+QcjMkzmWB9XhCux+nTsqwBeJlbCylBkWJxuUJNAlytvVWVDY+CpOCPJf
OZpOaXWLfr8RUBegemnaQvIE+FUrSUAwqn8tz9W6IdZ3m0n3/5sHSI0BkDaaFR7IPwFwAthp4FVc
WzyzXClc2jrewmAbIOfwwH/3yYrds2HUjGyRTLMPVx6UK1N6bVIE5A8XrUnq8QF/DHbhRJ3+6dt3
jVBGZzGlc4X+8LjjNaw1s+c3OyALRordeJAI6mNvWqSJO/HlnkBq0TTVC7qkUx/1R99TxRqWPuGc
qKWHNwptJx/i7p4e9P0ntJavTiNUABwJvlcFAmKDowcbVp5oGT9RK1uEE9JDukrO+8QPL1u217IB
3K004hSf1YCNwVMQz2iS6I3dzKDVHew3rH+ReDE5FAQaU0MD71s9gs70Bejf3XcdYd0Nnedi6zFJ
qPFoboWF2Yuo8V1ewlVMH/Z2LMT0avPcNGJJ0o3ZVWHpWx6iW9z7LxLoAmC0OCSNfrUGfD94lZlt
3hySgz4lSu4GK+seKcwcAODNUbrLGUB4xzJRnkrL9oAHkHRK1CYimrtBjSqbUF2dNOQ7xtoJVvlT
RJYeijagy/r4CRUq/i49kyc7lhVWv6lMgEI/RirkOxfedIQtRHKAXHKq8e8A2P8YaDDJiCx/aDXD
lkCJzusIdYA6sClf6lTX8aVHCyokDFoQruW1ezo9JwmoPnGK2+/jyQzW2aPOHACodC0d8rqA+6YQ
MS7Yo1wtUVEh6/zB3S3gvvpoQsct5XFN9mYpkSsPkSOsljdgoBg3jr3LYMMsUvR5WkVZvPSJkjHJ
CeZzzrb7oH6kmPmAhTP23ZP4Gj7nWLW++n0F1OA8//RREW6ifaPEBNGNHlE2BeM8xR12jndvLsIF
L/NxIsrObsMIBDk8y2rsT/XMBw/XJ0DlaizDeqV8OCASZ2IJH4Ep9FEg94vVx1PgniE7OvmAkjEO
b9wSdATB1YI+v8cLBeyhSNUuqjutFlYcnbEJRfVdIy4ASykOIaQhg8bviAjFH86mhbnOKmTpbjke
479pQmffaCRNO6/cEwRV+2zaF4k+OWxghefjCF1SEwJiD42wnTETst+5j03ashsMMmP4vPj/tMOs
XKVyTkyS41miDiCHBzfhBXBuBpppJGLA+2n2dNCJ6v38E1vvU862H3KgwBYSao3z9lrYJjC6iR10
3V3Sh60CKay61tOFfIYncRDQgmUYsuwrUD++xpDLvT+U4VPkYXfdpUmry+0oIZzKcYBaETuuiIgV
vFHAqE1ArIAgtnbrCsF/ZAsM7JTYkKd1Anxd60vBsYrpC4cjEg06drYMSgadaba8+WVSp7acjN1T
lViNcMQnv3eXpjwCHsrGokxgsFmtZUwXyx/Is7MQLO8klDxRsj1nVy5BVgUIFrXpNI+OgLXCih/y
Ecohi88M39NckV4y/Wjob1o1lJcqfXL687aagwRNApSRYumXnHAT1eN2zc3fzcVdLz810d0dfNu1
RrNxmctRuxgB8GsPhas1iuU9mZX6SFAIJ0cNjhMMzVFpxeMMjLYYWhhZIjQAT6HE3Ywb/tXkkqxU
LxHsweFqXYUEcApAHBevBVW43bzgGZsE7zX3yOxZymj/Ibzj+GAXmgTKjdUj77u2+11P4LvZVjod
7P+Nyeg5CxmtYqqbV7wOZ9b4UgJF4e2zAWvF+RlHNSnCU2EVwb76mW6vpR9AhOXlnezsoba6GPVl
0szZS4mrq/Ni16ssPtqn2Bj3PBBZOCSA8qZDhUgVdGQ2pcRkx8R0WSFxnPclKOfZJLdVFLZscYRy
aTHXJ7fXCM4e2a5BL97FZy2+mEmQruUCgsELMWBvcZLHDIA/E0CArYJl8o/ojZrvhhWn6+60PHZK
YX/gZsYP/2u0/flapbl5aNADlfotSSdBGROzpl3/7AXzBG21gcBztDAt8MWodJBSfTvLBJw3hwJv
RwJ6FZ3y9LSR+xGNrNxqxvJaCq0QLewp2n/XgMyVnckKEVjt+9TclhtLn2enXcwegntLS9ngC48h
bZA9YZMbBTCrWr3uAZl/IA2b0rWSQQmbrcVajbLtt4yvxoIBq5xBTWcFlYbjDNJQSat7JrI700jO
KpH4jm2JEz7P5dEmuJmZCc0y9FgDrqyUVSjyOrvgberrvC41GynbOa8eBZDWOxCpK6UszjM5KJoR
rfZ4YapNH7ZOAdQt7DP7GfDYVHHxXZxiagFtjUDQcgZOU79eNpMf3Fc10emiQ96B7SiWveV0QcnD
Hlgov5GG8mkUMo8C5SBuLahOQVqXWbzGEQxkk4QTPwmRvQMGG03UigR4+S61BEXAnTnUSatqKTXV
2aHgH7mRwstGkosg0HoXFLoXpKr7v0dP+Qt0wgV31AMTll5FpopyjLUjfZHXWOasA0f1WqVwPGhH
Y3vsTEIkx/Pa4iWhJiNxEytgU6Rfd+Zs1yxdCk5ub59MyG/WdJ6Fs4/ard6PIyukdwR1889nN2L+
VxGwOpYuxEn1QYOE2Q3LD2NxPU9MTkda0phlbFYEEeyGKjP25D+x+ittGoS178y8sf7qI4YkToAS
oXcVoXAefQuSDVebqTq5/3Q+Wjl2OWMhMPIW+kdwNZ/y15u6rdjJxAhEX4HXlHrOEE/YcF7spbqn
YjCtZjRN89I7U+rx36inXk4YfKqlZCY1/fRi7DuAG8mHBMnMcWXCMY+IzLPDwsteVmwpHpG9YAf8
FAzDvjtbUlE1yZbaVxt3IJKac8d7MWb4PeaFgP1J9WBXLu4mlju7U2pbVBivn7Zv6czYHJpaB4e0
bhi42ai9NnpqT8Mfy5Wi5sKopQa18N+P9R8yykw4oPDkHAfLyWOJ7ncEnNRH24X/+AuTIXOPgaY+
QR6nu47CqrQKTOg1ZJIHdmuaSzPuI5iWDDC2RxhcfUnKiR1jVV9rd2XElOZzxC4mbAwbkrcobpZ/
B3nK5YlfAiyIEN06WBqszYWo4x7LSnUXNUGXhQVbzfrGivUlV2FsMTuAeuuBuvCBtRGOutm+LrMZ
cU1+I6VhDskjnloYBLTIZHEfRBVS5V1OaoyUVPB1xsSsXUnODNJn1YQp5ZM8u9UDMdUF0/yxIscq
JJRrXJyf8sQBo10dMYBzi5TzhlbWx+y3H2e0HbRpqdP2LlVCyd1R3+DHZnV+o2fcv1vyb8ohQhH+
nzYWpT0rKqzDSj+so6rcAeRYlN6FdodXgxg7OhHOoH+jf+OAVJpbK71EeNtywvgmmiarg+02zbOb
/bCM9FtW5/gAATWN3bw4LjefnslMCJte3wmebKIJ8IeEKjxlJwMXxjsNJF+PUUHOc8zB98lkzBNT
suIAQ7pL0/NNInWPqHAz5QmPuGih4udVb64CdXg4Cx1LeI0QQwnWdu5Vh2UkhwkJYXy2ktKdnZym
iBGgSJj7aNFjWmfdCyGGyQSpF5mcfOtmw/iceF9X/LoLDF6IJ0cpr1+U78583AShtuATEUvqyetd
2PLrkghRK2S4W2OI0HA0KCVaBp9aM5MEvOhnSYgFJHZS+xHlfzjNnf1Hnwg0M7KMRzqMk6fYefov
k1Hpq6/x4PO2KJ3m1wKVEB1Ei0X8clRyIpj6MRoPLNqAks1010vxJM8yFSaDeqIVd3V5lerUlIwU
CQD+0tQkO+0VJ+2q1vhgA9TGrjp5Q8+Eg9jIIemzk3/Qjg2b13dngqkoBFeJIIui+l02LI9yA32D
8isIgJCSzQA+sCo2TpmB4L9ntq8jxAA9+C0r5wRLr0eAR4ida1DHZNfRCMJFmiX/7Kl07u1SdQzc
AtzfL6LuLAReY2QPK5HvJtLTbkhTnn71VwSfULApGyVB/VBXaOjVwUXkx/Uq150ZqP1sl7EWp209
y76WtQF6ttM0rnPFcI4Et/xL9jYVpc5CYAGeXDC4MW//Qt1sK9kvTHxV5+FAC9D2P8JYeLe7u7Ok
SYXQRHdvySyxQCTBkm8Iejp1o3q76RIP3UmPkctdUsWqXW+tjFMMrJSrtymMh32Q/3VNGagxD/44
ODvfUO/1SrNgHjsq8di0hHI0RvluWHoZW8ENPauZc8djwDOZkGBgWE+X0nIDtJ35IhvtqCerd+SR
0oT+9aVwaYdZp7jn5/aIWgW0184zldyThiBIUlfF6XgC52CoIbpbXCvqo9gtxNyUSxrdywwtDaLL
0JZjXcvRzH6t3RtUj2QWjgZEf04YAtM1al7XEH9Q8WgYPxKy0tL23oKR+shcj/JgsbVkaxTi7UDC
Zhnk7KpU0ftXISOJXbmLMO6ydhCZyu7L7rGnRrPdk8KrHBeN2L+XRoCwwzzYMBbSqNXaHak3b0WB
NCdh0AyGy7bZNUtGlCK5+3NQEj8he+F5eTSBBMGZCOpx3e/ASdtD48dg6dGA3+R+V+VqrE3YtnEa
MbbGs6z7YoQ7+0VS5XXIh7+VYHRA11Mze3qvyaNVvHyi7laZc4x84ZVMK9ktNrPxwXqXK9DCOPYz
wGhGsgAR9tYayB5wVOEPkoqomRm/tMg81xsIBPhZuCCNHb62qwonmKJCCZamngVngqZgWDC1WMqL
0A+NHlVk1OOxrPlOoYbq9s8EDNPgxEcr8dXiAk6M9g/8DMk3pb1IqkVxZpOaqmWYLFp8qVlXONtu
nkTv/aXTsGD/5V9X2wReyuKzG6Tm9d+YD/WUm+bz6avdYTUYCZZqDCAbJ+/I8kECBQA9sHO979FF
7uwSWxMxjvSl5un/AJr4YVomtULKba5kWkn8WsVwCCuPvocI5uck2B/2hU+ftDgwtqLNVS6FHUNp
uvPS5aAl0HRxiJ6J1987GpiIEFAdxEAbvwAvGJ7cHJlBsWetX6YuZ1OZUCRQ+Nx1nKffEW+wmRry
sKtiz8USEyu22qPG1UoanZUh40kbD+PRngX+dpOeTqdgEF+6L/LLFjmVEr7TMxHXRuk2RERZMtNK
zEKrgBgmfcodM3/bgmbnv2mia0Wzn+rQdCMoZe6jt+kUBSFVd/G0yPs6kK7p7o9HPeZKI8C+asl0
U9RF7qpQinjL8nhqBD2Av9mjQGvNCE8/l1xxNZdxLPOwhR7sAwG3Uo0tQRzH6damNzZ5wErzAlJ2
gZkgPECT/DGFekFmRhSWBDxVhMntG/ZRszIxVRS7OWTYTSEqW3H1Yde/m8zhSCwdPMB7arsb7tzQ
IpgZmy7esiFGaVv3PtJHzWrU00mev+w6WT+jCE0DSE3773jmtpxj3A6lyfw9xCLyNK0TwLYLwxLu
H7bUH6IPKYzxf4lPle1vdQ6yEyGOm92SnKKbXXTYNYi9KARKHpFs4QOBGiUjHp0N5seVAZFX9+bY
qda2vM54B52B1iG8k2HnOXbVfr2TzFEDT/SjICdq7u/m99vBMlK7Ce2gi4jHcV7CIIHGnLTpgVHa
Zh4d4tptYS2KgRu230ucqRnBhyxnhZ0CtQaFtu10s9BEY692C4z4IW67K5/p+fPei8Dj1mFrdRDQ
DOQFFWu5ZKsDDDKWH9+aEuyex2rnFI3oayTy9Fdb8KmmzPh9Rnnm/6hxTvEd6Fj3QMmf0XJpYCGb
ijY5gdfxRybTsBG4zlukj7t035f8EIEB1W3Keg/5bhAPsdn61vXgweKvEIEoqiR/tNzWC46qRhlI
YEIO/Qqhmo6qxrwfTv99/dTWPqS5B90VwyJzQM/CiTKo4PHwpBoaRJcytQ7D3pVPUY/HAqiz2PpR
yp2rwu0jECjTtco9U5J3RQwxLptntxNZxNDdDif260zufR75e5UKGPdcjSlzL4keYXv3cfdkm/NX
3XEnLF2tzs379DS/3+dF5t7Zcxu887llr1JO7y2uHYHFOi1pTto/Gww/o1621y1MWsLdxOEDKamw
TYefu/tHRS95xtIAG0X4IJpAiMn+SjlABFtBJ+gYHa7WZLm0fYmgXG8tO1gvan0TsAJHsgQNWREW
NciVGNswgWGrUTi6ycRhKbWVKZnnUhTfm8hOJ4EHGpymxvQ+GxtelJPb1xFSMPyr5et9gA3BzmkG
XK25kAvLnUuW8JQjv3tWuYPG7pK0DJN8AU8Pht4dPQ8j9snieWe7ayim4HyOYpY2qCGVzVmBb0qr
EcLwn+7Xc+CvwftkdCtX7zAz/tymcLVi8gFSUHryqq8PxbivWTpEgudNC8tPl4AG+deu0tyc5WLh
Ed0P5WPUPSl4ts/5KiyrrqMum4WooxolL41ZvYSwQDWRH+cZsIu8wYlG4P5wKPoo3UArb8wDLYhm
GsrEWET19LUu6iXf8f1r3hQLxJDYzZS0LlnHy45wdKMBtgZJGM5Y0S9jGT3AYyGhvXb2imK45FNc
tPZKtCxkEobdn/6eNwdN+BjS/p0iYLkSZJAcSi1H7dZbbUb8RwSHw3Xdq+kwWP7oTUIXJ3IoOSwb
2ZTDwrqPGUhYEf6JIrdYdzAABfVU6iQd9XCQ78uFRLDMB7HukrnZ3r1XiQQs5v8hXK8M+ICSXGt0
jRB0M86UbB4gIqRu+EMazwXvLnwl0GbZrhv9wa8Drg6Ee80MXDhWbUybookfEe90xrwKfeJxek5y
mg++vqtwbNon864wB1G9RzquyQwyNTkNbFerw2syy+IAfIWviXQ/862rYpjhouRzHJ92/Ra5Lwmf
4IVWLxOd4JgiH9uHj8dzc6/+EUg3s28A+/qUBe34xXY4FuiDpWgWAIb7mabhiBk6XbVhLuLB6YRr
s4ViZTzVNvp5sU1A+5+yQMWXpL3K3gr7UmAZtuk7aRTKcwQMeyseKF6OWVQ0tlqMWR5Y1GG/tqDO
99bLDL8NT9u7uCD2pG6BrdjPClhqPyh2n69BdVRnhQJO5GsBajRU+qGugJeH5HgbvKqQ7XoHgEc9
3GSvV7NZ4CR/pZ9zZPt3Z7o4uTFkpRkm1AlmWKFLcKGhcTE3KVpX9SMohoGV8CkKj5SJg2oG6d/f
M543oIZK/f5EBU74W29vzH66PM2DCcjK4zJbtPxettSFl9ECfEC+BGAlGmzTCGrkBTXZTljuIlSE
vaIS8U6zJgtqhg4o1SJ++1WMKEobTfW52NXQ9NpnWgwO2MY3//g9IEMwn5axEmBulKV15/v1oW9A
tiwDA3YM4h3zUjd1VqqbwQaaMyrOc6N45J2p+dLUua1vOsDpJW87k1USXaoVrOzhLAJj3DpGQr+6
4igVrq7alTPBmrk9DZLb3ftq/uFoIQXkHcHc0z55Nx9G9wGc31ET6SPkQPknqWNKDh8w0YQ7+Wtq
l4IwDOLHvqV+hQWQ85CBn2+EhF6HPZcYJOdaFg5IGGoLcBcIRBCaydenUoXSeu7E6aCJaQQ1SqOB
xx4uZ2PRXVlnvwWsEZPnLs/+JxPZsXRhcK8sPGDNHR9qQHgpyleBP5z3p3Haxr8909i9NkTOCF+g
B0r+4aFGIskQa210znG+Oc74+8ptuhisE3gLLRPi1y+4PwQYbpL6M/UY62wLs6FwI7ZOH2Qrqh2V
1m7SFotJs9W8qnj92yEhEOlKUYrMoQOPYeV+OdwA1y6FnXcBUcH0iFejYR1XOy1nLI3qY/kVhLCk
+QgmmIK96JNB5/WZlPZpP1l3Yldz5Mbcd4B6MObyw6pa345y52g12ji9TeuLMWamOrh1z+gqBo4T
o0MgjXg38xpf6YAqF9uu3o+SDGpyUVXh4VZOseL/DAD9YN8Na8zp8JmEsUiyAq1dflt1OpbMFcXo
uBfLgv8nM/rmfbxG86dxZ26bXZjnrzLv60t6cqgsTVuJRMlAjBCGznVTtcH5sN2vnpBfSClZV7lM
knoqX1ZgGMd5lQWr+Vs2+5bqnJyoI6rR7cxDD62/LdkX38hJvI2YWHhBKV8SjAbQKxybprZTgChx
6M/x8SeyxJ1tO0Yuz9M6QAAYlvlR7/ssl7GvM+2RnPIJKaClhFtilSoLVHVJhIGe86izOhSlFWM9
3EsTLESjJXJVQlvqy4Y70/qKHCDrECcEWLX5yH0AQ/3cKmqFZqVkKhOA5QgLpVpniZTcem7YGfgt
cicpnGtgN0rRP56ucGnxCa67qNz/3OAv6RIsmA/gkau/rPcjg8wmQ7FD4lcxUgvKHCMOBmmpTEEL
hMZsXh0HkW3DImCkpCeE9HQAqqfkpPfJ1UKRn7QBaTYkeQ7S9uvytwz8eSKk21JRcDwttx+S53Ia
rChdK2WNJhTWfDim3yKicHROv5davYh9l3lYWJPV1WD+gwV/k/qBYwJZBJu6GfXwsZ6W+uNuNFM6
7MyhJN6WXzh6lY0oAw6qr0KJNzrvr+uywJp2Jq7PFAlU/H7nXbLkSx7ptUeg4qOLiQnG2ct7ONM/
X2dBvn0C7wbYkeTWlmGXao6n9fyzAb0WwX+k5JXJPEiPv56YArlk2dPFgX6imTnt8MXU82EvUg/h
tDJNAXcj7V1DZE09Y88sWMat8IMD6jfGmwsRa2d+5XAWEsJIZYNYVRPvn/dYQaPtfckJhKr83nvU
Dxdp7zXDTtZ426vkds8o02xiPrsvqaIp16+ds8elXk6uKdwv2o+gEmuEqsQiMd9YVAJUVvvXSaKK
keFBTWl+/7v5bEAv3ynoodLPMZ6w2IkuflUKkh6QBwZaYaxmq7R8xeluaExFpahVM83NAms/hVhZ
hTc6++IgbBSH/t3KXHKAwC1s9hflWZYFmdr2FQRIoK245ywqAPfOWfNTegyfZ5NrM+9dIFF0H4zA
WOXwi9GAvsvL/+LKURSIBdjEbqbZHqm7zXPyrlj+2mviJHpT0AABkukSuJFV4BSSP87jMUpLumXx
TPfb9cYeG548c4OuCKIpLU1eQ3onyL7N3SMONS9g0QwXBQj8a8RpfJiDwsFkE8IDzUL+TmJcCl6h
9XBmYHDqY0435LqpflSVu5XrtEfbK5ttuVn5hM+/M9WQvvtbSJCNGrIEeKa4QKv1ntNTHj/9tf5q
kbe7SUJhrvRaCbV5EV19QwrM6dNBwqITXrJuZeu4WYjX3x97kvNP72Q4XipEdu15gZ0CTvHQjeFU
7giLKnNhjFrTChN8hcODshJ2Sewz+Be8fzOkWQ3XPBY/GQUdvnrzz3H4vyju6tDr8HfBW+oBoaPU
Si2KRDMokfBTDYkkfRr6k8dtTy8FJNVDI3jX612ZKkTxDqWO58PKEH5Ib6gTmqpqDHEn8TjSuWNH
yP6iUz41BEwF2WxeMAa95ZPAYEAvstWkNdaoQkfJKdq7UkPYUfyQeqJYn8L4SgN3LuroaVX9smGl
A9cnwy2XLtsPrdW7aojhVQppXywTzf3e4Za+vPm2JZzNxz2IbXwVtxU9PWEapNVU8ezvMCHYuZH2
368oLivS72t/rEU6cDHxjfjbAY4oNi1o1YpoVWPZp9UCWe5R6BpoZxZ5uBFyIiYOD3Q43/0+cYSh
EomtFIXG6HR/Q9+RlQv9uI77ZUIBnkVLccdGf4a767yrQdhS8pXVkZCHcSoYUuXFWuE5CRurpOhk
b+21J6XuLxUmVboSiS46+pPAZ154YHZJobsMxhuE/TFkD3j4IMNIKyYPlviUaYymAQ6Y2x4crbM5
4d6hh7LM1ZUuuf32zZ5T903O2SdDOh+ui8piSqJZaGaJLd40fQQopzkrmnuhb/1feeYinl3bhFtA
4TvEAP3yXXG62BwpeCg7ePUl1MrpxXz93wfmqBP2mXioyPYq1cOhycCOiig/CvpdOt1srQ7lZVsa
YjO86i6pyEv/wjYY1eQe+wgnkUKTaSrgS5GM+924uQKMEOPIDHtXnS5bPtSZ4owcNcrCqVriOAvJ
gP1LLuMHWjPtiRtsOM2PaSZe4fzIXNigQxjedDBQmFn6cXlD9LIb4h3nLckiNMWhkzd3y+4k7uVx
UiwB94EgLOIwdrSocei15fhrRdYPrKfHZ3sA4P7ESH6Su9Bc/lNWUv6eFPkFNSvW7VamzdRn04aJ
iuWp3pxc50EDzf3MERTsUvf8FhZ8/WTGyMbyTePnmJoiDcrOvgRcvmjqnMA94Q1pV6sRY1akoK4F
mz+EQwHQtZHf9OhQxybIqQhZ4T7kEY0fw+I7pM203PAHYIEYO3hws4UAIExR2+h6ET0CwyrELKsj
p05qrVBP/Fuf8nIxvKMFoeHCfMa/aQdKJ9Z+a8xOfoXZR+JJP/uMlcdynMvwfaWR2zKVwqkhMATU
6eUJr69/USBcICZsUk8TMxPTQWP2BudEt06mmMFlia/bw1LRuUk1jFsK0u/POjoVtsm1eq4EAYSW
nQkd/0T6CDg6CFeGfpZL8YYaar/g3apEjZPVzzdM/HRg8YAOUBIGjzia1dKexIoelPgLmh8RBsmN
BLt3mjbB6vOG7AX6kpHCFjPZAEgIZQwUYbtS3iXlTYRFnmJiZbKyEgbPdzYBWriJGPMEIJQAwZTw
x/lQK8v/Z2tvHECJC2JdqRKmxrXofTefv+jYiyQeq+HcsSCd35QQCi5GiIHoOq1B3SzIeiPPyrv+
hCt282IvuUHzqReVCVT7PSBGSzhk5gyvlkwq8yR7KH1ydvmtZAubTxR0wGwTqpIYjN0997myrTDK
l1hhdJGL26W5SbcGe1fDzjyOZDt8HFvkVBMMS/RmLZ9rW5PL7EruSGT823elVZibZDNQeF9CqSe8
WbAiBbd2V7Wh9hAIV+nTrCnq5NYMBCqV+3hv3XsY7MbwYka4jnHsOfsxD/ZPSrbYoj9PNrFUQPTg
/xhlIxM43alaICF1AFCufhGvY0KjKyls6R7TbthvIrTfW5WVpwSXEQkrVXC3CR7AX2mgH5r+fnEN
yGDoPbtgN08quHzjteF7Ci6MJAx9uT9CFAZF1purICViVhpYDB4BhKp0FZFttQBr/5+bcXX3d4hV
GOi+6XkKoAc7dNjo8nkmFH36T2VrrmfBkc2peMgfutpR+o9B74lUiiAY6MWTTqJWRv4f46dMmzPE
Rw0TgKCc1x0SFo6RpuAfVFH/F1J8DuSCHWUWD59WCN9t7+nPNU8Ng2vSal2jDeZLAkTegiZjgJBi
yf6EhofFUgdN01Ua6IAhpBXndXDiWxyf80sLwm3fD+NGad1QKl718ZOUIjwUuXqnIBZ3ML9Y+UPK
aCFahIuNstyxC9hG8wDJj5B8vMSprvCmQNsHszUF7lcTVSZuJgsfbW1JhXUH5r3SFjDGLEwqaMOQ
3bcjLmQlJYCO0urgmeD4MJL7Etj3I2sKT/jB2BYMaOn5yBcfCaXcgMjM7f8AZzfzdjOQOSBvsdJr
FbqftouQF9vezHPKXTlwZiuGy7Kk8lJ/+tXGRZl3tVSpOKIumqJ3fGgBKZNJEpTHbhZZu/ZL7sHa
e0BPwwJbXliaovu4L7qfj21noRjQ4ywj4FkQ1Tz7xhxf4/74okqR9wNMX5olezrU5/CwWVgMdj2t
Tav0I0uKhhIKxxNCJMCSDlK57ZpEBbCqA3T0XfR2Mb8zWFH/SdvISvKiPhjJ+cSoucda7r6nGmAQ
KFn08Kl5iREOzgaUMlE0MlT8alU98seCHisMZ/NXulJRFJ+oPrMIKO4HhY+2x5ZrL4SKBxwCXm1T
xaee4G/s2qEKGAHo+Jd3ioRT72zuBA4tmATABOnFxs6Z5gz9ZC5ef6S2to2Ce1qOIkpnpTOEKnko
W+e8v88e4FP+oad+jNl9Wh8+3j6xwDSNFDeR4dk8S25hy8mXZAxKZI+KJ/41KELuXLfreJtiOMO5
LvEc2XLR3LcMKNuzY47awvwh+DyZopSJ6PQBrATHuVdRnKFmLQuLElwi2S9YR8nPV6D0IbPDSbvF
mh3zDooeo2A++1Obg3mmoQInGp4jrHB/PUh3jZLGf12sQMuEC+oJHFqPtuSQspN8Hks7AfW/bH7q
X0zz/plHm3lCsetkV5dHRJgXoFMLM9BJ/Y6o4WK5kPtd7OQCRm/SNIQNw0E7qYFgVcaoww7LNJkd
jYqBcRwRXHY6uH8iIKAChXR8iWtEW1QTmQnXFNzxB5v0utm5pTjnRK11PllStiUOYzmXDkAkGoSw
SRF0ojNrqpDTTCzEQU8iKgmw3V6g/SiKNJMCukAWv7JKvBewvI3hGS+jSBXKNFLQ/l8egUbnSSVp
6T8Mf7rRQZp6cHNGZu+UlVpeROtKZh0QoeXSh+56TFaFSXWAZo20h6NlSxr/Nz4ruX88IecSRR/U
3soqrYmJuv8mStrSF7/VYXzTjYuNW86YSf/nheu8mt1ENbvejl7Ghm/D5qBA6CsXcdbP84uGdfym
DYiE/eGhjd3Qrrnh5fH/k+7p+FRhpvCkfBsswuBGafm0T2OcRpWyRPJE4QCUNNHhEgsp4QxrooOY
vIR0tkKzryrjAfgiF3AmffEBCbyYH0tC3bvBKvTBEGBxU4pV0wfWhNZwCQ94jvghHzumKzuvL12v
ktsDiulPT+SfpGIt3jo9Jl9J8WCpwI5YDqMKszQemEJGBBGobqAUys519T79orKJyjVvu+pvQCrk
N2dqlTgb8FH2oCrs+IUSdq+jJhcXiEHtx2+cV5LdsgA4nJix1g4JuO8PQimh0Q04aitaicVRZlO1
55Hc7iMKNVO0aoltuxyu6s13tIqg1XSAh7BpUh2GpWT542srhG6SefMp/Idzrrjiin56av6yvm4U
gK9vJKnfDV5OHH5AOSk0+l8JgNs8FdJA1hZwenpKHyRB0Tmke05R/5EbKqV7QC8fBXq5+AMNFnJO
7jAa7YD5ahKQ6Dp20yLHW6foL59wYuNmaBHWknmAzxP+Dy86ppCCE4ouMvI2+sJbShIxl82JfVDI
HjZugUaTU8lXnTVYZDdNLHYP/SPL+TUchF73YThByoAGIS+FOHXpaGr/UY6jO/vs64P1YXiZWQQX
FAzPGwBJWqIgMwktpXATGp7Qfl+AA4g8MX9UomxiC/qFfDYjQDRec80qqSRkwyNkGuFcsakeELrV
kevCPIG+4urPVj2ZSyA6IUIVArt24czPo0IHL6X5c0FlBjEdDg64Jj+KkgPJ1ESXbaBjcEEiiS+E
tmBd3sw75gdvXpEwH8VflNgTbEO2WF3VRn8brhlzEYb8+up4GPwXrdWqKpwsqLDlRGXKuJ/tqFR6
j1EzJUKfKL6BEYn4hwjJMKo3VRrb2Qa3TYkS+SLwPkSC6K6A2V+HONPcdhNvMAxMxpFJMoWZxQSK
+33OEWdeNHYUlkR+91r80rXriJ/4sSc9gZ6MkuPifWheK4xJ/ZREPZWvXRzX/fyBGB434IBMKtZe
DZiCtjAz7oP5KsgjcBgD2KSc1tGLnN370aYp3pdNAHL5E4nV4gMZDOh1tn4//Yl3FikO75Jt80sC
So2rCgB2/3Eb0QXqe9PUCx/JMg6AaxyV6fsOIyf4DowZfH0phW/361Fw1bC6GKqRMu5REmZDKYmv
XmDkpfINdKn3TniWol60x8ivdKdfsRa6XuSJyqBO+p5eSAex2veqeJCD1IJme2aunsnzA8Jr7vXb
RBDJ/Z4uN2DEShNk886hdlSHPGVZr4I0Enqnb4JVihN79NMQ84w6bD2Z8URN0asqXbCrJs1atmr0
oP4yTOJrVyJwVyuDtzONrd9B4ZqvI3W1+gF/fWOFOH9VMyAwGVv3ImdJMz6nAr3ykVyHyJPYTlYk
9QCdKw7l/vIBCPztwpThE8pZmjpHGZ7vD8oJe7EFm8Hax19MOh6xFj38N1PZ+KKo/ixdvo+dNlm1
iEQuclcPkEicagnxVl6hOxNz5MsZlzmdmL3q/A6rOgqtlo8375dUH/5PB5+mO2XtuqV8RRdy+oOd
YN7BzjLDyLqLDJ72HY+l8UqjmYtvJfDZiA9TVRj2DvVGGpzoBUAVx8T+TrX3NzkUC1jbLinq6fPL
8MX2a3Ou7QRAxHmq9Z9GYHLK02BlP032E45Cici3IryWa6G+ZJ2AFIDAV/iJAM90F4FEj9Tq3BO9
hIYDK8/fZHtugkRfSQjDKl52D2Fc8FlovvBVM08u+xByLquMLgucwMMHqcmAf7BV9DzriZsRJbhr
S4Pd+2d2DdSELq+ZgoAeHMDyveQdYeJaR0wauCdQy08Xk6pLRXhUAfKEt8sQeWeffFB51WfxWa1H
sOWPzuN76/3f6Ie3ZqwXd6kCgJpyCSmJqOwoM7On2NOLjT0oMlZA7BCoI0DcDsu09s2DZpdOZAoY
vohrS7ucgGBDDvA9qOgcb7aYweTcNzTC8h0c0DU07yYzRuNwrAGLOteWI5G+b0CRaaw+cHi3yuxs
hgNZFwOgTMKTrnwq09NUUyU9CIN33gfdpnRpeBH5ZAbxd/CoSaz+bm5/9PrXAwdWmdwyopHc/kyj
yd61X4NNXb+lEKcVgKozwrNhMDjYgzauxOHQSBNcDogDnO/SgoZxf5mAKhiBWASmEt2RT3xs2TZO
ZA70J89d5bTBwzZSCcm6fIF+FP8p6dBCeRhv7EdnsCtzUpMHH5BFNHRnDOaZUf0suZWp4JBz8gFp
nDgAEvwHv8VEuqkDXBAoRIwxF0bFQJuwFBvqBsAUN0rDnezr8ppypbpHdx+kU5lmDktLo4GECrRO
/WHQAFjYNCto2/bINlkfEKI6d2WP+RSGi0lv6hCu+5mCNINJ9ipHKOg+1VP4sTIHADBABH/3Agvl
vEiEtySXAoremA5jvva6sJb2/GW88Yex7W4+lugQWDcfMT4qosaIId2DoiwzfbEK3EYDfPrYNapC
0k+K4rudSXxwujHFKJVtqnLCoec/nXXG8pGjNiP4/ki7gdSJ51110GexLNsf8nrIP8/eYM3k/5SG
oDiqSC0U8k0HvLXiLhag8Q30tDOH3LwfjMQFt2tElStVmYJyiWLTPhVaddDVCUoDhDm0f8SonVjW
2Y7Qs6LNcnUvaxdBIuBVFK/7B3sTle+/DJvt0Qym2mlmUu1MYaUAd8AxYDGgjdJ6OkIomkyDpM9B
Wa47GBgiw8k5M0TqeK0QMesLqihDaz1/YG0mRQzuBudxH870yeRTlTmJoVuJmS2uXszPFecuOFOh
FYXa6jo/amuC1O1KhTEwrZ+2GPWtgHw54+IgXH+F+2+nR2IrlZNfJcYR+PmBKQf0YFJqv+T1Sy7D
SJstughkyIn3NCmXEMtjQiSr+nozvHQ/vh17Of2xohtRY1h7P5m8d4BzUONpxnzuS5lwYAr3ZcuO
NIFU7h012cKZRiqExo7EHcvDa7FilwVjmx435NicnCTlg7sg9LXFLlo5ITJx3Z0k2EYqfAW1OZwr
bJN7FvSY/17ZG9cw+iHLgOET40b3B9tYNqJLEpgke45DaIPnOfAmQ0jdI1s4TTGVvwpaFeuyHwTh
g7rFuHxlAQbxwIW2sTkr3QtaIQtmlLv366Tu8HF1VmfrHyyUjvrpAWS+02qyk2t3DUn3eDmyTOtc
VGt157UQNO4z6PHEO+8kBZqaTvAn+8cAna0Cjiu5MwM7vThg+kS/UGmlfNhNFLxigLKkp/n+I7tR
m8cdusj1UUYZXsflzzB+q1HnyAqBwJiOZjXEYnIVigeDtiT4FOQqUeN8GYNXqUasreT34xqLHpWC
evfdEIa5+E0vnaho8NXLroQmjfityc1dUELxnx6PjjpzPx1aypGmTmVpP4NOmkaTdsOlsegS/w6m
f2t54U+iKlZVL2IeqYOUcjyKZyZphD9IAVkQ85dUE1eqsNNtHv3jbjfsE633zff9Hfe2+JF9en4N
+JcmE5+U0pBsDWyP7ioMNJimO95SlFaIyAkhEsiIf80qUcId2CJdtOZwPWrfEE4W9JdxyfK8DZtn
SdIE6HKOJl2Qtz8PvbUItGhEja+8WjtEZUz7rXoFP6XLknrA57Kuz1oTEbwaLMWDa7x4IUMFxWCP
QjG2i37LoY0pfPi+5hwx7VgikJpSAPEZLkaP27xtlkUsB/zWc5gXU+AEpbsQl4WKVoOZor5QIX8o
JaIlgvMgSOhTtLIsq6MmLt7jpd8vpo/fEbgtAP3m6aleNhF5LaoAccY0tIdSJ8z1qRdD6Q4gOb6Q
vxnP8mkbGwdT/vQMqd0+QiNOek47ONLp7/YvAobo1nIV8f4QHuEx0MXuecQ1La1htQfQXvPAPZTj
E+lBg5EB1eal+rqJakexZ0mI4b/bBsR4PqisB/INTLzJiEsTKlCw/ToBsPEVj9y/kWsHIw+P8zWT
agufOyuHsLNHzY+jI4KA94qHCAvkErPi3u2fS2Vz3uytKMuHBdhFiD6QtxU0nFAtLripbRNNeVc/
s4QEB/gbCbcdY2V/AuVIPP5C0JS3vnKIo1Edk7On9OaVnKYqS+dW+RFUXjFPaUZe5Kx20LJm4+ge
mTJFoc+vJhdVeGOVLE1Wk21LDTCM0aZY6gnMbC9IFSn07croRcnHtNV1ygCCp5Es9LarV5u1dQ0c
dKvyTl+2LKhxauIXSFXRp+FpghRulewWthnl1jtLomFGvlj5BRRr/i03UC2oNlgmRY9mVfR2lNcG
5D1/42k1fvwr1X4lzlPKm/7UakLpBXibCAQ1Eyky/hTkdyInpUKzA8Ls/VN+hg968RRBBm779G2B
GIfeQPm/596jDwx5VH0GKvf6pgGtdaEPl/8V/JMRzXlYDsJ7UqxUy+CatFf07lPvuFeVBdKSUDX7
xYPNTT+Kv2CXttKNOIkL9OdWJokpehefQX11g/XtZq0scNKJ8ntP6JohgK8KdzOI7t0AVMLv5LxZ
0RGYM4fyWKLpF9Kl3c5O7d3pHiPBhROXEpwWvffFDUVnotieIiUst+uvG+gBMm6l9NDOMc+rQlww
qcisb9/TnyVfyATTaVaEUaraO115rzsPPGVwesr5I/D/5Y/jYe31W5WTKwS8sDlxd1nzMuUAGusA
Eb3UiJeceIMUXcLbSxlGy0WrREtWMiTQDErHbsRHu8aB9TrCUTzFedxE2zmk+VhcdwaMfztEtPwx
AV29RCzFTNQwHREWKfXihxEqeL/dbYE/Brg19yPmxLURmvY+TCDOKkxUf+G3av6IZsfUol5LNuFd
41GGHVNaAWj2IafzuTHdEKZ2eDbY1oWzvYc1qmF3iuip5uNYv9qefvfhFQa9crAPFIDopExWZCKJ
yqiQgOPmYuY2NtQ137yMXiFHjF60h2YskhRYJJV2dalPwIN1vxYMF080kgMZj4bsJyP/ULce+mvq
XP1s/8GpxSODG44MUJOuMD+lhWCzEKeUhuXquRNgQ2ulLdshnPS9+tcc+rkPMg/AbR2yzLu1tzDV
coyZvR/Eq1Fd7I5qkkJAHthAbUtHXEKpz16D+lV1JKCBpyuUb3rIK8qx+Wqd/vaoUCkGLD++QPZ1
aDfej3T0k2ZEsatOdUIpZArevmVfIdD3LVmq/XcRQf96c8X7TaePCFff6m8NynFWqsKAJqjs/nKX
AjqVIkXnZXNYBexRe3seAB3HUvDpXijjMENMwaMir5Io+chQAjIBJyF+CF4AAeWSWtdWJZOUz4mS
4FSdmi3WdbOp/z8gNeV/ckGmakKKExJ8vb9XwoS1PzMtPSAXFbmEosbmlAqBhLEmbf7/laB/2+Lb
+zc0Gc87eN67rApiIYM7Ab5osLfT4ZnEzSaYwy/tie4edIwCfHTSVG2mLoSKFaMIuFzDKru4b5ml
oPXX3t3uTFxzNx5gkCR9LWoAD+VfJGD1LhDNlZtIBO7ExeiiLxBE9wftJypy84Ze0NlN8QjAkF5V
UYKDNbt1qcPInywz9mzlvPHZoRi1ViCltqL6brVy8wCKk0cSrsNbd3la5SbwWMyiojNMiGF4qvHY
5h9qZBGGyo1UNhduMErAYPwufvBys8fYONAG4/17TC2GNN5OFuxfpT9Ao8J3u3eDxAVFxivJfh7z
3I4X5PLiCIsfu39oDT6tV1qKnfsVr4gecuQ6/kfI6OgPdVlp4WY6h0bvuPtkSuuv/2Ym1LfAhWFK
uOOghjq9+kclA80XuJH93UxZHxTTnShNOFPNR8RQEW5+eCK5YOtTewynnTiy74yCnuoobvAlnxiP
2STIAvwvW9L2gSJRNfv/7sH2aX78QyNkewaXSDa+IfRveDxxIS/6XIlX7iWEB0cXWZrWeDyiXtyU
XeB+dNRPjCyugcRNPuUM+GlIeEWiBIdSCO7ZfTW1qWNiBOltvkwBiHwB0EgwAQFeUmtahVbkpclf
MCn2Y/gRwuj2MeoXjhZ4JKwAcNGTDEocQoXpsP+kHBf3v54HwhAYoLAsDlKRJb3NBe8JR8M5f2gt
3hbogwzCv7Sw9y5OicSQyZPdyTctBJwc45I2obZTlzvwioUHU/17Wpd760PbwyJvPyY0v0NRo0h8
I0iRk35DHZjcPOzbH7A7OPLOqCxBCpJeEozlrzG/b/UUTMHFuNrdvz0I/qHfQSx/DOrzV8y/3RnC
sPa2iV9lnOL79S7lEKzkHkxRg0tP82kF4mfOIr0vHyiRexrXsGkwXgrREBlz1zNFwzs4n8F/cQPq
lGkgeMKjdiFQlqd15TsfmFZ2GScmyhzqX/Nz9MsMX0fa79K0L2NuuPY68tbpWiTxeF3TTwmERjlV
kFO+fWo/bWLBznMf8n0GeCPfgFw2hiZkwSa7/z1qLtYBiAyqBh4OsM2KRLhjJe6nOOfx1PLyhKLI
PItOpBAevM70j2bfXuioiSAtMCWK4NSg88M4IzrgZ4AxEsOKsLMMQKNmMnt1MMNhN6QbEmISZ2l4
2lRIdYb7qiz+k7I048//ttXuNSkz93RUVoo98o0M1+VeAeBIx4OG5MD3kN0pFg03f334W1u9iZxZ
6JtO5I3SvsEy/59kxXHCNewTuYnQ1xVsr8v+UjiPMaobicPHKewO8H65Di+cBUowx9eK+Ymn+PMW
41yWo7bO518hvkntlTYZbOgI7FGjZwzTTfPiEyeoiKOgobcBGVQNw1517FXPljnZ9+yYNZeCKM9i
mUam+jb5r9/ZS6G6XyAyh4f02HtUOmKCE+G61+TQCRVygwoZH0DZi40zp5wbc5ymmF5BqvUUhyb6
9BU/OTen3tPKWsn1bq3hghT6/QcXXLJx1t24eyZ3vSKS5yheqUmbaE8VXEf7PIq3hiP3OXPch7Dc
FuVV/Fkc4ndxvFYct9n4J9i08uWdpmLX7DIgKVKxxpv8zUmX64kaxujkZHLWAAmhkTYQDVv9r650
+EdXqDJPzfmOiiRNxsDKGAx444chhpUbZ/uochry/ic1o/HABVNu+wvzfp5AyAc4KlbrIAenYcde
s5C3gR6qSKSJrVCdLQwz8kzK24+OCzn/xjHnqWYZs4Kv89eafn4Rm/i5XzHuiWjPVjX4/HOhw3uj
j9mFc+GIF1S+73n896ibMsug6eJ5hlMX7uzUrdRjJsAIbLRW0xUJdOK2qjEtcM/tAJR/CFIncOf4
InVLLh9IMUHOOC7gOM1cVgpb8l+iFxpNq98d1V49RG27zFwPgyb2uNIwelgKPXzfoRtMADak5D3e
9RU1dmpv+uVDtkHAP8RDgLeQ3sGXUROtDP/HZDzfS4uewaCQl06TtuEYHPJ8nboNKTkZkpvhALni
50oYKvOGygD+MWU2/6XgK0f0N4dyWyYNLxxYBv57YPxzmhmAzVlDFw/a0AK2UP6TYuSTmElIeCFO
Bz0jMGmaWowp3Or7ys9GfCESFkwA9KlYBT8i4QiwStcOK4q20MVOahzhPmA7tVd7aC7NvX4MWFz4
uQ/JM5tfOiAW2H1kdzV81j3KOUdO7G4/DKpO6PTbMs0epOBKoCxyud6atuXe0APpyk5gnWzcNO3m
XSD7HeVU9FUtPF1qfBbOg7+osl+CC4wV4CzCzS3RkG3jW1Q5vlD0fzlvgydmqBFPXTBd+KMyTIBg
CpMjvqn5HJLsj7RqHLgagf4sLkirs81+FagUWjhpSGtOf+8e2Be4rhWsHrAgjH+B8fUnf9XssgCE
IWlOdAp/3+j7B1pUMWgIT9rOr/9DzzmiFAg0T8K8/BAGMF6ROx9aHPtGiINBDTO6fuDzZv3VzjdC
rnF0e6719P2Fp0rp6jnfC9nKYSELWKWhp4Xj6f8LWpbJyTs6NT2ILTdGt3cBf4E/eyR4O6aYKcpk
+N/zsvJHMP0SsZ724VKdWCBgbbJhbSP3+np/D6kPI0/UiusKroE2oAEUUlpWWpAbmcqDcNhstfJE
fX/U0zQBcDn3IyfoPTYUXsAX+ZSETUtXCxfqg87e6h3x0+qybxf/ZXWN24l1QbZJYXMS4SlNb6+T
Koh5sO/hC8vHidW8vSIZFqhyDX80JB/icsBYCBD9zel86b0bKxeZyFGURVn35Bq3MigeOfgxz3TJ
ip9PNQElgFVbfLc6CRonR6C7apOdxvX/Q+q1w4YmGNUfvrZ5guufsaEf4Gi3qEs1hvgY2ZtnEOGw
j/X3GUoYDvFXaLMJkIbeQnNfzcZN1/VpFZfYN8yJNRJNQxHJt0ZBXCFMIn65D5PkBOBd0QxYZ0BI
r3411KfMy6quMa8S0Wau8NOczjDa4vVp8XzCggY66Eqvzh5raYR8EGqcWKkrTMWX89pAcezRjEfT
uzME4JhSL6KLqF2h/mN2tb8LW5eHcvkihF6AmDH9/knXjJEZ0JxjoFPs4ZwypEIqBXYJn9hzrY2Z
eIn1qaTXgHk39Tt8MAyMRR2fz11lis1hfBoE8k/SbDg/boOQebm8KwaCuccbJdgdXxjjmj6bAAor
K9DwAFvktfshiBnO/LPWIw+I2gIFwcY4yN0rLwWnIYG731pTJMzveX1xAp4BsTsLU8LFMImCcTR1
5AG3sSoUT1nMp7ej7dAL3DGTKjamTz2HhvNJChbfrCH7kHeg9ZUoURLIAnZ8XieFmN86gAcRwc8h
Wgy1KYYZv/GT71M5B+3bXHhLfymsz0ggVuipJSQF9Cr1JbU8pUw3EtMZnkkwHBBqiE17dznDjhbs
OI3aW8A+OiRzrzckMAVVvSTm0sf0uhz+pzccE0MNuOWHUBosZFzx+/zNek5NCxMwSyrJOKuDi+KS
VzouR7LdR7dj4rZC23AhLz9IMgCn4Ta0oWB41Lb/dbFSK2AMkYZ4Ti4P5Ihs3cbW1Ssw1Ks6F9j/
eHkiP1/mmjzPDbRi+lC2i1bEAmXIk8IuUJJHEr33lT+jgPb4kFRaoeXpx855+uKvAshGqFDMM4FP
pgFgT6y5W8GzoN0qFp1ctfIUmDEhPnkfQ0I5WegtGPz+AO1ChqAhazmt295xkt0C/U9WLijBy1xI
cfSIy46rAJWtzfqZJsfV6jGMwNhQIbH8ktTUW+DsyvOBMSPCvlw60BgU3seuGTv3hZBKsb8VNHO6
CeLosXtpg1c981ybnm00Nxv6wn5i7V0Qa8gwmVHr3NhTrpyxaa9JrNUCRMZ/eS9oZq+2XF+ZaMbW
55N2CvF1ouxhzCwEzBqgir6OjgV1MpBa2evG3T7QKa74VqNW4OxtsikTJwHUhkFfAGk6pwGvHBxf
OWvMYweKalPuRhUu1HJFufkHI0TvL0ZxmJ0rRU4JTEDo3qOQ1TWJ9LcuFyqJRQroe2D4v/ONgZf1
YdYVYJef3swSPRm2wWofgwtFUwGGOGQB9Vc//A80iscN8JJYpMdMr1x8yt4CTZMPc0m+a7zLgbpq
jKZAQensFUFDWMORkr4xtilVqYogU+IV2C28N3dEshYJdFave8WrHuqzotkURTxBiJ6zPqQoXrqY
sAvQzWHTu2/6op7IzOWr9WCt/fOirlMxc4o1/6vRa+qvYlCWyvySqzXj98eh+7jNnIJu/jojHuwP
2cg37GqZffMTkpc2FrbfLlmHttK5ymAq2UifhIARi4tZ2oVysf9bCt00hdAekC2cpCIfoBvVdt7t
DyLhAnVC9UlCpsoHb7wASuswUmIjwMM9LzwC9cawE+B0ya5f0iZnnN02gi2LqZBoJHbf09gYDQt7
fUbr7w2Iku5B6t8qooGrTHdSez0tPXYbZfWsvpzkm3oUbITsA4qcWjzQ0K10BXJk3YIISbGEUOSS
SE6ZuFqgQIbxE7cxCOlkmpBkSTWBejeU+ScSC+EQItNyRfetc/2XSa2X3EIWfWbTUwT8+S7EQbgU
7hKeCSy7ej8tmmNUALqXOD8kENkLFd+tTa43kj+gk6z5ZkCRJF9STEW+grGrZa938ezfsmx4mF7O
d8dAUlpBWS8qxFNQglMUi/o449cGaJ8EO/tUTTwHi3cSAuY4Nmi2H68ggIxaBlXH6ShCruSJoGqT
vO4C0rmdo/VEz7SMu/uDrRqMZsucV2l+5V+JF726iRLAduwyKF2iX5YQG0TnALR+KEdXp1cthKrw
Hi/PgpgDetA5o9loaVBCgJ8rqUqPc/2zFg3pspuFrI4zRY88PB6h9KXPtVWpfurNUSKhc0SDFSUW
IOBuYnxEktDIkM4qpsApuYXZsfGpwEApdyDtUbe1Xlsc/kVsYb0Ud9eZJ6rCc2K9Zi3WuibdsN6J
TGOWITJu7nA+eHpSCiTFkiJiYUadiwotw9fXfyzqT69w1Stg6lIdAJbFIBqOx1pF28iQ8qBxoFnW
n9f3G57InMlW7qPuGN73vMDtEPLFstWNFziqtloC2MgYdEEwL5RZPWR1KGlRjF1CspZw1onBIP2o
h0Hcos04mfc5K8o7mu2d9ycp5tAXlGzArSkvIKPCjLpXW7Pq+A+HcIsjIeNw69sLIoiXgXAB6pr9
prOsavjS7HO/nqD/S+LMKNPoB0HPNOXmB1ac9KWHNmHqzvuH3Qf6VpDOYnpzc7D0oV9PyWGEoiLW
JrSnn4knGU6S5hwCrUHK9J4q6QamxUqjNlDA8FMXZHyzd2m3ulvRlBr9qDaFoUchnBul9MUSQags
Zy9DxzyMM13GFSp35andmL2UyLmU148wCmptE73cocKX+RFkiB9LcEuV5pKUG/8G0k3yZF7nOnNX
ay6bj/Ujd1nM/bovn/7jAHDlgKeFRAR9+Bspi9ImEm4nB+SDuLqUBzEmHkxbW/Kw9jNGTmBV7Xz6
o19ANjTzXsUeQP9hQXadPKDhmnTxfRbxqJIoijf8a4uZAqm3DwERIeO8GJ2oc8z64hI42QgbHFJs
VG562h7w0pOQtFicHnwwM5a2NvGkxqjcNVY4ADSehnp+d0l2nklUdBdCO76ehQTgd9pJbAWY0Mpn
PI2R+4I1eKCe0PqGHUNdatGvrZUJh90xW0wtyLN4KGKtIh4wo2fRiLRBdDZUf87ePn6Ocw6CPs0Q
+ZJd4662PdJ7UXlNnNk+jGKVWDJM7AxA7DpF68iM9iKi17bUuGTMxeqo2DsdTIUrzJxUlWCmagvN
S9bw2JW6D6fPcWkvnG9h8lmfSwcUHWKsQHqyHBZefBhmeuei0ftysWegmGkB3rWZ2ZvXMlIciU5a
aYzn8vKFD8mRa6FEgdYy/oSAtgjt+VyOazm9xiITXSTgq45xfLQ8FAy5ILWGsVgzmVjoMuozmHEW
wwePWreMRhWWPik/Nw8M1Ao0TGtbL0TN3Xh3I2mrmH0kew0b5X5VUGYqXnGUMGT85uhRLxrNhuKp
VNvsiQNgIhNWazazsLq7yA2Vlq0TARP1z/DiyVN431Core4mCbad6gMJVvvjwwfZnBk4hM9bWRr1
eVqMOjfPdZRr3v+/TcovRVHlM6dka70tPju+fAdgEjtClX+I54X4ot4mGwbq9RF6vMG5gWof8ZOV
FcRNEpu9v2gsR0E/5A3xDjQiA+pE/v7ifviWy5s3HtcHsIug247cYfqGD+/mzjKAn71SYJnF9m87
Kbw6LBgS/cK7AbGeqv/UJ8nwoFpkFbXVOfxV7qE5UjYw+h2SgOFeUvxkRp/rGGBIz/bL9oSzXO7W
oDWLpgBp6rataiJnni+P4Ugu+C34VQx18MGnc9Msl7rn8vtS6PBK/ERoLJCGPL5E1RW/5qvUaZbT
jNkuakUkv6RiZgk3RDENzg1NJlYym55wBao2deNqzNRgejBGJK0215bUgCMdKe7y3Juz4NrOKQ/O
au6FMKB7Xam/0Zu+3OOufWYTf0AApqpzx2/lhTHq6mJpKVX/ZM4T1UK96Ql93VDd9WjEMBV+KNfy
6Ccn7RTcOq9+TlpHko2ZfH/ZaVZllS25jAGmlMsSx+tcFcGABdI5O4UB8ZtWeF6xolO9IgYbChzX
sO1g/FYp5gcFBxbkPoA2LO3i8rowg60y6WevRvL8L7qiSAQwQhcAksIDD5nmG7YNJOz4vazpoYOP
zPtgqL2HYVQdMQuVbB4sMylVisMtWZaHXhsxP1+KLienbzds3EvU9J+zomhF/JLrI4lf/9O8Emsf
dcDjciqhsmDZWcMMT66KlXYDWW6XimuVvpQAc/9nMQogfd3CeSySYBfa4eWWsYReTGksPeWp3ZqX
lYWaWbVLzXsa77rkaPSwMUiBxAc0KYtCTvq1SG+0OAvPwmpAR5NH78caLGKmmrBNj2C/BXhVqRVs
amjkS+3GBvxZgKsn7bcolxxtY/fTyvih/JrTb1V7vzWcFyroTrYq1bcA7VoLSdDb8xGs1D4GB3kK
OC3gsJh6/nugu9K1Fre5PrrWKn+s6WeSOWUuB1+/6MTlBhSUCC5Pk8InvSdVCI+o1okqYThz8y7b
RMbJ0scZXH70xGmCN5ssB+7xz2XN9eyqFvc4XnYNxtvrdErjMYZ7MhLPJzU2BcD7pjRug4hzO2HI
I/YG8JmfF10sxhybuZOABkWUGXpigi997sg+18oboVObK8D3SYSf2cmPrmbb71gZsv09HNYM7Y6K
JJVpaAkyYWl5+oT9yWLbZFF824PYLCESMmD9G3PRBCrpBp/QFL43lMSdqvifvTwKbuUfiRObH3DF
hFWfy8ULjWakfWYao3xIGecsNx/1je5lzNROP7Fmq7jE4Uuu5+D29eo/3UfyoOMPDCUY7jB5OguN
69ooMUa7wKZlrTx4AuRVsXloPEumctk9NYCNjcqvjOJY78BXqWs4Y1oa4LN/GouXZHd9L41ifx7M
ssSqpduBL05aGstQdNbYqIvuvboG3StCv8OiHuSHZx9KWC3RW4wAhSGrzM9brdSl9L75h0cl2cgr
9Bij3OjeiV68h7wv8GyB/D87dAEmoidWRunjR0rtSLUOLCwRTvv9EHL3rhN4RyHpGnjE9CVsd+kk
rPehn1pd+KA9fqz6w90xejBqM+qJ0gAtIo8VCpfjuV4SvA1P2JoYtuoGivE7mY9tctb3CkPKhsok
L+0iX82cgGCAKxQxFIBfYLK/0FZ8A5MviGYmW1VLiKz3fEakW74qQXC8qVt8WhDRFzgvctXWXiY3
tQmHz+s3jlxVk1F8OUwMJGga8nxbhTaQpS6vponQrvO9g6WbwtZZO2Tx6sz+YffrAjPVOmrdn9x2
mnRQp6O489WELsyI2LlZpmewKUY+6OcHrMSo5v0GM1snxoGrO8+GaDlA77nEsAiAyWb//mCogdGF
5Zn8OwQGNq/4yA+lukCztpQuSG4B+i0930H4BA4MUiU/9hTmjqWLCe3nNfyJzrgg/ZdYnFtEBrSA
/LUvWnNSzaOpsNv6uJgylZL0xgtdKVLEP0HepoFLx+ePxzZPtb8Uyn7cNTXrFOMaJamP/MGE4PCD
IK9HoD60u0SlfTgdGmt9NlPbG7CZcigv+3AJvygXOvnnw0F2Ux7i/iTrE37xxwzYDRV/06MBKf4o
pMBEizkGYnvJURge4TB18jqofiVIAsHKy3wQFOqgy2ABAzJV+lR3rCV7jlvdFDktkwnCu9J7kdoO
l0nUnHDsIrp4LObtO2xUvTPFCIqb3MCkZ+BeVAaIR0XUtMTVc/o7aOqzTo+z4sE764jMduGDyVEi
AblS7vPys+LokcHl/QNpwqWOEXoAo1x9VXYZYNwgmqyj4PzIv6SBvRuyGkoLYSMKEI1fbf4+9nKJ
BjdoTaTtSiSYasWPDmO6/6tsdglDQ49zVbSTA9Yv7/zGXOcep5jOBjlyFRd4j7frGbP09+dPnCSc
Rp+Zo8T82/Ep81Gq/Yfoa7PPT/ikAuM09STnaUsWjbiDzPI9N24ont9Ptv0JCd0UtzEGjAKEUKqe
BYM8DhuZ3ZiiKNn8i3eCP3jyX9UcQ+UuFpmqARgsGwtOpNyEz7ChsviTimvajQMakzSaMzb8otBq
O55GDNg1Ddah6TeVlGqAwXnRJSxw6SdWLLjOSh0tuy0jpDvJw/CB3UNcbxB7jLWMLUVSBELRb/sE
muPXlUEZQYr+2eiSp3Ch6mggVGUkvW5aC1QLXMf+CR4mfGOnMQNidhyRAUwZBHljepU6U4KaB7g+
kApjktHPWrrIVUawpUICPnuRTEdSaAPpsO+rjav7+4+q8mxQCt2vI44C42GpVqf7oyfVHecwO051
Wq0SKQATHHOtdO/rBiWXeKShVT/dnrw3IUpeMnfsyfqbtFzwu/+DwHYsYQzzkPLdhDyQOxlybb9E
trN1omXCWtHFLUavFwxdvnIwEiFfF0TMOj2Zs53qEf/f9z8Vew8YkJ+VOCDmdCN1tLqoCwyfPwhI
VnfG0lO7a7DVLJorEQaLWLV79aGygRYfyvbOJ9cXQavcayRWZhgoDbViVMW20W+71lr4IVkgPhwo
9A5Y0zrwlACvPIOJpN1gSC0x5revorMfBaYtfsCn9mRPhIraiDvcRTEsCvzG/TY+RiYWavKjD9G3
NynqS7w7yDaN+xg3+14U6GSzvzQgcnqrD46Hnr9/EStzFwwB2NQbewrtXz/GvYoF3WdPyvQ8h6PT
L38OrRF0/ev9OHXAcUT01LCcDW1yDZtI7jorwI7eVc3oW4yspmNM9vmkX1RkCKRkndWomb50JMvI
cuulPAXLNuHTBXh0szLFtQ1tfvkfpIQMo4G7xqOcN60CiG3KSMqCr0wyvdJ48Qmi3OuWKr2L/HnZ
oH9DaU75ramuzLFuzTowdHtbot0y61f6sjvAKcNJWRvq83IoOjNCdmopGH/c8nqdF9E9SImMaQU2
2Dye/HsB3t/wKT6wGJg1d/lgRy/AIMdpA3zLk23kmDniB/f1MQcZEzsbcI4bOp+kHEK0afhxB9yx
5lIKgIygWHZcPmcGgflcNI3qgkg/h2dHM/38+Wd7cIeBUlFLRr7OviEVx8C3YXV7ReRfkPi24BqP
Y+ceHnMt9FK23BFfNXI3LlUCedg0297+YTFdog1nWMdXyEE/GdwqB+SU855SU3ngFW3Hh9glQ9lg
pdpV/7TqRmiVqWe3UDU4sQsD9+xh0OVkJSd3pQQjdkKurXAlUyK7y39bRllndHIKFhI7xtuayV3Y
Cu4OTNy6lKTKp1I5upH07RZqh0pN3NBz73Og4x0I4y+Ntov48s3HdLqCvhMmK9BrGR93OQQwoTzX
4NbCPKrm8ugyY89p9ASHTaJll7VddaqsY9TFd81QMsaWSN1cXBrN7n8WWlu8yQmL55tvLv0/VdU6
QFHmlBpbokwwXpBHDb+6CBmJ9Bobr3fJbeFuvgs9HjhzBq04w6eQh5nGE6yNjXL7SyQAxJ5bDwrS
EZ4clRpC7fAVW9u6Be3PT6De3Wd+baRVt7a6kIAO/KAM+PkiS+rIcUMR4RdiOPs862V8yOFO3GzS
NDmsqedgSW4CVf3ZArR8nW0XRS/NzyoReV+XhJ5EryCADRkjJkEGy2nP+ZWZSnbTtAwo8OB9y80K
eDc/6zd/Vo2xyAGibD5jTXnGwKk556Wni3O1p1AZY41Rqnw0V3L+M1q4OsEfSpWz3SUXuNeoiKRG
23SjYBjY5fX5KTEqwfVkYfDbmo/tTIAOIkSnpqFIuUlIDRogw62/8rhFzGyvyqhSQE2bT0Rh29MJ
eruZ/wqhDcYZOJIb/XWWUxtAz+tjT38nRPbKpHsRfUvO3k0Ps5aZSl5ek02Ao5QxeL9Oc/kGxxDq
VstbZ0uOCCuBF784Ls5MkyC7O+SQQ+5onCD4YShfrTzM6uhQ8qzeynpGlPvkO3c/sFnGUEPMOnjc
UMyKyqj/oigLfwIZnO9/FhqIJ6b3Vl35JrZZbaX2RcVQQ0fk41kulKCrYUofs3KgaeIbC4iweYN/
HCc9lUIh7xAhoMA0sQQm9EveOZZczbJL7LzYSZnFpCMpurtjbr7v3Q9EnZnLCLr4cCdkiG2NVnpw
7b9cTqaPPH9Evlx+zsFhL5E4m4yMp09gnWL4XWTtXYO2YsPQfpG2+wUYHfP5UwShgJHewjMh5iPk
3oaONTSxwbiPNmu65yNyfcSeHi+Xwnec+H8MxN273cw0yBZT1M6JbOBh6vk5X03tKDQ/Mfr/LJKx
y3BbVm1hD67nCWEaMQBfGQiG/nbXRVKRVycqzqnWZSSJr1wqO9Gx7sktRvfNM13VKTGscvpQL5n4
lek8KpkM1LsA+PD5CQL4sOGvnaTCbuOsRmGSUUzZUevih/b7CRPR4dl7TskiP+Bw7gSXlT4AG3Pa
aqHQZazLbEkvSzpKTwa1uu8J4holTmbOEo8M48J8nS4GO67cneChcLpfyWB+pf9Lq3yEZkV6gllh
x26Vedao+3DJSkKMMm0hhuA5IaSk6S+1bPzjqxFt8brDIyMBOTarnvjWEwPKhDMGYWAat+zjitU9
WeyWFYnnqi4YHFf0fIqJU4YolbtTy3zuXK/e85kP25N67778yZZH8fT0RT58b7KMZ5DfzuokL0UP
jlp0VK8Tt/2GOM8ygcl1J+mKVUoPFbwqMQg5RBQWPP+q6WD8ReiEQCVB1zF8x4IrpEywJiZywzJV
YS68XSbAtbcjM2TBDYaUBD+M7URHUZCSk+7gnGXX/BEXGESrm/WdJs6mBRwXQGzwUa2omKdtGw5Q
kDAfS+KuBQK9ucQBhrr+l9tokoDah1O/v995U2pOzRYeBjA47csw+Jdq8oypcsZIALJyy1xCYdad
VsOKIvPmqR2rpl1H4MYrAx8RM7YKSKaZT0jOIXKhKVhKaRbdO2vxUXLxLrHMmSa3TXqpqpNug3ZD
6z5okVVU76C6s22Awrtb1WwYDFydBahlgOyPO4g74YfGqhoD/qIRmIwmDLO8ccn0eo3CLVPKIkH6
/KTVY97W/XJQe9pXefNZfH8aCPtcPTUltOxpug2i5qBc6OEX1MZRBEdmG3xHOQyZCAbcO8mBFfsN
3GOM4Ptgu83JlLv3BvO20J/v+AFCeGMx89uGVpdE77Q3LyR3QrvOkUb1knpGBkqBOz1t/+TPIcV9
cviP5tn/4feGqAhbL4FF6PK3Q+02e/O3bLOfFBuwpqLoGhOQMfu3zqk+/0v43EUv0rPuGl5QzzAG
ZPsYkKwEpgDjxSNrW+SUEXUA1IBeVthH2RTpeMN02BCDyRyyXyVWBZd5SsVFb+GVqvzfMpaWuCAD
+Xmu69/aAh3s5PP0ZXgJjjfa/oi9L85XZ9dvR2yElfUf65oiDs7qZYR8u1u/Rx9dogdaJdMw3wfJ
M+7bM/4W8r0p8QQuNOEwBDMKZisYKEwj4GJxtZAU0AqepSh3heLVpNMYmMUiH3WJ1VxtbWPxIAQl
Jho72EqsngfE+eC4gRyhIT3ySppL1oirsEa7UXyMBrUFNwZuAmKJFxAfZj6Eq6xx9IZ8qg56fskW
wW/E6+gJA6Iu784QRe7aaCjUWqV0D9W3AX1YxeYzEJ7+nnezvTThC8EICDYk9vWqluvSeyGZOMRj
Flx7upEbVx1ccYnreK1PGtNi29Eybt9PAh8zG53QTCp9jli3PIildmsA9lxROq33/1541pLP+P5K
hPbdLTZdEMubzltI/cq2pyEVk7GBshH6Jvh1hTuNq7hOcMv9Fo3suCrsiTLYlrE9ootqTt7o9gWe
X/GXHFe8WxPaG1M/gE982gCtCt8CFJKocA+4Y+XJmeomvGaonr6g5JHNV5DetuzzNaC3XLAqt87q
yVttQBcl+vnzMUUAXzbkq30p6cc8asLv14P6/+Hq4MSud9KQKq7AawFaQZ2rxp93EKuVUeiydvMC
5oGC2rcC7qWyQsfZFbYoDcMs7rLgWs/q+ia5GBFfr2hAX0qyD7RrK2379ESH4rMvXf8GPY3cO5R4
h/MU1pz+9nrWE8qkCEV+WN4Vk5HiOzinvWZ4LDK+WWvzlqMyOiMxF4pXIVr9g8m3S25YCHp8ehuL
gFHgDgw9LFJEvhI6PqSDxpUu66b4UaLoVnIQVaevTrfXtPg0pssVPUXUNrgGrKr4nTdhQ/wD7En7
Z1gxeYKzMbX2Iu6EEI32fd8vWxmUUtHUL3Rw/7X8tfHfugwz70Fwrq2C40pcfQy7KKWipI8BYqrv
vm9J4oH885asbWKzXTkJKppSnBSAU0GS05wGaMm0dhdywyfS7oeeqLfn7c7zTOby8LI53u4wZi0H
+EdB/RdQtyBl7Mzmv9Nxyb8O43o0NMFnmRKCPmjnQV/QhUGQCae/E2szyLg/pJROpCKR3PGW7JjO
7I4IkiZnlSVcBaK2Uu3K+ZTkswxlonGnxknMYsYycTObgJN75sHJezNyWrh5JJM2Mj4DPo7Rfamd
o4wd6zLoimFm8lktIe4Q6gNQ0/EunA26Ckc9BW6dbysk3GYFUWtjJMHgJ7R4jtmYyiAIhS0Rp8ts
D9EIk0Nn4J7bVJ5FUnlbyXMR9gdsgcqKU0RxvTqrHEZ2XgFI/DZO88p3zrGKbmyuIucCaPN/H2KI
mlHo7EfKPHMHWUHPFEsTx15tzqwqhLZ71FlRJ6OOh21JjbQRi9z0nBwdvwFcAos4E8ftHAwjtIJz
X0PBPpbo1P6I8Q6rFhdJ7IP/R8IcBERNTlZ6T8KtA/oOGoxp0g0DQgu16dyIfszhi/5DD40tarKZ
3NvWioaPuc7INJUktefrR4vlcM186shZXMZWTeSWwNU1gt6qs2YojCh54qAQSARHXll7zFqCn5rE
wVSKMICDzS72E6WM/VrY27UT9DeOuJPRtAoyJNLiadET+oTd5g7Z+qcZkXHf3AO0VIjLf7cQ1Q15
H/I/hrOzYypRDoknMhIzbXR2gOdreP+OBpkbfmtvE3NxcOZKn7xMw+jjEYnCjtFEhn9hRIFrrpY2
/FWpAa3PncRF9ks9UmNRigVRU/sMTiB+bH9H7C5v5L78CQ+15iq2nt0Z3R3DiTQNA6WaLBkqB7FV
s9zc/PAExVaZOnsY8a/3+iYBnNqoiqMO1KDV9IJOpboctSdf0B+4ARQF8JQdNbXTcd54OJBCqQdU
hwTbtuuo7acERGXp8/s2Nja6WloEzB+9VKH0uQWk8Pa+HEZUKTrC2D+stGqwUOLD6EPPNi6RXhtH
O/rEcglnzI4Kp4wbek+mU3pgzFJwXOBQOLEr5OeY9XXUT8p+xwR6MPgIwW5UvULwl2/TOSUfVzGZ
a2D4YEqE/Rylgu7O7QyqJ5FJ7oB2DkpAJY1bXuSwP4cqu4mAmKcRgClPcYcv8FnJxk/wFQxwcjhK
eoC7wSL5SbsES+juZk0gaPT9BmjsQHgc3TNhvPsm2onmIy1LDXo630OWVWfa4g4qCcVA6BnEOYNr
DnZFIgY48KcWl6nvXszacMYafUex0FlZS5fOEyTwA/yvkFjK25QhRsl8bVymhdC8PONVyXtAI+FW
FfAT8DB00pb06j7erMPgNHqlf3qpFifxUAClz0BSllBGteo7kgqDQrQmNcjQ61l2C1F6vfEqrveD
+hTtoDaJQL9ghMMavP+CEzWoWpPK13OyH2HJOJEe8ourz5TD8RXbZfL3Sez9SKsdLuVR4m1hX4TM
MPmTOeb5YeSTuuQM0RauxyemakKWVhstBy1/kpMZOMmC5l1XmcNdFBGzlALZb4v7w4ucM/tHWbgo
vDR/e6kuM2YEHV17qWAVR3i0Cc0a/20D83NOiPeGB3N9c1pwQNj0GBaY3JgWt9ifkqkXxW9F5MPt
V93zdrUlzvZ0b/kPhtpiyPSgXMsb61VBrCkQpncO7ju4j0cDeX8QUuoQ+44Hi0nbgvHnemfWRIYg
7RFnT7vNug2giuJTGujxVOLwGZa3EGn+lCFnVJQznyAb5UTDOzKuMynarrEjYeSMb1/yve4KBXEp
cC02J2OiiEMsZaM1JhbEDXxeIwhfouOnZ3ZkSlmo4GNzk4w3O0YOW38f/1rMK7WjBnomTJR4k1sx
yiH5SJdpdxB34RaILrVjdO/c/BrGlWDXhHj2gp1rAPNJChhwpFgVwSnofYL1uYx7ziErWKuT8gLe
MowKTIDn7YJ64nJQAL2p+Lj3Yf2kUZ6ANgdHFQZ1nsuNMgvkbasv1Oasx5XoVZKSpKJ+CL7gcdco
BIUFNhwcFab4769vD9mwLKdHzsmdSIP+qvxFtklQAcmJzNUkX3evYlW3ROWnh/TUWALOO/tk3lo2
f9arkHNV7QGmfkHo5IFwuvCBEtEJOq2AKLvKaZOBm7g49HntK1xaXrLHfLOIDy9P24XKf6sem8pJ
puZoFP0iTOZkjColUQ/ZQ3RUSt3gfj+Qhs1a0pzvPcJ0D0hJkqPb50gHTqwF+7Y5P5tAf+s4vRbT
vVXpQIEam/yoYMP63C6DkqeFKsaoy6dSGX9hB9ZAwAZb3ua5sir/bWfNMzY3Rfd0wsC2Rtvt11v5
TMkFKuxT94H3hx5v8ibpVwK/gYcM9oBOag+PPWGKmudRrU775q37oFmYlYtLrM8zG+THFCQBzFh9
VEPru/uag5ibKzRkPZiV7b7VH30cPwTTwZWbrmUeCucGwfdKQPXjf4zjyb4qdN+l2WJSTkKqtCg8
0WvW6AR5e/y1txlgqZoISN+T5AWiSxvvdIf2VvKj2MrihEFUzP2FJQzm6zyW2YfOdRJCs4CXgQ10
XSvDvhdcbZz9cyemp0Em5ypTN149WuSnuGzjAFO95+BhMlK/L7CDpNd/98DUWdgFA+SkA+uj0cS+
v3aqs6JFpMgMEFkTPssfagbZqwtNrSpGX/okxT7i0GaqcRES5fGw1EVNHUxFuD3MGvL0Fuy+C9Lx
qTFnVsS5c3S+OL9eNnCeOfp/Ux+/BNN7aW+3/vMNaTjcrNqlqHNKXRazmv2yb9B9V3SVrXRPtn+b
G9gbo5GTJCu5dQ7LCzoMtrp5KXAoU7iHxHd4JarSkfH+gPf7L3hb7ELGUvIG8c2pJpyzzuYOMRtL
/7pghdpy6rxxWqnfzqzSm1Ou6dcWd4NhTFEwtiuaAyM51KEacUuQYOpOnYf0+HgCxcWHDZHSiiIB
crIrwSF8HiMfg/xjJlxR6tP1VVhmG+eWLn5UgNcJeJa0uiTREIkONKaZVjCXXGrRWuepEushVG68
VYNarW8uBVOAamc6d2++nQw/epdreLpBttcRHM+FDDKw1WhZXH16rolPf/e6teMfVftUbWkPFsuK
5daQFcM2aDRJWq72las7Mb/HOdNS8xPQcfkJjkq6rLZe0UhEUOrBJyyj5ASSTWH07XnGWYp7BkZ3
OVi6GvrwUgOzGYeMbuztqNXpVaRP1Rp83vM2tSNo1TmssmrEU/f3HVG3CO69qQ/8+UnewjbW+Gqn
YisntctM7xjN4dOKSoFGrnPmOKqZA+zDQAeL9BD/kwM0E0xnjlEI1y307ZVyNc9uI2MfoYyOHgDC
B04+luFegnyetjCGYvcullZNHzyaBmXh0cEUcVL/5s9lti4V0DX9V/DOvqBCp6X1ZzbOCTP/8yDG
TrJg1KxJhE1ikS/ZcEz/IgMzIIHzqPwwNSABV7IL4UAfoq4Ui5pE0qxphYlVskQ1Q9lSWDUm75F7
yUuOsS7H5TYPtVg+ucHIOsnedxqH2LOdMqucPRi5D1h5roaqcHBwC/TrkM1PAXqSyi9ITXbIa94U
oegcAG5BCPa3ymk6wvemj1S7RtDBOIP19BWtLkR/RZNe5+BtXkK5YZcccNIhn1hcd3aTcHaftq0N
fggWxGIb3c5yA/8At4f5PD+IcSLVVpyYC8X2Ndm0TcgZ6PoRrupv5t2GBIXTjulxbeh2WNA3lvUu
1VCaWIbSumWTYabHIG4s09+8SM5VumdkxgapWn3xdW3K56Idh5+ziXzVW3WhLgRGZATDy6PGjNiB
GwTArVej+PbLQC3nmkHLXouwZkq4jcO1T6z/P/kbzyz6OfT2IyM5UJ4DeNHh7kOrimlPjoA/oqaC
efoM0IB29t3t215t5hAbbRXR2a+ldS/Zn3x/bu+eJVNnsbTKMCdUWv7p0JNm6bTinV754t6jCzAD
MNGCcxluzmXddswkhNd5jdcjjrnoDjMRSjXeqcnIsGUs2AcijL9Rf3u2EfHrbOlIsuNZHv7uYubp
lYF2UvESipNfAzJXsMX/uExaL7qOULKEJ70Yv3XVTUwBdjgVG5jAnP5UvVANXdbUrggyZG2opOKU
jdqXaUK9mfBV6e2wVDj1o9Hwe/2/myhaOSBYIh7J8xHkKA1IBhzyVTnMVyBUEbA5bs+iZeS4iP7v
H+7nq/8hZ3pk2n0l1xt+O1nR4YD+8uzZzJoP6NxVlholSgXiH8qpvGpfS8UIVaKpnc7v9lPcjUJ1
7w8/EEZ5GTvcyWEK07DjMIeVrIfWBlvnxD92h0Y32Cs/AyEXpCEG4rXrbcZ5BM1IYpAPjB8E2WfY
Q5/3a7l9LjBKJlaN239yeg4fzcTFCfI8FzcO8CZ2xzJchYlvQWl86Br3fouGbU31JFiluwVI/ztB
zjI6i8GJoQLcwFpk7b20E0B1EEaEg5fVfVKkoAYst7YUYPZ2hUguYDCSCoht6pXl0KMifCkSkzNz
El46GDSG9m+KdWQd8KhwbSMZYodSJsXda07LHGJUzMSrUggUlbNUgJTff2Ssv8oL1cs8L82Q6IzD
xoAEGCJItMV/OE+yTMgmuoBILLZ6dSE1qUUE5YZh+93sYcSuIZ6f90fTKgFBIGu69HirCFVq+yoc
6bm/Epzo5ZCEMTj3t9KGLGY/mjW+julQld+V7jCxM0UZJq33NjeEfqACkVe/QRppw0Phr2zBb5Ye
/Bi42QU1VXCjG4s+h1QVvdP+s1GI6Uj6p5Zp3qN7bjaPFvp688qhs+NegaSo/VXpdDtGFMiaw8TW
25vW15O42uuibRAnDMYIdpNP0zxSgJAyJBdAizydKO0n5y7iGILaGd6gBKOSfkK0J6pfFaCWyRzY
gvUyuzjzR7b5gZqla4vo94ihtYwxrJyMDTpTJYqxo1k9sEC4gi/8auK+RzCYV+fvn9MuM6at11SP
ui0I4l4BhkrElLb8vPtkuqaaebv4ufHGFMgDDZv7nTfH0WsxhD3ixbSTxjFy3s9eJXRIjzqOb9Ff
E70G+xwmhLVikIOcNrJDj836ucgQoUFKktjBJfLxEBXE+q3lFAouxIbNfZsakUze5ISJ1b1fKL4m
VDAdM2mOJFRAo1OUTjLZPxK9/xXtKD/wsfQJP3w7LFNtj3EPE0+84nsXFlxQd097EwOJbrXLPNh0
30zHDFpI8fT++W7j4B+BRzl/+g+pxSIlmojDiTwuLG8PWu/Z9sYCbduNQtxQQINbPGJmIa6bWuCY
5pSZn642iCmdNt7ffSHNMFHN2+UxCR+XGV/bbB/h5cmSPRJL8/F1UmKC3k6TBNx4SyucUkDBWMQi
KojCVLoMket/+8cOAjybnPwqjXcxPeXF2FbQ+OmZ6RgJ1udR7jMCAb1eF0FynLtuAyMsjjFJgFW3
8DAXOb9LPg/oCWwdNpsLNGBEs+/C6OuTRkNov+GTTfUFIBgs6VD91g8Nj9m5kjeSFBfXsrTRUbcV
JGvgT9vgYP5wXBkObACLltbc1+313l7nUV4Hcj6/dUDQ8wxcqDkrfL6w/WFdOV/3rcv+vgAxE3uS
PrX3S2zh/VpMUbY53KF8Etbg9/x9CiXloYyxY9eCzRikR/Ws87eqct/Xm7l+yUk1GiSISaVDXnpH
2ni29KkKQtD+f4Qb5ATfZAfTuDLmc7sunz8WEsSdz1MMtZTYPlKRQnQpFBsqtnP2cVrb5qXtZDHI
QVyk0janqvnM3YHa9vkZFpMBH99W214ZC0Z1Trvk6ASrNZkn8ACwMzYxpDtGrkQrR+TeOaRNgD0q
DGG2esPTf6ZlsBP2QY4YNBrEGm3bTucHVM244CK8Zg9a+t633ZytxDYPC5KseIP8M8PQjsVRxYLp
RyWauVgnJWQSMFGXox0xSfyjF7cgDXT3ojCsYgzGMdFgwwuU0BiHGRdy3EvEayMLw4EHnUBK33BG
Yrc2lNaTTQRn/VfHtxTzjObBTQd+x68XMg3KmeXAd8PBIdKUOMPunc0OZvxrWw6NjmDWHMAmz6NM
56xXl3vVYwphebq7gZ3/mOfBLRQS7H2XrzvdqhanR115c03v517PyA8plJrIE2bqGkabkP4vwKsw
msr4ar2MG3bOyBgXb4Gl1aQmsfSFleduMlxrSNbLLxJoLu5s6s7UxdA5kegZoJQwjDx3sxgCBLii
Vz7Q3CVmCb3Ag82Iw+zFMioKZZbPXyf3sQgqram6t8B32M7VxVVRig0rlbjeFnspORoxKGeljJm5
oo3xG44QnL1G7HI3rwuI0IH9AURz3YNex8qrGjpMdtULHhdziKwX+XbnSafQgcUVRV9d88GWzYww
dMlyNcL3ttgSROl5TRWnb/Ag1Z+lqO1PMD3E3z59VdcXq1RDMdDTsqs+ELu9+3LJmfz3bjqP31ab
reuFEySir6uDWUfBp0DkigoFDb3NcW1DGk6wFE+EBC99r4TPDkt52bksZuHWRzuIz6Zo/b/vyLsh
D9cUo2eL9X2NU9nrDqjNxHEdttHh/CkzXbumAGMQZeX4bsmvrkd+dgmzE5r9ItdftFBiEC8sE76m
5eAeYmNrBgsEsale85KB3u9Wei9QTJW6G0gLVvuBXhCaIG4mW+9qIymwbZlAMyBYHQTF2lsKWHKJ
gF815+a4YaPbbQ+MeFD9oABVb0Q1NWUWD3Bnj5Jhz7VJN8Vf14jKn7o+6ODQxTBIO5sx3hQHDkQ4
+2NJhC2UCXiL3sgVHgKNB9j0EjnBTBoO1nqxIyj7J9uiZKXCdgMsAK5Oddk3MItAQQrrkCD/14VU
EpY6pDpYCF6zhwIprxFL0lrGBVD5d/UoitFpKrRRLD1riRXI2Nuz8IJqziAluhHnIefi4dv/4z0C
M6ZmY9+0Kjt2CzwJ6PgGTYnVXl/APO7QkHEW0f3brDreME8s9NmTidDnL/nrPLHoEwoZ6+yfR4nR
w0PCQroYvkzeL91fVxXwBVJgac4pCF20tZ+PWQEeS8jjfJtOekTZu1ZI5VNCffS3fRh6awZyDDgk
vxD3J2GZccNnAyXMKqHEq6pPgT4xWowQO9/LOt6k+Ku3VmLY7XbpA+/H/AAbzsvGd2IVN/hKW6ac
uHOW7Xxmb2TflatbS1LZlXD9VmiK8yKE0YMo6ABIUN31x/8y2/xZxyNDENSydWJi8icvvTIDCgkT
lMEE5uPCRiy/bIRB4sEeGI/fGC7Oyeq/KeRC6Lij5gepPlPo/T08pvknPeAOyt24hk0Tdt8zoYVQ
dmpiXA5JbAHElHcI54yG/Jxx2IsIVPj39F1kQf1SRqvyn3IVKv8AUA418iHPOSnKyjnOR5OWsMOf
Ga0XNrndmz9DS3inSzobG0ZEgDH3Q47vqxwLe+B40QhgYaSk40PPvbgF6P678c0GaNKx6iAeH0hX
iUBNZ92yBNE7r1WES3V7Ooj4fC9aCroFFFN8tlh9NdgxU6kDpeL7AH+BJ5i9IsmJLLzQMFR5gAZA
Em7OcmU0jEwr9zovuqjt4Az1KaynvdHLneCe7oeEWMcJvipNlaJ89xAszcTUKFL+wKTRbqWdVdLS
Lb3LrjhzU1f1DXI+KrcFmt0hfxCcSu0vjVMmLPrG+p5R1mOTuIpfzgIq6uP9He8L+DnGTeBUe8nj
Jar5gNXosg8YWWWCSYio8MhcKuftm55ErX+D9gQbp3zRdl3qYTlazzx/PwGEp+eztklO5tUt2QGc
djHD6YhXnGny0AH+ZJINvMPoniB1LmgcpLQHJsOZZR/5gREABsN3ZOec3bZ5IJPAYVCaBKSRTff8
n8rhpFX3aRMKnH5ARpWnRQX8NAjbsWU5lPY29mXcEXwSFMZMTk09Y7whmn3WSU5aLcAoY8bcclyl
+OhTt83UX5BX6vv056yD+Xr7Ocq4GrMHOLReGA9NU8rF9BcOxchqGiBwyYRBBeR9BjkB2GHT3/wO
9HIzv9w2LCKSChBgcrD1v9LYqQJ8YqBcaL6vJ1SG6Aq+2+NVSO4c/HK9x1MLTWNOgM3+LekfTjdg
9DowAIbFNA6U+LdwlBsd+uY1X87syVENzie0RuaWcPP7O8J0jiB+4M8Mg5gIv6Eck9957HVJ81l2
T7JIQf7Akv8vXi01I9nQ8LMe/8KuXEuDbKHrH2ludK+Six91eWaSs/3md9Gh1cp74atPvCRw6tUA
rwAYRK9Ar7NmdhBDf0lWfDimC4NpevYbgeH0dRzylqcig7SN2zsS1UDWYBaAaAJqHshzFZGAYqK/
SR7KoZJCglvlIxNqrU1ABZdyIx/PruC6OHVqtOsRSFZdVjxAlJI6vRDfN0r/qa6u1ZcqEdJxXQ/7
RKQacKrjgdirdB8LPEcgRfES4GTLX+46PSNZn72zPjrqlg7J4oU7Tkpob0IJUu666uIergYLf/XD
5n/fmlHhhShtnA0ay35igz2tJ0aVVFMDBqkebBxyAcqnwUPLonNiVzEJETMGSR0/Z4+t2qZgyvIy
rkU3J6Zm0lk0SzDi5bvZ3k2S/HtVUcZPQpdG+qi6biFUgVkLlhE4p9DagFwFp+Nh4yD7UPBR17hv
OMip04J65LZwFNEsuWj2NwUa384AWL3upn7jUK8L4o0iqIFfLpSa967IqxDufIqNLj5ujEtW6Twp
pVwNEPjOoKxjiV+XQUE97PHl8k922BvKQVqAQK4OCKDwPJ7qbeHzn7vTwbcb3++aqN27DjXT1+Qe
+pWUTXSe6kXI8z5i9tmSlJySMndZnjxxHwFX+z5JCwR/zo49WbuCV17H030SLhDoBW4g+Bw8rdJX
tMEoGPgFVL/ge2lvWBBjgTjNLZqvo9SUlRR7b9/DVekiJbz60RO7WrHFHrjiSYju93quFqMUF7ZI
JqEkP/HSfHSpYKqrRWxfE/CwLvJTF90Ja+iRCn2fvXG93OrhCDV6UgfMwog+fNridATgrGi5M3uD
1dfOsLJea3hkoIxpWHaBMG1G5h9FmkJ90IhPxzWML2dgraCiXYsIuUMmAQyI8mdMtTh8N2GLwbb8
fjg3vTm0BBXbaYC4DRtStBm8jqxggNnJPlSaJnIRa9pfbUrKTN8BDs2LYiGzb+7rs8QSRda0GRcN
HAMRP1+4upKwfP+PVS2Sm0cWyS8dhME+ISVnHdEqn5ONdE4IJ1uoo9D4Vw0Z0Mll4HTf0NmgQnJs
65zbu6wYlkxY6a3end9teiBH61mcuZ5qs6Qf/TPObE1PZ/1/8vow4alj8Wa4cNGbn15yi1WGz3hb
zDkJNWMCwWkGCfd8idpPYtBg0oQGiIGjYIVCG0wlW04gL4Ru9XlBC0/EzBb0nF3Y7Tm+3x+byDfS
gAh7KHzlwtlE6ewZEQ38H+QY/WgepCjyCo+To6NSGftUqvG+W/R/+gWbiDY8hkUWpE38z8YarViE
IxOOyRxSXEpvUhjfoApzggvC5r3Nlb3abjqQaKo7J396XoLt68HDJc9QVxokyiaJuT6U3d4esVEh
4q4n6ryjLeL53eI3T/IDwxJkuIxn8R0GJOSpa7Wuh6jVgngiR5tY8SBYWAGUBezmsPfIBQQXzgKy
EGKlJXAUEB1OZJedqY3hCkmPg9KejMoFQ42o3KRQ/+wLV5OMymjS6MPgCNtQCHa0W48g7AT/MgJd
N5rbKvwjtZdM58Q2l0as/+mZGty1S57SylEF7Z2yQq5Hvjl3VBiLwAzWYw8pvAU3r762kZPlUEtg
oXfzWgdtHGZo0ZUSaCuKn9xF5xkThsQGuX357/KKh4ZqWpjbCiiLQQcFrK79Uml0+BaCj4K+pbOL
bzMaDoD87V9cc0Fr9bYKt1x5edLJIUEQlKaQUnto/XJI++ijVccEgZjsXA4ZdDJgSDlT2qGFk+eN
tqtOgBKpKhOrHKHKoPEV2VsuR+1+1ILfzgseDr8lCnqtbqswQxU+28J/6TkYFrIya/jV6sqGOI7n
3i+2mnFeJONI+x114qIuA0vJpWfixPusnoLg41/Qc3UQbe4CKLg/but/1KsPK3jKZdZyFpGUwW1/
YkZErdmQYZvKXxB4PCmzJ/anuXTgHLhGwSRDFQ4nfbC8rO4MfXquZWoxmzHhDx/fkKwTV5lefgAb
taZzLkE19/+UoKxnXafNzSXJ5+sM7pH/wwHXiL1FZ9REpnq2hP0hZG+hktjowwFUnFcByYk4ddNB
NwAlxuYyd6u+tOsF+oBp4HD3s9RQbdk0o3DjnqtjQVAzv1F1cdG5zuXIIZpSrNzOUb5472hEV1iS
RnF8aWI4K2S+hY0SYaped6DntEK8o+vB0ONZUkirZa4XmR0bL9wINKnfrZFBt8qzE96noYFC7Eag
Vk9uzhNdoXE1joI02KvZ2s7E1eWS5/y6aNCRX6u11P11C1MyHzdEVRQIa/yJbs3zAVFNMsIyre7Q
8BkOfQLUUoPS5z/Z2P9tvIIREmyj6m56KB4z55d3+lOMSnnBh8UAWcCrVet1STi/K9kBztu2G4aW
aXwALSF1GTygnrjlQiMMlx40l6Hbqk/g87/ZEJsHvckMvy9Z74DJpoAziHcGEHF1rCefxa4I3rEk
gBNcZxT4MRwEl4smqlPX0oHkwrTq4VoU9q1/qPLm+9qOQYXxkgDqWRKmkbdj7hPWPZkpVCHpU3vd
jcd6Ljc0yXmZfbXJS0ykNw6raq5FFRW3V09WCfNtVY0XY9b6dnWeyxvBqSzD4NqAh1E/MrbMROBZ
tLwhO/hFBI+tTSw1AFi64Wr5C0PrAUQZx94hCVDlsGtjhzADOeFPKSpPOnw8KOTJbt0D2RxK9EfR
a0x9VwiO5gbIxKYyKY5UuBWOEsG5qaGShxEq7HH8i1gAB5WwgZTV3BkSg2NbGW+bKuPZ/lz1e2t0
L8DH69D4DHm1+TGGnEgo0yldWu4JF7Hwai+b70lTlWc4UUZKy91pQIFVrSljcTXOOFW5j1RRySbp
gquYVf84LOqk9U9X+2ENRbRLM7eWjNiF3NVijrkMp0MW0aW6MIaJlJNDWFvLAcKgbiXCSy0nL12S
K/jxju/iy7Clu0RuAtHJne8OZAciJDnG0qhHz79LgyM00OiAK1QCQwR2/m0gFfAUeAzQQOX/Ncak
TIP/G3v74OAGvKNSAsqz+0AbETQEYFTimDjX7anaafOozE1FsMsMh7paCDqnjtCJuqZCVv5Trsg8
gG9yAP67oPLWvWcgq5owkLB461Cp5MbEwBRHOSV+Vzx1c0qjOpG2vShqXV9EPuCWs1N2pYIdkWFo
OCSdi1H2Difh/CNN5MPucXQ+5amHeHlxbUI0W8fwOnRcMN4HDyxWdrDUrSEf2jR6Qyz9jxIXU5+6
PkLGhZp8xAswpeZlKezWPvxjLwJoXWKD7aTLoFIr5dEeRPsZUFR9gl0i1UiEdY0WCFcsvdcZzDLx
PsYfca67GdzHk2TtS/cEnxzHk9LIP3/NxWSl7kqlj0Xf7Cm8fi2tN4L6wdoEnloj8b8u4xzhbah4
P1ZXWkXlK/YE9lah1VupehatOZLneP2l4sOXlWPgocrufgmpPuQ64fKMIN79j5ULK6mfn79iAvVH
8lWDb/y+fphIszEqj5D5gr2qA39li4/JFU7L7CUDzr1OuqqTNLnBjPjISP5ECD8FcJl2Ud4WyQdB
5ePmlTtOhzfdWMy0u2Jr86JlIc/bJK77wap0w+G5IrtcYtHg6rNhzrjjt5DgQDs1mE15luGOVAcL
vJ7DloZGex0yGplA9YpRLQiCDQ488O3SMhs2hFuv79Ul7/7iS2X7dbAtqaGnlO3UNi/IxLFSzjOX
TYLWOyT+AgUe9mkl7sYOu1iNW+xsw7BK6ApVo+aKhLLfkVNvwRzAqpovk5Td+F28uSuPPmnaa14C
Lnm7hB4fb1I/oJvDlj+VpLQOawbodatMTHekJVLBk6iHfS8bjmUD6Q+xjb6oeSnkH4/3QLmOtIk5
S1/dNmVdrhlHh1Qvkh/MaFd+mOnXS5XkJ3cjaOPeVCXWmJsfPhaJaTmpwh8RGq5bcLZwjjGlK3IH
OZngYdrNJC4so/gVuUOc53qw5lNyBGsGr76Vlvyly3s53kWdGtBBfra6cGpfzBNkDeYDH5r/pio2
oxNA2QusnxQEZ+AnhS22iogD1VJEj0kv/7yH144bC+oMhIx2gTzJTgtsCtXlpdnxh1rL34XJslv7
a2avbs3e4KvJkFGBMLii3a1fL8mlk12vI4dY+dnRhOSkAz5FEKGux8U7Zjk2OJmLt13km++S7gqM
4bcmmqQcDH8UfWKRA/y3bJMtigAzn7aOEBK5WYsw7QO05RGdbl8ufyyfQgYGR67NgrP9/nrdcw2Y
zaekC9jgaAG8bAKW5exJNAvhT4uXFFutvT7SlVXsYEjtcsxKqHyXANd6KgjdCzWDZ10ZPWd6cyzC
8axjS1ntJ9CyHDrYfLTGfukKNkSgJj0NWA0QK4t3l9QB+yhY//APf1YL83Teohqc1UeHE8z1Y+Vx
iZgCNMeyroWBsPDUlddLIKfN7pMmkVoVdOp1ptgdBoxmzV7LCbx++z2a++zNbYOZ+aJUVaKJgWLX
KBMMYbMElB8Xs/RRoCuUj/oOSSGUR4LyC+HVpoXSCwirRRDAbm5nnqjw/YKMLBoitMGerocr71Pp
OT5Q/lzSKKDwOK2C3rMcQ2gBg6PYn1/vCec2uVGR+34XaudMuj7TEE16uT6JEEqfmoyNhK7yksZ+
4jX2OlmK1flaHKORIp9LXuRceOKmYJ8GTxFz1rVedb6UbNxp5nOO6b/aHe/Xa6AUZB/fRqbRdfRm
SyM1l78BRIGRNN18SMbwAXpUF6HpZuu32+FdP7JUhpTzbTVqbo9E6DL/m0NWGWKy856vvszO/ndv
Yn4gJsRFS8zdf2ulg95fkZUFEK+CsAT+5O3iQZb5Pk9ok0LpLhCjPRJmGP4fXi+p8yVGkpUvt5CJ
mKjpErsWxHHpQoDiVEJAuQ+s+WwApUzB9gPm0ARW2w726L4AXYcVYEo5TFluFg9bkisxkdn1oUTA
c4C1vXEwu4ge9qmP54geBAsOlXyznMHXa7XeWWqiKRvQtbB0ePoKGSaXvVYTfZpRPaCk8T9GJI57
NLTUOALpAKvPqOSP7B4FJSoCUlIUJ/iSDc3u47OZyY1Pou05bwlFt3SgzginljGGWvA1gPJVDTa2
a4g+nRlNw85v6oArq6gC9vHg3KTcH2diMT/3IilWXgRed03sVj4+wi/eeQzoh8GXcThjhlbkWh6n
xnP9kfxYL8pVLXid9jc2+Oe3wouFO66rwJqKtIeGmGGDNlOd2QyeWOjPgIMum0kKPbxvOJWs+cv8
4M0m15RgVWUBuhGSSe+BEFbkPaQKFWHMhFyKhtSfmLJpSj275+D9VIx0xHYKBWOAe3QnveDTx8O1
JFcmkz57JIMZjDmbGkMuAdNeBxZEi6BIWRzqSeOyOgoDWgNbJrno9/ah4nWvcezZJhFuK8/SrGff
UUR10Fj9r94X8s0S4Q1nk+BEaTk7B+9fcmBIb4T2tIe9kpgviT5/k9yp1KVf5vcWUIVtGwiBeiSz
4PpVAUMZGpbwI/TLimbr89Fh3ASR6BS55UywbyYLBKvA1H0sp4o8TBcLqUeBOShelN3a6WWjyz6k
EFjEikYl4BqW2lvTQtC2zsE1ek4YbgEdNLnwQwqpDvsYAqoWPC9ugIyL+v0kORrMcYVwZ3b0gt0K
OOHs0RshNw8b1n+rsJZEVF9VVCyOeIx+Pen752bie6rzEcF9hEuvGDntEhTQlgYlUk3dngYir1iH
UHdT2459jl3KdFXd2Xt9ZhmLbT+RSeKHraNg5CC48Y6CDoO+hIEnfGuGiaFQ/bB+OcWefBadZsHv
pG+m974rH8vdtZWuHJjiAS3TH471fT9IFrrfhMmFw+i4sKTU06n4gRVAWOMmBDwk6tMlCBG4IXNA
7Nzfe4RdAFm56FrKkNol9pSx3iqV7zDrRnoJdN9jm9ekaMUNfHM77/dy9gE8Kjd/wvwZXv7SesPK
0wZ086dwa2VrPsVBXxLeitLVmzKoeru3F6kUC+9dB1Qda2lx/xwqClOlle3z4F8xzJ/OkEfxV0fc
C4tUu9NfUotquIa1vKy5tZis1GkSGIPerOigIKZhZyKqG7K1QvQMA+lY+MIkgVWp9BVFay9bH7We
u3eodB3K7radmeYoRZgbrs18SfFwiQWlfXcM20u427SjRrG4VdEZ2IIbHsnt32OXPUKpJZXVrhtp
DPtt0+RLffxuY8TPaUsFaEtDfBQ6YofG6gN0Jt5KXkP6UkHpmpf4MxGOqe4UNRUd6gcLYYin7AgN
skkNsW5mx2dMM+18LW3shnajxirPa40HGIP/dOFTXj+V1uwlKuGoKisyeSmqAGPxKyOPIa5/qMWF
P+0Q9DmgYcDiRv8B+ugXI/dkzPcSrzDVmZbpFX4SYg8KfRWQOV0JhM1FOT2f4oBxwUX46RGj3+FQ
WSRkXs4xYuFxqGUUkG6KBbX9RrRdUdICeUFmSM2I4sj++wzHgBtnPDpigYSHvkqnW4F6TU1iPll+
/mHe2E4uVCqmRguuLgX+3HaUhNcTbVV6GFpnil6oWl7r3ef8Key0stS+3pwMWBvCI2i168YjDP4p
QHIu/T8FSnoHc7m72jBwkp82msbONd6sFCxlKdoIEX7JSeintgeQQG5oHnOL+9uuunbzOTTLHcsb
PZivB1if5kPPkJZ98Tw9+YNVEL49hyJq7vcZPVpi+NkhNCDFwTuwj7c56sNrtfSaOr4Qn4EN+gr+
ayEfll+9x0UH4Z1YunWROmxtqlAh8G0ZpyHpsRJ7XqMIyXTvp4HBo2vqEvrivW2k5m62MPq5tPRx
0b9wJYkSeyPzIRfJPDQpn53nXONvnWwewnH15lsadBD+HUsi5RnF/CrksDAnSZN8/cVbW8JMch2U
n1ihLvP9/zp+FlnZFApYH/R4ZcZ8Zp5prbTxk8RNDGGC8qbppffsKG5mB7jnG85EqhT1KEl4+Mal
Klxmc/mqlZaElOM8ViOPxSFVuatVyhDqdcoRCOPSzwNRVI96XiVJVjFoCDnMablieXlnQ5JR16Vk
kSfKddw3QEHdAsPHOUBKOE7yaJfICS44QxFXJINXzPtMDvlgmUeBYa9RdQlVLTZhauDQ8M5ntyTI
TzWuccBEIji6Z0CQytOjDL6LjLP3LjIH57Oysf918qkZEa0U4K02lxJzky/0v9TGgHWqLh6JHqfA
E82UnRX7hh1i8jXp794PnsvW/BSXVDOpnzdGC5vM6cbK0PgGLlpNWomAGDPpI5y2i37eC/a3dd5h
TlfGXqz5ee6uvEhedNEjFLzNhKIMU5FHVJr9QC4+q7HtwOjaJ1DziA5zG0Csrgwip8M4WYjWTgX4
pvvhEaEcX68arHNCP4TO3zKxWQw1e7/2HeD14rdc3t3jyujdfBfnwo66+frSBXNpfwRZ5iCERT3q
0XZ91h3ldxkyc5Er8byArhEVCVLrRdOYtMPMPA8Zk4ufh+F6ng7MtKNaNKHg2lBEA3KBhsn3T8u1
zvA894g+pQC0+I1h2Y89K4Tb1Ep+z70/80G3VFeqnrVvqRErCzFxU47i7WbI1Y3aJ8MrgTGyq5qd
fK1KdMF08XT0fsCG0GSwl3uJmoN6sI14xVwO0QKMFR6lg+2xdnHGfHvHHfun12EK4uV0HoYeUJEF
W8m2iXZP0ElR0z+H5MyjjkeAP4Vp5FyGkrTvMJd+EIkDN00P/vuF2/IHiDgM3bqWJJTwVRNcEvP3
irU448jAnHVhja4DzEe97mwidlwb2bZY/lsD/or733uSdO0Cgv6f24cCr9PAM7jvKMuVBSSRXxy+
shWUXSHC3yGBIf/eZi9UxJOPsE79+E+tqkYxd6xdcefWgsGKckpa4nfvtBZx8qnkFSOaJKST4tnZ
wL2j7MayDvggGLlNYmdy1BAxbg4mR89eIZUATJTAmy80rfy7/zDxO8WAqo7zaNawo/+AGEKKPx+6
EUWfPja/MqMXC9grR0deuox2QPLP1bQk7ebPb/GjvUZI0B3FEUL89i+dR9M3dD7HeCDBV/PNqoQn
u7xMi+i9lUWDcVvP8G+7o3n+NqB76FJ+rbyktHI7z3P4UVwWFx63CFn34ZqCYmkU0KkbjSr+ykzO
/tID2EuFtTEuaftWt85Qc1QRr5GxwbIBTZMnF3P2JrWawJfURskM7Gh8TXeJtzBq9zT+xCWFPEr4
G3ZWWBh+UG5+dk0W4VHdQhinqyE7JIlbHVDQ6s439MopgPQGgYTw7x6vQF6gYRoYv12ejBaB/GsT
xWjZbf/tAHbBg4ax1clCabY93SgnPwVJMdqvQov9GQWAb5mQtOII5pHMh+BlQviBx/E4kGM/fgHN
Mm63GFD4MJ2FTEUQRYxkyJwPjT7ruoO8GxFOO9t74b73cgTpzvyJ3qWNNtvIR2SAQC0eZpm4Hers
Z3CRZ8p92VUIiLEXE5sUDaP2AdUcFo5oRwFDg8o1AUMGtM5Lm/K2xWcffHp0XKcm2XPClNLvHrwO
VnbyCGUpmK57JVkkSOBH8UNZ7aIX0x/OlGc7QRjS4TFQLFtVXTrJua1dTtKkXpGKG0pqSof3b3D9
/ux5WJEJQxBhnyCwpHz+IpPV1Ssj+dbwTp0q648e6HkHul30xxjqJ3A7vbu1hpZ17Jz6d4xXGrqd
VlQrquTHf8JQzYm8gj45IROAkClbld2aTPRP6AVfamdsRRTwj1aX0SN1ygTnSPG1J6MV6WntjDMC
3mFtPvq6dxuYd2NNSOVBGd3YyO7m89/XBZUoPWuMgCP901BRQ6ZBVSke2bYQ+dDvGBa8Q/7w+B60
e7/xF/z2cJdN+NuxQdkJN2G75o7eJBcgNt7KcHZn8m5rXsRM+skAzQDJcZXs4MoEyVwD/K0LzecK
fAVg5TmJnwM+b1H2kcyzPsqlC0QWUhjXtPAiqrhO4VINDlu2Jwy8bXjjiK+nn78tiWpkkr0Z8bbX
mGo/JRHxTCdpoV9dpC3jCuDVgKjJyrgNWre2I8sI5/9LTon3iTNvJUatKGC73K8qWzRLQmtX/YZ8
FmWOM82YNyV9lnJUV7oFMAfAzxn7zicLFZimw/qnuaHP0Gj5bFZdlDLyx7JJKIsclH1pm9OWi0eQ
S8i5JVTDN9MFDhuPNE3d21ky04y5A7SYzq9qOCSguDI2taSMlDvXNl/swE+PANXEGLdBAvWqU0oC
UV1yZypLgMPzAvl6TUw4NWqbayiEjfeHoPEJJ2i8CgOeBTo61pF/aFRq8Fppfys2hytBBgfO92L2
Pz2+x05752a6FHrry2vycTrAWxxqAFha2p48d+ACzYJt4QZ7SW+ESlTuX3dgJt3T1xBDlO2fI5zW
jSO/OXMpRYRV1yhOcY6DXH6iS6GwpiYuPnQ0McPqcaV2i2LQagA6wV64sBXG4iJS6JJoaO65xJW9
WDKT+YncJkdk4V/bXJQXIhAz86i3UyMpyND5Mp6j+iq77pBH5IziK8Cxz+ZU1oau6bgLA2WOkods
baJsWv/XCK17+2/BSP89qozLjBsJm09Lf5uVnsAJV18eyF+9f2T7s3AI4VxvKvi5MqruJ7Ypl2Tt
jOSAzOIKcWwQlCtHBF5kWZmYg/HWAoyzEB7qt7qccy2FjWmYLGhX2mXfpYZZgAf3GOYANaLd1Yta
D61FIUSr23vFWrt92YH+lwC+at5EuafaSdC+XRM6XbFFdvVQoa6p6KZBW6f2PkTPBX72wtpFl/6u
pA2ZU3YZ6dVSm95x25l26eadpCcuDIJbgKnYjZQj+RhAoCVV2d74cCyGB42FSLYTjppMxSY7RdYv
xI6NwJKp1r+PifCIdYagA86K3xq6d2a7Vc768dwSTd2Q7pKgY98Jy9FAgZIaj1phkIOqf/oazmjN
MMIg+jZpA8K7UAOgU1Z3QmaI8fnyjVzPtgnt+Ycuh8kR5wqehLXrQfDQ1EqwwBe2yTa2yzllI3cn
HBh5JqYj4hvXRfiBZNRy/xs0Ur7U4cuMfn/GMTjEL18R4w7mLBrPIRa4Hp7gZTJlmlFAyhklw8Yx
VzC3dKw+A5pGmHMDTMFeEFCcdoBx6xvnnU2n6vob9aqo7TDmYElAQxd5Eg97stE37eI7Ii7Zh8Iw
OGyvLpcgl08OZe/xX4lCEVk38tzVhXdG5D7IqkQUCB4zlXrphyd4oifXgKoxNbAPLoZAnS+iQqX1
RGrHaTMU6qef3OCx0i5a+0+Ir5hxS1xljQp+nDJTI6p0nzz2rHfYhGIhufkf+cQ/LLiGpmpgKV1K
+p9zdKQxsPvGAz/FsCwCKggEAKpxnu19Mij2esKlrID6ClPG4+ou2i3LEB2MJruDxyIaRtpnG5D6
FkyY/EwSU53bNWBVlj2UVZB/KT5WWe9y2AjRjDW88NkyOvJIk9hNuuuDxHPnQpXuQIObIO+WaaPa
9rEHFi1kkCi6eoBctjhjz+CYlf6bR4DhFkZIisThErtAlr4trRvcRkZayz4Fv5qbnlROIm6cEp5S
2fzZ+chMKxvjh4gehj1eUMInuKxmDts77Px0ocmNn3xTo69wLwogLwfQrYupgBq/NfVx1a47KAAi
b31dPImjz+5fqUUMW2X1BBz01Vo6j/SZ2lOMDYSxADQclL+fT0N0lkTAs8or6NturpebJKwV/rkf
I7g7ayK2DsDCfAQCeY7o2XU/BOJNJ4kmJt6ZbElTPUADp15qbcwvJjZfG7H6l3VRuxi9J3/h2JVb
/bBA1d0H+cofh0EyWZ5iQrNev4yV3TroYArWWA7RoOCms8gacbR9d5QwcXlyMybLOpOiHHf6Q/v1
IhtgJd0BeNS84tMRXqXgu4RAaxccsdX2QBeYTjMNJN7Q4/306TTwBdb2jPb1/AUVLiXOqgoEtjH3
+LnbMKQ+34TMKfTEZbLIUwFgRZ07azt/LAg+ktgPauwEhhXxXRu2liKVdByzJxjyYbnEAoTbcSe4
e2Gjo/5wAPc3kZ+mRYFE1B7CmpWUXZQYLhwciU9v/ICbdgJPBo5/qpCX7VPAVpXD01ag2wpazkhk
CUeAdQOxKCa40xQjoJ+6U1ZmhdY3sGXOjgdoj2qOEYwC4OWYls+NtTXsKReXNbtnjjotr0/lB8RF
khc1uRC+27I5yNgXTtmN06YPW+SjWh13AbrCY1KpP+iXr9b0Y5yp0+LHRY+teoM3lOw9/ftHhpGQ
fok6LABDtdvAyFkgl4XL7rwfKeKa4uSx3WdsmhQKxGh4Yzjuj7A6g7c+JKJPSRlNlvyUom1m3tJI
fhlT45+lZhVhroVljDw54MMaTAzp8oVriCtq0S3kZ9UZnVQ9UmN6fvLcHTI8II/EVvFtH5gZiGhf
1EjA5D+bnwbjD5ALwL5t3JP8t12AG/nXgEAvtK5ySC0Xi+wWmipxrLusM8UFvk5ABYRndXFGe9M2
A3NI1dRjTwBCdbOZFQ0FAUQy6GjrY4IpevEZf+K2F9kYExOU1K3ndJz1rHnCaGD5knKoYdNVQJbl
JzgX1Pv2Ro+FQM4WTpSJswWD0RjGVJqXn9zR8CUNpTdbekJ7fOZykdTXK+9srJuDjyiXdG1RX1oH
KSeD5irQKRAGXOIPVHIpfl841CrrU8CtH3NSEKOyd5QWmI2Q0nVXgxXXBXviz/kvlh24n5iwGipZ
9hK1O+pdDfG4CeAiLqoMsGBjwTdYDhgbuBGFbIyS9WVMKdE20ZJTcILhlDmjngi/godbomNBmAwi
GHklk6foymTWnhJmUy0H7X+KTIcMDrgySJC54WpLgL64lfj0Nnf42S3FvCq0lOhhQKBX0JJ0pdTa
Y9LgQFlBvsNDj0K2ZfMj98dlTqFfeF7KW32lFpTej3SRUrSiHKknwBnnxzxoOMeSOF3kLrhWCnJF
uteX8VYK2BvZJIvlxxy88F2cKpwxAwCY1JgvFQ6Q1pSE+hZuZxxrxzHEBV9Xfj1BZkN9OaaIFqB1
oTcDufk1tYlo99E+iuBN9/scYEkQMYsUyov51HrUoldXozv2+T+MOt/sy0ByHaOIxwgDflyDBOA8
QnSlEyScbiEwoAwh6/1AqRf5x3sErCiuwqbbmTkghjx+hGKzy13shoKKJiVDbt/UB25tx4jf+AWB
m16dyxqFZkqNHOUQvCeQY4+ArvIhhS5fWC416g8tKxz8pvgYiW14WMdFk694PJrnSdMmdaTvuTEz
wxz3RT5YEjRnHSdQgVg545YR9nnhNj2vdQGuRPhJhHxnQKLZb6ZVwrQ1oOHHSkZ2g5ZPBTRS2UnL
RQqyWC7Q4jto/jpokBYidexMb88zUy2Es7+ivWjj0LNxDjb48Q+GbZUo/39hlCWW53tDciGnEvVW
aiiZfUzdJo+NsWNJu/4oCzHDJ40LNN/bUJMn6StmcTACN1smbd2LLOpiBLaoy0g1cOoIlL7gqDYL
yfh33jyWHoknmEdHh+ObRRBzlmIvcucGeID4YLPdBzDxgECk5ejQAiE4oFNNgC83iO71jen8qlJb
V/1ErCZ1/4qt1ce18i3CiRfvdw3nAtCPop3t3RP/3EezcOt8NxFNiTjH/8MclP3x0+WiG3ZJnVcn
JoB+c8n4UnIKwxy6NcAutigtDf+n7+xHWCWVutQDNEXK3hvig8io9KLh+Yo0p8yyKxQP9cRLAyW6
2e9g0LF+g0ZbtDzAwq5weQMtZcP3fOrRyATmj0mY/77LzukaoFsF3LQ5CY0ApqacACih8IA71TGb
sCvY4vB7uBdKU3R9P7E67K00KX0KE+w5lRoB8n5jFEv/SyHiY9IRkVUA/Cj/wCxLg/6j2Z7ZJVTI
Afm2PkQAv3KEfuJfIW2eTAktkEFRO8xvmTjTLQ/BCecmk22KQ0JT09By+CxzrMN/VTvC4o97fzg7
vPjJRDGA0/dtLeOOCe5zdC42QUgAdJmldXY4l66g7Ufx7YpeqasSqrkOxHEunH1kQmZrg4sx8ZyQ
uIMZjdDDqp36TjIGJXcJ/aX+FhbVVftROOkHpKAPaUGMI/0jzZTPlSqci7C2D/eGrqtciddqS9dk
2Vihle3sORes4X7dlmUydaMDBjms7l4DB3IM+gFrCstX18kPHYWLu0byo9imVOcp0lXF0VdOCFxs
BTQg837WzDlJJ3NQ6bJb4KlDwvF3EUrtIV11rdKbmCa+pETnVKPqMyOkrMxGNU2YL7Tyr4Ka0Lap
4HdeevpIe1elzze7zuZdVzUxNl7ukJ7LALBw+7el5QdZ0SOnQzjQy4p4VruCGxMBhCQfG0osaX+T
rQkabk2QjqxonhHoVttvZbwqABH2L8fABp4Qiqm1J3q7qOajroDjWZ9aKkRgAor3vT0+QhLo2Kqv
Bz2nGu0/93YOUtc2hcfGnxXCOxOe1tBjfV4K9HWjIQqiOz0Yb/grazSKhtmYHDW4UWWvLHFvA3yA
N55eijMlVsYoeBIHjjKQtGHz68iQgC+QAOUecazDHMykb4yzPvRK0tvNAxb+o25zjF2F2xeb0x+J
rQlxIVzllE+o5Xjxv9DBNtux6M2zzjzRCfLKFgb3AFCFftsZaDSK2mxGt1+VsQoSr1hd4ffzH5MS
xFKIl5IvbEJfxKGE3jKRBIpB9hdHpt4T15h3j6eJ8jytUTY+LZd2WFPzoGgcr2UkpprrBt/gr/nf
8U1SGUCYhJ7ieGAZTzUG7zQ9sMFUT3sPGDeSCFZpBrnQmLfKX9w3zZv5JtMNWeD0u3fEexIjCBEN
06Rha9ZA8zI0THF+nqU5lCuLtb+fvBV4panOvPfPrmFSYxQnLjWiIelT0JjAjVxi//ol+ay4xl1q
sVDbsu0LMYyXbX9Nim/mBTYr3TmY8YoUsVOT1lqUYAMLN8qsa97fPs9KDyKBsfhVKPQ9ItiDzpEn
y4Ppwgl8MfNCNxYp+qjEn2+peifPNAUSd+QmHMhEQfSu/cgfJBEfl3nQkePcA26hvcPF73XsB0+N
45gMVzwPKzEM6QdJGsBs8WTs5DD3/WjrclDkbHD8TjePyqUTeM1lWMrBKCiiJF7xS9ZIYCwwjjgH
F9P4RTNmqxSvzdKOCO6qnOjE4+7IZq1yoGC90pVVjX+X7h435HTBHVxpUdgGuQec58GNLLmczEQ5
/1ZgB+G2CUPaxyU4U9ZcZzDoqfCEOKqv8j/9pzrp72yPhCa6hkCzLC+YeybjOH7Y9QTvo/Y49Sq4
kBQM6/BFfm46D9zVee3DFrBfTVj52F9UTZz46ibxAcMN61enc3ALdshR1cuBkTWzrDxX0jwJjZDX
zueJdvBnJSuKeAL0YcYD+MyMZSnZ+1e2Dk9O+Z52+PEtrnVh8uKITRTolWhHU0T7yi5XQTh5g2V0
msGz0QZvyTSUdPkuVV9RGvwq1Cip2oS2enu2tZprnE1Z3XiRG3TSeUh7pxffs+Qz7G+PZiEFfMa2
AkkSooFaCZorI2AmcvKnYzR/weyZ/c8kHp8TBlJ/G6opsbqnCQZkr6T83MLpFH/la3IhdgtIWjz4
QYhr8DigG9rUwKxevu8BXWDrpccnMePPE5OcrGw7n1eSo/FfhPhFpZBil9C5hGdP+6M1UfhCOSP7
nor3+EUWLn4nYDYeMWDj3/eYzcm7+N48dJb8UupmtDltCItUouhHd3wXfYSn+u31GXw1AlC3v6qT
M5koR2Xm/GtEaz8Y7ZOydxJ/ohG+ETx/DcsKo4R1pUCKwcOReNfKTtlqvH53Krfnicr3wAjwHuvP
bK29VXmWpwN+VKQpA7TLIvqdoLtOzJ7pKIM27CbSLu8yAxo0m2bkJJEQIJYsW05S8YXzm3QZN+fW
N35BUea3TmBFhAj0Lmlj8OdUgCySgf7IOe6xrlSorYK8BLhhDXRjX7IYeSQvujrOyN7zLeAw/0nZ
3U2BS7Y68syGmYe4ZszqL8RgR6BwzB698ekiYWR7QQr+jHS706Du5htNcwERu6PikPCd+w3LqDpf
XPBK7DfpH/1rzKpS+s7aQTjibvi/UGqBLpXnpHcDNOYTbWYAw34m0nvWSboJn4liTREQMGsiUS7G
m6Zy0rWy17NJENRSx86omAJmHlQCDglZ+9udMN1D/SDicDnExOWuO/xCibULz8TCKNl4Oetmev3u
EkDtgz0/XcnmShhl7491pBmq9WGkNZi+ulxQYQiwgjTeDMUXrHTzCk1ATGUZ121RVqRtyrieMxXv
Q6YUs1hJ7Ceg0SLKIgvjjOt+zrzyTYquGD27R2OVtF+9T7w1B2bh9UauT6/4qkO4wQ7iqdeHLH2s
XIVHQVMPGdll/HfcZVIUdEPwAHEOnbvTaamMeiCxa1EhLLgbOrafpBMdww8bFEgA6AaKq8gGsTj1
q8LsacnuCf4GXLQ+N7+NPpY3miM+ef4NAze/xrHLskFfMNnmXAE7FrPtTaXtv261aIyfsI3Eg7EU
hT7dICjtny/b5lfkNrtlVrxX8gM67iV92xMHGWiAGHdve++h0z3Z7Jzmy/L1+TGbHL/oq5DccQVR
SkFwAcsYA1OzJFoSjYNx7L+eazne82l7u8Hzd6jpT2m1yD7RyHyMb34LjqjHQvE8brgt20xAtmmR
p1doDe86D3Og+l45Z33a0Ad+KFPpTlt5mva/sEp06e3ClJsJUtrsz2A9r+LUaknrgJ9tfu/PD9z2
2GkRn8MIvcWu1Y4W/4cKEAPNURSp5Vl7AYT5sPfxkxZBherx4zoRoXW6XVMhYVWAMaYPp+7pObSw
kf2zXt8DByiTN0Via+YmMzuXXNz5DKmWqYYwEOQw0U/8P59bi/tkLPo4Nbs3CeoaArYaXLxRBsd3
NSQ8391kusDT+BEzDeEnnvYzZWMf4QV1l1XqcFKuqWFuZc05AKBDWTcWy/vyKY3jEmtYWNLBgUGx
TDjQ40ETCHmEvMNUu9qwvGUH5nSld+/dlRnaaemFj2oL1Sj274J1AYtCzaj30Qbs+AnaKQ0AaSNi
jvTWq5GZ+Ynb/29PFeEZGMO8C/d5G2zL6NA+UBB0dTYgYmNzsTqqmISFo8WV6xb6f4n6eYxTgWjD
Y1T4zWBiZ/2w/Ao34gkjaWU/xiRkoGdpHXxZqX5/JS4aYN4MufvJnywV9IGhrFIKdJlz5cdzF9F+
b4wiHbFFM8LsjvR+9ohlX5EoJKZYyvVo3g86UHE2ggshf3YUTzwK2GmwK+b/oCt+4IyROI7uJoLg
pvLxr4iBn/nV7x8GpnbI03R8XwPYbIH1mPICgqHpCLVHRrhteRl7CbEbaTjKl5vUmbB1+x2vd/TS
l7uMjXsJaKxakUl5b+3AYSjKJI3TYX9USVaUPlgaa2Jr+GKHzTDviTJU81jkWbVN/Gq8CFJTkkrX
XAZI1HAb0iaee6762WjnqAYwDMit8Eeym1/kMQjvhCIojX40CvLB1DHLzUCReYDRo3fVgzyEPVZ2
1/mK1pjR9ErICtgPJuzjwFI4Vzj022RmzbZpPKJSdTdtymVhMLNbXh1rc4rgKK3pavRbTFFlZ3Au
QfSTRb1Fr65Of6+ZA8ux3FJAie15k4gUE84trbmSN6NKvYXz/waZT1M/vAjN0oW7tawbfhayWHmW
6BXN4JIY4J2zVyU1ZyjexZjjiXjzapG78urTtrJM95Halhs4XUMXWhBYgPLCyYqfLepr/d+ysqOQ
JHRuVqP+LQsvrvrqoMGtjmFoZ+PHtqOZaKWgJtLwMAZMEvTguAAKoa9H9o60RVGiWh6emvOkxNve
5SvM4iXJlr83Mkflfe4bHDbsiJuDSHtV+IhbaM3S454wRVHb/j3BgFepB0LQxwxx3oQZkG89cb9S
Za7L8nTzvX8Dt3lnVqzyzpPE8+5WsGzBSE0PByIo+eQV06p+eGjARlFTo0aYtx1Ckly1k2Pd8ajX
jmi6jjJdo4xlrhsw7eVOBtAsIrjO4WL71VfY1cA/Jw5vxfjPmWbkrBLapHGT6Fbi2ANanvEivNki
VZlul0Pei9HkXVkKiIVvk7pXLB/tjJbEJKkHNJMtZTJNhSa1tX35m7njvAM+uT/92F9jhmBGAPDE
Eyd/fhEwe5QeWvQwyDnvwRHndRi5qcA5MsmuQNjbieeGPJSamORO/tjIH+pM60XRNg/XkSFpqHZ4
ydW3n53HPII70KHkmWvGBDo3eG35MCiNVhZhuqUWxhJWAHnlMGjW6b/O9bEKi2fRkxkPpTdogWjb
GDdoqBryrDwUroJwnVtHIwugeT4tch934D//yWqWJjvlvHNN3hiEKxoTiYKp/6v//MFEZ0y1lIcT
HUISh8qJbout7s0y7E4jAZvLlScDExtuFCaTFDymz1Ief4J2U37n58yzhrDX6jDjW8jBu+tttCsB
kvL4BDUUYed7haoWElbx/boi5NynxOWkNXkqnl3ERtYlm4iJL565ESXx5AGdAD++ZaaK92n64Gwz
hj+O+4JLwsqUr42XntrZ+spL04GS7GegJsUVe2hGxkEa7Sxr82PSc00isanIahrX10NoCzpKPorc
0jKRdWv9RD6sRCFzecRNCvQMvgM359ofg6mj2NMc4//ODLsiQ+ehYbsaaIo78wtreXdJh9Ktq7ly
M5edmo9qF6ClD+GsWg4pvMmfysqP80FxFIvN4oSsnWuCC9rEqfMHqEYDBZ+RoRZ2yMHPqwyQeMk7
R33FNRrKkeyOHT60F/20Dq4lxgrXJgPa+H+C6hBMqVAZ6D6RFop8KbL5OT4pPC7qNgTj01TtYkUO
kT2uGvoaLJAac4m3zhMWHyOdFAtf/CHuz/PUPjF0ZA5wnf8AEgKqRyVdtSvTtlFBvZBLKsXbV0r0
AWoDKBZrtfIcHSj41PS6cAWGRshWx9H2ieTR7MgBEqWaD/zrRCkq/Vs8nAQFPKyMgDLm9+9MBGmk
yEhTmM0oXJl6YIwOyOg+o5cnuROJ3zqpowNlQ3RCDZo/iL5h0t4o/zKpvYgFNJjaGEY9pyOawUY3
Dv2inbsuByjNOTaro/xAoXwxphKZ3psFNNHBhpl6lHXxQH6rUTSN50YZ8OcExZlCh0kuS2Eh8CfB
5qs1/8JLHHa6oZkHOxtQrNrVABzy1PuQL86KPD0Ocn1ic2Uf8dn7u8/5aozDpCcL5pP0iPDYp9ro
dvn1pvKeLjUlMXJB9s5raDES2o8g4YRjfeFwETU8N5BqqK/A9vABJSOWvlyRXLFGMemi6+YfM2i2
2rEI1yUfcbbnu4TVt50JMEjQMrXRJKYwOC5JJuEqenBvo5ExYFRoqioLriZUB6LY2SCehIIuX4PH
xJwTsA9RXvT8WJfPeXZZBsUHZUyS9VWduLzizgZD9+nWuhi9GRpnu3C5JBX+xImdHMVXo3/rN4ic
qpEMSap6U1yHY2SxC4Jd/6CKVzzaO4e+3PxluL2Mr551qaAy9w5Z6P4UBNoaDm3gfyButX6zAY1I
OtB2g5+6Jvk9iWoIMFeh11Ww81HqQkrbcufum9whJMQWu7SVbUE4Fu2yRdH5+2jtVtznKo8vXNIZ
iTRCroovmGCX+UdVTEsZ4KmydytOqZyD/CfpB+o5EECfk2txchOJOXRlvbFxlCOKF3perYsOeI7o
POY+Z/X968Bg6X2vyxW0qxcgM6ntj+RtFzFvIIHDNJOWJ0g8ik/0yXpY6AQc8SL71v7OWe/QLrFk
xbPz1FwRBRp119jQttT+H8kucHnbc5k3n63Xr+cax+RTDzw3sZsdMX6RrFG7oHBDVa3LH91Dhk69
3B1C0+NZGY8KPlb/aPpXTYCWY8V7oaTNG77U9cMUUeyNr0i1GC8giEJq8zlIHUVfQa9A+iLSY2B4
mjw8QxaJFchGhmbLZmK51dJs2kBE60baLouKl8+rhqLd1aJctWCqzQN22i+HG2YcGvkY8Lhwgh0I
ZAipWfqHbq0J/lgWOklfhTsKcdM8nvhgtHOANTzAVMS59RVl6focJbliOp8WbOncA90Nn5FTgjIk
kpjgf56hB8d8UXs4lUPu0jsKhUoWSRq+pEbSmMDB5ctJhPRm4zkc0xJ7DOqcSrmXItuoU6JtTmUR
j88YdZTjRHYygOyYSji1x4NVvjrTWZVAcNcUNUHtiJ9nKBvFrcCKY4aZ3kyb4fb53+qbCQRAfzT5
v/NfjM30f5A2p0fu/vZcrYHh1D3jWkw2UlOf0hl3GfZRgbPgBp2oOBDP3qPokRcKeUXldHjYOlyZ
4dNGp1McC+0NZG6xJD3JyTHpsdXi3hUfJ4AzP7azRO8Lx0aea2zXTJHP8D0TtxOwf2faV/HahJok
riYPvieJHkow9UA0ra0fHi1/2/y+la1pAKhYS37zt7Ff9jKeKSOkQCMBlS+mtStgA8KhAj8LRy7i
sGwtQqMbnl+IUYTvjxgRw7lIpU8yYm7cOk1GeHDYdQxLs1yneN1ct4zGxVmzGkWpMNYWo4qFIolP
Nb6jhHMtLhqnP4exQY0EQ0AnwfcPlEnIyz9ikLvOWq3C9h2TbA7y/PJcq8e3yCzJ4I3v8rO1tCT9
xG7d/0swGWm+FM9zMD86qsITx4gm0iQesqX/gGQfDbAPlhyPC1xAZiuC/7//TfM9x0OkAOS2qVeF
VC1qYDqx51FcmizzNGv3qFArScKgVu52c7ECh4q/g8gcLBFxhZ48RHjcfb7r+aojOGvohm81SFTy
X4wys0q6MW9BHGQ2AsZEq11na9Go1zPrnEZSHCHAKEO8iOUPbBsRrW2NIIXtgOIBb2jBzdTkZjQl
gwwIs2/f9YpE0Bg28QKdwI0VBxmjTGg1ZO6i9ErWHewr43Qk0UdILuGoyeqyasY0hqP+fWEL2hKj
CS4Y1BbNKQpe+V6DH6RGrJBV/M4diZap7UQkwK+UiCJdZpBSOeOSY9WgFAy8byO1LiwyhWbjM91e
mdJDn8yql964SitBNFG7F/+R/UfSAqJ/gA0o8ze9DwkLEyQWMVMXC2Shdn6ZocYMH8mLpt/glGqp
GoM6faNiuaemdtG8c89e38L5f9AvpGbfXzlVFsCWfS7uHf6xQfKA/E+3vx9QVqOn4F0P6mWO1pji
uaTwH+rgF3Pvrez7mSAI4Ic/JImJf7SaA2+8Lrf4zLrgb1A9MB9+dBGPWTEtnb2XQ7yYXERoJo9d
4AHAUiXD4/ti2Ezbp2SsbV15kPlcPb6B+2Ur5aR+AdM9Vs7OvoH1/pAVC+HNAW6qFkWvtsIwWWQN
30Kzumu6YyJvhNQ3+XKxvs9H3gW+pnNUmw66uNroiCVCuZ8KpgXhy3rfQI5pLENsZ09XtCoHchCO
sSiXkw+0BPJJd7KC16hVFG/eR3nDZjkmOzPzaUuqEHwzUYFQm595BgfT5iNDmkRaZBtKGcRm43VT
WtxO+ICUCEbJLWnGW/wLUzzKV8+m9sOPXRZLT4JasBgwiTLl68savVz5XIVgbiIdwLIauUiqpU9s
MQApSlkZQ4jdYWhvYadwayy0yTfnTxvwZi5yKxYthccgiJbVU56QFHPLK36PWVWJCRSydbohT1cO
9JUzaygvFWy3d/zU60Yo6nuTH4GGq4cJYi5RIJmxSh6Fl7J5/wVa4gHiwRTsH77D1Qz3tL9jDP/Z
tFTIwRAHI7Gg+k9q8BMhGTZRLVykNsLe2s1p25nVX4UJkZWNfom7yMW+ICMrkQAjnQ0z0NjU2EyV
oDlTtL+9JEJYu7aKVxfP52bej9wYPybEyNEwHlBw29D50KTPSKaPJYJFjX4VOp54BH5TmgX3XVgh
4mJ2d9Xzi4gW/0Wn2fm3gXMG0qjt/DdutT99MUH4/0KhU0nKGtn6va/q49D4XlWj2sixuzmj6aeN
0GMwuDz6yVL0Ud8WWQecojufPNrVItbcIRE1FnZoQ+UuWGMXF8FTdMgZ4H8BYijsHugs9zMgClW+
27d/O3rEJdonTxJ+XLdHz2s3HhWe5v+S2YGZTuiy/mK4uKjcqZM1janbYwXPlfZDNPlKxAaJIBeH
EMPYjc6HOT+vKqFa0UkO1v9oYW2JUhUOESoQ5Km8oeuQNtTkYR+Ifvn4GcdkoTS8K/QSTqY9PsfZ
9pped8KrnLF6arOrR96FYOkEkQiDuQ0eBvay1JZi900QN1hYpHUNue7yZxLrwOsdleBdlO/sZeH4
qDpYTHOPjTD8oHImaHpYKy6C2ZWSCqrje9XYgHqynymbPOyBWNAcPXhoW3j5LNzEurDtf32sOCOr
BD7NOKcA3uG8ukzGs94cCcsr9kc+SmgVKK+wSQctdBOQRQnM7vuypAu7EGaj2WM+A1FU1b/1oFMo
+CFoJHb7L3sveu6/GVeu9l/Z7PdtXuyYrLxIHDvHHabcxDJRt7NiSH86TkY7IJG9IwKU99hUpeRG
Gb4FLiPAf822fDCoEjKI5276Ztgfl8nrS7FTA9um0VVDIhK5z/5Tv3qy9vncRnPWNF8D9XjP+ICe
WZrrb/GrM2EVnHo5r1ZkUmP7C/HPri7t6+vy6d0wRbj+Ycou2Bhhk0cRWEb2xiZHn+k7isbeuNaK
kEWgYuaBlEbF1WZxoXHM6ZdvklQ89YB4HC0qDQzU8q8ksG4tvpbTY7t2p5YyAIO7BkN6JAeaIoKv
ha4B3z0Ug2xzyTx2cWdiYwxyKb7S5LmowigRLajba9flRMFIGUqjo+5lU4r99HdK8WjY1t0QO68q
Amw7sXhgX0laoZX4tz71WT2yuENfCjPzhOE+W9RT5LDxS0pVNrEL4yeqAewPUSA9y/ejdF/X0tjn
abswZb/RleHb5+wvVqTxM8SB/FtjGuGn6hamHqvWUxVimr0urCwj2yQhcedbYGfW45TTr5DO2SxH
SSIWLyOV2cd+PWcZKWadMWQRyGwCSS2fmP3MrkCoOoZHMt42XI0wytD9xrdSoSXg7RckkR6LQW0Z
+P8GO0AsQPRjnKex/92P/HlICNloQrTvoS+NAAHfj2b4xRMoIeXbK3lIMpkZcfp8B0Z08nY34bvl
HWTnS1i1Y8nmenpzEjpzwvmKkzzbYrFQvcgCuMDx8Iq3+vwcLo3H5FdCIT/VP2N+SQCHkgXwn4oi
8beF/wcLEEfpkZ8VUjtLfE9TR7PCW3y8fhsExC2vqLLnnQV09y/9BR7Rz1TSTxU3CJeq9vBqVkdl
mQ4fFqgC49nxhMjUp+N908J+Y/VNzWGe5wrG4i8k9VJSsflggngIvKTexTOyMmaxURmSXMDTDCy7
Y/Ji/U9rqjmwadeYj/aNGY7XOVNcusBNialNuprDDg4M1VCnn2CLQPCsBQSxo0+5VpfmO05nM6Qx
nK8b4iHYjiW6kIWHIlrnK10yimmL9ViN8Nf9RaJUEtKU+yHNYXqDxOu7BaFrKUpecOBBkG7Xq/o5
6MI05CGw5TsM9N3jEZFiB9+HdCWnuDS2XMlXGlovwEcr4C9nnWjJq2ARSfdYnAaNX7p0tKuSE/ES
4WeUZq05DVVgrIwpLSsMTOHCbIe/AQLesKJgP2R+NEPOoHcgnKEOwPnxfyIgdRlBCRJ2aXmL9Wbm
HUE3KnyrkwMZjeCQNQzeXQI6HSjjwxGJR38C+pM1a0Syj+17aEB++7N0Kmem60oU5VN/lUv+YpFM
noVPt+3Xsx9BIM7VrLtDKxXyj4lMBKF5zAoO85GRv0mneQeLuCHYVh5PPq74VZExFvxqA46i3zeh
TJRZUZcGsXGa8y/I2FR9+InXDFPp8O7torTUhXcHbW577/Xecx7LGaza1puOp795ngMgIOPZRIWC
mdAwVjaRuHwrnt4xJqJ0d+ukOnJLs42ZYdjU9I1qq1vL0rN6s7ehGBSEEt4hgYKvKDOuUDkGoL7d
nWdMqKaBbehQELtCw4wCbBJFK3IdlylkXmKofKlJ1rnLl21dgUtmtXdsARfqw3ZLXwPjkeDhwIrh
Hxu+tRnpBtr/f9jj9O8ISPkr5vNa4a58qeLh7dq66D3nn/M12Sv3mM9pestPfLfIPP+Vw9CuTMw9
Jz+M2Vf2Sw6s2+hkEiMgIEDwHYVXVEGg18XbfT7sSc1LvZ1RObA/kUOpcSYgqP5PWpZxuFxDDvPH
Y2RpSnTOrVbdXj9G82rgsCMQNWW+0YCT4w7htmtoilImgJKcNx8O/MfISGSZ1ScK2ufkIeMoy+qA
iByKUiIxGtrh3FWQe0jLammWlnpMZRA4dHuc7aOLpDpFxxp9pZqRCnXFpU+zZLaTLwAtcFyA8AJB
OTzf4xMlWQkTaujKgw/PQE5H86DDwF6kfhoAv7Uwlab1SXaP/obBk4zdhVhRPdie0feTwEirGeE0
Miwu8MQgf8/mjUNnhAphlso2Cc8pw+NHd2AknOOvSLgEV1K2StzJPXz3IWWJB1znLWBSxxGz+dsH
9tsBX3AzYHWXWYhPKQlmmQGr4VMMNROB1YZ0GYEFYRNzjR3Pv8/piyVKmYmTHC4yL3qWf0paMMbj
U/ixW25UfzyLe2lFXl7OxIazu/LEBrF5GGGXFkBl4ig3wKWriyWTxpL1Uo9ZAb0mXWAycmcmVKaf
6yz6w5J73d4cAyb4xCWJm8hC5+gnLbtCXqteArCIwjaeYq7HBQEOIcrRC7cj3K3IcVr74GtCzNQq
XiIxpNEshGyRFx4DdhJ35LD0oYa0iFaqIvBkQemQmQqSrFGIz8GxzaoyC5dw6imk7j7sXL50LuUR
3d/cmVhfbll/m9CSnLbPOXqnX2t0UuOrmN3E3I5pcRa4MwXLlZXw3kNQoLXaj/deEaWubsb/SJcX
UD4rByOR5k501gQE/Ahpex6ZnZ30LjL0VkF3bqOyZ0tbVw12VxVEfoHfa8CeIvVjFmGtF5eSmZ/Y
LtDy/sPzc9NdsL7YGHLWqYIX0p2EiNCvCt/2hNquwYp/HNZ6RdlHWWIFhuEt+04eiyeUts/NHm2b
BLu/uEhEo1jiGfRhxQgYxj0Gi1DaSREA+HDHGfPiYddNJTf0aMPbMQ28i854qCSDyTl2ylJfV9mZ
oZ7fq0wyAh9e6z1vGQRUhq8DmzFP3naAwvEvabOI6sEWiq0/vv9l+xhW6avatZyEfuT+Ttl4rUGt
NsBVxiDMLMD8XJAcHDLuIFO/PxT3G3ZQZe4xWMDSxAL4bCEIXfZpdql24efx3gpo6llrsRuk+0ye
Iv2BOT9boOEYBbDdAO6m0hNdccQ6Of91S2m2pBxLg9FvZx+lIZVdlUrE9isOo6EaplLJJz18jhoF
uhBEo8L5+66NbFedIfRrCGwe/z4Y8cCkrsOryNBRd0a4/cWjOnJmMEr/0h0iYAeU5HrOlYnOcJ/5
XJZWuNn7ruNGRFzC5Q9lB1WPkNqRRmqYXb5jMQS1DZEJ5N+CQemayD+DjGuLlI8TzYcJukadUHJL
FxTB6Zi1MEL7+D+n8ccX9OjOxMew1PqByu5jbclrZJHrf5y4zP1pXz3IAPypyynOInNVFzieK2ts
gAfb7qRg1fleHEA87RwgRcnB9rOJqC1+DBbJCMkBzgl14B4SqvDMGHptZnI6jq+Jz9beduqm7Pys
i7Htrg2Hkl9R4t88xxR79zs41RLn8Boh91nhUw5OcP4bf/JcylPEqIlQCzk6QgUio4Zvbl2cc7r9
NYPzN+u4KaMChMfa0L/Flc8Hl/GsjoSiXeN+nNIwHM0fq8yDjPlCUOoEGJIyEDymWpj0/J3NUAK3
BmjIMQAkoo98kWjFJk4TL5QaCs0vipBfthHlTdChbPCXE9y0V90oSUlewEt2l6wCBY5zbIOXbeNy
OyDfWwiqdS9OjymOUC6raiqBogWT3HNNMAiNcHc2kHUcl2rfdl/hbEdC82kaXvDbvJM1oHgO6cZe
Oo3mzIZSyf2XdS4MJ6t9Grh4w+lICyM7275WQiG1b/hVWHNQ3wlQyV0L076ceUdTpQC2zFzYDsR+
hQjWtwuqVywhbpS8gglQ5Y3lJEHxN3Gz9mpAbbLWgUIVs4pUBRu2kCfUbNpfLNlxJSa8x1cC3tQa
GcYxlNY5YAIIklsDiPR8S+LIBhHbkrLpliFZ7VfvtCxQRkOdn18gMeDiNKP2kdkM1zgrKOENBqn4
D+dH/NCZth1pASc+wcVMyQgaRvaWrS7axHtIL2cMvCEFuyO1Nwv1EhiEWowVCGIK5VKXKNU7m6WV
QeVv4Fol9eGGEGiewYQ0gOr2PS6dwEIRb8o0C+a1GP08gpLdSFERTHkFAiQMjpee5kU84eQO4ZSQ
2XjLVt6aDIC6o745V2toXtAnmCWn2pJv0egyGjHj5yI5RxdRddLPvt+aGIf9EmEPE43tfHGnb2JD
5hTrn4Q6icxrP1+U8hJuLFcIyA5pmNeBuyJmbrdUxI2tTbENzBrPfVkm72PWc7Cus0aXiQII67YS
1V3wZUb58KFcLfZjjD1CfbfeB9TcPm5Afr9Q0FNy2SM/+SPjuTjtnK0KxsKKyy2srV305HcTUuu8
uhjsYNK/jshKfmAAABJdO5YrD7nrfge26hERtOGxca6R10buIA5gJRy4t4OZZuZKEU5cDO5axNgL
ivgMj/Rm2m3+aYOVzg0ZvQj2uhicwAfuMk1Vtvomc57jz2QV8q9PPSFSibcgmCPcXRGramNBhRKe
SF+1KsSK+HJhnSZ5sBEH5Jshau5bbKRp4+oieFyl3Bmp+EZqkTgkWzAtPoPzbk/y9uyuZaNy7qX7
Be80aTaGO1cK4PjkkOiLcmebqdNYm+yqatVCbcM6pnwi0oslLDfcHsUW7jUN7MCLjQPmovSOekpH
UuOzXAS5Amk6I3CwBRFJdJt0haBDeaqLGGSusJEmPUHp2bOx9B4N2GuNyM8xFfKugmE3x6yS+GCU
yCyBQY30J4RzJQDIwLG/AT63Ox0XIS+cOEnTgXluxRtUaoTx1CSgDoQ4Msxyq1m1GlrJpT8UyqCR
xo81iq4Z7/JQGDSlj4QV0pxOuAHG4pYatCPliRQGMZEqidieN+ia/DQeWvaXhk6nizld25s1kIIJ
ppVGldOnTfvroVycmW0zgB20pauLpjN5EiPhL3v4CqhBBLK8wrH0zvGEqa2rPu5tQQ2YImwS6hdC
3WgrCcr/202ffFGtHFYyyCY1s48alT1FHxInD4C5kYX+9MgR4orUWPEPPQ9zS9vujkSmcj5bjHdr
TDwqKUVse1JZHygKOAiXxe+nenqK3ayicsSiQRIF4mniNugb6/ClZtyow8H8NMxwdsV3qTW0dqK+
7Vvfp7slsDXEpDVHhBdx7Q+55BzOS5fdIH4+Vg5IpEvg69fpZ4l4DYA3/VoQfVc9FSa9AKnwdBEY
cEvWASvlKJFHQ7EBE9fTnc2IQzR53sdYqlplJDGnHI93BkWi4V/mEnE/OLqLKZSb/sp58pkmVx67
7B/xJSrkPPACfL8WwM18d7LLA8jpFO/uCr2/g146rDqhaMjBKxUahKTtntIaOzTnneGHri9A2H6W
cZ7gHfxHildLaSHymG+yRuMDXF75zKQya71E7/fKhykZMoprjsSpNs8ZzkqtvfGbEwDtxAMEaq9W
bSOnxecx7FAnAwS87+5O3VXT5yDTgVqMa353k1QQhxFPxPH3kSyS9cuI0CcjA2P7JTQi2CqjIUM9
O/W/x8jkGWHzy6l0cSbrNNt0Rve/T/BYHnDGjYLwxZ5uBzbLZnvgJz3x1zAmWHssBLYrQyTXnnal
2N0NO/nApofk55cGyCN8QNyrF9hMazbN9KWxP63RwMIZUogad5bhv7EDCI27ISfIUguwkeThuUIZ
XYmqymZtsVoGCHwSXb2G4EPvLzzWw+vENXLYFmxrCgqj+lPV50eSurnMdiHpTQuQnxvydSK7g6Er
+xfR45WnBLfhs2ZarbnoMfvKVdCfmYmhOJibDdo29ss/y+hs47NrSPXX83k4eYdPhMOoGG74Y1EO
TEXg6/AsELhqBk/oRYntq6BFCk6Jmfi70iWVXV69bJy9cbrQRNGb3QExUF9YhibDjCPcYlgrCTKv
2Vcvjlvcn/q+PRqb6IwH0h4MMMn4uMSfJm9uezsgtzLtTA4RvvI1jmryKASEheXHua1na+r4SqoT
3Djc46RtwTHi7T7GdByEzzPvqSn0chO9gu/nYpUnfEO8WxdkRyUTpvf9UT6xWt14sbJ7mwuow4IJ
/u6GYrhlx/jew4gp+1A+DRmAC8D9MIDkALgMpMBmnztfP+q3UkVX5h7tvDIG024emMO38QzTmyXe
rZY8m727AG6wMPYre7c6fyIcQ5iG8lkfeto+UYa5L9O74z4kuaCpH5fgUmbr43bEa/WouwP9QRCx
KERRwsFlhM+t26Lu7HJx4rzQJfaQFbsWijcQ99WvnVzpP7q1zFVrRJhUkRVTqeOFL26K9rsGpLum
RGW1+vKnifOlI32QLWxQD/P+y6LGRNf2mveY/Kb2MfEvToiUm/cvEvU7IdmGmWa2Q/sPuTUdzAyZ
EZlaxruxU4vZal4LE7Qig9UbQTmblH2cquVDxKo8JHdQItk8uI3t0MREA/WB4sAOaknnx4/VlN4Z
LKazpjEdP7761jya88yqgvbhDjwhs7map3gKHF7gOg/MetGouE2nqXxrzYRZY4Y7MJxiudEHql64
5RyC5HPmxuPL16a6nS+7Y4C3gNuexdEwbRnLO7Ixx4EdtJ/Fgcb4EOp/8cGA68Xp8xv5NdGhbP4M
N+P4UTXRba0k1Oi/uZ+Php0rTdzrHpiWGiOsRinaEpxaxKJ8CAE4hP5LtR/n2xTY+60wzQkUwHkP
PFIaUw0P7UIfLwA+Y+LWT9tbcYFRHoKnQ1BSkVeLlP1wgvHphgcPDptgLpfJJLUP2WI9sIRTjOHD
GOhnsh7PsnqcefNNz2IXFU/1XDmheskNkmR2QPEAziENRLteCU7V54cSDjgzjDyK8cl9Z7AMiMyX
ttFo9Miw4fuMJxE6TIPJfR8AHOfO/Qx1bzNV5FbpdVuLLZffejngZXwbR7V3IfUidKCXd1rHpI+U
EKNaTtSL2wyOMr2dgWJDWoxU8xKy++rcuDZ+3jyeFQxMEpPGYjHH4hdA40d/Yg0jSm86kEM/yZl0
uOz1W8H+GKjTzneKPei2KBivmr42YPmLhEiThiE+yLojWwy5bXN7yEBv5a53O+YUEXy25WlTKfir
AcpfvYPKWckmqnLnw8rDK9a5dfDeIabF3btyUtPrDgEq/bQI2n/fpZrdp4EmU9MAQPJl3vm5IAY5
M2Od2uNPNNNALWn5GTji5zxxKTCFcvwqu/ExAL72pL6KRNDkVNFc90KPLgmY79y98kKihcJquRjc
OVXbosTiZviHiVAkwDq+dPyFKu042zqkqR2e8u9EEY7GLEiLFPuBb+mkbjX69vw0e14S2k4UaSZD
H6TWGdJ4AQWGoiNs98Lsz2MctRtTEI2c2s+FYFskyyRlP1454cwYqNQBxJ6ycn15K1Ef9Cx5Xlbn
QUnjOqHcmoZBsaxygFzkeUMpjUCLdN4m/+MDI7cMFmdkCrRFuwzUWopF3Q6jStL2Pn+F2q6gU/AP
anMxZAPV88OXVop4tYCVAlIonqv+LktBEdo4VqgEOehLjSLN1WDUbqQJWLbdFyOtmo4tea38xtys
EoCMSB/DSvI12OL7ru4MclVSiq4HvBzOyHrNOHCRJ4E3Tbg+SzSRQK0a3sn8+ST1alZECezUIXjq
T3Lxu7cNPkOuPrYvZf/AwccqBp855tZAnCnjjyObbJgqS9RVWo+bSpY+8cddAQ2jrgRydQDupkRH
NdO+0cZuZ/XC79Swi+3KdPX0A7EUzocGBT/GfgMekLf4lgrKSZfH8bXHLTiEh+AExWUqJthQ4Kdl
9g/qRumo3pRzZ7+/g2+UXfnIuOlx+iEducAMFC/2xNTPE9PuFTAWSqB4hn+bzmKY4cwKTxG5xOnk
K934xemmRgnBHyH+ok/EuMq2VN4CgyCNGcIbPH3+mCxgMyGWpWsNJ9VMEKV1Th2dj0oveDHrjMeH
HIpgs+CX+ASKL2Ulkduv/5kUfYQp7s0VpOcbBQDDqq1LO2dsiCH+Bw5rrKvV2S/fpAQXMSm0Yv6K
4+d5TMK3khOndnD0bIoqedxMl2m7lvYpmJ7EpiZRY/RlA91RIi6UBZrKKSVSXuQuOXxT3M8b+gax
hNAvRaAJFgbHVhtcZxF4cdQC+VmnFN1Ov9vH/lMx/2qGR4zHrxNxYSVVf3U3XodMKl71rEMTXA9W
0/W4Ai5ztvPNaRk7WLoWe1891hTLa+Zuoed2TPXig5929B0sBdrBrZ+Vf9hVuABLhkaQ/c5wvwz+
p3IExw5B10SvCDKXQ2hGL3nTFs4lTdcXKJIXyvNqx99M1rygr9e0oW424awgOrBcgySy5WfCeQwv
xlQeX/qXAzKligtmIHY+E7pEXGLV2HSfMn2WpOhg8zVlnmCf9rwTk2xe+5VfA8uAHec+s8TGZl4D
xiqILMuNrakVegAlmuEnYVpBa6rVy445D9pedV+B+iMhY2Sdz3MZS7QEwxmKXvVh9QXHIvvwuBjE
qz+psRE0Q13eVjmDR+xTQU2FFrIPtY3C3wV4KAC5VfDaItVOKMKFwZvMnioqGEEpCAqEXIVTeMeW
wRA1eGwrIJs7vQ2oYtPCdnjL8peDKgY7EFXtg9fCHCVxIEOzYEc+RMlCbdtwoFU2aoOQJHkxP3Kd
TAr/MOWWoRRePasR3nMkBmbrmw+FTtlvRiKtedWU0EN233HGY8TGPh17uISe2seFIpaV482YPmfb
qeVXf9mWJ9KAeGb7tfdUBhlB7Dy+E5owQU5EGOSjNGiZpP6tugvVjJ7n+kK7F4l/bp/bglw4Jbit
vOxJuqfN0bNtuIvp3ZpJ/DHBj3DFRKSGsrlXyVRIPpBFAQ7K3znKgHBVIiCx7Za5WjzI8GzmHgxf
nlv1hZW1YhlN6IGjK1Q+nmmdKi/pa8bNUJOb5fza7d6yUXebwakM2DNS62TdygD5VsACJ7/uCoaB
F394ndWLEhUdWQU5iyHJ77UQcv9gg+eFo7cbvtKhdGo3FCQ6fdsRTTh/EsFUAAjvQObGS6KqWZ21
ZQlHkFG9SiwmpNHahQi6mlEognvKH5xQYMaf0tyymlopNfk8sJSdq7HrcNnkjfVTbTzCg8Md7/n/
ihTclw/l2IpCV6FOMwZjCceTYb4kgU9ZGgLS0f4FhFlFJFv9fPY7oOrGhZZ8ydixIwg66NpdxCoW
ni2sn9RMH9udNvcMz6sYw1shXykG1G+RcXP7IyJ3FERqN+52s9cyIBVgDNAVKyrZVxuvynLrJ+0o
eQgoEaFUWAo+AKNzwpjzeOQZsGC4YxuP/gecZdwGtp4884DF3zC3Y8c0AS3iSIESWAHYO+uiDbs8
yisaRI7FESKwF1pWh0UGdmSTOS44LIehH4isJcQM0ysOZwby43WDDan1ZHXNlHxIf6J9HCMFyj9y
+K3CZFNBQ5MBJz9uhIMtRkZPE0ensnEiacTjodlQiLUNKiV/+raubRMY0gOKkV/E+LzNJq2Sq76U
tkLiZ3LK61gw+UXFqLuFIIQixXmyj/IO0LiOGcwBbqaKXY3fpdXRP97vbYVD+heYDCWOU1By8afn
eUxYPh7OcyjBHfJiodj6vv3I2yQ4ShXidvZ+prO03cr+OyfnsUOLy38WhS8SCnfF9NIuh3MjAKS5
t4ch487BXDgR2xZQ68q0QUrY+OMkUR6PRF0osSt3U10HNqWk/HKKWAWERCcUl4GdS2KH/yl1dAVx
KiJGB4oX/XRXK3rls1ErXdO/AVhC/Pt4WN9euG+1S13bVaMIBpdpHoEnXo7S7cLZY22OYpQWt1Rc
kSmWdKtb4CFlh1U/YF61CiZX8XxSZxlB6W/XKO/4je6REdM6eVmNJ390fInJ9SmdXRTlM8QoivFZ
XTxf3zZD/xKzZ7qM4u+rpvthziKfgUHrtQCsIOrwpjdRAnSo8tRcFBTugwiuvLrZOBgIZDVNyUXh
i1AMSexf7UvNzolAv8I/nEbW7ip1Lph1+3HpoYBBACL6SyFgqSKJzZhd/KHz/L65FDhH0g26hAWK
07I3d9NEjjeXAyMp9XXrFg/P2pfupj3Lz7qDf7Fe8F8028KV3aQf8aNY6scuAGUTAbsk85ViZVAU
+5aHAfIUChJMDvONaFxE5aRHHVZatjoKiqKARDXP8Ed8RQa6MdydTLn6eU+f+OClGw/svpbrtqje
OMj8xBJtd2MgVH7vxeDglP1eEtqLwih4HwJO//LaGakgnjwTgZ5JYcvHhtPMigrYSNTM8cJfKxXo
ueknM/bMBMHc9+J7I+3ug8vuMiE7KYYRdgvS0YYKmmTy5b/aFkFO4cWebEAOSwcbMLt3oM28q+aA
lLWSeeC0Y/Sv/LAYbCVLOYrNnZBEBc+mv000x+GgerR426JyXPTtQk2rhiH86O7tuKsZ4J0aRyNA
iVt8t0T6mTEEPiRXcriK7/Pa7ngKWoBT7rY6I57sdbMmgX9hjws51s1qkrzl/J0oodjfA/6Cwb0w
MDFbNZfRsJmV4E1OxaLN9vGj6hYNMZaIWSHCSkFbZpQ2x7EuyrsqcUY0TfZuzoDajXhNxe1kbZiW
vz6t1Zi7TtPEL6lEQmBlKHJ4ffLk+SOgtSlrfnJfGxYHj8VV1mUzgX5V+5Nb1gO+ittiYQpYLu0e
y/PZsW4Ecof6wZsyvXKtQJKEyiasWwnuUrJb8/Q2YzfLd21FU4yuYjpQ02Ibd6DeSeL7aYDBOPQC
eEVEC8vyaiToFGpMLXCO5Kmn7T63JBWtBDHYzMbouU8rrW5j+TNP47AuIHGMW1T7FsPVs4ngI1GS
81BlrP4idDyt77fknYRNQkHb/mAq2XoBOpK9XQwIpz1ptJ+eIXVCTGw1Cv3JgbK0oXSJg1zMI3Kg
S7kdST+ctpDTgrPd7r8u4mwQ4BZOM24p29ILrMshkysYPAwwfJ2FDHQ4HRdXMNWgNEwXO5y/U1es
a1kpzOj6qJSg4CaJd8/iDRvB/LbUXyEpNPWSfKlICf1gLWreqBpZNfqDDM/F35ZFQs/QsToBZ73a
/16iNXoxHZtTJpNJZwjVOhmZcar6IPnBJ2yM301HkbsM7jxUNdLflz+vxMmnhf1LskFoHUgovMnA
GEKNxEbU+RgzoIyHwefMbZCHvYbgsuK9RiGX5IOL/AzR+lPUrrZq2bzI58ZH3vUEDVXWwYxko9Qe
yZpoO630SzQAj92hpMtrVRfTq+r/mjiVWNYKZ6vMceCu8eh7YACBNPz2uLVAPNuQsDy2eg+gJD5s
6m1TbzbX+7hjJdG7eQ3ymKUgqd6TVvFnSauHHPOGtLA77w77TVkzVtEOf2Bkx0i4F3rCWCXmhiO2
ApnsC6D7K39CIHI9bfqJITa9gwYlapYZ8w8uEAgSpOMmQxbrwj9PBXeV3QXkpe/vNyJNGsUqHI+V
WW1dFBqFEdzVbihtCCddPiAIhuqSzxgyQw7Y2EsHPTlb36aCLQaLcooyPjMIXN2r30pdy5cE8pQ7
b6K0fd20ua+rNpD/zete/T20lEBjVFfjZxtxijkP4HJVYzJILa2sIHdgfKboWXltNCQamIJu4rPf
/4BkWc37NohPVi+EbR5C2QIboEVz71m7/4D0BtbEgpn9WKrrQpVan1lpR11D+Q/Oi0q+Q8eXJJ4O
L1/aV4orrFymNF6Zn2kLExeR5ArSUDJSWzaO6PfwvRByvEBO0j9XCtl+6r6zpgQuwP6p9av/TK5Y
0BdqKChypvzywEO6hlFdXo7AuGqisJeLjuMX1dopyGGE+cR2DML6C9ZXon+m3gbJKSaWj+KqWUnY
FuJrkGppcZW8LAxNtoVMp2c0SYQ9qy56VaMtsGM5G7zvOZYkjpVjOCOYeJ8GkHpCwz+mv7QNQ65g
Ze9a2GnU1aZi9FwNSFL5fLMp1vjITRxmJ4APL+WaTVsZ7uJ5n2KOKNO8Bho0AONC7Dd4c2hDF78V
FJKExWqPvf++SEseNPqw9Ieopf/9DR2qA+0p8ggFh3WxNzjH5WMtJgxgX5X6JEtObGDku/Fk1yyv
zoaT1VOhzUrBSN6MJ9HwCUDmQOgblP24yMlmQCOHa+FhtMDH+AK0nSx1UyIaXJAiwkYhbf6wcM6l
SAgmV9EjmKWSDq4BSQu8SzT6KN8ERX8ZyDbUYqBcXJ1Z+CG6DtWUZSSvakng4MwfSL34QetnBGhp
xEfmJgfqgaeK8RTZGlNXj/LJjhWI8F1ppbsX1GO0XUn/4AtICpQ9MuCbZJ9Dgnw/OSJB5tKdRzm3
HZ3rPKvFSbrtog4eLvsWCZYmiRUD6mhmbX5lHJ1jsbThUIQ1HaM5a6q81fv6VCKabk4sQuKANJvp
cJ1g+WE1yoohMSzYwvYAxxYybmDlXdIqM6B+0iZk/o+sRV4NVA2bPd2mIVNbEz8cYY1rqoQyVqPF
2st/v4a4k3CJjo5U4bIfPixJzl533Cp5VtoU+IDLz/HiO3MgDcxQy34hksYwfGnDP2H4UP6HDcb2
Y//s76Zy9PVXj+prEJBQ0U4HlPyW8icZuHgoh9wekG5TsveGpN36P00Fu2iT1M6HTdt0Q6J+E1tq
WtwqcnTSxK8Z+7q98/0wRaPmKsNQcEu7h+rdEVZ5JeahrzuEqbGNGalkvZ81USZyr7sEHJkeJL9O
8qSsjhbQ+KkScr1JWBh2Ed1I85+PXKt0tE06AD+Q98Kf0zHoTWxz7t59iZkNPVZ0z3IY+jdnLu4I
EH0e90RhnQ08uDRUga6StdrxK70v4i4i5hCggnm3DXCHUda0XgUoJZ8CtJsv/TdBYwE34hFdCx1L
doPa8jEC0r2+XMKErwe39hFafjm+jSkcuaesiqNiKKIlygXCzBfVQM0x+ON0wNdSa4SmYkwuS5jW
B9U/C7KdOGbGlM7tXmpvtYf9OOTpq//8PZB07/c/5fxD48Uw7qvidEpCIHf0YewFHd50UQMncikw
NcGhU0384GJcWCu7W2kevd+kvq53IGDrxXTLIVqSPNNex6MwAscwqFcN7D3drjBpaAyMaHlPm0sW
0PbXuGlPHgDPwDqC2Gud9s8aK776l2bbkG4eJy3U5FNwUrwnNzcuuR9eINZbqYS0Eaiwqo88RFOo
7jqcVj8tvtSwJTXfUcrH1fnFye2KT2VgyuhsjpJN3DwJq4rkSJfQM0oWgo6hBZKSPppRHDF+sjGI
3mkm+Xp2sd4BP9bUaQtnKMMwnRDtUoFsZEYAi0APGAqnZ1E31xRZYhIvomWOjJf/PdCwk+bZGWoM
BSqsCbPioZlfz+AqlhuiaEeMlj8eA50L9Taw3kVuKrE8FY/i6wWE3H7o/WxoqW8GQp5ocoydPtTc
jdaTX+vqQIcenI3mUqvYnsW7sw27E1NkLo8iIBAL8dsTxJ1ghI+9+Sz0+BspBYlXsXXjQjfSoTMd
/J3BCcipKqDGbKUTsj+3e/xYsyq4HrAvJUnmNMJ/ku0PgnKNE6wFKkV04hWR1HJrZpE3fg73JSBv
fzaja//WcHgxUKLKMUVq4hPL7kC8EbFiQsPGuvsy5x9xn96cx/T59iQkEmbTkhOxWUFi9BQOspMO
UvbZcfJTRpSPpP1Zt3RvNIuK7x1unQsGGxhrZ1NfEHxFztQr/Z3InzszuwM1RyDrtt/an4EXkJLD
Mt1EairpE9D37yahGinIwxndlRWwHOsHn0EJEJIBjNbkILeOTj6YwKRqV7eZiOpSHQrAz5l+Cgce
7m3um+8DuUjdcaVN68fL6SnXrGX6cMJtFXA0ph/ofG38QmwSZK+aRBg8POcFCrlFswdelXxnpW9K
F3hoEKTzoyMxL9Elp8nSHMyVji0hnilvLCAkUZqMP8R5QF0ysWqvm57BQ0IjLdKHUKio12qKvDmt
7gcUVi7e8RWpdXHHZzA43LXirBp8VLc7KE8Y/mQSLjuI8W7j18tbZ9w5GgrlHB5sTg28Hh51ippb
zehqyGDUJvTidB2K66FeUN5PPwg+1+W4tDBgsiJCDPmDTgW+DAnohmrl9Xgegxw96Y4VDMiwfGKB
Wql8kZn/lNwLzhp3liDAYrDUnzVa+u0trQFXoIGLw+CYDzbQXHwgR0VkM2f7Mlk+LdqDw7UH23Qw
tRjVJ/0H8ToVwHNbuvUpaGg9t8CFKT4G5Srb1x2CtjB29K0OSrySeUVeY/toohUVxsrwa13vVS7o
ZLpJOlyq6Rxsm/1CNyjuQGgmukvVufe2ycyh0Nm6DbCnBJyUcqzHLubplLfC0n9TOcUCkx1tP4KH
uaKhTHSs2/hed455Ql/k6+pU1RnBep78Ipr1AnlWzju3O2UhQkHG45P/LmNFmm+5nom1zifEh7Uq
w6/gJ/yL98cGCJ36JV+ro5oM/pqqSq+cQF0JaBkTTQBrBhv2niWCYQYevV57dKy4eWuOSwZ2Cvms
VHfpUzwqtA+/c5EUIoI0TOxB3Szmq0LZD7LBnFQ8IxZyb7Dm2F7H5clMfpsiy+Pl0s68+eecOclk
KWna3QY2YeRJSkqL+c/F4iL9Tc8aRu3ZUiUI+/JES1CprLn0N2FlXwiPh6DDSDiwMgu17cY79eNA
hlOdth85YQSGigps5QazABPmvcfImyrwA/8e1zLu6wQEFF0HyQTjKd2HEr/+gi9jbrAvXoZdNEYv
MwOJEzeyEIIw4+t0DCYWWq58uqes3zLv5Ib94hr+QDB/wMs87/fRXGoDrqKzNZfR+X7823wRHVNb
i3oqIfFMDONz56yDtqMFFWrCBQl+UuWcvOdET/W7DohDNlQzngPSw8yIfO4UVwUU2VGib30+XLL1
74hDyuk2tOWK23L58AruAiSeBai2tTjGo5UqKGbD3032NHDMUgmgowVjJ53/YMbJ/HPIsb1knV2K
jnc2uvNSp9IR3WDjSPGmBJSVeyrX3Tt/9CtVV/a4bQg3BdUNAM3beP59dFSiKFx3R4ufz307EFX5
89VCn+bzwmZHrjRSfTy75WuOX2h7YGOgQru1+M02B1MQW6sxmOFgcxP7Yb87qpP5Zkw+5MYrdr3C
LZywwqujP8WfDSYcZxTuS9hOd7rgK5KekNr+z1R0hUxhD/gstZT35g515simc1rjG91AOBFfXz7M
AKaJqO8NiuKjtMiP8iirxi03LWTU5AKb/u/LaBLwiDXjsKcfzBNlCSA5GPzXLp7SR/EQ+O933Ehg
BrC+wY9hM1k8/ARriDry7KwsQOpZz00ysqBst83t3U8/WDIh0KrW7EvqClH6nu+AeW1WY7t6gi/S
7GtVkkq34MNenCH74o+TNy+B9SC3rstxfQueIeJB7ZNxX7tV24V/B0Rhvw4T4mcQGtKtIl8RozI4
+XioSrGm3TD8Ot6jqV/PgiJDsGP2MHfQKQDvNSJNYrvWipGyjyhDxTINoUeiDQBKlQVLY2tDMEcA
t9Un9kwYoMiS0g8h+iqdwTN0rvceEF1Homaxo5Vm7dDR9Z8ig6wz44uls7jsQ/b820K4IuSOlOBp
zPpEaJ7QRerr87R5gyXdM0GSj0AG+xziBufgf3Ucjv0xXxqjUMyf9O6TXPHb9FsS7i97kvMZoV+b
kiR4n06wl2y3c/UKtv0M7RFvUKoBxBEMjZUX7dAUCdT5FWlW8iuWcdGXBki6hGT8S3Q64N3UPziK
KeBwaXEynrR/mC8Cwh1xiEDs1nA2I/F0BM10rYcWuR+74DaBnC5eDriINzwdTugj3MaGrpWEShiy
01U2Y+PjiAsfFwXUwt3UfD6534h0YL4R90puks+vFWkxB9ukeUXmoWMZcztpcUR+NnJ75CBYHyvp
7GQupF3vlcCFKvS1wicNMKUD/eLqxysMuOmm5bZm6a5jn2XM+vk/mv8YgXNr1YSkqUxsNyshPOf3
G7xXJyLbYK0OibL+JKyXFxb6qkN2EGvvJ2FT1tBElQumdGT6bHnVLx2aLL6Z8tU1e4CIYnc/Tx52
RMnvleTTMO6tCQWD9Hcj6TGyyjs/12VyMT9FaxqB2c5zaMeA5t3J3ofRPrGmATijRNWaI9Aeju78
LfIYXxtyFdqVkKYOeJ3yLjvexty2blLCN5atGoRsDRjaCxJEaW623i9njqhA1UQwtUZw1k/DW95L
h0Q01txa2iA8GmV7o06si6QEMvVjFfcY1kBjSg4LlZfCRoq3mStz6rwSgAUfu8aQMHacO7NrNSps
E8L4JNh88vD+4pDH0zIY8AkI9sOdptOTCAfmk+N3Uh3TuHp0nNqJ6vgdSoz7wAhSL2xIFzusoHBS
hdt7SN+qVHde+Tv5pjeXpYkrWCxesfkZc9joHHAliTsrd0Fi7qWdQNmgwEpuH7xmR6IWKZVHq39a
fJRQ2/Qp1cs5ulxohy75w4dhtQkuT4ic0pLppT844+cDbaaOcDlfraff8lZN6DBMv/0zXTw8lVgo
zF/gUBmh+SqY3FsvLjClL7gVEuxfemk3binHt1Ep0WA9ZdlIWSEwfwoh5Zr/UyMKp0WZTdbUuEJt
4c+K+SmZA9ELODo153tN8lfHrF7Q6IZENJyMFmgLOSNJaYjgDH/xnj/Xj++26t4lJvjfXFwcnlQi
M+e9uwsRzvcDOTpmyArkqATCeQS/kdoOQeU4rJcPMfnLpZJAPHcSGnnrc36iXG7E8cpeWyF4aVm7
6WXbH+EQMjXmAMgRl5ZoqrBbwBXW4A3IkiAreDTqvjagDxGOopBiSWCydwLFoLVi7vqUAB6UL4nW
r9hUflga0spBhcibvScFF9zSwGaHs+l7Qd0R/njvRSd+LUCW2CfLZ1CNFQ014in7DXPnUBwpsyru
wE+Ca14ckQ33mL1KNiXNZnUhiPzgtVhAhieo1+HIS5ihtKibKTtgR6RL6KeliPREQgXUY8NJftwz
1aoIt+Jb4qaIZdaLehM5yMMAB7O7P/O6lYn8lICcCISDMqM5AIVyx4as5y0nBME2PVPkgRG0/6h4
GeFVP7Dpv+CJ3MBCD9I5gTxfcrWzD07bkFhc4UZKPLr9qqaxwQFxK2NnlitV6uzDfzKko+1RKTsT
3oeXp8oXFPxQ6tIp3jhCMnjngrJY2U8BlMIbDBMjQk5aObON4NTYJZktOOCA4zNYaEeidboyqVKF
dOpuCaUUx8Cr39v4JgTrlDDiM7yEXerzi5RykD7rI1MXVB6WKeDPmKFN474zDTiPcQI2pDbDRkY+
rrl29BCHNRyQ2B9WlwfmdSNi7UqV7wUwycx76wR/kn/HcIaUhbKS/TUk3mex6+ktgNj1Vm7x0zCq
BXWaWGo23MgaypIbs/oDK0h8uLwcZfIqc8xBi2BBlIBR3NUtcqQ5TI2broGbuyZomHxiOOfQhUES
xNfU4tktLTE/CpRnjHY21U70kApc4pOpzYeZYjCcPlh+vo4/ho+OHklYIGoQt0W4dUrW/y6RgNSm
g887GMzAClKTRW7rBIZtl2lQOsniTPGwudMzSgeJ75vhYuGFP46c9P4QzKeFmX3eXqc55bEw8COK
rhrNkQwJ1wnSwD2fjmHxAbfvxTjLneQuIDU5v+zqqwOccMoVVmFquKCh1+WTLVGQ4GDT1dz6Aaeg
sM6yGYTKEyyn1QBOrkQA/n7AJCTsvjWAXUdffDCqEKFBZBd8otNJN/ifYQqrzZkDYXsWQc+6cV5A
woptmmYvE+YhTdFab9Ldw7U6/wVxE6+c6/2+oBFzZ7QKDcaYqVFDsFEWP7E3eNB8truU1NjENqxS
3+jk22Gx7Pug1wRgwzZ9hjlEc3AMKHO8ExghavmF+4YL+K4dgnZXO9frRkHVsIlHs4zW/wtdGhAT
TRLHfS9TBb46PtijT9hVRqb1XcMRVWe8chjy8Djwzx3tMv80xOxuG6XA3aVEtZ5eY+T4/hHRrKsI
lVi/bjOJmrNkgJ0nMboIEmqUDDhZ6O+zdDJJYnwdJ+2iV9Byqc+QxB8FUoWuaBWAS1dVynR7Vxu9
5c/ozywdgezdi/EHhg3MOmLP8dsl/DIB3FWS//Y+syT51JjfXyIgrD6PsaSTocwV0VnSvJC84ay7
MxybU5/LJ7vi5GtNZ/l5DEA66Ym9EthC04dVMwjhBhqJLkbMxQ9/RZ0owcsykvPuODDSl8OOvn61
VyFKPeRo6/s95vM0NyVuYHg7y3xuTmKn74wTxR6hvcAEb1tzWdLDlRKWa+C7a097q8nESXlLm92Y
U0LkPVh4IP9Na9PpOin20NzqLP0ubCDTooIRUMLQT176d0L/TNNOGokoscevnYuW2Xyw9o/hfJNl
dnsx55NGArPocl3rPd1MH6pggvtTXwPUl9wWRFIcWsK9wu65/imw3g8COGBOtcNHsCrtRCeGQvr/
EwvXeJWmyunmqvgAWzHg2pnCKG/IX625NOj0e5aFikElccdJjn9r6IQ7wW2hsm6qdlPyKz5ibd4G
Be3giGJi9XKiG9XieFJ5vtJWV11k32tInSD4rGuY0+7ASwFmM7YFYCwlKI8ch20PYJbesJtfV8bk
NaIt2d9iuzsZY0XZQRfPRzaP0UwyJeT9PEbQGEkR1hauQAb/DIYyEJJcRD/YjBGg9hjao/dM4Mf3
9INMAd9ffury5LUaU1HWjktsfzj0nERiF/envQvMvkf9xpUqTxceii2vY084s3r0v896CJSCqRPZ
H/Ia7jgyRnTwoCiNAAK1VSQZwHc8LpGQRtLNF74ckrS0iBJuoI80+0puE4FyqL9Zk4bCXeBGiUhC
UAZfuVJrI3J+IkwDyukO9ElDNl++o4A8FohACMv+Y6jlUuwK6T8JBkoXtgqGYE2wNYs7iNxMn0SF
ljN7opSb1tRWcriwG2y3PpWG9a8sezYcvYmUCqgK3cGO4y1wZJ9M95VGwSDCWmZsVH6DQm/dc9Oz
7Nkh4v9RPVMuC1ZTvu+Z86gha8/yD92YUHSN+W4LRk+KvTQIHrZ6jtrXamZ525h9gbwfaweTaiHy
SphmMmjd1hqvuLe8HQ1KioYjRiqZdiKPKkqxzBWruuDx1l62SDrNbImgFi+SEnPRtXugXhTKW5xT
/ZQpvq06jW64adQ2h0dAoIrAl09DyQworpwoP6NoGMe1Vp0HQ9piFZ2bJaIptTziZleuQ/WqYL7i
KyYNCOTmQ5L9pGrKCYBnDYKhKaGw/PEEasl2GUP4KE5Z0PVz8MIaDnRPx15dn8pneVuZZj9WzDmz
G2u/7ZARu+YFoKQeeQ8es5oMPZ0r+REh6jv2jcY5robdnSp7/j1hsLIJAU+7QHFRn8HdHWQyWpnc
sqF6NpU1bgelmJ0JhBkj7HfEWJa5tSerdk9E6nbWVRYHN1yYab/e+cNdBqJ+7qf6Kx6OtyScgM4N
gR0vchQo/f0mLVkA63w4RYW3c1AWnv421u/XXVobh8RZVSy1+etYIKS1xz9zt/YQbp949VKbQCbR
fNek6bNZtdbNayvSLP857vTF3l0BDVY3vMRBNVgLWHdF0TylpW7JXv3YpghibTqjK1jsx/xHN4s3
3c3glvMBAds0lzmZRbuXiNxRFyNh+qJ4AZgXpEnoPBeoZqCSNyOwxcY/jvwZhqyJo7NBZ8aOBBiV
vKzyVI+g+4Iage3IHUiwBlAjYL6jkNBZQhtUVxiWSwC9b+orUqj1pKj7OtHJfu6M4QCJbYSJK1/Z
Tew0gsng39hybEHuziC/66bmJJj3+LPQ18Y+7kdkM/XEkUsU/b2LGG8tftaGSOSeERR58LdvmccM
ybGsypu0etM0MttjCgEhvsZ2/el1ENpKAxoU+/Isv1wwXypIgW7G/aq9yNcLSNB34t5YuWHgo+uu
otzsMv88EmMwZo43tUeDI1g2Ien/QRiL5s7CuTGvVfi9zqICs75NxBlwr14sAU8gfP9oBvhJHUma
zzI95L/bozRahLYIlHmFOpFdV68kqtfMw/Xy1nwPBE6CBYEDOhNdJkrrJG4qvJfA1AeEqxQ4ODX4
BGHlUsTIpYr7jVPTeXl0fjRAGGZk2lQzo5ChMu+5daRbcPAr3FZEco157TVIbh2wsYGicEP19Pi8
saiGnBMnBu8XGmLYhe9uXhMPfjUY/gDMxPjcFB1rVEWZ4PFdLscTB46FE6/KzfEB8vPxi7WAEEZC
7I9E+burXxC19U5XWv0HFrHMO12m1XrYk6JBXX/4dx3tXJyZiHG/yU14bKb9wDGODb3V8XCTk5ZM
qPD38UrFN9P7a5/dRBgri+iJZywyvtyH47I9AtPJWjQIM1RakItHN3YrPrS8KZrXXWkSNtQEQTW+
XdicJz6OiH3FU5KFmQEGWoeVMRUeUmteaKlqZJa0EKiwXeyp2fiL/HJ+zMgQ1zVSFXTbyJiCVOPn
Vl6zkdW4XcWeD1wVQijOVQ43rigcaNeXeNO6pD2R4GgdF4WwacxJj8d/0ngpoHFrjvVWLEiMxg2G
6KMLkJJFm9Yryk/qwLPICsIky6RLNaCGyqMA+DoZwYtDOWBMJrS1EZxIVG5R6Ogeuacz/m0qpDtx
CYI7e4Qk9/LdWuqD9ITW7+KUau3Jx9xhkSv3+YTJM8mhJadTY15XrfaX6g58ZSRT+q0aDQIoYU9Y
2iUJkRa7ts2Ixd/9x72MC9CXCpNFMmrgMTo6Jw4UAGRCKi73WzmhO46mnqbt1O5KD6CwM7c/EHRv
jxiNNIREBuHpXAGFbyVHDLB9Y3lC55JFte10is0jDGduAj1YOt/aajsNNoJYpPrhRax6o+s5o8Pu
q2uKGBdOsnAzXnDKKhLEKpJmpH6DvFKWVAucN6SIzL5ihXCbvW0PPmuzDt4sV5tV6oJ9Gt8Rj/Yy
xSIlSoKU26ESQxi1IronpB/8yZalf1PGSfX/QOPujuR6iOPEqVSooXp8ugCJ8nMepmEa/+IdhipR
OVpc/fwrkUUfWg+nInz2bRwEt5ZQwhFa1PEGq6khUplHo6pkD6nBs5dPulBm9Vu8Mf0twoY9EoeS
RAVblPrM/BuIdVBXVwVeRGzPwvJnHslWNdhDCyAZWdUTIUI0C//uTsr5gbWQn5qSV1xa9+ojet6R
CguiVuHZUsldKSLDIijuXpU+M4Q8+IugQTO9KOMVYDiBK8q3u7jLETccZ+w3QsnopdkDQA99ClTF
zR0CyLcyBvrwFxYEb8MPSh3rXVrx4Lc685cWY73xJEwPkPoqsOsDhgoJTmxvIV6l1BiLNj7POycL
RlaoqduNCOL4ioC2HBazMuHwODhx2vBMubOUC3lq/Qrtn5/ksCdjUi7ENVAc2pC0EBctI4kp5gMM
aZtzg8duO04oaFt8uAOETX4NVfyRPlikfhLreeY8wtVjxfo7+SscZf9glDAtiOiS10QcirRJmmFV
vjiDmyRiIwRUq1Up/VIKSn2auMqgXi8b4CyXxdjYxmM9BXa41fQTr2vYK55CPqTIvosirLHVPHhZ
6aNv5bkQ4LMdKDudhJUGyPWyOnrEkZhUJIm/RwpebrRti3ZumZLCUO5qiZyox8DebmvdNaTN9AZT
VA+LuKuOJGF/an12Z0zMOiRWS+/XQWS/XpQcW+Uhv68qdCaXU1/aIOycPdjpW9VJf25cjZKotKjl
IC75+VtTBnPvMmu8yP/2nGuiw94KOqC8Z9TMdeE8aSZwRjQ0y/I7FtbiDgxTapsks6QPVg/icxLE
yR/0lZoXWmMnOuhHd6wbdcYzLi6y79NDXuH61Tm+w8XgSqWrurJKIHT5LGwweVFeBKZqC05fAoaz
J//KM1Kbd2MbgZYLQeHpHgTR/8vyXwRNkPV4lxllOvyowg7c8OPWax2gESxFot0L8qROY/fHmfzV
J4HNG+RphBhuuu9JjfCwbD7mbSJ+47LMT5zPrxlLlzpIOWo8exEl+Yaht+wARzqvUTt2B7WE4eaY
47dFolvC0o8j98eisgO3mCwAhfpPEFz0w1Sgbs4iQcWt3smQoU5MtJBlD68Unzyc03FgainAKdwf
8crPmln0fPCWhqIXE1bDJQx+MI7MUt8uc8fN0iN6caaETDSeXgpi72mMrTyOe2p09dDeh3Y0o6ar
+XHOEfXtkN5K930RV2kwDL1Ilt2KBVQbwCaZmIPOLORbZnchHPvuaL4bGSot6kzL8/UBApp34FkP
BKh5tAqK9wbAPM6W2/rJDqVsEJDkkrkfcpcpkfJr/jBgFkPhMYVKdgOg4NG+c4Rl6BfPRvmuivIy
NaPR4jRBJpmInt/l2MVBvSaGqSZT5Ce+qx4TL42ozeCII+NGJOlhAzP/58icvG2DJRuz4CFFrd0z
aXejJpYb5kQAkFXpx5xTt8H9RwJB1hOfv0yKR9LMmAbP9TxFt9vqS07zecZAP51b8LrqPmTec8CJ
NL7FmoaIj39wFcGeSX91p5StKoOn1Nc1FvKRn2H1K1fKWm30G5jg3rTiT7OIOMdqEz9N62S2BncJ
rHVHnfthrE8KUfgfLMPa7mq/yjHOqGYkn0/Wg99ZjaNqBBUe1Qb8Fyw8CJSO0OR+TRdZJgk6xNak
mpjiqARApVouSeD2BxTXm5GvAuoJovaD36fp39DgnQepewNLpQqtlKFYATUnd8cdKbuVho3C3ipb
LcfPVRK3svxMJTDBL/Nd4SJZhkhTV/MZD1VY24L8s/ph8l8kGDhTYUDOzJ2YaRhCudqKv8Lyd38O
bxEmWx4kId8tlUdnzdxx1AdxbgPci2UUnPzThdnc1BwA4ZjRrKh91c3LZIUxMW4seoTCyxVwFlfb
Tffky1E5AhYTPl32t1rrUBWw1sElVjsY711jS+Rztn0eu6UTyTkm19zYQud4P7b2FMbTdzEq0167
XiOwKIXbHGDV5nSBgXNpx5Sz5secIj0YNCAv6/Z3d7LtlsZ9N+e5TvTw1SDE0fAe9OMRJvmSfK6u
VuPqwUR5HTrBXFz7APfmg1Yu4jqE//NVzPzNiclaZ0PlNnHD/JZgJvDWjdEbR4H9dMZhkr4aU2oo
VfEq8pDA2QZrXMQLJfMl2Cj5MUHcjrzpJGqzQfRXSE4HTUc3NZHMSpYwqR79HerF3nKj6Gxdl56k
kjtQkOvDAZU4l07L1kveJj4cPz50T0cRFG9cKV24agJ8aR4bJWfy7rXcwL8M1Og77bMRVG56/OSo
bmuk/Tg4GagTLHKXzXYjL9ncG2xG6lAAkNHdHcV+doHUmrcLmYVRx6aUNhEkZb+5tKpwYwV2zL8+
yisYAJOskVSkJpI2rnF2EH9eeACH1aWsvkcaU6lznoaQmX2Q6A4sEYs4bmIQrSC85sxvu0Rlz885
jyBp48Z4FchQcaO4Xzday95094nvc/hzznq22ZBHSWNYjIZJ5Ex7FN5Lyrf7gYyE7DketR3wmoUD
zFq0Otd19PVcY4L46L5F17LV0zwi4JbyXW2efNVI4KzAfbzCLwM+Yp1jVss8yquQLFt34aM6tf6j
r0qcVVD21r9M6tXvrNGzJCbJ9ym2koqFWdN5VGIXris0hgJZ8qZ8xIHHxzzqfNkmhepBInsy52qE
uw8PAsTokK7wpRLH7j6ljDV4osFYqwUgZweIwVsNK9VOuKjGi/iFiKn3j0CGr9IvdrrSAxTDZRYn
T2HV3uJAOHrf+nZxLf3d9HD6s8NtDX6lst8DwMuEXV7JNcFlaFMXUUYsxTfZh5gjjMXJRGqsYwS8
ULhIQ57rnIiC9PwEO7sWpMuotsxBL23GDfEOQ3uUQgPsQ93bvNwlWtS0cl/vlB9He72HVT4smxDc
l4muzgWSBU/Sp5QstbhKGpwdrbB3RsT8zUc+cF6XiMGPvKAO9qQX8l79jMvQQIvHBDNicO9Papsf
lhBiCxcQbMvIKHN1V1Sy2qmBfpk1VGbZjEvlrbmDNceRyxX50tRFAtKzUG+NsrXTvHfuXS4+itrd
wKTBz314vBViB5jo4LMZTQx+UmfEpu97NLsE7o8kxh4qeGNK/DVtmGKJ4YlRF2eybcDoVX0nycFx
nWPMiaEYHACxf4v/lrOd9nRkq1FhbBsHg4y9cGbRtyb1Ks/3AaECenOE1rscmgAckgN4a3mueLyR
dzApGoGQn3qUGdHu39NVF84P95wtTUXlRsOiZN69SPXAvwv9KN9uklx6DVw19FDIYi8IQTSIFGmk
91Qgtt/PeJjTbBeEXiCbSJd7ZCGSftdffz5FIKZDm0YRuA/zpYjSKvkHPp9PHFF9SmjlZ0vuWBax
HtpZ3ymafzvxMW2qfLW5QTV+24JV3k35gwojGcFVcS/foEdk6HPa2YHot6L1OlfYgGLE2/wt2NjG
5IaO3wKbQG+JYuRe3j64vJG4EKaWajEwuMo2X0agY5Qqa8EEZPPZA6Gp3S7VHBdLufK2U8gePSsO
uqLi7ftU2GN1uT8nffJNykk6M7gHPTDfEXKzCL4W76t0aI6y3yLDXAzZeJn5g/hqvsJRB+621jyk
eoxSahWxnFy8TXq/OPGUSwj/m+VqNSomJ3di1mp9jNF9y6NPiT00+P5SjJBAK204Me9u8pR4MeEi
X5LhGbFnjsYhtrhOKuUuNrx+imluHmM7DTAWAhFEYjQcObAuk8ZSrU0l2Mnjj/HIdRD7ff0wsmWZ
gb1m0yZUDc+UI2aWloHWDc1IlcT0qoyJyMc60RD/xaGSOvP2ttA2NodwrIH4z9BZomW53I/gyKOC
W/xvoQE4Kom0Zz0uh6xii7yTQ2qCtVolHW1lSUqjLExNIWfRwMJ9FaCTgwnNkr2xZaMC6EBv3TWa
rSzr70TNfmHUh3OZK73UfNiDkClVIkdyNj14rz7Oy5GcqR+UDGap4DnCSWMaRArNsgW39tWDeKl8
uA0Eb79ioS1pxiJ97Aj3bjf9pMZ7v81uUw1nJJzLsiJNDC1UT/00wYUE29WyW1MjRwl7+VgSugG1
FIa+o7CHJuoD4V2VfdO0fdc6XWNq7lcygQv+ru4x/E/W7tJBxDn7nzxLYN7DG1dATRqU0MaWHPsV
QqeyKLgyoI8X7/ng5BOraeymGrmerIXBDqrKmgnoLbMtbrLUNPp6Bshwrf1kb+dfMDUtArVSc8p5
/qxamJcpJls8vF77oMLj5Wdd3ROKsOl54D+XhmH8CJtUuhmxPqexYfL2mlRw9Z6DM36iz1BKGOmw
U5NjINlmnMKe3oO7HCwC2R9bRVoQvJGtS8rEv1qKEPxLuMw9b43g6n/GH1HRJQ89yYU3W5DBA3pD
rfYXZR3CZ+R3DU36XxTrPbX6Z5x64Tt8Ifrjl/yDSyAgzQap1CIASGrFGLii5iKbKjiMshSJ/Isk
fPujyQmN82rs6INiy3jgI+TEYIf5n0fvKGeHCdv4E4gTBi3SAPsY1AbKmIy0FJVkiVPI5Nt3yOVR
6b6M4QD6wMR0BcxL5y60HBXwWmAmf0/k1f+xetljUH1VdXV7hAGYInC7Xk6+OTUXJqxrXErf8UDF
PaZ60SBkuS5j5GqTQ0+0kJfSoTFT+C8DfB35hPaiufDMSc+zk9KxQ4czbR8mTCRtjSU04iY2o7/Y
VglbX57u3Dcr5Ztn1ofUhclKPeCsJ8cb3fbGPeMRjdaBpj6h62ik32ln2POUpDgaDNBBDdBIEt2Z
eR8yy+/pz9+EA5TArsZkFSc8XQM/z390BH6RFDONtp6mDnQvQgNfzI2zIZ1qpD3w9pqSr+GS+wKj
Lsp3QWDGaCuuNW6bIKB7Yg2pi+WJ7Uj9vn47z+/b3eQEnmb/lROeZ348f7U33mFvymnPJTB0zj8t
SRM59ZwO7hOUkEnewMSxXH94FtNJwx96FplAsaUHLFuwSvZUsFV9uiICMzh1jvv6Sa28/X0C+vGA
jc/VvOY9xHOT/2kSGFZFQexbMNPYD6+xQHxsUQtAVQVAmoTAyXAC0ocejoEUBKUbnjZu/YtkT7F3
w6n/dFJ6uyIx0TWttRckipdJwqT1TwKZcIAsq5C4Bae9xg210wXOV1uu4l/wmqKHsBUqf67t6MJ5
KSljgo9xNFdX/ADU8IW9fqt5MENPpTwOqNpqLUrxxir+h/YmozyleVS/fc9xMfWXMoUNhlPSfmPZ
Hd2NaxUU2YRx8BPQnBzLcOaHeNPFE6AedMHAQMAhEq1rmQLenInr6oqsOf/wUj6qKe2tTL5JmtQo
1ffRGVm1XMitKL253a6/czABD1Q5UT7Sp6cXos8D5iHCoW4F4GSgICT/IqNiTxmHrDJfYdQ7Z57e
yFyqK912nU+x4bUYGUostzide9U6YHFwVPYPNk/DukwSkHbKZC0vTCrwV4JDUgz2GXipPv33qD7b
qzTrwL/GNRJlOG2l9d+mVg8NgDpFIBepwP7uNDymVOMn2aXsdVHWYpuBfIkIbILBVociGpgNAC08
E591/SAS+RPFRnZVmyGhYV1iwiW/Z3fBK+khbqyBNI9/dTnXSyvy/MDpaQ4cKJzT+b3czVS7nDim
BBYjKnTMeAMP5VbJbX22e3QbEn96VJQTVFNJc1uwGQT4V3nLD8IDd+EMJGmbBSB/L1CCywfcvXyb
ui9ieLzvF+SU4l6zgAnFRf6pTZOJ8lkp3Y4L8g/WIQMa44vh+6w6S+WtMM3Ov3PNqCUz4b75WGFM
vENJwTx8teqjZm74ISsSWFXU4pJX74RO1p6dzjMQa+U6rm7C9bWNBaYQUAM7KjKTX2PEqE8paTLZ
M5NivGEQRIUrbsUwZAVz5XESU4HqV7BWZgMXGiu/oEwOieDzxfVWD6+yimgYwZjfXrFH7hHlg11J
eYAJ4YffelxWAJkG5fEdzoBayzJojI4FsgxrTPrWXtYTkA8B65UOG6PFORzGVgjt64glOH/YqAkh
TCJOCnbF+9/DZZ3ab5u36q0hmh4H12XzcL5MV6KVUuGY8jbVhu23fQ9Y+oBSm2HlM8fUjBUbRrsm
Aj1oqsg92F7++pZN7C8GOjoeQ/Bjkhr2tPGx6kkGs462vAHsplqTxWKO4Q1G5uYq0WpPWZ4KROZE
APIusvI5iOdXevMnxgpMsF8GL8MUOB2gacATl+y4mvjnpnRb0dpG0R23DTMjPoOL2pEc6UCbdDSB
4zPF+ot379eENvDpu7hp2WqMrpgB4m/U6C/0xu/d6z43Q9gJAIJejwgESk2RPZdidumefN5X4ksX
f5njh2/CYUQzGLECDHVCjDJu6SSS/Q9YmZGFUGJAFqVo2D0fvrJPrliSTZojTNAmrvPSDvUmvkUY
QQ==
`protect end_protected
