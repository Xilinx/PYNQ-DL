`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner="Xilinx"
`protect key_method="rsa"
`protect key_keyname="xilinxt_2017_05"
`protect key_block
F4DMIUBOruq+IzzSWgY9B+WKjDh003CtUayKKmp6KCPobsmWKPcB7q9xmJhH1aWojhUGMaj9EJxf
AJgTet/aIYPgs0vtLWvt+GHUP17FRg1pZnIfBNIGvDcmJbBfcAESov69P9ojgsJOQB0ISQz1BRsW
ecUC5xjYSWAE0v/yoeybYGcxuzDI7ZwHHl5XYUWztLQM2+90DSFmIxysDDryy3M4IcsGukyyh4BB
WbRwfbdkWMOL2kI9RNzRyYJC8stfRpUuxzXGPFadyqlibEQSpca28a/GOyG4Se1l0PnoEANCFnRw
RFh6XZi7dblG63f3zhxe+6Bi3NYm5NKzSrBJag==

`protect control xilinx_enable_probing="false"
`protect control xilinx_enable_bitstream="true"
`protect control xilinx_enable_netlist_export="false"
`protect control xilinx_enable_modification="false"
`protect control xilinx_configuration_visible="false"
`protect rights_digest_method="sha256"
`protect end_toolblock="Uul5Luuu8Srn/dR4dNgKDbcjqFZ+LAbFfFhIAkWHdGA="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2330688)
`protect data_block
E6sXewJSoTA2ZTY4s6UVs4oWc2x+dboOT2fR0dpSYbKWpFWM0Qt0wpnOC7mprnT+Rr8dr1wjryVI
v8OARw1MiFLp3/UwGWvEukahLDtvDC6c/qsZZxKrGcqgXOenXMQP7JYMH6/xbrvJCHFdhecdD1zZ
2UkqmYdHxylzMNl0XY9smlfPN6Nf+HmSCZzTqwT1vpZTYZqMn3Pbx5CPR3jQcIeV4zT7zZoYohRW
3BjyLPHyr+QTF/Fx9I8R79Mo+mgjYPPQRe2H/Y/2x5ZR1OQf97wD01pRyGoEbcODpKiaXPtxDm35
iX6YTgaaufosqMkN/yE2TziTtpsytbM/PJ/Wk8+/+IYeP6WEpGyP3nCt7n1A+FCrcq/rtK5n4+ZX
T+yZoi4R21aV6bBfalY5sETYLJAfrQKQiy4DgsdDAw2pAfeK81d6cND2y3hOcALoFMItrGNpcrnY
/IAwfSW43A43pnFqxjJx1M0m/M0nYOeHuPyJOsYLHResa8BbsLJKD+fhSgHd6wrXcZo/JD3q8AjI
qsV74VXxSM7TNhCA5ntur4wAIZ3+Yd6BHQmnXlISgEO9iSlkHPjvfCbraPBbiubnNi1pxCBb2Eqs
qwlOcGwu00blbqkxLhz/BzlmopV4UUHBBMb+WmgnuWsLHqsMJR/kDpIBvi81q9sdZd4yzp0TYf6G
v6uLNvCeZ1MnEYe2i2/6DLVXeX7yXFY9y7g6GPW+O7Xvny8JDKNFkQ5rI+PYO0LSgLKp5nf+iyy2
F3nLWZEK0xA2uE1Goo19PNyuIGKs25GrGrOZ6kekfF1p92+UhDwptHUdLEGoL/jCnY9w1bJlr/N1
/ZGNcL7F8Y+OELAxlU4hmguSw+x+gOtsukx0vkBuWpXj8BX4HKp1BAu7xwHBNpEqTpvpCAA9CbnR
Vb1W774ZRQN3Mncrsb5/OWH7EbulCGNxvPCkBj2HjFG9fEPX1nmGhLJ67UzEsgmjkd6Ixj+i2gma
nSpmh5qeGbutUAM31IFw+pK0goitXMDtok+KeMqt5xu12vti98iid5vgNn1YaIFhUJk+S/oEbBh8
O2pJTzSeklgBdvHwyATn9Vv4h/q7ClnFLJGCYCZFa4DkmKCMnrSWMiGBhjffhhU6Ig1xGoYqry9a
9zxJrSL3oWOkSbSkjKG9fAPPQL+7g+Zxkj3GvLZ6I4bYe7BZIFFQAmafVAMMKZV+ZIdLreQhF0Wl
7/hFvKeQ/1vZHBsXM0xZUYacKtgyKoAqJczs9IqTOaco6S5q5UO7kdQmUNOjR6D/LZ0KzJONZNZJ
eUIa1B/9aFsnF4+J/91TfCMXN9IXbh3oTqmh3Ckum0NUkkIb0PzsMH+u3w9x42/JpJQN3ZLVcILY
19eaGTOAKEaVEC9b88eZfLxsojwzuakvNvKObEg1160Hgq5hZIvHSIOBhteVK9tEqCGLvdXpJb51
IA7n9Uha0HoAQTjxsZ/TMFFmrH2ok+T8Oium/asYTB/k4P2Y1BHd434oo4rJpp69HHPfm47bRfQe
Tu3BzsOm+SCLhNJkvys6wRK84BrrtfHl3AE2xPbUoUq0VhHllvIIcIsxi3Xdow/8ND5MbtoaxHOS
pnOowaXCjIxINsrk788BtZ1mMmRdZ6TGMkDo8tQ/LsM/UYlyczA38JbDRECs/MMGCkfIJDD0/Yzl
xT/dPK1gGYC6bBpPi0Y57ds60cdWDgKwy90zM0XFn4+gHbqxZZQq2aRVcGFB8Ksa1LW8fKxhmeyB
IvU5aup8zcoM5fVpn8yyIeZranhbumyEDtPU+ixsOazayY5EX57q9LGjEUxmJpEgO/SLu/FoL7cA
KKzHlRAlOV/0jysiES//Z/vWet3hsN8gTp1DY3RbBfsnYRWoFjKGkwkbs+cYDYdxEbHRlyrtSxS+
UqEkI7YSCJU/4dd/uBatMmyVPImCPNcpqGMJV0rjqfYhrr+mqWDDLlOiNja/o5D/Q8HapfGUVrKV
ORC5FmhtTio47/vUXFQbXnFLRmL2oas0SJ9ozBM7Ytk4uq3T0aMp/3aLXws2RpXUfKid77RBYTCS
Co7DlLUtOvDW2G9xIXBJN293sYaIQtvB8z0ZS6eiIYI+Nle7IWZE7n1Q/FxN+tFsQ9+eoid32YWG
vsXJTWqL/apvnsf/p5BrT4PsQikygLt2wMYSpx8QtJWswIvJwe/2CcydBpze7eTayI+uJf/JMYNw
vx9YJV+q5A9hLHwsDuTwkyYL1vc9/iKxywUlRlgQ4wduwx82iiJ2KVr/Fh5CHl7he3N4M1kI2X7q
0AoAOpCIAIyaO8/wk6EHuM9LmbmmAJhejT+2x0Sy+K0UyL9tQMSdbjpWBjeLOICMIEHo23Rxrvj9
+8ETuMyt76gUyA1UHJfICLriNDrXYru/BwWPKh/yuK5uBzVOLYLXndMuUk5tpPLByyrEx+BdbDH7
PwoX/+rZHA/NZXAeAgaE8GsKIP4p8RwaORQpzdKjJwFwr7OLGm+TCgG416pgo6r8qJaxZAY27FyT
2SGVs34edqxxtskwjIxdoewIFgtDGWBQ1wkHvmIg5BgVkqQUiK4nOjGEXEihB1zG0aryD3HJk5n5
vXE0shH5LADj+3zRyuu5gsnU3R3MCI3pj/0sDyDUBGVevWcXSngAoihQbnfGjOuEySU6AKhlHHki
qN7kXRXww4hcZvqxBZ3T8BJ6RsOwxc0hvb/L8XQe19NReF0byVpojBWY5MaBIow9gAo9HIwYdOxm
+VHq38rHj3yV+PM4Kpu+k81InrKINQdsZZAYxjDbgmCw6O5NU3g7Xgk+d88TbRqUOs8uM+m5pT9B
QgiSNSIEIURm7WMtpsSSpqO4CV8zE1Npz5RSkDsrMnihWvUS7Xd6nH5A0Sc8tRZtkSMHPMOrD+xl
vl2GvXV5QvR+1iK2IYuMx3zEmi7VZVds0XRGgAP8Ji+xtATgoQkEYBXUzAvxyXYn9ViE1c7ZmHrQ
sISoLRsD3baUXXh+5hasXc+p4YEKB8+wfLPRa4suKQN4HrjwHzmErqK12MvN1+SSzb+/hi0afeGa
Ev6WGhWxzgmjl25PFPVKEnTIwOxUiGnFdYoN3WcvfbRlTMuPN/zP2+/VzhmqPjnomLIVY3cHgeZL
cSO0TTEFPwwAKXR/KydELD1NQgdgbMJNwo+PzdmDRLaObfDv/zP7obvRSZatyC9P6+D6UEp8upWk
d8WJ1wUAb5oUSxmDmrXCJf6pQPuwok9jVqd+9MPHaLYMvLlOqu3g89MmS2uLY3Sqk5MtPq90b2HM
dBjg129BPKW8ltmtC0bj19842TsysBOXXhPSQ6IrREq65peLDL0vuKVljVqXZg+sP96LF5AghvKB
exdD8W/vPxFhb0gfLdDtKAtepWzK3rdZTVrWAyoKVP+NK+tSOBPPV2FYlSVk5kPNZDWMkfqZSUFM
T0+S1Lc2kfUBFa8MwU8sPYlce4GGveyUxEAGKsyCD7lOlX6BjbYPb/nCKTBxtmnElI/jLqFtiCLE
qmDhS5EQgKyVcl4+gM4rNq+wu9JkM4XIOmv2rE7WVpuS4eZyVSlEtUCmiTnBBx3iC6RZWTYFWFPP
xr1V+OcbKHIL/iTtdSwEr82PyEHvplKzjnFupFm0/yIc5RwMmePIkV70+41S5woFSAsePSJAd/3k
hGXod+TTCArPfrgI2VHVTsKvBsQ9xb0qz3Jg1XsPSApyPcWS6rfQLdU2+XMniRrzRTscdZpc9qEu
fbBnPPRvDXhnoh0xH2l+CuxGK0p5ZnylUQw4GFF3eDoyCbEYIFHAsOlytj7+Ac1utgznVVnN+AIK
MHhHRpTtOp1VnEaw4CvmcASylBsH5tDXe8KWfNccX16DlTEL0Phmrvifq5huMoCJ34KuDUUpoGS7
fcuJ9kQkhlM8LMslZbg5pWj9x2ujxiGBEsVS2lZibw8krOaRIgyGGeH3ggbZw95jDnrUN1GBEAFa
HEE6txQKYWFSGb8ex2Oas/SbAwR3tyVc429AGEytjC+Jv5/AEwv/USTspb+FS30R0GuECP6p135y
mHwwVC5fIz1t0LoBQ5ZTimSIb3T8pnz/5wmNsIAAEZxfPVTIEj45yrw+igGrnqp8OLHeiU81K+Kg
ziBmW+/fYq8EcQfQ4/SKHF7FVQPXQ7vW7gs87CEjHsIxHSWFK5LT+1H4K2rK+OKubNwmjYT3ifkP
BYydkk9N3/BgyloNw+9lqcIKL9zrlJSP3NQdVAf80yesTLn/1bKIrWb5ah1mhkb83PMju76oCQwe
z7AkM5pDs78y13cT/oVb0mZEvqTsGqm6BcA67iTUUuOs81IJt8+un1Zz3Y3igNldPU2v6lNThNW3
jXXpJemVduHm6FCjGXM4eexmgiB4Dera7KeF7jcB2werZtWf6VoetUlIjxoJznHPm+QApkbZ1CNy
y8iCIWKVUnzk4KY7lFs+5UwMvDpXekH0vOBiMwqqvGpTMCQoNrj+Drz6HVf24WOHcZ2Xan+RK38q
VK2PPclzYwMm2IvrQKaXxzP3imKjtI34mgilZP1wrpaDlWmG9p+vSLJ2PMp76BlRCPCMwKEvomjj
h9XMhVFEjUDy/cfyRj+wEUKL+NfhR+yMLXrHVDCj/zflrg6DXLpWZiqhRUGmQSTE4nWXQMaOuJiu
LJcytyqnQzrrCxdQg6tOTarsvZeTCCwKy2R8pv+frRG6gUPQL8iI1Ln3I9hfMeTXBdGA2KuL0Gtu
NgRJAtGWj6FNkO8ei/zDHfR2N+IU1ois6q85mz8OXWcf4DHjIXbcgyBHbKLDxdL22nvk9YhoWTOU
2WIg8H698KX2gzqjDaGkvdsaMD+WEPwa/I1BhEuli4haPpJ5UXW/WELJkv+2+TW8JOR+Cto7hIOj
8UGfBc9ATcRqgjDfxbP+6ZLv65FxTIyBSOoTFaKCUCTcTBtdNaCidZ8W10FAon1ckdsC2MMMSrXo
7a/wSDR42nj+YQyQFqHBDLJTSti6UbEgDlcLG3DJYKfr8gAjO8l+RX33KZM3WWgahzYezUxDOToG
TBOVpmHZHZZW5dhjSTcGAC1FBqh8SEOkxtSyJRKBJ/5a/Nee2OIvV677sYJRs7IZhQWBGerUZ/Gg
9DIPiUKYnl4ftyR6/2P6eUr2aBUCTFOn85f4q6xF2FZSRIJtzdhGiaPPPSQHn2kht7EcD6vHiq3i
hucr0T95h4rOSkyhmN6nF2YPljBbn4KP48ksHwFn8ahCRpNog+8z+fdtfXOpkYFrXot+lzKBsJ8x
7viL3nQulJGYrbOTgpb9MmqaI+TS12xy5+KPDYWBQzCcTiNuLts/0+S46i2VxabWQtM2d0jMer87
Doxa1ChucUV58l5gymJx/f5aBCF2OjpZgazgGnYkXIcMsMJWYZnhNxCohC/xpUvGHMdKeZc+PXan
5OlUM25yjNQ9DIrPoUPzUFWkeX9ojJYwswxalLZUis1vLKSLyi/mI5bCuB2ePqoxLQSvC9ljRhVV
CtKY/HpocPXuFSvymFVyX4OlHw/e4565/CcIe6HdBpjgOVcaXzNHbXWBSRPxUsZRlmxQDDn9EBxe
XdbtDcWFEjFV1pt3Ht7DfmlHZfSLUfJOBCRuHSDiObdZFQ5I1vbPeOZ9VI6K74w3rXzc4NqTmFpm
TvX4rPC17xgGe9KQQMvrd7Zj4ZIXqs/0qTMbcG41ZCmN2+ye/AEfcsGFYms5aqYGnKDzrlmCdEnw
BZYUTiMU3r6AaCJhDr/p9DTQ7XqFAI1tFLkWwMC4tDVdd1I07EpON0Cb5wdMgrQ4wGCl2RdkhBYi
Us7Q9NWhDoDFQdV8NAvr+942EegG2txjWWQ79SitpDfiDJO3V3/uigxw8pFkOkFvP1e4gOUiO6Y7
qQkY6x30hMMxLkdKS7Ehme2zL+E1wBG/WHATN66dOTpSDD+zlPguVeC3yjEyKC5aFAQUsB5aC8u7
M1CV9VIbMZRxxBn09AM3qNK7/LSaCH6osGQlEbsH+G7FvZnA1moAalY/C0oc8MRPHZEQ5oDAfEBs
UlqwofwingxeWcqw4rDgcHuketM6Y3PgBSV6pbFhDvMMfkfC0CJ5O/001zRDzrLm3qujycKHnTPO
ytiyHEcTmLpwJioOIzHML4WKKHmRG4vcOrT3jbhFj1cPxzIYwxVH6VwwW5g0LL5yXV3N12fp3iZi
VAhb3fZ/m2sq/KDrHR/HpfUlLRjArshZBgQnLTY7syh0l8p2GsgKEnw2MoOrp/wZ0jgH+MyOGNA6
tEHuh0ObEeYY5aAVOAFOxG9lEW6OgINQrHhRA4LITFSRafhxTo798XhXSgGIe4DqawvuEJmBB0sy
ncUkXOH9y7+piV4h4Fuc8shVo4CoVLWJGIiNBVSufi2wBDph9vfv2t8pwpL9a2wnAsR6YE44Vqtj
TLKyJV5UOOaus4ESzKaWVaT7IlmMYZrLQqqRopn/mG/RykkMYdzES7EIkvc4lrlPCweqBVZJrvoB
B/GehGkqGfh6dMxsR1rLZk+61eg9pSNyV/Z/awbs1w4QXo5hiTpSwRQe7i2K261gMMLNy1nGDhNx
rlIZ5WrWstp7O9IrYJNILHbYr0PC8GZ/KR8qamj/Ms/tXav5OcpvpG9AWZnetuPEME22QIgJXb+4
6cSZFxyeRzGkMJOU+yqUhQjMpvfC553hEaTq+Ysf41OA2feJkwQyqNn58zMCDe/SbOVaNW8G5fx2
o4CiNvobq8DDrtxHJoVu/1VQcCqf76crH4f6CapBvgOe4DCC8esMZWYnpx7x/H6SAfNEfDA78tqc
IZ7TOpLKnsgQtQqSR6/uSscgMiRiBXKLYGZfhlSg9KABSVkHwx/ja8mZ2DuhPe4dlpXmmoLLNMyI
zJT0suBB+eY7H54l6rN5mn9iFH9+LedJEHQrpiIRhv5wmmt2WlAQHpyIUysD5isKApoURHwadBY1
WJ1ReFOepKrRT5HjMe5KfASnw6N2cXNWwHz0XBpckKdup6hYf5WPpj2OHtkGWrCkD/UcWOK6IYQD
rw5FZCz61r6XwKr0cc+yVtI26nqIMiaWVy8w+s0gPI9g4vVKiPLV+7kNjH5rnBNOFavJL14wsZxc
qjVHapsGTiLT3j7EE44f/SW1nJidboFs0ixJHYPBS7Ta59mxoeO8FowOJ2HZDuCkoq91W9CMwLQG
fgwZnWm9rNefj+uFp1d3jbmunrwdNhyeKhh6cxrjUvW0i12ekcNgxOyaPjGQ2kglWWKfO/l80wMb
2Y53ZgVCXWJ3laHzzkElYItkgw9CG2eEco59k8l2S92XxWzUDlB54lWTNjMMAfwheDd2qpCIbB99
DYzvrXNqBHpvcoU+mOzAWlCxQCcD0txZ19Q6KSkLl/f86+0/Z3o5+RI4PtHWZlb9EpehM17FFwRk
akcEO7GbHv9/QFFpYaY8kdcEw2uHf4rwsBv1IkK16AI+ryys7IwMJc0D3KO/5TgVI2uZxkECoL3C
45ecgTQZ6O9xYdDY63bB25hb2nz+zpDUmCQIx77BvXphp9CTEYkb3t8OolrAs1twHACTiGxwnnlj
SRkmdKOPJuZabbobU+F94vGXuEL04uR0Vhd/xi9iUpGrqh4kiuWfuhhfotsMtNAtlpYnYD5qIUYM
/7eWPw20DowOakFiQpjXAoj7iu3wbytX26MZRH+UBs0yPzPX6CFa+t0LMYsVNgmfHfuGspg448P7
wdb0QMWeKrn+vX7COyLzqMVONGRGIZWXvcfd7sAyUoSySCQIKRNH9paZ2Yyo08u63OdmM8c1Q54L
mlmB/qpl2IXO4wR9pmkfwgNleK2pFx2CBq7r+KDejD4uEM0p2gLPHR4oILTdj2TgO+n035L5FIyj
y4CUOofbmUhjrl9/DAQ0bVVYJoWKvt5lVy9bZvRzz8uj8czZEAVALeU3sjyASRglpcclqcj/lAk3
ERxBxIMtiyoujv7TxCoPLmQdHBF15p1lkjwz+83H+MH7OR8umTmIEp2uNeen2kkZjiZr0THpll0F
lBSoKaXIqDJBrQ8mgkVqCGzwqgfBPzV0HJHO+vHU/FqhDJRXNayTnS7uukxN1ff1B14zJZ3SrYu5
bWKPsFsXNJ4Oh+l2Us0bLHsO2r3JZJvduX1VPq6IKB+vjogtsx1UODZx+guhOWUczYrRo8zHC35R
lGUMb2FgJ3Hx5pn5bzoOqU0Yxt57HpxeOLVImLSQrFahBQPuepfkkmsXvZhgcfbCd+SnY2qXEMjs
KqUA324W/tXgskMwJBMH/7wPcD6iX7lXwj+K/JqdRNhTHQgHJwFWugNARrFI7s7TNgEgEvHw0XFH
JX+MZAKCz7dNoMMcv2KPUCl2Qsr214BmSeqgYFVebtuCGjKBgp0b0/zEOE3favWuyO6acmgiwFMp
2ywHEFXQxuWFqeLnSOq35ljLWdiT7LpXtZBHfIprcnDTElpjWFBBtq3Wm3U8xy/KDHVkfKkSRU5N
06pgvCARAryYf+uSCJaBW+OLqBM9vCdDCLEwvs+gDC8RYcWoOEvkv1uYA0N616CpfKrxjOqrTqcN
xQ3jue171x72Hw+jr5VwHdOK3su6MiqskzZBWlLhNq1EoQTwj/ef5zB1nm28XSbf1rUnfvcSmtq2
mf6HWx8IKs4IAMdEHK2EluNeFl8vysjWY2FOXlL0deD3f9fIeIa+GIvGnF4TFHXWwvtOEtd8fcL1
dXAKm8h+/zuxcAess0u3lnqAI54Rx+roCTyx1ZyLtBHaggagzNvikmvYOgheoyq5mnRWAIv7cG7j
bjmbV9pPrycZLyhNoNiO/8I8Q7lPt+mqFCdipD4dylLN5yfTEx7DNwP945MHXjHhYU3ZJtKPCFMc
ONfZVvxry3rUCEZpN1+KRVVlBjvySp6bYtlssl4P8ePym2TWoHW/eu8EXWqAi06RLd6d0z0x2RV0
6eT5arrlvgBVOIwZjXG0xRLQxXs3TV2cqPBlCKv2ACIi/4WVWYwbZK9AuptVAsQcyg3aMdh6hHYQ
RWwwgJ4Y8BEIB2OTUwpqsda73Sq44ML4H1JTzL9OzS+3lfgCFoEsd1gLn2S+x06Y8KgJpIZ6O5e4
eUuArvILg/7w00xsC2bAEDOSLqbVqXJjC+BziTpfSOTqSZVdUujejpn4QCRuogJmRl7WLcfe4Ov+
+NWHcq5brGDyquhCzfLkd5MMhnlLiMR/0JCzFOJEV6rEHH9WxyWF3rDti+TXgaH6afJBMVo1LSR2
jzKjiNyZ4JOblJMP6UzGblUjgxobE3/Sn3g+qlIsPCOcApUSN58AwvXiIL5PRbZNDPsK2pUXdS56
eWRs51+e16AULLt+eSzAIGkH6GbTH6qQSn6N3CbyQxTk+GyoCtVEEH365EX1anss7dzGeXqyDPUl
6iJPeg5VGT6ZGyFNBsdRp2XiwT22xAPXQAySnr+X2c7pVoPsgPrEtW+C3Av87AEKFtc8GMHUH7/X
FAcMqmfOi0kfHbshLXaWTkWOi/EvmEudRkC/GMlVnXT3ZdgCYka8ENYhjuunRXvgJYi5WSXlGvwh
FAYqZsBmJ2oJNuFpjPC81glhtjCfnNn9E8TjF+ZCb3l4xyqKmRzYa6k4be3g6HPFVoamHyTNpbgp
9uKNeL1k+wuhYSIueZMTEI1y9/pb/1/WfaIctS9XwRQd96Ph7fJpLXF+BhpfWqUcDvBEdZpN4Kv8
Ne82S1b3W0tzB+WzG5t1/wvbgTIN2LajmK1G4HFLysMx/wYkaH8LecMol0UEiQR/KpKDpDlwDU21
TYnzgXYk60LuF+QoVSbYEP2i3Sc7U/22TUxxDKmLhD1/6B87YecKSewMwo+POVBqka+PNfOAL/dg
ULRKgdjjRMtT8VWX2ncqNYYNGHiCsXBHHSob/l3/hGqMF6QdRjMAcJtcXyPaEEzL2h0I4JefaqfN
oeKw22qTpRvsPxpp993rfx5VdJ185R2i2Ace6o0aCdp7bbfEkprVZYdKS4THAaON2X7+pxpp1gSD
8cRspLH+UPa7+MCZkEU2zUwgw6eXOsGl/ZkdSypVkSZ8du3vCHx2okehCjVehE46UosMuqTb6vaq
FU262HZpMGcHepD569ze/dPTJYmBZpMsvXmhTHvMR3jyZv3tu4SsDdoe9fIjCNR6zYBgK1t2HYuJ
KqtRMIL2uW1xsAcfNJZT+KZAftrGuWqKMyfV8VXckrWFQuWpD9OZxRzTOtXaSc/RwvtN9UTGi7YH
yLRGv6tU98UjUn+ts1bPgwojFVR/8n1uUeIjiaSS42P0Fq0IgxV0nAycy7hQ2WqrQQvB2LI/ZcZe
a2IMXuzcalckdKkoQzOXwW0Nui2rirFEAfxv877hXQ+cZ8sHP78JmyzMlTGe6byrYDjeYStL7DMh
jP0bi1yubGwjjF1ApPayFChr1TWTzc1kCkvgtUb4xmMZluZ0hO8PQJ7vf6isaZ2E6RLuRQ8lozFd
HBuN1vNFHHujjudEnws4nYu/MErTrTkKvdG52L5z0qSCTLWSMwWD2l/LU/Qf7tQl68o5CM9Q1p2E
LM3Bn3XGQxXVNWgnVoLN+os2jgfR3OKZjUCqe9aQVqqNQAZN7hAuFcXdSmX1yv3oxsnMj0MUK29+
0MbO7xs55rqDbKBNSNGxLxB9J21EVTr9jnTqnO1Su78fmNXMQFpI+X0JT/RhXMRDn3J08vyeqjce
VsXNuocgdBOEdqlfmIbidAoc/0QINeRKSHfiyOexObdkFeWPlLLZo2jetwUogZ+2b+j7FH8IBV/x
UFDYSGKZAwa7QgTtDsDBoEPF6yIx479QqvpvGYas3ixazAas80RKjbD4iIq/ASmQKiarxxuwt78u
scWttdezXrrY0SkqfmTCjQrh05bHGs4E5jlC9D8CUB8TOArh168L/7ClNak7h5lwOyryQuBTsEwd
+BdZZRv47TljZiixfEtGunwctOl4OU37R9phgXLdpreBYcsvQcOcLcfifA6NbgJzhaCfgoYwExs6
L1LH9LhY/3FvoYEGnYFJnUQz4UMfZU00Kc3Bh0uK6rLZH+gTstxBK/udnX+tg8LB3qGopPYJvjZ1
f+b7tUDSvtMhTHhdKLG3/wsS67N1cZ9FW3XquxaQU4N5rX/e77Gnomh+WkYUXNCjeVssVZNEsQPW
IWY1S0xvXFrwzlme0TST60nXjogf4aU0+YasQtgF3AKNwsyDkWU/lmoS7GM8z8SBOSs8/+Zo9iAa
zLbBePmV1qLUEWGkLnDxPi2752w7hvdNVxEENBiwrooboTOLu4yd5S9lfc0T67E8FCzIO3i8ZCH9
qcq0aeR9C+CkdFy8fNhoiD2iL9VMERhM5ytLHT/EQ12ttAE39+4AlXdOHjjNPr5dzwc7S+WBVzOt
cNgKziNWuLK2jJ2bbWPl8rRZ4YCjZFJqmBEcMNJk+871eSm13Nnfs5IzJmlp5eCUj5Lm6X6tS0jr
hUpfwLkV82UGAgVmoJiF8Dt5Tujx4cVWfTmwTDyKzZ/MCaBg54xy7IfVBFXKVsuPDUJakkuyapga
0f8MR4I9aiQHdAzZ3BdYEh7ol8B2tiRC9z5hLGH49FM6be0GF+YJNRWucXdDVU0p3acoIv7TzFrN
Z+efTR3XSLlzDDKfwlCaLeWmG4ZHFe6LpaWOKOnVlGgM3jAIT8wUSwtPwLAxkzy+2FHUAX/wY8kj
3oWKPHBGSWWtabduVxFA17+MNKgDm+yG2Y+82YP/tWoIxUUksx6b2521ldo33mum2iF0LbbSbRCk
MsvH5CWvsiP+iQfGR+eez0VXtRjk+3ItAHNF8fRR5xk0z4SAcN1nZ1DO5G+sOburR7m23JOiTUhX
ua+4SyCu8ovU/jmpO5DfxxGColRigdf0zILBk60rAxt/EoAEiExIysONGtPLIvKMrtLaB1ZpbgL0
8X1tqM33VqMtUL70DBbx7BWXTKZZFVHevjxQ/0869HSTyY1AFfnTLjCDDGONPUWy/uYac5KSh2VI
/PzV3/7OP1yjav9+jvHX0YnzFNCmWAKhBg/++QlTGSK381MH3lZYmTqA8pHD3iGqM+j82ox1s2AK
efQeQWb5V03F6BpaMGNcnUVVYZdtPSCZltzoAfYksrRwGc7PNiGYi7UU5lof5pkLCe/E17ttHoCM
j/VLsE9amNPIv+yYO6yqf60tVQ4l0VA5vFlxdqyK93Bra6QfAZBgg4yXKlDBHw+iEgNLFlX/idX5
Z9sI2SX0bJZ9/qcZoX+T5wXWumishL8KLP/CNfOzkaidpvOA9q0x09n1xNive/D/11myWM29UDiY
0j2ECUOBbBBsyRU8GCwRy34Xc5d2DLC3dk2BHvh6N+k2kcLXec4EhcNTVLBn3yRJS6sKD6uA93f9
C96QanJGXs+ZbRGUQeDP9ssw9xyrENHQVE/uhNPi8UhdFmKUIh5v6HrGM/tM9l7tmlcarbu25L2f
nEXzPU+TA8J3uX7u5ZzyP6YQUrErSZCCtZ5Yl6EAezmO7Papsch/fuHc0S9dPwCaLuEPN0MnQcxm
SX08fx/vOM9LX3KyIGNpYlb8ysCXolJZtCskmQpRhVW6LjKGXGXOhdEbXfHCyRYpyfIm62XAXDgr
a0yR2E2WgL6SydbKfzqbRrnutolRtD9LbU7iPVCt/DqnKpIEjvBZ+O88UwmRdbaBVs3BSrMdveKX
8C7hdSmzI8hy8bVE5QSl9xv/HgDeA5b5WO8Sv7th/qMq8Rb7ooOh40I0KPAqR1WqYAl/fzbgWohe
68MOHFLql7iw95qQcplckc1lSnMZQQt+VvIR486LaTJwogyzRq6xK2OkB3v0SCWw+2TGUcgC8B39
AyOuyDALBMRP0tcDNum4crm36nIZeMYM1V8cZ7sgBVoTa1lIhztyI8xMTOalkoexbGCt7GZUW6Zm
IyQ1xNBAguB5EBCj8Dd7Yn4WJ0ipewNcmTD/ji149M9H2fwYqWAFEg+N/WiIBqUe5XCPJNulaAx2
goqBRpNIRyqfgiN6cQOOBuhuY1Y/vOOAj4BSvIR765UXjbDQo+8oce5eNU62fCGwH/Mw3W6Q3zAS
dC6PWTdkaxpP/pKFU/9WcfoJr1exxiTGg4nFzgppEOInu8X8vtOCe7/eQsn8+CKIaCQaUVKYYz1K
oZZ0wgr8VXkW4xnhRkx/jqUwuVoongoHsgUnnitFHMOhKNSVlKSX2P9BUQtU243y/41EApns8Puo
pAQs/dSjJ/488zK5/Hr2oL29dchMnXHn7XM7dGQLOjrGw+pgXyvrPAlLKHf9nuC8/DmFcfj8QSEm
nHe8cUN9+XEui9nHZEiBKdWDwqsXM+zhU2igM1E9It2c2KmLA2MppfE6nwwBCC/ug17/xMAVkNE0
3Y56ysLC4FCXaUueDhLKywnV+V/aBYvJsRQqJYxXfEpEoIMOdPnuO4CW6+dJwQiu5ADkW68ACwke
g3c9onbPasB5A5OV2hturVmbY5DQXj2ymKd/D0wS9PdL2ahmOYJ//OoaiQs/ByW+q3RaC4jC9WaR
QvDY1S3ZCxVrZe6s0R1Pr78Xj3gt9qFQL8lkoxz58NhHRGbQ3uaB9p17kUn0DqDjcFCXXyjIb3o7
T5NEcCr4dDWBC4b6JqZSMAEpCbEEXLJOcxShrUW4sMOT2gLAR06s0lZKGCE6D1bBEEgHdmF6xuFS
guVZo9GpzMBad5ldkZn0xqNgCsPi3BMzbyFV0Q3jWGvknfpcCsL6UJ/SztDRJMzxzQCzrbNWf/Ov
W6mVNyPyPj6pRRQig5bSMqPrJkiHg2/c6Qf+v/pM1hBXFqjt4p26ejc5LNixusLIksudBrqrHxBD
wXub7wKCtLVGOB/FSjeuH7pcezFlgOsELCGWLIvroZdJeAdSEN0ARaFPzFeNaj8HQrQueq7ZJ+j2
/Z+uNqehrq1aWX6ILx/JkZAC2OYnFqJJKAK2GaaSiMy241Dlh/TmbQq247i6AiAhdYHu4V6BWVeg
1rd4z1TSsPdXvi/gA3tpTrekAuyTGwQB8KsNZEHyt86TB6/ePvQSKQ498gIXMO4zHbhyW5DCi3MW
iW0nV5B5H3Tg5crOVxTXqOS7MLakdutCIAVA24GCCzfauo/2kcXbckDflkSuUpkEdIWfhvquDWon
kEbOLkaZx/f0sWDORYaHTA6LS+idZLj+rvQzeYaoKY8vzdo8Xw+oNPDJNjlTeyAfcMOlDEO5JIGB
Vh44O8XkaBSlmBRmTV4/DUermKI/EEUy7mCjnSSBG3bJrLVMg+5Xhm4nkJx6WdFIZNmbVs03ow8T
7kP1h+SCfRFPkSOfqIrMO445lPZzlvabN/btiNVMG9nO2IsAxUTTprIgkZHvYqFlOaQ/135NGQ6o
I40IuStkIBo0544sbsQ7DDLRnKxVTMGhATwANxkxllxTZU+bjFLwH0Mcjv0yV9bs6mUeYvS6/S2t
1CvUexdmfCCs1HXEFIi+kbkdYP4m3dZtq2QNf/DGCQmKMQH7K+zuIMzWB/ZmuKY4kSZTByycKuM7
WUmLJL/Iat0T9MnfiKD/mbJWEt6Rg6XkJtNbx80jgo90bTEap0HcSop3MiD03vixrMy/kxSsylgD
+DWJlqg1B7x5GRFZwUdwkhVfNCLzBx6o5LQ6czzZTvMKvLwSCRbPWsFDLCe5BGGG/7dwEXeOViqL
Jvmj9Ip21qhc0uRUhetEaPXGgdvZ5apB7IE/SIwzIFLj+KO8EBhkdbqDAhN7tvLJechERS3OFkJT
F0Xq1RbCH/YQsKOH6Qm4JtYMgYkWtdprtfZYUZfZ2bPI34fW5ymgE6/mHlo3y1KfFDxWPEwRSkm8
VYoSJUJKmFzBx7kvX3vmXK0uT8ycTDRrMjnlwDCHzl1dKbA4SEb4t70MK45Iy4R5hoC/njkB1DZg
dniXlxss+DSMEtSjlokSwcLV0BvU8iD1elP6S33p4I76IVLt6Dv1shojAhM7e2GkENTzVq/JXcJC
NtHZ63gvMrEObYsKCuNTXJF1ZT+U5z1BBNotZ7o9OYGzdSpFkH52mir5W18zijWAfCdgDbmzK0Mn
cUvzVwZ7BgHySIhkBc1XCS5vj3qpfzZQXVpH5v9uYIgzz8VhJfpmdTS8nZr1nhsY9AXaY9AhQteO
fHTi13PzM9q6ZZqRqrCHwpWqV1O170/ddae+FAVpgcL3PdJf1/iVxAqMHYI0VL82y25tFm0Axyed
NPtY9BnlIxMH1lyesnr5QjBaDyjolg5C9jXV7/cd4X5V9AijvWXEv+KmXvWlY7mPDmOwXqW3enLg
6e5bUaUTmx2bQpdbDqTkEoimbHq7TFNXW3AUMw33rAo9S6j84DvfZrEMCIlNrGWV7rYdr5KkcyjL
oLWq5Mcv8PNbVjQUwu/E4yztA//u362PQV7A0dRMf+TOd4mEpMkhlP8/gEueack72klKxoLWdsyi
vIIIHjOjDZyw7q7A6oPyTOROpPyeyAJLEAtRyOVZ6U04+kaoc+0RC6BqHDrUD8wS5vGgQCW9dHBA
qQk4cXOcmY1L+jsm4L2sBaup+rU64D7Bso3i3+Immvr+0i8Rg3PevnlugGR5+x/JnBj8dQ/zl5ra
t6CUiWzlcB8lfNTB2diJAeGu53jYVxxq465y2ECy/8tdwh3nr7MnmV8QzHORjS9j6t2yPDHze/Ig
ofBlrYsJdjUKaMPDQwSKVlbVHZEeRBFws61se7qbJBCVGirGz/aZD0A3gkUVF84y2rsAVM2XhbA0
AJurjg8rtjljIO+SBufsrT2w4XNofvgdVXBHTJ2XwbKIStDxXU/7T7ff/W/NOr0oIgv0qLNDJZDA
6jciaelZgkbU4B/DLKDbwNX/kmD56iryH9t3XGoVPptludxEhs4S6Oq49kt2vkBaQcCyVzfY0P25
aJ9xTmV/ZQU3P497QegQDpEOGYrqzhTZfDUtUpIU7JLyBRwtjgl6zeTB0LZoDy4dW9cSQnZDN6Cy
2ro5PI/6Mxz3RUVyXOlrEJ6m+iB6PpvOBX1/H2lhatywZMTxmxUmbVtd/viIXmDVsK74LMPdHghw
N/sUKBHRC/UlczyYnbDjspdoyaHu6Qkl55/TNySvzMIyrc6p4ouWHyj6bFM/u+f6g7HIoCvxLh0+
vaGQSz6uTjRmftVzp+1nyOscXvrmHuFcgyosJhpSJgCB2BvKHQTYM6nwW3zLjcnWXNem4cw5dHDC
q8VI1EbdiRsqFQZOaTQp4xQuvURm0HFVEUYtMAlG9gZ0/05v/lGrw2/GpvxOlXvdisrIHn5SP3EO
58xjxNJ5qOKcErzShfkUPMz/bHc1S3RYFaXsO2Ebu35aJN0vbLBRL/DynvFls2RBv+/sJprpT6Xy
LvZ+W+W7Pv9lR/dWf9kY2TeRFjd3eY0CcH1BjIDenz5JbEnwgPYSLF578vS0LC21iSFoLKoSXn4m
JHjCmi4RtF4uiJmv0numDN3Lz/am1lNEXd6VRHMIlOd8TgPkPFBGjkUjWxktsSypPNz8LrEPdpet
q6vfhnyVOCqF/wnPeH6Q3+9I+qyXpz6wQc/1nKtaDTjb2sEMiSz6hbI16PYcYH/lHxNte8IK8XU0
R6QqL5XRox8/dIUE2yuNN12IDQSRj4O87AtlaVp4Fg1hzEdLBK8BkOzMOOsQIVPmWF3dBY+7o4lI
Esyhn/DcFp+a2Le3MN2lSzRorWAXMGl/wHmHcKoreZWIwhRyRPQxvZGJ86G5YMH6gP7vhOErzVTt
B4IsxXGQ64PMI/EE8J+oYr0ZXt3quSu7xcLxrmy8g5od16jVMmycecSqWZv4HvLHUVPmD7Xa5TnU
UqqQo3oGcT0w6Rk4uP48n2MePbzjxI/y0pum7c2rnwzGCzr6H+uwYlY4G4E+zcX142eupJED/fD0
Oj3a651ow1Ab851m5n7gpHbmTsEVLTiLaNHnCRyrSDl1mzKkxv+ZVRfYppuJeSFej1VsrpwCOhe6
q0mepNiwS5Og1sFk0/uFHeXfmSOEmf6Tz1cBpB1NjT4XwmKBmPjaKfWTLADc26tikzxm5QbjGrw2
68MDKubPg8JIpf9LYcq48TXtxKmgUZCKsqq6uUpA0JHHgmtpHpt5vV1Mmrxo92rTA2AbrABnNbj3
zoOyzXe897Zv6O2Zq4PfyKt6TXPq5Amjw27M/3vE4KRmdJQCv0/YVP2QgOdgz0cMAqalQ84KlrJL
CUorzPvghNzReYVXJV4x9yh4WErOfB4CHxoXjBmlQtvbkRKCCtlXvtq349H3Tfylg9MpcKC96HeH
JqOyV9KjKkicFMoPFMoBhY6HVP9Cz5YwV3EraU/gIAIOdscdAfvf2bEREZuT/8pat0ReRfWoNfgl
iG6MosysbdcjoaiX19yquYAPDCBP7nMTWpLk0P50SlFJG2TMpKTS93IK+mQ6CnzzoDNVKHQMKtEu
zn+HIWUgCk0jf/rsVy4OTBUMe9ua0mgGHIP2qvw2aDsUFZZSgLMFz6bAoRJWS9PGg8t4CEFgCdnB
KuWtLwJd+mry/U+G8D0F+pUX5ntisJ7uSLnzxWnGwbtA91JZRCfUCAiZbEgOV5J8VD3W29wXVuuR
kHpUbXfyTDU4D8ceEaaYLuFI8lDHOSfn9WOsHK7cf91Nhf7Nx1Hvj1NeMgYAIeINNFU4u3H4tSDp
UR36t31sKZ+VsK/+mVWvc4uNN3lnWc1c8ZZt2ggJu8P1G2icPFYPNXW0nsX7/QNudghzXP/2NHNu
sBNwa+OYWN/hZBbzh2t/CDoHPhSmH3MgvUqtDSB+s2ekeXsxQns4NOaMrxkLIjg3NndAkQJHI6q+
7cj5rQgdCGqMUcYcMxr9terre99k6j1qLpDPxiHvcCOgKJpfJlqMyMvAcE/pBa9wJwyaqgEnG+kU
2qNNkLGL4lINCKmnCVD06YxWDpzxSwCjUz/dcSWb7mQUrJhsezyWeLIDPMPpU3ZiOjnbsDfYIS17
JCs+PSWTlRzXaB3bT8Dqdf9dEuiUo6J0Fi4JiMEsuWKuxvWFl7QkZmJPeJqKnaDD2mBYBaq7qtak
z8/oBRrhlWcmwe4QRRcO/FJJqvhxLFPF/GhmSDk1gEFnYXmSkPza4lKsPwvg0wSCaNmL4KaQMRiH
pD9jFBv7BgkQhDpQV3LlQNUWR93TFsR6J5S/YenHyjvwQoJlp053F/+Q9EK0plcLmY/RvI+tagDu
3Aeb+1hHfFGkyACMfmLmzuF2zO0/sM4OwM7kMpJ1QpH/aOnW4bnn7zj+wIJLuVAIlB7RI3KYULzn
nipjFbZ138zS0sA3b2ABeR8pfViws9hamm743cfpIOeRLqudqQQtu0pWUHyJkjEAlrp30hGC4LGI
wpobTG4aIijqgMXEX9I0J5wQRALTJaA2dioGUZeD3HfHhItnrjr/RZQbPhVQRufYcJ+t6CeLmBhM
P3ZMkMh9Rk84fXfTwFE5akvh5PEKxwJJcEyKTY3tB39RdURWJgmcngpYnHuX3HT39vtmy6gMa5Vv
AXWXiVDt7xBGUJFsBEbkhFToUvfUqVl2U+Dwt9mi1iCPCsEqa/+9Yj9LW43I05WlyvllUO8jx45/
u8ZMR7zFCrkSLz/uw0C+PTzKBfXoAAI8RBXFN5yoYQBoBhKGM5Kfp/Bi5n3RU8GSVxJVnIxdkaW6
yeZjZYEFJkcKoIjKlCgiu+H+1oady9JoJNbSpVWVspossX/42VmNm1MxtlqDlj8yCIUqFHulC4Fu
V6n8hPZ1BsdE9zkuR8flGhrbxovHKLDLznaggQna84VReu20g0ZNr/coqxqMfT682AFEsrv1ffuG
xZWmiBKgM+ttVkuapTP35OikFF5poC8CEsdkVd0Uvq4yw4HcqlxwKWG2RTdDU/oVW8/giD43+vP4
U5e1+RMSGLLCDIMnV6XamZ4VJIs8xdMAYXsitoCCk/3kQQtCWUFzydz2GZ+NmVr+yUDtSA2OHBNO
cpuqaKCJmj7u42pHxIWlP+aWH94/mU/YGkDEqRnSWZ0g/Y6+M14xx1meg7seIWFfHFkaWNYreuX1
Qho7LQnwwv6D3m5lueE8NLH2taIfhQeYY+oLG5fxc1R6ES2PZYiGWEZcwZRhlYkYDdJmaeYQrOun
D+N2vX3OaK/X3+l/dQoIQp5hct7N5iFZA5L116zq00DrZkHZyF8DYbghYy6euBEp00v+2ZNa0HCn
GukuXSQYgl3oJqavETy8hSaWfirvx6idNn1JLaiodC0ti8gCN6OX1JrL3dKeSFSLKq0QdCynWQAz
dqh34DGALghOfsGY3GLjUJYcUnwbINK8+gN0EFW1q1E/kU9/ewZVKO3m5BNkTRX7hAxpMJqs8UYD
adGAbO4Gz7U10/8QRsFJHaTKVlXP2VrvGlZAn4lAGbCIAhc806Z/EpMgeyh4/SkX01St9qx8l09X
QDj24sV25XetbQGm9MhIPWQjwUlE4Uxgzt+7DZv3VCbXdTYguAusQpab+bvO++skGOMgeUmwMTNK
AO1rqoQ4tyDMNVBpV14Zv3HocjdcFblYNn74byCBhBbdCQr9XHYz1tBVdFs/Cqn4+QYE6+XrmP/2
7bAJcVg9yge6V91GmQzOIMTZ2TIgcLZrkpYBVKQ3fwgtmRiBT8+sjTzU4yiHWaBQhhGYqBjz+tQx
G4wr44TC5AUuDTdBliQqzHaSHI4O/e4SQif7tHNBbSLreMFWJuO0ioGs8BjF5cDmfBRu3YX7C6wi
2Bz45HfnROF3JKepK/lfD/7VxtmiW9qIcvfBes8zLOHfZB/PCXLlbMbAir4LelcryqNL9g/DcNL1
F/hAj6sXdQpnjEelj0BVy5e8IAGmNfzI5t3Sum1Re1qdchz/DesJojxL9GDLw6o9x7AfeNTLxot7
PDK17z1qGs+GP8ncXEcF7ZYyzQ+VM/5FrEuc4NoD8TE5YvNXO0QLsNX/yweyhYdXxEYorcY6hWpn
J6FI/MIEbPl1BXwwN106vf4L12kgLr/AK3SYdKVfpLjQN+Z5mjw1CwhGWf5NJROnZPC2IpA/p1br
cPRgBIi7bMh13p4zzNozkxPNFSBaizVHTuN/e4JyaRCC083YZm9C8igX9UjN9K1WXqHavfshbo9j
Pmdkuck1SvuO1PASrq/kYgMaoaB3Ry/CwxTM8gNKoF1PJg6sPxJLVVZ3IN7VcqP/XKUOU3/vxUM+
gssSRmTCnpGN+IMbeTiHg2gjXSmqcGL7yRds9Q8ubz6ZoIJMNdLwZgLYcBAA5XBzFW0VZyqa4rwK
VVY5j0AqhR60PQmK+X38gmTWmkeehHfQg5MQ2ypvt8RCndpbauaPdqSbtWQOW8smIEODROSgFW3B
42xzIbLin9MkHCnIjkkPbtdw7TsZEtELXuO3KHPnUWTZN2qd61TD+MB5pDugbkWylxz8Sl74hyMw
t5zEalufo6pYj1yCoOHTG0+Hc36gp7x7hOEE+B67jjUu4nSRXPcCLLxlGVqGoT0L7TMlNi9oh59f
4KmTzyz4v1pWIleQvDcv44cxxm6LiEBB6/YCuMNxdgD4bR5J6iujO0rQ7ZbtB3hx19RKyiAj51Vj
8VxNrYTBXh53BMEb5MkR3xgI+qfpm9CoVAUd5hOZlsT6jSx6VX9cMxlmzsygt5Kbq48Dy/MqnIJI
wpSz0mD1Edbc7xlHN6CP84ei/ciGoKOkI05cxBdlyvXKkizSDweaq/GFDyrcuUn2tXSZXRWDcBVc
z1smvHXmRzBRBx5oPbH56Y+z1MUz1S3uMqCXLlKXLrn2p/TRs7YsPSNk81+rgPq98UmmzQ619IBu
wOLVPCh8sS49pB5vZ3wSZMNA4ichouLrXNOQMcrmUy6JViDTDJMEfOlNO4gqqdKmUg5u2XCcvntI
iZgu7cov3Z5ze9Pm7zmpWuk3S1WYvKxr7BexxTJH1WNj7wbTNU2zY5pswaiCQaVNjaSJDUEKmWXX
0RE+PgRpxy/i5hWXmSqhgiDcvluvOAwpbp3npJWmONXXoW5sDi7fNKwfrwj/RjaIk1disAVzvGHf
4OgEoB2arhEEbvl8UaWog/d8CfGy0icLNA5jbZ/nozDFmveoTZz8xFixOzsgaks4y3sgqhKAB4uE
+cUft7FeJ/wY0EOubSoWD6uNFLaTb6LwMZNW2uzIWUf/Hd2w8OzeGfeC/9FCEHs9Bf9AtIYnhgo2
ZT6KyaOBb7BG5JBBmrr2YaRSp/t9zORH+DPo2PAxip52f20BPOabBhjaCloCC0tk12WYtB4LKk6b
F7D5P08o5WXtK+q8A6sizk4InAWRcRxwKInzs77WY9bOo3BPkPXcXrytEz+AqMjGNEB2zuQn5byc
A3h7eYqaJgDNuUNzwbaYw8BdqwjT3Jcy0gPtyjTQ9ylSbzk80j1T3avfllPz5MppNUf6VhKA+6Mx
OwWV9ElThkw8ycQXzoqcwgF7P9nwK7VRaLIch4VCy28HtOJUuXRm7HahXIoKGBQFK+hqLhDJmp91
neMvziJM6dnHcDnHAagCHzVrM8/9o02th/sX1lfAb3sdg4J4wB7v+SJA5TrVzMTXRNzKJNQNQbA7
LqFG5kYVl6Eip11BvbsTSl/X+M5xTSMAL+Kg9hAgd36nl2WxejRU96P0gZG5VlGRntlrmdimp/F3
NiHmISYTc4XRpAhJkd/SY8ZOkpByQYNJAUUx3R2OcFRWNdNHv3SvKk5tDQqr5X0ZpV1JVnHJXhso
RU2SgK/dyB5ChG5NJkaiQdFRjQOGDzle9o8tJ8WgkgZeqREm9HFMy7saQxPMtd7az24BRn6EQMaV
Cpcbw4vM4VXRB1kSnnB6X0ar2Cp9eE3y9Xm0T5lhoz/ZFBodYuFGaAR63DL1xNaft0DwIlmkIZxa
4dy413MenjmOFpPuCxg1+G+0Hak2CFPRUdlj1LBIoA/5bezrRSoOqhISDM5FdAgcUxaJfLcKbuZn
Vs+JUbV31r6Yzwm2hrG7j9yhAhKHwt5c4nCSUJwpCB57FX1J4VgAvIaceRF39vT5mb8nIhcepRWz
5IyPrwEzEJatc6mPesQBUEz3W8S5HpH/wRjS4lPWFoInMjdG2GE/S6287jf945q0Gxm9mD7bQsVR
Tb0UmJthv9imKqA/NPXvcZOrADMAFzmeoEmHaDkdH0WGlVf2p+Q+zXisCdyc13RRAfZPHEXEHbgE
fbzo1oSwxyXyiDmRgw+E0hg2rzEIBYU+yT2fomZiJQ/kzS37JmPKn7j5OVE/dkp8wLZDcKgslZHR
JeXX4p/cEfJYWLGcoGvFCBgLDV2dHP+5E7MHaIadae3kZfDmQnhAdMciSaxCloLmrknnaZZ0SVUH
k/B7GT5PYvwO/77ZlByjWK2T40DkkH8aoWT51XOQwzHROucfL+C1TIVPzE63F5lRH5MfAwpIkySa
r9FysFjAftMox0ocf1/dp3PHZK3SpDLY9+CDiIqaLa6x4fDykJGF0TfIEQjT4ghDpNxiCWJnpPf9
RSvbUddm8zwaQIcZddiYtqqi7vmUooFPCr8HdBLZftMG0yU/4ljpPWOH8lf1w7DkoFxMuE98oJkn
OVXfw/HaIMt9jjSHwc3MdkjzzVwT4T+oXlPqfLNvaH3WhooVy4OITbhcMmOUBzp1Cm0XJktVE9jR
xjWwqNJXlFu/lfJwBn5y7hYyFgVqJm0e/WYxhWkXA0/Luic96JXq/0rWfiFWGgjRTrDjTUHeeXim
aFKRDrVHlA0+ajTvIO+ska1t2U6hygoRKxtqvrpELQwpkg4lTLZAmouP9IHj9h54RcB0lj33zP0z
uanGnrnDB+nAU+5rwbNGw7ysUoYIlK13jv2w2a8j0KrPl4fncVzjHEgSg9SmVNDZZ1Zw8AQ4svcs
6P5vDaiDVDsumzI79c1W1Uh/sjPJEcARTYs6it9oA/uuXIDL+OMVfaoumJK4CS2BWbIxHoKeFHGF
WGvvvGVSGlaHkZQOXu348lI2KsjUPqwOGbtDbybGMdrVc8l2BpzzCc/T7rnvhTvm2ZdGYuLgUksR
SbcdmWBgSTuCKhjWBeXLSS1rofQ0WfQwCERcDJstkbPnTNc+mUT6iZpHxEZ54BtnPdZUFH8A6eUN
huJHTSWIsfDqPC8vHvoXv5Zvqs+Sfw2LgshP9Cz/h/XANBZoKQrbotHt59xe+yPDSx1CDIfC0NEu
Ze3s+9p9+b1QZu/UZctEXpds6v60hHnDePsJpKq+R+n2c/Ca+YvT2F5BI02VATE60CTgsLRGhczm
gtMW/kqKxx8ZqIKMNM+Nys1xol10STaC8d/Oo6U/Mj1A/wcqs+LTfbkNdb/ch0wsGSCLKZcGoX2a
qFzc/ld7irlkEghmJiJww4a/+s2g4JXpG57bXKlDjNbpSse2+Non2k3NzuaV16pC1ur7GSR+Zbtg
WJFk7mmPRhTqc5Ovj06OIT2QYHPoOmjEPAABhVuvObrp+YhGGR98BRZju5QbQ2uXzey9d4sTg8tC
R3gG4u0lBC3Zm5qrm1WkxROUtH/T9TXORWE94rpcrH0+ev7uCbd69ThB95mvllomo9JcMUyy87r7
xeF7HatdJaX+Q6LEn23NGgpZsbZN54s4SNVveZ6Uq4cGsc2sl6uE0dK2a4pbT9AuICcnr34Ppeqa
3AMJLEeNIiHRqctkgg5CDOH3fo1lzFKjgSF2MNOFEj6v4cXXy+7OlAMijHgLeYzeLAfslKGeOczD
MVmDrov7shZSIglBeK2mMxM3hocnc5PlE9aAnDi0QATA4wNVC8Zzl6xCZ99bGAH8FcOKFshOh9yp
EsvAJHLiER1FD080bo1+xbT0Gs+hQqLBQp3h02EodjoX9sN/9EkvnKZE4alaEVFKiLBvHbRO0pQY
iSGaGXJZDh359bR0/trBE/HxyltOr3DPOZNxFAGMsBM/F6xJ28kmLJsH95N8D9+Z9WZFoWFVFfmg
C5FHrmMr1WAsqlyj91qkKju5euI4JVaGdwwc7G8yp5ocDEVistSSV2+NvBxwTP7KhnaZ0arR79/x
JPUhTRk2wBSFParRM6KYQUjr37jS712OODEmZvVhrC1iQcBRDQUbpEfsE57LcrDd4w5wDE8Hi7qk
NX/Z3aeDhgj2X1+Alf99fc4sRVraokYW7BYzNn0VE0UnAMN1qW3VTu9z7+0SESXxZvHXMLTY2/qo
Sri8qMJJVKLhMldlT6tCDRcej2MwxsWJ58C6zrDzArn7+cZSjG2pebK11ldMY1ZpAjDRAdXVvkJy
roc3iUSpI1rhYpXT+vXS6l9OKAmF3tcBRuFeaUcv0L09GNsEfnq53y0E9eZvZkzNW5X3UcICZziF
1PrNSA4fQlScdoZiOSj51SetKsh8sDQndM3l7TQpm/0vvkvaF6GN4VH8GYFbQ8222eJNZkMo9uis
4ILjcjOZvCTeayrxMR+uf59Z2Wplw/x2v+JJkWiag9F35DSV8nKzh7XxOh4NtqGkPbai2k67T6HL
vQenCaIyBifeYdwXOXXv/Ca38/z8j50BbQ8ZXdqHV4v1AiVtK3QHiP7cTZfqsKp5syZF648W+nBR
/X4UPptb1sriUasA0LmeFPZfydcltUrc9Uy6FiwboFaOaAuFWtS04ExlynvnETwDEMB0ddXV6FFO
Tf1MmISAg3d6MkX1/46S8Y3JMTtgCtjsRMXcnjDNEMyZY8b2TQAy0183oWH0AMWH/muq4GHSKLqB
viAU5GJwngZc3LWCR3+5C/18FzMzZt1KZ+cuojkK48j/S8KmSty5Dh8ct5aGLqGsMSY0UeGhNeDy
Kt1etagyCGbC/yQyO1pszObl2RTn/gKUYdZGJ8aetUWaKF1WIRqqg4C8Pjiep3gsGNabzrHgHQ9w
JxF2przdqD/QKzZWOgF/zl60fNVGapflDW6fYVP5IGKIJMcXAPB5m8WALJPyYHIf29sfgYamZ3D4
rEbxVoX8667sJbmBedb3wM5QLY26z1TIBLCIH6DFgtt5cDoHXU7mmzRx97/8CSbBxmx9LOKwZK2E
Phwj+4Emggzkk9XBCyIc7PayiIF0swmfANAwO1dI4/wvPH71t0BCYXlQU665QTenCEb47aMdZnVL
eev0CAnNQe+wDClR9WYyRiUhXmKQ7AowDmKXV+pMJshEIK2xGtWDyiEm07nwuFZESAe/mBS5EW8U
EHFRlyyE4onB5hhhN9d8KuKfNZzoF1FvzI+hXnyB/wtI2BFq8gOrVgx1wvqRa8F3dcF2guLoQd+d
KedBNVhc/NmcwYYZUaGWMvFWMzIAMAHDhpB9EKi4J1fgdmsFgfP25lT5XAWHloU25rZhL22EYM9d
HlXf0DxcwIy3LkaiK84Xnwe0JPxTEu+8kqWrEqtM6Wd0rOIXwAY7a8sui3g5gfI52PFs3DCN+byB
+KoeIsS31uA7yawUuKsAE6sPym65RYm2oxtkud1PaxBjoHR+kl2VuBo205uSHTmOpAchLbucBbNk
tchHNn+smpFF27jXK2WErmi7L7/CFcdsu1atMKR/zLOcR5KcY8muCxiPvXr7n7FQ6i3o2KqWX/y3
K7bNKaWZkuzvTuEWJse4wb+gFYJ1SC5lLWOwr8q6NX10YIp/5hXB7mmSrVcRhWRKbWiwmhyXNLpQ
czDBJJdRPGxzt98K+z2qa9A9P8APGRwQcYMOIc1078okKdKHBlrqEww3ahy+Zh8AOJZ0y4baD/dW
02MjFTONB8ZsmViASHc+jij9LDsOYEwu2vCko2WYx+mlppoujSHvCLYutrd8qgWcfaOSZLlqBLAc
RFVYqJ3CKjv38aXJl2MfSKurthZb64r83agfxuxv2NncmIZ+hDkEeqF82JXDN43b7JsWjGA2iYoa
SfRm5XSI+HZJ2Mizaybtmh9BX0GNglGlsAOqbCmNnIbAaRuO8LN1Dt98rjilFNIxn16WaXFIpTnC
x0e8LR483SSqaC4FDk271O8JCUIsrsw4B6Kks6Iz/xPL/ZckX+C/jyzyGi2jAwNi5ax9qsSYbNRH
PYDcZ03PEde0Ih3n6cXlpO9vMfmItAOoWZR/2GCa0mgGMvgs4DWv+dZGqIdN3UHIZoWxKnoN57XZ
F0QR2AcxSv08stkh1Zt/HKGD3TOhSpfgqsGFl4H2ni3OoN+qBKDR68NpBwN6L3iOzWFbj37UV2gG
Zy3pRUerObBQ+o1Lrs39ICeok4hbLxFchjYGDKGOkv3fnL4NcqlhI8wwZTy3+IusTn/qK8+UNNVx
Zs1UIx3g++IcwGodXgU6iyXJ0VNrv78eLz9rI9nYhxyLiNQgBx4M8kmrie3J9VXDrA0cj0JMtRrP
Pm6jwccVpMu4VI+BhoOdIpRv7ZajVQXPubk2A9vfuEgCjJdsNF/x0HP+iNAWnNnz0TZaTLlcX+hu
V4lFE5Qz9npW0te5VSvvnWIsCX/8GEKU1+/RtB2/KtbgrvX/XDMePxd1yGE+MeaIUm3AEXwA0NZP
sz24KLT8T6clvZYR6v3aFl5twwJ1Yc0WSSkr2woylHg1/FGbETyauLp0mO5pcbTsDGxnkuW4nYi7
Iub1uImsXMVUI8S6OkRItVj1Owx1aFqZJ70VM0lB8N24yW7EA7tfU8DF026tubSFvDayOBxUIfaU
aPEavOKmTKT5wGLruLFpLXRVzBF8XxvKQoz/bbDslcUyf+hphHCCLi4eTO7uqJwPZZ+tWj2hNltx
bQSJ8gRaqzVLBK/NWBXxxDGTPokdliHjADkKHqZPN1w5f0Z5/sTjUeE0zt6RT1tLB1gVlnp/8oBY
qfbBs3eWSDffmYd0VnrWHSf6wt0gtYRN+1Ej55x7hbsgzduBWjCCcBdpXwFdithTqMvZ2SL0JVoc
5GuZMH/IkxeNxR1N9hZn4raDyzV7fmvTTzYxlSUB8aM1nhV3jW8WXJdiDUYXj/URC7k3wuj7w2q5
JJ09oBNzfOvd4WPAciuFeRw+YhRpBvgGOGvl6KWJKDBTgikxkKtd8amovWqO2ubwuj1ZmTvsHwng
GSwysriDWZgLbmKD3RBnAjE34piDXUZ7ViZ3SRNFM3kADilGjKsJX0oohv63Ro/SzOuFFEbS1JoQ
fZgrjKIGB3/WpYWj7p1zyzMKVolHXVFncalADsRb+3lARQLkGl8I5xdvuXLdA4exjS161YWUBAvq
ZFKxUnnofi+iqq/Z7446s0uoK3IJUFuT9fKD8nas10RBQhsK1LFGMpgh6ZbjXS4tqwIFaYkXB+6N
61XsmoHlK8VdNZ0aGjinH9y5TG1OeB6zjmCTPJbjXLn67dyXya97429MY3lPn8Xd5SMu81X0Cg4B
fJ+nsex/5JsG9RJU80TSbC9HV2AtYDwT6a3slGUvzzeKxQFfcRa+L2Q55mVgoM+tstbHq4W9943J
XggnwXgqd4HmqwJedqL7dc56gcXb5Rxd2DtFPb7neYPFIlpLzTvDviugBVm5R2THoMll8P/KG/6X
m4jrhDNuTJm0aAElY69i35gLyD4oFpAyAURJsO/g/DALELkJN83VcGEAxaYkbAw/AqGuZHl7SK7C
y20aJ1QrsKk+n+7YcNWEK3Z9LhsPGCQd4cb0J5VqHTZQ2MqQ0xAzVBEAxCML+vqLQubsByn5y74V
orpMJuWiXaLvFc+981XhvBmLsmYLjsiT15769PP9BVG+9lYhNb/cXjv6ZBS0ZOrrHs4YUvgVPqri
J0K+MQpyELEBfEGayAqGja+FMwnFDykS67eTgFXm2yUAbfT1W2Vi+z0Y2V9NigBJTlcNPN9/wqk8
bIonPihu1ZksssdE1OeIgOA9Ty8OxG/bI9+IuXf4ChvQ/gr0Fl6ERlvlnTrKzeHKqnLNb4OA3PNY
g98pWjCo8lveAm4REeZ/IiRv/pyQ+vuSNVZnWoGV71WVAVzPaQFfiGgPo9zea6U/HzXkCSVSuGkj
JXcWhlhQxD9xqysROdUAUokdGeLYzkPEvCMvIN6dxJHFPyO9i9u/Wdw+LFKsnAyxWBkaJsuAABKV
bnguguRPHDbQZD/hjdxyR7JKE4wnnPUfVhDvtquhxj0K7j6AL58TpnuKwKGsmTQulEBGp6DpouNG
iYzyx4POz94Ts3yhc7PqwjGk4149aHSq2dVwq0tM4oXmJxPfBt3h0LyUSmy+Y83IWSDIl6cI0f0a
LPIYPzOq2wroKbSMyz6eARVrpR7HzN44ptilhYEAbQhLabkKy47Eckdo/OlcRqlQLUx8UIah9SXS
0FlGd7dNRLQkV3CLOfoo4Tx6dDDuUpRFg9mqV0xHvjoELblmC1zNKFXQiVXzt9+PybRgupuy6wYX
P7z3SIMM6EXMKSBy+AATLWGfVLoekbIe5qBRRI/gMXSqhKazUPCutLlvJMVzjQAt1zNxuySCC/8N
R4pDT8VmhGZSbu7snjQupOXhLuHjsnTtG/u7KZ1yNXCF+Qve6Zk2icjp/KnaNr/NdfKRFIEbQaSh
ZCr6yklQTkkqYoPLPuNYKzUtpPhBjaeYCTphO5q7IkZtcB5cvBPtyNFUv1jYorQct74eK2MGo/Yi
tyCTM+OWbz/d9RsbYGifjqcvKARxaweJuatfbwxVsmuvzkNVKONOpUZMgxJT/O3BQhxfciS5MHvB
ELPDeZQkW63lscoA0TtiLexoNMOzombTcwyOHVFhJVbCMU5CmzkUsIbefzJ2UN+Q0h/65hd+Y2nD
6keCDF2Bjm5mBalqwIa+3Q6UrI9wUUKKTsPTseezu+SE/nz6MvtlQYgVefneKUYUHcwaLlJRedEI
WzSbr6eljiOTOimtYWIiv2JuyMBxspqdtObp0Geu4VbDC0Tbg/QLl+ZNXJ5eq/88LAcQ+y39oizS
1pDxDcdicWtstloeXt6iuq+XQR5r0+Aj4Z0PtIaItRLwVvTDuC9L7bj2ly8wKnVdyJRCQVjZYOXG
e/1Spt+SY62mvLMi2/2ncQUzhWQDXi+BBTHqz5GOK36I2IGPVjTj3quwMDmqw8C9seuAnYMZr0VM
NytGeOuzgsH6BKXBtUo8bT5Q8gvMkrP8owCv4wr/59THV/TF3nEYhxBwe+FfE1SuxlLkZ9aqultB
qu/PJo/cZsvkmclKlToZoEEQq16GzgGW4U+uYSOog8fyNlrjvQ+/g97RBjiO/fbocaRt46SD9VcO
oYhAipBIi20el3bbXSDB5ojFp3jkZhRG7FdMpmCPgFbQ0sjoBVr7pVvSIm4ENmCHF+UF+V6Gu1O1
aIwYLXII7rqZ8cWcURSEx+yPsZhTqNtRetC5WjsKotX+5lgePbHor8/0DZGl7D65Ys/M9LO+xKeX
3dARpcB+O3OcANh1GsvOVcAJFn9zp/XwN0Fuxsd/3a143cC+ITcsZnRS3m8VGETh4oTx1s/YqBuP
xvaNb4ATcck6xRpjVKwryDIGrNinvK5jdCmVQZ7MQH3D9RXCry3Z0YNIhLnkuKUIUhdsjzXg7uFh
M0Q2UW+f7EwBnfdToBK1lr/QU2+OsisEMp5VbFZqaynlJ2SDdAV1vIwTUXq3OwfkHEDsJKyFETZg
6jHJd0DkNIBmmKnZGMd0gDg2v7mlx/DYDRK8w54mp7Gene9VMy07mPUCMvr6p+Z472sItAJGIPPm
h94PD04Yy/QEBmcHmLjpHPQQF2yly1qrIyOvj3ToOOLSfXC5eTSaVXSyrgNyFr7ZEohO3CsGfaof
HH4dUEpXAbzJ0WlDM8w6v3YvXGe5ZXRsRwdQD6/lIaqKTgDTDGwDtNtYay1+4xBzCD1I/EiCVCUS
7V/G4XO+ueeTSgq/NajkXi1cGpuPyCluuOii9JLSzEdg1R0tgmIkrHdU9FOemVKPR/2jVqdEdaBc
9SKG6C6HJ474beabnB03l2shDsijez6yJrQ8i3Ku9HgJBoePJZF3NXd8UOea7EiD2SMFjar7zMDD
mbyGHk4WX5EQzwajgZQ/gKEDFnKS3AohTK3bh0ldb0gOimdt30SbKl5zdyoJYISm5+AY6QZLmWpV
XltJ2jnWV4NLAXf1fbo3qDVVGIb0c4EiZ/BBaZe+e+Vcqj1cY+i3d0ad6f7Wy98pF0ZCDQcTwzIU
XCseSzbI9S9L3r1F1xXCaUKE2jqsdC9lFzmKocDdtxlRV9NMamSV/MnnJ1P8V0sXhIG93zW2Ge9D
OpzbZJxlHFbA0mB5EWvl2C83Jqe7QrhqLMXDJajXOHyUgFg0u0KSv67TNhGVLTDms8lDkeqc2/PF
hcD7TvwqP35ZoOI9pAhAdCiJc9zlhMFrusY8ldtkFElkmBOEV6Eug2Ku/Kfin/0se4EQ8ktA8bc+
xasqeQNZgVaBow9EtCXRBpq8pGIRg0T1ubw1x3tWDyWBLfC2TryX/W3vtusCRytLEYcrh/rymUYz
9+dbgC+OXojAZCRjDsPInLdj2AX8f/k0I/TAn0z7zWNOjmwUHUJPDFkSxJ6vUv+AgM3xrumRKilp
TYW27ajIDjvJEp3cSr/nSoVVqEF2Dz+blHuetC9oq0L3jSCafZSBkZy6W8RZZZ8431GhcnUpCMsF
QjKUkmmAL+ib5zZZIfMfd19bPOrZG4AavjFfYtcd5LbWEJeYrj0GtqUpXXzDZ33ag2E3rloAQOWE
e58U7OeOarB4JYW4g37+Er3gKUmtTPp3pIAKH+ayfa9gPPbMpgkHIc+CEP3xrl7CtUm+ms6ep07x
uZwA6PV3uPdfJljo4MjfF2Dydpx2tILlYAeQkuUM85oN807FCDWX87oWy+9G9wBN34mGhqLGhw8T
RXK1VG7aciGk/ozQ9DwnLZfNZOJe0Kcbmf+BPQG6U+BpG0aB/ZkgsQBFdT1sn4DJCO02Ey88+jIx
FPUva44NtFZUZSjo4Y3uhW8ykneWoiHnEPwQO6anpFxYXy/0kCAengHXlyYf5w/1dVOStNuFYlab
hiaP3alaLhXm1DtKmQ747fk4sl+yvTNN97ZtwlYAX+ECiMI6MzjzUSUr6Ye3GDRGQ19ApWm0zCP4
Gwvcg1uILPNci8W96t5tv5KUr1T+KF3kMjnx5f8xJ45cdV8bycpHZBRYlAFShuRBMx6tMIpo9Zzn
ubShAI5vdb962m/BalOL1JQfjXjN6tNHhS7gw0RcQtDLH3YziJ0FBl4njAAfuL5JdLh7lCWKbIRv
SONG2OhrAbbX19M/m/P1O/wz4MjGd9fsZ2vy+508TE4uCARMJOUePEX78pkhPKa12DPWhLWIz+OA
9U/CC4flVDynTI3w3Vg4W18Jxbex86EyRuwLxhxKIwTXiH0VIdxUmnOAAITC3qMWtGfzSO7YzTYC
tgZMzkTxbcIvcPPE5nyaRbWZmnHKw1QZ6Y+8LqYGpwToETmuL9Ad/5tZEAlcurxpWJWnPV5r6JQl
pE+jB8NRCgiVKdnoyaGW1sQ6fQFecnlV1nOOmX458CRKAVDE2yVk5N508Djx1x65ZgBYhEp+lUUJ
VW/TI+ApjTLTKW9Xys/y2gV0YlzQpzQZL4nTLYlm5JDpuZATrhXR2cU4y4bRtldD21bRfSexRL6k
bkhhwQaX0IlAT5npBmwyOci5HGoPcmpvZPEx3KcNoItWqMUOBDBw5UTVDBWwYDTJ+DB9lN5BQ5rc
ykt8ZvR6WRC+EwvlVYp9ojI1/+5m6TzuoDQqAzgFzr6ihCt7xkxdkVPQWBb+RDS8Rr82ZS4qH0MF
EoU/ilXOGdeo+r5IxdzOK4wTPTNnBGp7D4uLFHRezkPZt8nD9fH3QHmZ5ZzvLnd600ewDTMMyiaK
32i0vEyOky0PNSv4wliNFSp9f97B0MGfpL4BsoGMqc6ZRffUU8Q4UxOeMNDj+XiF9puS24qkFItH
qRDE3a2+q+o3JczPJ0C7N9tm6p5u0dqqNFZUSVqAPNPknqKbnFqtVSMfsgsI89i3w3mHTB7XenMq
9Ln1kcpAH+SDX2d6VZADQzeE/Iar2WeCimumZT+VFMFqvNRypTjcEklIlwTPl0Q+7JO73eJYMt4g
yK5XQw7tiT7FwBVpNpG3v39bz0jTP/6822Fuf00TeJShmD8Pm1/QYWBaf0l+zErJUYkFSTT9gcGu
yHhzAyxoAyMdYVKmJRlDzsPqp3GlJR2DnViJ8aK3U0a8drOVEWqMmbniCVL+WnwHk8rAGLcPd8Gd
GfORLBtPdZ9fW1mFc2TL1I9yPhpad+ww3ZpcBMhf24p4b8dI8/DmFZtJAo+TiuJNU20vm9gOsv4c
J15ylmIBe+nbCwy51EcdDN3mJn+vF4YqIC42EdsS9XvDBg9NjHznT6cqg1Tsr3uwysMSgRnvrpdT
sAefcPpiFHvUE9uV+jKbA1pT4Un3ihiKy2kPtLXBoyFahp6oK3y/WYpaNtENR5NBJC+GngBNp+Rc
Q54VbzDTRHy/oTn8HYQ8aJCZzPy69j0YG1F90UsXZg5KWzfKSA7g/wjtyz4TEykw8SG9Q8gerzBx
6Rbp7EJywDuqZdp3HdCCROONHxzYr/eJCCOcifcZGH5+fQxk4oE2QJbWJXhSiUqoZ7ibouRW+1qw
v5SgClK6tK7CKx0HcF6EUtQxxWd0qdQYOlDY1sKh7/fZ56iUtv3vU6yPwEYIMMhik4zyuNjFUf/f
HkxRnDyMvuu+/O6hh9ucgZXk5FmETujgs4WyHbJGfFNvqgxsbuch5PF/qoP+sknnOikByQFX77fQ
yZv0WQhEak5n9B5FXnBXhCD8V7h3TC1MBbNXabuV+Zy0iy4KRaGkck6da9xzcszDnBPDd1nFWrGG
7fkISQ5nkGQd7BT/h47FTHiTypzDnXCdg5utDjiedrPoltwUBLydWDErXfhDPL08g244HV/FREJd
/4MtP9tE7M+1ZWTOsabsuilEp1wv8+lr8NTAgt1U7aEAgkzxJcKRBRKwY70O/fP8N3Hyu5tmvLU2
/1olYN0vXOhhadOdFqFHx4nKN18qxufEJtBsN+n9HwekiC9/66WuJONyabvgpJY8+quyRxcT5285
xpuqPp0mSqVGrV5iOdiKkw2OopUNidjwUwjzbcP7t9Nk8DMaJs7lGh+/uBHALJIEq2Vhz2slnAL8
aG8qNOdFDwyWS6QI27evJ+3MDS/ocbRI0DujmDCCI+N/WtPBNolUG+kPSFdueCEeQLSlX2kMYpQM
uICRn4cKen1GR60GHTHM9QUvAkwBYS15K2PAJkrZq57HKpSrn769caJlbemPdQ6mOZbJTHdxVFmS
kA1hkHkC3Gml1VxyiQxsPy36qj6yuTA6oLlUx53Opy9RRcU/gBC9cgo6p9RBVDK+4lAWuK0HPYrp
pi7ouGzllGYxyRjCFLi513/taQjdaGeAghoUsIezyFQpGfX68Kz3XNq/X7ODdS+xFBUPsqoiGK/B
lcxCosRP8I57OLAFk3pX0BY15ltXfKRKJ7mr6i4iXpAZK8OEeZiNPElKP2+iqWNT1PPhs2nfwSMs
MWH6rXNX3LQp6jhRUyrEUEhye4rBNVizXtebbyDmGL6h5s1bYMzeZv7DzSaJfbUSHL4oCCQMsqqr
CEVqxaN/ZhujowJxUCMnxRpn/sxx694QIG+72lmN8p/b/lKbYntE5jz67HU3g3KsmW6wdcOetoan
tQvsRoKeQG+CjByEbpgp0do0VLQYsaqCqCR37TfF63XlmuVKPVt2b/w9Kxy7MXeLLO8h5tgnFuxf
CpGOvsYuyMHwohbXrqUrwXnODLZ6EKIVs9m1vYBON65li5fXpeIrRcydIKcoc9NLt3LxSNaZVj0X
UcKN1biSuHVR0CQcJAZS2aME6WdCso6Hi6UBv+z6yH6mpTMAs+eLayZlu0siDpAxsISii7TpF2VC
OcgJ5HrB3uSKNEWAQTMdCoMCaHcynWV4pxAP8ZM+xW3X/ZfCwEDZyJDcBvQBMZDcKzkDQ2GV3leB
FhFVV+ydVuMexMdUsbYSWAn9pshx5bnA/7S3HPdq8zfqszpoA62z+cFraq1pJEIefO6q/YCwVNaQ
hR0p76hOyS+FADr4P0qKLLL3LR2p6IZn9hR1hM3MjrOpTLqL0AmgaOFF4OXhesM43IhUpRwL3oKM
L2sx/xhiyXjxPDeLn/rziLHn4rNaLXU1HNDllGhJ7kE/yLyJX/p1JxzjV8VZgOA/hjFsn3eUzpEd
aS04iEkbXVOYxoVQp7Ru9bRf8FTnbTj418gcxoTu3J1Mp0iv2aEqAT6Wbz7gJiuq5zKzteEuxdMI
4xS35xPhV0/aDOD4JKrFsTqiVDRH7JFO2JowHZaAt5lBzjUC0ASTo81JO09IdZAukNKfoJM8C8oe
FKejmfywgf/i96v/BP9k7ne+uP922rcsFiyZnvNGQc4oTdixtU5w5pYnO26G46nHBFm2mnQYucN8
L9vsU3CuwL6F9c46nDU67NueG4mfaVK0U8n5cWVF+QtPwaYTI/jxjTK92vzDdhO75POGYxU6LDN6
kTPmKkiqqY6ouXokcIvswfyaaNuDjofNRxmveWlnt6VfV7gVfyWGQYMLlUUuIpCi+Aa0klXkEZiI
J99pRcN6wn65TyOg/WAlBtw6U6+ftMWTdW3gk/xkSnimDajIHXD5yf8c0vOOCMLq6sPk0OT8uGrF
P9NANjQTRwmq81aoYM2ecosn5XttdqmyjpgmIVJLoE5Rkiv9t/aYZ2uALX4sYNpl0LZu8oDOtFS/
xlfPBP19cEeudp7YmiiuH1zJ2WHDZCTZwz8/UhXUyVwTyc2P2BtAR8JdeQU2r3tK54jGK58VxyOx
a9dw+4QYcG7naxtW7DU7UlDGQK52ByE2ibnZsoO56PU8zGITY0Nd5NPc4xBJumk57eneFMhaanYf
o644bcjBYujVvoXnRYE1aFUG3ljwZMh/OBWRoMAvkT7eannUI6eg7BzuEJMPRDA5tO0kcShQFV4a
OmXmSpj5cSPC4h9KmHdi7m/X+Se/+PSv9kosAGSphwLi8KLDvwXeg/ixEv7eyGYZRXs7tWLAKrTB
3Qtt/2xzKc5yGZXIIB5Z7N87YnVgurZEXlebRC3W4aWjWRJfeyiO1tQJrM5xUF3Lmvsu/Z+Aroqd
BLIAqw03YZXzl2UwzFUb37wrlLx+VKyg7KVC8WemtMB1R+Cf3FBtnclRhWbxVEdYr4I3H7KTxc76
KQ5dcB/it5Jv/Jf1uaFqcQr368/wYKMyACnTtB0HaJ+kxRZEQG1o27dFAdAFOksXyof17GUNF9p0
N4JrbGvuGSC8RFO0TE/mvvW1u/qA0Ci8X6bob8XIeqfGigHPL9dFB29qatpnKiM+81m5NzvYZqvp
M3U2xjpxr2mWrDXG/v8VmHd7iLjaZsZBUpZVVzMZCfEFHoRsbWXKH7F6ItXI+gjK0x9HL/0gQ8XN
1kPr8XDN4dthLV+NgzQh5oNm9PNnspxvc31972XML+EYZMldRlOsn0rU6ZIgSlXfHpJXsbjdh6oA
j6IawFArEi6rSfLNW4bgYXne1sAfk4hBsT/jf9DPoA/986wVSzOaRN+fFrhoXiYH4zWE/Cp8i4lE
mb2NwIqwliz6vHXztgTEdIPAsSal78iCHj6pHyeuyxCLrieOv5mbD5T6PuBpchMdmtt8ebS1eA1n
JyWnVJa05Ly74aap5DMJ0C9bREqOFNkKyelAs55LZXJX991PnYndr7pAB+t2htdXrrQ2JdHT9dsB
hjMN3msNfDVG31/sB0QURRdqYi7SyHwTzYkyURn5sIVAbDuFoqnk5A48x95jQsrNTGEcyN1mF+qM
4p45OsQ6qUFDcBF8lcgh4iIrnH2gH5RaehL7BhYnTLk8vstpC5/xzvFOLJIqruKgUv96kiUg2Hyl
ExZsXzV3Bfzsaql+FRaQbFlQLGc53yhdcSoH2E/GFya5VYwJUy2oxBgFhn0KODt5LCXa05+A3haV
XbUkPILu61xEofcob5UjjW0UDvEILo8cuEOW2QnlM+By3iDy48bT4WCkCNKtMjQpHzSLUHqXEpDL
MaxpWnQgDxZ3areFxUCe3NtbtD22+pPN/bosWhax7kY/9WXzr57s9KAtBkSyLCy8HRRd+jhXnouV
JmbV1fFdazs2vCZadrt3FoSieAmwyvtBNyMp8VpqQbgSha4hSpYS0iJjei6RzmoseGN2XPBvcrM9
PDtf7MPrgkQJwJqiG4L7zsVPZWY3n+ydRMchrzauLF3NfsamWT/y60JWavl3A0J9wR8DwUI/ZQXn
gyEbAcFMOaRi9MvvTf13Htp8yJCAlgL9JvdAypca+bB1V0ib7ft7ExhaULMQguRj4aBPmiLllsUW
et1R0sC+xCPHJCfv2ugL+jlcCRgSKfR+1/dzaUtecpk6596o0H1Db6IyoAu+Wsi0WaoplAMc458U
Oc5TGGgueRp7BpXtyUUqcN4pEiSoClYHiv9dKyiJAjSP3dK7OFhOKyPNj36ec8vMR8xIIwHzLbTt
o7+Y4PFAxWikJ3Lyf02OXWgNcat5kho8Kx+NHO27wqCPFxD/wqjDbhFJ6MIDKiI7RzLj2COsljWF
26OAYaxZspp1nBbYvPgS55YtW5+7wvwldh4lbCqqlLKkeZTczbq7nL77mQpXZL3RbwwyBEHpiTp4
sJFPw7zVgIOQXzmcYyOJp+LiqWUFkHBumPQ/roStv+xelj7ZouPmacdpdZyp3BHuv2cccIImBkEJ
WuIl0zCZic0ym0rZmmrlF6iH7hjQR7XOsiZio4/0WIIVchhHC4e8df/kqaJC+HnO0jsc/gMRVkcW
4cdZie7mBnuLc6+gULYbrs28FBmmPoVDwaYvBVUsvXXMiLKN8i56qWW+q0q915jEK+fA1+gYWl3b
e9mb98K4xlJzMW3wh+yCm+u1QPvm9LU07RdTdvhtHQeQyjx1iYdSHwFoT4Tdd4YldVMKSC9vYTwo
i6/Yo9VgN51UVP4WSXZQX+T1x08yT4u/f6KJdK95PXR0fU+UoLVlZ8akr89hGgcQYEOyTM1pneQ6
+RS6wruXqA2So8t6s8rutv1Tk6Qw+SipJzQyd0EoRQgMKhreLCWxFrvqK8tiJNC320K4X01IyeC2
59Caois8uCC94WYkuHhqN0eKFuMNJmAGF8crrIYuFzxSIU4eZpVnSbPQRWKSvTMgJZlh+VNzFua5
DtDkzM/vuIXfKy7aoGVjD1Cg9VE13zyvws2fuTIxgRjgiimLO8ZJKOuazteMux6YG4Yb11ahGWJL
tl5wztCChHvRtDRSa2IRFWjR3FuzRm9A3xpavm6/NhXpqKmqeTzP6Dx7UTe+8g5/LOgz3xgPjhp8
xU21rV7B720ZmamvDIS8YPyxdBK0NyaA9FfREA5ptQkkXv8SYvnB/5z6BZHPCouF6Uqf54gyamZf
+2X9n6zzqFSnjKdsgvltuD+8/vTomfiQQKwj7FF3N2MAFgMb2QWqrapNgOXhC5D+yOO/4vo5N9qZ
11769H80d7CDrt/0U9BpGdIKoq6AXfH423F3TiNaVrvZR3pskOSNtKzNJxl0To+jLObBmAIwrTb+
qmqF0fHFs0AAK0rkHt6FCLrR33OvppHc5JUHU2fFJK2gNtrrkQNTBQ7/kMEv0GJwF4NoQP7ySDmZ
4ZOyBnKKcKaM5O15ri5PhKDiajVQ0xwe5YPtbLNXHx99cV8eFppxNwba1xk0JC8TOYubbbQfpFCw
rAigH5CDN6S1s3Xd2ebcV6+ngT3yIMxXMbyYDDKeg2CSi4mEZ3vELX0TUFt8NUYleOHVZ3xYCcDB
CV9bbvbf9BEg7Oy0ViruVGUQqFX6AlFPfwcCPIhtSFwm+Kw8xzlM2XR1aTrbcF6eX+3UXRI5qMiW
ghfO/Heir73qx1zMKfLVQDzD7C77jOWuZFk75wg7sC6do45gk2bDpnTlQaHUgytULxvJmv8k+Mun
3c0mX7yZLOVVHcG6oE3omWZwIJf91IWiwIWJ5jrE6Jtr7C9DP6D7xd00PVEaLeRt/GzQvgqAjFew
kILU8ejTi0wB3qYaQxbxEnZBbvjohcG2dVmZ+ngArMqE7g+boyqMpD0PzNVI0Zjk1FuXSvY+ebv/
h4p6RVQZDWPsjOM1oQfbeE22/Xyjk6qbOO9npJ+E7ff1WarztN2v+/E/MGmucX9qgGVuP/1YW9Fd
00ToeXFTtJL1MT+zSIuNjdjnxniB23QuJne9APE4TgQeZ30i9obaedt+ynKf4pLFCQrMYgbFe6IL
ntKVC5Va3ZLqXACLBPX6WYfNLvTBh8TWFNb++T1XQSXSyv4PV2PiIuGUrlmnYiM4BAK/Zc4soHKN
DIuRc1dIhJAqYC0O7wsaPnRBAupmYBKYNfsw5Q3t1b+xUf0tNuUwC/fTvCl/P4Ytjuvuginuue3d
Jk1lpz5rQfRKI6UH9L472bKgXxbDCD8Rnkq+e9X3D9bzv58ONOmAT5pHAuReW/jlDyKElReEkSFj
e1G8TU4EG7N0Ipkv3rPvzAJDx1QfqwL/R6+kCFZUUfJ3fMdW94e70cWn8r78dOHKtphykaIvwD/I
cq2MFgXL1VMCw3cvsV7oLeeD1hI4Wz1JR5mDK2z4CD655coibSU+B8htqaKIH9uAs8MWBGbCMUPk
MMyfJMAFEUla4C+PYlVEfuKOKvsZFWyhjWewUTZR+GGr2KdbdMGB69/h6GC34sPS6tq11GgvfOYI
2CWcDEN7px3FFV/B5ngVRMSYIyNgT19+uFlFfcfbiWhLjL6GvNLLPA+l/hOdvIR9MD2nCMF3ZHld
lhfyLdBiOKMakpdEUAwYNApL/9OtjoPF34m8sgvwfS4N7N8u9KBkB+KWx8OYonNK4f0PUSRD9/rQ
H0T7HDWV3zAJd+GSloY7u5qSJo634yoZa6jETSIGh8GV7NDGQTJGUJN43FLUfwKI+0vIkX2Btzoy
nvI7KH890/QeYo1yIwM/Gs+vPvt8x1jLjjVcMFxIWetnZsXl0Yo/pn7VtlkkW/pujG7011fBxIEf
YQnnjlCj3JmraSu8xo39DCMukzShvD0Z7W5Tqe2CUW1lAcycb0qSQ6LvlGTaXSBYKD9F5wIprrlM
QQAT/swDKkv9jrAUClhHhNhZZTwg2LU+Ba8wwR1EEx/O39rIPi+9159PCDCRmUoHR/yT0syECv4M
+XEz8ZyDg/gHbUyih4J7M2+hYv18qUXmw9lcdHfyq/2Qbz4CFO0y+72d7+gggXKvF/xPCKVGxJ7c
FPcHkQTA7QJ9GSGsO8e7T1e8/lK6cCZ2nun9MhF7MJwi+VsBrGB14i6X2OHti1cl0fV8JtEDQ0MZ
kcTXYg9q7dqEmHYI96fEzlCrx05VUZvgV3FGG5memDdkmdOQJ/cmpYPz9yVGOQbKoIfv+PzdgWJ4
Xap3dZUwgHaMwTIBQ1aGgNq4S91PnCDyVFx0tfDE8ulemDxMGDaoOO8sXNTXDDnjbq1lR3zdEkLt
Zd4nF3Sy+UjHerr2uEgLV+epFynuCJeZ4+PgwhH1mxi0mQWd7nXKFICa5q7ay70om4HzBHww8ZdO
YdiNfBV0JfN7FSKWWjJB4YwmenWGvgEDRcY5B47UwT1LPXOGuS+UBsD1dxOUHMnBGU/8iJ56vzm4
1R4jzjCIDgBmsm5t9aZbk5GrPEKZlWhR9LnGzkgXOmNhrbOwAlGaplF/9zXVj6BAge+8gC1tuFVQ
VspgaPOygePNWc9LUAKzWrdAw2KPv0wZ4w9UhOpA7jMB6JVZameJWdESZjsxL1L522gXnX5k3plo
99lGEhbH1eFwhB5KvzSG57sAFDLiI673DKWie36361QFy2dWYr72r+e6f1l2xsYbBNi3xzw6oOOO
9rkgO/3F7JZhyrkUeVvW4qpdvCmVyZ4o0iixaBsrjykB0RCKMQiuaJOQYAKqKBblGkR7qjfpWKXi
X/dtFvmIX8wa2g2uf3cIzlrBbE59i/IY9SP8Xop3gis/T0IRihW6FMxBgOH++izmjpPbWl4PCl3D
fUMQhLPnYO5Fy6EAL449Lr2efYMp2WJK0jU1jJu0ondWdZG0dEdWM36krtbyGxxdxEh3ErwG/QG6
O3St2ULXXnA54rhpI0gszBxoNnUUIibJNTlOOrSUG54lzz0uhxnO1L6xhUvUKSA6qAqgfsXa9bvZ
nkIunvaxAPP9FQMkUEvIJzOdaW/8PCfYVO18SfeqbcA2DdnjaCwJJAAPsxoYKCOCUrNozUw02jjD
Xl/i1igEgRup28VEOBMhRzMePzk8JXK7wIUEg7LqGIIwXEc8D5dmDTdr6LfWLZ8u62RgDho87Cf5
8cZg3oQ3W/Gvk3vxVfBwDByl67nId3TpbTm+yncoUuPGUgVa7t4mggDlpPCvAREByL7OQyYxSmiX
NVoSqme/TQvdkR3CeSLfbUx5ymUtmqH0IAyOxGodHFkx/mj0Bk9ixSQ9K/YW5E3IALjKd5FRBkNI
JdlSy8n0r+2UjWJSICQ4rdXntH8PxOtYuesJgQ6gYDBGtJoszM+P8dibvE4YCffoob8TSPirx3hr
rtYhiMSBlM+V93rKjPWN1+9kdPt0oSaZxwvkLTnC1ay8BwTz1f2GPpyC8oEfwzdHtXpe9TQ+khXY
dfMCfLG+SzSsGnHUJccxEkCbrDa3rwpo0iLemdH5GKO1hF5ZaCv8AFCrKe4C8Td8D05ICmvKHODq
hRil/ywV1ny1hRgetxpUOX4qX4yAAbECpVCijdFm3uk3JnlReeL+gXX10R5FX45Oejy3eY68VAdS
VeQVdSLvGtDyRMUgrKpD+hto3fyU+Ryl5mNxcWPWGuVbQ+vIKB8r3ZBDmDJkr2Uok/ED2ejDVI51
G6Zsb9FAXCho8z6OaR6R82C1FFIp2aJzlFztbBI7SPbku+JCCs/LCLeIOTFKPI+6P7F2ajDfRUWY
UonDA+i1Qr7OsQYtTAqGrEqjiZusu6GbBYfqOmZqE7/J8eNpCLRs6onbiWsydzFPLeMkiUHdknht
8p5lruv1EHjIIxl9eXOuxpEhRXTA/zD0D/YYlub6FvJJeH3LUSW/W4IFV+Sjn+nr1pobtBGdM5PG
ZDnfnJGwuvmxCmp55F+8VUGqN3mbFlYypXKjKKk/H688lJ6fszfpQXmXi9m1Xa0aQCbzg8+P7xas
Tk8zW0OHn6q6rLOHkTLGsQanIKNX2fX6LJNCGOuIpkaUFRrtDR3eNhop6doC3WWxPj2ndwfmyB1q
5/ooG2a0oAhwenZJAGsx4wa7TuQ0mWsnWpO+asra0OfCEQ1NUTTxcPnV40L6sFOpAupbcjE/g58Y
guKJpG/0jNgaXt6WrRKJufo+iWu0XIcAz+VVrfc79g63GlefQ2+zDmqZmjpBNWihBaS+M5wUsKcK
iHtFI5LVKZxh5NjDjT9Hj19DDlD2DoSaMZlaVYMoqPB8zP2zSV5SLzQnMkt4uQO5FbqMmCo+q2cQ
WbnLjMqkzHXEvvQdXHMJaijkExusaW1DH49YxkcWqc62ktsyipl5KYZmLN1hegHPyaIUL8/nt7Gn
Ea5UGhTJJicN7F4ZlB4/hw8WoGexoH0TL0OKV7OV2M9ij/piHLABqMURQRTpCxPmrnuwHmjwp0iU
Ewg8jMpCfkeTyZa/IyJmQqsTobwlAJqDduuALM+ofYS2MB1kBP71pnGZGpHHKl9OkHY8XFAczbX1
BJ3kPib4wGMUlCD0+gL6xZnBO6bpGzfImVdJVbvUXu/HCyYHubMQnbqOpVMfamY0kbHc8u0do0f9
gBnytt8RiQG+gpG5oKMhJKileSioB1ukjo9HyINyPKFwdKMhrZtwl1u+O9kYf621gCWvqLK0uLsM
iHlqlfs8dnOgg0vuHo0woPgMKtZuhrHvjf9hIqsou/Zey/md0pxwOlcKzbmzkb11vFEZJvFVgcZg
w918LfZxDcliInGTnY6Ya1nNt9RgpBi6XI6aJmBe1/Jzx8qQCMMWHKl2Nh6mlm/mavfA3+gBwUEw
P+rpqg3U8zpb6sTLpL1rn3IWhMMmES0iUKlfz297iI/O0//dUmwO6MMQGB4Td58BjhlGQkbvKGPQ
SFA0U4VvLtMQeKc1y52QdA/XeNgz729ZeNdhZUdR5k5hUJuqq71zhoZmro1RRARb2JG6B+dnGkAr
EtKH4ljMYrpvZCelAtVkSYECLrov6qxDiQZaqLZIP5LIisraV6T8Ae8BfyVTa9kAxVNHbwKSpooL
uIFuB5m2ruMquDTufMXg0aa9ePGeFjZ2pBHYqvG0GMXFfVa1SGItviMO2D4NpTExSZDrjHLq6abP
BUUJMG6VQcKIaJ2VUbaMZYBVUkUYuCK6plFOuBz3CT84HQxrFMIqxLdbSgq8g7+MnEBH/O52z4hD
gOQ8ngJk1ScM2afmhoVpoxzgY+DKG1GYeWVG5Hw7+dnK98LAvAnhfYIL0IL/jEBdK2x6Vio6tHeW
CyyUsq4E92yysMT5OupHRR0eYYihHkiOK0DOPXgNamHia36vYMMhWQ4TRr7R84SLIcvbNWW92N9x
JuSS+zZmxPFmkCO87+cEGSBMlsq9/LrQH6PNnBsuLx1rbELgYrL8OQCkdEFYtRkFdkFNwqI6SJvw
L/9dpM8T/vcGfO716fjIkGGkzrJlUdYvpJF5z+Myz9yXTl1qIKbLsq/yPQIppJOkxYZjz//ckA5E
sGcfwrJQUS4TXIUfTFdUAdkFmvQLsXwcKwGqwVvrtacB51hVW8GPLceJ3AGyYxeGaOZqgx0OgpmV
QDgkjUFa6yMnFiY3umw8hAKboEyXGSw2Y4EIhEzJpg4/amAVCbUms4iC9dUsEpmCOsoAQw41bZ0Y
q0FwMNrN1gqH93SVdY3AhsaTW5/XX5Z5IFmFhmVXIdzhnaxEQrkGIeU0bWeALz+qlC6tmQxb6Im8
bomDyw8hzBnDEiymUlVweqpi2b50ss37Vr4jMFzp4ZirdKGtkxEYI9XmIIPVbHkrsf9I3Djb1dBi
yDHqQwX5+OvpTS9mQsEbc0nJIY723RaWm2qziga6qxNlREQtt0qXiISv0AQALk99KGSNiKEh6kgD
0qOWwNWeopVpdNv84TqEMhPUN8oaKSd8NdhpwSR3LzoyyXJ/c2yAmJlHrm28n6EHoq4rLaGIZ3Tf
emYl/v/ROtGCLgJHg3TfeUhJD4yo6I38mSDGoK82noqGM0riEW40VSz6oBxv7MpGy2tfaBo93vdY
0z1GzOmRjxKJ2P+VowbC6f41E82EUYkgO2PjQ4ZvzS6i+kOBd4rhbte30fnmvQlGUblPXbtpcs5q
7/bdLR7jrJ9GLN3wfnxmEy0CZfIlRKs/BL/lKm2QAr67KQDnHxGp8xzUJkaj5qSpZ6YM5NKL2pS1
3KCVr0GdKJnTQzHHp5Dx8DRbuOoqWlwB8P98CUpEWZqWYR47aBTkSnlZZFH3xADJZkC+s2sQtuSj
n+TuY7gWuHbvO86I4b86ACDp7Wd/elkgV9MH2qj+hChu9To/UXdfi3SxjGCShaICIsNQA1LME075
utrFRgfl3hUZjPtxiaqCiXJ/yx2+3sXycLaJVhF6L7J/t95Qw2cWXQoGHzgNUqSYWYmWpCU2TJQM
a/VGaHIM/Q+siscQUtfviVhEsbVCHrAqjvRNQY8lnEK4uBaD+SPvW3xZrv1anhv0eoCHZmenATWN
20J+d5wYUdLdUPOrVFDiAuEnKtcThzhXpECF/8AmO3kYvmV/vPtbeNBVfyi/6Eq9Lj3tj4XOQwwP
W1n+CSA+i/62K+RgjAYrLvX4mKU7awGEWMI2WRMl2+SgDwlWgFRncgn8uolNmD26dtQing5ODnq3
o7Pj5uaXIzO84BT/cRPJfpcLU6m1sAuz2ggsCudK0QFHVzGPk73TerOIfH4xnEWQfdofJF1iApZk
UEp9oImJO3Pn5S/rWkyDBd2xGoSEcsv/K2RGoPyRVb0MU8CcoLbPNppOaJ5agyka3/zikWgHQoWz
R3KzZQ77viq3x6IC9rhLJeFgPg147CeR7oEZV3EhddKzieBI8rdu4M024QYrkH6ELFzFppYk3SUi
cVYXwOnUVaW6lwsaQIzg+G6C9Q8pS6TiroKLefRlvF/ImXmu4BVtZrGgNEniKB49IxShRQOjM4HI
ksTI1gu7Av0S3rrwTYflFA2pP/wwlakxe1r9YIyu6iJYushzbYwr8QIPevYpf7twJC76T98GgMXa
hjOQeO37pH9EzzbALgl3fGEdsQP5KfkWN5YP8uJeLm4UIQ+hx8n86XDiChgY/IHlW1qGwmBSv2ol
zW7IOOkxH7aC1P5aOl2RRBAY1o430qKIqLBWB1hmlXfjXTnwbnoQB4rFjPurFJ4Fa8BM+dY2zGqq
76t8Cc56zLqZxBmoNFQKvmYwMa+Ov8ZhmPO2VAdNyn2aRLmY449ZcIVUenGFUyMQZpjzvqLqk1vz
vagIJXaGuoxL0B6Ri2/rg3YXX4DT9XiUWJmmp2QKPCCEqiowlZPbP0ZeKCFu9GHqwo05soT8/Ctn
z5isysAf/Dqdvn5B8XtEtlTC6Roapdyvb5eU9rzKbMwBj3DzEj11V+smrh9xSxfSjN5LaTTc0x4p
uEGSHkXg6efrNakLerp4cjmS/G3PAYTBiS2ACY3VlMsWgNgxcnEuNwsDyjeFkEXzBPhwYd0olm7Z
vyc5GzvpituOrCRlYVdLQuIwPArJXlpYFfn106TH/UvDrVjXy3JockHdzXR8ndyG/UnUKUGDhJ8P
PBWMbsUd7RsAJNrPWRKosKYI7OMx649Yc39t049aJH7+bMGzcegraFT2ER7v5FyY6Lf24DbR2CDe
5LiEwljt48Nrjo2VUzqY03Vr59AQlVcYPlDkj35Q3R4YnC15098/ca1QT8YqMs7CiTCuE1Y2YRAH
ZERhV0SPohmBgo5oV66637sFPf+rww3sUI2iG89SbQXaDmQwzSPhKEwdxKKClsxzjSnhIymkzBHz
oW1qF7oEPsbJF8Umnj2ZHtWiI7FG+bLOyao1lCfm4suvzdJ0GptfSQdUDHjYPHwJt8NwhQeztnxd
pTbJu/SwWlqPqXka8asBaTGYu9SiNMHMU9bNAmti6txFsX9GigZwmodC1y6c75zwWKJfRaPdxU5C
hQ+tjBgeuIo/0D3WlMZoePKLAuIaq+kNxjtTRp/VRfcKEp5byjXXsAoVNqI3d/BKyvl3J9l/XRrg
BfJ8lXQQVz5m3XnXQ2choEGyW6UyuIVWXyZbellvWb0DXOdYcSxJUaCCcl32v34UkG+pFqXzrNRo
s5opiBdNW6l0aAEf3l1KXKJzScOdcKif7eKrqHvFy4O6RYl4G6P/jsj+iNbzhvRRvckxExTcvRy6
v3kTtLLbbwbpUBZPLY6R2tsQFmNwYEtvcOjwxJ72+SToWxNteArNWE7n6SvCSO2JD2LaNioZnJbX
sTP5xwO1ZyNS8ZulbW/m6BUe6HRjMRCphjp1h0zqHnE5GdZPzHz8iN1MtIHi0UOBgWh7sqj+CJ0z
ZtWDfm5Bblw4lTAwWePxx80Oqb8kZXgwlfS6CO0N86aMLE+lXCF1sB7T2bl5IsGbug4gLpn7WOdy
sWthqIsL0QZapzR4u9jSbMzm9+u7PIREm/udh/MB5Vfbd0ocnd5x2+HlWKZFXrRidMWeh5EUJYmg
Vhya5BkuHb1fFfsYEl+ast5it9ebLIqGjkgqWu0ZcvBCpGFD8qNkj1LbF+KYjOAf+Ge2TpAg7py3
pD6IsbC5aGAYEwk0J7W6+l6+fRDC4gZdt9jhPIH5+yBfhoPnLAxdRpE/d2R266FGmSYG12h+zmcj
lP4bhLVh4iSCYkVO+ndBJyKWcJrdZvhfBPNZ8vFnJ3rMQzfSA2s3ZsY5inbTX5Ys2ZR4KXKfnFWG
97+7N6xqXR5wuM4zK0Ep40yyCuWu0U99wf1u0fNdHkW/Yqbo7Pgg1FUInmNJLpT5jwIj/XzH1HWH
wD5RsFHbDfddqRr7PnZoeGDajvBgbXGAgds1/wSY0sdhhq8bfmIyb/xBOCHJcQyTrPe0nswrTjLb
U4nlXVxsxTV+X19Keqh+ZcCILSZKxyEtVZDYYFa28hyQ8+VYhrvVuHLIEpnkEWhNjwBGGkrvbNer
6jTbf7PgjgPkN8l4fe+ipdFsOvWe7p93xPrZFpjpRowifo+HK79mqLS212esoW2DaCLxnzgE3CpP
dLbyD4mKgBTyPR4+uzpOG4ej3iRKfStvsu0h+wL2B7AAKZEl0oLFAs2RUifZn43C1rr9GlMMW6/M
LI0fqby53pggsMJzaszLZg/lFzywsAM4EXeEyXhf05q8tI10iQQdaVKH2PbW5UxZ4TJhkQQoI8k5
fcoP/P6PcYxADlzcTgENYzSD5zSizrpcD8zRarxxqVzPK9L+bjSG8kZR5msCuRZs3NvWpRcyx4ri
KFQWuU1700tUDb1auAJovv+lClJ8+0UEy50gKxNSidsgaEht9/SEI9yq+SN3IcowUIXOug3ANSYO
PXRTTdvXqyOPx3GFc4de2KLsEMR9Ewpw/UQcabLkGTkqf0E+2130DkxB8Ealtq3X8r6LFN+IMmpv
K6jlGo7XXjUNMiiMLI135/CLPjLD1shcBQUNghWX5UPLA+68EbpwQhzCnlUi30jscwkyXuXZ24zv
wSuvVM+JQiA6WaaU8B2/uzg5f9kv7Z4y9TecreQzKAPiiTj3mRHXHOud5Ffk51AOixwvK0rze394
EKngW0BZRKTMc6v9JLVZvNfeg/b9lOftxaeZWisi30yGk5cKVkxGF7s34Nq7qHqWRJBpwMC08/IB
K5kNsGmOPqvxrhUe9hd7Sl5QqKDXqJXn/2d63Vo2kae7aWuhiOrNFoUB3Die1PvIuPO21X24QWg5
PGcKnc+b9j+UT4dE5VWFtWVmbbUfnQ3I6bmuntpDOnI1/w+GwrcffJ+AwJTfTxPzWe1QwnAg0H6E
PSOa8Mw/oOA4aOeTa3l42DLhYcBYZlzN9mqP6ZFN5QA9SYWlbmPXuC1qpvwy5a2zg66WkIMfHrIP
+oPmhxx3CV/LhFdZk5lZCpR0TleGgPVfCOGUtz4EavwTkpnhJqkw0hApSTGk7JamGScN1IZ8xh4d
Uz9SnAYa4Bq89u+eih5fNq9+NcaGL03UJkaEDQw4v3IAec0PMpNu0YrXYDzaEUwFwwqXBE45b3Ad
vsaTFIX1HO1hx16wPRH7uktaKi64v/G/dAzBkcGIwSODwSIku6IE0VnsZnI1A3NFO+9hSI/VVJgg
SVGQjkmiecb6SN8qQBIm2KP6KHMqmq66k4/qCmVFqAqNOEQF6EsmuG7yntax8awuHVLgJ+WsyMjX
Ns7mZSI4XHJ4gVD6s+/f6ze0Jml2v3hNmUpXvEyLz7bwfVPYl7GiBDV1vmyHkUF4oz/kdqhDECCP
hG3vG2rqn2sLDyxb/Ok7dkjlrGvI7PvzJE3g/5xmYbo52pd4nzb8G3nzeBcLXRtFSGI9qQ8ddV3d
vHV+EYwYeJeA6bnZHkNnrBMKaqaG6H6AQ/aKOD6y0cRAT8XWMDGgtMRPLBVrg5DyZIAJ8T+RVPKp
WX5GAPLkaF3Np0KUKFUwsWk8vZgeshS1hKsN+vbuQ6UsmvfIgz/nL9vmbMiJ4sfwULAld8EK9yE/
xfj+H+FZQqt9qPOEyjzkYXGH/bccBbhMAhbfBWK42ZOw6qsNaa66tqamRpV1O6UUV46C+a9jJ4iW
YjGL6P97AAeznCHssWAQJK1OMMu1OIvRHIDboqRkYAW1mIYyTFawHYr1nnxtnczfzXU/GQk+xwiT
VNm13LQ5yGTFJp4humIdw0xtgKaIDoNLkXbJjFTbyMb1t0eVMzR/Z/2u/l59b+VOjLsMRx9SmbWG
D/54oahTKBH9g/Fyx4PEMfTKlPZsFINTQJtyFsBqWBfxtD7MZeb79kkavvqAHY//5momHoeqAOp2
MLdEZQ8Xo28o97TFkw6S6j5WfghrRki9pj5uN67MJcZbhKTwQoD9xS5NoPCWw5hE73vwHH2F0/DE
agviMDaPecPzB15Ck9atql+dMabM+4Gek9BgBI3mMs1XUEZ35Qen9aJofoXmv3OQaKDSpBp0HcU4
PPXTTEE0bMwqKCn66GQsH5kG5rVcvrREPEKdFP3MmvURN3aJoGqYotnUG/FQhsx/D8mv48idEC4I
29VdHQUnCY+KCnDBMDRVyv5og4Qf5ah/8prEU9UM1pS6pXyp4JSbCXkxb2O+IM5tKxZWcd0UxAhD
vKt6JkErUobiy3FzuLX/vpHAplLftTZ/ZBSz8NfMUEue6ptb0cmbLz/rI4PNghTz27txmITKQS2u
UX2LZ34xWL/9M/TIOIiWnc2pf5bjR4d8Tr9haSpKSBWXsyslQP03n/M8134lplrWaU8v7zZKXT1e
cvAZcL0PGpOK6rDr2VonNd1KN7BFm6ACROIy4tFpbNSGtfO7zz8rNrZrYhc1/V955NPFyGa2JNJM
b3leGA/IkzZr7soMBQ/PzUJwxCwQtBhXiSX/L65RjKMZQjlcl4XV2LzisITL4yoP8fWVTgx6Y1bc
jtBpR4y7ksF7Hm7sBZRy177T5C7bP0yJPaZsz+QHPjaYrMcNLsloFJz/dANGiRwzA/bIwkGoh/M2
cZLOPvyYphb3SIMbeVHs5dYT5a4fzzCzADbexzNp/VhKKKIf0TAPsZFdrUTZHPr59ffPa3oGPHM/
NrBU0AjMkNrbrZ0Q7mmvz1cRpNPvJI9h+c/iNIAI/b+LyQMAzi0TuceL2feTAEbP2SyZYgI4rW+t
IidfqKcOQ5IJZoH3+c1ALezyK3lg/FfUWv7iKcWCT4VAd3s3CeY1Dt2oo9TzuH7bs3jmGyprurVD
dou2n82JhwTt+PgD/m4YCTGsOPo8O831gM6prh5pq22hypSeSBwgoziGYKdDYe6M7gUa+ZVnzGDu
/I983Zycl93BzS4rnSu1UTJ47mcpxtuIrQUp7OszEsMh3fj3GOEPy03cp8UjfPem0WAP3U9X/rcs
EeZPOciDMxXlOMn+NHl66FXtePqQluQegfIcHe6Joz3Mp2skS7is44aMrQR+mOk9Ly5mcDSzfyLB
ARg2TuhwGJC+n193revqIAXAGYEQTbkWfOrgduT9AQySg+7A/KX7y1LTBhKNz/xb7vJUnijPvoxJ
MK0En9wXtwsaYr21AhAnud0mOAmouzBsfajMo822eUWfXMoeb/wJj1d70n+nbDPoiCgVnffCPVpM
IUUpAzX0dRj3Y/XGRBNWael7O7q6D79yOkzuGQ7rdcxvlln9CzZpZgCtlU6dR6QpvJzyeMuELyZV
i1FLctWss7BsvIEM83CIeSrXZdEv/jzwCNRtIB+pIySS1E3re5Fkfnhnc9SBAZXwz8Yx0WPSnweP
MNrYeG1IzobPhMISSmf5olDZY3qD0+QvKBr2BPSlW3dkGydblayb0CFkL6WZUq7AIMjWjBuvCiGM
OaXFItNJ4kL5oqWJIPSTcX+B32RiyeefT3z78QeMLRYHUaE3xFo6iXxlSRktuSdf96bPM6jmqq8y
2zgB/9HAGNgZ+iZq/x+09oxZxR1Q6wVj47Pm+oUXvx0kwbezTYFICpome09ijXWzuUeBM/nuqmrJ
sf0badxFF43xUt9NKnUuV2BaStJcnV0nHHdjqY5Z1OlwqzXryNocMizAKpcRREXtBzJTBQlP6TZV
d/VzgkX4SkmfbJdKrlvoEoP0zrgkiwXgQt9SeKuXN14usRA8ydzbCnwz1seF6lyj4adzzBDiNOts
elhIeHOnz5G8OhznRablBqUb7EVgl4WgP+E0rChWpPgFmDA9zDVp1o/V5S8cMSCjqkDrNkaPZCVI
s8oVqUkhwFqr7a5afhfkBOsb2ckCey8YwrnsQYAAOWCSSpK6zW3V0K+j1E9czUZZSGHx2/9FJmvM
a6ZxSQpyBL9qxTkYf6I8y0Ds2erWpOu48VUqUbfOM6AWgAuJpxKSU5wtLtGBoIhcr0MbbA8FbgN/
60UxD0262Q8VXFCor9T0BYgYlhX0qrgXlu6tuGSWEACHyzqru2MIQIJdSPiX5WXJBkR7yHjbtvxj
EFzLHuWvQRbv65A8Ob/DpdxEKTwPJG368JJszVYYcvW1IkBo5PrtrgBLr7qEkFPZKw2spQ4ewNu5
3LNB/DYlQfnxucSzJVPvxsBUwqiBwQN7q/O6hlbZJOsnVRvY9PPbgy1Y3BhsMY0C8KU/EANw3LFn
UBpvjZxELSf7TF6cX6CeKSMUssSSL0MAsek/GqxBdZtyFBElsI3rgHJvi+G//PHf/CBw6J3ZVhQi
KbfxsMum45ZvjT3Exgj3j+bm0qWvzD7vRcXdROzKta4+jA9bRiXRb35oP0LDWzCefCzFbKY7il/h
keY3djiCgsUemqtUE3GsUPnQslG1gQGep33oI3R65T35F50n6ASbihfowZ+g8bJKQaKiyjI1XWCh
ZoukIMvzZww92TTc0vb3FEMi8qcPQKT9Qj42vaXnBlH8XN6CbAXyOyAuN8q3rgjjhtosCcAKZRRA
Rp8qw6rqdOfhLpBQ6o64/+Fx0RYn7jvlalOFYy43OOqgngVdjUx8Tt72SvzodDG4DcgaA+H+WY/G
qVIk4im3ocY4rd6THnUB9YxgE2VjbRgCOChMHU5I5xJxWrvuip175Pj57qp9ZF4Z7xRS3Z6FYHuv
roIPvI7gUvAamLUMhymscPGtak2qp10787IjrMkGIQYdN3I3NQmP0xlZzLPuFGljLTPYC5OOd7ex
C+BTK3BR67xBfT5TgRMkxPX4OMazSelgpy+JBTNpuChemY3ll8Yp60EowCrFLXkMpXXOV0bsdfJl
z7iRDJxL5TcAMTqPIHZc/u4NggnpXfRd1Ct4zfWQowmHFtscoF9IJk6ErKI8iWKM7pYtoKkTTS8u
4aPmj/DozZH3sjBEUSl7K1JHjykpkuVx+rBYyOZDyfD0Vj252vk3FcJALc17vnD3jmg09idxVQit
YyD/phpNt8N6QQnDZKEfAlSvSMZkUZ+BWwzOZlO4bbK0+fp7MjuTb4UdVdYevn14Pw15kT3MJHrL
wd/aR4g6JsbBiRPEpAUYLLRztEKZ50TVZ+sB2OK5901TWjXAvaxSgLBP1OlfXGz1B0ms/0Dq+ezv
n3Qz5f8C3R91PSbkP/IeyNvdQl7b03zf62GBjhP2bMjlW+Bs/PXK5aOa0jy9+VkHP6HdVFvfzC00
673Z+/Nmg7jpgqzcq3zy9G5eW2cDy48YzeUAsUyWMe+MjNSDHMhf3meNX6nld1dqiwX9kpH+g7pn
J5Ozsse6jWqjKqv4o28UjLxMCLCCekixr/KOFrFZNAA6qVDLBaNlQS5TSu2+zNJn0M9jl2BL7cp6
I4IEHhSOA6BQNe47ur9F3I+BfdGwSJsF9B2h17tcg1wF7qFRq/t4MSS0Fr48yOuajAtj9STfP/WQ
qskMli/dcltbCh2MDrFyFOj3SlblA/5msLwwG1SUcQoVemN4XbzMjfjeJuBy2ympSBX/2maFCe3W
T0l3GC8SWE2bnnrwVWY0VfFBLG9+FkQ3NiHEjrSxVMkQ35wtnX7pvULL024X4+oCkC2gRub1N6lb
AFZ0Pqz1/v2XPeRDwJmRQHpopn9EGXOqwvG1TD1Cy4+B2kg4sWc81nMXKpdFdOJ8P4r+xATSPZXY
v4OSPPMPDhG49emJgnA+lQshvdSpFvC5VW/NE+5YrN4X4orYOADabHNjlBbBAFyxG7++Nk9QSTiZ
8RVzxfRzWDCGj2bESI5P50qiFfsF2y91onLcaYO7ripRtdMwMnd2/99SfwTjx0QVsH7M3dUgbVHw
RU6odJfAS9IG8egNBvEEcYufwiNNowbic/II6vLB1QGDaeyvLM+8QLIfNkjefqIRjIYUoylgoQf1
DGNlKJbUop4qiakQNoQdRw9U/vxqQEaWUKdMrCi1dntUmSDIYjBfcHukwj+fN6Y4la4ejmMcB6LN
LSWfse00wy0UxYn/ZMiiLJjC/rFVvvsRkfC7GTB1vZ6xONTo0uWXvtNEzqb30RID+sIU1cNJ4dCJ
VO7wZGOogHMRg+Szq2/IdxbN7qtvw7Rlyjxh/0/GxObc8l2b2NM5qSjsBf0ragYzLMYLsMMnalvL
pGBsnb+xyN8EWNeppdcEDTSUAc5p2c8UT2YoZ1dUyvBVO4xRe5OgeNZTcyA5J+lmYqfq/Uw9aqcp
aTrfFsxlEgjUhkev3SmgSwKvMfuLOe1lNk9HdjI+0zK/frJJA56k08yPRzT6DmH4FycuhODd9u2l
dh85g/Nvth2U8CCnK8TMAQHUJtrkYA6ZYb4jxKo6927Bvd1DqU9KHr8UGE/LvJDv5L138sCay+w2
LIMm4mD1q4/i6he/z3ywalyB25LAQ54h5YzPZNj59HjTrYoTfCby+tHvqTT3jF9i7NsA+cuz4YUA
tathELMJn0J7Vpwr5TK+9woV2NPF0T24p7pnWDtmb6B0yw5gaXF449tTzsQAaQNHj60fmuKLyrhU
wclwCRAE8vFSpio5wxRSgN+7wn1Udt4wplSTfbk3503dgmMwi+LX4HVcIrfaZmA5Kc03nMlC8UVv
P5l7NtRDkI1JnS8ZVn/U8Boq0qleSLdN9zMfUJCUR20uh0xiRUk7G8JN0JmycwLPnOkiS9P/w0L/
DXxv28WHDTPQrv357xSbGsZ03xUcy+MGpT/w6MQzKpPH2t7W3cheL2UEbGe5sLXGaVfU/8Gct41B
rD45WtX1WUj0vrIUg8dormf3Eh+mLkQ5j1PwBK1Z+E+kLquQugP/j7yWYg1+y3wK6TqwFyw+tK3b
2COwnPKtV/oVIqcOLRJhudh4phAM1LxI4NXO8Rr6CJOqq6ZiK58dP1vwO8bRB1+gMenXeoRQCXY+
BeD0adE6qn0H1Bq0WlgHTTTfySIe2PHXyM90pI4pLwXi5NQ0OajOCFW1JBgWetqYoEE5H5g46l2G
HEbSLoVFfb31MIBhaOdmnz87BD9q1nLvgV0tvZn0m1jdphS/7PJ6VvWNJmjLRud48zA8dyDfJMTQ
xbnWu8bXhPbQa67tpW79C2o490UlHH6Tvx72bcts8aDr3m12qEkya469pxEj35Edt6ynki/+RGVv
UbL9TeNqLCtJfEjAsgEBXkDJvMoCLWwrUJj0+ML7bzI+6Mx4fTa6AldMA6qYQskC8y1MzPmiQk8U
y70Et5gaYrv263ovAZkgXHYQulRmDUVBaY4zKp9qHVAHeHn9qBSyw0xMyjubHa8DxrT6soDPLDnP
gvTGVWXpD8Xm2C7C5dsziax/2ucQ8sf6iZoW4I7ClrOQi0nthpYWflFdjmTpdf8tu6wR7Y3EJBSX
Z2bKhfTuPvdxpNIqSvrGw7d9EydNJOnraDc37SRLcyrIukUu9KMPxlNr166yNY1vK56j8sLKR9b0
vsqgayo0jWMbymYUKuApXOa5DK4sJqzQ7basoDCzS8I7OtzZbCqxN1rfQBJXEP9QUbaYncIMIxvi
D7LSImoEt30FfE2pJL2uaUZHZNA+K8/Vi1WW7w9P4StY1YdheXf+4aRoBJce3PsRJY6s0QA85vjG
EuLpXvdD1EUW36EFp+IQlZJCQtFcbuvjNWeeAeVGDm27a4V3/T2clHFrX9qn0vk57rQX/oTMDlRD
wDlY/adbJeQo2/gY1Dj/SQi3enOZ0M1V0L9/gGFPV+KWbQ8+ExfW8du2dxZrpdVjLK8v7Chg/1ha
VpOb3CZTLXtlDrFsNCel3AgnaWyQoxFSAn+1LC0x3BiibofPWa0I2x1bsak0p1hWybXzOiDWXajO
mhDDjNfd+CY62RKYVscktxG2tK6ieNIjFCZqSPhlJx0LXjbVjd8O87lb2+xQq4jmtg0Rrxi6ENDV
O1luFZ5InEhJeQR/MgJATzKiJXDWpMFtdHyGozR7ZYw0kCHHDOhDfYV4Uem1eEdLdmdwrJ2We8Gq
6Z1C1bWoAtpQUjoj5NwO7DDNJTJtAY7o7aBz8xmN1UK/o+1WexWyWnHkPRbdNlLvgARw5sZ9uKUL
A1t1jNDt2WaYUeMl9w7Ki79Tl67Ck5uU2iWFG6qk4U0fPaquTd3SoMneMDWoJXX3891z4+SGtGB4
6kHghZ1O95OJdOdnrmjRSnQJ5F9UC5/madZRXnK/SlrAUL1PQmroAaRnKGowIqFvGJ1NgoElTbF6
95o61E5X2EyH5RUIEvEhXECTR5Zy93u1IfuEGwZXXAWqz4gjRaylctwGDdZCdi70mU3QGjphlq+G
rAHODXqgLdf3IK9KdXzrTxpQvauvDLByQpU+EsoiSFeCxU8c3dxTWlhvd6C3ydqkS0may0Q3t7vz
XSk+yjDFffYU6GJPi6zrWAotZfoAQHEiVc3gzYdCeY92/YAa3t03HPlMQfvMQj+8+82ss8+zQsV3
Ccx5tlS0acFIqV0y8gCqQZmhNULZtedCgzpxaBMMu+3Z5eDqGiX5XVaKV8BHyM95G0jOtWXd9vL6
EZBZAcG8gYkkyvRBtEcKYCeAvbea7/mOyXRerQawxlNANqou/5GZahwAzd7kihEtf2mUbR4+qcL/
LwBeY+0ARpDnEyALcAH+V4mLJrIbmK/Q8Ort+4/DoNHIyWVuurdm6rz1AgibVxHQDtp6Re28/RyE
ZrSO9kD/dGUzjyj7hNEvqBzVnwr+x5Ae1mTE1CiOWKpidIGodd1gpp8YUz7+uYEmEbtNs7iLm5bv
D51FMm4HtHz0cUsxi/XYejr6CNXO2eX467hIxGKCo+KMYUqAGzTFcYkNY2ZDF6hWXusze8IVF0R8
7slGEZg2+PyWrxdqc6fS5y3F8nn4qrA6w7Ylot7uzFUfRFU/TesKt7IMg4QMeTOYBntkd+uqigPD
xK+7dvhwbjX0XEtmtFs95263ZQol8VcEgrBqSBKe9Xz3RY83YW/dVLNUvzT9Z5AESNPYI5Pq4dPb
FJ0aHNdpnyxdO7WGK9i4bIFbNo1c2PojOXwv3Dr5agCKg2UPlitPw+G+qBaOsxHw9Y8dVCCgJjAa
pfeQxW4ltS1rNWcUWOpgQg95bsfx2KFPJWrvK5OD1YHD5MbKnQijItdoZQr6LCUWny/X5/FmvIp8
Y9Gzu6nZz8qtx9o/mqgOg9pFwQW0Gd0DfUX8mfaHgwG8LI5JZZCtsBCh0P6f4BtlxFd4Svp4LlaA
femzo/XJ+nmVzgHZPWua95EYSP2wopVMuU0/UJuP2YXz/XBpXIVqtEtvpIHDbPSYIWoQYb2c2TxG
nepVTU1wg4iCEZ/2J9Rv8D/UuIHGPs3q57eB2nllpOdB36973FAAWrldQYJwg7xVcFvzdOPBOPN7
9kGftwE/P6bZxYr9Q0b+wd3FDE64tCKSYwKVRMXKPEI35FfCqshBz/B3tEpSFuE5JwGtIixoIbXF
7570GO1Stc0OBZivWphEwdGqqR/aiXoSvAj9DyTx+xHaS6OyKE2YzpxDEATvqa1a/XOySM3+GNUG
HTpFE16186DQh9GU/itO7PWZIOI/QtOrV70IPohF4W1dZXbiY0CdC1WpfnNGDCobP9bqUR6Z1UcG
RfNdPdQt7FcrVvMUhMnEfO+SRDaNC8lmxMVnESQOIfe0q+/73t+gm112KXJXYMdCCD8wRCJPikDF
BPTNMZzJ2pXedI4aaYEMiVneThron9GmCFy+jozzqutJK5Cs1jfRtcuboAf3sPSpONLZUvAP0Yao
xu0LYE+HillBnV9UpXaZ9u1b6Zea38op1W+y3FjZ71/B7e6f7yv/ACS/DXon932usAGOl3kn+svZ
3T9PinO0BS1Vj02YNCvy4mmLspvRhTDTHvISEel1UczYVaH7kEoZfJmPTkHecF64EdbnTTDvLgEq
RtPHeldZQIuuNLrLf/Rk5dsEvogwmS+x7pbh5uAOOaWAeODGXxDA60IVIndXJCROBTOY+8OP0Tni
avYpkPu7Ln2IF/P6Gp5IL562z4VFthZlos7sjuCHrvwSTvh+W09b6hGXhtNHsXQsyGH/PsWdMqez
oNNFxujCRzxlqfzi8INob9dTI9AKtu3xTSie3aUJRkWV4+yums5PY4DF9znZem40bGVuC59yJCeu
Egf7PLR9Nt+ImqPvUznYIlo7Zg5H9CVwiS6t7rEz1EYuNmiwXTlPB1z+g1k6ScLx5NxA3DZrK8LO
7Xs5JBVHiUZwro8XBpLdFjSwJJ1kDpLJVjd5am16u1uSrN3Zf2jgdoPYaP0EekbJCnvstCykwwWt
tC+oS17ICfnY0sOqCUC1K1Js/2+WQITTPEe+KbWHZAydu3dR1Y4m8QzPcZrsPha4GU8YbKi1V+hf
xH8CE2Iuu46tnDr9IBMWlbWowfiTkTQOYbOOL1y2P+pnUw9IjChdaxGCr+OXiSKtkv6XETGhb4XQ
6xXXEZAwsmUlURjlGF08lxb+Gp2WimXPK+7SMmrp/Kba/7qh1whXg3tikeChz9cuuJs/5+EAS8xd
Z5YWlYMv6e7ON1pknbrJNV6IcjFP16VkuLTwTNkvZuYThAHYOrDKdgPLfImIxbVbCK51TeYn6l2A
hPtQ3eru61dNEXwjvN4yaNimajslVvMvj6mruGSOIrcIKZ0uM62Px7yZhYLsuj+1RiTOLKtD8d4E
2UlZBrOZwPK/u5QFMgb/Atd4TiZZi03nIici5akwlI5lknLupdt3wk8HQ5vJOCz7hM9TIvrzP1OU
WkGA/SAgqffzh2kUV7zZ9wIT1EnUl2MQih7xrVqflyhNPLlI5FGxvjv8vqJmqizYDJAD78tAqUyy
nIeGtiwdtk5YsGlualpcMhJitBhqlGHxdvuCZuOHlr9tIYNtjuCXiST86V11enQc0TVy4XgVv1Ir
jO5N5mArsYy4OnFbGBcW3Iyd82ID5QeBpeA7rG6d1d4lU7ouYmlhzbsprPwOGD8blJCgt5pV4HEH
Ba7YiBaFlqRGkYU51jA4onFIMbqOwjeuABneqow6s8LsWaV6goKS3/fwPhBo/E58MpcSlsHcZyC8
byeFrimD/f2sNk6AvTBsRs0D3BsVmnJG/KSxunQW6zJK/Zd3nxk2pAZHUQEkav0KdCW40GrWZXn5
sUPMqvbXdnrF5NausMRe8KMfLh7rDbUZP3dcWL4jEg/eeGSATMfh+cjLPP3DEpfrGToA8aB+XuIK
jZXYQ4H/mCh3gKt5fEgSxY6YF5qXtTnAN6vxrQjeIUIzKIIEcNCbIXo/BDRZZi0NjGQtgZA1J0ml
p9a9C34GDA89j6IJ2dyPXAufzG+DsNg1N0doWawQEEuhbqOF03s9u8DdZdGwJuPcLUNWaJ7N2ssb
+AKPcNvrKKfd8xCDwVX7kKCuWAgPRDtMAEiTM3cJ9eSoOAUrS8wFIOzFN/A1eRah81yao9DOGZTJ
cdAYvJ/pCTi+5rJ0n2wDOkgWURcHMdbLHy6tXk1KyBGuLGWuWK3rfPKm4TOXZqChY5LWx2+2DKE7
qm+i6E6JlFCKEF2aOaIr30TsKPBb5+3b/WYJyYd9JefeHZC9edIfo+GqrXA6AxXfLxcUR2owk5sQ
6m0A0jBxN4XMIv0+FDLcBTeX/H+YX8enHnoGFQ/DP4nCNpEdmzFiPBAuuCUX+fBZU0QErX+4mSm0
fyyk5DzOUT7JYxHInlqncemw56cwnKN8TyMT26QU/Xx1+oh8WvpVvWAqPwO10ZN9MGEo9DWDlnnf
0UZdBIUglHNMZ6Nw46vstZg9DYsytbVHLqghYdJBmHBhqNnKuJ/PvGTfFXgW0IBVHoiH/diAMKRz
/QMCLhVF1qEIIbbMty1LCKBvgIjyF9rGRk8KFFEQW3/tzGVy4at0qCCIPwO9RzHlpgThXU2u/IAz
nGFxMgZX5GkZ9nOh1rn+yTRL5CT7SUj4QspXc/EYIvrLLdiJfbVUytQiwowknAklKON2a2+dZA1b
/5nZH3/Vw21Im0aMCp0lzsXm8WRv0dzvgT2GGb6qtPGCz1tGoDmVsn9XcknHjFSEutglp/LQmuts
gjY3ttHxMJkGpZsjo8QqjriyKP5o3WCFyrNhvzKCxzbElQlsTOuQlnhv+BOZ25z9rXq3uaMLqCyz
07Je4lRmOtjcKrwp9xT8FEAV4v0NtXDcobklv8ZUMzUjw88xZmwTBS4QbfVCZjOw237Nj1rX9GiU
2fOlOzeLQcMHSynOGE+vnGGZ4drhG4g0CvKUQgzObUIiTX/kpvuYh7R2o5Z9RiYevSQqKM0bYE2S
+HTWLlEOzgq9sh0Hg19T0k3z0KCCeR91r8LiFmS/kAF7ce9ZQsXwOkGlNMY/nyGyxJ5BSZYgWa0a
oHkhygMob5hI+kziECpyqAZdY2kCZrpszR9uOhFCaLiszohd3+wEc/CNR1daLcpTIUx2LCPoTgN/
RtdUTDtFhKWtBnSBBfy7NZLRXRZgpjoae6dbnqXNAh/toX5vTfTlSKCpO0wKZ/g7JJ0QMvqWeev0
bB+RDHDA4trSil+2VB/mzfv5g3t2MKTtEgqDquK0L1k3d4oD1R1CjvzscaKy7I6S+PFGmkseYT9M
U8y+bsfwzNUAEE0kFcvXQeg3Jb3RFpzN2Bsu+jk5G19+dXuOuaw4zzM1GXd3fm+2pRr2rpz+MPgD
3DImkulZj7Ld6TVovSTkT7lDzJtjOhZMWN5yiehtK4q6O7PUlxlRFCSRVH8QrXihtyH+3GlJ+crf
1x7fwRDhimXov1j8PFg1KtfEFRvqunEoPBdYAv3ImXKq1qU9Swm4S3XqJfdNu3Vxco2UdhQpPJl6
WO+nEztXC3jvyDrkh7qKTerAEuD3GrX2NZLDKNj8cdDbVam8kbCGacBlhQ/tDTYYsZebX5pGZGK0
dhCkdB+sMaWhfrYwY9l8StIPKNtAfJvXPBgYG6p76oxNKlOft3rRu1HKG/GdVbWE5JbCucDCx6kv
qaZehH4sqIZTpFCK0TECcjufGjEtgNfLQdauGP2ofOoKpzFwxBU4PvArdGWhx+bzZHtt+CVcRkoR
gfmE5Fhr1ve9H1vD4tlz8VoPWcSPAW7b5qncC1iCKGp1pEKaeAXmMvnaH+7VZYkDhtBsQ9noovbi
lhS5KOt53uXfRb4mSSlO3RckaXDKi/h2f3qBTMCcq0nfrDUtME7yZQR0/SegUbmVBQKnehI2fPz3
cWRR4x8YwVKgu65+Gay6/67pJS4w/SL36OGK02qx+BJtB9kSIMEl19VJ4lL67KYSeKgj+5hNMKRE
KkCNjU1EaQC9K3Xg80nxyGDhKi4ESvstyS1T7khEGAixCGWk6LiWPB1zcZSdQsgFf3yLs7ANEWlL
3rBfZ3OCP/YKbFdn8CDBoyFr/v4Gwu0hC2aiR+m+nzoynFGDac1oUyFQxUbfV51DT/+Z8wu647cH
Sblfy8eZ+aHUblv3f1sCsYXRQaUXsmAG5jdhp7U1igJlPIH0gklR3QE2jx1JaAP1BKXHBz+nZTOA
s/IqQku3EMZbBqamgG5ITlL7UFilB9DEt7NLKJmvy18EzBVT+8w4tOnQyFOzuXn36fBKMKqDM8zB
pWXmLsR+8YQJDP1+XIoT+lzMAksctuQlRRui/pKjKvwevIAjq96HmCm6gdCA4NucWsKycA1mQ2E+
X2sQwQEHp7MJwne/Q/6L8jjOGEB+Uc2Pwx9y7sxXLP1j1xz+nbcUBb7nxSGkVr7I42S4A8a9+vAy
b/0uxoYOywL3N/+QYPVsdeZOXwzxM5vL9c3yu3OkUDbbw1q5AAqWWiBvOT0jGVZIsoK75ElqfbnL
qDtVqNaRoIn5gbpx4hs0ZML1AGWKP14Fo6fRRtIdpH8h05fiK5GDleJXIGfFVK4V6PNMh4LRewUE
aWaBiSUXbMADO0/lLpvJhPLK/5bGYl7mhdG3AlSrhUnW6vjMCkI9A+gC7hRKCn7lk6jHoOt6u6iT
aQG7eyqmZIvqM91xWepT5RNYViZmOHur28FONs5HYEBOXaxvCybMn5ETdwJRVjFDabSjjd4M8zBS
KoBSYtQCGL2SKZqZ6Vh1NPU7c61cQ6TEBiUhSCnicUl2wvhp5enWJCh4AN5rjR1X3t0jSSq/sUuN
GhhjvOxRGsb2oW5CbzNFVd7B1985/PNQWOc7iFI+3A5t3XJX24eH6jyDMlMP3mf7RLrN2g73kMYr
h90vKqLk04OltdWsFXH4rYPkXgti0ejkPdZ6sIusVzgVe8X7Vhf1vf6SfoESM8P5UMVw5Kv5S1Du
LRmxrIKpF25+VkcNt5tcb4Br1YqwAVsq9ark425yLB6PFTMFkRdOGq7cAjZKT8Q7W5SUEri9aX43
ssgsRUZmCTFh/0TG3AblniVynrBBiWczKJDCO9g/IoZGSy2ZTu+29/W4aC4Is8AQkcW3a5Zgnk3a
N7mMII5DhN/W6e08q9Bdiusd2rxlq24OlO68BB9k50n6l4SqGZdlILXtp9ggnDClU+yDbDO7KRcS
CSwPbFTmMgH9V4T/is2DYCSX4jpiUCCkwWZrE/BqXOPARgy+N3aampU7MwbPkQeuIEo27OC4y5/Z
ZL3H2crBJx+vQ4nhJL0M53dhKLvtlbHAIoJlf+EeUk0457rROhYs7nJQdlmYBNMKRGcfo/Fc4wGP
RvZWm8CSBuyULIuKb6BjuGXEab1rIfc3A57ldMkVrEQR0E50GobKmzLaxoCJ5NDYfjYj8aOiPOQ+
XKuVRc1UBK+ZaxGTyN4EC2UcnQzRcSo7V1JIrDDvwk13+g5pnsjyLu7x2DGzZZaHpLewwu2OOEag
cS2io/GN+eGVNEStet8atdVhXr0sXPkGf+n9PZrt9JLw20EOce9v/T/1tff5FFQgxLyQNIDqzJvs
dcjduzYlqERn/l3TqPcfvCb29EiJxCOyp/XIAFh1V0Cm+6GyDV6wnYbKvixXM/gkL/CLX7Q7Ddl1
73pfANtLzzvrMlWgl25QPXPplT6fUkpksslbgFj/y2qziAZ2jqZDF+1RtEnIlom+JQJDBOUROzIo
DE0U1oPt2NmSg95Ilr56H1pbE00mRcHYBIPASKC5d0+xgL/rX42wpzYaZ3kJx3zg3Elt/RFHiMrQ
+ZZnt9YLGToPDucul1T7MveyjEeC++55UUef8OSrkOwFaUsUhNDMsRHkE88ehTiSe+Jj5hoECYIo
n91UnGi2jFL1zDmlT65WC19cGfqW6YMVrHNiLI4Zv7/+0cbOr6so0q5ni9iS9uhoe2vQPu+lLaD+
raBY1ceYvaPQA6eQ8PtnZRCh7ISjLixQsut6qKI8nyd9Rr8H5OqAd9FnbbLP+jslSafkSDdT6J8b
1lNzbhTeKQUSOQxXTyuZewi7DLf1UKLnkNle61ZfZDJj6x8py11eFR68/SIFfHEhnzTxP03b3UY1
HQJdIWU5s2+ZQx60dgDs3CF19dgEt52UlvbdWPTCnUl49SVbXlM095pa3SB3sLEgctrU9vERnKQs
OQsjCx070DkzA0/dSAE3rxuC6Yq9pSEAEg52QL22xAogcQYT1EyDqs3XeVi9vN/tEFFOEJOsRgI1
TN0vKemsh613OpU7V2lygK9ZOlhMG4e1nRezYAzH6gzq2cnjoxnVs4LNtL0QKRFjQZ4Iq87s468G
/bHqz75EF+WnCeXqYijGrY7rHMAHK6NWXjub7wnqXJobk8tadHBUJcdRYp+igLmzXjjb8r8T2B+B
isqG6cXcvoF809Pqvqt+SvMGiTCQdakh0Ga8qk9L/+BoiGXSb0b1Vv99qHJI5kbF0qfr2H3UJ6Ag
2RF/ULWSFzz7Vmd52ymg4uBbpOsOrPtcjmPPi7GlQXezVXQFyqp8mhv7T/wzhbDh/16n2ygzkb+Y
AOnwlNCfHVUMoklJ1bvYHi32pBrCbLO8JcSy8n/aFKlbovRhHMlM9bgHSe/b1sRM1bVH7ogUNOmO
ZGrKAGYuYCRRvIECt8t+EiyU0dl2FdnqdPGBoNyjshHfO4UeNZ9XbYEoyhYjGlQ7iqpDaFGqU+qa
ZxyJfnItHDO2plv2qxlqRI19nAA24iImc7wIBQqV0+8OVgrE6gTXR4GhXXv53sCjr9MLPB4JTxqS
M55tFhKRqsnFLtf3rQ0vgdmSuaadevcy2fMp66q6TxcQsNFmrhM977KOVQzvPM48bq0dFgEwBgJ3
4liWQ2lmEahcuErVMopOBcX7w4OKh93DJgJkp7yainJSEgQaUJfe21QpWLpIgeXxk1x4VdbA5ca6
jDdm2e0uZsAjfDkEwPwVnGuDVB2518lTu/2DTIP8q3RopMb1qWPJrs3HcpXyyxfEouPz6+ZLvjyi
BY8LkfW0TUhv9zRW2BWJeq9B4chJ2AFKDfx4gYNx8xaDH2fuxhR0j/9mcZCZWljcjFv0kFXfXx9w
Egrk00n8tcKKonemCRXPVHzzV4i2lHzFHSdJlTmmVDO9KDOH80hd7QNqrFqVnsMpnObeern5wMnK
akgRSmbDFE4RyqtK+qxw7UDmtFZyj5VVMsd7fHfkMh6JHI0uyfu4YUpyBBdl22Fhk+ZTVf3Dw7r+
Nc8pMjBqSuc201etwIHBFm+jBEyilecUv2gsBb6HqLsEFpYQS76PV497PEnMUvNAIgBQvKqa9UIX
yazw2RMPFSF9ejxbxX5xvYpTgvwPvq4IiEb1hEeBoZuXqx+OPrd6IQ3wlq4dSF0vBiOlYZZPa51F
53d8VhYvbw6uCZU8uM0nHrctDFEs9fxC4Aicp5xxjeAXBAHwQEVzsGAjFi6m21YEiUZAN9WFC2g7
YoLEGyES1lLoVjRy2Xu00rffjOmJx0HnkvTHocNPJUpl6PHM0nagxH/Qj5guk5UyQ56dPxU42lUA
36a3BdFNhDDPCULqSFxym3e9WEx8uBrotQfWPbRjRI++mJEmnPYEGxJo6K8P+Ay1Q++y2ngyqfrR
BaoNP2w6AzEmB84R84E/01/YWLMD0K1qusPRD1gqTbKWR/m7EXYzT3Lgltd/GkgR3AtP0ZV2QwWS
TI3w34NLTVcRmXA4Ne3WGjr9g9OZsCewgHods35q55oVxlNEYElm+L/8bjYePJblD2S0HxCLtVB0
vL9Y8rfxYPhMcIGbxrT9wQKfAi2e+glyeLi9w5Wa9JWPY+lnN2/Su6t8WwqSHIxEVwNdp6Ipz/48
A51FyiiZVZbOqJYdaeuDT8V5Hx6Phfxc0LcoZROzk6ZyNijBRf4wQk6Ot4nMe1U65SYzHyQNxJuq
isvdG8DneA3biLR3SxS/FKeeew8wJaK7E7b8SSa7MvK3cEfNZoFLALJ5fJT3jfra9iEHA9/jfbCl
gPLvSN/vzfY0sg1XQZcqglKAnBOr3iHgKyPfC5TWaSN6Gt1IcgnVrvHM0H9JCPQrGw9Q2WdMsDBr
3rQAMNTso3KLpWuS2HmD3pfpk0x99TTDN2bKqzt4A1WiP3bYcAhboakx95AZKR0YIBjY4tGz7+hN
MOaESEwFmwEo8dbP7GI975qsRSZl7QMMGkW2dK9mlgymap62qArlGNnOejKd5CR/FFDNoap7qCHS
aHBitjnlxhBbfJQ8HOUFakPhKlmgwsMESaKPse1tT7z2sKClF5ortHYkhukN7KYCliIxWgk2dm0f
T4rzxtcWfZ/G4spxbEhqIVwLGm4ruz96BUBAJ6itYTIXPf07Dbs/CnmFw9iPKyZVPca0qciLLYOf
NO/YxHssMfGSfUSox8Voof8rh17pK7mrYuV7s0xtdBM7vYvorwptXnAUQm0tCydw7w2MqB8gPfEd
88zRgmEOzMZJZjpD6b6Xork8smF0evhMbh8MLAZU2MmAezLjO1Gh7egesIMah7qmd8jqQclNc3RM
3sOX3gaE0/X3rIsrUHWk6sIh6bGJ04TO03O75S2mF3qYEg5N2TPEmk61lqK+ab74d19jelMZElrR
T9UhgILNq1gCvazV9BxrLMPPWtxHeWqTHX0FyaD7rSYrBb/BDfz5lPaDyKzSE13I6DDsP8Q/8oCu
/KoEE7cxJyS7h+hk+ZrszMzAXKchqFXrrkYjkP8vxzLFbEvUPsZzxwk0/JhfgAaaHPcgwGCQ+8+P
gPn2xH2D/Nkwqdr0096vj1h9/wJkLBEbI03g1zCJNtsOaoSyIe4x0PG/wiN6kyZTGClzhhfkcu95
PjXNunkfywXc53rjZfbFBpha29TCxwZxGA+tFn5korG4kHvgePoMD/+wdiRhZURTdQB2GF4svr8+
brM7vR1eGI+Z5fO+CImnInyebS7EQ7HyYN+Dji3NlNcAhZ+twR7ZAJNzy5qk8fDcyjX9WO8icXMf
WoPUCMgTtDCda1TWOcmzqzcUC2cNmIzcXa8PiUvkq1OMkOTvTrUXk2GsboNWRfBYG10YQ0oe7dab
EwhZDZp+13Ws1X8DRBO4DnPNxEK01klt3mD6VvvXhecCvv0oe3lS7Le505JWb1c5jUlYNmG3EAeR
EN2ZTlmotmnwY4bsfPGJLCaUFCAiSQdTPK953IjAQepq74jtgQWfKE7kT9tpxCM6KVPFz879NUbQ
fv12O4/8HdnRttgIxWNX3vrtOIqk8gKe7FN9WKQfJzCSb5EkDYoqOEs2mEC/ijMmlWNUygsGgd7O
vgKNbry63UXeI3MyBtIi1YQv6owkZLEXFsSOdI3D1gwi/RUhy8Jx1rT3UF+v4SKkfHfjlmndms0U
4JEq8hILRPIhvYXBchfg8Y3U1u4Ft0WyiDa9EPpOMB7G+e8m7o9SkPrzzpe/eGfMe+1fU40kzCSO
fRpDJZSDWTK/fmVzxyVdSrNW8ECmloOtV9qK2lcGkIv+CVOXFjI1/Q0AeKQZgw8BdQj4Pf2i2FRU
tsHyMPUXd4PLB1qvCoJLGrAyRiaqBBWDW1ae5546WZWEpRZ8zcM/usXueolssJvoHROsv85JRHbU
I4F3MdRUU8csdeTtCLkdQnG5R3QWpUurlMFjC6tTLB1iwFDQjydWcMbn6Gf/cTk6DL9YzmxKkcuL
xS5/ReElkA1c9qENWmRzL3FYM27xDnbaOlkxLJ0CM3JdI7UVypiVf9iIdrZIUsQwwyUKSRO2gDo4
rUaWyXhwBZV1Cg5ginMr2PEOpi7Z5YNP3/0HLA0HghiZyUNvpK5hoOVF60fwTDKOPRXSWRJkg3RH
j3ReVKAe8SRQFjB2ZMVxpeBX0V+v3mmuK/Bm+VNDUPwTRCvv3qu3P30XnFz2bAaNF6BjKkovmVlb
qOxlZpoEgt5JjDXj4XEMyt6Qwo75IJ3Dxubi4MAjVKXSYHf8fSQL8VrYZNto6xsMuONM252YnCBp
4Gqc14nWVo4Y/xvNv7nttyzDV5ZiT/YEErLsjS1/Avvo2/KcE6qBcbuvfIv1oTBjjlPh+WwN+qoc
Ga1w/Vmf6co6oe0uTEHUBFR1NKLyHHi3YFlRYYsLuyqKhc0h7cnGNhz5nFC9XG8sje277/171dEy
gf69Ya8FD9WEkij4BovjR21KNBppvFy0lgO4zlKvlAkPaGzQAiro9g3UGLMhyURdXMyL2wGdVxmG
qEBKCVVqRVxoRqmxxu1f/KmNV/wCw/yg74+fauolNVwQO3fncO+NkA9PyVsWbtuNjzYVrHaTq/X1
edV3hzj0R0UuZ/ScyVB+XmJ1dAavnRkOvQ9wQDfMkGB9FgUAf9w/onrt+ymevWOmXd31hY+gjr0W
VbZVRw7YwWCoGPGBkF1N30hWpFEJtVwTT0kP0BeXwtiodzUD6B92l/XRij3PJzJs5lTGNUEMgf65
cMrXs6akM/SjPfdffWFr9+EGjrvSkadtfEpWZHZqeID2hzHf7VKWMH4Y27pQXfsHS4eKxF82S3+w
yA003hPOsExUDh/+gjgLvRgrGqXEP5XnCVskvYUj8Kph93f9oAlJApWBG1CrLGBCYiKCjyTVM2ne
8f/6X2fArZERKn4M+sZvf5WqJEWKqngVLROatFoTU/FE3hiEgQv8lyU5v8jYDT5t4p2hUzh8d3qh
przdlAnA57Z8jicQ4o7mUWbu1EvxOk0ljX6n4hmN4w/Va6BFXSbnuAG/WJ9zkXzlHUsprtx+sNGl
nGxhapFWHdmG2Bv3t+rV/DJtNwXqn23eS0gELwFc1AYETgjYMhyfZyhG3vfkppHly5E8FFepD0QE
GjTuLH4wl1/1ISOdjuU2XFUNxFtcrV2LoT+VC5XzPRznWpBSD7V7QRSqzbZW1rHvIatqIcrj0kwq
L6YxZsAjXr3GZsoa/fa0x37qFViuOeoRXjRkw+ef1opMHN3ixKiNAzP7r2zSIkJWu0OLjDi7ToVo
uWhOC9Vhf2MgG0/0wgv4KBkDJMfwWRrCHhE74mQP4WTo16N/eG6MscgN1ulx9JoUP8cBDpOHatG9
OlloioJNTs6F7Bl3FnSKvmfyqQEmJJb3pzyVYmMi3JChg47jpIg2fdd/d0RabxqqbcPuH4nEza5r
fI0PuW+JI68pzbEcu77UmCVmHAOj7lEOIloVe/Imrh3kdGefSGmV5ukCuVcOuWCgbZYeZV7zCFfx
LfQI1UE65zXY47O2QvGipm7RnOT7pXAYr/8M8QHG5tNwyq+XPnrPG9fLM2iTa8gWhYUjOow4IrhA
6AELKOrh6GVaKqtUfXeqzM/KWMDyiAkdNCUfzDZqIvi7JRd6lrrhXZDrcxN9dhGxRKOp9VBIL+FN
Phj1k7iH+aGoVTTOBNOM1uqVEKBd9EdIDngXrCttRMqOHC5e9sZf4p1HiJyqMp9oRmc2t+6h3N7d
AWo0bP8UwL6sIns6KP/QnlNpagBprQ0SuX4+H+8LiwI5c7MJZOIEARVit077BME8FjMKsVVj0hO4
D54AGBmdmOpxoVDYjpBv3M3x2KmPyZ+5Eo/XJaXmnB9J6z00XQQATvqP7A6PxpY341GMlduh9V/C
si/w16sOrp3iTSZRwUeDXuGuxCTvsH5j7ofC5/Ehv5wMZe/VTzaKQoPZe+i1U+r7JNzae3+4taZV
GeiQvpE10oOVyoa3vZHs2hsAFwaxb+UNdMr6b0SIM8oVNmku/8CX1ngVxOdptiAXbizjAoNtAJk8
t9xuTdGNTUhzevS6xAxXrBH13XlCRsR6hs75HzBTrb+ONozZiMR+6qCNnPiorm48rySVt1K3Lfp5
ipRVOHh/nsh28gtecG0OJgyM5Wt0HoGeRkOP/NtCrICmZKs0txaHmdEntwjThpdeluhKL9Mlu05C
Dnd9C/uJbRomS5He1Djvlozj9A0AnSfumzxLuHBTNO3LuKLWY5Yty8n0tURBiXw3tKQ6m8iwMU4U
Cy/cBgp8EqOafHe/DWXmLf0fbocW6usHVIM8u0YGE96QhoFicvWuNDUO2aAsJgBalxzGh9EtbibL
LImT29RqR03s6eyI0lPLF12zWO8Z5X2mq4m8fia/2/mrnTWXQo8nDmRXoYug/oBZKmFy/Kd34m2g
FJ/3fbCQyqpHVUkOll1HsaJZFSOhfd7Ew1VTLchkqlWQf1nDcg1DRN/YOUx8gI9FmBZbuIpV3o7p
Ruhh3dYyIemPhp0ub9wuL1XzsP71SHvjQsX/c9tGkaUHMRmnuQT3+P9PYscmk/ONd41P4wWtimGq
4/A52EN+FY0l7Mz2qCsNCOIGnHFhqYsJKJz4fd4IoJEGe3iObr5TZND+n8SmAb2jJqzlRsZ614c5
YRHHrjPSp1Tzo8QlHWGDy6hmlGvTCSICq9n23RFGpfZ3+Byqaw82C4fwUj9HzFUwyzuom7/IMGri
SDa+lV9lQj6Cw6dKtBtj9SpT+bgdEFoW47aUMClEEdB/HQn2yj4GNMttUAET/Fd/mf6XEZSI5/HU
lKi10oktFkSM5n7Sr3ZESYM4emmAbGN/LpHqivFGvmAbNz9IOROhDf2HpYhJYBFNXAY3sRVew6YR
XEU9ocVUVfjuVrF0e3wia5o/y8zdg1QMGmYw0WLcmKPHaOhYZ0zotEtlSO/MdGo6eXiThIYH/5qS
wnvTu+iQHsUIIfUoCfjCASMim+xC3IChyd2R1o8vInzR1xUmMNgY9cWoY7xswcNSXytGTtmHCrxT
FdPo6ypv92U9LgiD61kw9eq3OjKx0FNKYE3aaW8WFG+P3P9Duu4vi+veMdPe08c6mVdXMpT4+w3A
hpnAtAo04dokhKc3GJ1OgSJ5JzQylVEIcr8xyVB1fWEaJ2QHp2xqz3aqOqlNaZNEViSOdFz+rnIX
kdeGbPBhcHiwR7jkM/MrZM0G5q58ivlEy2r5Im/sXN4kxymlZ/0WogOzSH2RXOolPuzTET6IPZfJ
9W2R9rd/9jcVFJrW/fg7B9EXgS/ADfIIy49iU/5enf4Tt9XxNxeeOezARErqgwEtpIRK+GkmM4Fr
2TuLkEr6DmfmQIw9GuT1tJ66DWkHBC/5VuTOcaIQ2pFAyk0OwxwCmH9GBfFfJTZFs47MZhSrK1Nz
5F37bN8vkPND0gma0iLgr2o3MXfEnz9sNQUJW8ZKCQAQZ2gHZzkljppcplAjiqexC+82u5s95Khk
sKZva3cSI1DjOi+Gic+ZuDGdGJSwGszlr+viHwTjoRRaTM1sjpQj4b01xPTk49iHKiVheLAHhoBt
u51nijAiIHnzIUCHb7VaWmW3nFMvu8U/d/m2KlkPSunyc9EXH3QqzP0l5JXZT76pE1OC99EVt69V
1pUicvIVvsz/tAa8oypx1blT21sHU8h/NeXm2ZVHR9K3q7Ui6WxfORCJjPWAstUvDWws1cII4vDF
Hs4kMZh/3qZy3zoq9bJ/YqeALWjSozm+QJFHdQ+AX5RXf8xxjAUv/MrpiGhU5ehLBv8ahYhI0DSO
5Li628IDmYEbGSUVVLe3CMrsefhsLPPo5myMb4byEcGiygXxfpSz5SmsQKBT2RmA64mYEi7QnaFl
h35hIKwvYqGo+6QLoVfYxrghQGyD+f64uNNdQCKugJgaibWHnn2UU8mJi/uGvXbDzbozPX+GBsc+
w2FPiUK7eQ+3loGZopORl6xHwf/qILWfuOSfmDv7/qF+3mO0CjnbcmBAXeKGCCbs/kt2ihlWGx4k
hbX3YUk/hbg/dEnlNTWEWsZbLVF1C3FfVQM6Fahz2JnYUFefj6rz12Xk/Ylu+TphfBe9p+ktfhZ/
QOadmNOgxSf/5aNCV7ETuxnyjTY93vGCxYHHKTV5uZ9A0DXwQrX75q0CLBX4mR0Q1NqqlT2ZpjC+
H5TDKysUXf4Kc3KaxYMR8dT4GozPw4OTb95oXcQ14b6Y7u55/tAUA3TyRMGcZUxWp8eNiC7L+fym
4UPwQgE0y5xELc/ZxwOJoBOJam32C/XCIie9DhIlX6NE2Dz0kRQt3qSGT+WbM89LRxo4D4tz4VWe
p2dw4+XgN5t/AiyN62zysFYRNTCNUx6+vIXqJ2Ll2ptatvgWA+wt9U87TGo72xdXzXlaxlyoml5k
NfTeJTY83SO8WnBl+HWsXxwGpswvhcFADzJRL+0HvvH/c0NJsmZTqEFY96QEAVAM1eAUb+hGtjH0
y55zBSN3uQXwCtOvUrtTCd9bxUVuAu3TiudBXGyZR/M7+UQrl1Otm3cPuEONrhmQ/iHCu99YcVRZ
JzAzmee486iAD7cb5mx+c7tY4Z73tY+bemnakuF1b1A0ezLsbAoR9C9f/lOIkfK7Cgb6k8Pk6M5A
1aYobzv//qBq8bijketfPP9gOBUquiYfxBVWu8W7Ewj3IXa0ejn3acjkLNaqfH1HWfndSxylz/+X
SYyOMBoO4KogvJ9jnVHOQUEO1jHfhSPQu9Ml59NEFrI+8tr9xUN7XubZE4lv+83wq5VZD6gqcTmk
r7pB8nRIhtYuPMNuC8IQIWQQmhOfUqshHNutEIPjt7sLvuaBAxpoPSz6/wpYhcaBEAaLuKm3uenb
+n4Jmk3vAw2FUQ5fh+mJf+Z7TDGW4AjDiqXNWQWS7v9a2RhC8je+8+4L6oruDNi/tizRADQ5hGjJ
in3TgM0Po75lvbroFy56myzOKNUwvy1QCt2P2IEXPR7YDgVJrTn6mURZyugk/FIAoaEnE7wu166f
y8ieoJRTDA80E5KVaBf8Ja7P1F2D1MDyq3xhEEdvtWnQN/fOtd4NFBlpaP35T90M7hkEb1XIVx97
a/QP6zJ7pO1dsxSwVYMKeRG9dylcFgAN9ZaLzArrpXQ76qOQMyXGK1+z/ECoB9yZIo0fPBg+z/ll
C6zh2T5GUyiBzWRVGsctxEYEQNiapCp24dLimr7og8KsxqOhtg2WXU+PYw0MjJaWlNVvofD1fbHE
wf7ZdkhmFzIu8G8znx60d3L1+N8+p/VLDjpAtUlKYB6OQHSlI3kH25It6kbidNkk3WJZ24tgowy3
otTBnqvk+dM1GQKx9GztHIKjXOg2+AlPljYntLyXjR8GIrB/buQ9lzu604Bml+YmVfDY/CQZYwr0
kMCgsQmYtUovLxRUlkOFCf6kRzgv1pne/ndbb4e5Kq1693+Xh61OR3RmE5EqEYsW2LAIXJ5rX/vp
SMR3k47lRChSsSosRCleD5MM0ETO2iID+ZKSvzYRJvL5EKtqghV1WRk3QeItM717dalJB+Iuey3G
vPALRs001ofeC6XdVcXtB9NB4ASIDMIhLW5qZ5H7KiVjFVPFnjsZqt7jQEDD4EWdlKc/b0joIbT9
Kvn/Um9oN/CBp2kqSWAvQomnk5W4YQdYaB2LtHxstUF/LRLZ2Zg8rI3g1Qo9b8x9xUYNsHslk+sm
1WKl053aKYXtyCmFU4O5g1otMufKG5LxxtGq9+5zXKygczD/pR/KVQbJNhMVMeuj9ODxrsd9lH/0
ow+Az+T1fAjzB5Ca6fYkT2VttVasmyJIaxOvr5jR/ZticbDeN37fWC4GEwi/ruDAsbVI2yjvhGIe
WFHy0BHm0SMsN+lRwI9B3oy52ueMeuSQkPC6XpnLtw36pmTH1YGc7Vc/tilvBWWT5/8JJra3caK9
l1S+Us8THa70CHG+7YD9jo81eskXq+pKbfkde5WkEIvEjLvkqR2WgwfnIO0WAZC3o9WzWHIxK8W0
+vS4Ue3qeUlPQI3nB7gYoShVlad69Hgwyzu23wx7dG1Tasz8c7n9XuV2fJbLFdvabHRUpRp9drcK
885HrIUuOD6LuXdVh1nwjgW/1azYr/E6ipfY3geeZQqeHJyEBz9dPupsjLSXbUImV0N7AF93Cokt
q42MMVe7g002MChnYU3DEGmbkCASviHf6pDOdU1QCofmYG2YiOxfX/dZAwbwwS53xyRl5WJruAJi
e1yNgJ4lFY51J5L50yOV5mxEzJvShdwRYGvOh5Q8KlPmsob/NTu9mo6MVXwwZsqyjl5J6+6ElXRk
2kfQGxmAPh3Db7lg4hfFVaZbi/GsHjoavL5fM0dGJH5mTwC902KXoHHsijEzns0q+NXsMHtOKF1n
KYXxnmjFSVtqg7oR10kP9FPPf23oOOiEGnauBrv9OA1gsyYqvHrUH8twjqXvi76gZ71rRwuDMETY
zh1dqSl9fdiEhYlWELL8tK/7fc+qGgKEFPdL7809s7bI5VFJrjWa7Cz6kRaHWVrk1Z6AaxVYIO1r
oh3cZs0a7tjJgU3G1Rh5Bf+6qTcO8civiTKi1aM9K2j5hVyo+/pINLhpCElazs36S8aaaGVI+z/U
JIjtDQjO5oK942ZaULUrBiOp8+VWNs/wakqavL4ThiEoqjckxSpe1+/8kfbZG7pSzYMz7PAHIiq7
sX/W6FwQycNRa+WxhV9n7LWBKtxFB2dZ6QPOvtRHAvBR3vcZE4N6WSrcKCbsMwlCEOSs8mgJlhSl
1q8mc5tuyo6ZCS3EQjkAtn9bFjybwP+vF+AXYdY8KM0aAbs0zz8b5scShO5EFxHwL9NT/Z8cDB9d
0Qkq1RITD0ijgAxBYWHNzNc8HI6XUL1XxdpBOOlig3tBUKluTD3lX0Fh1ukMAT9OIHH3kna8IaYY
DGbjS2aLLrbxnfynGg7dKjeFOoqR1Fs/tiH7oP5LVLw9s52KdzbzavaqEZEYjexVy2sATaCmom2U
l3bM0scDz3WZnyLOIoN5lSB7Oj7zSG7jSnClwga6kbyL+gZBv/snRc0n6Qqvo5A2Jr8AIoKywURY
FvVbG73pfcsISpkM6StbREjdobGRECejATQSsAt5EZgvUS6FcA3oOP5NwyG9oyQwu2CXiOMMu1dl
K30VbDXHRj9ORzfKQXoB/ihWrUP6bVZkDfw4YNhIHB8rLH02YUC7hZr6OChvQym79k0IG41/UeSa
MZjfRSkmfheyq3tC9ouZzUlwgHxt0DEIRfzL7XlS1REhqx8THbhfd1NQ77ngMhtfiNeLcbUKLCt6
u70IufqYD4zYb8+5rAbgXKVEl4SfoMXq/1ep6dlm/qQEsOPBw18UNJEv5qBKFZb1mFaXJzett0aj
SHELEBp5QVRzzLRpjVqlJji//+lK23/kH1nNjYQKp3l0FcKnKh9Izm9pUGAaU1711MUPAGqgfNHJ
eZLmdOlE+SiPrUh5nH3JEFExuObP0SVzvwWLHXNVftEod6qgOzFI8cWAf9DTGktLNGKuEC0Bs8IC
kZMD9/iiquu9CmNr7HYX4P1NOsEKmEAU9V0nxNRwKz8OJZlVHL2l2KcdCM9L6qR5TkTZj/rIV5yc
JQKWNRy0bmZShp1e4F/CZ2xS9CSEXnSbwO/GYc26vflY9vL8nGNGxg6tkPN9/v+hf2RtpH06MKlJ
0w+kk/Lg8QrHcx4jW6lT0EPXaPVoqet1W7Asqn1OOVUQk2JalS2lOt12++rQ3DTKvIpB0wREVlov
qWEjlzkXi+Ev6hwtGOTTldyXKUJJrZM3JttWavU8s2MtoqNEOYte20DQp6c0K7N37nzoYaKBvS7C
mwwyNPXzgX8Z+Iy6lGw3Xxur8aRl2+r3cKkv4d+QOQstc5dSuFg9GsiMiA4GKHhFXcE8Ouh60vPu
Z8jj7dDybc/7dKFeMyGjGPKnE9gVlhi7FhyD3mc5mBzADbN4nYC5zpT6FQO3ZTxnRgZvr7H3aAM1
8QeCo0xcskiI4HR8gpcNLpXLvtoc/W+tUCMUlyIzRoQ+0as/1HRFQQ+mt/RMcU9A2DFKB0ffF22D
+smPBXinEQA1zgIw6GdLCVK/YtOaDBuKNmQ7scx1FgWTxlFuMgHzfzIA6PLtj56HDYILjO+OcxtE
YjH7alyks3MhUn+btgEn8JVCazXx9q/8u6ApI8cBeUNVXABcm5Ca5I/8gwWd/M7fY4GZ79iqn3zp
ybJi0o+llsP25uTidokvSq6IQxH76Cq6ZYx5lNkqTjEdZTjZmYRYlYx5SA34zWP0MRX4NSF/6PB4
fX9mQZ3CZQjLehsT/ohwm1Jc0EA7V8Ovv+IIEJn+eki5IQ8lltrwyfnuEi5sfTYPZFsj+OVbQ0Y1
89PUuMhCjPwJ668HgNl9xIkiMSCI0lIVTZZaIdnpkuIrA06wkcB1nO4tGm3WId1v9bPZPFHbSnkG
Z1Jdg3v+8d3GLAuXn+DfC0Kv/pm30xf9nvG3Z+nykEHvRaOKwVZ8/AfL3vtXYkQnnqDheCjPU7xc
z/O7zQLklDXyO4QxyU87S7/7EPtuMi2BhgamXPooLU81xoz21L+qQfJetUZKOSc8WhXssZxSgzwP
+gYSgVX0GkQqJNB3Zo/X1SZS+Hb3za6Ol9gYxlZRDIoHjV/aWLUSKD/bN4VUYyscbhjB41nLrxUc
96UY+VmkzrRSgikYsZAQf7+zDvUx1sa5P0ikr3VAvUuCN2ka1ud2Vxvj6vezmtE4P6j6ldadxa8h
McWxTeyURbxSfrCSSCivylXRMWAd/jm+R6mZRZFJAac67jh0l5t1yPljWKF2Qtpypx/by+qdU0b+
nW6j23h+sKwCTAb/JobeguylHczLJHN/qHx5o4N93qmO8mf8HB1cfBtw9X9+MPDsxMzbxVUOQ8Un
i3IalQoTbmZeru9IR5F4RDHHCMTSrnDQ6O9ZNpV7N9D1Y4PkvyJZXRZqBhPVmuBpE7NqWi/cRuJo
Xfw+M+Pke/2DbHP9WFyQVhcHqENa9CRJ21rW7Sl0+X/VY1Fzk/STojX6yBiVoIoC4UagSDxc/X98
u0/6Fp1R96WdaWGNOE7GrCCPLPt5o8jhI6rszleFnAKdYtiV0/RlK1KStW6RiEMLb1YFYjr20hXZ
RmxM/RQ21FtD6QcNXHTU5I7c479Lz1TuNNmdIMQdXR4NRt43wT++ftT4BuyhJqcGZhQx93+ulMv+
VI++pguRE7hpBmg4BADsYBrM3RK4bKBYv+Nk1zZiPMeNKgzO4oJKtZBVkr4bJ6UN3TSNsZenpiHn
Lcz1Ut/D4fQ1J4iujiNYzXhDY4fCbsdXzdRC7oUybQWuPU7X5chbLetGVwqceneBwFyLPCSUYI9h
q4zeX0rxmOwl2pE/OZ8t0f/8Za7/VMbX8VZWPmAUD24GWFvcEDIG0DTMauQ3ZQuGPXk11MRn3OYe
Uk7XlDuLqhUCRSfqWbVdDbnUy25FmRs+2YZa9I33XVV90gxHjfYzPdkmuhyUPMcp7je1lcrb3BLp
hNN3NlbY8zlRAvzYw/KYBecDbN2mZbTu9VNa4/Dq3P2uz/jmqVH0FA0mLdOunM2yi8gK6L5Pl2SD
V50+jA42euJhp/e9m0cRf6Slm0aMNFoA46quEee9Lwv4ALg/UdwLC8Ut4izV0XnfXTghfsEzIlul
JCbxKGSF58hZ6vL2yh2NnKD7KqD8v1kXOyY+/hecfEntx6CuZ8tlMWaFsXsY38tgiTuflgiyOb1R
JWISHcrPuzKsEOuWMRqjkg71z6sm3D3hlgDuRSOAS99MKM4k4uhPwioMJEK6Oq02dogOtrlufXOq
cPRwwp0DeffchyW7bZXICTaI+qXh0FA4erpBtz/QwOjOjpVcPhrp9txMw+7sWzEgMwMVfADTvoot
z4T+XHFBADA7Z96hMZFzgrip7SGOlLVw7aNRZov8SLbI4+nK+hmPLnIm2+b/r5M5mUmLwh6J9hn0
kcV81s3x/VWdGgoQhcFitYZS0RSzGFfptAxUHoWDkrjtqPp7r+zXEHCicVidvdObfdBSbmhDEM0A
AT0BLHesIXrOSIJF2EHRfaTlx2WsuGJen/tr6L0u/fu7RWglkv6qHPWbopkzLk3NtFVUhbFhNVwh
XYk3ro2avbK8fRaHYNaL5B6mQsAL5lC/zH9fCKQh3Exxce16z8nsLy7tabuqT7OZttLdHS+Y/Lh2
27WKV9RVzhZsDq+yyjEmxCIRJ/xeOQNe03O6F3nWkSoxYRSm0FzhnOrTq/zznj6HMlWbp6dExGc/
HFgOATQWDJGF7m/ICZ1C8OVtvqsldKTdu0oE34T00PE7n9tR7/EH47sDjQEoxL4zLmfNsxE09ceN
t72q+gVQ7txzn0D6pbUAAjXHZdYLmQQSYBxNuc9BGEoLi5SqSCvCnnBdCh70qXkVtyEfpAA7lu9h
eZD5D7lXpGGhBY+uu009mfejOA4CY3D+1REMuLZfwrs13bW+pW7cDrEHmIKxQPCFcddA3bcY1vj1
91JgXzhfMAFiUj/V7OVPPID2JJT/TVh142INQBKNEsajo95CIXKgwjbXA/Qea68fxq6n7X53wC0g
c6Deyi3okGJWomWRuNbXAl7Lj8LxhiYInNEfzduYvQep2S6h405JrEfUHjDfVW16siKFZxuyaWnN
z45KE6JBuVNeCExoa+ZItbuXEITBeK+nDNx49/bHLCIj07n1q6yvh+p1AYzdqOmqUOiuJXdLnoo/
ll/EKZ8o4L/mY/Ki09qQQDdb5Mj8jukXokY3IVWra0Fhp8F0RRsZEddyVngHwOmwVTBioWYT7x7D
ITg1HzLTwynodYZezuE247H90uxktCBme3lGAK328cSuYS4HyrDfOGWJJMTWx/xPgauval9d42y6
XILA2s7i2hcBYCbnH1MyYksqP12VlVeYbmIqPsx8bPX3MjNaRquKDCWGrdXEw7/r8rjiyI7oCwcL
I+5g52NQ43fUlffGq5XgzCIXZh6rLqRiAHmLYMSZ1Z4t67h+b4AljjGuC2jJTHjAD2mhvPRDXSm+
iuGUIApC4RZ6zyQtt2/ut5aBSvVFIc7BNXmTErkDkA5QrBjhShNIXKKiFB4MbSa9p5nyjG3+ZYBw
bW5nytgbrZpbaQejnf3xZXmDS/XWPY+kJiPYnrzJVsAlAQC91UGC5PqDS3FtJUYCcJL7gqStlpcf
o5hYaB4jcL5dl9VTQzMCAE6iLEwXrZCxC+2TMXrV+pVe5q4tsfOfFJ13uJZcwcUyybROXoA6AjnT
+UgwLICujXihdDOXseVZH4+9jK0oHEs5drVgOUaclwV+FMqgQqZUjbuNJvR1QqPDH4Pi99pGMw9G
vAwupie+cDcen1m/8Y1FoABzb56wGnRS2oeEc6N9+eltX8kkZqMpUFRRyLuw6TVeDxqZzXSqG+OV
cPw50ytK0iu1MJIXN+nn9K/Pb8KXgdPDl8naJq5oS219i2o9mB9O72yOROB9mL1zE1m0sQtoM6OA
eNmJM3JrSfPQxpndBXHQDfOk2bSOM/uBqRr216sp84lylMYCh8BtwYYzHRuhBmjIUdbuVP6duC78
l16hiXQzymAvTtxqOcZzd2mSZJtj9/wG4/CeHojo44i2/Ia7nSKloclObngu0f9zNZoIEM4l6W0y
hn7AoEXT3/a0lWln+nAXL/mPHJk/zRQe4sNb2soixmNBysuCD1gjJEWOoLLnxf45fFlBvvrCUtKs
cogn2MfER1AlaNDqaJMb4AWFe0V8dOyRkvRfQZwMUChOpUTq8CB67Ym3IF9RDmmMH3TLGUIJSiRL
RdiGdUdqY7XCDJDaZzH0uVShy2/m8qGhC/pvoPOrIj1NQpJeeP9U3tNDzMP7FtWWm8DT7xTRPKZY
FbEhVPF2ZrBR5YJIGxjCMSXa7QsmSzYle/+Hjse4WVO4pNhxw37BKz+wWqrgknPphIBrOHNgb0sW
j6i8A2wO37UtZd2PpIHW/odQiwWFWmMeWz7W2ejclmRKgn9RlEcmc2hD5UI4WmM1T//Mf3QpHXJw
i/jpcUvQMtmr1Vl/vQhKXa0XnH7CyM74X6gWfgfESeKbBc5kyeOscE8Wi/kwvp7abFsZtvQ9MChr
Np0qngSbc1vcaQi4Dey0L1OMlVmzG0AznYl+6SZ4q/a0mXjNWjvPpX6dCRPSjD0EJDn0gQ/9XeTm
cp5lC9dNwgIPs5MakPZwXULFt21syVGQiPo7SnSXrnVZZ0RXlzKox/JYFMIaQ1GDfem99ypTmcBj
2YiPZ7qliCNcN5n8IgdZ+A+iojIFLTrGCOF09sn7Y/+0dNloEE81J6QnUrLq5190EJWBbPmhpkEm
YECFYhKl4hVmBiiMhc+mKXU6ZYJuxdCDWF+gYQcVS1QWGSlSYGTALhe3F7/utv7lrd/VeIy5xXdh
ZnNilxsBs6yRivU0PaiTEcT/BALXa4zOSGODyncRxxuTHFjTmk2BPFPFFMmUknhv2G9kSwOvMEvH
E5855MLKPMxyF2KNi06rFl2xgxTR/dgiCplxDNl+rOCYDXLSU+Xp26piP/kLrrMpReQC4Sj8zv4U
r4MlgmXZaVpADGa6q9tJ5saHAsiZ1/rprKE00V24nB6bXv602MrQx+9azAJvLWrxpDAKWP1XlC7E
y/pRqcR71sVQrewnCk2f7lKWihvGQzxi2nowhY9sdcO3ENOCtZYR+/w9CngKIthkoCmtVwttOh77
ZrUImaq3icV9scRBzYvhG/lEgkvEjGltckxjOcSEztXrPJEvelceq339TLkY68lL5TFAm81pdJSQ
tPXSQqrx4yF/kAunJIojGJbYUYtWtw/dOaxvhmv0WSCIuUWLIW136twxA+llyx8OlPUZukDzPZms
Xm7w0z628PCdsr879iqK/I2DAI9Z4Xc4Rn2mZ+45ZlffN0Mc9IJbehJVhS/nkHXrgNRR4av/FQPJ
Wi7AcV841xQCXXE7Fu6dFCHKF9m275Po9b0TBp0ItiKtSJoG58HA21iqa8t+vxFNd3FwMId3nhnw
uxkvJ9XI3Uqm1osOUtVhm71AQYMukrEAtro8BLdMjNtRSZo2kr2OAUIeER39V03Zs/FOdXa+36KI
bbzJ82B0OjOg2e5j1+bzkkn7GYDESiSu6dRBXm3Oz1DiDbC0U+PaaWD6GvnzEPilL5i0Dz1W5XXv
ZKpjCJNpWbiT/V9g1pT+wsnGKQ2fFoMwFxJo+lNdoI6+hgAuI6je8rBJmMv5E8lfMuG5mA56kQbo
/relBXI3FFS+Xjr2VXqBMaJWjHBpX53LKwOwdwt8VJT/09EVrXK2lV4uJEusZy6ZSHZHCvrvL7hs
88WICEyIdvkq+4cs0qiRP8cNY6AF/CjpOln51e9zEEWpS+JzwRGDVH3s7mdeN+TXjH7asAC6xSaW
qVIaroNLEJbaIN3bIbnfQVTpbq5o93050YOIO7Azb6hnuY4t//xpRb45RpZvrzJX67ugvdiIe8vo
E5XqLjXK6OSC83RkhMN859PCUUo2cAW6wNJd8yFkoYYijdNBsswZX/oqGPY4ofZscuQQIyctILyp
7GiwXx5pMs26mDalI3MjITtY4z7qZO2rGZn49umNNlwlwZXFH0hkLSBhlMfvfOtRsBA06/MoPOf8
q5UkmJAKiKDKKzfxmoeQfOGU3vNebEZyCaiTUfLX+Da9QhupVtwhiSXHEUqSpW5hxLYYBjJxxiS0
iA1mSpC35A7vscWsk+Gj7GEBM4wR/GUQr8nQhk5UwPFH4lfI9HZ2x83p36TNBJBQ6R1uKRhytw/W
/GgVxx8Cqfg+tJzl7g3MVPLr2Un2AK7wxlnXX4XnXntSNSyUcSunL7CBQ5X/026g5Km+59m+SPCG
u8KFF9/APlwV8Itc39ykBhAZzP7GMwfgglipCvZcZ1Aws3jxzR8lswRJByc2DZIO1zlD7Iz3IEj3
3k5jqZIastM2eBmXJQJ52ntWDT5xtAvRgiKIGpPkwvT/6CSAAjwkGzj8+vQT24u0CxppkOsPQ9e7
rWMuOYh9sDroyUnN6ZCh374HuUp6tAeLQyLOOhLq1/0T4oRtKe/syK+UpgQ2I3X1N367HWMtH8/o
dGoJm9+3MfJ5bJOGzrAJD8Jf4P5rJ7+yR2vTXmfR3J0Z3jPhGFosBIM8Qy4tNGkfuItb9Ig3/3L2
ZgaDcEYcuXRVa0Nqfo5kUJ9DHdyEFwNxW/zGbe1rei1hcthqsWvh0o+eh6XPt9Lv+/VHNMs1+usN
KHx1hb49g+fwJdau/QebVGKIDUkTc/8TxLoGy+GGdpROX61jI8QSePo2rHE6RB1wlKFUBC27xwfn
rGjKKekkNCingUe4tF94Y9UQ5MXxd+/V7aGazbE5rxMNCI/aanr22UgE+z8sht8sSl+rz20k0jPi
lHFcZunsgxZrOgUuKJA4NwN6rDAqxHc/FxBm6/XlGhAR0TZNZ2HkA6swzANe4FOT2yWyfFiwXEi7
tQGw2/GkLJABOkK1Fn4q/OnMyrzbIS3OQDwZgEok1rQ/Bvnkf6KIaFq4QV/ELrLbNzbl/t2jJPVc
RhiaPMBHE127o/Q8C2j1xhWQDIY6HHL2RHpCg7PIMZAQr5JA1wlUcT9BwjZ1NeAfdKgKCviMnEDL
Q7O70PfjD+cbvAqu6X1McBVg3JMYKtRHSbaprrZ1AkYcu22aLyzVsF/6AywCMZB4mHHN43egbe9X
n1FsMJpU8K9wyyAiJpe7PcIC8wqjdoCRxTiqzgJeEPSP9saOxQOJY2V8bKRrzNS5N9IMpQawfSP4
p7OF+BkyrTjkex3HOYkgLWvQWjxq3oL5jO7Cou7afDLe09p7ejAkkk6lyUrEe0AvvuQJrBXAAlQ4
xlFczsrYImU/HRjd6bJhxtiC+ymI1TZDl2gE6Mq8jB86XpN/bR0+I14HgqMcmCOOoibbPVmiaW0l
ryg0+LMZrqSD4xUF7L91B6IqCYlIx9JAfWlUl3EVAROhKLIJCCBefuVr+oDcJZrOeyzAdcr5l7bu
W2tU2y2oFHmdyzIQ4+UpS65ZbSkNq4Jd9xS9ex+xEUhXrxGMlrOugmp04BqWLQMbmI5tKDM1awso
2cn0lMWzG6CHQ6VcaXypzRma9e8WLcbOGkniMVy6Z0+bHp8IENzcNjiGaFE92XXfLXU2eSsm+Cpl
abtOCv3ukAuLkyRdkywCJIiC4JlbljC0MrG0HJuSiHp14Tx/Y7h9rUVeplYwIgxZHJiCMA/knx9Q
xO5ITHK1SadEmfkGOVS7zacfzyuy7HBpXnOFcIUzdBgkE1s9uarcSpdXx91F7LwmPIEi97UIKuyx
KrrOJ53/NhqZIaGu3U4Dhhbic487dJTmKX/fBMup03hVjy1VGeUl+WJPYzI4qBSBou5gTY4aeva8
ZbwbuB/bl8V+2FudHZREYWdUrSNVUQLu31/zCu3kXFX1ZsApc6Ke4ZKQcjVLr3PeWohQP3SwAYMI
Gdlz6rcSjTuc8es+Tobh9gWQs6nDzfQ7fL47ck/4jgJSkbrV5v60sHnWjPsWm0qAMl8BGHe4mvNd
crKz73sQFkntNUuCsxWavG3gqamOJuvH3FXcg4oJCTobj/Xb0aspXQVhYGFe7p5HUhXKXZ0QPBxk
WPz2Uq4kE9/tfVKWa6/L2Jmfma6GvnXlorbF5d4UelNwbSw3IZvTDTiRZmO0Y29haCVNJHZRrnLx
JVGeNMFdmIzXXSVwcR1PzAmarwrvr+ornB9XRzJONv0krlUPjxwCWhrX6BUhlbUIq3Y6y1qeDWrV
1qEcmoEUwCcQV4/JnGBXOrTkkzJ2TDCk4heOrsoaFIqIqa5ac5p6rZzHb2cs5JRjYEtjM62uDLcI
1pRh+va6qW1p+eOryq5VGtQRND2wZ2c/FnlHUBnISM+WGaDpUmMAIQql/uySle3yUudtogHLngxO
JJhXTZsNtmRaErIHV75CAT8rZVKF/7FKhC8obyGL3V6f+FG+hbsaC527RkpxFwJe1RkFySpP8iz9
exj6k22eMlNUvgIf2+jzxfu7Vr/5g3V4PiSCwA+k6jnuVnw0X9hOlrAFtG27sg4IoPID0oLFZLBJ
8yxAkrVf49N+6ZfzdbOSv65dpw1DGS6t3sN4AXWhp3EmcMvVE4hs9/CZ0G6g1w+GZXqUHw3NWiYV
O+9MGyRit5UdezPa1L8YG7+8z/IhViCvCRP0uUYEQcUMHpZD26CgtAkMzaVQqP0BySup4sluQy3k
8ylw34TEOKF7EbCoAMqy+3YLssE5UUkIv/ojXUPNtqrlnDsfjsO3UVHxT/QK8JODJRGOrw+p0A5N
93fcJMe9KOeQziIvkdS3Y7eTJD8PMW4T+Gre3JdxC3TDgrYQbdkl3nJqP6FpBoMrVCXetIG8ZL3H
9t5yUVgxRgPPKpgMuOGLdsv1yuS626oRRi4sGf6Tb1G1K07wlxilG5DChnsTivBvi6UNJ/eTk1fO
5oTq4+/N28SLXfLcw0w/EnxJ4RSXM2VXtKeFdmZjPFCFpyaJ+FVZPQh+o5fBjzUTIcbojlgmW9px
y9KhL+kyyI15SPV+NgyJyLrJDlR3mPvr2LOdQO6S3VUPJ4qd1xY/TwYud9/Bor4Z4Bu8sjJdttSr
YXCs+ETjQrYUx3yb0HiV3wdEkgJONPKzRk3Djk7OBpXlBgn0IeFfq+A7gNhHT4HQDdd6DYE2lJwo
o1F81fD/qHDDPytk4Cg4JYB+fNCCMQG95h3oXmPJnrurYP6QGfHzMYfwFUskGa7WZtEilaEOiri0
awvmLsrLYlDJ4Q4Is80pv8hlaxvFAUPinNoEVk94MSx7h+batNXh1+cG6L1olqFlSZ/1baX5gI0R
7KBTOTSb88AHqaPHt+N0wI8lu3kvFH60ymw8uUzWYzNXmX2ENB+nrHeo/ApdWmPSrNM8jjrkDRzQ
Zog9htZOAKWrZY34qU6JgVQywllWlSyWoU15CWbvbFYdXwQY/HTeU5Ogi5uwBA48KiRM6A32+PRF
ucUGAcV9wooXqF+Kbp39skDF1W7QJycip9Z6xvWF6s1XZbhrulNIzdAXi6+FeXG+k7FU3qZ5P1NR
113+SkZc1zyWe2ePaLyYjhuqThhP3to01UIBdUe+k2Py2PxQBbANvA0xex69EVWPYDIPRTTTNS2k
SLw8ZIg+/BcvXqjILG1c6HAn+ayi9sl2oaAFxt58aXtjxw5jd3ctulJ2KDX5z980EH4NzuILsrE2
Uo09M73tpOvJPtZB9ZheKs3yU7YrRRuksYoAbRA0aRtCdA3el/VqPNwanc6stKvdz6NkOMAYjNSp
4NyNGZopWMtFE4AXIRKMTuyFgfPfkeRb47nhTW14VMq4uHhNslxmNQcR70pi7KJQOzY720kD81cJ
0NTpmmelGnDkSXCqcfrdYlQVRrkYoufx/j4RkAIO4r7Jf6JFP0UtTnNk7MPaVtlEAXfYKkGQfXO4
kmlCglkw4H26rOBQQsxbRSiu1Y1YmUhBE3EUAUKrmYgF++KoeoARU6oi/xoca1yGEN+RblrMdFY4
sPbJRpRXUIpKybJT9EsQj+B6UE8bEOB/cP9RO45ocylUQE6SvalOPkAmGX0m7lLLDTGnwUBRPiQW
Szq8NPGV4Lx7jgCQVQ8j+CXa0lifRew0b+KHsc7/GpjIiivZkgdIItHvLvGrDq+wR+RGRAOfitgm
WufSJIalfxvsXqpyEQExg+CkXyhNtCtwPevdvjJFuYHpVpUuO7EfZOCHW5wb6g/nYsyRx0PByCiG
HSLr0bW6LpnXfPFmfY303o63DyfD4mKCOOt8pybcCaVIGiOCGzUqW96MamCJZgJaJ22b1chnPTbR
iNDIEz2/+43o6nCbkiliIInWbsl5Nd4M7/2daGrqK2PfY5eGmgGiBj4NmWRud56sq5IeLMD0ExVW
94WHBTElvYYbmw+NZiW8Q3huvNYxpsPNNHo1jLq0GJ8+wuPbObCob64lBeU5qI9/ox/VNuec1kaC
zKBlka4Fwsbu3onr3E0lg9/LIp0yA7XeE81la6CogRVKMfouicIsV6tL9tU0w6M8wEs5eXtDmJ3z
AK+e5BLgwe10G+3k3YirAfD7yOn2vFS8bQ2jUaSt7AL8Z2BBrduGPDpskKHIjOGIul206fSECXEV
MIBnjSx8Jxw0CxcmjScGBOKKdgOhxZCxoQK9IgIjPXbYL0BU3IHH3KkFHUgInrVGvX8jEjdpfKXF
7SL/TTb2JXHG3WhqV8fwI3c8zlB99qy2xldWzTQVA4bVlgH1fx12VFeD9duq6K7oBq2yOMbfwZKB
SkHjh4DPccisbEDfXNWr7rh6XvFbr16tag0YX4xWl01GCRwK2WFb++cjtNtfDSEoeJR874X/Hr80
TCDrDugvpikDOy7F28Ky+ES7A7yI59zQZA1k4Jj8scLaC5l+hs4r+Q5aJrYni6gTLlNsc+F/C4fz
lkxD4rHk+5RO4YiBUvcpVqaQz8mMlG5kBsdbDH5+YWLxEyVuXachr/0rV9m4K+dz8JRPYdG2ijRD
ddwyycm9ybBVtk1XEiUNIVMoZDOkJgIKaCys/9rKyUnFWPNWlatHyULyYPne+qgJDJ35jonz0+8Q
OVlDkjvB2zyV+OU/FKoELvqXQZn0OENrYl3jZsKnsu592ewOqfmXJf0khmg81Iguv1ChuHqD7RZQ
CST+EA9dXTRWuE2ApzkzC5KwqnJAL8+pPHRELz+aYOSzoPscIAEUp6LD2linLmc6HyKdwdOdYgmX
FN9fmh8pVCCRoB1Wi4jg0Qbln9yco353wUdBE3jU8QlqmrJSct/CD8JxRj3MbMpTd7sPNSK+hzMM
bnWNXxsv7TqkKd7AdhpQyAQGBk+2dG/uhpOqCYu5lhnaewBoicsa+wL7s/qUtdNXd4k2HKOsluWt
dqo3OfmZ5TD+fbktTKquBnw+wqORLxMTIWk4V1/TtpaXLemYXsU3Aoj4hL5L/MuVEfZsbnovHEtt
/7IQ3cOvTzx31glOJVn9a2FrGeMNQWMM371dmRSiFaRm0XrQGV8/+THJIk1+BR8eZBsL1ZrCddT6
t7lQRxsB8RMhBiFmu3ffbOpmeEYK5+fpgHP+FJo2FdHC1zmN0bPkGZEzofo4uokTNmr/oi9FLF+Y
DyX9Q2jAtmxUspmuC0VcapsiGYi74Xqq2ofMVvFnbV1LkP3kGXSYsxoGXiDfmb1Y3BNiUMkJOUY3
1CzssVHAxnZ+5kP2QtOSsHAkI+QE3JILY6UYTmAdrvEzzYJKjbrokF3iXW9a9icTnglQx2d38GSV
toB4NvnGNcJRO8qtuLiwRMbnr7r+3Fe+YydmOxydwTyzpbQOK5jcTbiGQzVrmNaODTaSyW4MP1tV
SC4IXE4Ara7IWbB2/eLGR+4Pxi1tJwsAEdpeEW/caMA7vAXPBRI6sjOl65/vvWj66UsoBUpimIGT
V0JD/DtY/TeHLqSSFQjBcfbXthCq7VCUA6ZjZCGU82AeM8p9F8VnsvH1/Ib0FUB/QPnjiCmwhb1Z
ruEi8YrRgN7arvqGnToauOIhXamA/ZGGycTrLWhTKhoNJCZwuhjF+IChkCN/zVLyXo+T2JPebEmJ
ArsXVCEKgIvRP9ofiNdQELLaXwtHljs1q6ZeGD8+SCZPT5JDrFLCBRATIfI7Qp+pDRol3q4rNBOw
HPUhhtyC3rT7aKmy/TsMbmTimqhQi1ynsNaNVfKMY5mZVVTSjqjhBCYmDB/tyu/HBIMbSHLs/8xE
jATcuSwjwpCCQ0zhBWUXUt+WcH1lYqG1yHzeGnU7VUKN6FWkzrL/Eyj4uhJi5VF90f1wDHQRxDff
Cas3L462aYpIyYwmL4SvfMrFyt/qFkJW9DR5/D3CMcfMaysSnB5FY2jMHZGT8FOJssI48fA6lLbK
v8jtvZ75b4MbeTH3WJrfI/AlawjZ/PiR9nQ+i1xkyyDqYKax3gsL8x4wz4SBqtFq346XZbdkh+gV
xVRWPKU1EftlEivgGce3QTgrdPg97ayNSSCTQ3GyCUdU7vR1I2kom0151kfwH7YZkcG+6PXRpEC3
Af/DJO0x63vS8REgERsQlU0tlJOXkGeFgDAUhvwAQMXFPAeTukJNLxjpS4bhmSH2UnuSFjL7IFar
2ltJxKjzGCPjOFt1PEtAfZFw2UjXrwouQAhsF2Fqvjgt6e/0xOTbkc+/rnnGQiAJjQlwfflKJ8/N
I/5Gz3FIMSbeVltkHcLfRI0nI1DpaQ1QiM/5ZRRcDzwt0vhPN69RGFTS9hY8Thhlv5JGIpSYTYRE
h85TX1TCz7FKLMKdQaK94GoRkW1Ztoa1k4CMrwaDBUNvo77ZCymir0cUMSSMT8wcWoPzWescHLyz
QzHYXxLsrCcNsouMo0suZQXEh8TZL5BtyaPtwk8ZWO8BUDkArlq8hNiVx+oKAzQXQ2EDS6xTInA9
TRq/qH4LDJthgEdvKxhSNG4439ZMkiqR5lt0BEOAEinmUzqtyRGlEmJiPpq4n+HPN6/6CeZ1s4Tt
ezsgE4W9EhQvkge76nApWlNZnhNT5YgPjy3U3JrtIyL4dBPyGIzfZ+05PNxPP43ptsNRCIEpC5I2
1khX67sU8GK2/lFDIzEz6Yh6L2BtQ5fuSYti+WjAPTXVqavOioLnaX6nLZdI33aXTQ7eThOvBMnv
nFCZEZGhkZezzXxVo4rD3t4hhPXcYkzX6fxtcDZIEVnumyvwQA7LXjztDvTW6jv/XAuc3cuKqaUE
QqkPAiXhCvl/37fQzEXwypelReyyqsewZwaTRgIKfFpdJrLvAdY+AXAXkN0BVGbTHmIW5xuspEBM
XoE6pTxekW776ZM2O10A0tYojjt2ALqfgIOhGhCpElGCfy6kvt8lGAfSsUyiaS0aQL+BvH8iBHTA
nRVeQOG6A+cJTaq3LvKQgZi2pQgj+h8l5df6FpKQUpplH3F9QL6twx49nEe7zCMLacPrgZeYl+DK
hBMvM85MI0joOAYIGrU0igFIxJ9NhLiTuWmaxrP8djsmzSdpTYIwWJAA4+bUBHwGWe4ZlFRXWZbI
6SL5p6M+77+R8JBwBEh2zLUfZMVyUYU9MjPmPw9ZYMT2Y+woz+QeBd8EcH11ZMjSTWVHv0bjmvLY
zrJpjUIy8D35xt6io1uOPm87K6vEz4u1BHRkAzh1ZWzHevuZaKph2Kre69w+tCzE5KVSXEtEDeQM
+l63CRHV93uayn9o/sV3f5FucCktfePHQVpfnQi5/YfcskzWRNmmgcCYVreuG/Wvgz2KJXBSau9l
tBDlSJ7y02T8I7YkzAjw+Gayvai0YHaVORo4gVeg6Vvw17r6Tp5OB3nOEWgKkhY3yQb9fN1YwoIS
MBVw/xAtUuUb+eV7SrNdaljSKueJ8bkd735TpCINjVrQdEleCnMQpU7bCAONkLiCmI5X/hOYLdGa
wg00jjTzZjmT2q89tX1UjfL/kZKnuZjMKkJyMqgZmN+uWXl2NkZ5JiyCsW1QmacECBXzzOweaDO3
MESdyYejdsUdEqne1wESpCIYRO9BJvug4sJXXuwLt/oxx7QGHuIbVQlubsZOhnoUlyNDQoRXrgm8
Xkfjaw170nKyXGIEuvJKMwQ5kbvIcjAlCfDn6HcWlFolSWSj3ihN7DJJhGHTZ5OHFCSDbwOsGmjS
4pt7nKWI+tlVxBnoDLNCBlwYfLeQWx3gZ4Z8Dn27PsHVsoIb6Ki/9KpdVMhO1/LlYezokslfDlWg
xsOU7RtBU+Y7v/qYQqTrcjy0jmScq+jRAFffRg932MyUj20ipXe9SJZgRCC8DcFKbPHrt0fM/0Yo
scc86BPzAWOfh5FdyeOljSGYNPxB+hQ+G1fMDTmdtzt9a0APU685iwsmSLa72kj6vDNN6xA4j6pl
cuDdOlLl1g7BOtkZKd2mBRNnPtS+nuBhZg697hspsUW0hqr1q6rFV9pIteLaWKwqKHRY15lB9mPt
XArTRiLONRM80mIsBbbSO5/eoGkp3WHI0xrYpP0reEhU08+k1ruli0WtkNw9OfarYRgl3KxcqSQE
I21Tk7YRHDfWSuFIO0HdfSc/ZK/RxRJ/DwD/p8z56im09KYQnSBGXe3AohuSINOLxioNOhetH6ih
wg6D7T9PeEFIO8uGFIMoCPTN4AHtTSJp0el7evRh8+Nf8CDqkzb8OoxxxT7er7zv1s1EgiUMup7B
vTBOMB/WZqJccdunTdOilKAu1Q9DwIbkKq5cPiKpQO9rIOD5LO2hXLaFi7cxX5Ce4jiy4YdbWlE/
e/s6EclDNxkDq+unkb6wSzynfigixrixFz4yfP3XSTyWI5NQUBucgLm6A2y/YrkCKrWjCPfw34w4
wp79zc3blTLy0G7z5+6HTphc5wa4PuF0GgUxEzzQOYk6VVaoaQ89/p1mmN+WtR1+giUiTpYAtjjx
My7/sWltAOPbkXGIKEX6fpB0ark0WPqEsqQAdQS0PiH9F5QfDaY7GuHbY7MFL8pXSvCA5qDaKFzA
0HLuQDP1kmaewVW8Fz+vVdcK7Z2eDWAEiXDHPEApZNn0et7ujFjVzOvRaeOpoayHcKuhznFKfqU4
3qs5SadtVliR37cXk35E0LD35DEt4X/oNNVRfZiCzj+ue3IWxIoLVWclMar+rzYn6GnraBtIMILK
yTHTVztvDN4NNMg7S17h6n+swxGE9+2GR7ntP9x/40TtWzthCcs/DX/cYm7ytyFOQXV1kH8L49F+
/v4EZ5OiQesEWmMWrMtjz0chDVmxyIR+8x0M+Tnjt3Q7kTxRGlDcM4pUI9weUqiuufJudK89L3XX
4Ya9XwuixsustOM4fJGSVq6CKxES4CXp2KuCwdoE2yt4VxvMTzFIlJOrwef+4GDJnJu23OFb7frU
CxHBtmCnsagSrILh+aJ/iXg5kP3omtON++/fQUCBYGtXY8qrC8dxROkfPb2MW0+yYEyPxdOo28ch
Q+d56QvFl5mKEZaGhwJN0tTSTs2bwUnWA9jqnnpaeX33W5/iQYFrhmlnRy3dY59zwEaZEzFzyj3e
2ZRIjMS9durwK44C1GqIIy06njXl/KvYWLs1pMHmn58Y+kMjkK/2FUUEsDbIsfJhepiiOCA2XVqs
hwpc2ZyNqZ7TTEEN1TanWETk+XXbtPqPwFC1l/PsOPdecY0LDMPon5bBKS8ty7L/L0xiq99/ylhN
g7uEKTKo54P0KqfE4alAJ8LtdfcnSJvy+VWQb8WJ6+HVcVDbMKoqS/BWxzwvV11iK47Ya44+7aCK
GrbPlmOj521hQx7TXdoNyECFkbhztE6r/o9EbCmGuUIp4ubnkvBGo2XKtC4xzZQ2HVSw+fzt2Feq
lIw+k6VUG0sjMhLrUzeigXZRBsUtjbeS9mG951jT50scgPsOtTktFWB+OWCk9c3uIXV7F//EZVM+
WrfRe5Ba2+vOybwshLrmqPj84WR2YdIOuwOxxMnoya7/H35L139pxI18xy5V+CH2WGdTuVu4seSm
SEwkQUsQm/pMRWc4fkPwfp/inijjHTh0Isbgz7OC+nTxioNAqIwq0BhGoipEb4mMtNY0khlkZdl6
klP8OVaFi86rRkOcTDhwvLINK1igK5UZUlCrpQNLODK8N9epAEEyRmEBeNwl0K6wScVf9vMDb6hh
j7qpceo4dv4Cdjsbe3LHTHRmmYzS/Dpk1KkbxNzkbMwfsxj85zO+YIsrPjMdVhjqG42q30kHwii8
43as4xhu1ZUSXBTlYOvwBTE8tttqOMCc8jIZTyuu+4NKkWwE13DmNuNQbfP4jqUfB1YJDM6BhoAg
JWUNxQdVYIjP16dIQcUEcwHH2yAImxI4j5WRuFLJgCZP+kej8Z0GU8Zbzrp+kFaGEcvGUGY0NF74
q1Rsk5S1JQWjq8pfiVVLWTMolswhQAVxx+gP+NqQ8sAzH0abn9M+wuLpmw++GEK42vdBaLIt3U1T
W0Ooen9PV5CMNEiKrjWNaSc7yLyGxxXllMWiwaFWnRLeBNfaJXgUX5vZxwjNuLfOwVpeR8jSxUoR
BpM0IcbXDLnvU9vPKwyJ0rFSBfW1lOWx0JIrvw7QoJf9NGzxnRzGsOB1fbfZU2QaaPxPvbYkorbz
ROUrYLJ86KuqlC++KAu2YdZ1fTe/RGUJapnpPq8w5BIuSFhz9Q3E5vr+6QXrAdYczQpHW8UP2jEG
pR0MwDuefbN/mQuRq4F/uIk7i9BQT2YC0Nf4ruu9IB3IXaXI/PUAco10bt1bt/Gnp+XapHfnS5Ze
km74Fm9MOqSx+vAtvBrUodeoOVPREjaMuriCaPRg8DQXXp6Bgxi2SOYfgE/mazySDhCCAfn85/he
pCAc2ljhESljfpJCoDE6LOk6FcbI7NIM4d0Pwgfm210x9mRg83kdP+HSwbP4WWvOGvipgU22kpnz
Tg9UslPJVkz96GB7+vZT1JraWo0kFwZYJiJD9AgjDKqzwegNIYyF0XuMsunEUdEUkGbfG7ODgFOK
CK60OH7JjUa3o7R/YwQOmWpu3GN4lgPbbWeUz7BCZOVy5xR/8e1Gia3fE0t0HbYJMGygEhDZ1TIR
VIYQ8vlq9fGZon2LufpaOmuB9vgw8lXBvURZzZDOheEaiRCTH9DvDwgAKA0NB7nl1bFM5h4mG93+
8Rdg5bAkLmf7b6c+KhQlMLIZatE4jpKz6abOD6f5EGBhMNRiJHktT4USUqx/g9HAA55nXg6K/hhs
H4BuhjKj2FDjqcOKnkTAp7EKDtfCgIX0SNNN6FqHhdNQShTllXXZKa3KXhef8QznUv2xXi+bJ3EV
wFqlUc/pX51NgDN6bYdX6hiXM1RbUasRaKOLU2u4dKZ1KopW3B+YP0A1tMQakpTGAfvFgCs7y/5f
0MtkLtgaooxDyH3QQdPkyCk73QfaApiTmNzJUgLAmlcWi7i4r+uF0LPkJvnXsVJ8K7fAAq4jEDkU
QM1tfaKdX9q/475IMyFF2TPoGMNFLLBeMXVcRLdAv3chnpqNa8hI+jpJXBQMvuxK/YpIfK7sljsJ
UZoPpSJtH3MZevfQFXfU+g+2L4jd8UoPpknciUP1LTlVdnIpP7G2iwsQ19w3gFpLWfqaqZaX9YgL
q2KZ7ew4P0mUyIn7vPylAryFRM78nZfezwX42ckCI2FMKjNLLrmCK3hVw1XkRsQSMfDYSfqKGRs+
znoWrcDwM4TWaSEsbDWNR79z9jK5lXAbdyIabcidSiUaXCfxZGsNYo990zApA+GgIP/bdJl5E1uA
YQ4XXURYspCJAEP9gvi0JFLX/IzsWBqAeN5/4h14GylMQ/x1xgJzpxrl1yJC5wdZgDdh4FbfbnIE
DzR4/QUUIgI7W/kWslA6oEX+YHBIkXpTKwca1Vx1UgOp6Ga8i8hmWdkLLq2MlZAUS0ZEKonrLX0/
AfWm9HBry6K0N5tTzSIHNVX7hB+W6UJ2gX2Gzv+cpfG/PhOrFASHguT3mheXWPPA1Eh3q6aaWdfV
+KWBiKN9JA6hcXrHn/g2ys0kkcihGIR6l3yt9BrGaDI2ho00cylJKlheyZxwFiCpeKPVdzrZ/ejH
uU0faevmu3I0jb1ZsUdZgYsD4GVR39CKkvjwahDCgqSkZ5z2TKjQgc51gIRsS7b81sxJ4wgsO6NK
angIxhh5gpDTGSNvTQ7nudrGuHW+62/ndmMgX/awSapYn0Bjul/tICCYTkg5WnAxLnK1TI6Rw0AS
vVJgjRuWRMwrZMixu1YRgVhXL1xlNfAUeiiDwM/8wouLnocjA85/wC2MD40M7VwUtflTSA9leAbd
yLJl1rRqUKbqOPClZoHV/+a2gE0WM1TG5dCCtXhGSHU46bTbVhC9LWLwoBSSQ+cRq/KGOiyvoSOw
2YMl65EemxkOp1g+ZZngxdU4uEF/pBhCzHWPZ2wT4ZsrAa+bmGPFxxVfKQONXuox0MSy2Xr5q6HB
pnrb4OhD55oHi6XlVmUwmiHW0dvybBbhm9/uVJc3H0vCOvUjx0lfNUcmzvJy/u4fawejIQDRQ9JT
+uMXHsW3hy6ebpbVel2ypvLp7wAY5eArZz278ALkLniZan/lInxvLzYxzsmCA6R4ZbsDjAuowW9E
lTLzVfdQ6/JPI7BdYACs/oA4lEoGOsJSdLk6R0ZmUzz6dNCMBbmRDN//w6/ikEjh5r1m1qLK9MD8
FqaI4cqOhFzraNbFE+EzB2K55/hfSUXM208tWurp82tFCyvXi/T/4sxPLzQ+j3tFpTYyoEFZtTJ0
VpWzLmIl2+cvqtFpp/zEde/CFbPu9kLZ0cOy2OC6a8LIC8cMRi2oThq8/yVibMOigAG23YVLVfLg
9CnJWptVPx/i3yOx68KKEOZWksY968F8PMMCyQQxHUCNETzvR6ZBSxyBvMpUiS2FvDgw2m6hihVu
CP28g/7T5+iG5uUZaOi4QobHalwIG1m15YZTZP4/yiyPFw9wxHTHFhrJ2+ZHwh+cGWfn0y7Yp5J0
7bokcGPKjy5rJhpxdJG8AWDf0EOZS4HKB4THSCEOKbdT/DWyUrOwbmjnHqBrpofJGQsO49n3mBNC
n9kkfZJa4IwFqV4DLAIL5+4aLOqorIBCoYMprvgODXJt68FquPCmdFQftY0UWTEwcZyiI3dyCgdU
iRbY8x/j3OElmIPj10OgzA5SJclf8FP2sOPfLtRyRldIJhwmKtEzVtUNU/XxcSIrhYmpio1W7Lyi
HAY34kD9Gim33kEzcBFlOnW7o/GcrRdgalCarrozTSsNoCAod6YfpYy0KV2EJvP3qlNnrv6uRH4Z
UKx34iLbc+Y0cTw2TcVbkYfaW0rYA9ieHbsUUuas47KkPwPRgcOC5hS5nSvcR5HCzq2lsNq6u/1q
XdPSoYYkhvMTTRBm2Z+AT2+2Ls9RTyq1+loXrdwkcLX1e/9XjjkOme4nbrZ482RuzSosjaKR6Ris
LKT/GcBXD+jWySITVsRmcuDlS6meg1L3Dv5Dsouwp53J+IBYBvkJ4oZbi457yizhv75MkXA9pnoF
TR1/iNGMnDbIUe+um7bYcY3SOotCa+NeRDvIXHR9SjRexAKPHux0wHg2Rz2+UUKsrdUBtcts0S3o
XZEy2WR7H4s9kE4eiHc1OPfNJnuchW7ci2mc6vWNwB3muQokkRIrKYhNE462YMZjvtnIlHPcOtu1
iElPNCc9xd/hRcuw/tWSiNoKMW/XgIRFfh32ZV1akvhK0HY3iqnesNjkRgVQtdcwqqQQH0NznAYU
96FF+hZH9464q9+5epbFa8XNA6ZY/VLozhvV7bNZyxC/guJSCXJVqPa1nUiz0HeTPqvlEoRJh63l
YBmH76SRVlwuZAGmLCgdH8kmTgF9Jr7Prm+cQNX4j6TyCHdy5Ln3ae/ZUr8AJ5fHafGBXPDI8dJr
qzzlb+P++kLZas1ZEamVRLqiJI/iuD7MVYNN3YYXv0CRvl22jip7SodVzUlLpvFE2MmCassJTsfr
ItqKyr2dNjfXPdQkcXKFI4o6gV1Rbs8sdu249rX7su++ULhqvs93K2Jd/IJchJjTtcxM8R0Adihi
rvquMXNpwEYWwkzq8seUIhgdGoPNMYZnmXcQsMRY1lraKQxh8cInupwNQpoXJyeGNZSWkw0bhkjV
fGUDX3mO9yC1JJ8ehQvMSALlOlgdD8h6GPS/kPiBul2tP0APrr/GVhx3UWdFadIAehNur3mG47ar
cEJ+4xC9V/x2uxP2JfsyVxEKq6M9cnOslPLFg+v9ky2iCxR0ao8mMYQTaVuErMCQLkkSwD7A5GRx
rDLyW1i/eKwn8l4bipl480rOFn6mYoMpyTghBNf4J2qoJw9KMaHrF5Zfr/okmVmq5NzPO0iBSR/u
ehFs4szMw1G+Y8kCnmDuvo3M3pS+CoCp+Q1dl2Avo43jHgLE5/GF2YI9fCNlztuqw9t662vHT4si
3LHPPwx/r+MlOXaT6R8TyNcK5cyJ1iAXe71HMnzxTGgX8yIET9evnczbaaE4j3RsENng18aGe7ZY
7r/h6P4WRv0CfCVurTP3vbt0OO1Zpo/dYnbDfZ9Ad9m2tllYMKFY47FvwzVFMF4m8Z3OFLd10EIu
0aSVj2Z5HJJhJH66YCD2MwNDOSZ9Bc4D7PCD25WpUn5598w4smn4WygtfGol93KAOhnkd/qwq3G7
BSuE0BOzkwqH2PaWOvayVV4Fgg86fpfUroqSzTCN50Fh9h4PbybUJMThAgg6jcsgl/fSDgY65Ahr
Z5HX6TCJuxprKTDmYbZpy0U/xDAmGyAkNMSWlZ0NfpA9vm6YGBvpxhLaP2QBp+zff1b0YJH/pCyY
Uy6t0Fm7YCzgvWlDWKnUk1aUqArS2pl+PK1jjqWMD2ntUI731XAlFCl4mg9vmeVZnPZnC0Eo0wKr
mEEenhz2T7Bf+Z1TLGoF/D4ze/Hb2C6x4MvJ/jbYJqAVx7aUP4cB5wnoKQeOAzXeYeeX/8MQluNv
s5X+3bNwGW0fKzsPpWPK9hUN3QXGoMd+h92n2yywT4J9pta9aADMRkrJ0Ngen9NmYRywzqVnd/Fj
kp4O2njiHkzNCp0wAobN0XBVN89I39BG5BRasq94YZPUZKqnbnYmEWpIJ6yC1XDGSVsoB3rA4YFM
qO0lVCrMzkiszI1P+/HhF03PzbWntW1M3WBy5ouxUY04rjMD7xRYF0zNg+dQxzRT1A/H6R5emqvM
zP1pFWt1y8iDNJbJXlAkDnAlPem/4XrUiKLdNIcNhio+vBfamcYwZiYJ8mF5WediOO//f2plfohQ
+r3UCKCY564bqO18nRe5Xqz4UhhGTj2YoVqax973tV4AydvnYwQ5KTQmTKtlURCAEhI2+etmI7r6
JC55BMgC7qTodSjhdlzFqkpCeAyFQeBzuS2E2otN4VP7Sgad2ru8D7Np7dqEdcUOfcUsfDn5lwp5
JKnLkXBQjAdaSzWYw/Fw4fwAZN4C5RIM8wq9rlcZbMvmSynY5tyCf+2mUtM4kKkErln1+ySz1rU9
GEmHG+/ydR+NyPdXnWzPASTmUmOedDcULDGoXYL/crLA+PYQYqEM42OYgGl5fdW+m49Obr3zbOuN
oStXyju4E6ScYWwoSyTbBbzyGm7aYMhfMFCO1PVp9oU4bdtrg1vhmqgV+cKT16OZyeb1vLAxqUzy
yds1Dnc8nyLiMz1tFgw+TWnUXVe25uTHCnNGVyLVt6nfVtwHmvUuh5p+uEu86UIm/o2wG8Wp+X3B
RAbrn2frdbXT+BrAKXzQ6PDUZh/e4wBhyWPnZQ2DlWBu9oenE8QhnGYkZ3i3aXoCmqWj0tvkO5yw
Al9S02DBVAoN6fYyEgMEoQB+Mp/v5CFu66+D/y3w2rRg7nhwLllczrwzM12rENOD8qKjWQVK8tm6
Wd1JwoaZi46jdvvX1X6K7qAP3LmG1vk/ACYpDI/ffb00m7ZFHCabHB5nJrLme1j19aFscuuHgnLY
xskArfgsjlPjE0eBkyk1YEkYQD/d1FJyimXZeAwWU2exxODMFxx+JbSYJOnts37rHqnoyWQOJMfu
Ad/Pd63Mkhot14cg9FdmopMaXLazv4NxjjxTkGpsStQ04PucnninievDpfZz0COvi1fwwxOjxyWw
O79qNgyQBlx17kQ3umPkitDoZGF6Gf13tHV7EZimFTTKVciX2byKyrDy6/eQ1YltYKBV1+kcQrsf
YdNsOyWTsHqQgObTLwWrTQNF6BxKeLexj8gn/g8gz5g2duk+z/3acQnyEuulsDH2wtI/sbJ7WYqd
oQrFCiVaP2CNrpDc40jQmGFC5GUpUxzr6WcwXMtGYubPNsKFU7QStnahw6nOF3R7CWeA1E5rP9R2
ECXDY1TAAYkXLzy1ZUEq86OjSMCbhtabZjZAf2HDJ4Tssd7ReV3CKdtni4dZXNk3z/nw3o3OfH0z
mxMN+nN2ZEQMNVi0bT/PINT3mhMsRe5SdOqFpGTaoyu44PYZ8rdHrBmH2OZ32j8rW4gUO+QybKHl
P2CFT7J1XYTsv8U2cfOtg0UDotwzrVUw/dS7yf44HY7G73HFN2BDxaK2BGvVrs+qwjzEnTS2w0I/
EWbuQcCnBFgAJw+uGVK+w9jIiRVTQjPbhTGjprVHDIEMSjReNLVCMiAQRVb/UsHMchzah/EQv1tp
3QrM0zemNYl08ERnj8NQwHCk5dg2a1E1LzCGC1hP01V1Iu9O1Qvh+hkxYFxy5r+QZsfAC3Y9OLcs
GJEGHICiqk3ISwZGuMo1zWrFngZBkgfSLd0Bb0fE2oUqMpEvHs8za+iL9xLwWjzap1wLAx98JS9X
9/SImkEvtvpL/1o31rejP430TEUZWrr/hHWpDNZTWj8lOIX4TZZ3oee202xErHcOTGrkoOzRWawT
uszTZ7Hu/pjiyOHJ1tB8WXL+mFwy+FMcmtL2gqwSriYIVeFGq9gl/RKwVVspQygNcWkaaBwWWs6F
UeHnX/ukdZ8FieBATpOL8yDcPhQ2O9YsGj+sM/vo+tW6pP9INORjRLeoeg7ixBGm10U6ThSt7D9f
nv0LRR2ezecOCWr94dcKbLWpbMFGsZc7/50ULnRYWBHC45YDU9k6OWut1n7yG+hTi4Vtmkh/Ptqm
v7AO9cNQgpKuMf+MYvcw+9ySOxI+Zz9dxUhAPSOD5HE0EeJp+6gxGuFUpdXpItLSs43zPcO3CB0V
B+Gdbdmag0WTVBVmg7iHmLJF911W3nVNrFI1Hprszm0uu1a+9bD9laA3sRLFS0cPllLcizP5XaoE
vou2f+v9Ig5ZxGTqvrDie/r1EaNbctUflVTAV7OSo56LLoEFJfDbET166CEkZ1KZcMa1KJHDTVOe
dA8+6n3c2LBfOT/fdLQ4eYXoUygxSZB6ZMiQ1+ZPRq3raGVqbtepMm2GBFbAdmcfCpNrvzyElHiu
ZZU66EmbYNInKstAZoD+SjJzTUHfQzDbLUCt/5Q5pyPTVVdLEVPbfEGlNe/iyih1AktaBkCO3llI
3EPOZA6b3QDJqfOMOjpdu3Rh15MxEXTEaJYTsr4gRMKGVPQlWtn8JB19KLI/aw2JSvO1usuyKj1v
va4bQRHbpncYYvpggZIwuZkdp+GlCTmEZLjFNseE99erqn6y0vHrth4eVsZj5Zo+PEYusoDHy7Zq
2ViEh1GHnxT8J/p6JkL42LREJHQkJAzJ4xXx4jJYxBSZRWb8p6/ZeLY+PPpM5mfbTEOH8AbY/db2
A3HlwtPW+OJwef4ridzPaBBTQ0TX8lZ7FewOaVC3+1+tHOVE+dMGsVrDi3nfR9XRjlARBE3o2gq3
DNVPq42SaDlRdOsJBV8PjfOIjEw9hVWO87V0P7i+jNjgdQ/e5N1MjQqdaS65aBB6z9+0BgMmu4cW
Kq/5WsjSWSk1+ugKTc1vMraM48H6b+Qgv9+FKDXzFKx7+tRFnDednsh0sdJj/gBTXtxroZGVIszu
CMlTfFgNYKlcnpSd9fYgSes0ICd0/B10CgOvQoU5qFLHocazbukLtYg8A7Pf3dMKEn9lRB9j87hP
9EFdhL1vuqq/+eWDMSPGJ1rhwAZX8Eppl3NqgRBxamEIr7qFR9vKxStyiCKk1F2QmLgvkVK94UYg
iiVu98HAaaoFlIwcjq92WRDmlGtbnnKCygoVZMfOC+rWyVuszHtQJIRpiFuwLyXQ9up2y82gV6Rv
e4OxH6erB+kLFiGW0THyvr/ak1rbQSuUIKIPHfAR16SYzUGwCpfpPJ9u8LqBGAC6L8aNeqPtKvUQ
NxJ01yp+2LaAnVRA+utCn6Ky7ug88VJodREX7umFrIu0C03j+cxp5MLCUn3fXoXZV0oexIT+7805
Ff+5fv9HSnr3FrorxjBvwwPVcuIh0SHto8+AQsonYjib3DE+E5ph39zaOQr8Me28U6whSKBI+Hq1
GDi762UHrGI3TuJ2imL912AVM/d9znDls7GWlymhNLtMucl5xqyUrzFIYO25ToXZLFDcp5xIUBaE
gZaixT+IoljB2bCErKW4fSsVFvAA6k5AjDMvRCQhtuFA9uR1s8VKyhsf+A0ZzYCyLU59vXHvxnZo
pWf9ZeZ8xhNvIyO/FxfsALe6FmeMzRdPh2GzzNSy4CX4zSM6FvIleZag8vgkVSrsvU0XzRNIU0ZK
LoAzU0R1tVEN9JTpZC70wpRI+8NxdchUkrNhW1DnBtBBWTt6A0wzdI2NKwpKNPnprcRaRSNBdi7o
89du6gkhVQqnevBY8Tzu8Wq6arafJ/1J3euho/RonXF/9DLSN9y3ovvYLRNlKKqRYLvnz07IqXkm
Ooz+NDLxSLXckVY4vFHjA2P5XsvX5VeeWHtS8MCM7kEY+8bnRsllkJDoKMw5ust/hKVUHJLZr3XF
yB5sixOPpIoB/pFqFcPKoQksvTNzoR51vv+02Ormfh2KdsDHI3r5/pRkXkhiGCefx5f2ufLIkFR2
A7YIOihaWmz1kJMmxGtGcc1xjnbZVw1per+F5DdVA09TIoJ5yUtaEpg0K5czMLZ9XA+etAnCfI3k
zjv27Ndd3pdAd0UE4ZDvNU53l2mmqE6bRfcLZ7e64+9/9IJ0SKVmfmtQjpgnbPQUASZoff9xaKFA
zYolfY1j3FQXnlOxCqJj6fWstkGXSvVGHjh/nNLwrG5WWEBBOJi2D5njSygY+7uqcGCwg3RUBRUM
ocqbOVtuRR5AC/Cu/EQxIjCLfdRpUwXhkzCKA7kiQf25Yfc1eSUWsTHkEjWBbMaB2zillXx2E0Rk
AaM2wvgdoPCUKiIisKqilFnpwhOVaLFOLSU8AG89I8SfRWo2wCQOSd+QXz26mDKbTfK7ay+1arme
05Bqkv6mT1HM1RTUH8mMFlr5kn/sslHDeN1qR8LtJnXdjQziw6yAb4WYvXak+gPXNPYDW/HXwzhl
jV0Ba2O9ONum9SJLYUGvCaF7gAmQqjfbU6CqDpdwM4XqyNQ5tjzeN3Hutnzk7zcUWZyuS8Mpdg/j
F1+YqCFXZXffVputf7kLnQy35V09RLNb53cbIl3lLGd2PZM5d6bXOS5Co+LVOb87FyJWdB6NVqIx
7/b1B8cn1OJAwA7LoOtruzPisIVz16dQEHIRO6iPMwbHJBiyDE4pgLYKXrSC86NPuFQ8v9W8gj0t
NFSeW2vdL4nJqaC+Gyi8xBTIg+bW/FnFyn/c+ZwWWP7i/4wi/RAaLvn0lEHM6t749K/Rz5oVLDS9
VJ6k+m9lKOePdnsJecHZSYCXCUBIY0yE7G3W+xg1FUFeEt3sinA8rdWz9z5Q/nwHydgDpRTAf4kx
KxfwBvMiBfX8wj2whJOy3Yr64etoYieUKrqeGr8Zs7r333GL/rug05P9MDmx9PI1skZ8KLxqOHOH
SXky3sJCwfvX5asEHjx+pygIlcpd4+2RyGAkjIvtC2TI2SG7U5bFVhBQTUXo0PylI9NqhP7NtVtX
tKLjZUQZtMAdSuw8uzSD3JXfDXaQXsblQDC88eIdfrNrNOEz3jw3Ww5EmFBR6g/8rp7feLZlepDw
YBRi5eQlnSVqWzlzqy1RrODIEiyVVbEt9FMYUjosIUOcWlezftYCAmRT+eJYQC6hpkjmHUTRbAQB
5BXhFOu71E9h575zWdIUJA33kck+6wILlZ2rjYGKkC+Vi7WG8soJe0ecuMrF9vhUILOo1+Uhgohh
ghpuYfRP1OHKxjn559X/xxx17TsIqSmHSVamNs8/zzUgoc0F+CKOehm9w81eliseVO/2qjc89OXJ
EcBjg+U52ZRnJ/wvwNYbhAGJEo4/0N7HflKANhbcW/UD31i0js3S2j/YwPA3s8I18JtQMtTiRm8A
CzpYbCHuOPH/M2aMm25b0awdhGIkaxtQrXmxxJ1EkuniWmCMtb30kGMtTgEPzNSEcHRmQlqvRRpR
O+SZ70/PXojaAWbzsiVHzH7ct+92W40epHf0/trgq0xoJ+vglfTIoGKG1c7zdjopTukRr/5w2rIn
KlHPZUXehGAokl4hbbLAA/g+Qp0mD5GjEh9Dn2fJeWjD5h8pAXU2uuaT1lcQD+0N8Z2v9e/9RcYV
wqiPoVRqK6Fy0n4oWF2qncvRGamQHZdltN7rD/ddxItj8tCuB2Zl/LasW6HdlGkT78FutAc+YxMG
QwYr7w6yQfdfU9+Cr8S3+BuMFzigV96rmgOEemRmdBbrnOe7wvkALqmYSTch5vzpLyXTKhukGrS3
pkLnTpjpIrGMSigCdS1ExTwr8UbBWSpEe4DtjNYJVC5iysD/z3w/6kWvn3c7hx1gzgDjNIkxleeh
m6UFSxi+DAn8PaRIEPkHV2WrQr8dzq8H/FfeEEbGeHd6jSXVPNC2X/3abj03ID3UODhPnYDYyaKi
W6X8uvlGZ6vUwqWTMN5fledm1OnUNhwYzFhmP7oKL7SeERB7LXKVHQqqK1BA7ZX1ZqclghXrWYax
glKl9MIlIpQIml6R0Ghi71O+2W4Q9GFmZKu/icNQGS3Z4q+86IwHya72+nqHXNUr7k83Z533Gyhi
yVDiUz9xIH/A8xnretsWBn/q73C677AUp4Q41p7mVxpLSU0Yx2AMZYF/0A1ZxhxL1GVo7IUYfEOI
sPUnSRvrVt2cG4cFD5Uq5i/N5/V78uMshNFe5FedFHAZ+SZ1Puq/+DUnNi4/MGuZg3A/w4CXZvLl
IdFGnO/DnZxUSnuESIUNVPOPlIA3ABy6vII0EZUOxGQn+ZlFNjK8wJq5eLlMbwQ6On+VOr/R5kot
m3B+YBsUvw+TJhxCMNv8XtZ3vRhUo5JGIJ3XnGOdOLlLdlY6Q+fAfHC1dRuSEqq/75wC/JK2wXN+
Yyp5hBWw3DbdMyLVdjJLhSWM8XBZvsfgukuDUbwtHQWLX5XUhbDrmXdtX63SvtjSHt9x5oY2vq/n
AwK1gkTSQ9w5pzLeN/ytsIix45WrnAR4NScUyrvloNMWQZWCsbu1TE1b/Ck0C/OMNjssV9HFDoXg
iAbES15VkrTK3uu5+fjMAklIz7N0GGFPT+OPkWK5tINg9kTFh/aAKxHnYPYGumXzs5evvrVFTqcW
DSd/pIq12E0/qb6OjIqJ0uOk5OPOQOSs7LhhZw2nAuzezrzKErIRg19AF/NfSn6FvLzTC5zvP+Jn
goZraaOCjy5qSjRgX3M1Vw7df6abORTRlojKpDF+FgTUgcIxG4XZqvVyLMvJxiYZhWNjEhrbjOy7
X31Qu9QO848XF9clzXNOpgrt2eUsP85UJAS2BgotInuLmHE7En9A/x/YpII1Jghh0pgHStXvRAo/
naQ9RIIhoL0qMBxMCqCitIAWGH/8xpqMlDkvNN66b5YroI/crupiDWrGyEW57kvnf/vofLwjlmYH
E7da+cqQGU/bTg3nbZapCIBC+Tl3YeGxj7L7DiD5+ysry93Qlr4e2lDwCBDIZnvj5lN+D7iI5cSg
14Cu7yLko3BJDTNOhirwcDEE0cP9OJNDlZei6bFkr2R8IvDBK0FeTRxgNkGPvnyWVOY8GBU9dNnR
/BKW6Vt0yewh6SDmly/4kSxVwpEfu5EdGmt4pPK7bWUknNqC43Wlw7O3yCQ57Lih2hNz1pgtVMHU
4Kwf8mtaYEp+o7uWv9BoRGkkPQQ0Psr6rtXDFdXODBxh57m5ick86TGmrPURyfW/52tBLciPgTDC
gVeYbVjDgsCgpxU93UuBtVXmxXnRj+AH5A6/AtbHejfuMeMCldEfSmzPGCsTYx+XSjuGwUJFS1F0
5mRjTdpjniaiauEKCeAdZBiiP1PnYHtOnQBhm4wXO4akQ81iLsQU3yvmMuh8NNZs4+NvARGnme/x
8AsH39h7Qa7rtwb/rt9vSDHVNyfOYoYeqhSFoVU1S1L172kRGJaRbAYNAiTjMN9i5VMba2C+g/u6
A/hxkTvVydX/r2QdK7WVVbBft0PKMRRhGYVaU7vP4Z831rr2CLtUsVxPxB0qcJoOE1EOqsOuDR2g
Dt1lmZzWLGPEZr6440DwO6ILspABPLhZ5rsXBCNdIeaZ7qQtFO4IqQ5wnVNgAgTaWY6T6MyI0Yti
7uYbdjJ5PDIqgjFKkO0zhjyv/rSO0RNoZaCscXfPTj4OmMPchxGeW4WRq/+XKmUYzsu2KSC6GcMD
MY23rArRvuLwX9rnPaTmHWJL2GtAJb3yPP8NW+Dkakz4yeQvwOD6qF01vq8lwVkjw1Z6T89ni91p
R/hnnicBD3MmgGehy99oyy6oky0SBvp8yuo6e+x/4uKl1453wiucIQvaFZ3gtrzfvbiTVa+kfIrF
YaG5+pmqNK1GUoTkVOC9G7ZFdty08Gqdr8wl/fER6xxzvoCvYh3ush7mQb4xpOa2S0qGqPBr0pjk
oiJN3CsWS6UX5XuophmBeDuGCdTMBlCR7q+TbNVDm9fziVCEGjo7JPsQKw71QL2KUAbC8mfxk+Yu
2zWsmFvu7WTxdf43bBlMXUI0vzzONQBLlIH9hC3R0C2yxMDwLtyDxzio9tAEK49gp3c64Q20sejd
eg8re04so038w2sk3w8c9l1U/9UCvyU3x2BYheHO8svrK/exAGWvme6i8P0896gj3n0hRPznN2NF
6Nu7EWhfQfXE0zTEkH2j8xXhzmLHVN9SrQzUcqpv8SHpjX9vXDRvy1naXFVA8X+bN1w345+GDy7q
KCrm0GHwzVhLEW+W8r0Ud1Rz1aK5HBQQgeGwOwCIyZfrM5CFKPGvJx4DPmT0f/qBCQF8CObu+gyy
S9V+KMmcTqWzutnktzGYwIeR7x9mM2gTpuFSPt0+amazy/t/WzbpGtDiTpXpBgMwE1+oKPJMAuIL
DzmxNah42FWN4ZNtNPIgENaovsc2jdetYtmiPnBqksK5tpV1wMor9XzOgDnLR+Mg8eKGUmXAs6R8
I0ejyGiH6ULtvFTThGj3Zs9NDnwWPmWK9OASnv6BILMgGyGyYrdQdHd17ogAgExhIPn3r6zvU88q
rHHLcnTFqfEuEIrzKa5rOsB8ivLfLNKhQcUyvci7X7gdHpxk9KIdAvYEoqhaNmv51IqLYI6l3idV
VmCiXuOip/S2Axi3gjHFgvjjDQE7ki3aEjsXJx5nvyHNgyhxmzvB2L3kIlmpmFEkI3DmLLHXpdX1
4EgoNs5ucuXe5Q3HPxhdwcfCWtlALn1yznvJEXK4YudwsvYAHrZXL7Sn16xW2lN5A3p9ARoZrMQY
KLXYOgtjuiCTeRVAJhU/BgU8Ow2xxOgTYaxNnlevMxKNEuSPhOxgQLegvZNyLWS1vK8OWJdMNTT1
LHx1XmnTx5kdJt58M/33iTUrfdZZkSj0fUauQoSXVDPoN4P1mfwdRrAGbFGzShTISxtA/sYLCpz4
d3hwYoWG1iK6iGR3qaojKLhF1Anjpdu+01dpw6FLXsM8R7knw/nAfGTcB1s4JLquNzRKkC+eG3be
8ryDnfBvJUwIR2slgtamXt2VH7NGUmRr9aqPqv9HVrSWcXsX7SJscslQhZTVj+6MJsDBQ8cUngeM
1dU1jHY2DCTpk0a/2vaTuEuml4GUW2BCyH4Hy4FMuDtmvjxAhdEwAaC+jxr/JMJCckgENq6tOX/S
9V9++cvE0Ya2zTLYkCv0yhWMUbFHRw9sHPJG8JyvnZeUPTbdJtahMbxizfMPj9/y8fFbd4dJ+RpN
p65Oh10qAkf0zPcS/wSWP7ERqwqqVEGsEaZuVBL8Ks9x5/mOq7Cc39d8LJrYvbpwpg90GdK0B7rj
LSeRqOUzAgsRPijektcCLBIpuohBNXibq0wP+gWPP1ysnR4f5Zai3JsZhOT+lii0Gb1S1s6WnnJl
DX9aRjTZaTmSgLdOppJCRS9mKzPIOPqSQ6fgWmbcO9/FkR1ablmFfS8pQii9Y0IvOfG7xuGQ7rvG
MwqONeSgTcEwbcUlpccmKSpyXBa/AWq7k7XloP1hA+vmmXrOY+C9C3192ISAw3YNRa/WspzidOkr
YjWdms6dboJ7HkzgAXGSMZbDtewlqYUodDQG+bGZMoqJVXQ9tIcEkct+9yrfayj3lgehQvztj/co
lhMzp1TZ2wE6d0LmLjK+e+Ixs0vBNebqrftCcGzLr//0OJ4KJEJCpXP2SpStX3hmkN46BhCeUX9u
rGcobwutIt6lf/WOOCcyQ5LoWL+X0XN9uHnyWAtaZ9NxIYYyD6YbAOcNpEj6x9QmDvjfTVtqMc2c
ufG97oV/JU7gM166CJ5LI/TN9jcu7s8dzwLQ9s63fIov+GY34RJ7N4Gz+itLtUq1l361ykJPyeXH
aW5TktgG4x2QF6dQ/kXwZQvHXB4Sa8ltYI8C+CfULQXymCCPMxtxRhHuhrGyT4Vx3u+OIEpBCfkI
1vdMI6H4xiQukei+/FsLU0gIMAFxvrqqxTJnaQlSSL4smZDLpDUlG71schX9iMHab+hv8CEBi047
ljugUvnqJ+sC8FeYu1efsfsrG7RII0vMngwBrXEl5cxAoVXPRbdCcvtA9Gjsq2WkEqjl6NKKrmKh
QW4sVBj4XrT6AH2mVdLrArEx67aKp5c705YVBc/8OJxo5RthXRqAa9OviTstIz3qCa7GzgWWDZK8
NQhZRomvdALSfcu9i8WFbX3PKdBNTMaJCC63f1RD4z6b2E792gZWYH2ZGQFMKKk/rhxGHi2OKnGg
7y0wbjPizLU6Vw9fSLlNbSXYNDo4sjiztoEbmsuWcw+qM5GAtoQkHovzgrHfevroXaHa2yUaX69j
zJY3w70w843EBYw/XgoeoAp7WS0LtKqLznl1/XxBx2+gk8VwIHyc0ByxCnq9yRgbtA2mqHglB+k/
mU/xnTEx7Q5jr8MMNQS2xEcnCEkTMu/xCd1XNklEWCuDy+IFkNCFky5rVsFAXNMZAkuvitFZJTOZ
GA6ow6cPR+ntiVcSBmT0Tg4RX/z2xiYIIdWCguDU2MyD0mhcyVZPj/ij8euFpGHioZ3wSteCKxA1
B5CVo9QZif8aSmuFAJReRsBVHQC36KNzF/KCNMixpz1c9A7yKuED1oGzYRnWkBngA+O60YRAjyoR
K7Z5c6S+/L1niPYoxJurkRkDDEUCVn69uDkC608Tf6nMk+NkjFGggO6bCobp/5dDbi+gfK2faJT4
3P2gG1uO3TCpKWBfsBl/uC/NCdrcSO4xfjED1bBUWG4u84QXyF2TcPgxXK9NFWH9qgfpIZg7zrfA
NqBsRDjfVUtZh21hfztNRg7ok5+EiBQ26Kb6r6bVPujUFB0OzD+pIa2Au7mwPoS3cuw7EPpe2HqA
21jaeS59FNFMlQjLXn5U/giXL8R2QwVBZ26dsjckvjE1Nwi9+dk4b69IzMEZaLYSpUISsdtZSxGv
3+sG357LuO20FookMCgfxHGTJqvj87FX5hInCQxxEEjmiD/m9O8u2pGd7Yv5nl/z1DFCozziP9yw
laG3Txt+fLKqMHXHAVDPXZGWLNO3/nAh3r6/sFy/hrSijhHLhiLHfjkn422PK8uGt6L2/x1pFBDy
pTrXrfHYWZzMTpOe3neRpyy7coqeeEMRvMvq/RTzhGFwIz3YFbt1CCnMUZEvrmVBLH3OjMl7m4fs
MvnSacVsg7xhg3if9PYXbLfWD/1pBhO3tfJbmee93dUGsbCWgA0mOBXjd/AqkmeBVJH72CmZPiu2
Kr3Tvov+hb0Rx/pPUwWmbgt6sFYfYyqNOF9tYHPiLQI+iBhkPNMQs0BXBiFlBsIZ28SsFw06XXdB
myRcZ3bhXQFTHq3TBBF1N4Hss7u6TJyRVQhhw2rdIyIVaU09JA5802YMdFtAcqPtoHi6ATfnjRjc
LjFJBJZMmG0z4h5iCljeEBE+3pz9jawt6yeIGHpMbMI+L3rqlpUw3d/Pc8RLeZSbupbf2345zYbT
0b1PUnleBTs33sLjU3sV1PQBYvztFHGrYyjzVjSLIfkm3Xa2W9BtojUv4b7UJvgUOqpIrdLb4P+z
1DGW+jBYjaRA8zL2m4Dbqzx2MqE1PjA+rgwmEUbwd+uaCE7JyPckB/2/4ZBWDL2gtC97Biid++3T
QpmqaB0N+xxF8ufz1y3naAN2y0nc2HaQ5iLmZvg1AYcaE708583MGxUE9XiY7kFZzvrtYopqPZ8A
XG94Fsh+BkbNeCQXz1YXhc+BN2xtue1So7emGacdHGYTLzz0aC/2jfSc9Gf1y8PEqx0+8Tel4aOO
D/EMGQ8c8LhpfPnRJtJHB5g/pDme6OLCQ0CVux4DIhuV4WN9dlyUkMkcful0N43kJOiqdJv6F9nD
qU0XRwlgGDHkFkGm/+QY5V5MKtINe8YvtZEjwyGDn5eZbbjcLj5sMEP8dZZ08IXlpihLMuuoxIlu
uCStB2frZI19fySVZoF7bP4RUPyplIqn1O1S/Yt5ldiWdsBoLzkKj+brh3unniCTAWOLAgZLuF3K
WivZROF3ymZCMSBxkVsHI9tIQ95DRp2Ws0XqI9vFmPgxfWvLAFg9eVDx5IwC4xOpdntZZADmaEp2
sWe0Jq5GHBreTidj/MOF/gpnYyYfBLcbIZu3dPW02OHE0X6Au0mzX9t/DtgjtyLJW00xXp2kA2YY
5u7bPrTwtcIjQ/ZahFy7q0x/JjIOzQ2zL3f+YvS2jggPGNE9FRjcyeOMn1tf7vjrOE9RadDgnukm
b8VhGfIuE0UCbE+AaHBSCTY0Lo2PZeh22R9WMJpzwd/sjraQ6eW97Q/8RHUKlrkqXsLwqOpIUgJO
ZCCDrkqZVctpQ8QJzzVB0Fo1K5mnY4bGlfxDMYNigbO54YDKZ5D85BWw4Ys4C3bs0LElLyLcsrpm
w2dMRegQwGKngTZBA0KesVCC2lQ2xK0+XwL+6hXWQCtN0JLReJu08JVnpwJmc56ZWv72sHdLg9ad
/WKUP+Ks6LZwtDOLb9W/fAObbInbAsFP6ZuaQBqQ1Z75dkCys1BT5Mlxrn0+g4LPB4moBOggOwtr
rHmMrEe0MVE8bQ5BN7atTTVKGidl28RLXQcLOzaTVAlG/Pt/K0m102L4NpmLGyzP9aoNnZc66Hen
GildQEuOwmgBRlWxwZdDX9B2zPet9ktbjo+i6YfMyjodmlvUnhBMfyPGUEZBnwvS+CfvA0ji5uqQ
jNBSa9oXXavXj59BEK1wLO2lKoU7awhaAoH4WXbxs0wYcN/HdJedcX6Ctq4JkpEMKnF4mbK4p80L
O7UsVJrTr9fYLnsxLCRBhMxm+uwudnYoFKMtIj2H4ZpqPGrHUYlQnp9KOMRqBU2LPv/X1JJFu08a
WqxG2eYQrgRaUywVR4Cz+J8uqMO8saZ99H0Q/iGAMHpIhES44ttbkbf3vKNx5pfrxExeIRQ3aFI+
l+LN+X4bxvrG1abcV1HrYY2TKR/iZOgRj1LAm3Kv4zOGJHsFMSww/r+P3weS8WIylp76LLJRWZ8H
k83BYo8xdQcADWrDDUi+zQIfSD6sggCeJxOf9G/5GYzGlzEanpdhT9X5GcpYfjngX2bbFosBVcpv
aAk2XONB7bq91t33cR9su/tgKAUhYIdxnVbd6u28QuLOMWl5rMcS1O55DTP0hYZmnh0xMb3nQAq8
wGxN2N0r6jbhvWgxeFwn2L7jIHT5KMLff3MW/sxPxQXB7MgDfXoatS/8NFtAjy2BFChJTVRi+tcM
8rDRwRZ8eXQFDcPN+h5BKpll9wLRt8O3dH1qKTKgp4gW34bpMkT759Q7Zf23rYQE8zDI0mR5RGeD
HAMzyBbdnWaxRJ5awmNeD4RQdS4Wi0g2ozfrR50K+0YYPVD6Qw/Fqjf+3CDKnwK8WueS+boXDwQP
kVmKN9EKnsLuFqiYasXXhOLuyvD4d38zjqcTM1hzXJSA6eSDTtqMtejZ/N1R/l4fyWYR5tcO5C4r
sfU0RRBaEtjZVhVDuBJsw28bxnlKbRPJUMv5mcHSB9n1aQ77hSGw4rhKFh1u7QelLUC6Bb4s4y5A
IhCQQqfc4nxUtDQ8nqNC0S+T5OAhJLSwsIVnk2bcOBhW5R+TT+GSQmiK3iW8l5MMWUAzJNxywA99
T2FerMifVjlHwSUtk94cGY+fpNVHTaMv2DuLIueMooJBVZgmNAZ2GVpcwvJYvsELPQxVW+GLXUOe
bZdKZAmETocHWdnAy5w6Kgt3HcxdoE53WJQm12Ho/9grcTInqwVm9fHXU7m/4KYMcxOizd1TkD+s
yMcs2JdG5Wt8QhMEunF0At2Mwo+RiYS2JgfqnsLLStkFfdays+3gv3O/L1WfAnrvy+f//hd3JSUQ
4UcuJzFqS3wsCz3V9Z3q22UL3OrIQtAE+hG8N4Ulel4Sg+HURucE/Qj5mf1GbI3i+ZaTEamWqMtx
jX2JpTccgXVOhPnUWpzIEAa9h0+10k5Bcc8nhtz4xif9r2QXr0TImM3lXrkDfFcYw3RS53nKHvdh
CpsgaETJvn20kbcLAzg8vdJM1sfWtFvqdxlONmw7QEvgdSPTHw2+BjvNxo5gDFZlwCwajDzWb+h0
kYQ10E5Angl+FbqF5PQDSzBIyE1vASYXYj+ShSizLQDxKRbW5/L53Y3L39Cr/RLbJ/qqjilh9oln
iU4yA2Hl+Z86aK3EgN09enSAhHw8U65sjbLREzSLteZPoDmjm6NNCytmCpA0onxhL10ZX5G9q1Zp
yU6Uk9yjzyYxS7DQIfpoYMspNAUoQ8iWzJ20yw2MmtuV+lPnJRBMGWOLHOBMZZ0x+TU5VCEVxT7T
kJqwVEofMOMPpUFfWdS3PCb5JyVl3mZ0OiY2DNLr4gx37oei8xFHzTrlt6kOV9r3pgtOkr3mEr0Q
1uL7EUz/hciL4Ky7nVX4bMR7NtUx/EFnhBDcDUAwXBcx3hR85ilyWmQLoeFWP7npgdtgmTZKo6N+
jMKbCw/0BQhO/IdfX8qDHFAAK1ydnnhH9LPXCiFiAPxPNAhI4uBs89sK1CeHVmP5aTS4ux5oGFhR
w7YApcXzVPLn7O9k3tRI5Z8WjajE0e+bwxfDa2rd0Pd8P7XvBtqNZvcZ3pQeZyIIJ8hRepBMLI/6
l0P165FzFIcX7qtKGECCAr9uFQFkDVvGAXUpGkVu5rEivmj7Hjrhvuz4IPeohsk+BDbKMAgrVyDd
T3fZ7RvbmPLMd2tVFPYjGjY2EFN1DuI5v2fdeg0QCU6xdlnF26vLISl2BhgHGEKWDhQDQUBD/Iha
wpt8gQ4FaIgbBlvMbCnGSnRGgAVX9cAs9meaSMsYU0kTQOSRK7OJ4Dv9dhvaxpZ0JaT67uhEJfhm
Pek5hoQkLUYiD7At5BPunjbfpWcOAiSrc+bd8z0oB4E6zJQrfqEGgM4j0KfjWv1n0juRw4xj7GHc
BdjwO5YgtVAXjFB1VUuMNZUpGVyjWTzHWMlV0bmytsy8LjQTONRmXp1w+g7LeAoo2MHI2FtC6YWH
EkaXTSCLI2xav2c/44boI6catzI/cgiPolnmx32w+QLVZeen+u9X3KIilGrgxFdo6o/fBT7ZUG58
sTxCuVapOLtw0fONxhfQzNr9e+enrYmtg+D6aPA63ipLnjyaSTyPXuF/YmMyMld1WzroOnsDSHKn
4GZMIJKPeHzQwqu9VjHKWvKnV6q/pfvTlUCDC1LRSFEdL3Htda+p/um8Z4u/i07pbKRXKMjZ6zYg
eul9NzMtV5TZwBSaPiY8PjAWCMI/RZMnRBEj2eyehBDtXLdMEkBFUlve8eM28n+omIBbateniFgY
OHzi0Rk8lKxvCpY65PuGk+2toyW1vcPue+lz/RQPVyt7mqISYfQdm4hNsF+pfkK4Q/69bpENpvB/
H7O9u7S7DtV/hei1vdCTpGvwJGla51oPpDPpY0uxCramM7y3XgPsVa/raxXaw8v/NWSOf5XkqbH+
DsVb8/hcSnR/pLfYOr2uo2S8OtdYJXGmPBLzr/H8f4klPTmZBS60XetDBId4cWOGwHgFNKHRs6G7
FctDtqFss2UoIPreMsav6TX4Yakr18AxjfXis8BOjODqsBzZP7bRj8pDn4jS+7ojDm6HXJbNDc75
K1M/kv0CWe4nzYRkyeCRLutPypBELO4NHD8uY1MR1NHmbS90MJRh9k8DU0qThjPUmETiUyE3dxvK
gRTctDz6o3W0wWnLhi3KPCdLflWDbDF/AbbCfufbGDCTTiACuHoQmVcqkxhzCRIYglVVZC2Q82tR
wi+lPMdlld3d/kkZwWomZ+iKSX8EWwEYmmd+JSSdPxK+4PbfGSGs+SNYn85ziguqpW/rEcQD3ykR
gyiChYtFUdasbcnT+lcpyyOJ/mTNplynSHrcexpZpGZcyf3ts0fNJeh409XsKbv3wy2hDGr7JHvp
lz58qKQJSTOe8r/2J5smm0ZA7D/TlpADjJ2ktrfW90X/wFFqyzkTW04vg8BbE2/PFsYWDQCSdsWe
y0mwajE/Ey+yMNVvGIOE7zInLJzY0pRX1VEjDzIa2FO3QT3KyIMQesf81RHltgwqLUiXtdhXbh5L
/DWuL4EW+cEZXRrlRrvxQhDsgiDdAdlxiuio/TNBjFFw+yaRqngR3FHcs4EqKu03Jiwx8Xv7VwnG
S/99R3JJivtUqa9XDgYeEicsgaquK4RIaP4fMHZzy7GHuGlOQ5KEsmlbWMv8i3dIMNm6bEJZshgH
0zpsat0QBFCO0uvOG6g4eAiFgCF3Kl6tfQCeQnwFDprl94/9502q03sLJ9kAHFMS9bzKujLeNTN2
3q3aQr9qkF4nOJtipOYCRbt+XvV/tG8XLSnqqEZInBDevRFZeiAa/59l+6nv/MNFIaBSxnwXiNbu
0kwCxdLvQXcg7PMb6gMKkiLVaofK16+gjsaO6F7vXIWVVXWaXhyaLZbYuc1dRmEoJzwFc5TDqITM
KbO86GSYOjWLRZhH6QE8ojLNW7PnTwi91GJ/RscZKChlKDHE3a6Q1fy/TT3QYxZzuEaDKZev2Eex
IEOo3VNGkcK5HxLpB3CPvW7gLKRbB2eHOMwR1BXF7j5hsgi8N3AWacE/hDuqbYyHCKxNX8qzuR6c
UBPNUFTkBE0hW2f+BHzHpICsuAuQwcB6OeaLkvzjx9wkTOoM+j3nYQdFmnQdAwYB+kmqkn0uhZhm
Ib5RnMMkKAHySYo/7urRJt+jx/SJV7CoenoNaeP8vHwp0NANz9Gb4FBJ7mmxhIV87jO5iUpVD/G2
vkYBsn07s0Gm/+FdIujwlF1PKMeifqA1RZwxqlmiTnAxsxliy4F+nJkSd0XsADVxvNmhYoW7HH+m
s4pwta/8KQn6EEnIkplqJQTpGRk2EBzZGgIBKBDt/HuVc1FAeSV4JQr00Tl/quwZlmm6psYQWFB9
kABZnwZ5CSMbaq6kFA2bT93vdZ7rSbvEz+LvWXfp4DH1EU7AzU+Cc7r8yYNUDGs407Y5sJNmi3fB
Nyha06464SjhFcjYkollW7LYmmsgszesxwp6i1JBbyv5fvXXt9ZP83fpkGarfkOw8axn+5EM9pLi
x8mTy5n72gKyRyNQ0e+HCmcTbhNH5lIYjEHI2r/j+RmjvQKcw5L3vMNgaVo3h0oVsF7EuluTHQjE
rCxr9q38hCdKM5Tyz8JvmiDgObKZNrYlAmTNpPzS9JhMLt+0snpCK3RnoM9Sgtv3CO9E1BR6sKi4
xVdqnM4r3F5q++K0VmXYe5ITtKifXdBaAzY9puAN9PHbM2YbNnTORikBDbL3Cd06OkSHadfc/xz3
RU4G3n1P1HfMti0zl0MC1A7C0Xny+i9h1vdK5rLmgsJKwLw9j1U2I1vfS01sdLFCJMv1+1ONxvhB
JaHL9i6dzoDlGt6vSl+f8p2qiiYAxvEyQDnupV4MijnZUyTsv+H/3ikhc0tSTujMyq/IKTuP0/bS
2R24PTTOGpnx246Va+Gz0gAHJlEcJD5IN1rmINpgM3xZgc71DqbrQWZII1jHpeUmoEvl92M5zXuN
Dus4b0x1GRKdaFDL5Gaq69pZm13AuB7ZkL/Ig9B4chE3WeNHz99HYSgVCbIzScR4Sc9fOtQgU6AS
d2OpRyeTxDm4c8wRIZoAPvuwYl3Gl0tQTL9WiXp9ckBjNKgXYSFHI6YO6i1UnJITzD1UHc4+zf7h
a/sqda+2yFZqEecxL56gO4iWv4+uNall4vo9WPq7RDaSjgCRnJ72qONohGijXmMzzwvjQaVLarRV
5ijLfgxZdHPasGKN5M+GRmWMpDz9Yz/qZLLBRG2OnO8xAsE7GPxecxtQwAG5WBUuW03P8CDuGOug
c7Mj5e6xgXUy4mWJovYSLxVjMkDFp6orYUjc74f0WBgU9h7WH2JIkBuLi9OAa45VbdVPjs1BZ+5D
n8Yyv2ud6tGipGOej2vOd9sDY2ZX+BkZTyC1QlzX8EK4/Z6PWwzaTSEPBy4hL4PbuCn8a1RGCHOC
RP/4Rg5pDiZWo6LbqhGY3VQwikvsbe59pEJF3TQoMiVjYaeM/wwlyliK24MmUynHTio+f3hmijuI
bS6kN+e3sv9YXn2tIQFNUgz0xZUfj1zvkjUmN/owNJJduB1U2X7fgXaxx0otuJdwYpZxIhjsC7Mr
M10WZoZ8pyORShPx4N+oL08NnS5RCxkBYKtz0MRqjV8U8M4MJPKPpN8JqFi6T9sJVkzxqLBN5Bm8
pWagGNr1Mi5A8lDDwCRQYlT4IcFtB9PXRi5+q4XZzJrK123WQZdk+rPo1JZt/Wf2UeX0FL4onEfg
KSgTPo2z3G7Sp5M8iQiowA/PRLEpxNbc2RuEoOfv7iuZA8AZCUTwG1PEk36/6ib8umfwkKTbqMRM
z+llBYKnIDpAQEWiMh889DdvmAzJm20QdFZ9hwhfesJroYqgLdp5H7/ND+iEL6fwACNLENHwyRfm
Jn1frGGsnaDoHA+2vuln+TTwOZagfasEpEn/ZkPFiduQj2nq6XvBrCEPaPssCqQD2mqoHDHt0wP+
3jsTvhNxCXkd4lH4drZDEuLsTRvXYlbsj101XsJKD25SpXGSIYD4robGMDGMwUuqA++KYUElToH3
CCz8pK0a3mo2iJne6pQs8Dn0/PSOqMBF+iuRJyAZ0+mcqbU3tTJJuIbIL6HuCInBSU4uVGM3YEE9
DBBh4os0SutDOIlxCWutLMNcnsGKL6K+OCKC7bnlQqo1LZFT7Larr2nLauoP0JWDJLHKX8vjEgjM
lDQW4pw+cmr3oqDaIK5MTuvRsBFo3k4EVZlYupF796X9A5mw4T49SbG5xcGkw0GDvjy3cbf5BtTW
kDmbp1wBRxRwLK8vQEnEytIAXzF/qxht5X5aExHVgBFWUd9GONp2bm/BAHbvGaB+qn8C5FxAYCh6
9P+1uMF8IMbh9QHtjp1w3jT/qzjQCqnUzp40qQgrSw3gairJ8hbNAzmBSmS5C+tOL3rgkxHE5pR+
WE4CvlTGqbz4dFfli2vlr45f1Jr3bcYmYW9BM0L+Ud45VW77y/INoiFcrVNsOnErCm1F4XFMrvUD
xAVzI68gNEdzLM7iC6RaTSHaT+UdE09nI8aAZBJko18nZE+i8QK0VsUoKkfGkgWicLM1KCqhdXiw
nyh8+iQkr/oIbAr9YlbyGlL6v6dBy5+nWRCrcPhwv7XozmJF6gzMuo5qUSEcgQpGyS3RNubQaU9z
z/eD7jIs5peeLYcIUCRXwjuTzl4m1RhhBB8d7zAigeFGGNS/OGBeh21ki4lwAMbju6fU4nqPrBGx
hIPF0jHrwIusrmaH2yL22ddBXpDciMMNNjRz763HnNF+jndeJOPDRoXFa8wTP9D3zFmOTDyT/rZW
x+cCUNaP3O6tpm7bHKE6JJ1UzFP5FQ6+io5XTOk4xR6VqM0ohmJMzFcywmY7UCirUWFO6e3po41n
eoomlbRbVDdNky5M/i6CxW0J7LXDVSYPHu3xHcXSFwbiOTY+itOXrTmaifj+M1EywLkzCwA772w/
eF3VTLR4ZHWu0sBzwysjTUbqw0d7ks8Q3XHhBVQSm6wJl5YvdvlXrd8vwdwhdPKh+fUxcKoqyPMH
Pm+aG/HM9sAqQeDHEN3kuroNv9SmFivSk4BT3xH2Tsy7zzffooCvqEieDkhRPK6Qdj4HebHejgxa
POY7ogiwpMQb0jafjF1pT00hKCSOOc1clsA6iaSIKRIOE9xE8LQ6NPsQtn8B8f0sfg4wY6F00ILq
YtWAYqzI8TLUeQErZlLOa1lChWE7sKVK9lF0MDepTNnDoO8SLyFQfUxpkwHL7H7g/u4CeyA5VrEB
RK75bzgIXZEL3TfixM4x+SIO2QhVNTaDXDwKV5Le7yeDuT3D17hb6KO3yDDTjoXvMuzr1lbPzpQi
E/FZvuq8BAipv8NgqjmFpUPpT1/nug4sJOSSAM2H0/OrWHj8XYHdwHyO1lDPveFfP3OEy54R3mpi
5sMZ2CPtv49VBoL5CGoKOp7hHM/gbRVZrbDwZWq147VyVF0SXBF8FUNoM33Nfx1JH6aYiPyB8rsB
mIR3G/VJyGkAMDGugN+g/GVfMzmYt9YNnu1rDbw6riIQNxVTttFFLqwJefszaHDxfQig1dkzs6Zq
JXnwimvFfzO0LYJVJIaDjbi28e7PnPuxHD98zDze84WdbaUihMfCze2YsHITPVx7OsIUcKtUpRYl
xDUMgAbM+alECkx/UHLSRiMDxhALLa7HAoD8eId9Bc9Ownv3h5pFAZISdIhoqa258qOlUHCcKe9t
xu29PlmzSABJYPJso9dMHGGuEFQCtMIKoKZFLEbbObrxHeQhg1BpcOB6sTpJ4Sun1aD6oyuU9+fs
ocy+iLvuZI2uGi9C7SR/xaoh0rOyJ1zYwLlSSLoruP9UB1ngYlQ2lu/BneOH3/pWYuSM1+vH/etj
m/EgQ9WgjS82dL4oQcAp66j6+wHNy1Vu9xqZvn+FCT4meuBfYl+sYnellTPOTjmADoKfhP60ab2L
/hZlKOfGCWjRW5oEruqwX00/bz4UBuCQBMpCfvZjCJuRyWqMkHWTuI0yff4ZmMH7BUtTLcgoBHGK
nMHLkSj6c98NQquiGuovgMHGS2ugRR/rISR2EEZBp/xA7dxkrIITEVtqOwkjdW0EWoGnQBu6Lcog
kQ9OLEy6xp9MZpClmkeJDUmCsamArgtHgNkaHTZpags0PzlImKiq0Zar++fwZovhqZv8EXbXeXkS
LNe7OQdRmcDEVUxsruu1OsYBcTzcUn/YVmgbXvv1N/JG1hxpb2FYiugSiyy2Vw7rEyO8C6iCmXWw
vcxtUa8v+71YrGkOsxNG6kBoAoa+OmlZSlkAQEUbVVCj+jWHuQx1S2wAwjVnypfuuWqdPsFuzzTu
KzZTJLsUoPb4BGEVLXOoblw54GQkq561C90R8JP/xH/sZmmxta0gZCRCBdWEo7suLNG5fAhBXaeh
+XGEJW9YkP2Gjwur0ytBI5vo8FX98flb5A9FWggsZO2ekBEaa93uvlH9sVT+UxhFigRLjE4Eu9YR
WyGbfeDcQroerm7j+sOpUTOow6m8bnc80fSy1Xl4rh34GhYpFExMgG/luaJj9OeMuNAooNfbJxxC
d7Mq9Tu8/BjwDqfrV4D4iUHZSZupVp1xFdN803LGXiw4s5q0NtXoSZ7bxml17hUlvQA0ILZW5pdx
Kw5irOgK4ZsF5VCtHMWJE8RdiulN0QzgboAmh7HMLAZ/iFTTf+xnGEfkiVaEwGL5X7b2JW9UNrax
RcrhH/in2DPc5O947Y/NwOKhx1vHx8qNqs5FrhiK9tvXuquForJBZcMXXM5s5cEexTEsXVd0lX+J
Gh5Brvcy8kX3PcH1BvKn5ACX5i2qFN1uakz3Aice7DjW1mwWvdYGPorg3mB1Y5jKxcbq3U/MUZXi
I5fkCCXu81/8f2aeJIV7HCy6W38Vp1AS+UoM488kZ0KgfLmnbkqPyGehQsJrbrYMBNhE37n06Vlt
L6owViIzgSvEVfbmPbuyJQ9QehvyXg8/YQf7ZlFiZ0hvK20u5SGvTtCke49QCParUC3oPm5fiRc+
rRBzZPcJFzYijcHbwWfyXLcuQHNOcVHmZpip+a8rQOlUL8HmfcdTsNtMI5VgzMiBMNe958hJoSjV
IXO1gIlF7SPpsWHddQVLIFYz/6b/n9yuNehucPEThmO1yKlZyFBebxGe8P6Gf2I/RW7CF6ct+j6R
qIinetUnfj0h9QkljAZL4v1O509yeQ+fHmNY/mRvrn8AzQAb+ilm79O8VlEVf0cDxj0FG+4WZcm3
B9AW07RcPAva2DR+bDmnMhGw0bCWXn8pizXflK50VmUOkuA7ZIs2gON7MjmOREG7wj4XV3Ubavch
ujTr174Mn7PtvHbuRiUd8BbglGaiFN/PZNIqVfyZarUqQoAwBi5S/oPp/59wailpXi5AAZNGi7Lp
Jc4LKcbzz51/pQEmHqlU2/JgSy3dbK3FL1tlVeoGwl2DTH0SWCS0yVcoHxNwIy0OdESq5Cbl31n3
rlZVJp8wsAy0ayJcCuEvanM5SMbCp0htxfo1eDHW/ddXabwUnFZXRhL7Er0UnHBS0xKFQVXbFOXp
Wb1iFZIoB2i/eqOZxydsXe7K12QwFdNPC7Rgfdz9TZNzTi2WlGR1cqnc/hnqV6M5BjmAn7UaumRL
4iBtiJw3524cqiWmc4A4vfBQxEW50eeG1Hg09aalK1++irZ0QA9l9vFoUwowzoIXmm7W1zneIvoo
je/fBJYwAn9sqfsJp5nifgI8L9go7tbrwWQwTC4LaaHR+uZo7HRFbxXHsgUi6ens6bOIfdd1HITK
aLatsseiC+qhtwrqfZL6ia5NnALeyow10DkEOKh4uU0zezyENT+wVLSgZvTWUj7Y6cy/D9OqjNVr
3CUQ2dDKuqwPeHRo06SNfGepuqF207Ii7VWv1PsgiQYauc2RicWnmtnQn8hhGS27hVH+iU3akXaS
+VyEiRniNuLwTEZha/xQJ9z9JOggpPxRTQBt9RBVWaIPz1P/fIH7w47Obj+GIxNeE/KpopDcnDd2
JTqkZZBvVFvBq1IAy0aJK9CkS2QcPGxicRQKzJS/McZcqbQBl2bD5nf7NLLidBYeR4KqdIPMJyFt
c/y0Su6vKBp3wVrq9ieV75JXUhNsSf50v27XvPgwOAHCqppR4xAHTGqg36kRNczsijY5BxSmRQEb
o4/ebo5djTKL8TlFlfpqqTGTh9uCdTDZ73HrWC0RndC9CzE2RB7TNWOMC7s5+fOvUebTzBHhYEbF
yxVW+/xZd6rrKuJAYBaItOPLdKRYS7mETjaVoposYnQJt441Gxkt4ULExlh9z52phT9uK3rNE/+u
KCjBQLgyU3PAJMAkmeR3vJXX3R9gHCJ6duV15PXS0Zu8zx1B5K7YaLbNw0JnJqb8g99+5pPD7Ot5
7hKj22VxlMvjdM5IZKeBD+jpADws6VjpNJOw6Z22jchG2HUwVakwJUUgMCKQMCn4hx6xC1qyw8Ro
937c9814NfsmafoWroplxDezo9xzuz/3QzOtvOZzdqE3F0ZYJftupjdaw61w+kMcUdkv6z3oOYN1
UuXucxTJ3Y3+Z2gqftHmumDNqOqF2Mwy0UjQdJfJRbTqXYCEWqNzYcYGb9ZB1FcPEKulr0p7pIQi
1M3no/iPsjVdIuZyPA060VrhWR9r0V7SkFub1rWEUHoM9hWFT3L2fpXPvP15QD3fSV/umsknXnRx
kgY7aJLv8pfb5sHrin7BdhGviIR/ArHmyb7QdqK8TN2t22wAOqsb+IFVMxzmQ5bC129Yl6aqRyiE
KKpcumBLWXPFFeu3fJlXhKC7VnQkjFE4HHh3FCSvzF3o31CUxqt+jdNeC2tzMb0mE9UzRBL6Ppau
VkcwY9FU1StLgSzgAltis9I4hCpL/K6MRlpw34zi3HZyeDsRJzAm9PV2n8z5RgEyriXhjDZwJVVj
FGPXs0j7IEPxwa2UKPRNA4iA22FkzLAYbd8/rvthArNVZ2++XVfjweC+R9eaRSh8DnHS/KAAUpDb
2JzDVhhK0E77pE+EfIEJaFx9H65RoxzqDnU9UBcPawWQmdMAzOpi0QnWKzqg/5CE7z8g8j0bpMCo
oA266MZi8CG2///sy4ZQEeQPb97cBimOAZxGwJmaijN5W8GhmihaswEXGgw3F1zPlzSA77GNwkEY
3bV+1t+lMNWw+zvHVnrb0jdZebcfk7zClEOFPg5pXu4PMa6DdpiVqL2J7h3y33Tnav+Zq1OMCx40
jgDpQoHdK4Uu32AU2Obx0eeQervGQXkLeAxmoKFjv8ix3wCu7OYLSVSxOB32Omq2BHS6/UY5gz54
m36BZzxGOuINbX1WIEmB7N970hQrr15HKXK6VWZJ/sCEtzYy8Hl7C2eX0ivDDV542Xj7UixN3zp+
c2sHtaCQorG48nQedqqcQDiIMUTCTGz4W06FCgOLBEJT1RU8eUTj3xdiGNw/o2XE8N6odIeZw7PF
Ckl1bv7AwIEnL15UFX4cyuRGQ/ICXKs0ue8h3+VfoBQapkO+UCpKqtE1THQjFZEi3Er7IOScCNmK
l71ZG1hmwXbrUTpvd6WDKes6cKWNXAaab19f/07cVSf27IVghnYwyY7S7AMxeE0j+fATti0dPxZi
nXjT/6EYtK91RJOkqA7DFGFa6k3eZd+CaM1vJWD6guuLAtXO1t5/4DrhgfJoEqY+74J/gEbXTWaS
hBBl9decbf8ODle5dJmhEwYVg6ONFGY0Z/UCywT77SaHxQbciriNM4FkeSysobYkzOK/3mDQmHAy
AboTxJJcwxA/C2qDF4Ng5GAQ8h2ND2jZbxVoYEPxQ+DJfpvm0Nz0uS6KQGATjERlumwxLQPwHhD3
e1ovJyQbWnvlaHBoGJXOB5VSeKirrXCGFaIRO09tJy+h4MTwrC63f4grd21xVIYm/Mwmx/DAeiIT
inNxz65mut8OPBRfSzOb/Zn16+qcHCtW05caFP30Cno8hWQxQqj7KhriheGLgAANFrQQJbZANjWt
YMc2UrxOmzBaHyeywm8DcPL0YE8Og7pIzcblzwu3j9zOU8F2FNGKJOS9HsU9tLPnO1Nnd4YQjXRP
oOpfpB4MK1cf25pfqww4bAU7/iAUH7yBRFzz7LKPi7y0X0zZwlCjEwHaA+WCVh85HIM9y3/6173p
uj3OemZvJqwfZOT3/wPf33n4z7j8zvnXXv6D1cfR1HbK52pQOljIjMs61fcYP/7v77HPjUqjcWa+
7GXfXh8I72pfakZTtNs3iPEy272oOZctf2OT1pmf/VCjEWUMSyVJHgAkBAiF6kCAsDvW78tT5cx1
esHnHcxQD+arMeXA9Z28ovazwsnjz04dk+F/2qdFLnmVL5kvkIbsbglyCKieEUKgXuKWerS8JopZ
+ggdQUPp+jsE0IcOE2s9oeiIAEo7bLv2h/eW4SeJ/Kt1dk05ocBhdpcdFIav9mKVC2bzHR13yJFD
KESs9iG+H2Rye1Sn0cIZGMOsHPdw2qqywjkBRZhDMpg9zj6lDTC4FlpiB/Rs8A2J802uvIDLEhvC
r9o5iwoZVAhf20mPu3NdV73QypI8zoXo9+xYdwb3pVydfJYpZCuyACgCbtgLcTprfyrQtL7Ye0/q
3dH5hT/W1JfI7Y3TwlI7rw5NFsI+6ZCqt+XUKx9oMCQh6NTCTH2JB4UmA2bk/4aqtmPisbbZEfl/
vRjF3c0QqEStoJAhr4/pMMaEe2qF4zjHxxVuZC4QWLoe9rzK+SUtQjcTdZwoNNx1LBGOyWyBojHc
KR7UvhBKmVUeO2Ozn9syh/VMK+29jzzCGbtK/bdP2b5BYDpT1SyjnAuR8PXJnIHxX7V1I1l7jYJP
j6n00yb40QP46emMhVQpBl33fvPUZHG2l8unxsKkSWWDU+s88pPx7PhEpbkvMqg1dskKsAnXI9bD
u7QlAdA2xF8c1IjIOaCXTI445vbFaIkS+QoQYJWUJQV09sH5CTwyLwf+nqVxVYsK8g7oXI8MdSDO
TUbnrsYwnUcZjJ54ijioausutkoNBfJ/GTzqUueEeVJLofPqPQmBE60qz3b48UtEwVfG42olbPY/
2Cav6pSHmvO4YUlAixuMIrBHlubh3ldQ0YpOC5yyKoZJ1DUvDTGHIGTw+3QsA0VaRhP1ZM1w4WAT
Q9CWXs1aSqhm7qBr8GS8QRan54iRKsVfhyFs4ybYNz1T8qadn8HBwZdY50D5bPNvoXKvFd8N7udY
UPErW/sF2/fzgHUXnSjS6eziW+WLkqn9jt6EZEycrr8vneelXRJnho+9gRHPzPhBoM16LhL12fGk
5HSvVfvF1XD2CpbdZJZWLZPDZzhQEDnEpoAXZ8xpakGYq3B1XvkW7w3ykLpiU9UcC5mbn0OOX/kr
gVAZfpgh+p98kM4btO+XqgEJT/TwSkZ7ovCrgiybMGhThjul3be1ABr218vvW1MSRkMzUrCbYihO
wTslL+ISxSy/hr7X30yzu9nERFn9pe18nMPm75LaNlrLzxS06yI6pry59SDnHYm8G5OILB38wlKY
KulKPCNVf+JFMT3Adq97k+lNJ0rWJC70/6whsVldTpiZIF0k6nEEsvdbMNLqVmyqdgxQviZNt9Qj
ku5nox7XE0qki5MAhHO9OpwmuNAOfXWa8Y1OSxmbIJLfAwETBK6mS8LTUtGYBJsxUDSk+GTV6boI
TdK9nHL1llKY8Nc/a3gq0QodeIWkdlhOiWNH93EyuH3fWfnQ6sSECUwPNfstG/SedaYbVy4Y4ZBB
lOzCsGY31U0+i9pUx0NFY9uOsGb9TQoiQWqo/Vj5/ceSON5m6npUrZQSWi5WObj+/ObRqTmDmRft
g9TBi+Nnp7YDMbR4Fc3g3yVSt0T3Oc9iSi+IQbBNFL/cSHmzoCOIZN2uXRRg7zFPGTg9fh7uOJPK
rQzmo88yOYxHaG5hGebF4xdT1V8Rx3Y+l64cvFLEBi1Z1pQi9AoyPhqf1tleg5U1Iylq6pXeIXJH
drLAD7BnYLAxMf9eXqnS9LfnqHWyWWHankR7bZ8ZJ/6Bu1vE2PAEI51sI71P9/4Vpwcur0RdvNgb
kZTQUnCklXfSorY8qkG+RzLrd5g0y1W2RZGWCEKDU8WPiXQ5jyCNeVbaekRWk8ZS4BFV4y0GkSsd
rd4eHeQUxen69LHmmCH++PSBSS47CdtHXoJfl0Es+ZT+PLs2RKPkGSzYsMjcX08JypbjuIedTeVR
q6e9/GZ38T04Seod0IzA3bBX01NYOs84dT49D4gzXSMww2/k5QzhXoKRUaOJ5s9inhU5FRrNoWDQ
xyl8z7ES1gwymNFfNaCnzzNgPGP2l+Oi076n1olVj1xSo06zHzjfFLRG+8B6R2MswPPaIBBLqDfY
s6hx/zut6BJGfw+j8+ZessPsP4Ij3t7G5zyMOMigB3qQLD+MKqXIR0DKEpObx5Fyjju+rxKcd5yU
V1ejhtzZ9EM9+hIKHyzCx7/iR4ih04oyF7a8tzEvUG5a/NmCiY+9MQgqfpXn7pi4z12CoHBYa2A1
MvwHq8smoXWMTLeCF0bcnpcL88/HF8shAuf9HSRVAOv6+BQbJIV9wBVsdW8Rf9a6m3FWjVz+l7XU
EBAEW7pVrHQnBfg1m4nV1hbEAn7HMnIFLm1dS0PrWfr7Fze6oE+i6U8YLL0SwNEu5YMFsSzCisL3
e0luLttyKX40GQMH/4U1W1QugFqiZcBvA/eNFe1fqmD/B/I4JmZWfhajJKi8nxBf32xwb8n1uv7A
jNQ7onZMZBWSB4jjLlyck+fzdzEPupcVzSjHN0Y/CjxYr/3lfcmooLuGIG4ib51Lla5TqKxjaA73
LzkTkyyl/rdkV0KABHzsSh6i/85zmlGQ5xTgC7kxxK0t8LkxXIgZwYGMSlfvokwGX5eZbWtCtIwv
PqxqSmxh99UQ7PH2+ME1SJUjbBi+TWzrGdfm0K0wlMnzscH7vPIY16EPoQ8jynRlMjCxPoRlhePd
BBUjjozIEF0R71RlhdccCvpOAbK1t+lIndt8Onf6XjswK72HOB49aLR3ixIKJ08o6/ZTBSy9bJEc
WlDET71EiYwuFJa8gAZCygAjK5RejGn6mxhZYohnr5q30YDK8GOMJgVJKdcslJq6zPczlu6d//aV
XKlqkcbyh4Uq499vP8J19l0uIQSgWFQvnbpeW2KKPYYBuA0DBbSoQqcKhJkZB3UTdKby4DLpAOYW
AHVTQv9CSP/OGTOq6vIag88mXbS5pm7VlgG+OiVJEFpwCLar782AHhzlCcWp86eLTNSqCfkiMW82
isAcom6yOLSeoL4zAIr4PwutoYpaVhYT24zATqAO8ai+9qXAWUJYMf2IE6e4Dp1jhhfapXlI/zMl
oyTYQUhcxzk3deVzAg28jkLGUHnp2iTC2ye6B8w6BDpCfXGdfzm4qx9wowAxLilcz0h3VjrU1xm8
VAIRvDIoGGjS8h8xSalw7HLmSdaubAIUHyx6putY+MHbXJB61WL9Blhh0/WGLRpfeyLmdIbuleRu
I9nl2mBbty2UzlhgJG3Ou1UDCIF5NtyvcDVP8LZgzX2tcqnLPJX3OlVx3L9MdXciSkXGAFDGwhXp
RbL0GaZ08VBLPZyulSwNHoRAEEK/v7uNtI57JpEbWCmAropzL7hWUDevo5M7gqIDFmeCR127+bUs
76DGpqG7k+DYONk/3vQLJ7XYMbh9BleiEpTRGM+JV5JxS7YuSmYKhq3wcZUQlc02CvRBZhZhX7qk
tiDR0R1CSBVhzUwDHLdyy1JtF4Wd399/60yNGBVwGh/29hT6ReEmBHaBcMKo1jZ8jE9LYmmnXk7L
hz+WfGoAE+T1FfWac7BLn4MxqRHfnzdscRRgzWMdLffw32dRvblmBjTarCCck8eFcNqfKYeWpxOs
FB8+Uwz4s3M9I5LlKotaMC1QiZMhSMt4S8A8FF3ijsVv27TdWGefjXsye+nxAxnzFodPbFq/3HdY
4xQFoOWO9bIWtjpycILG3qyqEIY6GhKVs+3C3vbu4y5eegJHZ4+f819KzzbvcnG29Asno9DACgZ4
+8TCR2m6JLWoDIFhWj2UV6gISndWlzgvyCw7SXpGhTrR+e/8zHOs4OMn2AuHkalLEZgG7U6PgsAI
+ww1YWMyenpViWvznjTmIoqSgLJb5qXmITzdzGlKhgDUEdwdbIsP9ywf06xDcr77eiq0pcuQcd4/
GG7hA9TPvAKyDfW4GPciGkINGriEmwIaB3JSapooTNecM4PkXOCSNHmuqCxHs593zmusdzhdu2jT
KtWHFSTR3jSBSyTm5s4frFAnGiDYB5wOsAdZWmmaM0QjdaXK8RetXI9RLId0/HQUebITA/7KTLOH
wn0JDK2aMxZbnhn/jk8P190lX08sXt37aolFj5C3ND6Cxzlczs6goEpMe6fOj3hDQrpizJggRwrS
Jog1Rat0391T8OQfEuW9LvKbvBvSC4O8awTDlUrdWgyRQ/okqS/ts0fY03zhMNKBNz9/TCsaLRKK
h5rSPDwxK4rTjjs1nDjEj5r1sIRKXNx2t2yoH8YwnWSvw3UeCeBuo9I9yl8J7jYYUIM+t2Zg2pXy
q+72WVZ5puRg5kO30cqo6NHfApxpfpGbYfSdrB+a68ItnksgfNl1KSUTXytbmMP711R5MZ4t+o29
KxFQa57gqQj+UvJ+s33To+R2M9Hacm68dsTMHQRF+rDrdozcGIXVqY9YEnxJPfnOo/5Vu1e3PJno
yhp8y8c/eoc6ifXrJB9spFfoUJCrglMrLtoHHtHt5e5q/K97yv8cj5G0ByeqG4dJ0eIwtJYdf+io
OPTqYsZc2+uGXwS6cmhpEpHr+koqiuyIqY9PcEXg6ljWL2LuFK0rbJ+YUs44drcrAT7iKn3L8BMD
gQ4fBmWgzZAx2fgzy1qpSQhNA2/U4oIUynd/tghdasx3yEWvVCwhq6qNclWYe2PEjEN+P0UtHQll
1Z7NS5m5Gmz39+qJXmciYcMAkAqCzKzpl2sWbtNdOuxMiKrqIQGgP9Pek4+IgFHLmmG/4r2mGk1z
+6irNHB2T8dr0oeBkFTlqK7Jfe4AATiIvvE4YZwF1/ZZjF2oC1/xNaSEAp68PFumJG4slOyq+eJM
Z7w6Tfn4SHgM7J9nVRCavKpo9+obHP8QH1wYaBQhw4YGQ7vjtBqBgSUpE3OJ15QPYfDj+BgmkF1t
OhE8uTpgHqwaVbmUS+LT9BX7UiXEmtnXHC5bp51UkawKm9NgdSA+xwLHWFDNRztWvVJ9fGGpwV69
CjwgIawsYQAjzfgxQIN1htVc1TEZ3XgFTr77/Yt0d8liqcqDzbpqnBY+psoaO+b6w+oDMc4FHCWk
n0t23TsMYV303aod0JhhSY/frrDmEAvW6C76pNsbYWXAMAVeKWdSAv7K4U4m/eyLDxmTyTyh/ElB
se8ey1SQgL+Na49BbAzwRG6lNyHndNVQZqpDBCTmWyvwXPY8Umq/zek5CaizXlf5u4ZTEpzJxdvJ
NoRKIdbmF55NC8UBQQSZrStYOTUXjb5N8kB+SA391+f4YBiaj5xSNOWZNjmAfzMNhXMnL3Ju6K01
dMCwHHWUrCCWMQPtgifqvCP3GrtwDXz6jkUn/dxraWiZ16HsHl4LOXFmb//IMBdTUEnGFPTuS1gi
iRfaa+sjgFRs8ZiZIuyF5DkDkGQGNNWlS/mgrP5BSDd/jzefPAOOl/K62i1oXCgf/B8ekCiaXWu8
wZU9YashFXxPZIKyDKzJOp0hnenLYLR3vqK+UPlsNAkebO8PjfZlRZjo/jcsczxrsGpPQGSR+ptD
rhAzW09jTV8rrRC6KUtwRIXFnkBH4XGGzKvd08uxCqc87iDXw5mjhA9v5U4bumqv3j6d3WLnfv4x
RwWkqAOCyyTyUCKUxHBf75SI+FjJSd9KcW8sRe9X3mfM0LenWt5DAgfGGD1ka+t1sC7JE+V4x0dE
9aVUVdJoQYm7eBKTQLKyTAOOhc8pksm2R4HMci1ov0zP+4Jh7X5DPP6OjGsUJEdxH2JYSHHrRDrD
ehgsKEb72lqFuA+ldmuO/oNCVNoU75cMFUCWZAQS79SLxmM1m316x/wDhOK7pLImbqOkuI9xIcDf
XxvChyVcPpW/5DCVS5gwZs8x5QvQS4+6ojbvwe3wJ8GGTSZArNQmvfDTv1kp959db/jVs3MPa/6u
7QeWzkzqk7qjwfQW4+QGqLgQ61Py8LrL4YmwAtb2rHVcAcN/t+JojEz3pZVQpj4xaDcs3b8jXS7z
GPVUDcLz31BLMP1gmnAqkZ21XgBXY0DaE3olnLY8YmK9w2r4dba4TjAZjTcB+jaqRKrMcHYimc72
Aso2cOehVLjUVAyrOo4xaf0qFq34pyoMJ1V3nTpXCrVBiQKybrwqaSxSaHFOnpQL2TFW8xZzo6JP
7pN6uOrYPw8uypYL2GvuHxzPdSS4jBzwyDc8APj2lDp/Q0wz7NEIBCa6xwuSBw0W3JAxaXzdOyt+
eE2ywf9SDtREs2BvGZ7WjaLQvE00lRrcOlw8UmyPDST5maAMSQ9g/LjIq/mBzF3Q24IPAxB9I+X1
AfBpGpjwo8enVBKSzQ8IM84eG6R4RCjmi02QHJexFzsF8hSVRo8DWDOeAPkyDBjNYI1Kp8+ZO6/D
w6xcbkUyc8ShSByh7I7kgpK1phlv5zG2NohgxdYQi4SP5OUciremzA5w8ry/Pk7RhjjEPHGhU/Aq
je3dpzVey963ghusSCzIKjauFkpWgCXhZ7Ii6Hms0QPqC1z5ih8+0w0elHkQ7sUOi/epuVbu0aVa
4oCAbv8oBcq0HpjPuvDPbKlE+6Yy9BPeFxbu/3NR0MxSKGfFciSlDGbNcTh090nSJi/TeDA0aw1n
giIdKf3vQ5snBn29tZCGXZHpDU89dqkFOkOn5QLyWqEsasinTw6k7DyBBCGfL5esVCQkZC3uUJ+P
6iAnnvCx5AytmJdYMB34CuRvLyDaTH7gLNvRHCRRG4/Jywn6J8p9X0RYjKeJUb7ZkD6CZPXx5DS/
p6pq/4Q1JCE8Ckowrnr56ZddjU8LBQIE3Q/obFdcKyMQImRQncdjrvka1FSemj1UAfpy6W4Dg/tQ
+ibjkwvBOokFT2L/L5gKLDM3Tv2j2poENWbps+rrvEQptj3HF8giNjWzZ1p4Jd3su+s/7XR6opJ6
+3FrzGIFK9k5kPijZN5Udtu0IzinqgEmUpTr4HVVCAMwr7GVxdj/Dblh6w+/kcCZVvN36138r2HV
KPLqnFWCnbYkxCkVhCAM4oMLEKxBNup11xgDILMygqMClujNO/gHuJCA9QLynX4on4ddJ03psmXb
Gvgn4ASKtnGQI45BDvYCZdpgwOhVIJzmJ5Gco+DY1vdmF9CUoiZTf0PkEyhQ87ccX6k0x9UA0xmU
995GEPsRy3sEVAkKdLFx/pfhd9jMiMDPcPl1vMg1Kf6rhi51vx0w8gWctKENFe5OQ9EYAYgXZxVk
yZ6nvddKUWETpkFiyqkDrEzHFVen4hZqEFoD62QETglFbfHg+gDAK+h3ySIklico/STlkhlwNfog
h/WiAhyQqvhsYtKVyREFMO0ukQOYcfx+JPOf2pLPrzgdp5Wf0sBLMN1wv+iNBOrdgoiNdF5cF4yz
tt+uOi3SlacUpULhNogXBNMS2WI5AkO09u/zHYbA59HHHBYLg9hK+hHR90yW8BA4n6kLfARDBcAJ
WW0nqBTsDI2yPCyMKNEXL33oLYdDawmFgqggYOB5Qe+5W1M3hexNNXjJx8fYa5moaBhk+jhq7a7d
y5ojBDafL3hWZ5BkJht/W65mEMGZucCpeS8o/JVnofDT7kms7a03wfJheqMOwQljuKamMhZANOtr
lnHQ2bDjbRK7I+9So8xOi1o/mbChM+DcdBCGsg+XeNrpIR6QmMxBlMrqVEC5z8MFK9ehi6CVQx5P
JA72AOqus0e6Bg5QTb12EgoHfmwGnk7j6jph4Ud6ahp0y3a6FXLnFrzSYwBGF8+PtmyigibCMoqy
LxJlAErO3VkWI5vyzeYPAuSOuUco+deYtv8G8km04I7ILwuJNiZ39fgGanYJR/Xis/bh9pTg1EzN
UmFFCheOTOOGT0dWEVdaAvc8ZVvNsBdZanKmkhrc55NsSZbrI4Tvv8WNyRONmHMb0miJHOepl17q
gI787lJZZ+9GL7RMP4c5kbTwygS6GMq3pbV1wNDKMxO5qph1LJCV3zO2RUUlWviA2kh1B6kiSezG
TcGgHFjUndTBsfwOoPTRXsrlaGlfb2uJbL+u+IPOTU+vvWRk8igqXVRLoSd2rdVVavLKADECy7kd
WCawi3RlJIn2fmBdvAfEkDnsN2DfSCc4NxR64E6oQ0XGH3keQMK6plQeFmqQLaeBqAw8YwHb9LlI
ZswAvD7I8d6vjlSVzVOngxf0+o07jXTgNDYbSudfHve+B5KYNOUADqF1rMsAC+KgySgg0QDjO8Dm
erD6Mi0ISGN4wAMvRM4wGqDUeRZ//Cyo3c9D/irCuiMxZV2P5oYicNDV4p1ORtBNgezFPhi7r0VG
WDgvSvgniNFVj1T6Ht0WOASq0Z3kNC1C4wgO9/5hbgrnt0CF9Wbs3MgLiPsClt51kv+MLlfQMC9E
mHk0BgilZ++SinwuhJnPDbyVGsVFoYSKztCSLeYbzwffcwNDbqUCl7cn3PMoMyYJ1dLDjFaQRcd6
TWq6NC3IdOaNYjVfRZOBsFQ4ypVGLSV2ibl2SUXECaVqex+vTjclGdqwNJciZWQyqSgTZDv+KrOn
covCeeeQ2rFd1oACQJ01zjPvrzLozEPZCYZeabM4+mDu7gsL0riW0Yaei6eEJU19UViXDWH5Otqa
sWh2vJnKQc/+RU86uUGKNGbioXS1PtCEXVrFGA6L2BT2jlhLIPEDuNXJDLex0IaV5lf1IdkuZVwE
/kwD9vqI9dSU0XdxlypCqmnQMAlKBV+s+m1vS363Gx6Cnc37YyexQRp/z3jaNQ8Xl1YhFOcCj1rS
PP1qSHp7tyw8INU645eyDWReCtFgBxgEGBJmN1aEz6UJcfa0kfLA05CvctWRhGon+E8Pwr+AYgTO
PNjD6f53hc2fnVpoYc3v3kocIqpam9b0cegN4V7wDrLEranNv7PwMHGs8JoiOt1ReBQooX//sGto
EI2irZznjyixCliZhYMiAlyQIxsGANMyiGyQV6Mnf9+ukLouSJk2agZpj8y9aHKA9+lndphZ3wc3
AKbzeh8lP/ZCdmUmas0W96+gw+locDNOVqERmjgBFuj9DT0/TXaGleybdWl+x1k2Rogt1likzA1Y
HfkXhIg3ealYYyMY8xeK7ZXslL3x+CWnI4VCpcdSGIv+Yj5rtwBQIQR7Zr2c/QPd3bvdIzRxdmYV
I4lBmQsX2p9UdjG03PMQ0PsPxFCWWOiULFKT7zBUvTOTdcvUBdE+4zVpTNA0O/IKjAbPxYgbDyoY
JlYUc1Wyl+g9P7gPNid8O7kvbi7ANW/tgYlyb5S/pPOewhjTecJwfjSeeyC7NNc2Ukz7C+3phH4u
MZp+/x8fgLoqtGlqZxRqST8fTvsSD8FNL/8D1gF+E6pSwViBwo91+c//HdZEW8A1tCPp5OkHH1Cm
xjQfASRieBZVu4+zmgsrJMkjnmlIlZpgx3LK7oylj8cqFFzGoJvD2h6T8LvZR1xQ3k8URgNxL9IP
jKiC2cX9KP8lE3tJg5iCJ1qkLHp1YTqKBaOg1t9ma3qAkLGvCnHKiaskotzvK/73hLuJrs+IdZHj
3QJ/UOhCMSE6o9gVqpmDW+34Y9Xpkso5b0uUIBgN48Jez8mtRHLU/bG+juONKIMJZZjhxhwp94+4
djTpX7ticbGs/LLmLjhs8xZLZc97nthikAsNF76ey6GxyiXkXKrAxGk/ETo8vVgg7LNa61YIjhrW
vGl2JWkPWB0+LXZzhRtRd+Awrkht9of7WwVWs9gH+heihFxaqM/y1apuVa9JgqtZPHcOWz2TeFnF
Uo4vfxiwjB/N3EE3C9d3ud49bTFFV0ttvfFvLOxT4eNuFYMIKhJ5WrTLogdNU+jhDmD1qO5zZniR
g740LRaeWPFFGO4vqXWJmt6ogb+aYRe6DL64svJClvLYTXPEVP/BlVLZ2mRmEGfKyI3W+M+1CnHc
70YBFW4agKsr9V/2RX0gHSUOWMnDCqeVPJ7waxOVNkNaKtSHgAtAq0xdnGTSjPgq7S/0JA6aI/pu
DcXkaHWNcJP/XxOaMyKeTczaHnw04GWJb/y5qQJbXrYxqJZ/1L0UVCsBzcEBEbRjWYCy/Ms1h0GA
N1opsC++gCvlhYIF7jQo1rt2cAXgIIgVuc68gosO2E8ojg4PZNVSu4SRXV5plDia78sUErh9M7P9
bAqpqeRuyGNokdCcumfMlcrlyWGmtqPlE9qHGu1/S3KbdXb48tA5ipECEfbqNqNIvQexJsQqeldx
7bGNJj16E5EgNdZtJFOgxGbFuueXbVHN8Nx7U5HXLK6RWzWSpnwP+FV0Gj9crGUnxbIpYN/sWNP5
/vCDKxS1xRnqxqyIcYiIFzslfRTHqCqD1qIfOlWQBJsayJQIZuxDjYxrgpxRH89SpQHGPruuAzd/
d+tUSMzIHoAK/J20gdz6Umnp1KLAYi7u1dkpsxkPo/KLUQWFwZNDNLCfrBRCnAykiSBvWJspIAE8
IlUHSNDT+EcW2Zdb+CbAg0s7WbfO4pHN0ikfmABjMXseP/uer2HSGUbHLtVnVN8b1uVe5srGxdmU
IX/j/OGue0nd1lJYR+YcUTeNDByFhENOwzt7Bd3QjDD/9asMdgxDK0j30YSg8b3+O724ibcG/5NJ
jx2Zt7ZARnxEA6odntdVODvzIyzJHpBPE44gU+EHiMACExjkMur3bmwFVRLpJeO/fZZHHB1bGTUA
4/Z+gX8MknuIBBSreAdF/DSYpxK+VU5wwag5X2/exRi3aM0v/HvthcBAAak34otMK/jIgU7T1jFb
9M0zx8ocZjSoztQiL1U7deRwlpor+OPW89qhB7XzDKZ4faCgs7dEzNhLo6s00XPlm+HyQRPfhhuE
dAJlzW5OLDH9xCJDDLgvx0KUx+JQCO3uyhT/NZ61Aknspi6p2MHfRmqiSUxuCxuiVpUIa4KX+OmE
0CXNj5glICoAMaU7BOC0LbAHIHiA03fOfIMTa4Qu4OoYUsMg0smRw5nNnqz0wwf471VvTYZ7QOeA
3zlfCfZMkC1H5s9MC85QD6Br7IHQiXGmLKGnTZ1ZxbC3miA6pTYNYX7sQU1w3u5IrY3BgkXlB2D0
u24gKIVE7ngbeS9jhGrlBrqaZ8LTvtsbkkn3t8W7272wil8YKBMZRmHPr6q5veB+HNa6p/hwx5eb
jiakJVdc8Ase4YdR6LMLXAnxPO/6K21Uc5zmzi9o2BEb6JMdZNBrVmTrHeVGZlsgbkZ9Nue4kuyc
AurxPQiTq7MB1k6dwG2Em+gz9rBFndSprW+DqiIZ7TiuBbbRxJhO/QBHK/FDiMsLwny9jNVchSTY
UU8Z79Pq4CkQv/uSYHHV6yifTj2KsjPU92j1rHamwLPyvqWaDlzAvUIkqUOaxI/0I3v6WfAJdAQl
CQb8BUpp86m2csWgtC2saf9wQ25kYAw5VF2p7sEJJgUau3m8nwMd0grXptJ1JIPlmSGxr95T+u3t
SHXt6w/av3Yj8OIb/+m8GkNVeMGPpqkvYGaC+vv+tRW7sTcRgAyArxdGhzaYyFARoCWTUxYsJSQc
wkFvtoF6RsIMIkWWUZxjpwlRjaiKir/0hjrvuehR/gnMBbSoY/LOitXHOchayBwQ6F607AJjVJ3z
xvb6tKW/+6vHODGGh++gQcbhbUQfoHc8tnVIhCp/VSc/zdte8Zd+9MygqRlQWQHLnhHunDYHePEt
DQdDFiEuO0TM4DbEj7APoBM9l/CUrLPwXsBUpUrrPAs5dJyR0Ug2DDKV0wkVZM6k+Y6iI0cPkI1Y
Te7PJXdhORs/Q/mirJeibFFzjdBcq+plOLVjX2jnVjFavSNSuo3js2hEMyuUgd1MiSXjPddE0Xp6
7QL94B6pRWdpVuCrUbxLBVYWQZTVGDk5uDC35ZH3R7rY5qWWazFgTp8SdjqmdIbP8rK63rmOb9Iy
IEp8SZS5zXq+blFE/UcQmzkS6DH5vPAeNjqihQ8kb3aA0UzobfdAFS2/BwHdGKm862Yasj5RgZ+O
pSLr8xYSTYr+EtPUApGlZu2wV+67Km8DWjJyhlUsGdc3Swy6jVnBKaCwW2mGOqUXo2WPPKpx7Ci4
dOzpGAzM2PddEG3k1tms5jw8UgG2Ri2uwypOAoGfuIl+RBbLRjAOgSVKyCSREx/teoEdmzgiSDny
ZzP0+IeZU2NR8y2o4+Y4IGGFgb61rOLW0s3jInxxsf7dXbUklZD5b+mgNcnMTkSLfXG/Q0eStROh
Op36ot5/PHEv9+Z0sDjg1cIXr8ZnhfXk5Z3nrdwRJlzh2NT4d0snumLd4CukY4wYqCisL2aMdaq+
RjC2ARpfmd8LgdV61pDqKw59scWl9eDFGidtf4+CuP+162k0sdcVCLRVS95sAdP3CzBM5QSkW+IF
k2UkAYiEWL2JzjpsLwavMb//XZJbZ9GWxafcS4DtUxfoEWm7npjduLse7yKke1fMkO7dOggZ7AAg
FZHMnkaFuq4fUsQfhH3urn+wodwlRyQ2pmMwenkSL6tgOIx3mnJrVVj/XoqJqkFrKWnSJm+Tpxnn
GCiNzxYvK5YR8vARR7Y1cIHhO0Fcc5zfb11ljOgdlH5Ej4hlN+3nWOUK88PG4nd1yamjG7MAUE+l
tKSL9/KlzhYE9jEdrQf26HYbDhX+2DrpXkhEOHrMnxecLRZidQabeXjK1Kz/xBs3uD59pf9pt7ce
jS9vfsXlGSQZ4WaOn9qptuQi//svhDEIxQG8MpVcOXvrftG8sCgpsJvba+wApQeKi37XkwTUQxHH
o4EWRRc/ZROJMPkmmBGIEyoRIoRtFIb9GsTJbzuK+NfCHSg2UoJuXBqZ4sAiPLkuisup8RV9CnJp
gWr06QrttFoNEDPUF+lNU2lH4AzAjvQy0vgpGxjP5X+NmJaFlDqbx16UGzlRvYHRUP2dAYtshVt2
2kpWQb7K6j2jzRV6yntVOzI8WHFEAcLuevPF88E1/OAxZAZVXinhNgnYgfxlO4wpVfULl7Wg9AR8
o8V/yIBlGkyE6Lpw1buBDmiXywU+xvbdusuoG7iOOMLG9l4A5PckaCsIj1DkoaiPltIPpdp1LO9i
qiKINkZvZ+sGfcMWAlhHvJ4xBwrWskNqKnV5ew7pqWy2vkIGSh50mGPQrUoA3IhdIKLa9/bDQ1k5
hKYxqRc+sBdc5sD4JL02vXWAF/5+GTqcxoQbBQigY+mtOjFgYB8B0q051I1r0XyhcXaDXwklep+I
ZlpUz4gLi2U/QUJgOKXr2QE186pAweTbNRduO6Ct/l4QrU2DWPjdXj/X4QGA2uvLtKAsFBhD/MBu
JOS7TB0W8i3xIondeUCGwAgY7kxAii6HUg/n4tWJy7kd7r0+3JUf3jfTNcxkIAlgdaDDR/d8XHUE
M6I0JlTP89AK1yJRJBcfuMeK+jImgpAtsczE+ZPoXfKYliMwnHD/HkkD9S8yQiCCcH3jn/pBY8Iq
2eVk5lWmpzwpEi2ChpjSfEg7fRplX9rM4DOd9b4Bjsl+PhaJf7QydVuS8/8LgL5HtQm8cUsqOdgi
U/SHd96P+9MBhhtHlypUnTSuhFT42iLrCnOmKTf3/jEVAmk11yzIIenV/vzQQT7OgrOvD+ZoHsgY
1Nhci0H7XZUIgXdTPkI1ErcBDjJADA4eR4aoKN9omq+xTwHOuIpGeZuxvgOiQvwIK6zIqltg3WhO
LXckdXWMV0cCpMXlqMsPNhLzaFeLQu91Rwco+ShfrCPGjx7EqWwAa5tklhJX1wYHf4j2mUMLGWiX
UMO162kghvEGbE0Oac0aQcBJJ38wzZMzd5RsfyqjSjdYBvGJrjKzgOETxuGEdHfWf+yKHzSqwsS1
XatntBJ33r6nZ/ipeh1nQqnlp5kbmtx81W/rQvrnNCiRtWk6h0P3Sebhoq2OrobCJUMqLs7p/0pk
0LoL2SqQ7gt4qlyPfRJYUjtMTOHW/jFVw4LU5zg1askv1Rq5R54q2uuU3eDHRniPjomiVdoXBdBq
Gy+PCmjVX7wKxwHU7TfLe6WDVZnmmbfE833lhCNPSBtKkWKAgdTBHbHD9W5lQY+QJrZXRbw8JeMX
SlzffDwMmiH6ucxHC/PVv0ykNK3LPy8z7TKHfx2apb15MGy9GENJuZLVkkdUzPavktjqKpBzqVvV
/xooHGRbO43yjwg+xHLd4iFyBnlvIym83LnaAMVNtfE7HHGFFDuZiNtRjzNEL6VszPNNamEcXhqu
6gQgOaYAtJN3EdOxYHb+Eiyc/O6bMA2DtdELysMitp/JM8/gUvcIWpQ2Bv9Ub3v+/Rr4HBwgCiSD
buY3WdXKrDVVW+kdnLvI+WO4qzWhZPG82nvjcT6Qqv/k6Ko8WvU1H208jeLSvZqzfA8qcukiUIgz
TkaMMOD/1nxtKqIZRnOpOwq1yFHck8POhCQO5rltqB1RRFB+jGMe8mYG8vqcovBOMyPIjAUdOpJK
/ihS7eZHKavjxKmj1PYZI8JMv8KCyn45sLjq9N3+pVvt3UM5oAsa85RKkVKx7nis8lkiifBn+tln
leZjZEH2YrBY/WO461n9OQ45uH1B7yFtaT4uXSoN/Zg7NsNSezGXjNHvljV1S62zswFcQe7gH+Ix
mpvMR0EaUJX6yBRzEGlBBw2gfRYvP+TIlge17I2Tc4eGsyF93DhJlgi01lq+ItGzU9MwPIoRZ6Tm
DOIJeE5Gwq8z4pZiPFKovEhhOzFGcKcy5S8FyWghm2k7pMyJqjmPriuz/nzgM8IMEGX7Bki6vGGV
+Vh2wFw7tcRtVYB4FPDCuXCayvrz305YbhzinfxArA0sDexdInSx8tBy2efeMVcbPwW81xn+EDPu
bajMAUmY7k78t8N+VC5LtTrgStKYGkMLfl2VILotvKGRRX/XW876QZhQTXoRbIIyWIGfOlR/BBcW
/0slFKXDtUmGDLhwWk/33CsppbS7uHg5vClGfpzJaBtaqj7tGr4kmVmgL9GkSLaLyu6vB7FGXJdq
V764HMYkMLnoSPuTXs+uc5PwOFSKGgNgS5rJxaoRR2+wIo6ArFQGUQkvqIUciiJP28/izehEvQnW
L52qSD65pAhipT6BWrr0wgyGmGmo7+UEbBYVdorpxY47yxTQ2k4p5Dx2ktbyiPeKFtsM/OLkRsUf
nMgnIaKX6JwxCsFWc7iayVjdvwaPRp4g9PQK7LfN39mp2zElldHy8IuiiMErXQvAnHJv10OWi3Y3
dvJyA1aI2oP5qY46Wo8wH4hSlgRQYJb6XHhi2FFhk9SVOv2ow3rjwQzAvRZERts6ShDe+smovVxj
KRATAejm5ZeUbBnhTi27cM+3t2VKIK1QCkeyuAWmqo4G8KNVatwIq4uzO4517PHfcAcxFfdXGbIp
SaSofZfEFu5LkWTVgOh5dyNuNcTTMb/u36jPok8I29/mvelu7YaPahCMXVxpNcOTRMPPK/XIfG7A
RVhqxRfTKoWwB+5SrGwzjnDkWIZNZKyLGhYKhyb4raqjuP68JSu5gC+yVnROPpc2r76wWVna3Cb2
+67bcPPqMVBE2ysl90tJny6YzLyrN0tOLzaQi6M/6L4b+bPdq9i9R5D6AFg4psv3X/PfsoFHeXH5
jQEyvL5q90toPZtmLF4kzkvPgOekQUe3iM9LEZwEJE91gMqr4zkzq0A27E+y7tYasb5jx0sJ9dDb
uM4J5GltkxBXtMpqp71SBQd9W+o8jHc3dcGVtXGGlamaYU3S1mXybys4cZRQNRKm5umrcANfamXP
/8Uhbvcq56W5mS3PKOMtf7Y/jeOp1jw4YTx7F1RLaYpoIzrVt+SKskmMoNlCuY42DN+7f5muU3yE
NsOdpeI9g7TGgxivx5wuId+KplpdYoHkIz5iOks/QOsigKadhP3S1eZEux17XWeC4KejQQfaMZb7
gypoTAhm+SDUs4cnp9PxbkfugnF4UbYIjN1ptdPoQ/rPFFXCHXqJd6qTcuIolI1XNFzuHejp+MVG
02LIbtzuVN9Os9O2hGS3/4m0pDaWvoxR3S0LgRP6zVoHwzaJX8FdiQlmsqVQmlhcByPc+8OhFfc6
+lmdlxEovkwzUj7Dq3VKdhZH9BD71attxpByu2Ix/nvUDW8EkxNph1C7ezMahDX5/PmGwJSrjqSj
iZhJQig70u0TKRQGazqd48MjjuvKzgbghorYT8mCzIVldCFNdsBx5Jd3rqSU/LHapFdH0fOus1hC
vHycoVd9RyYqGxNwf8BkwuLgrIvTaI15qiA4Sh01J0qe12RTn1n9YaFNIOaMfUlbcluETdvtEUfe
Mz2zdubkKVIRhMNd29KzmyTGaMq4tS3/oqqTqkuAXr3gc0vTafGaJVGwNqrsVPyeG879Go6Z5xHD
gGNfKef3KQyxb7+gBZevWLhlE2ntTSNXc6YEnpw8VeeVJzkhvNYoxaO1CBdUAHb8h2teHI/1f+L5
uGSUrx7w7348jJBphE/yd6+iQn3Y2j7ltuhNWyF+0QkGr8yYnl9B7rzpU+0LluTvtIgtM1Hui8F0
g73TbQyUsPT/1/cQspqlNFqzOoHHJt3PIEEXzs1UIMVBHqWsmHnFfw6VPVGUlOOvE5jIxTaEw4rc
j1uzTlauck4gX39iqq2zXGDyMAznBdbwzeNR7/zkmGVh+TGHFjl7j6ZTb67BBzEFCJRPwUi4ONYW
GWXcIaowbZuDHEIfTnLhZDXEZVygQd9NAsKJFC5Po4058fYkFtIHjKkty0l6M/SJtWpTZFgf+3HJ
RjapDibdhnIqqvHfJRJLeNFA5JWHGD+D3kWr9A4g8Ila8aq2UFgCRgHVogHmLNx4PXa5fC8o6YKi
kQMoeN0+9kgypy3BmlHblxlrAR1HhsVET0reZzddAWUMQe/8qL4x9XwfvBeUMNq6RljXUVJug1KI
MYXvef9I0oxKY277KmmEpAMJxrBKNxw+pHC2KKm5YTObjCUCp4DnzdPQmOTAlHoVXFrIL1JjJT2U
0piWxDWj6Ub0/7C2cW6PRF6H9zil58FP1hQ0lz5ebbQJXRdfhE6ZuzPrbZUZHuKxn5o6HZveYBfT
5l32t15jSwT9A32teqH60f2NoWXPCp6rUVZ8IHtw08gfumUQcaGvb1J+6JKcR5UoNj83EFAISgyH
XDXie1yjXTBDrDlbSnzwX5IK6tXfw0+isTADyUadUveoXp25sQiO9s7LMTBWyDOesZ8dORsoC172
NBYLSbhng/LgKfnlXeheexU1UhVM4rxZ0Eg2x/Jjf9Mn9Oo2nO254xWmkycanwOhORawMIifCZS4
3oRWAxE2mOafmlepZRgBcufXSiPQHyxC7bDvoWLIF7nk51F3InaIEF69sZVbEeQ/WnRIpzMsxra2
Mim1LoFPRYtC4gFpwzvderyrNZeAJ5Zfk7B2RZNYzuRTFTlVUz7TT2nnwbr5GcZWKfEtdYdxjwol
bLR82MukGz4NZIOf0stC4c97miWy4VKmYG926DX0KeHsziii9HSlm428UU7D/pLn7ZjUNQJe6OBE
yEaT3jMal+fnHHnlpsCwhMA09Dnry/hWrd8N4bXMI1qQZDab7RpqhGrRcwKFuP73sMSOByBjKU5Q
upzI4bGzzvFKX4RFcLq5k23XBAoD2W3/+eGfVsAG71+0U3gmGe5w+wjvnrE6BpjcaeM6m27536ip
LF2qAGcmhc8uWb3DLMjqEI2fhCYuYnBNM13+6Tmg1lbz/jLFOWTZ+QYi0XD0f8QlP/u+bfctSn+p
6ZeIBIQq6sej84rNfsV0IjqsZ41+GuFn8uLaJJZDcY0e8sPU2crqSxsBYblu+lbhA++r8uo3uuf0
IMQ4sF338XVFpq54kHWbikz4TkafV2kZ3fj+kK/gUC9+Zlh0NwfWUocYcHcE/lZrljYrKtEkJETV
vPPVQ0KSfVmlMc+Gud7xx7T5J/wgMfG+l8z8tNbgN+y/181XR8cqwtruWOkVqVZNJSeP4nWf4Ci1
pNW1dWNZS5gtpBJfJ6i86ywa6nKU/WnjzkdfbdpDiglhXQufONKGrXBj66gmWcfhxWSsZ83i2kVv
GK5S2lOTn0er5aqkU/QAu1YUnO3c0HJHDCHZhq09+Z6PBMmgm5fLQsJFLI7noTg6YvlPbFI/NHYO
+o7F4pZBI4k8RiYCRnl3l+c6S5cgor139NEwuevw/5eZ0bn/naqqdZ2StXXfZgH3C5pH4u5SZYOn
u9i2wG3IHduZzOV5i4/Xx/48EW+kRGwhrqdu20iXIFFaKuKelheg7t/xF4GAb8dfjulIITVwF+Zy
85k/6nXkS0XdDbY6JL9vv25aJGhCpIKyTGENrSRxa40KTepB1rNB/47+uDuHVjjWPwPR8zisTvdM
db/piQuWgJsEBPcWP+6ESfS1afXR1Uu6Dm/nNHmsA89JKJRNY7qNFxKF9CNxzfhlPQbTfA8XyFaB
hsk0/xDlGzZ3wAWE8ow2UUU+SS+Aa8180aZ+24jIue/O/KEbLXAh1ZfujQHhLhZfCzYqid0yLX0c
mE/cLwu526sNoFEPOEuWHNMdpiB1uhYhOtdJ/iz3n5KxIg3x83X8sEmmPJppptKigzOLfJA6Spr3
KFJ9mRzFB/IUkZCnUU+Y23AWAFQGMaBymNZhFoTADXicXjIuBntJsXfTCW6WmK6SUKuG6VbgcqC/
uRVxKGkGXtDzBz05zMe4qKoTZHsYY6hpaSKfEpHyYbCWlMwDGQcAhnTZMAj2s4mis21ivyEcGR+l
yCooUuSRdjmrOOR1SYmZUOgAbeZIzfb8h0thABlxkFF8CEgAu6tKzCzEZkAR9XTTb2I9EkXjTzFz
cRoosNiHUpNuWO0VddRJUZg1vK1tSpQ4JOe/nCu8Rk5iv3fAa8gPznW4AhkLi8rdwLjB03EE7Hk8
02afdkFTmMMgejJhEGAiF7ZWg34xKlBFKuek2GSduFELvzSpOJtGIV8N6Zfp2FHyJpSAwy96OctV
ib7ryVMTilB8Gjg5g2lIfWi4gOb4cMCQaILjWQt7r639iOdTdmuO8CMVV8Rtc0FnCOUORW0TAgmp
fSkD/ULX5iKYQuRxjsgg0nRYYNl5G9wlTtlPsPS8zGniOeZmkphy9yld599CnHlAwNYLcs9Nwc1d
rzwhj0la1BDfGKCIyiOBghw9AqPaavmbD5G9mKoGnKN15WuzLqXI6Iak8i3fAyBoLK5v1u5Sezur
YJuG2Nk3Nq9ct4rtbaePR8IbtrsDG7tRN4wZAnrRq2hmOEFc7/BXPLWRz/ByRMD+d+hu/QD0zNCz
UYJZADIJHOecGdFg6mH8dQZkPRmYDke9sVsvw+nD3nlgtEWNaCmgXaQrStDdqw7HAUbSr/h/vcP1
SEmgqdVLkhgv0t5eX74/3F3u5w7/mVqbwbWcImLXcydm7HCfswWnpWYGq47EmIE7TUwOEtIB43XX
B0HXtyVnLEUI2alOqejW7LtKCrHBWYZea+ro26uX7LY3JkQICvYpmV/rtDIGzEnJ8qTDhCzhti6l
EUGxa0KCy1jfVFIQt+nnJ/FxGNCIrPqh8NQjZUtyhQdQR3tyMEFvi/ej2JdY9LiM3H/x9Jk55m/c
6Quch7PGQcKe+hxUq+3wrOCm8vVw9Xj2KqrzYQQ3iQlz2yFaSGNcWjiCgUqj8j39w8SKPCIdOa2L
sy0Febiqy9/2RIdCIFxc6xm6Ml68/IlMvknV2Jk0TPTumy2LFUGmR6JCI5PgDcVqkvc6DnwT2+Wj
3yiZ1ULGTKgJeu1ThCrJ2kG7Rx7YM8eIiihWxSROof86zZDSthy3j4tUGCqzKKuHt0AIO4RDFMhp
dhZ/3u+phmr1myjqCfd1tz1iDMgF7Nzuazv6LihgSPsM6IXFbN3Y5DCaubRplFR6TcS4RI79JOhb
Hq+eLYnrW+GmRss/pBZyobhFIw/9JFf2MsVuLX1/TMc/mHa/OhQFOARPdeZlzoa8y4Ukm2DDheAx
Vj1StZQdTBK/UJi7iloY35p7VqU48NPHjGBnvI6oUuDa87zAb8ggA/hUieqiicPgBAN2cAXQ1u0e
tvLgw/AqeKDGw6LfOzdv4VGKSc0orcy49LGcFXEDIhNw36bPjo2i0WHJUWfPSefZyWRKqXoH/oha
zXWc7b6F9MbnWfmNi8tOJPUu+fMvbkes7PpdxLweLH8MFCwKCYSQnz+Vh6x8NGOnyOlg62RuSwrr
LGew4Gp2a2n89nLtX3VI7elAeaKHAX+dhUmlPuBCjdMu4rTGd1q0WF6o2YCXwfZuUfyeQlHmCk/5
mmqDrjWCdFc/lAmoSkbppdlFE7Tv5gS5AcgM4tvB23QzJlnGaI8aVAHBDm3WYpFKJcePmPzYU9jr
HMtTzrGPvi22h1Uc3Q3ViqOFAk+wG2+cOZW1nWa27BuhTWgaYq0aXyHFYN9MgQ343DM9t0XJO/pC
lNNdfQIEBhy7oNS/15k8MKYIrW9jsyc2AYa77dfEPYZC7kH2UorxYMCcfvh+zC+pir7p7B4JrxP2
7Sy57K9aEIpivamWQOIcvB0PpO9LAEpdOS1edlEjIYpm2jt0DZXD7OKqwuqdfKRL2KOOouvh5mj2
yC/vD9uczJB/PQ1lXvhXrfhSUZ3DyqyGN2MQc4FgwsTkhXI/aCE2MwSCXh8Wy8Iuy2LbZglPPJ9B
IvWGCGkKOvI53FMkgmGCI7f7T0zPbib7bZSWLqTPZDNQfpe9DNmEJdwYNt1/X1HBsTlUzMVpdtSL
ua37ZeeeaJjhXD12XG8gqQzmsWnb9tLf2Jx+eVBQwhFzYVIO064+Inf/6oaaRm9O8JH/1pSHI/Cl
Uk0ANXQqgXT9Xe2iFjFjGgE7Trbw2jQMWSGQADXO5Em0gJt78F5IeHE03QGkZcHikAYdjM2e6XAX
t+kam9+tYWuAThgAAOOSHP8s2PMDhB7MulAbW/g0siDDj6M7UXS+QG1ZtqprTSBB+iV/ECIBIMVB
YhsvUca8mN3AUJ6UHcMZljGjZH7BqtryA3O4eytFXhh5PNpw1qEO58WGx40BcOs+Kb8nZBd+7hZt
9HhxpVIC/U//lxUgg+VrcTIjVI9aacfZSxEjTECA8hKQ8+T3Fw++MzYyYRacPOSIHhcqf364d9Wa
fb/y92aXT53BuYLmM/oNhCANMDLAcLc49uiK5jGDaZks1JlvQL7/PEWHOhioJW2GVG73OFgNIZUE
i1A+G04hKG6zYXSQ/R43/yTmHKNYDnsCM1QiWvGZcYUKsG3ldpkHACRbck7TW/IzWXS5gS1kJRV/
TSmXLidPi3BciFih940bTxx1GIZAtgSDqHwLEJIAhsDWFoEbE088UFvI0SQ70t7OgAv6eFxaGVvN
2L1nmMm6RnF3isGyAg9Agwi8KzQNvY2KhEFYNXIoH+l0naQbcROOGkEwz4rZfgOEfdNOtBldk9i9
KI89vbscIPOYuZ7USsZulWFx0KVxSZSmUKYAVEHehAEVuLMI3eKrIU8oDhvKTA9Gg+2md/f+pInS
2oNw/rRxC9mVvv+XvxH9GWCIk4j90B5p8mspFKpKaVk7LPrJZ3iLWZ0ToAVZvWx42qZaeqVkkVcw
u4Z69cHqBCz2TiUVjSuZtfFtFru2u6BxUaWJAbPTDGpi9AYaTI7VJs3XM1ylSdC8+OpKuLYe/Fyf
20gUl3hAGOJCCcIDxg6I4vUGB0sbDSIRkeVbc1tdIeanc0qxR77JkuB4uPgLNIbW0h0yh5em7NU/
I5ZWQk25n7rnOkU2grzKbgxTeE4CTcGYhBShWOSfjWhrGYhxs0BSWW2oPOcfreb3u30vkW4Zg9SK
ZSi4d6rSIDoMC4sUVQ9uWjCMad7xwB50ifY5N5cqtx/wIGBv/NUWZnhgINt6+8CtDHMZAYQrFrkC
wVNMEIR2+JVF9Wa7Nkej6AjzETRM8xEa7X1XsAZDlaGpMQUKuOW+2jRqaTxiZM5kPA0biGJdNQsk
JsUKdrpsAk/nXNxFsprvpme67vuoIRDDGuVE2I5kRavYnmxoUFVgXXMrHZRUmYjHUCywbFre+yvi
Ks3c9PMAl7apY78BZyZWPbXnYvtXMQAQedyWJIupBbuHYBiDFOjrRQIy0v9rHHycDD3W/O/4ArbN
U1dVfjpALyBAQdsV2GFpNC1nd7jUtfhQ3QvWeY0jJN6yJXT3WroR0WkG6uiFp+j3jsACcvrQoJAV
H22X4LEuMCXCGK5Swf+qAAaPkeYWnlm+9++izrT9zjfHJz1eOe5acNmFlv+vyVGB9KiM49k8JuIV
mMW4OPnOUVrn8id/Csl+ZiRc0ALMHUXK4i0JU4/k4N76hk0Bl8LS0DxrPNWRPn4J/OjDptWh8rpX
Od/t/eiy5wN8x6+Oao10vJqQtKzI0qK4ex43Ruy5AyR6iAlGWw3KTpAnoMGiFRDme6yqtkkZuyVA
+0hxxmwFX9BJo2st57IQPoJaxtMGp9urCYmqHqSyv1CZAKPY/9tq5ykUwQw1jMZgqim9QpKThBvP
zkSZFhCG85Rjno3ZJ9/nn2nrgVjO10k6HUolwwyDmBV+HaQiSjhk9/qC5hGKL9DJo2gYJ3oNndES
MAd3FzTDUzs1097TXsqJbh7fXieJq1AzHwYRiwdn8c7ZxH7oGAM6uK6nwALdAT0eolKq7P9UCdmT
XgwdRktIVQ2+tJjJSMA8gwA2/5Z/I8CVPRHamLMp8JKEjnR+WUNuZy97VFhtSelpTFIvk7p6F3gI
4x6j7t+5v2u4eYQLEA+KFypZyLgfUIIFCV8bVQwtvukIbs7Q4eOJ2TIaAWrb6i7w47kYWFFMpcPE
Q/BvoSUrW8QNuMEMnIHZUoX5kNOzuEHujYclIJhRSNjwT57KXObJTQFXoM+gic7LzEaQj3l8lCWe
h5Wx4Ao0hEt1BMxqm06mc5dB1iXo9CWcOJ0EFOLEoBax02wTITMmx16l+ciSMVBer3Wz8ffjHPRf
ubx89cUDdX9nEO5M4em9T/lffnfr2STNcSkLA+K9X10SkdnMX6YX71F8TrH2vdOy88d5lC9MixMs
LThz7QxNYB5BgCojAA7KSvMrKR8qtiwVxYx19yiL3cgymjZ+75+EfdqZiFpEsY+0K3Cu7fDtvxGa
mBEF9fYrHyQSo9GyMIeD4QUOY1L/8DK+ct/tyf/nkVkrKK6C07oPq7bg7x4qtE68rXauMrVBOHrd
mj9pOSu/S5uDdvxsPzoaNQNiyQYEcPW+iN9zfbFkd7oDZuXtRQJauJeCIR3IC/YpVwrp0EZc9h/G
BRVfVAUSKuTs80Y71Ntr81OOH9478gPz5MZovymwF8wAbSTe7nzLWi3FVirnoR+d5MPAbBpyvxTm
UMWw4hMKD+HBTLBxh1U0vRW1Zoe3A608rX3DHpbPfYbqlxM85xw4MEtK4EnzZ256YYxA2EzmiyDk
w7uQnKsDOnvUX+Z8+nigkGNOhg55e8sUfUTOrUvuVEv9annD7oVT705K+Ofg9yU5dee6q7EtIjmD
rxPrSHdStCXUIeK21mkhgjeBrxTexukfPklbdFJfCI43j8QJWXg2MQ8dm/l7kuJhnwBHBVX1oPDX
eMjyhxRe+EiAzLgL9MldDS9jIDNrIrADV6YnDdyjglFYUVnKnXPA+znUzekHlX5RYQhZ0/BgOwDG
ja8Tl0yIEI07npDSlmma8Svo2eS4lGrNSaVUN/Rc1IcrAzkPj8Y/D9q1qbIjgJBiCI4Yhb1NUwSw
8Bp1GyCG4s2cvxPAr2mXN/qI9aF7FQkP/nut7Fs8VZvsYnmzBuzWLPhgoT02GJavSuJdifFouNTD
V6h1jAmRKN/0J/JSHJJ5C5/s/07VELYGpkhU59IIMDWZu6w4bb0f9zx4L6Bq0xi2SC6B5zBnIome
wKACv/o7OJh05vyBcSJdFSNwGKSjzet/9spWc2KNRqr/XEthytgI5Kbx2uiIqcQ60t8XIfZEkqNG
ewxPjqq8+M/w9QwtuSa2Mdp2lQdvExzv3qMuXzG9y9r0dEKGbkTOGNRIBe0eyj9ZKuec8l1IsbfO
4b7Sj735rxLbZkhnNA+YHGXse3kq1BvOwxpQxksAd2lU3RUePQknN5nPSZUTmVDXiHZKKjEA11zm
9jHOii3L6nusKMN5N1ZcCHy0My8XPeauMMCsfYSGPX1dnHi3A+u0irRx1gUMxpkggHcf+wXA6jc6
hbOGWFoSY0VB3Ri66Xp+ucGy+7GEV3Vv4RISqS9G58IinEwCR4GvHVP+/PCgjN5eFUqAE2cfp02m
Wlwt6VRjzRSohHPwsVHMNYQ3Jgxq/SiJZVl5HRsVr03pt9U9VpaLlv+lsyixQ/2DjFKwMXx/tkAm
BYSJiKNnZHb3S6ve3OKj8pkXUP81IFWYBdk1Y/oJpUNcVvM/+23WCWNyPonMw1Rl9pcqaZ7gQfJB
YaZamFbmiu67b9XyGvd5GALb+jzHkLNx/ltiTEVyjiUZeCr2aPUn6z7GDOvgGGqo9l55lYEcL95/
9R3iiWWMGol6b768su119dIey5hm4Q195BdELgm/CxtK+yyR6JWIy/EVb2orf3C20iZxg+aZt9gL
X8TnWGhhxTAPvi8wLOMJ53oNpDDhgLIZtr5twldLAKX2MXnQREt/YEL85eIA7VyzrC3QhpumcDU7
Sil/h22Xi8ooIxCeq5VCiyAt802OrkQHT8JBisc2L+ileG7wXTXFaO5jwaOsW+MsC1zY2G/Eb/dQ
kDbiYXJisswMccYYP9qxnYE7AQc4kSe8b8k4rf1cPwmyyEXoyzqVLbUY7SID7FVcA8YrTuFYn8TE
xEipSPr1DiJCNJCSmsnQwyD7qJodnyijaYWqZIKxFnqzsijMq0gD4qkvhYWACF5ARsV/KJOLLrA8
GO+pq90B3VRMQXscDO/yxsHY93xHDS85/DrFq9cKy1Cts26cOEN02/z0HDbqNN/7gVH/qDsPGlAT
NwqE0oSCdN4kg86pVvVHse7lTFoRE2ZE0xDe6pXTSgEWHKqvnkBeDdvv1zuiuOhwhbbaTNNT8sEJ
u23ctS221e15fOZAfb2i/9ps6TMgJicUHhCDoquZG4epcmLddywKvXTh4RvEBqCateOQIsDLbEdY
qyIFyomZGxDaWNdcPFN0xpwnCMjxDP1yydHt1vzoHqjUFpM+l4n3NrAlsSmatyTijzhjG8vw1gD0
EjzAB4ZEqrZUducchghToHJzstU/lfm80Jkuz4dWpKbljq8xeq/LWI4KGb7eLAOB672E7H82dR/C
BIrL+ZIGaaAiWm1SFDh4wa+3IeOxSGb2zzvZiXdw1FjDjSP/Lkdjyc6AuABXfibFtDRCDPLNmRTk
TeUY8zVr3LPavmw0mOqkkC0A5jxPATKWdKnAgDl6YW7Humd3Xs5dXX2CeG2yzCiIwF31ltFkanFU
ARIEuSEwuAW1DNN6HnTBHYKcP8pvjgw31s5IZta/J7aB4uM+nIBz7uRxBJsdIWYPaZafTB7phiph
rbVel/w0TsEJTIYx+St8BCVfEF0HoSISbfoi/46exgYh3OdWPPaue9l2D7BlQjiFjAUO2X9S+HMU
DrWiXj4xc4R7Vau5N3ZV4C3xq60ZIvaQ4DGajqzLP560KXx3py+6aMdWTGYEaTqkOOjZFW6uh9cY
9QR/0YSxLpzc7GmukTUhKOZKccLjQa5F4MeBySGzDIXSdh2rWdDIcBtMpspzOO0FVWxFV3s2ZIB9
bGhffPDYkO4BAxZDcBKJgZgO/6WYc26qFyWveHlo/g2ZxCSf/tSucwWlUaKiJgGD4Gu6p4k2H6xW
D8gazqlt1I7Rols2btIkRyiN4DQUxoK5KAMZssHZcHuCn3NudwAEEkublzS/QpyUiF62yghz8Uh5
2E6f0y/M5lUA7SJo/VKXPbpA9xtEjgBcFJ2fVyW85xH3qJS8LXdNidPMsuFFX8JzlKU5OFPOFw/T
cVe/P3owuHMf6nlwSTSrVlJ93CFshfSIYAwo+wzVWO/3KrSq6z3ZIgA3MedZLbgx+MIIs4/dzNBh
LHXh3EinxqJi3RWhrJcAZ48pJsXxVQI/srgh3KUIXxnHulP7+YUigT+JqaW7vpPze/kkSUdeTLci
fXfVqr7lqXts5Adz5HscaS+bqCntcJNde3IX9qK1gJ7mtLY0Wvrxwq0qRq+WdZJg4/+qv2u1ovWn
svL2HSCbP/Fg1wUI/0pvWYmpFerirwQoKKOeDLJcopVUzkrP8OgU7OdThhzx5ybKfc1jD4qWCBvP
Op5qMTz+yuSXeevqljR/y17WT7QmOv+75GNdbT29WL8n7/NbFNSITMfKY2BBLWC32EdfiKlZwHve
b0SD+ZB1E9zzWMfpjhhebhVWz/jCjlIc52Be4GjvL6cJ1en6U9jRaIS6v2ABQ2ICwj1rc504lFb4
+ecnckuBIfqlJ6sRO1CdmgM76AyYX9ByAGeOlyuTVF2z3uYnOdI/DxjJb9bwrqOnrTr8Bex/QM+j
V1zMxRA38G36MSZr0PR4cBlqBiAPgk79RTAtwv1TzCYQGagqRrH0wbXAGm1zbNQhJTCaY4x0u1gG
bz7+IdZRntrvH++0fvmsFVHNx2NyuCBbTUSnIrV9Cw3bQJRlHkXFQfQmZu5SHtKh1dpt/ChLt6Hl
3tjNNycnm7Qn+Pmxedk/KflOo2ndGa1YAPeL+t1hpqI4S3cjGlBdcH8YrfDHQ7jghDfO7nHphvpl
iOTPHh6f2EXYxFLDZjQyrQuSgX5Im7aoYReKPawTFPQ6qXOugbl+LLr6ViR2yH10+ZKHQRKs2SK2
kvPkJ6nwwgygG1W0PGylip8p1A1m/o70Qrwow/1JcIf9YeqI2YiRUoF/BPVKlia+A6cE7G8LMdtY
amON2W3GmCcaAqg4XTSsKko5Wjf/0UyNv9SfNiZxAUqhRaN6rpOBSWrS1EE/whE9s+Or3FEEw3r5
9K1mOpL3BG6F4GaXOBDB+hn1raVWd45nZQXmzdvAMflGwL1oUwbH0w5JLpUVzEeQRH03jPjqK7jf
pnBkuOC5/wpdD1CK+y4sN3S6CgJuh+Q23A3yQGBPgEKiOrLT0ABLrP7vpDBlkIW8DFzfd6oALPSq
5okYnazdaYou8zWI/HhYh9YLCp1OwL+1x08itCx99ro1YziQFB+nRElHuTA/2QlYqQ/ySTZEc56q
G/jB1bkSy7OdGivMXajlKvkbDWyxctuVWd7F8a4N/vxzGobsf7FA04K89FcpqrKbmiImMmOQGB2J
jH9tEhpt+KL9WRzrQwo874TUZi93Z3SBOjvr4cTfnxcXY+Jsl7x6eqJEPLjjuGoB4L4mWJPPHOb1
AhwNtYJvB++GnV4/Mt3T/F1v5d5vcXkLg6rn++Ec5uPPR/9NsWQaGFHmlx8z+nhKFO+jTw32PCAz
LnFH/OTSiCotBZBQ5TCG33tE/6D0ZLkzUhCJKtjRaZ5DERD0egYIUZ24DHuATExZp74DWWELK7QR
r2HBS8mK4bQ/nbxO7ZEn3ZWTDwWOkQ5sHyCEx1mlP61trdjqCtIWUNTCKWt/AZCNVqvx2SWAXxxR
t6oqsg1IPTEpF3wtxh8gaIEY1XsO0F5D6xagmbhQOrRk+iWIwpT4xf/iFTdWOlipvhSU1Wp8v25K
iEW5T2rraqd2zx7ttd7EKJWCP/k1Tc0pM0wbT/SYqqxPw8sZ3beZSEPeYkuo6k4sAXS8v52S52Tx
UkUw/t2IxBQg+A6kDk7AdeS2ewIkTPZBHDZUH6Y4Dp0OncEnLHMG5IT/iQR8j4gmuGDvCWcBgPd8
XSrkItRMCL8rTF5VybbffBhX8mX5TYdj51kA95n1fN71FOans82tEJW4VOdtbCOJA45sGPBW59/o
vhcq7qD9kk0NuVSjKN4OEJeIsTuGFsLbL4vkFReoFCSa9442k/+0AnhaouwnzkQjZfHNW7BPXV9I
0GFsST3ogOS6cYdBL7bPIHwz8edbSdH69qmuWW2lgB22Ry5gXedZx2bbCsbX+Ua/snMbMWosSv3J
DWFAdWRgUqXcwMQHsZyrtq0zVTjM8QqA6bdCwGVyoSio65i6rIBSy58alMLWH6a/t7CdcjglXAcV
fFw3Ux81vRgfoMHDijQateunBSrxPBX+ipOt+8x9gJveYN6RF4o6GOQuRPzH0NtyoYjkIDDKjRij
FxBtPOf1NxZBX0JJAaA/sh2fFRl1xo/k2HSZULz9zTzUWSJjy5MFOuJVZqPhr+lz19YfywDBhigi
qnxpPG8MvTcf5eBXYw/hKKjwc9HEROM/4F3bPIoOWvg06Pnc/rlDJggJYKxYg/m0xVxsV7HvaWt4
16oU4fGwf892xKefT7XNTTMQPZgMlcIWf+tgSLCbo1clWPBVeL+Am1y+w/xGXx8Wt6PfO+oQGeZH
MIBH/5AZabxdpS3HOexYCIP9dTzUaQfwgOPhVzoi5R5hGWBCxhXAXQOQsxbWRsnMgDWziKpiQ7hs
+Bi4jFhBdwjgHvDf5FElj8I9dofIAkEZ3k3YIQKb+sqfSb9xiY5NYXIuUVogWwdFk5fH0ZOwc8Z0
gVQIKTOgeCSUh7sVkAG6WacWgTUOF1LK11oE+TfKMXSExsCIjWKuRND1GNPCby3qxv8jAazFUBFQ
g5/j6kYoYAX6j9Cl+hTd9uPsP6MM98vFNGId2uidgcbLUkwEw/6tD0MXqLSBNFgCGQyHKCG+EUrn
cP3mfst0kaX3Hn+5w7sfv8X3brdVXwe0a+4l2WW+fVDjom/Fujy869TkayhvjPIWphkR2ETT+HK8
t84ZjEZOlAAhEci5oexLih0DOXiOfVuctmjVaGN6cHseiIkK/6raqg/FejT44fSaxrvC7jFvirhE
sSK+jZMBQlh8i2G5IWHhkr9Q6xWf1fZi2ZgYstjVkg5ESLRxA6hGJyAzLfjm9fXCZvlTnKCLfK0m
f7QJxF4vt/bPOOIFCsPuLJgjMqFBuz9SKmHbcpUsf5KAcmEjHQYYFrdC/ta7mBA2AK3zH40D5Wus
s2KCZJ4jaywcVij8S2+mfXYQ39d0P/NxbReURAwmvABpOI9bjd0O8p+VZRC/cHneP+XShQxyNWCC
oeFcUtjha3Br68HoOepDxzCQv1la35/xZb4s12uV2+riyF403BksRFaPZ15KhbKF2PkkaeUM2Xz0
73JRHIn8KBQbyIiNctYJcNJ5bp39CTnQaeu+M7NGQGoYZ8jUIvNkZAZL9w6ThGvteyPwkU38Svic
SxBfkbjavBAP8z04OrsdWdpIpemJgOPT8rNlCISub92DvWoqPqAez1wGFj32XEAzbqE/BHRFNI3g
2dNZb+PjogDzatEh1uSBt0VB2mS0tHYtg79CRJsnxStq8OfKsBpClkrg5EIXi8Qu+IBab2xJJS0d
aka1pSLVlHqwe5zE60qAstgk7fI7rJDr/MiPhu3E3FSSQ2tZEdZ0sYiIHMTBpGDCkH5XvHzkTwzA
k1CPjV1LKnwXBxILehSvDIn582lRp+rvYLdJHaDuD2ZJDU4Ei5BYQTeW/fDHeuued3LB/ABoz7FX
uMgrxuFmDLlKpTjhHJU13zX+N0jUmmoqS88HP8MdBlLjBZt2v+5wwMnxSxVJWi3licFGkcu6Bmp9
ommTkxF0r/HYb49IogqRJrIPbpq+HwTE9l9MSZtt4C8OqI11F9SewHIrmqB8FjrRGwHs1X6PTjzW
jr1V0c9Wv02mUvc2bqPNjtrvAOtZRyPXi6hMOmni8qwUlEDEkE+Otn1HbyC0dJll7mSf7weszGEd
MnMYPKU2UTq9cM8ts3Jj0ZxU+21Oa8GavSwsHmLKvs8yIOnRYL+In9fsn685+Kv3FpHogWRk7yYZ
BqB4JYVIQPGzIFndz3keyjP3F2GumVzcpxievMLqSZH6EivhUmkl9xIg4Rv9pXU11TteP1fDdaIO
cDkfsbULqhTydifN7KHNUUhCYs6B6ZoRmva4Mc3TzznN/QsZc5I3yqRGSLaXiCnRQjx+V0WmVjLS
3ORPwZ0O0qPZKZ0aJz5SMBOU+b5F/t1gAPAGCytqds8C7pWQOTH3BHxqKgn+kqCgzqnWimF5NAHs
vLkFTXNg/8VRM19ILFtTwsQYNJ/JO8XWJXFs/5o5tdMQnI7kxn09Ncfme7f9sJHEjwP+Ku1zSxub
BbiKbsav4HhmM+tl1/u6m9pdMuoU0gN44R9JmpFDn+Dhd4mjKO/97nywP6LlOXuJT4YmJf8TMYl/
mgkpeVHS3/52EpWjpU6OeVP9iJXSzRIpCfdJRIzU40BwPUvcdj55JvbQNevLfKH4LneYCPWLRmwl
457+J3RqeVZI04CPOUpW1mOm1YwKbqdnKexrwnIDvYoBk+On5e4DWmxoqpxpZnTganI0Y2RD0liQ
Wq10jpJuVCyvK6suTu0fpW4GKSMYUirklvFTjYW0xbYjiKD91aJt7oGJllDGWWVNKYun9/sG7DzO
5jv1ZnXHfXbagEadeEPXa4jRatja2h7Eq0jVYu8qhrr8e6I6+LvULpe/wlmJYYjlu94Ns2BaN87V
ndfyCVsWUfllLlLSITDNV9QlLxJ/2EM+i80l/4n2q9gaT04ALdllRf45OtREmY+awGHTz0LZvKzK
LcRudvLOHKJD81zKVIbTi5m/olcYY2Kj+pS9SNBOmpiSq3n8qkJuMJs9ADurkdVRUrp3DUqHXK60
N8vvdaGoG7FSP+sGfi8qitOCkBw5AKOI6NUmFgzqWHg7MLYjg9FVTOJL+T8axE5IYsZtoYcNjTbf
uLrPvKqX6ggbcqfnjqRClQRUwPcMJJfXE0vkfS9UG0MvlO+tC6PQFGeXTqHjROvQCDN5CtMgf3Gp
NwecrMhaApr1oB6vuLitBoKArg4A9Siom0ymTFevzjkVRUmU++CP5lYZSYo5guDys4N9IqLKeD+e
rJamll3tEu75vOTfMopuQh0iyK2jCZEoaMyK3yStq17jUwCThBfwIEYdQyf6c7YZYvbqGCweYi3Y
flrET68TQEn6cDi6sr+ThuSjESzNAVKAUBTC/4S8W+TYFUgHZPJWK3+slwK8eHiHc1ReMaNTU28G
6WU0S2lAnW4TW4R2SRnDvXInoTO0CMWL94Jg6UW5Oqgqj24HKzE2UVW5PsGnYV1nL3BrnuXfDVQN
R4GPkDxXwoeySNxz4f/lejP1u08N6BX7t+uVC9CLqDuM2cvznkDwvxUEOyBHM7KA7cPgq1+aRSS0
hRcL2m6RaGRBz8Fzh/ZkzB6W7gepsTx5GBkuCGh4/vtrQK8CIvAWygWgU9KspMHEXlvAOix2Yk3V
8tE3Ul7DwRf7Bc0xBY2E4Gh/vj3GRMeZB+pdojadQavE0YnU41ZpCzOWTK21MdUXpakvi9j1Ny7g
2GqEUwNdhJ5LS82DhSFaIR63UPBZe52nK8pKc5uB++kcNBqgoayIceZyg+omDur42VN00GwuN0sZ
ARfTRAe6fXbd/1JRcChV8hDTOL0RIu1VSu2S4NlaPDYBZYxs+dGJ9XgVu8sP/APdJ8drOuvq2r9r
Swf+g2xx/hj120mWvYR3WsHpnIRaL0xWeKaRDvJA3Ge5YrHxhjxkc7rq7Xjo3FkuqnWcIsfb6o/e
CwECMcXkKKm3vffY8uI4eX8Xw85HUQR+yU4eRsFr/LSCdtHBfW0nP6lTh24w5QX7PJup/FmiGuYm
uJy3dHEuLrjHMbp3NM6a7awC8y/E2RMsfYMOqlQMxlln6/go8SwQXvazV3GMb6A2vpjwrBbFW3Ot
ftY+BVofMBDa47DCbHJb9LvQ5HRl0SRpJ8sBY00E6FTOJ+PRmlbkjGl7tqN196qoxM5fh3QzYd+v
/Sp7qRndt1NOh2jEi3eIRU6tQyq/O3DF1PQ092U6PDTTGWb9HsGLabvASqN9QKWS9ecg20sH3BdM
zpOm8OewRaPTkzpKvq1glGHsOH0Lr57W1q0Z8U6gJln2HtVb7TUWkFb/1qLSDJXQIwIw3FAfpaMS
koKcTsoT4rNyGbujX7DfQeaOU4fQwkNVvltujLHSS1tfnZJ7WxgxpX1C4++edvWhQyfgOXqvK+CJ
zygxLEoPZsS8dzhJckIzNiepSCkeoXU1Ga3Ju71bP0W/u7i6LjGntp40k2r7Rw9xvbxm7ZeYWLrx
PEJ9No6W0c/sRowupfjBbs+btIORFdYgrrJXkn8ScHdh+k5psmGTKwV129aiPTB+mK2cjLnk2mDt
/g+FjKqWycj+w24Qv3f3roDEGVCN8L18iaEQuuH+cQ3TNr8GWbzoyTUFDCRzzB9PYd5Zm876GEwq
ulEpx6h6GMjQDWryCIvtBNTba1lr7jOsCZ3dPWENaR9hn+y4JZDWsxh3/8XkEostk4s4X6ImUsHx
o7BNKYziHUHAJnBzarhZmeMo0GzCorsSVmUSOiFTvTq7eMWS/75HGdE4V2uVa29mG4HhDGWzPSi6
5JpYiFPKg0PqYx5nfbnmgV7btJ+8OoXS0xM5o3/YLnSPW0c1VeOHPSkScp+oQ2/TLvq8VfQp+GmY
IIKvqf0l9Qqni+ikExU1nQaISjhzqnWw/IS1ONPwDNCr0xc4gYSnVCrntTuN+PD/vv1pqt8TEEn9
5hTOEkNKqJ1u+2m8zoXbyD7r1JjDYfbysPIgnOyvmMhl/qmM5t08eu42PQrKEN/mfrzz3lNP769A
0batOPuIrLg920JcymsUI7QAAp5nbzT23pwbkiPhYclrqcp40jNO4CLBEgBe157O1v99eWYr/pL5
d/SfDrlJxTdJ4msIeuUdXY+t4s7ykxQlgvXiLFefPn3oGb/mAXsxV+FIyU35MgB8QIKoyw42Na2y
xyAUT96ZHRAgGw51DDbHYkhjCLvGnj6Sdt0uxUBgoP8u03vWO2mSEsLrR1S1ceZdHngStJ3Jg3cb
UhRKcRwAuK99s+a027WQWrfzKuC66r3esWchg7tzHhqaA53k4BRUOJXgbfvdhT9lk8DbXj2zW5ox
zHUMUlCT7m68aGkiLPBDsINDVzFNH/xSC5gyWIRGC1C3ra2uwlxRciYfZPkUBa1qgqUbzYSr314a
Mgx9LRTEpVun3u3PO3Bs6LO4CobgGAbMygOuIrBU7hqToGlK1Trrrg/45i4QW3vAeRsILRSSuffc
g0pwGbbE1UCHbFmV6TkYhX40prP95VKShLcgwXhC8IKMyIxzeHkKoFNRDLRTmNhgq/gQ1nltByYR
eLLLwgyE+QWxEqYjs0R47d0/BPinbLM1Bv9jFubHyK+AN7EnuFqnfO+OEXL5TZhlbJ8hF/BLdl0E
zmNIpX57O14L2QBuXwv2THoc4bhLiB0AQ9JFfEg43L2JY+FZmAksy+SYqp0+yFcqtsflOQFBHKXX
h9o4j0ymcRjxU9FbtJpYIdgkrcrfHZm5SMI/6OHfcEPK/lcc++sMaFAnyXJa1We5XdZZYYI48f3y
0OHIyIcPEbAgm6H6htoRqBQD6AfyNabXnFyKOUqj9IQ3I0AVHKshB8MVyhifIS8xN+k0uaRaS/9y
eZrFGC9O6x2KEtjlmG9av+acJFjSawFi5fon61f2Y81z0V7MGY22NGG5tXJfmYGT5zqw2joqG5SP
TPBUU4V9HqLm74vcZGWlGLqMqzR/rYGmSetjETFzojUBueO6Yaan048RFws3pI3JCR3LvWnAkK87
uVjZn6xKgdlhnGmNkf6hR/1wCLakdsdgZiXkvOrc78dqr872JvaflkPxZHMAMEMfOH11I7cm7hCq
4boD2gT2aRgOsKyyhstTF+8mmtNf/C157YrYTEGfoq864fSfAF4nrzwXtibmFSir52Y3PHBprJ4F
JI1SFoR+YiN64cVto7Bvm/tVNkCt36c3dkGeJsuDsNIj2+7oXi2ESjpVvXKWJqHXE5ydoPATGMw5
Ix3KpuChFYYPviO5Y947kqSlgmCz/0ujaYZibKdLl3qdgySZSlTBt4V/STUf82YGrNt55k/BDSs1
U3jNofWm25Eqs8y/hRSQs//M7lX1j+TSosf5K+zAQCoMHsvXME4WVSWXtoKRsJc0TGoxfWD3EfiC
8qIRXAzTeJhXK+8rJ0xy83481rLOFbFBREcfSYH5Z1HGunLtptUXWajtEGyUs4SDYDce1fa4iEE3
epePVZQPSbICUfMj6NhV9dKdIa9Yl1GiD2guP9LtmANbUdnLU+JGvLpI+Qpc/1QxpTuTJbnCT5lM
IAIAeg4M6Z6BOoSo9CpB56KYs0CeDfPKRvM0E7xS4zjm2e5/QbxV+Mr1VLg5w2fN0V7zFHhgddGy
PYj3Y56wd+dP+p+qyTSTfcTFfZlPdjWWddoVqaHFTN6uX0WcN0VOx6SA6XpnVcyqJ/S6aLCL5IhZ
bC3U0CNofTYMzYFWiosCFY8L68LD3cJEBpqM0t5ec2GQm60jReWwxlg3Mhl/+342qOQMqsU4COES
PNSx125GtqKqbdc+RVEcY6xvRe8sdjqGrJCDwO25CnDhMwZv1ELGNsVi7ORnwe1fAw9yFERr+vDf
PrbZqFQqxlLZ1pwIibixZqf/PCCnAHZKN/W5GPA68jTL/i4duuI/B/0+ZXSnNp7LHBBFm9QuRNii
Wg9GTasJYJ9iVF0ydo7zIKdRRCDCFAyZYUzN0R4RvsaYXZvg8pzU1l/mS2WNr869U6c1XIrCs//f
pG5fsrPvWOUeHVZCOSPYe5TLhAmukQzfHVp6OxKVGwHOudiiHzUg2VJqePmLqeU6eRGcAotPmHLL
KZ+H/KVhv8szgj31ibQa9ow4resdrWg45McqbYRgMDj4CjIX9bsGDCfPXXJbRYisa6tN13FBrQ1r
MjAAjRHzfISXNJUICmKnp8YV45LSIsF8xWdv0EvqGXNgcXt2TIErq5TW0Hlcr0yd5dQeR61Cnr+Y
KIt6a/u1grWzWqt7+kpq+7vlbcdts0jMwRwgPq6MyzbHQtc/QRST2f7oVPs2xFSK5Fq8+oplAS26
ZAkvGbYe3kjaivCBrCPsgjbRmHxS6Ky7UFqrkJRhXgtZSnotmV1opFfCbC67KbfRxYsFVypvVPjH
2aa8GQ2lh7sygTZHmbjb3t2awIghOcELrLckfqVedBf4FlpfTEEtk4OYqpY7MH96OvJ44l+rmgao
7At9Lv7rDCnbm2+ba1jX48ot8349jQ9KyJmjKPKqeTcyzBctI44nYJeQIRQXwe8WJ35cGGam80FW
YPX+k/RUuTpMVrrA1SUaqjB5kliJ/4zOO5eh1Cb8THtbtTEEserfxoTds9PewUNxnQh+3EqskkBE
5HQJZCQYoR3triI1geSsbm/gYRuRm0QyXJbi4KzcBVGorJMZmKRWn706sytxK8MLRYcsf0D6sYtA
tTzMsOW2j32yDkM5c+bVIx5Z6XOMr38lf4qPPfEYLOyquX+PyZLxG7pNUohBGdOKTUiRnpiMqTwW
G/GymObw/YVJFh4js94N1mBmAT++YifJ6eryQZVKCMjOa3JM5b6en9R2YLHNBSjQ7k4dXSOwtE7w
cXcMcvKpAvysebB1xLJA7QrI7qL4yRa6mNvqumq1i+xOAgAv4nax/HHbMyoXYcyngVFjEr3qXSzB
CP1vrrebcRUfDBUF/mo0uEMY8tCCr0W5JRGHTKfeDbpFi/U6AUe/gJej6TzQZPw+aUSHu/OOduYN
PdgWtAEws3S2dXzQpS8EMckenBDMpoQ6RmXzA/R1OVJEMAaAKaE+650lLzwSKmTzk/06fl/Oqg3y
JLwFdXJxGNywfsITKyW8TzzBwmGOPcS0btuIgxPBW2Wc9xHAoxmDw6uTTKIl8LCvam1wRDrp+e+t
eejaqLOjxq9Hya/TdkOIPgK+xYxVFXPifsv6eWM13rZ6OmgnB/loCaIogYghhiXpba1HOcaspq7m
LQHSKtM3Pamzr6PymYpgZMJteZEguxFncMDG46iy7Uh1C5z5ooDOcRFnJtpnotr3pFSZlakMTXWI
6wHKBB+HKYuKCbdQW7ssgodUDAkkomF0p0tZiY/Fk5C6ZSOXKNcJARHT13eIpNJHM+kewdjclxw7
3VnVkJvPThTKDh9rQ+smEb9yWhqmouCdS+GPCJkpm1jBeCOhscDwJvorLsE5XLYBxSzs34q3dF5H
nze5vW8188FWp7x6DTE2xSa8EYmDwLOImjJvZG8mKIMtQVewE4SboBvu1YCpSVj8mp3k59uAveui
5L6q7zPV77hiHI93VemV7+1HRd013ctXXGDl9mEM8/E4Ndqywcx8EN7JGiQ0kDlYg8tHk6N6M8uf
WYySkc7cueV4Vj0jDF8jGb89Q+o8FGTmrQIwa3QSFYeYUB5sl3mB7iWywu+Zcd7GemN0ZgJI4GUg
62EaQLNUM/SvDLlXwTO5z2Ms5dAts6BDKwUQ+Ty1IGQ9DZYDcDzUAC2ibf15IeITetdOrN/x8SMT
VlTk6G/g2WtBctilutoCX+5ia1ydP8jgjBmbsko+26/9tf8nS8YV23J4QBOoa2NQZIAIN50nB5Hq
Ia1Y0lJsi6Hf3LUavyME7ap6uMS6S16dkaZ6996IrjlHpaTOf7uQoMghyyEXp9VvihuCfgiN92G3
slhhEbi+6/F12PRTSI1qEmiNSfXA4Y3AS9N0arDdWJz7XgIRqOr2m8Lxac0GUO+l/KI7nGomNOYV
Zgdd4Gn0L1T//netotYAqFikr44owVDQ/S2mPpSW4wKFl3LLlREIxYDcPhJZUCAPbaXbti4hJsl+
VdyuuL6IrV752orFRwMTKKHJSfKPuLpquCgG0BvvwcOSkJGQuqFoFkt/+VoRh5SC6yBrp2x+zJul
T8rzoR4iKc1RFBLykCk/Ir/zq1LYBMhJvlnylg/KSDctJ9b+djIqXkPp6yCwkiSSlDgNjEPa4oM0
VbK1P2zJYw+qe4t6bSVwgclDoq+lKGE3j0OFhRtJYjPZLbwznSh65COgwWbszr8y8mVCBMEFqQoZ
iW458Gelt9Ft7A0CV7CY+jhKUvfmTfmYzn+tDjfy9a3suMqJmwRslelfE8z0jboVKCjNzLMJN/L8
WEcYjOvZA8ZDH1PR+kXOv1BmO2s//h9esu2oz8UXzhPoVhTET6XmjbRYgi5Ej3ZKcvufS/MSaSB0
xjANa+hoRi1ckB5sE59zezr1HWKjH+xn2rOJbYDgy4gT+hCY4k0z3xLG/+yfowBttuoWXon4Dpz6
t3JmY7sphRRCSND4jUtDtMq2vGDSu1dRMIEk2BUnaASl7ZlE2V/dxkLiQuIERUqWdS3sHYzUd7tp
u0b66WT+zSMY7pi3UnWMkTwoQa4jV7QPKRlejSII8jawNg4RZNDjOhtmNkfx97sZM1yiiR3uaVO1
RblTmqmX6Yi2DQ2ogom1dX3DyZDz7nKZ9mHL43RXAxCAqCEf1W/jQPir1DHmKsizeaA5fqY0nNFm
SdVVLB85h9kRF85d7P0MJDPL6jx+DJsojsSofIUUKWe4qoJHNlLOsEhAGqMBaCodpzx8oe/54KJU
q6676p86qJvl+tKmebDxYXGhX+e7PcihQ6toph2Qjnqo4OSFWyBkX0+TXwQ5sK2hBORnj1nmc6EY
aTPGrMXDEcPogY3Wg2DMdPwpqMzPV+PUF+QLRqzb1UCu4Z/2whUZ7gY0mjvfyDwj+GHGKClSY7ph
kJ1HZ5P+np+o5aIpAIghp9dS2mE/TEfXQ6/+aE2a2KdgR4G4ky+k/LNpxL7TGQd+pUmryrDBGN1L
F3MzIWgwdvEdSGX79Q95YwoOe6OQblnXXVgQU+YbaSYiqMfhlSDT5jXAcxnkYG3KS9UOccWsOXpt
HFrHBhA5U96NW8a49YiEiqY77gvO1xCXdos53ph2SazFPGI4GQH3mkTWVS37R09W98O1c6y7BwMC
iMOmrjraRjQGug9NoM2I1VQnXTFgpp1pd++U1PcXPsfXKGLgjLMbw38yS0GIogVilMyr/7iO5PBN
4UMU+oUQ/FlDYCpy2QsNpa9il1s7SGcB0FF5Bc/lQWs/TZN0QtZigDXCTw1HhIsr17tSsWvQ7Cqh
sJipM/r8tmbYkTkRHrTEkVyzfMhutGvacu/RMbFCuaZwFx7W0CMsiTX2BuHSY25WT9u3/DANp10Q
SFiOoGZmgjWy0ppiZUtcq7P1guqU1iAPnoQl1yy2FUXZt7ZJt+z2DPBaiIwPa3iJ7Cgk12DrXYwk
pWAGxpeUPvyx0nDKdSrQunJqZvfEHuFmn4xQfh8clv6UFa/b84W1IV4ugX8CA3O37Oka4vt1PrAS
sSnL8CwO/6YZVDOhff+VAiPik6qgPajtQOYUUAUuNXGVdumYBiSlFgG7J9W+JUxfRu+0OhRcM3Q5
qgLVw8uo8NgvkqEIFXUgum54EIqBRWTxTz4PAPCE3cu7mnUE6gOO9s/xfZd/EfRGHhjdpTUqHC0/
EC2QbZqFLtAshsM/exyShXs58p3ydl7rkXYoLZ2THHMX5+xzFknJ7Jd5jLaxVOWfQ/e+OlYLdWo0
qqD2RXL3+KUuQFv2bHM3rmbRRUEHonJK8mBPgCSPI5r3c/4HxJfqZItlijz2slMLoCrVg5NI3Efi
cD3uo8XoKfmGwcD97swHD/tT+FlzC24+hLVryHtN2rKH3GCfmOtB5cLfrW1tJJOO3raaaoqy0R0z
lTKsAYOTLuBRjyvjkID/sNKUXhqYT3loYhe+XFGppIbMiR1Q+kRUj07fTFnfszrjESgz19L4BMUI
KLFqBDRHow9wsyASP+vdU5no7h8n2S/Y+QbkTXKMqgzoxwxa3TcTPxR8IgRE+C82lC262792vpgb
9LuzIMUTACJtU68dNakq/q559ZzaSXj1xRIseJRd/4+kFjge+dEk8T9D9p+AmVCPC2mrT1L/N1xM
/Yi1zI2eCQNjsnpb5ugLpKqgJs2f/vUWlvnccKjmGYnfL9z60f25rWVblB4W0zEfxF+ls/AMxuQx
LrwVcbBWIyxFki6tc2Xt5jFXsCtR+68GImwzjnLkkeLX0cezn5uTav4c5pKf7oh+7rbqzO0cW1Fy
Z3inlw1FkpxXE+BNe/7zx7GmVHmVV+TILIgOnlKcz9LsioXr4SF450LQRqrCRSeAfcU61PuG35qF
6ZuHm+WUJd/Bk23yJdjpUyQBkLWrxAAgqQTBnNWayYQgraytdoKj7KqDyZBkiV26dP4o/34cjhQa
+2+vQaedg9LVviyD3J33RquMXlzXzqYvPK3WzajNWbCAaGxDo6cZj1RnDI/yrEsp6rK3lGOuL78k
ZsRIGYWRBgWThzS5C2QjwKq0Mk8sAXhnGqW1hlZgFauDJ7s2nICnbqW/qbHBI3AgljGhIBn1vO/7
xRQ0uPmrAMLS7BpmhBgil8Zg0dvYhOtRaPxkRcpl7z6CsyG3jIrxtWTULY+cKp5Z1BWbEnYPlVXF
Z6ge2Ji+RxVuMl8dLUP42rpKXFwlQi2U+5vhG41Ka/vBcAL4x8LioWFSHo4nIdw85VkTGxI/P1gt
G/yHOnM4u/Z8nXDw7Pr9aJrLsC/N14neYbe6UD7O0Q7o1w+CdXDD5wGzgg0ayZ1+1+Lrtv/2P+mG
Qc6pt91PGI1/klHHK4M+CuZoVerSNCDGQhVExAb4fOVxagtpjdP57x0o/IH2oX0Nz4dLVrsB9GWf
8W+dhDEA86FUs5pBnQUCKN2JMTYzreELdBbgFe1ZNTuTz540G7EBiqNQEB0rESN/MqbDjuruQrz2
Cpan4GnihZc8bwnbZFqdlmNQhagg+KQFRG9CqOvcf9q7OQLKQOF4h8J/h0s5ppnz3xMOoE+tIAXX
TE05RIs/imTEol5wxD1GJm4MJK1SjvTFBZjSM0iNmT4/wZ2GQtwdcT9Bqex53pT9JbOmDux1nPvJ
Nqu5zE4PtnmEmjE613w3kqjYRWIRVsXjReAPyratLtmNcvYakNMxkO6D47y2wgS6yrSCcOUXZbgp
uA6p5vpv+BXDK2+mhnSyt3tDcDrCcYLGsPi4Bn9ezy8Pd5tE2t+FuDaQWDa48dkfz3ldFcDV51rT
vLxbTify3lTSmDaHe8eZjKOsa1tQSkkhchjSrG0uWSbp1eTC04tGCtgI6mSQ16rjdlahz3i2DXFQ
QM4bd20Th13kGZ5dJEMp3V39j355Un4rC5afilKjez5gon39MBFv6FXgDwjbN1qT+UasRZKYU1oG
x369wveo/u8v/ENO1jmSFr3IC4ZheV9m2q4YZzSZBFDe+RqVowdxGxojkMgmAM6kCOcZqv7hnSMz
WIun3/F+afYyrlnIoYmc7ZgDxaAoTwmLlBiz2pppbknyaVKK3o6+Hv4OkJ5kjhXbJ5eWz+iEo3QK
SKvHL64SrweyNxrddJZ/1G8N14Y0RNPNWXXIWJcfnBylfCBM6MC0mJZwxOTTRBzgEcg4GgehL/7o
v8L4B6xdeBpHlTOA79PCvGzljcgU5rT7+e+M38yiuXwiV6TKH0ScjwdwuuHvObLan5m5hMGp98EZ
Xvi20/DlRCyZs7jO+yaujxcCH0899OBIodL1Kq1ZYoekYQuNPT3wEBV7Ih7vykCcopD+/rRLd4Vb
+PDhv4PtX0NyUdjTyZVNqECkO+2iKTvibBkU6mnPN/alqY/8yJrV9og2O2F28NfXqGEqBwa4STnc
8yp+Vv1qYmUx9QL4SQOr7WMCqwXWR5FCZnbDa4cM1F1UyDtiqepNcuWmToyM85FNzxSHoDNd2wPD
TXCcpUad2m5LyXTntv6bNPr/GeIrttvnIiFfSLSOgsClRdxmIqHkiIxwjal5oUI50tZD6IR5HuvY
kP7JrVmmPgLXuNH8X0ygtfoEBhhtsxOzTqArbQhs2i4M+knRu5nZLkpPTHyTWpyzuU7vUkYS1avU
lPlkqwBVH1J7tVT8sdh/TF5kw8+Uxxe5KlFdcy0ocPE1QjwCHB3QQZVuxBL31J/L6VRo7tsktSqr
ezOwidlSuk0Iy0dvCNRMQ6QPT5XOhDuX4Nt+kuJA6Y1H2ZdCijY9TciVw2H37HORSvluFwma/bFM
0duATCi+4BDehUFoE43ocb6y/MFBvgATLPRATsrUkgDxZ9pji/teJZPr6ACRnu1WncDNVY9DGSWx
gAcWtnDYgomMRfqcrhgSWw7DhpZz0E7sG1B4tExggEfeXFIso/c9j28055kCHbrJsBrHju9QbWdi
8zUfgCEly32LOHkNVo6gZ9TrT5scDO8ppNO9g1YKHd8O7kP55dxsB+Jax3bQiRB0I866sS58sslw
pBx8V49OHWpzqFKZBkjEB7JYfQaPOKbD58x/t+wOnQS6dphxNj7b8voFEstUTIaJ8gyHO3CwO+Q5
WuORWdTcwAoHX9I2cwgV3Y4Cgzkz0Ys8obq+Zs9WleHtPpqec8XJ7/pYweZUdGHgJ1W5lSPs3J36
ONGMottGzJEGlWTZPfRAEkLyMMdXn0r/7BVc2cA7ExTv+g4yT9+tvAzBaoiUqxD2suY3bU+0BZ2L
j2t1CMqe/qmIlnpGxVmb/ge+dUFu7arAEEUMDS3pnddlmQPgjwg30e3L6v1H3tkRiTugohTdgLhe
TwUrOLaxN/vcU8SvXFVqXAHAfMLAa5oHAOSbIQjLm7TAjtX/0AIp8KP0CM26DM2EUnGeNtCMeZSG
ci9EfrUmcQxEt+gju/DzOSqWRva0Srq1nONPWI7KO14VqeE1wCpZ7z6sS5zeMLSBJv6x0lEpV+t/
RTpzE2saNr530xZBvefxPxwXLd/+VV+EVnB9SDrROePw/4QStkvXIChNcGhhBMBfNaa7OXcGQyuA
u1Q++0mpzYDD3gU65KkUlv3cy/on8UvnFD1ykbVnZRQrjPmzzgagksjj8R48OV4D65d6aG+5MYcX
UH6UDgyfeB13QIfjV4Bxnjfqw3880LT3cMVInyR2P2LwYKRM3Bg+r5o8oyGb9Isf//HvhD9pa8n8
yOZQyx5qlK83p7ogVCN6a+HZYf8agPMGiN5TiiiczG9Ywtls/CS5WACXIONYIx3DAp08Q0s32ZiN
hLXOy0E7R13l6MCTIe9UFhrI6IeSjocazY++jqplksEaJ0auOVDY2wInHORZwLgabfygMo1ia+3r
HFmFwlXwfTf6yiNRUZZ8bqEKRa7bb+80rmSWwlyHalTb6gYoR7Mg+fOOEqOj4+9nA680/0w3KxtT
ogObm9L289zSH/7J7wD8u68I8Ea7BOQK7kRV0wLSZWj7BJ7ashJ8UN9AjwrR7vMn3B9C+HIq+TlK
Vo6Fo0Ixd/5MLsSPWJ3j/9fpntOASkl2kPk2Rvz/HQ8VpPygi7QtPXY+O5B3WZHwbo6dJHbHvrNr
yU1ORfwDtkpT2O2iPH0EVXa0vtxtua0WbexJuPsvxzqzYXmt0fYLOU0z4MqFB9+Ahg5JZlBXLlM2
KomiD3P4s6dmgzAjybGqBJARkbNMgE69sQitD+bd5Ocu8r/YWg/HteDcQFYKidGeV215Yleh4NmX
jVHOeHd8zCQ0X481yWvrBrgVc8ZN1A7mvN1xbTgOfomrWI0JbhuLBIS52o0owE3RVV7oGrsEToRj
PBty5WRcLFMeiSNOZYwOa0GElC1kupG5Jqb+Z0O/uErOAY68Yhji8eJVU58UPouzLVmwlzi214cx
0gBe1dkNcgHIOZ13WJi1Q1hDqJEJ0xae+VlJDaCCv5OC0o37qtoTKOl0CWuPHWtqJZJazj6rOwpn
CxXy/sdXQSQ4TkBu3MlObdCM1XMnhRh2Cf/p+yHFUPutWbp8+vJuM9z4RFlpMtNMl0F59SdO73yd
Wcxpr1dkjlyeTnFydzsC+YX5KtjDziMeLZozAlcEgz0d1Lq6vR/6YXVQXzyUPEKeHOHLTlkQSvkT
s7nx8HD3kx4wURI9Oq3YUGLj3uVu2n0/kjoO9JhhZLIvTmdABe2KrYiTMcx0cSg6cNgsjD/+DYIo
MvFXpTCHDZslIFiLFy/nzKOFEzI/nHHqYNBOLBHOzfhX4YfxNNpsBOXasrN9+kzWc+u8pr1mEvAt
iukNpmFce1PR0sAJZIv6jB6Ntap6wH69W1suBf1x0BrpwB9VA2PM31QmXDD0X7UorxhpGRnv8GUH
6pMofAm4D80EqW53EGfmueXwWxhT+xgs8x7HYHT+PkaZQ+yCrU959NgvFBpYrdOrFSRvrkJQItO2
UdnErvNdwYGEAFR+ankHXMFAI1l7zw1P//IYvDSdp7Os4cecf9C91Lfj1jwLdspxlj5/lTYSXMBq
iw1ygH2/Rjvi0KK9rEHaIBkiaC8lOarzh3t58gjn9bpX2W1ulpuEKHgGQ7jUpCv2CWzm22FmP58s
FqKyusaHGqbi32Vqx3/gYJBNTKb4EHQPM9splEDxDJ2Sma0pUCNrhA5+tlZNXzHtDg4R0gl4WutL
f8WOi7g+BozLw0g1lVFkyLz02EhUTGTl/0+iYvt36uysVWmjWeltUbhQoWisHfN4OyLxZV8gNzbK
bWnjMSGp+wpJ8QPeNtJSE+JkZydpsH+1aXRJRDGiymGTOoAA+0ygdjTe9K+P67+zMyN7rKoJ324z
7Br/5NhJ/pL/Kc3L0J0sQg6zehsoT89VU0Wy/q2HfIh+RXB4ezdZOD+IbeVEaYj4IOAEsWBh/0HF
2bI4D4hluHfo58AkgYgR3W3423Uu+qo/QUWPyP8/BRzKJ/iFSP/NKzU2eBCGMfPIgXLc+9UUaA4B
FExThb0eTzqXaMXJLb77A/2oZ/6UWsiGjOiQBiJr9OCnhP5932c2QvQ2r/annpKTpO0GqkarUB9b
RZmMjCq0GPtpUU8FqCVBe3xwsC1vpMl3wp8b2rw46xjmqL/BTQtbuwk+SRNObNHWem1oGhVcvS1D
NfD567DQWqS5jSTRYDIWVaOASGDav3szOt/QJcKytPtIGz+bIWniLHZAEb9Th4sqQ6AtR3qB6x9M
IZ0HvdoIE5l7caRGki55EHXo3wAAuwj5ubHAginAXwAzoZOtzGHR1egNLROyO84xylK37NzLxvtP
RVL0PXCN3sOZcMZg6VYvVQVKgvUUoSuqZIlfOiWrd9eamzWTPOh1LEN+VLswNTdvqxWF1VhkXdSY
lAky3oTXXdCV8fTONorqFvCusr7Kr92tVJa1/vyjJJ9Ckv7Zfjb8IvgG68d/rcPr82HdKnX3dhKM
bXeApykDqEaAQp7FoY8yjqoDWkjokvaTqb0OSRRK5arfOEpTcVrkd3Fc7Yz2KJt7ggRcfAdnWGES
wvInyAyeG97DN8o2y7F59vZTiRdCgwvccERXXvQT/Vo0CtVhnUi3GDm7FQCeG4Nkm3ExElJUDn70
8hnEmRuwOw/Mhmy9MQQ9mHi5HIiZHGYSwiWykN+D54r7YL1cKELmeolWQTqkHaZglQjnZ1tPbIap
nZQlki23ToDi0jHuMT8eXaYR0eItajDiMre/9fc3oubTFIxHqSv39EZUZ4Lgv+tIHxgTlI0xG5gm
emm8rf97vK723ESap//uwCJfGtdvyQW1Lxd8DJtSAiPeQP1SPYXLEoRP3INcIIy7AdX+eZMIlb1d
mgRTSOHXMEMbhbcdqgJlmjiiZNjn8ojSa4WkcDAsbbZNw0HfFZ+VUPTwpvvgUb1Wb/BPXvL20gKt
3MZzU2QZsb90ZAjumQRP/N18So8tWKHx6wpRAhHDqEoxuYvJUfNW+46jJucDgc12+xRbSUpsCiGt
FSK23i0V7McPRuQf/AONhPJo5/Ncod2VNuPNA7QtebzAtp2FP1Mv76NZOpGNcZb2XuO1PKy5zynN
HctsQnoHGMNlip2B4FOlqMErhyd5xv6zkjG5A1krAO+u8qhpz46cdi1crJw9rMqw0nLWnWn0l2F9
8M0++t1GZnVcbv7y/eDlaPlJcOCaOhkmp6Cuxx2I69SQh5awXKD8ilStDlnHxUSxUACbgkZxPuFY
Fbn6jUfDnHlh+51XKENgYl00LJspuIlL2mKpydVxiKFz8H7rLAubZ9YNRf4siAKQ/DDq/htNoanB
jPJ923B6a8smN8ag9ri0UIqzbgm7sEwzGN1WzuXgjQWVsQyV+TciDleLc6wvl8tTcaB71+By//g6
mgHLO3cI137m8mDUlpG6pSM98QnYFp/a8Ae7VQbExkJWFq3iJ3Rpt3y/ry8pg/PnkqOrBk5Yi04R
XWKTzq7Un6ctCQbMvLfMRcQ1T9XQk9dwlEoP/8Yav/HasOVqGxZU9GTpnT5G+CU059KdUfYYP/xJ
ZMImf4ts6UJLpW4Smi4RnRCzoPmpTHKDMlI5p00Q5rUflknDsTb7jBPbLk4xGyhEHGsEqdcnn4be
fdAAycxBpybWzLxkJW6i3TTfpHGKhWqiJewsGEEbSyuL0W2m40qzROrBeQaGSnUcQKkgHQcgmuhs
Sf/9T7k5OMonhiF5NhF640LISI8AK6BnZ/r1eyssa0rdI4jmv5aAhiGRlQhaxEbm5jB/vi+5Qg7r
+GI62z22jwzEkW4wgqfvo23+LCgtzNJyg/zLxsXl9ywCyxDXBFIvl2mtIcuIFwUnRmQObDEmtN08
/yJqVP4AxC7q+v4snotOWHzWDKJVx9cy+0KUAC2EoyGlvRueWf4exr4Ksqp/736blz/CXIYFGwx9
sgelGz5A8/6ElGsX0mRtjk7VXVdUAHMGaZt3jfRS9K4pxXHvX1TVYBIf6v3hnp+CPZeBC8umc39x
dG23RR+jXYujka96Z70seoZOTVUANYFxZ8ng38fIQ/idK9TBlLgAW70/zzgHRSyoCBi70y0BVz4j
dmTzryKnTlD71E0YOgUYl+1faKrFNzXdUCyPiFpbH570ax0Aq8KP9MAVgMc/9fZHQWaHudJ4Z1VR
h2DzFm8q++twyj9X6UkjFiOW0V/pUnpzuJL9dzJ6Mmmjen8Lzjsmulv6ma732cwon/kRuoEbfK5r
Bza836eIDCPsgN9U3PkFTEWqgsB8k8c8qyxcnojlIGcprZWm9xiB5NlNCC571HGBl+jAjTd7L0dw
8lTmCIC1zsBVA7vaACIHgKw1S7n2GNnnW5jGgpNEvquvf+bv2weI2OJETJcryReM4IkjReptUleW
Ndw2B/4xbq5zwsS0WSo8s4Y/rG6OM6rp1pV4vtsNrkbvEFev+CJabed2teeyJ22YyY6dycULeoFs
mThfMC1xJjYb4IFdZFhlURSCmknQdQkZCBo5w8ACEAyqBsCx4L3rba289QXwBwup3bNPMfqhQTZ5
SCsJVaoZHeBI3dUUDaGcFBhTLiB1WX61ojw6tAjhkGeDc4JVbd566dgamyDy3YMlwh1tWnhT6vBq
NeUFK1c7WF1XoI10zmNCl8M09uQUKPnQDqkRpSlToOrH9AiSnHUz1PwctTRyb1GRZhRYHJPd4sii
tKUBeaMBiabiNxWJsEPHcOWo3Kq3o80Zvy5sNwTLWfWPHEZcAffdn29EYWyuiU00i2apRHKIofi8
4gH1tx9ZzacW/D/DRlhXe0+QlnzoTRqMYB9OSF8jU7nSM1r5u3OWcxlLAeTCOntBd6HnTg9MS9wm
+AyuyYaHR0Y3Xw0NcvB2Ci1Khbxx1bOmLGsbc01SPrNbYEohfyeajZJbeuljldTA/w2MTTp8hyi5
CNbxUi5YuZutbbz568qyIfupJVf51vuVVVnQk1QJn/6a7FnbIaJjS+VZ+pIQ2AUfC8PKTO+mmhVd
sHDAo8+hISyYX9LK5O5E2173kOgRvDAM6H51uwfsP8N/5j/yFXawSCfvV4/HhQN30SHncXBhjELu
5lcPbQcrNmQkZ9bDriN8gf4DKHIJIacNdieD5ZLbqNJqEdExlYzx7WpOtMgHIBzJi9sR6jynysYH
iugJQrmneSxGF/ZKBzfiqyLp4FwQ3Rof40n8/ktOmrLgJX5ALcHzlKYGPGweqLJ0e69nlSPNUom1
eJg+KpsebowKsWq41wUp0i2bWajUCNewoCrcf3UIy3iLZzVE1gCXV4pCyo5McDY3Acu6kCGeQRoo
HXGkBxdsUWrJ3ZoglSpwO2iCnTef10AtYOMO5e3AwFnD4R22EIPTA6T+QsP/Qael2Y7H4sHlbKvj
okjoAdAuUozRiUObkz2mO8f/NwEZj6hUbN2PzHeHauqCOQw6P8/+ZkktKf9jF2fqD2yTmOKb3jZh
j1YfXkibHsAg9/i00xPc13W7lpTKCTQ4O/7xW7om92Fvl+OeT35Y//9bp8gT+UblKZ+169HQPKeB
ZMxtujh/yRnLyy7pY0w3xH0ICvN2SUUAE2RVSaoqBqEP5UFslByQ5EJQbql5weVOJTSd8/Mr6jTM
hs153jO8Z7wxy32Iewwo9KxmI25FYwZTrqeIC3Gvw0Ia6vHl3NILmOr4JKmkXAguK/GMr8H419p/
i+duk9LnNJVIL5GKTwe05D7UVZTS8EaI9p3OKwCpYKfopInLGPA8nbPf+YqQbxFCs/bPqWzAk10h
sAfAtbmvcwzjFSayH0BNzy/r1a5mD8SP2btg3BNpEjia7P+SiQRzyV7gEQNMUGzbaMSMfQrWdhbq
3+gdDL8jkpL6pFBibcLQDbPEDrvrmlkEKCymKen5XXiKiO8g1ZmDjE+2IfsRntJKvuu90clPm8ZB
xiDqz3cDLwNg6x+heItAHy1zbVplW1khp1pFx6HiJMLd0P3CEHUebOZblrs58jzYxC5Aya/o9fg2
12bSLpsk/GxVMa4lzW8aB+zg6+RlWvGHOx49g5Wgfd7kDcRnmEO90x405ge4iJSP4OKYth9ZQ7DC
uLWTwOkWpu50BIIQr2Q9VmRTupY2BJKahPmX1zMaKyfbyMWd7BwpAzSQRtxsKh7g48qpeWfT6EfZ
fVidAW1fsL5feLLbusXRfqEA+sJ27jC1oaXwfGBlXxkCn37lySoaxq65uzoOJkeMbHdzIVwOShtJ
HfMJGjnV58kk7+NwBqCGX2EMkkzfgSjguA7L766zCcwxzr4I8ntAnoXYA1PnSeFAxaIbCzZEFP3Q
HTvPjjZHCqKByOT+KCv24J6b0RNntYlbxssEcOOOjQFka47ULSlyXYr3kJVvvsROopPquXiBJcyj
dLGFA3FkQx02MAZ+z/bv3KxnGQE2jwVwVXGqn36hntx3g/4JmEmf4eml9AV9Z6P+FjnXO5Ko0HDa
Wo3DECGz0wYZkVo5voOV6mLfZDbdoo2Jx5kYvUSsIq+Kgdmb6oSlPM4ALeMu74OGFIRbebVwHKhr
44+Rsu8bKBCkTeCrdoItVjsdo6J7P/a4sF5S+fM2bEYq+p3pVAEpPjz7oLtL+ZAjdoptA2KtskQb
4yOMUfJB6sFEgVbHBS6tD0dqc5FcJ1utFqbwS0uQLCM0aarh0vvr46eUguhTMAuVgXfR3CQ+TvJL
tL/Tau3HscXWIXDoEqdCfquTlYOp8fe5eTvSCarSW894qWcsx4JvgZsEYyFQ7WBNGkT7vt291EiN
kwNTx7z/ZS8lABM7OQTALzIWajBP/oKKhufa3avTehR0vk405Wh0O+KROEM1WPBIxGT2BCYCtn34
KdU2keo2Ce8EBKVs4QU2pSY5GtjfzFLOCOQKRgXZqXRQGyel9Hq6Xi3Lr51ndGNWz7U6FV6zjOH6
aKsqqqggMjTMiXkbpNWDmiCX3kiVdQPmJFd9E9+kCYb4BG6jlHbdwQWKTiREhJU9ivpxdYhtPY+n
SDCQfQDJzEgb5h5dMKxRBXc8R5HiTFmTKO7EjzukPL7SLhFge2B25Kg0N0c2Gd7MlrQT1BDRHmo4
EQ8OZAJ8b6WWT3nez24WlDjDBbxhS0K8D13QFh+kK2/sw+saxJ3G9muJP9rgSOWMe8J6E6xDnYRP
VJ4HF5vTEqpdwq12LzTV7LfVJZX+NKUb7hwRSDgBBsJrvojTw2ME2z0Gir3x8MFyGzLmErTxaujk
pJmiN0OQm50kpOH+8ZfvmQ4as/0joy4I7yyekDGcF3O3VSQyvjOFMRGNG8wcm/pk5orxxF917EZq
uwhFZwbRnhGY55gzz17DGVR/6l3DWVGE77f6oc+U2CbuZ4y02SWPG07fPR4p2hNeTWvvCym9ciuB
AXyH1taAMiwWGaPlZ299bO6BlkwShfXHjb2T8MRso0k1rlx7WAA0Ml/Zb9fwDh03dzjXcyykh1z/
KJ66+k3x63ReDOmgKBENdYwj1YnlxozHaaijgMqjI8ZKCLHgkv0NsBmFjIN2j9cGp1gk59Bt4dsS
GLEtHTDcTPQSWr4HSf0Zns4KXhL2OEgG23XQUD0tganUEQkyEB6zT8reoIT2GHcBV8bsgJj2ggj5
Y/R4otKNrvAwoIYcewCPlnjnaQ/WObfm4BusMxHXLcF0ZMV8p2AMxpwMA8b/2+7/dJiMg0co2SCi
EDeFVmeIM+Tf8L3iTE8wR/KAsXnad6DewmKOLWt5Fj3ws3agt7lwCD6EZsBUIm80Wb5tWIKzZu/S
Jlnj0gsi2Tmc7juPrmucFgq7FVVEniews7JZcluY8jHji56C89KoGAWPA5xXy4j/iQr0ZW+80LT5
HBghgz2fTKQFk0u4q8aXzSH0xs6jEy4vEVQmkCK+8+Guq9db04oUshnZ79PpjLsLf9AYSh6aezpr
YyCZoKJER9m1M/VZ1oz4AaTsjb2YUVt9vfwMsH8x2WafK4f0Q49/SaC+IDX4sj87F6H4XOgbupZx
cG5o5W/ui/+D0KOYk0PTxUpH1uBTsFDI+3znqDK0ULarcCIgdyOZpW1OAFNDWxWTV164h/kSb29l
X+9bGRegMXqXAdSYuwmce4F8NOxYkvLXayEud8X2h2Ze3+CPoiguY+BOFSvwV6sMqLBiPm7R6yhc
GyQ8KNmqtPr6+EjsJ6GEfQTwH7JuXYqPAEnub2xFP+QTrly9Hs75UYT8gW+DsWafd+3Usj+CTXK0
v7Vl2WaobWeA5fuGRnQQbzYRVSBYa1AtO5gsIaqDQl/OhxOPfHP61f0sN9S8HjLuhqko6KImSoTZ
yvtaYmStOMVODUnVuzw0/pICIhpkEdDvcZ86p1QwQSwU5t2Vv/nDfueRXfYLIV3rbPDg9bNJ7gBO
uPUY6ugDVdG1TBAJOCb/+oWApm4t5KLmuYUPYTwMwvIvfcuPUd0pMGbXbIHQ0kznCPxNZRcdLL9a
s8Lhx+w+XXEG2keyW9TQPGmr9XJGJ9AmwPAjmJq5BATMJKMuR27WxKWHB/kWVa0/KlrxLfVgRtyu
3fp9XmW0kqFbK24WXPYj7yTYuaEe3sf9GqRhVvhesHmO29nww2AZdAgpk6kWnZQjz050GE8lT44F
oCo3GTx+merSEgsCimp1VPMNnGGnjg/p9Cbeyqck8yYvjtvFT//mkssXLmAuXHm1xNrvPHHf5JfT
r2f93cilm0VQVs9ujBi0QZfngAVQ0XAweWYKwh9eNvUmzUdlLhysn+g59SDX3/Zza5+DDE8G/ABN
pG7+ycsg0EB5cpXf/ieKKunIpkXL4zz7mMvTlvxWqlbPNUiisijlaFEnH5jME0vFeDr1byvEYzHO
hbSP6MBAJgbLxA5rpPp/RJCvrAxPCMEu1Z5bXOXmkxMe8zPiHu/oJSfMfbTCcoJHW6JftKQX55pz
5IvCYPCSWiK+Xk48DnJDTxf0ould3IyBp+VoJESFyg2UGXQ/fYgBNZVsljbkj8SSRt53Hkr/S//C
RMwNJQUeOUNIps0ohs8+2AWgVpIEaiq7W1AKFin5c+3whxiltQnLbBVpNQHEJL/PEMjj/+fdH2O+
udkkKXjj56D5tVrOkO7YPknyC+7QchlBIuh9bADOiQZ838llJeKNmDC2JKD+AlDW5G9WYUCBj9qP
BYK4Xf5844vX7MNY7f+xJyPyLrVD6qZqhQbm6ahvlhzi3wc/5kpIP8j2c9bkCUDTqz6d7EVzjeer
62LHp4UTn9QC8ZAP6ynb3Fw9BpJI0SdWPLBZCy60BUhrg8uDf0ixab5k1c7OfDb61kGUpqfkfcLL
KLq51A4aJb83vFBkOTrUVMh36yhj8QPWXGyC8H5kEzXMtB16lDJazWBn3tfOii+/LGtvtgcM7qnD
GaR2lYEnqAY9ZbWYMqlz1Lovw+L0Jhc8HVTV/8IxCm9SaJIYjwbKTr2Vp9qBxRDwPdfa6c8xAS35
OmZCpofLNqLZbomLM2PRcc8zpRGT56WYVR3fjjO1UeV8THlPqpJvsk1KmlBQQf5Eg/qe7TWSyJpx
Rrx37P5Pet4Xh1F4kMFiDkGNSiTQ/ZP79Xsl78f6eDKjNTuOe5QV0QVhnsXt9gJ/3CyYyRlEA/C/
rZvhUChQkV6fjQ2A2dZWdh8DvdtB69z4kM02LHOIPuD06C2N8YwkRacfYIVTuNUQK1ELobaJCcog
2h3PFoz0LsL1Zl6OYq2S1pkmBwdi/1z99eU/l8GbYZF+o2vijSeUaw+PiNP/6ykBsXsNNVRVPuB0
CqoJMLtIjZPQOxlRcyVXjxXxDP1p6wZKoFyQATYaPPk3syaZ116uUULRRE2wwS0LrM1IxNbk0ir1
8q6LcCMY+h8cnXisQ7p68Lj3MAzXgSZdzCA1JScMJ63ykMOdA26F+Q4QlMKvF3y5YTO+B3jTey9B
khWtIRzesGgfo/iBOvjtZnWUqye3bA8n2/ySAB87biqZ1dQputTsYr/JRApLjujIH2vahmjqO0Lt
YvfGhJGJo0fT6G3xrDvpz2aBXa58Br3oXZn0So36PyQeiPPgCa13CDKYKj/hegn7OFeKMJdD8S+u
nBIdU/Dp0fikO/TIcTeP/uckx07NRQp0TYK6uh55ju2FZVV3uIpXRpQgUbQsXLJtbOtydNu2Ksl7
J1vAo28APs/hziiSC1n+q047uy/TluA7IN6zv5xkHclYGBD275zPFpZH+VSliQ71DLiD57PTIubI
0NovP/No5RXVxxOLGeuFiJk145hsxxH1MA8SquXfiYDG42Bb81wEXMZ95J1Efvg9oVMH0NWSUjfj
ybxNBENckJVuZNVNLCWOSoYLxgKBuPkJJNBOcnASrIDNYByXq2+l5oHfOEyUlWlEjsPc5SUot8mB
1ydp1C4lwkD5+zEbpGorQJh4iZFhpc65/lQ3n55nu8VNMjwgGu/SU0ZMrR4tkhXtJexuZs6tbqnD
CziliUPycAlzCJbdsF5BS/7qiaJsCpi4B51/U5v/dIrhC62uKi/tFmOwSo7rDwBRRxzKbIyA1G4E
S4mYif4OFt0VQHFiTSRMvZpBzb8fsvDakbuubp/8yN/GnpJcnhXF7L9nPSomzbylIneO3LU+Qj9O
MtILXWdSFU/uTXY/maCwwqSr0GkAUgnVWBBK++z3Aw3MrXEN0Qg+KDyEVl43mQQD29BvpTHILuA6
E6ebPit3fQXOkGBMGvcsXVn/+l8B9eAONQSceSihcpVuqGKpw6W5K+SwV0G+A16b8O+NiYebucMR
ZlZeOnJBDuRMqGYbAflOeHHQ5WgE+oqcDQyDaX7YTl53N98TpqwGjGmahwzI8e0tO/xcFa6Lzy7n
KvZopy63htKx+pF8H1RdTmDrTL2kwJTR410r6L45QjBNYnvkonYVHp9uhOuL6QgjgRJH8mM/UYlP
xqBfwHidRpZ0Kle0yZxIn6Vq6JrU2X6FZ6uaguPlakGrSCPUT3FuNyafYKDKapOhtlNjRQG221Wn
uRg8OpmqwnlMHRjwRILd+WASr3TUhfJMmYN+PZr91ro+R+QzXyA56nCAUnPRnBmlZ+jBwiGkdQq/
OGV6OD0Ys6iJNVz2376LhUW7ERdF2aC72eC7LJ9cwOAyNbLG9UzevVTUqm4Q//w16Ka1I7S+/IVw
zXyT9g3kcHIbushBcNMMBjZJ1YpcB9dEDgtkPeRXTurETvkx374h6W1fV1ghd+b4YPPe6E7IXeYL
lTZ8Yo1iwWpGNHT3lMJQIWu4rR8udyTNgI6DRTWR1VoIa2y2x4pOA6OJM+S+WQ+d3znrfySdx8WX
67YiyjocZA87Rxtc5u6uw3aGsehtl1xXPqN7Y+SGoZ60Z/eNWjp7ol/CDFfUOdi49T06WPW+tFyA
E98j7xpJ5w7ko2zjErI1o3PzLQeeVCkYHpkiGP9kyq+46jEviRZmOMWrdH93QHDzsng92a90ESH8
YdKLkp+kadapKirz9K5bUMxkkflZQmyMCMLCpuZ4yS0jtD87+BW/w5MBz10ahFR/lxV9ZqowRqc4
67iaplXzVcmBbsysFxkrzde+GfOkgO7kHtkDEmmK0YVPE3kmOnq2kYstVxY8C/rrW0dl+rSJKP78
sdOybW+3++AwXbyw8abzrBS5JR0PK6q4G00sQFPc0S+gxG1YrtPqBpYRtWUq5h4y8zgGZFfublXh
cSDqyKuRsWzHYCSbfEpCDSYIowyjp8IVPqQqc7a936DVeI0T6BjbOE9io7dth0ojT0ffRopp1lih
vh62V0cDJYAxFxT6Exa04dasmDdInhge4QAYeTrDQu6oW+DjAFinJl3PT/xIi+6feq1mSMKrgFS6
enh2Q+VCdLJgo1jNfWEy5mKHkfduuhj808qQPL+67yRYp+mSjChPnN11/y5PqxfBMQBh0NPvALpv
wGk71WBHsCq3X00LITUPW3veoZm/ml3T+4aAHVU6uJY29BsIBuvdGd57/UHbTYmtkQAc7UBGZ0Sv
cURGC1XRW6k2U3ErVe6c57/idm7tSl1GKWjnqR0s4QbCwqHn6pf2Vj7uqa1wNiIDfYVOepDpegWM
Jkm/S3fyZnBWlmJMH/74OzLP+PerkFTDGkWQf5MIeVlBsjqkpezPhYbxuOVXzmKfGZ+RsY8qvxA9
RrUhzxllDAto+YIKujnc/fBViU8JPpi/fLDKtEBrP4e5TIIuNk61BxjgAYwuaZywL/ljNgSs/FJ+
MCn5mPBNZTqM2p0tfQ+gzI+8Uh9JHWd5yWZDg0RtJoTr2BRnL+ab+OWC7vZAwLwfB1OW+bI/FdeH
Um7ZJFmD7zcuBqFsKkkYdLB6Kxb1ro0C5cIe6BHSr0l7pt9/ogyletj0ZvJUNWa9uzJju4q4ZFRN
6O8bdv8EZPFO/Cac8MzDBKKdse69Lv9eYonbnujgLKxOINpVKqjYrJXmVVBbB6Tp5mJ/W6nyjj9O
ajMgsSe7c+GyKnmNBVr87AkbngBRee1lKr0S3n679AMy7c6CYg3WWUEbDoQth1LwRQnO6X3SAoCt
pwxPmvWISm3OuM5O8r9Am3pYPrA83NFezHJMtbyITEvIO6dD7sy2C+Idr+A9dny+qXG2SYmnj3ty
DAie2eOoo4tDVzkZDjJU2AMeteUzzAVX67Kzp3BK05NmItQIk6ffpFfWP24D3c6JWRXXvTA3Bam+
LbJnqpB8P6aB+xnwY4YPm1mAd9KGLz7du+J/Z+CiO1nqKGIxlPmnlCN0jogqdoanRfbtHEEjQL+8
OadKmeH/200lUMzVDml8qMIElYnclZZgBWALWvgKQtoAwrIeo75ZiPi0qy9ehPosDFKAXSrz6byj
2c1v6gG2l7+HTMXx8aJx4lMpc71Fsb1wD30sW9BuntJSLs/D8f6KI2nSUryI7dRvK+pBpn2EXKfE
6wMdC28bBz92RurUpocE88/03NRLy/Hh2PT3oGrO1Dhsht1XzrJVKwqxpkDMTrzn/PQ+2IX7VV4g
f1A+ptB3z1qz+tZBTSIammB11Z1Cwr0sPzPeuOwvJZOQCMmOpZ/zIpdSCPhA2e3YBfqd83AXl9kr
+o51CMCs8XN6G35WkLkWmkbRoa9SQd/oWsrei/a88erafwBcuSsxVaTtqQb7FLf/aHuyX05ZdyZO
uJ+kYUyRIiUMfXVJVYyly4tluax8j8GZ75Ywk62poVrH7D2Fj2FeVkJyMZFe2Lq0RoFYl0n93npX
AohlpPeiRVpzOhu5JPUemmIwmfMbjmlorVOZVEwEHMaQKANPUA/rdMpIC5fPBsiYm/I7NZ2Sc9Y8
W7BFKSIjyVEp3Eg6U0kpdtzsJhL4CE7u35SlFpVtjjyfitKEFDTOI3e9X9/xU4nIx5RVgQCIG87s
IE2QArO1k18zCh8IOGRkpcSWpmXWyNWbf+ACR0LGwlL6ZaxWYK2C98iV7KRMDVEWwCJBkgGXdPMe
oda9LYgRs6OmQN3ldQ9YR7brO4iRsZOwkQBrFoYsboYhE5gnwn9w+P1anf4u5/Wk6ouNksHEYrL/
F+uLekblsTnJ2yinlQVS07BPT2fVKLBwsMLdn4BeBi43zk3yVv0NV1JsZC4G0ERXqVCpykNpdMMg
cmOBoJmnVHBxaFWRzhx3yI6hn597gAXm0f0hxWq4++jHNOifVsb2SJsJM/c1BSZyFJwFC5pejlZI
QNiAdA/YCclQmxGFMiOSglHf1pQ9e2uiJrc6x67bxUlExyM+PdBS07kB4mO39AlcX+YUzE0D7+sO
z+8A0gUhZPdgeSiM5YdtHyac5wOrMNon59PcwiidcY++RsF+9kXhIQr2Q9bUYGPjjL6GfmW8ZuLq
ag1l68RHuMrXgoWomkUItYDq3q6N4YPa54fhAQVaAzKxbKtORapaBuT6j36qA7rYd44lQual2lHf
i88YksXFxCnTF9sxfxxKrq9p1rBfG2ARPh7hQF1TZayQqLRAQziA+tzFxlJ0NdIrMwBXgOmGZ55F
/NlGCJC4BH3cWwMud2kRBncUehkTVPQ9vEpih6jQtfUhGoB064zX8DW6gdpriAYRWAKVX2Lu4FZq
6XPMA1CqftBKtXQeLN5TpNS/0jUTC4SEzO3cwN8drFfyBJ6O3TObDlcPVYqxKBgYo48LpOX1tRzr
S/WtNatuQBAp/qN92rcA0hMLwXN9Knq2YAp2aQBOOuVSoC8rE7fWqVTkwnWhQQ5xuiAnaKa/8GOC
gt6g085pJieZ9Ej+e/zMgNO0gqoEknoNFVKG9ONVQTtPxrYbrWfxYXeQNebXHIpl+bemdXI0OYGP
cvDK1kQfqQEysBFCxzYmRyVqAdoguRMNwm4JM3woYA2ijx3ipAmRXgIR5SCa01fsD9U0VOWLgmI1
TI/z8D4bmrmnicofY2l0MASK9/L9iiYSh8Mi31KMoiQBpYrZRBwnC83qDDcgIDYFWfElyUYs19Ft
uokIREoBiEUwqyO/WRD/S+O5eCt4Jm09IqM2Hn8RXkojkcFbtaP+1upQwcujsXL6j838iDDr+9Lu
AFaAUNez5yTzXeeB6aBwo90wvxDhvPxI8XLW0XfV9EipqygvceWnSZybxN+UV6eDADFgaplL3Q6r
JGNugMrA989V9YHCb6w0w+MDG3cI6auEa2zlqMqp+AgmNyzJyLKzeL13oQWByIgTaAJltUrnlU10
LgvIhjWXlW4TK7qC+CmoU3O8MrN/uzTfMdIZO4zhhXLVWQAojKhi8WQedYDZe8dcoI0tx7FOy0T0
YGO2OHoazJUeImJLgSl62kAhwVcu4KRbXO1VM1dB3aX4wAXx9MwsTEWY0pN73lEfPEkaGQZNp1Qx
OV4HSOBdcLUFb6xOQA4RVGil7h2uzVAXKPdtUce1ZLZudt5K4pDWg0alPJ0hlPlF637eTlPmKufR
yEes87eEHQbZkOJSawelgQt5NvPA5Pi1cXzsrN9cl+rDjiUVZjL5EfF0uUOQWqS0ksBYj7wktJlP
7LtnL+bVHZQnQcZzgFloaeg9wJeorrYpSBjQJp3ifazpKV/N9LPfmstO+aIY3+ks/IIJyD6rjnzb
S/GPA0Uil3vGnastB7nS4iyYrKT0cnhjxt5vrcPLzgXfkzg5kJSC0lKzEYjnXSJI8BP6pmqjyYsM
T1X9ElXpqJXgiSKzMoBDUMGEFj1+Gbz/NZgwI4OBR++ep0tuo4frQVcdpoeT1WkoIhz6F6eFbmCU
r63inch4cEwFNy0C9fqWcSsHGYa7U4lb/0fLc78aajPY+ssc2f94E8ZqELkolIKn8wNaqfqonWei
VX4RVrcJKTKfdz4gyBPzTubf7wTmNpZyMYIkeXNo26lrMh+g6M2EeKMro4vmopGOPtg18Av4SyQ/
K2/bk3hTPC0JdwtjUBvjLZCV2Z4umq5f579E1cb4ttTo3Ntq3RLvul2IZnx3I3xMqCFU5H4GkGqN
AVpbNVNKf5Fx8NYxKOdMdYtbHm0ny7hZUi0+hNXVt0/uwkuPVf3z7vNMcNgbG9wZ+nU0Clu1U9AC
Z6yOeCgRxAQe7GQU4/WcMeGmy7VS5XhaghZDef1ciR1J2gkQm5W9oVXoCjGJdj+GhD/c2r+Pcxz+
tryAcQuiV+3n4ubP8KaeSQpOuW+CidsvYfqMzLq7iMVo+/dO64fsID35c6L1SpX5mHgi1i2FwkIG
Py6Ssirxiy5tTu5hSXuIL3Qbc3MeT2iLmZN0fO+KyXsnBJZbZLWy4/dnDFus7Dm5yNaO62lbXY7O
OToGzCqX1RdD8/t3vt+FTjU8ZbolJXvRK09EeVoUgi1O/a5WZab/i19Wv3A6Yq9IIh9tVtaxQupO
21aBchP0aMCpdGFMc0H/94LEsUhpAu8w0qgGLim6X4l9AOft4L4K5M0puu1BC2sXypU9G4j0v3vw
L799US6aJfBVygHA37bf4Yecq7pekCfPoT7W32PjCKcOvafsYzQsfvLNISE3XFHL0ZZy9QuDwJG/
VM/N6KjqkoS+G9sGBudJB2WubBjbQ3y/CM6m1pMaQA6f55cG/QPwpxvSE5YQ+6x/5kxnCBGWne4C
DB4R2GlNYFnO1BpuPutzK1L7V+fdHmsOQLeBL6hS+CyhkeEIwK9fh9z2ZL/W1lmjtTgwsq0PPMSd
Ah5bwMPSVlnNZOGaX4bOPph4yyKTZtTIllQa5pyg2GJrxI8yX/IpMofIaslGQ0yBm8hWW3u5mVAB
yPAbIiqbeb3TSwjI9bvtTihmOYBicd2Ybbiau/jNhBPmzO7b1JvMFnVSWYwf2LG8UD4LKc5XhMSL
CS+HjgErqaPF5s4677dgnex929bJe94XyldWJOQvwitMq27wUnnnlGS55uB1G1Kwvr7SL6Wz85VK
jLKXR61WLM4Rvr6VwXQ8/gbpIXr0dWXD3HlITkMZwTN/AuwGALZxmJ76Yo55iRhaJic9zzJAysCG
6a/cjT4BTxp3RAs2xmVWzQD/4WxqmBLnl7kfnhhnlo3SyH7vc5HBS0teTCMZ2940PhMO1MQJvBXU
jGlTV6vY6Y5BVzCuJi+ukzXecBHZKZTjIz0LhrHb0zE4CXqEAHGhfmZ5P19fwDcj1qXvd8Ktec0k
Vm97ePYVHRlfq0mYAdqDq6jrrj1tO+CikBWmJMpd5HkhI1MiCw5IZR4uTom+IJOEiYfEnGZvCYWU
BsCJVUndUU1Nnw5XvE6f5GRuMJgYWitztCPZFVt65Djo+WIvRTm9gJloFgoyxW1i5bJXnBBs29Wh
fkR4JlI1F5v+mfPypkSKDbO3eOM7zmWaJWBlv2I4rggXKOl3FGR8AjhI06179juMUHVFkzWfeE8z
niJaK4u0dAatxiB4JVjh/yVHNB2b9+hw1lI1h9jI3SdlxGeoE0wtpdSWq1N6DGfVe5pBoDQeIBzV
l+F/B2NYKVpzCufUFHIQt6XT7xj9rW8xy1s01GrekGNey7S4lNEf3duWJZSwuT1+eL5eMyv5Xv/x
wKNt9BCUOTUpdOf1sfgNQWdQ3yMEC1r4h+qrw8ZBgVOmDiZhHrNNt/fYLHXfnd3tJKvfygeVDv1v
2DwNJREOwgUmOhItTENOSL7Ex+FNtAGk9XCtOrGlTqGgtKQqtfNoHKKa2rhpgh+ptzVUGAyj8X8k
E+AwDuxt6AkUJ7N0cZMh5Ri6AZxl2p2bGVBze9klgoPsXKApQXrI96Zrb6F9NsGDBu0DKPyzkp9M
7ZK2wXy6UfzeGq+dTF5ZsnvQulVaRCDUA6jJmths2LhshMMJ0jfyKRDogmKXNUnjUkX4X5lCKtSF
IKKb30ch2/Bsx6j+RSFG6lGynqbdF1k0RSWXyfHCj1gVBC3AKEEc6X8ZWR1z9nT8I1y/PCHM0siU
VzIQ+B76osPUlMKS3bgR8bDEWJdde98iHMU63ErvIIG6Vgem97urggQ80l1WntImJ5NL3E2WgdPm
k1rUzU5BpPRFywJI/BcI/XU4Fc5v1H2izfFSuwM1Xnncf/6iWRcvN/Q4ibiM8BiRu1uKAPte4/l2
UJetz2g09kMXBTnKil97kFaggXj+r4ynOrZTZeRZVcJAXw0D+U7QwDdh3Gn6j5A+y1qBQ1Gm+1n6
CQiTT3XOMPdORd/sjXiSLN3BrzAnHd5fFeNvbzy52jRmVV+m2O9vNlLZG6LzvPhUhHhkKNIl0Bwt
EC38DSh79Gjga8cnxhmfw99E8zXaNlBM+HHOICNcCL6oBtLWiRx+NACEr5BYp6l5TRSnVQ7QrFMi
Wj9MKjFuJ44e5jdOW4w7UgB4NthqytACiAk1tVvS82GND5F64R1J6KGQ6ELoTROtEvMYvJO/pDyv
5clFtjjQq05ica9j3r4Wk94FQBGWyyYS8yDALiEGbnmyI2+5WOlyzykFAjGA50t88GsBV7+i7qRv
k9YPAn77YndcZSWCpjL2tawYE8pAZ1iwPT6KM8S8K2/K2GzElcCV0g4VvLFcADsLwmvlZF3vpGwr
ihiYtgBJZo0gRkxlNBKJpRIXCn4OIXeQp7TMTb2oj0kJbiR7Ym9/qW0y/hjYf9ArH/3QNFVf6Bp0
WqJUfOG0pEHuvsyOMbSm4lFA6UUNpAmkOUhSg1czMZTv6P5RnF+rd5TcVKHEe6m5hOYFtVYKI3/a
xXgFmT6cr1z+t3Y6exnrGE8k0u+mIm3LX0kPA/YyisCgLqlNRa4bnYeOgxfVhLGK7vchbX5jWKs1
sFX/MEkRvwMBbMBgYfHA0/skrsX9KibMLNnCsOBgjPhxrW3jChH35ecJhd32f2R8aq3oGxyHrE60
HCFma1b8jV2TCBdGMRGajcOiWgcsImFmjiYZGuaufhFeIt6J0moAoHlcqFbT/LCUCZYt6lWSE5pd
D28ZAzk/WzbSKVb2wLQ4LtYw5ZAcHjZIFoK9wX5iotq2LZVNI8CLEpffmXifXnzNO644F5krHRNZ
6Dt1kn57ewz4GaUwSdQmSDK6f0rAbc95Rs9UsMGoFur/wx78rQZwwJvjkQ7UrKqFLYyKH4Wjbam/
Ui+c8XwQSeuIXlDiuo6zXW9psTJnPorOxGsiGSfroYOj3JqHRslaGrcLPSRNx2bAWfwXdwKDY3hk
hEpzRk886VHH4eaRDCcO1+mktBybYItIU4ZGvl+68TVmCDddwZVoyQJ6IfrevlCJ4SoS6/bsS9uZ
1liiBwfisox2l3inioAUk0r4I4VWpYb8E6KKPAzMnQALiFDzmhO8DEQwccuUzKerqcj1hCryTjfW
FLcvNA98tgHzSXxNT1zkVyjGxlJhjnkiSZ1aaP2HwRJQZal6Hq39cnT3ti7zjsyheYHP5tFfMMXl
Mv+K87CfocxazIXQp3MSwd6ZUG857Uvrxs7KA7OVCDpg55ygQbSAMOE6n/ztvg8ITZxCOxCa6g+W
yoedyASk312l5PnTexlo2+n20URwe65CzFmV7rsjrsCyH6MkJ5ogHYoufP423++SE9k4aN7Pwi37
7p9/JBr/CedegPYp/GWR4LzqHqB5VRAFh4Se+NmijZGN/K7OlFIXgi5t+kRQ5umZewHKyWPRxjcP
0zE5FDtttiFnTF7xzjTxfmLgeg4NOf3BtQpJqARjLANfC9vkD+tJsyDhoUqr2SXlWJPCZC5tEzlb
+zrgaw+pOk488zbugnXRZFHxLVietKAn6Ua1qoV3zQ7xCC8FoJkWDwtnjiwOLhZh4U3OJuVekn0F
zRHqge0hnedFAVnFkur7lZ5cgWCzOWgWz39hHmecWYC91PqmAGidM4ymuxo6WBX1IF/qt7Ziib5z
IjFwHZOmmFVcvIUYx51lx/wYBdvlSrmBH2lVo6HlE9YPtXkz3h5qElkErv2lr3n+ghLte7MHsAZX
ImI1bX8+ksn1eWcWeVY8Ftv1eYhx7Hz0hh1aeTYUa/fYm1iatX8Uik3vH3zqDBLVj6FroN1vWczj
6dSzT59lsIq2dzLQw5cKXSejQO8wT9Av2/eRAu9cjhZa5wM6xlhi1AIyzJqW6asexez3EZMZ93kK
Q1+3DWrDAceYUdHwqzpp6Ngy66rodAvb2TyI+VHFCDdBfUomdB/bOM8qVz76kEJRtd/t4SRSjRbe
HKfRIXTomC+YZv1vHpCp1vsm6Qg6+aRt5lWkXGZm/NPmZD0cQ9b9IQQGuZlmLUhLvEpsUouCtK5l
aD3xI0G6axdg2C5ARsRvHWyT1GgLnvRu0GIQa3p8Zk8tKinb2oG4Z+Ru6rfwMZ0cGHA2qKCcIR2h
Q7/bwhJuiKVytAsxGsdwB8f+v7rvN2pD8Cqv9hBw2Jijux8vl0ONqVvws9qkHZeraQ2hGgTAVCba
VqV3FhIC7WKYbsbOOajZYok2SqcSViM0s32LAayq7xF0UrQDjSz2SWP7/PgPiattAeQkSITta+jb
rE/1R9LfPQPheEj1W0VT9cOW4NnQkZyQRqbHNPR730mNRuklPvjj2Vi+1M7oZIleMAP1JFDjd1k3
9XKyJYlfE7f2CjhGuxg808ehj14tf69Rug3hWXgNpr/7lcxh7UziJQ9yi2Sn0vwzvEcOCxznoVon
RkPJXASrvMiKHI2cf9UEx+Aca94ve7vGz7V5RVBgCIlk9PEuMpIXezqkbicx1B2Lh9X/iAH29pYx
t2iTZJa+5JM8sGfWD0Pog5fgMcAVl/aogG+rxyhYdZqA0jkuI1X9g2P+9HGvx5nfuVlgTWkMx0rH
tYdTkJQLQYEPOaEVVzsBNK2BGgdrkz6jXVkcaDV9yFXcxnf7V2/JtJuTI8eA0/VtnXGxatQgwV2o
3q/jtGyqbf4UK7gJxjDTkdhgGufKM34B36aN2WW2G+gyH/M61X7qRArnS/D3NqgC7kJ7WQ1VRos6
pk5vQwpspVdCStnkJfDR4D2BDkf+4ckD9AHRumuicB31/HwzvOeKopWZv8Hj23gjAhxQpA+N4Vz0
f1td/qAX6BUCdwdnlokX3y8BcDesHWQYH1t4zfZjMtUV4DpkMhMN8a3qjaPq25UzyQ2QN2LL2pH2
LotKcERmCuk0ots58S8natetK1+qHewQiVp9Ttdfj+Q32wIjSfE01MOXHnWoDY/AUUoQsIkyTTj7
+IcKMuz2+rfPvHXLR4FEX7yDKU4ULtJhubXphnyTgJ6yKi2DUCWeWbRHLt5j+GLk/BgCsi9R41Jp
8jy4JRa2z5bxsdkYz97YDc9R27CvEpFKRHsqF/CODTKfYO8579zoXOLKFG60iE0H3yEhhveBjZNj
5vXbHkxotGvivVgBe8L18SvPCx/gtTiLF2V+1FRdc7UfmukbiKOssquqxH7/y0P59ps1utC+kVCr
E4uesmSFEx/o+gdBoQm9e07/KwV50gTykcUllknOhqshROhuRMsANl9lvkwqRBtuHSxzjGA8pJgA
kNNLliWuFJ94XOJiTucPgHF9IluGbdnORTr9ajxkByRrP8QloPhcbHohCiiNexc6cmDOx0exqLUU
6aADiI5X8Mcpuu/MQakh0NetASmp5o9QrdMILX5t45+2v5/rmmR82LdBbOeSoHvU3nUBts2XAWHy
qVfL4Wd3bAHJQDj2zrWJ1aqs8dWl1UlBSrPluwRYbR0yh0A3RWof9eNnsXryC5HTRnsR/Hfj5JBK
UlTHViXkXHbEQg7qQF20TUvjbD3gJrmnTR314zG8G0oN9NoaMFwgnvJovUCtXE53PRBQYe57gf8x
JEdUtCSUmxFTu39R/aDfJg6URS75hgoMnAfzqIUVbu54WUQRvzPe27871ppOURYtVWLeGjoz9Zrj
wBG8W35l3xPVmYrruU1pnmnrUylU+UNuvh7oBCCiYWoxCe4Lz73D5Fh+Ycojh5GT0Edu6op8wyDM
X3ymX1kf9eAXaB9NYPBoNC4zcXOWOfdGWjeyC4VB8m/J1aHZLCGsV3vghysO8WnXDX1R5CeFRvrt
rX82Q09sy+9fMxYAftpz5rsBfaU4ZTT3RKB/aa9U015DlZZnIVw8C0WhtfeFFY2N0sb7xQL00EKL
t5JLasW6c9ewnuST9w4NfNPZQN2POBR8kvFd6jZnqOkYCjItSpOZ7W2pMiqXDUUfPM9xSE80Kznh
xF5JV5IBGQFw9CPACjljZAx0PCSpLYJNVNjmem9hBwILG834WHlO33Vzzl7Ao1ZHVL2Lbjaeo8iu
oXowvyPBuSMLKbBhKw/oZ0mNuJ/GlcZ8I8bFWlWcweAoGvgS79P/eE1kHl+wvxgRVUdOwNQvPgKJ
jFT2LORr0E/L1urmEknweOoqaVp9HCpe8b/aIUtw9WYMhaBxL+9XPoddElpgXa0SagehfH1IE8D+
b9h9GbZvWUlqweFT/vhhRZpqRyk3ALDKqr+YiURPUnjFPEn1T6Z01cfGlFbg+BoTiaDA0qPpJj51
UM7uVA6bEXAuL4YP22gy76BaMI6HldSgtJxpGKiKXNY2uSJL8jsxNQdFJZqtXIVW1y6afltQDbb/
NvQ5lfKX4HwAcN3Zj/NNAzdvhRP0navnq2dLZctK4GcEWd0+4nzlv2yDJxeORxe92UgFOLlfE1A2
HPKoZdjDoTrQ/22D+Gr2q/bS/6QL60nT/cV2en9t0kZ/CIeCHQDvqIYrZYj5l+vl8scT+elTAcn8
M7m9vg22ZOoOxV8q1FMX/cnyndcJiKuY+g89rLlzqJyEzW59UdiRd4PYsREzo8Sk7u+OQO607N49
hokiigfEyVzUfJkiPkp/oDYtu7ZBVvwmoJEhBHfxguULGx14nuWeAB2nMCsOr+hGn02OKZ+rd8Mc
DF9Z/GQ1iFoQ4A7khWUZa8Q5nUG+GugZYYYmh7EgR3RbKX830A8uRphAhJzjCf59oH2OOkUFa7Je
1TnIIymv1tfGVmnQ7xIKqQESSuPDJPM0Sk/YUMO+b7WpK2cHUdY4urvxxgbtw/TU0pYZLNpIL3QK
rUogeETfWoipjpexEwmmJkCkqHTOOBMh/NAObKYmKVev7T+9wwwhs2k6EJelyz/9nK9WiFQ4zHR7
wQ66ksKRbUBWfG/PtR1yEUrS32ABU4XePl1A4eph9oJe5HM6NyNvWSomGzznVOv0a1l5FqKD2Dr2
AFdY8mnEcUjLWmUbHzl0PWCTINMV3t5UxK3iLIqnXOA6UgzDanpthvaJFBDPje4rBbso9s3umY0H
0MPKgLPXVys8U7pX+iNgUO63drfWXHolH34O+intYzP6lMC01axL5BUt188kOgpKsowvWZTQAMj0
KQE8Y5UlDBOkazzr33Pxwtg+hh11El+akKHEgRRscUN5iohQn9A09Ad6fOK7BT/lsDMzm+eEpTTl
a8NdNqegE9EvW5Q//bhylLHeLCGLJoIx6E8ZU6ruZUbIyhiRxLr35LWDXYLx0/QtY/Q7TO2R+no2
v3tOF/lYuEZLW0ek8FbrVUioohkV3tIzTQZNBHn1S5k0EY91ykUGYtTiGBvcnO7HB2TBymi/xGQ3
IL2w/bRi9Vf+kgM+Fz7/mG35Kwwj5VnH9Rq3TBd2Q0noyJW7pkgXpATFF7dQuGLsHwoDL9WXo4I8
GZPjisrnQ0RqMtrLeQ2WEs/lEcYpXLcTRV/14Se1eagwIDa8voWXYPpXdfRGBgISOwrEyqFWyLxK
yD3M9HgObgmJrS0N8A5AvkMCTajb9Ooi6muTYsD4sIAMZGvuewfJhMHYDT9P4mdmOoRUbymI9n72
laRx5FIloJDSUZXvC7FSlnhAsdFjuOIQOrhxcFIBOFbXcmFGQ35ihg4l4B5iF3LdEaXczBtGrZ8v
8QQbKiYSgzXlkt4ZripeSuWibIjJJ3/D6duIp1jtZoyaBIxwzgqh5U/JoZ0yFj9ZLrmlUzJ1ziRZ
+FUigKzqO6mCreX3pldb9Ig28W7uZ3r9Zhl/EU9YbE7QFAjExBGlVHdADo5oK1p3mc7q0BZDjeM+
ZhwsOp0twUo2NVQHmEB7Svsh6aa/hMT6S1+dgUvFiOhTLAeh6M9+NTl+bYZAfhHBZlcjO2QyN+mj
DwDIAoC+b6qX1k/9vCUnldwchOvt4unTO2EVgeWnaEa+a/1ST035L47OF3Wf+IBd/s2d4fFJsqU+
ZrJEoSt9ptdOVXLCKqbrcBJU9sLYUVO+AgBVcKZGcEr5eKshW6bLcItcXgL3Yld6VfB5QDokyPrd
YJNSTCy/1uzWMbixiDo3nLRBRU9nMa/06os3denAqynFeglsuQ5wTX1qwUiLV2Ihm7q0hUbrIOz3
W8rVLiULT2IVogNtVFYMQodycVdl/P3FC2FMklTsscrC4+NHV7x/oEF/dgpWUjQICB/CDlqlN2lo
s9ULehtyRzKaSjixV70K+mm3jNZQ/z4gpY7u1qYpaehJRV/g0i23MFkV4jXzuQokln2bE0aD7lCl
TPm9YyM0cT+EHxFsr90VRQ7QjPduxPHPGkXEHy68fhbOGGsUB903ov75W5v7Z+55yrmSR1bv1A30
A10ExKma/szfaHh26q2b05cQyQ7+yUOPcB8ZsA4j2NSA1lshaCxmIUBo/NKEpByWwqkn6jUneNdp
eHvVJ/Tn4Y43et4Gwm9u+9NHpVNae0cUoOKfmdNEygXr93MRlyEADvphgz80RwO1vPhx6BMHd8aZ
FpA7JFKxNZTHzAwfklcxM+nu6ZIE2L2/47JLqiCnUdRhVreruGhpaxP62MKY5C0tJbI2z+k8F281
UnHAERUJoZeVrbaHaapmEYXcbn151mw7U0DRw1GRRLN0OieLtAO+TYRC3+OHcNiUJLZ4dohabHtz
JA9Y5d8XkWHJwLVUF1hnT7YL5cc9M+8RV8fARKu2NXioaON3OOzZTFyDBniCAviflfZvMiD4QRX7
A8poY0uZ+7CXc/6KdQIx2zekuH2TH6pqGXCucLlAo0FTWQ46Mm9w+WZkn6Kn95v4SSVFoHHTrUL/
FZ57bx7xJrjhjEF1ArqT5oXe+RcbloP85Sdn+s7BK4qWS3GCo6blCjJ+4ECQnjYvLJX9BzAkoSUL
KDHP7XdaSLk+ESwQ9BAQkXPjDlNvgbeodtcvdD1bi5BcItcGDRCaCrQj5PK0v0tCVTOj1KNYevsx
jcM6JhTc8jhJ4cvV5XYLoJIgEWH27AkMeWWsyx7/Jk8/N0e7s5+0OSzUaPM0a2QEo8EZjfUBeUL1
PgswLZvz5SI3K433WvOU9p9H0xZR5evXSkNnAyEwomhzrU6Vj14ciNMH0xvn3YNTysp5c8Nyo4d+
iDBmsJr3gnfXkqRlHYhRgyJ8bXEsvgUGCQJHTziIkVlaopK9YXruLsqXARh+xoxO1hUeKOR96ZLJ
9emOKAhkcEkZ1CncDLtuBr4pkt95lgBJ01tmyjNaHxSJLdEJp3zGulH0jlMcHrp+pHhYZYr4y+qi
48K8nTUlBGb/qd4tUw4fGtzMYCDJgWINolwyel6eUnz9HzgAWelko3u48iijlIGyLTOVUZoEy44z
8DQr/72DxbgC+pClhTKdgXDmT1XAv0P5LCW528qsJXtK4gal1jmIfOazK0uiXb+baV9PsJDdDExK
IEeVdEEMCo/TXReSgKD5Bt7s/i3gjOWZrn1oJkyUpO2Pda4S4/KATeSjKTvUtfi/OHuJJ1B7aSuo
fFWrT5XQmdIUmKNhT3LJj8d47LzsOC2l4vB6J9hAiaDg5MB2m3TdFXAHri3eVxENP9lGFie1OZxX
5K9ygRTD5M/uWfv9aoDKM3meknF//Va46t9KsXZHGDOyEW994EmjzpoV5mJX3bMnhBQcu4p3YG77
vLp1Uj9KViFsv996rTGVgNw1POXd27OSWvBn73ydJ3jmPVy4hWzeYhxzIGWAOIv94ZEwtspQW/67
FalzUN7293Ff89pvTZf7C2yCSSfOYkAuK3OvlKtSLxDp/uRFZXKyRJ77bzTadCbpn923G6WVoGBx
757JDCGkNKBkWycIEuOCj4x9yIhGJp//mcxxwpXGmQdNpKL0f3V/eEHR/W5ymT2+zTp56iVY1zdj
Y4qdYfKFalW4B419K/1/QbPxZCV3qoPLRJAM+SB6NunOeh/EDnIEdxzc9bkZrwf+xHisujU79xAk
Ay4PeInH15/0PM2Y8uxx7YWvuZtTqCAHo/Wts1hMqlJFIGL2TmuinO0Xtx86KFfALJU++b3XLXak
pSp5LSDsoV2XIPS8D644RhzOeW/X+hJC2aagTaP/3WOIjBdTAlN1aUq1GwTJsOkNQXsSEnlet55U
U116ErWyi+2m/2WqpD5aeZYFHS94ycw/8xefBXfnVC70CYJlds7bugI9acVRrnl+Mr6fbX+H6QqI
lQRh4a1XCukQKpe2VjUt4VXFRwui9OeeVt52gMF97l4uz0qDVehfj370/Pokw0Owj3/wqxNWEWt0
jh4C7/F/dNbEEI06+ggrFaBlaEDkiIQZBN9FUif2RifmYTCWm6xOhfzgxsRS9brOjlstjLdVD0Iv
n10IE8me1Vh4CU7rwqwOi/MlWwO3et1N8JFW7izpYxBw5alfDumWU4hfEemEB+vC3IxM5Gx8eNdS
quC2qeTJsqUSEf+C99sh69jmGAAGpkynfFGUdkRB9DKY28WFjkxuVRK9+AVFZx7YImv+NgWoJfdY
ATFsXaTLz5XO+O63hT6CgytBjOH4u5SbJq6UwYoX1YfvBYn/TBAgs3zrDWB/3enw83d5SBPiJFZx
4wHq1PUmUPw5RFA59mPsogIFi8/nDLBGfdcgDwfW5gexd2q2IkPAMU6BBHrIHbVr5AVbX00RdmFd
byQtdT5quj0uowD9ybnNZMTMyx47y6DjM3MJXrskleARD1H/w+iESm/zERVsl94kfIf5RN0lKZXO
XtTydfLfF2SEVhs1gX/at5+mwVWmvx/tELP03gK7jVULwXPu6L/mY7/pzluUw+jvjB5Wz+oqOFnz
JJfeeMXgEeil+Lgd7gKmuIS+TOVTCnEvrc+wFxkUqdkYFK8ITkk2DyXY8ctPRSj+gIK4P/BabK+w
Ad5tyx41EX0OMBgahU2dEm+8ZUAC6cSZ5DdWbJHSg7kTuz4ynhOoLYOyHUx8TPWByzkdPMJ5X42r
sHIL6P0Om/cQSbT9+RKsZ07sKW7yMEEctFs0P2HXbBJS0zdG7q/kWOEBbKoWeFMbdFGs3Q0d26SK
ecO+M4VgAq+zpVLY73vQn2MAHCw4j123lQdW4R0NwmcL1m+6T/t1PtaCsUpRcy0R+UVwxE3HFV/2
EdwT05SjTzpXgiJPHIQN8QBODDDJyeroos0EQqqKpZ4+FHLpAF+p6e3uhspRNtifPTotlBtCBO0w
rQdkQGuGqJFEyppjky7VibPwRz1uFMQYfMAHrOdLz4+MPyMTLVatpFai8uWwIUf52WARhtyhERd1
ngfmt7Z7QVvaUaaxeqTLBXROYWJqPC3u9gxAQlM6bLIdgSYkm5sOHMltDGAK7LzYFDY6VYgU/tYu
4hjxeMqRJILC33QWC88+wzqDGBBSL01mZW6RMwdCgNKI0Kqcah/t83ZbFp8Xu2G0gRYAu1v/xuHg
cDxdwz5AcApcUNpMxgkKCaW+5fP9b/U3DlwYHvjr9aO2ZxP+5TdNrKDgM6mN/hjrvkc/wqpsiGCV
vZIT5thOSI5xDyINww0SX+DXp22pXgAlKz2Havm75pX0NK1iMYn3ShG+GwjpUPnyAJKxF7HcwrLX
9PJPzSweuAAFCIh/9wKBegOUUvghmxPN4ZBSFDh3kRr4wWXj442L+y3KWvruRl+croy6LIriWi1Q
f3gkQz7kcSn/72Da/Cs5+kaK+W/oKNPpq1rBZb5nr1yZ9ZXzowAXY4UOmC6iO+CZulCWMHyKstwi
DwBx3NYNs1/uaUoZg9+JPJ2r1gD1SChJeMM1F03xntQlU4qXTIZjXKdki+2+M1AftqSi8CjY7U5O
n71FqfGuLraYiOFZQrwYt291jeHuACUaGBTgpUDvrYfj2TdPJ98QE5Olcksqj6D2XK9Wc9C8gZ1T
oiDL9WkdIGOyRYZqd3vzjzdVorgFsUyxco+7woNwlZSwqxQiZYEDn1tlXyD/zO/15ZbpXM8dI9ar
Pv0A9ZJVxTW24MbPo3nWvrXAMVdCIbT1iR3k3h8YoXF3jaB5L30omwEThwNY0GuJsVwHdTRZHMZG
5XygBJ18CWKHiloNv41AaRA5OnAd3cdfQEz/S+5FMcs5CNemw9lsUO7pbNZrRdPkzc3APKzm+ddS
+ooQGQKzMBfYvVjGsZGJEMZG/GaMy5FvAJAU62zrNX5wdk8pc/e8ODOJ32TzWaI0PzHaf7+y1sGm
sGhdUF2w5ZP0JH7yCKGrYu9cse5Dsbzvppv8T+2mvUoleqQE2DoQUYz7HgYfQG18E1pcI2u8fve5
bkrXfisGokYAUNsSx0PayRLBHjNrBZmAF1I4vMm6xw+yf37Oo4j//Pf0toM6hPslI5Njr1zgB6lK
XDqtW6xJli2rq2S0lwBP68OzA7HiNtGCgGo7m+rN5teBsIoxHX/AAftrsEDsBMjHUTXCDn7HD2RM
9MCeTyYy4mtUw4cYl8mlO3OnSEhfl9VOtEH6c0wBg+JSDjDVoM9yJiOwIXzuks/76JAHNWCOPwDy
UE2xFn454nC/jj+o1P9QIYIXvI75vfchMTqjhd13URSpr9fh/+mSdgOfGWKgidcNQ/LZ4rulzLZL
4qTcuYaCi9WH+kUBpcrVYCZu3dVeKk7YNBm8P3lZfQ9zKzanHXMpl3XnIM7BiBYq3BNUgrqceQwF
W5JTTOvM7VKWEWXjeTpqezs7xZlG9P5lnA6e8UcV40gxZFMYz7XnpL6Kkvo6Jg5uCIuiGt90gFD0
viP010YQcZ/+9SSjWUJaqJf2D8CN8TvNrZtsBWdKdEw0jmSDsmqGF+o7+iGP7WtKwuJl92X2aeeO
NSZ6GckAjCeNnUO+wIf8Ym8nxIdw3fmpJiyAJuuX067DDayeAcUQa7sQaBRk5aP72owv/BQTMdbE
ePCePLoIMNyVLP4mFVPOhap+2UQA0kj8LE1DjFkRNMi6bs9y3skfA5igFtn9ibhtf/52JRXbPGDg
An2NBO3qd19TV+TOpvs9k+2Fxq5q+8zlbBDBi54voOtH891+UufhaznOT4I5QlzYYM5wGcYU9Q6q
UfkPK7daXQHawroOa7ddGYQKn3VwFc6/MPlk9fz0Aw/VnxF+0g9ZcERzjeBkqjBA8efzq8CdPkFU
z3YNxD8jG2wE3ocg5Yzlr4CIyhgfQASfiE2vgan5PerAzlYsYU5D7yyeYGojczY0QxArKkh/OamQ
GgHEm2J46PwruLnu+YJ8EUu1QAhEiNj8En+7H9jEYsSCMl9HLI5SPJRDpxPNmymZt479ezEKs7Mz
0SlbG8L2VYhyAN5Ute6DULeEyj/UkTmQlxcGRrtI6ozEWNMLjM+BYYy4JLoIjcRw2oCBeu5sUVsl
6IkUwWoeK4bXcIrvAsnAdnB2Yt8c0bj/WFH4feOctpDQMscQDSt1SgfhuRfusPAs7mlUpeoSqMxY
bEOkvv6G+JIZwTEMkPH9RSqTl7Z6k/kJxW3GmsIOFfpyz4Sg6vuaKlLCkIVaAF5klucX50MgtvR7
W0FZgZlZmudk8X7qo6aitzK9GTLfgPW8h+cQq7VRmB+Ij7xLIWbRhGqd6ys9JMncdu1NKyIPsaS0
MEC+TuBMtyyeBdTdQqFWF4AMhIjGsXcKGSufkhmNtiwFRYCUmaTJZS7S3rbA8UO+Q4zmzopxEdO/
OAzg3EPu2Yrf3sgwSqXekvwkHeLZStEPGalwN2pCB/la4zn+PYaBqwms6LGi4sjePaUkzDrd7Aew
JjHAkhnsONufQCu0vxcMbvCpkN9xpkrJG59OOLBm7Xig36YhBWCZwv2pmbwxYEbddcmrRHTDCEbs
KQEAEeHNGzD10xLXAdQkNDswLy2Q00m7CeeDtm5J3JfVgbfe5leEMI+VU76bkNj8a+uYLh24b2aL
AM+BX47GsNPlaYW6Uc0qU5ljjLucS+2H3yrZbZ50izhOJnHdWEaq6XHnNrOR73CQCeYYaMGIP0OI
QOetOoex0Xer1RNb2910BZJ7mrU1mSAs6+8RksRNEjTeeDrYvThactwD+ZA6Pc7UaAMx4Q7duO+c
PpGoQGuFRFvfhWYz1Ej+dNeCI40ir5fo81nRmWIaS++PxAnpK4F34lONEA6iFCCQOWyWmrvobFLy
wmAk0NabEdrME+0eKLdLo6/v81LJk8AZ2/RaFx5h6mfzEchBCEMgRUVa4aqMb/FCpit3BItSQSWn
AFHxtLesyPec+iaRNaxOYDkCFvVdM46ZLsw34qSnYi2K6n9onapIGajEM/e99CejJu/i5zrq5J4c
9KgeBy3Y1w1JW7mcTwe2AABifZW8l7q1s/JhoKXvOMDmV1+q01W0hNZg443s0Sa9iE75zNhBol1x
n3xeyAyJHYYbyqhQ8aa+vEu56gFJsIxfzkqUyXCZaFk3hoHEEyB8ZBEE7IM85iX8z7Z2yO8dd3Zy
k+vKMDdGG3tJunaPX/ZFLlhAjjK2BUHO8bUkjcR0FxPAF9RaBbMglRS3zSPGl/Otaj1MtL65LGS4
fU/Jx3ynPUlsvzXhqUSQqSNEjG/NDgYYcaFLx+xwWRvvQtrHUjlsyCPaTG+JfVG9ICQUbzxgn5m/
uECcjlwtqAONLUG2agarCEKtl73UCu3tgkD/HShet5nX+M1GSVEzJhMswYnXNYWbyytNPcn/OevB
4NCO2bGDxh37/JjCH1fcVjyBl34MYc1p4Xz77+J32WMysNXAIlAro5OxNE6jZIqeaqmqzxe82jTF
3nPzFWCDsoElxuP/+I0J0eA6w9diTl/aCo4MEJ/SMnEUqv+s90HSHYWTb0U/gy0GvM40X7P76xEL
AG4c13nAz3ySA/D1ljh4fGVKWDT27T+pypb2M0dclZfYV19A4J6HtRUxHJHergTrYs9ixnhmY/4k
71LgXCZjL2zXEqK1Y1ceYtm0FwucrsSnRwXblThedOj16NFe6/3ktl1b+JLk5E1V6W8UTaFSIkfS
tMrBGga00wapnMK1PGjOahEB6Gwyv9Kq4SJ/gBbPeSgCfMx42GOSFJ5DlhsI2pxGRCc6EtMkOwxQ
hHdsbt7pGiwhiglMQezC1hASJfab4oknOm5XKlGtZEawtequq0aQhmUWWkUVZkCxXXl6Gsaay0QU
iNAmQAM7TZNKY4RcaGYtCn0mnE59ZYmsQ9dWM5T6V0rGpR8OCpGb+OQCD4iT5DcNU9DnEvO9Pd7o
lZqHuD9DT3HkFahfbk6mpaj2pcHIoj6JK2ierMYcfy1OqyxctCj8r87+GaJ0o5Kuft/RYdN2LQN5
P3MSeoTPIZCkV7L97gl7l6qF+O6aep/9aB/RIMvXna51oz5BPQOcO72XPeftGVcLqzX7MVreGhiP
MeDBd2/w5G0uUcp7jacIEhnbnuaQQYJJIbh+kePZ7XU/fyRw3nXIvUP4Ik3gMMjOUuQjeRRdmjCR
zQTeRwYulv8FLawsR0cK/tj5ni1wg1fUrNX7tDgAo9I4kDcBSg0LDN3e3lqyrzIYilBz07pYe4dh
z9KZFxKbpFaA9j9A9xjzjexRBOmF71r4eZ+ZocoapcvXjlZ20Pki3CtVemEz9RjtO0xJ3ctpUHA8
JhOb11Vx1O/gfgISsCdhSdyScvpwFYfASu9mQQMk6NXZnaaPVP0ONaZ756mDEfvPpaEW+KBeco2l
IPdaZZOVrDIqCLhfwm5nUueMwV76297tUxOFT3NnZkff/X1ssf9EZz7R0EFd8kgbOTPjSfvQsh1S
MsOtmiXObga36V09pLRDf1MWNWCOuqzrjJO5VuAmHac+ZV2z7RqmCuDQIZj712QFTfF+MAvaiA8m
pBhff9PTTYv6vXjAzlwxte8mghFffYNqBiWnlKc+BOQQcdM5to3+553ArmCdePJZCQfEg3DqokO/
NXJp40pGtD5HMGphjp4AMoZ6s7W/hkJbW0CNg2gEVvVl1jlx6n7+FFjq+mZ2xcu3rhFex6UDK2IB
NxpMnYJ0pv8i6QS1arfMBZSylNCfl2GBkDlSDPBOXiImFl8nGn1oShhHJMsqe+9ZJbIoawVon+xJ
s11/tFSKGSkSTPsoPI6QXKHjmRFdEebd++uR2WpOp8+T9Mk2alJO3I/4y913ex5/6B/KwMDUK3nv
zS+h39XtaN7tFdHqtS33cGmQue6Xphlo4++Jzgi3dkt4+fhM2mxQ9ZJE8o9N/bEm2dvvvPUp0cjn
e2oLw9acGDBVYJkfoTrS4lNK2YxbWi2s0+oPhIhHGFazGvSyF++TG4L7QYgjAPn0MhleOA1GMbur
khaL/qQaJccc1XCJElE4hEdPQf3cdxL7LFIIvCQJy/DxzWlgg0KMa0bVtz7+p3azONssfApb9k/6
CKiGLgTBX12030zjKbumYsnyZBLzXKl9/86v8CST0VT/DFvCqdA6Md2sniPMfEJPhpMOJQMlHk9V
O23QLTWleB5LMkJ4bWrVDSKAv1X+dGU0bppK1+8AIv4G6j2bsa36O979Gup8T74Yk+1f8bA/NJ9l
w9KUFP0HJhO4FFYLXe+13p0J2P1A0e6Z7jKNGJoJ+aZmHMtWnuRKC315HOLp8KPvChYs20OqjEHc
k//Fce5rqJYZuIicKjb1d1kP+aEd3dkP1gisqQqZFZhJhhTG7UIVbpxhKdfmRMbAWS7b7GjrKysk
sYKND6kBSB4OVpGNgzOOi0TGOrvbn1JUpgZ2jxlV2oFP5OXfM1nWNA2kHzykkGz+XZi4fBrdsz7n
F1HiZE+DSPFqLgo4y5C4BeYqcMBlj6nOXFetlG4kbVCSwW1c9wn43GanIwVXUFZbgOGeA3mfXlo+
Xha/4fJYQLj6J80B4DHvRExCn1sbk7X8dL/piPL/WnjGnban7WDoVP5M9+sth08V4Z0WeTa42Zgz
VaOHxY6bKRn1PXouc44OaX8MBXW+GJget39L9bH2Q+zuHtMUYiAKsKmpnD1ebVVb4CEaSgCk+Diu
9Lvg5x064X4n8cSYo8SApfaObKF1hhl/k5/xh0gcRPOsjMl1GWD+BsOsvD0+ixTgq6fZwEkupmBr
OkKhv+ig8RPcJxDOmBhdkZFDDq0zZ32vTJwlJrDO18Lymg7UX5jFxl/tpc8+dcBIteK7pHfCwOPq
VutRuqq2O+WHnUtbJHlpcSVUoDNwYkEw8S/u34HxUsVtKNC7LercaokZDkursbniMrvfZXooasfy
YOUBk0xmTULrFVF/jeAPNxzJk3hRSrULqZVMhwdCIQQf/bMWslMz7IsjYyBJxLUOGJPSnIbqSaCq
r9a7qsNmuZJZ8YIBT3nMQZ6+yqczLW3XQ1N/4+KLRHpYfcIoIyshGy6+QcTgfiRjoVryuOJeXDji
ufDMwdegZKIJFTdKJSlSZ/OHtYQ+L/BptAQ9gdNUF03Hit93YbC3scME927FqmK1YNmbGXB1r+cM
iB6tYfccix6t+3PQu52BXU+r4tgJn1Q16pYt9T6EmuYGV/2Qp82ppknw4BIVNA4TKNjaNIf4gELE
ZWxm/YT/31jF0fgffFLsBtP0s4ZmjZjGhuq7LbNPv0FKpdDWTMf5GZ1UqqP4SZkbfZwJtFKxgjp5
6DoyupFGH7UevKlmw6yWYZpPbd9hNJdmIDB6LifMXm9xJSGvMIfBZwcaf81Sk9rZ2eAzMpr/BsCs
oYJZcDlD/fGNM7na4HoRoRDikE8lMk4HmOhqr8L/E72jWEjd/RuGZR0h8iJTV/tkTLZSlAW8BRIQ
BRlJLzRtNu2TlveSdzgYVI8/rxF1hS409YO9rocJRSStIukqH14skZ+q5BvBegYSoKjwTQKNSt/R
FqZZtBSFNYY8wB0c1G12pM1cOsssLXKnq9d8o/gzVHZwE87WsasGSVgoHqBTomk9OCHvy6muV7HU
RHN9gzyIveHWatDAUqMjUpO1IY+28qHNRhE1RTzv7fGk/ttcavzE6gaq2V9U2/ecnwxGgdplLrpL
vDWAmVWHaW+Yt6Z8TjQk39EU8UOvns5JS8ivkdkuTfdK9l9zyloRNw0WXbIakn/H1ufhqYy7cFR7
TgKYAH5IcwqR8Un/CibBZdwRGsMOXliOUQ6Ztgtxr+d/qWrnLK3+fZOvK4DeHcKstg2sHiVnZD87
D9njTKLeOC9+gEZiMkMB4DEjvzjVwv4bb6lwPFTi9gdAVBPWcAg5zUqWGSnmnUtfaB7LD3YIsVaZ
RwxkPsIUbs2R52B/9VoYVrvgS1ez16qUrIKRknXSpUgnpq5qscWabj5dbxrisZJ/9YBAtTIVEFkp
9wqb/FU8cYq6LNxAGbPYGwAik0hXEc4p+sIcQW+mooUA1Y5II5k2bDo/+9mjpB6wXhZNbcjlJ3q5
5qKIM8g62r9zgur7MRGt9+cpJoHV2WFYTJo/VrvQqALk8DJL3YZAgJO3e81rbJIcZNlTEtKrbo/J
pcXOIEmbeVNBKUu0IdttbLKvzdI15qaOp0wAceKwLv5KyFEEdSoY6lVAGtflnEaT+v4ngoUpBAHx
jf46eBxiwi/MhxXyRC0SqSw8Kb1Y6B5Cv0NXB8/GxB0e65bF+QkOzxzovwJ5qt8n9gU3PI2W5rUs
cAIBMqpRj3dW5hzpR8idee4e/orL+AXapYrVQjgNA408KVeqomBkYkTGpN+mOF9fqYfFOHQIEg0r
vicMP57wq37wpJdbJTmbjwWk8LTjr9tYsULFnVTy2T4zv7vaxVUVv/g9vA+23HSknXRCKN7KMlRW
fXwN24fBTjjL/9jiaL3AP0Q/YNsxW6iQUR1pRdGWekANzj0by40qToOaXEIIIN9z0wu1rWnLgprd
zoRi/OrY/EODc+qDF2u0ZmfYVsAhZqladWg6WPaK0w9G3Jm6Wt3SYPS0IwmkDQg/Gu7wieMGjtmi
WyolG76cBqxOfQf/SRxhoguVFOQgRF10or73JlDmHF0k9Sg+bdENDII2xD/nJmbpr/cB3k9ebsP0
FLpXRQyVgTnjSQMrjGA/fh46F/zZJHn5FYu5tBokt01q2TUdEu8ShzdnF/IEl1IijxvqZj9rta4V
lw9KYWnsbkiGnqGXDyvxvlt9HmF3PeKQ7oAuVe0U6RvgfJqZYcD54MBvV4IELCQNeGULDsXnMymL
jo0xqgOztgFv/ENPgOr46iY6eoYBLj5A3Qnw7QG6GBA3lDeAVJoMftIgiQxQP4zVObn5yIjOpgHO
uMM2vvKYuLKPHXxZ4ot4P4KITETegnb5Bp1jNasKCKYEMZdIrRrmIHigmQviLlbCa4+sp7YpyKYg
QSnAfDswHgyol4GDZW/N+lz7MNDd8RQyLwSa1Ra5HCeTdJAhSqhFGLuS675JvP/AitKAsceP0Zy5
wgVF5tvqxEtI4iT2gO1SgyTKTT+kwDRwsJHUlug0C3pcEfN0reY2hXDjWCDJiIIKUQAupHsrdkUn
m600Gq+xBYkjbcIXbdRaNEFC56HrS2fvm/5dCCr9M8diM+jjXTo+/+zSPF8int2GV6T1GBFX/KFh
Ak4NAWC8NyegyoabH5d2u3fFvSFFiJGWbmXYw/ELFoNrkJpzwgnzkCMK5/cYsGTSvdGXwQ7wV2ht
xj00sojx9ugWSN9dM4UAByBsv1ArJctVwMt8lZEUU3pqZYkvrXu+ty9p/C3SKujeBM5F9kd6KuxG
l03P8feXPCgz97pa4CGqn8mGyIg9braEDN9XjYguMVCUG3KErqfHf/W2j5Ja2wJH2TC+zrnbQsnY
anrkbQpoSKR7dHRgaxStEoaCWgGhSzgIdMuFjAHhrQiEOuILKN4ATRpuIL2oJT1cVvr+7ks0PHWr
HvJpthGuAhEXZ8LYn6xjdw2b4sbzbxB95/edRIBdze9mKDuHNMENLR/1e34LrKUTgIZRdyoy/KmH
bZP1g5+Y1G+Imuwv6pdqcMvWFIe5kN5nbCXUqBKNaL1tHk0Ym9/QHzSVAWenTQx6B2RcIU5TWFv1
IBTYsHEBuRQs2FdmJa4XXRz4jPs7DrgYALiUhbjzf+xpg/dHlDziXmlyx4ZN5+//5smWtJMsHHPh
o50WEp5X891atqYT+6x+GZXHIeMxgzwDlSxvBTNiGbRyZzexWgiSXMmbRQq7WK+kRjZsEqhXls4p
hnH5mDZdFVZsC3yORsLEVgd9aOVvKhZ0X+Mhy+F1LdZSx0kq/u+4ZXy/2cAHGYBLbQY7KVdLljCQ
dYQDifBxBLS1+DCi6si4Tu4nNVfH8KviAizTeLpRItJfQbEAKFIZB39BYKbXwPmgklaY7QUQWPAK
gHgX79M16M3SfqATRzSbOM/VMZU3w54kaEF/y+cN2yhdNHDo5vjZMWhUlSN7TBEv28sdyVc10JZX
c/0WD4prANM+aXs+rTWamTfKL4hEIbnenR6jfn9fHQzSc/cXT2eG2nkK7NKR/QdQy7FFecpc55QO
y6mAv5/6IyjIq3oDiKDQeXDpR3VYT7gpuAjqO+9e7gzWSIRN6W4icCh8MP919hbs78Mb5OYNTJ1r
LqxFDePlyeYN/Qzvp2ZcnxAzPMSG7m+QWLQkaq2bUMRsiH4URF19hY5WGPc03B1uHdw0wcGG2mxl
taUGnuihN7m52RARspnfNkseHupBUtuYrxMQxdyX+/ulQ2n2ashJ4dutyTPIoxQ9ILZR5ftAM4Du
IFRcsXKotcKhXX10zNk33BYtz5Ffr+HomOAOsqkxsjiXuU3MKk5o2rISZ6/ZqaRJZMTF2Zcb5yzi
SN19k4iYfrJ0Zz5a73Q3ryfzs69F4JgtyJW2FVIk5RPl+vYnYxQ1Fos77JRUQIDbsSqFZevI7VHv
FARB8Qbz57GkLeNfW12r/Zj2OUQjCYRyI6Z7BLuCkaUh38ERlcBXtTr0tXnPF3m9su2149ulPOts
V5U61KZwCzIypHdm8QVmoEFJ9xQgK/P7WbWjchrEeYfZhS4fMN/ZNIvFTb8HVE+Km7KdXrCNrWBr
x0zoX38He9/GFOOAIfyRfdntxO5MUx6AUdx9HWf95up+jdkYjVZkbGBseR9/zYnTnziu14q/GGrf
GFDqSeuTrlS+grG0XlwB2qP/YBnwR6Phr+KRSk8yz2FNKvhlmcBk6f+WuzU2mZf2+Yj2sLQ3kBP4
nzhq0j/aBsmryqJuLmMADPcxL1DHDlRYuxsCv71rmJMdmSbDxYT9zSQwB8GnNW4LyGtuG90DXPzr
ctanSlyXA9CKde6x1OLhZpMXvocXXtrICkbvU7oNKhbBMyyA0o/C6dOsR+wBbXUcei7AG4DFDspE
btYe7FOxGCUAuyDEi20JsI+yzF2z3J72ZCtkyxYz7gjeHDXzcxMZT1Ta4a18/8YDKGJs7+zMECpL
kGws7xUpvQMFWg7a1068FEQmsLrgG558GNf8N88l4huTipQIeM0D3huJVEJe+wV3XfchHsugtsNN
S28WQxFVw5sgLRY6svO07LzTZtk/KLhJuIPRf3p8MRuGs9OdlUEyQNgGQkyZ6RxZs8LH1tevqVmG
D3c8CBMlYeWghU91W9hLLJqfUfLXFJBY8yYQ3SPHuTbovv+TTwqu9nCb22dhSWCf76JVaGX+DwYT
iE8QKR1970WcSiqE1AdPRlIl/Tnlqp4DNMie1nY/ficcJxhMpiv4M250EF4u9252OvUSuLSdJpj5
P0Lbu20RfqC6dPf5tqhk5k6ZYCDAVHF2vqbMZwgGhknF8Xa3usi/l67bgYh8YugMNf6q2gfrSjhE
Dq8aYJeysvwLrq/ufTw4w3xGFvN+cJGOggkiXtsn8LfSjjVDd1Re24zFgleDap6c7MrcFZA40sz1
jT1W4wr6WzPCPhMlq+YpD+2V3RHegDuWPmM/q5CcLQmQ6pOU6wtAJrtDl0621izuYIgJKftlyd7T
S2/wWhJe6Pmh8fPqEC3SwWoYJTDaH4bAZRqsliXjst30mGJN6rh6sak1Ivw7uAQsyRdocfiee7Cc
5dPynwFBysCWKT3Eym8OHD1j2qFs983/mn6U5tFfIlw4JVCHsALl4qVaSL3AhskaZnGpHduDSwlR
ByvVBUx79cjEogCsuL/h5DPM+Wx8z6vdTQcOXK53Nols0uZ98N6YHGwmx1SM3kTwQCs9rJ3u4zNd
ChRKwISEdKjngOT0N0UoPLt1m9WUGl11O7+fLfLMLkNTrzd/XIyQhW2gaBIEo/AnkwWITTtC5Y+r
mTHS/tfRXykPxz1L1jMttFDOgD7Ni+SSpK42KOHz6pQ5mNo3UHZpQz2Hv1br1RjVAexeQUi2eako
McSganpCMNx/qWzt3s67XxgGN7xySCoYE49ogdFVx9IfWHYcAP8aM8+MtYEzbAtb/4KJjyGPfQe+
8rzUn+uuhH/ol3j6bSF64QJYYtwgrR0Zlgq5gvJRR2BE691E6u77fwWyyX8koWoHSL9yIk2MBDry
SUOPt6hv60fY5lIVuyIYJ2190AbooL/79kKVsx29/blzxrI5YSOZ497PajJsmidg1j3mxkAMeLvf
7jza4hu9dv+bsicsA2e5sbGnUEdGQI3gns532hgjsJx9en7WX2VxBaEozdxQyEcDdTbbfyT7hv1A
tJ0gzowsEQVYbeo/M/B/RkrpmuXDXEpYhhHMhIR8W6GbZdFvoZMS+FSMyUYqCzz9lQjH7aBNoHAQ
2VZtDDZRshugXVvlWxx9UyRK7O8hiICs/e9LEACBitv/9YgiQWOKlbh5cS4O66lpJwblAZTOZA1A
VVPV1E0vwS1ETOSXBZDJ6Fm5GlzbO8X0ZhW130dojDeIZslqclsfTIqKTz4dyhQqXFVp7Mvmy0gC
PY73beRs5C8xzuGiZPsCiWpFXwPLoFaS83NV1JVt+MglxzMcMRHdk9NO0rMttDusI7+aPbx5Uepm
LtDXdiTGD+r+CizpT7G4u7TdYpjFeFtN34gaoOjILOf6ZS0awtjuu/FBocfY117CYW4MzTg+gPmO
/F9i4W2ckzK/6rAIN0ijYzqs8isHxJ+E8bUHGy/2IrLsXy/eO7vltndFehlohTUaxY8Xr/OpL5GG
DBKxBVdQ0KIiLucOn5F4MU8yGJPWTq7Wvg04MKWakXvhKu0JnPV7nsG6FNv4NR6DfL+mzGkl8cPg
0dqhlwtdL73/Xsfsw20YgdqmjyASr5p52LJKHnwKq2V3R7KnvvkDhU/9UYDfnZh+sLIDiYta9n22
Or49PO3r4k3ihjyku9PO4pfJMJZPLMJvQm89H+FYmnCmey3USneDja01uuaXlsA0gA6OdrJiXbF+
wXVoIs2tN0O1BpMxdl5YIWwuMflm8E+OO5hW0f0H5A5vzU4ub/W4IvQJW64OCsp0LQBIgyp+XmCy
lmT785+Z3Di/fIBNVbBPqKmCEZ8ZuLX5SFTHSUePsSgj0YMHOlW49DME8Oub94mbCHPKu1IB0SZj
Iql+KCeqEr+NeL5PSyq0sMUdyF7JuTAlbm+dCjR9LlGiott1JKtnRhfar+U2bn8mh5XjBuUorgY/
F5DxGg2ohLtKPyZWA2CQ8pKBnQ8VUbXeCLN6czJTdj/ie1XIjp2J+XsIsEMwHaSampupTIm5Itlw
rBoxKCuCbEYXRMosd//+cVxT6dRP9iyo702kwE+1VDmJLZR1ZJXRYc72MmqowBpheK+V9oQhsJbe
PC77gdMHufuV0we7VnxtFuTAAZWJedK3idG7A5yYnmHAuNFbh/y5rC/E87kzL/zq2BGbsfevjR9G
INsKwREAqTfKA5BHqn11lhfFk3lBDjwm6bdVbbZdy/fiki+dH8n7EUb+JoeQO8Mp9BqPjAcOyIku
PLDI1pE1Fk2sWON0qiERP7z4TGUzGLzktRADg+P8mEQr/KAsgw0wyAfrMkbj47KNY30iKm8iw0BD
D/hMdSTfc5E0zWbGxjnK3slAGnDLRCM7Exfz+48DWjeVUlTkeWMDP0HNOIRNKCrbiJp899Coxfsz
whwYvyWxznd6iAyHxxYb8RTT3lfxLjzNQHJhE+52zV5uwxPSt3R/dnOkDnctKVLNeoP6iQDVm/Bh
3IWtyTckn1OogsyrmZ+LnvFkefJpZ1fcO9mPLT22hh2CgjSeXJOqR5mQ2bjJ2UiQanm1EdpKvKzJ
11gIUgZts33zuRPRS+uwZsSgoPKsmtq3EnVvvX4C9rnEOA7MwJxBNiSdte5wF2SjYAfASUG1cZC8
8vEtR1925xm7zH/KzMd5KIpM9WCMiXWtHRVC2lWXAzedjyNKrfkpk32rtfY4omIuWe7gT1T6S31F
IKooQJdzezVmjRtijbck+kSi75h/fV/6SG+L6LIKaMfKUTI8dUo31wTz+021oCc1jZvCyhGrHPOD
G0sDi6vam3YzCADgCmQ4Jv1sW2G4H3ubGIz6gWbZhGQ1zPWhcHtF0KrbZOMrJBBqeouE4cwITvl0
VSp4V+4e3nqh/2lcH3NbZUK12TLup6MjaNDdpXjrwdhz0I5rY6C8Ivp0nkY7WN+VBK/w7v343mm8
iGIa6gLo9jSWYjgvdA4/ap8G/gPkyFx1HMb63UJ9wm5g1QfTJ6k/XEzqAmuPzJt2u/dvEfE4JZSp
UEdNIAO/lGmTVUh5szB65il7d1wBqGIqFpacXJu9ckTX71zirt9Er3Yh1Ygvlu0sTkFKsyT4+CEK
OSlgGlXqkKaa3jwNSUWR7oh20hdhfjpdtT1VT1dpur7mOj72fnqMDPgtMNBbE12HlFU3uldlG7y6
nR4MxhfA+Xonkb2oKvmRF+aMwIc1jqmCY75snEnHlFd4cB6ztcc97J+FjHsUvYFkYItmUUJ/LTnN
MILTF+6lQBBHQfG+6vtOlLQ//Tv4tOLWdHQtme70mApjnNbFscT11JAupavgD1XXdh8ofHQLQKU0
RGLJw60H3PI/8BFCnskQpWyf2Hk0KdFHKCoJ6xkYpe4WrKLiiF+2Zw0Hvva01aMc1sksFRwSpIah
C+kVFQHbmKsnUO9kObxuMS7dOc36Os8XvWOJsMT5bN+8gK740Aj6Hq/hmE4Jf7ZMENJJPXytfB3f
OcDwYKZMvHL9ZPL/aZZjuht0yk7rhIj9wnVH8dAeJ9UJEPOLkYCrKng/LIku6KQDADDSkIZ49YNq
2QBKnJx838A3hKvwl+tZW+FJqLazpgcmWO/E4lETxNa4ccs67+KXiaLPVazzCFe4LqLofX/0q1Yx
8aQo2JZMhgzpMAaqei9+c7pf0F44heyWf9JN5PxnCvk5ai7jHvBp0PPAh0CCFGcSp15KSH5ZXFwn
+WAscaB1hCIOSkI/OKY6yEInvh2pqnKoOKCG6XplIMCH8s8Nntjy5Ks8qARefsVpPOwveBq0eXLW
j/8LJNV591xe3DWUTGjOOV/zfKtUO+r6UVpul0Lg6GM3d5JHIoC2JW6dnD8R3GGgUXWXgk3JRaxU
GbN4I450wrevnuQjBO59AkUIsAhmMzN7PU+G9FS2v4ilM5aWuiKt7sgmzm0+OIHoDl4EHVUaU1xZ
hNiQk3JbvQ9b1x7ti1xXWIVmRdZ6lUlsT2Sflt67Kh400YjPAq7JwaPvVApQje/FO//+jBiCfcO3
XACXmMlJdPzsMQLEb+N8wxz7nTBAqSGYtf5pP/G6AefFhlj6mzV/i9JfrbGcwAQA8CUzLCoqXiGQ
LSSHeoFMCpOTin0ltBYdfpmiOEF3BXw5zkEabvCSWA+Qhy1RA4zh1MN4gIZKRdL+sHe2wo0Ks8w3
oZ3QURRYWWvl2ouc8k3eQJCvAa4i1eVZsyqkAalMlod27cdbKH7XHMjcXjJb222xkIw8tDsaxX1Z
TRH5XmCw1+18iBqNC9seJyNh+z/G5R4/kfy/Wb+3TpMykQj+WVYjwykc+YkeBXVhQ21TyjaCHsCD
4OB7rirUGzJKptiTfFg9a4vrS/NtADzY6xH+6VDx0SQUC3lwR/QgoypQVgz8AKyMZ+AvdUEQaQ3e
unGsZGBuZTvJFhBz4NJF/Gm9jsaIC0Q89JwpiQNbBQeK+JIadKj9YCTjMByA6Tltut96QiCus11J
xvnf6lkjkWhh0eZDf85zSo93zLHqxwK+AElwWpTnKpZJiD+MSxQN0I/ArfSKjajbTWCKbnKzulfY
p1spKE5CgsFBCEI6e41cqFCCjCbgQc62TcYZ7biETrCbtoy7wJmfp4puydVcxnI+4htORqWR2YLo
0jXs3K6wCEnavwUD59HqHiC1cVIPYATJP2Bb8oy2trgay/14lstG9wP/g9GXAGkSpPNnNSrE1vl9
eEn0ZzgF/avqql91leMImilTH9nFKltrq3oOezF8Qf00AMyBu3oZAAkcy7LFoDIzkM+wh6wl56M1
IdGPellvOCjd0DO9mcyRS1mT71MuD5Nc3Fq0gfzXN+zf8uRsca4TFp36Kl8LDYRtZYj03iTYSy6J
z9KXyCEESzP0JA/vk+ZZM3fBjuxUwaoawIaoOvc4Cq15sT7xAAl8evbNE/Yw678BqgIw3U0p40Dg
PvnvGeu7Gxj4WPGlUf/ZITngvlBHamS/N/95V4wHW24yrEBjahmZ6xq4dkKAH3VYa3hk5ROrcQKQ
pbwUOq4CbBS/br8DTRq4SgQYhbZRS9trmW9v+pi9QseZTBe4o+xcnJklQfLnYVaFPMiuMAAcG8VU
VbIgXQlUHKmkX5FcqHwEAfdgRLbbB4Z6sin7lzTSc0MJAtMwp/TWtWUp9hE4qMQElfIYkhLRElMg
ZXCibaBmBUiKZ+YST1NXtkFKyDpvpcKPE26cMNvVNNsNtaBtERBiovJ7yQHb7bLdOwtMR9TVyzbh
8r0yb5/YFigtrm3xeEfrOWuVXau3x0eCEYVMrDEOGzBmpoHxu5p2UQ7Iwn/LzLjh88/bMc6v4okg
i29FEQugHP36xIqf+ahTij5kRekCPDWmXWx0sHQBzUfIPrtbsldrYA4BmLW19ySFfAU+1J7u+/I9
dgSYR4SLAmD2LJ/fJM0dyat/xLJwxhRvERqaUEzua4wHTdvXcKO7OJ/uy+P13rSyoj7uikEug4Ee
vt49V6i9sQbo5kcbQRDXR/b0+AYX2U9KEjWVIWVorYLrJzTvkEuB3cbN9qBep1Hk4oXIaQrYKtnb
NaDq9JqIfb/P3rYOgojOgN7ypnFqe1bs1+D4N6W0z/DdKmLADuHSglKULOob8MSMiWoi+51E6EaX
cVt1COkRXRJWrXg5RWjvClxe8hxKZTWKLP749rWNVMeU3cumQgnaL6xWWb8luRRV5GZbc6ZJ6CEi
918F/OZGryyOyHpQFO+bavp1J0mku8abfA9sAFHo4mveHULFZ+E0y12S6YAwFla8XGf4YTvAwJFc
96FbXdn/+HhKEc+HC0oHKhuCumSNaH0JsMNdt0LoD9UP37Stt5cjT4CFoMS046BA7oEiINeB7sgU
M0i3jCNB4C55J1NWpRbNo0jUK4acfGF8rcHLpVaexN0EzU5t1e/YqDPVsjx9cy7Rc2qr5f5ENWjf
KUJsVF8L3HyiPdsAzdj57nz+FyAtEC8UjVZcZZCyHKNB1IUgVhbH9PPJsemMGlL0z5GG4Ej0jcA3
h0LQsu0hfqnV8ctTWPZRpzOi1mH+h82yJ+X4zxwGglNB2ub7Skg1ss4g7BrjE6EfXpsYpzwi8xXD
nwpKxggrIOq6DVYv3JlwtziBPShn7Z58MO9GEDOPDMtlHraMaSgtiMOuL6fYojUMsqde39QahX3D
kCZEocW+3+LqFwaL1jFIHRH8DQc8jUSABeZnALC7XKvGYxdSgMLwBQEzY3IDaljJLhVS1OMrhHmo
JamZ28LzoxDKItIW4JalLFMm8kSVMqzlP6xrMbIMTeWdBc/imEHZgk0khMqyTNPrg9Rfb2AnnjYQ
+fOtWCay/C4Osir4brf6pjLhrjqdW1bFacLh8AObDPpFA9udrQpK4LcMHZ4nuJ7eqJRG0+QK92KB
jN52QBRSKwTVffRWdo9ZxTEvZR44MDx8IadptcEht3QAIVZiNPbynSKynZwk54r0W6mf7SZpwJxh
KzloN5k89ldOrFO2jDBCuPSLZER5dA2PRZsIH3ivnCqZNiTGw17IGvMus673hXCjoNkfPH2mEHqj
qDvAlqQujF56YqXo5ABZm9YHbG5dSJkXH30fgbSXURjcS7dR1H/n7GD2e2Q5/tmw4YJVmeseCIDN
ZfSOz4RFxFgI/9BEL8Hc5hhj9Saol6b39Y1mcCZqgyUUCkxaIUBOMwT85oRtxUYHWpov4kCOcDN6
peXkiaXY5QI+6BA1gCbmugZiXMUdG6N/LPpBeSmGnw7NffU2wn4S0X7D81irsFR7ND7iNh2bXuIr
coDyEE44d4kEWmFRz5Y5rBURPqAJ7W/wrYJa2FOO0IFRImE5yNVbbOdH98qCrGlhZvC8iZHGvi9P
YnjjDYt89EtuWYdnrZbsYUY6qPOwKyUg2ATC/oz86gwD2waYVsO9bQ0uUUbpwEpV7Vzu0gCk3VEk
9kqgG8dnFVwZ8IvVSCPnIVA6ow2YQJJFeOfoUa/vMLCigGFIfDeD9fpPh+sR3rxwSR7WGbe7KjRA
9hY01JaF1ocCUb+FRNL9/GXZPWMEoEDr5s+anBjCwjmcvP1r8kLbpLFMdnir47ahNIhz/tLNgWEW
Ggz4/lZlA+tcqCy1d4DyHVRdcXNKSMuLz/U61pK2Q0TYTNSU4hWMnxz97FFdjh3CyqgOnxorYnsd
kZA/DHvOTtM5+BkEtF3F0XIUgTvHyieStL6sXlO7B5DRSuURN4iTWpn3d3m5fjpZ3NTyyw34Kd+M
0qtR1kVZf5hY+J6z4YBeYyZdfoJ4o6vtP3Zh32YI51OGBAR2Aj0ICa/cUk95UEwj5JwedqN1xSFq
gtlYUaBBTUsL4FDnLFw1E7jkIERlTo/N7rR72uYNngOotQLclG4xPrsQ7fTba0XAVBCfBdQXYfpK
2/tGE2jgpPAblF3JZszrWMVVJBvihYg6MYuRW01qK8Et/cZjRDl3wMYxSUxsCdEmL0oznCCx1DE3
Rvo1dq0QOTHWrcIAGOw/an6Zlvin36v2inBc8KHQvunuyz6yUKxU5dsgcxyhtZWKL48GbW4rKuPE
WR7ZYDL4bzKSdU/80hs/Py0LN1dae29G3D4BPtlGCWEuRaZvydCwtcVnQXenyJtw1Te6EMuB+eWi
iVN22eCyXdFW8ckwQYCsdbLvWgh/rR+ZOANflWlXBBX38Sv4RrDnWFXN3Vkr53i7v5OfFq2rO+eP
WLijWXTISYc/nfmxIj1OznUkOkTAZiDPeNHC+iZOJoJO1+LGukCBrHlxL8/PTIEsUtcikO57CzfS
Gb4GRXgmlz+UNEQUzLRWtSDgGr8Ma5tySRl4R4Hdl1ohJgrghC5dCh44OlMVfQmTgIXSPiE5LrIT
WnjjJJ11jLGZdlIiPXRMMShtNE4bTz2aDWEW7c1ywjK3c0Ih12bohfU9qmvp4FQp5DVo6CoLsoEi
YTSlTRyud6fQuMp17SUl5bds085VAWKeJ1ABxGpSeDIpr0dZfVMTzzuWsr9OvuybmSS6AB6gNZa+
yMpWALLFNv8axmIxTAqjmw6fmXBNuFSaAwWKx3wK1UB/aIqKkdc16xkRia1scBQvVFuc+55I9UOG
EAfvA0zYtrYWnOFZx38ahpjuBp/wmIo3jKmjFmyVAUZ9AN9BDD8Fg7UKhdxDzOIK76RqtiICk3oQ
dQfhjTIGSDG3zv2+uL5rch+dq+5nO73d2O0dRHFOsk7O986DqWJN+sjrKzeaMJThAtT3w5U7+e/o
XC/Vc9177EMtopMjLNzxxWznomLKF5kP2yeNcRh0SkvOV1fB/yp8d2rupN/LaJfm8vo23Z2gMfkX
2XFFuE6XO93+dNfsbHep0q0wPJTj2gDDRMyGTr6HUVBVxD2fUC6CmzYB0YfDBC/iZ7p1QgX46rCs
ItFrLBYmVsW0pFAb0/Y/USa2WmEXH0DIbSrhZD2nI4j88Xju5A1EamLTu8WxSW5OGFo83S5A5Euq
SbbpVipXyNqOfGr56NTWY8TiLpm9n8fe73RvutZYwwtFO3kqZNH1fb4RTfs8EukQx+9R+KW1nIPI
oFls5GKGw5WuGIwx5FsgIWmSrJZBfD45f2vIOQUpo+YBuArozrrS86FWbAcWOSmiiiTGRKoMb6Ni
lI30PS2KyJAsz5iCc6hKe5A8AEHZGS97628Cckg9oMv+8M0zP0rN13o/c5E6k/wsdWvIcdho2OYW
MB71JOp4Qa9l4dJgGACL+XK2gX63F96I9STVDiNpOGdEjUwsgXaR1tepWWQbAXCDDLAVS/YtI5OF
b57D24ph/nYnnJFklN/BSjyXgYHf8M5Z3BZ9q5dNDApVPQCtSd9X2BvWCKbE3nuEDmwDC3aIWRHI
lqCuyORYXJR+czGUFUWddmIFIgYYm5Y90UMsHq8QMLGlN5T9LNE58o1rQzC4sYvCp2wWe4Fe3D5C
//e4CNUCScEfVMI4ZpUk9iUSDVwRje14tFWDo7iKsML9STlmGYnpi8d/ybqZe5tSCUdzLkDYE10L
zycfn51RbTLCWEPTEOi8cr/LUHXEXR1XaSEJYhTDio+ww7wN81kqToBITfe5SVWOfRWGp7YkS2gC
0egPTTCb0PtwF/Z6Y8bXM53tb6v6bUKeatw2XN8z3lGRbSMotNCopiKNMyt2xuKDRSW0uWsDSCmc
7BGckAxPUekki5UPxZydGDPQN2VXFtookpcto0Hx0D3MWaXYUqsjFpvVEHLvLhUZVusAq/khPno/
M9BPAq8No6Xz8LRGkN9A3Doetigm7Z4B92sh8ZKNe4huOs2wgR9w6tnAuIfRUhQPyFS5nDc1DFtc
IMnfKyrJRqx6Nb/2u4a1Gpuxvv7vntTE2pHpmmeNA+1vz2M5Zk4KjUXmc00TRAcFDtZWdVQlFL8I
wpdZc6IEOJe4F1dyuqzYIqvmfKue3cdhVLuKta/fEECdM/qoCloMG3oE2AqLgqpHGD/+ay4l1PmY
22GzUFCiEiOhkJrPzCgKtiy2uP4Vqyerw0qsNLSLDlepUO/WD5wFQH0r9APzsmSgb0mK/EMxa1IP
JeZoF4kJICEiOih+qFqyERGAzNIYry5u5+SsE9NHduU7DJ+3c4+G0ZCuXcc8atfXFHCd9BvaFCk8
PAF3QRej5z2PLWDlOESektX/dqnn3/qNQtnoA7Onj5DGkK8zcbyvf81M2iAMRJgUMmzr11LTguQI
bMZjPyF0wz3SgriV7CWQg56/oojEIfwkHPLjrHZoNxl/8Zb2NrZhUYpFEWLw/VlYGouLkqYY57wi
ixCar+uJG4CvGIEBUb61erbvMCyQiDnACd8oiiKvj84tBWbfIMtiytFGPvUY1JxlzhZ8nIuVW9v2
TrPfuvQWlxGrBgDwthtiKN873A2+s/7l3dSM1/es19WeWmcN3DM8cochxBDSsKRMYd2mPHSUzTFi
UkCpiTiJi9hrs2uTlt1WcejtXHfQsXFghNnk8zKYze/6BMdMR04ojNaDPedjkycD4iGXpqDu1Zua
3yBxkDlEtLRJEqugTPHdlQvVEb3VnNzP2F7y/veZC0oTmROujNWra2kkdGGe6/mMG5shqGNtSdRM
cYtGFjOYV170tLBEx5gg3TI654CA2ELeUJ1KtwQJBG9JmpkoLoo9Ff0SsudsT1yleSNNyq26vasF
C4waeVlKbmkacDtibTqlre4n3qZdpK+EfGgE0Dtl2bJEqJP3ZVBZAuwX4DhaxiDvE3tLTZsvBCof
kaf4zIr73YQB1u2z9N/uhA0QN7VZszGb8ylO8epi9bebDsK37UTRo0BVcOYZcT7DzoNAXaOwiMcg
96fZ3/0NuHXnNTBN8UKmtfoOG8Gwup413hx0E9juiSgcuy9ZSF5W2y0lzHoO8LTkvxiZb5bflWIZ
WFoJtsEd84+SruUYJlycyhd85f9q32d6LdcREL8GZR0+avBKMnVgZNGokH62KWgdtyl8LJZei8LP
UgJJMjzC2RdJdpR312jcc17M10sljIhW366ZsfpL7l1+Gfk6w423rL+rL/xYnlSwe8Dmh8cw5q0Z
flMyc3XsQvfgg3BEZs5GI5eIyGJSsxt/bhZGN3XaN2CmDRkalbggjCUfncXpIMPYd4Q8iwif2OL7
aiEQf7B/7nGldPGAdkhJYrg2IgH9Tt3xCd8jDYWx2iVdoymzVoTvqpeuwv1KrHkel4RcWsPYbKaX
WBpo3c0VEU0zrFI7nHEG0tIGwp7M6kRbHHOU1gnt0OjT0veUz0oZqJP5/LC1G4OWh2FKc+GKiV1p
kOF7SxhN62yW3qScDSVUZWT7hfrzEHehGNXUUKs3xWYUMYhkKXIu1C36FqbApxBY5uN3jE0BKurN
ply6YkL7h1QuMLh6lW9Ts7cXzodRrz2Ra/rjGSw6A72LyIVc9qqtA+QW1p0PT1Lyq4nwzslqfUpm
Qx5CCWBPpQuSl9QBTKWQle5XGQCzMhvwdwwM7BYHcvoo2x4xTC27XrS1wvHznbID4Bvu8rJ/MOGy
tiHNwj8hAYfA4dl3gVRKnBaoNJUDUPDVoin4ZY7CikD7TJPeAYDjuzq/F+xj69eY6k1YFaKeo7iP
/BFAzYEzKSSjaduNtK7YoZQwh9pcvAFu/bI4NVYnai0twtDJ1h8YQwbAL3Ar7DKIERNV9Orl32Vq
MXnioVtnp5xFhI4Ze7aEI8XSG4yotz4yU64mJCUg+38WkvIdOo4giM2aMjeLRoOjCCjlujkU5kdE
M6/4HZtmaE9HurnDz16k77h/ccC9+ZZDCKXE1+f/+YtbpB24+8yXdW1N3tptmDRg/Nh51vXDyDyI
ElVafZCJYfsKmS6d6zMpbfK2kNzD6mhTFzRcpLSM2IlEzoc6ACzNXbatdAanljxl9tnQxHNKmB3K
wvtdwQb6C9q080cd216HOZ61LLA6EYRlD1+ArRQ4WYqWTiT/XOlgCmhrIuPMRZqc64kbrL6xNgsG
UY53Zex/UbAzNHtKFtwdLKsBsyo6RRKOJlfVLLuRZg0M8aj5EJ9xA1lgmTGbiJr6QooGUrasUIdt
neblyOF1igWpr9P6cY0XBE3/iDQGrcPE/eudOCBcw4kGCT6AvxlX58x/Yniz2PJ5Q2y+iGlxMuXT
qEWXcKZlhLVsXEg0XMHoTsw+HyK0q0ouHorxyvGO9JXTEngkB1UPqreUc/f4+5GDQT2XiOaSuQXH
f+3RlMMOQq0RpnUSq50E154Crh3FbXZtMuqBDki3fFhs3ESgrVTlcXVswFpySCeP7wnwMVdzSNzW
cGGMB6W61JVqv4/F7KO+6oLYY+CRSpveXm7Q4NweTdYk8e7MwePTFBTWKwlYdOW5Jkgr+RMomzfA
Jw3rX62xupGaeAXI27+QXnsJo6pIiD+enlac1uRPIRH4+yVuqXfnfy774okrblqENuCc5dCridsp
R/QpXTjXZm8RK5860nPX3AcDoPCfKZqdwCTV2wKHZjIYZEuuEeoirt78C7LX5lplrjGDm1cS/h/y
dHaI7QJMHlRtC0EmaoR7fix9kzzW9PMPcyfKsL1L2TmLLgynPbHiCjjR4HWhHrjwj9RsWnGvCXBn
NeQqIA1hMBuImFVlrhJZonFC3ps5f/utKqjF2t9UXm844a4LgfR7wTwNNX2OB+yP8JwtdOPUWHYi
wTAINTh3Nh7EZBPd1SJqy17UbGDObtLQtYTY9PHsufL0RZ/Z7NTajQxHqyI2kvDebbSDjQ/bjfVr
qzbseO0b5l9dLgqIH5nUsyWIOfPHP2s1oWrZ5yJTpr40f4clftwQzG/OR3iuHxpkj+B1kCkLvVrc
mzWqM6NZQE9RwbfVDrGyNQXiJeMz1xsz44HfvoLM51TUuRmZq9Xxu2XyUOk+BnPRjZ22Ste9DWcj
jcIZtk+cf9F0O2uJ6MXsw3abib6QOgCDZ63cBUTwcihsfXUatsSpReKZY350Ix2i68FVqCfKVrpV
xdOVhdLHNrlKPnVXUp5T+8IPXd92w8kOjSvhUcJ0O13u76MD2HZhgkolBqR5Af1oB16A8zF48mQz
QGmhcx1diNw1WwekItEUJO0GJNay38FbJFeucY+bdOueI0P1Ax43RwjJ49T+O09VGKMgIfIJT0nP
IeSF8bgKMUU2DuFE6RvKHSEpaLy01PbtuZilnP2bSPTXqXrsP8X4LnDb/Xyyl95AAOQlRyhYV4+p
ifQxTaZOnG4j3m92bH8tqdfi5b3rLLZ3ulftsA7AlGuaLJrSX+LYnKMtM1ETjK3HZAw6ogC5c+qn
Wi+S+COsGZ+g8tLH/JcagpkjOjn6MjXRxU97yrVk5uQicqGWudOmWr9BcRaH3TMEaYcY8KQ6l5Gl
ERBDCZyfXIqQLkqOeJJ1Pkn8Y9h5upMGNkK9v2rBQZ4IvwJb5Amb7xMSbVxexuPkyT9Ifsr8yAhj
Fe9DluItsuIvLQQbhV6FQItpyjlnmTlswqLHKcOIOvYv1Kqoveh/M+J3QtDxkv8Iu0Zt4Tqh4QLb
1R66V7V+mQcvtZeXKWtLBY9EFXWpB5PPPCuaUJbdUjLl05k75F5zC+3rNheg8+Y8MX6WHYAU2OwO
A8rqeGTDmQd7PJkwY55D/SU8nYtP+2gTfhaIhNpfn/9WQvekUngnE5dsmrUoMDN8Jun/PIiEVfrq
IjDOiuy3xfxOnNQhR7zjNyeScoC5Jiw9TMoGmZN4M0tZn/IQc/QBUHpSevCJVTcGLuGa5M9OeMg3
eHB1nL+oIPBmipnKMvlJFnUPfym6OyGrVFwYdClyg8VLMEhP5oGThfW3jXyfKMEZsJzXt+VxnUOJ
AEmK+PKPIs6q6HvtA2cMxxoqxc2mhIL3KQqenA2JDiiET9EXZ/c1K240Dm4PuprIYb75kyA+Sxfo
fHVMcd+0PKrm8qkL71tnaUteJDpj0F97dXcwVJtuSl80dbhgWgG3JdexJPVPSe1CW6LB4Pe2LT3d
Mf/7ygq/HSLLCCnMEl0Y0lvKPEY4FmPcQW2DhYjwrIZ3kRb3sgbJfPCuGvkoTyM+V+gCtwNMDoXU
Q2XdGND0Yx9k46Y3C8jNROJ8FQpVPfZ7GUwL6+t0ViM3gHbJUVO8Xk/CemVi8t5opQZPbqWKVEiX
muJ419cZHKTrlDWBq0gAkv3zQf73vL+fzHwXCBKYlvLIVziyKpySW2plm+8PDYGFT2Wz0tHXiu1P
XTHz5b4z8lOfjPiFwKxLStg3U2ZWgOGLKW7HzU0ym28rEcOWH3CiulPvgdeS1U5vthXbWbBxSOrQ
vnbyghXxPXF4KVpPIGimX9xIud4d+3XvSejtr6f5evqxIwAT7SQpTSyjI2AiH8PZLXlsuz1G3pf6
dS22cV8B0yWYPy+D1xGvsIximMfHR8rgFyBSrSPvHF0ywcYGYa0wvwf+/zK0XlduRdhk2aR9+AzB
HnHl+fouoeX9bvMENySTOTyRDLohemTrbM5kxkinsZMZoqt7Rm8d1Wcqk10dxUvHB/VMmfYF2OLI
Hw4MQcGN9tG5K94R8TllvXROKGX1KqQER+uf9QTX7fPNtDVBqtg8V4uQDZgzAOMHO7trA2JaPNvn
f5dXjEVa6Nyd1e/Tn0kOPDnWx7Dqcwhz71tjFimog0CvTFYJhKVzfkEhOlA3KiWexlA+R/YqM61O
bbqRhJHZ4Ouf78WwDZrJQTf0FRDbOvNcArJ+SKbI2buip2PVN+XGs562pWFfoMVp20j0HQ7TxbW4
XZv9gPz7qCfPiRqEIEaSjFs4P/pF6hKH9pofyGXhdZcg4wbKwaPMetPb+7vmMnxuAaOAMj325Lt6
8gFiKXwujNBuaRPloMCkbcTmtKR6J0sczE0QdilQJlQS2ule4zh1M29V82HaWWz0AxAsCHXX+ymL
IY+b3eHrjORkhYX5bnRS48DqvIbfXcQJzt0aNRnnEzoVEGH0H3/9tz91wR/CqEUeJJARoy2+Cl4V
YKf7M6VO1AcgXp5/OKvTVWjJSptVG5XEfPOexZI+S0clSEFVrv+qrzfJA7GrTm5FyKgzjjuverBz
oDdKnHLc5IRMiZvBf+gjHy+2AsB97PmIlII5WTe/ZzJWsIN1dX0j4YtOLd3oS4vsggrlkGCVwsLH
FS/8lIplsChS0pgqyDKUeaS5lYqS6Hz9xrgYJqFI3bnjjzvzArHD4XrCG8C7GplBa1a6lxTg8oNg
E0GVaKNIif8oc0JnoUFK3P3FaJ9+ZEsv4u2x1EwH28kZcrQ3RQ7n+p+rAocSmbo/rLhbqJ+itLLo
aVe+XyX3DFzrgsEeDUDsoyoHcfGnsEyG6d4l55HSBXeF1l7jMbN68zK8YsGWHFiwUQ9D4ifT6fBr
aOFZzWtLLxMKzMKvLiWmeVLzl6yupSgFzyZzyZPboyqy2jvKhb+5rGjqLUn/JjkVSnlGKdspcMvk
htS/+uZwCoLD0FrCwUSnP5wkJ+XtjJX/Bnn0mzCG8O8snglQm/KqOKICHdHVMCfr4em4DAjM/5nO
GK+Ps1y9FzHAzfKfw1j08HaVqSw9zbF83fIlcqyCtWisdVTISQ0ujq6q4dDTYiCLELD6cOlW8jpK
AqxcxaP4+GgKhnKDuIKMPfgWFX32zwjLbxFoBn7acQV1HtdS8M6cBEMfAjh4emN4l0rfEnpSOtxG
DlhH2zwadi1EqoAFkc+W71DKQHe8WpkC0PITkT1wkxTakvWxMQeHH3UoSEb0PnaFTxR+/G7sB+Ck
pnVZQ7qr53plkT4u+niXyyTL2K2g/3YB8XDpoXtpWKjcUvXbCSwmA2t6JAHuzHY1/GW02vQmgJZc
8gJdSrhBXMxn/O3Q8ig9i02NA+bbrKuGwCVRYDpmBzu+iGQ67zrpImzcmZEzEmJ/SzI/kA7WhYdT
PFRRtReSfMEVdtgjVUh35NMr7C6ItwrBCZEWU98nPIChkL1O6Ssih9cuZnYpBZRyCY+5gXFXlgOC
nDIZuR1r30xvmaa8A04K8QESvaNphxYpx8Qu/pnzrjEww4mLxI+qAyTgYuQwePJrL5Mrou9PfNjV
2iCfaBL/1wvVmfeTOPQ8Hp7fC26/0+vGPh65lnFMDt70E2IsTWXJLXqZwJ+OogC+hjHkLUKRR2ib
LRQn86aB/zCCWoVbrCDZy+GmtS2f9oi3nKWnti6cCioBQ9MfNhOhbJVTSxIyJ0M18Hd6PEIcojej
oerbGkVr7eREHPofHu9Wx00AUJQ4IHnGQZRWT/jMluyBTvX+bthslLQuSKJwGN6jgLHNrM5WLDrS
hBBx6cUqsbIRcqck+FNFPHDuGnXwyuFz71MjWLMApppMCXBq6JApoAekW9vePo3BQirgOxH8DUSr
1rJfBOD6SxSY13FfUpvOQzTY10rw5kN5WrJIF72LXmPwu2/pMmv0vZfRiH4my3bEk1FGhfgKaL+u
M8XfvBQVVY9lAkwMvPIBtj/qntpjuqVU3H8EbFbxg86dEWDQBmC70uml+pD0kABeDR1R7g6GIOnf
FUWagiZmsk6SZNA29ovB0zTXX/ZY9h9W3d2hTEZgKbLNEUaOYt64+89477fIvSsxgapfIz4O1Mug
eDlkIzkDBlsLkZg3EKITFQbNwhcXX/p953EYI5RULhEZwZVlUUgjs7UIxqURLHnXLzacYeHH9QbP
BYCF92geZ5UzHKqi2Dey5D3d1xAQWp/YL691PAfL5064RF7huLjxRJklgq/Gjmk6ZgniiK+6axDX
cDPaTCV5AxQPpzj02C2l4vjP2XguYHH+b8SIXfxQzWabeVNwunvDTNWFsAIYiuKduNb+WLTp+v17
WEJTyjU0bQBUYx/bADZLzpzvID10cv5E1kwaaBa4aM3xueSr+NnzaT2lesErWrmNd99D9YThYlZF
HDNiXGaBamiApYtQPbSeDO9Rod/ZgQRNq2FYR2XOBPqephrzrjCs1zOoOVgxcu6X9zTm+/2iaco4
FxfNB2AfleK6QIZ5Fw7dhkVyelFoNlI/pGiTOeFWMrZq/9UIb8Q/jRS/hDKsqxpZqLyvb+AdzWIZ
YDO87bwvF6blMDHHYAU8pCJVIAq9VUQEdXuPnN0TuEGlMG7bJZGMtvkqXA4bQ39tfwKUrMSdGRtk
Lvo0CoxUKd2PniGikQuUjQaj+r+vb9mQPWLIqgq6XfJpAREwWfLY7+AInp4ujPUIB4K4NBc+TAFI
+r/NzVj8HbaNf820qQhS1nYV256cIUloh9WYmlAdVHgBe5bTlUFdVR5FQJLnXFbngFdAbTPtU1fP
sHh/bnUEvT0oJupno+pbG2fJy3gIbyylRJ2vjB5ctEV7ZhA5AhR1OoON+k4R1GegL8qGMk4sa5PI
yLa7yaqiHfd33YamBGn0ETHDKMPoZY+xY1KeVU+0Ck7fisWFl4IwhTxTRD7V3DinWY/nUXnbbinK
I8qHbM2GAdOxfVcF1Z1DVj2oL151QUippyFODqOZWl8Kf5cPsCsvqllXvQ3rc1eJNt7v6NEBDoTX
WDtVw9iYMnyR1A3/vQfsMw29oU/0NINykUWJHUHXY0iNKVGfVgiftva4KtTUc3DY0ipyiA5nbnUu
1rtlvzPAbcRQeQNK06fh4+nQrpOLwrgVgfypBL5k/05SFhfjivI4M+xkKmUar1G4lFRy/KyWEbGk
GEwNxbLYiCWL0BWrrB1n3T1dHMfhwGtxGDvtm2fLtofqEvIiohIxMKwwldXJEU0VYefAUWOpHckU
1/77Ho1+J1lywF/HOc5w4QAtxbi8QwAwCGfEpXCtMrm80msiXlccL7zRxMwcjJogeV74846GwZHH
d1vznRmPOjJdNrlG8OnIsdvqohHB4hyBdWhSIPGitDUxxs6l50Hhef/K+Y6Qqo9ATasLWo5hpiZc
iYpYsJqGaUKvagv0VbVXkQzWJ4pr3c/x53kHgGtc+IsdvKo8IKicd+CM4B5jlokoS4bhw2HLZ6cU
FODzTrKE87Lae87MqRIj/yEQ2BuVBd8i5uwyqvakmi+NSBN25JRagPLm4aGbd2EqZuHne0FgeIcc
ysWs3MYGCfo21nzVj7cOJZewurlrr0++JvfMpPPqAdB3nGBu31gBffeYazfbo8bU1L6Ax9LCMlZd
YSGVKpbl2GamZSvidE/3Tq+dV8agfHJsTMXwU17lqAiaPXrz7T0sCr2cbsCZl5a3x0mPZcdY8DBh
5rJYVTMHfyRydP0YUuh7WF94PUIk7mwLNVcgH3LEBHaqm/KOjaA8slBveHHFuQgmEugZ8ham3Opr
SMd0VdiJuJIzvR+aSp3LwZ3Dml9bEAP0dokNatkfiZUiuvDrkNkjA8adrUOYrsjEXDRXRr2o08Ay
BrTtI/EuftbtlPMsL3uiW78gdNH+sNt5KBZgsupPkLpLPFRZCYtNZSFZdFC/NYmwXmMEcetyLOo5
NhFlzHZQpWiJXyItoEkbAxUZQTGK9vJ6wg04QvCIhDdaDfXeTHcITfsVNdQwCW1fccfU2anSsHFm
ZHw7rTfc1U2BUXikeegRsIdY2gbRiLSoyVmTVE5JlHApFuNZEQfeJq9vI4HKOJPs6DIQTEhqO7nb
XSJ2RzFXKxqEdvxoMfnfsoQ8onR02gbrgU8Z2N2drseULZEQPxuijhVXwyHtw25u225jNXNeZ48v
iq8e77EYAD6Dh9Feno6y0OrH52c+Y407ns6hhLNJ8/zegVjrFkHl/+0DyFUEmZL+47YtyFaKR48x
2ijSW4SXlRTPDzCkCRyLsk45t76ja8G0Wv4k5+m+OSZ+54P1tEV8CpfqYQUvF7qxl4YVYQXjJjHd
8+n9jAXWvb3fMRpS+NSlce2f2s40j1SbuzlEz1kkcRqv9GD1ueYXb6b0MwTu6EtSDfSVrURqrK6m
fm4EaNtCVnue2W8K6psSaj4qPnxYASg3TbY7XdcjoWsmvgnqbr2vu1lWZdN0eITyTINN/P6hHAC3
S9flMD2ngM3UOWRbbZVF1rIkE5Aqad+YZcjX66Q/rQbg8c5VD/oxPy9if7xfpMg/NuLoU0t9giJZ
M7AZDYRF82yRazH4EC0SyQNAm5j6AEgvgtHMKE5S5Azw8wrOlThXeymwPKApRCGFna9HsZnpPXnE
aBj5703kcJBj2MaYF15MWbul2yYpW5iTUMaUmvL62vabpPI1BI+yb016gukYkeoF0gAMq0rVQZUM
rf8x/yWY5Bwjz9uqTlbG2XNpHNvFRWuIk2KjsKi73TQmI0etM8HUKve9uq799Ft57YFF513JNs2s
L/MSRdU5vRj+bQVdgQf0GX/y/hfEoM+MuV6Lc/GkCzVjl2fw6sNYLi9arA1Pha3+NGRniDIVD11e
E3Vc2a46I5i81lcDUdnI77DuCmOsZOvTXXEJXzxqMY17nMwAOgL6Bh9710EE1n8HUmGNzlgwIs9/
RqWk4k2jZIZNHgUWqL3bKCh+QkrXR51RgDzLTx7LvjrKgfiuWEX/1BHERDyjOIa0fbN8BKFGHPxk
hdSVqBHe1Lfmcv6tR27IVn7R4u8H1VxQ6pAGuO1eVueVtO6e8Nm64ou38mnWbGsMUMiSCWeqhkkP
kXQftfs0dSoELXxDiSAM0zBeL4wzwHMIduOD+yLZbKylUetlpHpK8q350dUVYu7FI9Q9xSaXK3ua
e6rbkJ5oBJa6loSl9rvGhuE567yYrRtXsPhQkvhcVv57OwAIBL4jkJqz+xxP/SV3UKZTR5xnhwU3
he35jNlqHXBNFFmat0aizK1/qmQAv86tCBhVZ7MWQbEGAIqVPqYg0yMmEStIfqan0n6ARIyY5xSp
deZNhIRRsEbcsanUwiBgMhOGak4v5aJd0ZxIFrlfeK7ecIp3Gxcrod+AndYNAzRu2MvEzcRFkrBh
jWACwXNO8o8ZnhX2AKxAuR2hsvRPdIdI6kNIzYiQXWdhj4chHuYOokvfTLdHD/WJq00FREFepzmQ
4a3uHogDsIHgEuwGGCE5hcSDoE+VN6MaE1VdKDUJYn3NAwHxrm9bsqNWxLVsxkZZRlbFqQqzNPvF
TLwQuL6xM/IaFrhWqG1uHJN22Z/Ptkz7GFf/rYfTNmhy9gsdJe7xHoPybr2W2l18gML6qq9g//Ys
vK8QR9v6ujHe2yJ2FEyPjNtyx+i19I9cDlZM1mBlSVu/2E322ClssbIAJcpK0frQJVZrjP/J/TBN
rUBU4QtoRV/1A26twhcEsb24uCRpam/Bvons+y7+aIWTNKjfhrZWJLgcEpceIwAndsGn99CoJD1w
H6sdQIdmnTobZHM+UpDgYbrHOFt6/PIpdOsiqsjbIbJsYGQdPCZ+qLAlZzO723xK/L2DgAcg8lgk
6w5E8jgCEdU1WDu3WPd/XRzMqXjpvtuyiQxIfB2AgNEUXJsb8U8Dfo+2OWYKZjTlQoKWawSPI+5I
YTytTCmjHye5lJT7/+uNMgI+93KZSWTXwYw9TLPmdmCFo/hRKY53ua0mgh4tc9VxeO7IJxI2346U
wVqeWExtr5DpRRjYIVPhdiKUHreQ5VfIt+3wfLsWxKKRJZuMrd+DKrpVqOFz3eBqQ5VvAU1IUkMf
DkbfVsqAoO8zwzE9quw/aRrt5mNodUeJ9b0vplzWemnW/M3PtWF9v1RMXESTmaQvOSYhCm7VD0O+
HNAdmZOPRXn2lc+7AAm8NYsRx3fbFDNhkD+dzX1aLhMhVPGH1wHo8PRtIwmM6HD+wGUEx4I/bNRM
x1vw/NBg3db8XSQSFgDf4srSptsXwX7vjRS7vY7/e0M4+yQ9GNy+rS685TDfrYXlV+iXMzzOw07F
CUXkre+sLm5Q4OPt7S/gQ+caFtMh8Cti7dXahn4gzy6mqgM9Rcgp7ZLDZ+9PrE0QT/+BgYrV1tk+
v/COVhtRAfwAltcvU0LCR9G4SksHhoowSNDMGUHQRcl+DZ1mir9AMSzjYFLrBpnHsVXc29/Iqsfk
ll6i00fa3cU2pCNHlNFlhy7bGUt9xFmcziskezzPZcuiHvqVNgsr4ewnZNGudTAyTQ1RYlABl1/8
VVo5FGavBa6MyWpk2JpPXslekeBr7s6Ip23SgdsXRkHlWRa2kKK0vOWT2K2luC+Ae89ruqpX/kg6
FoyGZ8S7+kgBnMgE0h9ti5rH/F9T/EseOTgYQtb7e1FULI/wrpWGy9M72s76EXivSjYRgLjyMupO
++PIYHffVRhm7w/GMN+loyZxmJYRFKu/L50MF/lHHDdJxiQF+SXazsTFCl1c79wEznyzkx2rAPE0
lMjKJbu+vLETJK9a63eCdfYFy0ljRkQse8sT+nwhNXHQ31XP2OxwXqNQa4P9hARODR5dTsCc4NYa
BQE9N9zirNHpd/J9cfS4TsU8+12qUpDnQ6XLHZRhGWvglzuPWCR+usrMeqx+ecdaSqv2MT1VOzKk
gmQEEU8LPAqPCWb9dXimDmygGTLBNxdMcWrpcSRP92b/7wHJq7CSVSWluSCStkfK76k08QSRaHXT
n+332y+o/PFD785glCT4yd/2GBcnKgUGW7T4YSUOXCoRwi5rrnUmmFecnUzPNV0sQHfEziwsrUwY
kiCzr5FNJXv/SAwGwRbcw15/fSTJCql3V+2ydBP21f94PdVQ/KjuYLkWshhQiAfpNcEW7rtDkDzW
cvTyd9YTRtIU1Y9QijZihFD9u2mSdO9xiJjpwuOvoya/DxG5vM7GZX7agPL2GgnApcgNp4NleEWP
YX+pcETrLqdvXXAF6N2jH2PyG6QyiRb/PWKRHOqwtiC/4gPl82uAK2nrOQJHLkFeUHNgyp7ZCc4l
aWmteoZDbtEWE9+APgVk9jyujb+BOrf6yTlJcIymC6+Ln4MKISeZjgLK8UNmfbCZZG8SonyoNeZD
DJYrF8hD08UjXn7quiTGO+sacJslCNOeu8s+5V6a1n6Q1sUp5C4AZsJ75s79wNOEeK2suCUil41c
z7jQBw8grwQzsWiYs2KJU3NGGw2IRR62oKXH2NSoJBIhmvB3ivGXAY2TYGXsJEla7HTAcYKt303i
Z8Q8Eb2rkd6K/zyaODUfl5ebE/GnBgcHpXZ5SHi5LCxHEGL508vlzS5salnQrmso6EoQACiKccn2
lXPBx10x8FS0MnHPT1yVejmoeGRBZzjmbTDuxxQ7LGZii7IRfM4aYmxxJOvxQXsVgh5EegMKgDVb
qIvk+ko6w8mYbUNdk8RuJBKwnYWFlHoYW8Um8fsu5eVJx7utI6dtVsOg7+RL86Ri4NOOBe290rmp
BIqxqIZ6dPYLUNvdbFMldxfKeWiHDA4yusSf00scyBHCaOEK2eA+sMZgwyAMCb73JkLCeUNjYBMH
U374POIL/V4p+8ZWiz4DsPHs66qvcmrK5DIYQ5rfhci1+HueyVs/ntrlzemgRFBJsBiWl1zWFq/3
QwjIwB0Ko0OEHTwXZcCl7rgmCCeGBZdXC9d/jbzTLifMJHebg5IMNxu5lmY/RnAWkCKVsrbAzUST
zxNMAs9Vs8+k3vcRr0cfkounR7KNEUL7oE8UmmYDQy+9odGYbVVgCEoA5zoNdXsSMwDkmZjOVsho
p2EoQwfKfQbSK3vgElsW7KsUg/g3UU4mDynozjPjzdpRY6oxQz8t8NvhCyJvRuLkSgNqsr+3xWl5
64FJ6hifPyshrqxAZKpaguXNGxPT7zYCguO8oRvV8neXSzzyy5ecUmUpk5iMj8qdzwlCv5tjtfQ6
M6FQWciOYs+KO4dFDhm1ppXKAKgG+pUp6aSD8ExP0kVYuUAkIJtvQZi4DpkJAsfADUtLVGKLlLyT
FYtd82cAlvtYQS1jNJcGtn/IaKLmlpdJJhsqXczj56mwzjvMjq8EL1mi5i0QclLYufOp4XC7DgIf
SscDB0klF9ZmflukOppcVRxSSFo6vhL9POPMf6g7BHunLbYqepkpZZJq5YF2kR6l6wKDefhrLa+r
Cv55uahZmY4eIuluQrEjDFeNvwDxRr/hnDOIW4cxE0mpfw7z7fQIgCHEr3PFVf2eKFpuuhepnFdu
/lIijpKlC+lRf3xqQ0qXQYt24rsxzQ1ce4/aS3jWjSkOddZ4ftyyhIyNrb3KR/MRz35iunO4lKwm
bIwdd13d61yk/lE39r39OiLf7I1qjR534GYOoVKz5OpYxYv4KCqBxm74ikFhxE55c3QWCyrbMdUE
IAx4lWBX6DtCdsWhDQfD5Ajtp8uP4+DXR7r8KGureeDdtutjnvaBK/YX6PLLolW/MfteT84hTQM5
YSnYwLk9Kuy3vsUpovnNEQLrc3RSN2yuFDncM3DYeaimkEK2tAAY0IdDkXDDgXjWJxh6eHqToWd6
n9VOxslC0ZJoh2QHUsm7JcM+4neJBjle3qDHniRkv+iEsT9FoHgkLCgGMvTt2H+feyPwyhsIztFG
r1/WS6i3RXbAoYxXM/WXlf60HB0DjO+Z0LJYv1ccsuWnekFBD0YvgVDVvuVq1xhCbCVKAar2LG3O
kXrDGlDwn/ic7AulUzCao8TATme7xqwXxoNXlkVGuBZ7w3YYtm6MZjhIEu0Sjc/dS01TZF9LrOPt
XBw+pWjYwfenTlkNY5vBdjINvSJCp4otVLFRVSfP1W44luoqw7mmS46b7z4NsU1CDRBLf9IBNFvw
e3iZjAdbfvFc8Jlgpuj0mBCrwfVD0w9t7yAFH5BIuQ6er629PNUtZxFIG8/JIzu2ydNIGXbVFQyA
CUiLGrHgQrve+b6wvbwZPMNrjEPaywv5Q+89L8VTsiXlA7Cio0ZKUh91ew/07BCkEi/EBHDvYtkv
PcS5SUGYyoiymddwnt7NlN9lFox5CZX3ip/K/Sieftc/ORZlEUg7odF8tqXqphWaiEbgUkI1yTa4
mVdGzJja1nhNs+KPmtARQEUoK1FO/ym7ZuvE6xzTNcXZi/e5gvjVc9v5Jc5wHvzZNYa9ZydMO/2Z
bpzNkpi+Owup/PGzADn8aSVryGTsr/1LFmUPNh3xJT53H1ulJgXVoYy0whG/lD0fMqqt7f+bNuSC
5b4beyMNo6VMufJvE/kXpfnu67/4z0G7psOWeaCdmzxGgUXu9tHV3aYrHH5/IHmb9BM6b8yVvHY8
eMWhLKvjYc7JRctny0AsWMcTF2DSv58NJJ5H7ezpFGYSsSQbnbuw7KldD3zitizM0rYTPiXB8On7
7vpDSNnUsJw0LqxUf/1F1YhtiPdlzVrXA99pTSs/qg+4pAWuXJ6DDFqPbsHDLCYOTuhTfrLBXDCs
SjIIR+PrvmnV7ehgmc8SgWhlZztU0z3IsO5DgRv06onHICRJa+hhdx56vooaZ6aOVrqM92OzFI29
/9I/jcdcF7RafFTzZZdT/9dC1BYGosWftYdoM5sh9MnNB9fqIpvawKH3kccjyRW7gyd3v24t/4ot
NwFQpt79Qu7SuQVaOwWbc3eyroLrQP5w4y4Zuk1EPHxezFbsTUAkgcz1IpeDAZaDl24+fa2JtX3l
gkkTapd7OWUX5l96hKqsqDkyRkzMR5uX4VBujqi9GGpnJ6v9ULyiF9kjZ9N/wCBRckx8NylunxAP
m/SLsZsrR0M/CBWrd3h8zNMD+K9cXXOHxBFwanWpMvo3k5nZOzND22Qy9E/GSgiYB3EjdCihsUEN
55Y8E7DSq5hiQNXD2pmhyRGlha2IdwNVUsyd3Dr+ezARriAnaVUdAcglkqtAQk5s5rPKSMsoPehh
eHOH0xH8upUHvhC4Ou5GNeTMlJm5mbgs0QU3JGV0buRQFcgEoBOSaVjCRFgQY9cf1RFEiH6yH7/N
9XWtY/EInJ+7M2+xQg9r36U+Rtk+XF6DnjBJ4jjcQIgyQ1bmlGVePWXbbD6o0xwGoFh5nFmbPlY3
rgmQ83yH5VT/KcoTGEFwt8F9i9pAESF/IFyaiRSFbeTyM5CxFvkb5yCeRZdOi7/koZocEUXrOXgq
14A+hhNcA/7GwOznRt2K2Rz5iX6CafBJAxJd53oQX8fosPIVuwzbzVmN20crzgicr6SwN2o7Zox9
fY89muydrQRnkF22bY2we+6J4FDtSpFEqZQ6aHkQWirw2xej8ClA7vj3PcQ3L8uptyJ+Xmxorg5x
YY73fgjEI3oQHIIjvejUVAae+HiMLlM7+QVeOqQPVqQMoeXUZfkTUm/SP+0zalIF3w/yEw09LGl1
Q7krC5JASUyT2QCRzACL1jeUCQntWN/LeWK2rSiWAVWt1e4qhrRyodlPlyXgdo1qgr1eYOHbnjqE
CMoiZUpeYD7aNCWYFg36o06YYcA4ifMKjKRWxqVfdpIZEm0TWakI7fP9Bnvr10iGyeB3UjI/M8Q6
r84nvgszm3rLUClO8MqrCrWOJvHE48uV8Vhd/rPEv1yyj3erbbEWcyiXcP9A+N4nr1oSmtxeLl1P
8FpOlOw9TG0QEjKpr/PHNpfYGpHTUbioeqS1y7WUFQ/AGAoXsgF0a7zxImeejDiRIxo6SOWu4l8k
295eSGOO223ixsNALZkBp9RcbqkTD4Xfbb37sUij8/ryHLfPFw+VKfeo9OpaeOgls4opNVK7XrSC
xH9cPWjPHdtE9Ad14yBfhelV7xOYV27i+SSKG0EUcacLZyKO6xqZP+bWadsglpCbv4t6/ewkb3+k
xRwyXz4mhKfmlNfHUKoJ2+XmrTrN3QCRaXgLjSzYZV1Vfbvzd4Nd19sBlSdAsBe36JS1062YTjsi
oH2Ttv0DOU4HArn3htEwIsLp5xzFV01Z9oSz58hGRx20sbbIcS5C1LqJdL420ZBGKeYM35Q1c6hV
yr+QOJMNSeA5g0rqkcrxhQEFBUieiwe7BU/TeTqUzK9T5rlBgaDxOcYXLBvdg/JQzMIrW7yJtnYj
s6pL3yKFWCXwaWAbdruLTfQyjOiCLfguOs9FsEORvIFvbusoTyCj4g975V0azYMUQLyAWIIjUTYH
ZAz+rklaybnlK81CHNM7e2L302V7YjqaLxiRqn+ECnQ5aCCcla7HeBcyC+4lZFk54o0PgzSnvAz1
lOe1rdC+/AUBpBGRJ7EjR3K39W0dDFyYh0c7JrZLo2phSDRPTL0JY/DBfy8UiJ8znaMB+yxyc9Uc
fgy4KIGZ107GdhHnmfF7RfaKpFmCxK6U2mWpNqw2rNj7gH0sgu6di8qHnQhH+MdUvx5Fa+sJslhB
oK2KyGrZNAhTFzwdk9PbL1ZReQz7d56tagQ3cF1+YwRAGiS7vJdn3K0qn1Hfnf9zZg4uRuBIh7ao
wFct18P9kCEML4uxFM8BS1dtdR2A1Hg4h+WUCFeLW8Or7SzXxHTeqdJ+C5Sc4HXEyKjPZS9pjjnU
vmMoPcvRYmyPXvjXEVNEpeB9LZJkGbwS+xn35Me0bgmpP+UVyJicz+0C0rtkuwtgyxTJSvQqXcc7
G5g6NStrVs3ZihbgukMsjQ5TZ2Xw2or+fjibLmEzTztbITHsDcxUolR5n/8yCEI3C6/CrrHmK8hN
T2RkJ8/+ymrcW+hqE0qk7leSAJU10EbHa7D5hzvKeKuQ4jS/0obqeB/jbk3WJgRkbxlgvz+y8QFV
AYejwxRh5P5kjKWp87TERx+T3qjo5RI2n2/XhuQYutPcuUL+bkGSwmJEzBBm0kMmpUW/t+Ww7TFF
BZIuoepKj2T6wHqEi7O9vjzDxDRTxEYmEB3BMDaVWpXyMBsbYcJbXp7dqQc64OQTOzRyEQuQkp0x
v1e+5J/Kox7JIaj83StExX3bj+/aGvjo1NlcZ1Anq0NwX7uQS/4bQq/KnUpmRQhxZpR6Wp1kF1RQ
PqnCEQ3GdZN1+qyUnPqJRDKk/Emq1m6xHYeHiTsfqfH1HDp5A77m8tyb4thSlqlyzpic9tPeNCAJ
4x722oR8jzMT9fRF/w5RJDNNwd57CGxQj2+a/RxGLwyNbZtZKKkuv1LHj9pKNeNgQKoBkJM5XUjE
oC0hFUZGY+5A/bEyvlUEL7pvf646yev/Zqgod26jmXp3v+8CYjXv934/UXDha4+d+IaLIznUn/+O
gcPy/J5gqdw09C4AMhJA3ZBxojhY+KG/lAd4EirgPxftvxkh8VQ7RsHijCds9KVvRUYG/dCoAnuC
bdNZy1nEtXNKgHmzgt5ld/XQnUgeHldIa5HbWb9yfrPgVgflUSKeSjTUnqGa833k1KTTZwr+ObkW
1U/g39H3sz0JvEmsXKXmnyUvFHf2pdrz9xR4KOlYMj01r2N7y13Lij6UZ/eD1hGM3iAGIXci1sv2
ybv64JmWo1MFDy5VmbE8tXXT8orFlKkAbOapruTKM20uw070WNA5oj3Btl/+Z66Fb2H3H4uY3Fcp
QaUsJ/gT0KBajhmgXX+Ke9CmN8Awafo+8HC8TOa+GVef/+72WrFsMaB0IQcBJMv+7s8nhYefSmRz
GQxjd+eLMVDtmCw6GmaYE6nds8utPaocyP4DP5o/tnCP0Er2L/SaFuc/YRdeY97L95AOyCGJn5C1
0+JHJ/wedZbTTgDEtw2lpe2O8sQZ0AAd6S1TeaPY5IVjVw7hfK3Dxdp1GhTFuRWnhGhcbJ/OJM3S
j9oHx1gwZf3w8X966/8GGAi4KdQAVMCicGH960YAJVNB7basKDrpZCy8jwPM5boYg5CuieozXH3k
+Ws7kCfIULAy74l3VnbvF7Bgtr6LjXrkZq5jmGMAVQIm9paih5L3s+e8gbRF+bgPcjqkMtcY6LOp
JkRYBFXYyovkBxwNL6JDye7zpQTti5OkbsBJw8M8v/cFIRN7gXo+18PLMT6G9LlPt9We1xurkBrx
dvzicUnHYxnSbkGEDhkIcP6z0SbrEGl4NoWP2KbQ7UA0bNbRRdz7hCv2kadp1CutdsU6JMvyg7YY
rf/PPpRpF7PLPqw2grmuEuZjmJVM8H7/2XMKCR2s4s3mj+/cvagdBjR2GxOywKnP0T2+ufrBof51
QYAFPQlrnnO47duTT9KkgQ3POKcM938s/qiu85QDlLsB7NJUM3XGkqdB1JcWKlPAmEqiVK42hyl/
s6wNCq3HPOmxi2v3NAYyfqLS2IDrGnGKkazORVTxCXC3uibYwBaaSseybCzOPayurrGe53PbHQGr
0x/Nsy0j+JhotUKCGKSvTFtW2aK0+H0upcpJSej2b82VcbLEs5/SpgFtCm+S60zcRzJwcINEHb/c
EC5MqGxnyBwrsWjRf323lw5D6SBLTbwe0A5wqMGGpApzIlhgJeR4OyHMae11z7DT1ohiAUfC0Rit
5GLflgeMzTo9jTJqR4Brm0v+F81i940qDh5JQudl6ZqixJoeB7roMjkoU5id9K6WTa4p1m1T5y6c
raZ5tNTABIQWS/lFRWcE7szTqGOnwOvXrHB/tVah5UcCi85iXMWB9Er2wtZ2zPTsPgCjdwLdICn2
Kmw3pXn+25h7V2htwwv9gg0KleQX1fHeahBdSX+WcwJQXCIrO/s4ydZH8hnGvJD1KThKzEyf/0LA
3VkGCKveFP5xxTrQJNk9DJa6QCW/DiIEaU4Hk5QiPgYmmPnmhPj0B2uOfkscpQVBLg4z4lAbfIiN
7nhQfGsJssnyVUT0c+VfIM+vP8VKOlVX3o/T4XHCv8y2NaRXTTTT17i/aGG27gOlm/9jhAk+P3E5
3NYFT1Keqdkq3dd/yNiY/z8mS8Y6svZMMxAmQHiZTsdpbTXvVevlOSlIGUzFJQTdpfsYifpbBEob
qwo3RHASJlP/Bm7JwVSfhbLo+7PImJTe9xF5ZQDROWTok7w74RqAh9a6cwvRVLwkvFaYSmu4V4X6
ZVrul9AUc20jG/Gaars8ptCluiscV2jKBIgZ+lKnWUA234JvmToNxBjq2V0ubpHVldjB97Cnthhp
LN0c9kA/iy8GlxfdLMnAD2AXlTbrgukR3qIeYuSrcAigG1Xm9BTNbnuVXMSjUJmNjJ407R1n1SDB
zJIwah06EqP55+2wqyDndsVLrbhiq+8hFoBVo1Q3yP5oOAkavgvD6ORJJLGryhR1ARvpAKQuMgZf
O2jN0fgNT97cunyCGOD6b4W5t/s3BFCtERomvyri74Skph/uQ7u7XmkhZFo13g3GehKbNNhUehMJ
uoUtcwzJ/KJh1VKZu7XSOJ68tUg2Dbd86eTk7/07dPzcM+05GaqnbTv3QzZkjFF4Hz6BWfGsHhve
fVqDNrmOGRJ5KXkoZuM5t9JwuhvLvPJ7RJwhQxJ5k/K62fHX0fIN30YL33j78ZKDLoo3KfOFEYiI
amEk5fuFWJEHmud73hHLM2FxAg55VhZJQvhav4MIzxed5Yegei5kkraTZWzqFV2o79RVw1QlVAvU
gdfX78lVN6bbO4zOokfdTI4yQXV2CC/lQYTH1pY2hYCT/0/uRpS8sjgUIbyaOM/3W5y+xVdvNuY8
oMSDjYBW4uKndj6G4i6mtN0TZ4Pal1GrXj1xl6iT1eHtBd4lR3tvJMMa+zn6hftZjl8h7mIRx7wj
/+GlPZQMDqUDQtNoBClvFKNR9/ciVczVnJcRXrx9fPDLH5HGYf6PxKg+1xAS3Pu8LuoyPQ3DwTI6
yzU5TEOwciawDFcRyQSrR0fjRZhZk4l/hHFn/JyfOTA7f7lKGD/r3MnYcif2WONYU5AcVMq7irDs
/P89uSneu1S2HffXJPP90jvHsrL1h1Alwqy06w8acCje0ZFZNIrLX+BIp66RHOF8lbPjRjSn9pEH
rcjCwy+IoAKz78OeSbbefVYDmNAUWUo+F90gIPWDm8nvYhvG0fPe2EOvLrAu+J4+lEO+1IWCQlUJ
eafWsymPJmbx9fzY4HZDfi/BKiZZJYQN2JoqEKLFfp1RNq5afynIneMoZIrV1Nwfd3hHiT7DZVN8
wiKr9MYMWpHjrIyOJgNINbum7XAS9oEnt2VKl1rUBeKMspER3Cdx+k2YwI7ifz8YnAOHTzUfKTPG
riAgeAqgWwQhnH1PxLRHbbfYQUIWwOnyyyb1zVbQB+yudJFIPXbtYfEGGwsAKEwkBlePLcTeCA1S
mvYtCtNOaGfyTuo6dJu5h5GOfVqrER16rtwxoooO/rTyj9klJvxV724OsGWbKyrZUwWN4sf3m82x
unHiak1Fm7g5ulRKtzRVBha+DXDtStFuKZl1VBuEDh0/KKvRm6rv9PQx6XYENw2fC32k0ujfgHuE
EWsrpTBJndWbbxwjEtzpoBRmXw72f9cXyT6iPuN8U7LnYk3b/HWHRybznqZHa8ZtS3bQsZMFNLYn
E8KaA89LTV9qWktoz7araSX35fuiB1LakOb4vRQUki+Qzu4IsNHc9oqCKeZPXlSKiL7HF0zNRBez
mJ2cgemxEu/a8FDOHWZ8ZQDtl63hSyfuX6hMjEUcEaN81fSBnzIDP6LLvhp0bZVa1R+ET8nbRiK8
6iTTVWEEYrMKoAr258NNsLI1gG3VmqLojXsnq8afNLCXcEyhsASAIsI2OLvpedhUqyUU5cx1D63I
yhJSoA5RBAxd6RR9MO8q2vHoQ/ZbYgMUWIZSrt4zqqHurT76TB79gLuNndUJulI0YUzf1+1oVhlC
3iRqgTP3zWAtlstXkVdm3Wbp1szlRlamW/opPmCRt/CKngDXODTN7EMdMplmGItSQm2M9XLlbzMI
y600FGjuL7Sd7gT3AkggJsati9umf+1TTeAP9jle2bukgosYcS4MWgIbSw4tfIf70/86htRcLg2f
eF2vihyJNRPYx6tP59P1gNv5fr+G9BRFCq1xQVIkCfHTbgoraPVhhK16htI9o96H70OyyTehFUfN
bO1lVUwemYuMLI8dlXsV7usEfWoAd3kmlA6N5wSiT88Q8O5xAA4rp4+JboCm+3Jy4YG4t/gljwTS
ln4IT979q1Ilk1i/PikbtkPzJYhugTGHWajCnTw6Z4PFAhgp4FVRzD3SU5pNa0gSsjlDQJFvFfx0
YcADn1z0PF1UTz04Z8YOvN5h7kFRK5WMjw+1HXqK0Ih+Z+JCmATrJrxrnNWcINo+Mr19H/ckBbRT
sobK5cnjvXs3tUyi7tyFZ8wEkBMWYukFOet31+HQTyjuUUjNysEBE4TQVllL5Xh3XB6nNmcFaC54
pHWmOMPmRD1QvNlY55zUN1mCSP7Ysd4+ylo63aVT47GUN9pvGjIzdNIbsilT2t8nGW+NngVvyH+v
hfXXGw5n7JExYRvmvUl4KIzEeyJRLGaybWvaHMyyn/nk9sWPChiN+NHndmngI+WmudmPXoHEBodk
34AZk65kE1Sni3HxNWQe8438b5ucIiQWEcXFDdN8X6VvkDs+Z9cj6+XvzXQ6TzsJ7hz2d8m4S9bi
Gk6cUbPIRWCMxlrWcaZjkpyDdk8vHkvdgDJxeR3q2WwbHixe8c89ViKnNqr3+i9e6JGQWCfT5/tn
BAoM6uiaFBBAMhhW08dAfT9G0tcRhRl/SoxQUwXNu5HTxXSnBvRzKHLDtJFJQUEDPRGM/uELUjZF
MXneE/n4UI1j0pf7Jhvt6ZHl8ZANzFswpOiuSUtgmN6itUKQNbxcDjRvnbbHXeHghM/jlxcM25Yu
VIBWd/cWXenO5dzo2pQ6EOLnLjrON4PkvnkhsDNs4nFDci8IsfFS2E5fTNsbDUACJqF9AiTihL38
OiWHdab9UCl0vVQKCdUMRtUEp+2fWT51l1DL6DJgqbzwsJxpZ1wpQf9maLBwIokFgU9Tn+pMy8N+
sM9NiQuFFbM+QT7nTxqHpTLbeQTVYk66e2lzneVUjG4cJgDvyQk+xCskNNHljgVANFJf3zPsDQnk
3p1MRb1kvrQq1aDmgII2tQg0JNv4KIswFEiadBRCtrK7CmJ3hY0su+RaBIvSbiUvj8iFrtiYH8xr
NOGnzXY5k3+uJn7PhJ+cAe0whwIMYAIsQRShCuuX44RnHRC4+9jGa8yV2eP95bkgigu0ATyhu+w6
QrdCYma1eaSN9zsax1cvYd0Wand4WeZEilyi5Mqo+fxFhtHVF3T5+96NVg+oKXBB/i7JbXfYzD0g
Mx1KKcFc3jsV/GqqzL+6UMDX77D3nnYX7beBRGsKi44op7sPftb05B/dIu61bfbOBp+3kSbDIE24
hDIia9VtfWf4mcCgM2eqqKaz9DlXhBcRmKxSJp0EOSAegSFx3qOw1VoxUnXcPIjP397cQVMCNYH3
fPWtb66FvMyhV9ZVuPQg6yPmc32y/33xnZcxUG/4PdTcYyeervfJX5PbwH7ozqNyGN4Vgbh4dsLQ
GjQv2cc3f6yFlTXYca7Qgu2sJoy5iegrcrmT28LcvlHAEPOXTMQe+gvtWaqv9/weOVAjbFzCmfA8
6SZm4LAuhPGMTVm4XEocjUn38uwxxJ99mO5ILY/Nxqkps6MsQCFfFmfCx5PTg7Wiq/sTlns9iB77
kIRIEJr1SPOcSpkHTp3sC5ixGHNswJxiSWh1bYyz4NhVfxabPOxTa1qJa2bKpmkkQBYRh3srRKA6
7xIG0gS9FBOfqOiyZWoXsKHhmnSFmYf7F4XlRBfHXWzXp2GhaiYSjHUl5vh+VzN06y1HEF7dy9qw
ILsPjzTXJz1EnJ4hwoHIraMtc4Z+vhbbe3WQOZFCRT6znf178fzePy/fugPqOGKXAVgFUqLZNHp1
cdPIYJdukERu0bSA+X0sF3EbzMlgiUglfuOpQIqZbFOhR6ny/TmfaqeKCLt306927WMO7LpRWcaT
FCUREQMvyXrD0GJ5OGRp3MbUorbcTPs5/PxI1awwBgfx0Pc295xPgStSbCq4zx4b2IF6NBGIrzcl
DPt3s3skHJNyOkR0/AiVs8eQmPptLxrtXq+uEkpDymxZC7TeBsp5YGUoHyzqFtlsEwr/KGJsp5vs
1etI4EA6guqQ+9vaL7GfDDQ+zfcToGu7bfQVEJ2Q9bVuCFStxyGO2pOiIJuq7FSjc49ykWnZsrX9
k3Y8WIjrxdrPTOh5cpVdSXwg/4c2N/2eVsnw6XtjgFLRXT04BbNCAABCcaL7P+Hwwrx+FIVbWa6Q
PRxO5QmTRFltCMml481syL2DBCycr/Wyy4PUUB1dUoJGt5F9T00eiGmY+WH4CMTWKd2+eBT9QGbr
aEMA1kCUmRkh0e7rpSs1ao1SQgZI59SDOW07w/8fZiD7BdRggkBJX32xEsXIHH9uB59zSenbZJHb
fMVD/Sew/HAVuHIipGL/vj4KsMt5B0Jj8XPzOXUe1a0n14CxiZ2Dwb5uR4dWUSyadJXDT0mZcH7I
mAQjLfMFQb926qoUmbnJogRqQTG41aXL8ZKUh98YgYHajj4U7RLiQAuv0R37RcYl/FirS9YpWNoA
P32iai/rOnySHZMbxwboMu8+hFYFqKnlpSQQ2piwRtzd7VqSVO/7rRNwaFoDfwxFUemb8czgI9GQ
s6ivwhylxyYKOOgRJi4swa6IQfml1tkdlXltZGOc6CLOEysaIrLBEa4nqPpskQuUfC5RcKW6PTuJ
uGQp7WJdwUMwLzxDfOXeUhKhvAOqIZtHkAyd/wMeKzpnoetO6c84ipMH+sfpaeOi+SOKlHndQ595
tdiA+MW7FITa1Iv6pxWuoCfRXx1ktbiq8V7OHX0CX3UOfWgy2uJPYBmJWiCW9ZGVkrgV7kmYe/aj
GUTkJuY8m4yrZCTGRjyRNZIX6fBGC3L5Y/FmCjqeS1vvVnaaRYN7/ZEk+okez/+QBN97caal4lJc
vOHuNJ5x9fqyXXYq4id8WgWtqucZqcd2YEHPAADsyk7ZsrC1hmXAtIdFklAJ/VoQORqyczgRiGNT
XqnQhjWqvZ8sJ3ndmBXP9IurVZmduNq6Xxd9rInoY5pFJg6+5Rcv9ItED6NiQ7uw8HQ++zi3/8w1
C47OsmkZQJF5sM5tVS4AN37wqJH+Ii+6XAL2cAqa25sZUdcXE3I8X6M7eBoV2k0Oh4QoKpRmkCiO
xxTGMDgTjTwuXjhG4bk0twItapaGuhAXwNXSOV2akwX5rhtDwbP7rB0bpuS6R0WO3guwFQLzpcCv
g/O+Ff/nJF//Zd9yFum1nz8tJXiBeRGvca1Urku0UBo3yc1Jd+x2fU39qS4iPHNEvFy2W4BxtrKh
0yfrCp3jaAGG3dGKBK3mt0rZXWi8NjXObvAbT8GpqwmZbn/sZYS6gYDP/l+F1oaPpAyLJ3/dMFu3
eqLxs1LZM89NPBesNV2xQlWzvBYQ1xbOIDWcphoY2KIJkmIECmMdFVHJZKEtkGbcBN3/Vu3LSkV8
wo5xf8d+khMH7I2MtioK1Bq4mJf577TTzqaID0+mgtUdMhA/hVkw+vaxAyTLQ8I7fg7vOSxYUSC4
oUhwfMEWpS/fliysveSzPu3uGjqqdlVpIXkCYiaNyJUSmJAT6OvvQn6cjO8Qz+DWAduIyCmoteC3
uoJhGn8l6S11AYX/9SOpFstRnKNaNTaLFyEmRYRtdHsCsZyP8kd6v6RBZKpiG6Al3wIm8sCacvAb
wO79rBTtU7fGBF87TONXX90ZRX8jLokWyD8TERLdaoWY7m52JJY4HEagFA+KFoSWds/pDbSdtXNq
qKZH+vy83aY24ON6WX+9USIo2vz6cKpWp0yN+kO9InFEeetOrkqB0HUNKq22GOfYXoV9GMSkTi6T
GSrwa0mBop5FCewFfNbtHcBdddifiH0Q5Of+lUahBG//jrSUhoykPkHND1GPZyql8avePiq00M+s
VWFCuKjhaAB3LrIH5QZmFjP+PybXunUCckQlPmVazeTMC2XecgCIBNCUVLMd7gWfrbaMjjQ792RY
kLufU2zIvCs9cQIPn/qmb2yZVvCOloMqED/FMt+zClktQyHWf2iT2i0TLvDL8Qd3sC2XyZdq1uEX
esSZg4CiEVYPBxyJjUyO+6t5R62heQ4qXgfECMscvLFO96V2a83opXM2b7gyCohsqPGP+qaTK91E
jLgcZcv338H2LfHwo8ps5UnWoHavJyYBY+wRUm85ZZKaZv9NAFTLMRjfi5D6vk39uAfGrR9wMiPF
ct8MW29EFWdJEAarfjvBWdkr7u3Z6egg2n3xE/gyXy5r/VQegSf+FeAntLjriWxMX22GLytku3Vi
baIi7F7pQFtmyvxKVKlc1USaHkw0+uWUa02gcTPuxBv6OThXEZPAqbjQoKP99cdhOo/tV9WFYqL7
va3lJpNe/DleggUZJEyPsE6jKTXbwZwdSL26R+g4TbI6n/igit1CYQmlwgSiORZa20Od8j5AMXNI
/8YD3FVhvKvj8yR/e1tlDdr/APRGVZvFeUj4yBuZ0oEs6wpuAeAkBv4pl56WDJERWfb0rQymY+It
RKGH0pmYKPH7ez8qHNkYNfhvVYvLhPUgJiyDaOzUvHFP+ts9fqBM4JBR1lTmLKAsB8NEjjp8rAkS
TJGd3wlhOSKuTpOjo7zJ6ww0znniqIOF+P/+3yAfrWG7KvqL/cmxcEdFVxFFbONSnoSQ5DJHewWH
c5MsBqLl0iOEHx9i8VMCXRbiIS96xKOeAyGitqNQx4hMH5uvFu7xr3ymFpucdysbGmXXgBpaAn2P
+R1j+7FYF+8chTOuUZmrYqYrYnSo3PS9ZEWpByskqBimtyRINtTyE0bYcM+5Rh+CDT9bfDkzZPFD
FkDb52+7LafdfdJ0F25AtDXDOBTxGuRijSCH0zSSumMUJyN85JvF1usGq+wEC7wvK2AMc+Qh+E4G
Z450fugKWAEpKX3crQ2v+xKSHWDqeD1DuiJxyqXm5z7mFaTcQSHGuCYYIGtjYeLdO80jMc3qtcw4
Zs687gxGoD8SeeeU69ggmrm0CxaDwJWiUmkcCZAnWQUc0IlLpNa0rN7OAWtRCkBIDSjqymGuge/a
rj7aQWxOkXC0e4CCoK4HQDvyw8zchdKRDfCAJjMV+DwEp25krYNMnjUIwAs9QYDpzUZ9DtD6zLfT
LjnMA+mGeb3Z+31kLXelN6r7Div0gHxV8lNkQgkqX0BXHdz92JThE+pAgbsNXWeFHbNd0eWHwAqf
YGzRzT2ePbtquD4RDrw+YtX4r6VgWNNLROOPQR1RbXbf5QORok0XWahVZoHC7Z7pK9BUrKx0Xe2u
kPYBVy+wAS+RrW6Nal8aNjIquXOnS2Xhuo5ny6gxE5lKLEnMqSiR6eYi1bvmcWIomJSpduXg6tf3
WP1IhAq1IwHwujiSZ/XvgSLiWiQrrlSQXCwcCo2fOlSWmHOE1XLXLedcFfZ4PQ7QYXEngg2cYqwK
21TA4/ALZvwQ6B8yIC+b/ZxwRbwQOdzoyXTw0EBniSoPpHBALTeCcH63RZv0p40is75rF4m1xuDd
YPFQmIiPno2JCik3Mi3G6bK7S8GSxX1rlmsDFK3co+OclGFR7PBjvyk8k6Xmk/wiStvPAkKtXhMf
q39TsUx4ys7Q+Q5zLeEnBpgwmt3vAEooufbEdrCexOp01Bdryz2276MRe/b/IDkMv9zD0WdwNX+R
Y+nP2sBD4il8sKsknhSXv2/dEivmSiFFRCWFnGkFZ9AE9tFkgM7VhGkQFbzTDkLV1FqwRdv/rgvo
FBKW3AHoozUcd7PgDw/AB6m6v3A8VksWYRV/f/V6P0dt0fY6O8nMzfNfhmMWNqs/afcROUD0ChVz
+vE4QkAXqfwnmtd/SjtQfVHapyxT3nLr0oydQzu37wuJti6s8qf5AStDq2S4bgeQBSNQ8hZJInex
txWDLRPK5hMuZTdxzH7ui45gVAwhg7uCQ5iK+LpU1q/krUI20NRxiX5l2PYPwH+2uLdYHjBNwq5j
aFmR1Hp8pQL2pxVbxhGtE2JHZ6U7MgKhbpTCFSWMYDhSbSOk0tWyvVgae1m0k0C23nRA2kpASn9g
6oVdaNOvMCx6mAcsj2UolSAMbpLUSUz3/zRwqBm/TeGN+5YB/jNuEyXswpdfRtjLuj90NvnNpeaU
Zk3nDC1uKGg4xq8ywMdcj6+LtUdiyrWw0+5Wxou5/B9NlvOIW43QknnCNHTDr8xxn3HxNHXRknjW
uDgP0Yd7v0P8DFhdXB6JRz12+1hL0DLWSL1e1tk+7ZGEaGK1x6NwJ8HJT++pkDQuQxodvroWdw2j
GMFjGKkH65chDf9870C7CYrQoqH5S6sIVgkP2kGgY4wEOIK/hgDig6htKGepCuftl0l38QnUqGmL
nXCeb9JF2aEznxNm4xCewwA9DPDmwNLpPl19woCy3M3aa7NiyeOqKv7RHv2yo0DsF3oDHLeZlezM
Zx9xoHM9DWIrXSmK7ZAtG6fwCIDjOGJ566BdNfixlaZhufFJhgqi6HAINxFhAGsE/sH2vNZkPQcp
0BTVdJnnipevKIzM6vENQV6U3sLQTjQlUnpN4KJXDwSEUG97Pq7skTMOsdrfNJUNTBCEojFmTYbX
6Rw02H9XLSOITAbViQ28mdNXeZqpnWsokRoc1YgkXscn7RlCpocTABy4t50SHKqJ3twT0sur9LEi
7eyYuRAOVtmbIJpRXhOhi5QoG5P0mdWMa0txmww2RsCvo4KmRLiQcZGzG7+iwQAT/Dlon7WEgTHO
UVc+RGwmKkgommHhwarTnrh7BCeu8XtyB8dQ1AZjZW+0/KFN6a573e7sCaOevJSALlrCgSVlr3uA
9Ci/tMKOr6g7lyJYGR1S8dmHZ95GeoVl9D5OBP0e305HhjJD4wQ5yWN3QwpDit7paifVdgIEyr5H
5o4iIW0CnMm+NTQDVTc5iA0KKQMZlRf1NI3Wwtm4cPKmkqYDI4NSHdZziPAlJ5SH8A474dQMvRlL
nnaAlSyC1Oxuv8RdG7cYRSc3Ajl1ZqXq05mfSBI++rSvqaGgFj/MwCpizHpp4EyieUH3oSAZxoHP
y/NGqdcJjV5HwEJ0yd/IXBJr/7Xj6gLpB7AhayYMA4sJHtBb8cJBtcOOzm6T/X3tOBVwaM/Qq5xh
5TrF74111D2WEnuuMrRG0I38ZKlJ23DMe5S1ABcMPms3Dz+AZv/RPKmvAseMd+K/GtOLQHjJl6BF
MkZLwHo2oXBTmOdhoilsQAkZy0q8uD+ukQUyJhV9Y/pa0kG7XcygOWouzoC8Gyc9mJZC178XEA9M
tTseSzs9vNrzQHb/vv/gXx+mk+hb1kv1tJXb/ff9jO9Vm3gu3uI9ywVcpUm6TRd+0+D5BnxfGjfN
CkjU654nKb2IMF2PHgfRIzFG7n0t5CNY72xLcpY0/sa3dThir2BascFEPbq3DGkT43H3lHjygBiG
5jVMQLg1m885eU7tXXAO8wPFHmNrCpP2/M3SUaksYoAlbzT7iYaQkw5z4I1l4wHTcXZlJ7y3lA97
9e36xyQYo5LHQYvoG15XMeSzRTBbABQ7XVgA0euqkJCOGd9amrpqCG9WBsyzbjLDzVjSFjgcyY3P
KmLeqjZRRq3Q63jokSa/FVmxsrzjAir3OqQgdiHIfDmy9vB/o2kkIxNxtdSTZhoQHjpVWKi7dGGj
zMtfrJPLgBc2B26xS8w2hs6EO1r2risNr9m0kpGeErIyddCay9sS+RWI8gRGqZd0FulkXN321a9U
64uwAjpKfhLT9j5wS8yJzkarG70IrlZlGB2pcxlwCvIs9WKOc18qqzgO1Yu5YLcPb8iK6PLWhd2j
oHHk8nS5sVYCqGK5aMb5wLwjn0mwOkl41BdVXJv8D1NV8uHUy2MNLOtgSuiaTpagbSt5GpZMDdaS
ucYeWM6rWYcydPqaZlriHB4+4zJvD0SWOk5cXjWkm1hei7hGusal6A2nD2xMNfZfW50C/o2drV4F
n0ppWdzjGr+1axbS9f6L+IPQc2JbmNpPhsiMMtYJIirZeWhnwFDbphbPS5v1coe62PDHzHoKULhX
XR3l9dVY7pbpvoWaFkjmYGvZ7R9b2ZVt8GLPepyKiLpeLrjcGYudhyYFG2+uc+Ufz3IVis9xn4na
JqH7F6k8tCNs9UyjwOw6WAS/VGsf/bKvw+cmaiyjhekOGVhoBFW9K6RrfQPFyExMOQwtAGuxt/GJ
sUxOlV1WMFfQGMXkMdD0HT6btMmuYsF48i06IYr7ZGWOcP2qb3Uzc4vEFTEnvf/nMJzbgWrLvlRF
aENFGsT1tsTMEK14i2QjLiiAYJNnsGNp0E6nNmQ49lid9tMlNCIuBh7OLIFHWidvlmghG8YzP4B2
W7aVABKdC6YSlzxgt52OoV19gtRT23Nfoa3FOs+ZI6KHdVzMXpe+4VnQEzQAeH3SqfNKHUigMiPf
0+3JXPbmb79mDNkvNr5h3xhnh+sb8FSZanrkFRZ5mwW+Ljx/ZhpbY7RtmhgViyE2LMK2ip8G4wWF
43qXKnl/KZa/Y9Z6r2u7UCL84vxgc7hPVQlB0S0DWGCCnFAniPBBtLUJBUCYDujt9x+Pj6mBxTkj
K945TpZ7P8nkihFjfqCeC+FsWahLXcC5y/fAFkBQSTE4aMqAIBRXqs7KIv+vFsNlUoFhYVZEluqM
ExQrE8EIWt7eQeklMQGLVk0Lu06hyRoo7RcI1jEpSEZ4TtMhS0TzIMnOFtZL/3kC6sgR5Erx0U/r
4cTBf6ea+ylbnDuuYYTL8zi47LRoFI0d8zHQGaZQxAqtWDcpTTMg9OKId3c1FyTx09zEoNCBOs5O
nhlkkpGvcZ0KnnBmEiqIExPPi22/8+K5i9s5Ohtiz9O9cD20Ns+z3g1z5bcmMtX7hAuLc5pQrPMU
aVL6ZHBL4ROiYk3QUh23zX7JYIQCkd1aNRDtxrW4CpWyYoJm+kDK2bRTmzY8q5AVBE13N6allCt6
zBnEJqdQlx3XINcB2nmAPamDDrfqg1xdwCNC0Tqy7uGqlceXGTB01n9LY4A7NfhkWPqXDQHDYrX2
szaxVO7UkkXAMrctWq8uhONRKbB1GoYZ5WPVxBfv7rUVPxChrPN67tEsxfofXsh/GtQGkLI6Ye3P
KQpsU2CE0CcpYmJCeOSGQ1qK+HY95FSJ4Y1OGnC86X9kHcaGv30J+gj9gUrWQX4LETw6hdzmfl3v
nU3rOEKqhRi5U71ePex/YRsHgqkTDemhoeADYUJhgSykGBj4HA7xgJXVzJxIg/WeY+9M7MbaFd/v
q2sxYCzQbBOwBBZi4q5BAmhWGmhyGvrQcAvLaN9gppzpY1llqgJO/qU6HQwE7lCRDJ/yRpoVJcoi
tkvJX/Dmo2nUwVZIF/vm0YkK705G3F1sCVyWqYqR8NUyPIz3eCm3WwllSSNUhPnGWrszkhfyG9Ny
XMx7ughEuQ6SRxqVtL/uGQr0VQiWXR5sH9FBjcmVcPGmXOz+9qyieFvT63N30zVZOAcWuTis80Ok
0O2aAxiybUtTnAI0NNyfNjrmvvv6Hhpe/WyO+ROxt8a7MipaJqkBJe6TSqUj7IwwF5CcQ4LkF3I7
orSAlmq2tr1l9QUUwUAN0Er+czuWAYWWknhAjUYQE5mKVia6RUh1V+sNMZX1FHLBp9swvvUqnDZq
xzko8RmJqQ8s41sqP9RGEPEe/kgjA4xsGEULApEmHPxenZ8POTRYxeztY8xpmTfG6JAnzV+dSZWJ
9h7kxrpaMrsKMsUxcZ0c4kss8GN7zLRyIzdq7y870DrulJqyAPaMyQXOx0D8FLZxBf+tTXBOcaio
1vHgAOFT/5YMLKeNfV+BRNeVrROKSshU7K8AjdWrtm3F48zw6pSKnVSj/48FKgyCFKtKZMamMyRT
22y/bWmVCN4+hL/9TlHMZu6P6mrjWXm5dEkc2E2HAjl08sYMVTUoZ/CXN9LJTddbg+m254DxIzdq
pYnyealRMID0ZFzdg0uSq8YTNoQEUQf1o4PFL7gTIKezkwi5YFDBuf6RML3GF5N+hDH53AZ4/RNc
9ECMDXigPkDyiUPWy+Qzh8JfmfdpTFouCFukPjHMd2JVBTksVt7nC0DEp6c9zFhXc6bdsXaL1/3/
OeAA3yrhqK5OKR3TCdr52SVkLt75YSCyu76txItIJUgvuOEMf2j0129Cqd3Rb5Vl6lsIPudtFDM+
vcxaBGxnwXiSNPhv4kK3SbCY8rIc9qdor8K4Hi48Z2cLfVwpB6Uqs5cQ9YKYy8cRZkQZ6t4Fg6S4
+m426EtHaY/wHgIPpTD6k/7/nn56xd7xZIB59r+pyCeOMHVrnQD6lCLDYgjYqvp/LrjCXBIQmRT4
K63AVUUU90Cob7AOehcPFL1Baf0rIPqohIDQditeUyIaWaiyoBkiffbyGbJ7PU8ZnoxdrCHP/BAX
0v5EVNqBVj20H6m+WHv0lQfPZBrT9iXYnl+RCdEs74wyCiGiH73Rr6g5kUbLbe5yhD4L6qi+RWeY
6XD6mVjDca2KBmrsdh+O/Y/3W+PSeoNa3vfJgthE8jkaanxaasg0TYOkrruyDk74a0C3A0baQAgf
Tk9F7LwgXo65dUm5f6Q5LJz9Knru3deWn9NsaH/BFfSg8P6HpoErHUnarwe8lF6/kUNkje+fvH5D
jVKO1cV630YxY11+iND6Ve7ibmrJSgC5/h2LrvGY//UCbn2x2UzRK7m/Iipmr79fKke4y8JG7lRI
2nzU21V6HqdZgcumS94+oGCw52gwUh4bUYpsnWldayKAd8f3dRw41ucIRSOirPO0fnd7GVpR7c1a
JJAtWkrVTdpLn2/gZGV8mIWa3pHcFj9inz1kliUR7PIU+J0eg49qWMtvoe3tk5fp5LIaaF+OCt3C
3Wg2uBnS7TYVWp/cSi5kYtamPtT9ExVfTw46QgCvBxOyHr6TAgRk79zng8NRe2nZGDRaK3s11YwE
jz+6/NIi9o6LmQZmN3WzaPf1xczNC5LgHBttzSYDadMK+cz5odPUHnmG1wmSOYrYoNe7PS8GlEmB
TYY0FQG0Tdm6wsxlEGK5fs4dV+Kk6XVmtKINRGExWDMwkykg913Y8DiSg6cXCRqW1SJYpo3J/3lm
zHtri9gUH99yR4fOFKjgVC7z1mdx4HVAfE9dfSVOz9IFWR3qa8i8H7acFRHAahFXFgDXMLzR9EbC
38GtRpummXEwlFjJbRO1BglNeVBTnVhIrneLH8NyELFh1vYpUqsIVuJrAOhoLnVFeEwLGqa5nhCD
ZvRuMkJonyNuX+JV0omCwEd5V/8hywXrWimdWNimb7dLqAQ8yHtSkRarGirpPgxZuhTAlqxPBnqg
mcBmfhLEvgNA3K1RIdIG2QHsz2C/8pN5YEUVGdmyfOYD6gLr0Xgf7smKvUejgZzTzYpvbSw+U7ij
T1gc3BAdtcbhyw2wzG6QbKo600+Y4R++QyBJOViWThq7AZf1PLnY+2duvkDa8pQm8PKcF1fkaKvx
kieY6xMS+4W8AS44Yf6r6rzDyEujnv87rplHMc76Fwhz2hfnDpIxFp92aQpcdIYfeTXxpTvbdhT4
SNxHcdEed9/Mcaphok+BU0LCLGw7k2TfwdBlvY+j0AnF2luFJkORGOUMhis4m6tC4A313h48YSb0
wVoJolohVdIZu1YiDvajJjI6OhFudQD0Oy21HfIme/PfmURfVXU49RLNx3HgFy55o52BOJbMWyxM
tyMQHCqDX8YFniZDU30wAQABQDCgqZBf+XnVndqJvc4zDoledmvXb0BbtYjzUEwHWQlB6Qxi5AIw
Cv4kR9EPBVje9C9Hd9j1ZzQqKGc0zzfHS64jFPEeRb6/HKlSHxRo13HbniJlglhNpj/S7HdupZEf
CWqXIR2mXf+wGps6Ls/m3amqZPZ0jtuA0yvIXofpztbgwR7vnj44zrKDyGnMroJ8ylHeDveM4To8
Y6dAUuyPhYkDWrPzwFVPRsZ1+AsZeOVYFvCu/d165iqy283N9rTc7kAQp8nluRwj7lKQGScP2AXt
UgiWHihIbAGbnVTPoy/dJRnbpkqgF4kPem1/fqKezwXuQrv5c9oUUfQ8WXklL95gK6DV8IObrYfZ
1SrHPCv8VcBKE4f3nGu7PnJsDkwKWMjIVQTxJirXjf1eKd110qyKiBePl/MkAxLFpJ2RmhWyK5Bz
oKoThLO29ycjzr3fPC1H5UuA2y3fFJIB0uqiam1FMC2uPSDS3NBhOU/D+ho2WpHS+GOdcZIEmXdn
JNq0Mvw5aM4JNltYoMif89BvN51gZYNLtIw374T9uP6B5RXm9BOzxCvO3vINdLTaYakVUgtSf1KQ
kJbw8xvrkEWMhXUUSOxY5ibXC45+jf0Mw6CFDgNA6zO8w14GtjfwcPBuLjYgSOaKK86Amhyw8NZD
hcnyCKGrlAFVKiYZNpaT9dfeKTwaYP5vEEXKfyJG9EDVLvA9UljCIWwb0/YdAaCr7jKQCoaQSJ3U
Zv+W66gF0tkG12qsZL1PIO4dXeHmQun1Y//KtZBUsraVJZSOxYntq8Zc+l1y6I0yzMNxOLFbUdiS
oHCBKxjWOneyBCzvQJbm9cwQRER9x0zzCVokyZdy9EHkDQkxYzdulqJk8VfedvJCk9636sEmLAuR
jbetg12bLtt2kHKGR9Mv4EnSBUnq0k9YU6qUw6ftFh9DQdDle2F3ZAY1M5Qji9z5v0Sm5VcvYUSI
8BTVS1A942Hlepx+jtc34pA6amqSWx5/gQ5B6eTzi26ns7goRNC5tP5G75iJr96lycWctax3LZWg
dXuWGCuSs7tvk78ntlMKw8tETQE88mbLJTi5RRnUdS1QmQUE+zdwDhhFQjjMQS+D+ny0Pwd0DFgO
kHOFLTq/OH5wW2ifyrrC96R0U6e5m1omYb7sIwQqORMqQykLJA7Zj7+5tzHGDLcW1eD3ZX/vN8+w
NzQhD0DX9ElKiEKY/Qao9NipP9tFfNZnreno5na495bL4Ynv2MyVlzqCM09iM/m1QG4OGgYlRItn
FIrafy8EbnDwBQcczR19/L/mDhRku0BwtRgOfbap92mL/RPU432tjPY+qYgCiLfHZohaUHPvcynW
dGFHUX2zOy5dzaMxjaLqga6SK7kbpyNZkMTv9sXfeALFQ8nrv0jCbGpm6hzCTZO+6Axkd77WE+Eu
zsqW1Oz8/5pDF2q0MHXdN+bXJQkNXU7WkY9JKQ/UrJDsS9DqKs+jQhhYc3aRc0Ud4R1lpUpwhjPi
IZyV3uVm1frOiu6k8kyGaoDoBSE/H9Xka1JqCscvOGcBt5fpC3UW8iS+xqbyRWLJCPmvs8IrwEc3
lRWr0dlT+8w9D+1jjUgeC8nt58WSJzdqrnAmei5laV4FdYDUZQLFcyIuvH1xBQKWWMikdZfPKLME
VgDRCVy6137raEkXZHoMcZkRoeUJ4kGs+OlaxnQYThkGO3cRhzHa4h2Q0bIqhZ09cUcoHNzbYfcj
xki1nDjoEY6u/OEj1z1vYIA5gN52jsc7wisVvArmq0rX6uxAtY22jZJG/i2dcVnUx45SNJcepQMv
CksREO9k5d7bS3k5Jj83CgL6bpDW1mOvCcqYfcn0GWJan7kbdPGT6Q3w3MVdHMTBne+Q53D5Ak4u
CWzngcpYQ1g5zsf512QOzosUIkBXCHf7+VJk6SkBD+e2e87aiH7ScSEEbKh06sVKFGvZAYI7ZSYK
PUP0aJLAtTsLcFDjf9IWAAaw6aL9FeFkm7ipgQKbUQ7rVRJf40+vLml+SRDipLsLnjbTiI26yaM0
NpxFmFXXbNr358vVfyd/GP8gNSVQsZuhNUZ7fSDnqcPcQfQJzneA8XLnNNsiBHcl8ybvUBff6tJs
/v+H2nZ+VNHIIqkQu6+Ku/2jk8ldYeFmlOOht/EQ8yWZMkast46l3mPNKHGLUo/AdKFR4iKLaPDX
/IAGiLd+mAZUueaF5E6COGILoADY3AOiZmg2qzSdU0iyTIEwGNGtj7iQ4rPYcSWZKz6w+GHGOfsy
ZmnQvGnfc8JKDuEg2uJpNDRa8INWtGkZPF6jSwDKW1S/f/MPcD5WawdZL6E5XK3C38uyTOcI1oeQ
Wj9xBdfXEy9gtXMrCaog/MuSTsgXYcRzwW4kc4au9ueSlEqi2SUdQPvVn+0aeLphxDyxLRuBEPwU
hVfkuOM2HSYzXGqE4lzmcRZXSluh/wO1eDPQByK/boAeRvw3dwhSs2NNaTpmqqQ8K5q8y+BpRxOx
sDSREDfxtSpJa2lEdzSR0Iat5yen+fbzbNXB/TAdmw2tki38KMGrodd2XNgnBZTiOOAx3wE0H+xs
GaQuUvY5z3T10xvZL4kEIEJ482TVth8R5qWdF6Yd59aq3LEVxncyMwBX8uVYFGnWdljMy4ERP5DK
GKVnB/5Z5BuxyrKWUCOJokrM409Fp9cPbyB+zakAa4FChO8rG0s6binF21Ltb+7gWMA7OMLa1mi9
+4YCK4o+TFne2SGNVs95LWib9SU5NQnXnVX/SjdTHxpSs5H0jzAqWRsBX68ZyG0bmx+AG5erstEA
DbWOpDCDydMnGYwtw0yJ9zGCDFyoN1fWkF73McxZrYLs40rC+xWntddmGSOaTx1c+l0QJShjCt+a
NUkY4J0B2uWOaRQNwKCXAtOR3w35Pqscd5JuyXHBU92Tund8DOYgJW7XHSEIKcMGXvDJc4b0s3nY
qDdDAt7oZarDAfi/mMcDJRbNZ+LCxtD9RtAwY905byNdVHARu8LxrQWLcPyxDeG9eQ0/J/Klk0Yo
kZ83qJ8ingC7aeAi5CnWT1LYTFlKJK399md55wpBLwy4WcXxjy8+bjmpLIEkvJTFprRYUFtRQ4lh
FyEt17svbKaDM/+eLk1cJU0HCu+zw0BW/DH6gEKK14b81z4pBUhJInZET34ta1iHaV3lutCQMeWF
X2RSfbZtRpNg7tmG7dw0Q75a1cyzA3eyPFPOzjDOaL1/XF5ZnI+UoRpYafaYQSbhCK5wV551ZC/P
eRwOzcgBbFMDgN84aygK4W9gPUydWymVLyxqms6PWHmWVrOQPzRVwd3w3KT6wpGPpBJ/6FPUc3NT
qd6IuVyYui4M5RfwDUB2R660Xhj9ErI0iQoUTjwksklAUf5NsneIGORtozRVBGGlj2rZuic7xD1F
SeWJxt+mMu4zNqKMfCy1ytanBuaCJz7bEc4z+aNKiIjvpEcl0nhEC7dS7l4SQC6BJRQC50UmdxSi
uyH3Yc0/IsGb1h9p3IbBVgWKkStRWvjyVhCWn6a/CCmvnQqpzsMl1ZZ9sszp6sKVu8YqO6+PtLBs
ve1G4cZHnOpNehFKqe9AtgzQX6XwV7M7j2LtUf/nj7/rS9G9dDXSYBVK7QuhcmmtE5bly0bQiTeB
4uSi7NLbdy2S8uqvqU5kaCQ8dLUmXLAhhXZ2FGOh2aC950VT8OD/wgmjXtXR0tWae9qvBjbz9VCv
HM/AE1vHxQvDGBQXKF23rhA+C5BKAEXJYcsDrybrbwCFU/1eBoH6pwpGO3cCVPUXzC89kxhiBp2s
c7w5hl5Udten1bn70E1XW2bQTTq53V16fitZZMQBfr9XepYp4he+pN+NBRIDuGIzam+WamiU9RYP
CEFNnKOA7W2Gz8yMMwlf42KpJEFgvJ6vKcMt9og8x8XqQdydAHf7paClqkEOPN/JoNF5mb3dllJf
3UytprWBQ1vA2uBMer/UsbSgjwo+D9XlteyMwGhoQlXJIpXaViQ+Eedou54ZHu6OTKNaIoPfyPQ/
6t1pxo+23u/Gm2FsHI/4PGwt7FYG89vsn+tbeIB9QaiQiu0AF31V2HOSdd6En5SVlG3e4G/N1jKB
qYznhDiTveIb8U3vM7GzX86+6fOc9pnr1vv3ltaxVdCSAA1oMTnylVx2ONNq/rhXAkKV60oq4Vgq
xfofq8FiXEFCWvgMgT+V3yM2FWUp8Uv09mfTlfVyFLbgqp9chYXMrwTMzDr0HxERj46A8VUPpue6
wuhF7PLBvKSCw2mr79RnKUWQh3qlqrWy4l6wWizbL0RKHEFlq8ODsoq3TxwySR7jxLlev4nspokU
YNgKZYq+pZ6ZD1EKtAQFZJ14U6P1llXCZDB86tdigejaz8wlKih0BwKeKr+8jPlBn/+D6RVsoyqG
Pv0XD4SGUdEQW/Ye6ffg11sHYUCERmCGmYCkOA/9TcRMHffSPsdPGTXL4Hg/D78ND6ikKg7Ry8Y4
2p8qyrTIC6m25jnZIS/w5Rrvykl67pvpPFDpGK2n5OgABBDE/u+bDLWVoF3dF3nNjZmPU/wcAHqz
VQL1a10/gqF2aIBAyJwd5H7CXb0VIoVojP/qrB6plCvpgKzjsU27zyqxcXCOUeyz0Y24bRHBLa5L
aW0Z4iNhG3bvtPOULqwI8UDIBefy9H5VVHGbAOhAS2F5JHlPh62UfxrqqrJ4gAZ6Ma7vroeVNzLg
RjX4Qcy0N0+AnMIxNzyTrbShekL4EVG/n554u13Ab0EKdpJzjneUHGvgpFq9E5LKLDR6LiHvACL7
DJ4gEDf9DzG5wroArR3yAijsqNTXjmZFEcuNlVzHizz691t5vDlCVvfZ3Zc4GK68X0J26j0m1RVq
xUVJl3a2XFXhXuyfx7gopA1pB07DRkhc/y6Z5Nfhw2//849SELFba9o2cfzOzk6qSL04rWjydDs+
2Qe/U2hCb3VQQRRMmuXmpESmoyNSCmSbwWVWkMpq+6btesJ2oHrAQUatN8vWjvIpyeaQLixLsrBx
mowwHdL0mGly1L6WN8E0jt8nRQ5GZFgFg7F+2EcrTj565vaF6vYtqLHW/L3vxn+zeLc3T+p/XxKb
ul/g4tZpKAxulLMIURTz1CdxRreHBz+ny22Vop22HyikRXfg8bKHD3P+RxnlJdpPdGJcaQntWs5b
qQR2COArx0wnSOCd1Xk0ZiTYub/mvj4DMnwzM6vf2/fSZ09AUbg6nF1Rh47lHS4OIO6qACnWvN0x
bkS7eHqISIOVK/AfFPJk5MjhtcVfYq1oxfLc/0E61vKIbLwJOcEbO9hapPGngJ/XH5sOFc/mTesW
HVC6BwvN/1zWGEeW6kBQEHRH+K9zF0p/ixCFxWpvPlugM6cPrq+enK70ASFzjcI24H4iIxqdARZU
BY74qydQM4CpNj1QVCRy8BkP+BD82P7p79h3GTqzJ8bcODmP39DvFGPslN1hmLqep1y/ITbszhXt
XQmI+BrynzKmiLJCQE4wl44DvFn/iyhnJkt7bhUVDPordJYfMZUeHUP9iZtRM7xiihXASxqZxMCb
Z/KItvTu5h2K751ktNpQAm6ZHLDa7218cHv/Mh7FycPVlpOPDtcgFmXR0IrBLalOu7rMfGqJf3Ty
mIzii0/RAB5DRf4YNZw+xkFXo/iIbNc3RahvTvUv9j+2MYiUQbFUz+cFBbB2QEUzKMrFMdfuleSi
OCQUERBZaLkID3VT6U3DU3GG0DU3KpRoXiQw8gBpbqdXUdXlVNzfvcSPNiFm4mYZ9/lWOzQWCWec
24Bi+jIFhRC8MVHqUyKjnjzABcq/FP0l2VpUeghioRaZEkJT8lmcZANwvwcxSvVUFivMffhi9khT
j3N8QMEcsXG7c+k/O3ITEY+7dadQSC9rb0ry+WvbLwfKrqcAkn3pCg/5Bo2ErGxIcBT5mxkMVe4F
4992A2wbWNLCL25jmCKO1VbGg0vhYdLtN5NyDmxYxjycrIqvafBEWo7Yq+mmjLCIZZfaw1PNUTvK
gdNCzm6OZe/riLiaWL2sR5DNYCpwh5wHq1gJWVzFBGrFqyd0C0eoY/cMdfP91qqtMuN58RnfdT3Q
3Dse00cYJyIqWby958/38qlciRkixofL2fiksItvTQAFAfw2KLhiCzF5ibIzG1aTBxtaubE1mlk8
5aAf600ohL4Hzgz2Qf0WRmudhGUf9SaWId8uX0LM00r/Prt7X4TMJwu6xck6z6Ti0JLvxzQYLprK
4dfDSBK5htZOEdMFc/1Yh8PnQPCCqFtrz22cvsxliBNTMNTQFPmxpDtwxznNCUCZn68vgmrFnNwv
9o35W6Mmwiovt1cZo7mchbn2bsMGrRjZdVVmHbpxoJbb/O3bksVUtkFyCecJ4h+yE3osQ8eOxTLN
N0cUi6L5YWgXxZ1muHrwGTDO9zIimjscp3yVaVWYbYMPcknmUeGlSvZ0zHBVqurE/8g5s7C6TfU/
UBGiAhFOVti3qdD0+p7X9vhcPw2hunfwrtSCGmNy5mXrqdUgiRY5F5rXZkgPxWR3myQCH2UFJ7ua
j+on0SfpuakVCZJitW/1dsV4Q+GvsOi4hVmTlmlGnFsta0wdXSFX7tJutT1+D4yjnkA9UlLZphQ8
gpt0AnlaGupX8AUyYIoW2VzmwGu+TsCFwniu8cCzWF+k/MZQPUKxCpAKfoNv/p2P8etkp/YTuaNI
3ixcOfJQHMPsBH9zZs1pZRGAYmy0/whurlYK4dgAWqsC2g5hMtKZ8MayIk0nQ58xvf045k0ja//w
Hr/dS+3N8lA+iwyA7AQURKeOBkKF88CuVm7vZ4NF3/6nNmo6oqTuRyTL/UOWR6vc8axypACtZcst
YIwVxCNjWLBh5Fs8pk6GQribiBV1SfKfF95Yuzh0oIHEiNOvfFZ6+dlTjk4nvfda1anxC+NJ1Ozg
MxMvVx5CvGV/bTg3ao9bhxtCMoUSzi/GvFRgdKq8I9mD9Ff3Yv/ZmwFUdbiahy5Caa9AQ0Wdm6fe
RjbzrPSmU/pLTrKN8c34BQv73uZWVpu7maDmPcV4a+PpxY2WQFqEwNoJUkSwkiU0gdTaWr0jPegw
VIqcBnVWxxWojVvX4Kr5YC6dlm78Pv5hzocWvE8jUwVsUHUduF7RpVeuFJcJhkRR/LTLDFFSy64s
TUf2itis0RSOBdqiN6XDGEMsUdGIgZWioLQRlIpvFmRWR4rYjB8Ys55FvPtyWlCdH5n2UrO5saqZ
NyZrsVlzkdQ0melLdb2xP9p/T1gxyL4X/Pqc6BwTwpoeHhDUa/cal76xFMIfDFpw+CKYodOm9qdr
tpfi4l7ECFkAuAhnYvQ4Tc3dsZBWHb+6rDu8+4/2pPNy8U1+AkAGPFQRoKtzgRDhq3tMom6ydVyM
B8NAKEYoOooSCl09TDVpiYJbLXV5/NCP+dnStp5KVFi9Jyt6ngSlTh8JMv4F+zYO7i/PNEB47pYK
c4mtXmiLtuGyTV3SpMBBmIWoqC5M1OAYX4LQoWqN2/e7MFn1Yi96gS1uL/CBihd0kY/0fnrFQMYF
/FESzqz0jwMz50QOQ/l7HGQmAgNtT2hk2AgTY9szMq7nscXEvRCisopDaZgEIDRFs8xe069eVeUb
F4Za45Oh/+tCb0X0J1SJb6iuBM0RA23icKNCP5DxU/zgWUKNjwyVh8Rc2fw56OrEJONgo+Yuq49Z
0PAQOIj0rRkLPgovT9ED9RsW7wVM7FtFblrLcjFKJQYF0FtOssHw0uTJ4AVMW7n0SxVmPl6MmWFX
OM12oep12EEzW/8KN5l0ujZURmYHGTDcgE/LJR/xMEz0G8/pZ73MEsR6DZTvS4p+B2vNJkc436ga
PjVa1pa2/BNg2tiRX0f6uymFUs1jkHHF8zX6lJuFYvT+MELPfnfGpYOq22ei6+o1ra6y8nwdMKZP
26dMuS0zRdK3XxDdvnpPiJ5wMoSAV7FED/zQOXQRIv2LB7yRfXvlcDxB2FZHnsdMYKTW4jco+olJ
UY+am448NjL0WzOSkGUyhsptbPmqIGSMdNzC/myUFvHxs33ozX00aTu78ePjHMcd3dn5Z2gkn/n4
aCoGq3hGVFJlKD9a7BjNQ5BxciLM5sikqyAr2c40TsZqGd/MPVVcY+btMhOMg/E3UyQaVhE1eqM6
O4nv4s6F4RzehAHxICKR9tnMT58/gvwKwkS66bDDD9AulTSJBsPK4eHi6kha1+LPfDlA73Qo8I3e
HEpzlPPbe5Nzs74IPfHARUWDle6Y1dqxUMT9WmZ9FAEHOfctHHR58Zs8CXCutqyGySW32m6kHk2L
0hArWLc6YpEPzp3jx/rNEcV7Zv2fjWOmlLjd3jfITqYcc8naMY5JjQl+HY8ywaK3xtm8FrbUR8LI
njZQ3ErfI5MDBoKZAl6HFqxTJ3LPOMGqt8w9oNpTwf//mydccOKrUBZRxYSBYZSyJr0tyKN5R8IP
QbsZesHC1WVD1/ybXUwu/AWMJd6ADvj8TytFtVsuuz681m9vlJmh7Rcu/qfFDabFZPCj37vnr8xo
DgBgf7cKl04FrW24SgC7O9ilJZeBvB/G/ll8glalY4GNr1C60aepIXH7T/JiPD/B1kVEzCbeMHWn
w6GM+KONC1sgWTOv13K4JVJltRFdYIwptIupCtlki168Soop2obwRLtzczR9Qddc/5ZLUSaqQI+G
VNrgHkwZAllfvk9RyJ58jwoOodlYMJ1+EkRt4MEjK02r1Gw32LTUI+CTAZ5aL4/xfrX8TMYx+PgF
mX1su/xNmm8/gXMoNhDy0Sk9u1wcTDHT53zUvrI6dXvOk8Lo0EJV1+1M5ccAhsOQv5Y+e9O6hvY3
TxpHpwMLtSGC53pjalfnNI8gH0Fxwk5oGm+VUgJPp0i310npOh+w5G9hFe9l/hbQvxPgfs9DCo5a
x6vn69iBRhGx3GBPijK5r9/+Figa31t+B2WFKJhFYj7Y0zeu5AmygaPedRJ7fOFB8D6ZwtfDzC8E
j4FG/g20bL0f215Shg2H05HDbcpdCSu4x1RLYJ1LqpbSfQzk/sxwuEV32ByDQg22K41leUP2yk0b
zx0obUZBwWB19JKje3CAioGEkzBTLsXHhIkoXDcqLBPgCY0Hc76zOWve5PhjWUB6i1YC7799oQHB
PYwDK8omhbrOKODTf7/kDKOUiNiLEpPDr3wyqy8gGzz5M9EKT7KmZYMMwJpv9VVPybyYKpqexgXq
ObLtGMTZUySZPFmXg/1dUQ4Ii8PcPklkQe4gloRb6ZtO1A8s8hX0EsVDtnDDN4Jwv3hY4BCc3h+Y
/2SZFBdEkNjB27roxJsYC4N8Z84lLwsQrTkOkneP2zrPTf9OTEoj08BzRnv4OsfWqi2Lh4ce4IY1
TfRuLFxjdWyicKWsAHWbBkKfInGJAVeWHHZiLYSOhRIl8ek34UlCe21pGeiYGfqzloEyCygWlSr5
D3DIRTEzG6T8QY4+d0vGCwqOlhhU4oqwlZ+TgLvwxihu3SkuOLGI9R1eGX74laYghqJinnkOw/fg
kNfUd9mE1lenZ5Osa96BuqM1Es04yVlNPMDsr4V9Qwxu8OmjWZVb/30lJV4CoAu0wLJrYE1ASYUT
zi8S8BjsuIcjuUiiIWvW9hGu7V6SJtVObFGBPE8jXWysklNkhc4zT9PoeC2Jk3MkP+xEFOuheh+n
Z3QfOvzn+FMCGSo9FCdEyTqt4R7xH6pd77wp11/tpkX8u2bvoFFpFL/m3DyjLHpkI1yxK1PPENB1
lFx3fA0/fV7tD0OAZy4823v56a0yibYL/5S57Aw8HSvEmFQjZwX3jkFqR00WvQ64mJzPFOWZeaUQ
XgWfpvBN54tkYMC75V0r4ShY5X1BHcUceK+8GtigqJ6O+IL2SeLbaYJRf6MuFVCzr2WNfqQ72QDq
qsSVuQZDMu+U8JfkBBOPp4rEvasOKcRYBEnQd91Q6fIafjDscgepPiWptQJ9Gm527LhAtXvD9C22
3UAVxDwSUytgBtjT9wnbR4lHn9YbVGB9DEPzbvIVgXQaKXkmAklx7hBSjRFp/N3+SOhIAQ/72Nsj
CpcOwTvwZmgYYYxlReRIQAmPAqfmOCCqcmZzxgpmHr6BM5+9Xqg2qk2U79kmkT0KlP0yNhWL8gHo
67l3a1rNGMpLqb0k9gomDW7H898m80eqNOLdYezT1IkKqjsbLvobUg7yGR2uT+2ml3tLTMzd59FN
sglZzQxXziydxeF7IILVwCdk542oZSrnRC1jdrtux+ag0Ba1pHOrzbpUPh1IJn2kjqyH/0nwG8sK
9ZeT5LjxWXogGc2LPoXIn4NlDHGvucNqGrrABTdETagQ0n77cxg08dGRM3y4jZeCQiOAhXpbn7E8
MVnlGAW2ujcq/VIlwquZPh8hWZxOBQxHJdEDBTiB55DSQJ9JGUV+uKzoA3OFjVBy1pUoqKds/jAH
2EnkA9H3qx6fY/hIJJIOCQscQPSP8C7i5UTXCdMfNssfVp2Epsvq4Hdhe25WRTf0ydswoqoE2gxQ
9jY5BYjbTUexlTS8T26C1qd4lD4rty1mN5yRl69/Us+ykxX3uJa/+Y+czuCrv/xwxEldMx8eLNqT
EJ2WdBmsK/2ZL4WVee+XUZpdmmj0+xROmjZMcyrNNmncuCzTvgHdS/yg02qBTiHFGorrle6Xa99V
CmO3bieNVlkoqq9SJrDKuPxtPrBOK2MpZoi7kCF5vMXoPs2MdCu3nYtnJHXa98KHQAu0p1TQ1NPF
+1c3rVpnezWjoNfN3yLDkBrHT/AEn0FrjwJLNCjNUEc+wdGDZQkE1IMjGzYIpfSxMSzQtT3R3M+Q
sM1rI2tGH8pheUo1TdhwatUjH0Nz20DnB0c3209pGdLToHN0DQtU5BpiDfkq9pFD/ZHGX9n+Ov8W
i8V/mhWg3kuFSytGoieqilydc3iwgtwDz68d4zYQnFcW3oxTQyzqjiwOrf5/Kl7tHYebUGcRGw8L
x8vd+BxAFvG7Jf6MztgI3gVfV7DUUXCikk0WdGI2sE3IuhlClPM/ry4Ug9Y3g4nUXbKKb9TjDuTl
RQ/xOtLbXz4g11Ywhz6/IDkCDYOTM4w2kuKmRbHYv5Nd6/zdCeaOBCn6srqeKAg7kBdF5iRbxROh
mW6zLVX7vwq/mgRhGuWZZG89Q495rl1BAvh4kH+5NGIaLIvvxYRBYERsvd2oE7N5b7j5/G4ndo+G
gJe85utStwBXKJ0wq7+cRr6fLHwtZv50lssEyfSVvefLo8IYWcYp55YlvSRcpksI3SZswP88W8OJ
/vO0Mys4LoWZo18Um79e8T6Ia1sZd2HPYNSYCPpqM1KG341Ehts54g1pk/BmYoaUdEKzz84Ez/KN
nTESqLGg56dr1GdjI8IHKlOIwo0zFf91wlzg71LPMZPqWZ9s0Ka+qpmGAFr+vXfz130hqQ5B3Wr8
ULS+GoRGByP4mQ/EHME0YK453GCdgx0qlC4sQ8YSL1VIeiynhqAm8RaCCYyJhjDjSelRdsru5pLC
TsL8v3/Tzja7db0NSNA5ajRxNZrFc3R4SxHNju+6gQK+ul07vJ6ZFGjJOqIb3lJ5xq30XhxvoHVX
vaskmljaXjoNwhb88vMQsT8SsI/5xDrWNlRtRE858rFxar1ses9hBSLLI241K8kn+j/c6ffqWmR0
rxTfetYJ/X/trMIjpE9SC4ti1laafMrSxoCFFqYWiOqODQhB8r7eOM3/U+9yHEICx3pDO03MkgR9
Ep8jkmifsU6Ur9a2OFF6bSqJuTRK/nddZZ83YLw4d+eN4+JKoutEeYktZ1CyxDc9p1cg3Y+mwnDn
ocTOpXw/I8s7YaqfdL5iVvKF23qVp2YkzG6hpin0Yt8KgM72O29d2hMaY7M+ifipC8gbRTJeSYS0
4dEAA16QgXWqHLRseJw3qpJPm5wthll1kldVs3mPeQoK7T/VfLiN+k8fTZp6KbYb5Hz4xaR6eg3l
3JABDhaxGmSgfFhVuIJLEpBn8Ac0+egBr3LDp+Fq/mANPgZBJJIuWZMJq/1ys5XgzfAxEXw/b0qs
H1k6sYvMcRcbTbseWPAZMHhzGxeb0bzDJ56M7ajyCDOppt2kQ/t9wJEtoJ4pC2X1uRPW7AfC5OcQ
XgTAAxd/aHnL/krNpnPQATy5+LOQpcYU0xFosy3LHT/NV3ZB2j8NTqg9+n2iP0xnCTBfKt2ZpibJ
H/kTAtU7TNOKje53OXKxv+oB3G8rVQ+L01gc9iPC9No0wx06EVmc5BzTXBDHnE6VLuDwpIrL1850
EsAgxAXRxzAgFhl5+mtZGoi+OU8G+mBDud2gv3FQ5XeaTYE3aCJvC3Ai2o/26NqW7YCYatXQ0wbh
0X6L9KHhtubnJRpjoY4BOAAvDh6uIiiqZGF4Vo7Qfitz0BFiy3QtkhutEjAfpwnHJYD2VQ7mL8IM
VV8SewmRzeNS7eUl1pXCU4rEk18dUtMUcOrOg+qLLt12UBf3J90q5BZi0sNVZGKYOXgktqhNtsz4
TGlGste8O+HeHaYqNUm4xRFB+B4ylUiHS0bjJr4PmKnJDCTvmCK1gDTylfD5D4gj6X5sI8+B6dWv
tidCLw2nzb8VL7pEiO3MIv4P0OTg8YCHtoJILvtubzjHXtI5Bl/LPC7iv8PrSUL/MRQlI7VLQQYY
PAZ3fCeQu2T1OwsT1AzKesFS8eaTjTNHR8NbKSbQs0zjY3WObQ31M5GBJpfGAwR0TV8Y+HeB4JpI
N5nTQQUnq0tcfN4KRaM5zYjPgUeCiF+kd2Ky+mAiof1nxcC69ZIo3i76be+VY0S73y1/HpL6AR6s
oIQFBFmDeCwINPLw5dOjdzmfSkrvWyDuNm/sVRddnc3H9AGswLjdcH5jQaYmC0P7YwGtnjjdcYQk
ftPc1OaQuSW+uzBPofDUOTjNqITzpGwRHsAqe2WeNrQDvHfhP3qd6N5u1+ieJwdMf89+XiDJKsRB
f2AAiH8uu2nmMVMqZY9RJrVPnsK0cKSQ0R8VpdNV3hDEirBoikcnQjA8V0UuChTqYUOQ204mEIYp
lKFyWu5wJAW1zB266H6Ys2iidnJuxmW0IXabaSgts9qhD4kDT96enHSos3vnNtR5CNbLQVrNf7o4
eHNhHXIT6FqVxHleyvqMt2Mrhu7C/YBKw6iXBcrVJ2MSkaW/Ryb2KckmjeySrPdbbLvwMt9ag1mB
l/0PzjevGbdQCmJM6TqHxT6N0vmUIjmEBCdg3IKxt1s2WvdPPzs95JnWrBlhtMKLTopa6P4c6qY/
G8iPCAd3oNY3MUUyB8IMaA0ZF6pGosxmvQvAqIe+4Ks3m+zptjp8NK2drLSH/IqFxH9TT7DW5EeD
Ro2ByvpLJzq30r2EsZ/yulbMW2VApn+oXWekgrOt5gwNJXa2VcoI8r4SvLzec2UaB5ewNROp1dME
QCPOmSTM1i8NOJ1ikBN8Ww6igpufSPkl04XniQxn/oIpFifa99cdM82MhIB/0lkCaQvCqdECzzL5
R1WAmgm7Hcv6QPq8z4t0i4Wf5KjO5kRs+os1A2t8iCynBqp6KaQVWwE3rVaFkh8nB/zyQi8KGuRE
AbTcX91ynenGFGLNdpEY0q4kFcI//gXfJgZ7vDW/BesDI1EcgX2/GBBr0dKZ546eiRVleF5PnuHB
fH2rZ2abUWHd8Bl2jKcbbRe9iC8Cv5fS1+fW6cOE97H71kwsn4TCtc8YIDYanNouyBsOqMV3a9pB
yJqxZWkVMV6+s2hTaey406kQRFfnth5x5RoD5XuiSZZtvBQm3Jw+FdgMfgCebfXXqSpsFqn7MuZz
fz9zESgyRbCcrsAX5RIaInJ1l1DzpUOGXt2qOov96druuPAlvLkhwvdTbgJ1pAWAki87rquApaZG
dMe9fDVyd+Fac8fI/q9BBp6gEbz7Xljn9IWijfYJnDGSp1LmPudZsRb2XZvV/1gl2MJ8oDEkvk+h
5kj1ewkhacmY6mQu+FUYx5vJVNQNWhKQn0pc9A1APssLrzFImtE+o+H6GOoDHz2+TqW1mgpUWK8m
M3Bcl9uzfUO9pK2KxElX250QYGLwTVjFCWfZxy0M5xnztgr5RMOdRwgFbLFaIE6XryUqKVbjosmf
Ozkz1p/vaMaPfF4nmHD45cAH4s0w6vU2M0jy/HwSBD8+QhjaSoBYY9YCB0raJWemFKvulSdFBr6F
q4w/UXwWdYmvWt8KwHEqsRlPxi3G0AYogT6qlaq4+oITstlayu1+GgrI5bo0nEzSvl5QJ+sPxCxx
ImQDv4ZC/wihpGyP0mKmqTL5qc2LnF5H3h5NtLHcduyHkWKzHjdgd7ORcweLVHXLNfxnyAYhwb0B
On/EZq6Vqda6SZzTLcS49mRO2TcysG2AHimfHiPwTlcBWPoVJFjR/VqqPulrIXMN1F4sjtLDncDl
dIgi7hfXNOc8tttkYg+MN6l+2RIGZ0semL7tE0jCyZt78SNT5r77v4PSoF8A/Wj6PTBAPH86Ei5e
5qCwT+mkpWr1TMeDyjrRkXmWux82+UFsHINxZiV5uXj6snZ5niX3ayA02CfIORGt1Z/YERftK+zy
nmtdZUTvJZCJeULVXSYb7XKcS3S0gGg2e8dqOrYODMb8KDKAM00tjEZcK279CchEkJBRjnRPlev0
R/fks0y6Jazlha87XSNmkbok0e8YHHCBxpyVXxIEHAUeOyrYjS0BMWDpC8sEfdErloPcjoW9H8yf
QUCWdhLZX83TJ+Vqo99tuflXBLuHOuOG3iQOuOgdMcqlkPs3AFuYasnRvZIInTF91KSrKNClQBIQ
2y30Wr6KcpaUrPrN7iP/7jkPeu6Z9CnANXGJGtHDcSBMqhO/wF+KKTo8gtekS/HdhSR6SBjZshiE
O2dGkCpyJ3Uf5z9Q6SLHHwPfFLPfouII53Oi+kdNtpYVY/qGvLviyAmnXczKuVj4vxLbnrZdOAIB
rSLqrGN/zvI74lA7uPJPmF+bL8JULAXUYDgx3S4B9Doxti8O1KpZFtyXY4Yr4TYdiEfp4wrtbNEb
utaQSB96/b18z08gT2vzTTsooSCTdmXBkdN8B3u33GCpFED5LVRQj900gAFribiF/MGFOLkALl3/
rA7xkO+thA0rEZVmZOeRjD9adoktRpXiVsvE4/uz/W5OpK47/hEjPuKpmq95ijW+EcoCu9woV0CL
yW83Yjvxe9K+mcDb4OrokB7ue81leCVUL6eniEMF1cA/tVvG9ekKSpuFQJT/dgl+7v7DXvlQzjbM
voztuXm7AM+PZZq+fUR/A0FPsjpxfo8vBSu0MrNIUOmVyztX4HAlcXiM9wkDhTujpm5h22+iRjlJ
/Lhcw47SRUr1kW02brPwEV6JB884yUzOaowE8zxGiU46LfgJrPOECls5PVy9vfXaGLdX1K4yakuZ
Q8Mqu39XuGPlfTkq6cMfoJUPyAmy9TU8SmrDwmt1ljKiOt1KdsZ2XlZn0CX9fy3xcp9gDWZHMO5+
retDadLQP0J3b7db0eyr/5qbkpoxWKIFFjTtjUZbZdQDHg59sSjg74OPYBRuAEEx0YntBlCm/OUF
AP5R7cGKnwYsifqk9YsodLa0k1IwX0g5/TOTtaBccsv+Ao+2HNtb1Ou1qhfKGdg+0MGextyXhYSV
4JW5bQKQkIWIH2mgTuoL67sIVSzIwilEbw/6dITRxfHCJNi3wFEP1j+KOsxL0nDyJw7pbVNf5xqO
PyF2j1Db6AJ/rUY3hzHDbuUt5RtONy0o2++UBjCFwNvitEz2bPQufQOWUWKtD48BaUQwSNJKtnyW
iRrVl2KySUwbnbPSo0kmmGli9Qk6H6eDqqpjC4S93iUAsjv50kX84gCihdhZL/W+Sw7Vh4FZBdy6
7EtXFApAw6qFxvteG6PuqWl2gCp3txi1tjS6H2qwPUFu5yFtj+Gc1iKMyYBeDNquMKjZMBkHWYjg
/yx6MjxRE2cDL4bk2Stcdx0BYkq7dxRjxRcg8fRRgc50akZknjfJ1lmZU4PhDR+bEuc/3v/bSVAK
ej9diOP+CBwGTuwxeYaKbhNWojaGMjr8R6AySm88D9HqTFduQXg+9jvE9ce+N9km22U8iDo9vJnA
PjPgW8lXgnVUkPT1RA/6e4XLDh9hU3vA/n4TPE3H0lkEIHRKECaEtE//VD8pnCktOrbueKdQSsAZ
p7jWWctQ0cCBBjNLHADZRE4LmuAclslaAfyUVNJAfb9URgqsrgyTDOkiqFLkaRaJUcgrtzLDJ+zi
DqYO4UvoIiLR1oQ+nf0XX1CRPwab0OJjJR09y2q8RlIgbTrUoOMc7uhZK1jlJGI+zTy/1FA9N5Dm
qOYcvysBIfGqI5yqg2QItmlp4kQtGSOh0YWdwcUh9DVgyQHMuprBsTs12ZwCM9V6DZoXjw6e3+q6
wxigJlRcnWBglHqQBJHFiCto1zuLsrfWEGB//8TyBTTVITEvqYxpjsU3x3KCYBmFrOXy8gWS4rtI
vWhxrSnrIPFqOHNsCbbz+AEFyIwe6yK8EefbK+LrWSQ2vrVZXJeROUlq3GxQgR1oHJBX/mH7dHIn
IeV7x7Qmf5+fwcmfjrE6xw3OZ3IWXZ7LjRjvFROGDlIhsne0Uxj5PrETAAxie6a3SzR6hbVupKM8
38yXMlnqkj+VrCOys7qExc6pZ19AspHJox7dt8ROgfGZsWWfwxe/g18ZKvabhGASVVbRpt+lvU4h
Kv/PsBDy5h18Fb+1xq6P5iUPRr6d9Rl1ndTEAvB+QTJpWV4cltW+63fMSnRVsJtkJm/uGlwvNE0p
vFHiBWSU7DTjqgX1T7hMBpHu55b9tbxdW6ZvYKl92urrVnRWIX4hrc7oTbhqq+jMvvW+1emNm7Hv
R3Yr9umrM96LbH8moYzxkXdG03IGlp2zjcGuXo+rX16rNThaVfczlscnYy2deY3Vr9JrbMxtyQl5
S56xbjYJdnWNwG22HGKA2ZZRDEjTiLONGGodGqAIMDzuSeCnm8tY8x8Mw5VYwwR2TSy0mk8z/MmI
3QtGT9gbgmR0sGe+WjvD1zhTZ/8v4GhtZQVX1T2xBBO/WAyqwD+kYCeCENA/m0Wluk1whRTDYUo4
XSkmQYDfSTHNiAHJ3/o3K9358lUjrUXhQPnTjl1dYxyHtOc/9cZpduGnBOtpay4RF9JMBW+8dAmq
tzz1+HWOD98UEAYiXKxBE2kF8C03bsOavN4ZtKeI9RXzizpUvB+2dSe6192+oF9rXDJ1pZpyj3QG
C3M7S2QXtA6V5MA2fy/H2P1ABBnWFWk3PhvwHBVPJrAqfXN80gJyYm0nWdHjPjXlHG38e2Tk1Ush
NiO0iggsBabwHi8QFIHnVMHUWwmFtyOtlB9DAM0j2cYL+BpwPv3q9idr6Yzz0sJ4AmrEcNM0rgej
VCLVnkt6v0lFyAsKegX7elc0VvI/WjlEfjRPwIKG+7JgK9pesLzaQ37BsdMsFj494Fa0/cMF6y9s
jxqOemXsPbqPEvhTv+zKCISAPzHyCKjjPH8hJQd36Ot3Rf0/I6egdMHEYbrO9T1rvOuAFyAJGI3T
BxWZwm2tBN8JGz8AWIvsQhJRsfyy6DNvOqgraYdm5kf21SzFTJhHlQOQKoLF0Qg0TXzB4v8u9QQc
gjHxCm+gL6thlIBuDQIUAX4a+qrOedA8BQAesqduwAPUvjLT1tgSpkPWLX3WS2OfTu5BwfNVXnza
CdTQzgXYfx3D3kxdmnXReHVMYCjnpLnuqZ0PfPwyiwkKz1wwOaHcnObRHJh5nYuWX+xgS5mvtDpE
umiXZm71tS3M09OBPgYH6AsWTtOAc8w/OnzIN7ugU0Q0bZy9Syo0oYgwavTiwZepw4wwseRzfo3x
QfIRvofwwBWC1Q/pSv+rHmhFtzbz5um55UMddGqc8c6l2c9yUnR4/ApMFXq3jkowSCTi5cua+TZ/
YAbV+gjPFTJQEBueaURr6gvnGAvTHcwCyUALvaPmYp9BLzki4EFwJ47XEPYkg7xGPdb8HXec6K0n
Bo4yFHumCy7hrD/7bRNquWNbpmONqMyOr6tDj7H4BaSo4tTfDMqAk7ij3zeCrRcjnOwQZ2tBqjFx
pJwpV+8ceHg6uWnJeBXsBrnKQfu97RHuXaC47kgyHMww3KrDcutys1t9W/I8yQJOZhTMoSedy6SB
wkm/WmgSyc5HK9fATUU3udNwDH3I911exkQhFVnbaogdVPu67M70CnPHsoCP4/p290fNDg6KYY2K
ytu0oojV+IRflOJElBmp2K63+GERXC0XkMjUrXvojXG6cOUUZTcEf+Goyocpp41ykVH8IHI1JcH3
5MiwjUL+u2ZqKZ0SS5lv6Yc2Bk8TXdPlYTLh0lBVofi9KNpRZMbOXtY9jtKnRht9T4GVuAybzmyR
253OQo2bBNXp6MjU94vdfRpgq2c8HrP0qsk7o/CaoWiFpvrX/2RHlYKnqHHs+4aUBXnc/hXK4T/G
qOVEb/v6G20uMHCVs1Lf+hLPcykj4NC7nCpdFC1xqq3ehLxw+VFhIeWqdChSai6qhrzRj4VVhlHs
I/l0l9atcuMC8ezbp2PYsnoA5PWliJ10oguPotfLkSp4UBV7W4+ja1e4gKN4FHwalG0LBH64dCoB
6s+Kb6UGH2YEUUit3BEH7gQ+CB1TYTHEfdgaUQtgQFnUdsc+0Tz1ZRiJRQHU0DtJXtinN3C3IRdx
a1F77+w8YZakGydKoIlIm53qRTwFVFIt/+sj4Z2D9nAtsJ5iw/L/9ZE/M/voLRQLTXRjlkHuhh+S
O147FUGTXxdsUbCRjKksAlmLoSJO1ODBaI0WZPZmbDeqDIpVvCN0Qa9lajnwclwDAUfhVDmwuNeu
zZNnhTb5UPRqkpL23LvbQ0SIol1av576hyzCUHZSZrdlgFWkCHhck14Fw3WO7htT6gLJCdizdn5O
CDhAVrkSi7lu2uhOR0GC4mxW+KefuRTSL6u71vdu0Lp7US3zlqyFEtCHMhna9QwereBH0yOTjDOS
Wf7BD1+h2ZdDNtu64O/yrwI++35GLFKE0wozTd8iKg4RkbNBYsJtp6zKrSkClFfYt3w60o9KpLRw
dH4am7mU9x31ZbuyIQtHciPkTgOKKSrOtcRwOtRWRwOiPS+xOYScRDUVEKacHfzLFk2WOPv8RIjH
RC61PsE0aLrqCjyCZYN5ghoQES/JYjlxOQ+N6cYFLNwuM1K53udwO8uvSff5xNUsc4AztQWEawOv
TP1lnIHHwfZmDKyEDRtBZYON+pGOtC6mOXbPm36YrIyo3gvyvXIcDrFu0amGwkUYYRqBhQIzdP5O
av9Imh9l5rCzSXFI/U1fKbKlGL2TVol0rGVmrbJUhJjrvUCuzZNCzYzGJcvHQcqkk/+6CYiE6zzZ
XmWJmtysUJADFGBekxeDJOH6Xo9avxONmCZc5LxDxq1nBvMjV+bfW0zV86c3QZXGsGtk0HafvMyU
01Iu1QhgKFzNh3jSySappF/7ckLX/UX/IPYVInQnaJQvMuk+lexb+sGwSGgkPVnDlU5JW3WGfVTk
l4naiObex1ZW4fJnZuRyBZTZkPMY+/tAFt3ml8fcyps0IZtdLksDymxAeTqWqcLSxIofrZQk6gju
SK3SMC5jgw38iIwkNlucG4He4QT1IkBvmEV1MD4+nX8RWMxB35n+yL3ICjWB3GYn36N1X3xryBlJ
Vx92pSjI1iRwHmjAewzaJY8DFpo6EDbsNkoJwwB0wZSj9iYyPAFdN1YPElfIjhmVBA6il3SNAYvK
MSnby978txWxlw98g3GRb86QP6yIuTNvvQub8tevot5HvReoxOzRk1AXjbFTIAr7IH5bN21TYBLT
kqgaFtOB0x92lp4pj0ZseJnl1pG8x2D+EvhYxcLAs6E9lZWxMkc3Q2324NvfPbaFqF9cUwK8urgd
zjJttNi3ioq3FhhO0i68t7gva1hgyZxPvMouOtn7dx1iUd/NFYekCfzfworr4I85X2iXDmpBk7mx
/tNG4juEe74+mU9KdzNyb4IEqd4Upmp4CtSuWT11Cv6QAEGZhdAd5RrW/4DH4mmY0D+XiRQ4Gtmd
e+yjqUIQk6ilecuVkD5gSiEdS9lI4XxMD1W2FY5gJWBedDoo0HwyuYzguAkfb6Rvu6aAQgymuJHA
RiLKWx94x13/i1a0CBPYEGE4S2HDCAL3Kps5t3M86TM3PLMpb9AfsocEB5+xoEFbWO0g0Yddsn7K
JSPL0KxJaKPIga0LsS+6GSsflv7Z5vw8yp5tfkracuH0Ur31UZ8WU9b415LOnhmXMgdhZ39nw9JH
8r/mgRSY7k9Teq22AG+GR+WQcs/d1dJJ5w50Tfnz0CTbynN0ZUSnx0IqJgyl8ApE6MGySqJwxCrN
DqmZ5NPAf+dGVt/luQBnJkalCkLcKp2RrE5pGLe7pn05/oFoMco/BebEbkJdxHxgn9QhPsU2oMko
C/uZ5L7KdclSlsTHK/MkW3Kag9QhIUP5Imq9M6sz7/BBskZ2BCN5x4vhgUBIaqp8tVDK3NDmEatK
3bboBLm6O4N9WXO0iaZvFJp3cogdZG73MCcYYlYFnUzU4p37M6gu6PDpj6iiy9QxKJNP5nea+GIm
u0/juhW5BrLS9qcpngCzK4qfUaS9Ike9wnP9xWq+xNjmOF9j9HGxwA3FXPnLiVcaCJJfdDhwJNj5
xWs9VD1sfp2brmgZxl0yGOUMU3pOvAHy4Zk6IyA2i6sh0jEqasvzeSWnBt+jQimSXK+ynB8a0U5b
JQ5GkSMOlLAoDh3Sx+ZoMKHLTrSW2hBmP4xwdGPWZxywwTDxd/KJTqJiQh0C5tmACsz/k+zuck7b
S4z+98uqs3tW1JkQGhlugKimHNXaHpA4il05O7H4OsESsG/Hx9ErOhCByYuGm+H4ZRCy8voWq2in
OkKtgoX2apO3KOoDgRKXR8dljKMD59j0JcPc4S1sn70QK2UpUc2KxQbqzNtNVTtrwmPyjomPR8tD
RbrI9m7IqD8igPBSgbnWEX6FfByTCWjywFQ/gG6aVMl5vsWGf/8vrBltjgxaRfoHssVqB3b6cG6n
79zE9sOA+ReMMnn7VlnR7HSO3qLiaVh+iSMZHDCKip2TgiJxlGnGappepdoLAa/NLAVDOpDt7DOM
WkIBuu2DEFpnlnWm29KBtV3lI79u88KjGDa/yRE1XF0T2UY7NCUg+hKd5pRNHX/mq63VK/7Xu6LZ
20VkmaUf/ezmnO7Slr9xDAjC3UEzck6YcgGdQaoiNuaAgd8mFMwq7O9Hz8VypMuf6V0xa1xSff78
1fk/jHwM1NKq9wRaHl0nq1MBs02Qs633DKEes5dTKpJqOa9fMhUieuBl6JPITw6RL8PC3Jaz8ePt
KlWa26nvA8O9dA6WJa/YywXuXtcmq9nIB5QLnHCZ4BJSIoAvZup3OuBoJ5hDQAY5lljPOnNgYrgl
dSX8RDxQOmf3jf1CfuleYlTMXgros3qLkvCSvd8hMRrYDEvNSFcp0yRfBeNdLLWEE8+jwc7T0oj/
9dtxoLs4ORdob+5ZtiXFJ/5kcSInrwrYciKq3qEIB34eVtJfk4OW0Eub9/38NKvkJSzq/VzH3RTo
RVdrcs2rVcDMtg43MFK5JbJznubjJfqD2hgF/yuO9rs46xdEIhCvcSAq7amxsvYSyIZWwyFhjpzX
fHeKD9k8toR6xK3uiRPwxjUfDY2khyvObdeVXPaY2oUDvIqVM/5q1TzOsOyA4OzQuBINWrB3Po/Y
A5PklhaNh4NHa1p/ftgRHuEWdmreyniH5aSaPjqKth943rMrCPhI9Gyy/5IsKeWH4iTLi3Rt4AG0
NI6AxUfeAUPKjxdaUO+tsP2of5djz0JuTSV+iFLYTT+DuxNCUSvhvQc3NdibYjmrbJN+jh65sXIh
YqrG2Irr2Hy+t5ZmI4tIqOAUuFKpvOfopnvb1HltYYTsqAgta6D7TsJez/75zbZWMfP4+rzCS/m6
8p6SVh8+Gt0iCrUT1ZGlTyBtZsmaV7xoUusl2Yy+n3W79KxXEd9GFhFuxDChTjIkXB6DD14xPJsS
WHyR3mkEe2MBx5K8Cl7zoBjt+XiJq5Y9iBRR2bhLng3DD5Gli7P7WdeoE0bTP3RZTyvziSsCJSoZ
nF/4bY3VCXso5cnV4insog13psju2XTBhZdJYoODIgtkGeg4cTtZJaShgYjvpaoia1/zBXia1DZL
QHpwJSi/4qosbo2IjmdPls73BbWvreAwlru2oZpOwH2a1OHh+CAFlP+AeaqMveRuee6QRFPRA0KX
FwqCDAQ7K8jbPfmoyNqoeOf/8N1uSDYkg/uz+3upRFEKWrtFy2q7EpBnVjG9242reFd2W+dHq+f1
rPxdr5gZ9lT+t95Tigtpc40UdxY0dTSaju7WrE6NeTDsoEmTMfrZF+K2AIDItkrYbvjrAfhDzl7C
Ph2M1uoh7KF/5FulflBkG0vjb59QOFoLvm+uUfsT26BhR1BqvOKOdTYM6C8WYEHxgIsC7aT9C5xr
gty5rPEtXtAk1ZZDufS9V7fFU93p6+k2cFLUXTwFbl3iOv/75Fked639zaTNbrFYqUZlS5PWhb/B
7Se2pFMyjaWjCKsPp/chwSxI0hXYxeMcGZYPP4qbzVeI4i05LMcFpmqRqbQRvkTtXiprmFE4jfZW
fG7tQtf8KXFM7bqQ98qGu3kqYVfOIcsQpKxBMVc3R7VGyFoWSsg0MnpJ/Fh8jYni3xXPGpDOTHUp
f5EoxMJJ6Pcah1vL67i/8hOKPV/+xFYc2RqahzWPtVKcLtB6cu4x2TWRCrTTw3sHschIQ55QeU2x
KKg9JLprUqgt/xwKw6GtMOaW6iUh77AwD88YxRHmoj0MRzCAcFIHiEl6OwuuojJW9+KywCryYTs6
8GA2oKhOMcvU7m49eBXXA0wYei9P8gi4g9rlcbTnXx8AgdyII2tgpJgeyBOVvQDbhrRaosK/cTne
kZhszUk9T1mOPjioEZK8l4ZMtFMeEzgf6ULT7x7NYJT0KtQWWTbUmT8wqag4LgxoP/oiWt+0jKMh
esje+r4r9wma97nMdtb8w8GJVaiJZ93HIcw7X53oC8G3GUyeCF3rprqagp95qQnmdL8VfqtagXXK
xaqV8fXoZd8wCNQ0rkKofDm2SkL/+ZzcPcWbqKdgrjX6jg8KqK5ZIHzSi+a5ooYPcMq11/BmArEf
xLinoolOk4+6u3Sulu7Xz44cA3PdnDiDggECjkN+VJkRej863RIkBv+0en3ayACsvOratjPDvRuu
HQ0V6riI+F/DVlqN7IkhDwfinS8bYeh5MND1PSwed4MWygTIL2XkDFeLQ5T42lJGtjWciYpXOFBE
GnOj7iWr74Ov9jyJyHEiU9UfZKMR8MkKL+EHMOwprrLivHWOC/Ttep2hq9VO/R+Syx3NhqcSbAbS
tDUqI5CHX76M4mf852ZU4CO9upcA8Euft+vI324BR4HtVPdfdY3Wa2nct7xyrlZu1F7RGFzUmMeD
lz4KV8ZNAwrLo8EJDCYR9UdfwokoLaiKBEJRIGlVnxhCyWGrnNk8MPStmSRD7pG+OP0I4ht39nHa
YfZ4fYcrKD1Cp8lixoIg1PSyjheY0eXGIDk+Ua/OZY4x2xha7rwFmPg3M2zaLCExqnxVezETdZXL
k85B5jUX1dCWrLyhxPK9XXxEyVqGDt39UEX9ilvIG91jTY6gBcpGT82jizKSOJjHU1VqfG/vpfLm
7obQrtGHZk9WyXgcY6ctiO14ky61k6x0UypqfX3g+WN1fDHceyavoXksbBSEM1yZE6p6jGPjKvcY
XW0sHH49Xme5MvvTDWla3/xi1+Xp54JD0674btDpVg0+t26jgvI2Em+S5PrtVhCnMfPu9812rf2L
Lif5wsER8x+Qx6kia9hwIBLq30f1M24OIZRRQEbq8um75U4jw7Rc5CPpVrHE4zpYt92t1cTA35Qm
cTwzOE0/xOoM+ShMfg90XCZI0IC7fOvewETdUIOShaWF8lMPSDMV6ZKLNdrvrn6aI5rkSfmA/Olk
lYa4dPdWNWyLPXcYIKFyNIEW7wjUxq9Qall39lau59Nbx7F6EDNMX7DltFOmE9M5bm4WfH1snEnZ
rqLFYqp2l29snJ754YHZ2Ft8pfy4dvYzQ7Z29MrozGP8lfWqCe53TsJR/CTkq0zvPaSPOJOt9CXE
Lpf4WHXksUAJ74iYt2ijCY+0JurfxLMxRSH4RYntjF+sjo1dQx70zbWS11epbe7xCzNRotAVbszf
mEGmPykZm2d+XjQEZi5gPmMV//l1FzEjAepezvwovD8CZwH1JVUSuiEL4Lqk7S6JLykSvaksUR0Y
2zQ+mBLiPvUrzN5DrIRJeDovVSF6nESQHg4EtlxyqYgAej8XSUomwnV3rfuAj1Ll1q8JO6yBTlcJ
pEU0RymDXNApb2RDteiar25iTAGGanPFwINrPot2n5agx5e9IwqixD/tUMCpTgUB8dF+q2V9ku62
Ie5x+qDfPTuUhhGOykGQrlWqcHPQgA7g90Ff+C24zc/+T0aWtSqkZSBb08XBq7DP2VwVUzuNDXpU
P6btMaxjhRAdsld5bARsNp5Y2HYKCUE3DAfiiCj4ipwt5Ein0SGvIsiZhTTRf6a13Xkf8DwiEcsB
pFXhA1Y9f+u0TEl5u6EKeYyGW3wbWM6lOu0F1DcgWy+3lFFp6kutLCMa+Q9DZE9uxa1WZUdvAdDx
jAv7pTUuSsEJ962y7RA3OmtoEViSJlWMMDUZCc57PnILu/aYNaFZ9GMZqCXu0v13QjNreMFShC59
LUkZFvU8L1McrRY+Z+rPUBy9Y2VVyG1byvnYpFT/DVrDIqSpK2c8ohHmd41SpED2ABaLpfSZKNIk
pFqHZzbN8k16zMfFOtQcSooihLUq5I0kfwKXI+1OzSWAnzImjgtu+i0w07edh9X3d9/uGQ+VyM40
VBiJXt+LZQVRm0H+Gx+HKFDNSAMIPubkvHf/lSmRbvNstMeO3UIkCfNse7I6iNRw6MbvhTlH/K7J
tqsdC2NvJ5R99TA6LN+owXnlyRJ7SVa+U6AtIBDquEcmPeCokze9mxj3x2OfREj8tyL5q+0Z47Yl
Gg8K8OjlSd+1mzGPVVV+gMgqmvsT1o3iW5TBz7ru0IdnJv9ABfDQg2zLzAuMH6KMWTO+I3UVyKVR
JPoePzGqMXpWIK6ArLanc35gxhKEOdx6uQAomXuURi3v17IPSnaapD/XsDn+EoVxbtrvWPAMd5tQ
9GJDeSoR8911eL20OTMbso+lpXaHI+59yMeawOyiuxBr8r3CXWt9YVT2NrcWmTm2IKK9dctTAp75
p5bD5gJ1kUluEEEMPce/XO7lTJdksgDDQEAN/HAS/Y5zIZ9Tpiz16yBQ40+IEpCodaOGb0gX0xLS
qoC704UC4lnVSseUAHnt8ttRECivWQzLZbuN4EQFsXTzYjRB4CX5EPyXEOqr7fe+uJ/U0Q3R+iXh
rs8B6Db7cfls3X/OUGmiqMNJY4Sl6KGGMdLMWhdhqIkG+dpmpV62VzHtjzFwzTZZ5YHG51dr+5O6
6aZShfk3lLA1gqfDTCPaICQPTFdD7jZdb/MAJ15tPjIjQmwWxuQ6NUNKkdXValmuMjzdZbr8sDsP
vDjJMl3o1JYYmLpzzaXwROcMPpYCBaveBuQdR8TQPtn0OCNQ0jWrUhh8iRJIT+Hh7hpcDZEXh0Dh
kY2wZLNrBiC/OulOo/onLJe9ZwP2nppEfikcutKS+v0kz7vEGwGmbzMmfCsG0BCiQfM/ilz2x3IA
BmSt/Is1YRlUwwOeKbc280glvI2DvpyeUW+5C6zVLqQE7QoovZ3dClJAuo9b0FwRjRB8Pkke0Uov
CYPBVMUUWQ7AIqvZjf+rd4fmDWKZvKouL+si94isDXhO8BuRAZoPkXNSlYbnbdFlbmnXNCi8MyaB
HBHDhdPJwEIfLZ1gI2AjKh4v4U9R4tiTUjOeZJ/XO06zywqrLY/DGN52LiGvWc+Vjjisw8Ml6Om7
2PxhwK5CGiiRg1gkR1OI1A/hh8XQIQZ64Ikg3ehUCWa7pm6126ZiLfs28c+9K2KcI5HKXs6VoPm2
MIzGYGtx/wDM7b/iNEJaWc933q42F/njbAlCfxBlIpnR4kgOFbAci2m2RxHJMZSPHhJdAlgYfxFz
sVccgAWGpQFmVvieKRn3eg+7TpWYGQ5Ggp4Njm9FJ/buQrz2muEkb1P1WTVzUGUDRyFPIwN7KLJV
/Y9j2eYbXC7HQTIgT5BCDf2d9szhpt/A/pkTN9njJK0sb9+dHDtycIPtaz5GjTw9+xNn22uPuWqE
2YoThnrKvQZyWQjjUovoWGc0WJEEnxvZZSdxDTTiWfn5cxCXoXd5FcD9Isg/Gylj9lLgnHe6V0DH
f4vnNEbsB/MqCp7ghu9MXmDt4aCJ8fikP6WMDLZyQa3JWzYa5DGxYPHiI/Hqxl3gYchJu1X5wmIo
eEuWLB4DmdeZgQONL/5sdAz/7o7hZWyA+mRhTv8LaG29o0Ig38F3AnDOOIXZPHJDLYpyhO8ySU/q
PvTHKqCKEtWmNv3WLNp0Z70zjF0n3eUuVt5mebFcDVi9N2JThX10TLAjivXn7oGUrQhUd2YNXMf0
iz7iUJvaKehPGiBnr1D6LUOeu/LQSfeNPKzIkRCNuJEXYTk2E8RigXJTD6cx4xqR05DGMnv2algW
QnhDJd1ipJ2w354Agx2v+s91xRDbCpQROw89Jyxcevh0qnMyISW1M9E1eKRfPr3tP02656nDHKEB
e1dhSCZPQ7QS6R8rhcf2kcWvrRGOPhQU5Y9OVcM9HYW8jdjpPKTErIw5tLH5C3/MZyZv0V/MJoyA
2zqbw4xJq8G2FaRIwTwdIGqoMyko0j8PZ4zymg0ev/VcfnwbLkz1VAA6dDcEfiT1qwpDI2/MuMdA
iY1aHa7piirOUePM+gAqESUQMe4BblF2ztl9TemgvguxgVxNNscGzV5lk80BZPqto+dwVevieCv5
ZU7am/yfrc30SF+4Dw2MiTRQRbVWFo74HSSKei7oxB2wS8B/t7kQIDju6ArpLuW7oIOjCyUsym1v
pN1xH7cMPD0AjNVqnoaHQ5UKh5Pjql3ic7fXb1PQXk0jOpTdBf63Y6/e/KWsdBsky0PeXK6TSp2M
xC7yiAa+6UmWzHQ+YX+ApAVC/kdcV1y59l9ONfdAxTscgT3uvimAhc/O9xzU72fRK88urj7Dliii
MNAP+mwRMohDHJj8atjF+NIx8eLd98uDdl7rRGf+zZNVa8GycILnSEac2GIQV2IQaccJXRGU6Vxt
6gFcn/rX5YzrwOT8+pduKgF2eKox3kFWUI5VV9Q1tqVpCV7uCRUx1gFt6njKTZX/ZptMLx0I4+AS
AtJsLUxtCsYbI4yUAr0VXHP4hH69y4/Q6am9Uvx+u1ryJFKJ1Vv/pWmM56SLzkmQTcNOEK9/HRRC
h3flbZfTpOcdwKFTE+rhNrwJKX4wXxQmoBUwNlOVmBUGq1OImVQfG2prp8V0tQIQqK7n+IuFSBiU
czRRTWnt3aOXLBN4pikrDzVZgo25070ZjppYadElIamVniJorlwad1EVTeGm6fSDyvMfO+bzC3IH
r8ZgnXoRVGBhDtGQsorgj6jCO2YXHu8dL6CNhCXshfmkuUHywMK3GG9+6toy7OYCEw/j06AIPMzo
cBTnnK7nRrzggluefIcyIuB2GRB/EDw5TNewowrVqFeAMT5/cJiKLmvaBKfRXj6LvL4T769+Wja3
rlDQP91aAqBf8OHPeqyWjAQKJ6+uNnbum161GaX4sO3fC97Z6/l2lnYngBo/xZ1tXhFGBeV2TUBF
/kd4NT1tsBpQThkO0ZOauAFlJkFrgPNPI183XcIqW2heoKziYKuI77vKQ+1FzT0DTefrkz4ISQd3
R3javAWZhzFiBxpfu8zOun1UjCfR5l5nbqFRlt5RnuTNGbUGjiS8cRsv88l5hLrzbnHm8Cp2cMyN
6ukDd0cXJAK3IoSsjjUOkQ31adHlXzTIj1flCN38nALw3KDe5AfJROz7ZMksHhs1Dn1NnD4nIFIx
TmU/P6HN3XHlJEqbTGA/g6GycoLg1ftYXfMYQlJQDKVbtX3IksRH0Nha8Q3ZAKQfuoNMKZBKktom
JTJIWUfwMPKoF54Mah5a7z07z+zpifsWYsr5HQvd5koOsN/YpOJ6wXC6O1CtZp6laXhGxtDLGxws
13PlVXut89fSDhIOV+EpBDp3PYdfEYqzbKvtbNLe54Ci4SEJ8R9baWCrjMzp02fUwCHaKELM1HDa
MkFham8PgnxsHakLXa5w/40UljWDad+9kZmypVHWdLXcAlpJG4eLiKI3uFLiPgg8f84s6GETxQlI
cw06NasRTq0Sp9GzkxP1uLw9qvqVMaPJETHMAA3GltIT5E/JPp6VEbxUNsLpe6Cq7kT4kJIuLP8H
h2cj66jtsUdMUdk9PkZmDtZomd2oOd7X5aDT+IobcRGc/IXqQ2aXnNULPjguUeGSve9d97hFBIVQ
W9QbXGpOVtMj23ffeZtshyuDRPzFrHyP6Eh3SbM7/+vDqS/RCEgXEHadV/5tjDrkSBGbh8sWsvOC
ZOUhLtAf+QnheO0u7g27ByfphM7lzcyywrGi2gq1DcnaOCKpTAltt9d48vNhupu+XL1Bn7ipQMjv
DJqVMlYsBKwW0/zCL/CfcnWYvvTA2Yu94kVhua/4Fek53XVHS7441MQkYgbziyScBgD+UA0xikfj
UivBcKu8+TxqOJJ45LCTuCAMArBp0STL+JQ4+RPZ/J/VcBwp5VJ8xhHzvVWiVgc4nFJpGVZPKcG9
t/ctl1okDY/Jlff7HbLNHyqkD3VfYsHTnWhOToSEm40S9GcqSKdyUwgABTcMx8IekoDfEqzKIH8u
WwOdJxS8yKPoKAxAQk3xML8LYijc9SigRyfkNABE8kXNvzySjvT+KVZR6PsuvwQULIe+XJ3m3z1D
rMqaRFUEGJdOybI8a0eDlHk4Jom75yqp8UVOnUm05zFdDT/hm6X8DuD1E5/qw/nVKyhA26zeg2yz
Aj++JUhWfakxULpC+NNIIGmfCdUpEcvFz4jsKhnN8qprEYjccBFNk5FWLIBtOXxPpAdLQXB+SpPH
Vma+/ooq0ey5hg54IF6aY91Hno44ROEU5STy4S7r2YWIMmSZA43UETe1Bj+P5mDe+iDsyOV/uZYg
cmED4uMFRUsMyb/X/qtwsElaMCM0GDq7uT9WSrpzkN1rK7Nw2Mo5jae0y/vEROAMhqnSSD/2EQ+X
m4uicjRbs4GIUAi4rmcRcLa/uPr/4JtCfcdx0yEECvY1ttCYZPwI06E/sa5K9RPWIRb7VvetUn9x
qci9YNG/hVTju2+8jWvw7GV1KC2lrkCe4BJ5U+uNUT9PRrcCNWwbq5+uNFPKcwvkC/ol+QZUQyTf
dN9tbJcc+fJ8b3jTMssPWqyNwelOucHvn5Sv1ewLoomwwcnUSB8Fh9v5AFU2oaR3wsA76kY+fcm6
1MTMcbI/i63i342EVrAi6kJJaEAdrAZuYkB8eQbuy6gucj25a/EVD9x9ylJOC9DgKKqPQJwYfImR
i5c2jogEE60eNdnEkZ4DeuQT3JQggOQy23daHUo/gaatjcrRTCcaLJrNzXaWWQuXW7sdKxEjszpr
3dghKBknUe9mdeMqJSqaxQqOKZgItEedQWQpesYk/39TPH5WivP8knWSUMgKE6tjZA8mo2Tb1fbg
nlCYQ4PtfiLX43CvhIIzi7HUSGL/311Pc/ccL0M2/eU2arWba+ho/ZeqSbg27xI77vB8p00N3L2j
qLqWXAHp9f4118PF8F5Tg1nu+NjDVSsT1cFtZBVEW6koevzzj8tcqoj8V++f7lRck9C0N05VMzNn
xdt0dBWXmDsl0Lo3BYgttWvn7tMaZGV9VgCis4QtBjEkT3T/Lqt+qeEc4nKADO6idaIrOaXAjGp1
oDzNrtJzBUX580vVQ+iUE1d9ufyOk0Au/kJ/UqkREYy9B13qfUBxihVrMOamxy9JyYmSvRBhhk8B
n28PQXsvS8AjXG5vqwQdtUJxrk7vOU6Od/2fwVIgYGE6D6Ydfv0AitPDzQUdFUsv3tdYfhLl5muo
/KUPZjHPVFHXOHxar71HEi0hUIm8iIR0KejRlu8BvzhppEnSSWkinWGvX1DTRZdJcx8VmHIiqKRN
BcYmCALtudAwa44pIcM/EavVJClQPzQNMbPNp5g2o7XFEH2fT+mOpwJKsk4inZAzXBLzS8coSQmn
n+RpcEevCeali3Wt6WpNUxQo/Wckvj39q1j5Vq8hVk6riam1Uh6FYYFFrwkkoLarsuKBEPQr0tXc
sNtqXCMHcYRWyrLVZ2DQwWkm+xmzLrAgWiQYJu0QoBYQmBP75GBDaHvJcEJpUYW1BvuF4anU3giz
TyXNhZxqzqhObCcSNxth1m8RbeylG+Y9CI0/PLrXvfCs7II5ZiCrLxLlQKavjauOtZLRzdjmSR5A
Qz78Pit+mkniDiFyA1RTKDkGIBRO6oChr4Yh+ja/+jvDXl8w5tCL6hs1yOcjMBmFWw/EZ6I1Al7e
GXpR4pLsoPmy/GTu0KKnY2YX9dnQgSSk7a4hzRIayghEYE35S//P7DKEF7Vcs4F5NlA50XVxLonp
2dUBh9OG53+vSzWjXlpgvxg5r31EZwLZLUeD5bSaAEom2A6k7LwYdy7dYWBZSRyIucmzkdg02G8d
gcoIe0QKLRNwcr50QGjSwJ/lDTLmXW8n/mo1iHFpHvqv46ceCK9kNmUZpslhA+zKWpW0rxKVfTyz
zP6Tlt4Cd1DRVrXnH7eBYL8itO1n/Ck+/dVnD5xIFfKyxvuIAhhD/bPkTkGN93oouKDxNcwTeiHT
pUHOdx6zTbxphRR7xEjETRrineJkPtcnRlKb3UUBA08TUZLcItB7hyAYFH2SrRshXskNgAnzb/0R
+D+/Ydb/tEry/SnS/r0ioAUY1aO8MoB4dm8dx9MLjOkb9kYuKHqSrNqwmXOvB+Ewg6D9RANxemf6
HhQ6fSLPpFebs4rDYlHyiJ8TbSk2hdVhao1ymYx8cL1TPrr1AlUwHfXwL24e6rH6gthjA+BJ9cbX
3rUVkKuJfi07AsHthTVolNBYN0CLJk9Vi3lH97VoeTsxm0O1Pp0Y0zEuGtOMUqpIfEQm1ekX3qgq
TrFdxedXRX5buyc9GlIB1V6wkks0SZ2QVqZxW8087LJZZ4CG/XDk7skGOhxhZavXMOohN1w3jGXu
npSH50ICDdWsju4jdbCjnBmkwwEMSYFP5PqiuZ108mv1t3HvbYDPY/vnLfHIpOwHQsFnH8kMP7mr
hHIQFUotf4beOInXl2xH9tdW8340yMFdParUbtStF2J5bL/imsqYX7dzAK37fsOgs0fL+t8iDWN/
7Hg87RDV2YHjMUdWLBH0A4SPmKufj0wS5oRcUMXeZaJ6y3uEYqJQvgfEjCl3U3xq2g8UYnGDl/Cf
j/7VErdAIx1gK86GDEcAbJgN0+FzACx9zHir8ZAsDTHcNa0i020i5rB7Hp7FGGaKM5cvoPwXKsFu
YENuxbrzieFHa4/W/BTG/sISoPH/49P3tQO9dZaM73SDz3Ndw3IFB9wWVdZac8n9xZRRtpb2kw0q
LiQp+8uJ74QhFr8qfStCPpeoM2bfrWOqY1dZxPLSlBfdFbWrwU5mHvIoOIImQKL/qmrxtWf2cMVm
syWvk6VMQ0Y0i3kAnEv5XgBpa+M5je4UWVTFQ2a+yKhKkGinUMG2n2MrxpTJ7aE8S/Ngugzg968m
L3LBfMl2vIEORjP+b7oCf6BEFQO+H/LreUSmfAbjD1sCQKDnHRyvSJwgIAb8FwmdkZ7+4yDwroHI
t3RN7W1D0POBCMf6x1DLExywT3OTuHZYnWfGhk+5GZmk3V682PJF3yKtdQdXkrunSi05pOYwWkG6
f7GFxRWc7k1z4qEk9ac3H+nN1ufmA0gmTgQ29OUXOO0V7/Kj/RUmuXOfEx5xZTGbMj574GdaowgM
yAvNneqtO+CqBPbSbIcf7n1kzIva5/vG+NlyF956qEZHvy23vJYgGbc4WXSHgLiSUAxItidgzgKr
fZw/Udp+5NHgtFget3TyPYJ4RAEwl5kpMS6Kzpy9wgP5mfyb6zVluNaAq5Fc/TFv5FWkrGN1TJ1/
H9mvkkiLm2hW4KwMf3JDXtorh+ovkAbDreUyTKQddM22Kc3mGCJBov3tak1aVNhIgIDsdHmBqsaz
j9Bs+/kvmO09wOb4SKJ4Eq3AuCm2Hdf8ytR7VXsYN51OImju0k1yYE4iXDJRbTAlVqU4lR+EjpwZ
yQmC5xoFz9USQIqNyk++E+rQlkby09ijUiuZIl7n5Y4ugiFfafzmSrR08/llAFfDbml0Juj+t55N
rwObeC9uK7pxyHN3cXV3La7a6gD3IR4DvFOOpPd1ef+pOfe7TBGAeei1L0jUGE/7DxlE4ifWk2Yi
UljA217iM/9nE6gorFe/iVVXlR4gi21yj8iPdg+Zf04pzxI0UBSeSsZDsEFZlljIPCWztxCYfHU1
QI9pAErZcFDtvhnQUYUt3/KBUJ9kFPzGEXlJ/9eSKX2IsL/wkrMIvZJfSRITMES0FnleN3Mriv8v
fR/43SOg7Py1wWR8AFEjErW7ZxG2LkNgIyQ2dDrtoSAIugyCYQsZIhX6JxXS0eBsvLSKvw1DrAD6
SBG4DVxZlZEdSbktcAcEu8nIK1L+4uIQd2DR1JfgSQZQJRLTAC6DP80isBwGqjeumdKOUedovbtm
IasUUq/RA0GzVxeYEXplBomf3hE0H2FydNp4agybiOu2zOmsH4W3cRUm/f0nQHIQJx6xNpmevAu2
KRpIHeAPXPj2HGPR6OO4FMy2+Si8hdwQ1I9OrFpmujcl47mkZ+Qp9yg6q6ugb0V6akiV8ni7GbiD
ithl950zEbVu91GcBAn2Pt63MEKtPQ2iwT8oL8kCdVhwBlTiDbPlSvcSLdQDdgCOxSNdV8aw+9q/
9eWgdXpv8Ri36rmqx6WLQNl813rCLdSy/o3NRGW49pP67xWb/CaPovh9ZSDe4bRCkiXSiQMi6VI6
FWqgfoauZwNmRG/ZYmMENIXCcUCw8TkUlG6J8aM6KTlCH82dO7YTSNBB0Crt4+dm9p252zp5RFxW
Uzmu66UVxwyTaiJvBY4M47KZcWInmxcXR4qo3GhuqPOG6+nBMJjklEAXDgsm+t4nEqairrmS12lf
vMjI4caJPg7HxTGcFnvMiYGMR5u89eNtwd+YVmAsejoV6pF7/ATN+C4JVRPN1J/SlFTKu7nm33+a
atAE9RciknuElcuAOq2fGOfHa/x77TDH7MzGxavwodkUywuX20V9lMaiT+SeACvz5vAKFAiOQHbM
P21fLDoH7E25shwPu346dNkFRHPTgsdGZgqYcldPydeTuRt40aGhEt9wvgBuc4lkmzchNzOnGcSV
q0NSTU+HZGPTfLNomUSGQRNVrRZvUqyRXKctP8FnJnFXBofYlIKu5ok9W157+B3scYVwkwDX01CB
zCx74FNVQpUn+6TDhhJ+OTdIE3TzlDK6my2S6Sw0VjIbDGOb3X3qRCdiPuoYMtLX/pkgfYdhonxR
qwOYZvjunFxNu/+HgSJyHRuw6dKIPp+cyW1IpOG5dEg4wjum694D0oCZVo6VHBCKPj/83K3pLgwl
uV5lQbKCGqko7WKj6e5KldBQOVNSuqk1DdnP2PETciJxtlC3XycF8eLvBKCCaqaHjcrsyyJOVqoL
mYW1QESlctBesDU3lyXUf0+GLIy95FzEI2HOwrPRqxvYSUJmBvP9SIuOHECbhwyTCPIbae+eZips
D4JDZNeRimGAH4Dq8t5FmO4zGiIA6IqbpbbvghsaI/g3IJPkxDXDNswTs/VliHQOETgrmqMeCYlD
BPsmnBmjPZWvErF1YAbH9qR2mo7UXdcxWtfl+948NbCjCv/4IQcStXaW7SFsK++bbBmj8EKDDtoy
Z+BapkPRGV/cx+bZqxPgfSnmQfAJoAwVu7m6usGguigc67OueNhJH9GMr3kuhiHdIJFtHOjbsI5w
sv6ElSaXVs4uxmbiDrhUkM77h0a/Ud/o+3xZZY9gY7mVNUnftG3JmegodxFifiCmbYm1UokoupDC
CYCb7ksrY4U3Z98c5PD7h8atjdze9qY0Vtj7CvWs/6QivYKu3J19tVJYOqqBkvsREVNm5sSOd9O9
JRgdgn8y5RipDr1OJSIR6GMgaQ/s/MH4IJs7/JmLqfbnMcDqSFcDgCr/3BTUEPLgzrWwLB/nMnEt
qN40QdejBkuG5awJQ0wiW3/dQDzgwbTnz1G4AZoQkPJHlMQcCYeRTpxMTf9wdk1F6WA4LCs+EdWq
FHoVgWs7thdAdKUikKBzKLb40Fiv/M+5lJhmIKdaruoBs/j7bazL/9QevqJUN5gdWVRDki3pCn/3
PxC2Ulqt1lbHxlZxGhAR+pG0OnpEfMi2W2EQWboi8zHi5bML+ZoF/vS3KR7l5LqtXIqyQs0e1PES
1Pz2EjfJYZXoYUkNaXmXGMzqoCq9kQFNj2jqXG5HvwzWbf9nyfrSIFzFpSZJp/SeAv7wL7CPacgT
8rWGXDVrFATxLmBWXHZMoz8Iv1kEuW1emNofnLznBvnKvOVR1vH+edvhD3vX/emtYqFw4VX576FS
9UlsQZ9850qDv1YmxLbGzRsasFo+aY6aRQxfV5OOeKCKXimHlGd5W1NDxAuy9BmljtKBQogr8f6t
UyBP+G+xDDLk37ZN9nfnvLYqEyzYHkMzh5rwNTH3PYhqCuMiLNS+M9hvsAMGlO3A5YTb0rrtx7e9
Cl8b8nT0NXlgPw2e2PQxjxht+6Tb4FPXCS2Nhjp8OosXMhmtCS1LBAXp4TDJnctvKvcj829GawEG
k7A3WeSWA1iHr/1eO1/N17U3gj039caWWwa0kiQoA5mx0OvfPHNJaLhNdNnvrxx105SlA5R7b/l7
gXO3aLZOT0q01AZQLD8Bt7NdhQrIs06wDYO/0sgGPacG6DxhVlcB8vqLrMxg8uO5Y2VY0+HQlGUL
Zio9yXjOtOZC1pat8Nb69gpkMyn8gwpOdzRbDHDjTmDzCRwkXqlm1mBJaBsWfWQi04+j8qsCaTX7
Q+Bmn86ZCc1CWDOA94PnZ17Pa1YKnf4BkGyo/bMo2rdwFle04tF/gE8NRDv5ntFsaijouQdjfMtM
0dblZUMvJobeCGaxyeymiUbjUQc72ToMUn+oT/pQydjB5oBnJiG0kTeT3aYfyla0cXcbVSmsLsY6
i0bo8iFo9ffxRa98IE42YF5G+7fuK44GP3cXflyNDLJJveyqvB4LDMBkMqymgcNTvAL/KX8xYnlS
ru9ryI0GMIwDlpCqA5JbrVgM6yVK2+pX7EtzYAjjvnDy2vh+n7/Di57NRuCFKQXaaivA7XhuUY61
uMhfemBRXuxth/mA9HkjPeewKIwQlRYAkD5H2/+6h0amdNtnOIYq6lBUkEKrmM/TOTTa5WUxPhDo
WKYd8Jn52SvcLqfzD4gGXW4m1VwgpbWgckNSrxXJwb2S2H/aBMrZTzBC4wQh+qNOKShRG0QYCxqe
psYENSAO0HG119mZtqgy138WnydunNXGdsblmROe0B/7fVr5mWqkGqIBq6ZqmqzYO4k975ETbTW2
wig0Ex9Zh1Mdb03a6/jv5HjT8rrItl9ERBHFKnFvY7bWz9Po+1KXZ9N7XjcEwSN24lF0Vallx4ei
2WCPI60QAnbFKThH7pvXqBpgmpet9x+JZsl7iK2dUB/or7ZYOm40tj8pPAVIbxL1ehnD46siXjxl
SuVZ3oYiQJ31iHCm2Fqx0C03EQodAs1VCUonqmGyMnmMg6on83EWAb3BhJp5Keb6QvwvEptGVB8M
Q300QOBYSogDG7+yEd3ynPsnQ13niKf07DO1wf1W4EnKKgkwQoZ/VIyBK4xAtdMx5qSwERpbJfL9
yAXyJ0uLUyznBfYLemSQ5EA/OcCEJsYbtVlwifF21XhlqGH1onuJ4oOarfXHRsQ274fcj+UV9obl
6L2XZSF9OQDa+y6gUvAsKRNQy6BZ7NgyiuJJp/xdgnrdcdZTUxh1FokiOPyPZ2vVjjssHZU3nQC9
F+45pJhpYjKb7fUOTKX7gqiE5cQjcdsKojPYsOPkue7RmN9MNuillYchv2fqGP4meorKvf3KY0GL
H1IN5lU2o9Zw+CtdaFJQ110bITwPtHdkER8jcAfRnjJ6VX2xiZBoSDfCv1M/a9hoFgnHVOQeEzx4
9JnK8ogD/K9W9MPa7R/re3Dxrzg4ALrE586hegL77oxdi19mRy0cE0O0gcBeZ/qhtjx0RJufmyxJ
4ZV+FqfHU+AtRt0zMwODQx3t8Jml998E6MRai5idYzqTKXf3r6VzB4yF0gTuSZS99qAgFmUk77/0
FbMpyEV/xT73hgn5RBh795AlW3j6aQdCp5ASjsxe59d+2jtuAhh/YUkQmMjfK0HgUYtAQdSKcJwJ
zUHY5Lkl6Yj7m1eMAa1j42z3ANz8UxuvjCoNmENlyo5EbJT9yEjt0SQt75rn6eE6e0brXT0NO74W
rO9oGeY4LeSv2MV3DDmEk5MV649uEnpIBgWXbpUFnPDZc8wEcDADpYN+BBZN7tMNFPS5UcnwB0Bi
6BP5am7PQ9FwV6OEGFOUwt8tujmIMYQWBLaOaGnbbr/nhUWXXF2bTTC3l0H35PrXSLiUELLLNEoP
VGo9hsUWFSmgQ35cIBFtsT/pNeR9CPLtdYM3+xrqDeZvuPYCLwDXzKEdeNyFnDjM041qeTuTJrjy
xRmmGJSjz1DuR3z+Ja/RtWp4CZPrcd0KUm4RI/kJOK9JBCdsUO2FipU+RKCPziJWJ3DyTkIx3n2x
09iRxiY0QCZZN7HNazWWMWe6m3ZN539+w3X/nu9L5Hqttr1CgnVCxbv25U016eEXpO7Wmsw6O8n3
NP1fECRUi474V+F1vRIG8Z+F4TouP0xH/PNbm56AO0j+PcfPR9wwGcvL74TnKZaKzVylJ2XBmV29
ffU+o1wlebK7XolRVNNecMjZiCbkqOzUdqOJsMOamVRZ39eh43X3FiGi8W58Iawop4pZy1ErshJf
l3UEqxGdJ3hYhOmgvJG0wArkO46hdl7aB4UCOXWEMSsN2n2MeBwt2kj7RPKEZbW7ddiu4hVWzdHQ
gyVx+Hf/BD5OZ0ttV5jA8scnky36lLdL4qn5FCnf/sarDf1OJvIBB7OjECq2hRi4RTOhswD3Esxj
Sh9BVesOUOg/Au8X92xXzsqOYvj6Mr74p0dJpJ3fyZI8X8+s6UySzuQ+N9yW+nq6vf+wqDzvCzc+
uvDBkMKbK/TivBYrDV6LjsClO2qU+KoEYoAZWlt7g1Sp23MEogDcQDPs+wD7D9sle4EVrJc6ZCE2
004Ow0kYtVfwE8oPe//aGd3kPg/y+lvWhsBQP8eOdL5L3AAI9PJQkeSovGmaK18Y6rxQNifTpF/L
30YmUaH6WSAlJs6LbVOEaKsi5+mxjH3g/ktxlJVNoCERx9f9xhB4kKqIfvAtDysrPnBZ//y7UI2d
db92dQAINs0kfBELJBaCNo0iI1HWKSXZAtwm0WQpZ31UzxkWuZ/QOORAgaieobXYtQW2okUcTncI
THUPy+/A8Ohk9y1TMwxBGSqZIyLRPRMict78+wux5IpTBrKcMrrWD26C/oH55TKS7RtvjEHuxWfC
LA2HLSvkIVrCQeQwFDdrg//EaZaZ7NUXlyJcUCxpMeSD0vkUUrexkGzx4Dq2uXn9UWDOQ9RxgV7X
zi9bCf6E6crRd8ig5CWezyhandKTIPekquAWm+Y4hQbdHWapkmGO5tIdpk5ECMWdaEFzsjrTAg6u
mkZEKTjphFCIR4hkQVc+h5hL7BhlxOSUdSYMFiHKqJM5jnZIoKdPnVXNtSdTVFCHGFFuR26jSd6z
LNdqRdZ0sDkqipKJiCvEObeNS9pFliw1T3rYHn7OHe8MyH6VUObiZHfasdLi1DhxJzCMKbTC/QJP
CceX9BLpY3HKroPAT7AVho9Y8q/x9Lq1Sr3njSvYZkDOBQ/vlDEB395iGLwufx+QcGHLYoSh3p0d
JzYZ3rc3A2a5C1HmpTQ8ZSc+e4hsmnVPrQd8UB/ZHZ20NfttLeeL0icrzZddA+brNM7r0VL7WxxP
xEUbrizdln6rOdrjx6b8auEgYtCuKVn1cHWjmERIuvwbzExO7o8vXwQ4DQquWCK2KYzPpL/H4l6m
wAnkylmKnYHdJyvNl/zZKCCPCgfI3WgYdxrShrIUEiTUBeSmI1BhLHAoxqfZjAFIMmP52L1PNt9n
8PMiojb7wy2cVBzwIWHY0i4GfhaOOu5+SvZbEQhaVc19N4C2t1R+01N1eU+2+d5ZoSRK/SQabkQz
uTzgS35JuLmRGNTSK5aNhmSysmuKxkLqRFQG7G7emUk7kZRu971UzNZW5hboDFw2Sp1gb1L+ze/E
KZg0vzd1cBm3BYIY4GnymU256L0FEEo9hlanBaXz7XvqIgu+g5gBZB/LI6Sscl1AH+jii6iaTLSE
cCiTFmiEtXDEWi4EqdvRSj72MM0AxKFjjzn2ncE69Qzdz1O10p9ip16oahLuTw3t+awSXZ3NPNZz
+f796PyBtTRsSVWTTjZzePIM47CMWIC4eGkfSMz/k7Qe8gXAIxIJPpRRHJXFuQrQ9vy3si8sPd+l
lhU4FDG0zLe81TxdDzXNYJu7jhw9A7zsSKvJs28o3rgNpvLwTl2dsUos6KFS2zhHVIA8KXmQOmC/
Y9Y0hVq81xOPKKX3UZQ9436Xg/6mfQkiNkqCnzjBVjYCt0Y1kbxf2FuMI+f8xEdDpPyTGlQV0uuY
NzEA3cTDjs762O7acLpqamv/QyNN2Nixpr5cGrsvJ48wxQFFZrETiWnZEv9rF6AMeTp+81L1VpPP
67b4bR0uHKnDuXBLcSCc6v1FkUQvnRnjxj6G4grR7DOKdJiBVTDZppMjqwAiALXQm3PIykA3LhwG
LRoBDNLMBpcq+qBdUthhu2856uqPeFbpXC56x3GkcR7sYr2V0Kuc8QsDI8TZ/mJC2SoiPeQWHXpi
vYTu0MgIYEQXQxU45yfbW+lu2yLsFvuEGfxVNli0ncwDs1N3YR5V6SMON1QDNLKBpB4IPhkp6Vfz
3s4wlzh1qn/+ZGRyKK4QD/tJ0+Kl2GfXYBZviMnxVERjTnSxNxJ3wY+zkIPiNNKXaqnz/iWVMiC3
HuDU+hWr/KAk/xKiLST01UMeUgJ9iXdMmS13f/D7Y2rUcY58WR6tMwx0McRdem7gVBhT5sR6vpwo
MuGgPgF4L8sF9yXGw82D6w0B/LSxI35bC0tbDFpwA6Qo8EsJfcS+/0oa57R+rWmH9UCeWAHYfbEg
vzPcISsxdQ0WhjNIef3Tg7kslbrMCJbZOz8WZKVQhNsfje2kzl16CGDycefH+m0aWpjAdOlO7R7R
EsaY23x0yGkJrP+4C75S8VIxmI6pZ5HgmhqZEg5W/wtD1BCoK6q5tP15XRSo16R0gbhbZpWf5zTc
GoQNaC4HADJ8ILG7Kb+yunLLz9OEJV2p+pH9M13+dVVEmdAhE/nMFN1JN7sgJpG35yb85hw41vDQ
DoDjm5j0QFJ4wgrRkfSTN2DM+PS0EM3yRPgL2iA8Q420LQJtanjpRt82UObLKKH5zVB4cuhrYpFH
dByb64a79RtmpRD8vILhMf57DDmlbN1b0qHEu4JhHp6WH7B7g807DZFZpgsArtEyhZQYhjwNNMoh
uqXi3MPh+ZK0rfb0v8z7z845smWvhdGbl0lRvrapswRhOiSU8R4onH7Z/Yd3bm4kpZu/MGtGIo4v
HnQj06dgu4sXpv7CssTYbALoWo9/Pr9AeZkWtgYL2YxHYAE4ibiLTJIStVlWSvX/1WxinUT+izzm
fKB5sjTso8Ilh54GZssfmIJNTnUP0rzPmCV/zpn3FZC1TUln1NQlUFWH0IlUD+o4jAHYsIfxhAv+
qo22pkgqzup1XyRk180q1fZ9n+UaDBhhnYRhYJ9EDDsZZgRrp360f02zKmGQe5GZ1uG60z12GFzY
N9zXtVEjE5B6bKGPzOZNdQIGs23W9M3WKXSrnj0135XPsevytdPljUzfZF7YE1c7cNAHHNYwW2zH
pA1b3NMsoGlUs+xWM3JEvB3R33sshWEt+iEfy3UN7bkrCMQgC3pEq3DTpcuMZ6tkawcBHHjx3UnE
dRIW/I4Ji0yuasn4qwEt1XVYeZYGKMWCWW1MnMrk52yicgh3lcLqfJzQ3FlAsecTQK8x6+t0W2Ul
YOjhgqeI3fnx1pSP2SmhPxtxQmAeXD7/pXmfzsxe1qg9sa5CJAzYYe/Cf2bPtsNZL/HBTI6HuYNY
Gdty9lZ7s0lmfhBcvfafXcGeyCDZ75qxv7tVBkhv5M1VBYfoVe2KKRYwHZGA0Aikr4i5uQ5kGK/t
+moywTdfQjwpSOFvfc3ThZqwd//3iKe7cky+2cK+C6D+QJmTHmUuUg3PfKtNF+K8ya17geTQWU1u
MwX6a/paQgq3pKbD0s04kydmd1jKUdu693382WADyat9nZLG7rK/pf0BGxRd8Fw6VvfX+L8byebR
8f80TL6UjkbW0W2wodDit3Pk09Fecl+QjycPWziBr00wsEwxs29hMFmXHUrHNkeBMIXUc0laXyTo
2c6C6TLBQf5Ij9i2QIBDQfPXboBr/UfC6e6PKfsXIlpdnNOAxK5zK4WMD1WfHIzIiAAqwQa3bq/d
COTNIsM+5Mvf7O+hGkm6eJsXQAjK8olD52xBNB/o/rU2wjefQxB1FZwnmGs5ytgilPehTIAlkc3z
gRDpQBCQu3WO+LmYYtPFQm7aiSBokw+bk83Rqmx56rmP5e/SOM/POh2PKJcHEMxYUAF4fInWCWYO
2bSZdj+QP5Y2JcltE0s8iJMcfHhnw4fh0zzpie5HAvowk4d1dH7iART4hve5ttdVtP3VL/Yd3+Vi
eFllbuFiyFN7fnMqnrn55Ttw4BMjmA+AVDLx97hXHe7IGfSRQ1gbNXB+bSHm4dJjgLXkr8ti55/M
RbRqFIywT6pXXBw4Vg/tPOTWYlSsgAs99Hl15BRtXL99IMyMTiXQc0XRYwPRO9/ydkr1Vgr8CoMr
ZL1hHvzwKOIUSAODbj4/iK1YyNF+7SbHvmnFgPAyoyXOSYKnchVGV9C5mluVhM2xqAE3UUUFdB8/
CI4FZS9Xm1kcNy6jZjm4Ec/+NBFEAfbXWCWLVeHZmFYBxa3ZIEaeM6bnjLWvTGTuzRlawk8Utpm5
4DoTSTXu1R0YqYVIme6SVkF8SlQY7LlCKXGyVUOEv4WA/C7E+8bX6q59NjWWDUJvaOre+uMP/2/8
bJ598SEu1/JrF2oPc8ZIpehUXmnGFmuZgBENVT+3yPQE3c1UPp3XJJppuwItKgmHVz3oORi4jcPq
k9g1xhbuM6/nYrKCB7w2VbYixB9hxE6HszhPVvqvdwtAStcGIlZ6jVOH5x08yPGgUIoMEfTg+p6a
9qIDs/nH7h1MeyKq99KrqbtN03FMaDJx+nb/J44dPvtF2X6va/peEUsM6dzjX0E+HJMJRH8MzkRr
Js3z/cWR4Chvb9LFF01Kxz+hNuVnMkDkZuerBqJLmjhzZD8aEMQXI+CZJPQ6wb6w2PpMPDmMjeOq
GDg525kYlNkN0S7l+vFQ/L6qkGIJZ75iHWqCAHZULFqAP3LmykYa1Y///NR2sNadBIoZdtK0R9IV
ugrJgh+UHMXQpmp2JZlY8rsYSizPAaRkWVDUhylwBzMoH+3JxHwyRcurcUcoPR64Ra0LkooW/3T8
vx9WXW0yJ6/f/5PV2fGS19XtRu0tuDcTtCV8nd+PYQIO780pOcue7J2Ni5TnDIqmKFT9eVaGI2l0
TZljXDk0wACfFvCfr2MchXBrF9ip9L0mb8wVWvHbCXbuL/YhMAAuKqP/2KUjEL0xc+ZebbN54A6T
3fPabxNd8xZhhr0s3Fi+cl3soBbOiklfH9D/PLv+0E4AHm12tijTOqGJGHfQt0v9GzjZ6I5fmsxf
ov5QIR+Q4miRiQSi51qjzwf/nxSUmeul0XaPQjYFhmGYEweQshaYxOPE9Y9WVY+MVjJAWrnEI6b1
6rZsR614tyEe/Kd7KaUlRtn3CAOkcjUn1WZClURyBAOE1e0OEyWlBy1J0+elQP7+pDn2Kep0AFnx
QJPlHUbNjspu8uYHP2FBpUSKt5gUjZ7YIEJUcFsNG8KV+RrU5ztrAQuXMX14lyNrJCF0MscYIBwe
4Ko9b9+pmhi44Pm8OlMiWxlSkVcQ6xOalScnOLvLMFmMjeJL4ME0zN3Jb10TR4iJ/D/jsWaPhAqJ
tETvRVu85QMak3N1+HqeIIUWqS1BsHSLQjp26Pv+v5VEZB1l8IdVxHBybT4TevWqDtzKTurIumhD
mMAQwj5mQgsQiyMettFAoAnvZ4wBRPMxcrQCAW/VwFw/Il/DAQ3H0dw7IC8VZieWcN5MkK5VcjZ+
diYR8hdbkOdPNKdEZZC2mj1SnbnufjxkrSlcAWe5nibwIrwJj2AfnK60vJvAqTeFXKOJiQ2iql32
76RlUoJwzfsJhDUZnigu8ZTbsM+vSWRFhe+ihhGASw1DebkV3CnAt53cb6lH+vfKINN8tyDQ0jXZ
k0B5rAqUWuM5lTM1KoBH65psI3nUApeIonIfBY3Unyel4dALxzCkHaSPXdfufMja6JQUQ2FCmE63
lXIQ3QhrGRkm1NL0Et9Tkk4Nz/RPF6kEF8nQgSkgTTYKjsmawbVW0dmam1tf6s34tJTgOgeIbV26
l0mbnel3F2kUMJMRtMn84p73oH5JmVCjwTnfZgr2R+1fRunB6UTr1iOdwfEvmtMyG6pjQiEj617F
LrLk5ba210NYKPHSfRNR9/mvCGxjvwaR4SW3yhSVfPCPz6oBPFef7wQUCoepIHFCQLs8HbAfVgyP
5Q9yL4mwgODPNle7onjAxhqMoCOBmC694goWeyaL8aWiQJt4fyFoFpJ7qeT3AU0mWLOdNdF2Fy/m
HRyrJzoJ+PZXG+cv1FInnY9QhRBc6RXGuajfSld8LkPeOneYrI5PZ9YyFlDpW3IW0AtiH2lqy7YN
0mhg/wCvCaRbNQ983juXEQtOjQA6f/MURSGukOixaUmq1Sfs+/ak24uwwXpC4hwsfIOAvaUgkV35
tzsxAaBpslIGKdxkyg7dWX7QscZD3Bj4CkLvzsAvKkSdUtxvfWTYXgpe6B+R4vkPIPQ7hQNwSR9i
CFHiEO+x+h+tIKKJrMb+KouRh0M7fv+2JYQf4axjVIa6ptjnH6sCm7CQWg/qwFL2dEhiXFiJ+IjC
yAeRloVNDpb8nag5IvZC/ZhzInJlCaHCi7nntGiq1ExaTje0HqpgkomomFLD+qw2JJSMcxzQ0GGj
L4WhhU9rmoJTXIwRQjS6eDtHnbiH4QS3Iy1B6nRd30Ndbl7Bha5rhuJAveJhTO5GH5c1+N2k/bHn
pWsXiD253+TxR6xOkUFRSA9OjA/fJf/w+bAaACiTJ3qjAGg7GRz8svMWSjWN4vh+LnejYzWFPF4N
7RK/GQFXECXtDEC+VyAW8LllMCELBSf6VNfKXi0Drb2/UMKTKqyBq6WiK8oM2ce8qYsXJEl3cOps
UFXsCZbTm43V59eDIZMaXdGl0jJT5CU6hsM5cqoTqznE9JJVh1fbA3Qq9lezQvxwLRRnneCn+2ij
HhxOnzRtYx92pN3riIgwlMZeURxaNsTqY9LofIw7kyysDGY6DxDIRfj3syEyOnC7TzZ5Wwpmt+4T
SBJFFKHwyR/y6i/3N2nkMoVC2xpuoZVwVW8fj1fLawZWU5I1pEiSkV2vBsXoZSGJjW49nrxKGjfJ
8jokpnJGfemZklSWS4KOqhsMIMMrMUqFFoHk4Og6pkEQ2Dj4ibv1n/4De6rRJh1NW2qg2/ZcIZRf
k9lc3WwccPEHbYKsBvInC31jlrin1B8e2dw4im5rYNpvckQO8QYgvOt5o0XP9s0eFwO/wDtaQr7S
kHPpqwVTx8abkvUzOL4r/2kJLuTnd3GTexjFh9f/8eIuUfdeGLtxVJByBLAAJWdUBICUCRwwA4zL
D+1ftVwooPYY+uE/IUHM7McWoYNM7U2ISKGBE9HeKdNV6swdP5Axl0JQrmi4LLEAeNzS6vwnuX8x
dSoxj0H0Gnf4iKOIJMxB1pYwvCdAVi+w3oEW38r6VhGBmL/PQfx07BvhViMWw4DxBrFuih0zfWmQ
XS/qYrcJiUibHaTcX0GQ8X5iLBLEwCwSPnEw/ccAdqZO3K5Z7R3z6p/RzWozPeOvKqJEKTpT35IC
Hut1fNdK7TuTam1YR9/A3P2g5Hfo2enmFbp/oc5OfA7+gg0qtuoAbewYhWfUyz2da76THJ0fbw7O
PI3HzV9bAsIkT00G7cVda1qbrve2RJ59R2Oys6vR+5BgeOYT4NPfMYFLArwTeKMwzYbC5UUtdoUZ
756ORkXGP9lS2bybZ5hrRvR0tXEsQBGN5SboX9ynIl+i3pyxrPUudYa+ropwJEIbmrTINYLVBCsz
NepSng5mHkCfaQAMRZWUDbDX/JhWcca2RMUY+vEIl2y1oEgiYRYoBVeF3m5AVRR88A/o7fYWSLbw
a1VAxr0IflfKW1wA44AjGmLLYJsnI03Osxzo6JLk2MKtfTGVdHomlTlgJpooRhrbyVoLQWuVHiOg
qBYlIc8FRGKT/S6WVHnQVrfuMa09F6ME4tQ4evX4vHU2q905ydnxM6J1p5yK8MJ7qE64cyVYXX6d
V7QXcKfX/IG0E/3QXspo4znRQMi6owuXKg16cVdONZ5LCrPcgOpk+nMznbtrPwRRJBh25t5CXLI9
uc+bhvkTBXUUW1A0gstxLFT+mfFcBIJzXQioQwiWM3GwkxaB8mNGKJPD4LNYEtSc1Cz8LYe++V0d
gKsBn92JBeputRYIXR5JAXJNzMICDsYrUEpcV0f7KAIQjpGOojH4BItG0MWKk7YW0EU8AMARt9x3
afbZdAgzYNEbom0ndQFHT/Aa8GVyHMOJlVu9G1Ffo3uT1M7LWrr68FxGBS3QLeFGmu9HCBEEDXY9
ZF9jMHSOHmz05m75kU3uJfrV2ag235NOoDCP3sCLnJLioxgmlR0MoWmnXcE5Xkso3IWhn/L44X0D
v7Ha+l7nmyEhA0RnoTzWv326U38Jp61hArDjc/l/wvrT/PAPV2h4QgQbihaBGW/bdyrnGl9dKqRV
F+ELM3tSrT0pMqfMB9kGFnJaBaOQNF6yxyJ5y4dObVopuxFDfwHKdjhDxBd4QCC8AGISBOLqgaC8
qj7MvshAdeRWT5GSIFWIpM49/w85EqJ55Cbh7BWV3ggjyZNEKqsfb6lnBHODUKvzsYLb5Us+R0yt
QtluLsDQRoYX9ePt7l/r/mBQGuCJcFbksGuYOshWUX3XTnkB+DdVTdOtZI0LtP2vS43QuURIPCe4
wsAA0P38jd0g9sJFc4SUtGXImTDnEtABM2Y9l3FTNSbILWFkJLvWxjzKn5NCXhAhWpMWPq7rANbx
Vf02h/92nJAd2y9+YVMXg8yuQNkcgG0srUwisRmQqMU24WOpP1+GUAOuhV63ajnGuexagG8TkXbc
19SNx+R7KT/hM/ONkZWVyvkO+WMGS3VTVz1fForg1Lu6AaU1Vy0PJ53GyJ/qWlVHWD+vYzrHPFkP
xiaFtIET2nu5oLyHOS1Eg3Gu19xeX1DBffgDTcsV6HnvvJaDtg9D8wivuyLmlRW5bjOHYnQk9IPi
vFHaHNiL0vrmQBAtL/OxmzpBjwH7HkOtF6JEcuZxxnVAj0r8XrvuFEeOauChK8R9e3Y43Aq7RMkQ
wgSuEc7xcIJ9nwIP5lNsdFF30KRe9JBeRLxDdwd5dbaVggFGFYtWvrKYUkW0Pg6dl/JdGM1GRwDb
2PTz4WQpGWHAOY6vVOADWh+IpF/EQQ6Zu1EatOoP+HwrTknCbwPJxgsDczPN2LZhSiCOp2zQNMA0
fCN4XgBYh/egpeGIAVwWA1q3Zhi/fVrfhD7rtSUbIIWZLqQLYlGEhzCVA+AtZHmtlGqo5ET5MUAY
x34iRvODXn4OK3HAH7rl5BoluyTwrSKgPH/SFAYdA0qlw5y9FOipOqycro/V1RvSS2MdRm3mPnJ5
pR7o/9aee38TIBMOfmFbYPUrrCBlNOI5AxVxFWJ7AFYp4O4dC82tIbTduRoh6uttm5Onm17BOIlL
pcmlWf0ha1IiR8suR3V5Ywf3sLT2rasTYMUPSG+Oh0VuhUA69RfyKsuisd5GK47ZJM5BhRSgLNA7
c12Ra+QeZjYFR2NrqqGsn/PDT1kUcoE8xHSE1/4QmOAPT7AGEM7ushS99tILgRKRXmSimQgBmaRh
cTBt1ZnTyzKNhtR2LfC0g7oi9lFXMTIHPHDpu5LTuzilIF8Il6/pqZlx8on8E2IYyNl4/VQqH783
PRO8WW3bsGYoV5tAR6VUVYSZvOQlyFE4L4mZDehB7E1fHMD+h90/NsDLJWjpn93DGIGpjBxaKIR+
TpZ8Kkb+kQ3WPdnHb3Ewvljr5HG5cKP2s22D712LVo7ulpuKylkz1ruJabEkZ2mW7JNFCiI0I5hw
2QgMGAu3RTHTJzndF/PhvOqgHYFNQRrvGR/i2WQ/5SASmsxIib/tR6pDkzcMZwpwuSLRlWx0eWSo
qLc/zii7ZSd1NWSryAtYgaihq6OBpTVRdi9rB9bPJ/7af0Nb63ckIIK3kUyNIdQDU5Cmt74TvXzH
xciHnym8RZctEk+nnzGmC4L58PhfVGu4B0+AlF7I/EOyu+b+isOx2tiu37fH81nO43YH3cFqleFP
uda80iK8fOc5tiQHR/rxqJZuJtY+kEmuxQDlGu7yxaodFPbvo9Ggv/TkfA/h9phJaCWR3KGRxHjD
QDAN/JQA0YwLKhXMbjZTe/JOIpTnlwBV46zANjG8wF5QL7DUk6BFyfOhJ5CXTwCyRa5w3iUKnliS
v/t7Np5kD6LaD8X9q94NwgU7sTDn3sjhAQi0AIjMrkgefgkUD355RI6q4/QBGwtSQgDmadf7Qcln
LR9nM3ri2qj/Ixb3/8ttsvFnX0AEB35OBiovQODWqoh/2Jx3/qLAUbmPetuo0qYriaOHdtTBhB5T
w5tHuwS5wNeuBWWXQOwBvdLHi9ab/I/I0HBaVpXB6RP+2MM6trPXBdnkxwxej4KL/bJGMMOi4PQ+
QZh/2VXF6GQ1E7xkgX8zP1MRZmCtmsV9+fB0HWWiArt/LG+cgim8VJYAO58odfTOI2VGenbNomVl
udoM7heE1ird0x9f90so7sViRGu3YpEDztyN7YJiGAeuHRgvdmSipA17TdExcyob68taBOFI4JD0
pMqej/IeE9ZWhDOTZQVDHIthT4rwkHR1T31jYDvsSNpioinF+tQzHzN+T+QfVwM+BB8MHHdsxi8N
rH9lmZE1ULdfZ2DJJXizujHPr+rb528jSAN+CqEebwdGwE8MhZypn3efoXzTGCVpMqNfe+AP/jvw
zh6Mqk66IIr37GhqIDkoXtGr/9ZFpeeNa+Ku2hE2vf+cqCS5PeJ7yBVaEQ48IuvSw8OdY9GSbdRp
5m6BaQQM57WUWtqzXQNaEGpWsIID3WLwNdLed47JKx0SiEZW1bBFTCQZTHKULdhhMYXRd9kZGsPR
2X+pO/ZHlS3AXvrEAPfdIOmQiYByVHlWRcVHc7lLyDhKIv1D5cnz52JnGs0FREuv+1ldg4xGG2KP
TPp+Hys7CyDJm17RSGr+7YUJkjM66tumS7X73EQIiXnq8lnD4TNsJGBjYwhekkQK/2HQ9rwaRt8g
1zc7KbXIMmKCOtKW0fJcIDMoAxAkH3pFcIOOLlyqkgR5bibLrgasLiYNH5vtDnEHO6hHF3559JEd
zBFtO52fnXczzDlVKzeYoL3XUt134ZQHQn9b+PYIoCJlKEwX4IAVpBoGS0yzO2dcfiPO7hvDaU6+
4HT84d1zKf90264iqtiOBlrtsARO6gG29kWCdnIEZm9smPPabc7aMoEO4vYZ7wjwUntCBND6kZbl
2xR21nJfptaD2hiARQXCfFrrzbz/kdIIBpK3oKkjaMXxRGrwOlXpXSG8a6aOLrazdVtK8pws0v6x
/2K6mqGIyWrr5moyXtmmpPjCoJbqbo0shX46DN+XvtrtVHWyYucsU2wK9iiTofh4RyJiLIcMf3od
4dWFHPNKN5/GR+y+I9QJkT+hksJCrJz++mCOH8yAvIVjfMsVipp5jccIPberZOPhX1y7PzCnZHZa
sbNB7dfVDnyEMHdmCKWF2riAUHNKr/vBSvKPmkPWDzOoIexqCJyEedC36JI5/p8Pba2r37edbZH3
zDvw20AMjHxGIUcoLcYx4kqunmDOEfw1K0zzAgeyPJzSwlvq/tkve3JMYs9sSOKUjg/HIZaTMlrI
LYqO+N4ZUfegfq5XLx49Xq9BG+YrOYokkLbP77V2Jw9+1Xh+E7xLPUSZ/DHyZbFk41XDBIUX5J/a
vfz2+x7PYBkROtWvclu790BL4OmZatQNazuEwErm34/9qqtdn9Swj+I+0wLB2jtRmsgGAVwD+T20
is6nprktVr5kqO4Ek7FizB9yOmS6XCNiLFcg7MEzeiBkTT5SS5KgUsOL2EmrUTuMS2Whbl3xRu/e
xFH4r/U/OqKjxWy/Ms570VBFgnyS6vsLg8AFWd27s0nrVHKm9rLTMxpenpJ5XKGY1qZCcTe6i54w
WRXf/hNSO3pw/B1L14x7QBjBBvDVu/HmTebZVDMMVPe5T/EIq2hr1k0bA6jGpKx9qydlNu3Vwihn
bJgIT1+16hD2/yMADOhLzJoeOTAVEQP/+hq/cshB9B3+FcFxlNtXHcqSHXGFfLTjMu5O2Xjx0juu
BmY8z/EXkojqyXd2ZBWjeAbjZ9WEwGpTKPAFUSIrsZk2CvzdySbusVvKZ8nfZYA5hVfcf/PiSiga
dcbLSTq0JNA4xnCBS9Kth9mPgFZu+2VAtdzOinYUtiBy/13T2yZadQ4p/XmGGvvseSFdW1BMvhjV
MIfBwMpNNB6YarEbCvEPU9ZluWDAJptyns3mlnSZ0uxIa0bqE7J7u76yp8FqbJNGas1HlRnWO5PD
AHzm9aZ2fWwN1K/SSIijMjDjH19A3j7AqzUvQOKEwiq+JesfB5WbCOg1cGV8CYypDESpelWTBEvS
2L3xKwqRCUMp1EeqNoik/FP9fGbPQYQ+zxwm4wM9ic9tUCILOY77BjeefcCisRvaKV/wsQVHcz8o
gP+OWnldMBvCmkQgdlzwLaahXm1xPBxi3ECgbPiRy+jPQUA2fw73JIy7o5N1Undqw8PRw7qaxRTZ
ej/wbcNqg9c2p27utLU1I1MSYSzNAxGPkn8dRdy4eViF1LaaaAqTr3GX7HBmJGILSDNIe4JcL4E5
NPGNcnpbuy7pyLffNm/NxPhd/GGOA/UILCM31zZiMRdITkXZORTY66owq7bEVGM+0C5icx601kgn
m+Reqi5/+1JhRPcQwmZmp+IHFwobwXKV0NGwX1gYRQfNBgfqxS7OuOjOKF7+HSR+WfH+tPqNHb7Q
eKHA+5CqHH6niOeuUkYJpp3atobcezi3dMylgWbBEvoehmCk/rKV79rQJSl7R2F4zKOWziZa70wP
JUsq1oLFvJQdE3HC1VVlHK0CGbAkj4CkV9QWDigWJCu3lHJ6h7uRKpw38YOlUBPXoiB3e4yJUUvw
50ZwvuqgwLsr0dqqJLrxcmv7wC5CfCj7CwvxT4kuWOa8XSlFAAui6P9FnF0zCQuTgXf8AQjSDjjj
029pc20hd2iOOm/Uag2hMyVoG+HHACxCu1GcXpXcuNPIIKsCH3Ezi5NkZGqGkTlop+0ms8bbphKq
Lt+ob8Bwqr3KIe145a1vXJJnchmw8IUySnLzTpBna+MAF05ImkTHsoe+dwsYWLVin+7Cp8AgxnaT
lYJz+zbRO5QA8fYp02uHMXyPs+vLT3K/zixX5RxXUGGbw9xA+BlN9trqcxhHRLayw/ZDsBJiJm+p
uCg9hA1/p+7mxumG2sgk3bAW36eKpE8lfBOghRv1POhgMGUtOlbb+MD/Z+aAzICvxkzhjjqyhGBD
Tl4E5kDdB310rXQvgQrRH1+BGW+ARXXQmUcLlaAe6Ip9kEaJABp9DxbEk5uhmuj1kEgbUebBQc0x
yvbeJtddbHB+exy4TKy2DkqxgjgVUPBj53LUSdJsWd3riQNRIXA3xukQ6zJTlrffbWjpNXiFqs7n
E6tVZvxiY/moo5nxXEylN5ai32Ltv+JhE8tpMWTHSWbEdkstwgUmsW+2s5G6Tgz5gRcQZ6K9xSZ2
gLr9JMWSocdmxTOC9nngp/bEUP+4NGdsax1BRDU4yfeAmmIDPGMBdCAaj1Uc0Eg4l1/WIVzO0mcn
yqfT5kgD71NvH3anXir7Nui9kDTp3OT5Qgpz863IXYr1XmoF841pimvIbJ3+Ug+fSAofJEg9c4eH
bKD11dIdeNrFlCEI78ROY5GUPQL5Lz0S9wcZQhXTIMxOUcn1zP4LBthzbSzcPMHwoSU1Va2P21vk
1gzIaiFPt6bqPJhgfXvgxherECjGAR7CsZ3z7pfIEl3rYEEDuFeutfqyBICux93D6XY5sp4KHbRp
xeJCEM41JZpx2UN4jge8FhSxK/KrZ7z4d7CNcFZueTpjHNJDo9SKEY/pLhUG24k0Z1kCEcuIFhA1
zlF66QY6+kMooPzwGSJ5xqqX1Douxd1i7pBpnq365gnjlKTB6sJPmCVErPncM3TNX8ItPEL/FSLU
LZms6gsxZhDbU75rVEZIEmqoDAbKzahnJcv0BCdIdrFADkA827i6MGQ+aJmCvubGy3MDy4fatJ90
OCqFQse1RXuVD+TQhnze5yGZ+Mn2mhRZIdpVACtPLzKEH+rR2rvWudIFtKrfjoRkW0J4FzON63Pk
n9/Kozze2d+S/FGmo+2hO5qOYByoSoS4ipoyBaXDbmALZFe60prO3hn+xfs/4iEWgm1q5E4fRjfX
FyOsLIkeWU7sESrrwtyY/OHx9FWPsc2tOy14aTqQ+Blb/WKUmtVcs42EVT32LCsavp6GmvxtSoOP
zAxfZUogXhD7j1u9ni/KlLFklmgJNRSeTh/aWgrXAicMSLHWi1WRLnx3qj55r3Zbi66CRx8M+io2
NJ0NlrJ4/5pGfurFmp6Hh2rvAUPbW/tj11hn6c+wzhgbLMZ7rUXOH9aZvnoGrjF3a7Kq0SBf1vYC
zUNt3EnsKHoD9shRrq/fcV+zvBj/nCIRcnWqgNLC46AfsTgtHU1QLhrfUiFT7pddRLzGlbC+2+Zs
7ekYxmVenTB93tGJIzotqqkmRPvA6GSDzrOwCufRm6FFsjuFSQ3qy16xywPEi4Ow5arnKODziyG1
5jA/aWwLAglrH2PkQx43IIUuxOyBSHeduagULpMpLIeml3HR56UfwlZ2FHTLqX5mmqSfa+bOIEWd
d0r9rdA/GQPv/EHwO59WNTq4CqaCsc9ZqalruygG8l7Xr+30UScV63BT+74hZWSYOwk6TrfXAVd1
bCgcvxrAFhZPBWIfGQsG9+9aP9ra86l0fglq0jEU+I4r72EZmj0F4ZNSvFCfAGQ738FKEnF8JQRr
9BwmSJla1ijdU4sWxRZzXub4OdFxmVOAFUeZOUrWRuCDJZThOlLEhK/bvyrlwi/brgOSQIg5eow0
bY36niYTIGl04Pzfd/CPmH2zfVIlFOjpYQasrVPlLq+2elGXsY0YXyGCrDWWY9o7vHOyfC2Tl26t
ZTYYyRtptA2g135q7ByNi+u5y734KNKFT6wxUY6aVbHqBVwjVeLhHhNsmkpa2bsyexYTw+XcvQpT
IKIfqoeEoaciXIlHVMlNzCoybdXA52olaOd9+n8nr0Wq64PjyRdGTWz6BxotlJu2eb8DhPTBTzMl
RLhvhf4ferfsaGcWvSApcZch+xGHlIPA582OR26bHokjIJD7VRbHIvezjCje2PqmouyWvJzum6Ft
TQvcRISsH7QkhjE/FU5DTC1PbcLw9nqBtmG3wTz8M092jxh/D79xwqJ7odYk04r2Ei/ic8U4Q5W+
Jm70S5R/gDsGI7MZBm7ADrejUhQ6w3ISUTYRfjfVxXhHYxEraMAypObGN+83+cIjHogJ7z4izeer
zpfGFwJUNZago4htBGz9O8S/kdY1ZrYWEqpbXhs+outP6hOFOjPtL4XaSrVE0FXUzIWnAGMxQuqi
v3QUdIE0InKr+CGJpwahAKXNioJXgKACl67TmDvvlVyuJOm3Eag5B3Rqa6Upvzc3ho44YGci5g3M
HTIhBJcZLCDO4eeCxVoRb5VzZHwyvBdaK4RRU1aNUTPlt6rU9lHSbX8g4hdd+BlOtTh9clkms0gn
Re6t/Q6vnhNAuC6NDoVc+JuSHq8dd4osgloBe6C0ksEY37yO/2ylY5ADO17NzDrRpVAVC9MT3Ove
8rIyoe/BZVGgX6iZpLV/ShbE6Tr1JOHl32TSUN4BHC/6IqPyyDLIFkJ49CHKN1+tRBiLB6pJXKkl
F+4wfOv9R7c7nC738474fCNUYnL/AW6ZKohHKugvTEzhw6P+Qc0OsYjtXkFQJ6Gu/azsGgbr//qk
fvU2GaLjo+pYKHneqvFerDKYW2ncPl7WvbHFcvY5WphJJaOoa4LB+8Qq0rgPKxO7c6WRET7W4ilW
ZIAeE97wwAftXR+TzTbFg39+ZD6BRbGaeuMfxky655bHHq9jfq2w6XIDhrTlqEJMVCeXPeS2DUoZ
P7t9530OVVXg4g92Ddej2gVXLgDaa1BucXjF8XQ1TyCdumffcQMEZKDuzYKqauzGjjLtOD8x646Y
CzwDmCWb/wnq/stmfvHHZmkwXMHwWoHbwdYDwAcDY2xx8hXoPrUCZ6KduMQ4xkcxq3gEbaSeP4cg
8VR4N85NoY8EHTJWkMwSLRYvg9VoRvz1i34KC+d9lA9ONPMyXYzYYhJXURXo5yBvVO7H3nBJvRVo
SB9D4znrGRe488W1BYVKvlP2lQswA2x26RmfsMqvPyCXAfMCRZHnR5pmEuLmiWxPlRbOKP/vdodN
XXjN9jUXn/WXZK3nVr8koxgoD4a7ohWb1Q3j4Ge8TjB+PXn9/Xo+yp+AFtgRpUXuEdTx0Gz3yrVA
cJvjL70uEWbOlptYFDyZ/Q22vGykdlonNxX72ox2TI6qq3/z9qiOnbJE7vZKz7m7ZAeVrhUFOvdq
EIOvIE4KhOUZe4sCniWYE7TXIjeiEcQr+y9MV89YWVLBTam+zK4w++OqgUsCZwKDbBKKc/iCkp/5
dDcmacAqY8SfNtlNj3mUYfuYN455xpyF719sQC6TT2St4zWQTPCABhiXTiGJud5LGQkOy7mUmjUP
F9Yn6FBsfHaEPWo2hE3MtvmpPW1oPuxacYRaHVo/03tgu4n1xwsOjCi1atSlABsp6DoSTXZEg+OT
NDxbjh8ra/WZNXmzlZZscwxeIvBGxDOHrUpZOyIGFePe1Pw+7n09jkgNitnFAOCk3fawb2ue+8nO
BEx985/XG9MwKcgW7SqXBZSMxtiL70AEmZB2bz9HJBVHpWlN2TFtj5IeLrhJpYk8uXFp/z/dl7hC
howaJiaHe89NxXWhA15skBCtly4gPeNqDH7CMIQtyKGodQ/eTVT/Ou2dLbi7XYDN1TR0yEnobmjI
UnWCGKRcfysDUlw3l7DxLpLfLtpP6lVQvctynllp1C9YS9uUKXMhcuDPKRl/jXiQQoVpJmfwg0dK
awX+qtvweZhQ7bByZrktCBFMH+geT6gK4k+R4K6XBcvAh17g83hVc3GONFbKW7fmP27cvYDD8H+L
45E3GPngOQCWi/LsEyZJHBHqbMYzAon9TZFhrd/b0FDlXAOhWBSC/BTFPVSCZzGsshWgw7Mr0xso
FuBwAj43dv2YDH5hZ+LmH7XXkLAignQI7MuScfNkSr0xaw/SKflID4eQ6/mnp90CCUv5KDSmIkkH
SWW//K+BVDJGqLhAZ3mI85znt+VkkQ2xlXiE9PS5MWcwckar6VyaetmWjv/m72XA0nSzKSOW41/7
nDgTR7wUT/cAMRDkXB6nPfCC9UorHqJFu3steICBTyVCTRz+rspJvhuWcVhfx1hPIICbhOm3lOl9
lKBeGXo11ZJOWHZN+90Zay74r3UTU6qMGPKbuQLUl136W/sBNt5o6mU0ALcjCjNAg94lyFlWwYvc
f01CfIo4+GbcTEbjzONZgrZO2ugowiyTa/lVuWqXzpe+ComjGsmXsBXj3Nd7orMbRWmfpUn1k0wR
7VxvDtlVNCyYVuUawMb9nbiVlqV/m0BdhaE0toaHfnQLKMKUlLEm0DS9fERbEv3NdDXaPAGwyYcP
AAXpzUGO2ALBwxYuPWxbcMTy9YCt8t4vALLSkkEgs+jApENrRBALWnx1UkSaNVY59okDW8Nn3UHS
97gYWZ73hm1ffWPD+RFMpEPKA6maevBvuadk+dIBu9sJUjtfhVBRDyQK8A/ZJIDEypNPcDpcKA8R
RIxrTBGEFrlH1sCHE+jYRdASIuatviUaW4g1wQ23d1wURDbIKoYZtuLN5zxPs0imExKbkHhawIzD
R+jUkD/lys65zelO2FPwyVishegh9L0cKP+OQpdwndbJ8ZjSmjdCmFfwqEPjqqAt7dX6DXT374uo
MtnSN33Nhj2Exdo+EDfRdSr3BOqxYa6Ty/OuNO8U4CIPbCvHemESiKfsdhPAZ0HcCXzNWROGU1A9
6+BIaKgtFQ2s3SajWYj98juYR1jHYr7NkEHCJV3+5VaabxauX+psLBn4/hzU1stk8tv8q0nl3502
6HiSnOFIKY3pmLZqbASxCQ4xCkxfB7voAbV/E9l1RiGc8SlXSer87abxtZtE1H1xIKYJaVNw2pz6
QMeaw4k0gumdvsmdKKSMCSG+joGGxS3OUurSaJfxrsA4xWm6j14IOyrzz5rQpb/KsydAEGHZMY1x
4lrk5logg0D4rxyHpl1+7BGB6o++JuBM1STVIaXJdeATPjiwRkSby+d3LUUUmKUYhDveagDMYC34
1BOEj8TZxnuvNsnsa64V0FQHRGkGgCylivf8D6KflGFWv0wF5GHQ+sAS6ra+gXV0HE+auytaqNNT
rzaaLyNv8hWOXZXp101MIMAniQbBDToGGMeg08knHj3Q6W8zPFIzomy99YIc5WeFheci9gk2y6Wd
ObLVxYeCBsfyxPu4dh14n2MfCmA4dFrTKusN9v0D7JIAnJZZz7LCiNCUySBWItMXDwJVIpeisCU8
Eml5aS9FOC/pu4xRcPasyQH0obRl7Dc+htAB/BsJPyVU4V+4XmMDKGU+Vd5AfcpIn9H//E3PBkE+
VlFGlzzVoO2st3q/E6nDRBFu9Njzof0dZD/Q+lc6xwPRqb7YVp+nfBudQ7fy+0kz9nJnlstkzcI0
Kx81atErAp8IWAEqjZpMTnXmVhUUNmRSdpamkuZITDxuSL4gOcYKHTARU0QHkR7wIHMQJkeLAd1w
hbHzQkXEvU2hvUJwwoyfmul5fhiQldbyod83a90ItPMog2/Z0KXXJGDWW/TilFONpTzeKtu6fo+A
7k+81bGf2mb+kMWIXrjsvT2BLhhwhiivmQuwrSfwWfkwry3UUx4gVK1LnpxtpBCs65VhM1lSOtng
c2qR490Fm05xCPjmsOqWTxaw11ZKOKhdb0eHenMvyZPKWBTPEI3OHnoCE6p+yw7fhvF1qIS6KcdV
Gxy4pYtrjuWWDi/A/lrXY/vUKXeYuS5wS3IrjmydoJYX7gRKZ/0tLAPMlS9MIUnLapOfcuGdek0D
kj9nf8OtjHlMp6EbtwBfhIeqAZgGwtKIfLYgorGVo+5eyGIiXrjxeP4BtCUbvy7S8oDZzcIU8yLB
x/Hul5MR2xRr+SK8dn6QKYzAZUP6Cb9VxbZEL9owDieYonS2jaMFQUll+d6J7EbGxDJS5Po+xYk2
DtNdwpfiSpZZKqrql30YQ/baWX13rgczp/lg6NI2nPQyVNMbEgk9RMYIcuXUWXSzYN9j3XGJeRyU
GtWpnrwqCMVTE9WbVfTaB8U13ibXpEau85hwRglbpZhf1deEv4QmroDHpUBIj5zCqizgdlcVnlap
9fOi4T1UpiUJXItEtEhC5/g49oSBuUQaRIiuhRrpps/jTtk5qA+s5lenDMijRZY4upEitLAoZcQf
UcbrRzisJkQoKqe8UBCjbA0JI1YGwc5H7etYv4LrJab7nIES1FA/Z2b7OuijhgJnXGPp+8gtGf35
+E+8waGZWd2oiuBl8E9cdAuN3evJ++Pv90X2wz5WggQpu7QH7EeNQF+/4c72Cxnd/Cx1HytPoIaN
jeRjykXafw2m9vn1hf2JBQ6ytbzLHPyi9hgjIaeEAumoN2JHiHWENguRYeRwuhGEPGBeU1ZialL5
v61Hu2ePrX5cOnZxjDwtnAyK1t6Q1pl11OdnHZcMKssAmLtSLU17e7yIIGP2kRm9/zJgQy73VNkm
rsQAVNbkZBMYpXB1wP46FZNwiCHlic9aK1PnttV6L0iWinlMT6TmH26OA7zX65bOFtUEEmdF6+p/
VXlfiA1oZzdLvO4eBdZoEkdMtADHadt5E/78YdcEE1BeYcNZRqkamopDsjYcDrJYurgT/Avp4fGL
izMb176VGJ3Bp6tFt4NYaRwonss/Dn1jG0r5xEmhY8qk9Tngw/kOeU+lTTpuhrFBwu5YjGbidN1K
92HTdqXje2MjEgy3W7vwcamc/1UVfErdzOqwE7cRFt+zkp9/N1IoOt33EyRQV9dm0wLFYPYGg4P3
65qrOu1PP7zcFxb8s1YUHeL64MQoKXC0iOLs3Ncr+94nznGrjcIVSLAcN+xqLd+kGJ404bkIlheL
nqvO6AkPx4S+jA7fRGwHcI6dQ2MrpFkbvdEZr1Cm/uuYK5FUOzUqbB+vh2yJsmO/skIpoIy49IWs
F0K9yVf9kzXowDamnGTf/0EwRqbN35EgvoOkyuRujWl9Qe5Rp+HZhjk+UiTo0zqffK3Pys9N52HQ
53e/c+CZ4yX8GqsER3s1N1mxiwh8YJB8ezv+e3kAihPHd2h7bhtYnUyyK6s3Eq8cZ03nvdinsbOv
V0hnZ1wY1ODeO9RV0QR3f+U0Jamgd+emvNr6IOetcqRGSI3/HehMTmRJPlFU6xrFF0k88xEEAvaS
+4XyApBHwHTDwnODZ98ddMeQQK81wS3M3ii+JXUjMQbQK3PrGnC9bg9Bafp30xTYTkz+zYEws+1b
fbVA/MUA9lM+Ok4t5xxmM+r27whx8xI7M8W0Xra1Im0Wk9WqXPtA5x23DSWajiIvsB2cn2K3bUbS
j0S1Q/ch99ifrUPXuEVDXBXIZLVY5IjFv4L9afZtoryiaW40/AXXJgEPJ3UNSDBW5NPYgapf/sz6
QcjnfIQvUamw6UhScj0DneM6rlX4XkNisB7vKlhDrIw7nIH6okc+3LscvZAfph/vfoAjprxyWq0a
mIxgcwl2G1P/u7U89YAbRSks9LTGvtxBO2lZkSVC0WqrtB7vrVhkdo3wnddpDPr+/qm0mbKrCO3X
zdiRhusOYIEU2qu9bEAOwCFuXvUFYOiN/eVQzinRwWGw3vhLmRBB44p8f7ePPz2YEX0zkxGpL9qC
L85enF/DJSytHPPQz4O7W4xrpM6B1FDgwN9uBtqkP4ihWdVJwcdp/9O830ORvPxYwlhm4Mf0pqLA
sCpytzK7julcYK/XGqIhKhpxqRzGOg2OLTBWYU3OM8e564t3UzFDnDiZ/rZ2h7zmvqG2Ci8jPskb
SkpwA/aM6dxZJI0/wiENOVv4TPN8ZTXaIK6N0TCKmSGSqEJaAbMtRhtQjoEyZjT96os9dvv+njjK
eG0tUxyz5YTFVbUTyJ9Ts6UHofeuwHw4ouwPFVcAE6eF8w5ttPNjXgONiDeEWQzekdUlSHnPjjlo
lZxKFU6ln1pPtcFgCn5O0b/FgA9WOirR0C3BZ/yh47s4tsCF0VJJBd4oE0LGetZhykJtv0BLsaiW
useFKAuxuJ997PY7KcUTRE7BUJyX97hXI1azMfeYzLrOhJMQWCz0WbLQ0ZkBhgQs14+rLnuNTDqu
5aGwrn2AVWlql1DNO8yTAoVGJhuO/0RzuRXFZvhkm11+AvzGi7GX8F1dgl8BHIK/W8zeyLblsTTr
WbapgtzF9QWEOf400HXiSFVq5t1Axao7f/MxFZ1w+qRYvn0YR1Z52blHIY6/by51DaEFpx8ZnqGo
grg6OPIw2HMEurX/wAZBXoNs6qw4vm574IgUnec0yykPvsUSIr8FpilDuKc4enxX2k9Wq2FxlX75
VybjnZW32vYEieFYi4jd/MVLLEjhjSmkmabuwdW1MLg/aApa26AwI/YPsm2Yid01nbrIcfDWOy0s
XLQ97u9SG3gPNmLdExKAC/kh/CVHKyhOqPX6kV2Se2sxiIZ+j8Af5M3O2L882STaTUs6zF69qJTD
zdb3yJsfgSqj8b8b3wsMR96Msc1/5zD3I3Xr688w/O2QZqCI9/xj80MzTgheAdoNbSpMBp3L7S8U
KPe61r++BX8Z9TNYYns9Xj3cFb/R3jc0tyEs9dLBWQy3BxARcBxdRucYhTncii+fpzb9rRyaMuvL
rpxO4CKeJN5YbSPvXpeBYJGjqHgOoZRjIzjkhCk+AUBJFh+AF576q8tf6r4uMhGeS5GD28SzANNv
xkuMiacfRt3b7cFoi0vyFpnMqlivqx9LzzY4h1DxIN9bVjZP18rZoEc2J3OSy9CtPTbVigU/wzNO
e8yGGiS0C3eW0dLgIkFpW6cGdDSDuUk+JjdX7UvH9a8D51VPQQAElGIA4q1IyCbgnHhk22aHTSl5
hcGsxQRc+SvZnD9bRM05jLZmJDbbviocKna9PAxwquXURSBNpk6yYRvop3mA0wK7WP2D9xu9iKz6
8jQ52pwg/Vf5dWvzbaCfB32+AjDiQ0RwzoEG94O3aHMv2gdT1WS1Fg/fZm+WBrc0KWHDwZ3OeC63
vL9bi3tMXegS+scWXqC8phXnHQrIHKaH6pjeU3fXVTCiDzuK+3LmoH7SII2WntrqLzGToBJ1AuqI
7COX+TqL60JHpHuPgmK4CbcewDXnIMrkIcnhQPRmpMCePenX3Gki3RtdfoFjf7t582pSZH8VU0Rg
5HA6O6eXvIy5hFGJri+mS6mi63qMyMGQevRuqXJtqXUZJ/l5JZDmnR0cpChmlxpZIF49TUd9hsNk
DAY+uhLekSjWPZ5a2reRWzTt82o1sTGkgYvRdFzC/oNBDU3vMoC9AQj8ph+TRuXBlFJFaUJjHlVm
5OOYd59X6AcR4ktsFNj0c6Hs8WLZKrWRfLEhpeNCbS4rBpcFt+QQwcrFKoRrgdwz2kA+7bzo0pKq
zsoRQiOT/dA7/El1MnqH015OjFMZUs9K6GrSiGP1yIAS2//YKa32osOJzfzRALN/2/rDAoWBEA3/
pYOkGzFZ7em+Pziq1Xe5cNdNR8nYwTuCkr8iMFDWE/ar445vNncBiVPjU5qKQe2ES5tJrIvY4kyW
s9XhzOqZAsM/PHluRN7N1WSD0nQU+GmqSv/fN+JVUgGfyqQ4j8mPWaI+d4S1zxhO+ob3vK0lSXsW
ImgTpikbkVa/8A9fkiVd+Tt1M7IIpNh9wY8nlQ06QD/ZRNm+YdtOtcyMTqwlglLfFVTJKhiHlOA/
bGtHKF6Yh5GC/ApuYlrerTOZCpxRhC4DKH/2o6JrVsjtIuoUN79JD8E03Vyi/345kdYimj7IEqjM
F89zLA2JJ70TRzemdrBFOR3qnRWLnAVlDojL6z2DTLengtY6rkDhD6zVc6L50s9yb9yITxD6PiOg
8DsSSlk1OTXLzLEhfXl0XPjsnHxxnOmeoWiTq7sNWBita3urKEleSajQ8b3SW0kUOg7rWoWv0TxS
eicpHt0/eqS2IjW94NOsTMxoCtT0PfnTyrpLEBGGAv4dyTDXkkIpUOWdHcYKyf6lVkjuNsZ2Uyr7
FPdtnnWhv5H8c39ilt9hSa1vwRekC9Bj0MV3FUB/Q9scxiQ2bLjtxlYMPj0V4sets8vz0Ev25kZy
OeWD5OE5CEyNaDnoXjJOE9G++SqGdGlUX9dMybL9iV+R5Pk69N035WrXhFOgg9fvtmp+Qb1s4N+l
/SAiXvrWXaRcwAQ2orpWdtfQxmQjCbA0kPYZd0x/Tpq05dT7ovThGqVh9Tjxn6lmQmJYIzrcCk8P
DZoU1GmujhJPJOj8VlyER4VACcTr458Te5wdZdRL1+U7MKFun5LRtf2AActRtDC6Kd91dvCYafgW
c/dxDylUsR0440mDJ5uAjcE2wfyIE1mpTZR9I7NIZLiZcyCgVd25ldG0jLJbgFcY19tILncEXHD/
IgE7AqnWr49Giz/hgDZnhKLAv2+VrDC8bup6fWjtMEUj9PBJdsPmAPr8xGo0XD0QavhGOlm9LBTD
z4a5sVVAkNwBhBSXyFC+jVieb0WKsPX0mkE8XuYSsN7zGI67bYCZkVrxNKPwMkKx7XMKtXJj/ieV
mOsVm/I4ltLxMTVXaNWLtacEGhwPQftc0Uw5Onlck/Hi3wH94qMshAeqNuJk2ECeDnZIcA4JLbwJ
47xx1GcyaJHjweUNRLQGriApZWirJ7LCO7uKgrizpaRvVg7y/i04PHAFgBZJXloy56BXwL8Rayq4
eD4DPPdYtvqHf39BGBt1XqOU9td8mmpgVNIPLWfTKnrazDNcyI0WCsp9AKxz01C5+M6RjREBOaHS
tUdQI9Un8RRpSeZRWMbeebQd7e/a4aiHvFyXQ41SR+VM40JVmEWSpEDXjZ41aY6OMqAjZHHQVdnH
zU1gl4+uVNdjpBQtyHc3XyT3PS+ZaCHR4QeiETstO9/HaS3lphWCisg5QE79n6KYntwB1QKBKhgz
Xh7Y+zvFkpABzLxDuj9x3cL8cesvswlytSm2S4lH28uLGCN/9DlEZw6+Umn1IOWJVtoAR9kB/Hss
TpeazTALjG7chGGQ0rZ7EsOUX49fgym+4RPkiJFDwnnxhYtWWejnVirkjHGwwZSBwz9LMGA0HpH8
D3Bp0vgZTykmITsSDRmpONAaYVism0iKYn3lH1SOpiRxQzQG+eQfVinKJE8jHh7vFygGZ7UsMrWT
7rdue3OXOtDh80iZo1BypO8Z9oFIGXkh5ZdAlnvv061wD/MU9FLfo27+75Jykhl/37Smyt0Z8yQe
RDrbGMbG0ZxRua9ZjEgxvzxG7HvvdfiKVV3ouZJyBNql44ulbH8AoR36VY85G48aODq4TOs6bemq
Tzf2NwDFV32t0bK9ZbOwIju0ItkeGXf16hZKgyFcAsSKT4nzjTn+s0/cBUi5PyFYbGarsX8Hxshn
CsCDPGjmLxAIJ8rO4RToYrW4hRqLI5Cdb6vzEjLeNMe8T6okjgs5y7xDcOHMtvIh2yysi0/fhTfX
IInz2MHHOJQHra/F4vwKzsmv2GFuI7HJXIFamAp53KXULLEIjoLR76LmHe6POOd+z/Zu/X6iDVN6
DJCmXSO4ACLRWOuIJv/ren+fNMdGNpR6kmTgjCqcWHqJNgdXRigv7pktdcbanvs9ew7hZr04K2Y1
XIdb/UYPtWyJ9+d96WhBRys9KTKavRpo0+GEcDfHZQ1OY9LmquUKaLVLrlQCz47avGmP8N4Ja8DU
8XY5Z85c7AIM2EIJYARlrs3kEzeNRNTHZKxU2w0BE7SlWYpucXEFbnnnDell4etmRe76pZrGW4zD
b9w/2EDOWEfpDhbw9DMiY5H9VTzUTmFdj5iQvbUtKAZgrfnIQ0EPdYUYBhu0QaqZ0tkrRvurtyRa
/7UTfOpl2cjQgF0pfdUjVd+p6AcjQE8D5vOuzbK4gs0/L5pHY5munLy4qxbDQ8hMdBvpWmTz7Va+
QkRR7hYxbSQzgipujvezTiQ409/YILl7QXqi1K0Shl3QVnT59MzOGhj/pzuJZfgRaQ45N0Y/R+AN
UChM82ZYr0sgn2oIcXqTZ22v/AJ3jOvT9glRCb2ku162Fpruw0eweKSzp55k5MebQ/BAPnNynMt5
myTqXBMYgUJ0f7GQJJV/I4JY2iuXbPY+4Wn+zSXHdYD/263uZMg1ne2TS7wrDB4mMEzHSCbqBWg5
WJmGIiwDT4lo63jM4i5RYefNtWlwVunwDmPrUOB0uqmC8t1Ph2DvieKagJvJSp+u+t4BfFhPUQq2
aNxX8xCFjadhPlm05TZjxAN7XAfeM6Rw3UHKVR5YPGh1EJHM+u7Y3hKYbGnLrSWuWxuKC4+L802f
MZVx+i/P5m+puJOika5v2D6Z1WZz7x/dvJssVVY1BOAqXNuwLgiD938Km4mjr1fv20mvuh8p2wU/
ERsMyNHJlwSOW86TZf3Xa0iOuUF/5aoq9PLaWSCTSRe7NdfLR9uVFpzOBQNwD1CCCkhJSWcPYjiX
6EqGeYwoNYR7rIJP2rV9qAGRKbKzVD7sCkNERvOjAAwgchPl4BJYbgQYPONZA+jsXD0WX2fuYwJt
jlc25WPtM43B+RnjiukjJ7nFU68Cs5OSVOEPl3LT+MjxmLxoq5xQCv5H+FSC/UjjtKmVr/gWY1lx
pXVFbIBbCMBGqNfEzPXraUp1me3SgS+0rGB3iogLu7dcwKowofJcMml4BcuMuU4DSq8fXduCto7A
Ic4LG5LSRUPILaOEmwzxjt1Z3ab4LazqL1gJChxXA3n22CsZqqPLLOTe8JODG1KP60BiuVr5jCza
9fZ7glv7U8vQsTdTI1JSlZGlugKu+hoKN/7+eBJz73oiNhpL9u4XwEa3uj/ziuEbc1fkFYsfUkv0
EbYTvHkkC/FqL+IX+menO8EWh3gUb2xrSxvUFzs739yuqXl50kMasvibFKyXN+71kaiZ1G3jkJIm
WIicZ3FkE8bAxRBqS6nQIldUnnE0BDYu+T+oErxoDXDD2KG2oRJ8wRqMQT1FV+deBNhwLNd+3ubc
0HmrHQjoLa+npGHwJmFWYHrDfudCy9Crjd85fJjIzD9ICTyikQbIS/KWpQHiDge0rWPFrsLvDbQX
ngXmU8+qmKtbtP+QEsB+gXatk55S3upvkjNAgyzGf2ppSmV+4p5pEropa5lihH74tEDTGYZE5x9z
OjJVebmNXFT917zWu7KbLn14sy2G8Qly9g/4Lsp9ZZYwKfP0leB22YoRpGCh4ACndxaKtsnfyP9n
2TeXwXoHARLn7DSGme230v4zdythnnG4UqtoDgAYGWAVnRGn6m5uKYWIfo7bDExIV485OK1RfR+x
/x5K/mJBSRt0l2dKQL6Xb5jIFa40N9yDDaWr67491gHE7K6+XlCasgG0yj47XRBF0stUkvIcESdw
4mjX5baT8ngZZdiQVEm8O9ZqGaGlNalkzY1Wl1wxKOvbb3wxe6Yx8wZZ+rSyv3Tjmi9FX4ZsMC8c
+DynjCfLrZVb2nQASeC4l5T+iBQqEsJ6EWbXoQdSE8HE8RskRGjc6frKvZN9wRObfoxsJ64EkgTj
YxCgMi3XwzZeAaKzUweyHfyzaPg5G+BtgpThZtj7yqu2qjFhcAfGowKVYdRAAarH0WU+J8GexSOv
+cLwXc1bCQDx4NBO5N4ScLagoAnbdv4rkgAU8be36W8Rs5f8GcmE0rlCyT1en5kgFR9q7tEstQKy
QYFGc/Qa4myI11foDdjU+NAMD2AwGNESFnAKVGCFNIXtHnnwhMJD5lYKiUpDpGipvxiJVY1EDiOd
FVRM4oRzoXrySKTjT368lU9SEle8WxGzWBCR1b2QTo4uPNGzpHvpBSus2jdrrhS9xuY22c0Rden7
VtTL4ABQBBiKj5FTVpyaBAwi5WWBPF76iGq+5a6AdP/myhaE9uFD0wkoD6normoJ5cWNv9UKUmql
fPvshwnxBL/neXuHbrGI8aSKMoTMskyA0Dmf65x5w8UcrFPf+1j6Z+e2IYiVNDiiIxW0DPxcyg7Z
5KjWEFf4QtcDDz90CwXcz34dMpmKyxhVPDdIOBfdonoIxU8UJt39UNBp2RbWg9Bz8rXVISpK4r/c
mUHoyNZ4NZmgI6gmZxe48ZLNxA4OCOmMKVRJsxs8t7Oe6lfwmYM+/Y5sRYGUIxJuD5yRu8nIZV2B
C795Q113rzmsObKQdTrSpT/jK04T28vTx8QjvD/yXWBZkM7EtyIVkdyhtPm/iT7PV+6wLL1XuoFb
hnGDZ7K/Jnm8j3SKSD00M1AIiGQsw2DEoOTjg8afKHcOx/Or0sLa71c8E/w8ECtBO1BM55pTAHg5
o+ndZPxRaLWANfEdW62J5rtlDlVOzSn95Dmvt69YgkGB5Rkhay42jrneBm2QE7Jga09JFdF2K6Un
bXgG7kVPgDJml3pJNtRWqUaH4b3IA/ft9uSyNGrol6ybD63wNK8/UibJzOgV0UAQFkqFKrMYEdWg
Ol4b91FC/ECd1x3++YB7P6GWzceXpBWz10iE+nHwKUG9jrO89EQe3p9oa0TKYUXT+fedBAF30U6u
nFZCzQhusRtVuKrGiFdFwSiR68k9IlndydMkw5wfyn2Tvqo0Ef9lZNMDDTdJUwNeRTY3I4lP8ihP
08Tv7Hua/BjAoM+AlW2BKbhZMhrGEth5o5MxJpXB/Y2DUc4nWcUy5fNKbH1N234YLGg3KazRIirx
g6gDPoNhloIW79iSSS4kmhVE8z/xNIl69pQ7DWyKuRoHemyhh7n3rS8DBMDtRBwlP8OpAll+eFal
sSrtQmtnGq4ODf+s5GlMZCocpMVqTweOk4rcj/SZxNfOcqrElz83BtTmH4IeDhgiBco4GOcHWK/5
QfS+Vh+xm70+0ui64IX1lEtG3iLiI7FN36gp4DW45GsfXTmbt5/mUvYqasM4mn8fnPvlPEdBGv5e
sk/NkE571MwHiOUOBKGClkEufwAOlq5HIuLRRz/AzLmQKyDeEgkEXMDhmaUa+peyAVi1f706QP3J
O468cXsynnNWGb+PYHubHGomeMVoZ5Fi6SvhrQT6aAOc3VlrRaqsJ/MHwaF7ZlwY0aMwuDqGCSEw
E9XshefqbzwkztPOldRpOotEMh9IvSfBlfAfMBU72Nrw0eht0G734I8M1tlJfdrt3gGzTMZOqhQb
1HbDcEONzH4e1tqvukvuZkQQ9BlG0mI67DM4trkBcMw0CMp8r1RZtFkIRShg9dltml04fIG4YgcV
RMet4zUXs+0yxiRCjBjtbYOxqFa+MZDBiL2XYbNRyQw3oRBS7gz1mFXW17Sx8Jkm2KWfbV7WEN8s
PBj9E89MK8GV5kw6pioCwWaZJimVu8doIurTpP+CMPha6AG4EThUjQ9TpbsF+m2QLg9OTs+ZNwLx
w1PTT51YpVu62jRYafYJ1EqD+MwNLtgqzjaqSVUAd9E/prXUBMyfcg9Y6LrxjtqmbsZDO8zJTao8
SlAO0fCdFSqfk82AexwgMr+1QmAvbp4NZQGeRX5TcquIbzK8agDXUyMEEHc+1UCrGIWoX2xVYeuU
JAFGROACDlw7e5ZwH0gYoghiOqNAI5BNEMGbgWbaQyrh0u7LoP+BNl7uA/0131KmgPMzJTfnHzuJ
NhxDepLce8npspP9YEZQo1nLtxzru0esgOtRtW8OpHLmzBK10Awc3juVbbaHOozGte0VyJ2eTXZe
9OeL4ani/Bnwvzzjv8797emN6eqZdToDy+c4jd6FpHckRPbMF0NvbiZcN1ENgpsZRtV/20LCqRhV
r2hPK5O+r42Vts3/06mXPNvSGvO9dzEtTy7eRHH6TChV/ABG9QIgUcReua8NbJLG2dVI8OStrQ68
EEsOxHnMxjUHk5rO5Pin130lbyeki752Sq1wToIjl/t45jEtArZBGG+pkrmu6VvBqvrbXPH/WMOa
c7sj30vxvdESXaHC4PxB/Fy04v6vpKEwt9XVwW02TBqRdv3+jL2/CYQhhraDAQ/s5m9zLUrnJOWJ
5DkwFbdYJo9q2ZDHA+SGAKLti8aYcplv7HYynN8Q6c5WhT56Yor18Y6SQxPvx5qHHImI1TQifmGl
KDjYQUw9AicoweThRXzqy4DVwpJL/ph9p373HvEPVwncx5ukjWUf1/e0CtTcL7bGQcgV07w8Agrf
H5MIj3ViMTcXLurscZZAf+sseVtuNPop71nzVL7sL7w3hik0/JwqAeT5kI6wroh+XB6/XSiY7ZgJ
JXy6/g5MW4wb+o38A5l2/+be1UdHJcV41kOb5nUx8EZsRHrAXzib46Wf8P4HMD5MIjYHIAHnoU9e
hiRr0mx3z1+tQI6ONMQfMyFCqw3zFvw0qJ0cn7rTD3pAA62pucaQkRIrnzeg36JmcOwQ4VGrg8cv
TzCCMmpOgyz4ld99YKYgg2MFAu10u3vINRO/VK2O+ld+dKMHx73ZklUSJA0k1j/f1LZNhkiSCT5B
/wJSZIgkheScotiJBIDk3x3yeM0sc9agoBr9X3E7huF82Fbsd1Xi1dLUezNc3JG6eLJ4f0Y56mJQ
F+N4Vc96u8wEcKzANOVQhtP4oMXI2jkY0WxZbODt9elbs/JfCLknXfZhU6wayPFx6elwWCWggy1f
p3juXHZcqKrTflZR0IDay8UOjEvsXd9z55SwUiZc8wJx1f8d7B2GLb8g1M3Euf2lKKczsMLWQiFU
wpE4TN3l2BHs59pPsNd2mcyzRq+15tGqsw1Ob5I5gKqZOs5wWIYvJ5Z3vUlnOMQzN2Q140wYXLih
gipkVLaltOAJfltZPNMENcmFo+hKnfo0jPMjyhQI2DyyCTNFzp2BOI7eS5nBwvbz5dh5wlm7mNuO
nFlRZ2fhVSEf8+32+8samJKLROAzaVao440NpkbdcFpe/BmH4jqTMxBORhM7WC3Y4pNDJ5OOoOZe
NqspXQEMxa8WMmK8vyfsRpkVqe4wrgaTtb+lrd2s8CbC25J4mvFD7loAD6ozrZA2olgUrZDYm3LK
jENMtU6ZGJzv4+LHeOlLklWda5HdAeVIDMgUHYkI3qfoSMPxUyuoaUFYNzxVhGEIUfkJHMrt5TvV
9u07YaiycTz1z2Znu1HlVrHnwq+/Z4WLs84p3+ox2yqI3I0E8G5zGGAB3k9d+Q3o805cnD3x3NnN
O0K+jSMQRKXJ0GozZdLXyEHxpTmrVSUuTi7aXdKuuijjbNI1vcmE1U8ePNB6KSyOwCLxBDYFnQdf
VjR1DMGxlr6vWJsLfnk7fT7n7pd6Mbyt5yr0Q2CDzmKg0a5WyPH+/VgghhHBhpmuEYrDg1D3t6/P
ALX53+qdHw+IsZRz65GORfqyuNPFteWC0dq8uaoaXAy2cAP9R40YgQ+yRq24f8qqqb6NuhZ35uOQ
WcJvMSoUiHq7rbhugg97gtSyuYZ95IlbmK3IWhGb1qP/qDv/xr0cPrKCVgs8GlkmOYB+ZC7BgvAR
neTEfPGc0nuxMM+htdtnMLjxi00bKLSKkRLL9lWa74kiiuur8LQ9h4UkqHN+UuEroKJ1AuVlqrZ9
ThGuZcoPTJjbZJFMhMfR9RJslWi5fy6qwNczwd5Sc7fPK4EkrFqar0dB5cCApPoThzjCZBav5GYI
qSY+chRcPpjf1DzKXry25yKMucxE0EZjzzf8lyaCWx4SYJyACDVPNpJBAJgV9p9OSbLq8ljZhvXt
QW9NxcSm6UX09NBUjRhqbtQUkD3MfEatxG5wDDy+ATXebYl2mkq+LgVifqU6/lBH+eoIGjy0rhL3
947+0WEZoHTMdYmXlQor9xo7gztogJVBnB136JeB9ARegYG+5VAxQ2e1JH6RCLg0uxhfo0OJbCT2
EOVAJvLgCmDQuAqTOgNBK0TDlgxBPFhYmBQU8E4KIKjxjgB7vtMrynBM4ygT2jLVrooORQmcY3rg
mJ0ofUsQo3A23XpS38c6g14kQKl2hSBpKi8XPcznWS+huApKdPqxb++/ELhVe+zangNsJs+vVXVa
LtGOyJivHb2kpWT7mVXpmdWPbKIapJtzojKCJX+mLboLyP253fM7DkCne7tAG2JY8bUEo8fIXJAT
R6g243g8sq+ZNoCmVAmaOCPVInPtOUYieSpkeLB8HpWQLN7sjE29Cilotam/urY76rJmGy31X2Kv
7MIV8TSP8ArJAwNGUGsVwqS+CbpPHMr/ZjYMKHcHdNYmy4wFsjU76tgE3M4CheAnV9o5A7QBOdtU
FoPDlGySoRakBbeipiSAHJrlYmLHM5jvvk92IEUCmTCVjia0E1k+bNmeGpmM0FlWoAx2eiaRg92y
kO6+2eGuqNzkT95r22d0zMBWnovCPAkfAmpo2cr7j9L+Pm4b839737LNPnb8/pEI6SEclS27EvwN
UwZ9OtMrzHa6WfaTdL2HcB4BZI3CDu4wpsczG8iYrIg8RzfAu1AF/W1ICFhk5TTJdk0kNVEeuxYy
YEvD/So4BvEFLwu6ZkzKxcvgjZEE+p95EFyRjvtxtlNWzJg71DtAlLvWk4K5IxxrMCaK7s0PFUQc
TULzB7DoyWghGJWu+RtuQ/IvNTG4+89F9YP8rjNg/JxO4gZ0WoLgcJwsxXTZROI2rUNxopw+0TVc
waNSv+CFjrY1ql5TPXRogw5AJiQF6vldxPukNQpxeG3jj0sdKOpyradN3YYD2vxMDz0m8BYtu4jP
bk/w3hcbzI8LgmmTm3X2lf6kYy3L064mQDJfPPHqMT4Ozj0J6iNh+oNgoTY3bD9b/8dCRYAjBXNC
Hh50eH16e8NgnXf3ZOsHR5gpQuW4ELW/igpPOsOAm8gQnjNe3WVxhsWKcUxHi1geMcIDsZtLecEM
EmvqxXkkRTEXT7x1U2fv93bqdKFSrXceJQ5Wr55qTsB90e91xm3Kce/RnyQOT8S0SwyoysNRidcd
tlha0cJVvX6tzc8NetUActgrSUSU2EJY6ajM33joLxBxplRNUWL2S1d6BbIw87bnhDHvx4TK+e0b
ls2FwGASorBEn8PVIFaFoIgQs7Sv/nFHdBxZC1+/nNtN8HAhXi+bjKyTZHckQfpK2jXsCsI+ws5v
IeH5BaTIJ3PrkMb3eF6j/vBQB57ArKv1w/ZUT63FT3bCc55Caq9gRGkm8mZjZ+Mi5MSKr0NzmTAa
eejq69Lu6qvp8ZDalGqDkB/YuISrt73fZPgfViHynJCudkpVvr7ZkC5/bUG/t4HURN0tqWLK0NJ4
CxF8CznsNWRJobx0hp/dvOCiwaRWjXnu4vImmA59J/D/eB3KC9g5nO7rsAQ+FL6/Nu+ZezTV7Fho
8D3LbKb7UxXHwZti92szkfCyngL6r/OiM+gzvMZy4/mCxhIoOK0b8IdG096kvsjGAEXMpWMJSnsi
AClwRWwzCj4D83ulXvU/psw2pG/TSRWuqItXfV79N5VqWLvi5SDSDAGhuTqBsH7nt4Upd5hNqWfU
7AdLTAfVzK8zHttc42VHRHDiNzWexgsDYetnL/seLxvYgUZnx5zA5PIV70Gzl+fSZpM8bAwUyjc1
Fpy6ZdhZMKi7sLlhLo87F9kIqHRLGeKrojWckKydDwg6eKk/19i4VXdSB2UZcRzgZDXFLdQ5GEIJ
9YHotevn+glk4kDDHbKNSzfPoyllRD77/t6GhqG7usFPNAaQyO9nzwmjuf56tVZhpQ1RjZJwvXDG
mh1uwDqSVLm5tsGcuCzUUnyUJifu2nPJXI3B9qY6MvkUG312eqSykAOSEIPDYbELsOU16kObXF7f
rYynrOF/+9m9Xx7RQD2bT2rfF+2OPG57PZCk5XlR6lsI2vrn9nqfyD0UD78DnDO9jKkKQdPW+PyW
lYrz8r+Are0hybUjfjgL1Ta+uPt4o1Jw/Oc4EDm6EnUDCGPEsbGnRktjbWG2+1ZzUQpqLLXFqhx+
FpFE9vj71SdigsbZTs7d7wIYu8ZhJ41gb+L0cuUKZImNK8kBllxniixYVOTJKip/WHTslb95/EHR
IqozJrM4f2C1SBMTNT2Zl02nQeeBIZ5xn9rO2qrg2Sr3eIbYdSI1oJRVf/bE/C7M8BD7bGaHX2Uy
ns9BRcGKj1iYAOw2/7jkWUNku64ywWcg2T6qAaEWPKDIPcipFhCN9CmIuotklD6DHiR5KHaiMt0Y
BDpHi8dOKniUi0yJsulVtTJwghIG9ZTqFPzCVNQSl1R8sOmz1XaFjLR2mNReDbx4tTZS8RAxElNP
9cDZ802QtdkUJENwLMWDW/yg3/FRpFG+A4nkbBW34mLYmeLFzIAXl8GdtpDZa0gb671ETBYpCzGu
DNWgmF5aXCGG9KAO9+PGedfevGMMgHAKHUjq3y01WUx1GObWSLEXudg1QtskcYGX9fcriLRVryBu
A0Xz6033JBpE92WixHOfwPHCBZu+0vO2C2P+wSnbrn5+BUbB3LUTZ2SsMwT3rE3GztUIvP0r7dAc
YfQqnWl1RvJfYmJh8RSDrNGpBuu7HYY2JzXBqFDOh8y/GUG1FJ1U8kc+a8I21Uhlwdj9zNmqIlIH
8asuZrzdyGJXqDTkYGZ7/qXDVFXf/QRldZc+UgvSkD8SCahF0bwTH7ztKqQMgnnGnmbMIfAC2lKA
ieKVIXvsaTW5Q3s/n+79A4tODYl9cPwFFxXflvzKTcrNLlOBkfaSt3kEYpPhtNddG5bKQei+VlSS
Ib2qES/9Sm1K6rsYd6ih9kj+gNM4KHlGe5nJokguxhEETYy81300DaUAOAxk/ZcUV1sRd/vPpvd0
gfd1bXyTy2kJOdkJZWQFJKYPXgDIwon/aAHE+pwXyYNxlqtccj/zL1iu6vvI7O0vH/3lVMuUHAx+
asIpYzMwt7YQfz5Wl0u52S9PGGL9GFmXNOTR+SN45e76ONSYT3SerYL5L+zum6PfpoBLQ+gvtDtQ
6npBjMM42fqn+IlzVZIzkQc/NAw0YSV3RRT+RJ18/8k0S/eSNTHaZxme06IHFOWNugijO8DWGFhT
Cfg5niKMSXvfhR0iR4wac7bWmmxNw5xy5Kj+6B+1zenzI19s+sRz8Y8I4hn912LZ6QhDY/XMfQZx
dIUvbjU49E7iVuDeXcrqgTq4l8GJTuhlAIS5BetGjQWB12pg2sNcJnYx3VjC8LxrYXSWh6y1+pQa
rky00459YCHxQx0aCkvEeFLdsl0wBytcEbb5Qno1uDkgBEDfUpKP/WJFbqgRLVWBd4AI3pgZ/cun
uOr5NPH0HjWW0DCA4HM9kQSvad68q5ns8MKbaHuSzH8FC/p0lcuOX5yD+T9TnVkwbF9HkH0OyJ5c
rQqlLSXV9L9ks1OXHKfXFiZNEhq0kJZit1ngvQ9bnJz+atzlKHUqMwal8b4RKJKPvEXvq+3Z4Xzn
yY35cSTxyBdRS0suW/yuAd2EE7tQdho68KHaA00aLTzozCGSoZRY1dOs9SS1IHq5xZoyD8G5sbtM
gMaVyZi/VmsoKRKSmkxqe2MHTfDYlOLq5+IfpIPIbwRU4pTHA7HLZQISQKrWnJsHbv0Q6mR0RYLj
4jBIg5kvByyUjOqS7/DM3tVUWjsWSMGKNVnpB4EytlSKj/iWJtN4VpBTWCDH8a5HVIQqrP+Y+yEY
cfGNv7cCPTvUUcbyo4GhjKZEYcIW9ovNHWM+jpqAqPGA+HDdVxRb8zK4/ljQ8BoEVqoB8/dPQE0k
i5yyVKj27CqnNQpteAibveIZ9fWfAfk3rr56UrSHuuENPwdCtQRV4SV1BVs2daKAfIo58/lY7Cmv
lswG/Bp0Q2rn2crV6AC/FS4/T6vrfR7kRprKYniZPcF4P7TspFTfvbZRTl/TyC0GHLF5F02mk0Qy
nIclJlCG2/Phy+ZNy3XItT/XwoFPOywO0d2pUAabQFdUkJMrO8Dsl39kq0E5aCPPJAfozoVHPJZp
iaBgA0fOty7F7aMS0ZLLkO99YO96gn7d3L6UqgyO8qYw7W+gTE2mObpe3mMfsmAJp7R6VsFiftYy
rAeeLfH10jfVMCJxtllq9TVW/H5fV+Z5xuRvpdM53+mjzChlV7fFu5wIC36bCL3VOh6xMga+q6+3
CcxMLzISoUeR3HGv8gd8i8E5Ytopcu/jSeCANyiJEMUl8VGsw/TPg4U9oQJ53hNZmdRwlC7tC6j+
31V/puQeebpEUaSojpPcY12cAenAMjZ7Kxhhy4FWIg1NM9L3hQF9AGApwqpHCv0wWqRoTTo8lnLs
dUa3MvetafH19/DI1sQCqt2D8qfVmBYVpHGNbJDkkPNaXSFOwn/igduIByyYurulOPbt8KLtzxCD
WACTQ+T59Cj2CvhltBVJCoV0l1K0bB/XI1iHnqb4W5ISwKerOi8Y6fvoQClpqaaos1cRXqB5u5ah
YHkHMIGz9w9wv8lSankThDiP0fEMVpHpfmRMGpNTSZ73P1HiytKQADxb/eeSJIg4N5yX6DC+8fTu
E4sPtVE2q1BymcjcBK7uzz/ZHSOwKUT/0h7iCgAzTBRbPjc4KNG07ixbcaNF51kPMIhaPeIAFbpp
6jwnkFqwwdaUhLPrqIPmFi9H3WG03RTzdoAOLzgRX7anwQZJlpkzb4HUDeA0lZk2cQlOTUBPAFo4
oyIY9HdQr5/Fqi5uM0LZKBir/6yAOIB0uGSodkZbizT+LVN3XwIBVUJiRD2V9Qb+vWsQN1w1FfoC
Lhxt1eZFzRMIirh5YfLp8n8JHqAdzfcO6QKZQEeWfKyCVssA+SmATgpOxhWi+mtTyul20FNPUW8N
9yd3/sjpgR8vJW/cNZP2rTsDxyj1IMU85LFLF73eC16orjrBSvntH6BQ0IcYNl38/d+5mrQqk0TO
hBv/koMwtDeqFgba2rWNf0GXwmVMAabUF2OyeGhAm8PrXUjshHZi5CDIqZIXGn8I9pVn/nq8g/6K
1v3CjMbMIKXutbTqHXQC7nwqwu36rOcJYGs1qNujDxw9kWFnIZu1do4iwOE4MsLd7T4RrvScav7+
cF/mTOVpXe73tqePwOvOXwGHX5g/iFL3Dg2uxeEwu5ZQmrDefhsShRLgxIJtk/pxsCprL6g1V0Es
dIDJUPl8mP3RkDi62dIG15HGgjs2KMETzrSYqBTGyFP330gsl27noejnrCUouy78ovgCFaMZQOis
BObQllefol7bQPbx0gyR5wiWcP5DRHMth8xRTUgSACl2O6k6q8KefldOvpf8sl5NhCOfYvvy/dWV
v5EOwix5PHmJEUTkjxkQxIJPQd+na6y2kEdNQh5XOLRKNVEUq8y5cwXCLLili70fhLriYmzgkyCS
LB01QJI4LS0FPHicXN/+hnBTfX+GPXCt7PAK/aq3U+UHg36JS5t4hrAMdMpEqIVx0LsAtZPPt/I4
7RJPbDS5DuAwfL49wZAIAPG7IQlX3kP7+qpIqWKNMsuAh7200u4ZLnsQt/ed5XF6JrH++gcn8ZkE
BTaEp+2BPOcE+mz1ddyahFuxBCyFj/Jt2Uf6kdQaMfrBvBUYxHYk1RBMYMATuNJJOWgMCXvK8Udt
d5V1039TUR2cqo4ZzpXgSjET4Dqfy43JI06zoAvhB5JuyUaNnk3HW/gQ4xrK6fzYsf4PhOobjeHx
cScKWQVRpppI47/Os4r6PidhvIVF+ZyqvfdCFbnx+b/vUfIh/C6IOqh19b0JlnaovDdw55nQFtCK
Yqs/0KDU8wn62a0AJYCN8kHB86RGddXSNc3G2teQ+/0hMorANofr5Md+OtrrmXzIMLDVoGSgImXs
rquXSVIdUtyLMn3dp6QDwngAWfFRHV4+5j64TzRj/ULWEqfrybqwnMlPaJtM6PaOvdAWz2tvNVH6
dOcOD1DNF4nzA3wg+qB8LMWAgShc3Qoqw+ot7b0OqiVUVuZLT66yYQcuTo2AHQYOwX8T4PoHDHT2
OPhBIIE9mj33Y6X4neUqrRMIIL9DHKbPemNrmRVCz83P69QXbFGHba8UMN9oHQgH0srf4xiwMUBl
Xw76tWMo7VZ7ZH7JZubYprd16KE0JsFzkRt8oCBT62dffJWTaMNOfc8IH7q+rLQ9gsvaX2d8Zn1e
8FC6Qy919ILLVjbXQR0fEXXxvMavBC2VoeXNaEN+rVTUaDBSLPFb1BSIszzdPjFVWUgCv/UXtBSL
A7ZII9j+vSVaGB1PUHUSMcW6fJkwN9jCBYeOxRWrOfqGo4SzLISeY4cSSMaLDswTRM4/uIIBntH/
ZQYix6yZxFGQRMyQcgdHExbBiGVJsK+pvKHPCTsMflgQx+aOBI6ghuAqqEk+/c/nHSnXHksRCoYD
JduKr9ZNWJLwbnkq/7HIKfxX+WvdNVvmFkSTNBix0WQ9L11hlDr0KHCQ57bcRhCPWl9vtTeFUQVv
y3EaZKcni2q67sBXM9oiOtjuLwHviY91Ijk5qCZS5UC47yfvdsMwR7bd/9ZhT5u0l2SH6bH5HHwV
SBMMhndVIxPYbXQ8mbPXKjdB60RP+HLGqeBBTYknxo19BaiAMAC3faBOmv68la/geNDm0xd6nrZg
OAbpJ/HjeekyT4oS6fqeSdfdWzFzIWnw41JSddItMUHUWAXYZUrnUzLQpR8nsXzb/vlm4k8dWJVT
RodMtC8sI6rou3MDT/FfcAidn2XkWtllyX2zPJ2OKNLprFXWxvLX/8UYSY3Vt1CzjDw8hUtmREvw
DjzcEL25972Fx3tahp++6jhrjyS6f55zl/E5yy1bBLgvlrmmqvXVtpQweIXBJ60XZgU4fg5aafka
uAEdk7lPp0z7ouPZfvCTyluG1Dn9LvNGqrYgD9oFnAI+zsYUeVAYnMN1xS7eZicQez1yGSp9deai
SUXWmT5lvO+jEjQ59vzBJcCtGTbrTVMqQ6YYxDRxt5O3CA4FhvBa46gwLSKtmsfuW9lEkOFmRV0Z
0wrFlW0GoA42ROTuRcQ46sTU+rGmMyvYQKn1UbHhS+KVUJpuLYULrgJj76dNxTagDvXxx7JhuHvF
vmedj0lNfxc+8EN4gEp7rCURnS42f2lkDs7rtdj0Eqg8kBR9fHgxOMGk1S+x4P0XOWEqRMCMNa72
nr58FEGmvM4R7/iGvt1FnmCQd/R97oBRO29gfNqPxtsBJyKM4GAYgX4D+/3Cxq6k91AID/8lLCUE
RnSi176r23rUscZNo61OCTAcxZ1FzvyhehcbsVXhYyiFgOjSPYCDSvHT21Qa9UvvFhPXuDNmh7fU
lx0bZfOuz0ENxx1hyynVQlMxdGU/a0mTbtQ23ca61MV6zGr9h/1FKkw/bNVDscd6RnxLT+F5w4zf
eIYfqtZU5//SXuzOv1tPbKHeUlex3t84YRCbgf408aEWrHrdtuJTWoFKJUwp7mbrKl1AqYBMfZov
U1fyYsytrBuuvoeb9ZxhRiUWNozaRK8FrGWPGSdDHX4gt+jo1hTBWZuezKnYxuXTgeFgZdfsp9p2
Y2HwWrHFUVWreZMtvcEZJC2qO7me2u8DAZy0DPXYg7S0jhlVULqiBwPecn8BkjXobpWnq36pbm72
U9k3+4BTAdk6BFJa6m61obGDIfKVELfK4+2pjGi760m3dl/tpBxj040+uFFBe+//2pFRNfpV5juC
4agQHlQiUebDF5XiQL4CQ2TnAUJ+KSJDfBuWDdXeyTsIVA4ymgBJBQZKFtQwwqEaXuZGIhVZpmBE
GpyyZi0dHx4AGGIz0hwsikR7iGfa9O+/qbMrpBtZCh0F/oXju+lBh86QR+ymPSwgTU6356uiBFpf
femYgmJ9xHbAy8sdcLQbCqrqC/nUKy68kskWwdPsL7F0IcGviaarsTGuE99WdzgNOpwrWly/rXM7
7rjoKKnrapxALASarjlLjcRlcfWpcVR4pT7ZeUmKkQf+fnDkCYxzzMbeP/Xh8EZ08WyGA8zOa3Cs
ODkrCrHUOqbEyuTGbgT003l3Iw0vyVgts2EHRQkwAqQSIjwRd9SBf6BKcFOLuIraQAhCSZuiFqYl
OBTcyoS+KS8SGvVtQx/ecSUscD8SLWMYHM0VYLGfW+hHpFVJEx59uJUKc/NH8/jJ//JsgbGJpodc
E9Mi6QkzO3IuFZvzYGGp6jFINGm5McLvXQKYv9IpiGE1lmlxXe1YaUuAwcQQBkZbyKIB3Xf8S1Sp
G3FZO0bpblreFOD9oMiEwSyDyyAfQI5Vm9g+EeOcGzQMNMBcBLjmlXD+p296dluyNjQpO01CPWbq
ao2tVHpHD9RiAo9vucs5vjC6Kyzx3CDYltEvyNRX1xSDQXqCziBlNbG6Okl0YeYJAMCNNLOwF5fu
yMX5XnlOl359QKO+NcElwgSR/qVgJMs4Ok0TfUW370yAtZkBlQ7zOAOIG4YUeY0FLYBu+bCNQNiX
IpPtyNeq9QEz0iJ17tM++J41Wy4bDADhZHBldFWvTfyxsBhhTxZHOLES0dnu5tCu9TmfvNRmOPh8
NGDqrFZxJjSnjahCDQ30YkPZrgAeQIBtk+9gViGhoYpNzHUX0OffFmLp4BAaU6Y/uQemlxsF+x70
TWOT45NBrEFtr9YpRy0voOgyWKJdiUfOL9wi+fT+jQdyKUZTI6yIMAn+pQ98oWjgBCgRnUlMCl1K
K9o5kuSUlhKsTmzp8rN1FA/pKfTtEIDhai+KZySmI1jFo7dnhfRKXlfAvbMYCXI2kdAj/r/zen3k
fRmp6pqUe5Vsym/ICu43ZHq15mmNF8doyx5VJjNmWz7LX45hANbwqnG6d/T9ZgdRUZ/hsC6/r9fA
duONl93xx47Opd/NILs7vExSFIpYxCDPnaF3sSGV/nZAWCbJtnw9lGqZf+UXuR+1SAfWcM/1MD73
YHjkpRvIn9QoMGBtEyAOCMwmfvsJwJphu5LARSwTv672J60TYJCdM4exSgwZd0FJuqFmqbldjnav
Yw9CG8hGc6WVcGmjbnFrtlZ8e+yzPq5ux7WCmwDYt3thmbuDh2AjkpVCKyzR2Tl+Hdg4NsI+1rmj
/yKf+DJCq6fTwH80HlajpLd/zdAHR0NTfAyoOzSi5dc0czp1Vt93WfFjl+bk9+jK+r16k2EUL8sY
Xnu4v9ss1p/37gVoXKn3N5jvXNQk7jxMwUJnsB6nEiekjch6lNnIxGX8BR0qo8BBBi3HWrp+oZ+P
USmeqLsDP3v5e8zY7/J28wWoSb5kcDx0OJPkPFDmXLqkqTI1z7qSUytCq9jufyjK46SrcEVMb/jE
BdON4BjT+IiPXcGwlj9ZMKIYfXgxX0xqP8CV9xoxI2z8641Lp2yF0/B0nQJikFoVAxplmFPeik6K
HY0zBo6l/H80wlPAVzo2USlpn92hmyd/EKtd9OXghKHWIrimUlacnoJpFKIt6Ff8CeCtlb60JkEY
lBGN++9gEOyaQNqHuvK/f+0eQuSqiavT8yqC1xOsneBCyJ+4DpyDIoBE3vuS/z/vlUwP6MGTwjOj
OhzY5VYj4aYBfo17iyY0fkqnxz5v4iLYE9AMb65Isnnpy48RR2bV+9alIvrLYG+UJL0CHE1S/D9t
DtAz/GJ/tDoE3Y82LmAhTd7jr4LuqJaijFOz1oulKhjyY1NSlC1Uu1UYQtfaAQ1jCeHbGxEfowhr
lq83PjJtt35edkDCWVWvr+kL2Y1QWPC2NdBTuk1SvJjPq+7kbrmAf2SuMUt8LJN8hw2aDtBtYugt
bvtQf8SOJtEzwBnjLNiuz0blmGDlQg5xpwWjRcNuIs7S9xli+lNl+s1/6SvkW2rb8Qc1jhdiftuh
YKqq02t6dSJQFU6xYaG3C6ydJANfssp/xYiZPzXMtWDaVjOt4te+g8xHAboFX8l+zuNw6uCAyP+8
3mtdpSMWIpZlyURGiWgrPfemM9aNZ0VjxEccOTuUDW/xpFvOHAvC7KDLNWbuTaGFpREG5xZhy0di
dTHCeP+E5xec7MqF3iI85+q0WxftLP61UiUfZ5+Kn4C7juochSAoNbhiWPPpgJKxkIuJR2zNh8Zc
aQW6wp8O33Dp4OLuNz9v9uxPViU+TZ2xUALz4RHY7TP/vNVhAzG0HRyh9nJHpQHAuEAHx4InO7AV
eGWR+Ehzytwa8qSua4kF4ZpJxBwbhY+jviIe6iWzcVjqLrLgJt2M+apY2KN8r255VyB/vvfqpxEF
iwlwb36s2ofWBretQVf23hhIy0MMfCTHVuIRp1Twd6jDFHcJttAJ7MITF/lz7/1EuvPPnSVdMI4C
pk6LFPgqgPeCgwWnXjnpXWPJiAQRRaGDToEz/6x/2zPxhzGhReyxFKmIJu0yZaqWRfmroMDBVlyv
NHkSEBtLH8arBjMB+7k4MjLOnU5iXA1NsWmIhC8ElaJb2xKP/cJ1m9z4JCafCu3NjbjDykqYpHZ2
VQnwX7bzgyeKZjlxjgjSfyViPyFVJCmwVcFJ+ljWb91KyK6P6UaYpQHFbao2y1T7nS8NSmXuwKSG
LcCPz3pA1cqeMVruJwhJVzk/zFBPbBKvFjy/tcWE1w0GGkClxaZub1VnQYPerH+4qEc/2j29lODh
lY1tykXTH5g4fE1YyZ1lgd7NIJOn14IscFp5Jq3SkS8tF1r81coQiUfkfZNp0APDAbxRbrc6IsnR
0JNCOf72MAsNPUMWK4WEu0hFh5oV4wNGN5EZLAW40qAbARXEPs+h5GySkyIxfzoD3x2UfcIsuWgN
C2FyROEFFIiMt9jW0vgbUODtWLIiulUtnkA/dFRmTqjcGTvkpJ3YFIk2UvADk5lxXoQD840MIBPM
PhcFRTsAWwkDooonsjkTK71ZDc4dWwGP/AFTTqEe2oyRNkrq3p32+R+9L8zGyUKm+bytFKMYe7nM
FGNue6tac+cypPQaRWCw2cs2aZNUXBdIrpnH47NTWhjKiNXX3Eholpnv9DmHWrvwNV5f/KU43GaX
wf4PA3hNkcwDwbhGhimKsb3dHgenjZcJ7RFmFsL1skbqpU5/X5tHHNCSDuzeOKM+apcjucn5mHFu
PjPWt4/oIBp1/km36gxqylgp2z5IoDxQCTZj6rwysB7sboghMSNYze/wWa8z4Wfd+p+m6m4cZmFu
PgBqs3OMQF9pemZ2rCyCyyEcxrLuxj2qtPVhOab3sLf17cVQJvD7axU1ovO3IUoIM3MhGth6dpC5
CrfYbXDayi1U4wujXVlwrDMsvQhV0N7CHpg1MuozCvWn+Z/TW46sDi6gENUPLiyzA6+5rtR4zNEZ
lL8KftnzOHP+oYiDqG6drIBb+75FDZ4QprUK1c6dkeQF4maN1h3COz+uRdj81M9c2TAuCucME9NQ
nD54yO8Wm6GwQ7S/9iieQEVvZ5D8vb7Lay4YzPgLQjWmml+063YeN7MKIz2tRMQ+JMQ5ifm9XeBA
bVcacjK8J4G+4L5SIibncFePhOzG1NJ53uL1pvW4VR/kStGc6UuzNAcgBseGcxld+GDwjZYilyJo
8jLxt+xeaCWEoClVCdemqE6blM/HjbOqO7t4bR43cnHkw90te0EY87+h1uWLbVfKh4f2Ub3gQXkY
/AkNLdekuj2sRDgIEss0eOiazmEfVXRmgGQdyMqwGR3+X9mAHZ0xoDK51SL22lgpsTfErPzZz6IF
2WLizd94/Llr+xiBuG4VV9yGcuRy9UzvpkiX/zKYxWg70bExVnX7sWN036zH5+77E5ZF1zt2yX+1
8pLTAawbhrzZNFWK+CbOsBw60K4QnCFEbbzU4PLcpoKLLFhDA8B4RrKw6zeYTIuIShWbB4E2IhC+
/gMAnS0BfwrERdwvrBAPWeWJfPGOI5M1drd7AF967JP8SC8KBkpgVWCkZBO67aUWtTPju0jmbLxs
1/DW2AYRWhKmkjNtTBdMqaHJ/sxScXBb59jZF5gTwaJsIk0OqdodDP0X+HGkZxcaOcPQZVjlVAPV
XE1/JrMfquWkINRBpihJYEnKrJy/OgKecH0qmWYTJKNyJT1IIUa1BsHAFlEheGaFvG8mBG7RIbJH
bS3YWyMIELGjEXg9Sx9Lc1nYEMVmhpfAgXaEEGUHES9/lMj/swul1d2nd2Mw100xLSVF9H1VTCfa
VsCSh7kFc+EdCsBdMA9TtTPcPg0K/nRG11E4fWfofUwI7DkxInvbaTf2u0G2I/OIJQocFdlpoMlJ
zcGECYFyRFxmsFawU5fyD+pn2VvCXE9wvsitM40kWFTwMmxWP+sW+pLyhmVYQh78kxoaCqbuLROK
TUpzW1UL4Yhf+5b7DNcIJEMpQKvdw0INTCZYE3qnfdcQX1oDmjyqotSXkbqtAH9Tnxwc2xKeRpkq
gnC7rgjF+r1Y4KqyH2khvWgbG5Fl7HfDkQLUWZV0SDMHcWeQnrDUnoXqoiEtvL2xhgYB0zEwUmWK
TA9ufCc6bB8wBs96b7qW4vaTFSukkVUA190iKVqv5UI9z2uo1MWfLbspe7hn4pFa7LeW3yEUEtwj
LQDp/bUpeGB4p3zk39jcaaJrEZ16ro0fufy2YucRz1uNUEyadc8fFmU6MvRagxQLw2xEfaLG5VBm
v6MMArvP2rNkJjJi9JRwJWmLyoqsMpyf9Qw+4zafHxOvKfEQTRZzBVL6MQW6doMC+elRw1EdNbjD
FIwQSNk6wcybb7Dqp4hb8XAT2QS5xupCYYPuQUF+QJcfDcrU1v3CQqmOEVhFvatHNsP5y1VyQnWN
j+Kh/zxB6sJcUQF7TECE4WyNoMygDsB8OR9H0GH23V1xha6MThWA4FrA+aUdhHF5LCqS3XAd27Pt
hxuRne29b3nyNdQ/DYzWmaGUaLd2oczhue8b2PQjfzG7NVBgr0VTiHzKGwvCnyEoinoqJcgjvIDx
xNJmYlcX/LKOfzx+D3Q9mN//iL5TOQX6Yp/UOu7RzKWzBpb3ZmzFvKuy6TcTRF34UoHupKPhpFRi
6zCV6JbBCaYjaO4c303G9GKwH00XHoL3A8ZL94/cd8xL9V9GRRyj0glpu14tX680h5N8GIimS+vY
Z41jrzDwaEObX3mixa1c45ToumLOP76JiqxVo8T3FPKH9DORsudPtEDhGvLoX2/t9Gy7hfi4czzI
JgSh3AkLZP7iPnpQx0DbDU+We46gc+mAJ/ofEhuuI5fbygDNmhB1sSBdxJMHiUwfu0+HRdsZSASm
4OFOd+kaFnBeF9J3rHhiLa0AhM7+0QURwpOuK4juVcete63SoTJ/uyyoR1OyWFinMiLbG7crymFV
BB/HRAJ+pJqMyGREOMOBObo+hOsLErRdIz5o2lNoCX6MT6mpLaMSPfW2V4vMSggBdvoW5ag/oyvd
BEPoVhyORpGvT/lPT+0uvflZYw6PbgQ8aGrLSYDmIoxTprSvvYIaEcksQumhDFYMD1+9+mSx5zjc
0edrEO836tRdDZ8uCiWO8vr36RNF3e53IWjZrVT+xs5+RyvmjYgxUYdsN1EPdgGkOMLtX58M32kB
BMOH67sERecuMCde8P6QEB55l05g0xlGpdUFLpWhEUzhSv+VXL3pVnldnV1cNylW/Bd/Igjdj+DL
xTrxIyIoB4H49D/vvv8kWNBv6tkq9IeRJ9960rgszipWTIpS5uPGusnsl4MofxNLKtHBgnH3ED2a
Ra5WTt4ajRptXxGB4JlQx6/rqFApeqvhLUO0yPO/NV1wGFT0S0EsRdbCC+MitVdKmtMc6mbZNOUV
TJxyKSpXSpNSG54pL4iJTuLs/0MYw1MdKg+J7AWDgoZ5843/lcUHRVe3HSiiBggNnamn7zdTSxNV
G/+1A6z8UDfMkQeACrL26jFb05l3sNBhGjMThXZhePYcBQqLsDzNdF4aEsiDlrtaO2b+CdpEWAcQ
FV9Ic6o7wiziWXN1KdizzZ/GYjtwspTCiMx3JWwV8O2Pyv41mDVigo4ct6KmE1lVd14htA6Z7diu
Xjp/goSohI4qDsDJWhd+Tkqy1QYcu66jJPtHdo4Fi8Lp/018JPkuX6MtDpRg3MovwPlOz9bWAlh3
flV9Rqv9W+Z8hfFhrXJgQigaNRDrOVW5gzmRvCK8XJzQSQQIzoE+Xj/Y2kuZziFJtRq27nVaivA5
kH5tTWwWnjSpNgIBjqecWIZ92gmTH1LkIwxqCIM6ublkPkwBZX0P/zQv+Vj4BdaPbR1vsSSZqPq2
avtt5+qje759m6GRzlIhXSnPH/HKo+Ja8KyT4dbJY3v2KJBDBlNXWPtabhqz8Djtq4TBheHaDK50
ihF8pe7cYRJZyJ3UjJf5CyDHExQEv0pPTMziUgxvdk4M5/BKLg5aIBNtNTId0zaxvtnvZT4Kt7/n
la1TaC5dgk0KQCZp02QYjF4eE3DMLcZkvh+bJEFDOe5ecaGtOnUYEf2d0DF6ujXrmno7LTC75oEp
MwyXSfkNvqNIiINLaw1K1hPAkYIrpukvcgDeeC3c4rPYRUaOxP+8PwMS8HwDUud4hkyjRxv1EuNf
CRSO0Jol6FBggfOlVPZf3oIUzO8AwRtKAJHMrUtbAus4+fy1C0c3GnJg938M3u6B39gae4jCPJnb
0ywVS63nlQ5gzzyaprBY/s4wvSc3FICayj3rCmb5ZiiSEQ0lQKBwkZSzuYZlEfdZs/F2F30RMLej
ANbYymSc3eHbpzqxHgr4XkRVah3YCEo7OdJz7PDYHehnAI/8fY+8j+1VP3nND2tLCFCMMwnDi2fq
DV5+8bA/XhYQyIjMfRCsRT+c+XZMz9po3yczTcqU5So9nlVirO033Izl/eq9rtv1pDqNdzknTD+j
Iq0VvQSeoMzA9B71pQwvGZ1DCDw1uWmeh5f/+8LO7ZNMGZrWZZpPB4fmIeABn5EVARoGtW0vvKdO
LbHj62EQpVgZ8uxbWmxuI4EyA/vUh9cm8LyZObq8U7s+4FjSY65H2xMJ/vuvq0BWZxBINIoq93K4
UiSxiItfzSUsEZGD6f6VDweNQvI06yeYVtLPWb5a7tpkQFJI778+D515V7rE+OgvZzUg1kqAWe8C
YW/8YUh8Qk85Zj+8tpLioG8rkKANiHyxmTyRix9k+KPqYeTbGQKJ7c0Hs8jne6B1M/cVSc3OdFt2
/2JoqO3SDerniPAgenBGSk+sVIFhgkOmwtNU2nJOmMg15IIPTc5xb/s1VNmojRdFN39UZn5wns6Q
5fhxsKoUuw1HyRW8EqhS4eHxa3p6eio3yg6O60Z6htMtD4nVoGPWL6jUVzE0sf847gQvvqsIS480
8zDuaQZu9ofEywyrF9XRTxUjupBUZTX4FZgjHbJByCGWB66/l2bXAeLTaNOoPOqvz5YgGnn37M6d
XRlDW+3opP5UYUzCDVmki8qxz9N4T8yoRXvnWSDuG3vJdPBlW5ggDdQVnkb75o9mZguQRkBg//nF
CJjKF6xv3gdoYfH8fKrxLJJl3mffKHSdWEcsl8Sbb2/tWJE8hpBYr4OcIOkeN4TGSOTNaIvXFy2N
RpTn9o+xSHzduX1tyndsG7ejvPP0b7kTyH0gZPlPl7cvrJIxh3VPXpMRKA977p3jj+6MjGrmvKj2
4daCfOz5Yp8GrGiY7BVx2GXNy4ps3dvmUE/MH4efJIWBGUz50pwElxteBSQv307Pon9q0a37eKVi
drmAuq/T0O76NbPhftNi/A51bSb/4fSHXV14nufrAgqks8gQkN3PCMk6t3XLAQ5wbEQMhDH/hn/a
wMRgbMoyU+T/C6TXfXj1oOhxJrdvPBUEboght4fSs8Abl7uGRQTsBF7WEPkqm2ZqzuWH59QaEmin
J+RCJTHvZtqfZeZqZ5ueRfwtliN5cQy6BmUkrA/Czj8aTnC6k4lo9gV12Tm70hi7DJ+v9H9aKnFI
pFaLJ0tLgaIY7iyWBMYA9Z6qVA4tzUdkaTj3U5jgUHG8937o2zqSqRb4iIHXDQ8xQS9O8PzUAo+i
tC3CnzE3C0Somjlj+BfqGEDU7ZnSF40S/Xl/0AqK1gWFovC2F5s+3qu/vWzdHEEEUs2sgr1K2EZK
jZwHhV7NJN3MJ33q7phW1VyTDcP6fmia4wLhEttYemRxaGdl9ocVynFElHY2Wh2Lbriw9qeICcz/
LZU7nn7NPqV2K4N1qWRU/erQPVZmfUw2jAXcWgt8rZmhmjQWm62hjneoYc/jqOKhlPiEvyCnI3aN
+1i/9W0XJ7vaE5YEEDixyPVmB2TsC2C3Cx35Tu8A6hv669eVem37+/bZGOfed1XUk7yx+YuOI6T9
LZkMhxrso9gdTfeo7U7g1IXDb64fqnx13SZn7CBSYR4jvFewia/dBhbfPYq0LvhIMR1+3PZmeJQW
HI1+ECFkMbhnKm4ZQaqZhIs2fg2wBy6MPeWZz5MqtXdmLKIwNxwBnkxicNqK5gDIqwVJmM/PQXqA
jeq9TDMCB1IlaISxOhZ5xbcvmU9yu0u2T3va7ziDVRBsPRokOfqFKkw8R8rj5UGk0tUidkZdbKKG
fsCKidBkWs0mz+QK6EQmuK7jrOjmR8N2tVhuzDExXKWKjEizSvx+kO2s5gY54m5XwLYAeGat9zqj
RRnjZ0YB64iPjOn8ykorHOxazgA9yrw9x9PddwMmJTw3PJnF6tQeHVmPFh+Xk+s8qVzxYBjtoDK4
+efJ2ItntLXi67H2xcpFHyKdimxBK0rctYLL2AZssq+1/sPMm88W2vmJMS6JP6CYbhrPGmuK85Mn
oFhF6ehGQmoN6yKSL2p8BgrplISlLAJGKRL4qHuJbAddIXWB9+4j3oRuHf7J/0UyiQyjKsoMSXMA
Vj4G4tdrFOTsET9C2DTrYSa0ai622W6/WTRcJcorkuDBTa3Kq3b0+Iha5Yu1we1J4VpLZpWFsjV2
tNYnsrVPr/aLcsCh7EtrCkQxUPiVBkhmflAc2VXD9MeQThn7lizxqkiegHJuwKRwUzRDKVhSedjB
PXBjE1/ojFpMSbSU/pa3CQTkWk1Rx7BR8l3ZnoNBd0Tq91tnglCRoosuIYzVu01yuRoXA1wbO8Gj
ncJuiEOeU2vsZjXq8DL3btyre0lQq0G+r01ZjILHjoM41fojBFSSEQQDo6pQrchkoOYHgEIEwwZE
cTxEXvNRHYVkvHsQbowkduB7dbM7RvPXB/zHqgfXjheCJCjMYImjWfkJdRiG0Xno4gh6PflxMYJ4
MyuoCu5QGOL0cuqgzH7T3L7UB+lh3+gWAWi0NunnZcIZ5xrxyaFWaNMs8mw9SCxBlSRGZArWVFde
dZZrkgIZlR7BtyoL7BAkS4kB2w0IopL/XonhX+kU5VeY8ivnojs3WkeR7FVaTyJLQbMuSLoxQJvu
3+o9CWe1+m6oaBsP14ber8v/JHM19KIQ5vcjZwczYQ7dmoK3wrCaBPKv+rIpFidPdMPuCVdwJc0f
/IuZVpxFSTT1rbLV7QnHNBq6yamOA2Fz0YSHjCdDlGJlaeh82YWurNmVN1vp6w5A7aO/RBXjVuEv
3wIQb3DjU9RuQ3ts/YrpvkbhUFblRvxRgQNaR9HtsX8GT2mdxepREKj6k37xZ05tgpOB1Sg5ZEPg
3ccMHKzJq91FBwXgl7neXu7IB/ailRlgaQpG0eMYPoY3Gy5PpeBUEaBrODNO6JlL+Sl9t/QfLAwN
MJWuHzoUiRuzO/Sm6E4DyV1tN0USzcFy5RL/Q45kAXEV88zm9NWwSOQlCnHZaHkHHinEYCWOaMIH
/2lUMlIILPs2uMzEGYYASHwIhpUCJIKdV3DcSrKZoFbEVGL77O9BmmQrt+nToa4G385Wo2MEclNP
f/lxKPUKPcF2kKu2OfxkokLtsnsUcAZDrehH4Ram94DqCX6CFHN9lAcdKmqgwFH2a3FnacknR88h
MexL3fsOtPmI7+957F62HaWluyumIGpc8vNozdTbD6XNRQQtEEmCWPR7XywRGhKl5b4iWqjHTLHn
lAjwyCqhqs+lZvpOl4gPW2a5c2tCRONbIbsdv1KWEJss5nXKp3SRRmwNZ5Swnhdpck3fSjYtoSYL
Ho5oEboZZ5m9ncDFd6cFvW47fffWywNkkp7vsGXLjudPyniENwjOA8oDu0R2BGqpBnIWO6IbzoOX
hK9S6iNxBNg+2TbFlLAKnGqoKKKE1FrkjnKPvU6SjalWyiPhhpobzCc6Zqc5RmYXXJ3s0O7Q4Rgi
rEWRO0zgUT5xfFDZFd0KDOVVQ/Gk5GwW/VqvPK3rLnHFqNpWhwDKCY/pYe8g3543K5059tJJ7/m1
GWzXiC3RwVladg0ed9Vw/YuxezYPi6L8YgJH9VwfGNdd37At8gU8ZqgXZCIONZgb1WRuW/+C4Ahf
EnU1dyVKfF1NUI7Ka8M5X9HH8JocNzAeNRLMlDWd8qEYe/CDr1cnZ/yDct14hl8GD3SMpkcBn+Os
yFfgsWSh00KBoTm95xScLmOgGmC2mCr7J0lOyceHAmnV0y5Wy72aeH6taTUVZdHwCooeoBH/4HRk
AsuaBiiGWbX95r9a61tOgf45nESUmbxxnpvOJsvHI3wcmR4Zy5NRJvIkZ/D6WE/es3Pf/RE0rd1q
ZheqDvox8ySjl6r4qlzwh1bPAGMzGp+IjzsZVwnLBta66eaSUGZYbA8m/b31g0INJdreyxNNpKI4
B3pdmFmxD7gxBMp3R93Rdmz6IbmI7j10lD+6ROg9kc4Etw0aMA1SAb/5ExK1RXMJxZ191v7+tFT3
4Z6NChmploF/dGI45+Z0/lE0W4QzcjOujk84GhBRpfF7aHmJqwgwLX3O5YEej5fDJ/FPe3H1i9HQ
VwaBlFDI5QyBJlPQxDAzpIA3tHkoAVntZEWJshkYPXmxN/4C8BIQsT+tZ6MqWyR2qHDhSUQqy4LN
5Ich+kd9fmebRlsYcLAVRueRP8TcXs10xRxUJZVU3evyClPLCcm1ggdPrQehNdWCAUkFOhnV7CY0
ODao6V0dxmJUuEE+7smAGFP51GcaiEud391MqIURnvL33l5wiBGn+mxrFp95fM8nU69sDOGE8NjY
XX4d4CmowG+ms/cxwEPc3oNyia+D3l6Xv07BMMxC82MrL3FSPgNF3x/iofMt3z3Ukb2kar+GD/t9
BtxT3tdFO4vxuzJ0z7PibgbmEX162WGKkMBD+Uq63f3E9ZIoDLVSDm9pFmVpVKbFjAM8Z9o0DoAx
aAzq+ySU2gdJSO/5MCzh5X1GtRKSOteMfu7UPvQqQLpZisos45wD7yL2vX04D4xSNZUpYm/13An+
vN4HgQ6darTiZyT4XifAC7pFxk+GlWEhSyC1ZMF44OvNZcnmUkzCGRJTcg6O3nQIbbtCGkCATynK
YJKCij1GhRhVcXF00Z23T5iUNlWxO4AKDiEBH5MBh61AHHbY5JVRqOV4L4K9uobttmtLFnbCqWoI
EcYu9T2wKy9At2bBW84eHua7nJzGAND9jfT/A6p6nKyONJuqXlug9NFO9G11jG0+4s6xpEsDiuYV
fecORj4YZnzf1Wf6vGTXalikiFOoaiGx+MTzd+qgNCoNs2xicGq+pQ7qfQqLW7wTCYPo6ZC4o0qP
DAGxNhYHVnOqEkSZie1Sx9uA/htwN8uS7e9bDTxJAnA9EftV/k0ZgYLNfOCMFmi/01+KQWRGQ4Hl
1xvKsP1bLqJ3KwLLzAP3VsWwHfqyLIyLViGEWThu7lG7MnIQNI+A3r01OMqSwqOkcot48Hw2YAdr
YFdCpeHtoCDWxbtbAnVKEhsauuxkWWfua/SyUbmLnSC6S3r7HIM3Pv2wH/RBogj+n+4KMSE8dmFR
ORHbftphjAKH5iSPysTroozPGbUK4F4CZykQei4OtfJLkERnUcGnaQ/L6Fp3DOCVvP5eVw3AMITg
N0fN20Skl1mJPP3xKLrACCSJuPDamSXkQBLsic3ROT0pr774YyBTpU+12hBcIaQzCH/HDtK84aOK
z4qgTSXsYnF/d/WECdsfQAL10T1dANbaS7vpOnqwxqpzBB/MdWeFsJdf/ZDpJGQ2e2Wi+4hnKqzo
4dW3R/PMMjpXwjA0h6nw/tSi7K+F0cA26qE8Ts5uTrp2Fy043YIXgfS+eFG3m27ZGMNZZo0fWUme
XGqO9Ik7+plVxBW52oLpEnnqMjrQ0CSx3cn6ZmyeOrAslodxEsoVCps+d1fshFd2cYP+Px8rKpt8
ynLWBvbgk2xmMG61wNUp/xjlGZzITd5AHbrWMLvof/xyEFdEyRxAElPrR/dALf1iP22z0Os6sxtq
OvychBcX8i6bkVktUmCX5O21ZTJIK+XTdYl54Gb2Kg7js4vwzBbptjZmthrni+AfR9N3LNeqXRsf
6orZPGPzvO5JdbmznHbDXIHpFmfjzw94os2yJQDROA59V1/YIyTtEA1bKt9CBNtfKmAUCuqKrtVM
ifNfhhEtn94+5Rnt3DQbts6Bo6NKpDh2jw7uV5vs2ux/JtxvsRgav1zJpDCxCKQm255xVgvm+hmM
mqUapsskE9ecRGn8ODWBVHLtV5htH0KPlM3koJsM8gYU8lZPRaXh8SmTJdUM050e/WjB8VKtBxgM
7fhsT7zeysn8UoXyJ4JwsLEqeq4gx1XYHpdhplL66nKE053iaOflQVhLyzJNunXTCITJHU9GvR99
UQ3nEdJSDRUOcTCiEL1el+DJVnM07BnFe/datQzMEsLQB3NQAfWIU6Ez4wmRPum4KS94mzHnoTHM
T2pR+Kn0gH+VxfVFjgnSLpyqANIEGFOV7WE/ac2teHDAiJDwL6NDM7gkevndJKFKdOuiE5zxq9Tk
qE87wXI5EqNkArYfh3+7V2716cvuixUzU2G1JbU8qqDjXBU30tWzGemaP/9TZnfS4YZlUBqdy51/
bTgUGeb4pWI6ORsjfu8Y2VoJ8tz5Qj+uwSjpvwLlH2HbCwZNfUk/hx0KBgcd1R0rjE5kUgni7EdL
rAIkHVqqcSrR5Mc8FpR46e/b2GIBOHW9ymy/COfs9Wcfy0RrXYp54ke2yuzDcmU3U8r/1z7g4Kox
nneeTsoEhO4Ig1k8AWPS3V8RrD1uVH1WCnORbO5P41B4uQbJCCYp9hVQXEF+DlD8mzA1RgtoXt10
AW9BSV9hFX89GhuBTPwSHJgHGZgPeuLWsncqXNA++OAuk4aZWqjUKphaaoRX7oZ924GXGTXVc5Rz
MSlsmJY1biAfLuosjdpiDtyudieepA/utTP4bOe2K1uHl0oJyTQAM7QZf+LG//WUso1q3yBISlnP
vYxc27GLZmraGKt1VeJWWMPNPQpbidhvb5VxmwqLXaUj9iNlQjPV4FjX6zhdLzpaB4Rcrsue3ws/
O8sXbbweyCDrtzynp9HmJ7qrVp728EKNgFmHqCLV1+xDU8zDrBkPDWB1MzxvlbBTr3UiZYRsjeKp
rSaht45RL9Z5aPtq4a2ka3pJiqGEYCRVnWGFezY6qxz2bLrUIPOYA0Ce+omA78gQ7B2753JdFQOr
iuCH2nt2FKJkuWcaeXwYdpFzxFEwaq41OsESF2Gra8La+bjNg90TEIEBxnT3LVRYiFfjq2Y0mKLM
TMmulsXhZmVuR8XxN0Okdu6sctbrK5OtjPMjvE8U17dyELlAtWefZR5wiAyJWnNrqd12udZ3hQmk
3cqXNnl4AYN5nKeOCsdXzEm7uYNCE5qu7nCdHmGdUjR5y9YeZnoHu15/w1m13M3lQCBgbsU68fnp
b54VHmS5hUfk0/WE008Ey2XiJRrVbC3AnoJsrToOJOVFwliCAjLdQarq1EHLZo3Hrf8x1emDlOKp
Lt/mwz8J2d2+xfXK88SIuqMBiJ0ie+nDL4AaonYMhwxwmhlpPurBWJm9rkQY5YnToJXSpPu5EXRT
xjIZRBbHl51yYSU7l7+GoeTq50I+1WmPj0LHrWiP1cgl6drnHpiMnE0YZfryc4T9p08F98gCscaK
Aoi9t8h3bq3BbgS2BtyM0s3+kJ8rLyQRYDMGjZsmlxv54BBxWjvxvKy6FdM/MeIOsoujzFlvVltz
U7Bh0Wg2IwpEeYC32gD40Lb6i7KXwfUs5ZMJHE1yxy+mn3AEcHY/zn/3aGmsXSfF7ZGz6+IS93Nk
kZ8nB3X9ktrn7u6TnBarJCAOfvWvg4cKSnQkHCDieYyTvB8zp6xaQjBGHsmjySvJMmG2OlJCDZCc
TgMbP8/SoyjwwvjWdDVLG/zPSUaGdyxLWUL5swMnqz5OKDfe8QcryxTSGMYa2gq3uB/qlK5vfY7N
4w7JtUt9zqPGfRvbB4haqPRZ51ymE98hZxHalcCvyLfjokVYIV9bd10KvTl0dVuF8CfK8WblI2HX
SlegC+T8ZbtND0A7dlkhA6AxKSemq93U4OAw0SfiXTfnnuGUslqZM1Rsso3dBg8zS72UikJ4sgek
U6n4rZq40BcOmI0O0DEKbBr59TO1XvaIJZ9cRS2G90oqlrBUYgWhhN4amxaNEpzMtddvAUesRVPD
N9RVughYoyr0+Bbv5swwAfJT3NguaZrACcxpCB/DVtaCMsKeiBLfHKKx7u7qk6AlwGOkhbRuBCfj
irSu2ngO0VHwzCBGeIAMXVcXa8D2oXkBL6m6TKIAQeVllUOaIl1Swqo55nxAraAvCz/annCHeQZ0
Kp4gOo8oBdn5QfjQUPJMYOT7r4ufzheQhueFLxhqCsv1rv3WVAATVo4u6LvB57WxqfT/B1OMfwga
BR7H16A+zlv8FRGt66sUb5mjvuh22V7wOgusa5F2Q3wau1LSukiHFzedJaVgDYEhrTOpkm7vZnYN
5jgRCPeRIqAqyqlbZA0/woJAUZsk7r5bs6Uizt2V5rQWz5SEXIX9uRnlaV7KTTmt2sOMQCjI5t6k
MGQtzBXGCRy7DLOTE2NVlUsS3OYFpxPjERmBJYLjBq4Nkzn9Mhg+nU7ldW6KsHCwerlm/LcUqgTg
3ns+dXdUIU9r22duAM8DbNPFAJ+T52LMlF+VudWDZJTQ+4GkfHHCtR+qNx0NZkHPsTExIdb4EbwK
4tEdioGGh++PitmVkYOEmgtkEab6053pIu0ebc1tCVPNSAV6I1uAnK1QXNFu1NMTz47NnLY0sbGV
loDoqPEsZZVP2lImt/tpGEWGCy9mvGf1g4iDgfbWl127+Sr0AKttFsUyUpaZxaCfo1qNTTFGorZH
tYKBGhc3HXBG6VR2BqvRBCYXh44zOUbCB1ATrNN+uCG0MIesDf6GB1hA/yjcOBA5AgP6ttrQzSin
rpdq6pC27X9azxdI9xxMcBidaVMRNPlIAN+zQe7ltTYuTilkwXun4WDjU/QCYv6R9kP77wcXcIeG
48DxFDinVPhAU7lVTrfQL5bWtIBa3rJaTPIj/Jo2MYO0x9xe3udtzukmhxZKclgCFQwwTjqZanGk
J2MYL8UAt1FhWpO24u9kN2Xs8OVfcNgfZVW4ibJje1RxC0zxmVzdaC5hO23zR3mWM38i6XPtk22N
8x2LVxYYv7eLBvTynn+L1672WzMlyjVyl2yXWosjbfdxGwkBXQJiBEBdVkqe00YODxW2cfIzGR4J
zLPwdHdhTpa8CVWXbnqdMH9b83ueE4TDs6FLU1dXIi8A+gLLh1afsbD3tJJtmtqNOCIFWwxEjghf
gZKCAt6aj7hxcolNM6lHlm6oRDEppe5BYDPxyq/93D1SYc38mSNbOdWVaI0aJTG+A+uDB9OHS6pt
gTFZ2GVr4IWmiCIPwNEYD6wNiqx9Sv3NR45JOgZAhpQ8U4QUdh08wTzGFeOcjdOmyZ+qZvYnZnPx
Evq42lyYZbzL7fU6HdCJEhwo6Y7wZ+kt5/qLbr3E0JydltpU651LTeFCl/mBqLdJTBYlBSGcJmzW
81mNI7/aB2+HoRmGk7K9QMwO4O7Hg9f3lsUWOYeFTIHkjBdv5zRFZxSDE07nECGA0yV4d2/zkBOb
agSbYhh+XiGk2PQ9ez02alMnG97mRufKSHxyJohsUCNijdyUMszBGUnWIcnW61LrKATahUjlckr7
NJtLhhZulekJ4vLuMYq0rEPRrUsFy12PuiFYzlxqtVuO9EhzS2osaTS8ux5Yt/FaIhluXa+lGurq
UA+yli/9o6sY2Jx3we7Mrhxiy1Xu/tqyMealSjJPYXHlUaWDVQNxCF52o65dlk0DUaRyLfCQGwJM
MqCGVRZaeAAHOaafPgb8A+GpVHdY/z3l6kbCR+JJGIJUUSdsNqed8UrTux76ZDxvLUElbitx03HC
X6mWKOC8ebQMsvmW1RBAj2aOMVP1WXbpRn/pspuDrmD7da2QdmPQWA0QhUvRjoS58QMC/t/C09Rh
0XrEFz0iI27m9f7ONJt2NV1HyHJCmTiXQvBk8FdiioqSSIFEIplvIX3rWSXU4x06MYzWC8h7OPbx
WWgzF7cS2C4BVbufEy8LQYW+KC4NzrHpOxQ1XqEHejNdYBFl25FGQYr8ZBYwnld29BusyhhyIZX9
WTx2qqGdPfxHbFzWNDw8ZzcuJoMmnPs6IN6ErQiWJbn0brrclWh3WDKg8P+e+yIQuxqvE6+hu2UZ
uI0bgM0lbzKa6zTGCGP1DgxN9kFJJYjqZSygkwAD9aK/AxF4FarxuFNbwpRLlR5dg2KLmrBo0/3+
mqVh+Gu0PnY/7wUgQM6zl5NmQgtts3OyhzCd/WROuQx1w6YQ2YamwrC6/tfR+0xfuaebje7beESf
iARy8/ecowwYF8CaionqBpeuy0k2bk/etKdWO6HsjQTVhbSCS53fQmn+v8/eNLBAGOG1QwZUmzdO
+SiIdlAx4rkHCFyYcGBgCGy/5HAwlJ2lU3bya+4vZQTcklGHZGHlqXXFobjY/UQwbN3+QTcl0vvC
JssyMZKFTVE+afFFsFzCkEDN89KrMHEDImDOBCnYSis+p0jSwEOr6WfWSmEbGVeAFGWp+p1RNBmq
jKsJ5zaRB1T2np/ZcqoX6OBoWxEW+y07GND4wpj6D4WdJ12dLxjZSBuhDshlkRc566LkmRWL8SrG
IRMsT9tOJlzWAGCmJ7+HgJ4l6nsWKPSoqb9eap6KMvbX8lJVzgH7FOokOpBCt69+pitC9Immbmvw
hs3UpCfGmsCzH4Fgog4ECEjTt/F61O5uxZPRY6rnJNlcnuzizcoz4XwgbJabVyqi1Loh2XqvTsC5
XQWMlHsHrGnOz9ooINGVM/k1XSb1JILbi6VM407W3etjPRNzRaBNWOblk1lWNikYpPtkQSl+EAwe
UvBmPEEm24pe4Rov1SmqpoEb5ZNHmcX9KSx2dWNyNrGblxcJiIfETVoS24uSC2s1Yvj2B8By3DvM
2QRfMcqCFZeAb2HAgKgxfj5R5/Noyy5bY4cQS3PUsUMGD2dcY6Cd/HqmoXhd907YOaqv6D/T2Nve
CqGqyhWi2kBSlvXqaDWfnEotY3XWTn0jC0GXhUulI+77GHfYFpRyQtdUuS0hTX8mCFHUXvoN4tBC
ACBsJPBzdGbCCW6XWrn4nPAJJdRTHOF9WJ/5sd2L42IuNxQs0BkPrEvaoaHgt0vl/rF8dJVo5Cv1
D5EUEm6XmvoPproGi+XsAmeKcpZF3KD7vUvvixiJKzWQZtWQ+c1bRQIUbffPM/d/kqO1pWTxGgwm
m9EMyttlRGoMUqiHH6xxUUzq7V42HIqz8Xlht/CBn03KNQQ3c0OFbj8HCCAqz3czLFaI8o0wwv0a
bYhvzSRlyUPyUBvgvbZO1/l/o69VHLJ6u25DiTGISsqhBFi9qZu34gg0Pxk0mhnL3ESxoqNyV7ix
9iJ9s//h26qeulP6dk/4rSi+5p7G6Ik9KYN+A07C9LOJsVr4NjoZgyGs3bIbbMIewNA/iulpGDll
YqIohFSgpTsR/VIUp3lKZTSCpUW5HhDDuZiyodERiofNUdMD+b8fKQ8RR1u6bEgCuY2AjewyjaXC
vW0GJKDToLIXaL83mgM2s9Wn3TLOxtXwNGMmG+OCvBFvAqhVSVEH7BQ7m315WpHLjBt3Mjirw4Z7
PIf2iANrft+G/RGbIJY41uZjZSwnZxyMe44QxVUOERPpyayfSknaPhdjzcIvZwH/JQ6uY1GBxsjD
ZXk196Uz7+w3pa2pX8lxcmrvnqM2TgI7qFrDaPYEWJr1hsJtlI7YbzUQ3zS9vSvFc6X0CWsJh0ju
NUemsmBlcjxk+DEdTkLfD59JGyNlGoLDx/TR/oaMecNbO2F/AbQ/jJXulShpPEhPjROnnzUUCeOF
WZ59YgA4dR/0YPHAs2OTH+GzzevdkyFEoA6PYoA5a2rkdtZucHRSrkupF+nWFSMtOE9X8Dcg8eTq
xEF1mnGWTpYtJ2va52sIpMmdBvXrnPGseHzWTdfhFwKfP6WhXEwT9wTpNcdmWiFIpENlR27FN+jA
3NRgaHzLK2YYIf6PeIlocou7iS5E9Yoq3Wej2jhkBvbF8I8DM0yXK5qql7YQFFuunOXmjMds6Hdj
/jn15qay71Hvisl5N8luIuac+N8fgKPVpC6UjjuMKbXRKCaN2DjTL2zhuVB2TanPuYdLevshpdas
30IqTIl+ofSy/e5OnRq+ARszJD1A3+3mE44Bv6rZbmxC/82OoghCJCUH5PTRjAYPXZoX/ayMX6sF
MScSPo5jkYfido7VMo5sEH4iX1VVLdwKwj0MWspk32AOjjoqEIaqNy9kqFAlyQrkeEvOb9tFdlKo
PjNQpPh2GEXzVrbigp9zSHP66yjXTeln/lInkvxXZTalwuX97xqxu195jX0p29Tm2O897izOgU9/
jwsAbmVjS7VjHiw8Dq/PzxoT5Vno1VxDek8O4BbUfrj76X53iwMIxHOVp5wqoGQzQsmZhwCbzErW
ifbEQGNJk61SM+lZux6BwegvFGdRVzkHukB1O6/dR4L9MF5N5O3fCOwPHNb428/IJlKLYzLYxGz7
2IyRD+bOZD5Pd63wWUNEDZxhb2kAG6xgsO1U26aef7K4f4Tx6ENUK6EB1elihUYjSkjYTCUkwv+0
lAbGAbXrIRhK+e40w+wvdy7UKYhOhszzo5hJpPLObBtlq0otemsosrT9xc8o5kSKaLjnniGNF+0V
1dO8CB3zjdA63Wd1AostpdjXIPg+b4qPKcZI0z6pQ48JkVPtIc/iVtoT7zA3Kdjl0Npbg2eo4NkF
FF8mR1xy68VUvDPK6liVhGc5cqP9+f1WopLavhH6RtscNOYCm4wK0M9DspFkJ+QZgh5sEvUSUSy3
5x9oviYOpezw+e8w5bKe2g1DtIPyfOP9IetGfIsWg5GS+KgBIGnVpUJVrRnOo3yzt9rEYemk3pX1
tMemQESw32HoXTen/4EsriHrEKsBp5bncEunXw0o12KRN9IYKby58Y1f7wQHl+6h9FRR7AyH33o8
s+YoErHkH4ALB/b0EJrFhwpLzEXWAfmdCOSZ8zkRINISdbBxSUWGEPBQmgIivxWxOfFOA+K+FwQT
EjQIk3QycU1xUoGu+SP8+02/q58N9YFURG1exBkqNUQQJhbjEYIKyiIrmi1DqiW8nrMgsz698VuN
X/BrqFRhzOUqXBKYamL3KWshj/a235TkaMPsJjWl3x9asYabexHMCR15AD9TDuML2YnLkivsviLw
sOdwGc/po/eK5RE7bN5kIhd23S2zqghKYbjkHMdvOLVDTr7U91ywdl2Hw4MI4SqSxrWShGVREYgt
l0J8IdPXAglkAHZJMj4WKpmAEx44+J/kbeeKYbgJozouyGv0GFjTU+Snoa/rF6XMxqulfannvEXz
CRpqjcTD6JnKSaor4wKYZmuPxSswzYh6K4AdO8VvpLkwPuJG7po+RrNMWO1fXtAe81BEVauYT8qf
ilcM8TD2WGzL5h90OvTKQVMAxYJDEEzIkhreKr7an0vUtEIx+kFf01iFxZudXusjHYW7JNc76dKo
0YVJ8s0cfjTXENX7ve6kAbe1lJ0evHyIYzqod9UbJiq+2G1050LqIQg2/abfbz17rqkldX6pkRfZ
fHy3CSKAf8QA/wpeWhOTkJvH4wTjpTFbgarnbmHWE4KTOFbl3TAPwci3HWVNQInrm+S4ZXgJf7zf
tA8vikz1LCcDUsR30DmespzrQMIBlDX3xYtTy3xn0wXM2ioOIr4fSYZNoKtadjbQw34UCg890LNe
WH9cKiy2eL6q9pQ7mBkMreWILMtgUqOsHbIjhbnVJvMhE+AdIWgFiw5Qog3NKzWnXcndp5dQ3J4B
oTqNXCKDqXXy+baaXAWL6z9uB52ZILpGRuPR67Z21D3ypJFVxE8w52XAlHhw+EsBjbIZIXttMcNM
t0z87fss+TvlJvnppQDkS3LE99H3cQvopDDXGOgoPigwpv3LDT9FUeBmhMXWsCVVExenDricuFiH
btfU+RYdul1SiDhKl1HLeXHQlsWAN0/IKzLSQDiyMkVwLKw7Bk910ZHEfMiC/lOSG5hccWn0sMXS
DN4jR0lqP6P3qmO8iMlukDJSyZekbxdL/rH+lXL9E4MkEtv48o6aSHEBbv+AhihJHwpNkyV6B7n0
J7kuy6wkG5atGWJCFtpJJb9Bzc+6rp3PSe1L4sRCNN8Cxk3FAds2Vdt6f48BNqAHimJQab1WxOXu
pnf+Z0BNAs2NcpkGEzy7v9sce+9Srw96suBxky4GMfOMU/eMX+rejA0rXRQ/LikrBfJMmJpEE6gK
zDq52hORirYqCz4rfC5JtioEMHRWPrtPk8+nKC6gZa3RoLKG38SLHX2Xr9XaMZeRY3A3FPBZpwVW
4E2eO2IPP2DBTNXsA1USCCeA0mFZvmBEqXUrbIxcSPZ/lUnmAhO1bsOUVmbE1qFYaLCkeRke34oc
kCEmy14O7C6Vb5p4iURf5dnw9ZXPbMS77iYEiWYxdIIGqgPjp7OrnUkkv/a/OCvFXoe+jOVFOPRw
YfT1RNpq7E1Wrvb1fGshTYUJosbDgvS5m+TAQNnsYPLtJAQCn14bgR96pv1YiHyAda6cjv6WucUP
Ey6dt3KtFse4sVzNhM1qiC80kBHdIpfv6bORY2QoAgjstnLuJt+U7FLj5wImnYMqAwHfgHMjekTe
XB5HbglgDXrnE/VH/6If9fGjEEqBGnzeWpgYSE2rW3hsLqN84vh7bbsNjIb7jR0cFueelWG+Mzxr
QC9KJg2dYsRBx2k/4eoPDE7QPh8KxHYr0faciy+BLlEVQSiJd6UEAFYsIxJ7skndaI7Jq3BFcNyY
IJBlIQPOGuBiyy86xxWcvA4+tzoxGuqBKrzDobOlVxp5/1o+3b8Og9cFn1/0iJVcv2D6KMFIYFFw
nBKLvhrgzBg/A4faRyqPlT7hs7ixfZhx+rAgY3+167LvBa5gpJPZcGlH54RgoBIbIE9GcXpMUNgN
JZhRiFD95fLpSA2KveZ4vxHW/Tm7TQqSny85ZRPzqmkxKBeC3obNr1iIa9AkMC7/Jp42SuLBntMi
aUTyUT35RJ5wSk20uKiTste9maAaiobSH9YvexTLaG7eXBfGfLnDpM/FgN02MuXKWp1SK5m97Xit
Jy7v1wSnmBLaZt2XpKx4WxPO5YO96BftJnBqStgwx64MfbbMVIvogwL6/VAEJk+mDFd2FBUC3g28
oUsoveT0K7BLutQq4s5sIMzdaFE6e1mBo90+fcy9yPiAWIgWyJAFYylrpik9hW6k+1PM4KOvEKe0
NNfXZLHQEaoAZly2Xs7rL2fpFITov3cvFWC3wGwGrhoz6Chkm8v2b34jBsvKBD8xEQ+IhYyEpRB8
ZdkTZyTLcWEda0981DvmLul4u/Thz1nwmM13/nACOex36i85gdjm66U3eqDk4vdRq6mPJnlVR2w9
CLXb/PnwqP0tFyjYHW4NJc9gGCmj0TkQ9CmuPoU87oQsKyeqfNg/qdEL27y+BYTaljb8Pr9lf9Db
C7N97jpxR2H/NB02nVfMQB4pdr5qxnGzntPKcy4UJ2C/wx0ib3uic43N4AYhWV2GXPqlsHoJaZyw
BXPugzLJ3SygZUj/Q61PJgVvJYD5JlA7VHBOvNww/85tAwzp7JVDTjCNAvAwIDfzkAHL2smXA8kD
9TpqXiYKlueIOy6wOl32tw1ARhdpN4T/uIKiELWBiNlTynbLk3B8nOa6D4BeoWEk0fEkCUGkVrOo
msPxUZGa2qjMhXBW4oYpBinSwyRr2YlQTzh+hB2KpBlWa+wCGsVjPp0IrrZ1dFv8AJv9jSm2Q+WB
f3zFvQGhMzcVjnT0/dVilrqBTHCNTltMLzsxMfAYHRiLg/MtN8/wAZlm4N/o/9S5QTH4kLQx13NB
Ja1uYuncj3ChOWkgwAT3iLfwe1KVm85VjhF613NeY0U1qggG4akkJSd5YJ/T9AYfyAGSY4mDvo9C
n5CjGMsDXcqbCQPR5Ly6RfsQS18qCvP8P8v6ZMq0uMYskGb5nC/u/RdDOwa4ta9jpNRV7+RXyUKB
1SQf8/ePZRHtgw3jWdiVhd8IuR28eMnruEBQ+ZT1onXD3jupET5lI3Bx38+GHhXl3j9509z3noal
/IbXptj3r60VTlBmi1KmlXbL0CZCmKzmk87cDy6qCi4f3v0vhTRZ+HLqtnzhLfucFrFzNHnN44JN
QXJISEpgrFYJtqmFlg+nq0XPGCivDJ5YFHD1qJkT2toEaOKzVNb0PYNHcN3vQ/hPRnGduVEc9jFP
kMuYCBNt+/ZOuTxVPOI4TUZz4VFeBbqM1W0hlUhmDjC65ZKbC7fx49pXd9q782k8igBHZ6Rf0mCZ
n07GAviscooya87dFkh81USY1j+cGs7O/zDT3Q6bpOXUi55i2y+ZwWG0SpcMiY22gFCb7aj6FeWR
vf6GW8gZmuQbDsfLhDtzR5n8TRHX0gL1MIL9ahARqHgSF3BmLAH3ZiiD/jgPoAUjnKLpvv7sR6GI
djpTg8ZACaXKwPICKguPpeY0k0GmNI8wSZyKLF9S2CyfJKNXSvoUn4ltNRFi1vO0RwCAIcIW3tc8
xK93+Me4g0hqpM2eGihzYXeGO58VxGRPEF02UPXOWZ4Nf8d+wvveUJdazefCDzoQIr84SUVB5UWA
gy2IrwY15xN9OKn7jcXaj5PG8Q9UT3UZlU0ZNBULjHr/XffrnrTnQuaBLKm+19YJaPFZsHd70nFz
v/jST7Hp8aJohSqCfQGJlPMAQB/fwRFu5/2zkFFHkoRglFQBrsc7ivHG1q6Gk/VYPcviLEIvmluo
GUEX9mCQxA5YtOGsP8k95xlxblgUME29sK6SU9wc0jBY6+mzvqhqPVT9hd/dFikpY2B3mFTo1Qne
tTr75BwGXTPqU4JzhvUkFI8xgYWE6kH/02s3m79E6s3FSsat+hmHNdPgzq2xVcuxA94jmg6RRCig
gxvRra8hFCOG8gkzd4008IlS7luzD55NNmugiJy1+k5/s20CVvfVYfDYR29g83Z1rXOcyXUHTy+U
8NQqoB17W+svhfFX+sJ+kUPgshP460ddYkEfepWCS9JNVf58/Wcu83xXo2LKYTSM8AG61SdyL7VM
hRZLUI7+2KhxU315NbnzHIj2TnUbE7n4VCsC1LAv2Z6e3ZJa6QoDh4P9DEqcwOYWl3XGNrXTIinc
zUxOHmOCgHopcbMzA2Bh0LQhEiq5PrQ48fdO/3ba2CjOpSvaoV+wbWvItpI52oIaRjPlWyipINjS
ImzJcmi9L5+n5v3MXJHvzo5+z7YR8I5H1KD2qUfCK9oEj3vbZLbsr3yo1cJJGM8SbhwVZYlN5snx
3AkPHb3JzYApJtHnPNZkwNQPqwUh903pRZI3XScf0otIFpj/dTBW1pQpvZP6HWNAwdJelLYfBzi9
PAnTUzFXg6iQiLWARsX6EH0gsq8zzR6dM4yjHdnul4qRFtFo/T3cltWlOMMtTxNtWmtrS1Xe+T0M
bV9tdrBuDK3jONZNY1JEkScQ+v/OfpCVPJIwblzNIz4gNvxr7c3a4+Thtwhwbasxd66KG+/FuJ/t
NRxzLnt8j3kbdbcG3RG4A64HQxg5zpqcWHaE0qFaUJWFwkhQS9BZvwqMQfHpCURpSAARkaPMTE53
hclpXsbFje2LzTbR6Tk19gJGX4zWtt0jJYS/4gd0QiPbXoybYV0rbB4KxeOwF8HpMkjPolRKh+OH
+l81AZ4iB5MehEzz/WO3djSfHQC3kL+DGBrQ1JuNNEb+zFKgmwUaYGNr2h9v+sUP8aE5MdOY3e5M
9HAF3JV8So5qXQo/tk4jPsVb8BoxyoVs4b889YFLeBhWR0iwvJ/jUKOLylTmdlHeEX5ge0myAalG
0W+pfNxQVJ8r0Pjw+1+AL2de0q5UUsmS+fV0mk63o/eEMx6k75xOnprnD4ebA5FYTDARE7vzIrJY
q5Rl+iygs+cXXcfNLExAXE1MoBH/GdOXG5DN7ve5qcRMqepakbzH8WNkHNmVdLKWkG8UPmgXR8Vj
dHdoNspvO8i2gqDLlfls6pmQkspXtUYVjUTbwdTUwteLoHsu4RuqZM870IFcLNMWe6zldwOwR5dX
BnN2IzK0AYNRZ3rB1ZfnxUQUp2lLCXInhxHH0uupc4UFWD6+XPgteSG/SyIvpsDHljVLDg6U0lvq
m1kW87MOVpa7EcHqRGs5KB8ZzXTxmNx0hxG0wW3wR1PcliAWxig85k29WTKSFlk8iamxtrWVVGbE
5Lot/yAznvKkAdJklw83i4o39g+e8kYfuaWfulL7CUlWvie2+7xk4ukORZMJHKm7Rx4is3KOYFY/
47NRxG7ZsNZ9WO5cZycjnzjj5qVSxd4QT7rfmbOjxNvdahXlFOD/tcLZPfXoFWr4wbUQmaAX0+rN
8AxjV+ITTdVj9YAWh15FyOVA1SKXsaL5JenlJeHXZz88H9U+Owkta6gJq9BC2b/o63T3/X9EB6su
12puE7EjSV7g51sn6hzKCTORx3o+w1uPYrp7YflHU439TPeEx6RQaydhnzbOjb0O/Y2/WyL5pYSy
eFjg+7EoPT6klszjBc+vYSJW9djwAW0/JnDRDy2+znqJd1x9c5HWJsRxE2tBH0sULeBSMwLAzmkm
0TMOiXMzZ037G+KH0qNlfM41VH2a/QkkjkDMupXED/snZ/7YiS4pXxgcQ2cMdtgz+FAJi6PKieyd
mcE85tOhtl67mHIBgWPOaHpxd+7RcBv8TR6/f/udeyz/Kz519GQ7Ey2Vq44VyVCSGJ2AspbOUmUC
Wd2EfDoXwXwMFJD/TX1z83E5m1jYnitIOJuyANgNPaU6w575zUM/4QkIpbLXV+EIJ1fVVtzVmmJR
oyAO0QiEdj+pRAVfrDkxNHRjYmNlGkL4Is9AE0uMowlvavm3XQtu+yonOeHaz+otUp2W6TP5Jnat
T2dhPtOD9w1VL+4ZrFQvSk1nTO7oPChAFCW8gmDK+gngoSV0Q7na8ZWy+U0FANI/063EQkP9qSyK
i1Y8EJKjpP/hhOU6EAS3vOLlKK0iOlcbEnt1bK2mG8M7beDZ16tIeVM77NCTtAUGL1+R8f7F3/uk
yRlOAaNWTNafQfr3kUzoOO2e1ZNHFB3hIF1RkaPVmxpqIUMawlCQ7lteu3qnqLXBeHVeNYu6vvN+
KaOonrg0BmBHw6/Yis0snWUMoSSwIr+5OQbke78J2AJOzpUfa2Fm5tMCgd0FGOOPl2mUKv/OcBJT
gi5iSu1Hk2/jVTgHd3fcATKiAuTUb9tvBswLeo/hLc3pXCxHjfA6opfCi7EvtIL1GKXnxBrlA+ZW
XO6OFp+RAvRUxd5NCmyD5zrcfv3qPAt47C5pAvHxlcGFNUBHB7TqIFmNH6p6e/29rGJNrti601lV
9kJRXbRcUjvL5fTxfUcjV5IjmZjyhLSVVmbPa0E2Py9HOYCnL4udrq7th61uIPkkMGP1J8VEArEm
NHhy65F8RR7XBscsfV3kOA6bbBTUXOdbutS2zrF2zUk8YLZD3UaGNawQeFg4oY9n7dHyPTe0zxzH
Nx7/V7Eez9hjGkQ2kNXMyrYWngM6pSHU8fUtuVfP+eVD6FnKd1tJr6z4l9Rh6QFySe/RQTZ6WBbq
AFXzmbf3zHhJGbHiBKTKDHskM5LtXL0yNuNd8nwPGq3JzR1Td7GY2+RtINwBlBDEiKjQ4kXCUkWL
JT7x9GEo9RtnMQ4hLK1clVXu+4PLrYCrGmMgdGaAzrK6SFDJK2xcGysJ7iVKxGhrl7f3HzNLFtNN
xAkMgfy/uKEe3ig0I1/OG0N/4g58CmsIVhIDEv0RErd+vRlSVHBFyty/As+N/JVs1GrIJFkcuJrc
rXxH494hQfGsTRZNAA+k5t+9+ODMeGnBczKJKkeV4V+BP8IxWY52Swftc7+NPP7dyXX4UEfFfvh+
yNfqhEklQfTnYDvvFWVpi0clM0ql3/E65ZxKdMLGRsKBjr9/dN4dHv9pfIREYBVWG9GC2ZEYxra8
xjkn7DXy0r0my2kROAHZOG16n2EtPHYJ8psW4jvfq8/TfC3qDTB7zkAWw5/LdJl6lQgX3/4B6gI7
M80n+WSQXrMXedcTXe3TUygVP3UvcOVPMv8ADhrIOjmxQhu7c4AmtaMc0W8jDqV6BYdjO0dQalMM
KtACBuP+yC6nC2jn4BWfDnF77bhlAK3RcOezAbl2irAGUL6ul1mXbJaI3iwkcSM3CJqxk8Rr5uU6
P9Az6aoSLJAcTghiVmQh9bJRmTWQMqzX1a5+sl+wUxGEq5Cks9D2NM+yV96y2uf9OYKRG8UuqtG7
42ygsX5pZAvXJ31/DsU4fbhXLsf9xgb28yS9JCpUpQgLfRUFT70ikWlfkdhfFcgezUG1mU3Y9wPH
r9zJ5jMxYLTO672643jaZxJx/kEcfspQeU698ZsokKY9h/Lssp24tknTPclU6V07sKLHyokwAc47
DvjZoCPdIFIYUAwENQC2QVHjSn0BxXM1CdLlFL01vZE8WI8CcmOTmY08smdH6O1wFiQD8v/t2Q6e
6s5tDPRzNxd/R02lJa8ijbXCrl2WQ6orQ9QKTTCe5SLLuNd5fXPeEyPA1feQZIuVs2s9ZVhehS2K
i6jhlHleloKGP7uCxJY2CtfqMAbgdvd4BVg9O3yBWA6LL1IkG7uKbGQ8QjwmySWQnMfEJK6sTcZV
Dvo5aYbbk3aSrdREzMUrt0mhnE/vCFUi7PPZ22jeW6hid0u6j6uMU/hZzEv4bX9VE26+RFq7ylG0
UtospxXzamvCEz22voLKDb8QjVUDanbWbyaYnUqtk7Ep5asCgw2FOe7BwUz6++TZX1s2iuVHLTlE
m2VlD26DSlfTkmB4Sk1eIaBekgA44iyngEopT1Aq+RnM3phX/yoaZOIhKvo23kC4RBHkGs1xLWOZ
NaIQdGHFBwgZ5TRvA32U4aBlkaX8xhU5R99ekslVUydPoKKkm+gtQl9Dm+9677AFFIrp+MVugeCv
CDlrw7wFtZyzpboxL3cKpEv4KRRQUtmPANLD3xlW/ha6irXo/67lHSVErm5/UTNauvWy2Yh0bE7E
QhtjVxehSe51uWiICG4/6yjoLKy/23jt/eJKtvRi5KhY2tm1F4/+e9fl2e0S7ChH1yxWOqbwLFF/
KXKBBsFEeDOMSVbTDKRKg78AU8OnVb9r37Hh5oDte5SQV4sLPl0mhids1o4/Xwgjqa/ksBFPZhQf
/QAOWaM5clB79ExGBXYOiheJDZ9FK1rUx/qac69wStAXcIroqxMm0LfPvjVJINtLAMObEZAEbtWA
iJNqKlbLA7Tqs+h5HcREVUDZUwoGpcaX6Y7GwdaJvLbE3JH5Mau74v7q6PhxIwDErSqS5NTtsaPW
D6QegFSSzfqlnxcquueNkJ+MvSfVDnQdgf4U8jUWlR5gmcz1YaKzvYHK5cV4kbsuWLaPH9wW0V1R
n81WTInJ8CBBMOiws8E5PthAGoNMhFX/GaEIGbsLRLx3w7OsyUk82abUbV3Xn7KKEDzHH+aTn661
BkYQECOE/R6hurGgE9IkfLFmnX94/tMt0MB1CB5tpgLT0ypXPmKkXcHsVtG+jEYKvT2RXCcBFHDi
r3K5w7IIjLGu2BsCJYWJy7SjcBSFxVBhoFgRkzy8uzZ3H1CRubw9D//YUiVsr4k6EgB4YdE6x/2i
6aVD/Cy5VJbdovcA8orlRH1+/mO6eiBGc742cxdg46vEBZ7csSVqxdEq+VGTApbjDV2g5hkP+sSh
f6Vg+i4RSVR9qNe+aDkoXSDiPiIc3ESN9/gNNHJd1/od9X6Y2ja9n+0wjC18n2WEbaAmmVnl/jIB
V6xlafqAjEnikgOT7BS19XAv9Y9UjVwtR672lAissXOb3CjTNCIVGvyJ3Ol3goZBZYQ1VIiEjnKc
inZiHFyKvESg/nIcWy3DtaQPoCGIAR58kpRiiB5Kdl0Hxsf+9wcXcaR7U0ZiRjz2dPgb32p1MSkD
g7Or8cYweBx/ACuc0q6Sle17evOot4B15W3Mga0y2M8wWJkk/NV79UM1CMANsDBnsrbMjJpSDew4
lbasis0v8cS90DR9tBcoB3pcqI5g2s3D0Nru0yYF4KOFBSn0tgDm45GETLhCR4coGX9oPQSCmnAG
YeuMMxykiNzD/YW7w3KXEnwZTOF6JqsDktdBZbhR2JgoKxH1Xb6sySG4YPk8f+sIgiVH4YYVBGRs
WMtOkpxYtblw8Nisu9zw3Cjp6Pqf3L/pQmQdwCLXpoNWpI4YyyklSfvA5IGx6MIV6npXLr7G9cla
Hn61wLF2RSuV2qYrn2MA1wMl904lKxnn1/E4o3skCrWbtNrAjigkjQFuL9LRUSD7Y3Pu+F3xp1Xl
YUlcK0N3b5F7WX5W8ZeaxxeMbDo/9vXRwrnW6EApRq3LBFl5xIY9MMEt2gO/liW5o/cooBEyK7W6
2jEQMy+ab2kCo9iOm44m3sRxZhO4kHuYQ+hVb9tvarg2geEoFxd31Rft6FDsKlGCvsy3bhh6gsmx
mwzBp/cn/jPRlFyPCXHcvWHgkbu0qvpeJ+f3CSoU6aaw2M3xcAFp9u96Jc8afN9nT0t6QcNm7AUq
CHLbFqrdj6VxyP8P+CdzCqasFMxEVhTxdXenjkMgguQxq+UdIwJu90c5jyXiFKRIkpbOGFfovtpT
MeZAJ+7enXzdc7PfijeT7J+Mfj3DYAGqz54NkeryPZgBUv2+Cn3RyzgD2JLVUVKBZ3XUPM4fVKYD
mx/9GSmE1c7l270gQ+vX3TN8B+w6/LMoLPdg+5F9sICkPX+uFUCbbOJqfRS6L4iDkgsl9IVRokNI
U5coax8jGjajYgAjeRPQM9XxRcBoP/Lkrsp9Tf9TgiLiXUDDZ6r87ZX+jf2XBCLvRA5EZCY5AhSX
sJcA7Dr+3sx1Wz7dFkzWF1D0Wr5dGwiBAYb+uaGLL8vqx16Urij8tPZF1pGAUuwiS/mDtxyzGLFp
NpgZ7XjmusFj0RZ1v1qs19fEKsIRJZhnmwG9nFh5/LMWq+gRAJh8lFn/1xvVzobg/giCRShYuojW
tvYi11RHYuhoQOrEj0634e1jXJSbiZcFLVUl8VhHcq6JH3WgcJrsukWuf5E06FPt+Is+g+Gm0aAk
1dr7VIvo5SKKoG8J8Jf2DwD8cDcu+TpBNa9TSRghoHO1xgT82C/OvEZJkp5N2aUvbDDdyq69s7vs
XT1HIlFSNTjJbu6oU1RpGFrddZkyPJSt9F1xlq9o00MxyIFd7ioz7lulIIjx6d365/dQ1ylcIzAE
VLJWO1Zfxon56La8CCpxA7GQiQlVCeIPpTFDajf6KOUZ8RW2nU8hbQwItxB3/AG/AlzXpBD8agpm
ZHOPqNIyiTxmBSqZx0N9PUM7xu1+aX2NLWxk/d74CyqjASk2XwFXQ1JGWcIiRLNVkuWzF6Ul9k1r
9q18smJPE6NLkpngCHMUlhR+dyzMTVRM6fcXwSh0ssLp23f2WcUeJIz1i3SM6mN3/jyXIiZPITKF
nJUs40SEg/2LxtZYtalM9pio8WTF7049TvQnRzHw1IF36fe5+sWSI5Bb/qDF39xkcun4yV949eVv
yIJZ95veuj7eJKCDHOO5+0MyJfXWTfPYPat1zBtBQFSNJv0fjazGcEkXfO+1Vl+WvMw1zM9WI/XK
4FSyuY4UfoygvaoEduHNexy8eWdtze8OvzUx6ZyTLWPR9hfMeBW7LPOZZKqYu0UlcCRcWxMTPeyB
FeXN04nNagRrEP4VRK7326FfkctRzOHV+XmM/XH++daFbFYU/HTHRwWVvcvDGE7LCrkRMWlsyeWE
N+1/y4ieRh9e4dvAHyTbCZ2R1Z60DS5D4kNac2BxReOrbvr8wN37UJIz7jwNpt5zzAlmR84gWsgU
80qmrBTbidkY2eR4JFFzeKEP7gai2OzOmYEOKsoyL+iXRntDt6FgZUctB5gneUt3oubNNdc+xi0d
DA5ylZAhac5ES4y5Dmcb8ZGVPRsPDV3n7fDvamNU2ta1nqFi2fE4etuqeD+eFhIEuaXMzxtUbuKn
uK9z+y/uzHA3dnrTZmJZXWdUK8c6ffEI3u6IU4C8xHrrlOS6k5AYBvbeBQUVKSGzx175JkKXW7yh
r3bObGH0ahunH26U9f9y5SPKE42plA5gQpgNh9MSWyveOwsDLJuz74pu9ITkODEddjpl2lDiapt8
1aMAOcPFhS9Vn5Bb5HB7hFNoFnNUCdt0liQDHdBi2LJ4Zsq1Ihn5UkhhFZ/xuFBM9tAhxJMl2ox7
OK2ugx1N9UtT8VpfmYf1pmUzgFEZv5d5WXEovUbbd3+kiXnUxpOiUpQWQJ98J/e4Ql6xP9YrMm1U
vpaEmAUS0WFWN2Nu5lqcI33eGJ7NeOPPnRcEVi994oYWw3D9MEK8I202CEr+iRWfv6wC7BVLyOzz
nLkKmpBdFrz7i0Y1OQnIRoE2buvmmTX6QaMLut3lHx2s7uJChFZdy69CCraAMcUq/uWkcAH5iB0u
sjbU+/bJjitG8cK3d63Ym4UhICSc5ZFIua0CadAoHyl4aRwFMHzySSJz/rgQeEhdsRRdW4aPct4j
HuMkIEgqFhFNQ6X1PPSwX5DcRPvepSxeo/rDIjdmVRNoZ2EP3sJMQ3QDupY/hy9JsYZvSm9KMuhr
uZR9mHHCwA4LBSFcNedlHIDJ8aM1FWd/Tn8zPYud2jTf0B+08aVRD0He9dSIj5S22el2YBjR+br+
4W8+Hc0T/O0oFDroj261ZE4aoV+wOQdPJLhJiJEJcpO5cBrVeTgqG+a6l4Jxx1YHtZT3oOTLKSZX
PhJb+h9n7llxlRzxJwkCKpVEcUGN9bWR1E4ssgTeC4V9DczDE5fx/Qp/1V9t5vwq5kMlre0vOE/j
Komr0FB3kH03tVe0U/EWh3JSqL2MYKZrcCXkrGMXhB9YuhLqncH5L6JX9yPEN1bXsvsbBDi/dN+O
7RS4sU78ad1bF3wTKdoPhnnnl00D2KlfjkkJbT3/l4midHbGfdGhpwzie2srcBIThbU/OK3gZ34D
3fNV7cWu3q9lqhU8pRGBY5TuzTsPwgCw/CqarLsryQOMkUd3UKYCgcp4EEvaHPomWXME7YDgbd6g
pw9wmC7Bma79WhbuTTV3EVByIV6YDf8UA9n2FXuPCPcrs7VmfPKSWWtDIzC+J/SxihmaVZ3z44dG
4+oPzO7YkEyI3vYmvFwio3vZtobmtk9PopgQjF/z63zGVGDVbqQog1fd0/yFNhAie+vjswBdkuGH
PJr1yiLdkCvwJpor0bQ5BmUxE2sHRKiSIJ5Bi3yJPOpN7GBU0ePZdEkVYv+9ujZSjXN6ykDLfI8b
b3ogLx2LXEG6CHUetk/y+JuaLLdJiUe7umROgI5mMdhQZ6jQAFaKMkvCs0TSSPCohvm3t8gcx7WQ
icQ+0bnFgwqYj3/rP779/jivBHVLaueb3PrwGQ1t8ybX5DVUdXE9I1ooikrurK0BkzKiVWr2viT7
7bokQDmEpyPGeuKn06Dzk57lxUhFs+QgeyW0KusKYQgTyXkJJzPJwCGcwHDna2F05SJAugZ+Ai8f
bkwod6iU7h52UQoje7u8Jnt38MPBoGt0LbsS1d6l2kBO3jNdljGfYnZhNvVPo5Bq5QUmjGaGkeZ7
+02zzn/XmNSpIq3RJ+YWpH/G6vKxWObalUeUEzyA3bidMsf4gL50j+6rK4aOnSGnojOl8btYLs4K
mt9xNdCV7oGh4eXY8JcYK1/gMUlxvAS7axdR7i2CYCd1rIKywioLZDUKtibMPPGSgFmeQw7Pyghl
mtVw4k3NVwhQjKtlrRN0cr9uA6eI0o9CGw0TIinTM89JYlaoj1bkrfV9VGHbvumz7cvH4GXzQzMy
xcw7DFloegDXdh7gJVpfgfFbx3Wt+LLAyXd8apwuUXbTUyPl82nrdMcVl3ocsEaFFUbV00XtoTAV
PGhcF0pd5c+aFkUs1rIAq0dWhRq3ntyG8uDC6u0TOrTHjZPHYO43+psl9j80fPOXlfI0qW4EGNvt
tb5dGUrAbcka1CVgsi93NA2TBKWbA9PHMK4QSy97bfAS8qkEvtc8Rs5xB4N4XIojVB+aSwauzmzJ
kmdHAK+FCxf/qF4r54jRE/T5onArX5706IvvIpyEDM4I5ucyU1ZGmZaVOpEngIBslt/gIh+7Ft7/
N2gT9OrY1OzWqox6dxCQHVfSq8LyveSnfn2LW4Ah1qPL0OcRkKgJ3oLRP0nIP+m6nGbQ/lu2WTol
cYZi4N5qzWXjuKW7QJpVqYOt1gm7BrulMpasUqRyhQ//DyLcXgfRgY62aNIRetcuRtxhd8tVzdEv
6dr/Q/YhMcYpbSL5iumDxxwYrPntH9/DpATRkq5XsbjyAkjFPtmS7bG1TZ1c2OUxol+SxqHGSrNf
Xi0ZkFJrLKL2Ytj3PMJsEhwkjWVqX83xeyymc78EBUHkd/I0LKslbvjQ3IS6kB5itlKOLs0Mi90W
t+U8k06aA4Illya+fvXhVmWIFYtBynio/DrHIY2fslxhsXjrwyjkeSgu3hN06So/QNbp89Ab7j6x
ja3ry7c4zEEvZLrjkoZUww3x8if0Zxl/hA8TOlRbZpJzR9vj37TnYVcnD/BxvHFY6pkAudgub0XI
oRreyB1orDQW8pvctwyxEURP2h2TYr0OQPtzn9xJDdt51gNqyMqJQH6v58at2MBRNEb06Ya+mW09
rTeE+HyQgkhrToCgZtMFbG+RLrmAciiyWVZgSDqrmUW77N6kU1tcrEgsA/atyEuZ17nFwep8DZo2
DCG8aP+8XWw8wZ03TAyQrLZjyWdl8C+mdNT1T+yB7AaHilFZS4zoRLbv0vBFCEk2UmbDASsUAIck
Iq+BznlPSy2x94AGVgzL4I4n1zCuL7PQda0tSMGP37RjmoxvjqvBubQOyfJTSHGpUFpSu4tHr4sf
qnWxaS8446NfFEXhDwI0Xhp5xZrzZl7al0t7N96FvYswnYQKjlOPIX6UjsPxdt/cMxjA8eLx+fPO
SuEcwFm9bK7GeuxVoROdOHN38mPZFl7JP8oT5dy7U2WEP6rpZYYzhwbHW6Clb+IROZ7VNZNbh2of
LjbqXqpaMLgag51vBbag6dO86/f55/kYlyHZtaq6H+Rrg8LHZ5zvEil6JOgOO4zJS96fXTqOBC2g
ZN/ZVsrDSBpGbICnIBSNnCdCKJKf3mMxXaNl/ZnanARVk0APAMCzWBAwdXF0tLz06b3SnxqxxBP7
i1eJ87oEiLjLd+JJ3s1A9s4/W9vBU5nbLgdXWRVdu4KZ5jdGvcJh2v81qSzmDQNOylTaHCiCaV/y
4XXPzcOQLa230bTERDnNQE9Xka9lDcrQsCrKzlTidaSvLbx1Bbgf3y7HoHR0oBQbjQ9sGZ6R4AZF
3xUJ7jvRa8T2eXd3XvGm+yYnwuqZNGQxqWxb5M2EA/u4sxT2mrujXSr2EAk9LrRVbZtJ7Hf01a23
TwnVnspIawUTrf83w0q7IJAoXiGA+dMaKmrfdSj5e9N7BpCfoL1V3UE+9eNUei3h828dJckgdSZx
vtAqfGDtm20djgRkjPk0JvLTOJyPYGQKL4SmRoo7bA+nbe3bsSgWaiUvHMZitcnS+7X7gJDtN7a0
9w28gOX3sarzlI3id4hPdxM5sqd1jVCSdXI6Tbp+t/0CNkY9fJuJuldHlywhZelnf288ptQJZbmI
vdwa5z8A0D5nVztY1fmsRNsT54W1oC2Trl+bVu3n26nmxQIL34r4R7ndRqaH5keFfjSYKIJydRmE
R852CtsW87DuEh87NWISFxouWGW4+dkvHc9futRzgwsVflCrVBS288e8du4Z9c24HhT19q+12Ap+
4JpCXnUGCMU7q7EGQSXRcHwx4rnNmWm3bl0Gd3KKsry25jvF+MiAPxvsyyYmwlsEHYyOk305oA0Z
Xhrv1+gwmAlXheVgzEDRtfge4/RfCPeA6QFlmGr8R3rkhuE4jcOsKfk5bn1OJIzo75jICqPEzlo1
qKR/Sin7BeeRLbVQg/rNWnIPAH+VxREa/OtcH8TBAiqz2SIfrL9k/GzhfDANYRcqWnJyxLoT6Rkl
nPHLVhlKFhT7V+yREYh7SVBLZJZGH7WqPTOhfhWkPZpat3+VDkth9/bZWWyfNLiAVXUVj3jdhUDN
UhVlaEl05htkWHfnf04l8wUJiaczzf7jn2ana+8O+nIY4GVT33S4aU5oWEkkYATQQnTFmwYMzjIb
G7FC2jjGM6jmPlIJwzKl5DekcLyri15ZW2gsCwfy7O+fCQQUazCAk0RcNHiA/tiKUh9y1qdWmd5h
Zy62LcfHxSLtK1rgKQHXvwlBcRh5E+zVbXoeTqIIKEywAtIaKQvfAd2WZv8qiFSJ3TauLX3t/WZc
W7QrXogLg78s1udGuzIFc4K3ey3B5Mv2+GX5MNr1J17LHp3NOzyg4AtNJasrmCk2x8uj/0O01y5a
M/8HjJppDtm2RYKsn8+aHTyx/5i0ETEKgYUNWtwje+3rdmB366soTqprfiyQtd8kLKw7YQ/ndkcY
O+JvG+NHoCecHnOn+IaIyi0Qf6V5MRRYlzv+LUs6XWmjc26aFLrZl7XqFnWXaDHfRbtPXFWFJ3TL
xssoLbigLb7k45cE4xt8oN4RI8CBQUOv+IIlsmQ6rvNbuk4PU1tCdtM3BwDlsljaVknNI1dtll6g
uXBrM0fg0tl46ReTYUtTOBcX5b6hqpvzPFBDOU3AD7QiE/xgH06uzSesgIctsoN8E63GIDmuC1gI
zPI5cddsOiKV1Meq2swsnMWJaJWwODscmViz6v03K3zl59bFO93WWC2IrXIlcYpMccO9sbhz8iN3
BlcNlOZDRwZrEcipH+um33TC8wDDAfZlt9X+9BLnRvIrrf/fELefcQukPG1N4DzIoykjZy4964ZA
RZrTmkfTSzaTR2i0ktuvmjK1kjKir0Tn3RVC+tYu4aeYI1iAm4Ery/SeE7wQbdB0V3RZ0pT5cQu1
inzER4DvlihfW8uTs7fok3ORh3e508xBtvH1/1TODyux/33GouOBYFQOvzg4q2e2SfxgVARGVHyU
4kZ/g3zcb7erwRjSxt4NoF+TiN/ROp5K04NCzOxZemSJzCvnjcx3UqOPESlwiOL2tQ1pQ+dwiQJs
JLiexvWcjOJpiAbJiRV/rvyWbZQuGP5BTSsjUfFYlc3mw+bom7phHDO7FCGOQfHxOoBMcbFOzNWL
qywZrZuYIao0IPUoO5BHxTuVVN8o9z2okpqO1ciV3v5UQ5G4jGICMZSQojAtYNH/vIHlSO1Qjelp
Cu3i0jp+Oa+Lx1Ip6m4kV6SN1MPxfkAnYlIwRbdvO/Ktazbd3SdQLxJ74zfRkYDmKkXfvu9GLPOF
xUNm0bIyj4Q82oKdkYvx3duWok/k0sjrhGZp5VaSIwEwMbguQM1zpIyhldr+MmZ6WH/TNY47YZgO
m30n8ypNcAwSn0Y6HEs6GdSGgYBV6IYuygX9tx4ktyoQKTVKd48oRfUZ+si2Cft6TmSng+uIEXdJ
YwYkYfPRX0HPXDp/tc8Dr9HjqqEiR3QMLP3f4VBOWe4Dp3aak1VWQlbl9xzrv/xnP/PiTrgIvKH4
rTAvw0UAsUbw7W9Tb5OMs3KMST4YCqrzz4cyqzzbTashwcH9RYCp+Acb0RZdhBUZd5Zr6TbE4wRq
vxoj5ZEPtCyrqrd4BHmY9PtemmKlOx0TDQJ88vnwL4Mtw3L8v3SVBONYfkJWIs5GQfDuRj8dzvTT
DtuA+Nxcx4XfVyZuOGZ1F0PMMAlV/PjP9Gd6O3sZ7o6VIOZbiRSgDjQPqFKRHKSoqTqiLjUituEo
SRYXXRxXVfRtlNQGCo+1mSXRFqrsgd8ibbweK39ukpYiJRvRBAYIXszFDIN9StnycBkgX6Y7FWSg
r/udCQpclH/2fgqrpgmOoAc21NLUVG23vPLt50CG9VN2pjTcaCpUW8KPwWMjqWp8yCWZvGqxWljC
REp7D52q/L9SkNPE3lb0Vtahv3iKxpdKTeP9eDoM4UzmlYZZjKo1S/2e2+aQr1knnRsrN3i1K0Pf
sFgZH25HWx6A2sDYHb7T0pkn/lXNAOPZXJPuP0kgUisdbhIIh9e70xFVz26o/JNM+s+scmZqwrGc
j89v9I0hiCKtaQK6T3ZL53CoWT9pyEmUXNolPPHWJ8NSK/ZoxPEsi7DtfHyFF0U0ixTnWhyS3W1X
M1mpzBThPlfVGA2lkEx2MvGAQqogKIyWqTFP1tMmjZCx6bY7t6Ci2D66+ugSvA0mAubUe+y7AjcI
1EGq2NzJYgsO7osfK1o/1drg3PA+cjaAPdSBcZ7gSRXBH1SDrQM495HhBIGtnETmQFuDlENMhAyG
Wf3yD8cZUTOCUgppSctmkt4zY/vGS5SfeeoI0FOBE+e8AczfwdbuPzytV+ojsUHNtcbBHaZSFMSQ
jsTBdV4dwxwFZVn6aIW1nFU2eJnIMu+7EHU83j3BGfR17Lds+TKg5jcMFwg3gVBXx+vSS56lWsso
Oy0QbOfeRGaORznJabyueIvjmRYdT9UxxahFlBbtGB7FGLIc9a/ffabhblLNc9ZS8eIkQKxwJYK6
uRHJmqnJFVavES1yxhcowXlI93NxinNR6ktFiGH1c4NEcXxUzu4nX9JRwLh0Dem60zVPtd7e/5hU
4lRxXGqvDFC203T6cavfnh8aMAJW/vU9oiHYSmO7EqIN7W4ezC2MZGOjuBP1VnWQ52eXbhN59djI
9+46u9TspR6yWBBwREoXhf++zsqx0ioRovbf82R/alKDhGqHPzBxMmj+d3Om2cJGtnqjj9wrC5jj
eo8rJ6toNHPMB+hu1WRanMrOJ5TbyhEm8ZREXZFzFzpkr0h3uVgF7RhCLCRe61X28IRmNq5B+u0x
QJmF9p0SaZvgXiepIzxRTKDOYamw0q6mwcleKA3hLRYy4csgevT436xnLrAn12UI0Q86yb08rGOm
3g+nLAhA7t9ju6l2P2fjtTWzQwZVgBggwCi8AA+3LWosqU9MsB3CE/dN7WrZaYMPj9TX3ogA/kwC
FpS8GTpiGzMvoaOka/uHqocrfB5DKlL+FFGLYtptxw9pSA59drEGOKVfUoX/fM9PXH/7I3pp+1bT
CCT6fx33gSQ3ARKT3jDra9VV5Uq6KWUsXyMY/IuoLXJHA2tC5QOM1apyVqF/R5fUAHhHHWtZLlW1
3iHpj1mI6P37qEbHuuvVo4G95EtIOjP+no8nzamEr9ijeCc1IjDgcOgEj+gpD6Bp88moMwbeAO8T
adEMx6xQxXgulicIxJEkbFMtp0lHjy9wgVD7yiVAu/LimAc0e4Jmq1THdJX59uFkNpUl+q/LdmZr
tc+uFvhtVfJG5Kv2R2LvE+3PeByc2bZa0HYhlfXovvJejmW77DtSyiNlY8L9JruIDaJ2TIkN+16B
Jsh9DQXzu2Y7mRDQ+fgzqHWYjc5sRkAQ7VoaP/pLBlP5Uq2EFyj0nMzg2IPw76H/KZAkqtXU9Gcv
arPbQNhTiZMqw2bB81JS4NiLqFEcGqXh7G9XVBiLJ/hgipXFrPa/9f89TJaHFfMUJ9atBwyMnHDd
WZQ43hrQbatbUv//pg7+Er7/U/jOidB06GFFwTsbnF+J5erWla+JtdhaxuK82g7cgY9CMVNQlaxT
nSZoEVO7Y3bylvd0B/37Is6lKGCXluS6uY8OzMYpoyZY8EZ/21DlB1IwyFxgM3OqZRUR01rpR6oE
gj+J1B7nxEPB9wCvCNwzxqqB7uaHDE5WkTGQWcmXcg1JF8VApgRBJY0jyfatIy1wBDH9ppkvnNqi
t6bEd/E/tBiJP45IS0gnxQHuSjBhp2B6vlAbdbMIydju0atpqIU9lqNfDykUlV8Ck6Ucnj3+42Lv
vMuHrKsoJpQaa6mTfjFGXOjrxNACeed0W5FOiS4rBrCzHbq7myZRL14XqIqRE20lSSROPnpEPwyV
99dHksB9oosIK6uGyX3dRQFFujBfiuzKZG+ibHN0zspgNi/YqnHfPxarTpZeApGbughO+yIYN5DV
IbdOSsDpD6gsW6gy+yE7tYxlZK52lvJBhNSHGtS/4TGBuLntal8Z2AtESr8C0TePnWCphTknUmAo
FHnoyHPC081HfiByDwFOceBG2exu1AjWT/6Mj0c1A/PfdP/ETymhWz653udvx4Tf57MH70PyOE99
YoK89uTWzUdBGots9A4jtyqlIPCH5zUgVAlRb6hBz9bb9jSAFwLw2SatPaOpxBQnF0JwufdKs6gb
Epi/ZKCawxfbw9lgId20BOD47z4F9D6UQ4qaFWOK1BXbfVqPu/7oG2G4MJsS8ACksItF8oGef2vT
TNccjFdyiH3goEOvoA7axLSNmUL2m2hlxctgeCmzhqsdpyc/aR7b4S8QOe1oL0irx9W8MCuk54oJ
VR2OsVkb6mfIvLdHgQ7BPEfkHpRZKIWRBsLZPkMrjUpJOLdapfKe8iIutsFHb+vNJMuvUpLwzA6F
z9X31dgVWXstgryx/JtZdZZHmTgr3dVixo9PBOH2Wy9uYrOhITDA3h8vVunTZoWYs410jxqjrnK/
PFgTlDyOkHnmvkbApE8wgQRVaWBBXuIUrRxs5LCgtUeqXrFysWzOPxoOeDJlGEZyALq8pKZijiHK
jkdVNMhxUxD6YJfVUx3F9+DWYYt7hVgm+OS2+hNRfxWmFkGa+2yvrEIE6tV93BJEwEdAPDkRL9mI
VMPUs5TKsUFh6OauOC059sDiyeezuDZw5VZtU52AwIWb9CvhFuX2zToR3o0SWzpaff9ucc8jOhvd
eNPYFCufJrYBLuBvTusSP8d5iw2S+BpQJYqHshWxSv2AWoSIRk4VtXfZOQlw5peS5SnvOBD/SHeH
1ZXv6Q3NgDY4Bf8PLzMaD8hgfI7nRlXHaIDOhRmry1lq6OdHQg2e9q2bv6m4AgoGM4XmH2iI6Vq2
H0ffzbTKgKZQBr5VYBqXP1Xg2fOIDs2B6RCY2PtCvYB3ePokV8SL3VqDJFFiZ8+sz8ko9LiqjPMF
2GY63g/GbGh4LKNko30+Pyumd31k21pB+hID7meBQqAwKxJp3AGXtFsDldR6B30PBlP6dh4NMhEd
1wzfePcthrIUqW8xHB4xHeUn5f6WFQNH6UzJIplo5TmXljKvSd8z+SXBpQ6O4/Qf9wVX5EZjBWTN
V6pdSuCeJs8eKrHMeGAutQfnKmiw1j5foRwdT9THfCbeAvQhUSyKcsvxVjyVJuT+VnUMFEMu2S1k
SgxS9BF7hPZGqbwuTTs0fSgtMKwfM262rPRyJORtHD+SSlab2dNvwJdVvEf1mYWBdWixtL26nG8m
ODypiING9d+sn8TgB3Wvev1iqx4nS9axjtZcqJgpiM8wpAr4+TyKCme2KbjrVI21qRMV+uJbfpIl
Fu3g017rmDGPtYWi2OiYj9xM9f/53oQDB+5q6LtLhVgVKdUyCpTX762p9M1cW4+pxItnRLT8u9Qi
wLZ0B/aGOFnVBTbJNvIkJc+gKa3r2huvOi9M/stBZE4ibLVwXiaijQswYoO+k5u5i0eZWC1ExLcj
fyxkbxWhEGqBP0Sp9ytN1da2bUdKnmuNReGdXwN6gHierDc665+T3OOuPaUm+gcpUgcoHuaF7aT9
eTaQLUN5tzWQJmQhxkUWsAU9SFo57Ju/+BhfW2spjDhdyuDORsEe7imQykJegcBJ5XPsefONBCuT
mOuyD5DuCjg8+UHZpPyBI9ruovRIruTyDWTU7eifJm0/dk3jT0v2RdyXlsH72nY+TB3az9Fd1Vxg
6l51l7hONabxezp0jpfl5GVYi1rmQJEGJcupk4BXBcS5VvaVBq8BJVEhzSRSiL4fvIhkgbgK8JEo
HPKr6L8f+Gk8KUNUqxtw/A2LqAMVgGoz+ElLZz22Bu59NiSLeGTWGb6wD2l4Vrj0sOWXMiGoK8c9
NAyIIRH+i6Z2GWr9pUAloxBCyQgDDKzgP7ejAop8YqSw5KOFYkFX01tWpvQwY6IET9ji8K4lhnrs
Pawpl+M+PKjkEkl/l4ZUkWSZCX1JRbn+RvY4jz376UZDaokgtYrJVNUyHOgvLUn4qhW29f9Zo1K1
ZbpZSCk6jbH8N+0lrfToJk78apBZ7gtkZyNC9TVWCI8dxWfsKU4c5TOrQdlWFRduL7cscfMx/tkQ
QdaDD1lEkHfoe2+Qq/BP1IVt1g9wvUyrYwq+4Wl9wzBxSIgEnMDfmIFwpbiwF2aI1uMEaAtmfyun
9EVHte1AiazuT27V1ycPGkybCFiItktq1AYP/x0Hzw5y/asuf8kgXGQD/4sHZU185xY4YRb2d+a+
WXfsrT521lgADahSjw+jEjfrE5XNHu65RiEWpEr3VWl3oXNRDJT4iVv9+igLzSW/0eQcZtdF1rEX
b9i3Az4ZueCD9ZyzGle60G4Lo8Jy31lMcQabSBzPYUCMVW/Xvt9si9y0hihGs2JjaRnRuWKHeqxA
GxXgP2HJFQ028DXO3T3cp+QchAcD5+KGEShB+Z6iRdwt6+Y7Rr2kYqs9j3GOugnmHvRrwWfK8Gxg
kODm2UwngzeaKCRsEmDWecXKPlHgKfhKSXCjSKQXcpfGJ+tUkDANzSu/y1IzCTVsNX69l62ajp0r
xajSsUfTkFtur/TMx6UJfB2nHhtxEr8YNOjMorICREDjLDOliNu0MdBgj52IbqMD5gQyujHlW4R4
Yc+UkcU4yk1vfe1vwc4chC3PMh0Sv8eEu9h4iBiO1ZpXz3yMEj50212Lw1QufKPCJFxv7zxgMAZf
WbuFjBgXGSpG0Nys4+pzHoVLcCimlUcskcR0GbRh+HHJLZhIrv+qdp2f8088zABkY+uPkGGaT0JY
q06phoLZ2xIv5Kc3xE9Y5ZLsmiBNntBR9Hl2MdzqKTs/Zx9G2ZqCDxIfeVj/BaQ3+PMNgFqREBVe
rQNF6kQbCpTXRk5pnxK9RecT7oXu0Lgbr4eBcds7a9nQpg0gVEL29muc063Harr8Wr++fF6gYXJ1
DaQRY227XrKG3bpswxkd8uJqabPkhrl3WdAH/fVykxA+D79RZTeJ1rgTumeUuOsplfau2/4pNVSZ
e/iiFaH8nP+vAfzErYK6h5g+muuY3oTkBIGiqUN3tRjGLd8b56eHMemF4putcbYEdUXWsbTtslYV
GzHnLWENllXQeuoHqcFrZLm6PUmK3BYUysYCkzNd0CFr70OLQkk7//0Pmvg6ljbnsArE2zaMdSLc
ueYlE3zLt2aS77tl2Y9SwkuRNXD1x88xabnOVQAkoSdMdoHk/sVNec0mxSrnsmnMgYVgakCzFzaH
OGlO/J839DdwxJVK3ccpvl2pyl393Y4T/ju2hnVMi2QMf4S09r1CbKq1ycdhti+e1CYL1YPfR6oe
9iVXpVc/A96iYcPilTZUQku5qMj5hYbaWT/Z26NgWS0UVyxKjcghxSpZyOnWpkk0JabbUveyq+/o
QCTP8MfNF4w7YgpKrNgGO+YH2WymEqs2d7rfZYhI0dG+TQgacyJ4mMVat/u3oTOpdJmVtEcaW6Le
lYQtOstXU6o9CkOiZWSdkQmIC0CSF7ahOpkLZ+mPfRRgJejpDJODM6JvJKHwTOxYFiXbww5JHbq+
BbNgniR27qnd7BC72Dy6xasOUtawc2EbMEA7KE1O/Oig10mUc3WQuyJl4jR7pg+XJf3FOrDsFR1w
JEEZjx9RN9TXyYjRbIPd/l+lp9/Gh2mcoGHpSqLbD3v05xRyJ1d+Hin+Co2DQb1Pbso2uMkpNrWd
tLNZiQS26FL2et/WyWRXL23boHeBI5mPgZoBfLhxDCNcqVA9z3W4Gx9rc103YRHNnSd5WZan8uN+
EHiurkcG+QYqb02EM+lwEWwkFT3gIgM/8SHL0j/9FAgm/QqHo6A9GEZwMx6o96whOcSDCOHt/pRg
zLUdq1fJgnAFaoDAE4M8Q+c61vqAC+2ifC0Ih/6d8eMjvfnwyn0ACAC7V8FvFLbS3YOKyo7tIYPa
tPyl7BnV5SZo2tvMOiGfk+XdJhmZXDDakJfr15pBiixT4da/evAA6HCBnmHBuxeFrNoa0kp/9fze
yUOU3JhVYW5nHFF1jQt8Immja/VrpwxW/NeJfybxC4ll7ph4+v2wsWs1McENIhHVYkXxtzdJnLQD
E3br2tzz/UA/ESLfgwOo+COukT5nyEIEsv37Ng7hloDJSRvb9tr4Y/YDrLqp2CKi+AENRO3x1ktl
zyGYLCTZitopOUnglkOcOdqLH9WWZ8iNOTWZ4jxA6TGt6mIVgB1NkqhhsCXEfZHqFTxrGo5zV0ea
uBHHxDDXcOzKTTYtsaQSO/VC5dKv7DslXtTwv0l/ZkvxKzBI09Ce7EUWXEk5hGluKMAb5EnCPFvF
r65xRvynlQBi9DhoJbCuzWFtWC2Pxg8ywGYq2H7wNpqHxZvjU+4kAIWeCcJQlUTW70Bo/aTaGDYz
dlwXtRcF14elE9nv9Im1EUqgSrHcfSxKrSIjWmGtNLV7xAtuFb95zKlhuUq6ao9FmsV1XrY44pgR
KBkyhuN/ttS6XbIGsJ7VbzQ49AQKZVfTSnVvlHQXk+VcEFaoTBHTovhWRSi9iX2B2vDCh2pUNwrP
FFlU11gQT8Ebx8cg/t6SGEjvX4dXCYcbQBACkK5ke1CAntbrCjlwzfseSTy0X8f4KYnbkxWMOZ3J
vborn1MIePHhhxItlUd9WDtaLUgs5zvrGDrN1zUuXhrbjYYODdaV3HBoUfSyEfbwVmsA1OJi9ciy
eUoShxyNASLFfF7PCOzemxxzZ8RqPwJ4Y5BHTLJG98uhkBDzh+ERKCf0fnweeiz0hLCFmaAV5BXA
ZYPI+bZu1zpseIUCdAWzy55g4qzy0yTF6z8Q7XO2ZvcYzvgYiGJRuWB+AqcGxr6mMBbErODHj3oL
zlXG6TdJAXY0rWAdInYwgUO3w/EvLbojOXTo2ch48i3pPDcmC+Rqf3EZ+GVsGm46jlaQoAypSmVy
q029worx0CTNMRCVi6DXKEclwWLrQ6UI+zJw7xYuENVJ+xykkb/ZqeCyu3Y76wH9LjIgAQFYKkOa
YA3phxkkl1A1ZDeCoV5ObpQXkDZoOF3R/q0GuErMuF6qEX3JbcHpvgek1UoLSbErPFuytp1kWKKb
dR07VowbT3GYC5XdWIVMd55MK8FWA48HOZoWV+9L5+jSeLJAVPVuCg/gjVLXIohNGu6iiuTxrx8Z
CdrI9bl1Y6GNJgJsOYZrF2Sad/2mgCfcZYRn2ufKMdKHTXDd9dbh5yrQ2EfRpzs/89pbFrit5e98
k7nk+RCMtgfsbfD5ODJMSR3tvFa3ty/vcJRHvo62RRrPlalauUwdH0NGG2F6oMKTOOSYtzMWchfi
wrVVMVq3qnOi5D7awVJylZHMzPaoXrP48o9pjKMoQ313y4G5mp6zXQaqD1EcEf7gw/r5DM5NpODw
uyyxhhnnSJ51Y8qkACyPnTOSDWxWEkmLtUL/JXcdw/0Ic3SKLzQcnlBQ12vtypmqxAehsnKq2HZk
6sxDVKO4fbURp71wTef8LpM1GvGTl6hzmgbiQF7LK1t0vJff26Yr5lgK+Z92944J+TJFWWzesddc
I982Z97lrBVgb641S+8B16dYEQEyk0qtg3lyH2twoqGcj9ZZLFEJ1KtOWHD+ARuRO0BvZlx/cceS
cBvyBUk41poEjClVeQIlxvgNIOy0iFvv75W1SlcYOQsnq/wPyxDUHv4X+PsfyMpFjAQCiWHz9OEY
PXXg+Q5+spnlefHFAfLhRaES/dfU+JOGri6rItv2fAWbe03xBcgyHssLZVk9QsCPmmBulGunIqEV
8lPf4ysg5Jq18j2b8Y2M6uEo+yTwq8E/7uOxzHlT337aovlXJN20a0vVdVgNXM04ZY27/z9ivpbW
ffToz2avapNTBZCS9pmXhM+ex7g8T+XjRBLJtZho/SjpHZRPeuIai47sxI19o+RNxf2RIw3spPla
v/0bAMgWNY0rOVZcaTknhNcseSTqTcnBv6AfMk9juuAnTtL6ulE92/jLwNnr07+XigrTxcMtyunm
N4aX8QzQMl0aDfcfvc/4r14CW2j0AMwvqj5MqiIuJeMG3Kxdji5QedcWXw0kuhpL+sRFx1tHO2Jg
LV6q0tTEXSCogPrF/G6b3dZlFZl51sXEHqOB5Ds7JqdN0Vj1UDpwDD1smalh4A+e18HDuoXa0TtO
UNvtVZUuT/wkz6dU0fw7CV0b0/wbT5/5pYEghwLNNPQSPOtsvooPcZQnRQSmOkYAnHxBhiXTckzy
iykOrjYte6zfcsPAVSK3C9PHkXeL0zI5xkqbtjAVB+k7E1n8TjHgL8ztcloRXkWXPe4q0FY/IAz/
ZTQBJBf1bAqkzCItdDu93GlrBqvSuuff9cpJFnmXMgxSduLlMnKnhtMN56S07DilCOjJ6r4WGPFR
ke4tet9kF/uK/Xwn3LhuCKdTREO8STtidp1zz5QIhSGcN8mVwUONVLpLDny95evzMpqav8RI1paA
eH5j8LVSWn136GiFW+SHorgvIM0ESM+cYWofFqhkxXqCIb6Qn7/1mjo5Hmn/QPI8eIKc2366T+iW
F/i+xkHUxC6Bjox423SCRPoGUhjORXrd8S56/TNP5iCVmKsoV2mL9NGvXx57YvXSNy9Ln1Bz56T+
BV68fSaFMYE0imSp7ReamST/KOq7Ru37E+ZQfXFWafZ4n6IJFZGtgaBs0zYBO+scX21SLnsDpy38
K+jB+5FMnYLRWgEwGoSm/wbgrkxPnFKsyIvrmhPb0NHnIvOLlwsNOCv0VhG0vNkyYik43+jp7hAf
/+2f0TafwkHIm0aAHsNXEzmC5r5WzbU4Q7by9/m11bf1eG6MK0SqV5Xey3tsS9Zb5GjN9L62m8DE
gcvdzLlrbcLr2AEklJ0dHpyiFMzl5ivmMt9q4S5LpMaagT8oKZ9BrIVtsAMoFZN+qtdu9iXaR9Cm
GWb8GaWpZR0giZMsL/ZbXbnK8ysWrOZJYCoQc0zt/kfQ8a6nH/HETka8AQwgV+BrAVK9/ikm3Fje
uGb1yJprLFgED9kDrDmR/incoE5Sqr0BbVredDwS5xEqrrhWhghAMmdRxFmDb5P+qjJlsTC0SQpu
6HKYsSf8jllnrcr/EFzg78ivx5W5B7x+rMObhbUPeAvj7ax44iCxP4ZJJEJI0Do1otYxAMpfjrsQ
7WikHJJQO6A48r3DTtaPi+EXXRR5p6aL7JYuO8VCOgCpvRAW+wiW+ULPuNjYUgZ+6bftqVBpKyj+
CaEBF7NyguehNdyacVj6wX3kNArL1DBYagDbWOJAGFY8BoCzKODp+6Fhk98Q1XBg7KhIhoX9li/C
UsBJOihSWbdB2wwPiYcCHfqU0Hrm+UUG6s0nxtKKA5DSGWcgG7v+aSubmhqoxk5x/AFpOhI3a1fj
ggnmlY6rTfINv3A2UWQRmQkjKEgpbjq4/AMZGPAqv9pXaZW8Xu1DOkMLKfBhkyQUGPsgR/8vVtAw
gKQEPyGZzgQsFHg8KMTK9pgPYfzfyWU3Pc8AX7ISKuFu2nORmn7Zz/fcFw2rmQ6mk58ISJKN1FMF
e2JjXDRwEFVMi8er4QsqT9cjDFLntCC/g0iGCkVXhJ+G6oKtv3nv6k0z9HaP9Pzw0y2yca1X9ibu
BKAwOg8JLom4UXXTqfdaPSCFoU3Uo3OzY7mWDRHi4G+CBd19kuD+/2v2jym5DtZFrocvN9Nb/L/U
WinNqIo4oHfkNYdCRT+by/E8h8T1BKtkzzIj3MZLjr2/Q97ptcqrEhSUy80pQS2712aMGvtO9RyW
MADh1MTDZbBkJ5p89WQnldU3AyuOwv1KycNcw7pZBqjt7M6E0Ft6Fjigh3yf5n6WGXNLze738hI1
pwcmBIEujffi+yhjc9BlhS7Bf9VWJG+E2paBhuwKCKZGadXDK6d/gx8XYkhXLFrOSOcSltkYwtti
eb8utQT/BttfA90D8T8Gj8axgEO/09VVBlDZAs7DBj0a6tMBhV6tskTJ060xRYl6Z96IJJ3JrkWM
xxCoSmIKNGcg5c67AqoL5quieU8IxaOR3mmb4RSGGWWl0Kwi128yx+JXxvzRt3vK6PR1aWu4cGEK
lUWML6WIlHwTiySg0ResA4pa70vHblFQ0VUQHU1nFN2O7aJhz5fxjBRBlMHyJwB402tk6GZRNxxM
cukfPbWH7STyQG0d7nfjAmkPxnRuIbIcRTMk9yyd73R3vl2hoOIcilbYu0wVdZmsKT8bp2J6HXss
mELya297U0cdnZMsRK/lZgDKvrE1bLWjFD0RdV7B0uhR0XoQrIYfoL9YZTUMgUjKRiAJy255V4ig
dgnxOM8FMukjP21vyx8CqVTmcYvWz1igK72xlseco1qX9G6ziuxkQ5NZYHxSmSQWdmkLHJARPXp2
YrV7qdyuO9HRgCJZ3ouNGWfDAExMXy4Z77WlvV/gK10CtykzjLFeJw0YC5+KCLcX+NMQyjd0KBvU
1id7EtpWRsHl+w5GyuP5w8dbEmn9kGAzggVqda7bxjRvqrcOF+vylliof+URfRRwRilWI7GE+iES
v2SlMX6AhrQPugMKfV7zSB3hWM57NED48Yh7wXVyoWiKlsvo0AkBcPP2ZeKnbnh+QD+9V0f22Vo8
6l//8rKpo/hUJEz458Vj4qzB1Gz0h8l7WGQISuG7R8RzhL24EVk1Fop2KpjXLDv0HhKXFpKskbP4
2nvXVR4dTGVwPLhr9Zo1God+qZ61iKq2JZK3jcItCHPEweZ/gU6HW28DqjqQlsbkwUh+HX0EXDSF
E9jmqREOAqwBFvc+GJsJ3gu/2UDG+/EHn7FiPgcsEXYgBBmJbZxTvLZZX9WC3/QNVGUmB/CETuaM
n9KsgRVvGZgtki2uNWu+ZSQ9XUJGdJ6k7cOTZgEmHrw+bhNFvY5HjQQBKkl7yt/qi9/Uj9Nkrddl
04GUpULR+5F2frqSejMn3srmcMuBp2f7o59PsKc9tixAoNcQ11HsTN/b0El8wfF+UYBpC/mDJkeP
Thfjxwrl1341Qo4YEBwMcLc/iS4K/qK6/Y53m54svyDUmS21tn7FXiMMXvqtqCjQ1UWlKpEsQiJh
Fp++6ab5eemhYcPcT82pHC/bVGFyT/WWBynemYJ8twFm0CwaCbtsJtVQxLfTwNN1JkYOLf/t+NPO
AbGNEuoxZXy3Au3HQK8IwKQJUS4divn+WhTiOLtclV3655Bb/zZveO2JBIz6bMWiIv1VgsrB6g9/
zdEuBIqZbu2NUrFn1POnyu4lRmVxy87f8K5iOVtZoUDf/rdDmwcRDgO40NUNX6l5MSCXw5lYwhOj
qDCDKAKVEMaKZJkuQNE6ccsRFOU08wf7RCkPie0NSR+0YJGLeJb5CJaP3c7r6L4pJ2yLBc0qV+tT
njJViQ6w2tiW4JSvBIdYkfKYEbOnBW20AastJNB0e/G+b+CPNqd2CsYl41SMO/A20qF+3qhejAIf
aKFv5Q6hCXsVoc2RGB2TQg5BcJxAM0J4Fe+AfArlRzqB50lQbqjyckYt+BTPW2uroLsJ4c0Uq+So
1GCzV6yXLo1o1MLVSlkcY6mRvv4sYecU80qlNLO/wAsByvD2dZzt4h59dVXefH6h3mAPofoB078I
v/Y6O1ekN8n83uV+KfS4aWy7TRWh/tlXYKw5C+yU+SPNP4mP7AIqfFAv+Zph2J31CP0SK8h8U5XD
HpEVU417uuenRbAABhvLDQm+bVCiPtU8bB6kPFynR5g+XcR/gq85EW8rfDtGuQYDCGdGzoBR/BWp
g4fjKEB8/h+lF3l4Y3WkEX1Unf2k3T5DOjX8r9DAs/gBsCWuRydATdEo56zOTG10mReK5OREMaGQ
n+uJT6oqpIuYxwRgRULOP+JHy+ylsMtTRYekVV0zteILX10l62iD4tZMoXbkFd0/I1nKQm92CYsv
B9EEsziWp9Rda9/v2MAjVssAhoV1+jA/Cu1yw70oPcmGrDpFsEJ40HBbYt8/9hGMlP0bMzQhcNF0
9uVABf7rQMfZmoqHT6THXCbg+aToLHapNDyyexFXc3I0kw971DkqHERtd/bu0T2cEZcf1qhqYs1w
5cfdBj02llZ9J4DHqxTkdehIFhMslcFg4fvQv/axWjEdsnbtXiA0Pk7dUu8x179stPkRc8sA1IoM
jIMp/bwrZY6iQfj1IQ1PtmDu9HjSArw+ZwGuhXysd65Ii0OoP/EXqAY3gex1Ej5HvKiTQFg+UzsV
TiHGqnivlAyBc4Dp5sfw3LfT0eC03mQJGbJnR6Q55gIIlzbP+sKXdw50JBZ8jx+dKNATDSI+OV/F
WRf55OGMxwAffoyKp/RfjjLTP3gby+U/btocpYn6WdqEvJ1h9R/6c56s1D5iNdSsA47i1OGGNTtl
/8DiZtu8Bdcv3yrjAujF/62YnDpMgaeXa4RLHO70JEiFLVgK+yTbWc2FWQAzA+osxYyvfvAAQxNI
1bUVAo3bKQM/VzHOaQGu01Awi8nEvqM4aQwGGbw2HYUDXBai2YxtFbHQSyXqYaF40AeadrQ32VIa
tku9QSjeXSPY/n76S+tEbUaOhdV2iantAGLc/l0BGoYkoPEskEv61VtJynkn1tQBoW1dVdJ1e6rR
X1jSGsnUcjFhIwEX2NSbv+wXzZVBt1958rzE55YjZUmoHm0fYqDrkVOvok0jHpypcIfDVE1TA894
c2SjTt4LS+CN8mCF1ML+9NI9hnNqkL6L7NRe1X/9a+DRsdWgDgw6WUMpKS/NEQT6dLCvk7GDa6Mv
5ULuPLNPqH16Q+gXfGDGQ8xyREzMy2IfbupHi+AEiGExWqwzfZxwfolzKho3F21fNC1vr1h8xkme
8XgO5vdve8zx4BBD2yhIX+rWr2Wkx/0XM6rgJfKJQ0T6A7pNa6NnZnEpSgZT7Pb0S1tSgPwuisTR
M48WSyl9RNPHkhGSW4nXUJ0Xe7k/dpd+t3Ggmv8+jiun8jsf4J5TSu770tp5/XLrZGVjISQPw3uv
BNzprkZ0EePZrduyTM6v0xm5CFc40GOpaLocUhakslt5u5WLJaT1UJ79xF85cneWgBIy09frv0+7
n0fCTZGdvXPpzW1dW954zmBASnMXdUzGu4zL1YEcDSNrmfvOu6PsHW887xkQ8L3KD3Okv4VzHy6/
0wKaGvWVkSrsftD2PhJsCeEtVXosvTmGPpoP9VVA5utrf0ftPktbWLXIWvbt2LXpUNPFo30Wuq0W
Dnm4yTa7iWrCuDyTqKdnKoOkonrFaMqr5I0Sa9E50Gn1UxLi/FM1C+V+0k4KYNXVJo/TnFGs/X0U
eCMO8kxDBOshh9u2B6OVE0/Im5NFSq7Mjsvn7HHZH1nPPEUYzo11kRAroVsYkSwzgJwVZNYgvofD
S4+CWVSAW9QgDdK98qcU3JfjBFnsc/bkx3PUM6GbvbninPWRo8v3YMiYMkT0GZDEPfnfSTLpjLAc
/GTU/nytPMke/epgNNN46I2ZE6K3INtFbg3px3+A/fOjW5LEjG8iimJYTlL60r5tlxNBIRZu465J
XWlCuXSAZhqRhLyPEhzNrYvutAUq73VpdzcV+v54Sav5WelRvxXt/EC7uMAqpKQv/wR2RpoAX4ki
g9KskDYyM0Hf4ruhpQcxCQHFnxDsP7qNzftdyArxT5CzIsuHxQp3j6GkZVdtg9avxTeVnvkrnaCH
LKww5KvKq37IVoQ5xWJTb7MItBW/JBcMMDRaUQVrWiIObt/Nojrl0dPS+WRVMDLajnOfauHmqhJ9
TCZJZ0Ja6P1Mgmk/Xgb6YTWTyT5XSjQX15lSTXtAklH5Tu/QvNUItUpfsF1RGOY86lSCRHGQaHhq
28VjCSs6yCQSgjFgsQ3VcwoW4LmrXOl/q3W6woxscLfhBvu5odtMdCW3W5aVVhF/S83q6PZwTzoP
OShqn2W+lte0BMMdFBZvq8rSxe6h6GYeUakK31P9mpvWf1aIC4nO/Hk9Q2nXJ49XJWmtULjfcpMt
Xar2sZP8wi5wsgsuIeYz0poJxs6tTruhNodNlh9I8euryyROsNQboXSP3YTzza4pHedLxAqGBQwf
V5LDiaM3RLzBWjXth1jG0nho3ieGJmDTVzRDAV5R6A49SNt4oqW2w2XFLFaLqCqz+esSRxR3pUeD
W4OnjSBSWIjO6AKNWvXqdoonM1lUPuUXqAjCH4kVqqsntaI0KEHO7gjOqr6a3K3JswG61dZdYN1V
l59gU5LA8uqDGSPteydP0lJSUf53lVefx80Al0vE1OsQZkAiAKUb1opOHf8rMqZRbgjujln7qQFb
Vo84WULP3kI/AZ8lnGgGTRxJmjJj8KUt44C6ARLwkasSwTKf6n9II3bbPiVHJV2UBF5R+ZwouXYA
79eDKlZKpaFM0R6H6zKlpz/9TKTJjaPTpcSYkLpbIwqa4NbYLJe4iQK8uN6wLLz5YO7DuBacA9Ou
/qEtNypZ4x/EGslAHoPvlQzIG+SbbDyl+GNXlIuF6NKiliiOM8DHywwpSn/q1fKJyqGgijv4eNWA
rBXZzteyBDP2gbTx4mgG4/npNxz5x0nyqFwLMESamBTn9+jhw3it/T5zWZgHgjZX5pyVCG8iExlx
lus711jUtzxgoSGXZPExjEMeALGGlVuh0kt2VPZ5UKypfRI8VfrpI14oclYKBAdqGwjNhBDfl2Ix
WRScb4KFCWtP1TvDNSnM6xDTEhXMNqX+mBUYlRser57Mv0JXclY+znHnVQWPbsRNvMIIJryIfgV/
XCSqEktN6tvH8snzugu2D6fBVljmF+Lh2jINhimATLRbicNG/e9onK2X8meXaJ3qjZK3ZzrEPDZk
GPutoZift7KXOQ9tmvIZRT4x4Yhzs1gcSHhWZT92LCnT4sMuVCele+EXIz1EGOMKuVqbs48n4qZ6
D+yjU3h8XfY4fJ8OuM0Yrdmyu2iLkSgn9guiU9C+z4DPwMummWPRAvI+DOT4LRtsminfznPjJUf8
W2K6SVIY/+T58SKaLFuhD3yjSvgCa5YcreEv/Npa48D9ziE5Oi1kdg6u8DheVPYNXeXAUrbKNTu5
BNJa9wqxX+y9lXO2mc6HUNUQ1wmrrr40ehIX01wTKNywypuxQcXIKGIxgEH2tEYxFEHCF9lTsUb3
6tvEdXYD/Guf3HLt40cmbo/56cBfHJvl+0BejrARoXqDBaJUuMGFgzITXaQrwnYaIug6daFai9ta
MAC9ZLWcBLNa7mng5h9bKLoE5ksAgj9qJrxvhrdtmA7VLeT3qsUsx+Uq46asxc4CnGaFCLoPkGdr
tZyl4dWpkZZck+4gNKBbSLbwQABF98aFPeBA9MER+k5cYqKD2epONFYjmRsy3fdmbdoKW5Lg/NuL
nTXSb4FMQyvq++G4yVu2lL5Ef3Nv93OYiVuwjzaj81rGCkNk9fQpQPAkZwebCFrsGLoahkDKq8ov
sg4VtOiTLCQ7OQRGv+rBa9wJXxjoqMcp/ftbISYohEL30dwK2fITjGg1FfrVs2wBtTXaet+oMYYr
tTt1b2H1uSP6i5Eezh+JN2fwHeiO6pYpgN2ZaVLbDUCivv8hWAQH7158lus3iQrtP/AgnOVIJFD6
yEtsYKTSF7h/P1Hg8AP5YGIZTrXpXE9PaeyV1vN2avpEe/30gfFq4e6Keu3f4VidC4cM1Gj5nxGg
P/hZVyQlSwxD0anZd/vikaewV0WdHCQNOd7ylr714naOLMYgv1shA3ocZXjqrisIa55Oe/JTh6G5
4V+0sMt92ZWpbh2jqPe5Ia7Tel7Iexj06eFQMQQMcv8WcsI7H47EwkQHDuVeE0pdt61bDQG1E7dB
dXkecTV+iBHYw12HBAESgdZXDRU6ln/1hWd4udlXmYm7C3WUWAw56P+HULrZLkPExHMPNMEVCmFY
XCqwBh8jwbrKZCjibcliT9FbhbeJzoLYyFuAfGyIN1a3DfybaKVgPiclWSGIWN+0HBkS7IUjY0FM
q+iIjzukf5rwDf4D/0cmLewhQS5xAe/crLovu3CmjJRD3MGTWRoPYT30Z6QW8HIuYUN59H4ewxmm
I6xwI3aRGa15k4hNwxcgq5aL524C1Px8lsfsT3iLgRBiSgXIefWEHFyCb3P/UyTofnZsUUaPzjFa
sVZoniXZ0Dgfp2Z0DKmnAS8H+xPzGW2XCgVvgdR9TPbhy9Qin10TdEG1wCrsvQEqtn00LJN/mEkY
1/isaO1W5esUWrq/I+c3EV19AP+0Ho34gi/oj2zRxuWnmxbtHlwnk5L50o91eBYhBmbwba+r0WCQ
2Ssa6Kb5ZaLY3yHWFqNKQxZDG/kbhgjlzVG9aWhhTuc9G866f0kaPHguzYuyVfC8vBvfFU5ZTMuS
o5t0JvCggnRjqSANs/ionYsmTWbArL2k4WUmtYAqcxrFgsHfjI1eeVXI6AxCEncYYEqqB3a2yGQP
vsgU2OGDSWU6qfT9uBqLv3OvapC01h9UZQIDOcXSnIw8isxlJcd9MXb2rAR9sbkDyqk+4medqkYW
MbIFXYsbrsaKW++7mgPf7MFKklpvWaEwpdjWpaMbR7VJbtShuB6z+yk26fWLc4WnmHF0CvCVyV/4
v8QNtaJkbGqkm9hCJXnbuPwt1UahZ8FKXWO2nMIS1LDl5PIm6abjPOEHZvWZPPCaYYDtUuprt5gV
jApwp18YDMNwSVEJVmIO7frAtwHe4iiidOZun+SaD2g9Z756CzeDgbGn63vGJvT+UWwsQeH/K5TL
VqKMKn3bCxhM/4YsMzNdvbOzTEDUTOwT+oK66yia4nyB3yU0R5/9o96nD/X4aE5K+Yy6x3KXKdce
WVhAG5zciwf5suMI16h7L86e52udqnVu2CSryyFOYt8Kf+FxJrixnN38/Z7nRGBpcvS/BepHAQDz
PXVfmGlQ82WjUV9eM82jX6UgRc7Kak39D3KQB8hBrSCc0JGm/xecTStaAAv6F+71b+BQDCXrvs4r
EGTmeuiSd/kvDssr1a0UWwIMub/AqXf3zLNHYTViKG6OAYrf7BrP/m2K3UIXeBjKGkBGTLLEoViR
vN3eKArGt9/j/16AIur9JrljEXa4m2UAEaz8t7xNBW3GKtuVyVBX51AKcGGkd6BDfhw6R3PWGa3T
DaPOJMo+WrDns2iC487B0K/hbSB0Rcg8vUAwFNMwrkaV52Nb8JAGOFd5EEjGPMSjPQW46IJDNcfU
dJXD/KKiHwDzWnI+zMHGqw2mGMXKrjZ8acBUkIEXhWCbDWwm/Z+JZmnM+2CcLOjsvY3ynKNxl94M
aU1njyRfCoqlgPyLR6dPZku0YgWzme7O3Lx+t2MdC8fpGqcdRxN3gybViUA0iF+W1EKCow8OsKTn
QL8fvdMpF1Tc2MU6rN/QgYwLOTx6Aw+iNiGyrQuoS95s/X7DzLrtjurocEB0DTmDrROP5vLxNW3I
AjVkR1JIsWdp1QoSADY1H02bxFLeVGxTGee0xwHGSUXLigQCMmulE/+vkKdksOjfdHem7wy/U3Qd
J7edNx3K2fbjA8v8aF00j5/Bb73DbL5j5wIoFQ0CUUYor9dxCHIr6Skn4QxW7/PTCo5qPgjXfMOO
GC66lb3YDLwWLGGrLTBKzCpLWg0UjxBmLSee2CbyFimRIEITxa8WB9b2UxtuVLALwOu9KEKPfgB/
jm5NCnAXNDq+/4hXRK7KiE9JlM8YD0/MJT3KUlnCC+C8kNDWOmxtn3BBhCnIL8p1sSfYZYXXQ9XC
F7N807bYpO1c9tQ2IcGRb3VcgQ376UClGHpyYV3qRJqGKkGGMcx9EEoJ1bwXKWKsUn4eOn4+0Z6n
GOuQ7Z4XkJBdWX+o8G2vWNdIyrwSaHH1OciaC6xah+p/5IVYfFpD+gQ15rCAlfpLpklkGaD06Mto
fGSosrUQaOI0sX7iikUmLihfpSU3BbEcNI3Rvq3g/lR/zzWX7aMyagdEYKuy8k/qY25Vzw1by0jt
CZeHIHG0xLAQ90SJxkvvsMlnPIq9P9vp/bCLT984ZpITUwwtojMG7OjN02ufd/V5MtH3M4rjmwjV
utWZTh0bydI0Qzx5wkM7xept4MRl+1nD/VqWyln9QvPmxirF/iPLvPZklIIte76bSIV8w3cjWKiL
jmh2tOAqXLjD8jZmUaHVr2Z7TJlmilM3IhAugXtevOrG3c7fke+isL0wmxzoZBBqfaBcD7fTBPrP
zODs7OE6oDMRcDdSUgJA+8gHB0x7X5yvh/NyGjEhfLfOpNhZXQAQqjKbsJWvJX0Xi7InME606s9M
SMdQGqeJyU18MyHCPSxYfC37qcRRcF42vKQM70RPo6xUOBlubiQcuVH0GfGWT+3bmgV3oO4/aEPJ
UTDcAPu1cTZ2fDXAhpF/Tssk/rZU3bc5oEGKPVLUuyjzYMGAF/8al10vd7jttKEfQZFzz9Vnjt63
ogeQi+fjFGfrdMqo0ggLuhWG+HAcqFw8Uw0LMGYf2W1NQpp7OFWmu+6HrnS2siv0EsRrpckZ2HyK
0flCrfNkrMyagmyHxgbXA9R3QSV8ILSK76iAG/eMboEjrNP1BQNJSxtriSIPMG1u12QQ9+v4LVA1
RuVcHCqVClhgE+h59fw/8FWtGeqOjEhF/Z5BZKhi5gX9bFKTlW2DTBBF73BBaQaYFROWRsbM0ka5
Z+Q21dQuifAsP+cLUbCui/aYhtmGIN4zWUoIxjMPggRSwL0TQzEdTGD5M1k+qvMd4cnywWYMz2H4
qq8zlhli8E4HL4Jb1JN8vkbHDtCUCzD19O6kOxLJ8nwq/2nHM+2kWogXRz2dPulgnQgFOK0dCmS2
f4XQ1eN4TQBFs62HaKSmWaXq+KASoEjPhw/pQHnNIM0K6eEeb4LzipztPa4Mth41GCHgtyvWeI6p
EAYMIsPUdicT2UgRbSINXYiEjY6oEQW8IYQUddD3rPoYuRI+JDxXPVcaHGxe8tCtDvu6TsGkMGlK
AhGsoTLKnGP9hRpCOouq0ew+Prx07I+TE4kJO8ZPr8fslZU8+03udnFQh4FSqn6iS2BY63n8vvec
sQsKgf6SC+FGjN78cUZsT+azIx0zetfkPlbL9AMXOe/81CNOfzI4XjYP1GcbGSEKt+Zn+r9lnifG
ljrZATCkW0wTNxYznjKBiF80CM+StziWhlJgg1jZ9EBpJfaiTeW6kbb8b9Rn80lnfHY0lDLt1AV4
UkuPAQPFBciClpxY85Cj9IDK4O1i947OIpkXNisukSpSASedZQxi0DDxfJI/CkD/ZvPXxNIzaELy
5ccEywJ8w8fRWah/4GlGZC5Km6erXfuRCTvPMK2Iys/JMxFVy61I/o3bLzvEl8hIozL83H1jeXe7
oJfB+l1OuoZ9HwlqQtXqc9ddg1zPc4EyjvCD0nhFCXPZ69oqU7UWH1N5vR7ZPfcJ0G6Rn9L/OJ3T
CIOZc69J1jPOeVug8T3ptvMHMsC8iU09gStLAF0s9oBjWWNKdPbuT1nPFuFiejEKX+h83WOxezWU
42R+FYoSeT9QId9sWUx1d0/LAv692LUIH+27jDws2vnymyF75yRUXMumbt4iuwGwmG+xguV7PR1G
3CqwdxNF6hqTkArzHLEXuhTikXpHaWZUld6wNo7Jwql4dgl5kkjOOMj1mYwMqulVQzBmPjTCTDxB
cr0Qj3fdZut245l64lnqFwdyYwVZ4yo3pLrAI9H0ASyxR3LHum5BLzhiJY2i3Y+MMnm61jpWXABw
FIdESAHeTYafC4EGiT6V5w4HKgXYkNySWJfEtsK1gwAaLi3GSdfLyIu42Zk0a1xIDDP4Jzmovtpd
bWTcNqGeGlPpP0O2SJwOkFo93fR1JhTGfjPto7YF0fsfIlVxmgIJM1flQrg5S26MY8trzUktNuX2
FwahWP3OGpjHAHVGq/vEr1JwtNUbf5ntG8rO00pqkKM84MdHOYcG8qfoXISvWqDk/7+Yi2Wi5otV
ILj/vswaTX8umwadyZ3ksUmN/XctKD/86KtirGatRr8PRoC9JTe8XSIovitlpunz920iEuVpUaR7
4vNOPY2t4n5KgYN1kU8CxRaK5rjuuLpFZUmsTeSkP0cZqSE+2CMk1Npfk9ZtN/jV+b1nA4mavyix
xMKCf6OlM/yv0Ad6uBxIW9oxekT+uNgWHqK4dwVWb/55J086S6j5FrErQaKPtH39HWXxRk6KLvQP
yrqfC3tqPsOzxZ4ekQpuBjgnDrIYVibQorcIpNCsLxZhMHCYwsA9cWFJfndFhlpJm+yRfsx5rcQG
2QZ8rJD4kphci/oUWOWZWBSq7SfxXlVRDEKVU1+Q/HwBfaqsNrQDMkRUEuaDhKiGbSvHRedKxQtw
ZGFKSe+djdCZHlwKr8TPT3/eEBAgEZegifMoFzmIDgriGDELKUKR14ADYJwtMQXV1tyz4Nl6E3MM
aMt8nr3jfO96e+EF5mHP5VOLSuDzFZKi0ejlQ5Sez8TLS1XjRquj1bYYRWRgl47qy21OKGogK7Lp
SyFguMDkKXYWl2lbtQtNa/zIk2QStIl/VBBidSYIcYpDq9R7xFLcyT4sbsnA+DoT2xCEA87rvArM
51lvg/pjDX3DRo6B44t7jlyqgn1JowWRy3oBL6JRqlQUArbm4NBFX7KeiCZO2GKxRzNh1N4u4WEz
U7TeT2ab9iah/BEogZJa6DiDXRqOKgQJcDUrup/rpTtrb/EsvtmNmDDs8smzzYFjhGX33H+ZI6yF
YNMrFrfMKMO3rgaBZrzQQBGbtgsRlYXViai2Q4xAhrqzDBnaLWvURC5yYuFeKd4HspJdvXmakdD7
UTtC4w6/dbR1BMfw3dKW++T81pAbor/c6PSqiIM/57WYFA/b0AAhed9CIbGEj/2dmOWO+FiugbNP
/iiu+IAryz2VwBVY6H1ufvbMmZlDF/PWmPHkI0dy2QR9wFNnXERizzZFrnVDtHjyApsC8JQ48hsI
isEvDpO5eRa6GxNJFdzdSfuVR44KfinXsGKYbR36JyW+fE4VakJjlRTO2YbBWURAXqmhtQOw0Bu9
Mqe594up2GUdC8sC3WJeQNpki0H3uhK0c6VCaTxTtf9XEZ9EhUsKvLKOi9fA2pXy5EIALDqPRA1k
ERtjVk3WQo+GTwQOBU4BqeoHkh+/PcKR0VCJJcEjeMEiEKbmTjuQYQR03utn2gehzdhnJGvJNEXo
mkpIEr7cg0pPYSeeb2oStlxk50b+vnPYDvTigxm41ZUkI/G3eSCv1441AaQmnYGWGJyvsMwalD+T
eF1nRDod4JYoOwTeyIUUIFOZ7TjRLpDxmdpCTewYyAXrIzTiI80JVN8jyVcXQHnMsLpw/bpr3NQ3
qN8tFDCQYxHFKUsuP5kqfTnDN0FRcINkuFAXyT5xqpG3rDNaruBx9dPi0w+Syzl1i89WaoqJco1v
Ht/iIOGJnUOzYy13jD0oAX2yryBOPDRz6QL+vUK2NedB+bDNSvr89w4roFhJbG5XI3mmfUWUnlsj
9tLZDg46tym9uvmJmDX7VVZ5LIZ4e1w/O9fqgrzqaUFZgBaL/0yCV0UcmKByEcOab7GBtbqFbp9v
fG9fDvs/uu2lmygES53q+oDsAJDpAmPbSasJcDyRsRbUsTVc/VzrHoV17VGl6No1FMEjDCGJduY7
w2qbF6uY7mlvZU0q/cNVkxQDymeGfnK1rGEC3S2DoqPQW0ATPRJ8FYrobWmL0CjRa9IF8eeP7fdC
Sfkd3c04WqNyNx78Nr+Pus3wwvAOtgA5vYppdvld1YF4DzIO/taCIxDJN0I3PX6kpHarJi0O0hhf
Vf7cAJclxIibFe0V+7kQ5uVTKUPuGtI/dg4pcS2v8eJWA5LJQXke40Of9ZUday4BWC+fToGcb+qg
4s/vJMw7V06k6WalD79N8uaIBpziAdo4LCII4eVEmpw6bbqJWJxY1Tp5D80vPxCi2pql12Pup5TQ
oJwRXljPFiYRLOxzf8qMgKXR3n0ixiOnBtHX6WUk8ufWWxBfm8vX6nP3MHVzfTrgtmoROol8+Mo1
3uqw5FYWoM0gmR5JwgK34jUwEDZCHvI+q78zzky4wBJSueu6B1WQZzxCJ/1SYRav3ls6y+pg2iWM
n/B1KP/SY3WzaNxddvz+lxrIdLPWu7YqWh/mQXwlY7JezybNyHIznPn43fK5r8iAd7zrN1jzqQHO
0XW+5arp8xKqCuL4W4+knU+J1vFdP06Coqcwa5SR6LlnEv9cMnfnZ+LW+MKIXmJbJ1ajy4Xowj2a
DbVCHzBjlioc+WZF9sBLKa6ZAoEvCdDb1NPovGPNhlENNhq/x5Jxv2H18JAYvDqiYYbXB5ZRm6Yt
uzdC3XhP7KTwbtV1tZ/HHgTTYLwJdQ+jwH/xnSGdN8+Atz+bOh6GiJidpygCzmSJ8c5GAhY5ckN9
rRjW/s8/Thmox0KJGk7ATlWS+7pvwEvFro063GVzlD+fPKRY1z741W7YWrhG56tbmqjd8qvdihh5
/EUbku5g9XmewRcbH+SwGusxPByXWkHSLE3NwA01fezn28Ix9T3D3BRdqeGEpEP5W/c20WOtIRD3
GFfFdlujRpEmfvn1w1t+Gqs0EY1q5h8UsEUjNntYfTfe4JMj1+gMWFF76wW0+mf3AVbfWA0DPtm2
xQrvZJ+/qlKfmPqRImE5xbbKsgYe0fBJcxoxEcVU2kqJbI9fC4p3kAc9WMf6S8wuVt9cTvOFamsV
Gm9PguZEfB0WwU69zy2/SOphN9L5Z4a6V77/JpYWRLCHW24+Tf3qz9/g186U+/xaUxWhaabJ3jpD
1yc9EAzLgDIQgA+FhkFuBkPu4fE+YbFblqnec3GnWqpiW//uxc8eWxQvyg2RhIvmDQxRBnsVfQg/
nprqeifan0V5Q8UyFJxokuYq74hyT2qRz8YqJZcahkGq+ldEjRpN2ZZBGEnTdxn8wstHIiWT+yrE
rxyTDB6FxCINuYKmkEXekowIbp205dzvhqf9b/7McKLDV1WhcwpMyO0lVoKYp022dQQknf087Dj0
P7aeM7QzBOdZCkkEipvjTjxN3E79wFxl2iKROwrkkALDav16qz0/opP1/R3+HOnUJ5EcakaAJ7QX
deiNIgotfvWRPwKWWP+pAXmWf0kPduJD1MuJV1QGmyblzngGcmeBJE+l67HUwzfFl3sDb3iK9nWM
kdps/d/VoA4601yWVg7eCEz+qTr2dgfXjGewjyscriCuIuUigVcfFR30rG+VgI44lmPXZcFzmAbu
2cRXWqwBHoNAjkZ3VV/UjM+SUYhPauTC0c1cSbbEqrxydHJ3oOHlfiL/xy/8/nug+sLhG9QyOQy/
XR3AIMpa5jW6jqsUR5VtY5bOtxKctDZONd480JwtP3TPtJ8t+mbPEAsz0pHP34dF/E1Y4Z+q7p5o
zj5Xa8VOGhA3qVst0Ea56TG0Y+AUs2MXml+VLshcm6lujVcNQSLwFTXFKGN7OYbmfDdL29np2pSj
vBNbq6x/qb/EvPGw0XWndgAtIg+TEEhY+a1YHgTrw8SLfS+IsO4dB31IDEvTAtu83Cspa81vStoV
yCjataWnl8bBAPKE98iQe8Wzn6YeiQ44YF0DGghVqjWDo0YMS1/jNfaEeTcskyS7tqYUgEog0cKd
loVXXRS7XqEA7ryBi6Z9csGnSk9kyv2zyXolLTje4/LcDXm9qrKqP0eAWeFphrciDfW5g5lKZAy4
8Kedz16OCwBRi76oksZtnH0zgfSBgExT1t/uaH8fD5XVZBTuIjEvnFVLHmuBK5RHpkUN+WuECAWH
0WRTYUyiKqZWvuFLauYqQEHE8/qvM8ZZqt33hXWQDZP4apgQYqMEQa/q7+cOfO8blUPtcRBFGMJP
kYDv2tzHH46ZuzS0PQ4iHn9E6BoGS5fAbPkcQQUqMe3/wdjpl48+XLPVfCrMGz/Uqq6R8S+2tUA1
vfFUNFMewyDkgTSG2zqBMFJHyEHK4efaNbQ7cvtvXZK6K6IysImJqVV+OfjykkPm8eFLEOJ2YOV2
Wug7zth0QYIhlUyfeTUt5xtR7xfsz2h0aUwoIUuZRvvPb7OR/z6RlrchPMSpD6r0+MRpcg5KGTVD
aGUxUWn1UMwyzGmHSYhEm6u1beqCWFFwWVsIOe1U4czVbpRB1yqnz9JtDAeoLG5AASHSwo/exlpM
2I/98bunG4DqE95zZP74JdDMOyQV2g2JRg4k8YwSgpYxLwtnCCOPWO2UtdPTdLBXD76kIwmfXiwN
VBMpcFxaar7553zwWqnleuOAwBBC8FCnynuo17mFajoXFszn/lGfE48Q4FWGK4OsF08CXqyC1/nG
fSu+oiMLC8o6vF12fzFO9TwQv9gP5DAzqPexTqS4ygFdl+aOD8//fISdpUt48aK4VLx7P2wYOTZL
E0k2fmohGqjjrToOqzj26XnQbyf2tzfZYLb0jvl/utLIitwzjeY0O0ACirVSMsoOjF3DQa1ljV0Q
go9dF7n7xgvCIeqzooYfJWIGJ/wtY351ZOQR+PBcj+ZehB/PUkio+HR3MhtLdTlD8jktGuC0pGkk
wf/RZGsJGWXV2J82JrrcyHQkuKvQD+9gF8id+gFgV89t1b4mux+AlapR8oPx/wZOIwEYIpoKiovd
vvrrhS9IcEY8IJZWzcjK1G7wGFkV7VreoqbED9dqK+tUPGQVXbFjafck/Er+G8JJV7OoGbMGQS1P
7Hdb6EXeQGek+t0wHEj6spubJ0Txmm9hycpw6B6vjIVAMfcA8KTO1O+qvchxm1/vAeUsaDLmAlf6
5GBXklR/Bbe03dXc8oQT1Mv43d/kr/Y0Aw2/oyjZK5H9gfJJg+xiwcp+Gl1ZOY96PufNh8oIqcQu
LtoQI+En+JBSBmTnJ3Xr5ODeG5UChKcg14CoRIIX0Xkol0zw74vk5yC2Tlk2wiUC6nwgUeTNjL9D
B9JOt/BfVHMYuZS77XCG2bvgE9pegRfeyjmX8iUDHEqYWxsSMHIPgmWnHQDQmDP6XZUvn2GWImhI
JpCZzjcZy4nlZjOTAU1ZV4FjDOrp4f2LKWTXcC3I4BaLnHZwOYkTb26N5/bNkel1WoChaZw5Sw59
tNvSY34MSWSIupHKFvW8DzIsgNyOzTyn1XYdggDgXrpXPCIf5Jg2WlEisAp3DAej/3ZisK2/JPg6
ZWAwAdbDhXG2IfvUNy/lPoecP6YHodBRku27opeeBCYH3yETVAOO2P7jh2UP2R1MDlspsY4QTeum
DUplOkRBB0jMFpn8iKoboHXKflVx+H/RMIfCQbQotdIx1tuMHI1CWM7Q65VtLUbiHD7hG0GhZloR
reVyRk8YkxwynvvxVBjPkUxmizu7PHr06PmSA01dP1pfo0YZS2y6uq8xlxQXPaBtnt0dRd+gd9do
A9IX/jPLwHnAHYHwazJcAMF7WipgPK0pTL848t5XjJWlRm7Nt/JCnc1RymyqdvAr3U9ZHqfIN0XO
DGSbvW9Z/ttxjOTJAGKH3Nz/tasgK+mt6oAQ9r3psU59ooZouWWwukGPs9pqURmb0Z9GKHkT3IPg
/QllQnSEjx9w2Vbo2dpYDNNhA78lblL8Ob1qFSTlNQP5O3Ij11O4dWiCNBy7WYAOwkzgH0TU8ZYf
D0IqWFRC7XteN7u9WMYp1eYvzghYXYynpEivopn3Sv5nGSFDDSamxsyWx4CqgQbDHECAvdHcpV5N
Ql6sdQNQ1Gn684Y6/W4ZaIRh4ZnLO2PsuusqKMz7mjjmKNCtyaW+sZPA59CcDQi/w5taWGJYUR/f
IInh42qW2ISuzV/mceP1EWrwO2g3KRVmsGBr2PwVl4nSYv8vRckEiDJFpBRjsywMu7dRnmNTRl1l
r4wfTBqLVZQcDNPbLbvNyvrQySRhy8yvJ8IyUt5+ueaJNR64WpSY+CH0pbSQvGNxiHBFbvnd1w5d
9Qsg6+kfPwaivycDqpnztRLzeq610MxhV7CAStoyg1+5M/N/wGqFRMCkke6iTXKVdER/YiHzrTxj
baFZiQPYoiqCXDz9jQU9tvz2qf9DQHK+WJAjLo6ygROAhYjxqTEgNEjzb7jNMBcWl9MlrXnWslkP
O8TDbl5WJuNvxeRafp2fP3pPa4XeZXlzvKOkdp0sFMlU9REmqpXdXavIUu8SAohm89sGy7A5BlMu
KSrCDuEUFcffWf40ITYrr2JPG0LQQ52+rcLDV2RZMFbSlSVR0K29HbIl91aaevlpN/hoTdaoxHPE
0uOjfmieFhOTj0NHIcMJOH14OgWoJ+j+hsgwHksfscDRtts3VOMN2pk7C5PEXWAU44PIKAfw1+c6
BMOGgQ7B95BjKlj+fHmAWgb9i7hH4RXFQqroLIVHgA1G43ncH/5UvjyKrzPUNgGAP19HApL2I8Os
lI7V+wwJCN0hshn4z5r8CNpn5b80k36/41WY52dGupD4JsJ5EV7rFM+/J3ulcYb3p+AMlw1UQ6KN
tpG06YppfeRcGeO8Qf9L1zFY37QY5/Rk7jnNaYu0IhrKFaEBrfK/9YuJdzCWc+WnJuRVo+k6FdLR
8wc4FjwTNW+KYSDyawkDsfv3VE5ga5bOPm1DUy4T92lJHifKEU2wAIUilM//kn3uTvg5SULvZuu6
G6iF2uhd11R+lxT0J+etv9wuAHao3p/ePwDHM7DIJpAPpR8wwrYqDIlOgBkvpqLim865TZTFjbBT
s632mAH/GI5gVIay5Otx5FzdTaSovLjhinVDMQc/hoKE4NSUvM7CS1m3xUSGtuHLdmE4dRP7k08R
iDDNY9pxP9UQpRGuZ0CE4NLexu9wtDy+z4yH7I+wnrcKz5lc6dNsRrYfIAZGLg1s67eIOGBB4Y0U
S70K5pUQHrYRhS6GDUzVOdOdV7G6/ynSgz1ILAmw3MurDa3TNpyHRBJPNLMoZS7lpR5rWJybdYe8
fdup/irmOFB8e48psLwv8kKlLqihZPjcngfmGTyXnZq16mO9+OjBbRvyyABxZdMpGcqWSmt9mkzw
esHioJ+eBvpYM1Hjh6LgygVrfn6xPHt/tqiz7D+8jSnvjPpHwpKOfn8kspKDT5gan14sXb78jI6G
6JjKeaIqvjaEekNs/TABw5Pa+JxQrMpqZoiyVu6k0MA9EUh07WIgGNN+bQYff+WpU+r2UsdNP8dy
5SKw3KWQOi4WgFxSCOf2wqM4FIHF7EjC5BvRzKpDZeNsCDRBo0adnL+UnJ3xPAH1lwUDOxAuhC4R
zhkDEUclhwbGCfmd4iC7lvOoyZgx5Q1xie1lEwTK5QJ4431sltwb5WbyqvpOVw3XTkFUArWQ9QDg
IumW1ZvmWPVBFupFcu1qZoStVxOkOfAQs9N3OAyO1JjAWg5Njj5cykkxS1ZbGaQ36f61lKJlS/7C
P5ERMJBL47X0KSit0tywc8j+tFOPUAx8BnjocXj1aX4gRvx4/bBB97k3uuXqJarEXbs1WuVEhliv
YEmVnsKa9ItcboUkEF/lYZrPW3AzYn8LQWpMefNsoKLEfVmbLPayo57jrY+QAHA7Ze9hZUTOpsbE
tDdRpDnm0M+emgUCSl4Sl9+kxZYbef2Ej4impQ1Uk5MiH1KBDu29HBLDlCrwGycHJd2qsHgabb0g
Q8zXMICDW5G/7TwrnmV5LULsAJloh9newoT73FUjIZFJ/vQ/fuyLF3AnrWJ93R0lWR3ZfbR8vsLq
HHL1c464nvymvgSUL5hLCVwuK+mYduad0XWzW6Lf0zSrkqrt2tq0zCWKuwFGzs87EGlLX9RoB4ad
5TgHKh9VLkb51VLq7A9efb85UqFcA+xkWfx3+g6Lb8hkNkFN0GMeRMxvyR95EpTUgL0wITpJF9Iz
YsRKQdYD8utTdFflgdgIC1owXdvuWmZzcD4X/G6kMt1RECo/Cf8d8n8IpbT6OioHWqaUA59wXy+X
Y6/Rhwu2sQ5k34y91lPWxj8AihoGMJfu6D9VeRAjt+ObZmeMIGeHFKtqRiDS0k+8xyZSEVR7Lva8
qlflkSeO8E/nnYOzfNi9B8VZAMJnWyjUsKx5ojNgancr667GRZGoMwY4x3JQIBba4FHl2IfcGH0X
VbK9Qsgb+nl7F5HRMbL01yfHlZWAdqMeLLxXIa7eUZQUpotJ686TX/MEyrH+l4CtjHXjmVEnkIIu
rGOz1uKyNdFL4fmygN2jsqQy5ja8UJn7OZl5aS1ggK51sFBE1z8+bxi0dhdSMN+Cwjnt1P6rvnxI
7rSv6MUtLdBgPiKVeJYvpfevTDbc8OqP3PKjqYeLQsKZUSie0/L4he74v7ZtGvrxG/TCKmIxAv50
Eq4DBaVle1dji1Wvk485EzLER4UcZJbZWrQLbM/LuRYcHp9ZhORXrnJyVPiQp31TlKBvxOxOcVGz
jJ0RFif8vADoNgNzRgtQpYdgNwmwMXyRfOKSrbKZCdoc1b9zudnDWsfnfrpk/j0Y6vKSlgthsFz8
+tcw33B/saLgJ8k5e/f9QFGWGDf/Gq6nS7H2WlhqeeK2dNtnqYUtjrluTPgryat8QQ4MH3uw+J3X
VzOKJYD5aEqWROGLK83P1Z3MVgcpbpER5yx4/5xPmZtEcP50f+ZkbitmPYrVbnJ46gTF+iAuhiBB
MYrHkCVC14GemvOU5O9Q3YEqAab9e+3rF01yW9IQTO6n3q5wy2RmEHMWMxBztT8xJOTE4eRMHLEk
ImHRnylNOiabv4iy3eyzit1oPR1NSpYGRyos59eTfSR5n1w4xIwWk0auEDX2uwdNWuKjKdm5Yq4q
uJKC6BOveoL2oVCO/YFU4GFQmhYRxo/fTiyR5VfemisJR5x1e32F/tzz7faQroxBU8N+8isqH+bo
tKdnR9EY+tTZxhdx1FNfSWR7ThG/D81zyvpScZEBXE8F/j1Cca7LMLyju38RGJmVEVdpb6D2/XpP
ZOtCUUfTAYDngmT8bOMHIweuq+HLOmw30cE9l5qdC7Fg5IidJ5XkVeSgStdJKyZvA5RG8Ub9ZCsa
WXUNZwJ76dXt6HGsbAlM7VUFc8LHCgNEOypRY7Jcx5FHN3CVKT6ZOdW4W+hNje9pQXH19EUfd9s8
OLa62/YLGgKCB/tEp7n0BxEs5t0Kjw9CYtJIm78tK2ZDHwAtM3Stdup5EJHnimQvo9ayp4rzsLVG
6QegvG37JjH1lxnOEc8Z/gtIzM00ZenM0cRlP9GkacEWMFldVQSRJpHIgBSIky+prJEHOitk7BSG
KmHbmguHGEdljMDdD82Vf+bx+kt0w4Fq+lKXa3T/+xhFbg44dwEJ6/SEofxwadzw9xmxpE/y+/yK
1vQnWgLNcVCAeu1vR/FgmkI6jfaC9rrzqohUBBQmB/wUpyxly0CDCgZKoSewHoeLtUqcCLzB9cGh
7LN1zSJesjQufQ5ae8RFhBa84M+Sj57WSHhVP6bzlYcIEaTg66W9EmxjQqobNnUAHPeyTKJYj1j5
+SVlxyUcvVc6PNeJC75vYjsY2WtMkyu2aV5e4s9YMmYTdjYdYajKf3bRBqiZrQORyd+XNppuh1fi
8zXcrhBrM4F/f++J06/me4F4g920d7eZyyQKfFHxBWAWJQUhVMQztORShSsAvEc498MFr452zcMT
P6jVigYk+ZW+snAo2HgiKXCVUCI9shFSYFmJ4fA3k8CL8f36nnm3d+CduKmwHEJg6mIttChgvcjg
4mjycoi5NIPc2nBPqOI8iJecLE6JfxRjZ+iX4MASBxrwYWaDcIS1EzxU4xJMW+M/K41ndHF9EF3P
NpVnMjaPDXubIKpVRK7zp6nYHtOLmbCLdP5XloC41CH2by/hSC8kgPKPPjPmKHu7FlQue61isLmu
Z0ZGyrmx9Lr00EQJhPejOxFcqadpNDumStC1Ros8TXIl0mRFTIFTZ2YLk6ygdqY1a3tJKoh90zTn
L6Npy+KHKG0jtcb1mT48AOgtc7WfxThdLR8e0o+NyUOzReUT6Au2fF9terARy6Qhpzby/BVNu77d
nw6REEJ3ED9l/b6gEQ3vjbesSq/hEonGnBT7eYNGzrqnmn2GvCpI0eW5hSQg7tEPyDnkeTfDHkVg
Lngf75g4Vt8//6RQqUsRqoA1TkkoMM5xMkm3CfQ8SNXpvsibiUJsydON5MEPEtxDVwJ3oDXO6s+G
PgskfHwcEPLZ0ziwYi3aMI0IM7xpbVJQXBK6SMAz9gwnWmlNanRDsdqJ7zqXErGHfCo7tm+5kSqR
YiS7vue5nqtMBHgyes5iB23uO/SBTxVh+SFZQJZeIfi+TCbGNAb4b4TCHk5Wq+n5yeDqTQk6DlWY
AQLWMWmTPFF2lroBqGudo6E1C05XcZJ9JB3rtHMPLlDaSV/BtjQAO/zTpvtQmZYblsmp2PdgA4hn
jCSaigxVntClmaHiD8SlYRP2lyqpKjgVgb+XrLoWwux/di8lfiYG/L0UgzPxsfnlIAEHungAcxW4
glAnt2e2kop8cq2P7dC0J8yRAPJ60UdhMBRjV+KjqSnn66twNuKEUn84eRF8eKUnSkS1Pv9ZPjKl
NjbTdLOpy+p8xo66H/1JYWVuRe9xPlgC1O6s4rtBCZX+q0zMQ0zTUTkIZXZvUuYttgBGsL+MuoRX
x0BK1JUF4GI8IOpHy1Ke57UI+/Bl1FKIWurSXuKKgxxy00BQA3vXUOt7vURTjoRw1GTzYXHBj8Jv
pbHYSB01jnDw7aY3ZWV9um0BQgpYugcR7xHSxDvcneVwNcZPENZxllKSRMfbappE3pJT2v9lXYAj
n9K9lP1Vs7xgzICrXOX7QJxuANz5q3XighM4erK0ZAxLFHKL4gjpUa+U2aCK4gZGvyHMFUv9c+bG
LMdSkPSzhZvg+ITszL4ukBYOJfHQJBDDdnvPdZaWydbjrHts+u8dT6vQgyajq4iAO/HMPy6S6iyE
y6nt9VZ/vqIpNFP2YAW74bQN2i4sLw3FviQP8Tbj1jTP0yDFZ/KuczhFcaEkIctQ7+E5/VL4zmP1
egvVrTYiPtnzWARc7edkyYKuih8AdzminA3R0eqjqaMfrtc2Qr/l4+aIQzYkGsLdN+1CsDqvAshH
zT2RgCUqmA3VkWKajyNxgm/kZ/ytOMHIPD0lhNxTlsp/5+JgDIr0HHWbpDR5OqclZoxL/gI2I+pk
YqR04+a6DAZZeyBvGPM9UVm8mpE4/OkUvpYhfJACFNUBzgR4bBn86mmRxpWqamwX5K3Im11K2oTg
lDI8c2pYO11p5bvDQn5ChKKCMqispe/GhfI2eAScSHs2jLszEgAlTHrB8MGcXnjJACLabVNWLWUa
GMQS9YuA1ko2XBX1cDWIN18C8xcyRx2ua5TbKAqMPuyeWo7O12zvESl2z5QfDpdH8eyT3JfdBtJP
3QkYqh+n8sT7HpAn0rursarmZ7JLFl2YmYpeGIqRogYvzzNj3m1YYEYbeAQbqeXRyV2ljB2yvzXo
+slIhMfO8NBXOYRny9c2enoiUghxQxoD5CYg3o/UhMJWtkriRaF0wxUcgf6CZoCwf3Muq0lWPMyV
XJTBbXxVMECBtlMVAm7auVy/fS4T6Y+CVMICX+lpdI/PuM22XP38wbtuOiHk702eOa8yTEwSB20P
r/G+59COR9RMbXcT2hRakrOEeSeKgGBZZaGMaphvwSftUfQkaehOVu/9ARfkMpyHfeZDCJVWYJaD
DJvi6M0oyUCA7LnGiIZfu+3vspsLYsr+gyrcaGD5OorvKrIO1Xt5mzr5804HlOu962sX0ZOam3CN
ZWH1K5QilAJxa7N1Cbfl8uLN/cuXqDoI9YxZRKObQU1WS6u7q0vp3K7SEKFFrtx4R07qEzOy2M4p
Z2ctg9F9henZKENQ0YYMAnAsp3YkYf3btPZD0QD4lvVqgc8BOxIncdaPWGNa6a07YMZZjiG20e48
ykEEWyCufRY2ie+bcPXMeF8IcByei7hEXm2VUyDy4jbmaXj1V//eYcI+2smP7MJAuiOiUM/8FvpQ
VMGkLo5biMA78DtQFxCuHgODuxF/z4uLmO2GwNsgP1l8HZEb5p13B5MkA6R9zYjM3wfqUQUKgZl2
2tENs41cJCDOMnbQRGNanLilgyliYAfb15/Xu/hwTo1KRt8znCnwIDDY7onBjus2P1kGyKB4Qd79
SQ8O/Vk8i6CsxD0sIVxWGbQ+MrkD3kITWO5XrkSMfSMbhfly/2ahlAVC6ZoQBaojWhOnXYnYTAZa
aAOhGH3WrY7UxAeAeVizWzCJwIA7LUtDJ2ItfYNNhurDiyq/GIa7+CBjJlYLMLYfl7XkqfWffeGv
TKRlFXkA43diI4Sxm4J0560KUIj289aqDiBhgSJnusDdrWvT/iWauv/ZBjkvttaKpScLsRK8LdAt
1S8Au44k6uxBUIVr2gav6MymTNoXnpT1qC2G1INSN1kKxokoXdlhyHugpcWNU5ZDlsEy3RDkg0ND
bIB/SW3hkLP+zayQFGCAMz8uLyc07V9+zcjlKHbnyK8wX0oDEnRl8KfK57txyTIirDJB05MYSpaq
t/Ff9yC0n7NfImx6PazlEldrD1+aXHHCLmpkL5MRJm4tVRUERqaTOsTRp657cGwmYjX8WwDEPIKq
G7pO2H5L+I1HGspoeE1kMmZg88E+r7K39R1pOIBaWCayL3I3PIcya/l8UkIv86ezBtnqIZdZiZgV
ENEK4b+WnBGqQajOdykeB6mYwDFe08saGA+ioqCsLjBlWrKxERbrAbF9dfazT+kENOHTSwwK8jeu
31FlyHQ42WQxCJ2Y3eQ/T4qzuJAia4q1YTaby5cpsBr6qHJkZSWl4tV0/O5jtp50tGCzFxbzVZO/
Tq2UwEGBfy3tgSK6UsbkInguGZuU6CuEChXu0wP5U3s+IHwv8emX3hLDKji93DzkPFF9uoO8oCTT
QMK04GsPIahnXgA8fC2eK9/yHUaSh+m0I6nhr2abYUcqvYwtf5DASnVsq0A2nKmWI2ZxJJPR8zCk
KvwO10rQBMFsltswVN6bBXQ+zZ6+AopHHW4TRKyIUCZeEUA1tbiADH/M1KkdayeyT02/nsQsZmny
YTmRLBdSPKALbj7/Y//5bx5M9cvOZghvIwWAlWNq+SIFZ7mOz9hrahPrPzZ88KpNLuVW1U5Wv7xT
ggtTs0C+Ongpv5Lfrkr+wAkZ+H7Qozuz5SQiVmmkuQVQxSNf0Rj61ldFf9TNszdp1MWVL5m7r/Cn
VEv0gEKv8IchL33gwhsT4vnm5nR+cV1+BVwqIJAWIhgs/7eZIeCewPUmopIcuBi/GUXHaIgEN56v
NCZ6jbUIJLPEscNs+kKA7xO4vjWyQSLLkto7DfT3Pwcm5pChuAXKzAURIgqMzvkxlPDmvn8uI8Id
wMFs6clf86p25Zu7HqvIGVUkh79oT4TS1Oi6PjxMxNAdyQGIA5RVjMUdoK0YqI5sTnFgBBLd+heV
fpPHMvgtxGG5scuSeAa92z5vTGWGgudtBgUXpboF9em2A271IZj8lVwHKPouCHft7u1feNwM1pL8
vYXm6zyQg2y8AEQZy6mI9ZtGfwPPjqebWlxtWmw7WSKLZLZMZLEn6WI0t1JPC+lWTUfKD1u4y3Xd
eaW+jU1NGnzNyjGp88lRw6es6xD9U/JWbm5Asm7cLNPwv+UxBgYuEtUlbs2HOLGtPGcCJX54gxv6
yisaQgw6fFeKcZ/UW/YzG1Zq6qg7dJ9P+eJAw9eDKwgV/ZWjMhoQek6EKclryQXQZW2BnrWf7q4T
XpqPbPf3k4WX36e7Ddi3y20GdGqQk0C/FALpKbwXvXupPqu/6DcladE/2ZTnTlmn14/0glcrp0zn
VayqiwY7UGm1aPiFNk1k4CjvWKvwuU2HqJdZvJgSf0Si++SkEjLwECDLSjt2R24PJB+WDHEnbLdF
trD7ZmSvvliq07ztCaaGAUDBNlq2c/bZa87n0KRkF/lmFalc955c4sJgaWnH/vobEBwHhMjIPXuG
ZbzTeqiwrL5vFxdBb9w0KpPTH7pr63UWamDrcfcKXC2H7osDOLVONVGtHpYiLfoQROh3/3Ht/fo9
lEfmkMAUF/DyVGINocu051+xfuVvz+8QLmusaPEHzVrooe6+HI2Rxx3+zmUSH4mny5c0tYvSimC5
4z5JnnQxzAyz3BciUGI+r4w1VesuX41SvrBzUbt7qAEb/khOwfTfGTVntLh+EtEKy6WcvNHTgqZ+
U7bTFj+W6nRz+CapcsffKEzKnwWXGEOYkVnh0eOLhjKPHAGJQhfCdUiRGYm4ZjcUzjS6ia71sQ9o
qyL0Nd021NpOkM9rHoqRs32BjO+AhJdCe7yctLUzTThcBvYHt0XqUUlGDIuWajhatk11jrx/95O8
Y+rXkHxbQv6levT3PNSvbnmAvqFkjYJx+ujesZ0DeGF7kfInhV/u7BHGFaPilqslqpW1/mTNW1MN
g8vKZeLDrZIx0t/sQI+LxQHsiTg3ARevLQH77jcyGNFl2MSzfYQtWDhVORddYaLPsy/gCRyA0VZK
Utruk/hyAmNsqOpRkCUmJPdesb0Z0fY/Z0Hb+31IY8EzO0QD9LsGWwYNJL3Z+fEaIT9PEo0M7TQp
h9Zy0MEwRijX0JUD+w0t/anwTpOnmk16xnFpX7EKz3isZqEPbItR8pHNrI68co+U3oE0si1WGu5+
6HB8VObctP8dTezWWlHMuLrjjUArQS9n733hx62Cx1WlGGub1/6oxz3Bl3Yk3kDkraaQEYmlWY6u
DEXaeT3ELDthkIJev+JzxDwoS8vz7vuyIOdlZRKdAkOTokFFXTAA2NPEdMRBXE3eSyMHHOTKPj/c
Tl9l6XvQWm92HIQdYe31RChzN46mGojhWjGnDumTfwsFzUFPs9uCxQNYPKxfjFZzZqxADS85MiQa
kjC7JVlFpLgXEa1FRxbVXe27g5l1xTDjOxCPX9hMxEFjzR+0lPgwBt4dBunpADyUBJuRXX4TtpCw
eje3bFCVGeVXXvVw7WtChfFaFM3Ghch18gGW6T07tcfVvDrKkGWtyI/2/XCAX4rqo40xi/z279eK
IgVohnRJWwF9peUuL6uMf/mB9LGIPyKeRBsxlrFpMiR58MLGn1z5YgcKbpO74UFlJjXNlIhix6hn
54lH0Q3TQW+EvvfOTMc5UudBlnmOhnGoGl7i/xMuy9eTOlGZavQABqUcdWB0jSb5aVb8oNIO4W0+
PUOqYTBPefNwSjdSymz6xKpyHcqleC/kRw1Px4ThQJ87m9Jiv1m+w9Xvu2MaTwf6shK1KhfFO1NL
jsPtlf1sSymZL5XjJ7XRZ7JZ+w7c7/Qp3YSSqN+XI5nQU4O8ch3i9Z8EOWe0tUkzopgWEL+8EJ8S
z7Sf6YBxt3zV/RBkm7gBdGuRdgJQGeCYzftP6ycZ6DxVr1mL88CziMmQ17JHSMLF7PkGYzZzj9lr
VfHy29RXN+C8JQSj8jOgoz8toBdlQ+fXkJVqrCQmC5K/sp9J86wTjJh41QrORnId+5vc3GAtk1Tn
3NbklSf/rNpe5UTo0dmjDYDiU1ZmjRvH3pGbObuUvBtNn6M2WjeQ+GadDEcHpTCBls2uVUCuU9NB
KmKzTnPHaQlZqbejAOu9JiqPlTh1H+Ao0QOKottetrTJngWSM+NcyHo4TDEIJUdJtg1A2oAeY3ef
q1mwqEOK5KA2UkbSsA/cT4391Qq8KoykmoZeovffrjzHDKbRD/BpDFwOf5Dg6nwEC+b++Yr4Ehn3
8d28uXiauVo6pm4PcwefzHALN1ZD5jZsvJKDMM/WQrHIWzFfqCeyFnAKmfSRpOuQhxpRl3ALZz1g
z2PbsoSgvH2vDgH7tIzLkcfbtqUGw4YtpwGmDyadDqRn7cRLZCDVwIWcxlC6DA+cdbJTIYqIs7mn
hYmjdmPhmP4022aips+xl5jZWWYz8PV0NJ6jd9QtGPi/sB7rcz7ZF+Uj26YwqC+gNGolIFX823Cv
+9AV2940ImlDSTj1z1WN8ZNVpIOS0IItemQ71Mw3GS7ywFIDpx6rZXPAyZz9z6fdw1fPQf4NUPIG
7/n7+sWR/PyEiUOfS/JQ8KBhmriUWLb1C0cJEDvMB8t6xyiyCNCTEjxS62xbvoYe3E9/imqiYt5V
pkIaPh+vVDPeKwTEZ88KgMK6otSu5OQmBTo1eZyt+t9+6FVxiCmykgIXRPxxxf846a13IbbjI9mp
RN2t7rB9b6FPKHsMc7OEMFN7O2XB9ZH1+3htGdh/uubWCvWUOrJMgUgO7y6E/troADypvfPZ4BND
RxnetEjSkcDsz7979oL5zMEoYqVZUHT9XFlqOUHgEO0SZPDVEaNmtFj3UAIyyexGkN4/M1Q/D9uT
FFlc3QOrqsrGzq+Gq+QuIUYgbIxmkKU4+4hkqRNVSQM78/VV4CMmpM5LNpcuLEamaTUymYJwakVM
uEwZb0oMLrR4KJKlG0VSHSfnRn7Xl6VMHeP76WyJk+p0HWJrA81j2+jssqgyM38w+9rfiTcVsKfg
4u0l8lhFck1LnBT3oCtYWrjr3OAQWz7QUqeAkcFY+x7bNBUgGIxJ+Cm2PdL8eGTUEkSnO55k2rfh
81ietGrzmjNr/4fKDhgBDqSqc/VH9A1p2sACh/4/L0OXyH6pucf93ARGRegR1Eyl1h5a+uij7DMZ
92I5qgSheZsUTLVs6bcxjNpkalkFDcYc3tP63Vb5aniTTC2GucnZZEuob9aYsrkTmGAVFsnPU2/5
9d4yuop2jOQy5RKgdtrtvcVJVkAahKscjp9XJz4fjO7MPQV6RV3YypY16pq+62OleqSRyI88YYDA
8aKdZxvuo4WpX9UHPnP3T4d+WTaeYdqLlzttG0RhrZ2Wj550ioITz0dG8/oQNA5g9jzvxrQrUCod
zLpdF/LeTgH598B9mpMIq28xvKzXBvJra3/aH/cYoHYY/sTk9++vGACi5xOAWxJlpjmD/lK5sWKB
xTi6MNQF+lJy9/Tyg/Gl/2oXhA8TBAxhvHaUYyvMd7XMQnhiVaOMTqQcydMfd2vE8hy44IGfGYv7
VSBUxyPSgmtVUtd//TksBcSGzTX45hrCA6Meb2TTTAACEp3IJlDsbdXFhePTSJMMVLJC2iH5MgmE
70qXzKklZZX9EBbko//0BjEodAewLaCz3xFDitVyo9wQ792/xCAhmkB6NCZQWOHoC54T4JsHeKyx
MIFBTTGeH4gZ+82rY7+uCtsU3c4EDvDZqgzWRUqxqmFvqFOZ7V6Gakkk59LktjJTAfK67hE1+6WG
lDBHxPrlv3blkzIDjaZDbkMUry3f8xgRZLsqF3AbnGFrhRNuv2ZKezIAl+xkE/3AjUffYlXshMMu
Ki+9EaLaJzOBzoBI8UlrPL3idbarwdoVZz553jdnAWLjWEbploQ1zr2FE1i7oSh+h+N1gcsghYEX
a7JiomXIDYFfds4QSQoeB7apzb0Y/o0gQukZVdtd3vFg8oQp38EC1anjW9jStGSS5t6GbVGkyefQ
AMQRsn8S5HB4tt+/nIkAskNrW3S3Ubcg65Ksdq6eitx82Ya4cfenfyGd0Av1JcQqMp0kobfmfgMl
xS80kIs0596587qC/8WAFEgrqOCT8A/Rz7U63CkCwKRTc3C4KQGiMtnqocTBNMEYiyvytuLfQPIs
RCmHm5stM7WTKZTY4DorpTS+eHGUKtZH5B5ieO5FRWNzuBCVjms/LSH9n8zv1hqMbX58u2P+I6Rw
otanFkR1XwuuGL7JfE5hWyLH/VMMBgIpHseJhna7O9ZCnDP8veJ7VCUpwII3kTrNhU5z3VtY5GG3
DvexDsPZJCgJKvUp+4TuHp3MR09hYxddLleJOKckU73je3aiOVB6NZoKgoHWw9zar4rRSaonQ8r2
rtlYCMfbqUF3dogKbLr5KR7VVrfqzXzz4QTueJA60IQF6Zw1hVFFJhZplyeA5/vZqRVB4NWJRQ5q
reZvJ5UT5Pte+pSz5de6G8ArlOJCCiKEVdSwj5TTkphl0xVVVsPwzOs52Q8mlenIiXlTkufcqws3
V9YoCPe9yUJVzF8BQKon/MZLGAGbANhpo4nsQnI16QfYba8jfm8nPkIE8GnWTRCvPO5yeDUoW1F7
DDxLXfJx0eTaGt+Kypx9f5Ckbhl0JQ2CX5eGKyXqLnWXE63KCXEElLHLvKDnYiNlz0SVevVokXHO
9RF9wdJ39eyLe7qNhKWN4qIM3Q9rBNCCxRpdHRE6uIwNpVU/jvs4/vdVZJxyL5qm+q2prdCVIGbf
WBo4L9pMcGRXtamjjHhmYILwfmsjnC/XZJZSNCj7CA/TIo4B8A00b2w9REbIS9lbN0T8OfcomIkN
/1GDwcbdkAJNZ47Qb2t29vxy6ZjXruH05aaqYW0o18a6H1aXGUrJYU5Tq/r6djv+WrO8z4wNxZAr
wyR4EgyCPI1wchspp4e1hbFoTdJURhd6DDcMELz61GEufT7HQMIbKvTwQOdqFi5kxxaeG9JNXdbd
kzSHIE2VeIPm4qpe+aLCAVLnXEevbNwkgACRXRbCNXw1mGzVTp/Pcb/Q8S+Sb+9LMB71pejwGkBC
VgX643D/iNJS0rlsqp6kJRSxuZeZgVGM/EItG2iUiJt7bjY2YgPvIC1GyKbwKgKjww6SaTPOXOdk
EwLXxXRG9cQcVhcF5MX/IK3rO5H+iuZZSo9hTp+6h9KlTaTMhGdVzLS0nP/dO9q1ctUVcTItN7Bp
sfHqGdY3DMVzQ4Gg9w7/UGgbol7LbXQwlV0rSFruVDru6Z9oB6fu+K0BCJrTK5QVsamWOlg7PO9v
+PTZdzTTsHXutynRicYVJEXuTisNmwke3D3RMSPnRnzwz8N6aDXMdu+bMNORikqmrX4GNHFPZ00r
XNNWRuVwWlmB61gFv1YnBsite0rtOl8v8yQ3t+RYLgmrWXZc/2Gv9OEevW8DZft3kubs6zg5FFVI
j+NDt5JlMhLoR77c24A6g5Rjzucl3VNsbjMekLHcrM8dR9FuyKppNWTBi8vyo2SGOz64oFYGBCjG
wGT5Ursyeovf837b0JkiWfhYQn6deH/8AdtCUnr8aV3oGl5ue11puE1ooeuB99/FgPAjVEo87c4T
ftHWPvQBxmfQYdCwtvdtEr14g4t+xEQdft+Ca5lo9IXeDTKnKOmUMfN+HJwn84U5Z0tNwnFgTYU4
6dtkjWmyW12Q52bwjQQoOkrFdZfGFaFuwSvy95Usp4X4MqSEGqBNUpvHF67escWnsaAXr1pDZJvP
bTntraZ2OsEoywj1eDW5MD58cmUX/Y2WaRRdr1rldK+x3ihE7gs/aHoYoGK4a35S1c8ZQig0AGFE
E27NTj/DicxN8s1CoNRT1oWRQ73ifl0Czv+h3Z3A5ZFsp4KL1sosgGHwiAjayrJgPZn90I+S4UKS
3jyamqoQ2z4NA682aKq8QOfMq2KofhC9ebl/MQ3WRVoI0dCN5PMioksb4MuqoT09rzOw41ORPHWX
/NKDCOnS4GtcKxLyzFN1/pikp1W+/EeVEyjTaldcETtsUZgGQ4j7ih6EmJ/k27MMBHO4rnt1q32U
wehLN1VpdSKv9FyTM4a5AW+iuWmdlOUi5lIJMppzs4C4TIRcFv6V81ds88yG7coHST1XnEyKO61n
H3IP4bnDGGa9uw6hnAZfTyROaDqMzPnwLjt4Q3QEG8ia7gSvPegZqX/uxA5mphv9H1k21eQ2dMwD
OBr6RUwciEHHm/0wjSsc/wvAQYqOZATYK1oKRwVmSnWvyZaPv4Dc0wQOSZ8Aq4nnTNcFfuPz0XUc
FGwYMW0sYWP+E778KMGswK6YsjuR1NXaEx+TyBkkdPwSCSkS5MIGkbh/w9AxJH/6MmecKma7arAn
3ycKVSG7jkTrLko2aEb1hFFPkB8ftwGAX6Xtb2t+toD3bcMirrEWGETyBA50Lp+j7nT3TrarLb/A
X/JrAQvvzOGBzA8FLJp8PFRyre2AzxQYeGJj48K1omHun5Vk0KC2JtoUhdyGSOrZaVbo5PCiE3rK
OgLOR6DX5AliPXxpTm3N3CFBP+C4IItZwHdlatOvGD9nC9xtvgl4KDKYhD4glHEigmev13T7xOpx
naxwBGoKsqeTeJGY5jD1XWtMlFlptyVcOhRbd5+yirjXXNVc7Ixz71zMF+Ei/xG/5M3+/kKJiSha
LlcZMdxGBK2OGHnipbXnbuA9rHaQqEZCVscdUQ+Szx5yIkeXAwcOAm7oD3D9L9qBBYYLrLOH+rEo
LSdI3vj0B+OEJYBasBXARzm5RJwJ7Q5upKOembSW/0kGto6qBzSMEfGgjxYQo6dS9f9dYGbJGlzS
Cg7lzMrKIqmVslVCaYlF2Tb3ufBI35aqyx6ow2QMWsVrrNNohHL1P4fFnI1p6Hn6BS/J9Ntup5nq
etyQ2Zh6yvZ4y32MXuenE9X8YZ1Gh5qsieB0iMJiJslxbIVeMZaWRTI5NA/Z9cfaeUsjYG8rqIP4
UwcNLt1HXFPfq602JHD0YrVSed1p7W+Ct8BIOj2+Jjj/BfV+HOomBzBWHDo1n3Bf58YVm3VLlLto
WU4m2SNaF45corfuSE3BUGrG2ERCQb+M3LQaCjlEcZDEMHx70Ee+ehA++mUDp4ocDIQ0I/DhVWrZ
1Cr6OYswQiANWfkrixvc/sYF5y97DQvvTvJnVFIxsNVqwowR8YNRGyA8SVkONTtdon/SJXMVs3eL
iFanhH7k+nULoc/sUrGEKuMY5aBOqAh0JSwXN54DnNbUR0jrgNyHaRfO5qvBWTPpHJTZEwvP4tzi
MclKe/xUoDQbxDFFHCuM/LSsyXzL7/PfWLXxFqwWVGMJkxZtvNXS5TNKHCJugxWbYDrDCxlXG4F7
rxrWropBV9tcRcoi58wUKcLUFfeVrB2NdjiMkO0M8NrtnmaKuK3wllQeQERv18Pd3k/U9wIIVofA
4CO/DBHVNUGVal7dk+xA48Wzdje9ooBDwzdYntZhrGLNCXcuuLVqnxsh2V62gX8qPDkCLm309Dre
O5A6Xatpw6fqWvudN02TbDq4DhMjYp0rUp+d5oeGI9SKHK1BTk77hMmq2quoVWgZGEEDGlvMbGuw
cn9+B73KiqQ1ENAnqOwW6ZcZdVIvlRciAO56U69TDOI6Z4+8fbltQjhhWKO8E6/ew01tgmD7ICC9
HtMwEZAafUDduL4n4wo7eoUjr+OUBU7VjLyf4p3nLBHn1grOVAyuQnCqD7xL4RIuaynEelJHbRzF
MGRieZWcso02On7HZN1CeYCWoyAwIv464P0Ujah6IOPtRdBe4FKQEpB4z+QtJPs3P75ASqul3o0n
xUAwqt/WFdS0Xm8/VVpc+BGuDsRnGKC26I+90OZQeJ4rx4z1t8l4oZoZNDiUgnP4yU4ZolQhN8cm
+gGPoilPKZ1qW8DHRgXGvR4mtSurVJ43xPJrKhI6pK/esYk6x1CvsVlpgI5bMmF2hiHH1Q37Ob9g
d/2ovAJL3azOZ4PL11Slku79f6YNNYKEfGGbMwEgvqQ6jwgILfeMoqz01EgUHLKEXvvAYVlOm2X3
chpbwmsrPSzMA/3PR5GoMlvN53C1oKiqNKqrLLIX4qKMXlFTEC2WV1w99zJl1rSIxpAPU3yqsj0Q
HZYEcdxxVLwfY7Ofr8rl9qfhIUZsA2P27uUHXOouyjWEDfcb+Dxuqzhy6pVhjGzqP5gXr3A4Bk7d
591v1qJKYVykv6rXMYyW2xu3MAtfDbocD5SKhzvFD3f4h1puO99Kp8gW8y1zJpuUtJ015HUw+wNo
71qvgyEhaQa1XxH80LEfLrzowV/o4z2u1ugKFp7yflaFyYDxdu9orNq1G27hXZAMB3XBON+FSs3p
3ecZNZdI/0qRHS9QPeIw801ucdihwQwkA0I7khGmTZ2tRAQ7ZV8xBc7HwQJXK2VjQLynYsXaGxyL
VtYknOMLRlh27gBwU0qTnNe1MiFoUDLEpN6OxZWdHuFtIqAPVHlJVuphrL6qyDH+f/xyPkq5HOcX
esEpHtFjSrB+rnRGWfiHvBaW4qc5iwztIs6UsonKxflPqUiENswLo8RM2aGhlQZCOTLXPCctXniO
6RRKbQyefICh0oe0G5NON7T5T7YiY3dD4BPiJu3rxxAb90NzwfGUdRPYl7TgtNn7zaIMJujEpHnD
CvTFRBJ55prfGiHp1cvVvbYcHMi4v5HbdzKojo/5Pb2yxnl4iQs3JXeRjMwi9vlQ97b571eqfEHb
qkhUrP2LnLJpjjYj7XZYtbFOBL9n/SfEPm5MfOB84IlU8kI6J+zqNcHeG2jKznVf+mXYJhC/eZh/
NDQQCVfBuSxQ06N6lGbyBNAE71odeQzL+5gF9d/zIQr9mcb8SScX6ZLmTgO5SQaRaUO9Gmm9ZlQX
uovBHROUiVLMjOt1pE6mAUKwNKF/WWaO/vl8QDsMr4cUrb776Jw5TZi1jEbjDtP4jekdsuC+YZWq
dA9iBG0jAyv2wxxfjLZHzdE03IgHewu+8/zie6ti4SHkGFR7LfrZKq5ivsRx6uYXsnEh9iJ9HtHk
lZUNsBt28EhyjvQxWR1R+7A9CsljuHnvZPk6HFpLS1+dmSJShTaynvvHxukusPZ68gxEW8NugKtl
o3JpbbdJ5R9mYTItw0LrkT+jBujoRnWf66qyOJxTPG5iQ72ccp7JzLg41oJaUiuu7CL7E9zQlN1c
pTUs4KGGKhpXn/Y/bjQQnhICkamefyFfX5HdXNtkJ9PQ7ly/lGJNyEkhnslAcxLUOwyA629/kMaN
xO+LTJnyViZOBl3ce56Rqdvga59yJ5O3+G+Doi2DGAO3pkIfeQoUClpmW13im70LTHeVycK2NxnJ
NN5wWbXmcES9tzBi1P7BYr9j+RuMa4iyTXCCUncIWnEhiTKRnTfIS8ORBT9wXVLGVISTm7L0DITr
4Gln0z5dTj22PKUoBPIY20kp+wEk9gHhvRjrLfD13GXVhpvbV88ZRjUz1F60qfiR2dVR+CucSHzO
liSEwgq7W2QUWX6qtSMtkkUJV90upUpMxeCFKPH9p6bMmNZiTXgpB4HV4sTH75nW5eqwm6lYgmqW
2pXuYcKVQWDniqB87jb2vEj+L4KqRmcLjkez8agskomDcBdo61DpBg7eBW3uTV4xmqQvtd71TTc8
rB6SrtucxpJWhwQEFK/0D656nlq3Su6qB3UVqrwxipQ6BYWbHOsnOHzOzulNTJm9JM4cGXkT+TvZ
rpuEpyFp29H4/BiGFzPP2JZ8pRCfN0+pY+daEd1ML88gpMe88n6zD+GT30TyAFHSRbC7DQdix7Bq
f/olsbiuDd2ysaDjxhDgFCU37xE5ZcClFUyA3p+QzovSqT1Ab7NwNf+O7OWBbPe3yiuTUj6lKN8d
9ZsNPSyaASfInBuwEScsnw2Y0mH9dRHu5zgKDa/dTDv+A0UirkQn6hXB5U4RxgirGTIjBU2hQVpK
jzlsbksPNbWa5wtDOMPKZ6tRviu1vosn0Hj0gVWp1oYLARfbZFGhU0fHWd4bct3dVW3F/l2i5dXc
cq5d0IoKnBDqFHHObwpxxyefXXncYxCAGsBu6nI/xKWlQba+A9MC+9aQwX6xF1+LhTLS1jQoZpOj
WEK/FKUiYZbEOwxgpdeUMn47bFscfG3BYTb7a4gLp6FrkT7RukiZVjfLZLjSK4MUZuOVjziST7YC
4TCoEYBtk4XznhxhSADgQl/VIrBFKAFUyZ7KoWXcWv92E6yR9th4oVwvasaJ9afKxghRXHkd6SF3
UfoVB3ese0Qm0hKqoaeCC7d/rVcXOf4va8bEIx01gl0JkYU7Bed38vqGKV2ehpM4XXNOlOAaYley
h2h4OzZlZGwK6uDXPoVWlDm+gNENmsuQChylcy1B1wrhjlyRy8DLY6u9n8VIMzbhtoaWPs7pCABD
VXdGQd/E4c+Zem61qPRoa4Hx41R558G+iff7i7A3dAEuuNf1DDSG5TOr29Fjv5TyueUw8xmAy+nO
a/AnbfmAWFTrCAzvTsoYMrB6IaW8Ai16NP6VFDPpPOqxIyri8AEoxwQvhgmFRV1e8+81jl5/dN1w
PmzYvGLxlNucqOuTUPYiGhwmybWshWTWNK7+QzeXHRPnbf/buZHCXrJtJnastjdVXWnhAIgAFqpp
U/cAUb/dvX1w8LprvkziX9unJAOzl2b4jTcRuY3ARPSbp5nsakIfyt4l0JATijJ38tz4tBRSwrXA
VVFR9kXaH47TN8u/IMNUg0yocPrb5gIc9jBU+57d+gALxp7HJCdk69H3/W5FYttBnHELICZsPEzt
oA593yjrsS05YsEzDQY4Pqlki0VgR8mJuBaIuljoj4ks5jC173Bh7hA7j2aHQjxIGXGGgF1tlSuE
9QKoXvP94dwATCJGxmpFYFY2fFN02CM8dgz9VTojugGe5vJc2P+QnOqmZKQ3EqA8K66sBNZS0UVy
97FfZKkjUSfY27gSnrHXjTcxQUD0cs+0t6UMlzKztkehf7yhjDtVawlL2vP3LmpnrxcEW6gq61XR
1KH87QmGbThQwuMneH81nXqBc57tyz9k6XcAmIMfSQ8VEDsMKZkyiR6AnMsjSRDtqYknz6Qs2uQK
N0SG0cJMwy7gRAKfaEsLnCQoM2B9vKnqmqCzsPHJM5RtNFbUJ0QxQ0aaBAB/19yV9v6Gsn9fUgRI
gjfW8MX/zik4j7jS4K4LeLOU56VeihalZHtEVycuKPJXM9um9RX1Q/4NG1E/6w9P9hFDnjnlnfgr
PxCDXDDx5lI5wQAygvYZBItzqSIge8AJI+iAjLYVuYF+rO2U3+4YLDajQs0/ac7iFHeHs+6B1ene
vz6b8nzAdt13B3Y3zwQAl/bfPnCiZyGzCy4ZDM9uXpv3Keqcel+TIlVMr4fLDdz61NlXTbTgrVoN
INXhEjIv3g+H58rpdZ8dgaCthFcT+dPmwtqeYG16ZXjFSEeY8QsG7+DJW6i/OFriyCB7bmDEuAoP
GcokVLCxs8HjOwduA3svB34FlgbDunAaPpFrN3Z1KZqlfvYHnW1O1S80U/bt+ECVi89bTUTa1KZe
1A888na3fcSqSkYc/4ZvSagq2FK/9mpKuA5g/gGT/GlnHDIOnN8uhs5PH0apPwgfsUSpExkCrhSw
5yghQErhUrenddLZROI8sJ7XNvzuLLlhiOA7lsShTDFV0d0bam8J1s3BK5834cEPdPxAamlLgttp
bSGwCLuTlK9ui2IJn6ewgFFbrjY+5pYj27aRbgyFF1IrWXzbXYo/mUzd3YVzPus15oZPJlFB/5mv
khGIemVlExTYXibClMUzlPbx0/xj256Y4s6f4zxsKy3Ar6UBOs++WHJQgLiQE6dVGnFoiIS2tcQ/
HoTzvnSAvxNFN+fGaycVsNWxnTKtXhbBboO9k6qKaSx6Otn1xPazoLAtmg6sz8G0wom/VA7JYWZ7
grewWskEUVCP3XAJ9xwwETxOgcog77GaXzhS52QQsdFp6LwB+PbKBoTZwjO8MUEcthPr9KQjYvhr
feQlXmEOKCQKAbescPHAXCHFqOpPB6WKlywg8D0egXG6OL2NDIHd9Ovi+iw13Aeu/99uFTa3xRID
dZ9RnXNr5rre2Fe1kLa14Hztgg6QRhCaYG13Rwc2ju/qqrPjrRd2n632sXuDItYBxt6pSw5Y6du0
fufDLmnN0GNs9xqt/Yf+2RKGaSV48c/Mxqe5lUH0xQOYnvIUw65s0A676ctkuJ06G/Qr57SXu9II
zd+jdmMFGbuZsIYHxeNH4ld3AbG4ztVsH37p+tlq0wr1Q8dK7LhT/Jey0kBHV8CzeiEEu5+TSEu6
RzLw3/Sh0msZnKz8WkpgVLpFkR5DgXPyqDzwaH0uSWsjWHKQB5YJUszVVBWuToCKlCd0lieRFaOB
yxscwR2X6kt/4HJu/rJLSSMlDjRCcjdF5FzUmjVEq4Pw2E0s0+HIs/1BLfmbslXVAfEV8EMNCbut
0fop9W+BNaw2rGrEQIU4/4tkZzM14amhAVtaAtZej/deGXskmnpsS346fQ5zzxUVfMMJsMGqWBMd
dzlaI57GaLupmW2yjSMEPlgYRdHJ1MzSz/C3JxrRz6VqOV6juGk32v6NRdNoYLd8cNMcJXQd+mv/
+2kA6uLNlzcHVsReFjDRoUn++UmzwKOhkK/qmqv0hFJEaA8AP5N51vZHpNiOLs71OLM6H24TW5Fk
S+FV4qNWw2OmVKiSJCsmjSWydHYduTcFSRT6v/ltnPgIOxck4egSs9QNLlmM5EMTvVm9kyBLjFXH
V9pxd3aEMs9TcQfRtIuUmZjtWngyErKiuvAL3xoA2vOXxPUL2CP1Coa/VT+uorlg7+9swxXeanKs
Ny8k170nOtKhitHDD9Fm5V/n/65qpDcrxKIpvWy3EWv6Nr+1MY+VzGcQOsp51heO6zr5P938RMlJ
1adr8bO02lcOCGQfPsGIcIJOxj2OFzVKYAQzLZEvadh6bmWhvqncCG+O9P/f6jNRfpLdHHAfodEv
ErNN0p3ARQUlCdWvrhxK+jdl8X29t8/rAaIEeOV8bDnddCIHHtnsPFeT9rebNRlwzGoCo9PAziD0
cNFK7VG7JO/SRDLM3a7mj/ZCsWf9JM/V/ZW+XPHUeDwmYxSUpf3eVId8JMSrJ+eutaevDvDNPuG4
Pt5WnDSmnopxuAW+Tzhf7v+kKbLfsi0WQ/vXRvzWf7ymMwhzdmFJEKYjOX6ZgC/a1f0xrQHx5lXy
Za8gez61T+6EWfHJa9KBrEq52j26QU6lTwz45a/175ixkU3NEdDgmKKnm+l7zOMA/GmICGOTSCKk
d9+V0/g7s/Zf3d0THyPP4Op0J5NYfm4sbh6ceBKgpMGSBYiDna1mNWqMt3B2r94745SSCE1b5VJj
kw1A4LP1S1UWd4YsMIqGYHPcVEEOr60UNEIWprMN5BjEFLS4PQQLxgIfMmYo+qWmE/Q/zmcXjvl4
0GinIm0Lx1PwDuNBJlx563cIwu9IznmQagAAoILzx/8c24P9QYXzehBnsp2DmQjSculvK/0yzVNt
O4xoeIrCUqv760fJTHmzxviMDGl1w4PikzqHYZEoUqj3u9N/W9d4WJA0IfEtXHAGweF51HkcD+5q
J7/1lMB80wuEmmPHwH5m3q4N4Pa+D9M/eKGqlrkTgzRHH3UntqO+K1Ut0xDfHL1D/e+I3XeQP89x
ygNLq+AZLITm5Sgs7Voa5Rsbghlt272Yraz/U6u1lkf1X8UPBK/kl/7BEp1kRcF73trGyJtlMJvh
PCzVN7JkE3if+2/8Uvr0FXXGW+6DRHiTPxsI3k4pL7aTU9usSGVijV8RL63xBZIj30qF0onLY62K
Y5vrhN1ZktH/eGo+qv65RyIEm+YHKV6fiGcPWu4JXCKXwV8IGWchOrCyXKAbGCdgaZjJZYn71sgP
eCqfP+l7JPCg5uu0ArevVeU4uwWrxkjJHhYxxqe6QkjnJLEp1EY7tn3tFXQhHt1jP25SLo1LSWhR
YjHr0G23fsWcsrGLmcuNZeBhqX5rL7q/NQlcdCd1NUsHDyat0/yslRk6dbkPKVe5h6ioeZECxdoh
DnxT6C+akBs6Hsz0L2VlN+FJlCCNp3FI68PlknvvaBE67+MbXsvDQg8ul14jYkfvt1UKg5zp/rt6
Tx9kqFTNCvsAy/bBNMgX8NLOVSVxSIe7HvI6toTmc9ztLKFyh2mLK7HT9Q/fgTurjh6HmC/pfz4l
yVFSs44BUYm9ytIhEwgkJfk3PvBqpedSav8WFMfizzMSSJf4EkXUqBmAJ4Jv8GIUANH8Js5fcZTW
jtivjbxr7qN/+UKKlxIS6TzBw0cRZOQVfDheX2bbXwG2wcgR4NFdUbaR7c5qhfffCO3plDMrmzTc
xwBtiHxUcLV2eiLEP8hnpbpQybgN3M1hAzTJZgrzr1AgAaxXu6AO+MTplc5YyVgzR00K9uyRBFtx
qalXKiwD+ReMQEUMWxhQYxkguIMPZCN3A5UN1tpxRnWl79GJexssRTX+hxZvvp1RZ6jOWe4jhZNt
u+NVX1b6VZR5Zz1U+FRdZJC8KAbt/FLKCspAPIVrBcWbpvzI6+YSC1dA6MHU31QKCi6ZScG9td8s
1qUHlfNK42tQ4NXnBHRCWb7b6aa237cg1tfY7pxbB448srW0btg7W7DDuSzD1OFzH7ZF0P7jHuay
J2ZTcERDrNTBv9lpDkNyQblRBJQV/ZdItOAj9lW8S+QyqsZtPeHNYQD7j9pvsg5BLMijX4YzRFN7
sAKUh8b3fwZwbMEqfaS69PHx+SmnScHC/0QfhdIaVrDsxUr+RKKR5YEeaAXIX6lBnnMKtciWR+4K
YbLaM77Bu7wJDg0PVVCOhBHiViXErxjjCTrpnphyj+aVogmZ4mL7Xa6HZZBSr0XvaCwhkiaJYbqX
ZjZlk1Q7HhpuFzbOdeRl5JnTZLd9wbZKGHHSPayc5O9gDz1JFZVQchbEXH7weL99bcBKVBpIzNzf
BWZJUvRsm0SlauzKvtVTwk7caImtgfRVukHvdHUVFreaR1XuNDiieYN9l+HHGKRk0Ur8noCfd/4j
dX3GxWjXSraVfl9FJL46chYu9bAPC5EK6D643l5djoUFQBkw7Mwf/ffMz66U/vgZWe2LlG6GitSb
YL1r5iro4P7fC2W7VPc6uSLlIPou8D2soQx8gOdJHsYDIT9ngZd6C+FvjWuE0EcHif++llj33rfg
/Vaz855swsUq6XEZzdsZ7yN5P6O0LXcNWf76XcZUrdUkUZ6EFNY1MgF7ro+HmaIufKQVM9jUpDkl
+rpMkKlSykX7EQakGIIQy9gTP/H7aMm5rcDwZSihTGqRBXKqMFa3+uRCdXowvFEHF7Ulxg+kw04Z
F/uByY2wx1J6biuq5fMa/T21miNMhTgCtoQ/w7ooHWMZ+Hjp6XMawMGMtr3X6wwSdiEvWv5c4T12
BFsvmiYQlgWBFwj9I646K24RIX0ljno3z7xJQ9bOmQ0hNYhjmmUMtFcg9JE1XcoaYvMPemY/T5PV
SIflsjWw4ySos4PDklzYGNalTFOMYMe2mziDCsgSG6Ji+oCzpMyAyUKNl+5k3FZWL/ZSghVxMZfk
gYkz8xsar/cAuXiULPdqAKxgssdKBUmOv3VKObCh3CNuMKNfzJNaOnssTR5imeFdue7gQrybB9L/
0wrQb1gavAorUB46/0DnziA9a0BxKSZpAzWTA0dNFLvMq+m8wlqPIBqMZniXmVKv8MM+6Im6Vk6h
ML4q4zEVnXebiQXHuuip7ZxjXynCb9hu1NbJQJ/t4mpJ8QC06QxGu+y6ehXi5pWteYBkDpIfGorS
/o+/M97JyD99+N9aaFoWsp3azxQApN3xeJ/3horfaXmMW8Refxkrfn9Ldf5ozxvKhySoKjNYOZQs
/M+XJbwjtdPn0XdjKL/a2+8fyUMjibeHQNMUlu6ySzztKJOc8HU6t3sxh4o5IZdl69VhkCpHuWpl
pjfFbe5xr7kGyyx1TRJiMRemmBYQ44dno8QEbdweimd5HaSdyXEtlGHAtw3uSxW/eTkuELmoQF1/
59qoc9hk86kqfJsSVMbzaX7IADxiyhlX9m2jTk/AZaUSR5pb+gUgMiTtyabzqwPr4AcwK6sZya6e
vNUYLMkZn4VTEacOVWBZtllK+MPc6gMalBWbA26xsDoAJG5pGubAejm9Kj76aSz+7TFTj5CHvP6I
oLMuz9plhxoEKU4/4BjFx5ffEt5XE17nku2g/ldBZRtZBavuN+Iso3M1vAKMaxUOxOjJ+aHp7053
5dRjavY2ZEFluJ5sn3LIhLG74tBFDNk8aFK9rkdi2xJz42vtRL1zQHopAp5QARw78ZYTTgH3CKkW
fP59n8Ta6XDoOTKbFGrjdfC5c+2K3EmYR7hdHbAr4OeNJKoZJGDr8RMFQCBNlUl/aJgJuz5pizYO
Qa/ZmF1vrpLo6OokhapYtrE9/vmAKMxC1ItwgK43ZxbgU4bhtMHDm+Pg4eI62PJyeyPWSrBU+9of
PPwQoNpM/bChMKT0PyOvUYFznPKrfIHFgmWafvnfXlDNu4fmdISuXSQ8fZT1tQtPv2NYAzsLlQ1D
nLfcVfUFUm80mcgf5zcZXHKin+HMjLPlvp5i5WOTgJ7PGE25hE6Mj8Yae6AyZhSjN4wY0C9AKub4
fhnC8otC4Gfe8eTzjitu2XsU8tF4zYpLsRd1qa6cOuKkwdOLFa9fzYIN4Hxo0yCrMSSlLeg3fDpC
4ts0mWoR8buNF6dxGw9d6iiTZtivh63vqJWwUJdAfyto6h/0Y8v8JQivbmu7SFBlA/i9gyYjjTuK
71G5a9slkJ+1becgW/Ly0K/twpThmXJCz55XdiSfPz7QaFrSNXZBiNdKfnU1Ikk+XRjLyHpCAxwa
7RtO9aVNdndavbK8ooaBxyw9Nb7HJ7rDN9q+lOLM2eEMJyKmdIYL8AmIZLovfoTFYyDWKxU2CtAr
QZUOhADpFLAoEjtt8NROo5bBnVI/byPT9/w+gJTbwhmq7ES39Mz8F8Gjh+zTN58qYFE8P8Q3kil3
Ds+3w2YDsqo2xPLIj10W9bPgIejgQsvsiWNDIwKZQ5QOzVWWZ0ueehRxhk174xouqlDq1U67palc
DdI4Do8yP/rRq8mD50GbcQfGSQIInyy5hNwtJaGy+IpKZF+6m/Jv7+dXsoP5d2fQaZDJ//dPH2nf
6vn/PEXx/kk7WcOmXIK30pp2NKhN58fiRFEOSqqkF7OZjs1+V+ePBHK4/LJez/iZ30cz43X7znlM
YFgpbBhTnvRMXWWUnIjOmiAVQQM7EwkSOA/OKq5BAxl7My49VrQu2OCU3B253I2yChmK+43KKSuA
JxjNVClNE1KtHx+GkZScqNmuTYD/yxr3eJpUZc9tRzNWY6AAWADS/cvzDKEnUshvvKS/PBVWvNqd
bQa/QsXXak/11lCJ5ot7vC6A9MP3AJomRiD1TV46e5btQ53nB18amj/LGDwpI+4sgdAU86xa0AXi
WYK6PA4Bq08s5+48gneM+j4ZpLIgethfWTCnesaqcL/y3apvm5Iqs1Vd9TbEB7+uAcUczV+C+vdC
6Tq0I4pKsqXaF7uAC4arXFH4mQ1GAANdfpHZZpLrRoApcGk57hDCGeKziTyV+XeA24Kl/n6RE1SG
hcAeMuN0wVXbAzdOdCrPC5dWbDYQGbITdosbB9HTGHv0PKMA5MUkmfc9So9R0Klb7BKoVeFZyFJX
ziC+7ue5jWtrM6TpUhINGg7aE7YpGVfppvWqi9s1sGtuRLqd4XcTG9YirD8Z11YOSptiGmkH46Nt
rj/6rlnvXZRUudZF7ldltdKC6W+NbxUEApB/HMy6+dSEg9g0N+Mb5DTd1q+SzWU7v7LeG3mvi+48
aKtxn0jbWzlofxn6Y0SF48V1kx0Guma8oTBDVDUIKIAUODsuJR/Nsz3LsYEECX8HcgleR+1RGyDa
+nQSWNurtkJ/Mh1r9vfadO4wKZ4MRsfp36Ad7wwt1x4Kexc6h64UPWyjC7AagDQnM3DxrLa9OKW+
BeLo8trT5NOzXQfLxe1AxEdkm8DxdAy0UL0HHdG/O7Ed72LYnIHigarmhtBcOGDvG0/+xIdXfqka
wu6+4qEsBffr5pGK/uOGq5I3jikhEBkjnL7m0yrdyhdECHx+NFaF8LnD2o+kmfadbc+5qSHiGnnt
zQqUpTHubnEhIqJVemkRhDZy7tzAxTJ77XFxL/IC3bxCvOtVLcWuy7uutw+Ij3pvGZEhiL8mxHV5
ApAtUC1wr0qROCsmLtQO4AYShfxjfDJSGS2wxWKrsSwF+9s7Js0+arR366rWZS6tiUn4PR9ZCIpS
m2BgIjWK5czdvJZu7XFu6FQdQaZnyiOEx1/P2CK+a2jyOxlxbVdZxgPPbRkoNvqtMxgXMY1E8NMl
xhyeajdzGEz9pwCOp6owF0qMEfBbIv/4hqs3+gam7uDX+5XhTPh/LawbPV8oA7cyXjsYDrpTSwnq
aHcutAjMuKh83fPBPgR2WYtsdJLwyGpjM6dhtFmV2erL4Qov29EDQsJYZMF9IbaAL3oAGfuvGdAA
nOZ4l7ZCoC7UAPHuKWjhFB6iuvIhsLl75hCOEkt+ArWpuHbn7yyrCT9sJNImhD8187QRCeRJB2/V
Lhf+eesovUKfNjYNeZDp9QU+/tS6qbyacPBlwtfwJWmYsIw99i3koa2g6ylRTyiYFXuj+aPsZUvI
RAgd4KGf1GpBv6EmknRggJM2hvmLhT99+ry53VeFmNm1GEUAowFGzgJxEWEjUAq9QTCCxBan8pao
nvpjcFSf4LAmTHUuppydSSPjqD84uNzfbicziY0uuBtq+7V8zN/pHR5RklPL7lHeBGaNeuFvINM9
bttaSTK7o2kcxQDNkUeW5JszPJBQ0knW6zeZOXIcqXzVokT36hVLa/k9xhHc0wayzH8uH5Yi6zbu
6ZKk3HosT6qKuN39QMRc8mCtNsNlgCTWcPZSwURIda5GQQcT/+wjw0oUmtD9fD04fRTa/QykuYLe
mCKIUE4gyvls5l4Dw9kv3zjRjRWRi2S5/lPftXyUm+M1EdembWBLwKRxhhYzcBY4TnXJFSnYq4fW
z5Q/O2/kOuz1KzVjdDO0Pnp+mclyeFNk2BMTd10GtHccREA9ScbC6JNwfH2R1f+ivfUXLAk+qgOf
jDPQJN0AQxkl4ejp+ZES+toLjOLVLrqGduVGiUaMMimecUyZ5Ho1dWjf6kOkkg6At/zdv5S4oJL1
Ubxr7TKv4KODlCSL2WYcnrY5RNncW5eR/yydvYVQvEbYogHdrO1To8PHHNvhlk+lpAheQxxM3jOF
/PKrvTGKpAPlS8ocZ3KLNjp/kPvY9kBvjrxxbhkJtP/hEnIQRfIruRlKKS1K4MxxFIJyBa+iqiHW
MbUX8AcNqCVaN7wD4HnDV0SpuRpznozOF221lzmDZUXQT4pJi3GjS5roEofptq1MPbn4LFVcQZYk
VrdIYTOpnDGl0nMk98CPBlLdKR6zN0TJ8xcJ/5MuD47VpGTsulYOj4zmzVt78xwcED2gzygV9f/s
jLEdgjZMYIBb7E/nMhpVvXlvQUvBojT6/KR7DMYg5GS7gF4UQHLYBuDH+yKjDIZYD9pJ3OgoJLK1
gPk5x4FUNVS3XMpbQmBQp62S8bTUiHRdV1Tskog22U99Cnll7XOqg9o5ZFlSAT8oV6WCz4imVOCr
U2ANJWwBRl2IKw9n2uu9S7wDdkqK4iOvK0L6bk6QVStmltEg6evH0QpzMTXBatrM/gvOwSZm7Ok6
jmCPHfV49+9LMMeSyrGUhGBhIcQXvsZokKj9lv6guajlmoqQHsTqUu+XZkmlrdSpZDnfVYPOreGH
/M3uVYixYfML+mfZK8pTjUyQpng+cA4yYsDbPpKfiqyTReIC1ydyPvWfO1xAhFRXm5ebe8UNcaX4
8ode87LTas69NJRYYSD1FS+C2buU3CW8S3JyW+xx2917OcS8QIaDpmhXT39CsX65J3oJRda1Dk+4
LRx9TiDiFXqcBTLYOifGOY0cLXZpNuHxWrLlwqUXXmU06ngpNWpuFT7i6z0AkKXjFpFC894LZyGN
wL40PwYATkRooZl2fQJBPZbRV366+WxfllJTu9k0BkM40SmSvzNn/o+OyATm0codA/g9efH66+mk
6LuS7Q4vYCl97MkpBnn8XApupAYx2VZL5m4Gk8xYiKCRvkXZ/BQHUdC18B/wURcmmC8jfTQyMBuw
0isatXwCM3wqHnHrwn9uG9V4GzudaKH+GNaAfWCv3S7AuD4lK4uu3F6HSMOyjPg1xliqs7D0cYeb
YRzycZZKK1mRq+hqZt6qPoFaKHxws5nm4q6dult3IyKLTP8L0r+mEMmwhV8MMTXeS6b247azluRv
WM515dVyIxfG+gZuG53RwuWlbpdsdsFzGWpYlBh/RjmpTQ61TuOCfBK3HDU2r+c9F0lQg8VX87y1
OLZ0yGR2w4gF8PmDA5wUqaE3HnaOmFoyYJ3zmrsed+ncgfr93s8pyYXCQmZMIuoWO/D8OFZQD21y
8mq2i9jgQ+o0uMjvRCdzIhqooN20p3okgf4U1VdVqDH/dMVqf+X/JsjkvAOStV5oPzIW26WVxnyn
R4Ub/1OrONQR0igGqWx9h979+h1EbYaxCfArEzvcEkXGyaOixTDaeRvrxrcSrDrIip4LYltQ4k+Z
1hpbMfzHv93TyX2AWuohinNaEr2cRZ6mWUc0qvWZMhoPynZHqyBiALhRQ//t+93C2VVXNiGGNmg5
zU6EX9dKYtnu5O/fdPMcjFX195DBCdjYPJfjyAbvHoLpy8JmFFQn6fl3nHWJzI4lHOW2PS/FO5lc
X8S4LBMU7C6AAJZuCB3CkXFUyoHMthCLBhgr+lCxFBOvB0v1HEiBOoHTHjRt3Ah1kBsWin/F20Fm
IkfAo/BMvKcKdNC4oF34i9LxBRosyXCz5UhJcrWLbsZOJE5irZgOyeu8ElBztlDsi5SUoOZnmBMV
AfUsMPE2SJVk1Lv/lLnIoK/nFE4ObmQigF6CiS6daYBMRUmESyWaddCCtKjGLJ0fEKdslAwSYxIS
vvqt0HrZC8EcbJIEBoGr/K1ei0KTnetjTO/ETxByX0l7b7RRTzoYP0nwRb5hl2mIZ+h9OqFVDv58
c1dMC1aq+nOQCjzCGqhi6Yok35rH77JxqAukhdybyWMPW8fmaoYAWJTFlX5oACi3LuvVje3mg96V
wQ0XtxhbbunU4z1mcji9g/a8m9h1xZMPJAePvEl0Hgccz3LuzhlqpvHnJBITBkbUT8h5PKKYuQEa
B9Udm0FnIf0E4nVN4h5j+LKyTEGfPD/pZCOB5qEV1+KPwP4LO/vdTmFHsan7qUfFO5bY+u64HZi3
+BvsWzgMD+0k2xW/RW2CjHrqU7L9RvKz06bFZFkfwr0ZhfQ2A9EKdsLkuBduR5mkh24kATjYAL4c
zWZetG3D3kZ9OK7WfN14gfBAIClj0mr8T8OHo2IkHF+sVl2BpgjUXGTSUv4NEYCWbM2gntPwcALc
3Kz092fxa9G3vdfHsOmNvLFwTx401j9WePb9fWRKjGOE0HwiyKl8yPCUXkufZ9lR0izzsKWiMh8a
TYvqIxN0zmu59l9KDWiJMii5lPuuxnWqWyGGu3+X60+AR+rLYVxTXHE1JlCjV28o2ldnY5Kh/GvQ
YRh08nphviqtKRIaaDtMtaDix3WQLzL1NA217xjh1fH9KmODhX7PGKP49L4atakTeXh0Lz89Uktj
At+8p3cyv7srHLC6Fz2r0Wa7ao7mi8QT5nWaD+NwbLTEcSS6icmjdFArLvU4TJw3Gw3vme/2iNOI
8VOME6++glXcageFKSZ8BkaRhY4GGEl6pEqk7zAS4lmiTI2UiJVayNvt9SdBzqyQHwPtx69SFzWR
GfkXRdOPxtCnTr1h6GarXoS5yTr9wFQDYK++GAihQL8Ok5lOXKYedoCGEbZ6mxrKYXQFFRVDpgxU
jPN8TCHCdVjBVbZeckIVXtKO3CxEwv3sqExWKrTTGwPucB+V2sxXjVS13NOgOvzVXitcE5qAtQP7
j9GcNjcqMDZ4f6bufSl2hMplHAE/JALpq54yz6/n1Y0xCafqLPSJDbftDHhNKqci3VoE2ymfWfsN
+EXhwYoNBTqiGVz+dDuLg45QRZ5uPCt5Ed0Rqp13qNZtF4k0QjFkprMPzNNcAuwnXZADjKhZDMUl
gCODeecKS2737OOo4pKvepHZ/gdDeCJ7VDYWr1Gg1lPjlY1nh/jSGD2ZCFymRm0VlJSCcllmoqhM
HDadkvlPd94RJIZra5rolwvsaq5Jju/SIfbRvYZ356D3l3NBkiFT5fez/fFcSIVpPiDa41HqSLcB
XgZJwHuQ2YvIp2kufMvcKhPVdTkJE9iQ5+MHcDHySDOzxd17TWlRHbspkd4obWtAEySKRKvK7vDM
2uJttpNmdnnYAIg872vHmxeQ7P4w8+E5oWR5TVXolateSfUMWDZv3wYl9sY1hD0HKMl5RCeoE4Tn
I0o4vdJnYyHXNshDCLWdqugzJV+OJzLdZg6ikQtb9tIHvqGPvWoyRjDaF+F8UOU3dJFU7qJGLu9P
s33MuMOQDh3gk2m+b7RGJ9uKgtH05bv/AsTyE4hRw5b0OebarAtNCUx7ssctAS8c79bZ8I6HKJyq
e1CvpKiOorlxGKBoKwjAhgJdDgOc0rpHQ8+vYxbdlsVw7pqJ0OnuqPiQclNgCoa5HKOU7eBttYQI
XoIJ/ffwW2sZcs3ilIZ7Q/A4Qy0CR7D54G+kvPlODBxBUU/UJ65JnESpF3bqbQAKnrrdWeRNWS8N
fFdZOEZGPy3ssxsoqo+F82EUcYygqynROkOiTAhIOEhT1a6zEJMrB1LZLG6F/7Y9flC+RngJoGGs
nHHzsuxyuFqgweiQopOSqdaKB7J1mxn47OeQInNbkiOoMkjk6l2L+/cdRbx1uiUguck+uygsA1CV
mAhwNX7im9AKEC48OkMx6PgNcQkpOdA6aTV8QG27yReYaFJIiFgwHqfzCPmyL76x2MAm3FYUHPWV
4/ZsEvUrzTdUxshbaVAXOKVRxxRvpSEI5SIYt41MGGaAvqcQYSUHnCymkAX38TaN0U2n1G/5feGP
aGpOlyJbc7aReM84wQWQ6LYA0ii/0xH+zAmQV0qC26Ao9q2sKF0MerdCJWZ9B+h/0NNJ0u7AZDvj
kWBLFsAi+yJB9l3qDIQrwBflipU3cCFCIC4zAPNgy+djn8xTHnXHJKMeGoOzM5wJOXm/vZH3wE4J
w3T9RDGPs2WZBiVrpiCmz4/Xv6I/3/yHhbzbZacMuk4jAm7jAht6jtRca/CVlrcQ5f1jMSkkyWTI
SKJD4jpmPgVQyn8XOPFZJqB2WavS20FMRTHuVVMmaArboztzb9CCYEBx75h0cQFuEd8UfuNL1ysD
Oy229OmRqX3VJDlQNlSlNL5MZNFrTqU7eyonrmTMOlCSOKcJbWnn6h+MYpHUCvXvFhhtiqUEkILZ
6W8boe7SIjWL66jyXIJL8qwRG4zYpr3IuAAvemWCxdI3rGPO/Zy6sw0s1Oyi0uSicWp+ubs/yCP3
9sUcOjKS5NOVSEyKolQK4AGXPigo2pfpEHy0AcuDEzn7a9nrdSeYp7KnSw/pkKKj8D8szhWuR8mH
EXHTzMEAhah9P08dZQoH/LsgavNgsxYD86UuKKRqsAA8lkezTsW4BDMhwY9LH9ozYFzUmqgfpX10
DCX2lFNkUFLA/R3jm6+YzOHVqqm3o4xpbjmetVKlHjtTInrEVWVajVNrRqSLC9Z9bTWdBSjS1JmY
ACoKB+J/yjwH8vvDqoUk9bYYGmN+05FSbHS4ozXin2jkOnhlE3TUTtpIE1ZmA4poBuRYAOBMG/Us
zvhLop1zYCBnqwECTxnx6lh+qqM/nFbizo8uVqo80HZGg1e9HnLlC88Rq/bn2VbUYXxRddrYNbPR
Yn2Q+Ffrx84zBB37G7wyvtsrgiyENH8dOZq/IdJrO7idwhETaoCb/Roh8fn2Q4B3jZzuwc0s6y4V
f0zmkEyXfnAFGf33TQwJ/MRraBJgi7ZQspDtQnCEmWp2KG1rxNpYLREMxtLPDJZA0dP2vJQH16Ft
HKtT0rWN3NpprzJ6JkWcBVpqk4Xv71oFlAWHNawgJS+Qo0gqLpJaUlAHwnLF2BGN/hi4ZBclYrvL
t1zoILL8ZmQF2DjdcMNDwBJdjYXcyPLIi1TZQewcxqSEj7ONml/6toL5JODQ7V6yEP48uYQETw39
96D8d8lICKBqVF+02Obj3HVqemYScfQ6NClESnpz/oOjM24GuI4EnrGTt1rR6XPSgvsfVgduNPUV
8EWEf9ANstJiaRr1yqodPYtl4fpiof/ZojpJVx8YmjxJN041mCk2pjRU1zd0W0l0ocotlIpk273l
UYWQllKHdivOmrQwQ43yYsO/JNaDIVXMiGCj11Y1gbJCkDHQk3U1mqOzJWLfWPbDaoutijFxo97a
UAW49sdP0JLfszc7veelVB8SspYbybSzK7XoypXP4I36aYVp4PX5Wcmoq0JaG7UU2rdGX9Vbez1S
ef6Kp3pCUtmA8FZ1xNkMjchVTxqq5mhhkAsZUbavbcSYyfC8wB5C9KtklI4dl5jYmPO/tm/Efh/y
PhnzSWV747z8JC/6+nOoFtugK4WXTTf3HBEU1X1+TtvgH1AyGQIlTUPIKkzkatSjxpRbcUnSsN2K
9mo1xiz89gdz9z48mCBzqklMSnlakUmO4WYnRDlRoOlbwVHX93trEIkv8tYHelwry5IrdnKaYllZ
XUaA5kX1OWH5iQKBy6G4qp7dwlOZkWtRXkBCIpj6APkpADrvjLSsQAhfuzhRinp7r9akNC8YQwZT
s8jJI8SHBxms52Nbd8UU0tJNEbmi83vx8x2hUtjZU/2evhfJB6khX+uRPYbQ8DTkp8+0YlgB+PUe
SvZjRRTqrZvwqtapLZdtxpzyB4mR8wV/PjgZrfTxCSXyXzLbx7zi/5fys4vMyq5n2ncbfwo8RW5s
Fpx07uTb+MbWrnsu+f6/PuUjFGECyLSBgz+YCMxz5cWgqmeQPPB3m12EPCxMrnZBw4256RkV//i3
4Ky48g0Q4aR+LF4rypkmvY23HIGHswNeqUs3O3yfFEm7dDdmvsMXGNB+O48W5OzeATD4KIgmW05b
rqqGns3IfyE31DLY9M43K0Gf8zbGFja2+xRp5K+W+gqafbGil79RpRtBzSpEL6SipW9WARwYUoFb
DMP1dvatQuy3aMciUDTmK2WjzYGY7WHVVlegXkdmlapWI2swFtvFnGuytufsET+TgArx2ZxgPOns
bxJS2TrS8+HVIgSzpx1jwLYBopPjeTs7cTqdYjRbXtkESbo5+3raoGNp62J8edWVu9ObOxMF1ENd
4yd0upAES5VkFvKEfvb4/31e4p/PvMe49ifaKGiMkerG4tXcAWg7A/IBpMC6Cs9lI2Wjhf8uWZje
m2smMO7qbCawXJ1pyTPxn9YM3jh0tMKh4aAsOtP+AQ5gmUTlaX6cd9kjz+Pe8GTyiNFr8z/o0TgC
fukiz4zY/GY+vzBeFM3Cj2AuZ5SuitSqc1dHsoGU9UPmI9aeHGnow3X1zpz1dIJ5vW79Q9iLZYoA
z3KZhKzP3tlsvhfXO/vB/t2eGeEPgvSny0Tk8Vz2nQBKWRIJ3Ay2hfER2+l30Zr/FoIUC21eVkxN
LCIZkFqDJOwda8lkl+tk7Vpud+rR+oLDBrVpWMWVDqC7khf94sbEmdhFXw0rT4tSi5OTFcrrL0ZP
IHIS1otUfjPhE8R5SpBzludMwB343WuUtJrypMvAH4CaGdbWq6Jfv9E49m4sRSdLlUKUlIFusynP
lddulQioxkkVewPc0kxkMWjCzaeMdQ7fkBIUpvQSIutDCx36oWNop8kCjOhGoYBoo7LwolrnDy74
Q8TFlnC1i+YXTP1pp5awoaPqH9xbi+Zu8ocAyBui1j2WBVpVD4Q5wmzG8nRoQXl6YyVMRqlwUPhy
WpETFuazFwd5MlEaXN1Gfw2uIMa5qaBPeCRdlHdbuWPdrOVZM4hN6by3yENlNyz4N2cOehAV/mUr
LSP8AKO7HCeq5bvxmRGxJRlTZzoEeoZGo8sHjmk6rDskUIieTb1FQIWDqtjuoEWfi4PH3+dBgW1u
lrEkVHf8t/CGK4EIkdRmlg+gimfKN4q1W3JDxjxPJTuIICzj+TK910dUc8gWt7NrvpUFgKrUC7tC
Mj9r4d2onaLy8wrQh69ulyWRkm+h/UgYM9334EsBdPt8LexfbaiW2y8453RJrjYSujJ/S9vXt61R
NYI9m3xFbsvvEqKPGqZPUI8erbM7lOE024nBg6KKi+Mh4+Sc8oR3rzSQOB0+d4Di5eq0Dgv9zH6Q
6HS3IHsEAZ4zwak6kFpBFZhPRTYdlyxtXXpMfOJ/axzPQo1s+N4P6G+oo6x+4dj1ERCjqiGTU/XL
56OJ3IRO1OTrOaKgYUcfHaPXzYcHFwdYPzOm5GnkZ39ThARfb6s9RN7WDZxmixvotZkW/Hv5rS+t
97vfKSlnYaIUkmjB8oIAeuR43xoSxcCznwYyKpxcp8DJN9YlropfTmoqyg9wkEfd4fkgHDRy1cPv
z6A2zar2Qc6LZsjDcSMGSBtBAdlHWSZG8oDA4Wt/LdnPanG02Eu4vylgLNvMGx31pvO8a56U8hJq
XYYlxQlsmyL7lAgpmW4P7iLnd8Uw10InyNecXjcEEgoR5ITJv6Es1YQi1456VbvGQOJUs3NoL7wG
H6IqFz4latscOM3XxS6ribyIMfZNGixTCCJpVCf8GzQV4VeDoL/wCywQS+vkdLYAN7Srg7vQJJnf
lmlq4aVy9l94mOYi0jMJyDoxvJ+82GNwlXTY4dsQgFB6LS+0HI0epwhz02j8TpydBnFUy2OWX3nL
ADDLipW1fp8/Ny2y3gSMyDfs5B3fn5oT9TQHqNzqiUufv06PNO+zdXSrJ+Ykkt2Vm+0pnUL1EZK2
d6bbAADMiX2ZlP7MV86cof5VPZ2+fzYj4YzOcZTSS3+cv0XzmJCtw4PcIPZyNukhxdolcO38Y6jq
lTrm85zH0Ng63J5TufWq/G7TlzEQXsEqy+V5mpIqs8TIo2pWRAV2VeUjRjwRHXhTi9BT38ZDXIi+
MB9wijJGUKD155x6w+V0kDScdUtzXw6zKpUt2itY5YWvmIvb5zB46aE5s/FbHcnH0+Cwu1bxPy0l
j7zd8xlZnTltOo9cYSTYkB7zmkHySUSkEyeLNu8fi3khfXBAqzF+gOvJapCtVN6AXWn2+eXVmmwf
WBrXyGvWzFyp20CvT8eGRgeuSU1wJr88TNYr51M6r2I+FFpo4dkntlpdjiGOApJAinrhCy707Xsb
GxG6FPhJitAsf6ehYwt9qNZwwGMIcG+eNlwhkSzRWLEPj3KahpXLiPrF/YLyp/wuDfWkCO9OfnGb
S5x2nduCeG4Kaj+pseOKxvFsv2r65jggoX5eDm7UU8B5bMT4ku5+HS92R7Vd6o/60GaNDDHTtBsW
VMhX2ug21Qafc4eFoXkcTN9NUOmk98XvcEq2rF/jmhdywYikwcNeXcBX2gJe5H8KCKjZd9han8Z0
o+QJNr2KoDN4XOis0e8mXfsSaCfy+c+0Dex8HD5+pB8mv3L0MtjMkLBkdo3Utj/Qy/a3I0xJ8nzi
BD5ftmex0Ds/juLoeZMikFhgDnHigHBVEuvrYVmMJIOhPqwzO7yU8b3/MpVeeVusqy+iNGwGFgr0
gZu+ncocdXkCjZCw0o75KAqXx6DFKw2fvuEprIEsvF+lP6Jb+f4eW4EjO060K7cVCVKqYJ8fFI71
VdCJqkDRSmoQNZVSTHp4EGbhnV4SyQI234y2fo+B4iqIx5lFYy/88boWtkNLLW2M8mrPdHUGyU9b
mtWH5Tf/0mnrrXJlgkySyhFerPCfnrJHQ3gLruDSnHccM9BeSb26L4uc7I2Yfh3B0omfjPzZ87n9
sGq5RcAFiEJHvyjMexFa1zls1au+ETr7KZKrvxBzCWX6C3QBI9qXjMljQbHAe24q8wWA2Iq0v62K
v8dhah+BcVUSyOKu4niqJsopMPcysSbLRofpTwKQN7RG5B9t3QfESq8yInOXkPqvNnonwoKMAX7e
Rtp5L7eadDMe/bX2ivmL2P3zFPN5tfZ1etlT/3xom+5+WDEbQjKo+giuEyK1mnC6T/FsFcMYEyav
yXn3AqZ0bX4KSlAosUdgKb1sccr456WCu9bOyYZ0cGlKGwhXGpovN+cqHtM2/rDhIJSUjZh0nAmP
4zNnH0R5UwdD5kI6qUzP8zgaPKQzREGuohersqrVo7fZFF/TKL+E1k5zs/klNW0QpzITP7tTGwCP
7q+UJ8P0Fh6mZuDiN/qJfNcSBaEkjvjpCOj/nMVBfWmTuAiX4x1iAwNSOhQrlbPoL9CYJQrezsrx
dG5g/LcOuhC4pXwiui7HKAXaLwQ5dt5nf4THruk+PGXHeukpYLwgseF5wxYErliS+EhwbWHDsKFI
vgo1ZPamNov/tiFSweh+6f7KDCrcBK7Fv1ctOXBxxU7JqJhkvsBZDjsV/k+Fpcb48881p3/EnBNn
akzDrfInxilgOooE19Htv5v9Y1hZHeuFiT5Xhm0QXBQAas0Es7RyEWYQJF5OGqcSGmNQkYCO7Htf
UXiCEFf22LcBBmg1aOj+tvpqd6J5gcNvW0FbbVWve3vSYaVJTCMEDPsqORGxjNHIXIn7VDaxq9pX
4FNcd/aivYKyKP46NjJsifT+OYFbGk1UZVK4ALdnQq6lyrpPAZBuzEEbx02zua9edTlEjffWn22z
xK+jj3/+ydM2Jng9C6OtkknQ8V6EqcZG40RWC4GU4nxjRSlvUvTFbfEQaD1Hf/YACXAxDckrUeLA
OxH9kaw2YIFvTanK44HIxH7wKA3mseXrFUzyIejWJY1GV7DHfKvZL2b3o64ZwuTIaLHrsETknsXe
ThmWVT6TeBwodL3oR4GZZ7Wq3ySo2kkxoZ+m5IRVzuduVNwMnefYWafaml88Y4zbGZPIBmqARRKb
cZzYBxaKsZsGqCUG6Ofsh8f3XacPDRiCL0N5UPCJG6FFwr+drsEzEn8bPkMPdVT4dF66t7loGCmw
UUrfUvteDV3iCSJXUfbNeO/0ov5kFHRKRrif0HUh/Z5E0QLGP6YC0x4a5lQbqbi6/H70ecwvNYUP
/SDIhTstUnWEWn2OQwVP2ERh3gLrgtwwxyGGNLRnCmTWI+EiO9cX/Qw5Dw8ZcLu6tjimVAJgiLoa
vTxNOWQKHeKIjQzDmL+HCHLaA2EYO8YSrm9QK0ckiOEkN6cldfkmVbJ6Oae7ByfGwVf+OJqKEqBY
INYt++yBacdz9Tuuyb+XvxnCNYDnTk3gSyQT2aN3ka7/CDeqObNK4H4OhYqdhCe30/B8fuOfBBxw
D3z2p93qBl08KLZrxmZjjCtYZA8EnT1LYMEtLHp8vJ6FnOol35f5obP2Zz5ZLItFtfw9PRX1mDx0
JLTlZiRirOXr9AMjaTi3G5VQtdsDW6ZOzjmCmGF/jSg9S1bxdk1f9/yEaHNDA/AYgvcGhgaA38+A
LQYrhMhw6N1i1yZwq6EAiovqIyHO1hwdKFxsu6CtRmjJ44W7ReQnHrvmBPglSa+RJVLdRRk25EVE
EewENciyVlz6f2+QqmL9X1NiTU+wEVpAbwZu5cf4Sp86dnrUE4N5euuE9UCEsb0HIkglZUa9wW8a
GbIjCGUNVJ2qMjXQWrfidEGzl6pO7yvIvS1v5xxfZ7VHdAEu/k6q+fVe38NomHoe3F23wVy1K6zq
JQukhEg1sI9wNKeXgRUk/Nkc5+3mAOS43pjzBUXhcRMbtyXoS+lvdCPEooB+ysXNaUWeH75ZQIX7
flFIGnSNOVosZ2Avq6VPi4p/rqVBKBJ6PcDR/QRM44OxvBQPtfhIRpBfoheBji9aA+Jp/N6AK7TE
qpn6NhhTz9UhMeI7typYqqDJ//1gb2fxr0eABgLfSc64S9DgXfaEbx0Yl7p2/sxXwcznVKMh1GwS
ydGPV2xPzQ7j9KC7i87bqhOnepfBpdmJEMY3QrA4RjMbvsaszi5QeFp5Exc1YkgM29AP5ypt2uvQ
io7Jgl18SJeD5IwCMmI2iBULZ2L7RrhIV9J0bhKpN24+xGm5TjERb8eg8ZRNSFthoMrlmAbuz8gA
+Ksy/tMx/r67UUYwiDe2r217v9dlIqonZ6M3roldwmqwHzQiUiJyxmDevVS/DIK22yLlAYubWUia
pB9FLK+0enG6K50ddKEt3XyGjMWrQuQs39Scg0rEgD7slzhYQlBjktQVqbFEXojTb+dgbbhw2qvS
/DOnjANPoE4S/3CkJp1E4nwCHDkAwCAz0yZlfzzzGkaxxaj848eLE39mJRj22iAob7MVJoB8L03w
VkQA9qrEvSmmqXGpUqOsfXEbMUv5LVI5NxLZIOlTcGexhOikmqsM34OcQupLKoougZBKSbnbklVa
xWy55Kt2sZxIivY4UIpainfUu42VhontnIo9c8TnJ6NZJ+RVLYxarG0CisSxg7vEXG5VmhfZa/5C
B0izUWajYZZae7B3Mic0+BrsEyXiJOD7W0inZPI+xW15shRdc1gIMeHXMVdtu4rJOJAU5QpZuOyd
FHKqQnjxDCndUPfubtbG4P9Qp8f9FFdoNwK5sMvXfn/r8L8OdBrA7dJD5ziiN9iH+166E1pGy75C
xXv8Wdf/u/XRQshzezFVNcz2bscetu0Annpg/dji7PeNDF0JENmYG7kKq7w3c+majInnpTJ5RLcH
INZ14JNIVTBq0bRsDLI2H5CbKwfsnlbbrJ7hlFWya+8lde5hkhhxj3ZKf6et56jinM35hhP5XUfL
DGWLRaseHbQO1Jyx1uWHG1p3iwN72JZeeQd5Pnkmgt/GdzJ45kPjhl/FL2veBMYE3Asxw4VQwSS7
wzBRg2IKOxO5MQ1DiJAIvQUbSSkOd8RkeUyfeXBwoA29d0VlDytD6+ZeSieWASlhD2JMM+3EMB1v
5oy6v/Nimk+cf0YGr0eorh6QsDv6L1CrH3YAQY/aoN2XTR42iJKhVs2BQ1u2LA9dWuE2HYJk51JT
R4D4Q2wR68y69U6EUvsbKv7OZUitgiPktfHqmwVEALV8JeXzLY/OlEjtU5EG22iDqFFvr3J3T5iR
FZMGV9+nL0Jg/rMXt9kUgIdkZ4Cdah0awh6B15qXM0ulUdYN6jRcrJ3G51bZSyFYS3gl4YdiWIR1
6e8d0L14DztsKh12QHmyqbXpVX/OrPGwvYpZWhK41WLxfch6XJPE34L1Behm+I+GxcOkg/UGXRjV
Jl1C0z3vphRhjUW469hWFb1QpXwvE8RqqUsMksI4qyXFVtZul+imWIjsYIofPs0ZECyn4CLqcbZt
PioIZUs0pxC5OVZFVOI5z1BKdFGnLinrNCzYBhfyHHq3DJcSkaZlts1AK8MUYkUh19oGGGVnBi2r
gy+yh1T9UZhFmgRMlVCWxtxPAaN2Eu4MXQDf1kAtED/TaAEFHiuYGNY9kZCVUYhwe8epkbq6TmvN
2x4ep2iaBdQfJuocedATy8L/e6KZQTCqml2hpPCILFkErG1jIyfLHAjqXb/gkkCca3mE/oo6sIYX
AF+bmYMVCpBn4NVr2tG+vZ4epGqt1ZfWpU5KNdqJ8IJtUuEcuxcVrXo7EXNmS462ISKjPJynKGw3
OKioNP3IRVfkgkyFECVq5ktMearUK+r1sqAU+HU8lcJQ9RIP2P27HJN2v7ijLrgOibqAPULypmXC
Rfp8rjXompnDc3FcCjgbxJEtINOIbjs1+2x0uvWS4W/esWO+giVQvQce6rfM0wdKo2ZxHjRAAI45
x87hYNr1Z6V/5m2/5AX6pHdqYDwwmTix+ZD3THnZdwqCWlnsF8jj71CG4AKSrbhYfwcpX2s//OXe
oFpCkWloaV27bAK70tT8Lx6KklPCKfOky9N65YKTihVmuNnNaDzynOfhf2fbOMf6QaFo+jYALN8q
ZP62nCv1EtWnXa+fF4XXatlE3JYZFTgzlhbHif03ih1G/zhTjm/oP4FpYn2dgU8K5z1A7bMwyxgu
eN90J4WtbnFeK4ah9RRs/ah9zlEpiWllkgPG9vT7fYOo/7ZSLTkNcqjZ/yQBLkUdHWyWoKnHirZQ
n1aCarjuFcoTNoBXzbyV92rtayzK4IgSyxJlUV5aPDC58jKZQAECs52iFVJ1+sBszcKMZqU3UO1O
NuSTEDvpdtHS49jq67UGa7b7HZ4T9SHIfCWWE3V2cZmzqbtIveNiSYUZpDbp+5OSxfNmCl+mLy6i
ba0+7UfRLMcAOyNfUPBEbjgcJoCXb7Tbz5eTjEoDUPAyMALdvumyoZ53g8J4mhuQNeoRf66jtjG8
WbURkWhIr1pg9UIXpyqi0mStcih6Y1Txs+ko8e74e1H6WhXr0J/MhGFva8+z+8L6XnF9fzJFXfDe
SJqch5FQIdC9hYiQgI5G4N3Cz/cT3edMBaEF83gINO33t90TPEqmVTIhvocCPf6w1cAiccPojTcb
Blr2+DvE0jdhYjlfCceWPJEi3DQnZQiuP/rxnjcB5lpMzW9JFvRjihsgggkDNDcreFEbY3WyqLnE
cm7xn91g72e1cTC0A1yOzPbNFpuj9QnHNiilySxubJVR3qos+V//0BXvm/u2ud1O6YaHTRoc9edS
vsZgpVbSbgyiJYXOZLgIHyeYmc4kOBad+SxnIzoWTOU9HD8KnUZA9hGtu97EM6tMXpQy6+GA2yQm
Bk/Gbpwxa4Nu47YylMgzafp7uRgfEVHOTcTDp+pHrCIA/JZHW1NGsSSdNNSLDdjWTLI1aiQLvIUz
pn0qc0rHiwig8zrQauJpT76MnXEYUZbCz1F+6de5rBV7ekfHDyBcCdX/dPNX1gDMMSjpVJhYxIUS
gHmd7MPLma+co4kI55ooHekH6XbAVir2tyIcbm7sweHk3yoc7jURjBaEHckvh/J12VzlS6AzdwvJ
ZbXyXsjkAJc5xLmeCB3+8Hp0qh+Y5CWwkd23gGTIUv19ohE+E2eYBriR3qDHOKK91/UzXMMd/J+B
mNAnM8bq5U0YY1rQhF66XPTaxgTBbo5g2jkK7bs//Wbt7LBc3s6IE8BHeUxQEFg3eJUFoRk6TUha
/2ZrAPkGyowTB1L17Zb/qFwPF0Rf9OzpT3KEaLGJNV/fHGDDukQuwgnhZ4Z3MXB7P4KLXoYpApm/
qGrUbwjmCZkhV3K5NdfyNsORaFXgVqSFcbUx2EnItJVreU1vAW1CdaoZRLUsDlRykxYUx/eo33b6
az0toGNVND3zfw+DaMqBufDaQOoXAlmh5utCVrozCKOdn/BFRVWcrWSyhXN84/vLHJKOAq1tIqdK
L525mDow3f3R+LbkDadQvwto1q+ahdSGYMl5k2NmF6mdObN/VWkkd5yCwa9IxjEYgQ51cxGff/ex
PiX/Ux4B+ae1aM9r3DAsps8Q8GvPWBLBOlZ/15DgMnpEd70CDd+vGcBwQVq8ZwFYAce2SqgAqQ76
gcqcXHcN94QB9kZQAjGVHxJselCFPvYJ55SWSiS0gipeXHVIdNMFV3NpH9bgZAr9ELArHHTU+F8b
7Sqa65CISV393cKWRnpKZsM6RrOo7HQYv1xcsvXUtzfLjb1Nf+TPoZrNzUpbP2+U/ARhOT4LYjH5
E6sJIgHtvOqVi0WPB/WBlb6QdG/zNZ/fnCb2oQeoD88IBvU/tTSAbs5UBHqzll6cPd7vpe0LGW3C
TkURzXgbUJ5XJOGD+I5O1cuduottgNfkCwe7SSNepyzFeakVY4hmx75vuKOtAtNDqpsEHylVsue/
CGTp4EUBEx7XRrjKOY4oS1ptYH2nRgb3XSik5ppU6mFu8kLGhrx2XVi1QeXazOHfRylEM/GJGBBY
OeSyqh0huhhHAUmx6DKNjUMy8ouYL7SMUIFTzP7S0izgNSzk/mik41C2J//dFxKgf3GpZGdyE6EB
3slWy9h8YXqj5xL/vtwRdyiFCsjlLGku7El/wo0MLs6oe/Io9oVAr44YmKmM6ZLmzdaLjbRLZGoB
P7cpM0CfVn9W6mARTYdYGte/xZvykOR6r5aBePa80MoNee5Fh7yvQhlGcWGG4y38Y+akEE0r9EQq
IqSoldxF7DWjT0JeEarGXxWQnSOmFSsKGrGbsksGoEhluVQVnr0Cy06wadqJ1LAKYRi8tHdu9TFY
VPciLr/A7BaJIvyr9H1blUaOpUSWCRk3OjcVpaPcYYfS53f4eR+KXubiWF5i2JhVgVxGD5QUcCW/
D0Fh9TkyhhRi2vey3hw3yJf+QFWz+vDOCqPcSbEBevyXVCOc1wCUi9E2SEeHFfAzahSR7nQzgHsl
0+G7XYUik/EuKQuAHbOLJ4YWLxMYCnJYHlpYEs1Q823B9PYs2pw2Z+SB/sO+HHrrgOHoJAMR6hyR
3E+CIKkYJVum96f+JpNTDx4XkWpmIVkFLfa175JxmeGa5hBiDld3t4l1FybeeAIUiO177nx+kz7j
0PYPw8oyDhtNr7K0eTg83+u93x0pycPeRcTx4L0yAwy+b8cHZnldUop4LpfHcYl9LVQ5QRcX+GHO
6RFjDnB9Dp47Cmcv1pzcptnFancL2xQxSo6gOlAmQRAFiC6fEuN5CjpCnC+G0CNgegzGFEVMaaaF
niWhYiMrjkr6k2qoXIP8C/SW8YQVjVWEU1BQ1ru0b56R59Y2VpsQs0pVhkfaWX4RjeSYEsCZOQvF
UIG7RZfyrV9eA7/O1rWbvWKCySXSN4MKedmNDilGYjs5K7Sm9CvGsDH4eJA8lkQRVFD3CZVmPeKB
U3PiyaeCqNJ+aaSo0sZ/rbFy6UuSr5sUEa+ifJJLKH/otOONFKVvhgTGOEB5u/85x/+Vz5WreTHD
/zTqorBpadXrzbUPh8h7uUQbeymIC8fi3ibMIvo2PDVNav0WSvzXSCDjF3THylzf3Yeze16guzHx
9SOBU8S8edJVN2kOWszPj7fpbQZLqdWRHov0pgrZxYrs9FOMMXmj48WoD6fr0WrLvp8czH+tkPCT
/bEKpW2awKY8+EmJwKFMXRHc+SnWePkAQkQrGwlaN4W59k0PZFkehzBqr2SjOyL3kVZ7b47ATIL8
/uyqSXCEIwg/ohJWA6w4ocjRk+FRNui6PYvBxLFBtezCicfOeWvxUnvtGfvGBq4k2kwnDzzOFtfc
i5/qWX5qbDAbvKyCLQxMPGMS6ZiJIQSF6hYYkARmMFTcL6jzioTXL7Nev8zE/yy+NC5cyKF73v/D
XnQbCmFjTiMrQa/uuy9mcZiE21Mw31ajGrca8mGizuLh6CwT1NQeCesxFaLJr3ZDhUCNK9rLAkzX
V7lrFwqbgzWaSK6zCVNIfHqgu8QD6YQgaTLkUruQTLq7BAtMeo1nD9TO8ZLnZJaXPSuB1zyfiMIs
PispSuPnkj09eGKfs9U9rm/48FYlOEiDDdwE1m7WF6yWj4YueFYwTK8QEgRIU9SKQ4SBbxf+AiCJ
2uoZq+wfuTQaWCbmMRrfkNpYBy8YNiHz8kFUPSo9EzWBBUGPkoMzMDVUzvoewHZjjb0X23+ZO8NX
/bVtT9LI/+9rkVBArBf5e7bOlPitI04zQMZDgp7S8GQ5jNnqoQnKSqcG7psHuIsuhzxxukVH8PM2
YvZGj2NjTD5PpVvmxhgOJZYejo7RwK+NRLelQmmSzNIsMS4i/0aFcBb/TXFdI1MO5zykaqsWhtRJ
py0OUDGHRWQRJc1PZmhSvrZT4O8Oeqfsk+aQ74A5lHi5cIudQbRHb8ac1PmDp2lWl5iC/mU0L/PP
RLsBXCwjCvCDJor2J0vznCyopzU99uQfig1fICLka/DoJzi2Su3eVRRJBrcTSZw0qGXRayBjvzbX
6cnm+kWFtvMpEl2cIit5e+fsadjRhQXuJYxONqJ4qqib0SrnElV78KwQwshokOv+IPtum53liZcZ
S3tTeXJs1J1Ldawg1YzbbfzVWy9qCvNhUoTkpWvgCNT2iwGuIm6ovNdy44QTX7nfu1wtBf8/XPnO
sSJmM04L1O/JcVCzbPhdM8rwKErWu1zn8WF2e5ZvRZ2nXH17ldPFEI0a1W/xK6Tz1nbpJRPkQQwF
ZIOB6013963+EGlTwV0ZfU4KnmPxY5F5Q0TTPAwRDUE+hOVd5iXKM6FELTMZmBsfbG0tI4qvezze
11JtqWIqJ5NmP1lEEQi16BovCJ/kLyxdPZNauCsinhDMuhdgZVGXqPUKNplY+tS+SCPTwN/Oz3pa
A2GfvU2fovYN+Q/u7izL6s1gqubLfSeAhyl1/U4uQOUHi3lk3s73RQS5hC0dBPtraNG3DUxtbyda
Nw5YcWPT/GgzOIwJJdxzExvWCKeUTjxE/th0dR+xbTQp6XjbsnSUX7x4iPXPhb1R/TnZVwtGsGL4
5MZYv8SMaO0lU9rwp7uO0RQndAw9QSPVpr8LJjHhYIUYm9RB7TU1iyBi9WShpxwEMIw20G6iNBSB
D305RSBOZXpMEsKbfk94CKlh5buzO3g/FyoAJf/WL+aNm5A6v3x/dzwm+a3nBtAvZZYTA3Z6XkE7
PgTi260sUQ83Zf8gSzx36VfNixjcoS1Wk6Oyx0lffzgjB3av/gto3w/LgyniDM4DPsP5ZxmJwQZo
qPYySZQPS5kxAatn40q6XAUOc6fPj4is2x2XZMTy5Xv7uphtqsUdQn5oUHUy1NkGM5FgvMxdX8Zz
Ysretzg5+LK/GOtXrWaHp8tU/93EMXwdFNX9e/q+GZpSrJRkT+Qha2yruj1G/8v6u2JNmNHX1+IF
Tt8uOgNBo3ROGafPQcX/cM5b7jIh/Tjvi1iIu/xlDQlpeIMzYRNThXmeWrsztWzKBR6aQY0RUrxd
v6h6bVl0PUr/G0i5YG3QUl5PAigSzs6RJwfZKJWY8Gii1zrLHefTVBthT9sN48NktduBDU6xBMHd
NV6E6yns14KyqirBcpI1BT8/DSaYBQ4B8kaf00DhSdqH9l+Z0B041LQGf+ulvp/gF7X6Z2925aSA
aFTmO+TAn+rW/DpaW0Dgj3RcYrFz9no2G0Ttj6EZYNL2Le7q1jzeUbM76WGtRPWsoBRdxKZwlFHl
hjsH5wV4odZeP/4uRxCy2oH9xun44Y+KvhPXNZFQ/pzf8rWpHAp0MH0n/f42FD4FitnCE9F9fbTk
2nIq3+vVmVRGqo2BneXUN9odS9PNeebCcmgufko0bKQ47VyYMK9zvcAmSVs7Y2jC4bFs8U5AH77+
2M3SVnaSbhIs+nYVcwRLIaRwcBDGaKgyrxUR0D8mMb81rYI8vMIaRvZa3oZYkCwFUws1fbzM2zmZ
JxqNx9kC/gospLDxVSOc0uOYcTPxf7gbFKbArAabk2ajE+4rDeq73aXHXq8GwYi57JTVQJrqElvM
bxDNF5O+43zBV46WDy21AS11n8IaT19futOk5rMWaiXWt94VHcpGgZbyDUNqJFl/TAx5CVzegdK9
Kc6A3xrvUwn69MeXR8b2/uLnI04Ezl5wvRL/rXPdGpbqDSs6tP9opgT+NQmFqr02OmrnOZNWx8D/
JiCKX0njLAaZXTInPWmj0znkGwFWsan2juw+87FLNz8R9ets4W7UmiXCnkotZPPLNlSZrDCLz/qP
n+gOCDZuiZdd32aJ6qwmEvSoX7O/MJdS8oqUluBwYKVC018fPE5pwqd9HLBKOWYBOBOiEEkMws29
w0jbqZEVKNEE0xydcp9uTM7HddzdmVJXdvGPmF21IqLdjt/oVzUwfSYvFpyvEesg2ePhWDwXX+mh
0WKawlJ/nbjjKzBN1fuuI7pfwvzcf54zZqvodi3QGZl70NCWbEq0ri5520HjLIPKRk3tZ9SiqznN
XG1G/RQGws2QoHPM7dG72zq4j9qnDTE+CXidkPFMaF30h0NwYicJcxg/G3orsGaObSRFOnMnkXJD
CNMTKkG+FFldTp/LQ5cOBw40Y5S2qc8MbfZ/uVlRIF7bSZ8aDj67DnsdILjcqr1LSPLNwwPk4KL5
f/lYD4RkDUioYXMhxyRDpm2NgNC1TiTWAKyBde+KtGQQvzTHPwAHryzFLcfzZcdwP3+6R/ybm5jV
zKgjY3gTcSiyO+f00CoDy4NoY+TRkPTImdEpgRqSegUqoN8a02VBdQZy7sKeXPR3MThthguelpkE
WBvhl0uDTn9tSe7dN/7H3+rrBNIlQ0LWSNhOpGR/U8i8I9mCMDDZuMaZSAnrE6R0fS29SSScLXdC
d/V56kRMZc9EyVsGFokG1B/JuhM0mi3d697cF9DuCW4SRPaQLaIggHJSAYeRzTb33bpR4fZGby9R
jB1aec0/+ia+tqFhtFkVDWMvttemGrQwyia254Zw2QPoBVt5M81S+YzP7D87VCX1bliMTuSoG+/6
GiK7YspG7yQp//jY7peyUSVE1463R/guMO7C//6ZT7XgQhPVAVmhRdo48SQlhmHrbJr+w2+9t9EN
EPWETpDzngtiBuSG4HhMfBhF3MRN7On8qt2JON2AGk+vE32L9XWkq3SXSTpNaPGKxDUVcAQ2iL+Y
bg1FXlwhqh3wJTOLaDzufUutBPgCxkjLuIXZuGS42eSuf2eE3T0Ocw3alfhqbVrL2Ddr5zH5Mlvx
ItzOTwjw3Z3zaIPH/hpqvfmd06likPJpBA2beME6ctB2ZxicRF+OK2tGSDxWAIOXdGHCV61j1cjW
aBwq7wV+L1P17O9I/+UalSrkp5lQFqb+vvWPWFfizETr4Ysn5v5QVRla2q50183wDkdhP0NpiJfw
mdCXhB/vBL0Fn/8B7kzDDplvKjlynWESwD4EMiNTdaWl84BKfhX2NJPZetn1UlWE3+rxk6zEB+Fo
BA68dnfjEoQR8tbXVjnfaG5cN+nHl5bT+9ukCgR+U9uNcatwqkY5srHHtIWzDd7bfsjtBz1eoj8Q
DU5eRcLmCMz65/YVjwOrd+kthNX4+uV9cySyP1NdLA9AgVdRc4yvzlKhI3r2YRSR/woWHEN/+YUv
WK1jHiyB0ZkSOHUhuzvSMx2IWaCJsF1a8CcAgwDB/7jjv4k3vphy2A+FCKditkw1YXiHY7+PljdU
WjCMf6I/qOnvyxUyJA6fX2rLyAEgxhuCHyKU2ArdKYTPzfNSNMH+kciWWpgmrnE1JNPx8Zo5lQ8a
e3Q3M4isbkiaXTYF5e3K/3UF7le1+GhDI/7SmLXgDqnKeSAC5twtOSp3Qf6jj6CxorpEdbeelGel
G4bbBV1Vpe24KuqGEARz+6C56VBhzj/a/KSEdyWwtRWvV7IhfufF7HiS4rRnrrUIdAu/JpVjojcl
Fm2ACH2NO2aEZ027F8d1ZsID4qdeTV9GFlx+qUOIE2E36jxnxW1mOPfeQ5q2LbhYD6MrUWjaMAY7
jnyR/9iZGN4g0yptQ7ncTFQWIdWidJjLG1dtL+l+thwmHDskK6utK9ibG5dV1Y3k969aApEK5O33
df+mB1Mx9yALvAYK7O9+w6TJnSl7LVxRzxZq2PINMO52XpZJKb68O1akgvon5lf/2v/kyKeTC5oN
UrZShkuBNyhZ7TcSTJjIPk4bcIAGyMI6Cwc/QnKjUop00JCIWwjG7XJTmhyih6WYqiJuTHwM7itT
btK5+1czsKkA9dne9q47byDd2a6ijuseOARcuRY+J7A7X0Bf7W7VKbkIsCelqMem0SRumWn1SISR
bkfohkxQwtRbJ7Jgkj8B6v5wynVaJoAvaE3//Ak4Y+Q7VC5IwN+zgiScXU4kBL7adb/axaqFOU1f
WJSXBTVlnAv9ur1s46xoNERb3Mc5xI1ykgi/Xhsx+s6O9OaT+KPgZbppsMv1iEm7yYKQ0kclTXgU
0NhhsKZ50/OCRc2TSykbvnJ23zgepGQ26Ed9o0Pmm+Sv/1+bTdONfGh/jkFo0AxkecgN7OhgqCXD
ULfrKAqePJhif1zdLS25wKKkLNZsAeQ8HZdib6oUq+myX1YaLTvt9LfJDmJa4GwIjw7NQPFwC/T2
YmZlD/SshGHfGStQJA6rkFUIRoo7tegT9NHhnRHeS9hW3gB5miG6YJysrwBGA9/Og1znJ5ArwxI8
7XLjZDU8vwTK41JSteW8HiytsNz5aoucis0vGkAEX6rHMBe8jzpjQFsrCfk+xp1EoZZju6tsI4Yn
O3vIsTI6d00QUn0oW/JL0u3bmJjdgndU+g5KQ0Eo5+zZGdW0lhpP8jbhoVr6mrctowhy3i5MvGM2
oNmU7zkX/Av3T872rclPrJW85yI3wYB4zMrZXNVCVT5xozZqhUJBlL3jyT8Z5u35o12qNuQAGM6k
TMLumdrVVrqL0JB5fNJSgmD4xxqkZbMwbUnOzgGS+tY3G+3eCGLD4FY04fqDpRicnYiSwLZGrhVN
dbwkBIGVPYC5dMdJeHUU8ngEwsP55p+jHSZT7qb9By4Yqlxw+NB1Q1nm+bLt3tpM5LQT2/wjRaPz
9l4eigdPunwBQsMI7BXCR/8V6ybBt8JZUsUhBbWGXiG+obc0cGOvznXjXVwk+zqskjDM5vYEDrwT
dpm1qBBwiLiTu7BWrURJRiEDQZmR+8qSm48R9qEeed+bKznaVQvTOB4p0Jdz24MRSAHWH26ReM2w
aoqA1eGmg/75dQJed4RIBfzAzL7urtQb6V3b439objl57nEiDoG0Yl0jtcsFlHwBfw5mi0IDK5zt
VQ6sclkJNu6hKGKsrdM08RfHw/hMuXZtap+k9AGfaO3orgGLTBQxXp+Q6P/chEjMOYZpnanrbGd0
LCkfp+hcD2EMVIqVrDgZzcQ6w5twfV5V/jCX6O3WQNb6sr1uaMDd0/jpR+5vIPJMPSFrSQSYY2wq
x3I0aVf+eeFauRu6r7NX9ptcIs9/1XUSPlHs+nLd2qNvdpXfhr9pYZlsggH0nuqg+JXS5EomwqWd
B1uQGwvD8A++9bFo+2h8+ai7lTy1RAmeEPBENkjYdPoT8dp47gpnsYO/vGiaxq7WAoZw3zpxRveK
c5ToMtKUqa2gbfEeZBXO0gMkdjsVSf7rYdGV55b54xbjr7DquSBpCbyI7vj1EJDFIbCjC3+ocfwi
PiDb/AIOReGib4Z5gSzfWi8BSfN0ykBxU4MpfdnYUNN3DQIQQ1gtzLYnd3xdojX1/DojtfKtrT4w
+7ChSyVLYJP9RHV6nx2Wx+gWcNYqcDZF5od4N2JU4Cdg2Ppkm0Y54HMSXkIzXGIS/Bf+ILBC9GcK
Xo59+bOxKci1ow0zi2JA+6dZ66tAP/2mfl6R66V3P3qL81v7gRFMksi2sRN1c1LwFuC0Q4q01SiU
FB/QJTkXitnSS2emQmVyiQfJt5XxL5mZaIZVceYEJwNMjDl9ilUiQMbYyTW0XtXgmQkbZbqamNLA
wenCY8LLqVmwLf8dYHEP+8bP05sdLpTmrYRbMS3GiueNJHNMQyNgpxa1+d1jVn6QFB1rSdXNv0ev
5LQSFl/c9VwuoKBt+AkomGgEDUrevfbY3iM+t+ygMzdMCOquLhd4NnkjWNnZqKiMOGC4VbOWExwD
Xl5o2u8hJE3m5Br2/qiVDdX0Ml+BHpzqr5mYReU//gfWwUGK/KpfiCORF9lfNUAa4hBiqmqtDDrB
IbNR638SW4nByAhw+B3JTWnERfBdECH63AZJbZ2cy/z4URaP1jmZ39IiID+eGzuDCI/rrwgKWkVu
Y/wgjQUmBiFpJkZOO6DC6TckM4eebea37FCb6yvEg0LLs0VNqoJURPuQ8FcvgyE65Uk9I1X2OCcy
vij2d1eTtGw3qNQ8u+AHPxVBfNd0NbHPM/GzHU3z0oDMLVSrd/SatYVrct2smPaV/BiPjDwEQ7lG
GDzQpMbGiym63Mu2buawMwJGI/6JJpIQiLtgxZIzh92g7yto97nwajEiw3iijO3HAcqXnVSWGmV9
lfgFetkpM/VEpL4QAC2esIhyYuKvFlXceb/zzbk/SmKXUpGT3Lo40M/VHfQp+ev02MwEeP7Brnf8
fGtqoE9oodRKE0qxzvYuhFSkl0X4PA+ApoumzC7HHS4KTj9ymc2O+SMs3JISCOqG7i7uWvNgWbX7
0Isa0Byyx0gRPJkK6NsBdt05J0dxwcLpOaTtNBytOaSvE6Hv2Il6wAeD/mlRR9HESYGsCdziDEVl
YY+Mg65CdDs3JVksksr6eMxJQXs5uytlG1zUYhFSK8SFJxbPkBV5FQ8iAScJWZHOGKX39JI3ebaL
tucEQ3VQgSe/1Ct95G3RCl/eIxAwmfbud8dYA//W9Nibh5u+BwNYxKf5n6evxW+PmQYYaFDE07u2
RZWADbFug4MgqP84TBgHr8AHrqt2YzWmWIg3Zfih07Vu119TmiAElhEmZPApPXqsAz8I8gdHQbub
QUGeRE/kIhZC5Ft2l7GOrQsoWaBTOqXciaYmF5OkC+6Fey7rbVd5nu09UBAkM0q7fTS98g6kB6a8
ETnl3oq7bxg3zRZxHs1SJFhIypKewaNLr8gGAqSF+3Xe8vSzXRW8lQA5ndSsRwqStMUpcPlko6Lu
CQYP1uS+HzTjHQpMvRMvzRj0n7eDfwh1qxvrijZ4Zn+gUwbe46zhRghGMqxqLzteeFZtZ/b3HX1K
bqwXn9+DzcJnVzjzUGHVbUvF/g4unr8OYQVdcsvkC+G0hEcPNPzwO3rCBjPz36r0zLJGbCiCxNXa
ZBHDxvXxtYebNe0AecCtz0XOcUOlsuC5Nnbwww6x/j/RFQ8uhWZ6QSHfk+21akvqo2zgHxZQ2Rla
MhkO/eVyUlzWJ3d3JN8SxfbAh9rt7oHoQCxQUhk27JwmitNrwySN1Kg4pU1PHjVyV13GJ/3Tusa5
d6tkjXlzFOPi41LInVVwkxDvCTM+inK2FGNTe8E9pL+YvPrhjat7hR12K2HeKKOo9QDxAvPi/2iN
0PxLXM8ZSFZ4JCQsuYoHMDgQITlq+5vaffnbi7H7jUm53vcBtc3/trPKSk7ieJlPM9RDoC4kOlA3
AiDyF87W+EQCuVxSw8eKRYmi1DSrMo86Dr2zoqOg2MvhM0hI9fVQn5tmbUEKOqnheRXZmXXdOC6j
QNYEabdFkrvDekLINfGjga7vD1+FsuwerrPqFUPGwVAh00pxeCWfSF+0J/lKoRB/pBc/af0HyvjN
0iYADTOqVlwWjxfqjka0RPpa1f4YQufg91890ONyKrT70G8T1+31ZMNbQB17TPIKKaV/yW58VI6C
YQ7lTcs3JPfzPIoO9phxQhETBK8Q/WL5vsUpv9ep5/1tnAFmy3aybzTlb+BY42SAJXthEgNYbZPw
bWGhhR91xDk3/aeTJTeH3Kl9pNrHRX9ISG5lPIijW84Yp1FBv3P0lDrubYzq+9MRE5E1mlX7i2C5
BSg+xchLHkyLYe4dNVdYf/jZ/PXArUDkEs4nmddTgPlXOM5cXphX+rBFJjuxt5oltShQY3o+30gj
sP3VM4c6F/ddhRzUjezB7u5fxxuoAgyc2fy/PV2gGNRMA4ff8fXDKkne5vCfo4G/xexi3r8HvEXJ
HWKli01Ek5z3bKh8KDpnm9AD78OXq36N6Y4QvsQQY7pfyYC1QWvDYQvZlZYDeoHp4mueC3dUhHcm
3kxiZaINEI+kBd9ZQTMTYUbTQ2Nr8eyQZg7rt/jgxGsWxHYNHgVTqhbuzyFLKpeg0in2EN4W59j2
s9nShHW3K5exAQmIJdkiTN8Pr5qjbWUpNs7ixGQvZ61mpMdFCcb8vKMpQlJy6gOC8qEMX1kDa7gm
6gIra+0Gd+SRwbo3Jg/2cBqOMCQ4izijolCJn+YVcNwu1ltENcVKDnCbkgJTVlL3Vd6yzNRvC3ey
uGqjtNYap4sMBMJg8fD+B0aPBRgSup++8s0jbinLo9MeIic9Ul2B6Hb5k/ZDLoN7VfVlomXNp0cZ
zE/QL8t1GUmB4Zl8I+DUR+YThQS57Ju0usYAtt9gkor661+rx2ub1CLykhEp/kkkBTtjUPYmXeFL
PQAC3qWLLsl4+i9sVVM/6ny4Ux6JxZ6NDkGZBGVcHnkAchz+XotlOwiXCQ+z1Cwysr5M1tnFt3+L
A0D/14/Z76D8XsgOU7MWWvjHDFs/6PYmP+oBusTQ8sF94w9i5YutVzdte7hZkl5OChq95oYpcxka
gs7KqCRPdd7CiU+mgqHQ3yBZ5/VF3flPZhcE4zSI0HhlYSMODYy/+aANUSGgColMr7Ec1LAlMFpB
ThSz8nqVZGqSO8sBqahR4kcFDlCrpgVgp+yhUQeNcvxTr5Vd0HKHAvheFn8d02SifMY9+VXoQXKR
sj94iOk/Jga4PO0rnD0VmdQ3U72T/3dEPiXHrJoFDN6iKDBKKNGfXn1U2UNqlM2PX/BYQlHgAXTR
IB0g71vH1LfWBgTAV95FyIkHb5WvarOpUKkgnQKVJ6Xk3AFBlH9aC+SvuohuwsWVU5fkPnnjzPOJ
ArXzsAriEd8Yj5Zp+50rB6g3Hm5yLP5e/GETg68xCX4Gk05yMNv8rDNyJD8zN9UkJw2FXMSnlwCX
hWCKbkhyTy0Uj87z/UrNXxJ2Y9j7wLFyk1YJnthjpxuuKeA7Vu+VLg7QU9MC3Fy0zEwCQA3XVp+O
Q04jb9eiusEMvmGLK1KfNGVOb27zX4Gj27bNA+jOd8o7UXQj7Ov2zScgmPDd71KGWWn9yXqpDKuM
D5/kZPuL8VRP2cnZhgvvZkivzioYJZRSPnqOBdLloW8zLYLtMjK7SZSHu/Ngv/9Fcb7z9uMZ+QDF
YhW5hRGm6HwvQPgilSUxIxaJpg540d8ReY9h1MAylP37tCKpMuSHyRDQZVY2NMSzn85tCYX3nvuq
h2tcgL1NSSZvRYzgqUKkqqMNRdua0XHDM4EgSm8qQ4HUHlshY2DW9PAzkPeN/Pk+uKYVTtoUq7kp
+HASjvhTdQ46qs3QhrWkeY3qnPdVvAU+ZKfJemo1RrXxtuxCpivTN1Zi0tv/LR7PSJQ4Igh9Ygiq
Gg/YPngM7itda7XsuWLj+j59x2oGrj4iFriqIj4FLGt9d4UdncsiO4u4lRb3spH+kDzUOm9Ko62f
wzpYvLYKthEDYOFNxQOLq4V31HEdLCkTrCqP4M2klzgmibeDdtqJrP6gjKqyEQxiwjoaTR15+S2C
2IKca5tl9KDZaCgRNoIezs1odtekv5JiHmwWBJgaPoxxtTlPZ3pqCxUX07zRmHOXMzTey0oVHVgo
39/C5LFRAyjgG2XngelRWv68aYYvSXr77MLQFceHAIz+KbqfnHPxlOh+cNxvAWautgyQDtUnC+Z4
ix6AQzfwoURqJg0vsrpligjrnuOgiX4m9o313xLtgq0AiXG1iDz4AIH5mttuh6zgN1iBjel2c/RZ
8EUJkwp0NZ6EiOOfichKh/eVfylwSf4lFZmIkIx04EXq0YetmFXq2MIt8waGp9/Tyr24iJyV1wNO
gFS2G1EwfVctXIK6HXPGFdu23efQ5AD3BgfidHFcHONW+vZcdwcncRfWZoWwM8SelAyCKu1ciD8I
w2Vea8zvDl8djK8TSs+6bQAO5kQxqWxUrmGQJMPHTkltOeYyXvw4meX6OZKXpOkbpsJqy/xkZzgG
w05m6ubw3UU+y3cGrC24Y7GGQNLyxB+75TJ4LqKAo0nXRZzOgBYz3KMBldKWfWjrd0e5TqZldq6V
rDVqPXxuay/IYdwX9cKLQpDtGfS/SIPqJOqPabHeKBXZSHkAKbyY52Ml485UGwv/y572FQ0dZoPW
p0bn7E4OXMoFZyFcxOmydippQAEr3IWFiX4JURh9rbYmV9Ut9esrGpFe11YGkz06p3xsIga8/gbf
WRGG8rJx48z4IVIXOnQGEMC1EQx2Fe+OZJXS/3GnTGFHTtdYMzntx6gN+Y3p19cu6zv1pOjzP/ZV
IvzEATZf14WjL+jHsnN0xPukJ7jckFLLfgBHwgVWhV9ZjTnbb60k82aDarO74v9s2SkNUjSPBy2d
9LBfX/xvW2PDFq3dPvDDx42vKrTPojiINZ0cpKEG1jbycH+mx9NWJMZPdAt8OmKMlTciPX6cSG/X
RI+jH1K3ZsFl+8pPEWAy4RZfchHswlgxhHOSxZuMn2Gb2WyN1SBIFaycohkJfVLcaSarNSgvoQ3g
oSKNe3AA2qW3rGWTySYvixUffCDNQvE7YlZ4G+ZbPUt78X+1d8ulJfz7lSGH/Bp66VLWHDJPrAID
DhzCcBOszjgffPZAS4uYnijXZWdDNjQ5H1vfPAQ+hTD/ARu1HnmAFygi/uhBXdvT21eDjobFXuWC
swwz+yZsZOoUBJ6s+tnJuklCWgLY9YOAF2F2cpEivqvsK5GxVmbx3gRLn9RhUtjhNGHw3yMeVO14
GlWMtRps/+agzFmbpUAwrpdz6YFEBGNneuVquuezDQxvY1D53BpB0DzKcmLKlQPZXH8J9mEwQ4t/
Za4ebdgdojoSFwfp2GB1kKJ2y97ijEJL1LPe44mAskbl+ZfiZ7CbCxpA8DlCE5xOhBTgsKPpa3dR
senuDavHyLfVzqx9WaI5n13C4YQU3QrLzLZ984zJER4LUfOgLrch2dFgMpioyjdmbMpOfZFKgVNU
O0geD+fzFYtyO7IPl6UhQMaA3u/yvleSQAITyv9j8zNWJq4l1HpqHI1IxO/ndO8b8INy5QR9sxCj
jyCvMPkOYDj5MEzoxZfSmssUsLtpTNP2CpZTEPJpKFOsoe/Q6SV7lkiIrDx/g7si4fN5ko92RySa
xxAZP58xE2LMHAB+EFZuHhdnG3N0EoZ7w7LYUOe9H38RROn5e2u00WIi1JQs5xld9XV4Dmh58mdX
gdzeTCpX6aMSWmkl4Lo+JndWuroweCBDLl318qKmUwGvUy1R7JlVZSiRDBRAwVQGrYDr/F8KlFVO
3eYNk60o30/qfubEB7YS651FNMwS1W9J3pxRPyevinIP5WXqy/m/KBXSXGdtR/kmr9i0RnvyBfWE
nYWK+FesrvVfpqIWySPn9pnEhfdyvE5CE4qhdJ/kH9wFn/FEr74lbkpejsJVaa1wZn9OdqE0Ngs8
LEy93XRX1AakMRCRheABFEC9OANa8o7K030i6UTIRzx8GYXdMeB4qnw+KW5wgDuBDs8BXAp04l9I
NHJXnOS2UUvzgawlmwvliKBQhDz4Oem0P+Dap0VBzqu3BzmOkNejqpSTEBjuWq20gS3D/iRiSxXT
gkffxD9XBhWxYwtUsErrctq4bOOObtakjciRqNlMvFmIQCG93NFPoJM7OqAzRQsPrMEhCkT+guNS
Sgv8ettRG3D0PeTbBhTTwFCposFYAexI3lggW7KMnk1xvRpRky1peJvPW6lVUiz8R+WP19s/QZfT
ziFtx6jJIKunkmQz/COwygMb0ncfgZIRlLR/iFOYcqA8/xXeUJSKC1eDg2iR5QieS/nl8f8jP4Oc
cspKEf4xbNUcGRJ/Ol7nN0GxSC9mouQXfkE0yRZxezK5QEQYsnUexabVa2XDHrdXnB9KdKCjq1ki
OWdURh5S727WPXkdWsK0NUz0n0YJLGaW5AsOpRrJtuTuy5x4/LzWV84Dqp/wRyvU2Ct85ty+61+o
K2oYoNK0yIykMrfEMpYMFfObgvmyTyHpVJIxrOHeT1Hp1sJy/bFU/PoRoew2CGy6LcJkYrETDysI
vflOoxvFX7bNoajokYd1uPfNrcNTFV3c81RxRfzJ9UVVIvM3RMM1/S2zwLT07K2mreI4SPyztRVo
ziUIj+5DP0CWA3wLEEpvcJCVRqlbZaoAMVozUTHivaDDR9JTzAjjhUwHexkeAuBa14S735LaIylK
Zr151pI0oFGdfuH4vS5bXnNvM6e+2vZal6TsA1xR+GA7990fk5zN6JKm6SMQfQA35dlNoSQ1F9nT
An75k9NwPco/kxonyCrI2WPZnJGb4j7cfQtBwGstwcGE/Tyu77Yzx10zJx6egORIS6SYwjNfISgg
Thl0Sv3VYj8+6exax8Bz4HHOiYWVFXZiXDPa6jI5xuLk5Co4YLxe3Jt8M77MV250ZzFz6wch4TS4
rrZyoxVuWuawVVSz2m8tnqLrV7LmjiVrlhsyufAeOs7xToIjb12EGmSrD84SgFAts6I0flvIYsu9
nsNTKlqxBB3evqY/bCnzuQ07jlmbfrhIoaJU3RKeKWelIfHRpDX0MoaNBwyvTlKxIoPWkSsVzwO+
EM+z2LG1U24g+IobTlEYnoyFpMUPpxvopt21G9lwqoC9N8Y6v27+fy7lWMVnTDl5IwlfyN7NoUxr
4Sx3wvRZYy48v9YhdRyZRgcBEuPTtu1zW/1yvmwSxwsnhNaILSF24G/tBoAO3ufBfIB5CCuPsOtw
LFftb4JZFoj/W/tc4Caze8PSHwTgGE7eK2cCL+Du03OH7nGKpkbCZokGfnbAL9ZVgImV9HPS01Xa
Qh6ZNFkiKc6tPbX3vRnYz56BMIwHEDLP4PKWgdiKJOzWFNgjZd45B/R3WRY5pPk32xh0WhluJmN4
oHo14NIO7N3sWY01ICghTVndOOocQcwwfHBayp/DwKnh1vy4XlrZljLSX5ESCUDDC0RZd8CYZMfo
KWyyW66jAMMKb3Gua0qBq/Ia4kvz4WteBdHphV4QTnq/Z/JmlZHxkG/QFikoZn6sHfiwtJjq5SJv
C+rC9c9yyAIVW6kqiUXbfAyn5A8vq41sBGPITbDQoZl/MiO5hb/uUoRQENpeHVW9hayCcMKFYfmA
mPgM1VrcJt/gSyCE+0Qa/qM5lpoTGSkZRR40txlmIqdjvUP6DXc1UJu9ja4T8zTk+mhfcxkleR1m
oXDQgMJVi1NjHpX8HyXClE+Stvxr2ukwoyhUhgyMzHU0zD+bDRIqXur+i171ibf0Zcizh7zSQxZd
8JIPH+TtLkUSdyJW1CSFl24nJsbOS2HSn2mQzcnq7CWQINteNAGcKi7R2U1FCMkgtF27nELLTjfX
Xxav2COpDSro/6b/VY2KVQty7FWdp+uG/5SM5F4tKzafUFx3o1K44zBJseM4Z1aoXVAFnanjSbNU
EyzwRXY+4XOVTj/7Sk59GA/wUyrh6C33gOkyCn40LRTw453sXbNATCgN713EeBlcVwGbMxM3vAav
ZCxI3n8eUNW7mS73/abMBuW0DRh1940yhyza75MHxpDve/T11/eLoPeBLke4pp4HJJjcujoiK9YD
QhZhNpDqcmEUSq6oRq9xp1SW7mLXc1wu3iUSpQPvk1a9lngx/Ywf9kDYLb9PHoVTIMcs9G56QsBB
3ZqUZF4XvQT3O2tQ3l4LWfa+lrU1entmCmCvoaRn8QKmsCmrMChhL5oAmrQAhN55Dc8eHV5EdcJD
D2Cx157YDQ/xOEbrUtMgWTJzYnfiYMs4BdcWUyxc9l+VU1IFh852XeGJws/tdcuYC8YwrwcCwT5f
lTZu936IQuhD70F5+ajbQMbaKpuvvN5G8TXcUzwS0t3/yWHBx/JoRgODqj1lp3ywZg4hhopUBxcn
KdUs7usLw++T6tSfNKapa2yfYOMlV7GvJEjJdna1IKeuVTJd3DLIyxtUa91u2nMIpCv/BLHJjn2C
txsb5zsrKQB11w0MDcetoP91UD9UbdB6Xd9GtxSN+48B6rkgT47vX2gfyOk4UPkoGy0HSfIxeo1L
TUcbmQAP4Cg4XWkyAABR7yzCPEgeCzfoIBgUz1ZjBsUUAZcErLhmt97mS2/gwKNiyuFMtvloCcVf
SLvZBCFIC3SQ9p4akT3NPbxEPRsWAvpph9hpvgNr/Z1e2N0KU5+qpZDsmaYJ2xn909msczJauIlY
zHlS+JUpp6hIxQ5OVsL7V0cspzSYmY/5LUhcO2fwH/Qcw9GMHtVskG6EVw6aI1jT1WRrzTL20vkz
opKllGJ8mMqj4Gsg6OQk3qLmt2Wgx2Trwf5nHWvNjbabMYT5YzMrNyKbrO3BCEOQLeew7AIG2gA8
M4rJ4Yqohx2E4tF7s4H9fueCcla7zMFR5WE2eOMBM0myFRMkwvG0ZIlXZzK7kwYczeuxnO8PtUV8
bM88t9GKVMArHGS88J6EbmpZCU00w+hN7d48GintW/BXfSsAtsuVFks9sZxSgMtMWTngV+OnTFNl
IGTz/tMSQ6O+pJP09DNZuDdBt36ZHQ3KGt5Gxa9c+aKWQAOLeYslUlSpfqSOYgxSrJJxmU9iNu7D
/httslCMMMGb1LKQ9N2z5mjM8kY74mArkgGkL0a/31LKQV9Wz9QFZO/LGrQNzA4z4t8xxABfkjJ4
h6AmaGueIsAe9VLj7Qxn+kbXgIFklqq3E5/swfzfhxmvtP3XD3GL4WS7iK9f2RwxphTt1RViICJG
fJUXsdMCy3Ya2jgG4J8k/x2AUbBFr8/FvUZt6URx6h0/7nIjtnRaPegXAeZXjbSJayBLzkVet4Tw
/xts59CdfgtgJHh/gNZ5DrJZjpPwcYvmcLNU88vRroxMWcjCQRfjcjX3jHjQkta/KTiRPjGSy+Z7
Cmf9PWII7x1Te5TCP8h8Zcm0JZTjNX996m9+77fodj6Roj1P9WW/iTAAHRqQV+cQMvAu/zWF1FrW
Lr8n+rNO2wxcfz5j2xbtIQY3cRIsTvVVUShXxzgqmZbMICBXJPdD36MDv1KsG7gbbC3ymPoM5in9
TW+Sc6ERmton9HcHLeulkS20lWyYs2k3RH6ipbKUj2n5W05TaGBXbbqPjsTYiPS4oaO2rhNNUcG9
OGN8TWU136YGf7UR+uAzDFWg665JRomtnkpRhKb/e8fcQfOP0s3gXihfqtpdKxhtt41zBBcEFAI0
uipzkcXqqyW6GCxdmtLjHcjPEbMErbWKXKg2zpQJX4PGV6FO22m0lIR9c5rW0OPUNt81qxTNjKK8
xPnFSV4mI0TBa2qIid2dsMs+JQh2Mu8zgMqO7R5/UqLZxbqLO5x1MIEjQxCglirwYqdVBwb/1P2S
xx8m1FOTQmx5GIHNhzzko+jFTfFLeKh4bZKf02STV0jDH3pz9rwxfDgwED2JhDc2KbdAL07Hw1RK
j8r0n0GJsRmzo72bzug2HDvcJb6H5dwtuluXnBGFwVo+Bzxw663W7zrJJ9v08NuC2ARFQYuytmMN
vMDphPNOkDHi0pbLfS7a8uJCDaXPoK4wWiHvZTxg6GUKbdWCp6XWp/pkEQFhchzjk6rMhupdWG2B
RB8tLHC7DAu3CC7NhF28bJoqbjbdldmki7yw/AugOAIK/DdLFx+BWqD/6qpwTfK7iBDp+ITXLjyc
HkLxcAU+NGe8Q7EjsPKTx1IsFkYbCRntUwQzWLE0Cm8fRsuKPAT/d95dxRhj4JIpux8q18d4mkDQ
ocot7Ly2+kXDz/+LMhJobDr94fNul3/gMrSlTo/jSa5XrkFWYXLA8CLv8ZwsBvIim00KTrV3bLHt
HsBVzCgBBUOE0aPxiWjPWmBxnuZqNsaIpYd32O38xd07WF9WhjPBB8LEndt/lbCeZkS7+fmmobo8
uLJf5kWvLbzE9fnyVBllKtdp7E496i3nBrAsRBxbEGiyRyiNqKylOk7PdqCvyk2/4ti4G2UhCBDf
AcRW3LNxzX+JCjaKg0ylIRJcHlaO5G3ONBtlICFbp1wJjXFqnvXToLqaQJFJ/zwgl54dwdTnrVdu
9YO7yoHSp4jORthuiLRYqt7AFUuw/XO+IhlmCsB9Qyi1caDsGlXuR40G7isjI3xEuR5BM0GsxBDN
8lxvnDudys8LYLAHdmi12Q8mZjNGY/MaiJNnF1mLD1q4hEx89vIiIY2bqX1uIOXeWcO3CzaTEvNz
OMfgbR5lv2NkC/BTG/SGKyvrGJ3ZuUARoj0s9vwgQexsSQGVs+2VQLSRsA4eWmrjbPtfbFFOy6Z5
XGVo3Sgq0uOWpfr9O69MNpzoErXMD6cLx4z9Yene9vg6AIpgjbgCN1gDN5+nx1UMrioppmKghYTU
QGsuGjUiZTT/Dji+WSR2XcGtI2+UyXb94dudLEAl2VgYUcaEizcimW1JfNNc+ijqg4faAr8XJgZa
By7qKB4LIK8HtEzp6zejbEY6c/NDQK9otQZG1kDCPDs72aEndFI7sAf7TLa9nzd/dMreV+Be97hn
DZWWuty3W/uyE/k0Bc+eF/iWDI9acQm075ia+Bykx7FZ1g7v/FdVPlD+fhKbcEZvTT1KhJftToWT
LGcpDb0hQ1vJEr2IvzUCMBYi/BRGNBrUmPwdb5AHzwLDUIi7zFMNhueub3Wn3pOxW2xcJ7xCWnq/
FV5f6q2qL4PCESWRs/6ZKJGh/+ZTek71nVTcdRYHwzB9ah2CyV/60SAppxWXmLUo0hxwvSwSfDn5
TMJGi5U0c9hVelyTFcq4QXefuGpFMdgeKqwZip6ZWMgyykIJREh3qWJW07XDaUJSQV3QdxEa/WC3
B+Th14fzwrAM2GrY05Jn820MQ4z5WJfE3I+7n+hQhomCOr/CJkdRf7R8bH6RlTxY0uLSWMi/KCDp
EFtK46uoigCvkYFnUHyR2uhvTHS1xFm87CD1x2yHfkQCHNkQSJmBYI/NEmqCJrVM6//nK3OnT5AB
PaZOnLKRsANS7ANHVvaCzQ64Mv9WlPZY4tEtYOzLqJOBKRoX/eFGJU0X5oE7Uz67gVCtVx9d0KDt
OSIiNxeD7/0UaI6M+sCodV0ekC5LTqvB6kwCtc9CDy0Q2fX8/p9ptO/H0o0Uk/Q29p8nUAZLDc93
jEUW1JCt1NXcx6KAptijv6cIrSGuxVHDviDd25ZcATjVUbIFIROv4gH5Yw2eClEyc/5SrB1Ivxvv
uc+MKbwn6DkrBXufpalcZoK7YmOoAe059XkI4kr2LWclG7gE3+kA0ZcClyhE/9IZJhLYLVZiN0Oe
mlFHXm7MWwM1moZs1EpXa6BRYXdoCPgcBMwasQmuPSaJf/sJVc8qFznirfBX7v+yKkqMM9ZVwpqo
IrQAl1GfAAVK7oOfFYpgUdQS18A21Gw8NJWHWOQ0UtdHhqzzjouSaP/1GbkBWmNjg9CIitzDc4X4
OytTzOWoJ+wIgVRbmlUi4Gl2Lqedjj0C9qFR4MIGZkR9nyjUUbLWj29Y7d1hgSC281VIjaCElJhK
5LtfzNSuw8x5fONJfl+X7W/xUjHwLC5Tnj7hc/S8TzV2OPcGcmInnOKZVRqfpvwBjP+cIU7hYyA0
Fwmi0yzMNkORVcX5SId9FRDgrv0KY6jqWdIfMyJvmkTrnHeZRaA6bVv8KhlbBmWMr4CmQO9BpvXd
nY6g9o6HquSqjORUj/TRmfJfijjgZDte8W4jDhZYV4pMJ8EuSwV9UmW+G1YPOPYMRtG+keE2t/Gt
34I45/KTFxk9fqDEVpXVP2ehGoAMsl+WhE/l0g57BL/1mHkuJEMp7eNa/iwhzqWzdaPLEQsTLe11
Jm2I9ndXdYJyXwYofGZMjFp5Avbol+UhbKsKWni9Q/o3PI3L++hHveA3ZKeO+qatgkhH2HaQxpgV
kMRUnQ0iKIZxmeU/0GbsVDrYD/W4YhL6FhAk1MFtKVKUYD+SuIGysJk7xZDpfCCZw/o4R/Kvk4yO
LK34crhmbHq5X5VLRG3z0iFF1CbIbA3SUyb94TQc3xd1D6ET/3c6f6PLMKHbVza91TcdMdsQf1Kh
uNbMe8tQBBtkq7aA5MQOamZy75P3F1PT32DtX6wFjGqSy2WPa/yfjbU82Pr4afXu2BZ/DMg26GOh
VXXsDaIV3XyH8PUwiD9Pm7ROr0MOEDo9XZRLxoFtRe5UDvvz+OAZczbrGUOcyLPOvK5zf//X8vRt
G0u2ZqQkRP/5E768T/aAe8epuKxIbR4npmcA+HeWu8fbIECMXMpbv1eFzrAOnHLdOHus40VWR4cg
03xift+k8hpTrNMx9+p3YpAnnN+rdIFRpaZ7F33d7I2Hyq1lguA3DUai0hLcDVR4NgzyEhnAyrLM
pNecvTNLJL0LnFZsUkwDs6DBEXG8g4Lb+CQ6RM9qUwyfQpwLm9wLAt0xeG48z5PD1aUSCX2BOcZT
cuZ/RKH0D3W+ghC69KqS9pZkZTEQiqSlFviFtUTuXFOGAe5vqo13haxLvO7iD6y9D17JM+41TzQW
zPyyXsOyYEzaThF7hCoivO7AP2h+YKEelMJow/RsUfWBGKrzF68K+IPBRFGJ+ntZNiAwp6/0U6zr
vPtXdtZmlV4s5yIPUsVdJRXKBRmzAaEXcrc4yruet7TnXMxDVA96ke+9XEc+PR2sR1r8/wwD74gn
ZgmAq2QCU4LXUJ6r2fC2J3AL56Cmeq5552A+fUDxhBqGRmzuRnJm2iUmBJqS+dhBaeZQtajmpj3X
DNB+GJOsHhoaVWGXlVC/oqmM4UzSGJwT5IZUqNQfAjj1s5F8Xhy71QvbVrAr5odPdRuPQcHwH+vL
/bVaH+McZzsPo6cpGt67uDYcKCTS4OMtmuA45XFcD7W/alpf3H96d9DK6S9kLg16TRFzjCK+tViv
vDt38iwFtb5ebRMWrzqsATDeTF9OaEm0uccrhME6PO7+cYPN2ZebbSyVo9J75TQq7yv2mqCck+rg
jiFiZRYqyOtKNXjEGPTLGGXLGjPkfObX5t8ry/gc6XhieBBzTIUEOrae9+ciyTQr1vNTqqegOzlF
xmJbo700K4W8UD/mwTmHIwU7PjjtP4X6ZYKuwjDBbUS0JXW3jBUVUGGhh4ckSGa+Vcr6N5ol4l/S
JY96UL4T3fP/w969lQykCetcdkAL/Fump5O1AZCk0gnqVJe+z8Jf9yt6rKu9ESrG/iGFVfEVoPy9
6dxOrIIj8BqqC/3OPnlOoioCPqljIEhEg8B9UX+kvLPMw9wlGpzbwUIe6zdRlNlbBjTNTjUYTS/l
qjaf0F/vN+J5pHNGKXqvHePJ+bGcBQEgfs5VkgEn9K6LJARTLS5LeT89dInc97mYCK1Z1Kcm/88N
yn6W100e1Lnz85n7VhNTLK1nQV6f+juSKkR//7p7m4E1gf8BjIUGfHhQI4xZIEi6HCP2+u7Iv2+A
bXTDaiVEoxV7uUTfQ2y7MILN0veF2BmUxRLjEfe9mT3Pfej8SZRAVW1bsxI6p3KbYjC0Q9GWKXjl
w0TU5vp4grUC1AqZ8EQWnUNwHc2UVhWbIpDV8Wfntxe7zgy6sj9YNz72D/Ai90fCq2oTj2O7kN0S
3BpAgg6HBBPUjY415rZiwQfttGhMd3r+wlRDDUxMyBaeFs/wxAUdpu/AEFhKFftMRp8b2dyby30l
XfT1L9Pu72mb8XVjCzKlKNWqWvM328cpsp7vfdmI77X0Qopnz9Og3yoYucSmndTaTU0G+xAR4WFy
9AALHlddauVGQjreVaBhDmwcDRxBTJ2rADHX6mt5L1RivbrWjOwMtazLaZyXnZ+n22+fcFhRhNdv
pQ56tSolcRNlcq8wUe43G6BNtNiZbLP85mcPZ/pyD/kZUOlqNEzaC4m8tLLzVkFMChYNx8GZUO+u
G4jCJD9LEmF34bRZaVjFi6PGX9ZsgX6TD8k5upzm+to5ZrCxtbEX2c75XJsv6G8oMS2r8CilXwpU
Ovu2R/knn2cS/1kV5XnkIw5LCxCspZcFnBFc4QF9+6juhzd9MiZ8ZoyXVJn1o2h+nbRwjNUB5bgl
Miak0gUkCZ0UcX47THaypn7i9VONVVJmA16SzGnXfMd0lRYPyWiZdHFof8LzjWGws5ANbbaEHvGo
pHIDLuOtlSqyp3s/7hizsWo0oOWZm6W17wPAmP5K5GzQMQEf5UlC/8ipu/3bFitQekbJhYPF3TO8
7HpmNxXPD/AbcWHNY38aHwsPXJaWZgizITaDBSngnG33mqQA5MZ6tbgK3S8zCDjahNlsevbdVQRu
SfuBYZYsrbr1bSgJuX+rH3lrNUGX8UnEEFtJYNimYktQTVU6NRTOATDTSotbdUzkca0n9MKli4oS
BZePA2LnYwwMyrVfeizVsZWxkBJ5Xxn30D8Hf7qsmsqELh8POfoZ5K32Ri9VkHvBliBOberQAwJG
JBvVfWALl4vyHLNp5qPY7MySb1r7vCGIpD/UZlEzNNRQBPmPwTNXs7s1w32fz1w/7lotygXb+RvJ
lgLCVF3N1+dtB3V2KDqcN0uUX8LxFl3H3tRqwfxebixk+4mK5z1NGezGAuUGgKAi45RGmMBdRuVJ
rmW9C0QcGsPKz/sNWPo1atmrMsgal/9qNB6diEM/s/GlPsYw44q239h5YmR09lVrxi4kuXFrjqlc
IE8Co6vXihO9A9l7+YfDkedF41FBLQl994BVX2AD1+/iS7+MjSYMLHetYbQ5lB1evNsQt5PCepsI
gVylvP0V+b1ut7jYuffSHMRZ2ZHDMqJuL+euUfF7cTjogqWtjxyMu6SVqP2wK6zvg2M9ssr23nnI
nJvqgiEIwP5y0QJo4EnGbsB9xDnfpC/jR3L2cAnFJMEKK/J77D4nKABAfDZ/lRIPgZzxmJ/kzwXo
kKmTrXMFgmWJWKNoxDd7RD4QUqcLK3H9A6oiWll0xOGThebDC23wFYME55SfK5TG24E+VQBSsGjI
SDe7KYUEtYENaXofs2xOqfiELAMms83cr++sgQ07MxVdtw2Gh7P5e6u/llv7NkVvQcQWJUlm9Sgs
BTzah8h6dO4NM4zqVFeSkZ94xbVUk+/zL+gfkXzjIM1JrmHwkFxK7g8U6XY1OJnuOySmzPBFH1xY
Cexx9FBvduXJJLCnyJb6iI9/RKNgEJy2TaJRJf4JgormGFqStuuuWZoT+EVrYEo6n9yeEYfJnwiB
iS+EcR/czOECSIsARrHL/zO6+k7XOowBvqeFoDdv6j55f5cvPOqacKaCwjIjJTEPWqplY8iuoD/k
TEfmdafamMHd66gdGJ/gv9gPWjwvdicIolk/gw+PN1R1qh3b93sbJgxqeJyxHR/M7I9uBIAycw2R
mmuFXcwAQc3NISVfQzvHHu8FAQ6+tPkDrbuJFaEKt5eLhNxbTpnFqxHn9kgtKvP8Wg5WgTGQO2mH
sPlk9wREX0ecNfA0/qR9p0zXQxlZ2LdA8wQO73xiUoercS65ZvFDuYS+WLkvG93bJGCKAokYmzXw
YzgxcBCfnFPFljtROdT9N7YFQTHLjJplnuP5mm8nVyn/laFo0zyLhz+cMGPAjSsmhaUt4FEjEmGq
zK2edoMsLMuLVPkuevNyelDth1afE18+29ZLDeCwpo5fJiL3C0K3pDM8MXKkOUM6LwQPkRfOhcCA
NOLza28KNckdoVskO4cG949CRLyORQ3hm/+qE0HZ4E+4a34Cm2vIxUWa6kN/g5GdZ8M4lEqozMdv
AxKasYZoQ0PgjZMeBQXImsU++GpAU+ws1Sto8j38lacXhSMi6qlvX0pazmeoL0NsoseBz4Gj7tZ/
RzyP+7vj3s/qw+wmo80XT41NPWBKa4n1RLt3Iove1N2fgoQzXCykHvb6HaptIEHw4WfWN1OuVGIu
S0PZPsD1RBftYLTRB0OjYFhlLS32Ow50kLaXBRzPf4eqsEEzRFB0g8iLeGvcs+I9YQKL+kd1qooJ
gLqlogXF9TUMA/WxrXjvOXHjVqpSjXjy7KCEnayx+v9oyKS4uVXoc0Mu463KACHUGrBbEMW/XA3b
jfE7blqrbgVDwWsdo+icBlt83tQhjTopY3xTdnV+x2Hxac9q4SfU7gxbnFJ590F7J9PEZNr1d0qP
gi4xfqna9pEz9Wc6LFl1yggWT3j1z6Fg9WW0tVkFvc4CSavyQyGneqJopMqSUHnnDsak9hvIREYi
aTfWidAY3B6NDjlcG7UV6uOTlS43acXwxiy7HSANW4z3mWC50VtxjRCCZukyKt61ulucJUk9Hl5w
/PWhxAr8XbhKqKIm6UetQ6gLSTR0TsoI4ENQ2pKCcle+Y3kJV6A0SPJG/wDjBPdiz23fPv1BuD36
I6RGicDU2ZA/reTNGFxAKvm2ySBgEIwfGHoDwL8TuVmvI7tBEUYtxBmU22zFvCvlubbRlGoF0WC4
ZHSHrWtz+mV+6JIOLcB7E4UAUCmRMuWrhJHcpQWvaMB+1uKRRMr+2xfFVbwMWIrWV5lnwy4DZPyE
zQq9Vx6+Nt7EUGPXm8cYRPc0Sv0EONCQkeEouwOx8or9xReZrRoQUIR+m0vhEL1j/6OJlEwXXyxy
D0m3wLGH1K96E9TQf6sBVT24fUUSTlvlaPokw7XfnlxyU7hkKVI77X5tnsBeOs1nA3ZF01xTLwHy
mFsocfBWS70QC5BrH6D1qejQmoy61nvYwtKijjF1AEgj35kmTrifDkoGVvfu2vTUKtfWgqlz34wn
RzAF/7mRwUKAYgWCYmiGIL/Zx+csmjoog/DPKf/BeTAXHTzclP9LUiNslBPCS/Yjik6wWh8o+bXF
X8y9j0q09ABDhrKLiWtIYOpi1lPKO/wBlwbX9iUfyx+hha+NCdaSynLaig9u80Rh6eubun8Xojtx
+8v0xtg5Ol9hpmBUTq2SlAIqqJRhItCG8DFFZ6Hzdih724OKUU2DhczU/nHy0JKQ+CMHyUuva3ua
dG7/ja7YLDhU8Fd/XVe2QiTCiPqN7PFL8lp1WAdEvSVNcnxDGo7dFerltlMyfF9eDdI+yv9UvZZe
e6ZfFdM2RFQETQvtyD61y84YgbhRdxKnnxcaGLwhWVLxFEHH8tiYzzORAjLloYgCwyzUzxueVQng
XgvDXPFQ4mT03sUPXV/2V/nK9NmrfORukUmp0PY7xh9mfV9EqMVp7Tc8JfwOEuecRjCavhMSoImb
kIwkTvszy7cXkFTnZQtn+sK5OHTtvF6VJoZ66KW6qEMe0zfbkbBd2T4JQVyQ5igV6FZ6LJq6M5h2
zbmWKt79Zo3y81K+VD5SKbQ5nVSRi3WsnJPINuUznaxktC5FhHuheXbwdKYS3fKts4uIEKwojZgV
WGUDFTh1CAITjDC2vj3PI57UvBpEcr9bbpLlImelZ8hFUaCFqf9WAemfIlvITDzLimtPfZCl3c7d
h0dK1HZrvbyridbHshJROQVUm/Vo9KCpz4MfFL77S0TxE6q4EHSpphan5uq04oYTw9B/c5uXvRaH
kV8xMC1ILAPq+zmVr2Tnkzro4gdV+PmY3KP5k5GrKv+G3+Nb+hdbajEdHXgTFEoxoWkGzdRav/VJ
8Vw/MWt2h+8PShUHDz6ZnFdmsH+BXphZdWcXbHiaMOIFLRsd1tkx+MONv0AYvYrryyI7+MDvW4D+
RLNQV/kJXzFgqEqnp4AIuGnrhlGF0BF+sB43+ckq9yJ5eT9jUtuVTFBxEf5UllzPw7jSGc4X91CF
U6qGg+h+rRhkxlK5VNsTsTrnolkXZT7c3dovRMvQiInScTVSGXdRviKFX3MovO79fx9QYkbeXj5s
Aju34PvItfqEYPJ6bRipuOYgPGg5KPBBafCbZHvgOMsobj6USRmRjNUVpL5k435dSA2z5T3xyxgi
P/uGF+XUaCUOqAYqRqBQ1x1AxpRGIDkCUSVd6cIPB9u9VsixYbtu2qqh+1hHatkbCrNcJnkWZV63
QzYOohmNz+OhOdTYzYF8PRGDM0pJrio/2+oDY0xUFRp0xQSXS6ztZuABjgrHrqZp1EScZT5sDUPT
sjR8SMcPDFISE/+k1vPlck59kC3WOCsyQgqJbFpCZ1OUoHaMpTi7ck5OGzuwaSKYgmrZvkCkk2ON
/GphZVx7pBXIB6KJWKnGxYSoGw+K+aXFGC1ZXK0Xg/in/HZpxONEGmO883iKg6XpdPrwuaUft+S+
A9XzjqCMH1iNK/7qEpKojWgHJ2YCMxFSbQgxej0uMcyt6owejZEq4XE3UhHc+la84qkN4DCPhLQt
NIlD6ht4f+Ts9maU9OGIY2S4RKGmNvSIBEFtuDEaFLfeISkYq9cCb5a0qctQuPC4kBaDAKtKTBMK
aEV/cMEed4Jy2oTGTrRKAF7AK89OuY4jCKArsJL0EeitJWpFIp9qGjlZdRDOiFTfA71+5K09zFd2
9ppsgluc2NVD+Aa3v+pENMVWyGVRXGDLOY8oG29nqPxP7yJiwV/N46svcJSSdZ1sQN7npT5SVPde
GUIhKOLoDan9HharVOtL7BHnZQ631pzYelm1KohCOamA/eve/oSR5KLKEGvSpa17aoMYJ+H9+v1v
sXhLg+zrA+P0BCKyz9zB48Tj+fZ+uIGdrhLr2Qpej081H8nR9f+rEcEtvhwOmd+z+bd3O1WTEDrE
WEzfqGFbB4pEAWPZR81pHHK0m4fvqxHU93QINcqeENPX6Z4fE0h5iG15SvYNlWGtPmPFnX8LY9/h
JpVlTMlUffVbFf91ZCCa0Ms0E1hFxzs6orjEcS52E3Gr/21pSnUWtY8P6zM1Kd9eSPtxKyiYg60m
XiQLzvQvZdAnUqzsjnalXWDJZezQMKZXxxLx0Rh8YUQdLD23SDWrUoezVWUkQfJagiMsa/2b2KfM
kzCiuojE5VIBGD28NTRbhHy1NeTcnw8oBh5eo/FeH2SvGV/BEL5teKW82Y3b+NkXyc5sY4IeK8BT
zc1ABTD+yYQck6AKWHf8UA+r4Q5xLSwgY5gKctzuP4ABd2zKbFuwIz8YrKyS9Wnd4+vBdBq5jsTK
HkAWgkXK2ab33jNor1Ps8d8hEJXCjKKXFEM02b5ecq+zeYyCV4K7OOYfolR/uBvKMTzV+MYoJ6BH
Yj7MjgV+39IOYM4ZOhRA1hcMwbVyTsLagegE4SYnf7ipY/n/p9BoPzjeH0QuDt+VOdyyfJQoTQTr
nqnpQOMzDzOmbVj5iKjtB7iFgu7e3pMgWbyZuepCgliykoCKJnrj3ERJKFkkLfMs7Bf+2qOVaVHg
Um0NeqMbWKLbgh+/hgw6atrwfosANhPBkRkeaKzwO3JG8uMlnomlnyMerkPb4by75fbNlRrlgT2S
V6TPsXNXVJonmRpANr8vLWP8oJwdXzILdGwxRjSlcr9o8VfjjP4gcoBveTYbg/RQL5jl8vKtkR5u
tH+4QCrHnXMCuCDk8TvORmFUUfHXKQC2nIpRMHod/bzx4T41Xd8UOcvmfRcHIz14IFP3Al7w/Ya7
Dd97qrKdxiquby9nqTeUvQuETMwZLUj8KRFxqbg2lcJwXCmT2d61RoG7R1WuP5VD5L3a/q4n6EBX
6jxYJqRXLb4gZjqmLHiD8DEcXnK+yI8c7Sne34YeBCpwELJgEIDpqRHkFU9m0oKKA41JV4hBnmHr
Yv7arMCIzg76LLHZ367Ff/x9O9bDqQmDGfkHvBTsrm/FzmUGJ8khC+q1hEm8xqdfVqD81sMA7TmP
uDgSrq1Cgzdav3h8JeRfgMHk+h3QPbXmPTViKZbZ5lmijW9G9NGLJpaxz2c+84Qhdl+YOWK911RD
Ltrq1pLmGE/IpTO5n/gcq/NxtrE4R2bVp4QP8/8OtKZ3BWrcRuXlJUYk+B1tuWOjlhutug8bRn0E
jkhunz1qcH0XJRN0NNMwSZRupSRVzHXbQx/Vg6DazHhHaXXUyKIwiKZ9L6cDNJQYZ1mxj0C5Ot7S
FkUP6IBlgt0CwVt8bcahds9Og1ZX0Q+1wqat15momf+/QxxaJYPbDcsaUebyedByrYmvtZc+7okq
jOMcB66fV6WGuMK+tBaPbnb7EkaxgAtDp5j8Ur/WF2DBDaTf7iAg+Oy6LYIRYW2+4OjVXQTF9y6a
jPI+lR841kVD+Ak9VSlgZBWy9etXJz/si/AC6YtIYA3NCw3MxknaPMvJ/jwOFcKDErm58hMzPuYP
wSGIUkqlfxXhp5ABQvmMuogVR5aldkruCEuaVmPX8+VPpF5sCYbDju279tnLrwIXZdQ1Bv4Nx11Q
iVOh07XR6Od5GDAw3ZGBOUu5tWHvEh6GcRpJ24RjwfhR7OQ1Z2/klgJbhHhdfFP/QQOEkdxSgSEB
XeicaOo40WQvHC8iKiTmGLm8Mu24h1CwK7RcouCN+ijlhFX2jtIdXU4xOh6QoaPYJhyl5L4KyxlR
ZqjU7gproT0iUX5900gSATP87OxVn3E1Sffe7f4PjLx8iX+P+1FTB4ymZpKeTxg5GFgJD2tv74r1
Fp7P0NuPZvSZsvsXmlSrlh6hPPMY4/JP+66YBIwGE/ZX6oVs0F/ygZ65JI8ItsHHLsfTEEhTisIS
HRs9usgR42NXq+1zMwJlLDZHy3BIdP7V2AHdfC7LgffNW1H+0zL8ot5fLwXWZMRuFqxKAB0vfNgz
HFglZATzJ9XbTAt8kZBpEwildpZnug1cBdhrWFFTYxwC/t3pWXSZwGx3c0KNljq18nw6NaJajF/8
LQbpjjVUtX/qCX5MHHgJQfs8xVMirGXmm8jIXR1jgYtRy/GRv43AB27uxbKne6E3a0VqW4g5NFKI
nwArzx+00zRu6BOjYPNes0oSO3aHzz7KS4CPduX3WneCRZ4yp6eYqzwqrjoC3+mgh7GYyNvGzPze
e5ZYa9CnYhUjnLFEo09/bLBt2bYmOnHmt33xzvIAg1AllDvgW/VRGTK0XMH6wPQ6L+vgbQGZ6qOD
d2fwATPV2+HHmRcWCWWjjGii9tlmyo4irDc6nZbsHNUQSs2Fky5dxw7RYR/zJncQ5tWsALIwd4v9
WT4zJPIZFRwi6jkWTEzcW2+t5yrK4bl3Tt1fCmjLX8Ru0/5zB0DwcnXKyPAnuNHRInyWyNUEeNTo
s/p+6iZ2UwfeiG/rvfoKbW8GHdh3N8KokV3Pl23GxXBjIFKUIKWEPtCCCJm0TvPDjHaAXZRssTJD
8BzETVK+L0Bq1clE6BQrUKdDKuPZWaRY6Jl4UQnOyg52eYV/ypXgZpoQFG/yGxU7ftLCntMrW1Nu
YD4u4jEzaAshpL57xj2nlRctBpp6lQnFVq8bNnXQQO9xUe/PaOqdnPTD3K40y7x5Sq1GuQvMwm+O
wfjeTVDctUWZPZkgxicsYnK5FNqhxf/kiO3HsjOn+2Qx6pKhovCNAoEthnbtqLFOX8508BmsIobi
Vkt+c4shhwACTa6nTPjEfV0LkmynoWWjP0nT7mP9kDyBcABaFFnprQQLVcVMAkjMAoIJTQeAE0Y/
IfASsxU7Vehiramqw2egEBcnk5/akrctggf0VsvyDi7gGYaHPkjbuTW9bfb1YIMSJI2iBkJ926UQ
zQc+bKzTkAxT31xkAP6MKuHt9UfiVLypQmR3S8VdvvvD4OCk+Ega9etULOCi/3hMQJa8X3DwWQ2P
8+ce4blByJn+VCX/Kj3SQA+eNc1Ha4wQ2OsWTK0qkEe6xO5CUUN9gMOHzaSEg+P4L9t+9YOCHqIf
8r86dQWbCxHys6McQiBH/EdGXywCZVoGLTowuT90h0npTN/2752hbO52tc0JHj/HyZUwHl9Z5X06
RsWrGwMO0ODBDZFnwe7SOQ1wnuqBvTZoTJoZW8qCiQmKTrQVt48LNg+gQRkG113CXH9x09JPqUOY
6UdUHyNQv66fUKeYXnVr96R2/JnCY7Sxjq1AFbVtdADKVmqn3TPhnk2Xh0DaeSMWystmZLqjK5xX
RQICsEqiqmcv3I8lf5TpT0S8WGSD+0Gr/y1P+aX7+qyetsuzM0Su3N1WPayTdge65TEr3PEV7NWS
7FuCdHm/wa+M1wJwFKmwCH5c0JnemkPDEWW1fT+T1jwClFIeVN3RPbP8l6fLhIk37LJWp86DSjs1
NFamRC2ylkyaTO4JFc1a+C6XEqoWxzKpjdAUM/hcE9WyLeqFeY/newE0W4OJSID0IJAl4CByOlf8
qGrAuL47E7HUQUnb6k752FL4DciCWHbU8IuhM5e8JDyIyjeogC01U+PmoHSXekVDhoJwQNEOnFQo
OjOvEYNSB2T+yCc9jZ6gdvXxfYj/UxLPZI4CQvhhkfITwZjUzU3DU1HqirDKYnDbnsHEN9xg9MLR
6AsuJF2VBNPOALDT8P7uOSqcqZDz5qwRoIfjMl3BgHhAaNdA2vxfIsYb0O8I8QDmXOIKz1drFEKZ
L65HFxb4iJH874R0T+yWtd7XHFM6A1mkU5cz9xDn0rJPIj5VBiqL1MSQGLvaaBQfzzMu+i6hPaou
dzxYURJmDC/oISbDHqo+k2g2bUFCPQmEUP3t6ExELoUSMZRmfvFb+gcWyaoQnGl/lzE4e7CNOY+7
ilc/9VEjuY7XIeBeCM3culHL5b7BAjpKgRllVHePHnSQuyPvLaBsc5XQkd9TTYO0s4VeCdYW5zHg
p8TkiyGEwC9dy6Jqj0xKLx/mQVe1Spiv6A05QovosOmFRftRiUSRLZR952Nr5zj2jp1/w7lfUe4B
ebmnXfRzZTeMOOiN0f9hxthGFCY2RUl1gFcxvxH8sJDsKsVEXyRr1doCpjdjQnYSSfbZ9SSMFjLD
FopapuRKXo2aE9DrAztoNH8RceEGwklAbJyA+lZlWXEZ3cquhKtobupNwkKQIGiphXPo+D8p8QGX
EFnB6OBUCs3bgFE1Yz2KuaAqqUzvzl67PwhU3zsgbpQZde3OSuYp5BJKG2V2jKuFza7++7/2w+No
hvD193Tc6dFsvrveqZNFEePrI9MBDyseFNRaAzeSo9peuIkvgNi6HRx+iXUj8HlI7zcNE65Gch43
9XI8jO6oJ2RMOYXKP2jpojcVOrSCepHQqtKsXjAbxxgoTNez+fmbC0p+Up3h9gyf+pOeokYZ2xSK
ubty3D/zlwEM0FQNA6SKK70d0gyDEmJZENpeBijbjZZ/Ot+5WxqlmwB87d6uxBWocBASsGwTRoh/
NSCTkRHH124OnA8v8qBFpWTpQX0Vvjfkg7bUK8OMBKyX6aylOUJlgNBb8UyghLLgxRvRGLgqH3gi
QFL0p3e7a6ZThvM9UBNO8VIyQK89lZT8vtBQ7g45wwPEoCh+OyeUemSM8NVMZ1an7wYCRoONW/GY
4Jf9CO8ArkCY1bEWpZA0xk1vQvc//ejXcqTZT8jbc1TL142RmX2SwCZNOvunaVB0CEUEBIjhu3y/
jm+qVC3kbQTPgOVrz5gTVCXs5ztQf4H2D0eIn0rVjSoi7F8mRHKVnU00DAByHHFq0i1KulpCnEOp
zeea7CnDquszaxXSxZYDJtmfL8pvZq5QGHFbKofheX/MSadn1bZ49bvWhRIsqKzH8M8uPhBymTkI
BXqKoQzpL4h91HpkiNT/jY0QgU7Xn7SkIBqvaiY/pM25p5DC3aG14HcoKMSvXVAx3W0Y04DU2qot
Cf9ZGS8dNRw+Av5wn4TQSOfaCiXk6DVufcfESPU9Phi6gLNAIGXf7BwGpF+x2Tr64E8mFx/gL+jB
RvTjmiHZotKyb7QXexiFVx+83TaYlZUwE5AWKhPhhuKNn7LFfDiYjGvHigbNcPcq6SYKgApQku1n
8LOlP2V9QdaB4BA6shArxJfhhfP8L2Nv5MfnryR0grygF2E3j8JHDajcHVd5/kSp+6HXmI+Uzzjo
meGn9XqtJXH6AApAAORNQHMJbhHB6nklfM3qJ6BZcZM1UgE8QFRkDYX4Dwu1yMJeUh/J7+h1ZQ3I
FbymwTtaVUTE6zERNXeKW8twZx6Upa6kUrHu+d/R6oPO1ONFWf/4Etm5trP8PWnVm0y70zEsqy+J
b0vnjNyWEZ3X4Lk90VnwRsQqSpRVcaZJYZJICy7dB1z4XuMwFo5ywHsBoh93ZZa/Ke81r0Y92s4r
hxK6IZkarM7MLAkjXJy12p39ThEZ4fldycas8BDHN8X5Pgo3D1RoJhxKv5C4O9ktgzI79+6c2Y8u
3DW9KvNVTDCdSFWF6uLNWxkFk0NcJPx696kelSn68Ou45rmbN+kPr6TR9U9EBcxkMKkc/5gPHq8P
FkA2G06XrcbMq0RmYmzdHkS5IShHdb0EANgBUxjNTrB/fcJhqwAiF4jaWPnKQEdScwQB21MEM8N5
TAGgZPioxRwjEpAf92P6nuYLH7nM86bLJVwMaejkDLb0PCC+axR0KeqLpkF/pNRRwA7jMbzfnCtA
uK/VuqtK8ItqjzJm/5/ibpc6E1O/9Tx3T8igscfVTtv2j/QAGjpxPAPp5BPx5YxOANXxa8rtFClJ
OUoUJP5zjt5ZkdIVgGPxm7UMJjDjTrjr/BxYs6QnE5QeYUomVz+sz2LspPavjuXKhQmyLZRd1Z/4
H97bwRiGKuUXGOYIEzKXziZ90PNQ5GrCDrr+G/sG4G1dwMkKbqjEdSzwRL8zPz2JUXz8nu4/Nq0r
ppMkkVEsBtl91erhQLUiicAiU+273GhemI1aBtJZ1NGvjFN/fN7jmPfktNMFys/YLv9AcrAm7MS4
oaSvk+czFNTsAeQQ2FESAogGlzVeWx0Rk8Ayt8udpY0xxZrIm3wvuQclk5OX2zz2/wvsOcS+JVoc
4HqwsUIt8GF9GKXEJaCXjdkYEP9IWU8bybNVwcWmHGosI8X3DzK12b8dNfF+bCZPyA7to/GVhVnS
Pyd0ypxNmvvKEbtBhHTp57jQ0D34Ef7oT7c/sA6XCHb/Zac5kuF0iQN64oDJ0EMES/tM9i9uVS6Y
O/82ibrEmU58102urAMPQZT06BHL0s4ffZAqMLXaYFaYlF3yJR31J4NQtPMAk6ZV8JIXHMDG4f1d
qHCq7JNsSrLH13D+lDIT4JnlcRwQJHynm9fBeMqZGM+c+b7I//e3WGqtEEDOe731yBJCpCWNzMx0
ylku0HEoSkMSWHPzKLA5P6Aw51Ez3JKlcpUdCpG/MYL4BKhM6Psbg5HQ+ZkTnCKUe5hFJtcLWo5d
twFSJn+Pqt1YwPYCewOgcKoju/aRrg7yVZvf7wTn4BznT60+8hv7qbX6oYMIpmAAL4Iki20IvK6o
GOSivtmtiQjdtz+xYBu6IqeIYdwxoXVsNGA6YcLPzso1gfaE7ty7rtYb8XxCylbSfqiezXPisGG4
nf74tkQ/x+OrgFa7lYvsK46j8S/4iGlgfERqbVOF5u+KZWdzypHXNCWDB07eW6k4rmr/rIep/oD8
BAg5k/XbZeBWTeaYhPDdrLwH3QxZk4MLOcb0wf6iN4OpkSU6CiFBWpn64Zdpb0D3D4n1qxXcyGgY
wKGT8DSeDv303pn2n6mfW2h8s8vxIt3B4pEYZ5sSoG1LX8tuJeYAdop6DPeoJ7Nb11ST7IcPBZLS
wTSYXdDtoW7FO+C6pGWIJ6EZGm0kbG6PbuJLyx2GDMyZNqIpR8Mxv2OoRrijApdJlCLEZ7xO96QP
u6y4RToRbQP/8B8tNYg1T5TqDm4YotTjrXg0b8J96G8rx9zb73j314hrTL6CFyhUcKrpEOJZpZ0O
bHZ2sLZusecSIoDOjo2L+A664OAFAel4JYombVZXZcjXahHkgOFzVonLCPq61qzTN+4FjKnKpEYp
9KLiobfr3RyqrD5FgaGC0QjHm59W1SgVg6rtpehwiQZcvSs69F9bNiTAPdBlMwjaSeqoVY9r7eKX
vkEcFRlnzMFcBjUZQSYHXzBcIW7zK4VHguxVp7BC9BiWgssTGbGbnYpeOmniOLzfytss/3wQiki7
idshCKREHlXIylw31bG1wxRx/EWetFJkWaUTTB6XVtozFdfaHpD8PmN4q3I9C8busKMg4RGKg5sO
jhyBAvmTKaYzELbHM+c06/uZ/H5+X+PP8dlb7aHKe4NRTChjdq99JCN1p4CBSEvA2zYjpd6G781H
2Dn4J5CRh1D7CVvoYBQfJi3zdjpgp99dccZwYa6MICQpHayZTjTjw4ceAtdPHa8c8lDj58stpZ4O
y9pFoMWUaFPwpwRgdmdoKqhAovADF34v/QJPfGfOj3pECOywHVyb1p6jdYPAe/d3OMyiZArOzuoN
/Fn1DnAJdwS7YxEy2+I9eu8/XpaLjC5DGUhb2eShdLoEmtvpcNT03X/lX/6OQu+Me3t1tbUwCEkd
8KjMfQwF47BdLQGYapY+xmQQS1kpIUBAn5syJnGVWYr7Yv4qjCJOE/yG8oK5JuJc4OFu0Jedabat
xmUmQGGVlbJSCpMV5rAEWSrTVfPgMYgKJiSBDRC9M0F5ET8WDTIEUYsZQkjmmk0tIUP8tLBU4NgW
5ghiMhdm8MHwaaB1SR44arym7vzqy0Uiws7DxVJVUOUEvLw5Ts6suy6waNU3PaKW16Xz9lrvLbgz
vvJ6PMUDSs1Kwmnw7TQcFHfy3bwPqDxtli4H/f1d/qFWHUiOX64y+51qqYhDstvigS0922mMSMfm
3+TxAiSO3GUNF7hEyxW4ZvC8wUEIFozWGxkLsFmtr0SBA7sOt/BzLINv54hbp/EnbZVcs3r6Ihfn
E0FsWjfPQ45/pGeTyILYYkuPFG1fGTT3yDizy8HvnJAtMjcYJZvy7zm1UTT/yQrBb6jcErIvK8Yj
2JE6VDDTKyU7OsLq5iJ81B5ZlYayCcf6rXQRLar/8jVyGttWngfqgpZw7ziezA1HJ8w4qcmraHQ+
kIumO4KTH4NuYSSaSl0yxbWIywZwqHowGII4KQzpcICxBT83DAPu+W/CuLrUcCfiDU2OIMQktXxD
dNTqcN+ceifSI9cJl35jRWWD/CVYzQSkFcxwAKfGTINlA2lv9SUaRjGU+BslpWopT0pZKTHZjBTL
o06FzSlVs5hVQQsPuvM+OQoxuiwsZSj8MaGNRFL+OLK75Ch0RLaILiCWiuMmTvo7v4VPj2TrA0oC
CaCEdfKGF7oOHMk8GX8r8qPxhbf9VRuJGDntknqXUv6SKeGS5dlZD4+U2XTcyaBSBJymEQVKm/Uj
w8QsPpaM0JMh+Zgqo0NTRKFA7pRgZqkD3flcrLUzXJ8dNFx7tVyjc4Na7r1z72ww8/eMuhrgrcR3
N+lxlz1zSEYW+1xzRkyy9lPXMot3QVNGBjS/fk/2Tz2vdaZscqlGDHNZ9eRToQvV0Ii8Q0SGR5dY
ZQYmHNKyEE+6AUvE4djYcL+vF2bI503TcALwGmhEFChZPorISehps+Y0CCqG0xivktOxtTdTTVvL
g+pnq5V+4rJ1Uzq3M5gE8Nnd3H/tH81mUyYbvLpCGVd5iBFXJIC0pyWA7Jhb5+55VL9MJuS4u3hy
I/3Cux0tyR5NdxHrQQyvLEHOWR5nH5hJk6PfYuPxXua/FGvm7/WVogqDtsK/coDNnlKWuePSjFYq
fPflIOrx7ztIVPIOePVqaM1f5G1c7Dp81LyKXwH1h6iSeEcuqfdmbhwvK0vfdh9XuXqi5YTDYqEp
3F/9rPsjCBP7OXDDqp+CNG2tpdBY7lJblcUCJCQSGAlqRQlHa84HgIiJrmhPVvKWwusjcxLNlLm3
IyGj75HAtI7yExOfiB9lfCNz/jqtcDE+c5Krkb69+u9RLh5afa5CxhMFvg6vz7uPopcyZsJ/DVMU
L/hKnP0a+uM6+hJtgFkKcVpkwbMwRiwy8twk+oi/6qFDGhi5XBVsv4zmNYjxBTSgtbE7dPkXNJtM
HNjtjrCO0nxVOFipgU7xa/k2owWlV9VAU+wBp4EJ8ZG3CXRbDx5rhxr9zzaQ/HAJVIbD0bywc+AL
co9bXWBfIDWWdSUu7MNmaLyq/umkCU3Bk222m+Cc5JoYZlHyb3cm17wIDUe+RpZvoQeHL4rBV+PM
jJLFMP9h9OQ6j3G/MCnVC7rAvfjI4EM+E43QgiV1rkcOPVLqtk8uWNxL36uclU6WheLVtR4E555d
C+0SCp55YH6q3g0573SG2sLXBlewq8IqR7RMuzRXrH6ggfTIVBtmQI7SGXQNiWArKAlIdNA+OJKY
4KimUAupJSdQxSg7tmV7B1G4bV9REBfMhEudkWxHTq/cQDqyWOJM31/lVI9Q7EuCwaZHQLJoBd6t
BLzJIS+j0P+gOxt2vSEFxvgAen/7dyvmYLJ4VeYwxeD1HBjwOWb20+s//ZhA3MBtpgRy2fnTb1yr
BiFjlVSsOr71W+5q3QCgY33Ikil1F6JlBsGiiHViD1HlLXyCWyKC8aahkq/FlKu7j8fVOZHWUAqR
C0BRhiJYJYgcm8bKqrdWeM9m9rXV54Bt6Q102SPEjsF8Y4GipB227c6TZ743lmCOZmWk5/P7vfbX
RJOsLk5RJoW4jifUxRfCynNuO0F2K8rk+7Q66BlKFjLpB57AJ2d3nDXDz803O7NTV+Zq5KEt72i7
/oNiEM6kGjMmLXbABor8xdqBuM6lWg3/Ryzqn3ASW+PJyf/kpsEPZxOBRHLTTFw7vxt2M3PIcikK
RZfXm0ibIEEw/HXZH0v7Fj0wDnfFmoT0PM+JII6DTZ55A2Jq0oQPbju2bPPJih4ofMwVYDWZnbd8
6BIWKF9tieqzpuYAcIbbOHTUpFxua2dQUFJmIFK4/ybnLu8thKowH7fr/upSz0v262Vw+pYqI9sC
l6zlv9K0HUJ10RmWHz/CTUxjlDydf+J4Iz6u4Z9wOUFRaT9rN7xMJJnI23IXiT+XBGO3uMnsLgDp
wuk1qPKFddXiQAbB5Soqyj3XTPFhP4hk4X0Mroaw6zoD3ObqRJuBou//LCRye0AnjkX0b8YAy7Rx
Yy7cLrU1aFKFvBPKlLzIsMRQkECaSbdLN9VEnDSDVNWHQw50w/pzf/4ao/RTFv8Kn1mCpsat9BKD
pbYaGFwnuNTbHBX92I91AM36uFzvBPOpZGw1IMUhWEB0hyvOzkSvjCGs7aK3Yyx8H5z3wuAwt1t1
vJVArHdkvJ0rYBSg4HXApBFg/4bEV732P4V4AiN27RqvNDJla4sLre/X3zpnZK2YwX2C0vEzTKwu
TBe0O97qJfbroTD3Nim8/PGPNUXdtx5Gt5SOus2uwaxDOs0O9c9uIndrOhFMHI60ajTINafQPSyZ
OmoeEz2iOPAXWedu2a9rib9MGriBt/iLzsavDDkPcCOJSfQGyZoIDFxXEVoeP5oVmd1DOfSrEX2a
4I4W3QzTX8vmiEadgHTqaPVR460ylXpuBQ5/Vw1pWgjwPUPpQxzg/NZ8Upv9YIKjCcDAG1ejaeK1
DsUdWzV+tD46wFYQXx4AdA+MyadhrNeeJlyltlPY2/Y9eHXRtna9S42Vqcws4x0BnKx7c4j/FCli
A6Ryo45y0+o/256VdvfihnMlP0uF45iN0neqQKu0qa+tKxdByd23Kes92YH+8ZX+r3fT/eGjMt1v
Xfnu0Wg1UVE0HAbZ6BH4tyoWvzSTiE2r75zzsntr4vViqoq2L7rg5Oe0eY3tgo/f92qSzQddnTno
F9dFHbBug/lH5R5kTekijvWD2DKEtqaytSGBMyfEiY6r2l0xziDY7KizhEWsz+OHY8+B+LaygolD
vT5UisouQ+NnNnFPuAjukIu+Hl1a7brrE0GDdZqDfRJU0mFT/msar7Ls4PCaPgobf/NHuTJjPNQf
4Q/UWXqtNHwNWC2f7FpZp4yl9PLki6GlLYEyt/iU924/6PmSPd2dlYp9jcX3UmtXPoGuwuVijM9x
NC422xLv1UnCo3htS6msYC2zDpzcmIqr2L+l2PNzLOo63k1pmKVI9ox4knbKB+VnJzwILoP50t9y
1+/4zNEpXbngDqbb+VjQVykrxKTw/z8zlx1SRmUNoLqsktLwmIcyKrZ6mJReD1BqlOHuls8MUB1D
jLJvkoa7BzqK3rn0rFLaji5R5azsXEajSrsEpRqfD4/RJzJdmfwYFowkveLOyKVk7pnwoR7EfpG9
IRAMbMuz9P/yQjUUa6vfy3qkR9WFp6QWbTcWO3LnOnoA0fGTlz47wrxCpIDiLNRE7KR7KgwIBPq/
FK/2EGWcHUofxqane7W1dEASK+SO9+44/K8IUyRGpDzagDToeO57YKlhsH+5Jiuma5QL9cI8aBtP
DkYNqc3wzLJc8qrN00PGh6zgoOKUy0VMc45phg+ht5chw4CfkJLlFBJXwYF0Bi9mufPIRBxYJQYW
6nJCPhRZdUiF2M2o1j5l7lph/s+mzwGOsx0TOL5UaRk5P0/ioLtCJMQa1vTJiNLmYVPuxwcUOeLT
AaDtfCXIIebmYjHSThZxfPrhcsGziKDqeF4Oa1hORW3XOX4CuBDEBNXFmirHzGYC0adUBhIYBdAE
ZHjO6+8DcPhHF9QOZ060NcjXBrXWAb5TCQgyGbXc1f5ZKqGvv5Woyb2wz1ugrK6AyGlfeSNKQ25t
GphwXNgBpm0rlnkCfaiEutfVCjWeFXfxrwMcX3eBBr1V8ZazVAum11AToButIn5tn5nRB29R450h
AKxxZ5nSRnCKxqdWUFn4EcoyixzfR2s/lVMTa+GLxL2gQ8rHNfoXEyyS7RIRG0GK4Rw5HH/iY5Tv
yNT7EPqrzOa2tBFXYs1+RoC7qwbURviRH66HLDViRrBSiQQccbafvF7iv6xK0Nh5chNoCl4DJTkp
bfjymCdXiQMWHsygTUzJYZpzr755Wr0JL39aDFAVbkpnzhYR6LRuzSMDawKKWspX5Q1srl/ofNLs
WCQDkDnNpfp42fhzOE95t5wIXhqaGgvpQFiec1Odv3oFi6tjXrmw0IKZluXT5z5koHmgEQXeDiR5
CiHqRGlkJzoHdutYId/EiK7DG9NmGT5Ba+AGaTzpctZ5cR12pn6RHFK4fV+D7hCyp2e1WQ8Hb5us
ONUoUqtePhQyngob3hFqDdZeL60KZBSICIheUr1AthPZmPEi9bcPZ/70YJ5KQD2vEaUIT0w5uay2
1em0P6evgFi0DqkGGydpgH8qbMOsCGfa75KijQYNUWTDKR0PrLkmLhDqoUfgUSrn3veE9wo8GuOC
L3DHPHDusyVyjlLCo0Yayk/yD3jms8VLewuPhjhK7OSadvJYKCbBkTSUyCgTxPwc73AGRQTriQaL
8dYWwhuy7lYH8kBXHsLIhwnsE2Yo+RcsYWFMYY4HlDTS0gM4QXaqG/6daNf2Pr/IHzwp2EAjDXIO
3Z6s5F8deV3lBzowox3bC09xwK+PHj2pr7/uZcwXST6nxcIboZQXIXx/Ci9pN+uQYvXD9XhnPspy
tVBzztjJlT2HJaMWydASLuTeGa5iLvi2zhsbqaNDNUIEMKpBbrfSgY74uWjJFO0ejMzSVagevglc
x7Or/+qFtUuVehqrLLmBbZ9HuKVUvN/AOB1N/XIjYv+PN8Ws1tdqoqgPoAiD1zHnP/1yyry7ea+3
2CqvYFWVWEZddX/3SwmGqq4v6OgEznUypV4WdpawoY4zSdN4BkNxkEBL+xY5uOinOM48LcCSZPVf
QHhqoIpcEhYLWsq9YHYozpGdjancUc/Z7FmRqkLZXnKl00AgHjywID6pJX5ctBWJt0V3IKrNzkDC
aNzdO7Vc9CFJuq3OxhNFWGLeeIA0/Y9+7zYK6MJJyghS0F64WF2pjSNvCBu2x/wBZdAAJG9DyzKJ
9SMrOG3MTscy0ZXPG0Mu2jShiOKZ8454a2bUIlyLb1KuEv+F7Wkcs0Ews5YvIHrV1Sp1NNFyGS6X
mo4NyDYvEdIAL7/UCctSdYqbg2oVrx1kMHkAbBKRuHvymyn/9WWvEAMmXoHpbaBUy+h9ARw8oQ5m
oTlF5+e8kNm4H7NAy/HEQPXuo7eo+5NXBuuabG3kdbgdB2csLPwLum7qpeWJBTuB8MNqMzW59blU
4L2yGgaw0eutMrPGmvtSSS2QZNMekiFNe5uRSXLfFOeVC1idLiTj5SS420aJeixeHbxxcL9Rg4gR
rk6afKTheo+MKeTf1R+2fTmo35E4Bg5CpQXz0UIrHJWcM6e06rR1dDvZWQpbK5EzCWt2VjX9ISfo
N1JN+CJCpi+TZ24avWFyJ2hd7j3nOEySZnRhqp+rjTstev96wKMCxs/tbenWjuY94KjNo5Btguiv
6fts/Czm6DMr/neWuP+i9OfNHpDx0+fzCCRwIr1LDrFSvd12ZgnY1AmiFJL5Fbv3dwsoWu3Sw0AK
Xei4zvCs2RE76bq1W80JlZtFHgs0p4E2tSAlDbuoSK80c5RNLbmHOz76zyb4dnt/05yh39iUYHza
KEI7G1mHoejFRmjBiDIRPeZJGZjISsPVLhhbLlk5IrZYVjd5+c5AxGTXtDoRCKbnfTJXnYrBWiH8
haXvJQHy8gAN5HhsD8T0wkQQGwk/IgMaEc4NuyW2NUE8nSCYMxZRx/8K2qWwbBk3KfItZOTrNN4y
8C4DhrtJE4vVpH9ahlxUhXgWTB0WNFAUoLcKBNJNHraZxSAz+eI6xyXr55YWQCB/QZyNt/tMLE3O
0GmU42IJg0alv8j39/6unNoj8ONTCZ4VOnB86/w0YqrcRIA+wwrsxNMPPdBD8qvEuvy5nXI476t0
dp58MHDbPCbLKcBifsnGaO92YcX9DXieUBLC3fNpeqKadRLUCdKwdgoR26ltc2qFDso6CxYcZ2O8
LRu/YtV9zBAzl05ANvEzwb+o9SDsCmpTcypv0Y374SmysX48S3U6JKMqh6+VcxOWoj587O0drSzX
qE1U7NbVfGReiLazk58XQopLxfxZ9cDXHz22B1PRiWTFSRJauce2chMsiCog7gDOTrGQtCl2mkGn
TXxcPo4AqEH/0uFLMzyfXeMIzUqpa0g4u11simxwKoHpB8OkcOZWtEaaDpxh1IH7F6jK1Rr6zk7N
gs9NnRshC8Z73UUmc9BQlmH0nYdiCVXHVFOavn0NvKUqIrE0kVoMGCKxikiBiYtj89/DB/DzPVux
YlwGR0BHBmXPGwytgxlV0Tooh94Lh9cIbHxXIKN4hvL1dGu0uOT3tb4QKMJph+e7n3iIkP8PWyPF
Qp5nE0k8xkc/0MULz3yhnojYfy+or27XqNvhaa3khxrS8IWELEmXE7nOrFxUXt/sJOxsDhZREIhs
aHlVltOnf/A5/HAx5+YFxTNFjdWF7Lpnjv1uvPUf42pIfmsEhqg055uf1RPvqms0gViPDbVsa9vq
dmUyLMRtRKdSe2NDVnjl0+TW9jj8Kb4T67HSCay9xWO6Od/eNKQl8/bSTKu3mxDqZPHV9GqBbZiy
3LQD2/sojGiaKyNooScM1Rtl2jILFXgImEbPibejBDrJulsobY1+Gc/xyBtiNpDKfnc5tuMfMlSD
HiiedFnuRtu/8N+sDh9jTSto8VId6lkZLpG75A36ksiXXbIgrP8hL7FLb7aLzpUNcURd+lE+kc/p
3j/Nq/9ROAGURjSPNJUAQDxVH+UhbIOk1twCJFr0oOLg1WCCWioYPoGYingRfa2ksVe3IKZ9Z/AN
BusiqRc7VCbSsDuOaHebtW9q8TD41pHrHmp4pZVewmDM4HICBliwX0D0qBz3KYq7N9QhJHlKjWcI
Nr71BYgRUbG1MRb9IlLsLtdK1+3eKnP+tEnkBO6x8PE4rAhycH473iup4bXK1cHx1ZINTHcLLgJj
iwp1uSBDj6SXO+nsnVCHuUQo37UKt96w+vz9OY97lxmaxMsBPpIBmVJc3guv3VffKtRasNHT9usJ
nZxbOTqL7f8R3Bs4Cv23mhx24aMawBZEDhz4Pobvr0Anddvxwz1EMQx/5evYYOoES/K9sddUH6xG
3AHcFh4apLHfL2mZ7dmWhmIf00FQlWkIXOcOaHnH+wSMzBV5AG6NuGlO5b5wY5/BJzKh33y43R4v
wKwB5estOhCRpxZ0+N3wPdgEmHx5KoKP5KR+DaxITv89R7axKcsL9AXjUDuOah6jZ0HuSzQ5N9+j
TRHIWbMFLV7NjT6xaLEcDkv0H3XXmaCrEnfuYZv7M5tAjG2hZstcVTXR81B3q+2UmRaxb8U14CZu
Ar4kQRqkIl2DrGjM4rwQXbmlGiQaoE27x1xkHYy4TBckQ8tNMy7Y4SZYlbfmMfBT3AJ72Sva/vxs
NJPlIXPLjkxhRBj8RSrgkIFp3uJKeWPfemqPyo3aBsVZsEYJcwRqlhh0rJphhmMmeZ2WjiNOTL09
lO2/DfASb56UYQZWJfu1Td6HhzmkyLo4dU+RRGrQaQPwck+Zjv1SJ0upVsasTrzCdM4EC681JUId
TkV2TN+ROy7KeL4EuTIUUEg8Mb1UevN0SDWrykuaPrgL1p0Tbja96YPrsbC9qEDNvbRMi2BfvQQq
3vQ9f7t6xqUI685hbU7H1+kR5Q1DhC806wLbVMJa+QxG/o1VPGbbye6RYYjEkNCaOKNnz9cPO7pC
XkqO6H99PQ2CoexMh1Coggwcam+5BpBkPS3mw1k/3vQqDqjYBJpmhx9LALQwDDrQSFT3qvUxqOTm
K0mkLjY37etFSFzh805wYQbgJxQWpebaFfRKyBzUpkyBcSuxmRkDyeyeMCUjmluA677QP/jarzzK
zwbWLZudvgWyjYPpEDV3lHGUH8pbPZDscamwVYYeBIlPwuifKJMv/ZjvSVu/ssXK1f6fdESO1BS1
99DngLiyJpnSVsBaTLRaVBXnrTr+5RW9qnDE2R5jjWyQhEMiFPObe5EP4N1y2dTAqjzHtP4EZ/Iv
QY+3f0myB2vTT/JsP4vuMgL35Ql06klg1YScdfo3g86q1lH62lHVt92WGIEBxiUufXeBVSoFhD+K
ZrNtkmW8ErpHv5cD8iiCcJcZ0CvZBcVgS3K1MN1Hlqc8xx6aDKZH6VtTDOkAhqwoCJ+8gCEs/Rv3
QDckCSBwL5MlHZQ7r9ABqN43Wjs1citrYD9kORMkS9KsJ2qtUgCZWkkGY6GGl/XXBftTYe0KzNkw
utd/vZXuITbvpRlRYikHDfAFVAZrTgH2z+vm4grS6/SYJyN4uNyJlYgtjIrCqM+Xz6neYmfdE5xh
UvCZnauQzLKzFoaHbjwo3zx1CCdCO0puOcC3eiRcLFSBD8VukSdW1L0jQowGlhuipzvR6YqaV9rN
ed7dWfvJy+KoFmLYUqRpw5F6enjZlrtRGcBJ4zIXb5z7tXqol4LxR2QPaBA+k7j4lHBPEw0LlsMx
LLHJ1d/1OWMFXcesOgusUimfSaqOEH4AIYqCrtwUrEbipcLKoxSHpjlp8RALhKl8NnyZuvoWoHgk
vH9PLk6dq1viu7Pi2bZCwcIRFFxxH266O3wn+pHx6RqAdI282bY2IYGsduLVmoyOuq95NqlOVtHp
DIPZqqtKGtdM7og6E1J2Af+P7TZl6grC8W9T/BU3jJ3Cqlc+/TL/D7l2uYobUAbvoj5mK3MWCXF7
cKsY8+FWYiULfZFDHx82K4OJs0PPT+CDCBVtOtiFGRAQpQ/tlN4i3f9SFY44knPHpkVV+5DLqwFe
7FWkn2FwdeWmJ2Y8zXyJJr2ewqStQExnLdULXPnzxQjL1ANZbzwg1o0E7w6d9a77/mQI+goHl2iL
RmWqFrdZNbh8AA19ZnLl41pWq/ay/Nuv0ECyD/MPjpWhS2LsQQBXETz/X/vNcyzc5vA6YqU2Uw2h
drKj4rLEwSd8oNPRyvyG+VmN+wbskC7dVkqEaMuKzJBx7dCVhaUQ/8Gf7wSgrXqBbpBZdfCiYTGi
iQPhMk8tHnr5yZesyT9gZfQ11DhueZpbfxnTP9Kh5AD3PN3e45m8gwCaKk8tx210CBsCex5iT6rb
yRL4ASqiZGLcKXsSAw2U5e1LdJvKFwoRKQc6XnONOwAkK282xwoxTAjMurJeGYB7reoU96FP3kv3
IwK/DrnrfYgVbAnYEI8D1bor3mb7Qq1zk6hfAQqbrew2zasaqSOwm3gx5rvqXd7+vLP3JIYVQzIq
OKK4Fc4uGYz3dXg1caQdjRpPYvy8T1K066s+PrpWSL8xdKTFWDf9NesUarNZ7kgOM5+RxTe7j57Q
WHRl5e5fTWlJ2m4SJjqlFHy6faVGoIUPPgRT5dmsTAuDsOIdjXnoBhb4YNkLEuF2Y++ldAb9+Hqt
o1aCFmIjcvndwNShJUP+3ahrssPRoYKgmDMl4RJkehpqRg8ui612Qlqq1fuKun8Am0qBn0py/M6y
1u0+yfJXKO/yo4ou5TvDZQ+NR/rRLCWdPyCko4+QLNKfzYclQ5MXU0BhpuwwHgUASEDrwrDlpua1
cDaX4c9a5NAIi9OVPsawDemPQbkCsPFZfKlk//sArmxVa9rguhyxHNzy/d4PnTptbO+uSWXqaUIk
vgGVkzMRQsyZOe9jQPKEdkYX9ZoJv9uRyXASF2kUmEfy1cU0AcRCN/wfMi1Ekwq1Qc57oSBDm0es
AJl5nZInWviMQaZupWlZiUL2Qv6EIubo8PEs/87owL8Ai0Pj6FCxF0XbZXjL4IqPgq7+q3+q5xED
NEiYLKQalGLNnfOSHPJljZ+EBjEVVgX0IzouJINlH4u3fGZRkGpzDeZGXc5nT5t6qRb2gjKkVMWH
r3YktCNaHFzR1E84BXvaU3HkncJQXVok7z6ZfqbtTe/biBB4aGB8ZZyj/JwBz8ejj2YNJKgPty9Z
zwkvGWNt+lILIGiWcMdhJdeVGluhle5JCGxg5Wcvmr6I24wuPPcu3/kUj2fXmIeNUMDSxfS5RmJJ
oGyhfgf/aaxYZDTApk7TvB3awEaLbmktl1x18hAjL9OIpZn2JFv+W+2PyCTGYe6TAXwzKDzw1IAp
39BhSeFgDTjLcJy221J9pgJP1VXLE2ZbIMCeI/3EgYDnftPWTx/qAPJedr91LHiOnzRzyc8vB/n7
bHa48MJMj2pAyzeAH93Hy+vz4lAp/s1hkjyE9/cT2jyAKKJDDcM7ezr88aHPtuhwIHciFY8c/6X8
tBrW/7qTtjA8q41hSBZ9BYpoNr1XkPESeW2I/oBz0DYvoD/I5sQLOprMCloZ36I/z3Ii6vdPA9Oe
PRxqbum3+ko24U7pRDCZzqgeyi6EVHafAmZ/iy3EJ21XSxI9CcNpS6zzYBOyGuySIWEfHgcVmnHG
UYwpOy7HSLtlfWr3jOfuarmyTJKSrXZQokwnLxAz6D9EkMI+ktBRxLdn6AXuB5OLxP/B+ENjvObr
mJocB7BCpCAkYCbG94ROW4XtPEeCs8w8HDw3CA3fBNPRXmbND3MkIjeoXqo1X+jGCFgNSON5nIzr
J/LpJHPT4pnWyr+4HQ4nAOCtCP0POXEdSb5EtRRGnDWOojuIqzvv2Iyzl/f+YVMYv65RU/Hpz6uC
Zkj9RY3Fl0thKXqVx/lM0VWhDIgjC6nn80uLkxwmZpafNInzxH8b52oKPHmtPd0tf1bG7ehPsoAA
k0SxxIrRFPf1V+MEN5Z1KAjfW39Gb3fji6MAYgdXoNZWRw8Uvuowcc/uQ8xasrziv2LPLP4pZ3Ay
it8ZV0Is5X/eARGxXC608etXFjJDDGt2DkZl1bl4NCy2XUc5UZpLS/n1dThzpeSSrsrBj8mNxI3e
lfEKn5WlXNzHHkKErQsLFQpunJoT4wwAdZwvH6oCch8autVIMDDVuE+7dzoD8mE/lP+Q1aTX72WC
UXGdWv+ertF3v6ZCXkmqZ807jhvfsArK9pA+O9PopcGowiF+0FH0Apzao4SUHjRoHzwAnhxmvsF8
phWufNKi9YVbonPx47KCAXSh588vMR4IcxSfLPw03hIFmr20OK/gHS4gNzlo6rxNKm6JY/ZUV0XI
qVwistbhzYSSRpg8cehVnL/L44e/k/svRgafHlaKQiYaPRcDjpzCT7czSan9z4VNlIq3HOev7Ndb
BRBFB/20tdFA63RyTCN0Sp3GIPy4wgKADcafowXTu9EZvi8wB9ugsJWdLZ/am0c01vCfWgdLsJ38
VeAY7Eu7Y0DGhWVtKd70ya3A+pil11J1AMFG3GtKLmeH4wITs2XJa/8EhBU5RkUOVP1WVS/Lkk0h
kaXet75jgO2vPFWyDHfxdMKCI7VgDl41zTJxT6ZyWWW8SCs7lAIwfvMkNVyqp7c/GyZlpt1bpSih
SuHyANU1sbQKYW8Lnf0hiSPbz883uea+PV9Tn+6Lf65zNSTkNLCfsuVQHmdtpZmlrEbp60ZddTTt
FnU76zJMNkb+Ez5BFE/hPxRWMk/gQxiqyyDD50EnzOcLqYucEXl2Gen8cEYhlkBSC2X/UfHKlXbl
mb96jcAS+1f9wUcFFHqDUCQKK7Dzc3muKIXbfPFzODV1rgoh7b3s4ns1rmdQn3DyGWyigvc67MBH
ie89vexxvHDrusWMdMNNDZM6UdL+T6TVrOiY77UM6waU63Gysqq00bSzMPIC3u2k8e9Gw48HOSFF
1IpXR77QmaDctxOSIbpC3fPb8jop3NqhPFLj6gc5TgxHeocbUxgmEBD7ctZxoaS2CTktv1uxP00K
x9C++VRhmqGphOy2RRqnQqxoGjTHZiKsEY/eiB1BAtLCukEmQ/LGws063lGBtFl8lnz11MLeePcJ
AieembMFvF3ozBDL0wcoTnCoykslMIQk7MvcCqaIWzXYqApou/8jmUZlpftOFnaBXrVu7jEFpb28
4vGa0zTPAv05q6PjdRGGMOLjA8ZBPMGnnvjJ4DRHvdmEDX6q7aZGEkOE4OPrQu1rsAam1dJn0sgu
Gb1p7geIuKpKKuBQQev7SUTtAoOawqFwTVB0tRV3KFYdvyYssjOt5Y466vvxsCyJ0vZ0LRHxXJ1T
+bXAL9K9Uo8+XLs2DxtoS7feXun2d4BPNQm9hg5yg+mTyBmNYXE90uqNygdXFN9uuwioA2fsP1g4
6P0vi0obHSFUWilxh4F161HE3fsSJowhVeISMWf7yhVNltEJtz5fsI0iQb2g2uuCkyY6MWMt1vf8
j6iuBNyKjsKBGDv69pu0fSkqMdP+fbXIy8UMZ4Un9YyQgLvVRNO6Z+XFWYQHVWr68w0Dp+K97bq5
LOqK/pSl6U2MLP7c1LEBFpYKnRRuVMcUMxZqAfv6RokP/vSjqBqv2WsfV3PLF690Ywpp58cJdUbj
XwGIBoM6JgFGOGx5UXY/Hbghd+uYdOS7mit4eNNyvYcO1wcm7Fzkp534vdMwskqlWz+fl9eJk5bO
sD9LlxcGV/WDL/fSCHOkULCUScsPdIkkwvzX9O9RJWIqa0u5m0hC6PQrACZ/p1Iw6pQu1o31Ji5i
kNRlxhDI7t3LZsXIbFPLmnfA7deNkCgZnAymWjkTRdOAy8C64HYEIXHpzmS8brWWLWeY5nlFj2UF
dGJfBxN1aUvhXvaqynhTwTqpdJ2AWXIVINA3l8Vj+gNc4VE1c+HZTvOWRG4b3frqX09jqFfVxfRx
ZK04Zawa2SqFbluq77A6DrATgb7AgavbFAIhsAZg29sk9Au6GpwGFnl4DjAPuow83PqT4U8ZNGli
apyw+USuL15z3jjeIIPrkByG8l5+eWoKylXjSaIEWFbAG5mS2gMPPcg04/C5suq1JXi6TmMdAzAe
BTdumIMhPuKLnDj36oruAoQ87k5HilENJJHRuc2JAvREEY8g6YfbHgBXCMiqZ/+TPumuOeV4MR/V
jA0ZetAeOLVkL/6Z2Ox2oCa/DlJs+rEP3zab2Uuc4BP84dzn1rxMx5TWumX3RogiU5lDwBwlDOy8
YuHykzFtFjF54XRGNJ8tFAZGXEgRgt9rdNj0E8giRiBOGu/8QEETJ8Usu5qXEyUn3ZVxHfs/VIQQ
wrcWdu1Fjouq8qjBbU3bgSXuJXsz1ygbkNnk5i0gUz8rGuhEff++2643ymA4fSgSy3WXcq5UynrD
1t0+flGkARJxmlgrZr0ECXppYSp4aS1noPKs97BYn6y4ubxxxYJz3wHVIXzXIgwoX1+mfzBQb8kZ
cwanHaodt95Ruaqm3lXj7Kob8pyGg05al8uT5Owmbhdx/0Ds2FyapP9Jf+Ea8zbXLwsd1cn/tbZo
tQRSCQduL2pbRta6ZbhJL1ILSQT6vulDzcuE0Ia9h8MN46Ad/6H5HHlN/qflzbGbV/llW/gLQLUR
g1vqx1zB2N3f7WihZtKvhQrzyxbUPi+HtOxp3l+q+xFDouFMZn26IvYAsw3an9brK0+E9m7E1TfW
f7uji7Ns99Zq6AhRsIeNSu7nx+xRuvdXUYuaGEZH/OY+jgYiXsnxzaSnKHUMiHl/EVE2JHTKhQHz
9AlrJewVh3cCqvxR9YkhtZ87v60llLoeAmKD5MUI3CK/gpnlvUloClCq+6sq4IcVA1AWJJoc9LDZ
w0H+CNJYo0pC9MwuWqSuMPrVYsJZEOuAUVdhI8d18wrSJm+WTla/G0XUMAyvtBPeNK2waev1Dppk
3iUE2CoIvL2TwIDeUf7ZDmMvzTEAG4jzY6HBngMZGJTljAXeHaWzufZt6IBQykaT3BExvfkQrkch
yy87t3Aye0QOKo+RcPlLZ7KfdG1lT8aP2UqoiyrvlrsmZWiLkKWcIix4R3J8HkI8ezSg8ClJbydO
gGvH58zT61RNG2OocSiBZDSjMgZ2foJ/Xn/6fG3B37dkKCBD7ugXr/VAnDbGYb9JrD27uonyo/nM
LymX2UpO+c0SsXx3/Smwj38B5vHEhWK8ojDk6yFicvkTcjEkl6/a5bYB/pSIMZn5uHbVKa7TiIlY
/7eOHjzjii7el8iTW7ipYQ38tlMRkSJ1qPsq1MCqKXY3RlyIQ+ozj8YYfnCTxRIL2/nkmADnsMdt
6XJVt7XoTytQhQwqByPQZizerVPA0U6MItsuOmYxX7QEPCAoo/KAUR2GqN+aQ2RRbb28nDWq4Jcf
jR2YC40JxMYb6kVJbSeJwAQrwObPLkeGgLJptMhJlDn/TcyAaydW8BKSxKCjw+ML1dogQ3qFc+pW
F6ChvftYHvavqHXgBuTlk5D8pTxaBPl6UnhK1z1PX/AsJzegnNoisjABNyOceTWKuJthB9Yw5VYK
D/DoVcqpSDutfxFVF62zc959eHCoyhZ4Jt23V3DjIeCHnMLdJaq/nZYQzIYc+0Ipmw1HqH/hVRxQ
fqymh2sD6PLoPicvxupK2yQc/Y3Sqd+x8ZCdys5RMmnTN3Z6rcmsHcAWmkOZjuRPj/BkIw2lF7oO
mzdbq2QC56+Pf2kL7geigHuSoBHBmutwTx6nD6I5DConCli819NlgXK5P+nz6uzLZdwG/Zm3+5k8
KhWTYVmHWt6v5MgbsBfGavPaTBU2PMr/E/BVtu8zPNvvjL/IMhJU8/v+Op33XSOOtELK63+Xup7T
+vniYw3ApicK7rnVtsD1GCxbCYeUeLOa3MLsAoBNOIRohX+cGdqYJFA3VeuU8FC9/RFfiC6LbnJd
TmWpjOwnDxNV8fHnAYKMHnrfOAcS8cbv86IiuYpWEgUU2Wjhr2trImfffoiMIbXrppJbl77x54uo
ZYR2wzGKtiFZl9FJsp5qqDoUjHElAD12uTKRXj0X2EDqrwKEfENfGjiMt/XwrVhCB/tRkjN7JPZ9
4ZCh+Zsgv5T6Ns/wRvdTDSJhc9XyC6T96FuIzKbf6gSEn/SR26fhc3ZkKNkmrrhUovWFbfq9Sobu
MCZksTmQPvuvR6V1DUxW/GVl4Ao+qDcRHMUKjaAqAYj0TKTlzWvvcbZo60K1ERiB+V4/0HrlzhUA
WZWCn00ip6lY46sVevx3qUKt2e9GlmTl525/YL98qO45RoGyDGC+vkRBbvAdp2D3SKPqFXe7EjQD
yjXGYQatbiYnIqSjx2DWMRrKdb9ebnFUpx8eSQOzfdc8w+9xigX68Wp3SWBIgbVRNn/U9Exhw6ev
zmk4Z/C7gIPS668rd0mcgXoyRlXS6qTBssf6SxyfLSAaQgzcxqXXlw6ZZAGGN9F93RdesKNbHaOp
igAYTesv8THoPBOQlVC6BE1c1xInL0qsYAlS1wyMFCE0jES71UJKpQlQxPcNOmVlKHX3oemiS5i/
IjiwKUhud8ybvlQQkzZXW0YTmHsCYNehp5RHnFzhMRhac6ZkM5t6iTE/5f223v28UmJWgdZdZFie
e6AsCTvsggemp0183/5aPh3n5gR1rvQEorIfnxwG987vGIjBIuoRcLuChLRlHrFLye8Ix2g39IlM
t0yN9UMCOsVSuOWXbRLwjESvCxsuLjLTEeYDb1FbpZbXd6fgJETcYKjbI2OEruTDIlASGEel5FgN
zDnmD3oKGn7aQspy1Pu4bWPi/cNFWAtw8zSUEDJhgV1y6QrdInJCHwBHt8Tc6gAy8xltDtQmmpYd
ea3++RdJQuuV4pRdH3vfhz9Jzvq+7DY5PwxmbP2ZqX3qjbUCKG0dVV1IRRQuVY/ThsWVzO7CIs80
wPmGMAeclbW09IofxYXZWzFxK8FUosEdRjuyOwifnCrC1J9wdzZVpESShJJzfxa3SfSjvS0vLhRM
iYWMPZ6Ys0PE+L+6PDcvRah7b393p2mhDZZYpAPVEuTQe16byYnlYKt8uDO8XS/muPmRGwZzF4nj
OEfyq9Ze/+EHBe5q6uWIBHT1ia/88zyVvn0HfyHO95W3dJAKyzUFUoaIMJW1FVqAZFXicgM7Hm5z
gbx/6aTUQ0+BPc/IdqHUBg+BVJWnN58iKqFxwPv0SXRDQPXjqmbphoIhT55L3uBuUjSMnpVCNFlW
mLwoESv0hoTFMRIsgMAKGOIvOHR1O1v3/IGXDfSQyov4yP/pS2pKjelc96R6YfUzDsOZqEcpHP9z
t2I9hF5f9hTiKYnZ4J12kMfZDDsRRWAOaPKB6OjCshS4uDUAic5kp50SfpKVn0Dw1Drz0L4qJ0kS
qhvAL0ftRGFr2vYewB3OyF+e1KzCH6ZJeeVeUZdLxy5s/cDnvBbtsOz2wp9xWfa5tdN9JNzhb7sF
QEKOv5UTqg/FauVL6zZeuOew7f5w1ja9ExQx/dl53DI+6f6KRn3Ws00tkXfXZBKu8cugPBiU4MiP
khwWxc7ty7zgSbip0IXq9EE34HQMvz8zElFFzx1ozMZBBBr2MR/68RuHzi8VCXBGYOi6a6iddGM8
wLBcB/wpN9l0Cf7px30sjbCqfSGnih0BgS14ZUmLVesqtwJhBv9LMRg/b41+Pt8uwEgMwS78ujCl
OM6s2aRFm1oKE557lEab04o7O7yaDA8jC3wUHjnmGNjMphX6kZFoMPXKFRoU4WcvakT7O22naOdN
j/UaEd9J9GhHQWqAeU4OJLTFTtQJtxAuRyFdgoiAZdU0wNFeyc349A9nD/IAeZShppJjdy6nvKlX
SQRhpAhufHj5vplHh7/wCQ2CLT4qB+oNu+BtHQE4J3BXlnLd+Syq90dsfZJH3679pK37DOiAYrsr
dKZMFI75JfDMVwbQRZoyhYUTZnNDHcyBeAWHJrVOyPhJ4squoq29Nk3ajHI+nOEbzd7Y1iyWRk8R
o5sOx0JoDTiRxK+XmdfB/QJwP/NGJElyaSJ8+Lj7rkZYmbDxu9CA0GhpzGg97vXuabARjPjOZ02N
l/nPHmvwnst1wyC1D6TwWafOTovuhpDRZlm3UgRbDDAppUZT3qNufVziqsr2CtXVCoduAHTNh+Ld
+n7RlrR4Mts/yIwEdqLZTM7VB1SGwAyffkubkAImr2r6vFoOPb0N5BzjN+anzNTesb074QzIVt6w
75T+R9Bj9hDgVWmnXWgX4G6tkoBTVF8xbT029Dzn0aX6DPf+XuPcMxue98q7M1W0xuomJ7aIt9Rd
PtmF36EeL/GTNFA2TgkDX4znQ9NhpdKA5yfoVANQ8TDVdq0r2hM4PS/Zc0xzjxIBFQgNtEiumPVN
kts2gEOCSvs1IhlnJqLuy34+Cx8kHbDQMIIpzFGvYTrwl0Vb5eD2+NdloZgsON3tbRKB0ZHQlayv
d0mewuMJQn24kEkDeezDOxqxauI8ejKePyMFOGI/mD9D2Fbne60Tp3s7av52VILwABmF9yt33BbQ
k0m2WBxtYJjARGeAzXaBJ5Gz07cfTI3dYUNFuE7yHHc8CaZ3ZPjItsVkIY0F7jnLYT5rKyeiOsG/
zIjEIW1L/qhKSLN4G138jxGf8aoRReDw3ktVdA/3fVi4laGwrSAf5ECr0tXzgmRfRnQJFPGmWwqb
KlqdD+O71TdpqBC8iVHGRSmbelbcp4aBbJgceoaPx71P944Sl5ILG/WA5ca6PTmQ7mHwNsIZwQiH
UkIqWDTcF43f2nydXjBTdEg0GFBpdEFPe2j7H1ynEW16wOpKEfArC1K64Kizsy7i1RN7mDPtePww
y0Wv7pJ5kSE7OZdhBjw7IHCu3zBNZ6A0Z9q1EZxCCJzo4JYeZ+rlZT2b93um9SjVF3CmFWrPkpBs
j9a4No1eNHB/ZgaU5mwILxSFC/tMjoT1Uq4dAMLvaN2BgY5km5IeKcPumwzwMLROgPrYUZdBzJB2
P5biBFeIpW+J0SWe23hjyR1owik6DeiQKfTNFZeHnihG6z/UdynVThRimp73g9pQ3kOcglECK3IE
eGWsRfM0GaCDDKhb8PEsZpV9oSTAWwmJSauwMLUrG2v9L/6sQEjXQiT9g5sOytK250byKV4S8D8T
vwp0Nc3kX8i6+ZjHhtdIXdelMCuSn7wRBZhVF5hDAhysXZjXghSUEUuUmOFy22gAjf2nc2nWkrdW
idq02/wksFvCuP3IjvevBfYqYuZ8s36m7eyB9lOci9H7CjkYCjqL+S9IDDR2uHmftLEkIr5JkfKg
kK7ZrBr8PAGAPOpZa7pttqKwwo62P0USC8lRnxILVzRE+lfeIlwDyKCcLIcpMbtK12kISzxEKAwx
gY/2rM2dDm1SPE/x91zGNA49xW6DN/gV6bsNb1TY2teeB0LkGpVO+M5OJNJx8/yfgaKCUr4/E1hM
wTM+ovCHg48ykYXCqLFFraHDDxfbVDmMlbiKc1r5wL4AhdNQIRcFgp2ynkc0bsYy9F8F+ua7YYc+
gULuuOhdE1K7ltP7VGND9W1hPKwD/rwcdXt6s7ehypZjM3XDB7tc5ARZf5P2h0ke2qAia45wwCUU
zPHxeWHe2z9la8QrIhVQRLikJiOW8VHQ7WO/s5zNQtafXfE/+naSZT5/tqA8uhNe7xyms9AvfD7u
lvx14ySqNF+zntSJS8H8avUB0TuKmod8QeX7+deUKK3mBmuMlKKKNXE/tYzE0CPiZ3KD5aaPLutv
9o+uIz8o7veEt23dcw8qVbboGwb7ayOe769CvORot9KThPq5+3jiV2PS0HokCUDgAXkM9QE0t981
gUum4AvnzRV0PyX8ddwQbwrC3RQ7fCobFgNk6aHM6uCOoJITxBhJPkR8/PE+CHZdUJlA6B6UlhYc
P4FpZZCZfCPds/W/HDuGSRvFaKH8+cGRUPSfL/MpyLjdDM8eRH8VdkcujJbJE1qZFHaj3TMVwlz+
8QBWV21DjYpa94c0rf+4fhbIy0CVjLAvk2hcwll6uyilDezZu7kAA8GfpZGu88kKqFAaIWK9gT7E
+NKWP91xG/S28g4SpI4ZUguRMIBaZfURfju37/F5I66KwpwcP+CiTNzyhjlBK+vLKWAramWMley6
nqlJLdCX+6b06UTrBWELpDnStisKlDIZqueFJDFiMAu6yuWsLukq/xeMiB5hh6Ew42gpibM5ABq1
gmhcdEdXmbuEta1VepmfahNVDK5jDUiOEn4E/WcDXf//dMay+ivBfvmRmrN/eQXxdH8rKyW1d/TY
V0zMkAPJ5/5jI02a3vcdYaCbLrtHynjS9dKEQUN/itp7aVwFmiX2zaFXE0gpm51bLkoPCll4oYUR
E1o2hoicbUA15KLmS31/5coFT/ECwMOp3bYXM5LzLCTY0GkiAlPn7oU7VnQiTsyC0sMZ7WiV+fXc
CPURxcVqOgjoPjvJXwhR0rytIcUKoHsv17e0LUymz3wZq76jykAq5ZAMehI9OymPFAzfPJ8s9m8R
sdr3bhncjndGH/FdhjFijWP5PIyrrrATeeZGb5RO/WpsEJFd4d2ZDF5SncNigvwLdixaWyR89JVG
8LGePp6e9kI+OIVgDjTIL1c23Mkl1VnED04YZ9cPAMZeeTY5NTYqZp+swkUHW4O4jjXcFtvXcHhk
I3cr/8/45J0+2vP7rTge410wmTkb/Je6fLqQSEX9S/8wqnrh8WTy4TMjf167sMSnxq1NjSAOkR56
CR0W0oof8KzKzUD31Un+PVUwOkPqPs2N0hjYVtuaqjKAmGrZAHJAZvaVXRMV1doKqZJZ+kE7F7c5
cXHD751y2z9RS9PHuX6GnxBNpSNZ3hbF4KuC+LyAmdnFfOwCmjM8T7dduc6K3AU/L5XR7PBUccGt
qvgvYKHfbFRsPUA+kBlwtCGVXjCX/xAG+tqb5KF7JRzzpCMpMxdyGf7iy1Sa2t3pUhJlaxGjVjwl
muW1XgRktbRxBwyDdukiKW00lxeF+ImucQntsWZGPn1kKl15+4f+toCsKV46aIVmeAdHuVqMW5iR
ktLWKHFxYbY9gSjTS5fgzRHoMKoXHKb89hiu+xzjdcY8ZUoqFKqoMpC8KvMY7U8ktZ9SQrYnSTWv
KuFpTBkdOiOI4RG/t+IvGyCmAIbshcfbpfMkzvszypfP6EFUbDh8Dv00Gb0cJ+559Znevgod33sS
uITiFBEBluLzAh+xH45pyFDY9B+seTCiQbGllbOxJr1tFUphjVO670Ic2Qr0yNCy4KVqEzWc5u6H
FLAjpAE81mJb8vtMi4xUcVLocm0JPbmiimzOxUEVv8delav5vxsFqYYC/N2vS/Iy65GO5Ow0zDMa
c7QvlZ1eTwYnFRK3dvz/1HakV4bdQhw13r2mafqpaNISOqwfX2N6QE/c6NNzAqMN6vL6fWJEnTzo
Bo0bsRoeDGYpeZc2Smx66vKOU3cDaWMBaB1yxJYnD2cMdUyiFcYg/37tR72iMcLfvglyIzGRaggl
cwgcTpIeoLfOuncG3d9hxlltGn4ocXNHz7g4ihNtDWrE5odpr+Py21KtmPDYPQwvfFIFznOClCtU
ABB84Ju99NO8uYDDoLnXlxxRZ9B+Hi5xEM/3gtnWe50RJG/m399CtZfGJmkOxRcmPpl/I4Ni+3eA
6MFsMTslZEA1cLIEc260lJfe3+OUjwJFu06cfnCzthp95MgyAQYffQg0saJnad32tawA4kj4qbFf
sNyzsTGQ+tMOyznJMe5FXufVsBM7DVU4jmHKtxqheQtYc52XZB8VtOHnvv2vc8zwzKGX8DfaAG8B
UXetUwSJUQwZFWbJgOljkK3wlC5B8SY/uiO0cDHMGKZFjXeJF4Y8MKwdMPLBKCrQ6SZcLVLoHs9k
TXwWusNUU9OnDy58m91IoQimposHrkDLsO1yiSm4zjUIJ53AZV+NknSvZvgrLbZs5F2N0z5eMeHJ
V9YkJDCroXDtwtnISQUgVD2sLQXdtj/ceTvA8yw+84YPrZpD8VyyUsaxRgkMjByXDHs81AGrtL1o
2YxcQszFqlfPXDLee0hhVIRVfSAIgogmCrzcO9dybAfHYLg4arBdokuNiACcNB1iiW4fQPqStelO
t78t5kpywNbWkYMP1zTxswdM4PdPNn0BXcwiVRffWPuarFEo+zakU8/UBv5+5HSQMapEvqyUZqe2
grDrr+dm6G8174cXKESL32Ewq/f8aO0x07yqfJ934nXcqxtRsYzJa1Q8NtMqL1lrubCeoQdFGjNR
Ku83eRyam+X9BODvmtYCIM5XbcVr9ZXoMa7N9W3JOljNeRFlWpOv6PDqgTqJ1qaFMlGf/pph3Nl5
ggvFV5FkKc393ATBaVTY2pDdiZBKo9T4021Ilqodkp6O41dIHkMYvtBvZCQtgOWFOvlQnT6W4g3R
7wJljMfz0rg77Ds+3x7ljVecOQqLPN2hxd/ngMeQhCxilOh8HU1Zrsq9z51TUY3/kEIaHZc02TRQ
3f1ayB+s7GgiOp1eQHcWzKyp5sIo/YmZ2KNoNb+aaAjKz8t4/5g0YtL3QtHQbs2IJqmKZkPq1LxX
U0ZukWpVIFPrJ+x2UotNtsmgcZP+40ySMGXQ9eISPtEUb27/o2LwIjNCsdaiRGPH2jDRDbHH8+wq
cd/prtLPZQSRNugfNKWUNX5HWd+NDyNdOALG0ruZLPIn/lys2u1v/thYJ0llLqerwnZdZek2QJxK
1crU6sI3ABWrrnklEm5FgqzGiYdJMKf48JneJ6geqR5XO1+6hdcJ0udcppdF59hmsy2zcHH8FVcC
0clK41nlYn5sleYhg6gLvSug0ueAc4KUJVN2q5E7jjnV+NyuCCY9LnIZOfnz1QTKwCIvtT16iTrK
0SxLmpSVPhlwg4K9LtAvZIgglZHmVhXG0XSYriwsCvdC6wc/nB0ZeOYxh/NOEGbYnM7GUlgWI1rI
NDcaHjFqAm6N9qDLenMrBN5OsSiz/ZU2fXeQzCzBUAUPQCHvFAhBXqbRA1sDRg8O31xZSHbtWUZx
RoXcpagj7u3Ms4nXq+0z3J5eyyyUzkZeBDWocU7tBjTg0GH9eezT1gM9Zzfe8GY6O0pxHO6NWVR3
Xd/fxrNHSshi6z6UlwjFfgh14X+fitER0dJki6O35zkrPAB2UlKhkycNGVogBazlHX3o3Zd1cjyM
ntWQshmZ5NMCfXzirM+DnTT9p2dny24n0onJBQEbV2gVGNdTE8KefeyDJFZlXpFWmk5v29tViojB
u3wL3HB/W0LOnELtEEpfz1S+/5YSLxo4q7E/B0XnMPZkD6F4yMXa/k+Jw8PebWNLKw4SPn8Hicwt
qy45+6ugpthgJwEHiyxp2QmATaHbDVkAHvr/+EtFBhLQTx/qaNQ+Z5wl4+VikzNyeMbIch/NheJ1
d4Q3n3hSy6URcAN847lPOsYhkNPtclTl/4rW15sXjMx6bLx/RUJupg2I0IDaK3iDDyLlcjQ0ds/n
RxVYmUk5nKA32xFEBtebJDlcAl9QfNyMmI3ChYKTuH7LPy2WA+0wT6sAjAv1aQhu1pDVHo6D26O/
3axfY1R6sWxdk8Mk87MJTPjhw42icm5gWnZc2bC27Ka4upiO6fr5xPGRJiW8mmUL+Ug0jc59ngxi
Ln0m/kuQQQV4p9YSdwkiRn5esOd7QVrOmvNr/kXKIuuhIA7nEwuxPshE7Ox0MQFfl7mf3yguFOjr
jxtIr+EKwzX5ZK0kVNyCW9KGNkM9+QeG7i02UnXuJd4F/kBdFaQhiYsIzfKRXK+XmArpkSmdZalI
0bg0NGeIVVPaZrVUFp3zN3hadmDZj17j20eaH8Qjw1Mrz8HTMMLCNjHFiL5uHBguxpJznyfTHkRX
eT8+ww5KGs/NiYzU2oftlRnQ+BRp/QkmdmYajOg2kYsAEl/pzdKbz/lDGIwl2lB3UmcpBjQmvSNh
9WU9WorLp2l4vdjZu+7sqctTCLsEGKjEzt0Sx7s+9DfUVPrX/TDWaY/Z0acuqGaJ2cgJWKZd01vi
HPer/v5kPZt4Gw3BPi2/sAtP6uh81fHdkwMoVhFYQv7nIvbgwjsI0QY2RRVyZMW3RLlxP9B1ytN8
Awdsd2pBbfTnS0+rYT9soeCXDmujemh6fCxs8WZZddkhvis07XoLdHW9gLNxlu4386pzpq0GFinR
+tWoIUYwce1kUAOSGATlZMgphDd0dfmIcy6x9PqGNztYXqU2AMq6c4BCrcJBjAYGYK7mZzy9msq9
mCSFOyNzcwXyeTTIY68XubY8TE2I26En8wdepbJDzBam+hGWMDJUCbraM+/tjOwg6Gmr6jTAPZS7
eegWWoWxJwulcujjzyq2MoBn0FCwlAw6L02sSQDOX7n0oeuOgZUzZ7JhoKv+WqYvI+nz/IcJmF89
Vun8vzcHU+c3CeOBGhY8DFnP/ZRqrqeA6sf6hbJzaUALtmFw64EGEQXTdMXj1HJqborueGtcBW1Y
V7nG8FHKGyYoDuaVo7ziagIWv8ok6YiQhLVv+p3DGhwvFclmq8YpjsbqiLC7f31QsW5VAmO/Oh5R
nDtHlAJaSTplK4EFRLWsPjQpT8lMby8awpfz2TAqVzJe9Wi1peygBlZvpane4xoJwkbm12vreq55
J00hf2sTWXo2nqBZ7QiEW6BlEiXYbOdnrZa0uN5Sbw47YfQLA7nuzk1pUhyJmg9uB2MqiX0G7AMD
zZFkCWBfGfLxxTnz7NEfHxOzt6DO+VpZFoNxsKG2XYsNff4gUI97BloCSsWHYSplmDNB7+uo+lGY
CTD4cLU/wfesfTnoCctU2qrQWxZieHFYQSxwNatveZ/igT6DEMltkKLkyQh/Le2lKCKNsVDYX0Tk
bNXniSDgsAimHSZm+x6hCz9FhFMNxtxHxRkxz2ldvRepVTtII1lzIACl0kysRuEajs70GsAtBFhi
ex8JxDIWqFx49EABgsJv0js3oOfpkKRvt+QKx+ZykIS/CTsZpbw7ToFiv1ImMf0UKYeO9O5sfu0u
siMRdQjrmoe+KhvGKznbSkAK8YrMHv0U6nY88veQ0ndswaEuGJl3vV4InKPxIaJmwX0IT8DTk1ML
8knn7w85WlfJtfMo8RBGI/sSKyvzDh7pMqn28lJ6NMZgCFZauXY+sM4m1jDyXviQdpSqo6Zu6wdC
RmfIDFQuwwyytENrMGpeZ9y8zxpLlVMc4QB3y5H0LGMopkXkOmpnRKjQwvUfGP3hi3WCJ3Cn2Ypi
OnRvWfhBQANvquybzL81UfrXzFG3yrlfQkqc++Ob0xWUYqQbt+ztYTPgNXRiGLZCF8f1hnjlKRHg
oUWN4wqk8K+YJ5xcoh6meXIpeCuJJy/BPevjsZfo8x8f5tIPOiidrH0MtYXJtLH7jROjnGkMMuA3
fQkBD0tamVcLx3Y843bWeE38b81m5ZojDGe0l0WT5Gwl0nJKuAjEZsGO+3Su4oLVT82zV3UmMf1T
ypdta8Y8hw5ABgjA7WbRO+wTGCiL7VaMGPbUTyyqGevgWboyxK6ChI991LKO6X1eOSD/cfVef3x6
4VLOrgdA0lcDQBCRGR3ppn4+8ADIeNCrtGvafpIOyI+O8WXMN7kAbcxU0YvGY97ae2Baz0unV5nZ
Sjfbnfeii09vAh5PyQ8B5ifTj6ssn74A1HLR5MKllKf7V+WM9tBqiMSXe+zhaXL5fEeEB4rlfddi
OiJmwU0pH1iZ3ZGepEhcZX+ddR2GO721f2DzftYhzV2MRHnD7OOJM7u/iW1gQtqw3Ct33USMGPI5
RBba4++N0QcMzM7MLwOeygWxHTh95DgQWvUDoE1+OYFAuWz6+Tt5F/96DN+Q+sJEtkImc6C93oUM
A9ZFptz5Dtdou+tFIGWfj0jr0b83YdF6fKEmtVtz4L6JKdB8CPf5zCpvfXUVMxswOByCaIAmiLVa
rQYHHc3onuUkomvEbYqJsqKjWtC04OERjj6SuPCoaXxGUmzigJkP3NNzZ211bK2rQgNdcULY/sLq
KVrQWZKrRm7nI+tLshb+n1vIP1JBLx6hbLVDEk2+c5Lo0/rbubW9RxBPb3u/OgHwiYV9v1vVw+Ky
hrUHc3Of/oqIh1FLLTghGt9ILajIUTKYXb51yz8wpfkvGVN9RSb2NdOEmJhoABp1AXLhB/lduLiy
lhSpY/yeIruVv8C9/ds3FGSEQhH56D99iuz6T1o3rEXAG9eyQ/nPhK07pSRQ4SX50pLOzSx/mR6y
hM43s+CxSMZQ+bvGIpK6ncw+fakDLhgXs6aeTStJvnC+Lfx7eQpmjIf3AVs644wZUfBALJdGag9Y
wLdFp5xFO1eaYmERjhbn93/TvZ27uOJ3XmwdtL/UyNstcTkQ0ZwZB3oeoquEp5AOpwA82r5CtDr5
MYoyhPrUFpBwHd+RT/eiUJC0iZIafgm9mfHwAOqID3K7ulI8uNSGuWYZBLuD7m+b0Y28r9GX/n/K
hdKSQc4ma2HI4HMB6l0VVswI3kv53MHY7+IAyhwz9zi5YjFifC+z9B/kl85MdRcjPeIKIt1XZr+T
tMD8juBuIjTntbweiimsHI0/b0y0DU+iXvvHj8Os4iUQY6Rw83SKijShdxi5Pwkny6dWxH2H0Gzt
H+EHurM5dVcG063SlWMQsSerN3Zqoml0CObwAlAb4vi2wjw34fIt2NWXhlZy6n0irF6et/oMB7eQ
1YeN5JVwjySdl7RnKgJpEVRJoP+0t/msQzpviCQgngz95OxKNof/jZr/5rI1GjNVMF5NoeENPCkX
e4bZx6/9B1D5zaAaHBbz85Mqa5lyrthO49y0vUSXltX8z5EnUmSJLicbV5ngn3p9VbrHuw1IRlje
ebgNeVSg5EjH4crTmXZ1DN+n9wT3dJGCKKrxZO+LaGuU44v0j17fei63ajRZuQ26L1ND86ODYmT0
Cr4kCXGtfEGfGeJ3+FSinvTmHiPzywQu/lZy9YPn2f2ijWBH/b0WetrGS1yvKx3zRW0CQ2JGU2Yv
1uPVjx/Gvm4qYYX1q5wfn4+j17oTrWm/gsx+LXvQ5vplIxxI9wfbyut8j6tbxpxPRayuEKlTJP5Z
TAG6YcvRlYDIxDjIXjhyO8FGf92oHtKpeEZzKOrK9/97Qibzl2efbUSu6vEn8/0I/P9tI2FYSgdg
NKftflg4Pv4wbUV3dYLF9c7QSxLdBTN+sT+iNj2KovJoiK98bSfjqW3np6f6aZZhKADPDXJ/Gl9J
JXreO4H2eLHmbAI/AmkdHIOJXhnpH54/ESBq0Yub34cUhDrvUUNGDaa1T43bwYJiLQz5dJaReqG+
iQoueijhySxGtaZ6/tnxpFt92yQlJ2B32TwrfKZ+0mjqk78WiYrlqCX+jzI6tvMtyongNflrInuU
Eng2ywZ21S0VfKacFZGCLoE2O+2ZSXxm0gy/RpQ2ODYGJu4iPz/M2M4xFnsGgv+BvGO4nCHp305u
7H5vvDj6FVIRHejoHjkzzd8DbqtC53RGX0x458Tkca8vs/l4Rt3+S6+cRBK+XF3kHckyAghAXk3R
omYJOjUgwQKi2NMggvfhpqQLwgIdQ+0hWoMmgb+Xy2Sx4OnHDTOjgf/1QPrIJa+tmCSYX3zH8gY6
CmLXB+M3hOVcmlBze68ljz7RTx77NXOpcHfKM5M4TO16ZQi9pJF97j5UKRUIjW3yY5pbPwajqgfG
i3LZb3RWHcNAFyTBQRt847Z1u3/nDVEGPXGcMX6nHbJx0iv7yNg/dyWBwdgsKs4FVtAioW/zDZsu
6AvauVhbm9BhGv5ja6vmX+iMnGu3Lz+Xv6DzbVMhH4RYhXQxL95z900p5x8o5IHZTsxXaGf1L18C
GBasnVisxP87EE/tFfGtPT5i756P/+xLLAfyzH03ikMivkrk8URZBMXpA7BaldjkNWlvRGyq3lp/
kiv0xyWuLgV6JR4XdrMyKRxUkrZtpHP+d+UmhqQG5pY0c1TZY3vnaCs8jGP9vBdf6/D9W+wbv4BB
T6gRpnx0lqLqx0IcdBlaJDQQ7CZXc1SkiEJddKzwtup/p/VZctyqigsZCwW8iPGlDpoI6+ecHziH
i2jqcBDF5oqa6Pa/bs+eiqCxyQgQRVOzLkJLwVWeVR2u+9i4M5fdndgFSMsfGn01nwjCu6HnXo1a
jVf0oicAFpw5JnsED29BA7qiXKaeDXNvzovZ74274izKQ2ujxnuCiFGZARHyCSbGHN1zO+eVjrrt
dyTnYIhaU27iD9yZwDrSbCioENg+dDsPUr/BAACjz0Fv5QZHVy0l20qG6RJuUpB0M8OhBAN5IARw
12EaG9VEwRwAcKC7TaojZjdJtpXLCh0YOIYCzSYbgTUTS8iXzkPpknsFkf/v/RUiviI2toeiMTFM
qO/oA87LDflLpC4aWb+IoygVrRIW2gTATe1mwfa06caUjT0XUIf5CfPGa3IQJil8nR5dew334oie
jHXO5QbxqnI8JqyLLEAW6YhgGKs0NX8ov7UE7JzA+G+WeZLPVtoh+ZefO94SmhwiGNZ5FXjbuvpU
56JXfkRxj/UartqFiY71oF6mJFw1fTpfT2V75RBWXnAzxtNXI2WgW04akX739FVxWjTAzcFG4HBo
5HKiuWBYiWkL0G4X1q9FIdOvLe6IPEP5wPRlgHtRZ8xE0ysf1pClQqtR9HIWKMZ2M1JZhKccqngK
cLJ8E69BZ357z7RLRp0MBicAhDsnOVX7yPokZRMYRgeKEE+/GM17yZ9fN4T7exEpWj2ZE3/2qrSA
6dNJADrQrjN7LrrSOPVaiPcNG0Jfcc4NqYKxldnFCNjWI/GP88H1E8a/8FtQLnIbIxdHx2ZxEClM
e8SnzizdgOpv4AS0xqKLhrqPPjW+lqKEHe3J9AufEx/n3ncYYaARZH4HOeRsebizW48SwvDkm04V
ZTy7axMY9c8MXPq00XXs/o6TV1I+iXcRlQfEiWrRXxtigbEtpiXiRsy6w2VpI8BzapKc403R0O/g
hI8IvvbdFz+KHYxO+vJCn7EPi8plyCkZMCLdOqQu9KNevqBuxtoEyctKF5W+TojnUKkc+Yyr/6Zj
6OHOpwds3R4v+tjQQxivnH+v0SxkPTaGwgKlfe4i1dyBE6+5BpE6LrGp3k7+4g3aabsV7G0edn/W
kKWnkfJum4tOgIn0CUtHn4nUIsuo4SBFnVSWElavkrQWag4WOVOAN1qWfPLZvxLXKdhBra7W97Ug
BgNMExQObBblqpWW4OgXZWhoDia0h+Vzix3Al3dS0xGTouU1Hui0qRpYRm+Q5jHNuIM3XOrl84Wd
NQFFqPydcClZ2k7t/TgpCtOCicPOhrQ6W7cKP7ZoBdlyd0QxtamNpmHsXzP34enZJ2P5dRkmPCes
abV141/EhU0LFTc+TYRCkBdtCrQHBMhazv779PMxTst9KboAoK1jVAvYiRLaaZCzWacszXcIYvX5
IPr5yvkVG+2tRMMubHAh6E+7dKLzoWQDwXpdx626AlI8wcKUx5xqhEsUspkev23bUVhsgkOPrwIh
VY/1qxv6FfOxeRBQUmCkOEQDCD6JODMNmNN9DNdG5pMd5na7vhGVR8Jj6CayxlAVciqnK7BmaXMg
gB5Q1E79ywoqZ9kfuBzmotjRU+/7iLeTIqHWKn90KmaD4tZJ7OhEWdBteyZ+QWJafAob03L8ahyy
qpaA7xDP6mw9W/EDOW3mH4E02PA16QftQDksIBa6JjItACClU//hlkX9RBH/38AnRzLj+Q9rFxCW
fG/gkvNaK7zUui3v54MDotPMLJ8RIJba9sW2fTEgmcymkgdSDqgfLzTgZPLgZTdn/7qJE0x5ihY2
/GiHpGNmNTnF83yxhGO3gWoGM1WRMXVjgprX7Meed2F1e04xYOQ6tsmwxTHj9bLGuTkRGXZ4+wXD
nUO+rYY0LKW8coKHTzUonVYqg/jkAG8dUz0NDs92AvdKJiu6imx8PQNMdgS8z/urYCYiBtlKtl26
sWwHcZSMq3YRRcBZ0fHHVjm9Wa2uCz/InhAYlgNENTK315Wl3kNykjSRs18baYFR6EreoJMMzo9Y
WR4kn7n6TKtd4Tsz0uhNprhRQhAzqvBupo/Nk2fYV1lUN+0pZWP5Vehgzfv0D0qg6jK49VHkcxxq
7srCqf2TPPJUjU1uRCUFxIIiOV6f8sKjDdkuKnPe3QOw4SkOtAz/YSBgKQm6IPDFTr9DVdkrQOZK
ezd2JRfwQv63qXsTkMVzUlF+C3ai8KGO8T3THaaRah+MoknzDRSEgN7VLwWJAqfWHfdLnprxHGxk
B+BIQKNzBMLAyJPUaEx6+RToNn72/eZhE9r0OWe/KTOsVZm5yns5pBoDVrZ8ot120sI1X3qIbKcU
ZKQh4zOdYB+PeU/9HWoz5LO1x+GpCNvGFgN3A84P2Xn356KN7x5J8+dinDJ1yi2R5YJQq0D23tVD
xvLGCLjOK2t2lh/89yyOwPacpLzU/SWHbpmEISNihG3gpBSVG0L/sWA97q9VJxabhMKLo7yLripM
dkQCYRc1Ew/q8DXRPZiudhV6PMbtLTzleCAAN4OZpJy0mSg94RSXpMV0ogNcpn880mvWxOFff2IK
WgaFU9cBFHJoQ/g1R4jzsC0c5M/spVyyqgeuaB7/jUd8r9BWdTMvv7M5Fw7xLuZ5qOFqBb5dMTyx
cd0GKxNaWG8zsGz7RluvETG3q/ZimVzC7OA4CWjPalE/zpCQOhlNYAaBHraHdMEGmlZciTNRggi2
OV638PWlH8FPzDXCqgZLHtSEtVmtOinGEcjOExxEeRoZGiBvoC2erGs+7LUAKeSsr9iwzw1/zkS1
SRBVLIkMl5Y6JFsg5dCooYJ/BkuxUQU12qQaHHS4FgBOiWcwxTybSq481lvdeNwYxl7qPDPOwFuI
fF7ZkRjGA/84bC2djDdToUcdaHjzWcDOnSgMlv7fDrgf1RimNQiEqX0HD/M+h+ukFd6dJh24UgdN
wP+aL3KK3svxEeVsyuIJ7BihAQRR6GZp+p2uLRPnzuXtHxvCjf3yjkIHi58XwIFsv9cfMGjxdyFL
Snvtgv2GBJc1ivIYoscP4kMN42ifVzgIBADW6PZ7Cg6e8RAsh0QcjtOOotVh6Rnq/eWuEnFgRGvf
qZuDkAhW5p5CpdjBDyKcROIh0Wy58SAYve+asNIaoFpNdjx/XwvhjjnINB8ugKPn/uRf2kIJH909
9p46rNqOScL/+4W5ymj9qeD4THdPgKBT1MwfUAjpQKoCSKMFleXr5RwiEumaxEeskjOG0ma1xBUB
g2H0FclN1rQ+DdurrNo0wGxKmhULwNCM3yyZ1alDcCnsukRoiZfl8NoHxYMj2wfF0tLuV+orEzZ+
x+okdb/mmzu2hvJf9nGS7GD2kzk3OGPDeqhj0qCvDCIsrcz8dHjWvYQZpyB3ayEoCYcOx+pRQs31
RzBTNLaPrC8lD6pRQ2jhZl53Zz6Yv2lvNpidM5A1qyB81ZNwQ9RTErzaxGEWYwpJI/ouF1Y677W5
ymxIXVDB4MYIb8uYWhyqFozR1C8p2Qii+IrfWEDy7uslTj36uDvLGMLZfDc/kSZBR8HaX1cPQjxi
ThNOrEZARiJx39Gopt7vk/qxL5/73tfCe9WpnM2ayTrjSCq889SieXgrD+NVaKYWNhQiw3PUSviE
MFS/r2vRvVBDMg82Z5KUlWXJ1HQrJMpEBGfbnmjHphl5i5dmuKTq2c2DxJelZEH3UkIT5WCCkIPa
/VX7t1SU4yP1cIFi6g9LX8lrqmxkEtZszGxIY7LgUoHEmsMymgKKBx/tsOBaARbVZk7D2j0Lv2dD
NxaWqCX0qurQ9v6giOXLlGC5YTlq15dBlhsmemU8t17LzogWOjoIUhtms2E7kAVrnFil0zvEG0uE
xD8JwqqqtiST3DtPAEoEhtbhRQKiC3ossXcka8IUNcn/VxKI2JVDo5YHPucO8u51eiWXEMdpyk/W
4VbXwXL+XKTezGeBzqW5ZpAMnzHx/YSFIrBKvu22PB78uOedUYbm57C/lRpr9AcOXVdFytXVCIJV
7xkyxn2M38cmgbiknsIDLt4w1iDOuBeQ6oWv1CWbWcqHld/ItOJ2Yz0kJ/yfrLVwWjy082gqqbIj
v6ijKpcr4p4kbmvqrS2XLsAIBbDjNjtQip7jOgRTkvDscVHa8d74X4nyKfH7LxbCAdtoEtd8Xlzp
ny9ZnzXKC/RvUFNxThDsDyrPpe5w3WqNvN6SwEQjNOLjgxczT5HsNFHeRPtFj1pTXHE5wcUkfGVk
iIdi5ZPHOordv2J+k4vnj3V57z8wDE4OSqxw6UVUXK9wILyhnN3TT/R1z13ABr4b4f6E2PiEp/Hy
sphElLWSsQD/3r+Bb6qyAkKpkh01Ye0g180sQuv8/f18QVAatJy4KJ5zu0zXbQwHfb4N/h8DZwz0
mQ9l1OcEhapgZk2mV5KmErIH2TUISegX9R06kuEqv8lSxpoDvPwoa7Baee/Aih0JBZTgtyQnrybM
gn1hfW6WUckXZo5EV7uUlbyqkx6IkarCbWrRG0N+5nCyWPzsMF6bnHCfOrzGPQRNULGKoNxM9Ttc
A0axvpXVsvTV0KNwcIHd2kEJqrbtmJZI2h4ZpTxAIZSLZM3xLuwF1HdzIZN+/9MclI8nIE96puD0
BpVVO1x9bPX+7eCVmMuhtcJR8VULcB+MSKL/Icp3XblO16b/OwFddaqKDzV/ovsrFeaVhUoHaZNk
w/ah380U3BNDXX4Qyee+yZNYQDYzsWdkQMQaV8bVxYEHZdtKnbJuNnyioDgxg1tX3/MtMXT0vPJx
/lok0dePOLNqGQr5lem6Ry2droyVMpK/3NYZgNsxUBI1M6SEkpMMXMkAU6Z5dOpkOPS494JG14/R
C+q0YkQ1jZJHTgfl4FZool/J1W/Th6xBCK/RlRK7jyYny2YmDIEGc5Yj2nsMNJGTxAAcBQSXK/or
MmSulhK0/IO91UfWYIAlpBqLjBXOWSf58If66y7xpJQzhsqo0dHWd+6azZUi7DbtkMwZXta9oqH1
4ZO1mQByp5wo8NmhD0UaB9Cffueg2MaEIiE6071BLv+I98Axj55hbY4DYBhc3KebymUqn6hNP2c4
Ux6xvX88C+8MSu3rf+38gsW+nCXx/0swKxnJ3Pd3a1rDXqpafwFiibJ0Gq56mumwW8ow8znBeqzI
xHLFaSwgMnx2N4ynGBs5bSL7Wg9RKmCjk1UzW3+CCMVkuHA06G89OD7boVHUe1+0qBdRQwrMtuFP
Suvi2+iAl9XwWhY3+6Qy+QbvEpajCsGP9e8CMUCKTamM2OxyznGf/r6Lt70dVG4NONHmIFKUYtp0
QSyRcB9Gjj4OCBmJtcXhaQyvN/LQCcXzet9sWD/RGKBBitQoF72gPICInr5aZ1ogaI577oBAQmDH
p6wJ+OznhXNbISmRNtsGDKOKEVB4oPfjL3zpEu+CR+umUThXHf4KZ/e49gt3FEIejs/FzhLao/bj
DCfwqSlV+odKK67d3ohvfVt0KX0xSJYF09A5hkICecjW12PmvUhzum+nJFiYhsaUPRS3xSmOcah1
kbGgzB3MgGrChtoFZPG3+gFS/RLulJMGEu3b0iIHlP5YZpTyYDJH/JKVW0yY4mpSzL51HVWsMWwz
CU6IIJF88cOyxSZYD4y3hWIEytKduHeuPsAigLKe4TI+Qt6JU/jV0m8/zbTMBqyIe3lPyXCy6Ewv
cOsH9lZWcZ9OWq5Ko0uIVOP8tgcbaVppWn0Iy9jqYb4VdQCchbJ0Bl/4HyUQQJW93PyMOUVOQ+DI
t6mMirBuTO60lIqfipY5y7XSQMyxz+hypaGmwZxRVwKDULz4jQnS4Q+05FTZ9cxtBy3aFzWfds67
d+TA4LqXLqAlAHFz1pytye1sgLslMUrZnmc2TwYxja/d0LBNkGVo0FYYXM5tlq0iqn7Xwou0GeRG
cFkq4qrfVRfDmr8p3QlGW9ac7byLMHQPvNZBFw0uU+E4Vz2Iskbm3Z6nmg8uXn29kEHC043UI51G
rMsYeAV4z4VRFkH/vSppoij3lDHOTKhfaUwd0f/V3YAfCZai4RKJitt+/tyYCltCVEtEfZmgdcjw
GlEEi5YMxbJLPRwQWbgjYV1ZQJ5ZWPkABSR3wn60DlWBLXuUAksQ73CuFvnoXKkCUmSaSfEa8Eze
hv28sIXcT3+h14co0kyTjdJcucgGJHeXM0QUFgTdBet0AvpGYEzlZRNvP9oE+jiLQJ/kg/Ddk2BF
StRkMcQIjpbAAMPRqa5iD/oWzIqSHsvYctkxdbZDpe/h0zJHpW6EUGQEP9HKV6eg7u9OZ/oDsRgX
ranaGoCEsqZYr6XE6av1zh/BZMaVROub8i7rsVw4/l8C74iexXuBOvEKhnFCOCDLBqWM/gqn+zKn
zQJP14IohemSN7QNmPpRv1hzy6xH9mGn2SxsocZnvm5mhLbK6dtevPYyWdb7tXCf7uCAwdtthI2z
/vTZk8VjAJwlf37JlMM0uc1e3Ms15vSTMcKs8z/ban0+Dkkaq+iuQ2A7MVZnCEtFhbmO4bA/EQxI
KYP4CJwwlFxzajqYl8NL4qZKfL7NRqroup49mJjsyvHTQM1zUedezpPesfyaVKAKfpxMeYaESQWK
MJDO9Rj4cMx6vbUlmLPItKUMc4NNZDXmKRapJFVdyRLH2DiqlBNc/DX0tY69RQexIYdjb9JZZoU6
4/uU0drJG1R8nexA6KWCRXGC+bRtghMOuQJdrtnw4OnB78XyJmLdXS5vTGFiJRIB3fGab4X6TJcE
zQdt0Bs1Z0XNiVGUbmTJ1zXi4NmylPqXAJ1JPjtLwgoBCaauTZlEM6BdqbHapO52WyETf3lMrwzg
l56774nGUkOwRosAcUAJXafPt+X0UevpvZKqyhvpkjuNTiAe1cTysz4IWYgJ3s4SfnU/HzrOx4Rn
PCNjl+wuVQdGbw85WXXDnBDosydD5gstfSXz5/Z13eE2UK9HW6NwZjpmpboZiffaV6v+wPW2ed6x
pkCVuVLI89Ulz2/sKrRh1Wkxxu+GDGB06GKjsG3FQVDATMVBsdZcSETOjfwJBN+OxoVWQmI4brs8
H0QjeViorzQ0GlEUiIPBbcOsH5HokPoG48SZOS89N4yPTlyAM7/mKb+Ub0wsI3Rh7bhnNJh25fEi
Yii8+AuMlMJyWJWXgAXW88bTH8Nu74t9VnrY1lF28orjnGt/ZOYGzperOFi9SBfvWkY+KpLxsTbv
C1fl3iNd+yuRhrgEzQ+K6RGJQxtscpS9UfNSwPyUMlLjBsfrS3LAaNEmsYoaYlgjHfAf4/FpQdaM
pplvc28PcQx7Duo6ujxJKwpus40htRy7a/dRcxGIb8yaGRDC35yZk3f1GfdTRYS7I3M1bsJxmj8T
SazR9fQh0Ooh1+2NFaYcf6laaevKS8ocGnoa+68t0RcaEJQJIFw6vAShmoWO4dtOJ4MtgpDk1BmI
J3TrNfIQaadMbbe7htr1D0PBXiQ5rMdoClSU1Ioc1Xs8RGiDFr1zn05eAjrBP6nwr1X+1DSIKeuq
9Y7ufFCKftBuDKNidU/VFudzmmvp2Bk/+g/5GFLSqGQLB4/2Ds9fl/UiRHfZXx8hKrAg+muVDBHD
GBUIKFO0eqpb0VaJc4/tXAPGnVQr8Tey5jxcgM3rd0XacEkuuId0S50MtU3zPq2XGSPah17ERWph
MBR5yGGhKQoeULSkBTG93SQxHpH3tnT0nqI0cJgXC2DdLmUDPkSAHspLojVVgCwoGvqa842K/T/o
GRbO6G/DqnVejKfURo/XUGNvUDngl6/Pi/MyAGHzE7NsScCJ/MNc2aDbSR8gt2KTCoicBNOIGWyU
MAJBKZ9erFxdmSVfK/y6Y8NbCzl642WMYoF5odvwqReGyPXU3H/LbhVXXr1RbhAML8fkqReq9liH
O/ZmVChT18wt4j4L9OodESM55nq+gKTX2mvORRHfstd5rL9RgLD+t9ZL6j1HoMt5ZX6zVKJGiXLw
E6+vMc+XHMhkCALXaDSGjLAI4YPDABHJpnTQwOuURGEPzc5mUPKjMYpRWp3AzLwBcqALTSmQNS0D
Y0CwyIXpXfxMhbFQcBdXtKIRq7TYOYf5g0wrKfC3va2UIZLyfxLSn4c57BiByJ5M14yRayU3870B
zx1GbKZW3KS5ZrGXjOxGQDmWqDAOlrc98UboN9K6S7OcRMirAZyrWtdi00dN8IYNksiM/TfCMccN
bnsDOumwmiaN/umuj/ndHaT2qt6JFyAYbi76E0aDx8s/kbxu91kzTX8ahkKb2EtiRj/UwA2ManKO
LdThqC2qnOqh2lZV7vkruukhZwgPquzdg5p+M/2LtUVj9SgdvKf3xzET1hWWUeonpUMAwF4/veDE
INMOvnkQJAowxuO7+W3k6MhxjwRQcVFbyn9c4d5vF1ChDZGFAGwFkDf/9O28dCWg8UD54b2wuFns
pvZfInxz0jKmaVy79vOP0a6BPNBc+seTFrCezr4fkl23HH+h6NcwouMBKi5FggnzNKVn5IfuAkKp
6x5kyY9GitbnLnZn7l6nzj9gKQnki6yyDMHwYbaYz0Pt8KWLjnJ9OW5QF8cxlsycFafiY4fgz4qp
mX0O6moOmOnZrsFQ4Gm06Rflv/F3mGmKgedcyI5uY/YdzdtZTA0wwqyDpY/sXc+aled9f84EJL43
f7Xfgqjo3XOtZsoC4Zv8pF1APInRIBSfoybZMopxYacP7o0tY0dzu0FiBi69+EQ1+0NhmfW8UGhx
XhrpDTM2DMZKtqT+PGbpV0/OHzjigNvFM2RUmHzbhQhn38BkDsDXFoPn0/QX2aUFXnpeKdP6N/wL
yeYFUmnkGYKunLieeVEThKRp6dXm6z7Nyak4AjleZGdh4Cc6DG2Xwyt2PEm9Z8pUk+qzjVqsG6ei
70mkq+x7xcNMJLuHEeN73JeOYB6hCxkw0NrWM8WmfEAXsqI4HPA0T2mK+6RPJxgn4FgFHbKVYjEq
swrKMj5FJUIo7u5qoix7Yp2qqz3Xfpe3KpNQYDJKMncy6/YK86aayu6Rr8iqWpnF4HRVG2JB3wS3
ppMswZrfuy/+Qn2egxW6V3en7ixuRT+YhzK0WWdbnmaM7YOMNQFH495MIUcSJgX2yftB4yGDOOwg
p202ngEpjhBOmcOdfsM4Za9TD0qEHwsMPAI1ILi3fZ2THMq1m+AH+Z88VPTSzHlreQV5uosZF8t6
mkgikdAkzBwof+VEv8kUaokdeJenpyFYnjA77x6PcZ4h9dJWy3V6eqPj8+gF8J1Vp/cI0gOfO7Vp
0gAX8ol3ZDc802rfFhtuwqb9//hE4LXEhZNqNmYp+Ur16m3b369tYMIQdUOlbHTWtUKr2Z929atg
fXegTZMlnJ7Jial6cE+hSFEuODqw6lddOkEG7IdPJOELqm9lZe5Jy76QMQ1MYbTZw2LLnOfXjG6C
AyrYnFgAHRd7dSaXXV/F86DWXPiAcsjZs3/Te3GCFabW+sha59JDrEkCyIQ6u7MzOLShm8A35DVb
XvXj/GmMGgPLYOgkZ0P17bcORnJ84vEBsZXQ8xAFoXakzqYfeN8Te5jN/JedO/xWU48WAG7xffVV
WEzul4zDLnTow7OjdOU7u4W+KP3KxeLlMIa2c4W0/0S7UsVZfTDQ/BEiwpvQXHPHTypjFDDFbJXf
9vgNczAq7YgHy/5LUs0XTQmRYDHcarAcOZ4TGt0HxX6HnO5/N2lrh/MiPclphShMXP5TV9RHshwq
brBsRfq1X1HSB1C1Prk+7BIldmz01Gxs0PrvAYVIgsbuqusuF8GnDU21DaDXIQA+EQAnI1mkWxOf
6IjEI5FPKQ588PW4YTqkXqJUEGof+CsVF3SStzrNjJnfzAd7wxof+ClYE/yvk0evbKNh8KSE/inw
Q6ZZl7M8PhbC61LzMIRk3NOk8Zponz/TFqyGM44i+AdWG6FKkhMPuUKyLB46AwtIC7ba8Xa2MplE
nzKdGVldIozr368yWH0St6iCm3znkEOfKzLWfXk6eEERvRy4mdH5rMZYZdMelwsRvehZavormS1T
ELYRJ7SLPo/zujy1m5r5LTCr9DQP9oBnvxQ5lKJ/9Q8sd2xiY1T3hbrnR6YHo14oOCfmAviURwgN
cSzTBF3LMZ2jZzphGmb48dZ/WU/BJciyMjIffN/Lh9R9xzBgV5HvUkL3BA99YInKfZ6dOCOzLJHy
n68y0KG8e3BtGP42MyIt+jrZUNnWLpGA1yyKlLN9slmCcPyg3q5sIC0u7Sb4ewFaWcoC7TImb0LS
cYROuc/zEYON4EOQC1SvmVW7Sks89RkII2Hj5HJRC9YZlFuWIUWzo4gKm4RL3PqvE5VFxk2+q6gk
OvJteRD65/t69EuHl/w+8tWIF3LtNFqqM9hQ1J+qlNWCh2IHlmWk5mkcB/DVm3YSy1O06s6OKX2J
BoqoGD0ThMBHUbV7MbjHPHpVm7MClpZqPBEknIPSsniGdnLqBP+p5HFowW0+6e7BnrF3lJg0qpz2
b2LW2bVHs9zIjriV9RXQSaGprNccJPWaq8YmW7OL0u3kExP9haTbwVag5ObxWsvlZw6/OtP9xzlI
Mft3ZcIsJL2uCBAdfNKA2mscRLexpOR9h43XQsFFk7e4Q9jllq9+8oKYTN++3cKAskxEBqVEr/pB
5ZjBc4W4CciC0lguF83R5IYiK8QPlvQ6N/6DoH8sAqMommxhUs1odS6vLB3hPTO8ivn6u/kB9GZ9
hMhRVGSO2Gfoyg2Ibl74E03H0F91ctzEFEe6GTpYc6q2BQT2e6hOzF4yCzetVtm7GjmrV3U+o063
1RBpVKR1MB/Vej3Qm8+b3aeQuKnOq6qRbZL0doJHvaElk0u3vCRZsW1laNLZFBBriJnhZYsghr0X
TU5cUvgiXPlERovvK33s9nUHLUp5/Jt2+Hh6MlgQN2s5405ng5nv8ojCAw362MZM5uryBRd18Ku4
HhSlTK3YaaxaiAf3iQni51aV0h+ElF58koHh32eozOg+hvA6B9pTAUXYH9PT/5N6q8IbFLyAh8wX
bBoKXmmDKoDIPNpxWUGFk+IEvFShzfMP7BZ0rZhxIZ+RBHHWeCuoethmVEMwsvelPSA8LRHfY1WH
fpavZFnzfxI4kw5h/TcX69zyR32VFiE2GwGz9UyV1B622wEEU04tO0nnNJap49/XqobAFwWZbXes
YzaLwCW4/6jyGJnvGEOa9V9XYc7Z/rX94yiGudizgSp1l3+9YK7kMwlqx/6pbP/60IiLOWqiUar8
VmJFHZMEqxWrehUX6NCPrOMerL24kxftx7oSTZenXU3pnO45cpQfNexBOsMzZgjxio2XsG/d52VH
ptw6mg9o+eGn5xPu1foItkmhm9prTzEoJ3j062vuUWWYtUZlM97nmr4Yj8+7yCIJWRQmCMZc8skE
tM3ks3sIFTnkPopFlmAxpiasn3ZyGE3I9OtX0W6m5Zf4f0i53+vyRuquyvm5KO95YucQovaFLeet
i1Oqi+hsv+ZHiR+NGm5ZcQUDRjGB9ThwQ9+6fI5lqNvcOGsc9+150QDLZyW6m4zZFWtfo/mKyrOh
94LBiuXauRn45CsI6eondmNxHfG30JAseaM3FqUouSI7/3/2SINmRHiYVVGRfPvgNSq64ENNoYwo
M3YdMbU2AlPb5RZblRe007lGy+ZUpvfuzO2m88uNQ8XINGSITDTCUzLELX/0t/bICcgW+w0cD4F1
f6pXuRtkOk+SqhuZaWy4vMn4MjyJzdjR6JxXiUoQASneIOSmPmDDZwIoJNyiVsiGN5st6PLtywpc
T6ZDUHH7P6OWZxeMY25k5e+Q19X6vzFrbgpKRrn/axklOMnlv7QvJt0pcVk2V+oCH64RmnPtT8Hu
k+u9pBv4F8sx+I7iElmcpuXVAZ6Ok5P1CP2CNqhD5rE8VEH1u+S5QWPygmV2kEyPob00vM8mpfQ9
M+MXoqAOwMhHar2KGK4LwLPnfYgmfClaAUiAtEzne2Pw7/S3/YfDmGTyM4c0N5dxzfqbKJVmlelh
6KF6v3a8UbRSHPV4ySeetQ6w/uXP49aMgO7j+8d5R8VGrtk9iihE493AOiIlMdTSsMSrkeGz5+kB
GZVbCX6i8ccYkVr2/N/l/3OrvDuFkrI93r4nHxB5jpyfGQlM8ayvbcaIujwb9zhSVLf0y+vaeRBy
nVsNty8NqwrSXRiCbG6eAP6R8ldhExHhCxbsDpbScEmozcxptrDJ0q88mE3J9padni5eeW669Ip8
F8rbJCY9FGhkfl5V0O73qutkJjWG9NiMvmbWd2J5qXNFWylsmHRimJrqb+5jKqCfhKTnhTpbPI6k
vf5fKnYleNNuvQlDzsauC6baf2YKm38Am5ZkttyVIYdNr3TsFo+6+T4u3i4NB5dfdP8+L13fZmK2
QzB+gpUfUiY3cOtZw8pBmAZgusSdjjp5YlDZ7+Kcb9HgCNTBiY61eRbdPRoSBYETtZFkh2ACtPZz
vR2P7xyyFSgXBDEdgmrIjluok/L5dr4a2XkPOrWD/RGIxAMTXXfxHdFMuo/uM4FquPi5Puir445W
ZItoa8zBQvJbRR1ThkJFjr/ALL2ydVAu1t+2nx4LYok3Nb+2b62WerKsqHatT0fSpSU3B3mE7+Fw
LCUam1bQeCI0dc0G8o8LhUVoivu7lCU9ouwRSsQEfeGLie3TwrJPiAnwN7SK1usIERTV5JF/HgR5
N7toEf7CKd8iknWAQn3gSMx8eOCp9QKapQj3Ffn+uYeSbc8fhhvNXoS6rmTsoWyqVyvfoIKjN5jH
gXy6x6B9nEanzB3sJIBwIJWj5WLJ30EZVT+SSHSmX7ViEN+/MHI3t/gTBJOZaBmqO6iRLfgfXgrQ
ILtlHxnfv0JSmMcavRDZ7WBvGjwXkg3HS9/VUNHAH9m8fDYKASbIB/mUM4jthxoz1Ib3z74GJGW2
qEUCELKPR3Fr7xTmez3z4VOu3eYCfSXvFErYkx2hkLIbdG9tVuLOhvEb+DDfyDM9mbSGy8s9+6ax
CeY9xdnMuXufZp1Q/8GpruEBodtn4m4r2wqV+M1TwIlj3UNmSi/ZOdvRcPnq4zHQmnn7tzpzOEnz
mFbCiwi6ODvBtxgghR/tBEXltDEG3BxZKB+kM6tEMfABTzy6XPsgaW0xkCpbIPEaY5UicqbrnC2V
F+Ek9zbJYqduycSQCo0QlCxfSAJ/1zcaKnVAvqPsBQKpjI9e949jQdlrHdqP78suzKxnjEE2ppgk
ZntqkIi98gHXY3XY+g5szUP1ZlC6A4xxTvF+2/ynsE5KCsBh/boHlAVGOdeITa+VehymFHBKHy4Y
fqH95ONn+E2HQ74fPPuGynyhFNCUcnxXh7UhEu9wFySH7bvTDYUc+rDnncdFYnqztUDjVWA1aNXa
tSuyjD3QkR1b9AX1ypiBjNN9hAl+XxQlubTOpXOiUS17mbed2TzW/XNvrnkag8/fpV9D1tesadTd
ZDOpVBNikBFb/zQZMC+T6NfblxImjdFyoaTRsVNFWMzrJq6D3uyH5fpEOYweMro3H3+oLTNCmnlQ
B1grB8D2bpkvL6TQY0j1Ov37pmnwNr0439vpdGDSTl2EuIjjFvuUi+0rvq0L34QzCSH9KI7oSp0d
B+vjwfPzPD0SxYrpI8J6mIf6BdKie1ptd7zplZZIEyTMTZjfpGgNQJ4QPp0n0k7IfzucrcaXi79w
iVIYzFSQrJTQ5+OfkveVHj2eoFdqNTEGfqtO+uXpaw9Vet1/tOb2twXtrtuLNBEbYN6rnSujEWHU
TnAA1GMZhNMeuoR04J3XUrZpFX9gf9CuWtm+8AX9I+84ywktEW3vp8vJFLftT3GhPHTPzCgBInRd
jHK3ZGnAGY1Qet1Igw6GepXLKLmhI2SyAhTPU56h8UWJg3IyPqraADS6KJE7GRmzjk+IenkceC8X
rU7jHHtCCy3AYw/xVUHrJ01ycFr3knCuZBS0fCl9D+RBfWx8bujZzKfBr7DIp2GdED1ZpWOyvIVm
w46Q4x4Gy5xrkv7FpH+wEsqHIKVf7Sj1dwBm5pkihASUPApOJx9Zi2wyi5AytptOwJfK/goQG+ah
EXAp2p/ZqLdwylLc1qBW2m3GAAytRSl+VlANzyNAJHjx1Tb/ZwOPKv19Lw4J2JRtTZYkmbZ+Z+lP
w7uQPmtktlE5M3zToK7MJ0nehkBJ/7PnRYlfy0KVE1s5zHphldpMTUpdJJiM6zNKsyuETljd0AkV
FA4Mx6iGM57Rr/FCGW3B/rbJiF3xrqxSDzMXD1/l9Te4B6+77yzRYSdY7LypJEFkTxh/nIzHo5lA
VB5+9XqHmmSVlppEqqYTeIBy61ViLstDQFcZuyrnrg7eRP0NZMdsVSA6crzlYmEqPPn78mlGB/Oo
pFr9YEwbgLizRZ5j2CzFIFKdBmZQikOHyADoQlq1olhL1nQyHOcGGB3nitlp35eAOl6MZ7IIcmOt
MmYod2l4nFOo/i01Ykc8W+AescMDyhrHJUXC3kfA9qx5tGTbie79A+beregEkXZW0it+IZZKJs6V
eh1J4578DVQMge/1WawU5ySefiAHnKCFu5l7J708JWjoYIa1yfJch23E/xcjpDzyFzneXouTwb+g
aoJLuPIAYTBLLYrOmH2a0s8rY7DJeJVEBmf+MXC6q9X8TSR43GMBlXO+8Q0a5LQz8n0/4WKtHhdO
e7l0ThG1q6FCQM6bhZ28orlkh4b0Uy+0J2SyQ6AlFLC4lykcUQvRe2Z9n0ZhF5zXFyyvGMhSHQsC
8E+5Ln4gPG3frzqMHh2V/skPsiuZSAbgv4yk1OayoEWA6wDpC6RDzJ5FDpfTgCIzHdKDjgBxUUP/
9dB5sJxMGSJwv0yt/q350nxBJ6LZVhWenQir9FIbK7YnlYlEi3qU5kpymYC1rrGoCLGoo/X2Hzej
fe9kcR+PSuY2m9fBFEQcI22mmkD403lOSwSmiVHh8pdrw2VuJR62YAfMgRBfzb1cWOmYTi5lIlg9
tProT5uKKsuNzJdXz77+Ql75Z7gxJS4f/PZG/TlkSLCItIWCmXEVPapB8yfk8QntRblY7b+TkQ4K
1DXySmvfNSIvLm2Xxud47Ryry8grdk80gOJwFCZg4zzCBUXP22wxYm78CCdExRcwOB+ZNKReISvU
FR37wD2Q7QnHk4GFSwDbPFENxdZPficD2gFzEPl12Ygkjrs+9pIRARbpAL19zEMD7ur1l4UEv1sk
rItku9Sy8Qd/ohQR6MfzAzOB9eBTYEcMrJxanLsjGS5GkU8u7XM1OKsxooU6JoybKGmjAYEJc4An
cB5RSRwQAsBVp0EY2Z1Tr3rZHstVn1wO7RhKRKBVnzDizWrXLpPrjwg//R9neSijnJLLPA27YKsL
d7gIk1y905PyVY7IIahfZFYjLDlxCiv66mZ09tr4ZmaZMUkMrLzEG9R2v/d2MtENfsEHUtmxaIwO
P3MgXtrx2KlDQ0FMpmp9kmWAtRsgZ5gt7YW+HAAsPTix/PvddwnSVqAQagdlgp4q0i+UoWbooGSH
WE1Y0JgWJzm8DWWB40OhezyU61vM00+Ti6dbihjQdtgIcD4d6XJeudsBR2Rrru+gooC0NsHhXfH8
dKkHP3q8v0EtcvG4eG618PiZqXut4SWMYjZ9pYSc1dzOq5X5X6xBxXLJRjdb4AAEHcS7s6yZJPTt
aN7k80Qlm7JJEDOUo7h1KTQmpLdgqdSovNRLX35Vg4hmksvz5AallAnkRFGlMfaU2XtwujFRjgkS
QvnckfAAlKlNU0ZC9Jkq0KnPaQJoKjZWBUwJ7MCf/ENJDyZnVxYYhVT3cn4tqg6k82BcYX41k3dp
PUMo4p2xT5MJ4vP2M+MCIsRIeydpr76Ieur5UkGYIJHwnk1JEBhf90AFMKSFsuPpN69QF3qJIRk6
1fQa8ZJ8ILGa8w5gHtnuT762Xy/NOE64j+e2+45Wghge2kXIFoqzw0zhfbmw1GVuxxxLhD54a0+f
7jXbKPMAXg64q2Qxk0myKSBLkPedqc9lPTRKcn4xc6TweP91CjmhPrY/RZvOzzlhq3ytGuT9U+b5
6WDrr4sqaaTuDODNliectfcr6zzn0s4l6gGqnQiBB1YWvUH1ur0lV1PYgIsIPmY6awvlECA243D7
sY0JM1VYhC4JFtxDnlblPQ1NTnmbnljr1HxkVFcJyi97u/7NyT7OW41312qEgplHiEVTPuAx0B4O
5dWkitQAgra+JAe/ELxTINbAKZjSbqTOIGuWcn5IreFAAMGcEL0aLGr9YX2HYhT4OwYs4MkJ7gsT
sCpwi/wxdWOgPMwMFs1hm3VPC+IR4owR0yMWvaMY1kXm0x7YepEMin/f+VANafgvHwdIwrpqwtJe
q2KnlVPsIVvvx43aP4J5rjot4wE1hax6YGorIu85PKT6oQDhStzym6pxyvTTThtqm8ejxlQnAX4C
OYIwI+VRFwpELlrQ3uKKaxnehNGDKFMgkHIixh/bHHDT30wfOfdwlT4z+wjBE/8dn7UAdQ1Vyjbp
HWHhBHy4aZfAfuk/JT1U+Irh247CgaeIPimoWtTPLs/Teu1SxDaZEmJDXN3B/gyBvEx+KQH8D20k
H2oMC2hJR2Fw9w/TtyAJJX7OTI60pPFG5rhNINIAJS4cKg1kKIKTISjTvq44DjybVvjgbqsFzTMo
ldYKDoTh+0lNAUfSVNdFTj2DHW605Eom8C+QDc3s87qRk0mufyJY8w2TVsJx7uZd5O8P7yg7WlWG
RjMJdTh1ajDhd8MulnD0osZkVoJUwB4Cn8nokdwCKSmkzBdU6BzFrqaN+Fvfz2oETgSJNLj6r1ip
tsk9ijJr5mgkTB9BoGiO7Bt5VsynpCY85W2xP1ulGBV04lMiwIFZMUzrDwJ/2qhbjtz3h7JkTn/c
P6M8jF2Han+d7lMnoK19vg1PDc4DrlcUk1RJCMw0qET3PmUX3wXr9Igm/m9dYl7bzPg3O2T6DLwS
lhcBHPHqigdEjCIrrGfkM8JA49pdX9yq+q5YwIzbr6LO1+ZiddzT2kEDzALJbsk7TUAW5XdbpjDz
CqA2eesut0bt4H7HhoYzlQYpOSpIq9EikkVSRwkwywaU0bBevr8WZH2XydLwNYdD7Zo1u09X9jZk
xQrgW5p1u6N3waFr/j/HSlY4oUa2iyyRHtf48yGS3XVBk32YJ56DxG68OvkQdN4yrNYZcSm6x2cn
QpTmyFoWGFINiM5OW/B36CpMdsdLWr1V8zSNtLoLZMdPrVPQ9SJEArnAKRh7MK6Cw7JhWqIWiJ1i
JjYFxDwdNtYbN0ePgDF7386Z4SmB0+d28nwqpWVnGkdh3K7HzdKX/+61DXq43SZZwC3nB+cWYKNU
AVNLG+RgdSay4jxzXtVHf2mwNxrcnUzCw+LYCIxTpgR8AObXfbfvyRKlLPl63Yui0Uuudeak986M
UwHbpcjPGJhcHI+ZjDeQlWNlB9j6jBzUPc2lPFgrCB/aXC0C3gNHJ4+FKvK71q7VJg2/dpB3xXvB
cL94G6/pi8pYb6ThGaZHyVMC7YLG0WMJDKTRYg8f5iOsS14BcF3btx/QuHU8AwHeST7BgkCsPXjB
AC38YXqehoWAIk3pPhwIyDMPQ/67mdr3b7POdcUTXDfwpp/qwWkOTnzNUNXbjmEgPP1pZ/AEkM+k
U+SKH7nObxJI29Ip32DQ5snL/mLnqc079TvprvREr1VmiX5X9pDthN3H5MF0bxrJIlRNL9BNOJoC
FCBOSHKk4QOvl1wAJst9a4mB9hbmaw71ZNcT06SMry8mFC6rK87pC2cIjWLlK5Mh/tctZjeYaZbz
XaO+F7We6knF5vS/3KIx9pSlNewDiDe1FZfwEbOpwJlAUL4gHX4jw3PDOYzWWq2Hv/aMQvM/itft
mecESjt5fS64+8IKHWogLoYekblOJLdFsNb3LfljPGaZpNBOc0J2hgPGOHPkTMA/pg7XWJlgyZMk
PJX5TpGi7xylPJCiohWBj84+GVYXVesHM38Ea+wwGst/1/kQBqbN1OycmmrkL99+lGP4273Ypjxx
al0L3fRmQM9I6/xtFNNW9d1bIOPjG2NH6scZih96YGVqe4V8YvaijTciHg3xbJ6VvmpD0hbHmlvD
tG2/t/j/NajXA9i/iSj10RkwTGWVSro5Xxn9a0eTPMlqIBrof7ooBnehBuZ0feOz/gKa5HwktAoZ
TmjdPgVM1R7d4WjNkXRKof4UKY0v6QPz46lfjimufvycqiadlCAOQxESsx/MF9wROKIpWAjdsAeg
4gFk5mhakcqyiZeskn8U2F9UYrI8BTaJqrNgIJ+IEDYZIfLV8XLT9vr3zb1rpGnte53Qs+LFbYM8
GKkTGAtS8M4KhsV5Rd2/kukWgHFKquV9FUg4AqCRz7SfSIdjGDoB96QTsm5wRTlqFZMGOJ9eaQ5v
W+Czk0+sd/nYgHXi+pNros3Zib7bRCWCvzWaeg8JjM8y+JANEA0/PBBmLLZ4bV9VrI+nqpFjLMnh
iySPZ3NfBGUCK8Ohdg/F6U+ZAG1b1GZ6H1kLV/+R2DmlOs+ECYyaIc8swgjDrnq50Urq9RKqRBOP
RuEXIQrHaVNenJoj09SxHlzRpgsAt1C1bz1BpgCGPaxlRqLD4YnEkpkbwGeAtKr2FkvWBYY1O5Aq
l+Jy7r6lXETnNa5uUJbOZc8fR+hqnztEv3tWvlpZqF1ckLaqTgvt/HVBn27sYcuO0jgWxomqB58U
LjGzvIeiFfRoOOuGrq694z31cu9Q2DPQVq0k4IgVx3MWQLSqAJN7msatnktBx9QIauck5/S4FdLU
AXxWHgcziDkJR7luEM+phan+NxA2LndX7rPGalYIvsWeO7kQkvzhdvXXkp4zdks5cQzt6k1Ey4dL
oefnTQpK5u//Fmwr+g4n5oLgeSnAWf98MttuwLmmaFS58UD1/IabuRukkpZuoqAHFC9pJwgiaHD7
FGuKHu+QHvkB7Bx0zpXs/oeb/ymSEr/PKsJDoXLhc+AhNgF/MBqkAT+QZUbnMZE0qkA3psl2gq+9
G/1CchIoGx3noFut2pgxB1O6VChav/lr2H8Rdl1vdJGcd2VczB55BPvNw46UlFyxhfLB9JJf8iMd
8Hxk/kFdYWZM4Y/f8sTXFYbZPHZGGIAbMxToMeCTUkz1vaEuklvLMc0HXLVWPdXigfWsFBYlO/rM
Ql9PD2RFCPSJpQqdYlOXPD1vdOd3gJ0Qe2RhlXVVTFg6ya+AKeaOPPxiiBfcAbWkl1tDFaqndA8i
BGtBrdpbR/DAI3JhscZyr7F8JN7UmKsoVr+OHUZNpOytklzf/RxF9l3tr3H1hO/u9CIQVR6tExdl
6Yra8UEyUupFJ+0DgSo1mnQdpXc8Gl6G/FDMXEpUom/D5fN1WAd2yAnR9UFtD6dbk9L0y7Fea2eJ
kEoh+OsBOrsHG3+IBeaMvXMQI7gsM8qPE94hplwb1VjeMWjY6ItahCRpJeM+uVPnCmzoLqHk3iGS
8Li8nYRhSP8Nu8OgWT/pRNHOVQWRRHyp/BNPAYS2+9Dx4Usn5Yv9Ig91edeKHyEILXUz3Anhzd6T
68tB/9UWcCVAStDNz21UFXOtCgou9MRxAMn2yVXbrnVDsJxYt9RhlVBAh6YL3RA3Z0oDLVuEgAKU
0v94UL5zq/7nFiywBJWTh3N0VXB/R6wK0wdvDNNwQ6L2j+70VjWSFMKkooUbT+nvsH25d/aSqyb1
KZHdL4HgLX20mmSvCL4n09ujbKaTlj/EAX3V31HxsEKEhue9e4Za8dVI1cT982n/GrMmqSHwp49I
PxAjobDVJ3LYGxoo7APRrEEN9Z4k6A/Qhh3oLOioq77/MBNLwFu0Zdhqu8l+C7ydjH+H+Zvwlpsf
crcRC37Xo/dLpQrgkJ0y84N5ShDsC63B9usmDf3LAljUZjXu/oTaAGFIIK3l4XtdnH1G6V/9W51l
zfUz5pNEL4YYEsa9YP9k30FotiCOgnLmdnERF7kAZ0zB8QJUKVWjnbtOJn9nO/0fY4SNkfkS4WFg
pegDJF9AxqRYo7R9XR5NNyp8Fs74oFHnixPyo7+VFJnOkj0rQFsHQ9fPefXAySeYHxNL/BjNW3Nu
fB0Eg8FYpjHwFhnPW54odaZrP7IUg8/YzReNOqZl0MxLYz/fYJakQE50/tf/q8ClEm3QdL3KzmRf
t6tP8VD5CdKZ0KE7KLQHH27GZjYnmrLKxy0CBD4vDHIigF+z2xqzk2YwE2XKMSTPdHlqvYOB7Gab
wKCYj7k1Llmk4u8qJEe+YIC+QVViJKK5Nri8jKta94kIlvV5h6nZoAdHagRVhXny7W7KCZSZ5h9w
N+pgDxbUiSRRDM8N4nLk8aERSeA5Of2YS52CYAbNJ6Z2bm8MrtRyrqNFzSkY7k0dMYh/fFMXB7dV
n665dsm06mxkOYKuGQ2qnqz3LHniDQ2GYlhYPiM1Gd/o/EUNtchMMvsndrRKEY01R+s7sN7/f5Kf
IoR7Sylw7LFzmQyl1Cm8xLHiYynNKLkyPiGyaZ+CIygBfAOLBotxHh4i+Cz8DxtSmDuochl1AV+X
cWhYdWkUXfNHZEoNtphBLepgyvWVv0lu1ekgr1pXRo5BrIgdttNoTKBkb1IZR7GfUviISHXV1ejJ
x8qEXC6JCFYN4Au//6OVTzg7O9IZ+il7y9vLqawjHfAlmHTE8ppOFIhbCc+5nW4X1WjhaiJtnp+J
b6rQ/j8zQYC3DQQbtH+DB+mjz1t+odCZMdENiT7Emh2tIMUMfwJ+hYcDGdIzvoAc7FqZVfj3fjk+
25x7i+pNz+w8u2afuqmNN7Mnwndjjm3YQf/LpQPC6lvWPpPcTCGujx/kVgNo9zEXVJRPpuNz4XTn
5O+viiiNk9ioqzp0/0TAxqssEs7ni5Frqa5dqnretUm9feqjIr1xRD3u+w0J3f+FT1T7Us3TvKrO
d35z78dplXhUPsT0Hrkfj3aEbtuZMpqYt8by5997tTAHES3b5r5vM0weMtDRbfB1ENkulqJ+1o7f
onDHWgnC4ZxnP/uoB/9Zk75BiCJlRvivHlNB3QjCNLuf0EenFp665vgRqU9mtwX0w+5RcsOOwBAZ
n9TFC/QOr2ImRg5nqelicmPrHZ41ds0fGeAKhktY9s5pCWh2PzE/F8kD5IUro3OMCxITgL4vKKr8
XUuImYd1Fm4gHHmWMpSNMRVMfj/np2vvE22W2kPhnhYXEJ09Y5wZr1w4hioyxwDwEi0QTuN6Uolv
88qlgF8u6SX058PimKy/XNmu/E4UwdNRCQZFOYU+94ztYrxqmuK75buB9kO5o3b7D71zcxdVmfND
LPNCuFwGXVval2QN+PdaNFGDhBb8buFhWGcXLfmPaPVlcnGR+hRhfX5QYjd+gblA15xP+IekNwbn
AKAzUsHAnQSw9xMWKLwWSkTLBpQDbrqha55pWiteNIBB4ennH2zGG0KIUOhpktMCp4PbH3JRW0oD
5ztN5GPTftT4Muf0ALf0QzBSOKWe6IxIlH30uMWDNWBcrdh74Eqz5i1oj0sXmKjjcBzzMcpor/z+
AjtTbmpr5gdHb+X2Q6w1VySNJzIrA9zSbRg9xd5Av7DupUjaBtGtm/S7024FxPQcrbqwDQ40E5p9
grzb515Ed6XJ+K+sI5InSI4g2npVf8gfgFa4Efvi6PgFyP6qBquvqwyNWc8RIiPCCG67suuNG9st
wSVRY+7wcNPKcFwpl/5fB7cGxp0rQsr6gidAYGLlk9E0EL+na1XFpai5wZmEaKjsGwONCNq6Q3Jz
WSf1J/TC+62L1dsoIvo+z/DhtxvmsNZrjuslFrU7SvKjfq663ucVLLzCqiICxd+x7wL6gjeR47Jq
uIMUf5CyXvir/dJ3Qb6V8FBYLrzLuIMEixiNoFC7P6ZwaBy6BPdDK7wOLu+M/DZQ0MLXciKkvVC4
5c/wprGU4nnAk26wp5aI/NiEbmD5nrmeSua5wDapJcGdx+H//yVGeDogfHkWrLHMavAehRtNkxFc
+43O1dTGhprTlfwHCy6DBSzq7qUniriHMA3ewkTNod1P12rqEfT5mbbx54nwQqVIZNyZB5d8uhyg
6O+me8ENp3+gubBLXP1Pv+s4W/HxxXYCqyTRk0HjB6yiFMwY7suQBfAvPZR7ZlLBKupaOqAWqBOa
gBJR2DG9Zspz+H7FB7tNgqE4MYBFgIiXh7xQrjWjZ055Ziw4RMEY/cUup6z0QPEnXbe4nmDPGmNT
lc2TXs1HNtBO9ZYn/pscD0N2IGe8SS6LJdCkSJxSrE5XuRtGCJzKqLcM7Hp3NEnWzD3t1NWB92u0
pMSzCTHh+bymz0aWECZAGWu6oKX//Q43NQUVgkSbb7ZWwgA4X+gwp0ltcOgGOkEktfOo+pl0SSxF
hHI60KfXWobgMOvqBgsCfLTbhDAnP8XItrnvhtFxOIi5lXoj4jqYNFrQnPzZ3WbEKtgEan7iPrje
rhH++EKCPkG3U0+P839j5jI9DCXaJjLdk9jU1TW985y/5qxooXXuB6C91jKf5toYJRG39vBZx7eg
FfB0cGs06rRkgXWgO8KlNs/k5hl0I44P3572NH3oFC0CUZtPzBqCXplxeXePolyrrfU4PmRlzXgk
5Jiw2Ghnh0brpiuGxHL6rJtFjl2+zquFRYXFcwBU+bbpP8z9XpSKBTKBZI4NaJkXLmFXu7lGZpum
cl6YqHRqkDwf1Kle0oeGumUBjmUxzZtiGm+kvvykBXhxhfYY7F8GNJBcppzaHJzTn5RdK+0b7Zbj
crZR6vmHq2XQ8FCLjBkAkkEVReZ78RxZq8Ol1JJv5kabJh7X1o4S6fzmJ+/w3Ut/gVdD9JImGlTk
zJP8NNM+u4b3ld1fmeGWNHmzvMUkI2b8TCJsUr9J8N1WK6W90b81dtEPPf8bCy+WJ2zGC5DCpwI/
qMreSyyuEJW4V57SeqSS0iQlQV1cMKt3nC9n7jE3RdUw8oj744yFo1Grw9P6dgXycea2sQ/Iavmc
d1WQC5GfUJpcQzxtmeVj5vZvEGq6CUlNNlRHk10OV8f7ZtwzYJxxgcNxAJE/mG04y9/r3A5dC20q
jfW0h10Je+4CkL9DHCpfn9mflDVhnYKFVq10f2a7m7yMSYOarFFZxHpFVx61Z0Dv65J1THFifBPU
u+Ix2wSAAUJ6hcnWuO1s6chm/VZSpdqeHOtcHkrfysQP5VQgeacZyBrdK/WvLbux9x6ST/ypiVcm
fmxy7XGUYTEDtYzvcFH6OmvVqQIBZ+L6D3En3cBYSMw1ohuBF4Ke1s2fjGdjPLLyBYGpohnl2vBJ
lj1HaEZ0ZDqmlYfSjOapbyLHxPtZcboOC9de59gIY9g9YzCGCiAC/BesAsWb2Y+cIq1ag0R9k9K4
1MK60ZoZHH6fsPSfEm5xUXhxoDUrsIn8VIDdM3e9T92XernrmsqLB0mYEv7XP63wTmGjkQVFM2tE
Noz97RlhVq7+WaTnrA1RmKt/HVRI7WDAWS/Fi3hpDhp5oN/YJ1yapAayLijC0uNR10SQVFgIBwM5
nIrNGrxdwVh4Gw+J5ZzY+wMsSg1az78ejCrU9WopQvnMhpgn29KPsEHRkbMZs7jlNT4ySQPV6x0c
hZgaZ+PqKrmcuTERmOfN1jstOeMQerwgXH2OdXmzVnm5N2YaRO943djdioLV35fPmwJfUGlwOuX2
fuNceeirZZtL6kq1T+qUqAOFanNNWBXjGg54/vVYL7VkM/5/MruFO478HXObcroW0gc+45JHmpAX
QU8oaQ+a/0v74b2HdjvL1zEi42UMUm3D9D2Zc49yzWYDDjzGwlPQ5Wmc1uyibAaY1X1rSIxULes3
8ckvaRzlr/QM7kdjq9P4V9xn2PNjaUkT+uP+5Ixz24CXFkx1xbMLC/3Vomm/2M2Obn6A13e0zwx5
Ex9eW2zBvXbMjJxe5jvRpcWtpNcFem0ebr8OCLE1NUc47b6zbJZ9VCxz0ygaxBt+Ha+laCFirwEG
jAno1Ioqiw4z4Tx9VSHEAf9UAzWdeVgJHCge9gQFUPQ6vsWDTFMaI+Zme8OnN5SUbzRnN6Mjkgea
7YkODibj8A2ohTsAbMy9Ep90CASD5Irjzt+CiyftOmNBdtf8HcL5UbIlfxS98h5gBh1NbqfrvdTF
TYsrQeWhKagG2ypkMH5YBOg5YNJ9xEf/alxTM5WbeIU6EE6Ug26ZPpDECXkYylnDbG4VmkKyFFgr
azK0ReYYMapCP2+ewncr8SehQuqzzvpLtMlHgJRRUwLB+QSRt2woceAl5iE8ymQmVuR+rS23QlPB
ZqHYpF5Ajpnr274G48KHXjt0MkxaVluLD8b2/exYvCk2eU4iNFc1eSd2I1ibc95ooLRW4AlgOsZj
QNgQ6PGzRgoYryeC1DW88zwWEWrpBNDeq33TI+A0leGCA6/RCdNhFEhHZltF/2utQdQJYR2b4H/z
0HuqezzdtrKwJZz2YT3HRrj771rshX4bdq43GC77QKYqnEOvajMMpPKXgCg2Shu/AKhGLxu0mgWN
HJlg+26VOfKaqmU6NUdNPDe2lqh4m+QKRBjMt4a2+AJFNQGVjcCNIFVQ+EsPdQqlFH0/E2UZfCjw
eEAZP6EgxMbuTd4W0/zuUS2aWYWB7TgGxtjPvza9pUSAj72whLDYsIlLeu8GsXKke/JfI587jbBK
zwnvvkCUFWfi5jXw5jM6I198uZFSx6o9FPqI9RfaBNv7ZRRInNGs/dVjvFbF3G/XqLs/z3S5QeIi
NbKDoAtOSZawpmefGVKkUFg7YHx6Oz9xHY+VO5+tOnLNX3SbqrMww/lFzUbfx+Qnlw5N06Y1E3G1
61Obt4VewRAs/9Gjt2HLO7AyFszIZxlF6ES3+JpxYcV59NjobLKwoTiwFETyv/KlkvzIgm1JXxDF
a6UPxXzXVCIepGO5+wG7vMiIiE2Mt0lPUZmCYNXKGTUezklVX74UWOjA3yE3a/ask7P2UboTuCk1
pmTxs8OHQY5kEjrGygk4jTPmNAvhgcbNVk/ZqUGwP5omGLXsWAqGzrwsBjevz9YX4D/kNyJGUq/h
3p5VLnVbKB74N5X3g+Y0YwsjzwiEx4p3tcXpXh6D5PuYYxiwYEIiEbJc5W0bvtO8ZpMWopG8Gt7v
RLp4rZFO2u6cYh+54rZ/94YO6mSp5x2D/jnrVvvuqD968ZXoXnKd66mSFPEe6y8grd6hl8aBWWL7
ZRddAwK+mRDsHk2Qfo488Nt9CaBh6iGZrWAXYbVHS3KRHZnF2fCF9/3XHvzM3jT554UuOijUF4cX
m3OIkoCpiQ2AF3VDsjqDiWpLk48hYYwYDHymgXeHh7VtSsbYsQlkvJ/+G9/ADfpC3YNiY0Mnns09
V9lFKMHyFNnAoBBkIQ7h03am3J9oEBCNaQYAmicIeTHyi1bKVVPwPoa40oMy2PokhlmOD50cKCrS
cF8igk+mcy6vZC01/CZvSnkI2MR4JHQzIf/Iwho3k3yblS2b8KA5N4ymxGmLdWCvRV8tDiB15Z3C
9TQyVlLZc3uUbC10zqJ4+WZvULSR77O7fASxirA27CD8crCNtQFmnJM+xIUwLmdA1v8aQF8a80bU
jRjSXyNsAzT3b9xuZKKy58/5f+Q3gfnmoUbDLPdeXD7AzfHLcBrL5eH1WOABFxL5XTldbeUJiT2B
AzOHh4syg+kB8rnaKrCNSw5YOvsp9y0Rc3dUlDVPnJVbFSJLk0h6JV4bUNA9qHMRWtbL0HMYjNxv
wJuHuI6tSRs9llPZuLur4n8uC/EdRErxrvYbK96SclWVxIAQvbCoj1ys8gRlSNsuJsaI22pTdXTg
cl2d/lZ91vnZdMXB1p2xCD3j0C3IscJDMq4xDb/w+Si+TcIGiI5MtisOs/O3op9+Ej79L+mjMYob
rihAO0GaPzrYOTwxXeIKYOjSnSPOLpVY98hdDy0yLwgXQ9el6MFoRMLbJ0GXr4xLljb6Xxvk68a7
gm8WKzCzrCB3NRit+waGiMh6yHb2trbrO/GcehJ5RRpV9IxSCTq+VmnN60t3eolkx1zfN86BPNMj
086Edtw0vVnUObZkKPgzCsf0uXFrmYAEOUUETlxvRPpzz/I1Lp3fIGQKZzrj3XILO9TUIOjDL9UB
fJcQINYQnqvzoWJkkmkv+se5JZUy1HgN8Hf/5RH2HK5IIgcuVqNMrEgfiMu+3lEXiOs4rua2vdIj
OtQt+QDSHghfUwbIJJB5+G5R1OdQN077X/Sx4Cx9eqcANDDpH/y5Gd6nh/alJNum7GO4saWhlym7
4jyBb44r+uEwQyg4hqXcBcH6kA8SHtHydX3/3i0HR0TtbVfboM2GG3sz7p7ylllhOAzjM/hhAubR
EQF7iye6u0eQmoQfbKAAr/E0LqBpalytNAAoibwu/fOzc+wy6V0ZuMrLwGnScvvkHtVR2OUFMHYb
51twI44BmGRVqkwGoSbjuboqvIKc8p3J0726UPgpzqGZMACXTiighkqiTB8LDi82oIxLI6YImAac
fzDqtH2HTpdisCLGurKuQcQDMxWILhFtgyUlC0T3DDvO9nmAIWfJ44afFze60dRnS+BjL8IkR3DO
y4ylEnnYHz46VRbnVfOyGBR14/06zsA5KxpgX5bHlwt5JUv/Vl899b13SGWxowPl0IhKxZXV9CeI
eojF6beC9bav0Ln3X8MPNo8/hOKEOgbmA44hDmzty5gcsYEBbCKADQeTO3ZV6ZDdk6BLwStqcR2k
0Ij1yxF8oCtl5FIPkEfLlqtNVyow4oGD5fvY7Sp7nzsOoDfhFROn+bzJRXwDfksGsYxe4GdyQxfn
KaaHoruTVnvGJSssQN4M96Yjgh49E1MK0Z6QMNIJJhTDxWOMebGheTF7qRyi4kfKbnt/RfY8jVvJ
c59QtNoTElmdUhYeL9RYF+d4bGo8+pQpXV6oOyuIuMNYsv3sF+sHsi74Ein7/Tt7IAEkVUkUctNr
JPh3wUcKB1VsKYbNTUD8/o0ltL9ygHmvIYylUzTHDwxzRZ5SGwOeOtuwRjAsRuotpvunoZG5MnkU
RPLZjQWVo+OP/sWrCpCYQAa4cIcuiYi++vPSv6Z2YgDZ0+pudUYw1LCCSlutRUaELCqxyog5QxH/
DGH5S8borrElsLqvGLqikhuqvrBs/7pqHXaa+CU09b8ocP8PL+OtO/hDUl8bdeAmZNV8+b93NDKI
l5wr+khwN8tkSGg9nICcO12S9QgCVUkQ2OLIoZLo1Ywgjo20dmQF+PqbiFBIVBihHD6GuAeGedjl
PCbsXkxFFMhDPLRh7Ac7prUx67zZUCm9IJRvAwHshjECCoSCVw5osaCBkqFsk8RrZkSLSTdPQYa2
LNefiLTEdCMBqKL79Y5UZKxnSBDAxti51ffPR3e+K63czJz2C66XjE4TB9ppzEcsrApa/9pWBbEq
tuIb0xUQS45bcM6uWmDVZRQ/53DvCS7M5YwUAMDQAaAGLLWkvECrG+xeo0lfyl+/wspNIYlF94th
JbepVVZFRLB4nCcMf/WxPCBacBCXFgOYqmwDHaBpwiNok3ifnsXiNYm4odLFTDw8/9ZpomT9q8yY
nlqb6PxK/ffoPhdd8wcMtjIGsE2xhBLDJjP3XdsDDQ2z9umUt2Xn3uEmwWY+aKv70x1fm6XZbMqr
mkq1hI0VWv8SqhHd0W+VUqRKpmS04iDyTEGCt0FhJI4kRCLB4GCjWeZpRqXLozpgQEJcYD78hjDK
SlUoEqvhQiBVp0xd0hclrr7ZAxVqClldZLspGo1pLsXylVYy8yZPo9erhNSQLjfGGjV4PbHYWgyj
BahX3qTmgHA3c8AR1yucEK9ehsFInA29k5nLC7nVN8haSMIxwCCAGbvkndRHhACCsCrhLOkEG3OJ
JmVGn0sHobBPZEPEsmTr7j4D8rDkFZxDMJklrAzx+iFsf3PqTYKOaNmUvDF8Q6TO+TAUpgt2Pn8E
apo4+PPUNfPbfsuVgFxqb6WrEmiPUSmKuCPEKlHJ1VGkzN85xEK+nreZPfWnfWSBHgYjuD0tYl3u
TEIdx6JqFnXFL0nSB8ie+YPWdodcCZrShA2h/0AaSTtzXYMoOMcuKazquTQZsHgXKzopJ2IIoZfh
lFykTwMoJkrZMIdo8selmQfk31pXwXfgbDGPPHeSVa6p5Gtk6Zt/ARSmyl0TA05+z88JjMB1hIG3
sFIYUCHyctImVnhvjkz1378M4wyRY9E33/EleHg+cO7ybREAUjVZnhmYqUsxjc/naM8Lqc8guJRX
601nsg7Ios4spnGUNCutkPd57HzGX8rzBlIg239rNKiR34OkBOGDOYhwyOqUxYI8p9XyHQB1wR1a
W+UO2KUxUI3SX4GITzefgycbSGvHg64t/e+HdubtrZmWpFC4t56V94cAtWXYWtGTK0xYo5KZclND
G1ngSXflDRBdVvccoN1wD/iGKLV2/TltmNiva7/zf7NqmF+tvk44eQgCz1oTrGK1XBju8obaB9+z
JnSnkKqD79IUvszeQpEnCxWQYpZtxRF4NO4TPLMt1/Djoqd5eNMVxxiIkBC2nLxjTkMsH3TumWl4
GyHursGpErhYDylD1gQLYt+XKnZnK0hxmAIEU988vioCl36wnvXflzjX38yV0jKV6BoQch00ZxCC
0Z9Gw5k0jzyx4DQYluQfIs1TMoERmq1O+DR6IEcZyIKNR4DQex725mAgIhNstIkFwty0IFck2rha
MSSsUKyGVamjwvXytOczjfiX8xJKkDphnkSNrSNkf81jvYtGWr+RIKHfKWqd+ApZP2UbqVHMVqiS
wL8z0KwaQdCoLiEG3D7tToXX3pdipOib/o4vVKEmBgRcCNUDGoR7JIKf6A8Ombx8wAkKwj55VH1I
l5XMtqkdq3Om0YzkPfV1B/VIt4CSpN2p+UVrLxOB2jpEDpM+HKM0TkIuTFt/SPtyNfNAFyWhdg55
Mvd2enzpyZP/zmWRN6+zC2V03NUFhU8+Pn47JvOcs8Nj//OXtMkG+eMFgn97fgKAvvXKHv4T0t60
ulVt5+fBZulBI3La78UvFOHW0qX8e1RuB9pemobt//7qSJRqUErmFxglUj4XbNcCbCzGWeW3y8TL
SHlsi/XeBffFbuZF53AJypac8r6VC9C96twkGtSe0DBmMfK5KihCRXnSXD/JeqV1Of7bHCme3ELs
Kayea5/U9Sm+bjZmd4TwF0REUri0ilA9dxOp+jUJI9Nd5lURnnEk+W5kxygJZDai6lLnSD8lwZGp
dwfcxb9mRDLXw/a42nOcfmhP6zNjILq1bsw+sMjMIEYFJnly1AxWi17Mqva6CR2OrRliYaVuzcKb
hnFLkQg3EbL5t4RP5zJuOAsOsgwgnI7NVrdc3O1IHRjLAl45DFdxGo4bM0AJi3AAzYqtajQukLw/
qBDcBj5QX8XQ0hK8xv45UfHooXm/swyNjxmNntP79aZ+TT6TIPL83RWfXL5Q2qzhdmmFYSG40POb
8gcNpqRlkAOibkH1ZpdeKU8ST0cvTV3bdjlzbGreL/zFazFAhHQJiOGHao712+HuvZEWb3skEOn7
j5nTVhmoDh7ZVnd0OUWvxFbSGS5BAtozxiqyTY4PSIFnJp+vZ5Q5Wqmi07ghUdYsP9kNX+IA6Syi
ch7lPZDXbDhI4uMptqAetGU2AuHw3ioT0uq0NMgcVmRr7fONJhnnKZXqwV4F7gdOHS2mY0mZH1F7
yQXmXcfrCL11wYe887Y/04Ljo2iVlfWaoyxrs/H0/L0F0bI3y/uH/y4zSSrMEYX/tUWg4bwM5YB0
wAMsbef213z+Lt07ViywOI+spQJ7h3naGFTikkArv3YZzK84WZoMHY7eit2BHEJS8mMiDdADACnP
3sEiijpD1xnIgeaF4PockRV3oWhsBonWtZhewznKDtJ/qSRxEz0gSXYTbHbmkzslN8udb5WjDPHh
TIwZ24/a2hUxscvViYOwMIkQWVmkhIzN2nAIx0fid5ctfjb6vQxFjloQKkjexV+oEMj4i0YUi10K
sNY0QPS4ZzBsqwE4hVV5GghHKa/y/G4J92GHXLW1plVxJZan4JBQIynu3JrxJJxA1xj8tBAfYpYu
YNIaEgvD2u41+P8J1pcG6YvKGkh8QZpvd8GzUZ7f8x9I/Ore6r95IdimmEvo0dDZZBThGHLTKTWG
2wKL3JzbWZO/wFJzywz1VdiO5CTdEWqny0U4bVNCopaHAIWfZEX53YMyJJiLgyaaH2vYsp9Ocki2
5QlYJzR1eVeSXzcbbyCj5dHCpiC51RYbXI/BcQlrwA7dzP254MWfuaO3Jmb5xIwKdVPFQnm/alb+
y792fp/Uze6ELQBx6pStu7HLWpQvTcMd35va8CLYTdzhr5aZiQ1DJS9XX8D+i3ixzBaVDPf2elue
dUO9pGv05fq5eM6RAuGbEXHgNmlpokAobDyl0oyYhvhnPB/0T3Nxr4QYZtOq5aCtV3BOoq9nfzbc
NXtNqAI4aKZmzuYsm4uZ35tpSjk7aitqMytgm8yLmNTZ8KN707BIKE0GlaG0U65wd2XX0cZ5L34S
0uu/aOq6oYjru0O11DGkB++tAU5vir1JswpvyPbLYjBKz+Od0K+YuyJlUvzs+1OLXTB7Pyp32lGZ
D2/kEUEWvaIG34CO5WAscKY3NFd4zcSb+bp5TiIUZvMZX1Z09CT/W24VnaF8xDsfczpH5agluX+j
E6xAWxAMaRhS/ossgeHMcoIkNYfb4g2wl453dZ7r4IeT3taKEuFZOSPzcEKZUBYonlDkzq5tqIi1
Uo9CtA8ew+bE/1JmFuBt6ba77WHQ0lJqwukAo7uCuc3g1T3IWb+vfa5INxRn1nMEDjKgNGNaqmeG
4B5v4hhrzacqiXGCv0NkB8F/3fKuoOedwK18oiK9w6XGYuUR8ilOT0n1Ad0GjVbdlZFzaGkDfbQ+
Yr729Gcf1w+TuQzUWsFbJtNczO00IkiyMADEjAFi4DdOKVjHbELu+2u7CESVV5qXtKt01bIeIZbh
yCRg2meSo0/gcygcDT0qrrYCkOo+oiiSwvu41kUTIxQqbUcvTyip1fWmLHPwQeCc6GLb1xaXg4wr
bbUsmQ+85ZoQacVZWs5N2nglvl0OQdXGefzTnT5nSf8vogDoN8qrjIGt60i9iQZAlbbcvEUy6WAf
4lypQvDLyUBf9ySG/vHdtfp5rzZQn8bfcElSJIlpAcJqTThJXl4BjW+6gawhjNz3rlF8P2YwRuLX
55Sl2glJcVyYVGCbGOWycwShp8MSs8MbLolO2Wczk2QPq4otnNIHP+9dabbJCvhKzLXsHpijYhCi
3v13KPmU3C+w8G9dtOKHNERWCs7eJoJrIdy2VL3/c3svmuixJIVOGhFF9ABVMn50mMch2zAllZ6Q
JevaRZfZcHSWJzoUfQGncimMm/zSJV1xT4n8fGEj7xPhcD2A4hBJMzRqUNNITnQWDmvfSs3Fs5+Z
hLztM9YicRUdCo3sOEsuplQm7zpfKqvRtI3EdOcu18sPIvFVHaXyAop3eAD8QRk7lQXs7m5nxnQ5
DlvVaPDaYrxsIhiCGNjedZC3Ayp4S4PiuKFZOfTGVUIbGzd/66xamNxvuNbapLdKtEDMKJd/CTX/
eanA5c6iuQtR1AgHj7Syvgq897FBhXEDaDqLdZMyeQVCRidqir5bgg5Qq7ZA1qGh0zKpsdqp6MP8
xCobwyDbzWls36Rb27g5akju2pEkKTDNK5vF8EGgl96JHw945ICV/l21a6bYyiT4jr2K+/nUPUOf
UK9r3LM6QWGgrxNCKuBNFEhtkyTbPEr5PeefCk1ddAaZwWkycqTbEdo5eQ9yKhHGNiluSaX5H7ho
goZ3zlsg7oOfdnUHw5sGmO4Kp7WqUR1GynjOX9t51kpPePfwSE0X8HZ2Z9nJQrFvnISZdHPTL+Yv
eOkqTmxp0HG71C9Xp9xB+tOo9I9sqQihvVf4r0K+bLEbqwhT0wPJs2PHyrI1IaCHvB5gpNNYfvL3
N/7sbRk4Jx/8MzLLgR/nJpVXR9QzGPV2X0gP4QP/Ad9GetVzYrAniKule20YjQ2LFGfNEc1KdETJ
O4YHBUqgm4x6XAECbk+KzDsx4FXvV0xyqj8KwL3JPywG1thWEtu8xe9v2yXr+pYdl9kdbgrmrkJz
kAB9alQtuRsv0m1WBTXdbkfsw1SKFsWxJsFM0uoZeZ242cUn4rnBW7L0KqvF3f0eGJHvY/B/bvwA
qZ0UGJaODMLmatxwLwWJU9ksgBtvZ4jofXP3L5ybfXJbMa21JfjxS8P+xympLf9ZWhZXEMe+wS3r
jtMcpD+rL+W27FOmDeM8t2/vFYv9dkklrah6hs4NcGn5qEZnBmEkJ7IQ7+PHMV2HI1VXmmK77B0F
0XGhJueu1cIjz+TaJJsu8Xa6m8ocGUNQhg5ESNRqKrbq+ONfQsyphFSwuUUvxrP5KhkCicypz37Q
Ea9H/RBFhw+6UI6KpwaWxnWTf3IbE80C/5Ous1c8ic8fK+//+6VhvjNISCZdXRLk2BWa90gwglrv
UeRzRc95SuZAUIu42EyOklPWzaMY/wmXBmhDLh1zuUT3tz6CMx2A0yIXnJ+fTLBM6K9R1Egv65zQ
6nUamEi/vgn+p+eWi1VvqkXKDEnZ/gVWCoqZNpKvwmQZ6Z1JS0XIjWybpKF3kjEBUozu3br8pP4A
c63bB8TG2SHMyZRovZDYZsb0xVyW2cxJjg0Ny99aCGIseZ168I0PQXgkklIldDdmbpc+qR7PmMPR
fQPAlCRH3nGlD3cwQa0yBp3huOdEj6/gTZPOtaIgwwIwIZ2STEz0jxbajW0tIju2badTzbcLZ3ua
ceDdcVckLC+zHXIt5HADi1gftjxVQER0GTCDF1W0kvVtQqm6tKfPLQyuLdiR/GiLJcmVhyvqpL+g
dpje439kmz8MVDXM+uDokjI9jtEsqlPuOys410+4WXWPr9ekRv2wToo0pUKsJHcicTvUHWukyRXh
5wRlSKou6sY+yHRQ9tVNn9KnA2sxjGWmZ+ZL7m2CBtuLekRuAi3NCpYYN47oRKG8QL9gS+Q4L/xb
Kd8i1eP4nN5Mm+l55iOgOFJHNFtWwRrH/NTxVoMJWiZ53/BN2umauJ9qyF04Wk9OhNPSRZyz8POx
D1+Ez1VQIvj010OunXS5pb1FsJYP8CG+CzRYTdJrIGYP8qUuRW1ex8RKELYGEroieyI7kct/BIBw
flxlZS+hGlmn873L/9ZkQ66chCEdY7lZ8oKVrK9kEaCDLUvBjOQJdaLhVMatKs7fLMcZbaPuCxPT
6t0VI/mpT5ZgAAXa4C1ONuJH9qgTVqEVGVelqrTPb4Uho/E9OEoR3pdN40B1jn8U2cmnD8nvVQyA
oUZuVJkKcWyf00P55VqIHEd8/JYddSDPuyi6uwvO2wOxDvb+jA7U/rhIQ+wHyHXVNr2QYCsJvLU9
qVZbHV5SLieNfXxK+KJPHQy7vXD8OeL5SYw9kwsyzgrRsQI1BUP3kFQ/9fTWsHnC2BVbhyOIHF0a
oxKvvbRX5WD6eAlmIsYRryDeR+dX/rjM6F8PCDwpvhc9R5hbC2X/5L2uhdqCGrls9nRqWxLk55y8
5GuOj9pPs4lNPgzHQHacx2uBdoU8RpT+Fe0Ompnuxqte1QcpwSn+UJv2Oywo7+lywvujMbIymbTg
V6qxJXA4NVTnYZaDcTiMWJKmPCKgEonPOeLF9T1w5/e/xlrFKWvGMmKUrjJDF7UG2T+ahsihc0nc
q7oKpTy03q/bX0mbGYHt5ix+aSNOJ2Gr1u2t26J0UUtnDA4VR78S+c/FxhaslEax9IoFWQyw/Frn
9wWaswvskeWe1Suqj1cjCCK1mF79AvYpfqdcEdDIkQK6s80dX1SP6LYAMqSFVc7nF+9uGEA9jqo9
QKpMy0CTRSDF/kTX0rrg90ngKo0CMciyFT9TPBpk3+dvfikDE5U58rxXCp0ANYJ5wJNcfHoLIgTE
xuO5fejXhPNag4eY3Uex9Krfs8rREViLyhJ7VOAsWQEZARUchT1Q2QOalecesTT5tALRP1WySwiI
IICXy4syroJDC+oGqt4vkesbeNjHKQCq3OxULgWu+IbPGFTFPX1GbEcBvIc4uiJF4jpSsvLitvuS
RWiuSkzdKM+m3GVf4SzkvWZECfyr9Z6sGlBmUHJJVu/MH5IXi8u/qfyAFNoZTbGx1PMpJcY/hHJr
3JsujRLnevilWiQ+n8AL7m+8JSTrhY4hq0qRsM24Y1C/RzJ+RhE2Ew1Whk1RIH8AxBzJcNw1agwa
RMq9lo3V5MojMwQOJtwWcSHgtn9K4dKN/E9URVHC4IrPAIojY5+isg4Z4yM0EInGAmE01hUVnDSd
kZys8ePEFnBYNlbkDnbM5KQkBEKwCn+/GhEDAKWjBlImb/22Rssjl/XkV6SiTvNQWD1AoWHhvtxD
8OEQ+8rgvntgCbVJKAeL6FeGZK5aGy4B2SC001oGUNp16+86MTK7ixoIHSrFjZKuPJCNiyNmpyNQ
enEGFQ+XRelrK+vKRt25mndTDiEgMF8ZaFGX8RaJjeMwbmT+r/dJPYB8r5DDtYVWLNuYeNquyqDA
P1t0bvEki0LykIKyO/DbcC4w81xDzZ8PHJaAuo9pc4xH/0Xgk3Hu8jg87vF+mRmKYLOBb1Q0pdxU
t3w0GByAqq4tfJeti0CNJ29VYXF8BgtZC1GvrKHB+xBRA8ylY/7i7OCvHUspqInREpaIUZATWyCK
C1vHriLreQevzbir0oFtdPHfGtNu4m+mBXcLO1nIncAQEYJaSRXsJPgJsa2iEZuE+SWlEQqOBy3c
/9GIISPzmdsKC/KNr2FWXedthe1sL34YTzEStySaMw2Kf/KyAA8fSFm3Lra8PsIwt94UtINhzE9V
/YOeLYR1Ru1TngUfqM1ZntvvPwDEdHPw5+vH5zkGesnQKMMqKaqV+WjhaTP42z79IXUF10/RDW2d
+A+hECn+3hJMkOX9k7F/7zBlltk864fIzUpfxBko605jqclM0R4FGyhfYnlALRAVVwsmpXp0zeQq
1KsXdCJ5CzUjhTRtdaLNyLx+AjwyjqcePI9HOaolDwt+D8KOc9zTfzqU+Bw04gucKtcoBKwEJ8ZD
3Dhv+2Cf5k7jysIWIbp6MfK+swzPiFkkliajk/ZMwdqwg0XmMJiDrWIrCwUs9d/qSnrRxkt2DClM
tncWi5vjdZM9vKOGpJFW/dyxWx0e1ldty7QaVGhCp9/8dgZcGPO/poi1Z9e3U2Pbfl/x1uDkUtnn
k0yb+VM+TR5ueqdwl5NvApjD83CN56AkJxgzdmBAVoVQ64gaB7BdTHRBrgB0/yz37r8L2XC+HGOB
D9DB8dC73Pb3iVaROG3d8XUWjdrfFUUjeT47jfICJvu5Vupr+TZOO2Q8Jem3NhJkKx/ZndEQiE2Y
mpdreNw/Ik4pTEimpAXpE2MJNCUABJsYNKC/gRYoecoISZE524kzhBxc1e4ABqJqi5CdkQEyL3Uo
ug9bNpVJCFVWEigb19vvfjifAA7EUV21NhAYfOVx9ND2JPiGmHh+pgYwZNYGv6/rF3trLp+pSWgx
W9mA0YmE2MlMDnfHafuvb8dt7JZ9We4TetN1t6HHyJ7KtgdDTLSLuX8bcULHMj8LbF7EUJDCqFZk
l8eY2Daux9poV+4uigyySsvJMR2qj0Bbqq7LnbcNC36jBr042cyqApkGgBlTUnF3JTlUviGqBRHP
pVr/gOpsgv4PH1mcukg7NFcZh9D8J7u3hNrusL+eug3HBf9joMiLO9xGkh/J7CQL5EgZuCJWxZDs
Xs78sfvEDAFI/WASNZKAs/GtfKRLnPaPcLNvpuzj8fZwDTpyz3s1MithJ2VL+L7ySPaMKO5Y6DKR
JIkewrhWdtCPbQQ9Y0Q7U7DZK0llM28y/3I0RUctnxd6+2Oaqdjsa70XyereHuXeZNhDpx2jwuCg
n5tOpRyayHW2k+0ZGM3Lwfx+ZYrJNC768/5vBvdgSEKp+a+ddJqdVQJMg2fdfs5lg7Qk5ErId/SW
v+p2+oSlpuZKiMIjxjnqyDQkvGcFZSnOGyGX20PStkbacag4aGQNr6wKrIj4tMl4eMrn/mcEuATP
SXrEGogEjmPP3jKODK1zfqVclQZHfSafmUTUYts/sidh7jxwSfYGEfjFiEL4R22Lcbnp87NZ7KNT
3qxgR0JOmMGsxUyO8g4tkRb2C2S/mcrihR50pjutUhRYt0Bz4AcgKSFWfZZiP/jpQIc7jpyuSRgG
KKH/3vIr+x9ztz9Fn/Aq5ziczwe3qpeXYGU4JH42lmHmnc0osin2ufuXMIG89zQgNuoyQOn0rqwZ
6XHskantz/OO8OSWipcLskD5CNV209sm/Akr3x5AC3ocWtIX6lWBfcUj/+7UgAaehITVi4Kah64E
oIDsdzCyAO0WhgVj0UA7C7AoBR/jqqGA7e2TbXbrf6x6Z/57KrZFcEpKcoX9gsQvuAonEXTe9oR7
OYPyITzdQsW5Dwm979y2VFW6ceg+GSnoN1n8cDtC5rIbD87IuuT1NohaE2FkKQhBJzl1S4s4ndRE
wNW7JDONr+fVreQzzulHSmRl+UYg1VEHz06ObMg/Y5l/cYRrnGQ0vHACvcS7FpFhimaPK9njzw/7
m8bVjJTKMJvEAa0rN03I4rEf2zEkZUCs1aWVidvi2BeW1g9D+BoXmJfb2HEXhfgapjx8la5VeBw4
/uW3tWBAhz/yjtmCyN3hsJQSCbN8d8T4ergTWov+DIKVYvCeucFULWA3saeJdCuTrzXsoKWaiq8u
K/x0C6KnNi4OB0c2zXhNBYYhfLeZ0bIVmUxjJ+Pkuwp0WWhaIZO/N7IZpPbLPJxR8M2qUk6XHmGs
0+WUmO7K6Bfr/rYRr6wVVKt0Y5OANIU3LUsdFSDpGAZJb3Tk+qddcG72jPh3IOSqLNF6zw1ms4HD
cywdovQ1IWo4iQS77H6tmDkuimTWkxbaAMLlpGM+M05/ALjM+cMigX81iMQqskoY5XbZeXVFJnm3
DJ3oW/iyIlP4hK+XopGF5tGgCixmeixsP7p8lxmKiDia3QKeBW85UamZ6+wwd4MUR7FZ7YrHBsXY
v7RScGGfws357Qwz05uq+xn5OU9l4LmYmKburLPAnI9g2dBd4hZRWub7WKbnnuKodFcChXYCP4h2
/Zaangat6C8WKa0qmvAhYp8KVEW/H8DlxKjgsMOV6cVHiVVSb5A0ajM/Fm8fS+iRKIsxfgbI3T3W
+2ssktVJ3AJAs0lMBeA7OiKDmFn12/gKeM7RmN1C/RIML9xG+3uee7Hur0z2CYIb0sWf6NUN6z2L
JdWfRllWaxHEuQZXCgVrN4m3sc79oqZBapOWFfUx9GS+3L4yo0GMLS4aVPtluGr/apNNKFaP2kPo
OgTvLz1HjDb77Cz6XsIwl04cmCil4NUw1pIW/qVkq4lV5UE/zDp4wZ9iRmLz5+aqbW7baNKBG0zO
nZEF3uw1vuUFdRYtiyf8jd4ZNRvHGK6hdTFW4ozLna+CrHe2XeS0ew4p9NLY73oraQjUK5BytvpW
en8IM383c5uhfzD0XW3bynLbJLPFlDg9PhtRjTS+xUBDOyrZTQlA7YLkruyKIe8ZwocPBUeY4v8E
DpHZ0uSJGaznLg0e22EHvMq8B2SKfIr6FVqrazMrYrOSuGtkTMIzTj3+2NNSa+1n26WypRPEuc7Z
wfSygHYaynme8WQg4p+d/t9BtsWimxGfHsX1ZqnibjAm8s2bqDnz5IqLVC0xgf9slBuf+i8QgLbw
jCbgDHGnYgqf1+vQIwKmo2Df0fi/yYWvWpoBYRElkfqUw1wL0OFu0Kko9LQXCr0HVTQCYKBN1FsL
cEDhVq8Pf0a8RoMfb9WZoBjHwvt0oyuQBEOgDCTjvpBsHXw6Jh8ns63wWqGfpeALWTaG7fs+B2Vi
BsulBFztvA14q+yoRl9VJ9k++HnznPNf1u1WxLVoEidm7PmuU6H27R6wP4dY9Z128wauVQ4mjM0f
S4a/XmHnK8FI8nSc2y7yub1jx2T7UQfY8/xAP56vXg+tZTwZ4jm8ozBZZMiFdTG6w6EFWcWNhTES
pnLDUmF0w3k9usghzfHGABYu/+ll8z7235o25h00L3GZBQclU+9mFyjqYyPNV+A81FTvJsZgMZZ4
QO4theHoFd7Zgvyei4Zhi5e3ZNd2RkDK4pxrZvFngCRoDHBc0knUfH2GqrK5HjB/URF3VnY20Yxs
zT3JeUxd75wO+Qm0dvb+BGz57aVLpHLnmTcOR+ny5yuezqKqaXHa3eeMPrsPEnJrnuwU7rz3N2/2
0ETl546X4vXqzafAdHy1TN8oKUl2F5Xpiyqo+nedHLx2jAW7N3yj9wDHp4ZN9mMXeEieI03pO8ah
pHfR4qsV4BAK2PqU4STMY2QR9XuYWkKjZSAQtpNx296fq1qI5Gv54Mghjd/7TLVvSXNbCgiHk09S
payzDVTxeIjrmnsHw+mtAgjx3U9cMKBMRnWEt5b2q+kFudjEMv8lniIW0ynv8rd94nE7gB71xKuk
k/mYSwcCg6/a7oklHU4Slb8VPrBZkzEeUZ5GZRaKXozs8jQgkU0Kmk2cIvqSxvc24PHZ/wRr/KeP
o92OHaTyC78vF7f7i2dSUt9JPSdW15yLmvi9s+RxvYCEPglPIpnsIwUnmS2knXrEo+ic46bYzfGa
HclXRgMvSsN75/n5O7nBHVii6AnNgOW1ha81pivoeKipylSdR03EMNqcHr+xxKyY5fslO1Hqz0Qt
h4Qzo8Jaf1QIq+PUl5e9RcIIt4N9Z8jMqrfTh/88tApLm9hyNGHRNgZDikk+nWEtOKNVi5TrXMTl
UVJF4QaKpf1Wo+2Dx4TkV+QMyegpfxXplrvROkeHhoVO6sVnz3ugxU6Yz6xgpjCmrIr4oJ2x0jWn
3vXplvKjlk23sWTlOWicKOaNPf2JW1GLaaIcI4/cn//g8h/dJIYwkOfBi+N9DjyzlB81HSzBsqus
hP8SLd6BvCQllIUV3E5PN+d0/689XZ8PXWu0rQ1xrl0TkZ0Y0sIb/8ROZO8v0qK8k7dA2biozWjS
5vKFGwKtEr/KHAtXptvHMF9d+JSodrLGKoU8qppjVMtnfYaUHNjciMwZQLby2VFP8h0M1vq4llWi
Ek+gufRH36KypALHnZl6kDHv+yM2o9kyziK/2bKBmI8n6x63UfBwmoJhf/TR0SRQ4ANrV1Gjng/R
quqCvDxL7dcOOE/oGgHZ+whBj2qQvmlVDIkhcq8kw0h9JGElkkwp3GR0t1VwdyhaOTghfeiL3hcz
bScg/w7W6QiVmKGUuY3TBUvwAv7lubGZtABP6Il67B7d/r3muUyhU+6YmPFCXCZyUOgZ6WOdXqKL
MqxeW3wKzQNAZxB+0e4mdGZDSZtbza6m3cp6xTqSSQZJ9pu3oHexHsQuzkFth45OzUB8Cppsxc/+
2rj2mnZuFQ7ZOQqcFV4t3zL84/MvukqbLbyn4svLBafZCy/rr9D+6wIUlgiDGd6gyssUdoelM5Bz
iBFzdWEwsy3gfnsd1QUcwcmme6aaPV/LdSbk017foN5oFxjJGDRYN2XLKuobGVKI3GlQrcMfSV/I
9b6OXRBtu1X1meI8kGJQehCZxduKhTcaiin2/3blGA1sS7fIISH3rbOAPjBB89DgthyjvlxQvt5d
kDDeGglSHOqY5yPb3QONw3tujb+5uJpzXhtgznFLxGL8RdI79aS3wvnXVAmk6GPHLe+lff4U3LRc
xmn+y88QxLFJ3Gkf1I8ZnVIDJo4kf4u6rBvUuY+JXNHpmL7Sdw5Xqp71smOakPIAp/VXYxwoWHO0
8ZuEMwyZqSgIQ4kk3T2zrcV2+nKE0Vu/JerBLFKkBA2d5o9TIeLfvwsiE/53tQQLlTXrxSBaCeGr
PldTVUcfXnZhDSvFYDU+CHzX/QdhwDSNKCuE+JH4VlMdNDeTY5Je4GKpFZdiryIFvFGqw4BpcGDI
FkVJ27p2bie9B7wNCb1yWEozdsO9KMuxbeMMZfHzXjI809o8XYeks2o6gGyQxA6zMBmJAD4rLQ7t
VNHomtKjzI8d4ZvSbSMMLKKS3BJbfb6F4UTNaAtPYMJSJNchV45iKOoU9xa+ayPn5nKs+XQOyEMf
QExHLQgfNs1qXHuGiEgyatGzh0YaSTYvvC6iEDew1nInQLt3N6ct9xs8FEJKE+7ilSSUFDjSasva
KBRKjzBZ9VHvCwq6Ap7JuxitZ525uGmoyt0VmOUGpG5srp/McNrDY8EwBVV/ataFjOs9DRhYkL/r
sRlm9OJYU9k9qhxvMRN4lKpCoFcaaXDe4JR5O5VI8HBxF8S4T9qnKz/nz5GIzhmPXMmHDyE25wMf
3yPOtPMoyNhdL8WSuKG6NxY4eBOF76tu+pABMuWNket6w/Gv4S8C/ozlZ/g4O1myvqdHIbCaP7g6
F0vfKTJyqSySZL6A3uw688aLvYQoPjdnA8Vu5GRRx10ew7ky075YQbZERF4tjDZR8H3CtZViR9Bt
BFiPvjdgiRLAbNhM68JjGCr1nbJi2bT5ndRjDO2nlO+btFGQX9hvt1baU9t1dT24dqpepGGeBAPx
degh5SVZON+/W8kEjsQbRa2ueRWWFcIsmGCgRzInB2y8oYX8uG6ZH1kmZUTi81sDaioG3FdiSu0R
5nxuSZveiITwer8nFuH7iqC2X6yKhbUdAu/fm7nnNAGP7i2+LrF1SOw3KRVk3jiCBTfOaa+8knwX
UlKQcPdidnqYh2hDVtqvQ3GTbEmRkHs54SR0RSU6IxFNqsbAzCR1IIeQ9h9loHXmb5D8/NgHASNQ
Fe3t81AOyqsy0SAQrYOJR3VmK8fBBBtEvKe5FYZPiQRdwyjof0QQzmmv2lKpCopBOK7tDzBtGxQa
TF/WIDYlmRVv0IDJJ5gXDl4b0PfRRnGRM26yBZ/OdmMLuSiGsB7NWqte7HZRv5+91oYU4iaGlWLe
BiCWbBmSWn86Q49u1cowM6EeaScwjaX3NfQ54A+DHqJm+j2FQLkQ1gXRqeR35RmSER9m9UnNLKle
c2Td0ThLIfW/iOJqHPTmxGEXO3szB+E6yJBVMHQAwGtVheQCvvj8h8JSw3mg/t9TTxtAdUhs5+4C
70DZ1McrYqMwdIdrlgHuzoFAEu4GS+hp6eudE1ml2xgMYH2974ThfYcLw8bb+tOdysMyvonKmwx+
ZNYRFTIHYlt3UUaUx02aWRfs5ZNnjZ/uZHzWZKzodVk/JDWi49p0usOfqj4UkRJgD7S/jpyQ4Pv+
eZ7cD91x4PYtJDaEMHarGwRqpLLMf2pPG1JIbxH3yeUIJGoGGf8dCW38wdy5Bz+FOIq5wfZ45rK4
M0Y6GI16UylmyPn3n7F+wdYBXZjtr6kAFw9s8I8DlUyz7czEW+mrS8LwVNxUbKMvEKb2vOwcsVPq
TDZrKXoXDxb9DHNe3yJYPMjW9vRD2og+6dakpXgyU4vHfHFAGISTXyE0gR1utXdQy5qpC7fRz9OG
344tW0FmrGmR4CLKTnfTxXparxkzJXlDVPP95uyWpX1v0vIn5hBmkyjnYJbYupzNp/OCSqul5rHg
XRDg+RY+rmMuDeORjWWeDt4KfkocUvfvFQ7wMAjU5zgKHwpWRtVabShDSLJMxr6a2tfPt6wcAAs4
L8+UFPLRLDv9ptAxvna4Ck83t2oR4gUo0QrABfnx3WNNGhmpBZDAcwm5qgztD0obIfbOsLAlwP4F
rVxxfDMW1F5FdnTiXDhJNIhRF0rwScUDMzf5460nsS5UPUbkNIToi3m4+0lPknrdAd9hh1y+D4E2
+kFmai0GYnCcciqqD+GS8kVqpJBkBUgfBSpbVBjfGJDmJRRbJiQwBPUInRi6FJUB6tpSQd3+QAa2
bPkXeQmZ15dL4KO2eKiKgk8BKqAfiBw5c3pkIAldKj9QSi38mZDk5/sTApfmrWTUYcyiv1zUYIaB
m7BnmjFRdijSxMD/KRPdErWYyBfID5/z1P0KZ75eH1aD9jqgPGngTIyazByjOQyMvjRsPKSwKIcU
mkWo4WVSdrk8iZck/84JMQ+aZ3uVgiK2bWhqFFBhyPaiEVI5eE/pV48GNnpqvVFW6orLJh6o/b03
dJlzotbhg/wf+7b1BO0SV1og0ScZm+h4zU+er6HVhuQ7kGn/8zbWNSS/e7QfVTI+CzIdka6PjId0
Kvn1RP8QQvUHH0PjYyfHCOE6iYcu/9AFrvgMjeb6QbGe+GORpOn9Wanqy0bpb4JoFUhxQQ7yzsQh
pYR68tEOwxe3lLak7koy3hKw+2ePQ0PId5W6YBj5S+SnDrhqS4k58vmMCMdgu49s1fqtGY4RV5/F
slrewj56PR7/Ikw9VuFTf8AdajoCs9Ock8jhReh082k39Z3UBVdlJdTqU94vr5DytHxm/PiWiWgA
9ZZxyy6Wrw2Is3XeAIvKDipgsieK5j6YdvnOQgcClH0HXWdsIbrUdFeXsuVOnoVcz9VJ51uiEbPV
w+Vofd1fAw2l2P1MRPmO5oWog7as23CpYYvfzLS5PtPT1sZvCpXs+XV8OWlQD8gA7q9unu3FUK2m
RoZ8INQiTh2hopIJcnpVEKeHdFE87FsKUkioQL0GyNR/VQPu2kcF2nQcKyqv2JmYojJzwFGjk3lV
2kdkfQCTenMDk6PEqUcl5tcO9LBNRpQq49+bUzVL2SKVSuGArtpA8un649nwOcfoAFLl+PSH3Jib
d9HQ3DV3FdjoRD15N6wNVogdJV8smHI4+9eGx1jXFfvxvFf12NmFrGhiFzOG6w4S4ev5+O/bzc2N
Q+wRI7dWt4wn3mqt1Fgv5FSl8dylQNovD9zAhf4AGQwfOvkViG/PFHCzLAhCQNkTNr/BVdoD1D44
2HIht369R+ONYCvvyB++FbE7nFTUFk8srNQwN5SokXCm/pT+r29X7VJydNnqgFI9DSHt5eh9qc/u
uyK1T10YMMHEzjgtnFHBOw1p742XAQxajAxCPUGzXGmqI/ZWcJQKead66rsSsKKXd9qOY++wmVXH
KFVEOsLsWMiYXXJtr9fxk0YL9Pl+Qs2RPpvSzZUbXAyJRdvgFCZStSYjS4aNYUoS6u6J+icx6/6B
RwY1WNgrvNKRfK5mKGEJtxuiUQOCtv5lFcKkNjVcVd41+XapOvt99/xMDeYam3vlvVsKU8AwFgJS
2QCLs2EN2R1aW329qA0CS1GBf0cT25K2Htp99jTdD0sGXNWaPAeIcHEke+uA4z0ANHGmqYgW2+c6
c1HMQHTNzJiIbVOz4CK6Yl5TMWzDinZjy34EfFrW+EqYgbJfTGCLWExY64jv/Gtg3LRB1Dua8mtg
EwQUYpzEyfkK/0zQy8UeaOvF/ewGUz9VpSBD0ka6WWGCKdzxzwgJpcv8uMCyu3mAWZXqvdyNgS5N
JNcayAaWheZhhKhV0YxizVCbwW7otssyMOsryepVZYkfjYs+j5yzSU+i5N1LQMh+jlftoNjJ0APK
Lr08yJ9U6c9ULhLjlSDzJM4Zq0O3lT+XFRGet3jsqzq3GjZ+VhgXi3P2bmQfMAvEgP2MhO7hfbt5
tlPCD+McOpWNt5IGjbAorZIUGac5xTsNdZH3WSIp8ZJLg7qBz3+01SEsYHimmNKMEW5028CqyO4Z
h+UNuym8QX+yjihf6vQkz7ZfCOlxoTyDbW3/odF3O7m86fU/IauppwcuXCpPz5GrUERzsZ7+UZXk
bQcJNlBpXczQdjRjFyo3VU2fehQGeXrXpYR1wCoaj4Xq+N+w8pSOk4vydBsUdd97CKN7yTUjX17w
oDFuYLNmGQGEKESi2Zl0ZSFx/XwSvPZw9y7EwpPNjMEDjf2nafO12t4/yP5fc4r5m6uWynfqzjZJ
5gDaE/mARJaaZQi3kuDrGr2mlI2xGz1qvhXL+Y10fLoRLQwqDlGRtep24+Uc4PkL6EDJbWFhFmp3
z+udg3SmEc1JJY2fzXzWrh2oJvSbpO0Gq/SEAeNolKm0jRhsppWAx/Ue/FWMyEBHbK++VvHsCvcy
uuHeT7DNsjIOkAc8VXLQRwprMoTtWE8eRqRVgplRuHWshXtR3rXPB2JeRA+9/PItheJVT51OoAtF
uiixO+FN70Dp2s21gByzCSbgbXOuIR7dm5dIMWCmIo96hAb1R8USMa5arVC/Mme4auXq5kG4uPe1
af8QIcatk2rGC8OVFIfF70bqyX68LK8FTkfh/tdaqz/0btUrj9zDLx8az9pei15LSxwL2pfPCyR8
8BEwi5tNP+nSvoEeLaErtwiS6/TkpYQr/0aFthF001HiNsLMl8zZ0ndLBq9uj7ukBXv2q/P9fj4L
EJBXV9hl08mq45LQ7amSDXiqh4M4T1m75k1ySTpxXezJnlcKKDKFPOuqneQ9IHqavYyk9YJXLf0E
vR1fWJD94v85jQOrIBGkN9Waa3AAIxWul7ZvQNEoBuX3IWhv28uwAKWJ3/qqERyAmH9yRhtru15m
QmoKPt9PE+SyAiEma2VuBXcJ6Em6tBFhzBZgN4f+XA/qQJ3hklNkacM/j9zvjAmJavh/Ip7HOUNR
7QNgrHcDahg5QtOYqidel5iq8SaHz0dUYyxC9oRa5JFHTlManCCW2HquEH08osfyZfuDsdg2I1Vu
cI9lVF1EUX1r0ihC5YIURUalReNNI+BypE+QNti2OpmiAs9GpGwaMmTdokj176KQj9BwfoC6mcLs
b2NbAsN2Y+udA/pdH/clYXwQA1SqRcWcP5y/KysbZlscpPTbV5RGd+trgI9QfJbWFtfeq8EUtqf0
htrXinwn8eWmQSl30A2yD9HiowYkbfaByskOr/11852Uioc0utpSiSaGkn1K86nMxti3C8Nk18/N
5b2SLbuUDhi6oQG9H4KY99cqu7ggHNBGH57Mgsa9iJeF9xVJb5lGIuzeBhdjfHS07AHmbu58b+AQ
uvx+txbL7ES/6Wza3StICD4dGfSOgH7/G22/XLMD8bFv9LXaAoqn5Hv742VIj/DMaorTl5aKB8do
UUst09r56gaiAmVevnKDozq2F8MZ8eEeyZW7nvIa+W1JuVVnkKTcugi7Z3SNkHz3nlRiHWe1hcQ2
E1ts+j1hayBfI30bHnonqChjLF1G/iZDBZPL/Su3zKIm2juOBEdHjsMXgwdyJ3XFag6Az6ihxaTs
7QYKMVMOJelsFnyTYxiyA4jeKQ+RyA3uEMrqXuyIRVkTj+xk/ML4gDaJveCZo7fgiX3/fRFeS39t
gNvXYCVC8PjKhUfVtedCbu/5LolV+DdXFocxSGhxrBidgNFKu7qAh4kNMZsY/crylP4Wm82DEjrY
MZjUNl3RYNPett7itlsOjsdcXStZqI8eC4vj5agrVLMzDNt7ZKVPc/Jt4TUMRQ4OWGx5pWdw908C
eS5BREARumh+1w0qaxe22309MbEAOauytwbrcz4pSDG6l8Xkv0prM5sIUZBnZmbAv6/HSGKEERqE
CqZstkFl6qz5Tg8nlY2eA6XTuuSFCfAwEF2u7T81H0at5hmLGpuuu+5l3ttUOH4CrIkbQONm1HcI
iYSOHNuAd2LGFvphUn5tgcfJ+jqKtv2Mt7MOH+BZSPn25D2NvwYgYaHe+0ULJ1PVeFBuFU9iJ+iI
xOIGTWCBvcFIhXYJEFWdbOYFWFejJVRlprBN9PANDZfYxFLXH/MhtvnDkWs7nXF16UdhoI9FivbQ
qUaxeu7QsYuOVRU5HJ27K+m4ylUK+w/8SqwDd+C0YRkR6eJCqYj77kCA1X7FOl+WVmzauXmhjIuN
jid7s0oewm161LFJBEAjwkzv0PWntPIu39tG7epEjE7S/UjvxNl7CqCnlIvD5nlWJ50vpv5/YE/p
eiUDCo/ByBf2HUSpIigrVKItEfMqw2FwHmyQCkoVvlGvBPZ0jluvX8GYAqtPBSnNlDoxcxWHac8n
5jYQBlLXFZZ96dy5f7euPNGguy6ty6SVFjxWQArPZzDo5FmxTj8nGIWSyXREqHrxSpRO5ww8xzN3
zobm0pUVZeqnv3IPYosi82dC0kqAhSRH86I8rcCzygLfs0xGgImPfm9M5mtj5ugF414mDI9yBU2c
FYGAT+PpmG71dvoZ03RU3zDWRazCkjNYxpAAYglE6d5c8+V6jDWsNIIgsxE/58EpWMmx0lZZQlzk
ioErE3j9ti5H46Xv8+XAjIJO8iDrNxrPRPAPTrj6F5bh9GPES+ORUUq5pjL6WK99/xbnPCwtj9eq
hCoHF5HmgPm1DmUO8X1xyBOi0k/imh4119JDoMJQ5pCNZ+FFvAVbpFkFARwv8w0GtGkqHFJCT1+R
g5LqueVUvOaRd3bMHxTeZHOeIATYrxxqgXYuTDR81GI0fslqQwHZgGS59S3HLWW16y0eFAwRCKFA
ZjOJ2PCzFvKNYu1ESZuxaDXLn37jvC11nMXFVI8YkZleN75Zgmr+R6jlSebsMIBUSwz9nH6Dp5Ol
shRAHqKNPaEW8PuUb6VVA4xP0hizUWGE5G9VTXHb+BF+++y2dmMe2Wt/Zxyh7KSh/HEJoujmGw3X
KVlQvKvVKtjwUCySRLbdFpFpXEQkTsOYsKX26jt52JOgIlVrDVYaW/HpXaVJF8Lk/ii0dhMJcnox
v+sUHdkWztqNL+OVDILXj5sAtVsZiuOAYJtDVVD7FLZt7MgBiL9GBRh5HsJy5iCquHSSiE//SInB
wWrYaSt3jDJTFA5gAlz53xcgtjuPXcYuYURHUosbt/w+6inM6TmNETpumby17EBr1wpk1+tjM8Jf
jnmTT8eQQGDTS6ZMMmVav+pZT7vPvdoN4NLT0G9ltb7l2zvtAFigUEg0f8A9Kr0khMUs/O9DLHdZ
h87FmvoVPBb9R/yoeT6SuNPJzurWCxYdOk9v49aj8eukH/ohg74NFErvQ0uj/Yeo/X7LMUo2rw2c
zYwLkSF8Jci0KWQhsoAO/feoxfgM5xsqgYjihxWREbqAV9eEZc4JkL5UeZ+IH9A2m0vioQLg1sDX
MvGDQBzV0vwckDysdQxyDNwTqfStKc2TA8T3VQemP0H8bVOIQzFkrdsf83MU1LzqKcHWSCNA6MNg
Eaq6E+sg9QG8E7Z0i4FjL86CtXTEB4xMDO3QjwRNyVkNjPuqQtCXSaRFfcEmKYT/DQ9ioUOFaFVi
Q8S/e0JbOuToYHGxf6KMadrHcaABZ4O6Rq7LvX2vl4knBbUybr6OMY6nHAGED+9UF1aFSpmaJ2kj
nY6WjPtNaaMzyNeVMRCDzxTnS2Rr0Y2xoCeT/MLMwM0PpZLfAq5Ml3usLzJtMN6Rta3shzhY0Oz+
avD7/a9PnqMdAlUyg0i5o+9cBjZa0M5/AsB9BcOLx5nFeq2YTMRJ88QrZHO/vGozAYIF8IwQP8sb
7BzQ/4vso3V8RZZxYYkj0hfvHpvrw74v2SiW631hCnKGiCvppZjG1tUOs6abXEEGH877vYsU1ieC
uY+3PZ+v1zSatxm0/klG8eLcMam8u7HwFHe+ORZeCoV7dNl3Up8gxvzlHKq1sp2rtjswR9cejFL1
BLgM5s9t9kN9OOpGHpiU7W7CPvG9bbXqWgrvVo8Q9OpA4hLGZ3sHJvFvhHGqGPA7jH4hanrkRr5S
U0QMfVrLnvpANG5XP4rahadMdaNZSM95tEtXTGibkmx+VIjL/TD+qHMVN4nZmT3GRhbDznLphTJo
5aHT/9PU4NxLOIiCdYYgi28sesnfas9uU2eeaufjA6PwSDuvOFnmoUP3RssbrldsDgl1WN8xvata
aV/UL+UiiOEZobGbCvjucqiPiQt2UZZ9S1anNYvfs6YwAoRTi9yvd7oWYU3ZaiZRwHDHKWF+CDZh
1txvYTxMpeT8JVVCnKaMhlksh1PSscP0q/S6ZuyVt0lj+ItR43f07FR4wvY5NqXjAhm+VxK5qsD7
kWZe3CDv3vEAoXgwormhuZgP8s3y9i6PSARuE4IDS2dQCuEQN2FltrbPj+s2ZoIy+bb+S5tPkSZ1
n/HbMKf4jYKqjNaOrc9C8UIbtWr5KmM6Itd5stwRDWNbxlYi+AjJgfPkl1pp972LWwHqa6xj1Dzy
G9Ezoblc6dFrZkOET7LwSis2K2Sm/w16cV8pJCc7gdLfheXcJY6w6N0Pb4XrrTXegDTbkbFYbRNh
LPJ04HeHDiPhK1X4KceJRVHq1H5cVQGlh4Ta2gapVcJxZUKOvq3somd90peSrllQSa+LppcUIFWU
1Lr7Lw3wy3Ufb8GCybwHmJrHmkOa3AAIRNdpzDE+2fgMpbIu5nZpYOg/1WYxVtE2LY18N1rJ0/1W
7TwmGWqp1a1Ihfrmp9Op5cnh7WoTBkjhQ22QSTyY5ni/UU4etTCcq/In15lK8OcB24Nevz0YOPpI
wNGfIlFd6UYkjNqykgDpumD78kAcSFc1Y85Dzb9fe5Kce1+wwIu3G0LK4tXYfP7VBu6H02pdyeeR
bHxMk174EnP9+e6M5NytwhklvZGDCkrtHUAiD/KfqQWrVL+AHt3Qvc2f60P0004HhB4OY149p+rH
5Ek0bc5lDUqd+ASFprNp7lz6Hsv1G1M8YJormBgtlIYThl+j6KrZ6coeYCmsasplfq2Lt2d76zxY
3uglqQ7+2EAnQEv50hB4c2rxEWmr+Ali5XBYUHEj/XhvjcNavfwciPHrkOO47PFN8aFxquv6Rf6m
9hDtuh7ESpHAbc/zhQPMDmEG/0u1+mKmn66fKptILDonvQG4Kr+mKQ2hn+VD3atR+UDuAPie2HS8
2UCj639tQpJdxP44OxVhr1Wwyo6eY0QBJAOQM2M5D0b2xXxN7+AtOJ6d366WtX8yqig1m3IiJEaA
PzuDxaNq7gImbKFfVPllVKXfX8eKKD84jiw0c8H4tkS04rzUahgkxjtzZakEAIPWY2omk6Qy1doN
gXX5h1OYX3pujvYhS3fHdLs5cvUvq9GPXj97yHA/pH73Bf9c4qxyvrfKBS08MxKdaqd/7MQQqkE+
9jzb0rAUzZvK82AcUdRAHuFzWDerP+ZkWoRidhCUEcOuQ76SRAdAYBFykJt7NHlRMe69RcMxDHGF
tkMCK+X2AI9iobF6Mj3nKEZCL17hF9+Tg7wY3jHdFJmV6EQPNp4duEUi6PIFu/A+5FDoP4R3G4+7
Bgxz92F92CFZahZVaJlUvVQMUxt3TBFNr77WJ2p+ROKjojn6H4ffR5dnMDUdtlLdMqUKqHkM8BAz
JosVJ0i3rLEY1bwz7s6wD8/QRHDQkkM+X19KLs90RM1zFAn7WlJvaOLWZ92qohLmQhRR4kY/2Oh6
6aIcj9IYTqUBsdJFadJIaWDUwLntbClJzAgRwPb+1RNjYI88Hgz5tDd8c6tO6wmXm/Uu5pxBG6FY
STzDSpA1XsPchbw9j2nh+tVnzQADa0Y5aondwThR07pbv4MR1oz8/u4FQqMD20bXKe+oV5Mv+tfe
3+u3KBmkMwRYALMXVvIm2ViQ0GbAMVP9QO2wmzVfqcg7O/gR9QGbb9mOIsN3aSKHxAMJi4e/EH5n
oi7/ZU/tKw13jbo9pn9R2/2e9+GMKg6ASotO1emL1LUgl8YFCeZOj4sOZAsVa97AhJlWcom+Q9Jk
AiquPuq7aBEP094o8K2RbabDGDz2kX3No6FbGHYjJQ4gwkLBngXs4HnKiI7ydRAH9eXljfQhNiTV
1etpXhR/cZneSpb1yTj6sRAoGekclxsfWpp+ArRciJ9iBmjO6SWtT/toXoPWPPTZpddxLYuI4JtI
HEaUoHx5GUuBLOuLSBnElghXIfriKzL9KvDxGIzHjp2YOvQ79kRtXL+wiG2kZOBaOjH48dWBctRZ
AOPD6vi5bSZ6I8E6oVKuKWmYJK0l0AGXT5KiT1DYRB3HDsAesoVzQZk4PPBNMWFTeiu2VdR1clfJ
c/EHQUHLoPOwT0gTF0cmXxhp5eeDwg41MufxyYCCcrLY7YusLam9+z4YCb+hpsRLlSgjYxaGozG9
4veImWV5S4hy/x/lPeEVxiIHc+GMwMS7PwmLnuv30NHp1gOKoIaV9/YXyKiUk72qDefNypMoeIm0
GI8bybYPMaDPou9IAHMOmrpKD5UXkJl033T/0QYtO3RvHpNOo2F2e4RkH7jRnwshG25d1hZzGOVE
3l96P53stPwQ60ypfei+3Szoa1tGBK7RRZn16GSqHp9BvsmHahii3s/ZgWMnPN/8OBDq5NxiS/Sw
mMKXhwCmRX+u+LrvWtvXC7Z74GPhfd3X2Fbf4hiCN/h2pk6DgdIPkyVU2FRuux3dTkRS8e7rpQ2a
zMf54tWWk1kpskDrQIeb7oGWpjRhZS5w+FeEIDSdFh36pQbi0shXfhiZLK2P0p2GcnOxnUKk2swQ
iDwgJ/bOB/q9ol/m3VwlyqreNFZx68HGRoclO2foaSKd8ZB8YZ9pGSY5KP8OKQG9fEwr892wrq9s
VnxIoM+7flgn6d6rG4Zail7HcOo0F2tORrdcMtDlV8CiSNlMyh8tNKJU63adOSdhvvtqPKAYwyHg
s4kENNf9RArKVNC4cSe1sNZb+KINCEbSLJhflZvHsZp6ItRRdNzARQOApUytwNVnnf52POReDfxb
ZRclzKwW+EFI5GJT4FYV4UvzuJY9GbRcT5OUIZd2wsu3Th12MErX4t8kU8f4UttHnCaC0PFeD2sA
rsyAfaFp1o4BvJGiH/xjoiacKPCFXX8jCx4WYRT5+c27RU+DfCgPKxsj6Ro0B702NjiPNSZ6k6rn
jibKZqY3IqP98MtrOi5tXRP2PKmpcKcGxAGAz+inSDGlZxuS+R6tmOdZ+uQy5nYdVGPHdeavFHeU
mKqdMuTkHho2g9NVKLW8DN/evMSHXTFi+ebj4ITaV6ghFfT9fcFFcezqbrHGIlfC35gJ1dVPgHRt
79/wo1JYm4tij5mcl3cMng0l4LcVqrSXzB5AqH24JpIIn7gusaK3JcbD11Qyw76C+H4t9ESOgdvY
6hgRKQ5xGOlqDL7lDrVvtqJUIj87/bQHKpbSA+2vgdN5w1e6wBRdsM+nP29Q1wZOLp8d2ZEa0U5k
Jg+0PhEuqyCDkX9Ub3/nQj4zsGfNzI77RtKX9+dzSYoVelEIpipr1SIvAmjqg+DVGetVEbhSq947
ijOSbEYbmeDx/4cYGjVi5/evXC8mv0829MBF7VSrNCDVjSlP8gv1qek/DfjxSyDgJDcJfUa7XuaJ
LqcoFi3p5q1lJCyi2UBdy/eD8jEuQ3J4sTtWlVTja9LCtl6cNCTyUAORzPdcpPYXdwr5a9dCp3UP
54++DiOgvgJhugMUwSM2u/JEJ+BVAlW8n2Ok1pq56R7yRyfUAL1HjhZZNMWptty527/VRUyg6OLk
9RH0pX1JiqgnyiNaoU386llgPf06kC97nlKvDlC0BRqRrzVBZzdad+ijEgTpTaBaP5dRMOZ8QBq9
mpBykN2v46+php0ehOEm+AU5iTfSDfdlyFutcFOB4FWgexx+mHRVB96fTiT/FRXOP7FuygEECbAI
noXs1JtRYbfowxm5JOwcZnz2sKhuPfHPYYIPP5GIa5Qp4MvgIiH18bDU74L/f/3pZK9Dto6N5zDP
FoN0RGG/U3bMOLI+40O4bb9Ei6PQkKvdObGZbwYn8kPeLk40N74gckq5GG6xgogOtVG38CilAVGP
l1HQJcap1igMaJcGfC4yj4QY+WwC9KWBg6WeRVZeOrqt9rToQlyURIIZSGxQZCDTFC3tOyB68fTQ
rG6DhMxDtDgWU0jdyaghS5VtHNSDVd5AzzXnzL9gAd83jNrSfimO1Nqm5o2LJ1gg3juns72Q84dj
+anRyHguoWvLtYGSi3smJHxIL7g0thI3+BDhcc5CaPdrVs8e6W0/Q1U5R0PwJx1ViY0hU7e06Jwe
v2lRJidTrGZz11BlfpuyiZU3E8vcsdkrs/j2eBCgLdN8JSa3vjust88QiD1kxRWyJIOVKfMoE2Vn
hMdjXUQHNgWKB37Ec1prpB/C8H8G/IeaneyC4a7WNCczdxWgoJqeLQvj0GishqyOQXPDPIMJNyud
GZYAFz6tz6HY3ODN9u90N/NWZk6uGzcTcsBNW7UND6i7qRuD1NOzkI01bksYish9AMDBx07XvaZI
MkkVLJTBh7R9bDIRRYWY72kqGWbFEm6yQcettJR3/EWPjMCUejbRsihY90NuEei8VRakOmWA6cpk
tXJazcEGdncM7luc2iyLvuwQHk5zmp7nDa7Fu1HXkeiocY+IEgkDaglsw5QLTVbtNOU1jtLj3CEm
WObkJn6KQnkfGJ8CqdeXhO1yYg68CNDhHGJISwqL5gAE8aYkd9HKk5KfYEljJV6oM0FYaNMndIIn
J0FYmg3hDUyadpc+wHahBWA4YtiTLjGqoB/hvq8tBkyCJysIzBAOoQ5he5YALI+caVt6mgxNkRWp
26a3m28cO5WqWGlxXde7AWTE6ZZ8T9Ge6jjhMyXG/3M4sy1QIqPvbGUL7dQSYjzbNfU7PF8f8CB5
oTops+P8iYXGP0ui6EGtuokitFRBhggHLDOfOa0nnr/ya0XsQUupfl5L8FnTwnLhPThyVSc9RQv0
a5QZp2FZYHiSFN39uNknSGR+MPH2xEPvpAjxgcCA7Pa1vX3wsJIdrrN3JPSaI//kpaVb6hnbkktb
r+NIxVEcoARktRffWAQHo0vbHOphdLjWXzikvQnLq/SSHI0rI47NnLKxhJc3KsybQ3nhDAK1O9TN
25/dOco9YbxLXpcdMen2/9cakK9n+sH9S3g/ijmTRjmhzeeuyq60lVEi/Pvkh/XEfqO44lbi3/TT
TgEISZXe5/91W+9MTCh4n3c/KZBxfBhiXoGXgEH6mW6jO/b0Rux90Y9Bhul4ha5F5NnOJmpDI3rt
3FOdvHLlWBBUHDEjugu9/gt982B/VUk8AVLglwKOig9M/2wEMqRcxBt46vAiTs6BdWvXvjrK1Vlp
0pgmSMmqIqhUqkHFXTaAq9TcACOBXL5DRmefapn//OWhdIN2dVImNZSDY/+zIRkIrJdGp8hrMD4v
tVRXTRR3AH7pHd9zyK8O3ookZO7N5VRwxyfJC4EAV/gRuxW+qDvm0wAc5ZKTVThaCQPaAaz34JxB
nSdporH1nKeODmMxHiN7MAQY+jqjEdX3DVJig55BpBC1wrOKQRnG4DiKxlLr6dxzgeJfWVOMdTuG
YUzMA4fQDKuDj+VVPzI/SoYqf2mH1UZk7wx+VMBor7SdC4pybl/Kc2k6PRHtcE2DKvOBZlkf5nVA
iwsxXXk2yn7ix/N1y85mqg+1hOYrxFg6NCsVfqV8oKO55Xufjqw3kcTR8/TLcHzJTlrMuCpb8t/J
yX6Op9/w6nJnVmTKpn+7ZxNj3IkbF47m9rR4tr8maTZBNT4aN3YX0UGZiYbLvGPVdanUb+p9u6RX
FSDUry2rJzGnbOaCRJCElFWIIx9C8ZAHtfVKfsX78G3RVSdsJePslhD6H+iBqERfnvhubbcu/6kG
D6VT/RZV8SMCOSUE53x2kWTEoJyCkJPgV24KEhNoX/6xFbx5cHZwqhV/FYQSqE4aCGHMUk7ggIz/
gZlKCX6I4ec24Q57N0TOK41SzoRbCu3HBA1DCPtG8omol1Y4moHzyFlzlNUIoYG3K84fPIqDQw0L
B0+tojJ1eZOUPu7e0L6//KuMkmZlCRfT6cwBDeTfPmsrADbjrXY+LCACMPHDWxanP2x6mtQaxubD
6H7fXNrORU5UpoRiZQwpDGa/H52F4FI5OI8+4yMULYm/WliZh+Qjl3CPUf5+5UkpeV11S07GarfW
RIRYjQunvFpnTJ5llFs5Bw2NOrEm4ff/AyRjUzPmiZuzgmnQdSdrYunLGYEhAEh19O+t8Mb5hBiS
i3tp8UT6W+uf3MeDUCSEPGVJtjjiU8rV6H8XDWlc1EerUe1w3F1CbcGzPBFy44w/pYhbnaWRNZfA
kQ5EugY+Dvd/0mlm4rdv/QvDP8FeVSFxiFWsr/BDc4GdlNML9az4swuIGxLyshpzKaV+NJl+4GlY
blsoBUxIfihslQCKFb+84FFQvKuIgp7ha/muVlNwRyoE2NT0x2DK/YlPRTjjF6ibrYiTzHtGuEKr
ZwABSI9IC241c4ev5FUFNI869r7aS/Ylll9Ny8S3nJd8yYnqswRQ44K0ZGB2NK27CaUI9Z0Pv4tE
pC/fFqVSxa7JoLc8gU0mxbI2Dw/TMiXFeIML58KVGxq2swbQ5oN4bfPNvet08GMOANbhbgMqmjJk
xxaupSiq5lwubC2m5JGV5DYNFh+Qljfksxaf6+ewXCcNMOpDQTT8El608n1nu4vwDbZs79Z7vlNI
8SvQZSvkWdnuqalqHa7+vaJZyC8AsuXcY7fpxbxcsWIniU1niqAn5Q0tjXIFZJb8/3fFsxBJn9hN
sxGct1NQwrTpoSoK3/nJUimyUm6U6IWoIoXw/eHsZeugMpmPubdzwITvu6PQFFknzm0BcDi3DzGC
tm5KcoRdtSinkUgPqxhIO6ZoBRXjwa+2fhKq//t70+s4Nc9VoAkPCBPd1h7OF4DAaBH4lHgNHN6T
ImQJ6m8D/NrK58IUEzcvZdcprkju5vxoyjMxWevXK6tELjrDOBCE41N9lJ7/L9439mG1EOi5x3GE
n8X0D6p2vrq+RhfhVtRqnX1xvWwGLdtqx+765atClZk89Wt423tGrwBgavB0kchGynrOcG/eo2EQ
jLYNrHbmbpdb7pkapsQYIzcfCun3xvWijPVh5VDMMFjifF3ypKJ7opEor93DYlZue1NHh33RYp13
2ITDopkQCXCqy+CJOwmm342ZRPvPYa1sscKqyzLPK6YhqNtvlUwcHvSW7LGlt24kckJKD0fW5fKq
7ni84uPQ82qqlu2lxx0U+p1ta2v/7iwJ2dPEqfrz7MtOBIsaUR7uEzM7cJ3HYhM4NDl92xquZJCj
Xno7gBw/cisTRjSxo9N/qjmviJ9TMCvct9JFO03wX80h2+vsB3n+z7bMBQJbaO7GcyV89AOSfxIn
dqdqawwWlnH/Zu/6VzUwque2jlUL6ReqA+J7FfezhX6FnA0Q5GVQbYNjs3EjkiVnU5nW9Gez/k/1
uqTkJYy5rd2Nr0k5eGQ/ok1Rr6e74ZprC1NDFHhEg8lQCniZvmpAYwW+K0moIWaj4Ox4ilOsm7Sa
ynxqb1EXnitT/u1XoAZ8EVKfE4CoQ96G5ytPCVoLhTJvmPHnWp1Eys9/SIb91ty9BeDGB8uPSj04
2G8V54N4sYEXYsiqJuzlhMxlxmlClfV8DW/mWVM9wDVsNExCGjFciSeWkS8aUSe5NkQZ+pf7KfQd
Po1wTrczz4L2ZgyiXz9iDFRLbn/Tqjo+RnHVW/0w+Rg0G5GbRxyWnpZPyk7kBvx3wvf4Mei6L7Sf
2OhrDVpNDJDisb15k8dm61TmGG0AWUqNcyl/1nMmx05HYXvVws3zB3pcEifa9hdv3Zv5AHchRjLt
6G2VK40cHHWRf6GCXamzQA8lcgXvp3E0vzrhJW0aomdIm52DHDPqttQ0jT2VFxvnU+wdhfA/VfnC
iCB0m8Lv7R7OW9c7bkGNFXL+cwSS9u1ZYRy13ZVlUSLeZXU1brDGZIHYiwlS/L9bBYclmGJ/fhSg
ZjA9FNV8G3cIViwI98ddnrW7+0rZ+Y9ToAH65eqaKIMNLMnOIjzvalFmGjBpGGSt/9oipXYPAOvT
8UI/9RfISN8NKZB40D18mTLABBhNhjKWXsxjoK3dwZS1rn+qyzAQCzRaKOQ9WqBT65xqJEp35wv8
ogsA2YOh1AHcaWlgsjwVP1OQ2FUIxrSojw7EV2krZ8opmU1Qu1KN1aAaf+7o8vG9DpF5ZxQQNKP6
vxkt3PgULxkeuANEewZWKiQqPzHB8JilnW0HK6Ighq5LeJaswqKj3+VXClwXYy5SzJt07otgEbYB
x3T/fSrFrmWW0Lmx5cqVYYCr+VVqqjR5oy9VjkRQ7lTl5iJJEgsaW4u0u0i66COjU0sPBH59BNba
rHa63MJmj9ud+yTvTTmsOpg7yg81APZeAm6OHjctZLWg6JC34Q2DsznZ01tBGGC22et6AkOD5QsT
g8dUcvulR9pqQPlhX+5zETvpUMP0XmfvOof8NwN/SQ6xU730ECIRLDVxX0Df0nkLKN6RX20N12b8
NHF91N4+teNe73U75Zk4Sl0dYjX8FEdUoPcBgHuFMdzRChUuA5slp7FE0QlJK/2klrfqL/CqnG5V
marA3BFh0HjlTbL3VBf+4VR4lhvYy9u4lhiKxcczgbjevTzDMXMbZsX2GJX/CocVV9/hncFRaK4j
R/Rty74537dIPhYzSFL4yHoh6dPLqR/v2JQf7/Qn2q1PLWa5FgHGGCkkPnUgKJLRfNqYzbfvZkYJ
D59vl1mnfE8j7DMSHlxkJtpKfWeNHs/ZmJ4HaqbmPE4FFJJs2ooZAkCTllF0VSRiGS1CY4OtGi3f
JiPfQP5ileOtoR1z8FWqEz1nv7Gf6akUKxZ/EmvWkEkVaDRLQR/pssSUxGbPCMnOiII2g93zQShd
fg+ynl+k0KsO37A9AICk5HFNn2IUz3UyOfJC/n+x15bUHEX/deqm4s/JQQ3QuduQIASaJ6ojtPuP
sAJn0svPDtrm4X/mdzIsl8hxMqEzPV/a5Ult0ruU5OoR0PfwZ4llYIbOHrGPzA6u9KcmAKBO6u/S
DvZRCd/dsJJEsbY67uvVQFmbanF782qhbRP8FaC5vwEe2G3iYir7+o0GrMNCaefxQ2ENmGARNlV9
5/MDQmbtOM07EHJqRsB8/C/WdgXaY1NXK2miE63zxysYEuBq7OJqyavR/puQu4FYP9S/KtlQoqbq
DydmXSoeM37ylg0eEJ+EZspYBWlgrGpXqZEybDChNaZUdyfsFYVCAF9/YKBs6oWtA37yUhV44u3T
a37VkB6VlpN2Xrw2l2/1ecM3PQIrEO0lpht55GfLirys8OVDB5xXtNJNxGRt8COSjFiKo/uRDhvz
BCKD9iHseztAonKkrM/LO9aI6fhM4R93Ll/VUoig2eUUpPw5OqZsMrq09AESiiqdH9BMIzNixl67
r39XaY9xwDchHWDsINVRXjVx/VQLK67Ivh8j+R+PYkT2QpsZi/NTc5xXM7IMHlagsVfdIguATWkK
y2q/9FGe0dwdDyfxJ52mFxr0MWM5yro5togpuUedJ9gzQfdxJwmsn5A+uFt/bfmORF9yMzcl01h1
5zNlagNXWOJxA4FhNpuEev4qkAUNxYlwYbuJGP+04H7RyZ/MphMgL1UwY8s6vSxH0U6KEPF625At
Ov29QFruuStW6WA/R+klvPbPB8wX2+8wfY8hRr4TYO/1McDZetk/zoSuaJiEaUZwL8ZpFcqrgG7C
t8ceF1+Mu3v9LBXya8EwBALQuo/V47vdzqAqoLQFLnaw4GwIlPK6QAlQJpXi+wyeIYw6etzdyXb3
3sMKodibQ+1jOtpZxyJLwzDIOY1DJ0MXCHrpf7P4GbDM91vaHAxKyon4oAfLca5Jw71CqAAnCn+M
f+6FyRJK9h651yQMROoL9ZAKdXLukjoQC2LQWAOB2jtF31xaEZapJFrRS8K8HYpPBIq8LlmvBlh6
+ZwhSA6QUH9vvLm9Ma7lZoLdWnepBNrsg4z+O9oZJSHyQVoV+biq5ymIW/y0/MD14rvKF6YCbzug
5wFBS5upbDStLz+NBCmqgaPR7g91sFR7Oo4Y4TriTOEsBkb7dpuWZZTT36YEEacUVxojH1MGglb6
fcQwKOzI/mqA1Rdumg7SlKl4ZUd705RMMX9feMzlr160htLUGDD3zNCkpuY54RP/MdCE0GfCgVtS
78fvzklrbEjDx6NIoW5WjOUMpzQ2P7GFeUInOVhY+mWEa6dBREvDLY04Gk7HrAEAT/Rk8Uen3TR4
mCaFwQ3b4tWpQBy0GO0goWoNfeixBPa8UlB7vaJx1Zdma4XlaapkciNZLLMpLhfsE5Tq6KJUqEwH
9HzUL32/pS31fg2zcx59UzlHFcUGvBB2665dZRHDD8KT/z0bnOR1Uly90hD5EIZcWhmWZbvFZkM8
ke7AlQYfoOqHKOx9kj52XBCujIdb35jZiQziwd0Hsllx7YnqrT6KEoK8K8VhLNBtVJBZVNtVA9Dy
imtUCpeQwW4tjuR7tZubiU6rbLh9LUMEFNTvL9bMBi6zKghgBH9KvAuLExvTZqILkuLqSgTfAcsF
NkyPWcQTZgPq+3PpUCJmYBo8Y6kWe5GdRe/ArJAn3KLyphb6xTk9PSOM3YiSX+nW+N7RhSZNZK4T
W7kxs08zs7ItfKN4IwEJ0tpgc808ko41MODv2WtmZ6Iqz+0f804r+/pwpfyBvzHNybBT9xClexf7
zS4LsXOGp4J4NweQio5WERvor1gd9QQ++IcZBpNSOnSll2uCo020JorY7V7pssN8iHsg8Vx/NEI3
LSogKqjsZ6OIV27kiOwMl7rdItf+/BzbGv+kn3lIxFdQG761NbxqaM8AttImwxVjwDKX8lChzAeX
8iSpQoBNSE431sv3CECtbMvwTOBD0Bs/qO/76Usi6ieDXI4ffi44MG92uL5dHryJlIYLvaa+WEFM
jX/4UUFMpwgZkDnyfTu5hWfU8Ntxi34d2PQ2S+4Tocxvcc8Rdy6xLs1Tzk1QbCdp9vQzLZZW9xbH
tXp9wCpylmaz6obT/ffnsSd2Hriolr9gCMsLzUnrK095ZBvAhAtDZQL6IXXjuIW+CBGas8jZ4Ct2
B7tpNZU7YIvQJicuSfix8NLNB/bXzTkktIN6BhvIE/rj3FELBpoCPzVI/VrQxiGdj1Q4gt0MyvEz
W8RjUXIelC6D949FxxmkJUQRoqxFEheNlO9nM/G+dRzfXGhQPTERnBHKKTM73wE+bdgZpVOC01uO
voZq92SodjXVxsMPfTTOx/CPTFEtDtpAaJ8QbsaaJUTUeXGOU5r2Lto2/N09AppdhBYJxwFo1aw7
ApCFohyuuA3VqZO9/xyJKfX0IDIpurkgay/HRE2qGeZKdMYP1g7Z9PHI+mtuL0H+N2OiR0x5rNXr
//QxllXR839RCBOERUmDd7thAnsz1TmYJllei2muvRkE4mTEgU0NeYzi0swyIpJ8nojsjsZxuC0D
up4sxCK6c5XJdNrZyhvexqsH73J1q0e2ptWux2kfxzp4LXyKLxsBe/PDhlU/sRyUhBDxSsPIyOr3
8kIDYUZwuPvpguHv8oY3vQ+b3DA5r9uoC7DsQmVZvd6M8jonU8UqBL2hzLnD6Ce9x3BApOP2djUb
30uBoa2XlWLgRB6g/HIklefB2JjVGSz8y5Iyh5l7M9iQ8RH4zrvtwDEqPScZz7/JeuPrYUMEBhKu
QzPl2+uPdfAeBxppxYDlFuyFrCauw63iUeD3uWcfsOFeqccrBkSVxHkUvdJNvphQSORwo1UHhxvJ
IS+BgJJQb0t93AzxTqh0wNJlYczzj5ruaE1EKmBqKPLTrXmJ3FLuJvYXMcy2BaRO4rTm8XlOmxro
pfzy7UYSAx9LScIecB9AbkITYT4yVkv4T0wOD+cPhLtBBjj3XOvF8e9Znaz7NU82xlWsLHrjOiBY
P2RLyXpXDCRKTXZQXs+luVa5P8XJS3mneC/SYR5zLkB9GE1BAJqYChf9wOqhw9bl7CJSsYZ/rnlv
0llUFCqQSqCZ5GCggfWCdU4vIEuN+5e57tnY2+T4I6zLklfqtSV8jOuVLYKtrNe3Xm0oq9VJuwdO
XBkXiX+Bf5SR3OM/1uBvKTIzD4b8QAtmLuCqiBuK3Y/LMqqxuwhDPa33uZTVJejvyFAlyGqiv0oD
b/rO6tm+g648UYiO2kD4vqkQtUrL0HDjXR15ZOcG5c81OigUaqvWJ7x6ZoFkzwqrdUB4EI403HS4
LEwiYyvQBx0xU9tWZaG2s8Hsfc+DoHvVqFswXJ63S3fPppZMsYYjWLWIYhCeo0K0cPTfIW3M7rMs
QXYPGfMRQoGAYjhmJJldNxWxdqnW7Bv/71QgIgdjqJe2K8NAXHzdBwlXkHaL/nUpSw7BbAu7jzBc
gh6JaFCMcShq2RS1f3LnwHImI0RRtnnhRwEkjEEG81HtH3syq2DCI3umWPNvgeicmHLIxzxeYVWR
oXNL4URfvUHbaUz3T3flAsnmBiKUUyTtrwCuI/kg1757jrOjzGDigBkka1A0KnS4uspEWVnwx5Yo
iy/B/iMDM/4qUvKADD/YtlyKH9dOhYNGgYEjHA67cCUNVT5E+vTXQAL3Ups9U60DtAK05rmAOUeO
zWcOeHkjGKxUPTYx+n/ywGfOTpuiE71g30Abdx0Ba+DNQ0xdyz6xikxF757mfMnODWUiF19l7fwq
wj1fKtdYT/MZejuo1uYuUmbPxt3P2dmlL0UdjzFRA0E7O3Ncp7fKd5Gzysu5TNMVF0MeRQVGLqPr
6Ci+IFu40bpMw2Mxks9EWJ0NpdteaYJRwwFZZcz6HzMSatcr+6dtGnpM3L7BsCUdHObFygsYHP8G
oZJ+QNMsWlDOkcoC9v9Ltlb6m/aO9q6UurIE0B+OGTwbbb1twLG+cntbdCbl6cPOpSca/R8rdycg
1euGNMvkl6f/HN7tAuQ3LR87Icm2hF53FCISXYj2OKlfZGfHcsRU7A6bG+5d8bJ9dftlyj/U8byV
I1JBbWGwefz/lk4PTlLJk8rngzUIOSAu6nGE7wySNdK/gO1HxnooTC5Wg2SGwJLYZpcJU74D4M1h
cVT+u5P2Xt4/VEfzIzGrNjrs0KLbpdauyo0ZU05Tdk5gvbMPU2+wEcQf0xH9eVo+CITQjCxJ9sTn
W940sCXfNvoy6pcITvhGdp/F1d5+GEyi9hotZnsBaSnyFTwwfYLyq/ut9hIA1iErkFDjjZkMNoXd
27312D1iTDLbY1r77kAtAUigENjj8mDDYFedxv0RhflOFGbzABGOeoQZGgowoK/e63dKoPbxx6DK
+3ujzkDhMGIxO1w+Y3/oi8BXEbjiILSucTW7Dc2lStZsj2WhL+k9jnDesFbZ19DYcwrCHoY3JY3+
uIbGscchmvm0DkcwlXwddIVwGc6Es+hxD8U6zRDebSYWgxjTyEo4+uwqnAkwm0Hfetb4eK2gdcSA
9k+yf6Qc5ysKUwK7g7tCqe+uKI2jaLjvh3I/4wYmdEHkgg0WZn0660jcY63txJMy9FIDAsSb06OF
hRZNoIM0NaekpALP9RBQlgaNgIYB6JMdbhlOn4z9k957IadB5mfrnDnwwDFr32mY7Z/QVpxPVur1
NvuEl6VhRtjZgu485Hj1CU5ty+sRM7xqJABt3mEyK0xwvflbZ/8W7h9GPh2fvXJe6kWXeL0u5xku
EMMmpOSbRqDjNa3SFkaoqgxJ2Y4vEAKtRtI2VDerQ80KwPQsQ/Bzv1mdRcmdxGVK96j6FWNQFg2k
S9nEZ5URgkzEit1IHZ/+jfKP1vk5L07pDd0Iu8riwD1ZXvwsXFjdVezpKLD5lNGmAWAeLXC1IUnL
Y5sY6CCAj3+XijweMkFWs79HeTQpmQk3CgN6WSZKWgp6MFfWlmWkKQb/GW/UUY3xx5VTMlYGENab
4Y/Cs3q72xcJX9sY0MUqs1L6yzKVXuoXxVNKqKCbbRZMSoWkYJd0tWXkoj9iSfMzDNQHlv4T9tYd
swN9IQmenT7wIvQMHZTs2mGYFLCjVvTjH3k+TYdxHnHca+ska0BPd+QQJXUBqubdi88QRFliY0Dc
LQ9dDIxzRV+x0PlM+MGUFU6ayEAUhutcOioELypbYyfw0xZMXdKO6YQtOK5ixCsLHMOif2HI9inS
AbZ4GqkKMnX/2qESFub8lWiSwJToayzXqm2hfj1IZjV0pgzNmOnIVQN+sFEapF3iWNU4ZIQALqUe
HSaEJ2cY2E7Ky2KkM8WOltRx+yCgYUgFp7IPukR3ASEzrgDTahEvvFjLLBYeHUGagt9oM8h8fprQ
DE4kX/jbAyrJYTApNxgOhK9vSOfRN6SFYHXX1+p8OWjogk1u0BOgy2LZuJ82jSbXBShgVT2Nr/wD
VqBgv4y5cNX/sSigvuSEkmBToRDpZAr5DHhjtXNcGsC/4iM9IgT0eTOGKCilhNcWoxxJYRI0D0A+
IqUHlIbyjdnbjGTsfBDdXSC42Yf407OV89mQ8SgHNWFCeXdA/Q3hXpVCjAz1zydBqJg2TYOlli8U
97tsFN6tpZ4GY52b5j4frgYKfkydrDqUv5PH8KAHmMA1jkhETEPnfY6b8iXyS88Yw1Usp7ECE/vf
ANZY1hxfkTIhw2U+74EIfXqdwVEcEP6JXRqR24LpeoyJeSvNZr9YGE1FyrQEDkuVSONtj4j1WJZu
2XKgePGKbQjWkh0yZjt6vTTnMmH7QW0oZpFtL1XTnksjUiL92SNY2Y73VaoM8ocIkUn4KLRW7Yfm
uvLyk2NzIuMjljm4EacC/hl2znBe5+oH1PRMPSIPQmzwewO+VfZUgPN5KTJxRgWh4G5shBJsWy8q
oTVncainVhN5OtNNP0aiVjr+NwlxRBhzet7akyaPCMp7tDLnqLPVbZ3OBDyVJlhAZ/Dm60F1KGUu
7u6Rz05OPPeevfPGxQ4SyZvPKR0jAeW2dcskHXvg5Qg5JZbiObFdHUXIqMtQsqfqrQoFiYm2wC8t
oDxeOboBVA8q2qLUFJmad0hbd8gziAKuTKcK+C3ox426J+pd4TOQoYWxKaQIbTlZQPKSrcCorgAg
wAR9xY/TjXlLm6/gSOH7QgGZ3cRh6QefkUz/6mMYz2iLsOIMI3Lunlko4pPp5eVZOkyNXBHJFPUM
OfGn/tRo7FUxx/U0AzRikswqLQ3m0xvNG+c10Pwuk0w1TJNA0seqYlbystTRtmRckPzVUlfUT+1t
yAxHgmHmvUu7wGf5oNGVK9HzvYzN6DbthMjc6V/ZZhpGZXGPf1PxXkBTAikFIJI1iZon9hKLASNQ
zXCDrFJSPeZx84r3WroVePrqv4qeUCtmZy1qwQXyJmfleqSZfL6HUpweV9iI4nxt2i22Y9+fiLtj
eg7hC7s4JS/n/UfcYDZqPtKFVFxcTIUeLehObuTBT22TLU46zvXay6hgkxUXCHP2pFAOWNSW5bpz
bkymcyFSyKfudSPSxHn4Jr/l4rBJzIisZ9v6uqgCh33Ob3Wqhpp7hpgjClClPicm6pnaonsUc/KB
7GlgG2fkaY4f3C9zkB7RmXrxWi4r1ke+RVbfDcsT+mvmKXtxO9rFlQyvzYFBkvkDuUYDos7OD4zX
9FFmlyfuFZr8x5kZehqUu5YcvlwdNm581SFAlDLMiSZBsHRJBC+A1knQcnuNiRdMLtYriT6SmsBv
sF/0QDuh/CpZux4Kv0yTiNGKCt7b+yDnaqPbh1fwjsaLc9tilccrySi89I3/FUxyJjiREJ1C8ZE/
9evIcwNxTKvRA3sH+WfOc7/4iFlQAg76VgxrlXU2ibnI80yIanupIsx6Hz3XbtCfFRLncPcmjJgJ
D9f4HxYpnC0FED8ujQGlu33o/ojKQziGViZIgv87zifexx7vikXP5bOQI98TKRNe4SduBrDtuSfd
hOjU5AIajG/ywkPsj0zaOO5tfuBfUI7WNgxwNEKg2FNDUFqhURjMBD1cw4RZAw1x4xsKsrEFNjkP
sMEmt2unpM7cRcNxAmkt+qS6T7+0TctWTzZj+RGUa7e6wIyT/Vz2pW79YjH3cOyKtC1ZvNFEOH70
ZV2kvAyGNo/QZWwxsRPMHCImXtuKxL4UN+m7CseiJyhz8s/buZAc6PvstvArfo/ip8P5z55OuwhS
xTqZdGAYzXcKEOWHXHvh4WnNIlNZxhggWgeZsyUb1Hs8NFE/fJc4IEQP+6SzDf4+jdlj+7d8ExT8
R9UA6AFBA84AXyzNFs5L00iOfk+GELXNs6UyZciGWoazs142X0qHbS6tcrDe6aOmCrhARzY1y5nF
MFmUFlE6vt3nMZcUFnPDuJ/3tdSfHpQerVBpcZHdDxooiy0ydJgrhSNLSzNnosXKpNdoHz59kZcI
fmPFYXQutUr17O7VYLzSxqZrQJjxSUJO0FBcJA2JKFdSnxcDbCjtbZJgm9dmIV06gKtNivWYj2kF
pTHtZhtA68+exa8BoG3PCMm0k2K7k9x2jb8EzSxnIYi53vvp4XT6TrPKBzCvU61FyQYx1lVJuZ2h
WlEmxDTeLr3uxuDXNKWWlJIuTRKOeUeJ9FOaleUWpibO8Aw2YBKmA/1/V4wJb/ar7SrUQkECEiQr
VZ5qbD5ph12jWu/1EYY1z9CjiAZwrxd9bPmA7HDFMSP4wvcbgOhoOHGYGXB071Tb3MGZVvkhATR0
mfXH+8H9r1Oy9pSZHaonWRJSzMzmeRsVKLhAKwta43uf0HLsXhoRfSNiVKt+rGVpuQjuvGKVoksM
z1XyioKjCR4lDwDtzM7AIFysp7kqhtlzBCHaAkD+S6J/vChtX6nFYn4d09BJ/6xIMzETkTGJbRS0
4yb+8t9ussQp5pVT7zLAlqkFdaabAjhf8bvWblmiL0CgsHrrm71zMNmx42d2B/yYkXfdmWstTrTJ
tjmDfIp91+WIKkRmsgcw5RUG+G8IhAOVhg6teLVmhihPXjtWsR7SyUpiPHkPuvJCcWIBcjsiP8Qa
fDU7nL2WzG8/C1ih6VhdK5R0lsYT2TNMrLN2KrUVGCFq+IDtZM1npae1ASkoo/n5gUD4cBc8oyxR
4luXkLBQAUcC4yIs0DUrsHZWVv8wKOF/OjWOuWR3meMF4cuAUmbQ+jypYfJAxTGsUI/X/zKhbhK7
6QreM/hEqnkqUQAMc44RJ9KHE75Gz/thsb2jThJgnncVKyx65bBz0dv9ktkOZ1k/dzNaN+96BYP5
cjM9VeA10fJp4v26Slf9I/N97WzjYSB1l8U+GQ7ndbAMDUDcHugt5j4UwyyPJ8tn05lhhYhp0Ng3
7lIm0d8ex+molnQBLB2/ZUX1ltPkk9pG0KYGExD1MuV97Tml20xGugHkhvFV/d7PTpDx92folL/R
mJAuD8nk1ZKuvPoJeGc8Lsgx7P9ZrpOirvsEpMR/UdpwkaIt7+JcDbOabWxe31a0M44J30zpLycM
AFxeJbKV2x4ZChZrOAq+m0Bl7n7Lh1I3BW3k9DMlUivlxEz7lnWWL0XCMiJGwTOI6e8MYvmhzQTd
pOyD+w+UKoIExKKkFO6yfDQtCQbHMzefcKeb/hz0Qc4tFPzONuZvK6gsja/o3VnxWOmXLeFhvLt6
MgPik3QU+QyLhb95L13IpdKVnkkAWAzQn/B2bX0gM67PcMfhCJH6+aYD9OJQ/06fzlzrjVIgDFQ4
tLoaN0LfdOx4ykWjdYKwNWIl8M7uoJST7c97/JB8wJMzzggXJNG5bDdvutOLka9APCyjJwW5Llx5
b+w2ZhDVjUDe6vHvQBejBcToVQQGx5vS4vFt7fgRMcWoSz4A3GLqb52QqWeVwtNn/fUz2M6E2Kn0
EvYpadj7imzvAxNRm/ALI6RM450ZOFadGUOu8JnZuIiAo7cwCW0npS+ZK6BH+ni7TxmogLswcfYu
NCar+Rbp4HXRt0ZOqgNos8HQe1og3+7pvX78ei3Rv8eqptyQJkEKMRgbTqMg2xePgnetndC7gfgv
HAqEMh38gdd8DhXIJYaAYWxnhMvz2Nmj6aMuiEnuXiSf2rzfmzOrAYrUOIJENYyp9lC5suWFDF7J
/CGluX/WoQ6autRfZ4X7ywhlH3hPCrjgBKurF/YnfO+kfhRaLyV0oRspBNd/0R7XJXDPUVOSl5dW
0wFAEdBvVVe0CrO7e9NlnCexHfP5KOXBoGQhkTTcZbshsMbKSXU2nl0jI8Tu/8XJR+tPb1Gc3F1f
G1szfIBlwRyhvNSHPeqWTb1Rfl5T8UktM98cMB1ejhhgMYVXOVoN45isSUonQ+bhGZ5ygzVZDmGd
bA8UICSLG1cuhBhnKCPXXCoBJN72pmpTjqsaAPJXSZ3sOr3zFZxHHk0XDdWkE3RpL6tKMLc+hDf8
TC0GlMPVGfB0jKv/Z33admvM9PDQ/PFozWZgXkwfzq4n9Ab9HFKzRZlw3A1b8A+vQqh2BzOpeOcQ
BhXmZ49/QotdsDyqBqn55Xoi07uA5TOC4K4pzPF520zToLOYwMcNc8FZMTSZE4SWF8kqEOca2Q/W
RSuYnOWI4OsifB2DKgZoFhsf36ej0+gFCL/TIf6+iMcnwbB3Xx6w8Wk5nDEajT9kfWT5UDc43NqH
+GH5dJFurDfvnmPwekNIweHUWMCxTWvWKRHeucbVDKHmFHhvSQBfqxgxJi7G+QyDdSEJY2bw/kWT
NutrUHE73T4C30af/ZEvIZ4mDC/t9H2N/OjPJbmEyRw/95Yu2+D9JS2MiXbsidZyyVZDW/HqcO33
AR2vfzIXWeOWlt4P+SnF2Mmn7gQ4FH8dSYb5RPuAdBLtkvpVw4rWqsA/gYNMhnsbz1N/ecFrQmqt
ZCJVqB0J9O5oLgBSLryXkp0V9GSFcT+0UmzP9/qLsbidM6dwfCZmbCxV7oAyIMIMSX4u2MWt3iSa
nkltICYSRP3MqzYpQFPiYckusCvK+jETPfKVWShKYjg+nxTykWxO6UsruXY7D4ifZWIQGQkM3JGk
f6JHwgJqmd11pAQpkGF8ep99EB5CZ4oAEIBDuOYePCUC08MBsUxEFampnhC1x1DOMfoZIN3yQmGP
yDF3sLe1bDSOSqGFdiNcJx10RY3MMRXzugNNDZhI9YXVTibEblLwE2FMEiJb/By+faC7iesaav/y
VMmiOjvH1pQ1EjmsUxM03JeSwityaDmZ1+4wqVZYkaStAdpDDW2tUrGCJ1EQlRaEY/N7u04yzVnG
sUPdoWchDoAYhFDgSXQtY0HTweUueANjZQf+DHonkgLK5yK8mxgSu0nLAkrPAa8rjp+i/KLRs7LX
ThBsawh4StkzH1s2hagD854YOm5byPyHeRi7LERXU+jSAPjBGFsO5LLV/OaMIFmPydcMgt4XmGeH
d9N1puIO9X7s+OCVAMwKvZpEcCodPsdSkbsbZsbDiFohtazpqp2oCLBPIgSMa1oGG3eBhwCBOmMC
+2l+dUsdlM3EcHaujnXzSvk51JxPE4r9hnWskGj3L1a+3jVI9uK83Wf1Sqv7SvA06Cwex1BzNoBX
VrcMuIZdyP1QFbOoZUWook1OgkLo6VyGFyVM9BHMGgueucT8p69p81wYAL46hu6/VA8QYCMo6CLY
bU5cz4DxV53L8+LLNruZApb5+xnOw8nbJ2BBFPBKvcHj4LMsu74izJUUzAKFbA+R39wCsd01y07a
MsfKp7Rd8O/pLHt1fap7eowNvT415c0HW0WNWG6gW69+1H9XQxRx3LRYtFWhAx9CBHsqL23lMnOu
0IXTejT4wyD3vaHi6It9krJZEjXNKJYVEWUvZCb76qh2LED6ycrZDbEv0LRHkSRBwaJ/MrP2mEDL
9bVmwFjWhJnn2qPsxLGLchTnWOjmlK0Rt2Ephwn+tj/k9eQ6o9VoE3qoSY31je8Yi60zlCt97U86
8GcmlxnOk/gxSKBZnmwVbZ4BiHhtXZpt3pndFLQ2HHtRlzPY1Zk/zP800E6WFM1/MtABN05m7aiv
jIiEgs5UZZ7rcJk0ymVh3wRbqVkSaKKIRhfxixFBQqH2GlaZ4Ir9aUex6QAtjDqgZY9peDfvffVn
/Zq8Dhkrhw8gX8R6FlAtElpoluIRMcRPXN44rV5f3l9FZ+JMs37naUo7bRGdJyNlVaR0qC8zgLIy
FOtcaxpRUCNTHytIHHeD4peqI3g6WVlvncg22kXetSb5mZuzJRSKi9k6sfcsLMFPbUb2OXiJEo0V
rdGclktTehsptxAcixK3PeDuMQGeNfaRRGEOKrGaazu3U8qHF8VZL8A9fBopHKsOLrzOx8wOifdV
su3hfTSDGVuNMOZ8JIi4rY6Tq6aAuTS54qJkCzf5XiU7GLUfnuh4dqJxWyn5VH1thiTaN6Y1y10r
ZEmQsjh28bMz9uaXAHgdeEZO/oCl+6z/N5mjCFV9GSBzdARBTWMUVg1NTl/RHEKtFQyRQeITXPaN
lI6jofFVieBC3Q7IPUY+D/nStxWMWnoMQbz6h666+fPv1eHGwrSYGzmTMoT1C6xradxpLWKF84Mi
KytzK0eOYBQm5lg1rcm7S/COWVCTERGtmuX2vncC1s1c/gJuA6rFrrAhPvMiAwnbvegQ+5pXhTUp
f2Rx/8gv7SMp4lW1YPcJnjCgWEsjXD8el4AT6qIDebQTJpfl8cou5E2dL7GMEx55cHakuvAqpVz5
cs1EeO6QuEtkksOciTUdzshJ9AqPlUUmc0WZHFWvjP8ZpkYgHJ1kqjVgRhmrmC+6Iz6HAWcMymvk
WTt2fAdycS2zvqSpijj3VAz8yYGHx0ZxDM/eWcJI3bfhwDurbYQ2w4ahAxvUjeWi3D7h9z71OI3R
crM/X1gEUb582nxTeJudHa6tJtkjgID/6NfaGBEEcp7b/ZZnpN1/DnZC2nJLl0p0M1ZFFG7tu37P
0686Oxx0J+JKNioRniuAR/TEOn3ZtRz0WeeGEhi5EnZaZLbfm/1n34DJbr40JrhFJeAALfM53CPN
QuY14UFHLBJySFkHHPFkbLcWMJBbrFtxqzjYAMup3xd6FTSCGZ9UJt+pkeZLfP7F0OEKRT0hBESI
eezqcK8IKKVY3n5JRQOFz4V07YqAFFHfk19gVkPcJhQImQ2KQeocp/6NoXxgFk7SnukyDRcTqygw
m2w8uzjWyLqD+i2+n3ABrLMK5idCXyO00juZEQO4TVCmc/NPbHIC+3oUhKSdQsqtWml8xTqx0ZTs
10l39TFwwZNVYB4xrR82JM2RpvvJZb7GLRaspBboDrMJdwhafOV5kCvQ/EVBQgn763ce9H1A/5fn
RJnSfAPGck0csR1nRLlN8rXJ+MSNhgw8UHZm2UH13M988YhPnKPv6U8Ary+le/w6aj0JID3+l+G7
gks+GhzoE8YrvZuTMuj6PqtyHYfmLkbbAsMC65Db5Ul18xa2X5DMD2VqjWUO4nv4qbpAmx/FT1rM
jxmR3ipUDP/0hSeJj78FPUq4CdFaKXecQVELyUfSK6bUdqGpJtlASOPbrMuK8XRHBN2QVUg+bOvK
5Sq5gFqPePN4d9qJ9YlRwrJyxtqMB5fzDrgQMLFiKLx6iDx0Ri1k32pQqjH42pmkgXaRUuQKBTDx
nvfbIUJ7ixKQKhrWnr+x7cSsQ8w2btbjoB4Q5gPkFRwNFhdrx9xIXMKzJkRlrDoyqizIKMfqjblE
ubp8rl4uoh14hk6M4BmoxFVYfKWlWjP9VPIZJa8T4H5mSG36mpW+B783vZ40BkRAJWWUxEFLzD7Q
P/4PvnrGyxolJaMtRW8qz0gtzoi4Z+fFPIi66MkOiaPAqd2eIeBGSB3Ao36OLv5oXb0bZnQeyo65
DPdn7KigGQy0Csb2+2Fi2D41CnEHT3h0n8gYgnoK15MuKasbD4eYczy/WrSduYsoo1JFcOEdkPzK
TlShd4Fg9j977VcCTWVwMQQEaJiNa74IlZ1KeAZbVRRovc0+13T11/Chh/5+kNfoiI/Q52khr47W
5K4zS+Hlt2vzLK339KnoNoUCvaK4+zZwIyCC9CzQg7TnWX8xoFNgQfe5ANDEN9ee+X2b7TZO58rd
vhBLYE4a9S3jOYsSU9Y1IxdeBBs/Rm7L/dundc36gYZ2DKa0FDDbjBW53QXY4hwyWzAjBvRCdRLX
AbLFI6XeNkxNAwCZGZd8akHnoK2VtEIK48zej6yeCIBeXatwSLkTSAt9Ck/SsZSlf3EakjYQnzrZ
KUp8vl94m3fUloeZATKargxlyKMDhZyG2i9a+GACXkGf7XIpi7dJ6Ae/6PO/boKT9D9tz6y6Hl3E
60xC4LtvgpD8dHSdu7MBHv8OPFnuYS0aBfY9otf9oyZBXyGkuhbseEBQHIoITwHpx0QmpMtobGOC
8UjnG2PzAdh5CL2wtvfAd5+UJVK3SZ+f8NAC19jJqft08NyO/G7pa1hOB2iw3DGDs3QTS3YqtQLO
9PfZWK6jXCTKUBhO28aNtYDDJHLq5DA4q+KQ/myK5WOs59o8Hfxhz8jPSGdaeqMq7/3ResWXhlbr
pbnJIytsQ0XR9i+eUthDGLm1uvmLnHDY1tOwW1aqNBDxcVc0GFWWt4lRUIp1ZLI9jz4HrOHfj02H
3os+TiW2Mo3WUKF6AFcDtDSDPHLm6Fi3GWFh0ZqJDHh811EYx3zBwFW+hfNxW8Ubi66+SAuR1rkd
EHCgk9BZuB5FeooiICLhbvXBflGDr8z1PTZMYtfryVLw59u2SlF/b7GdWFAQQ8DgzU1w/ysRjFyZ
OB4wKMFjOm2nbBOQ07bbsxlJXmWAGFsVgT2vkAyWdvG8lai649RQ9wHWl+tpHiaVo0v9Id1sn2iI
5V0mYJ5OVTbBLVN86/G0+z32u91EZwo4Jc44but0V4SffQR7/zNMrCcc7w+/KIgoJsHOY+wo1r+2
k7bRrV/QLDM+FgwX8dt02wMND/tuGipRddd+Jk5BONFlsAd6NtyPuRLCmYChBZQd72Xfig5EIfeb
FDouEpCCApvNTO1pRrQ/biRBgzgSwvPuUD8/DV5YlvmKXd3D47/cF5dQensuWdmHnjxnqIUjXuvP
EThnle0te3Mfnav+L9JYanGEvJ/eqVBLnmQU6yWB/GthwebQ3YcVizQBiM0tq/UusipcVXWtp+Fk
0mbq0H1PaOxkIVWtoue46jsXs0XiRRKKiADFGLM9em28hcmrCC90VJ6tYHUBqegY5i3K/iT4plAF
qIQizkj/8sV4IzpZlO2/gCECKStOCImXCYSqEZVpNUN6vfdBOFYiA/Yq8+Zgtf/BCC3MQmascATh
WJtX9bMn1ZAqqbvrs+pYGgxaytv1CHG8QFZyBTtKxdxmXAxcKv06qQASpfCPa6eJM0QJJ+tbnZTS
EnsdVmYhobY12hQ0bCmoAtQ+D44LiM02K96SCf3QMUx6u6jZBje+/u8EvHWyne9lG25Jv0NsxQWg
di5V+Uz4Gwj5paFEu+L37WEnNGvtxbZJDktUK6LPprzRC1vUWUWs09iMvzMRQoTJwtMDRtLrghsH
7BgfhwPdQezdW1jZmurlo5JeetM4iVowDMZdhyJ/C4RrhiKMmZULATB4+P1s3Jaz8gzWCFghFdBw
MKmBScmiUHGPS3T88UC2JZYCa9ZQtU/yat5pXbbXsyEuvJYd4vVPGCZ4vErnnPkSYqTGfO1ACpsG
F6Ur6ZkNhzo9RyTGmIZ/uqZJnsteLt+1De3Zk2UTSN1IaWI2xUrdqL3rqBGV8xxfVeR20DnPzrYt
uZ76IQO8rj8GemN8X8i7BfgIgQMdrU19BBfbBzyybJDbLM1dLfjmVEQO2lEmB5igg99pCll1ULwC
mSe+CEP89UokTBib/zItC6dVVuaSaBLiZtWpHs44kb+rFUJcBjfS2FpTuhie/Hgw4dG+6IbLbfBb
qAlhkmNmB/eA2ePjuju6c5SlH3mnvmgC5rO2HBx4VKYsgrY+o8Zq8gCCGbIZNn+TZUT4lKj4O3nW
rLCTg3pe8EfcfNXQo6Te/nwLNcYHEk4R+E0HeUotcHJHNFtRLlQ8jSZ2JsQdzNI7YgV5VqWqG61i
gBAVqK9DiNHHxD/mrYBcTTBXnKQXcOxWdSbkklAKDwkRVOpWfFR9vh8Xiyj1WE0vi5DbNzGWDoOH
HKvBO4ss3TiXGycwv+yPZJPi5hd9DBdKJPSDjPvYAZyHZWb7N+KCUEtXTigacTf7fzMlbncZq3yv
uQqEM8qvrPtxxV6c5qDREdsPP1hPptFOeFXhK9+LeyEnFG8aSUJrSOweQsD3ccbWpGgltKlBuQnt
zamv9cy4MxGyfA+nIHWs4R/9BPgCn/V4s+J6y/vzu/UPN1cjhVYBS1HIa1ZH0QMxOOoUl+OSINnL
Dn7WCSjeBxlSrenBr8Tfj7Pk4hGQuKlhHS9t76c8Eb7n97Kr6XpJkju+Y7RSWhpTutXWjc0KL98I
bRhC3iT/jmnXrzRZE4jUwauppZI88RlS21FGOd0hbtVCEgvS3etMMrITP2QLBJ5t7FhJvMy3GCQq
v9OAJt5As+X/321O8TABJOxJHT75KJlIi8KSoksR9atuDwAo7ukMIjv4jzlIdxdKbXSsSP2aHE9E
aCuzpwkNEY6Yu6VxARVoJmcBZbIIDWiJXdSIXEreDdHeQmxnchgqpyqX77RwqJN78UwutS1UFI7A
vEy/WiL0LCDpqSTdpmMv9Uep9V8CKl7U48zUz75+ztrojOpeOmIAbxU9E9noy8pM796B5CRGKrJD
kUBznL+wf82qb/ssEHFPU3AbL2/cwfEcwpYixKK9rXDpJ3PsbR1XUoxuuuuyycoODTZ8u5LWgSDp
ZIGvGmm9krpeUYW0N+7AhGFTQEo4llKD9M0x5gAQzNShlxXyGqLUejbbZn7hh2YpBdCwU26XxSsT
zytccvQfA6L+iTGwDZaBAIEUgo81gBieSjurDZXYPCM4GQ5gtVOV1+yytR85qyTJcUCIbqRow24G
VB6Lpktk5w6efuvcvWXYpwChW9bpJO8C+bHAoX7A3g/QmtXUlL6087vbiz9mp6jauZ67EnZ23iRS
ZUMLsSfLzn3X+jNZ8o0Wjogx/FjDT4EPleeDU0Ut+SYtMcVeYPJ55wxl+zrrLVouPNJ4zJ8+no0U
7hre7aV9rBxL7P64QhGEIazCFRJhNxsnkOUVQturtpHSMefaZVDHmwKMFJW0asXfbVH2Nxw4smue
Aq84JLWVkpu1NkepoOYLjfDM+IVrdmMdGxsfokPOZdCiqAs/ceH1jokz6bwce3JTuopvlVUBgLYZ
ZnZWZ2sMK0+WZz53hMAF56GgRtqqlwK4xZVu9+VDQ7mVIAVAADWnxIRW8i90VUdI8w+6/mWnpTOh
NvjHOr7o+CNVGDQaq49DSW2QLZ59Uje2PabxmuZBcUaobROTE/WZUw62n2LnfGzDUm6Y356shj17
PDLlUZvO4WBRkUHEuTef8pLFXKHJMWi7EF8IAIZF6l69mCZQ1ForHnSO8iyV7f8HUNLgIb4VQI8K
1wHaSLbMg9YA88qfoFUOREgJy1pgE/YVqehbwipbNjcc/dy5B4OdV1aFOY8OWd+zMqE9+hF/jGfn
34y1e9YdBocBSQAc/XXTr72vjcYzXpBxR71cTOU9Hv3ZDzqNYpfw1PvUcCJrb0jrUqSC4FKITdlX
8mMfYmNo1tjKZDThS2SB31zzCok8P6hCz9dE2aBllcl/TN0ed6onXaE2MMnwY9DdZqCz9LhcWHaw
/kwQXAf31GciPSYML8YTh2gzIsEZtI1aic5Bcv70wWyG5T5FcuezkjdXvI6Mk5GmsdBHL4KdfIXs
7dMDS+JlFZD9bEWEdncb6UPtZxjB1cqgUEcLzFCMqHtbg74H8FpvmuBLExKcxIQBrmY9Th1jCKUE
4zNDEspLKKtetklBSqX8Qw8KOZh8zwK9aGWjEtReD8qbjl9mKvPVkBArGI4aJuRto0w3zHISBSfT
oFcPFIlK7icG79vt/i6lgJ87tulBWR9urtR4+FM+zA2OQe+IehGpii7N7Or5Xcnbu96qWQgXqiU6
tX/FThnveAD5P07gVD7dofqIPFH6Q+0Y0GOtoYg/p2KX02i2/7oMvutfUkuPGVeo0R+cYnzt7avN
FDa2gpx8wrWjJCsSZZ9uxiz3txC9jNGbagmzQI1zAicRryMNI8Gf3iWQCPwHiIdrQwO4PZltGgvm
vX0c7yfuyUbVjh+ncNBISa7ICkldkH6X1YaH6bNvSZvPNbUyczuI/EKFMSuwAGXyCM8u5TQcrIIO
DADjIJyo4VS7+kBsV82flSMI4tDcWk7jjaCvCbeZocP/kf1VJiKJG0yd6MtfFn0OXPZlQxnPycmn
gxcG+X2AbKxUxdCDYYMvIfIn0PoSE0drG5GK2lEhiWoUk0ahlaWY9abMz89hRJypxsycqBEWCKWJ
tJJ7iUX0kAQC1PvOhTGx9IS9r04RrNf0jW4984P46Jfh39rjXT2iP1TfbBNeRvXZpPrCxpa//VU6
9QBB+Eu+YB4LX8iH+ORLGlclFqzFpWTv6Foc2CqkTIM4el4ug4198QQMwvAKIYhRUX5xif03EPZk
Vtm3JaUhM3KwxI7/BmfVegpctiycihXeUOGzt69ABLO0mLheX93l9CSMlNGiL+R+yvPxQTOofBQ8
GSIWFi695XCEZ6vbVM1r1oGZaOjWnEhH0BmY5RYWWTD4g+ye0jaUuMMLg1QC2MYy06UWjMxgZwS1
+T0PSOebg1u1g0Qb5gDpw8tfqKLzZgYWYf9zIb7qrTsXKkRDhxYCHMeVIXFuj83VEPWpzBQ9iSpn
ZspPJAu0/DRzFCwQTJev6c5jL7NepfAE5gbs6dHtCfT8cNFoIl97+Aha+R6k/fH3d8kICfdT5zn5
fUYR3i9WQt7VMj6kyl8brb7iUG/ghcX5oYXr9G0xuVgeXPx+0Ol07b4jcf+zcnaMaPWeZIg8EBXy
mVzhD16ZkFoyrJlenL86X3fb9PGVnIyuCKXwHreIgjW3ght/c6PansFzaQh2A2JBpAUasHS3dLYX
9WbKkVPO0AflYYuh49GpWn0oi5wBvRRCoJAGMR5GVuvdikWs/7X728Cwm0IYyO1z1F2w9/iUgM0K
e5OoDbNpUMh9QLCkUmz51tX/86eI0U9GzQtXBXTWLsch6J5RNyfCOCXco3Dd4RtvV13YpGiV5E3t
gPGOzaRHnrh8ZlnZxPdpewItr9M7Wk38UD6IAr1ykJYGOcrG61Uv3YJ+9/JH5YDnkU/UvrawHBmG
TMdi+3J4iGWoTTM8xTB6f3Cn+uxe6xUA0hrUeBLGw8I2rXQ/iglgD1bNPYuJ3EMcoytTfMHROyOP
xnoRQirmKIBeCONiN/er0v6tIgVAdWMQCfyh9xbQ+8yzdIJtZp5ZQAOdh/yKci6LpEF3yNAHxybF
o4RLeUMas4/Kzm3LiCJPxHxJdY+LNdoreH3GnubI9/KibRsbzFqh7CZRDHaTdyLBtHQQFZeWVTVj
+gpAmkww5hPcg8qIeYhtt1hVQRq7fTmqNvxNgd2GFCin5z0cxdpOwF6enMOcfiOxVnAZbgltqJlo
rpt/lu8lqjPXfABdmDudZvCZzcKm6X6fr9W5uBxYDWGYLxvcmi6eP6eUCWbXJNaEsrlh6BwlFMVe
nEKDWF6/2lIG5ReaHWqv76DflvJPLmpU4R/ffrylN/EicGnbuWNVkwUlU3HWnyq4gQ2+iUrTEega
YYWDI8Unw4p+uqKgK1P+WSw30BXX2kqZqN3fNNRMjmk89KMV7ZNFEb82HsVIzMq9+/l2xCgdyncj
T1n2jh2jw697yV8vXFK1H3oTG1eb+nUKfciWjDc80LcoGQH73aXwhaEMPsohlLXB/qSFYRLgVo7I
nGwwtxkDvMPWEjFdOnO6wIIZWm7nff6gYbVFf3FIxcleNeFwFA9lMvtqChrDOFD2Patdx1tq7rDA
x1rnvVXo0fzWySOUBANgutgnRQ1jCnApdcrkrJhSTtBeWK72/+x/EZ7AXWTI/y7GUqh/VOJPX81E
9uP7ftWqeeo8FFKXMCuZxSWID8ez2aFGZVyYLcvtNk4dfhOQrpSPsVG345QRfC7zp+qaosOfh/yJ
1x3pd8KxMTjpUFxx/gn1jX6pEsTG8HXqE7XryU/xPNpAoeRmDEEf2315kT1SQ7urge1AO4GTcgHo
IV6OWyzFcruSWKOYkfrUhOc85EZ+6MqwQ2GXifi8JsvavnrJTXIFrsdrF6fC0tOrMBh1kRqE2Owh
t1oB0qdl3znmfzHC5JFPxeg4Bw/RMi7G7N3VhuIB7EDKmv/iSqQvK2tT5PAkZ74vt/2NAMksdR6O
Q24Yfi21KA1qt5ee9EjSFD09R2aN2J9cKjokxjwUcPDHCwvJOzGj40CDsT6SB12BICKNOBREaqBM
rDzg4B00WF0sSd4etHd/Lbtd+v3ixSGr5Af0sFxhjJSroq5u5xwkpdvXHvM/AcHqdisVugB1FdXR
FqHwj++6XSWbsEv2d6oBJ5BgTZKz9h+NZi3cy1DOpWueusAbFkjfAWi4uEFzplMD8Rki8juxSUgI
fO+NKvoxAp4Ukuowd55wSkF2U2lIjQhY1y5232o3VlvVYesNZLPgQ53LCX07tKxQcRiGYd/0qnRi
Jf0uAAGhCHvyo4wdxnkVMlCCggopY+pqEQCjJrX39ryzDCOptyu684HojVN6687U+Wm0hMEDUDF8
1b9VVU2TJZYGst6Yptuju5EkA5SBpnzDEoooTq9YDgSChVcvm0dlAPkfqwXD8KuE7yrBk6MK6J99
067ZBonN+YBVTRBuSYqA8sYbbuL4pCrV70xiEMIRC8VxOEQvJfIGn9wJIA0S4Wn6pViRTP6Dj2rx
daTCRG+ulli3Y/40JSQG5WdjfwVCAokCyQCwpoJiE9GAcg500oMJ/Ej0m/VSpc7HZqT/7OEEgPP0
Hf8CYpCFztnDEbzglAc3cBYnn34dJ1OLPSzIg709dGs9jPl4MP93vS/stKhCLK+hjguFcwr86TIp
YlGHK9pg21kuP8pdZZ1xoWSd6qpgvTyPez7dv81XvOCVKlPzzgaBHSeTI7O+GPUAGay3UXeECGIK
eFaA/CzIQ1gHz5pP/eBTEpHgu0cEQ/DWNNjQEKBwEqfgTf13oh5Pfo0Bd7XOW2tEeD2sUuEBPZXp
1LyoJdKHm7cFCkgYPrNaeNZxJ6I41ihT1Z1j4CkqG++6FeLkzxwrqA/QLr/HVYsSQAFtcgn/+cfh
nMCvu7M+UBx2ASlQ4srITdjMeMoc9RjZnFMKa48LtXvdNbKpwzitjhFzYXjQ7yrhj2JbRD7oTgHQ
FoQSFwdmlMa8+xxCJCwUUj+dNQK+SUfZ/ls/bB0k9DsLUWwvU+z4UdX4WZ/QoKE5OB1ULGL0G1lS
onNkdF+eLqmvvAdJ1jzItqvp+nwV8cbLw239AZWxo0Bh/RxHbT+C+Q/Zfz3gqqALzdNLTz0GciJZ
FszpsaysKQJ2gRWCDGA6CiXkyYrSAqv6Ny6eYy7YANSfv0lzhFxyuWVtz3Q2a/dN85Q7GFm+l2Ct
DiKUGB4pSfwgXhGUHlK8jcl53+KBufy1Lwsxy+fefp0/bTSLcRPulb9Kqz2UA/11T3hfGuEGdNSy
InF9BCFcAYABPR01LwibilbvaWIEgz1fhq20Nv03UT38xjXtodWiSksQK3Vd8CCBUbnGPZsGTBPN
peKcGFQpfU6qbNkeTShV+oCuMxknMaerdUGAQPg+kbP502z0GezmAILoLmvjTUAxh2TvPBv1gLt3
+DonolPJFMwN3YLgxzqoBUgJbyzLNxGwq5XMyfMac/K3oPPN4XlvclRJm4Uj4QGjbNQgbfkroYL1
nc2eBR6y3F25Cd44JWRJkPfU2tMPf27gsepIg7vD8ORNhvkD8EweJikfUOkHjEb713s6KshY91im
gunft4l9LgWhpGVnP3wP7TOcC0A/SI+LkTzoBfchimH4d7F1DoCGP78Xa90i8PuqBaGIcSAIhIJi
zYv7MV7xNwS1E3iZfqDsy6fESnScI8WvK4UiqLVW5ZiLwUyzqc4x+uC4VrwD4BZsXi+tpB7JsvX0
QsNPQqqkGx4n9r7xAuuxoPwoFkBzYmh2h66/4P3UtqjJK+Pij8BPK1kxgGhS3ZCIDnlpen7QWUC9
upl4G+37DR3IPrieTxKS9WIwMX1RTqjBkntSNKkkc4qJEEwFo0DKTJRSgfJDcDnigC/6hJ9QnBFQ
xm2OyqGNm6lkR+nVzWFfZOUfyxs9DWz/3tu+OPYfMbT1e/mYjvt40S1hfCsJ1PAji297F7cdetVi
JF9lhECtpzhLJsscrW131diGw5sQYutr0DjAVRgdYPT+E/z8Q4MeGKCNxbXF3i7oKJyGOxkvuPK9
GkFk6Yec7PD6fLU4OXs7Umwm8avRjz2u5AVuzh3SwyT/AB7EBUyScZZEQeQosk6TmiGvcjvyIRsY
1Vb4dXxM0f8WQXtRl+JZnQw19xgWUIJogiiLdaUl+wsodaeiZdGgat2Yh1OVgo0Ttg8YXAjDkmNn
nYUQvMMURHNcH4KKwQKBkFg1S6/zyshjeOvecbwx4/zELhfBCZFJ7hiCvplwx0lgB2EUuW1k5rJb
RsXh+ASlnHLQMSUpk1lgxa+Wgs4GKLcvnRQBmV42vLJ/1qkLMdzUGC7XqLInqboj/E1b2auWGQOC
QCT93wxfapnMTlcXKJpFIuMinwPCxlwyrV5NgQ1vDIH/yNQIOzAAUKyzy/sSAdfXEhFgOJRzzxww
jTjUhR4ArkwRM5yQk+sBxvtgZIar/8gQYPJVbkkgXf6Z31cD+eEQDE0N+Q7moausMXr0wQQvsPpb
Qpx1+PpTaddagyN4bjIvKykZuYrvu2YAxt8jBArY9MLBVDDZEhzBM0/f22lkwWsv+v1tbCbZofqi
uE9ECuMAn5L9Xr5oMo/zvZRZ+n6ZXiElpDgWXoblrQOOUz86uon8mWZyVh0REUi9daW3g09zGVdr
g4Ujbl9T2hfXN2jCxc+fmP/nomRy6JNyeo24b3lZ8PYNvPKgeK0WNzhcVNuMUXMfnr6m/7+4RUY7
yp5tJ0kDHH3pttULKEm89C1fLAHTBcgv9PpkemubrirT4zOMtsuBhTWDH1ZgPYqRCLZRmISWX5Zf
cWha5QOCcx6ihtUiQME9aXxDwGgWBmhzphn1T6e2P7FHaBhkYT3zV95cAi4XQS2qqJO10W8khLBG
V41jHLr17Xk2vUtpYfmvxs/hJ/yDxuvkLTBQVPB3MowWjsPKjBFk848tMxsth5w5R3UiyIzTun6+
MyYA0jwOSohGoNbyLCGw/T+E+66gMphEwMFOJjEL8Jw6bGFvOep9Yq9/Ixv3t/MQ3NcSdrT1lp14
tIKhoC65iptFJWnd3PEf2gk5+yBScwSdom0AK41HTFluACW7fkEpFSJWad6agD7n2ZyMtsMtcsXx
PxUobDY7io+0NO7rCbj7WL1Z0TazT1nqm47Od1RllL+y52D0hAT9sLvr/nx1G5H3DI1hsij8nZ5/
YOZIVnEkrCvrg+ivOn1/psg9RfQhfXVXYoHydE00c09Zk4lfYimRAdRuhpXhzz1d5j6mD3Q6o4O9
RCt0yQTtgXd3qAKskrQ4DbTZnQKL5uJP5TxvbX2qFN4GHbWpmKbTM+bDTqlyi5Llw4vgqnQFFjxh
szNUYFQh57PK6MpFZwqgF2H1HHDM7cRPyHy+T9prUTtud+M5IZAW7LrhL8IqQaygpUC7dnvk1CyY
ZV09U7LXky9A7g44gr/IwrvQsuKsgXWF9IFMK4SdQy4Ac9LWBnki9QRq19Yi2exgcUaQvfv1soZh
uHp148EsYbnfi8mJoBhbXBcOau2KKITIqdhvDTeYN3f2N7NnVMZ2WR030t0GWb2SAsXjrNcm75T8
5oovnibHGGRjqIPalUZdLPqaw9+XtCCv5mf2GNMthpdCoYhicyzmmIzh5Y9USWihijZ/tsyHh9oB
QbQlQJdgMlhDT2djbtVcJ+xkRpwihv5u5B1ugHSxtVHm6Wx3hMFtvKXMgclWcoIBWwkCGuPa3Wix
/ZAGc76IReVo6aA0NJDa/YxeTiWOMbyhdfTAoBNRTkgt0kqPSLzVOpb15GiH1d2xXU24CVGs4or9
EG5C1WwHcJjuwD2jc1MVNv3kHCPv6EdwSVxgVX+4ehzYQ3o1VMf9VgRmwhJeXJnw6Q0fmpRx8Pya
kB07RgqpJLGmXBG2jtPi+XkB2cRLdX+ee1v5U99PO9DbY8Ofenhx6zl4lJghHS1lqIQ8Qyp64ekd
jIh40EBsizAKnncbZQvPoj+09OhkaK0pYnqbJCDWSg/u8A30NOgetme6BVN9ylfll3X8MlgRllBG
p2lCnE2NiGd2d8lO4Uox9N12JDC8idYOjfmG6fkOo9sUkD1d0/72Lfx5iLahWRgNvnDTXG/ODrme
pF6gPtli0E3PkswVX2avB15/FXYQvUVt3gbDvsw8YoZOtt8j3jPxHYPM2xC5epCAwYbovrk5l5mh
zQYQuKEjqnldf/NN1ZPAEkM6WJxM+eeDT8AEC+tPuyFbFlBqnQJ5eNVJcaX9Y/GwdsBc3mkxGGaZ
y0zEzzudvXv7pu43wVKBN9dH3KceE8bz4ZJwlMaVSbh+Ox3MRou5G+RPcxgdklFi5IOcStLcqQ1p
ueqbVgB854eMwoXjC3JacpilCswtZn8tWvhthlKCj+SAKEA6q0hk2q4sCdAW5LlapSunto6+oV7J
q0Dy3RkN1DTojWDgw5Utyg9j3o+o6VIVFpa/JcnCQzukGp+GfWX0w3qNTsTVI/UynnRJLy3bccpp
Bt5987tZrwZdWnInT1LtDsNWd47ghNWfW0OuPctPLZfMrC5Y2PT3VipOr2ReHthLpDr8w5u3BwIM
mppCA5U4dque4bz896RW071N/mAFmwSDaD2pL5lNg1n7FkrhqVrFbGlQztJ2bLTcQrZARkNcudcX
A7e+9zA5uZ75/oCeTgJBIKL8gU8Ym0ArxCdR/DiMQ4ADIWsAgLMRe1MBaxXliYwBQHVFQ89QiVu1
naBd3HaBprQirtQFf2boQu3N0nsM/UAjtfl3EV0WVM5K8xyeUdFOY2TqOVt1hW1pEvNeGiV2Ytoc
kNAIyDXl7czSe2OkkBBvd2w5F2XNYX8mGawmrjSlxIftOb5C+sDH6bXNeEofV2DfTCT8vsdSYsei
OHcWEfTwzhw0hS/46oy4AbEzC0dO/3Edm0baEjCfz2gAryRKh5D6lYKSm4wNKo2NPHNoVoiZj05h
z2/VO3KzXaw8SzZe4rIViTNBVRJwZcCcInRN9WltVgXq0dKjHPQDlpRe+ZxYE6/uTAKrqOQ/OY+m
PFBy9tFpeCFNbO9br8hDixhZ8uBhhDV5WterGmOsSPWRlCXm8WS0ZcH3KSFx62/F0FhL0teJX4kz
C0Kn1t2IOMlH+Y8VFFP9X78YZuHW90vTTJv1y5aBoJM3xoWhLqO40oqDId32InpAqp6FxW09M4r0
nsWY8aKfdnPUsXsrN/K+Y4rnpuLruSKM5VTWZlZqnt3JHZ9LTckyqagWN+Sf9XL9YRqqtbMZSTIj
zNN7nTKVU+rvKLAlb6emYm2tDBYepngWbnUn6UOUG3QQbs7Qm5f17PC3hRCMSxym4xcXsG0pInay
Ynj9VSyuzY88xtXk8oafFZzkwj/h68i9jXf5MBIF+1FtoqlGQrf2JLtvfmRMegY0jLq6XcWV/qiA
9Jz+cwmHtatMxD9WXjSMo1B2z4GdjBL8hDuolQGkVaHFDiGJTTQy2JmXgPlnOSpZMyRJudpkcJ6a
uSOZtA2q+lMiPf814i4RHQBxViRlfuEzGr+2DoAFMWpSiq6pWE0jkWVI6MGazTSvddww4xZ9pv3n
l1WIO2MntU0moKyIth+eA4isP3UY2+NEqQHfcwFPtpNNgRsxe9ERRIiJ7rJOeXtOopFV5HLfu0AY
RRO2reHerLJTuarWfcOSieJ/dx2PFqQdyWx9zdep7R8N8L0GSyb6T1c/UXOaHImpbfYpyjIgO0Bq
3i9O92A18DSbRPIkGBP2sJbVa4UgWNYLVCQOKGNtJYR0DBX0QL1iGkfJOD+MS9JCAzAuhEaPTA+L
99LF25AtXiywxBakfSz1KKr7U5u51ymQzfLLFEjXlSvk1CKnL89gTw9uY93YNL/dWUb2ZBwmiUpm
L8lFcFUdemLG6nAfAhuIINN4El6fLmiD5gyKU1yCGfihcOErFrdqNb3tDV32Jqy4HJJjiX+MWxYD
hRDXpgyXTPeWhiJYpzxlSu02VPcgxNVLWXQXpNnTzn/W+jUSZLAIZjZr8/f5uV8xXpFskieWgKLd
SDGSjbevhevHy+kptDVVqmtQdAp2mH/9xnN79jZ4oceFKfSxE5gkQIBr5zWsnOQWq+ghpwIw3IgC
h/DjkxI2R+y5Q6qA2c6y65JQxZBZ1cJf+31+vK0eeWnRqlg0oXvgqthbvh6OPQuD6fcWCgevJ8TQ
dYpzaiH+Bjsgp7deqyVV9R//BO+Wocb7ydTsKZ1J3BGCDqhETEqnkBuWpOMnCwl6yXugQqotw7vf
5decCOGWcxARMdnbT47kq9L1mpgCtgDVVCliYOBNdCDdU7u/a55155KAGZax1yL6wH4QoT8FGShJ
lAvtq4tBJ4xjBEV0Kn7nKJG8ZOrjQaChWD6Rxue8/HturTQ1mYmK39TeqCPB7cDi4Yq2CBNV0ZDG
IJrZmJM+MJuba0D4UM/pEm7wOWkNweTSbpjvdgrEfI/p2dVpmwAU1slnLUA4dmWOo2VOohQz3Ojl
BPt+w8vvJMJ9E72AYbAn9IbXuTqGqtYiK5yVN35IXnjooXPx2/vdVttjLeHX6xxVDfPXEZdZMG90
1VkeKBYba1t3iyZCEkvF+sVIgXOosTqrYufEk/emb8gqYK48oBBn2zyuxMxJTCAxg8RFQX5NQusi
oNFIjwxkRMd9g91tt2w5w0iG/SrlDYuNVZutUU1b4yB8ehxnTJfE55tdrBIWf7hkW+viTdcOy6tQ
7HwsfKwtUVPJLmeym7OdiaWfqvvzde5ZiQT7xykvlD8hv58MzFyGolt4Zb948kChPR131346tLok
9pjM7iUThul8sLO1Xit9Ds98pyyZtK7xpBOuaMKA65OXluX2o2Kl6JGhND+GGFf3jwXUy12FkzJ4
G5rHl02j6usFV58A8Q9zrXim0wISfQMuWO5ZXRB2vAUrezob8SPUpNvA8sTKX3lpc8g82Aa8wlmJ
chqEj6YZ3LRa2m/jexlbqDM5D/mDwZ3Chg0NzGmP7H7K3vhTgBYvAE5FgJTSUsSufOlNVwQK3FMO
qWMPv4DeA8HMZ0ivlYltN0+MqJjYJ6wvlGLYPnpIk/WNEKuMsa208pmaKpHMr+/4axpdAexoopSM
m+Emc6MJsNfRPc+qIKeErIi8KX2DI98TBaBX5mpm9UkOkp3YxCJ/VPkQCGfys+9bCSPfmQdFhwzD
RH82lu+APuhZrDLjFpPjVl2GG6Oo4r5aMpXigk5Fs9WWsHWpEVFaiMnVFa9uo91WKW23MoNwzJON
Ye/y90nH4ezI1xX8uaB/GG4CGNDtOrKbLU6hLVe6VEfcGnudYb1EzFH5owSgp9g5j24Ec/NuDPN3
7THQiA1Zui67ncYrS5Pe5XFo4FPiS4arq9J03ke6EpknnkZQfVJ2zLc7Ztt+LyoH6pLcj2wfrHN2
XhJK1wAid/YrygUDM91Nh7kuGMspjiC1Q9OxMGoTgCig66B5WZYo5KQznMrv5/Mf4h5wwPYRKbtd
zlus9tQd6cfxuQinMgpHNX9iO/Ost8ukPe1ML2rcar9EqDYu7wrIJoctp3Tb46Qb8jo7C1FMFh8O
TV7Ha8lxs0ufdN9C5y+7LODqld5Q3h7JEKL6nEAf6HXs9RpYE5bOs8gAmsSn4fG9vCRaKIqnz732
nXQACWn5ratorgI/Wi9X+t8WWJS6tRXEjvax778ENE0TmdqZkItbCKHhgj6S7OOoCFyADg3sn3u6
ukFz8QghBwYPzGl/MlHCnEsq75BGtcIGuJ1Azn/rFGyZqDCVEOOC/U6igq8qsNSWnhtqutvSmj4N
GVkW7zfZg6fFewNa8JWTL/ciDSS87BPnrIp5T4hVRrzGKSIHa6QMhY2bMvYD+qp6nre8P0meM6S+
RjS1Lu8vqdJCOC8tONV5rnP8ilFRIcq1lEYP8shy5pZwBoGGGLSa6T4iJ+Wna0Z8wws1zGH8Wu3K
5FtsU7GN4YGDJp26/6uC7t90HrdFQhJ/RxgR4QbkC5yjlGgI9OuXiQPgvwsUN8m9v7A2wmCUvh0L
ph74Zjt0R4OAZgdawAdFu43KNQMthvyAevv53KADMrWznpRbF2y9XdnSeClx5FB8jzjB8Vfg7342
iHJVfrwMt9Ez+dntsHCtCUtESCk/pEJ5TawfBhbIwWM+MeHAMmFsJ36IncXFUB97uoWbXnCAJtPl
ynwEv0muVQ4J8wezFD8ZdNIYf6cPQ2ksYs193FaBS1OVyVAzJNXGGKwC8Ed2s7ncfenhIeh5d1V/
P98ha7gFh6U66RUcyntAnwTDL6RI38UhpNVMzLGny30m++Q+mC0p3FCfNbH/WprwRCUp59+53g3+
oajcEvMKJMdNdddel4z9zYI+UXEfbgJMTzZswAqMUj4Bqc8wXWmWxirZeCzH346gpgw11JEuhzgN
nAis9Rinxfs1mc3u+70sK6K4DiuqDO5uL4qh7sFqFWwSdEmZR5rRcF5GoF4AUq/TRz1X0pLezktD
Y6GGGfRDKV81rr2NaiGcN7F+lCCVl9CmL5EfBHHnEvpvDaph2aU2rKAbUJCnx2lrUzK5oWqsXbLj
Ka0aBe35pTdqYiCd1tQN2jLJRJ/BWlNPjJNYatM59KmktdIv1gazabhXVNBfB9bwI9/q2Ft7UJYM
FQcbf70aUggabCzvHUz5G5s23LOROvtI8obwTrtRh2hfjZMCFkBM36hNQBZFbspf6MKauNRy9bzL
drGhgvlBwv4RitZb+nncrG63/RbTxPWyzSf+SDkML3hDTd+vMrJF/PdfvjFPUgcMBPXEqnGX5yW9
WsbXQU4zK7wXwFBIve3tpvXLomRH2eTJ6YToVtXujIvVPdff9GJ/WDQtvHBupb8Lu2M2UAxOowAo
LgB2xBSwp8mbx67EuEzqJeETWjgXItNJGAEZvkliOrtAzPTeAWVMF9zOJe7SdqwmsBtppmc0fn13
dBl/H5KhMXxWCSLo7GEUGwbrbg/OJKz46DsTaQCYcYpkVbJk4Naq1Ovq5kK9z4IRuQP+pqATAFG3
Te5+PQLU52KtmcRoMqz7g7YwkN9KaO8cp5R3di+BpnDJYBSS7vtGeLxQAI2zVHtdhaySH7g33OmP
O/WXrcC1aXCh9J3tROtkSJ2sG+tOn6OS1BMpESIoStF7ggbCk5e+Th2OUPizqLUGDjguKuDauCnF
9Fp9aIOLg9WLtgv/siSDGxvth58GZuGk6YVgOLE4YBez439bpymQT9S9QtHW47BxUN2OQqwyoWI4
AgtY/QVlLq0utYrtKwRc7BUvMjuZ6aZ58x7XfniTJ2nEVKzd7+v3XZoUKkobEVyQ8fQLv/EUYMNM
zF2fdAxYjbC5Z54/lOcA4n/ViotkdWNiN+JrCsfz0+jO9Y7j9KmEz7mUHyql3QOX73iJCZuyMbkX
6bPx3nMx6Jj9uVMD5gqu84PYvblMRBRfEyeLv/S0WXrUqOgk9eXznaRdDy9SwNR/ElcY6W603cxk
mpSoUJC3Vu+yDuC912A4mth4JpsSMyejyCrcR8RnyYCn1nEhunF7Kg35oVlyq+TUL7+y2mIa32xG
aeEIKKM36/OThREtYOzic25axPfCFZYe7rqpVMvdHyfkRodGfkm/V8EKRenzjuQiWmPUgOepd9Yo
dRdE8b7sSBWwht0YQv2kLGReXFAsBIjdZLPbvwtLMYV5C+jyCWRI3Ccm3MeTMUZ/Rvleo63ykZn0
o43IjRYZdwK7Z/Hq+hOq7cBJAk99epb+mO1LAPlPBq5GtMtEDQMKugB6g/6mP1rjfqA8ZG+442QH
588vAgfDJonfvBq6nsQ+ztLPWxAmhiUHN6xA7+/Vcca8WbX/xqKRC2UWx06neZzsWWBdI5eYJ24s
M4fBLyT32+MQTLO8TOXrnEuVG7ZStZN58KAbUesey/P3jugdJpJZrvB0Sb/eEYc9igrwb+q+ilrd
bOdMlLJbgBCp5Byf3v9ncN+FUS90TcuUKamAn+dtAyMu/N1X+9VvHuIwk6UoiBYlHvJUY8Ti1QZ7
g1t3YInZWXwFwqX3fcIvrb83FV6SWVdJ9NAlh6jDGHaz89lAo8MSMn47MxFcDYE0cXHRcskTrs8Z
tWh/otAYFkVyRbBOyshMfywZNFEbqYYUJbIbqA8ysS0Gb3DMcn9ZF/lHJcQCuHCsjvPgMlcH+Rxk
lTFlEIjkEC9JN/PZBJDsn757jlYuN/K0GyScEtUxzAO6ygvDjg7FzrcdqC1iCvxmk0SSQSOeLu9u
S8l6jjjOu+4npcfI8kBAbDZh0sYi60CwzFR6i7iezClCFCADiU9fKR+3sZH5TubGsHQ3ZFJq5i/T
NCimN/JUrqtTSLYpLXFkbn1hFFb53mrZkYGlL404j+SnazyhjM4Zis5UVWJXQAcMnoppZ5KlUHwV
BgEM0IpeZv5D6edLUROKvTCQ0wpNhNrlmZES6+28WPhhBd28ApmWREslCwkI3mw7BOzh9uT/StQw
EJ6C2cTUQFFDDecumSZhzsGNCxHQHPZf/utIG33PtdN0MWDSR8+LQtOh1di+Q++9icCkZ+AH+Ti9
5Nl4w/Ez9i+aFYXxmyIGNTxwS0uk+epaTvOz7e/gFdsC9TULaasOK6QC4yjREcGJD1t4UG5RO4bW
xC7U4pUI+HTDoqxhTg+m3X3EvlLRoEVznYwlsaA3hTvJk0RMRoXC0GcbGwidyPpI8RQhrp7mUikK
xtqzAcvxJaSUKaCzYyVISKwg/HbVFONr6seCdFjEyblzf7TIXNwwoX3aLdV+Yz4FnAgRQA/MzibB
9qERvNiZpGAJcNpwXeSE1fy/YA9jHjtR8lPqvU+otaYrRNnnFar5W2CfBpgvXnPrv2NSg5RIwkZd
/fCDiqMAo1Z1YbieWvqX+n6YW+27SQil7KxoYNR1TVUE5mqGmlZRrBzmkyjmTT3iOwJrTJQjhT8C
2sMoTIWJC96gYVlv55C+yWtJQuz1PQqSEW9auGy7q6HMhSUjHBSu6Rf4oc1jD87SvDOafk/9Bfdh
eB0IfX7T7zA6uEL0j/9stSk7yTktdfV2JNDJbbqipA0+QqYOMcN8l/QGelYSqHIc0YPaXjDkfFx8
+1EPvSgg2EaTlT2o5PApkfojjB5MZZCm44Y4vAcLMXc8hQCuGDQUseyjNcj4GYdb5QS7q/2CQxDK
qQQ4rSzKoCn6/Ui/SEn/Nii05dArUISumpCV1wwXv76585+bdSiI8WORCfGmvbem+vhb9lZq6HWe
XoPNn0RgLPMeT81mu/2ZntaznCqQivIYZAozhV4GkcnQaOosT2K3oLjM6sew7h5D8jmHDxzfYiGq
PO93kq5hu4/+WawDi+DdTfG1cbevHIlk8Z8dK9eI77jWFVZ7sryAMM++3jkmgtrdRfPjS6p+m0Hu
JEtpTDhqOCyZLAxNV1xs6IMgJZmeBCQcXPpDSHjpiX3ujxwkeSZXfaD0uHwYQkoEtuwx7n/09892
TdhgoY31n7QHQNXMiAqMvfFJC529YTIr5ID7yegztQzs9R3hO4oKJQk74zeFVv6RdeINmU/+RaU0
tL3l/PhGZGaIX+41lGAntxBWOOeHAe3/7n2VPXea/OXxisIjAweSWUtYTb1fvRgZozReXkMWo1l+
MB35anjMKVeBW93iMJ52Lhm16onjhDqv62h5bkMvKw91ikiboqmyT4lSj9BO54AwcwJnzOl9uvio
I3sTcBqdpz0WAwD0zdNkWz1USemBlS3ng2wYScL3ZA0v0NQ4eyXG6PstLaoUaGxvVOc0ddkfRW6j
58alhxdrJkTGn5TkjJ25UFqWh7vGzi7oKm/28NKLj1VTWYAIgrycUr7BVp9bAxRHs6wNCOSdMef/
43WG2rg/lRbUNbG+dqDixiMQ5caL60ktyymome7wqD3EgBIP/1BklsP8racA6F6SGOMc5Z9d3ghI
2qTpSLKgCrCWHbjI0axkqg5y4eZLKuT1D1vJoiYQ6rH7iK/hw+fmU+dnxKKxSZgixa0+TAXBPmKy
d6y91sZ9+ySunDOlc5GYrmrWvOTXar2HBTMndUuwa1vsWOy4Jx3xvCUCrY3JwdkXUixhLAM9a6AQ
VOFjkVZ8glO9wOjAWEpLIpVEghu9dxcM6WHExb3IFuKAamYEWFpGOLj5J9py+hDkgLaPWx6DF8KN
FdHWZTGAW/bTr9tyK3nifpgw5sBmxnfwxlW6nisZxC8LmYyJYDeYpbwwXPWo3mVWNMcQIaIDwFS3
j0v3km60+jd70CaW9C1NYA5JrMY12Hw55+Cu/XD/CcfEmKDSIKnIWyamX1ZhbjcDVN1Jvmvs0RGe
XjzXYSNjbznsj/O/Sl6/Ie4lMh1fD6rN0Xwaz39V4AtbHalGrDMGNsRzGH/XXzeCD+jywv5ohA8L
tGxzgvMN5nESCJtpVQVycMprs3D28J96V+sIIJIatK0HpUVYvEnN5HD7d+Zet6eJ8a5LhsHkWodT
Pkw3eJ0pokEE20vDuFG2cTLRcGvShM9sFjh+iTs/jtaJI+xItx4IqU9Cr25vWwzgPJ/f0jP+FIC5
f1GIZVpfpPDZxbkF88T4s3vPPWQSSE1TXpV9kcZV2tIMBhi29UdQGQauYyV2l3hA84MgS65Rvqeb
Jd71SBT9NeKJCrkvFYY/6Sazl6t76/Cj4McEqguve7KNZAdvMlRImtv1Z5S9VE2tGFhdC7XdNe0U
CsT0dGu04B3dVKbeKTeeImNs2Ya6XWpfKIFpqdJiTjo0fp7fbYKyDVcjOFvXcgLAaEG6fHxnMIuq
1usZ428vK2hM4h7iOMO/VHXi1TyHUnbuEIJ8g2s+9EqFtpqR6TPoTWN975SywZSRiWeLfrT/5mOi
C/d+Sb5R3iZQztg2a/eme3mjj/pcWQ8nHg+iSpqHkZo9+HqXe+lQjLa7axTHsBbR7Wa+PlFXTXmy
4fb6yfnIIDk8sSjyfdTpj/2WvqjcZQ1GhiDN5PpQvEZwfhklBfIz2LsS5fwXkEZ7kKRq5Tm+dNNM
f6IVylSAuLjpEAMM4mRo/JJViHBUwVaw5jpK7CiGhk/8hltBGgAXJubU2A8MB4m5Z2nm/68ufDJu
9lKmxitI3IjCljUIw3TbB9WEJ/8y5Al1Ob2oNzGAaJMdi3KPLJ5Eg51zFTJ140sq3TAE+3Bk5RQC
7uBAbdCQM1XXU0Z0T+eTkmRIbFLCXTyFC4+oHGOfhEEl0RRqeX7/BrFcL7fIf2Fym32RxcvAXtFl
6iyRwwNTIzZv0hyERfS76kz8H0MN/Kei1pxGRS6LCj73kcYRTH9H4wFBNj3Ay79im6Catgcnrnqw
Iy5FWk1Q7D2yLPTa5IJzqFW/0hyLTZl1IJFN+EdMytX8xSCsqv8ulM9n42HK4ylQeImoc7Q+T1xr
iwych13tHvS1zG0n9DNa0RnFvR5vLvY9KVaZ34S8Whxj1SB3Pukm7XPk563VdKU0aTJliX9FdXHu
zC7mZwzFhLiAA5oW8lxIAKqsb0ZJ4vEn0vEB1V296AkKw/EgfLYYuL+874G7PmP6d/hh/nVguHkF
duI8cclCLo14L2SYqNJlCggVdpls6uf5syWNvHj9chWOMhUDkoIaZWGiivoiE2YYpl74k+DfNelT
NbWwOxpREpVSQ+dEPqW9UbzJNLJ/u3IeRnz02nCyYk4lyOPVQnY3RWNc+KIbrb322zWHTVnIb8IN
JrlxgM6gcWQjbHj/8DNz851ilasx1Qivu9Wu3CNNvUbnljx/RRqR+NxO5b6XYa3kPyXjIr5QF6g4
7GUI74Vx6owDEK6BQ5+hFCHwwfVIWST1aIo1PnZVuTFbljkMaZ4NPpaI3yAXdKiiANbRQfIugYkZ
XISK9tPF3Yx+PpZeJFjieZMg1094zjoDe7ApEaGgEeImzU/FGKSukbqRgE3cv1eDatdX1zGgjB7l
Afyaok04E2apS8o2eR2kmyxy5iOt+Xj9mb32IuaMGXnD10VsUGS2NkInPsdaMwSf9tiT24v9hQ24
oT9H4uFNLDr33tuuraxRxs50xoJ2taY1m5VSujLdyCnp8iz3//MbLmc2jgMdv9qw4p9Lfj5U2lfS
kk5d5gDg2CRq/qBaNYVMLhDYlWKPmPwd9C/mnfH121Gly1m9Lqe9akpc9Xwb+5v+Rz2Dyk0CD6LP
edLzZbP8HJUeJU10QP/5sqbAUNWCvB5xhv7WeckwOXokcfDU8zbHP+CYu1nLVhlmlbOx+sJgT45B
eEkQ52F+cxcm3HVRgNS5G438Xl7xd+W/9h+TMWDgjLg8nwYHfZTQb8dRv7NhC8/L934T+viUBF8e
GccZ+anFyUokBF1EX15vxdOy/KgeFSIkJRr0ZKTMqJSFpPrUfX7QQuSaLEssT/KQLRAUWcHQC4PP
zTwsRJeNFWknG7R0ieJRpQbxJxhwSnOdZbjMkiqlbQ1HyHOLzR5vhtRHiudysMcFvoUTAV9OkBpg
PswngiQgDXoId6j017IvxAjcPJhYJAxpAcGePmbLXNgI49Ym/qsjJur1Y+rDa8Vof1N9LszO0oOY
o9g7xvex+PgiuaGqjlUp3XKCpFmkR3+RvhY3x5q/U0dOzy4k2pLzfGGoBghA8i1kKoVAY+PrW4IU
Q70OsOb8Xex2hv0dY4bf7Z0t2tHQCuGNcw7GIDk7YWmZ8OtAEaXMv01ae9oCWUrUmsGqccorwDrD
nZms9E28UVbZViCzzE8TCR5Nbgg7OmGpkcTCJJtDyGo/UabLJZ0YOwOLxHP47g4O2yVBqKHgolUF
PKcv0BYVyrwe6wM3YFx8WapnqJlcGhUdK5Ns0BTvbZEVRq7gyLhiEElW/9r0IZy09Tp5cUwU6+Y4
tFruH3TsslpL2RBlG+v/ToNsbgehNwkUldkLljVlN8Nn1Sibri6QdehSDP218YflTvBA1cE/yd8G
6DsUonxEFFlyYmWXjKTn11ksaSi3KYXvvV+sF+cUYJ/hO5bc7LqhGry+c3mVn/mTO6EzBj4eV8+7
k2+TXpUojD2pmRLiiI+yFPFcLvzlzSaX6LkQJaP/V8FCdtCLbtoVvI05xitLs8KzgodCKrLPfRGg
UbwZv44CNedp7Lnveb0o3xOsHNoeKPP/BRiASQ3JDuLaJVTqqXp1FTQF5L02jyotDy/ZfzHdBjWM
+hL8XCAxTOV7Bq5HK7nxv14w+XgVpTzzimt7pYnxusUDtare3FAaw7g+hVgBmK2a2TMH1+v2t2mN
BasA+DJVThwAyiKRJ+lIQQ/fU26eFx3DOnmX1iqTwKXcHLW8zTBfjEDLEKCtcoiaJ+GaW3LtD+gL
1GCKDxAs0I5KFkwSl+URs4bwycDf4qI6rbl71dZfdC2nXIPvnJfulEmq7jbj/9Hvqqkttx1gWute
S025DcVnLNZCMsunmi0Ae5qi7cRIDTv00sp2n5dXcn/A6/1ypoxKY0gdjQ3pyo2IcdxGSM+4y+FR
LuAGV9sLKhTwBCOO3xgwIyv1iA+cAx9FL6oJ/W88AotgxfrNAwB6kjLMCoXT2vPOsMBj6/IH9Lf2
ujlgld8x0rEVNmeHNXSfZ6h7JU00rwULpBzSUzuoeSwJqawJz0oT8kp/yqQzlnqeuNK8mg8gI6H+
IkvBLrHLIf2ObXhjFtAFU3uJBOpFA7QKoQf5dg7uHlYFR/5TPRdIiK6V4NJL7esyzawgv7tUWMaD
nf8UPVaYEaF76fghktKkLSqMFr/Y224JwJ76htjHEyMx+AFsHwY94bDY92Ov38p70oDU3Gu05jw+
E4enakuOsfUqjifynkMK6l9kJpR2A9XSVsUu/wCb9RxImUEK0uIp+FNfVeeXl+ukNE6FGWabOM1M
V0N1VofY51oTuIATCX+O+x5paqJu+V1CZVKget7hEnqinhYsgCbIb6Bkx1QwljGrSt8xrUzbw5ea
bCMBEwfhI84Q/zhj8bJ4mZUk4d7u1Ez7UX4t61W0dxnihd3tIfdMD4CmZhajpnEGb+vNxYb61jxI
7V5VDo07fTyqKAcSD0Y/cnt1p9ASowJchcS9UYrb09z4kEs+JW6C7A2//aCmkKtBnex76F+CsOV7
672v+VmS9ctyrkzsWkAy2v+W6Xtubi4h30XfTFdd1iUz7CaM31E6/CAj7iXPun1d6rhsjFPz8oCb
hF7in4os/vrlGpSif0cQRoCV0CLcFrme3q5mk407tMh0f/PlVLCLfGoO7yTrIp7VbSp5vQ/8XYsb
BrV1Jda1QUbDH/8Xsxy8r0iJFcj5hUmGDMHW1afLkW8UdtL0RxmzrQf7bTr9mqfSuglv0+WrC5fR
CkKTWbPQUBPDpziMgJzkGrI6CZEdqkvE0OQYQAoPO//CzgcNCA15sJr0DUQNuNQykit1SbWG+1fV
xmpz8860kI3zkrTBx1YUptRb89AUv94PGJhpNF6RfmP/rPmSy7cBnu7a2wMSYEWM6SxNMUbF3JsB
sEv9yjJlhgyATdSfSaa1BHqHa/BZiNH7jnrDvaTqRh99fWs555QC89AXwUEbkBZwsmbVgLoZHOaE
yp2ArQmglXtL1vJdD26/vB7XwfFOnaZtQUPrPIiCSAOl3+NAJ3IDOCF46cd2pop6rsgBAOijQjIo
oj/uBz23VZMfcir4obiuplXKo9/7IkF/d0ZoMmoFvyyoFiFto0hH/c1qj1eHqL28sj0nF4sLxs0N
wMIyxPmGChG3l5ck0tU3oy1OAS1lJBvWqwWTN/TLlBsdn2L+Qj1fLzpsN+yo2YPDa3jpbYHns18I
RGQMHPaMTw1k6d/33ASoSVplRwZK73Lh1Ik68bGzUuAvyqRRI0unV6Uii8fCGO7aePHFgLpNGLMY
CgUU7kRiE38Yl2yR9l1/6cp90xU68cIM7D8ecRkijygoOYY5sUfTXK2GQFy0WmSdM8acJUS3eMrI
tqTlxzJfsNu7pVikm3DshT81jZjI5xPHZFIXe9i0Qlg5FADLiH4Oj25cis09eu7SgBETV1cZ3xdl
I+Rhn+h+TIuicc/c50AuQHZWoUk1CYHUbqfQth3efc4k2kcCeoeZNTNPjWLMnHYDHn0fPub70hnf
pKAkU7Z3MgEIompHhnD2ugMIzKmT9qpd3fwSCec4XjZr/iRuf8oZaBnk3OukK9iNoNUwMe8EBleQ
ItOFp2oE9Y/dwz8ofio3SMw4MCljMMLe/DOpINnS2mkO/+VvjqMAWOIA15/dmdl7WztsAzwWMDNz
vlo5lWxqYLGJOxgqFTA2QUft8YOrNfcEYdOLPI1VQhecuiRpK/fusF1ppKuHJuqtINJU5KKWTcTU
2H6AEcjXwxPrNZjpyNzucF/086eEmBBdVA9NrNk/Xqo/2ktDihewEYMkfuq8KMyEA2e7tAB6fmVE
BQnUeUfEhkatI5ZwXcqa0MNlseUODkskxtzrmquHmDMDwdtyK2c42P46vUL9y4hGpXysWf1698QY
04RILbg3f8NgDFfauK8nrtU71ln6lj+Kr19XRiX0/HepIDrBgnnF331XAf7n13vkZHKZlgNqUtCG
89/gdI+xxot7gFsKAjMrX+/o3tN3CzJq4akcv1Hrdq2vGu+HY0/SVeTOncao765+nqNX4iJKn3TK
bct17o3b/Bih/rOlqhGXM44z0z00wMgadBmeSwrrkJpB4c4UUEon/wT8G+hKSESPs8u/JDPL3FAr
Vztsmz6iebBZBZ087ju1WaLuHF/QsWkG9lFXh1J25t47bMpL/D//kP/AvHMtxEq++vo8AanUub8s
DGw8LoZT1ZzsbptMwD6r2F6Zle1K/Jz1Mzg12Q4bGsFf01RQrerkxw1w7sCOzUS8Dy5dJb7k7Dxt
TqM2NwCB84iYFw1fkCYZyk8BnUlgFUmGyHCtwLQYMO8LGljD1XtUX33byn+ZA1co7/J5ELcy0nlE
Af8VpoqAsbGJh4vmbA+lVSOmwRuUdJoNDWhKk8ciPIa28qvNu8j+C38QZ4UmPnXabayjNhXtmINj
3dORUqRL3QHeupvRVClhGjGaDrG2+3uuT/ROlotOpw4vC+vdbpbdTedCgYz18cqjvlVUSJ0EgKI0
4xtOii3+8mr3WwKje/aGsVLipam8mExf2VLfVasRbav8dbNaHjLV4MpzUAaeSdt5ZMxlDoBdwXhB
RV1+bSXToL8CRXsMpECXDVJQpq++9V3KbT7X8nLTh0a8t4tY6e+HEqg888qHPJpZBctIDagTMRG3
mF5wQvzDSQhMNLW+i60XNIHEDuTv8xy0aYX8Lycayvl8HfWLLFtND5zmukjrEtuewgwtudlJPrNB
ciaaP6Qdpj7nbdpDp/jD0eNLdRFpIDiT+vlWYHmETEyey45EVW2sSukSDihRrO7cV/Tyzx7ey4d2
fZfl3IS+gcqZgYnl3Zx6x08JxNGgM3cHj31XoAGgmQAt0eSHf3Aiu4s+PgQejgXYsIvE5uHlf3p8
MHj0qkvamP5qvaPice2tEGbYNCYXkrKtZIE4wEs2quz6s7yrUvRivlFl7sxHMMm+9irOp6MnhGe4
G3E6L8VksVCUnyOMf/8TDH5sRjcn2/Fs8u7daj52Kx5OdsbaJa68OOSXGSWgKepkfPAEdCUMmOvr
hhjZq66eFnmE2JP0ghdX8zQtMXNo6NlWXjTuc02RoAYZKnqKwb/3p+oC3cXeBCDoTvJOfAR0JHAS
o1BJ7jR8q37HuBvXD28UmwQG8490yrMlmjIwJeAYDgpFNrX2qKCgJrv4A1qreeE9HWfGWz+tTxsO
kB8NK4445rXkKsCWTcvNIF+MVq8AqIHUem2s574Dmt5b5ubWZEp4Pcc9FGviFSjnyDh7X/LfDCRv
nXWLYzQZ2c3AOMluIMU07IXkrt/MgOyTDnpkChb16/sm9zoZUbwlWp5Tt+jx1/OLyZ+Y66cpx9ld
tm0K9Vi9n+V7PliIMBDA38cYrU1XanM29O6cjtZudXrSxsVaJ/1ctgA0JpoZVn+mHcNirj2V+nBZ
2YGMBwFRShuhA43z11cdx0mi6fg5mecYRHryR5yJXTvShh1xJZ0zNz/gsQBeXXEeoa60IKhqkPh1
gx56sJ/BzUkHK4Mn9vne4/q2fUXtq/IzMgSwzb6XdHI+kCUhrFwDYve7ZIZnR47Whoz6orJ51ZXy
SoW6Rn7AiW0M79iAU98PV0CARJu4yUZNMqvaIUljP52DyxWRXqzvKEdxr2dxewcdxKmAYaLjwf/B
hOhowNFA8rWIi4+SsOzBrSeOgJoqDmpWCaeXwuQ+vyqHrPTX5Bd92irhKGAlAHqaCebBRx7SDNkn
0EqBR/GloIejwxTxxJXcQYCDZ/2xpEpNjt14RboA24Re1MUzfms4bQUfz4zsU671KTLqB9brZ9S3
KYXhOSBpD/hj/ZICHgiLkUxwM7TqyiawLceW2JVGSwqoN/BxctSxEuXMlgy8MOUHHsfihGqDPJ/r
uYmNwjfpsWRMR17FAhQ1vlvolGiLTILk/8JdyzPHe/t8fjbBUrMhN2DvAArx//rx8frQgw92KuwX
Dd7ijYbjIGb9sxI9/egxo6r0+EB8kwl4mgmzhOXnPO+nuVvz+4/WK0u1S5CJU0VFA/kpZB8kDZba
/okXWcJiGovLyuQZzUtxVidFqJ7liNHX+negO5CU/s7eqoHEwSrViFnnxB295FfEfpYdotnQ0Pmc
g4TnfHvln3nA3GIydaInuQ1XK0yVh66ytLcu+yBgzMdG4Jv7CXn1gazFtaTOnW/iu5kHYGfNN+vb
x+1mzK8waQMVfvxbEjUwug7VKKNhrO4ZSNLNG59fRECoHB7dwznArweNZM28AP9jj+5BEI2b/IOw
4IHp0GkL7p9T/vQhetAhaTrbneHyaTPM9HpN6xIkHLy7JRxr1QFZjGZFn2kfP3UqzY0HEOlLWPFw
RwOzcwnZzaHO9lAiaDHwipLo9D8K3wYMd12zVTPr8tvOeJrbqquYl2xeFFLMCYnRcw0Z9c1tyzM6
RsmQIuDuHU36bmU837Fl71afdcwxQsk9E9MZ5Ga9vyOHJOGKikwsYJPCruOWqxlIrobUhBkXJ/BL
p+rccQqy2sW7cJcOlcpbF1QaCBZskk+Pi5mO7sjDJ/IrLZgu31ARjMzMOqy5ycdu/df81olDJ3Bp
6fFE/RiQCnk7fmbEnfC0NIP5DGpt+j1LgJ4qVnEnvmkMTQ8wjX/mNnmSDUS+j8y3n/MrLb9WGJMw
VvvXoeCTToydKBAu/heAHYv/zuVoy8TQhuvOyITR+NCHW57wTI9LCKer17ZRp4/AEjS6eIPIE5rZ
zLpFex7Q9q4yuaDi59etXeBeuCdmhXgH7B5NfLOnlwj3R83l8IDYlZbUC6s02WhNmc6/GuJxVy0I
qkCM0ZnNwrkQSe5xGpTaWuhtl8CFTC9YzvbErWDij2DaeF809iykIjQHfdCxf7iLk/CTGBngEn1w
yoJm6oKh0h+lZbzfIyM7O0N09OOW7yHhQtteAzYgiFUD2BaUJIXgeGByNuDznKIbkkV+g7e5/y+b
ci8r80t+weMdpCjHHIzbKGinDewpm6y3xvRwHB0rN/cet6v2jAGap/pXUt2g1kdUDohe/duvA1AS
SWAzqoQHtUigJPoH+upJ6dy8nz4rZvtp7suCBtdnvUkj58Kv9yos4A2OH5F/KI/tJohuWh92qzSS
8M5jM37E2QJzkLWAAjwVS90knRq8Ov7S0kKInYO2+ojVz8p+Nadb+GRTo6PKG0a8yhpF7ovrT6Ab
FucAVP4bn5sKXNQrcPEZLhV51DpsNtpyIiNPYcWRujNVyEYjibluBPAt5Q+aB7EHRLWEfzEYVp+7
XhSKtZDj9FxHW71prQByN1j5ubT+7wpnKYvOim4YB7LKNY/7IpV0t3uTt65PLPqTV7aq4m+9NrUk
P/2JfoasM0tcI9VYHiB398sMQ6Lu8uAOZjdHygSWKAdJbXig3kNMUkrbJZ1HHZXlRslqtnD9+5oc
rLDydptq5JQZXWTxirWoIfr6g8a+8dl/3c/ipRF773Ki1euGpI6ksZv67xXa0p2c/GTQHQiReUdx
YS8WsrBkTVefAlhh9f9obVO1DV2u83TfV6kr/UfMSidv06NiXcQVHQLql23btPjyC83gpcvCXEzN
AWiukPV51BpkN782tPWOYgHxh+ykbtmhDHS9wmQYooo/2jIP5BwSgQrPB88q3u3CqeuCZ3TWiHbc
0bQXMUe7jl0Wzo+yDbIT7sMhHWPpzC26U46iPXTjCCPGyJER1r95Z2mMhle0vPIaBVt4siJvxqQ5
l+G9VYGgO/WC644Hk6xaaev5bWRj+jNd8cs1E5SkiVratFdWczjJ3TNXO0Izs6GVWocubGg7f3eR
q6v4koQ9ZLVCtCvcT4SXkX0OZRw3JjpfE0vV6I+pjdf4LEeEXKPRkvTQnHB2IKrTUE2zx5iVYGOc
2C0frAHI3L6UIDMYE1x5+7jyqc1DpNbj0xC7SFj6ukdFH2LIaLzs3d7gaJpzaZmdqjrnkPsv6MJA
5of+jb7kDLgGIKSKK2oYQ7+T62AuB8JjVYLYDcKweZZKL36ia79Z0A7Hvxvvhuc+KF8hNXsvwMO2
Sct+apknRLy0AlOiLZgBI4vDz7muA9uDlQwMBbLfT3cjeoYod/ln2yG4ZgglLzYJA3trV3y/66oN
sXzbzi738eb6IP/VhWYKI5kTq3YgjTG7vkRoOEumca14jm2bXFiTfEM22Fu/CmtfVlTCnVsbF4p5
KmJ2OQKuOvnp11Rg50RMPBB4eVrMOV9WVmjYIKqeNs/JJW4baYD5RetkbQtMdYGFyATI+3eXw3k+
aNPHkHzdiGltcL8ze/+s4Ei387CsNN1bwG7NmyjsQASlwzJjpf8FVOt6ciN5zGig/SpQ2P/ZYZ6P
FgRyXl74DT7Fze7F1lqwDjEki5YWHILmQrxLTMt2OcWAMi9regU4zsA1/iK/CrVyf6UqtfNUusnI
jS2xqRRXComsQdh+Jgvuvt3+ZxCKfr/VTGjxd5wcZTxU+F+cy18btyTDCG0JKe88O0nFiaqfpOQ9
twsyR5aV2SqRSkXBWVK2BZUZfAmvPP0kptzzfX1/fJbGS5E5ieNmjlsiOuAY4jFvEDHIbZ5nww4u
bdfskClr5ND6EUCGmBso4mLciUTPkgAxkZUViN54TePhiX6PhkYJomvsoh9eFxUq8+93gJc4tnqJ
yNs1FoO82p8xybJHVyDaZaH+QWGGvp9n9petQzs0qPiaXPoWb8+Xix9ltXT3KuZiM82F07ftKO5p
QnglzJjEYa1nCaYdAFrULkEcqOeNFUNXuizomJwNg+ovR3MB9sToZ4WSLKJDfQVu59+MFVUz96mD
5rbsf4KL2cjkfqcykgaBEgnVwEy50B+BJJR4VSLGqfxUU5/xYwgNE+iOIaTQbwi6HxJQ5ymCYPDG
7CqYkF2ojIvgRR0Er3KGPETp6KILQX96pR4qET03O1AyNpKFeQlC+FKbpOzmmAGpqwuCsfN/yW5M
EeS8DrXU+qy5dZl2mDF//wLwxAmmfGQQX4Z1Uke55NWRcsPpEshjvJEoJb8hNtWGVwm3uKdLRDKf
uk2vtohgPOmyAWMbGc5eRnLwLS+/qwjbrwtEh8A3dKdayCxlzXHA/f54NqKZsKJcw5YZqxoxCU4p
Hr+yhVcHPVYhIwrgwqDfihArJ/v/voT2JOZCiQdTZqz0ctyULMWGrV53UYcxkWMvba734SD9brFP
e95OAycH5zgRV6McA+Z71ZeAn6Kn6UZ+pLIe7/saHKcxPYrrX0jbfWOo36h5M+9w6DAU1rVoLRr2
8cfCVvgxdGoTrH1YFaVK0F47B8W7txC85ckkuEXGlh7LeKBgmBWmXMQ4xMBgfzsDyIbhze4wYMeN
Ll6IquWOM4IiA6fyqFJW5uNcADQsQrJHwwCp/fUSY6QjG++bP0PU46wNk+PGsBdbqgk7rkRzlu0g
3DgPhR0/6Uo6+ZZCx50NAWW7YnyViLGUVetA/V+99G2Gp1IdIX1NIS95kx6OzrxiU3z5Dodtu7+j
dG6wQ8K4QJMuaVzChSxIWdNHJTuojrWCqAr9on9xVkWvgPuqDx6RxjgIjcoSaTJ2ijEO9hMI33YY
u5wD2D3+npyzL9+cdEP1HFgnL60oGuzv5ui943/NGgkqSAyNSSPLZbwLmzCTn1XndeQEccGecA1j
MBPje2LxVqRscXeQ4pJHEoxix9X872taS3yaMnN+Et6XhqxD0HX8fH1PTlv3BmdjJlpsT9KvAz1l
2wbMQdrRW3WBXJRiHRmHCFmEF9JBwdOYv2XvfoTsp+69ucG38zPrh8ZGt2UuRG6xGiYMs9Dj/Ybp
2L+MBvUpq6uu5msVX6CjT2OQqicpPSbapFK/BfxlZzKv9Ev0epLtj/CFCj+yBOTmcNOHnzSc6vrl
iqtdjaKJQR269I2c7Imnm+z7EpXheggtW/I4SsczHKeZ77BplEUm3k8YKNyQJNF3njj8X9oxFvZg
WAib6GhWe+sX8Q3+wV2kaNhZ4Jk9KhQxkS2X5lnHzLUbAslofe08FI6nB1Kpvgy1DpUnGXxEVYO5
5nt11strevMn9ZZq+d+DbFZDn4lOlNEukEj4ON/r0JWGbl5IImSJh/v5vXuj6aLFvUfDtNT8HfPu
eGm358Ue8wMtV3UuqHgGZ1nL3uL409KWc8C86CVApkzfDTvrxWllwN6mCy90CbFncwQNJarQaPMO
Q4AMGkWoZyxO1PtGzP8Uzt20aZPySvzpEuv6vamdyWmqpWrBtwdAj2wEh5e1qNWRP6mOuydKb0U5
59eEwxZb2CMNTgp4YqCCGAimodtoxODKk100mvXW8JfzaUgHddSJ7eBsYryVSZEFQUBC9l/a5Yne
PDn7vxfKl6c8OS4EiJdLbrpQVMCOcqGW3Ii+2bAKeCIKpk3c3UqriGlM8q4yODvFEBshxHLHZejt
6JHjydLh7A4TD9Oi6xO/QR/oxxkicvox1YwJUPbie61UUx0MQn5EqUKp5Ffk3xztEK2GAClDlRrQ
Hs33TByhYe3dqS0KOTQSwmPWdyv5+jfYEls7oMV6hKGDI1WODJHEjdz+FLErWAjCkqEdgGy5FgQt
aviTg2Fg8ukEBm3AXRoEXF9QRJdWCSQwXctZkOaHRinI8yH2aTsJRx64J69MyXgyAFAUH2PmEJn6
ibcJNRaarYzGfEoqNHTLpN/JTxrrqSrhHxDBtWydN5IXc+zQt5MRXDuVg6JyQCJFrdt3pYcFttNk
cRxyW/6qMj+G72SFesjyC/Ndnznab/UecGAVOM4WgtXgca02ls+AZWOKkpw9aVIRQMqTkiR9t9AG
na+N69AH9d/UkOpbneRHsYFI4XbFAgTRTIcSqZIrQiIUmWG0A0szCEWlmP5h0E/+qPBVPnKCAJvL
hKDK3V4WUggDYWdkZJqe1hX5SLezpXoMpB5eENKPEnM+gUfvMAuvdoGGThExOG8mvR/yZcWqqF/p
ntSUg+PIHMT8vwZtlLHdn2PiH52AEcBJp3kTS58idnLtwu29NY8B5m7SBqXU5Le4Hd8L6lZKieVX
XBHsBvwx2JEuE8sil5UNhVG3IgHrEuic8n0FY2ZV8ITBvVhQQf8aK0c3/ZUd13CT1h4n4C2waJPT
CLh39BBQV4RSk96Qm6Aut+Qkzs9R/WHMbRaLOjs084h031gdlBahl6c0lApBQlwYJH0Z86HHhwiR
fz/p6hzrzfOWnJXmskywqpLLshzcLPWG63GPUH8kiOXrZujuMdtKuchHi5V+RzzPCP/Cu3SH41zd
nogU496CWoJD7zV4ebNlvy/J6KCnTEY2I6FYOLUA+Eah+MX2JY6mbcUtLVpPpF4O/1Q/FlQ1XQAo
AtLaCxGFVwIZWoygAOYrjxQuWU1MYAt+rdYSoioV9TIHCjuujxYuSRCx4cMhNCyh++JhVl+cvNOQ
8Y0h/Kl/hRVF1Im3ODkfgokkzpnZDoBG75SXS+vlt8MQq0NVKMzldM9X32FfVHsP4AyBW2fOhx7b
aEoRrZ1mBnUPwZNlaERB1XlySlbDPeaQnElrhpHLlSmHOnDVb4oXjD33bjiJ2JZ/blPYiCEuFSwA
mq+SpSIHm2ioi6+mckRDUO+K/ScyEHlm+xZCZ1no81sfhueKYc/F2YMEPn8/fRuutxIfY/FNQfIZ
UWnCQg2zJLHGO0qAsKAKZc37riPgzdJU22OT3ov/iPPGNhNek6WCvGN1iWL/f+BrfFJPIVsHPBYB
wWEekL1QrYFmVUyYzzMkBo0hby1K/321T2LGAD2v+ZKXtEKT+XFnyiCZOZErfl/OFSNKoq501S4n
MEUzU0Hkb9zJMTBnFReex2DyPTwkQ4zWLkEFi2pZWDuNm4OyNSc/UpFBJA8Xa9YfOEL1PSOcPR1f
k4Mq1ccS7wPKHO02+nv/Ss2S9W/t/WvOc3ItFzoGM7yEVOHsL1Ed2VmnXgeyoNikKQpD0ApyjOOB
nqLsHhyk0F9qOts/UOtvTRYqFiBKA3BQi/xCIz/kekt4baScNmf86EWJKx7/qlYrlY7AGftQclA6
ThY2pdml2XQT2/IyUtvzACMBN2XXbVFam47n3+EpiXlniEecja0ypLc5suKTXw2v8p+QmUUIs6Ck
cH96/5mX+P3wqLqo9Qp0XU2VZlmN9LzBIP7H6VB1NQXzaABaCwl4GeQEBS33tVXgikUnDHGFoU1j
PGw9tu5ZkJzQwYnZXDnd6aS2EWjUvUeqfaQfzCJv17PnmXtqtqqUeskQERHvRnMOMWln0zORFxVJ
RwPAPBJgSBywcp7gurV3TKa/zExdUbD/VpuLFLJIMBMk/3s4XkJ1alM78n3Dh+e7yORBaK7U2Q4e
4qmF6OIjFlctaelIDerIdHPlYHQkFJh9hiyNZpwk3hYDTW08K8kTrLZQbrTwiYpNTLvivahCLfQg
vsDNSdqgXcA4P7SF6xusjNSULxqbkMjPiyWRBnRASYF4zWXKPC2h/RwcqG8507RqAwV/eexhDTek
oZesuKNleweXn5L5OZJP/WwE86eKVvaSANfUNG412fLrl01Fg4NrtWQRKKUPsv2ht0o/no0OvUMm
p9Tc4t7VXgqVsWLIT/gVUMpHoP2a+f/1MVUUg6+PXBdZBWD4z6XPDkNBs/G3di82bxh8icGMqpLN
K8eCs4uhFLyfbNTg5iqIpirAT8shpM7s9H6lovAqEUV0n6RwUDCWy4dFv0CuhBRR9QM8qpatptdJ
IeKavfy78SCWTaWcSKJ8A2KivTAUTs29s6Qv/FgA6LWztB+4XKtJWFWXCvtb39/Q+9EUz/sYgEgU
RxHhmhNY75O4aBSxdOazBgXMvqcUD2eKInapxFNbcZDNjKeuQm5nAUnGS6PSNXocDhPvoXbz7AdW
FvYIAuRsH5IjKUieHl9IdsFwfkSZz6blB9zv7qc+VajNoXS9sBetCt9DNnIfNMlZ0dL7Z0ns50Aw
muoS49nUM2AmRTk5XwCWT+0t4X+XqY99n7IFWu4ChhpMCZ+NmWiq5Md+kRnLj1AXdLFKT9b+4PUw
4O8ayjgYaSZLMDCj6mNbKDJ4/5B9KsyZkZkw8FuG9b0EW6TAGmgDVZ4k8oDpoF6JtLsRZH/XuRRd
m9sT/eGDqgJxEGzKQrSEcfYsx60+rzdnLI2MZT6ow3jjWtOttjm7UTXU+gBIu3Dlt7STs7tJKrSF
w2KhsCvXFmx136QbyVlr28aV8JK6+g10EIu+F2MH6MA1y7MNTgsNRjo1/rqq4TvgOedSJY0E7lJG
2b84eETzRNUInfcwENMU2YcEHXKW3z9hnOSr7/969d4mCNh1SiKFLPScXfDZOmJkSqbTIWoKGDJK
owm0GRbPta2WlJXqYnjlXNSkTg7y/8KpHLNmkJxKBcGgHh0MrjYLrkCxkwEj58j90tVE8cggwE4W
HoF1LJsEOgvKHIOJv6pZnyoToGgb8/+/OK7xSbvtdi5dfYx/VLzpRvti3OhgP3crCIxOo2wAw8Tt
mjGD6RrHo85Er0OAwoR5CCLpuKFKzh/BmqLWGai/+crAf/kRIsfITrPZWvAzwRkyrqRg86p2fFNu
5qBCO1hLTrTgqjoWGGJkO6e0e4zo6wJDOcFeyYYcaHbAfJXhJ+fFDboBU6PkAnYwEq4mFwlfE30w
3BPnArrfmwEMQD8G1u5bQkNXsoviM4TuIb72LoY7udG/TESKblR6bJauCukeHWF9/qrfrszD2KLr
mhm5QtO5Dc+DFHA57mTqAuoA2cVK0ekyOB0jibGVnCF1SMC3hPF2Tum7rQJdomVn6O1qMS0OILbH
vNJTBlBwo3fMS1Mm0e0/msInbDvMSaeEK0GsYStjOQEDHvddeEzZrhag4NnEebj06IrbQstg/KlW
xHi8Eyd5K1g1W8g5tmYWXvphxuTk/7MvVbkFscPcarFOtAKW+xeW8bjAh4VXnhZOeG2+hDLjz4Yz
S9kZHUDSUf/T3sVoNQavWYC9Mh2nP10TXuXPE5QvKd3k9xTjvSPhMbKV2xFD5KFwVy7qDeltqHZE
61+03rovJEw004k2T1pdlYXKvokVWCWHhWspd80SwjSpFvEw6ITK/D2ckKzc3wdjHTm7GEfMYbVn
FT/s6tbKgGG8poz6oiAZV6KBtEGhxAAjHjomap2IZtNDygRHUzjePHR51K4P464tVVMzIs8g4Z9P
WqMQaQQc0sQujVL0ZcglZ9RaYN/+1h3Rn8k8IdMcKiNLKgoPufLwmaxL88VPT3riAaBoZWjycSbb
TEt0PGqdcpNn70v8ST1ghaeoC99jp35WUF++aPcxJksZawsUF3M00gRMGdZMcf3OjQ/enSXw0PPL
d6xRm+48F1psnATe45F8DzBo6Jl0TY1PMqGQxw5k/aJ02634lcbQJPr8r2dAVe+N0dmZss3Ji634
BzyfTfRh49X9fCQNd5VDFP9bcYBNe48mNKBSjWR1ECAjqNzz9oNGGlc7bxyBCp373zAxfVWRZMA4
hVqkFtYlM1MBnQZww+F9dYej0KWicd7iQtfQDal0qRqtFWLGgIKHAKiO7K633C5OWBl5b6fRZwCl
qGQQSzh4KzNGysFISJ4ifAbxdxL949SlyT4u+Rh4A67pi6NwaYXPG0fR6K0xAvXTEsGMmtF0/cpX
N4hMV+b3A4gFOFxruN1I4uIYtDnCh1UQG4ZjJoWl+9rzjk/ekK3v0lOm/8xf+QNdKcfnRGaXd5WU
Dquw0bXw7mZEU+GcgVphR4g6IdNny37aFV5KbkaVmelUsGjIPoR3ziulRmil2o2QuGFUM8SAArZG
YNRuwijCf4BoxGxMdd0aHL0Gkv9WuyEdW+MIARMP1Aj8ZaDzkPSaWushrYvAjPmc7prfN+8g8PPE
FGP7/DU1Afq0ArB+pLCjGQrWUT9WMPlPp/beGTg4g49xnc8rJTVthNwbZDg3EBt+WU33M1eD4HhX
hrJ6385DQzmFaN0Sesqz1QULaDTnKLCL51tL5EU6hx8F3e3b9l27sOwjt5mqxVWknFJbH/Rdv/f+
XEM38hpslngRlqyQlwdyO5UJMrBkH6i4RsfxY0WSyxZEjnRFcLqjoth45YPs9wGviXluzHSZC5WK
MLg/ph7XBr3KqmZfaFadbv+9WjH3RuhXomijvbW5X3kGXOJR4dnWCz8TjlS3Ya5kOkrzugtZ/TjK
0XBHS7DA4Vsf/D7zriM+ieqnRVfZwrNIu6fUfL3I3pjSX5KlA0Cs1o96P6X07tvmp5BO4uA8N6Gf
Xo9oKTZ1GpPvC1BrdbuhAckeFzavDH1yiUL10DTXibcAxO0lwCn9F2BwZWVfm357hGD0jA8/Jrod
+91DJRzL2znD8/FbBOuNS71SgmhpgDrruNSfd+uOBdI2gFUe9GlGLmzBbMzZSdd259fTfCvsQQtz
xprnLa5KIWe3K7F5vQMMbQKYiwfFCNFT92TSxmw6x/10pa4HxEQbVbj0HjWGomZ3E0sD9M9mUXBD
JJ/hss8xwTKdS/WwyVpHrhOSEVqYAxwvjGQU8MSzpH9if5p9kUFoezqy7XXDTT9u8uLGNd6TyUzh
8R34ldPLwZ+oZNCz+AgaXJMy9J22vCxLtKore+s6w+M0YQAegkQkCnOzUGLmoqcZ3B5Jpho9Am/y
CPddR1i7R4i72TLLY8D8rwgDFwaEx8Z0TE4ZnYoSsmpGp7DyJd3m2AqFb98v2D0NyGwS6qbfYhP9
T4uh4zrd9nHKKISE/7c8xkSXyNXq+Rfj2q8CUgU5HDzam9QwbKhnFMwdlJzif12C0W9inaoi1g+b
SZbSIULUzzM8EEdYwOOWzVmVzYjZCWRLvGU37G6crLRNvx1Xsnx2ZjZp9mZMgJ43tXed2AvmkfxW
i5vCjjzPOa1itOTbnvZJjhBgsL+dugt+ackdkx6Y8dBvg6HUgqSgFDELawAoJX95m3shmxDkKsfE
YbmK4fMxkjT8TkzWmDmd2pS58rQgJcFaadk2OICDyT0pWYt2pxV+UwRhueatHHMLO27ffDq+U9YY
GvOtSnY4/6Jjx5CiNvxHZ91a4qi7ZCO/ZMc6QcpWeZdoofqYXyhwdGGNQSwmpMqmQtQFgk+I7Ii6
5jlLXm/ZRrOJWuhSmWU52Ult52wIIGsOouhQhyMQUOK0165zXDJ3r5Da/tT89N1m8zN3ygE1liz2
XBjIoA01May8hoo86d3lGw1uqSt3DG34rZFAH1YnvdzR+RsDI36wqJ4pAcWfKkpQa5tDKooUwFBD
uJw0d+qWaS2UciXsbAfYLXUOzT9F8h3CmCb0NryKdjutZvo8zx0QDhepKeOWOdLjGyiOIqeBvxSt
hureeGxrilOhzLZ2GYkYPa4kl9Afyz5U35out18BMtEIp4ia5k7jjWnpxuhDjgghOgp8qgEXTar3
A7/0xU7swaLb7L5uR4AKAGyUMIYPZOMrxp4vmBmNprrl1oJC3vhDszuY4j+qqSo0K/dnO+m2DNNR
JHB2jCA40umbh6ufnEZN630ugJMCPBm2X31dPBJKwxEF87fjv04V/QgUHvFab6ICGIKTa9565MR3
fkKldlIb9bIGaBZGx2PnUbWa2eHbkEvrFjS+kGUkyNhr+cg4zT/ucN45S0A+FLEGB581AmIa5171
LRx5P1G1KBelitR1AA3vdOWo2/NxtPvfj+MYdZkykbV7wKkiIN8doiPr/xE73w3LETcXOtZDfZqf
IS3JlIyCLCvMsPuzqe74v2dhXr6gME/RuUD9fQQRTwlnRlcThi94fCNbsFqB9didkbv2kwkGVf8l
gIG5X0WrKsMU5vv5MO1mEPk/PUthug+BtEd8ZmhTKA7PZJ2FtpwVbzaoBcYlF5Hr0PgSOJG+CeUe
v3XntdJ5W2vId/MEgTSvBKO9NGSakTYP72PAabL2b97GGrB1ww4SmPQAGvdIF36FIuX/7Qx4diLl
ki5WAg/yLmqwfeu1fVLElGJajjWRl8rm23YhM2PljYwB2no2sp/ndWz0cWlPlmavTgQJB0bg2r29
ZhaQqDLat2oR0RGk9vt9UOC9Lq2g2UHeQW4s0KuPRBJQbKpfU97wXws8jSVXjiMNYT1LCqwvplki
7y04G2wf4nodUm9U1bXNhqVfnFEocGkmjX7LR+OvtiJzSlCqVI0JnsNR+GNmlqdYXQOGOn7ox6V4
WQtbjeRyNdv1XA3wlepySld1Zj9f7CbqCXERXn0DWuH118tNnhZVsMNjyh7agRS62Gkujmkhx3rF
2r3Amp8Goqr3etGr9F/4RKvKb1oYASTkjbvwKuQy7DaaF4PU1Eu0Zkiz5VjZG+U/rT+Q6rXViMn5
J0CjAd06ghN5Ql6UaZJgoeSzAS1XJDf8GT/8kBhLUIIK5KyiHpYj2iuo7UEY+MpfcmqZhTZNoboN
hfThdErVJxR8A2wRe9FJNoxa/buzPABGbig8GbtD1YzUF7SWitIVq2syesXPBPbQkOOzy1vNFk75
SvgwW5LdcakDanKgdFVTqPW5xRpM+16/wqS9A4RzwdhYIkkP869+mnjE/zSh/1cqVhmQ+Q/U5Cm+
F9Im/spvpc7mAgQf10Mv1hTS7q6qgnhiFdAilDVwgKSCTA7co2D/NX12ilMQC00B/nFc6u9ZR10f
/9qIVnOt0ykqUASmM3Wags5wXmI4R6w+6nlpSi0ei/B17ZkYGw7I2LtKZSF/2ND1CHCAozqYaG9F
S7cgqIv8S3bngsfJA655gtf+pr0zfkFOMAPGivi0wA7iRy2lejaGg13i6bIemfsg7ptjo2B1i8Pg
wwQqd70mswOAjU1YKqoeehRv0iCiNP3YK6XU194x4oiBM1v0Do192zkUsBDQeakfrkNwK2qC5qWy
a9bQXM1W9g8ZnkeHZ1E4g/eO3obqc7M07cy4c3Rn5yhmsxLsY+81WE1Q+rLkUD3LewDtLvlTbllD
AXthPu/weQEW2+rYaRP6/7XqnuljZb/2/xq8tBSgcs3B44fwI17mL7hazhy8H3Ija7VsWK1ySv4D
Otpv4h/8HLb9ZDdv1tXBHf82eDXcFY+3xjpG2WRz8enIIf2Uf8r7j5Z6Ir/wzDAe8xcrAhMMf653
i0ZqVhmJJgNpc/uWO+bdp8XcGmHPWhwycAwMXSFVTFir+vQ8lsEoV1znNjBR641VrXfjqGyvYEJJ
E/NuzTD3as983vcu59HeL9tlMsItMckZ6mOOrUmNMHEJLPSUw9GWcw1tEdTNaEgfxpY8EuqP25c/
uywi8133YKqGhM7THUZY2Wf0EvVWZAS5s1hKkPaz7JrTEPDNmbWIyJu2WL/gWEUkdEhjK9Q/P/Zy
Ro6LZzPtQR8S8CUFm/AAD/CnftUYiHkQLBym9dDTognL1lT4+ZLV40sVytirpr9uPfmxjcSa5WSc
8uS4iorR+UYSDC5Qy1IupJDtY8GjlIm6Qf1+1BJRxkRQAHd9WMiAwuRagh9H8VXCFxBqf+KV0GHb
LZ1JH/vNlnsjqDiga2krrgz/Zyn7X0/wabPOzATOh5T+bjiUF78GmpAcjnN6jl5PRpqMTw+BZrbp
POEGpXMys/5jEWy0tQ07oqrOpYHZ44xwDlGFa9NSy8rEMn+ENjep7B+QPj0QCuK9VCl21ujZRIKw
FOShlU7kQhXmEIFV8inWEzujG61kfeN/G7WyePWh9pQn0Bpe6rHXedoXRidv9sOxoACjSIEM4zai
CcblEi97mj5QNEMrvvPrM/vf37J2HhV497air8YfW7CXOPm+BGgqtD8A4hxuglIEMQ59+lNc4KNP
F/wKC876PwfWhNKXI8NDSLGd2JNX3JO3VWu0MeWkO5VQj3tBrmHekobnpiE6wZK/r3vt4IE4BFuP
90glTmoEuFR7a1NNjTiR85xL6Q9lH9r5qM2ssvOO+225W+KvLMXclyMPAJZOS4cNo3XeCkhA52rD
afUAST+wJxIOZtb+FZ+4V3WNCSZeZbFACDiV0itVilP473S09z3CzTCTI0spP2D6IAYvPZDQTTxR
QuWlO7XdZ8MGbfqifo6C8I8NxbwzA51Q4dtMIlfByEMvLPbDIE/LDzBrxSwhV+VenZrwEThfH0Kk
9NoqsfLwG3/65ayiAXs6CLYJr40jNQl/v3hvRdeTaWub8IZxkQPRXOkMC9It7v4Fdvs6+JKBGM+f
+CShfpMF9JA6HHmue+9ZJlQJrGE/WGs/S++inHr3F/NhnXurimV0aD+t8D3cLBwC1m6t+N28L27L
cGv6/qCDoD2J4Uf/pLXY6T50slZ3LtXNRvhh+/F2iPzb12j+PAfAyoD/1jaPlEB0k9G+Xjjql4gL
E0/F4wUR+pdHmI2mXpVAZIRnKS9DSDO8X4RKH/6MISUYyziPPdHnGiyLxizu4Fss0hcrUd7BiSWQ
7oExNO2y9oh4u6WBuC3BlZwV8d8xwPdJS/yDD0yQZ9rOCjTjaAxm1KDZkz2BUc/+l9DjKrHoDsse
81ykO2MkH5WSYBv/ynYchmB+5taxvFwjFKyDxW+b5wEFwXH+FBOWLtbmQfahGlquqYeCsu2ZX+tm
NGKmkjnG2fiYPOXDa0IW2mABQDyxJXdkXAmEeHt16I3chs0oPSdhmUzEMBrQeCTZLY1XpYK5Ivxo
lm2ug4bDnnePH8MsvIsZ9vWAu9hH4F+YvFlg7dVBZWKpbd+2CIuRPW+GrQy+9Yh1lqMkWj2iU2Ag
wATJAg2JZcSQvFlwkpyt/6OAfB9mvtCGtIMSUpLH9D+QIxFXwP7b3AUnPbEGTuQ2AYBVaLwAwZS0
vtIJNTl8tjlhn9pzkWTaMdTfrPbLuMf0oreuE7XqN7n6VXnDKHoRF+ldbAFfxtqrkOkKqgUwLnZK
vy7lhRnCrEJ+aQDlBCe4tIKnmJ8ioCa5Hl1U1oXZQWpVH615LsgMoM72gzR2ZbiC+ppKhT5skzeT
xeETBisJfyEoFeDFnWR51gG1mGym+wFAac3q7IwqRsTV4qCZdlRWZ2iOlPpIwwAQY+uUlU1CDpiU
0NrQaY/clPlaKbmz5kRheHfKoFrO/aHwZM9EgcWDr5mnk/nvfQK3qbETvQpUZo0fMZTQSiFeaeip
+Ov2ZKqnpHeta85yVKNYP80Tcv5y2QLyNq8Az+wugSmphA3YZ10UOX8mLA6ffZJL58hSouekA1+X
PFi+h9/Z4AHYwQx8Fg+rvqZgZXunwf8Y9X4VsGe9RqGkw0iSGr6ehE+C+g1Gqc7QIqenVdyy/e3W
QE6d2Su+SoWd/XouFxuVpmoJHm1RDW0BX7KzSAl8O3vBGX99MrnstLgRbkx6w5RgtlhwIaQT7WXY
UM7rlFSdPWUssIAE+amf4luJdf0UQ0yTA3sjndGL1gjBLEKQMvQfJ++OB7OIbykacX5ix+nyl5ED
0tWM094yNFntMnZU9Mbhr+ltc9TUtdfhDUlU16FG5uHDPH7ZRqTShtFwpE6sHqWNN0iPyIO5xC6T
t9MQLUb3HKky9L0Ier6fmfDHmCApiNj5dvNVeDBPkdYZEIAUPxgRK+TmiI5fkXEG0t2Msyl/iZCP
MSI+8AHWpSV20u7CVpn4gRfwiIJrxYrnhzPVkgNrYZDX8W7DUFYStjcQHyfcdDtYfbCnlPECENhT
440UcaTEVIspF6zNkBC5mSZKB6V6P1urtYHXlVJmkINp/SE1l4tvhmWmSGw+0DlsrNEYKEiLZdSE
roZ+9CS1y4NAlVXWtulqRMMfV//Oh+UuyCoep+7I9RF6z9CQ6HAt7Y8Hg+OJTAMTyRiZ+GO0xV1Q
oWWeQJD8q9efdmRnSLgpV+xdt6m0axloslJQY0Psob9v6t6x0Bgw2+oqpB6a3TH9tKfVilZVPsjz
5RDzbAIc9OxfyEqB2GdjO7e7ormmW7jeh9239AB3xgipYas9BLjJQtKxTFmU/b1HB6YPX0Z1TcZ7
BYPfV8tFQjk4+MlAK7fMOTgMRq7LAmIO/RXZNL7Q77HO2Cq5mvEbzNMu5KkcGIc49xgxmWiRWpJ3
J2wrDyA+IHvroztsZimncwT4jS3YtaODGAs+lWrABv1ZjBBvZqZ+3bFr26DU2guRjbPt9DroBlRX
KJJlCtJZaczedJ5wC3UEh8StrP86QBXteybkB8txmXry86Ycq26KAmohqRkU6O6pMe5YeeFPsHpg
Vurvu3CeUaVHWkXqhVrphjH5e+uTzXgV/2FhQKq+72T/hjz9TLsrjkviQYs7VmeIGPqqUHQyKN5l
fhMYLC8u1CvwvvItD/wOFn0pqP8/ZmjvbmILNK6qQK/crbr+KOGloPu8QRu4iLpbf5hwNW+kRcFc
l8n9rI2emHZxdkmULm0FI565NmOMvPtIGZOjvfi7cqchZgOhs4ikGRLPrlyir3tGGvqrrYuRj4Xl
1WOZeyJyZY6tUrIWUPOn9fVDddIuMXKQwMERhPzits8I3dYLpMlKiKGrUnzjEhUD6xascR2npuUJ
2oLQjjkY9ynQbTrp8vMXj9LZ2BZEVgDYvxuBdci82HhBN7ANRy7a+LZibUpdA8O69+oMJDvIeRLh
/bBB+lV/1/FHKlhJI6D+ujZs1snzRJfrdSVK82YMGTwuBJVoNRvhLqZfY0/7i0xGizkhbnUFVP1Z
bbiq6Jn83iKQKXShsSdwlu0DOozsG2dFsg0hg+sRDUURdy7vFPXlgYyKLp93SLcUnZaFzVEBb1jD
pluTD6wW8PAbjXL5AdjvbEypkNltsGywco5nmzeLakFn5GxddkGkeJBFUgKYbgDOnD6kFMprCzvc
931JLa+GBaRcau3HENHWl7UN32RQnBOkN5N6opYMihFEF1BD1xFnezy77J3s9AUxzhOL2E2MriMI
TsGNTeO+sLeG6jMHHJQKaZ93KknVNgUpX7fADRdpya1yvJylUbUoW5kSbmLEylr60eq3t8hiup7/
EfbLaeQQu4x5mjx7mDArZv3i3l62ouJx/z7K5ZVPQDntya7aVnAlJKdnzLGLWduzEt+OwSogK6vu
m6OZ9caApyGHKEpv8ZZOn12Nm4fpjSIYP0fUgF5gyv0jcsIy7fWGhnpU6JuhNjVDklhVD/3WRvwR
+LbJ70aHsExMYrrScPx7pipH7LevVwhp6FmyzGYs18HJ2BSTK7fPFuOeOX2j4xRbTQIO6/0EUO6y
bYXKmBvcW2+mR/q1wsMByDzP7d7k9fe+4X/LdbCfao8CDDX2eCXQfjp+al9iwRb22nTL/sNMwtFD
VByCucDYeKWuEoC++gjkKqvfx6HI+FonQGUpP0ofkHSWmlfwZVxTeB5f9UCnGFCdyT136y5UpDlT
Y5oG4BLoOeJf4swE2N5+0h6YR413OYsqIyHKlLG4mpfuSPM3V3sMGMqreT7AJ1hU9ltZmt74yKjB
432sKQ8U3QRGBr3jEjW9n2BUbK4I0aBJhotLLSAjn9V5laa4vSmDKcqc7rZsZiDO+uhAwVwdI24X
5jXTgtm90BgB9zHnQC1rnRuvUR0t+0q/dt1SbJ/FFciNVYIOw6gQZyzZPLO1zn1Gb47Gr0hlN1I9
guUlQ0gOJ25Nly7w9S9XQoU01kWV5OF75TZTH8vaG+qGbdFYJiYrQZYdUFl7SxEg9oIS5DUEjIxF
28TQsABmylV91kDQTTVxJbZ1oH0OzccdKTUiXI20mR5g7dsrbO5W1fNoobfFF1ni+Mjj6qKXzvTY
iDiywQJe2QuYJcLEPA9qD9QZsuHcv5GfNIjKu2O3n+91VCcSmhIdsRvuDHjFuNR7JFWAJ6wJg3E9
stRypAwOOT4up6TkQ87zSlntqmD9JrF+OD2hdLGJb9FRXOl2vt4VcB0bqrFa2BuWBkmb5cEbEdSg
A4Y66BUIldtaZN9KGhXV3++YIMortdAMlgjqoe92y38Ubaa/9je+jkI4p77tnT8vXhGUZ98u++pk
0rVq4EwdFYmEf1/+UeEyu/dX/Eh8irURT4gHN1A6cnl9q9109aGqFgmT+hKjT9TZF2vC8jx72Zfb
eXCgVUmUwM/ApM0SSjBrUqXJia3PVFJP+0xVYUYmBTH8YWmGVbmpeAx/SfH2ADc4wsobeRnIZZ/N
bPJX8MK0OIgQnrvK1BLATE9zwy3BovocDQbuWJujcuZCju8MBuZ5D1MGyd5qTxu/uvz71xD6LHcz
mMKfW+O43UcxAtxDvvOgFsBV2wkcmRQlUFtAJpFDPCeWZt8eg4ShqT1KMmL31YrmuE5DTgK8UlWd
tZaQgVm29TWDrUwP3bkxLaVZbgkWxeBqdCCevYSqctN4p5uHh7YprecWlRFi3ZuB/uyJipwqasrG
agXyEQIVoJMA6ckIq1J4KOlGmZwTv41Ivhk8/Eko9WA99PcmPMJPzkz75Lr7LkdhZH6P4wbmEuKQ
/C+idu7YDwl7D16ZBHLBqqxlAgmXOqswDKHc8iFWd1gTO1WJRXCPVV1Kf5Ij4+lkiU/oMr1xOIcJ
TfabkhOHhlNjSIJF/YUFw7yVzp81cSDm2kqEmyfAKaBSWcvgHLvg2zi+Gp7OS/MxWfjHQKPJqjME
szfxEvci7hJZX0qEcfVim8l68UdY5lyghRZatLAP13tkAbdcKjhpHdd1OJeaeYcoyN5mARbn5U7B
nH6CLeokal7+P2rZDBGJFr/JGrdaZzuj9IU0kZc+ycFbZYd/dbIMRC4XPnyL2e2mab5ZDA7nfZRA
MC2Bo/9qp4LWbaxav8p0CZQdK1l26CuPXx1YkXtxPdB2GgNE8AplFXUtLmAtCc69Gn5WNJlsiIyb
mREZisbkkuH/NYouDKsjy1WlsRYLPrDLRKlv+zC+OkGXz5T57K61Zev8UPHnv35znbxPLuWk1r0M
jgCDGXbSDOxzaEdNuv0yLh74xCYazEVX+xhuRKAjxv0Bs7KbSFIVhxWHEWreu1O9IZuAp5o4/Qnf
gESahfFJZ56/nCYiKvyxKcaa6MhyYewbUfnhpW4AYCUTbesYP7JiNPLJClzHNvMROLMcmpqHY7BV
JFw2brS00KHBTj4HuQIByY2xQ2J0AWDyGwueNATyUNf/ZdNcgKmeB8A4ucbGoq3UMYlvfo69rUXW
/sC/jetcm4CR/pSSzQ5ii9vwSSmfhgCkgWBQ6Hqha1N4KoJLr8c32RMqHSycYiupqQEaDRC+R/bZ
fVDtKAuwpisHUHa/v5SiQvDOaATHce68Gx6p6e5ZnHViMgBskNFQRf9+U7Frzy9hkCVtbprTaivO
/p8J3JvVDUYsMSscmG0Ex4ttzo0a+oqoR9HFFfAHspwwsE4cMUbVuxvimXCUkglcFLhncaHFyCjh
t4I39B8fCR3T9mkXuPETIkxHLUPcv0nE8Uk7qVjIcFnvUoV3Cc8h3OspXFxA9/xc8YEgVOkrw5MN
r6Gl2rWzvsOs7T7h5Y1I9Lgc/EHV0SkzKByeY2xQpWTqxEe+yw9doIRFu2l8CVYBeY4+yCZBmf7O
Tem3s3oXUYbkIz9O/ipzvVKuxIfghaO1E6Y7RdrN5An5OfDaFWXZvGz86QNURKrrLsmjx/ky7X0W
9dD/MKdIJPZjc+l4X4sS/t1f9PkUwRU6wtVkPEQ0CwNohW2J84lbEq55ULUOcC3tBcmMrLzmM6kq
mnvPc3o2XDXBDNOW2gYA61WolIkA+mSiBTEcBirMYQO1aFSF6UlqMo4NtXjyD+VKqZIam55ZaJNS
ZHixPmgxnm3MOJPFxO0rd4RWN8RA1/ndbqcUoHk2i2xFB+bl3ftRaDrvjhHlVaxPWfdfUTnZFQ1V
1o+jkwm0GmgKfn0FPhIDXmom9P4Ty00LKwDbkJgzJqb3zIrQP5SG0oH7noIIiEhJdseUUfjoFhKc
8HmGsNvDY3SfpOsUpDuUoGlj8Oir8f2ubi4dOs41EIR1LHsFFLOvGNY5bo+oc0wgbSUBLL3qI7AH
7yuductasgZZMs2n1eol+vZCVi5kE8WACzBCjvkGmN3wkdQP9/7yY+V3wsZJLXJrnLU7+Ll+IjVs
GtbRmGvjnUSVg30M/qshap2g5y6U/AYNb0ml6NWmGOuqyYewiKGf10tYOe7+MlT3VjiFRHwb/QCB
H2dkjNBZ3++wmht9lm2MVyXcNw5Ddh92bgazhfZMLA/hffI8tV0jGSQm3kPjpweXJXoNAYL1IyhV
roKT0fgVmY99VRuQoqIO3AqpYe3oo45qvpINjAU+lOfQqocsX16s4Qd44C1atW031wDUvFkjvLfP
2Df4FvVFHGcuIiR1KJNDUFeYzJVaMGY3s+mTKHnyUCq2OUyGqfL/AEiKL6UkdzNabu2DgPaikV7u
gdnoYIuf3t3QvhV6k+Kn7qrAHbbdTwqYx3gY+Z3OY/E7VzGM9XEEeeFdtjNjVe196c5aBs+AIaA2
QUBXSXY/a93dYbs/E89aQ0AmqS6fsVO+oEoE31a3jJarkhus7z0BqCyKCmcudF7pUdjOGqny5stB
Z8kQvmEavbpqSfKtft7WrIcC/UBiiG4USxWVLizUUTx8YBiljxDLWATNCM+h+7gphMVrjdlGkYW8
/EDjXQ/APaei881ucDvOUcMKWEhZ2zSQAVQMK6QPoCiRxKnftirsEfU/dNZL2F9U4jgJK6xJBcri
U2LfEsZ6vURQmZ0O2rWv++tEs/s5ifM4Ezzp56EaIXnCtqCQ/rbwFnPvhe2vRFknWHzGr5cH+Wub
WKLEe+6gFzHBUfg8/jy20MFFxiGraqnHRDWeES8CUtkL5wy8B0q8aUZHroletsuohq5H1sFYLBte
rGIoWe5PqNQymb28YXLmSNKwwSOvRskfawi5V0qnZQt31ObZkoZ2mqrHEZ5gIZ/KqLyOKd1Hi6E9
aNKC8oGlgl0oiAwvSmsEhfYoG9MPl45W2cRKFInN7d5NJrqj1kIWjW9yoBiNAKKGp1KcayyBriV2
jYTr1RmYprwpYrA+33LE/lPaVdKLWG7OP3ueV8AhpSWJrWYvUHT69m3yflrS1StCJlsxmUGmNykY
S7nCAEaQRAx2MmsEl6MaZTNtWME8dGuVZe1g6kfG59a+Ljq1/FqAD/z/xjwMIgps9GTSXaNdgh55
9r85GGP5cx70c5Mo6BbNjTcL3XWfs3KoOlZPpoA6VO//GNS9wCgTzjebMkya4Sk7qR3tsFRpncH6
fKdX+wV+iNUXVmapCh+u3HJWWINy0bXb+F0xEIgQdfxDN5jSpOgR38RQh4P6odCSoC9tjTJ/Hcyn
NTTCoH3e1xZ2Q4Ji2s8iKDsa6gykosXQ9/p6L6ypytqqXSSrq8nxQlYjyp8VZMSKBisWo73iw9ZC
gnLHOWaNtSjgIxIDFmX3+t5PCw7FQTeX4sR4RcHM+Zu8WwVhlgf1/xj6cFVGTi+Ya9/CdF0sKCds
1ZHl0fJJAzzY0FuImfxOJkue0HCxo6AZ+rZ6c8UX7dJwx/N9fkNqAdzJ8VI7o+ovrkKUinjJOCrb
OXkW/IPXlFOZ6TQ66EHgB5ys+pW48iQoO0iQaotfCcUxnKqqjQjm24HyI/fLkgM+f7J5DTE45bPg
IQjhvQEc2KkZe8sLzBIpLcsKxkKl740a0GKZ+VUnc1m5raLFSVf8fXikNdmLvNp5pRivLjgJEZvm
g/YfK42cYyzITHej9JdPV0xfifC/AymjGzc9nUxdDnp9agl2wRFICZKePMrnDSc4NQD71e6jG/pi
4+f2O4TvzpbCYeymuXNTSjpmIJwDVPqdX/+eKBG6ty1tIf8FINOBFBWI9AD5j+sDwgZLVcRtHzyW
luwQfGuHwqjVucLHMLPf6O9qDLEMCJDKOi2p7vsDhez8yptaKEiY0mxTgK2Hq+BQT6mJlUc+Clu0
9pBXRe3lZRHcAfmZjUNhsvNnGf/wUNQbXfIRepxlrwzkqMx/ygGSlE8uKt291JwDYDi4GsZeM0hZ
3Q6u60mwHNEJfykc7KPk39yADbimNDQWpr0BwVgBWyX/fgKaalaS5IHfuP3u6nEB/iziGK6eigFt
QFfYtEpP05oguaF8NXwEhYsJds8/uLU/5c+xkUhID9F67EqKiBcaAP+1u7kV5IEmLg/UoZdRjiAh
kyUJUbt1pXGRdLv0+JDZdjJSZaPU5dyFfAUTFP81qotb5MqD0yYfLwbl+ONd7BMBr8ZqnAwo61js
PfK8ftSU3PUwKVqynR+wTJnkzb0er08W7JaAgZBemWsxM0vFEoFQkZrMeVskw2YxTuEfX0+ImUJM
0pmHaJVkRGXoWuYNj4FTZxmUVjsbV+fsoG4WcvSl58y5QFBoa7g1FQ49HnhZC747y+xqUDdh9WOI
69NgC0wy+O2JQZ7p6J6vQxw6fHGSDy5W+YgLCTiUZJUj+SzWL/NXiy/kVpMf7b+Xy5jQ19sGnzQT
IP7AQrj5yyv8X749KiyMDPKhpiO+WYLdTgnaYYh7VLfetG0WffZmhuDQwWAvtKmzWkdCE0gNxhZX
j4fMtZPU1oMiAu9cXqxh/cin73UANAwYked9Z2i7Yv0r7Dh1FAVBLEc3dKUzvHosenLHY6SzRmtc
84myfvJp4e8DviFx4lTuUpnkSFbqd0dLNN6I0eRlk4uXxSJOC6VeYPIZSTRJugvTK/z5UDipQO8p
xuHovq5KimHU9uauRkKm5SE0ytb3lM968Nc91edSy/VP+pb79JTjhUP12ZUpyQ6QEqHZH3/W3MkX
hpdbp9+sacxaNOsmyMHRDMcYq4Q8hUI7MUkmI4gh85JIvsFnxuR86EBTih2HDK4RhsHhuWY1Pvce
2mtNiHkNwSffoZXIEC2Dzo4I3aD/DyWQyoX4HjWtENu4kMTVIdVptQd1xlPJckoh89WQkHjJyPHV
0adPLnHszjWLND9L/ZKM7zzmlbkD5SktxQbLb/fVk9IeE8Ms4Ntzk16OIGSNxbXj3yR260kzd6/B
5rTs6jWXITrNDpZDcy4treWuodT/Mi8Y3b2NCnWSEhBiR/pvNUY5iAQciEajPPZOxN1/pUcGnpx9
YvMrZL9OL2Fc95GPFJHegoA3oIVRbz/gRM9AYpBDUUek67LiIK9aErRFYfcaWJDMP1up3sLv+7Z8
JHSfFZ4A2JO9iK62yUiw8FFel3whN2WMkFuTAQz/EF3SGiKFjqlBA2cI+GJxgfjdVgCs9aSEG7EE
HQXT81XUgdil1RhztwAFxDEX49mj6+DUGvh4Wb7dfkWxl1xst0xnj2owFzDY16mB/vtfR94fxlEU
r2FgKIU+z6ZLtKzcn6A7iZGTkFGwhQuznnfZ93BZyXZMVJgCoFNxlysPwFO2NyeeOTxd89FTpCeA
o1cKW7BDLuznOUN5W4p0sFPh9B7PKq/zAJHU4k4E75AgCZQhh7SQcaiRRU4MGLdrycMQhErNzyzk
f9VWgBEnxFCCYcTs+fG151yrlXjUxNsAdYo7X/L9sM4ap+KrCFFTaTln3PBt+IjBkIkpMOyQb3Fr
axrVd9DulN1vlzuRhbyXqudB7U4eCMNRu50G+Wqzcch6HJMsYtdJ9amg6kvDSrAphuIN+brZgvQ0
GYFrrCsIkQQ/+QnaB/YJlyU1gpBFt9JzIsDm3Fbx8GC4R/3PdoIkpRjSRBSr4eXrFv0rx6xvebPi
MTjGTyo6vCt+NapkgVLbRyXkFpYVX1Ucuc7Pc50frGGkYFROFPXimaXIH3b/oyJwMTVP6mI2gdGU
frEf6iMz5axm5vAsuh3/Qq/hwic0yh5Pq4yme5ehGmCILN1uRrOedoYxAJDKXGdTX2V1GHlLOSIh
qTCai7sFadzxlt26PbWDLGVl0f8+OXC+3mT1IabDRYyeJcRpA4g00MK1Ed3peDWZ3U3dVGHHR9v+
HLKcwtITptsoRqhnszQ/EDuczVPgRoiMvZFMdl9qAxxhfLbcaMYF1P81r/gMkrhKLi9VhrnCGs51
OoD37OmgvAGYYMMKer8Sxx1BK/pVMqev8ORGDie7iDHAlnet3VWvUz9b9gvGTCpa8OY/stir7bhA
+Rck+etLBqIkgIu6tMHQoge244wSgOMaqzVvrKEFihmk7b636rL3OYP4zaBvc82UnTTdTIs/kZa8
7DuSoR7wX0ZrWHp7nwpGgOlwUEPliziiHigrY2MGqCKGg7g3sbgI8EXwtHsMl+0r5/cxGm3w59rz
RGE6mLR4P0tsfvABw1nM/7ywvD8NaSLq9HYIdtZmDzEYAGErG/8CrMcLTXfu8p23emJEy1AP5/xJ
sDw8oJ0NslzujKEXES7R6FcmSRqtYjTilD455hIfwmEKKTmaZ0t9z7UWW1DzhDNLvpcPo8ejk9P2
2CQIqkScGJVqt+CqJEQT4oIHE0ix2kBO9MTpHKevrDztHx/Y7x+XJ2AFLdZJX8xmtdUQuuUXFWYx
xHAjIoaAaVPO9GK7Tn4Fgx2RCjjpVo1GRLS+upKcGk7CInbOrgFvfL7KOwW4D2si2MW3c8hzzryV
L8jj6EVSOV+/UBO0PRyXMN5uJQARYmmV8V0l4pB8lkmTGKJhoRh0U+CFo17A3+/XTKVomLy3Wc5v
JdAewkb6QfAifS6tHV7N02a2rgyRrw6W1PAnY61gaev6bAkIC/jHtcvKocA0JpBd1FNlt2t+s3im
/amP2F+ydHaf0vEhE5KVlKmbBjcz/TVzf1zQuqGHjydSM/5qfY3jwWNZMAkkgcXktlhwufP2fjuB
YfFWNcNZj/WJrFzrVGx9iedGLhLNPNfvCPHEDV5hdBp3xuLdRBI7BRApcEllLC3PrbCkSpK+IjgB
tGGaYIHWGpYVgiKkryNuBqfySt/IB5cveM0pgutXlZ4npCuUzcFf+cJGuTPdw74JN/ygtn7PNCGc
wKriw7ZKd/JF6TNILO/w5/thOObA0wiRpeCMEgyTGlfuvd5sbOpfud4VkrCP2uvnHtrbhAjkKWGQ
xhN9LnH3upv25k15v/ZWYqM3RtUnVsfxrytl3SH8n24ZLDtIg9cGgbDCZHSCksspb2R+7auz73gk
ctdwiuuxmskNqL58nMTEAWV2jeLJsSx1FYwtXVlCZTJAMJyiHf1B+NMHN0D7y+qumUFoIfZCKdkE
mLhNZMyryXcsxFGWfR5xuly6H1NmuULI804y+kMsAzcEAtR7Dy8u0gklcWFgDSQShmTD5+CXR5jR
+654VTKr5X9wQ/XyPdnq1YK3zcDkB3k45gG4uCyZX+2JcI5LFPYij4qtxDk7d0ngLx4JgZH3FXVm
PhEkrXWPMeLn1JavPVzz15BJ2sg9idQbnYi8EA9n/Z6rXJgYDrDPrR9IEiiDeRQ3fRx/sNBLY/bl
Qay8aPqKoOdSrchEuGKaeDNmRb488cjPzwBVwLnhkqHmDrJKAG50kEpEINOhGGGesqyLPZfRrbP5
s26pPwvsZF+7U5jwK8shR7ifvlDH91WbvujiqsalcB2QVmg24iAr6zplf4K5r+FCEcQVdoZWh0vF
wobV+xeQX9df4Qg7ZWGHgskTAkariCpDLHGivSQqyGeJ7kgC5VIzj6/szkuCFTCSh60f+gUpKPeK
NLADZP67abZ4VMDqvDJQwOD9h4RgKeBfmUk88ICFJJEfw1S/pb+Ummf9HD/1ZHmEcP52EhOcPcJe
Kso0DngtKG45MhDpyON3R4lWBZoZP4HPqBP0UfbO6QrRxu69iiFBXC9hSSahMHWcYPDKIct3v5X0
kw2zQgVVz6PH6UHqqVMTyr2+6AWJjvHzmhPza9Xk2hEygrrMxIEcl29gmdoHNzBM4+KTTQ+plS7s
+Nmoz+Apm1gBhtPdra2WLjmwjvclgT3ze46lUVzUoHCci8ECMGK/jUXgSMNTjSFhbvp9EBNNHzfG
PYCjp9jBAycpmuBOQsv04O93052ICKKIZtQq/0pTUJPG1WLEy6PVjSEkfmcKUhdLMRHd0xoH9BTL
za7RaomsmtqbmmcqLL7AAUTZV7VQZyZ1Ze2aj/h6rJhlL4A9xWOebf6kkpD0WNq+D3e5xcGOZzPp
Bi1/D0mpbFMXoXKsYRMSoLDjTPrX0Dp+AusXGGb/c9lfPYxs2USTOxhIvY6Xx/cHU0oGWYGSqYBI
tV2GeXbTy4EsqqzQcwvnzLb/NzAJXt0B4fPs6MNgup+aetByJm8qoqwnZlcXrjNL2Yibbsi5yDX/
OSzHJs4opKsUSjsH79JmpSMePeL60T+PQzjDsXCl3r+1TkCQoLKkHhrLQdTxlG0+umvyFYzZPzX6
U3yBE/Zs0eoqaQJBwi8umIFKByWt4sIBo9mpwct3Xl1ox8VGGTyHR6VPxSCbUyIJcTOMq5YXlggg
WilpNZHmQLUfC2ZLcvRz5Q4b29y4UBJ1MMe5Pt9FYoIXk0oFXaLm3Ru2ScT5v73jWidEcVYkcfpI
dbi7IT/D58J6yQK9hot9+3MWn0TiKJBr4pusWgmez4SUyjMFov4vmluwF7D8NjX1sr6qfp9PTMWE
cYrGNfXMVYXP4cv7FmjE2Lv4aeCG6wbyTiYPXOOij12aTGhllvl212bWXe/bAz2nkv35BcfB8rrh
wfZ/VEha6RwwUfl26didtFsUlTEHuE3+7bU7owO+EV0p7IKmwxJ47WotJaGicFsfol7+GtVzc7eQ
unMO0XDZOlHxBDlYoRWsQbqabl0dQG4EPAOFlVw2rWM+ey9ok/V1E2iU5cPbJiNC4jOSJfrcxbl/
hScUvGFYHDI9Xc6SGxNcM4CuoPZaqDCt7zwmPKKLxC2kzIME/opiYAPOER+w9Pem81+EIoVK6R8C
XqHCd6cYt8Wf+tQLOyg0x11DLrLOinyiyWF9ku9o9L+6U1k8//hCz+sif9wXrcQWUUR2GTbzzm5m
iYjFz4xNcKvX0mFfbfPrWvlsl2p5QFvAqY2liuQU8dJRjaZ4oXmo1Ao3uQsfuCKDJW5lokmyf3Lb
jS1tgOHw+YwDLzYOsvsgsgdpjoEx7g64YF1oWvpjeKjH6PAxRb4fjPOZn6iq/LQqR69zPl4AwrKY
BKK7KPpv+LEEmuOq8iKSg9UpErcbUvKFJ3W7sQfPIPCm5JeT8x5EP218rpmvpVS+AyMvAYyMNmvo
oNjPnsVRbKrcvLXsCDtJusqmgxKDrNm7DWWwUdc/OEKYWoS+Z+QzAgbwUZW5UK/LOL76icGMv6NI
a8/DB5ou6AcdPLvj5f8acTRDlU+8knWfQxPdfH43/7rhA53PH8wko+KX2LU2tWQxp1cdCjMjHL5/
ndwXqp6eRpjEowbVEUwD4ShIzFCo25NyX4iFfuxnkKNKTi+eDU66m4rAVEZh5pZ5m/s23MFozsNQ
XYWM/D9w7GW7Nf43Jp9m2QileuL+RlyzhehDnOXU5fj/MsbOzWJgJL1tOpUgrOi6NfEEbD//0Kdy
ugrTWIPwA16HDMMSF3iAkKMSCQ1Oesy18PDl/dOq2/mr49/tJ0OlAFmksTWU4gct6lTDfkCFSjTa
lfco6QpS+H3T6mxRcacnlvvJsLpDnoAyrXARuKI33wy7QdOwmpC4ZuMJrSFslXO/4pxoSWhQn5cC
T4GpkJjr6uPSegrtCGknW5ZaswDkRms1aeiWMWVCFxwOopIZEf+ubFXkujRuaEljFsNIK4XjK1Vf
gTT/Q/ok2rHZe4IzhkHBelNVLUg+2qf73XNEDWgA+tDqZf0nQ8F9KZngdHHQBb1qyEvbiSYgJ2UQ
+okXne8Cpi2T90IMIvDZRIg42il/BBKRMZeDLT0Qjxcdt2HBf8nyE9Gly277R73e2jpXELYezj59
BRJhEmL3BloZKBtvy04vKvVmm4//A6drEL+j0eGI7mMOMS3/VU69kz4i+Aq6/5u6w5wJZ/b2A43S
L1KYzVDTN3n1GTWktd/c6NN5iUHix9vJM4+qROfQ7Oxlc3fapla5/XzMz372D6zFRIKUPJcoavYj
DYv+ZwyVVqaJYLz6B9SG9GyJF6vP6YQZOqol3S8YTYvSMpnT7fXeHrUBKEG+iPAsiVTFUe7ITPg3
R1vjkEPmQtOpxGqaHJ8LIlloHSMKeZ864bMfgMwy3Urc08VTbdNNpvmUgsY9vydfeCk0DCz+oBxk
cbZzW/G8rcL9qSbKdDGrUomYDrVVtq/ltTJVDlL4vWqOP4C8VwEn+qg5alPoTwwyY1i7f3G4UvBI
FAVR03UgEkt0+e1N+epaIBNsqdoIqOfJjtlzp2grS2eP8v9e0zBGc7HzvlRQS+c0cAt67s9k89QV
ejSnHBcOvmi9jF5AmveibZUt5IOVkSTRbiwahRNoYFWFLUIBD7j+vK0hyA5lhGE838oQfiAVVW/a
evarPWxyOdK6dykgE5Q/LM8Fs9+s1C+YBxcfP/4IdaMAeA1/yyzsg9V8XW/U1AuOM3gYWw7BVnnK
QSdjmT1EanNMgH49MDLZcByLn90U84R5YqK9mcs+AaQyek2hlT/0QFeNf8rTcszZEMkPBRrx6ylZ
5urYP6pEzjHRumcbQBiXtdKoHXeGCVio+Fsp0FNMnZ8fy4o64vPX6T+uYEpr2lSEYlpge5z4khqs
S1rqp+FXqzo76SS9wDBcpQ9N6UwwuWuzwMmmi9Y/bZF4AH3Ugx0OaPfS0EcMOIuxTfJwnjbFOC7p
V4L2iwhW6qhnErED1dmnCNeY9DOZuIA0N+ea04cd7VSG/QC93YBgLuDxRORmyv9VCiEB3RLJQP1U
cwJ5wJ2FBle0tLoAIn9jsl3m+FXYueA1UjJ7Cx723Yo9qzy4/cfMssP494ZaZWgsi9Qhf2mygHky
Lr6NaXYRp2aszG1SXRs1sxlPM8r/q/STG1f767pY6FlzfU0yWZEqtFs32TRiQfyO+8JowEmxFrZm
T+qxpkw60DIaVXxwM0akD+Y9BYLNv2OH7ZzkJvdPoiy8ytG7VrlwMhXdhcnq4OFiYmcVvMTiTr8y
UJavjt53PNBO0wNMFGaR9PibpWfigyuhG5NRAYDI9b3O6rg+ZcPdxruF/pRKQkpFSVlXnJIGKOFi
tXFRXHR2blOxWkLDOqt+AlTXoI5/zKzb0648NK5NCtGSIDGUCkJVM05FBMCtk2RXtd0Z6b/RT5yf
+xvYvNhkKOefaIeJAW6yD6RTvsYnL10yJMk35uE8/cdDFQFVAACV0ayN44g+o8GhFxHSxT1RUG26
9t2kR1M0n5YsPu8TpKHTG1Szw5myhIBPPl14PxDIEeQz/xf9JIOQq/PXTKqsppYoii44Vh8Tap+v
U6CoKbjkUpS959j0kWZjvtwAPw8eKd0I8awViFuslizAgoKMDhb7W8/OEfnMo+5ckHPuTob1iT8z
9n7onPCnRasLFP37M6EH40SPkXPA9VReIzizf5lI6GVOIOV6eMOGh3eI4ni5/0057Lpl0lcLKF1U
9Hzwmiwjgf/jr0bxciAg2vfkNr9J11bOJIAAe1dxTxGkaIfgrF2LY63UjKwI53AQ9Ce4g9h+PYfv
u9uBHXXFhYnjDb0tVsoT7WoDDNMgeVV3i8MP4I4UF1sxJiw+HEFiIDsy0HU33dgQoUhIglqUJEFI
NdUYEmKlB68dVf0/UHKDIz+jA/30dKk0RVZMKhhX6vOEoi0gABMgNyGW16kty+a5xakDTfJPtJfC
sQdj+TOFPVBIm/5xlpOXs5KX7NJRlkEoK97BEKCRfb/ArUIwp9DUxAYtxV6ZoChErpVq1wkoGAUU
67dE/z0X5FyFMroTgVi/0oY7bBJ2CJihb7zZ/2OqpK2oLNt4mcfiYtp0luqNM75Og+xjzdUn9MoZ
IxGTzmBl7jM6KVKTrOSrl+MJ906g/bLXrswCNLUTSdh1D4PDQX4rU9sVHPXr6zHXJKAUqhDAGRxu
9oDdxPe2E8sXn9aADhPajIxD2pv/Q8FAd2GixeeL948XN07+8nuPLB/EweeTbVXwhGrTcaeEsbr9
kQYBC0Y8s2vVmyvWkFF83AA/ht4uHzm6ZjjPnai12sp18WJ6pO71HjEDbt2dZ1NCzlY+j4kl/htv
YGcDQFbuOMfvraNkv2sp7C9+AoDL8smIZ3t39rSfY9sIH4BDpH1jC/T0qnYkAjJv1kXwsYm2gQy/
4W+5y7CCN9Alx7LiQpdaBwulKiRtO4mUzBi26fRuF+FGPDAJF+E/fFu06yn5N8TRc6wIOKB5eS1D
hs+aDvUFTBCNJoy8sDBHPCbnBVSlxsLRnVto9CvvbTtBlqh3TOQn3pjN3xMnb9dsLnvd5VrDjQ58
edsc5lHAk5457g3IrC7i/wrnE7Ncuow3dlXirjnVRGG8W9ikjRap65dFgxPTLkeW0fvgJR1Hns6j
M8icjimmT5/zwW+IKptpoG4hvgETY/D7H52MyllKJw6OGoUJ9v/Szpf9cjwxEB3p+cb8Dlg1TIwh
DGHJ7aOjeaD/Vc2KBUMljvQXsSgUugDgWsuzlaBI0I4vGADdrm8e4dNr2QPw9cIB3Y35YkrAOCY7
bJRH/RwpdNkbTiK6Y/EJDb0Y01QFNphwQ8IPvty8qsegWWATXaKe8lnVI107EEHoSoUxAIN/9V6l
FM8lYl/Zr/4VbrRA4+cDKaUuxTEe19p7RkvEXACvk00HDm+7l/ASaQg5VJrwslzTJb+sgKpTVeMm
VAEJVsDI7wll+Cn5qZPjfLUbXmqhQYccwyz2QZr7cNDTRPuGMMWc9cKfCOPzSCffm2DmyouGCGh+
+elgT9cpv/xUjEKY6hotKEykGex120xRNTLfJfVtePrYLhxmAIFFhhaj2Wll+H+yDPxl2cxUx5oE
0BqJ/det3jsdpapF9meFMZ4SaM3PSWvnwWKpV4PSHRBJKxleklLdfD3SqYwBiK4l0HStiwPVTn3z
8EkRUC/m2gWyaMcmYp7CFpaKe78DxEj8Ba3Glaah/KAUqtTnEzZbhAQEjuq/smwZibpYI11ytMDS
wtqEuM4izRfHSEwkSgqHv8YPRdZwVKlGZwKZl4L1szZG6wQMBx6JhJDNww4gpwdABOgVIJgrb+cS
hCq1vqyOOWM/fEcMfWUp7vHapGt3198RnjpXmFcSKyAaJi5mQx7KK3VVXVl9v6eylliISYKvOlq1
hDDdXgNjYPcIL/e1yYwaR3/k3aBi+AeDOGIGPTgqC8EKNWn8ehmG+PWQSeb5Thd49z8wmKbGTSqV
86TImVvKS/bGEMbuP2KNsj58XeTBeAART52ePyshE8xDPJu9Rgo5eXzo1gEDQ0kj8sh2zl3dgAzo
k611eKN2igbm3Ofrd1EkVxfluIEBXw1vX8QK7BPco7+GFTJgWxx3sdzbtSgqdJVZvFPUY5kjWz37
fy/7Jc7lUiutg5qYQOERO5kO9q0yusPFBMqIzJLJcttMJRWAO2oV4l461j9q0k8PsC3cwhBpoT1f
+Xbe8MmrzFxQc7ZAqLp3j5dZ+GY5j+KeWDsQWO1PUeNQpB99mIjXehcdY3IqJznlJI7qxYzAhaHW
466eavMHE+q/86UEURKi3EkUEydgKRmXGEMDJKMQtCLtCBhryoTE/5rTsL8NCpqbn3sZ8Y6Sj4m0
5JNEsq/ORbw+enD4TKwTzIsjkxFLi99QcxPFEnuOqff1g7YFvM13qZcfU9QjVDFvn9FaJuX9X46m
3unGM5pobPaiinXHsR964t/4pv37LSDoOf+YPvRDB8hLfo/DUXvvlCkqRSBwnTr1JDQMUZitGGla
IfxLnzH51T7tnaP2D44QFMyL8xmfuCh9NRXShkLP5hQV8Wl+dNfRuDeLVCU8rH/JDt6boYpfCtvk
jUto7sdTTJuOIGpp/5GtmE1Hlid+EfKkqBeaTsDdNA9XZ4X43BTs2Fh+Djx9/bytBqeAUk61yRwV
yCbZ0KFf44N2ylBcmBRvvtdbAmquNgisDScBcHcHY6pG0KkTwuqKahh/Rqn8yzUpNzMkbWFTV5b5
XXViohZ5/dnZhJ3EZskcoJP4FelTvAcjHNGtnrlJwrdclO3xA8vFnMM1ubTDITgLc+7dZhrquLxC
s0NqbJ74sTwLmDjLhPGF4r7X7TPzFw7QUbicDNT23voXhUosm3lcfVPD6Wj+tXp4BIQnlH1Wnnn5
sKdXCzuwwlrUHHafv9FmLFg+zNOnSMuxJnJqz1+i7TvZMXYPFXHAzf+TMMOTGYgorSefLyTxvubL
kDrqBxfEs3SCjCvocHbtSLIYN03c1GpnFWU2MBVAN7BPSLypIRiCLstUE8h+ZBs1tEdCzse2QTv9
5ZP4G+EcSeVAsYugNPoMvEAuo1NH/qWIEGkdN9Opk3CWh8WD5k9HdhwVudRUtTeBB+YS1r7oZRpb
mnZG+1Q5ZeydK1I+xdNyeFk1zm7AgC8ZqNF4FYqRTyXZXxEfiF1xmlUs5LohxVkx+S/90EHn23Uo
QVKedcL2UgeFrEjz4MpPH7RpEW24mhNprjB3Rceo+VSrMbCSVR5KOjMaCG4imxNMH4Yl4uRYyigG
dDeylvgVvXNS+hLGR7MA/Olc8qZcKkY3XqsPjauxPlUajVcBSCM+yyEtsPxqR801pMekJ2KeoUbU
sMQcSs9angQiURtolxh/sGpO450QwsEqit/hWdgzpRkmhQQZ395FzKTSidWoGmAIqY97LBkA1PQv
HeIWi214BNGgffdmu87YOlEwI8uLPCWzyLtpfFQG7N6vPK/9mwnPtIg+fdFkFZ3gDt3b2Yt2kjHF
mROngRd4SMmRsn8aEn836ECNP7W9U11WSc6n1j/wl3M3TreZuh6KFdkBjf/COtv/q3PV3HCCPpKC
a/m7YthqNl0h1RPHmtRpkAP7KrRRd0httHCWyMVdW/AIsb5Dwp78jocImUcYeTwUoMvqzdX+L4YZ
p6EjL2YzXOqsjGDDaJp04aLcX8kL0+u4rA096E8JVkmj+vxHVYGL+bLoIttEiFC2tUKiyYXzOFYc
0s41mZc1iOSRGcErjQlQbLe0wmoPYLMEO2oJVnoZ9Pj7n7OJS3nT3HGVnCD0LH7SrY2aBRS70NBR
P3pnzbcoZJ9ruX2J4k0vpIisUhsize+Xy5WxgRK1fVZPPLr0pxdrJpHR52w5eSQ3GU+jDHVMZN94
K/3Eb6aXA7ntshdPhern1pf0KULAY6gapwiNFSitnQ145gP9dguvfPBWh9IcwqxT40iZ3MZXfGBQ
Hx4S51dwSB6ca/37Hm6AhL3ty5SGur4Ks4P1yXmkSqKCDTPuboa31yE6hik1frGt/khiw4hbZ6fh
svZjSLB8VKcB4kEoOepECsNxDV7CQivRZMZeKgauNTb5y7L+iC2tYu8V/uEWQrgAS6opSJjKPwna
unRiTdVvYbEDMtfEwgg2hAorcucBCtYc+sNXnc8+S+HNf4FZGhtcjsnDu/nDJ954Y/SmQLu+Ir3B
DgszHImorYCL16SjofFckIa59fj0TlFTfaVnIXrkXLujU8fizzKL1EnZtCrpRtgvDGkLKPH1wq9R
Qy9SWN5U6M/AE1JAuaA4EG5hcXI6NieXTPG2pY26VCQG5VcYtuuRMQVgmcPPyXBoFH0smXbK/LD0
J2Norx3IBa1TVR09lxs3vdX/Sp/yTlG/5n4LEymOuDbSrXw3RR94mUNFzOzO7M64tc5d0Pu+xaHC
ivf+AZTxM0d/TFO6Tz0lUBv8W0sK0KkdEi1ElJE74UYR8p7C3OuQDp1+gagafmb2aszdbR7HgGEY
G5EeWQX0uq/z1vXcGT+NAWDYxrNraLIgJSZ0kps1QlX9vToo4u25rs2XJXKCN39Oz0jSuUlmyeo2
qrBRf1Xi+kxF9CPk/0IetkPMG/CjvAKnrDXABtWpVQ2oVqPcBdD8FJxCMSRAXflapY1VajnNKKA6
1FC0vDgKvfMe+CHI0Log1VQcciGhMivkCoU+1RzQWJ3xRVgBgdI3wy9DY1hlnvu7z+dG7q+avPF8
cYL/t5p9XKh/PdKP2EKa/10SPGatbPh/bv+iGuiGeQhuwnknUR4HndOc/5o/Oh/1CUK75vcwO4Jb
eYk1soywM4dhbZHAzV08vG5vbFxSeBt0vmhIyRbwxD/OE8cK+p6lWmCl//55i5hryy6HSMbz0lV2
BUdUjRPvjQ2q5bpbp1LH5sVIOPUf8mZ8OvwwRKQhqmkJowrnXT9mRYit2zu4hI5hA+RMEWZvM4HG
cTqIVUG4WwFUmHAw03eRTUYTrEkr0xCU2j6FVCZPGS1PwP/8oAc1TViNOr82G4KliUAv++exQ2Xw
8LpvRIIt90yTSoYsnAkXwFWbWSSEYv5vILTZZ4hWA3PoD97xY4hIhgU4fB31YTLm/41KTZhKzHS1
oIAoOz6SG9Uklv1YBunfEGwi7nx38XAvKzGm3ezA7uLU+3v8ERmMUQCwLxedkODXxgs3pK3YU6za
sCsRKIzquGDOhUI7Bt6Ija1FUj9aLQmRk4BSv+FvVGGLMshZE8PGJ+dwJ5BH4J10IkGisGXZs67V
FbO9KX9Kz97onodWpf71xpSry33nK24sao326uZmtj4H7rXa/0MKXVUxsBKn0p4nT30cOQXam4w0
lKVpynguNM/HR0oHeiA3igbdUQ+59GFu5grbEES+B0dV9l1WCX8p0oS3hBGvfftyB7tOr99CEo92
7oNajQ4NZGMOij6NcwSfN+2NtBXFxDMIa44IO6UGqNgJTsDsQFXKeVDqb6b2ETK8efOxpP1fRqYO
BYFCzx+5/d1jsvOQRzt59Ra0fJbYN7QCUrQKXEH5BRj2xEG4lVi6qDcc00FAIiU3Tij0M+mpOq8a
HF2Vbs8sU1oMJUHKw4Lh1t6okUYZ/eeTAsZOiHnaT1Q5qm9kWiVxfIRt+k7QufYijqZLVNuOX1Xb
uD67dInURVe7PfcheUz37ByWMhDYCtAKzC3FhIXEcDsXtkhR2g8G4du+jjKi3CmGVQYN88nne9/R
ki0O/Of8h4fxFtjIx8yH+8oCIKcy+AU4RhscHZzI9XhFFchr/yrYMZig9xxdZye4NFOT9ra87bam
c+Tmqjz9XaTJaK432n9q0ShnorYTgmHCBkFBpEjS+92f1XygUkna546Q6SQYQDH02dp0X7AjSJll
g3Z37bE+n8I+kixBf6cRis+MZ2YLJAlpohASpEhxpFbjbbQvi8AEzpRcFiL8dBKT8g8eqRyRoGXN
mB1mWkmxl0inYUfGqC48mEUQi6H5U7War8uv7ND5zsviFfhaI3wRd5LYW/P2Z3SOZ4ND07wQBPf2
qTyaeBy8ykaxa0yBx5e+91STU7KZEeAlKuhlM9cyIAryuhKdBATtnuqSe7HS+sQhNX8gchNiErzh
4aLYrY48DGjxSvgTqgZ3cNkXofqkTOXp8OqM0f7r5E2ABkzJNRkXOGpqUT3oGCX+RTvgBxIRSr31
0y3rEIRzweMJjr0pHpnSXIuZCyEdY6e1tsszPv/EXBaQIYSczFgP2QE2f+NX/P7h1UjWzLs8hdp1
RMqH1u9k0neMRtkHVtfbAGZMQVYFMqIwXz9uP842gPGFLc/mR6+R5+qUa5j5zySeZyzA0sRjivx9
QsPzI1PJWtFitmhzzGQDgU50TfgZlGapFpoC9YLxFA2I8MCRJxIUVvkhTRGuPChRiiALxB62EtcO
UrqZfrpx147VzXh6Cvq3RyLh567xMRC/li/gVY5rvFVL7RPO33+YjifDrkAWhnCARAKlTBGjr0ux
rcN5iFhI/OIxUqf0qVTaHbEpaJYjc8CxFDpiXW/JqZ1yLGFwfQ6CTyYyqMj+jVCrcQZq4uoeZt9c
Nd4ojF23k/k9rJJzUzhYWU6tM8SuPCbYL9m9uFhm8piszGpngiGk2BNVq99Onl0Ua3WSfKnhld2a
/+7A0J9KGdHeLYImxld0XBPJMBAmiQ/08ZglNk6ju1ZSrNuOA0Y3IusG+N+DmAY35qwV2DwDoKQl
IkiOG/2emPHLBfSqMjCLNQkVh0+9IOQNgPY+Fx2Cs/uRuOr0G5v0s1V7cLvpoUKDMDW0RjACsvop
TSq7Y6tt3VuOoHQLmPxDZL2Cye0ssZ7tAfNCmoDrTttAod2hx0rC+LLG8klUxnwS3ufQ3zPfgv5x
bWERSQsXObp0pAOg8ds1GxLzF2K8c+eB8pNf3NOOagLovIbywTTS6yAmFsxD/ddfFdFrkdXumyRE
1R8cGXQmq/EFp8rO0G1Tjsbbd5ahAdztdyIR5/cTg55gStiRjJRT8VlprdxNUTDlai+1200P5jGg
dlREyi6T9fPEaKNE/f7cIfOpUt18WxenVq4dyZcbXul8twSC8QQ8+dLpgOdrut+a3QLxJWQrwl/O
bpN+Yk0I8MzZ2cGvLAOlCtbwwkTqjA2T7szq5x1vI1aVb1YIqhiEUGI/J+yQ4UgI2RsL3CygHFFJ
A/c/y7XHh/cwH0Kv2/CJkr9tcbUk7CLUBaWGDPVRKxnNfCyTla+N0kqdoLGRJuRSTStW5m4PemoT
lioZvPeTSuI/Vlf7873UrSsxXYtwDtzwYKzIbAFz3dWDu1AWEMzBA1Z5ZZ0snRrGckp9Q3DBY7I5
Om6SyvO4sI/t+aZCospj7h0hNJdZSNn9zGSFfOGikZuKp+Tgs3VEwhDcUvvtZfR0l8kHPH8ISpoo
AbfQNIe70pHsgIvRAI10ZEVjoFPr+rTxsI6RAcCbL9LFS49+RRc4wOWEZntT9cOk3AaoaMJRK4G2
KFtO4Pk+2EWJCyynDPQOvbGJY78fqGep0zBNpCE+fPmpiWoEUKAn5yd7r0i7xcGkyn1/9XXK121M
JvIRDqDpOwuoK0Tr3EeNkhgtmz4Z/mTCnxt+7pqmkWeocsbN0ZVrCSDSvGz2mdOx2Qu4HyTG64Tx
5yx/Z9ndlp2C802ira3/sJXCZ2jJdKKufamBu8R7fz2Ohi4bywUezM/ra00U5PFA2lvL+jpqeThy
1NC01mJXqavpr6oE2GJBDeGtlKxoirzARDUAzi18uMr45aHhqHHI0KjJUVN4aooBSJW9gHW/zCmP
cn7X+CMsCPjvodGK+Tjo7YlILj2NnhnmDwLIn5f/l9jiUU5EBBGX8wpZVgzDfOiqW1WJD/1U+c+Q
lJ85NTlKvPWbwqUjnaNn8sjfLfzH/5hN9gnMHzgQRK+FN6rGVMCRjpyOKpKwK7cWEv2neYNaz2ww
YuAphrHKx4Yo4PM6lqIoZmpWTLQfKjOBvZ7DwaXwwGWzOH7mvKmgBfxvMNpLeIDaOMc2kwvK7zAC
gR5nWQfO7ovQMC1Tu7CnzLHXuPiYNaYvQm8+qnnf+bibMJjBED9AjH8ebTkiFAhwfC2FQF3sBmWU
6moTLoRhfyqPgNDe2Rzd8/l6/WZFta+nBWdq4/0v7kQnRKBKWB+SO+a0mR4HB2hcbn9Cl7prPcrv
rCLNLaeLuaIgS/1GooXYBPSHQz6Xf9P/ovFdSlJmts+rd0PvHVZeUh84eHSD78b9g/WOMxJBJEuf
IR6ZbYOclO6HvUhFkYjooEjOnqVoLDxM330xg9Q6iktIRggjMkLFs7OFiOGYkz9r1nNp9iYkL/hs
6tonRkctJ0OLusm1JjvGr7NrmMhhfSW8JVUYmvSVNQ01KsXox0NO7o/sgFiv/YtyE4yCpFKjQtaD
ZymwWGEMSavy3LgEyFu+7Zo3QUIbbMEro7vDwP4DY63rX2yhDq5cUi/rV+Tog7NXpwq8HCYchr8k
bC2MY5b70s5W2tuL72zaSAPtXw1nf79yPd8jepaqcokMBVWWTjsML2Mb1C/cEJ2PLfp2HCjZrXZX
qLCASoQlAzfgOq4annDGQgxh2jjGowIai7BGhj3YpR7lNKFAMBVc1oqB5N64dJviIN/6WoBJ+0Yf
CHKmUPIUcAW63AjdB2gv+ZfVftO1Z3+Bwbwh4O5wKf1iZElgG0i3Q2HbZvPtyWuG9myQIWLUOtXS
5c0VTfI9FnjbfCoYeqB+Yj1EY1D6rgSm0AlzvNoNamWGXC3jKFRJbmQ2bgPXAD6Zydx/v7beexaz
jNgofefrQB3kcJVmoLxUkKLCXKyWKI8J40u/H9nki+1/brg1DR4uyFOwB92/BiW+fY1LtYPryRQZ
qWVr/FSzs2J8hUYG7LoOD7mT8H+7kZCo+0zq+jLX6aD6Q9NshljBML9hP7ltyra98X9rWWtNKLhD
2hv1JEAVP7hUCuGEU1aFSN0hnMKi4kMXy77iosWwvmK6PF7bgaaH7enE/iXkaQoW1t2zhknndbjb
CgHgkzj4/sDdjElDWnpS2fU617D1gkEZXokJV28kTt55H4Edubxuov5DnEgo4Qo8n08pjBAvFspE
qBaayW/XkKvg5k63ERY8ZN89dIy831s68Ipx+mmdibBSud6ulFm1f58c95nOl/s3cDIYnfOH3E7s
/P4sKr2tnCmgTTQEdlJ7YAOjiu9/7LcnhJVIxo63BwPVqhc+oBlEo+Dir0P1aPvCUuRfNK5h2x4S
Ev2VQdOcyudYd+1ctF/Dw+JThAMCKyKd1sIevYd0wY+kN9He/g9gHOmimJAYoPj5yj9NPdvCquRi
8jscErKAX33ihAZLv8H/TWf00A4YIzYLSTEtus57DersSEH2zDvYoijIZr4OKMfjDS5M+lWzkNDN
BlaxcHQsG+Z3xF1m0/1TSZARl7+/59GYFbqUf4jFnSd7JeTktPjiqy7crhre3/+w4TD5dHDCl46O
v2yK7Oyeja90d/MhWjriBVBAoGfGmrrcF9ihZXB/6yM5VsD9cSKelUc0MZ7eMNeSuuZ8+dGFZ/dM
BvAWmiGvoTWCFtGuZzSP/gcO/Ixi1PCLdgdRzcJ0LExEGfHuujPyask0R/UjWVvhzyjdH9Xs1/gT
/tREdWsuhK+BRymza/hUzsZMg4oUEOlRae94xtMBUYuvPxLdNoejGqcZ8HbzoqOI4TMxizCstxpl
2NRihTwGXLN2Z903swxlE32RvlU1E/SXXZRBlRCyhcZTgJWvRQS8Vdt2ALFT5T6jtvw+YuqzEW+p
Y62vVUZiGbL7OCiUTzjqmYGoHaLhenV5WGuYRZZ2Hpg3DMqDmt8abWZPiMZD13Q9T0RtqqtOhQm4
3dWFGrx1bR2T/dF8gFeQN7Mznp1d0Zf3JBKyTj6L7rpY8wMyWVlaT6JwGBjekGn7P3cb3swJW3aE
/ckHPVUvFmtt+OQ7L77+EyqSM+JUvaLM06wApINBKmQzhUbfOVj6LnLSHYoj+XCRuU42bYermzLx
kil2SSJYG9MzaXNuff32s3YHgLNJ3TC57YMxbDsl6ElluxDzjA9IOGYsZxRLoofmLeB/HhYWZWnV
Q2+Z/3ksaOz7jgWiBzE3tE02bU+yo38KdxUivn+RBCU+2uGNpHwYmd+MUKvTrYDtFzOcJfEFLTJt
TOgXIl2t1d2OyQC4VIE1USNtNzqCqx2HyX/7rmeeZ/FiCmiySqq2zUJeWsIW9eegHfjidMjiKr/m
fa0/xxzVNZc7sYY7O2UArjheOfYueGQdcDcUtlVmw52exPnCDJ5/BP8YLpwG4KO7FOoBPyV75D8I
NvEIeb5iUIrr411u/EZOD6nqQ015bJYViKzKmXQ027zMlzytMuktvWclE5qSaRdut+xEfkELFqJt
KM+g2GMv8LSgeyAbXAJfAqg0LxyxGUaF00miO2/NZnahV+QtgHhgfnXIJ1cb/zrc7ZbNpceEzFNL
MFnApWq9kyQ9H3OLh6BQOhf1qlDdhZ/bGUjYrg1AhPd5BKiuKbiEM2+3YKcLT1VgDZbHDz2RGXuE
dghOaGAySuKWbEaf6PqpuSthhZEyk6hP1er0qHp28b5KRZmdRpmPD0ENejTWBRile/onjv1t2bUs
JGmtEGjEc0nHJ2WErdcJWyEZ4PBZ39KzfkTxmv2FC5YSn3P4E58Gltaqv3kF8oE4GijbSsO8Jh8F
PttMw6f/3xYxcSiqYCHAb0yMTDNkRlDNDDlMXMNoyrB8vSFKPDPVybvl69cHUhKTiebxhkCIrqbG
RfGqhPn27eRmpWO+fgHWu8wh97aW7Zjq2iVtXRVCdOvIdUBBAvr/ErPvT5NvnBjEpHo155TS9hjI
GSLOlqPM8XFQEYXVWzVwUZcjOI7/nwmTe/mP+IRqphkhwgnNWMuAW70u7OaSzy+gohEKSOHUpUzb
tekILrX+SXAx77lkF1QXZi8WS5orHIak5OO8QJqyt69PW3eN4meiYxZ/rZc6uQINA0FkG2mcdk+L
XVgzvYPW0SQ9KYtjj4fhcM4/YIRKcikgzgkiXq1mD6QXrUrSvHUQoGDpBX5P3B8d42DyC3KyqzPd
Wt/c7KxQsCRLuCYeK4zo/exquSiOdFebdqVCxrW7c2+nYQswlqRE3vTztJLBocSlt8hD5QcCxGml
YB0D6oQhyx+ZjPM0QgZZA8pMOJS251hmyZ0Faue9G0obdVwc6OdqXH0Xuq/zMGUDxLDT6B6ccxlZ
izZ92VJPff6X7DiAIoH++0r5uGXR4/7L/eBYT2sQ3j+U6eOO87NpytHrpo9zT6ozz1yDGZzZO2Be
md3AZ0QzZFofFdWxlQY6CZh2sPzSJNTtC28g6xgwB/i6FPY0EhvQYv5mMfYotIuIyJp1kO8PpfCR
ARLDtmxuRinIovjY9oA30dHN5ZXoPNjL8HsH2J56LqDA3JSNwkUAm/6Qx1dG4qu9Zr2IQ5sSDCRk
koDoRZREBwg9y3pUHPBJoLM5zP6x90oAvNptVfP41yTA5UAEl+ZFblHhtWVWar+TpUu2E4PVel/D
6Z0F1uKFrnB9YTBt0XPsSUiqw8q4Jth/obW1m46Vq1GK6UNG4u3XVv7GBYGd3TefIbo/TpFVI8bc
Fjod2ZWPOJ0yDWuwV1AtsCCgGKze5ZAGMLMH7CVdkFQXnAtAGic+IE+W6+Mg1wP2PZVDQYtOmMZM
yIUgRganlZ6AzbI2z2L2KMSsZonv9WPmy8g4ReO/HP9dlz4j8dPDbHsbiAGifV/b/ihcPUAIoXJP
EXUBWHt/FngbQ0hyptH5VWoQLYJqBqqRXlrW/5pW4n13Jbp/DIG+82zbCO+lIhuXr7BDzD4Oh/7X
0zI5JjWt7J8dOUzGg4mT7s4WM+blMK92Rh/enZE6MV5n2c53Bnm/ZkK77FWjr8VDdeaccoYdZ9kQ
sz0MnOstPxID+Is2N71qRhAE2ZaIVMlboJgnmnG7wQRC2bnj1DDL8+lstbSbmLkNIraD/rSmUrDv
Lk059UHHMLUonOW0XnRPDnHIo4qDiFxpxTvWpuebNm4nBcx1dLMUHZ0CqOy7ANP2/JsQ2U1YQtW7
CRzys3XJsUkIXaZgTl8RyjpR66eXceZ1GcmrF+xb8xHngkbsbl/cPTMaZQCCtZRpHNXpC7hAED1N
/bPaA7MrBCuBvjD6/EGY6XEczniugcDDX72es7Sb4/5FYfClr5/4F1mTgkRWJV86F2DAB0ywNQf7
hxXkXKzC0k0UZBsRFeK5I1VvsGcc6eIAuLGpB1JI6nLRLBXamS/biQ6LEcB3rON2/Tm3jMNpxJFn
8597d0PE34teOHQwNNvvLCN3ICyv5GtetW+ugBECLxcBltj3sPLLLi5KmcsKYN5mL6cpWVGC1vDF
tYRM6xay4Es5PjAYN7mnCt5ioNu7umTLc+zuzrXH6OH/BuT3LcnzcyDunO0dHPpb4Jj/NfP3v8OM
2Al6E4MdbdCzWWCGh9b3stwml34TYsqGIWafV5Uo3Pd7qYCkUHbH0YLkvFlhPMuCwSEmwQPghEgQ
kOK4v9/zbRtadmjBXMzYiusOeOT2jpjiaW3kOEjT8iU42wkBo5DzYzwb4yDhZV1UjK8iNwasqnoT
ovWOm7JLOOygc0i+4nFifNuXugIp0i0lU62E6SNXiqc1NNg6DNbruRAJvUEoa7KUVOrllGk5BcQ0
5SrqkWk7QJM2ZrmYjWa0V4QWfm5mqup6DVmq9COAfN5BLiPIXYeukAojFQewfSoczXgg/dtYa6fU
gGLX9w4Q4OshqVtzlr/XOzUpDSmaVw23ModFz6bI3efi4irunk5drGBrwFKIl3zK9I43MrUywdQQ
zXLc+UaY9s5Xdvgbbs7Kvmjtlluy40pz6IRigSo0P7qDfCN+P/Yd88ZruyQ7WlSwtOyd00VJOktH
dPS+Cmm//+ABvLfmu5jdBd8n2vgYc+LgFaC1WL+MadoEPa0DcQHzpwZkxARGnecDu86EtDjbupy+
Ojtd/pkgtg/83e422MT01OfSX8j06dgaDRZPKoxrvAilsB0hn+dpOMMcWNNQIhohwcOpv2KOkfKj
Gsby9ahPPuLAytpMFfiVYWx3lmZ/EXM4c5dRgmZKSSvPGSZeXEjy6/SWMi8xLFVt/0rhqaugqA08
441rUmOzUXBQs3sw7GkVlXG1e+5hUoBEfZKDqRkLE7HIzafoNPKAIEyXc4X2ImErx3C0+4o5YEIC
wQycuL+YzVoHaFNcM5FGoVwTzaWW6miJ+OD5K2lpq+sBFGz2YnwZV4w7B7d7G/AbtfQsllEdWzfo
nqB233oMql+UFkuZtEAM/qsR0h7FCY9psKkQcacnaqDH2h99CJ5KG+ZO/f0FxbxSJf6Zbu70l0Um
2s/AWWT/t1bdsuqo+hbOoXjwm9h48XGaahwIWsOrnpCegdALbENbI6WFbzut+D+pmq3SjCWX6DPc
qm5m0eT8lkel05wjYCMJx0bwPBHRXe4e8egwJ2SkybiQHz//UvQYl+fo9NHoyWtQYZy3697IJ1cu
XNUlcxmGIwAGNgcToigSA5NmyJAgiIjGA7q+XSK2lIgP2rH+HKkK3xV/TQeRYpLg2icEALD+tYQ+
SeOM4OnbMymCdBkTVpQieWgb+aq77sZv/yEz236fV50yllU8bIvrGUtta1Zoit94a6yPKQ3nn5s5
LwBrwplFwZmc0Op8DNR4Fz6CjcG9Bj0nFFmzhqBiq/qgO2gKZfsv4dQ26HKSRB7G96/kgFS1hqYf
yOrYJUi7NgHdCbzSLuBpwsk4/k/Bgp1ahDy2CxxGz1X2jwE8lT/W1yCbhDKKD7Dcq9AhMrlvPBuU
CFbdCbmWDoo4JmZ8XV6lEbBLSbjFutccC05jWXdOMq5LPNVkkBfNx/rBhBQeXALHgkIgVs7iYmSc
5SlvNtzi/dlE/i7Of+h9Dj2Si1ZDSxIVcSi4sZBU7ADb9ctXCxPsFZqYwu5f28fNWCdQ5H2BEg0b
JRLc8dClsDievVwFyYjv0J+rzLLBPKXUmWz6yMPxKFSgOIiB1TBy/dG+tXuhqk4hYjt6wFBn8W2B
uLD7BL2v7bofNI6P3oPTRQhq4RXL0Ds+RMH/RrT9JM8Krt8qP4ybL1G8rVGtQdQSnfdPFyQs7vGX
YJuIMf3hoBDB+1PPyylzONrGILtsduxpcz6rvTLok3ayg4XLBh+2o/k5wz2ElAk58sjjmVr223+d
XhCVrNIo9bwg/38mQy4uYz7/xHWPOc12juuz48WB6cBPzWkZmCojkiBuebMEp3uvqEoo3iXCHcgg
bnLr1rdHfbkpdMOHuFEubuPR/qIH6hJM8gviLpXX7O5sjqIKSw/csc77DWF3/Mz3nhEsYt1LgOzZ
XQTRzm/RT7xP+WzxKxNht7R5IRAVuePeLZVTPqHfzeoOt2d5nJ5qQuXj8TZlOUtkSkyWpOXnSBCl
7XTgxN+zfN9YUP5R33+09QBNEXfqvFslSDYAwRQNSet1E/qrK4s2pzDQxu0TllGrPTh80S4sGUFm
1jB4Qoe1uneF3RIbhoxnFkQSbXRpiyeFoR2G3WpO/rQOnLsoEfVWjA4AdKkxQZ7J9vFuXnrczjxw
FCh3mMTxOG3zyEMbkgXy36vU9mjA7bi4VKDt7pnceWUnpYiuV63Ka8bFO1Kds5PZ+JVb+hLFC94P
XdOYPvCO/Nwt1enXJor7irw8Eai3H489iMidAHwqRsSQbKHGufFKlFUp13UH1Uy6r5WOI2FSmkCG
iP2lmaRYGDn/7kt7DMaNo07w+JUyDSc+POW/vLRgRz4y8dKSDsCnfCas93dXr22dvjlNHGhpXfp1
2gZMDfFmEHXtOK/AtsmJTwMozJMwpljs8gOlkrBJZg1SwYO1r1Iamb03t5kEFQTaiTIazDVo+Q5L
17MJp8ojfIpdRHHS0QyyoPiXrnkj2O452JLG5AAyMy9jXz/6CkuGhHgwE8Hc8/woWhQD1tr7KNZs
yxQJ7eyHHSFlONoD+PXbjytLf7rZD1cGaSnXk7h9sQfqo18qNlpCIfCH+2pXatjU9UlkaCZKjk21
Tpo1y215rVsXw1J1CxahU5MWyxNalhIOtjpD4H+MtFZMUmewUpEo8e152LbDNJArB8crAnhPhCAQ
BjJ93f2lhEKbulAmtOAc/GiKzUn2Iqf+T6AakddVsZgVl061PSufXSHwHI+dryu7iqbTA9211Xfg
exiCiAG7jIZ0r3dlDIwUljFhtf+BgOIv+QfMlFCeB9zJTtQGyKG7qNn4zffSK9AZ16EcXy9JVQlC
u1d1dnpUtjQRQgY7jFxrjYB0EhcbrGlZgEEABw/EPD82thYDFTvqbMMGr+J/q+wx/HrZxyppEmZa
bGMdGXepmIqiqFeotLjg65QQutjtta0gTAByR0LwqlKgJiYeXQBJOW896PU8ox+eZfambs9yqvGy
iHRl6EeT/cguKhOKfA7OQ/Hd3n8+nuQzH3Xi9RP5CHnlH2xr4IGtPXrWlZzD98gA3lfe0J1CXXON
lMOMiJqBhh9h2pVijVi5t3xA27AqLwLf0hybH+8hRe96Y7MOOofzJybm2RRvaUk/cVy0lnx2kG5J
QAFlkpPnAorB9bra44giC19S+VIBDQ/1GdFErre1SrZj435DzftsXlK3dftldF+vi0/dfeZgtPVo
651qb/IV2DQ9YrHx2cUMPokASvhzVS3p0vYHn9x3U3RTlZVsUxKq//ovz7qxu5xMrke30QuZ1iA9
O54n5hAUdzDuHII2aRIUWLJkmSoB5f2T1WgBn29VtbxrxPV5csTeo5zkT/NlrhUumY3UnoKTeBI6
olZmojeb4cpTSpSM05nqqlKCtSN/wbI4A2lz3QxfMXgGv47F1NPiUg8NmFcoRUWlnbSlz7kHqUDQ
2h077UNps9E0yGzwW8w6cfZwfsPNvboLWjkmqu/MRRBBaDdDIMbR4/SlIH/uNjS0fcEp6AboYiOV
D+BThCeox0nirnYLP3L9NoxtLfMKeGY31aBOJGRUK6LGscINtltakep8nWA6S52Rl72GI7fpdb5O
FrA8qdfYMY3wTsBWLugMjUtcnpigbx5ju6GgTicMsLXOy2kTvQMi1cKArSE8uXVSpwL9xv7pKEpg
MdyAlW1GLoXgovPjOlMUr4fz+b72yXMAqrEb2+bR2+FtXnTXdi762qKgeSJKqTJt3M54um6BxgCG
mmSrzZBvApH1N0oiHNrWahndUphGBsb5ScRBXP88EtGmZur2NHsH8yuVCZLiYoIeO2KzaFPr2C6a
MTlc3aotAH/sDsXn/4fTZFkB9lNkl1OO11YceYSvvj4kPgmQciCssWmqDFOvkcXWjN2qead4UTZG
ZFBpH0TAh+zgTYpCUXovUfmfLtEoIK7Jy7GbU7VpbYnniTqiRsDYMsjNVWJiBqedO5YLjBKgB+Rb
p28QOYKWXHqeBjYhANUPZR6m9prd4yFZrImA/zIFVN8cq6z3gGS8ItpKJTSU3rR3UJSpz7oMPwMx
7ZrGtwtimgZnQqcYBLPXZwOv0nnDlCGDre9yykzvEn4fpiEYhtSqikgH/eoLq7weCZ4zbfhz5qPy
4apgJIUhBuA1eRSA9sUHE6g6lPbTAX+vttaT2tzb6z/KFOyCV5s+fnZXcIAU1XR+MOrBLOMx03oy
xnrkcFw2wVkz5rUqgEJpWo2oCvzLP4lVuDWFGyjeMxZrjjUFp2BXkjfPdnww6pweaqVQjqCGmuG5
WB+307C5tJT9yJlga78uBeKx/VyUSGbxN3nd119H25p6Y+420up/u+f9yCNntBXC2DNbgbeWjVgD
9nRAVWXRSpTl9BaoziPe/MPwbJNydqDOz2+NbCEp5hyLxvSbhQtO/NOwOHzKgWAU6bZSWFZWBRkx
xrZgutYeweUgUHqZxlbTcNIoeG0UpzFUL89uExDUUIoVpJqBsalaetnkibU6qA2qF+lpxPzaS9DZ
gL+sFUX9OlHyjQotgMGJyKXJRN4Pr+fRXlTlVrKrmOTzxyV0rG+m8+mYmhiXa3KIn50D7R2Zg7w2
3JUpN9frl+hYHAkpKMJieEW9bzxmP4BoXbX+aWRc9I4XjMOtUPNQZRQRqv7dlqN5xA8oYimqURSC
WsBsNY/q3Cm1aKx/kmV2o3PabszOGSr8F91bchkwhSlR2iFSSPfVw967yOEUe0Cq5K4LxOccO5SV
dKPPPVdR3i8Fdq+HRe6RpJsBAq32+rzx+ikgiEZxID1Rg+8IpK9cFe51OFKRzVqu8ott+H/p/ySo
0JJMjF/wa8hSgRxz5g2rzYWwnb2NGqu+RFZfv9QSVAdCcMCLor+xgEkcJgaP3r2hYQZrR1HU6v6k
sk1kMoIkF/KJRGPIHgEic6JgIkYmUODIrXrlro5a8L3gwqFT2fUQZRLZLfl70ccx2+ddJeCZBTD3
XBdSX+hyeKccEeW/8oHYOYBMy1yPxfEMgwwNrgwYnoocugNwUztasn3jU4PHa7nf9PO9fkq5SwkC
vLapUDOA7W77J/1hxwY1mhR+XgfRwf5BHl0f+bVClfWaL4NQ3rlvw+RI8inOZ06ocVPBexv0Ym1m
vLy28XC2nAB3UQhatG4SmmYeMIm1FNTztzLTs2jiqWUez0Vpu704luQpxQCieX1lMC7WGZn3IPP/
b+fFLR9w7lgOZnAs33wTlE0cH3oWML7W0rXILONcsAqvcMMimX78e0bf3MauOGJp8XJ+qxjnsaj4
GAiFYUzLfAKYk1T8DG6ZYm8pStSgA6oDfC83lRgpuNrpzssxYRMXl/BeBOcdmgLwbYDQD9einm5g
/DXx/dqIXbO9e39VU/uk5KI1FQA6jKn5IRJrNuFGTdHqUF0pr4m/HtVL+aab5df7mz93DGg3F2k0
a7uc335oG0nXSe9TDcHAhs/MISmBpJkwRzmx4+1py8QhB8CLTWElNcwLWN/bxQ3ddJbKWucqbzWA
N/1RQsIf8R6sTAB5DKzMDYH2uQHoFgmMbUodRvhcUfGPNZi90KQ/Yu6iMIvYSiXgwoQz8RBW/kDE
auZgqCkHd7FNnjEuAP3rpJndQ4vVvb9I4Xe5QOnj9l8Z+lWIJnAmAJJMbF9h2y3Ut8c6vUIjyaWP
G//VSLO0jhigcPXoeUZwH+91R6JSxq8PIooGwD8DGpTo4mNASNfSLTh+kBYsTn2kjUcm0hsf73K+
CRDoBalcQXFmFlt2XTH8qRNl8cPPITXISykW7nHcA3muAXDuTXtyERN6UgDtOS9zwAg/1G0sR/pT
rdzQTHv+kpUqNqmvWfPsHcH5Zjn4jvYWNMuqdAWM7LAr+R/ElOfmfFUu90camjyxefjJJuZrPpZP
4ipEcPAy93z4fWNJRniiPWFvfEY7An7icwLSiykpyhu+jUiZpTNBJSt1wLkuUnq7SNE2TdyXpAb5
WC7I9kXtjqdiZi3gqAZH6p9e1aVAtqO5Op4KsavYD8s0ZkkyK4uekIa8UvRgxXhFI29NMcJXfPA6
0mMHtfCtMsFZm9tUpx9roMOdvlHMCJzkQjC28/3lTlOfVKXpkkqBQDMY28z5FJ5VXlIz1HaPbEQG
SDtYhkBfG5UpuuDnFv7ToZSKT6gA10qWs7jGxzhio4DBXMhBBGI0PIwIxYfTuEscaJ9lM9HvMEP6
ZbdZ89hRGUGtS9Is45bfWh1z5+kFdO/tKl//i+qtxtCeaYaNcui4mpQ5+91f/mHlve5FLL6Pie5E
cfHbbvDY/NGVTtSwmmwo6gsxjiYo88pGKAIneDwPNCgbpHAjSUQzXMOMxk9VYnrmPP+c2nxqDB39
7S2S+6ahmbf2gsdiJKxowzd1v9Ly4zS00GIyczl7vJx+hqDutNSRbYhOX0R31RgI9YoatqavQsk0
+z2n8wDliuuZ+JapGh9EgvbfAXpO9cbesr4iOpCWI4L4NjBaqSA7HUt3RoFJnUNlGFfElJF393M2
+4zv9yt3aFVI51a6OV7uCCOh67aZlYJhug5WD28DFqxVg05HddTublLbqdM4rtKsqye0OxYbZqQA
lxfnZMtVX6gm7gGvo5d9WBqYn0RdygFO94V89Gc4R4UC5lC2u+Bm5lBIdNr1+SjNHVGSq5Ijmcx6
cZ1qBXuHCxGu0EZZf7pO3b3WzuBKIBy2aeB9BrOGndoRtIgKv2xIVWh8MRNWIKKtj8+pElCh/9rF
NMNVJsShFpOQ0s/SljaYqzvO+TjZllY8pxRO5lJoXeZ79OzSJ8mfqMp77U2duAIxzkyid90u43cL
vXMsmhFKrG0XH1MKqs1AU47uIRBrqA1xg1TiS9//MWZTpgeqS9uLFWD9c5WUbt5xMkXbZnIldH0p
XM+2Z7uMTssHDZatqMRwnxqQLH4GpnHLnzLmUM6YrNSAFjfrTgwMOKa0CdN+QrfCRITja28afTKt
ncfAazZAoc5hupN/rGRd/1oipzsA8KQaTym9D6gg2p2WgaKNff972OUK4Oi4o1HIcjb0Ppyn2orz
6WCJrGI9oWydZX/CI++yx+2EvThEBisw4oUXZ1da55curf62QvHNkkX1NvSUZXCXzXyw+He4XnS0
yHHhZmZseF/29QXirbTRoRIG9cuNUBjlGNINqAJXIkDIR5RqjYs5acfpwTIUH8677qAsqBG90LPn
IV91GAXl18fuGZlhM4/y1Rkw0K6UaPdO+tekwL8nZ7QlZA8udkSfU2d3w1VXG4k5plqNOFdZMr63
ZNS9pq44NP7cnJcD11mRqWDu3J5Ya1C5GZArXZboLgzBO0N8ESIdX7bqZj7rTBunIYSNOIfyQatu
syGfVC6be7oWAXofjHksldP/aOo5buP9KhNV1obokFmf1OYBoms+wipbFlqDM3iwwCbWf1x8DQ6s
9iUnzbNVQTzyDYegDlGj+4PCAfQIGpVer+7nncWtmJlXq6PJ3ZU/6NlVgA9f7rtgeZB9JYwMBI1A
mpnyVoFEGtiCTLDx/LtW3jtZfyHqYQGrqfv03FgEZtuRs/9euSVB87SmWLbXyZLUYI69JAhr06S2
B4uOLUxpvzWuT8EIeXsYWtDBA+eP74is030UDV7FJHkhrHCjvGZFqwyq97RPFCOJuesxUAVP0N3g
pcy4I1NAxqFXh7VTbE3tiWvOyqwo3uY+G+3QI7GtkPDKyQtIE7sZEJXRc+FEsgaXdc0dLB4y2LK2
8cF5+7YLo1ZPdpenLfzBCaPahuRyAMk6XAu54R7d3JcnnzFdcHagGzyl6srIAeXWk8ci9rDqdJ7C
hmXY52CAt4HmJdWHn449zHdzqaarupUAmnZ7PXCamxenqEqpwNrLQ2PejwEjoJIHUmHD3jgObAjj
kvOoeGDAtgvuMZwrxN9QLKepBWAuzblCCVWJACI+u415fnO2T4bkURmneKwnOjmesDoHjEa6JcXM
lMahmXD4u0E8TAmhB0Zi+M7iYImZOIhbfTh+OSHCAclgu2D11nKzvv2NmuvYXgcOwZRou2CV4T1z
Q5x9gG1qP2vYSVbxrBV6Xa9WvMv3nTL0NnePfEWI15JSILeu7+rrdSpt2W3MmRMgy3KJkTNB5dNZ
HPbunWZt0Mx8S7QQArnxd5Q9aPt7UYqCU/2eAf7PvsMP9Zw/0awo1/o9o91oah5jj9FM6GUgyv4V
9rJpmLKxxkZg4/94zZlemuhKeA3dx+5yBYzYZvvF8hEw5ZdRwJ8Jxk2aTwKPq69F+LRQ3vy6u6dr
6L7vUzFaRO5VjCfXUYgHbkiv9Cc5C/8ijM66Y5weCYV34nB8RerzAzmM6M0W/87c1d3U/ZloI3oq
/IRfZbHYq7czQiIUXRgbwusnLK2Gh6hHgkplZke040iYxor4PH1t4+hBhEHnqypPfXso2rhscjgJ
f94bowSK0Tfd2r6+KwlTElxonpxphSx7H0fEwHXkuf9OXXwPIUM/pFa6pzG6DQy93b7OKygCW4A/
nF2HfEmu06oDQBmVb8XInR+9QIGdJmA2RFkSDNMKpBzeH9byyVNU7LxigJl7TvwhF4CX9oQF5d2j
fqJQuFxWmFNPnWewkghfAvWCmPuKA/62LGxDu/DQ9jZz4KwoUbG/Xhp8SkAjbLohu5qOx/C5q4yr
NSEMyLlRIM9cQBhCudgznlNT4YomNCLnm/tZ1jOOTQmCvzaPsPouuSlxj0C3dUc0vPsiBckV2bOE
8n8TXpFzYFBNzJEYy8HcCZZcfEYCjC9KjTQjR5LhpJHlrfA2Cm9Tsvlt446pO8B6bPGPQA/i7kMw
TaAUkjdWZlhRk2nSEMY8zN1LXQdK1Bdwnv47nlXKH9cb9srZNDnKdqpr+vtKoAj/rHRv4Eyxrq+u
+89vydaSADxVa33OLf8dnV2kGaepDaKLp+YHB++XVToe57Ta8aXYVNRGe58ge40ce3voy5kRJWMV
zCzBGvOeoLJIzHpi99RqgmDRphGP8iCvGk3Ut28qVVTWZ1P+2k/erob8VkkLLnt7Jx6ZunhCRUkI
OtQYUoFu1OmbLj66kHEokJ2cR8o8VteIpU/MViZMZlBvp+yHHcl51J4nOAz+IL23JGBt4Bnbuiz3
vQL4S9mee/riLXbSQDLIuIzbNUAT2Db6oJA29ZSBI4+7unt2FkuQ/0EAKBb7BfBm6d8I8tTwr1WJ
IboJUEQlL3K/NEEKqHlHVsvh2qYjHQhWYwOm6/dPWlBDm8zMMp2fnVTuxugsUo5qKVZL4/2plNkQ
FBxrfFzft+r/BURGJ2S49bxJVsSQoVivCymFRyAJKcycDI78RaWWfkujmSzKsBXu9ckNFHYzqB93
ZHKDNtla90/6GOjroYN1JeCzlMPZJM2Md1zSjfqkiyWt2lKtpnjoQ7lOjy4NjZjhwzmRzgdIag0D
nyW4jK/m5Nc04OqStbVkIDKu0Ueo4Hm1a8zq0Y9SHRIBVCao2My0YsMLxypFsGrrh2XfFBv1a8by
zN/KR1jKEou2I2PG4PCqLVzJGFYaICXfOz/IxLjEvadowUWy4lvZhX8dyZY1CTPgL8G5FkML8xIK
eR1few3n7N5dczUjfvkLNTIafZSO2p4MTpFchIfY8vYx32QCJJZjTL4Lhn407k6jp42wL5Q5Vl9+
vdaj5TEGddG65feT2SVCkN/JUxesLvm/nuxT27Ya/0G4ZEVg/R2rSXMyy/6KduPPvbOSsbYvNOA8
gDajgUUcCbkrM3ZFJ9BmCGpEoL2F9DpiZxuqGRi+O3Ex6+VjrvWtZvflpgnYAMXr7nRVBPDxBIYj
5ACiV1V/hsmfMgEJOi38/iBqT+UC766G5YMIQ2Ipdo0MzeQnkfeeMjyLHafRZq8AIFY9vr9S8ni8
wGPT9Rt9Xjuv2hUPC+ASPaMOUutCWNKvidoCm1L/F+yrFW743xHtJ9phMDOXTtZYZ/X/9Tn2y4y9
fVipEl6Gu2KzcEKbGUtOweSLY/7gZi4sCGZBtVt4XfG+Bs5YLAs1DTNVKHEzSx2gfnDmtC4Tag2X
CbqhsHHMZS6ncKHr0fIIYFi+P79pdvuTqhXhvy9l+V/t9yJT81MKA/KXKlDdTw7ZXVckDsrhNh2D
U/Ws/ZBxfjAMNxrUL2xQOJuH9j8tVpyrnMaZ1cB+WqkLolZW85cdSLk6R+gf6UPdwuOZf8dB2v97
K2LYvYPiyuS3hXMdTDMg3nYPxzmVQx52IXBpKWiTyCuSWKuRqAgvz3MMbyrTCK6aDZmCcIJNqXx7
mZr1APsGEbtsLh+a+/ZQ7BY4vna1EspMx10I4rxcImFiLai9OlXZL1m0m7xkP5MMolZNvuSGSMLT
WqoUaqxUqMaLOkoOIzCj/LzTckeT6epyjsyX37cpKNcjv8NbkiU79bX2Zf4aPVGbxNCsc++3wBVa
Q2oqvisqOf0SH3AhWbp2nQk0TA6C3hZSswMafZLcslr/gJojFDmLZVS7FFp/9PcFKubz83oil6Tu
1Q5aQSFa6gqOZ4MPaSxRQk7LStskvY5psYqVhAnZfqanku9AdXEm2NEdGhh58Qw/kmC/7WLOvDAj
oCMjGOK8tOE4ip7RyWZ+l+5T1o8/2Y2FzG0j3CTl10aAS3WE/2APKecM0boL4FllnNxjCPuJHaqL
jTxu8Ukdk5J45KVxRIm0O/D/KtwPW5d3peeGF2fWA9xtjs6wp7A2xoxWztFPJbyreYTBaCRraBUZ
VoG3ygM1vfidhEgt3CBUfO1kK6sTgslxZuH8Qq0ZLXXvyFNDwfmsuglILszPsd/MfwBouq8z9i1Q
q3ixNveqYax5KzoKmQfOTK06R0dujcyC8CR5Xs02c+ge3bXnoKCwWe9AgcEHsu2DenIZJWDeOOqj
Xl+kIjRJQOcT1HDvwm1YBvTYTGSmhL6zmKqqUxgYHQn/i04kR+9maPu9ufLkANaWOfgY4SLno9WB
HjCCTgkTw2coFcppkUkCDnj/DzE1QLw0RoPP5pRoAmPUR0+TmNCaPp/ujeWyHIgl7p5AydwA/ehK
MXEKT/jKsCX176pLOr3z8sx8zszUbGP+efFi/LL1UnuCfFGPAfgh6ULMZtaEF6h0KcXwVMp36moI
YK0D2rpAmo1n+uKrBCXgZbuf/OdsckJzl+D6Vj0TRdglCfblNxKCz0p+7sHf79J4w0uulcGLEcpp
I1EsV9+AVxwdHM3k3qwdVlfk21+G+r5Lf88VSitK2cnguqTa/EEYuKULxZNNNNNDBpoeIbDyhGyI
8LWtmWOcBjrz+rNSltUriUHpg3Idma6kvycgv/s4kRuWv3gWbjyoPNf0hfjIfOxDU9csK04qf75D
wE40v2tsSrKdwMXUMT9h05MOBsz7uCrnMpKRaJHH52govM7nyog8V9I1kKLK9+045v5jBOoKby1k
jnfeRyKv3abrPz2qlT4W4PRtYkWVjopXVVblXJO9UfpZ+0ZaZEyRw8MC79iF+VqK40ACwD4Ax7kn
TH3Qo8b1VrxpJ9Z9Ou6Rqh9mH3Q3boa8yJaoJHkMcoepjmoxrvRemUlzOT5hxcmJmMFtf9k1ybp2
spcX31jK2qjc/A+dYoJmVw98dzTGiFIFiKmix7JYpm6rrCNUMqkBqCjmDiqDXCdImm8hmjvzPTKN
eYb7g8kQvq6rNf8K66VYsuxk9kvl210Ou5mcrbafTxRuOtraoQonADw8KgEy6Ma588bi+G9XMUsy
HTK152b6aUcSjTYFIRIiZPSETQD16/6XFfIgi9bTbEV9yCHDqdcdQyiFuWT8eQz15jyyIVZgTlMx
xMBNon5CW46ugoInCB7VfaUdRwOmJZEtjVk1vRGTpKqm7jyAK1fbkfxp0WRJa5pbzBeSiVjKteTa
H4dtRGT3LcKLvspKBlsWKIcnOJnvyI/Y19tDqjG4f9O2M5MQcWve6mxqjzsDPOsiSBceJen2dYNr
jzBZ2PDQucvEVjHAUjhgiyflZQ1ntDPfVNxpE74xpovgNTrSaCrF6pO6gBXb8rAjYaQeMbTyCVLm
p898DAQGSJwXr3fG3x8roTC6L3n6B2iqRIoy2BjiQ/+2MHA503kUy3IK24pZClRj4FjP2Z1KCtYJ
nfEP+59PJs4GOUSMJEhSZNc16gzNGbhrprG7LcMAhY/WNL+BIaZ3IukwxBTpxB7fmOo6/QFLy5CP
JcS/Dxc9a4QeZD0KSqV9wDdGgnC8MjtXriIE0iFePjHVKCRDNwn6yvvUl7TMKhrr0EYosVCKkpqR
blbSbIjcLPV+qlAgonFfI5Jj1HDBwIL4C4NhOvgmuOFiox0pGUxkOIhpCJT9Gdek2P5sGukOkPcV
9C65BA3W3qjEWzS++UfCqwzpWBdIsBMUmNN9xhu8HSU0ee9oKBJA3kf60uV/yKKJi7mj3WILyNfG
8gjzoLDBQrwmV4b0QZ65CHriwjhkjPpP+l8WLD7IjMc+p+9z0WAPd5xwmwJwEVHoU1bEB5XTxPX1
vxbinxJd8ESlmDI7xh3cwwBdK//YrHYg8A/JKzxrL2alC0oUrHM8o3Ovm5a+OzDGr8ucwkto/nlY
KEyAPTZbaa5NlaMnbieypWSk3EQ5rMI6vLr+CB1xrJ+MuylHKmpAokDM0YOD/C99dfWxaKeNr+d6
s5BJD3wEAlUk9nN1B6pXYhcI1Qj/fpVsyNz+T3pL7P279ogLZybA+uScc+DCt7alqdSajWvGMH5l
4rLd27taoZdNyT2+1O2vuPJ/1RW9pZkGfDxSXs7f6CPcN/AveFIHEan3f71KeHIIk6U9jBaezbiY
yadZ6HboGIBBDIy2tV5Aojo+lR+mzdxb1xvNRzBogKce1TpkICl3nJBrVXK6G0krQ1VD2Ahk8Tdw
f1T0mFWIByYgj12sJFRciLWO24LTZT9cIeVqa9fhbrkFG/5LXdrnzlfdjLJqjU8KxQ1C1JVszPU3
1GAKKl3T2Vc3VxMlSFeBusrIJLGsGYJGLNGEZEoPdfzI/3MkvlAnI9nvjb2IdYc5bFgY1r44JMcb
jUzwgmCbCh/68wYcTPgu122uK/+NX231sYDPhr7n4q76qoneixi5N1taHNgi85euMnfN8JEQKuEq
hEk9yKeOLmBuc8Rv34w0PKNWR5hlc5QvKa+4+1bznN+qcKGPma4GRMpeY5L6YZL5Ic71MZYNASr9
qQcmFTweFbjsttx1XW2Vd/U/krzocs7kn+j83ppNl1osXSglRxi4sXuPKWBaoitAtA9r7O7nPQv3
OcqtGgF4QjOMFaMDz3ql/pC/F7m1ISvUjHnzgX1w+qSeS+taFE8rrnlu9v/xcvv57FhRJZotUUjn
8nfBhvD4pRG5W2rsdIJaVf53zmysXiWLk/34lZe+ZddRkTlbwOlJ8FHkMUvcNkhX2i12YCaAOX8h
32zJQYG89by7hidtHYz0sSHAsFBczDKVQQy0GAbwj0Rc2XxCtJDxa97ZrKBL9HkIVY0UHYjVOiMi
uPzr09HtNf9JWxe7TYsF3aXTb1GQud6gjsEMtQRt4Cc8FNI3yoXs7WYRnoYoiPnIPLknYaHV11f1
7omw0X8puiXjvADREv2jE7Luhi8U/e7Aol299CCbH0ww+s5fkB4dSrz6mrIK3dkka0ENMR/Xps7u
szyIsobhmIu7vgX+n3bEoGgSRR/FfefELcy0IAfbMNzQWyhFE+O9fEiYxwjoxMcguSfd5ltAFcTK
hsxKjijJdTloqMPEIjW7y/OkW2j4nmf/jM75gYVD04WpIGhzGUcHWvxQfOcds5NaG5wrcwJdU4MU
otdskzUeP7Z8VoJcysBJNavoEwsfyO/sPOnHG8SUdjKn3usnw3KLTHl29mNRir83n2cMwtk+WWgr
j0BBZRnTNF/QP8Vyd0nfGNHF6LKBQ0WRGUqs3progU9hTqd70ffp2jWezOpegTnGZYt7W6cH5z1t
IlqMiX9j6mEvbLOaIKgsBtdHBPcLGfT+/DXYD/rvtfBwaShOfEZxhGNjIfSjH2mtHQ9yFy6Z+zBs
ocVKXHoAMVE+d/hM+TELgTUJn/+txDuSJGBHkc6NOFt+cvdG7YdTi/jn+lRJLqbnNAnZ61ysvC0n
f9wFGNFu0WYv8Mi6Iks0OsyepY8+J2NO5aHt/32ISHdwjiyj7duKwaSxqVSmNwg5xZi/EcDpnkqA
hNeBdWDV26kP4vlc4X2Uhp62nPcjK0l+tFRqYlB6jrTExd7LW8Q3Ul1Sn3teOaINPGUfp37zClH4
HuhSRLZGNXrq1dvF1VoL0InmtgU8pcausqjoQBiasXvWLlKWgR2HhsOPs2dqDTBnEj084D0T/O55
n3wTCXASdDdijMD2Es+0LX49t73Gc/PMrCoGS60ZmRKzbINexO5Lxk8s6Mn6er9zTHWASkQGfV3W
Shd+K7rs8/4AvRwKdkoTNLiYN6HuBlqCo1t+gott6lxcDOML2Ul2OZeICA+741ukycLWb2IjiEdT
FAWmRWLdy9uzR9wp9ruFSuHdCGnm3e0/MyShJF+/4tZgF64IG9T8RF+XgSGtq6QJfO5zRvvEULh+
GP0W8BDbyQfjXk/wZVpwtqBMP+tp9Le8JAJmyC/kmx7msv5Q1eUDnZU3gpWDi74HwX9OfVXjb62r
dEkm9i3gUYfWNRRBYbmHTy9b7zt+Ud3CAeK1A/ztpyNcxsvIgmnLfbBE04iXEQQpYuhVPIhZYrcD
o8Azi1TI2sMc+YZuPlte9RG2sfg43dRLfDwlhp7fm/QZsbRxm1BLHOElP7ylyyzUXcg3sl1OQvb+
YRFIulXYyhT/QzwWjvb9oS7ERgkqqoytjhXK3GUzSdlUzpWs6XYmKMrmLfFtKL+wOrUjEnZtMmnf
dDxC0/coSQKJ5gXze+C98uicT/dsAn6nuatF2eRFhllHmZ0nMvQdTSWw+bjaOPL9U+NFxg+7ZWDi
0+/G/BYPfZG+ICxJG/pmc95rk46FjxOxUim0yevFKF0qIFWJ1HxOZuYTLbe5J9XzfO85zxB0AKRb
0njJfLmWX11AJOwIKxUheNheQsKXJT6qUfz56qhIPe4C4XQOuJhqs940MsBrWLsUYTlvjtnAxM1y
T0EtQYd40p1Ydy8x/i6AfT5F8Gn2ww4ot+T50EEFo+zYvN+Spwky+0XvV+nHSnqDPRgBVIoRtLPT
br4t4s0fm1NbgZDMx9lKE4DM9zcwL1TcAvKWIJFMmwE72RdNMGjVFLf3Ilr7huuUCV6pTNrx44Jr
BUz6GnJgqmEyoWm/9CrTS63VKVzVJ41nARmZpyRL5jKfnvUOPfJ6dc7FAjZrXC/vzTUyBZpigMCO
u5/40ejdVR9d9F0D/c0gRLYTuSLFD7jFMBZKU71zF84q7M8yGdvw4aJezWgQOtSyf567tkXpNp9+
fc5lp+C5Eq/3RhL6tQ7pCsT0xqWGCSxsHrCwZ1670dlMLp745VVLUdn63e3TXoDgnEpftgf/x45n
WVcfP+s5obW7JcGwOFLoXAKITYvSRS/60aDgBSw6BSSY66BzuXJ1Ry/3DsnSvD2QhqMAvVnS4wrB
pqMXDUSLYgPzlqdV+9K0eoiUroKWF3xmSj9P1ErJDtIAUlbkrNhMG587aSPj6WAe7S5Fs9t1YInb
a7Qh3ewqdsB18Uq6haEhxx1+UweaS5QKZP6/NyoTScM9+YsDA1lcucQYcsLNO6lhaXwBCcSeSwjk
NPLNvOwfXBn2rDqh/gKaVVZ8K0qcSBzkOlfcqIqGYZBYmBDDFLqe7LcECpmwFE18+MZnVkglbTzq
HFuaDEOikQBp/OPG5TkUVuaQQUcddfM/sVdM16nRd8kUdr8AKXEVW+XX+YwnAzXQUHSSltb+4u/K
jcPKIr7E4ZDil3xyRfa7Smc7zSp+E3+8qFCKL+1gO9KlDPwB0q23JTCTaAeIqtR4vGyx1pPT2Y9z
rr+K77NwY0pByXsMIb+oRy1bOIgPs5AdLOwZYC1ZMB3GfHoPo0CdhLlEIpwp4OEALQKkOJV7Hdpm
q73K8bl17gb9TK5VyHDkTx4BLJ/9mHu9BAP04KLtRlKmAeDD79XjS9eSgMRdbfA0EAuwqTX7/CQa
ALM1pSsEqtUmWeXifN4VsIbIw+Nap8DDlUEoK/FvTkwAsfrXmgs+ckptvbMef8tCSLu1vAvpqReO
yoD51oosTp51eqL/8kgFToj2GQh5a3Y2eTjBjEU+nHaJ1/X91M8VRRX2RNqgM+e3dfV00H6aLWGw
+q60qxSrGcKG1XuLixldhlrjCofAqMsz1OYR6015gbF6CUVzX1ry8rbdhq7nJ9MKKfBe32RHP5C4
axT/otPxq135YaDD/6tsACfcA6joAKSb2RoZM9vH7av4LH7UurNJCcB4AOWMB/NShHwMTzJtuMW0
LZN5jywhfzi2zAYA1X5nenUju2GjPoUhSS12S+Z5sN3NOL/gwVUirXOV4r/gAC0aGoeEbKNg/GG3
Fu7m8uEs2EXOUXH6KH9i9cq2WvVzjrcLkgNDpluLBZPCAzSlLYOLgJ2iHiRpfCkxT40G+R9q5n0L
N6JuXYlBE7gVAcJNppSrINZuyoqgaRDD9EwobVJqsafuBITdXQv2CqxCJ/xHAbFd6P73OnjVeXMA
PuW+YF0Ab2jGBO8qnbrgJTpqh8nRA/31s7BHsFvhwW8yIkRtgKUPVfgXG9yCZ8vYhhvcMvTTOa3y
USjmzvCFFSP4tbXgky8EqaU+sbC5zfb8ghmnPQ+YXngkncPmLEQ7JCoRaJTYY013FYO+bkA62Qi0
Zj5xvF7EXrG2/DdzMCcgNoCyG1uTt6KDVx7eLWhe7HFJjuDXnF0r2fPsOhaWhzICsAMHtSANpTeL
qKW55gcOikcGfse9vqKDQOpdZVjQJykGvJ32Ipqh5FmQ0YgMthIiBtP+N/pPdbYlrq/LtNt/hvlM
EIC8fGC3xKddZXt9CH76xZdtKz9wpX8n1wa17o5+8Wkp3VruEtJ4VwWJMsU/2CbxDsbxqHg5pnEp
lTG9OCgxA9wmftQwkSnJg6d0qfWBuwPN4L/oaG/LOe6jUHbTZyfE9ljR7bHFnpOrfmxpC+lmcmhh
fHOZzaee9cxNVL49yFmI0kbLNXph/j2zhAde1bNkLu489zpYK8gUn/BxvHOk6nvgTu+G5F4nfG1x
PmZdRRUxWriyCv8IywEpdDuxtCxz2H2cuwo/xSiweVs44v4SkKG07fy3PH5qae6YT28HTfDsZDwj
SmgVt/BC2ka7W7OyiIRl1w1Hj9bMjAgRtUk4E5EdUy1WBEqt3wUJoF/BO4sh0POEB63uWa1OKL6t
O7uGLH/vTlGtQ6sQ6GWOtpcM2nTKnldOJUpfX1nYCTZbYoRWrDhnDp8XqHHypU3CPSaXP5J0sbax
xUuDPeMvQr0lVrCflpr6F0pFcH/vLjfENLVo5GzzXqnVQJtzTYtYD1v/UHAR34Acc1f3/VR/F5e1
FRMbwRJVrSTjwpbLOEvXELKHlWN6jbkkYigJ/Qub9oSWl1fdVPDwQyzWubUrvAOA6XoLcAtuENQt
vae+1RAUB91sTqJhMWsHwK3k3nEw8Hgdpdf8ZRI365J8aW4GSCMWR1Pt5ixtzAsv2CEFTCs9ZxeK
PVhe5YsrqNAXJTs0JY3dIz+0rl3F3NFJDMloH6CmgMV//0rbyc6h1sNv4yEi03mBPTB3yP29KfAf
k3nTz2KDpvDoKHX10HclGwM0AYsserWfAMg7EUovnBDBKVvgsVeHGV5MH3i8ah4CLPsJ8knP32Ni
T3ZWSfPz2nPAARQIAJ+19ZjM0vNecm/lEanMt9Tj86dWuCpeHakX06Y3qaWM9IrEWEKN7JWj1yFy
Y/XYJnc6GPLJ/gdXDW2WbBnXrFUD4jy6ZMGmJGJl1oCxu/RhJqiCsnD0xkTRTJ4A0cN1hTinvQDR
3OIlKPv9RvaDHo/XpGPXH20bq6GVjxjxB5r1wTjFRhNYR4CyQTmc46F6JI0FZgUkXQDyB7MIGrV1
+1pHs8OEYh7b+GAj3oV6fUmP9b6ZRByE7Ig3qoDJgiCVCuLUKsGLBXb40tsS7gn6DYWd6+qXsWFJ
r+aJ+fGdLTCxXKnUoy8j++yr9CM49UBK2vi3G7FmWLEHwQdd0ArQspHFB39lfWAcyAKVI+xdRLv/
AWJPOi63MaAggYxTAV2oZjrj2+T7kdw+/XZkrQLL3N+Sz4s+zSN3K+lB2IQa8DIkQKEQtoX9ED2c
WZClsrEjZowUKm6xrQkzOjnTiWjC75CSRSSnYya29V1MuAN9ScO3Ezuav1p+mIizxyyH1+QDb+fA
F6bXMBqIWNey5s/GsniJVTu2sZSYxc/Gp2c3Lqf2QtOlqMVbfqJAQYRMPfEU4VSCDLT5twLf/UPm
/rnDWEnd8ArM46jxNbIUZKQSxv7OpzRnLaPeCrC4ToHeGdx/YMkO2shymcu8WA4gBS0CtdogjE76
wvu2Q/dCA4n5KS3aqtCVrHsVR0WYInadS/syVoAPmNPTBjnurzgbxP2PSIk2w998fRqYz6ulBjio
vVE2LWoPNoDAlPhOxcDjpiVVk9t+fYqdFply9JW9PNmru0NuZ0UjETCJSVo959s20+9ASOhpWRUF
Dd5tyxKOwLMf6yH/VAXTG7LLL0NjEL284yQ+8ifFtr85BI1bbb5YosFZaXJqT2uBuX1s4swOAvJq
8+B5v4TYk6udSXPQh88Bd0veKJDKSxQnjs5y2k660brxledbMCgkPbf4bHIQX1OkLMLkaPbf3XaS
IeOtYH1WlggPOtEB1MKbDqNng/9upAN5ztgjEWqcA1iJyVm9frjlS6HDI2Djs9nVhAyJP6PfF2AL
nBdRFhTjmao3TzixpCj2K0JIRAqU8nALWqh6YKpcf1CBHVtRJD6eii8IDhcu01jpfXrbQpSBGfWg
WM5DyLfzjmg5IbVHDSSOPy5jx2ivgf+ajbi0nsMB2fVVLonrnzqR5oGhIQk4UIjff2sfvxdI+2TD
uru6Zyd3yAaItPQvfrGa+X9u9BgmJkjXHpq2ghuwErLoBvgaC/jEHTffnsL6/IZXmVLpBFtm3tsr
E0Sj+VoitLAf/ryhKHv3UqdvQM88fIcTG8M+i1Etl7u89y6IcI17tkHTfzb56Cks328MSVMsMbfx
FAUSMRpIYCgmK8rf8qVm4TeE5AoHv6DxEimLP8hXao99vquQPKkwrHZB6CjcjGStqO68K2bjck6m
uSmkTV5maleA2CTQBQ6VXXf3TMfgnJ5cWpJQbDV6IfR+AElmsZQWsGlFUlM9ut9q0swAxwrI1Ny0
g4+KGBvVL0Q5sZROa1Awk19eSn1uxOGAry67Vn2SLJCbKXaCazRSZi7x3L6omfcSc8lX4/Xb7/ll
SpaWQI3Pxoi19b/EG4M2Mq3jPwZPv4p234/DEvh0mUp9Dzbyv02BTjbJ2GZfUy1LvJwen/wzU+q5
afwkrQnTw4ADJGqx1MOfpCiyrBn2x8foXjXiocISUcZea/QC84N/j36PTkK3GblKhkt06qSQlHbZ
DX1a/ibwlZAIp56gsHM2rvdIPcehYusYfI3lzgyRfkFI6f07ZHHiKvTT58JBnaPI8ai2EX0mqZrc
59IA40HEg2taEEi89LebGNoKV85cpKk23zbqrjUJmc3i4o8YIdHWSm0qJhBhpIGb9SuQISPTEWpJ
FDlvP+opbtKVikkbuY5VYeljCQZ2zA2e9MOSGj94wkvDKqcZmOR7A0LpECSe54QIO4UeJ2PD67AI
WzCUW7eSmGJp6/HKEKi/PLbsYXb/TzwC/4NSYk1zWUPys8+t1c0EIayHOQ//F8pCLjjhaQ1iXR6O
D8bmIIWzJ6CoPVkXJsCjB4Dr+196kfTwj+6Rtx8q8GrSi2XUmxdN6hH6UY4nBEcGNVlUyUC2k1tn
Vh0cldAF96ykNCtzmgkSU6V3Ev71q/dNYIKW5t0QsrSrCdHFBM1/BrHdkM1/UuPGpjXEj5dG0tVM
rtPaETd5iRKKGqOF3CJXVngJVHaODw2YMjwQPMsrc+3zkEctufKCq6PBUho6l8KtoImyZYzrXM8F
7E7ARmzKpEJuMNG7L/pW/Y7u9xz2m/b3xugKTWe+CFmRdjJn7cofFQfXdmTXfHio/aP4lDguCsxr
ugAloHspmocSK6fvQYPVuDpozQFVq8wcI5ZFMxSFxQg1i0MwP27d9wZ4mKIUn8VdTZ2xonr2NxL2
S9FNYKQ7RnH5RlsevZVF9U3hfOiwkxh6kJOT+fz7EC8xeCN6VcrRyQUg4xARtBN5qXlLPtEIfBNj
FVw1hx3NXzApErbzZbvEi7HKTGJg6njY8t3J9trZ9ZbPQt0PlQnpWaUFm/QFhOSWQEkRIcZYfgK7
7pthnATS8lNavYCAyVmO5D7GZoB/s4qiOsjnBQ5FA9tnquOt5JH+CAHIbt4zIz3nnUTxkV6YK6zQ
tIsQuTDdnVbcwxBNOZck08YcUAXQPLTwSz50SeZXu4o082cynzhZQMGlUfuxk2HhjqF3uXuvcikA
wCqHZDyvtAoV9md0+MO2FN4CvFTgiArcLUOaKxCxYjgHsePTrh8m0zGdftb9pj83/+4LOAoa77e9
ZubJgZBcWCPYzcegcqJQMeXaCP9uMytodoPJR+sY+vPXMJsihlcooMNWgFFHq1+OUG+pODculidk
tnggcFeI7MkLfqlODeQiqTTlsgDbyJdGQ7f/0tjlDlwdjvCgv3G8sovkundCGSCVgTbolQ8hHDxZ
mEZmUR2GhNoEtFKRnXpIAA9F+KU3OWGGEYbScct9ymPaGJ4CncytIiLwzM/u1BDQtI1hiUjaKBA2
jI5EurRwmury9k1x6h4WzpWrHUU1EJ9jwgEfe85mPJPjPaKbINdsYXHNvOd4fF86t91V/Cvk1ulc
y+FJzQxfDZJTDQREXzBhrUeE7JpRTSl8/DtzknONGFW10BBlAgJPCh4TwSinjbJmcZTXEmbcUsXn
87HEXUNEJR3qFgElgS11ge+HvNqzfEHrnR/L9hgNnS0kQHE4KWGYHsBJVhyVn6Z5stPzzZe+RUYr
KilLX7VKrLlMGL9/HASO2mTLmPbEgLUuajh207YdT9sxnO/KSZd//W6eEg589j5O+kDCgD4DkcG5
ZoUqBX89gsiUQsStDWTIsb56/fvgl1zJx/jbN+6KuwITkLG3Zg1Aozb4SPu1SPPB1YLY9owrDtHN
Zk+2tSuKqGKK7MLGOJ304LzyUA1TEje1DL1rnmsbo9vTlqKDfpzNcSz8CPhCRqy7k9/QVToDgNDr
f7nImWqiAcHqnVrbWfdZgSBCgc+TWq0YSfOD8fR0gme1TI576U0t9bHqrSwvSrhuX34rNS/UTsDI
pb6MwLQ4+rrGvbw+Gplrj/roJWFGiCePRrXvgHH57HD+sMOILHWkFK487pu+m3Jwk9p3bdF8p+i9
9fzNvEAJwH7rIymRHqTJZ7zCPCC0CdMHTpFtdfWJZKCq/Wu5IBVQwyaKwAx4I2qnZ0tP8v5wdoVO
x0OBPhuAJcY32d+qXftyjeRaImBuCiriJboKvAtpXEw5uXeq9tbiHOX/UtoKtNe7TFULwC3/EW9e
TRo6rYdSRCiIqlvx/yfZJVIEPNey3LumOHY07WUP2GIP2yYYpuXTXRRwRI/v21JcspK2ppfzTp5n
+QA8e31Eb89gr07H5WGQflT0J4AsDQRzbLnWmtKJk1yramdYpIohaZsOML2Rpe+fbwTN1vcLBiyI
L8W34rwfHNvoM0XBAtVBQvxdiluSVEQm6VSRf0yLVuVEgYSrQXDr128dcyQEZoKkfqzQCcS8W3CF
T1YI7jG+H1IY0BlM+mxNIEVuyz3V55dult2QVWVuDSr/siXfWddpxAtP6qLOkha00q9wyX07c5u8
YjIICvoRBfhp0ONMPH+EEYn2ghSImZr9yV0x4XKv+OJYpeU98E8eGTbVoD0mEp5OoN5BieNGogHw
Ml6MxyjuUyVCjuLkt170DWXt3R14EuEX1N3rOtw04cxY5SxLXmI4hu7IdFNXOlHwysTfUBN9darC
wh1H9hq60imoGhUQkkH1hBUE5BE49Z5k/nDcUQCoLN/cCrXUZj5LJoVXhDUEgQIYPxwtC8KeOvE0
yACf8zQvGLcvHeCJkTtOB/eygNZxeTcAFE6vuVEP02ypvYyo2EocF7Mnh1kjYTdiBMrLJLp+oBD1
gopnigV8AFcFZC8XPNptyIUSexfJebgchhCAuJLzC8uJMhKc7uixalScEC+PGtuJuHuycD6Fx13z
51WhLq5cwLpJ3Idp9NmtA5lyw6WRCvksWtgBU31ntSr/I4/o7GedRBtML9CTVhLUQY/EwEH5H5ij
/Nf4347cpybBcJ68OQh5G6oN7R4sY8B5sKgt/VCviHaBrFbrDuCA2J/2jUlCcRLT6pIkCjDeHZCt
aR5DfFShEs8bhUC/asM9D+J567v1xC6QO/tk9VShNgEuLnpan1qBB6JSVmnyXXZQuoQgjp6eE72s
i2KRoCJSKRQ069ESLfyrw2AC7h/PwV6BbDsXQfn9aEQ6qI1uoqncoMl7mQ7+I/NEcEpT2qI18UdB
zRkGV+X20ep/MplWXRrV7ELGTNmU0PRBIRHrVf38Z44jVHFfF4C+4v9gvO5GmiKZFkj9W0qZonoO
0xfm8cqPsJKaABk6gJ/a0Xx8AlmWLkueOJ9jrZkDON73NWsjkLX2PLirABW0iDqRv0k6Xyov8wOg
cbu5eZziPrbA4QdPoHxv/AD84ioCuI/+Fh2zMqPOmE8vgiUwzcewfr0AL7b1UBMF9Eyj1TwsIALa
DCUNZRVYkkm2vfg3eLZDWh9za6fCEAfwuNc4zYA/NjUb+vYSo2NptAhl2z6l76LLlo2qORw5wtL0
I91lyHwNdiUhB28Mh80OkeSryvDGrg87lk+kopKJCV02+SIexlfF24O/VmFEJO3lfl5Of12AmjyY
BWqXJi8SgQeaihCRapX9nvgw3uPe+gAdr8I2Sx07x88Qfc4UoZuu4q9TTFDkUSzsRKCMB4w18ySC
W4NZof4s3dVSRI1XA3ZhQTs9CjpsW4P0YPfd7KqmDUWDCAEyHMN7b3O4qXxX/pnNe67pwUD02+rz
FZ5TozYKzorFWh1AS9sKkVyNoMClAUXaW0BgCsE+US1jUFs9gO7+8VBKPIg+5Bb5TYUwDIHG02gj
i+kq/tHyJzpBSOTiAF+ZGcJ22tGajIpBtcn9uUzUEqTEhJFPsCwW2YVFP2gDMLrDvE2SKObMDJMh
Z/k1Ev5EPQ/q6h3OUbvDD/tfyAaJIdXfyW0AmXTOyXFHjtx965U1GzZAgADst20VuUdL7W7LSai1
rY74j+WwOj8wT9ThrVz3FQvueboSrnqwKWiJH/e0hhcwpIRfowK85SNPuIfN8ogKCOdWSCHy0V41
N1PuIfJUcNKz99QyLjQ7XwpcDoilgnzpNPIVDaAEO0yZJLOnEb0qW1XewS5KFLBFjZFyXCIMe+7Y
oiFRCujanT83L1uVeHo+aSO+879b1FxBLRLOOx2vUNvU6Gmsv0WCRRLmEoDPuovuMCgAVAlUiyZo
pYtO027oY/rPTk1Hlbx04dt29Q167xTRaAm1YKvO0Fq6xzzPjGcGVKIx4l4X/oSKpWGme8DYMLp1
IFx5vueW7f4SupJ0E1O5LwUYbtu/IiAAYIxupIACz6477kvFNj4xGQYU5sRQqKvH02XI9SoueL/d
TFnHQTxhs+F7hbjKIowpps1eJlq4GoHS4tDjegPY1XVxZytJMNXcriQWDds5KkVZCYoZBmuCEsDA
C+3UXWbwUvbBQP8TxFdUFljpd2rwvcsoTTLtShYOtcdOUZuI6LXs2TzKILmapqFf1VCrIBPxTZX+
mwJioSmAGtH6xeJeraVoO1xsJByFN8b/zBUWzeGuwRSjsJlV13cwWHoP1LsN7OK0huUf6wyOfM3S
5SNnoUKzUpdn/aQ8a0IrQm0UdrJiQht7NhMwifww7PS8C9nTnIq8vk7S5sMURYCgO3Hg8t3ESgIq
w8DDgv3JzTfhzUYI6jmJ9KoAGdXRF0inLQXB9FavXMid4bVyAn9YN9n2Qx6EIxsmO63i1etBbteZ
eaOcVlopJmqX3frffXZcA2FLinIfciAqvFCxvYpP71h5emjQnEZFMRIKiu1R8w8vdMu7Uud8ed1N
IsnFxr6WtVcOB1d6DTxW1VOWTWxQcJi92vseD0gn5g8C5tdo8SrCCAHF2xCkjejOVjOleVR3fy/M
tkRVhZd/732GXMQKrx23ZQRHjDwR46/4rYFpL9fID1AuIiaUqLEIstQgMXQL4x+/JxpVYca4prz8
E2QVeWZ9xnxEg30LtuBrLEXjdAiZ4cD/VLB6LAdjpVKnjlDKNM153ckPCwSNLcIgjx2Hdow/WKMS
2Xvd6nlDnXjWhBZXE8Cw9/HqlgE/k4Oi5c+aj/XI/G3nPGuYHwYi09t2MNhZaGZc47KRLQNMUbvN
PjYlznvdmnL9kkd2ZX35psZMTsuDM+vuE+OqT9SynbOz+JtLfy10BDLzp1j+1KalB56RsJaAbvmj
wQSJ5OGkMWEQdP3uvDZbVbLra4rBNs0zKe5swaFcO5qQQThwHpv5e9hvcG8oYTvdNvCobd3VTMX+
u7JAu0MjHJksfctaJHmgfp4y/LIcOjgqMXAN7/ze6NECdbEgafGg4tP4wwT4NIniULHmLQ7oaCHM
dtALpC0i1qj2bXcyWSmdlL8oTlFQpnKm4+VyV4jalqCcUDSQMRuS5HoVswOc/0R//qwUfiVEsj22
HpkJ6bArizXpzC8Jt0I5BS5MqDwmFC9s3W3hWm90MWbdGSvV+zsa6KaWInZs3OvdSpz7VvxMyjW9
pa8OMu21B+InzaLeBjB/AYY6/UfCXpcgM+Rh4bQAXZnKJr0CcG7uvk0ytLZb6C7eNz3xrUi8jLj4
0IXDNF/eLgoQ+yzE6XZRaCrQmCoshQdoqxIGyB2p5bYCypCuR+s/5FNf5cK5PWVDY0lI9FiEpFYJ
HkJDLKDkhmm9GFiPc8QSjbXg2nSOzAykcuRwnOeWy4VQSP98a9EvMdTOU8AIu+jdKoOrHYICnCcO
jDMYohJNhb0YBKC/xBhbUgC+TvR5eYfHVvvRYpzHK/a1Gwga6afr3a/LFFSdSrNlMkDUE/QBpbR/
VmWU6RFSx0+1NZocjxP77dzXASOf3hpUaFxC0h5kyzDPWasWgZV3eom834i2BH0sFtnV7OzcmkKX
AJ1CRpxRbGspyU1lYDNmBoz0FGsMprKqMHMlSa5Sy+t3VrXJlVbPNeZzDzUakpe/rlX0LiLVCErw
VWxCua6bHORiHUUetugAsOYO+WbSnC990jPQyArod4sWRcTfGuFiKHeu6KjuiUPIJtiedUF2CQHz
AdAq47Zv0yjnC5keOrVn+HtDrRZ9iaU6/nnQwXOZRRv2WB+f+AzKk+NnEHkZJmq15VDR5bRcf0qT
Cm5z/z2dJ9ETsLGCjhrFeungwOcFmAefi9Kfkijj1aQ+9XcxCypD1Dp+GupmbDeOjFuSQLBY4tQB
PHWYQcgBVWwC6Czgov/LJwpW+6Ml9eJZlIO3CgMQHS5fKFkbJy0mC5/md22WUsnzFKJZ1/Ce8sqQ
J8k2GGF36+Fqs78Dc2uAtRJPFFGmYOK5kG2U4CCInyH6trLo1xts4eKTIAUL/PA23vSuDk7v0Qia
jeLUpjsLo9zQdLIbvJiDmYwR6pcv9PXjnmBwFppAVDFlJtzf/4cy6ZXKNHTCtoOoJrctYrX9GjY0
+UPQg7X3gv29Y2CcZjFz0PqCpCPOvslY2wnfgznNhhvwOn674KmAydM3XcAsazZDm2/K6iCA6yhr
kNbIznqQxHRs4/+Y5HfZk8T9wcRCAyK/dGIs4u7nxQ1be8z7nldjjgpGer2RrYICksE1giKWPB2s
x9enF4vLoRk1NI4WwiVASygsUp7Ul6LXr/SEkLeKLxXVfisBwmlNUTHQzVl6bnz4Ts79QebdEB5+
JVDSrS4hWVhPuOpGWGVG+pDR3f3MCL/ZqlidobxGXFiMtFXle0kRcHwVEtIkPIkHxGJw2GK64lEJ
eMmm2vf1zWdb5QwH2EFyQWnO5gw4cWGcl0xpkQTL95Vfppi2f6Ve/fUhbzT7uhyUI/kMJMMjh1UW
eP4JtGhAoA99CUokxD1S2Cx7SmjNKEOhu8T26dI8yOXv2pgSD06CaQkhc/jQ0XldGzLu8/JQnQgx
uKSE97zWUatxNue/r1+GMKEPLXpDi1aTHBGY5C33mg6T0xQNFwbnQzCmt0QGw+3Cxbeu2yy5gZ1X
jBHKAytr7oID0SezZSz75kXC3z6GHaM292q22Z6W9piEkM2qyFo+bQl0I5kncfRbpVOdE0vRzTTA
4qcpHb5l+3gkRfIfeobivW7Rc8UtFJurFKlxoK6KWniBwT4xKYl3IjbHxqNSu8/gDv0/JDMhffOc
9FJmGKdEPoC8SG+TU3HaSWYxDsUQxtpDKY6WIcuhcJJbMbZaUQVRRX3uQ/TTkpYffjc5z6AX8i4j
cRJ01s5kK1Ld0zNSYuj8mtS5WnU0ZRnDtoh2ndBPSt+qgjyt5Ml+/PAjgXRrdgbuXmT8UqBoenUl
hhUf+WBfG+Kauepxzz/+rjMDQeclXl5nD6WG4cP7tez4TB1pGBufNiCdWt3ZRH8GDEYhIIhMvLGA
ZJmYWj352lFm5N4VdJ/fkMzaFbhD10yiq/S3ly1c21czcfGNIQCzDYjDdGklqbKFnTyeFsfG8Q9N
Zpx+D3WCoXbb0yM2QmLR0EwovcTk8e5n3t133ISfv4U4Qo2SJsxJW1kvX/T+zLZRlbW49xKKIVbc
CZUKTh5d+5DotysRLao9NfESPC12/EhuQdS6dow02CcrJoR9DhkzyOCuGmw9GMX0hQFm0tqcRSLS
aoB6Fxd+Gc2c8t2ttjXgaF4fnYq1QFXLOrRvocX8/5SHv0FifRmotiJvc4xYdg9U2C+bta6z/Yat
UrATzL16HaJVdkoNkky93HtT8XQPxbZemfDBqJ6zrYEUkfTX/5eWY6dc6MP9/e//NEFmCn3sIPP6
URPWnSyc+eogrsfosqrbJu+IHEYdUSWJo63v3k/Hu+ejUFupQxJA0cUdkSjvM/KAsaHFmchU3pNj
i/6B0EHgTHdM3yOvHJ7+uo8Ix3U6TT5exEeDL7yKkgrVgfoBKJiGEgWPN7iqN/M4sxtzKtQDqx2p
vaze1RVg9LFUz5qWl9WIYv/6wC16CAuyGQ1um2CQgDxlZx6wK/04b3FfvvYQ3U/Xlo30AdZx1/9T
ExBGOYb1QafOsgwHIxbePyIzfoUTJTcGj4H+Ya0YY67P3r2t/U+xrlHepZ3id+t9IzRsvPBcnwLN
ATq/4Dqf8fI+m+bDAxE1/1INfkBAac7hdeMf98Pl8DlYXRYmUNlR58t729nSpuf0wbhdOii/jApr
7lyo6myXOAuNoJw2i+Qf/nYlfL6/F0yhPvPXq32o0UjYlAZUMLUQ+vyW2A22taSLdijU0DfCJddU
AoqrVeSxR3gz8ir4lACLNj1CtUWQG6a6uqgjE2Fn4PjOWpQCD3JotL8uE/1VqXiueBib36sBO/jF
5x14kke+Tfy9s8/HCw7nH+6lWwmeFMS9LIoPYvO7odoQ5Qk/+X8Y+nI/e6K+QdCdoVsARJS6g4iV
HnMrmHBevetCqKQ3YiPpfEswKAS0q2LSjNqtijFLsckC63BWZTd9fM7A/vU1pD7PIwJU/6LMaRFM
oiIIjq4e6Rk0FdolTe8FDuXdRA2CXcryc2ECQpBCTPZtnZM3jc7IclPLbK31fhOLZtmztuwN27Xf
DJ2VT1LnBg4vfrDp+FV5Cl1G8QINdhiTWlUG4bQi74iP0+N3B+YcvJaLvz3Cj9ho/4oSOaIlN3xl
f/UI7y5dKRYJJK+WHjOT+ZBcXFjeR4zZCsaYr+nhzeWLzJBzMFJfUpufuMN1afjltaZMcU2rbr+u
p9xs8D0b5K7WZXtTxm+FKs6UpYOMh9ky1BVqJxfIaxLzz1vbuPFpF/sbSVn9BIsdxc9cVCrN7yvM
wLUhtmrVWUTS6W3SYT5sc7HtgoLM3sLQCtJfneOcjsWidwO/HKD034A0hzF7vkHeTw4sj9ZaOjIp
MDfXkbpRzG5/QZlmhVNrglllWwc0JtiRWVHV8cF8IW1TGH9ib89D4IU3KgJBdyWk5X1uN/KZD6Tq
yJQXJxxY4kngUwbSLESBdh8vda/k1mWfFfF1mrnS6XnMEDyLVY3ig4nEH2eDToFQtY0S2fxGEYig
I9g5BIeQuZxAZZOhj9qQDZGi9V22EoWarusNJd8zyakUxtCk8p4twFGQx+aIXh2wziZ5ZER6SnF/
T20068os6G/nA52BSCJzJTD+PgUiFL9QIP917XljoUn04bU6Efrms3A1e6rTgMSYxEvYTruSbSzD
vY01uhF4kJcv6MyeLZRRTxG3D6Ll4XTG98x/geRFBGxbSOLMgUSfoziNd39iGBkqpBISiOlu5XeK
khHf2oquynp30U6FXRB5oRA5oCsgYuDC+VcYPrZfw0yDmcFnslVho3WzVgz2AX0dkfnn1hlbT1Xd
KutL65m0nSQqVKPd/vsrc9WiQGpKmOHaZtTyit4V/UeQu/LU4sPc2T97LURaHgZfmHQ+VwnmeNGn
tRhdNErU2WwJrs474Nx8rQCfiIBEl4I0yCAHR51J8G82kOqzqljA1gDdS2SFCM1gZ/GTBdeWBkU9
z2RER/U5gVGRtegRyEwhLuyBiro8zHMgm5CAh8ct5x34DoZ+oPtNuxbGsZ8UaUEjCwHD0AAyQ7QU
6qXkZMErtCEWuv9V1czBXWWpVE5eqZWQDxyaywKCJjk9OT84covZIkYarZNGE+F2KNDFdSyn6TgD
MhJnT14jJqaWXMvfPOfOZO+JQV9aam3gRUsVcQ6t7+am5x+RI6uXr0cXkxAoaT8/g9NDygq2Mioh
7694wti751jihHay9aU+pjL9PIbMZfZQETtaUBMcVPub3whxdcA9MHyN04lHC4OVDYsa7FrUlsa1
oTbNOrWXmsk1Xf5HOIrMMQEr9NElP5rjRQbBFM7CaR63snfnpp/a+J3qjHbW2OFWKDCcn6+M55C4
gFhLMPeHcCRlzZCc6m16ieTbyttqSLBrCY+r9ypD8R8pbSdtFQ+m66Srw8eNVoeRIYiP0Q5rDeiX
ZT0yAY7NNqShrMtpE4W6SNgiE4Rk9l1qiFNYfPCNmodhoOm6txCDPmFPKQj0kojcGlf9/s5J2y2F
xMQzl74ofQRDZyjA2xrj97wixO7OqHySPgftCrF6QjGkyyLQSuWhr65qtZifidwfbMHoX67Rr8m7
R9W9n6Fjcqp8n6L4dpDwiR41nOquiMCg7ZvCaL789Y2U2JA2xp6Yk+gOExq/YZfweXzXQtuFwmb/
lSS6HNFnAEESapEcKRErrEw1SUkTVzZmtHlanFMbyebG1WSE7zZzaiurZgdAE7Ku7+qtnbf5vKqW
lD43Vc6Egyle59bKRrtr3Nc1YVu+3e9lvvhDhmy+OPH3rBtBDtV8Ha759XrSBMA1Tbk+6KiX4GXA
vS59z2F7HRH2Hq5gc9k2w7KORGhKlaEAT/gGuJ7ATH0RPvIfvIdk8kFZzq4XL7yP83HyzOWL08MN
JzXRhroKW27YKMXuMf/X4W/i1+skSF69UVkThskHfBZAKBtoDd6+bJdhwI1AdOww9HeGmwdmyYcG
T3DK614/smD0WbHxpR8SHF5xqQGc9No5JY1+I2thjMC8sFtvNPXRelXBagAH/2hrXdyqcsXBhier
NZYyIIubDZHcBMZbD3VJ1Jsfyom7U41ETHCBhIcLV5dMXUi9XTbgtJuWWlhFfS2u0kxwapLuiDSu
EOhdh306h80JYHSQR6ba/GH5bRdk+IVoU8tQ1dfPP/QMcwtHqrCdJPEUlSluVejZkJvPkWKkOaKh
N7swDufuXhR9tJh6lrfViLd2JP4qF1VQAADRWRb6W0CclzVxxGOWXc6o/hVblTKdlC0343nV8GtY
lkUvtv2N/no1aLUyFXjNevujuDV3dGgajq3/Txkd45U6NctzQYbOnwpEfsYIDRoYGghbNAzq5TRV
WKyf6/8xYsFFjlYeKmLcsRJrrIpgYJ5Wh8m6lfgStrA4E/lNJhGz5uSiJECeX6ehXcAs4itW/qmB
FwV3oXcTPVX32BUfgkRqXTvzqHX2QOwacvcnujglfAKmf/yiVpUH+TYbN8AUk+QuShBc8iY+v6hh
XZIdGYVsKcoeOkafBUdO8O5PRENDPT+m5gF+i4SC93Ci/icWyVXQXgsSemZFhr7WcFvfWz1iVVYW
cgyUz1GKjo1vMzg8HPRf8rPe2SVskePsGj63txwoqQn43VEytg3wgaKkAw/7wiuOqWPcoEqz3Jpd
fibRdg+ovddQbEMfE7mW5++wKX9aZWcKoHla3UjGc5c3TyOVJfWniCWJdszkGniUGFyUXCv55hpX
ihPstKkcOj6XYcLStJi4W4b4pSAJgF2LJ0gzGJyVkOK6BvpGotFx8ltDiFaxe61zU/VhvnG5/hhj
WzRM/Ccc5m87O+vPmcfzOyZUxbqPVxr5s3CKzNMWw0/vg2aDV1DclDv0mZIp/ezG1dxJd1aZgP78
c+WhUmJgmSSFUQwccnDnJMXCnvJEKtiMOPV6cvfIB/3Eg5vdnywnkOKkAylI5HvssOIxUeNe9v5g
ddwh6dh0Rc+4CtTKSxK5O/WI4AQWACtlk5L6CsiZY2H3R07FwI5ms0iZoWjCmfTTfFl1cdbq36Pk
kXprJOpAkrKmaU/h2Bxrc8NvS3AFfu722Vtde8p1x3gHTwalMs8CR2KJ9FhJMC2kknojpQQzncjg
gZW5MPAi/cB/sFPwaeIJOt1xSrsI9c++KuE9LVgsWK2HZyMrvDy3yCQUOyCiPyJqaeFZLl+/Xydc
vsQF20NMKPpismQd3/0Eryj89QoZsQdHxxCCoR2wAF1bK9DutlrlIIVfqIFdBFjDOEzDlDSBZLo0
qdQolwKBXBXiwOy5p1aPwu6h7cqk+viNI94Lt79OdYrpE0+CIC3zOH0IRG+5W3RGbL2NmjU3ayle
eYfdvH51M4w0MoZvuPpcaw8bsbVg6yss4Wm07kijimckpzlJZL1AwWX0NLTItO3iq/9EwRCg8pyu
VlOVYrj6GfQWgcEEMFzu/rVjEpmtAGGILPdk2EfR6bX/HtjklKiJlaEx4qrmeKh/Hj43WyS+vjOz
KBW7crccFjxWBToOiLBRzQdE9EidgOqT0qh+Bgj0XwLNT796Ae5kCDjM9NgxSHsQ9+tF7xgRw0Z/
zUHVYF4sUkm5nNYbe2YOMPpNBbb8ma2CCYAqGTNEB20gN0ko6sFN4CLiIHeOKJb2XDZtzdim64ri
1dBwK0Tmickgi+u1/NamjBuAvbZ4kflt8cWzpx0B0mHSLnLEg3yCpNEIybimTJrHKmt/8G1qOxK4
50OlIw0Le/Wr75lM2B+CLpov5WagJYXoofFxYxwixU0m9gcvIXSCI1uaJNevcy/zICmHdgCedLnH
/LhcQNWi2NKVxuZm6RREvYvFhaG8N2f+CEvxQNlvf+kDQq07LnfoxCZ7pZ8/3iSxtrlEParzAtuC
3InpqwKhMpG40YukMKl7WFrjuSEZZ4o0ss5wbSiq+Ddkl3EeMEZv2LfoAlRHjuqcWzUBZrkgpX+M
hcr7SBsldlVhbIEuUXgJUi0eEZna4UrQwPv4uhwUrXK2rEZ8M36uPX7F/wDZ/5xUxQ/+FSYFVaoD
SOx4W148b/MzqZ4BBL0aHoIsIPLghPp9w6sP8/RngPKl1S6ka0NQ6JKf5SiottHAKUDsMzs4EqMT
i+cknp/L80WSDvpbbgGsfsDcmJx/YPILxqT8upbZDYQSelGmayUI8HuzYywmVK0MhP4GAiBdOENx
TOLbaSlvnRFWnEOgX76/AJMaERCFL6zaefYsTxn4ywTMC8jwP1W28qjhs4oOt8XPrvoJZUMj3btW
wutRjaTbwCK2MA9OUsSufrJopBBqi+S8xzlaFiTWJDP4FQCEpLalreC8bJ8IFY1We9x+JNAGu+qn
v8tngUFG8usYOEDR/8vrkvDZJkxacVW+pdGR3WcE78zWUj0h8dYlVfubBEyLMXA9TEH7Q7pTgymw
lgdqkwW7919j7euts1TfZzCcvflmbMNnrU5AND8obsR1zogkZQnAEoWDDxwz2Kj29XtmHKEA9lxN
CYH9c+H9DC2L7b6/9v421G0Z/fr7SurzSKW71GdwYXl7C0uTqZK5kAoxje54tdUC8i2FvbK9nJRW
QMvhgvK6QoRQIy/VlD95OTXKSwMjizE++x0uRH3VQH+HwdLyd11OPJ3t6H+osZu1rMvMPAuHnoru
aGKsjyWz3kfYm9bhbqh/MzkkpbX7Z4SHPSquPYSVArBqwdaFj/Zefgomv7Lcqv86TdB+DIWTfAZu
1hPfH4dyfY1J3wvkzZLBn70zNkexbUr57z79vwKT+SeX23t5Cf6Hi68BJYwJs1cF5PIHXMOLwKcm
EBt614MEWqAnekIYjz7ks33UErChAxIXKZ630OZTwilTPJHBbLGZnDfK6sR8nAGyw6iGANaLe7mt
4HXWva8FQv3/6Q3L+hWStCL7iW6nqykl/bYhcc6T9tI0pgydURrHyhcpenMZHnW9d1Cj/EN8GkSw
qk8LqusEIsW5eb354tg73feJKEqqpOiAacRhgzaOVf9TLaf9KQAZGr0PoYW+upRYqOIVyC1sUfBj
8JCj4/NbYKXuyCLaGsiQaDq+q1/bAtyKQVIc+Dtk+eUQMxluvINWd0V/G1fjNtxuyqdjTeWHhaZ9
tAEI9Q2oX/ueRuhJRDS74N5xh3z3PIKWVRmP/mIvIra0lqJzuANdvmp2ltBdvcubJrbiB5xg5byZ
8CKuUmHVkaxwOvR12lNyNrdIqxlA3z7WNh+XOFK0L7v7A9PMMGC0afR9PxqSFjF5bPwY4s6pY3tz
GuzlgfwzcM0feHerlgZzpZZu94O7wZ5u5j3oFV65/HpmiLEfLLf7zT1o/SAL2ETHDMztk/ISsc8f
K8+m52QybK71IuF9mtdO18ricmLSrWanmkAto9hOZA7G855CL8BfIqRR9fFh/EpQgS1UEq6ioS5Y
SbTOgXXTNtMhV6yCQspAa7OBx5zn0Yfm7vxCmE2cmOdJsStCpkpCay/+m43o/7ITm7Ek2vjc+k8G
UpC+9d1q+a8M3EDNhCro8/DylQeuvi4soMh+3iCkhZAuWce1xaUBPxSLYDN1hbM4vJMiu+xJMpjq
Rn+q1PfgN8imtMPkDDx8r5qbz55sNk9bipB5f4DGnh2cXVfHboSguExQ4KfBj2BaCw9iebnNRme7
YV1jn7SAYTkmGbze8qENfKkEOSXZrKi/jStjHTuNigRZ9/gxkMvsMUcBzKkb5J9IYazApXMha5P0
qJd1gEdjOdMN4icDtLgXXwKPTC+3g7i6e+/cSaoH6DAuHL5pYoaDfD6Bw7X0R/m0b6MrI6kJhzLi
lGlXr5gICbbNjmygXSvlqAV8sfr75mUpSXxyCEHxjFNCJT1axqoYebfaFXOw/VrH2FH10R0gmNR/
xNiOvKc90yMB5oKB0lGCk93fQL9U3Yvh3z5OuOtC10XU1PER4AaaN1aWoGZ/o65WYk3GbS4bp5ov
Iv53EuhNxbY36UJNHVBGj7jWdLZMWDsEBQjCuD41vt3cpGiseI827t1CSxdzfFCjX7jXmMOPKH1g
LBfow9MtIBrs1Jk1zM+Xu62Xayut+ZUBQxL20FpcxjU8uMuQMPAIbbigb7ESMmnEWCAqNlcpfl7T
wflybHJGuaXTohuYYs5uhL/bZho9RYCCEIHYKzo1jdBmQ98movupADGGYu94uHfOW/4YZx+SFg9U
3RtTWpUUpmG49+SpQ6PV2xO5ZEKKn+gb8iYB0kyWjrDO5RNgdJP9G3hUu2mVl6oHA1xgS17ABxZG
jGkMpBXjphbMo35BaMujQdjKVqZkgFbJSAaZPloywZrZngN2VR8pom+6LCJ7IdBvG3DTno5oJA3d
DW179V5zEsunOmtxEYaFKHQUUSZazTBDXx6/KixIEQjBOylM1x5xia9TPTKD881iGZs08nNczXZD
catcidH+o3ypAZBd77QeGW5qd8u1Kbl2xSfaQ210Rsc0ykrqTYVatKmfqpEkVZe9/untZyceqZIw
TKAJrI8YcZAHXnKFfs86eC+SfGlVb5yQB+5M9uYKHD5SYgrXwES+/uVuf5FJuUSaG+NYEp6YIRUi
HCw0lb5V1K3mLoAKP+R1ckJpm0vZgS6eQOeodEZGH+hvmd2kaphK8dbfSI+G7ZL5rfXUNF7gxdhO
iPkauRwRav2S/1uWVM04p7hQgUXUXm6/HcRlTxbq5uRp63wDFJf9Cq9ZxnzXXCiu0FOYuZBJSiif
n7mounY1gjN73W8nFlMKu94qDSGUcweD2jw3ge/Xop9Uz0OF5IsRgNsaPmdGDQSpgmfBdEoCu6yv
phlWId/PhZasZUrvF7BBJpYqZpVf2tMv+D46OECxFvGGEZ1rVoJuiZMHTZXH/y5RShebYCCjYVpr
cm5VfxYp9Jdt5RE6bgD+BvX8w6CqgpEUOC3fov3Fyaz2z3Iw+xVxRrE0U6ouSYrXKpJCJ+RPcI3N
QYeptgUhiKu4eUypZ2S5ubyDhd7dIJNnsFbXd05i0v3znb0JFN1lP479KLV8ilH1dDkKQYSdcxvP
bi5v14EGsBdqCNGJ+lGSvRvjnjCYTok3GH+DZlH4M6wP1pqXtVqSOPSLfa9qeWML74BWqUqz3pbH
Q/bNx6p9XAEeCCMFv4+VDjnNeSJHnohq1SeWYaUlOqQnON+pD6b13GBEOe7lMuNdiTAOOxxs0qpr
/37/sRcJz1kBrG3QLQSuZDrba4Rc2JzA0vwmaGMq3w4CA3vEcRdGLeZsigVTMMmj40gRxvPjZuSa
9FszTLPfhZeWQntqBiWq2IQ/uKSS89MQUWFrseJ0LiIbHwAHoTQh+Un0JsMhYP+J53TytGJ5Uk/n
rb/c/pAIrW0Br99EUd0D+pHq6xk1bc/7+eAAMMQYng10HTf5Mfx8M68JOItqtFqd28trBWAgZccA
blD2zUPkFIgOAzpTsAr3d48jFXtSvZz9cFMFvKW9qTH2boJf5QExavKNvN6I7i7i44rL/mGQDZt5
tavF1RfuosFLFK5/lYAo4/g5+4LufdQOlgXjtCMpZeuy6b9ldhA9H2c7TK4PfNWi8CqgVSC8EZHN
sFw2Q5efyYr13nVbEPa/X29w7EcweFpj9+Ff8WS0eci67Z12NE6SPISsFChVigL0We81jb4CbNoC
kXqjxdfOD2SJtHsQCH1RJbUi/IDHph9ZPMr0fOdaDonrajyfZHsTY9apPWkrihvDfoK1T0Hc9lRB
ONFAXDaHRc0h70496o9AdA1rPvqaXVMyvAozzFIMVX9nlqUeFGsMRgSh9HHsIW2CKlKgtEhnigTH
B/SZAQ+IJo3eh+mxZX+5WRJ8HXG65mlxP2zKu5Ol1tgJSc3hnG7I2vX3rNNj2OIegxRQ9+aFm/lK
dkRKyFjbwsXY5Mvt4/jzmtoSg9h+dLk70N/IBD5oyvIvJmVJIkbpTGj5W7LB4nVsTKEhBwfBP6lC
QR2yGneb0MuKZwva8mTw1wQ4fC8d92gkHFluY9fI9syHEI5wkfpLeBPKmZI7JbE1z5yeqqCGkA/v
VWfkkbHedANVpERUHu9nbbikuVfRwxlKtj0OXubN/vl/ST6Uh4MzwuwLrqa1jw+5VLFrQ1NCsrvB
wbPFkIYW+aobzImICUfroS4YDrxAFfCTQ6dt+e4+aK0SyBwZMCSeUVHhLtCbPG/SKbm8syE2tjdc
cY6BaNgnG6JFggg+5NlZYEAI7nYo/uxomqyLJHcLG3fEEhAJeGD2A21AyEWfJnhbE3BcZKqTBd5d
QEGT4gDncRgHH1DWgN9LML0oRLlisRzB4t9Yeg4Qi1qcb3vyRN1UjP4x+n+2yRe5WT6kJoz7eFxj
0cHrGtZxIic6VW6a8+OW45RZDV7N08tno4L3NKtHA3go8Rq35SSdVR76JgrlvmmnJzhR2U0FAqUV
Kz/gT46nqAt2UOmhPZaJQXCHpn/Xc7qEAtupHuFfcf8YbQA86nGT7ZWUJark43aI+voE8DVDYfEq
v9F+uX7eVr5XnDwAEVkXsXy4GspGikZODyWYfesPaVOAdZiNy1y7vtSsJCFmn3jWj0ytPnrynj7B
APaIDqECDEJam7SB8+35GPpYqhgWsssx44P5fl/qPwyvUO4KMAabnAh0w6kGTJZetCv25IgqK1yH
S+AlsLO0OyehmbzHUy11PcSNDtdwN+G2A1O1x/z5ygRtN3nUCk6eTMbi0/nqTTm+iKucUuo0mFGn
NsOo5CdaV/WW4eh7AyqrjR+GJVyzbs2gESRr4sjLshX+MYXJXN35cJhpOn0X+yvgbhTAQrWVJpbi
7OJqwwD67p7EF+XCHvNaFQKckFWXi+ABb+pMN6iH7705Q6lLw8FS6EzDvocSE+nocGyPXiRhtOF3
StSgQL+hK/1QFHO6XPYW/JCSmFCfC+rhuviElNf31gEQPRzqvghbuR95n2QaFjDJNyKRrREbQvv3
AfofOK+ixNnYnWX/FSNw1rZxVVROWt+do9RQGspEqyU+Fhp8e0iw88FeLuqJpX77xINYXUpBbseD
0diIBudV6IOoGPDCqBeLiLcguBlDUEVHXDXZUAqA68hGBYg1MLdsaRzkyYdzkljBrndwf78QkbP5
0BOwtXqz+mBtrD/9vImxC87/McVkjvHDyY9+sCPg7SAX8vahmqJnna98jWfJX0dYGXQdrCWKSzT6
EAPfTqrZ6G24+5rR46hfMdpO3dWJxhMAHF0BPjmrrtyUb2g4szTTTX5DV3yMg5QewPFheaFW9nXc
b+Z/8oBkK4aizH53RfanHpQ/MieahDGfQigLNKAwvp79GrP7NKI94q5/wZuCA1i6fuuFD6OnyCdi
LSLPexi3XsdEqYyuKY6ST6uB4ea0L+roFDpGs/kUiXcbn2eCGoh1Cec1aC0i2d17p+T1yb4IVlX/
b7ED0wNtCpRQqyBCNFkgwfmUo4Cvp7B3Ry8OGNfYktzbLUZ/kv8J5ErXXrC7VWAwd5S+sPJyRyhb
rl8PXozqdQACS2BexGUp4AM8RFE6YgpQA6QhmjsCJqn36qhMH0WHd+uAYYubH5EQ2jEBUJVb9HQ/
waL/iTEZeSKmjaKvIa+JA7EHMijlL2nxjTA6zyiy0Kp6oxFGyFgGx/crNCITx+OvR+Yd11PxvwbZ
trDX9TG20MtUuYyi2MZQ9Ny2I3xwy4iKmcnbKz6MhRmj54TDsjUiBa49S8qvmC6ME4J0aVuCmPkH
7jtCF2p9H/NT+k1BrURFsHfx81WhSqDufUI1Le3NLY2OfVt55IFCSD23qoTB9tTeTMqiYimxDsD9
gnrWgkgFsuWeldeFMn9YmU8xsxG+MwGAp5k3yq6T/auyoOc4JTScmuFFRG0N2fWQgp2zB5GbfCk0
mwHh8nRXl+TlU3C8rfw+nJae/xsjNYUiCL+bLb/dz3NCuXvI42cqzUv9rU1nRlAq99sh+VzgCfbm
151VfbB0DlHOCPJNQ+cYRkYIEPMInFlkxaY3p7ZoPloSlzmeqlkuASeQNZxC3LOKsDlytCgIP1Iq
nlPFcfqTOodztXpwJcY0yzP9NViOnHDMY6T3miqSNLkVqqGJJYAJLEG/+AxNpmfqO8lm/W4dG07a
KCDqG/j+tNp+7aNRSSXhNe0ouEob1jT5VA/yrXJScR9DMcMUBZfv3b3gjwNNGdetb3T4BgPqcJNA
D+Jfyfwm4JLZ8l5J5omF3iMHdmU2n5ggD+d9nVgi52iRrac+Lv4cXFBuczcltfJ1z0HBTw8B5g5C
ARNbRNZ3kjMnEsq75tabEM3jJ1tzU592vX7izvJh6qJ8TyEkJX2/j5WZthHh1Mzb9W1TymFJwXXx
gOxhBFTQzHEY/W2Zq9N7cGC/nelXwyYjlKPxIArI8dqyWqPfrDVMUZ2gdWFvrI+lQwF5qOTWZrtB
j3K4MzmfQuYF+OWFejjg7nD0otp1dfOXAixD0ECvag287FwdsHeLFSbsSftxyZtUp7xo5yjz7OfX
YzGXWl6UNIlFR92E6ESNYnNV1WPES5ev/ve5LHa4Z0G/qD6ROd4WXqWaSGeYbyEP0H2MCCkW9xzU
QdSP/lbOnecJs8UDWsBuXQLQSEew+OJNV3FOv0zENAT7G5XL3HYEg6XGpPDcvjuVTkxch8eLDgHA
LaHZcN/3Cng3Ybnur89wgdTh+IafXhlhUgqFcmORzIKY7KG60S3/ZDp/UaLxqQYLgobq58Qxku91
4TmUCRDCef7YcdI4VG/ctyHA75HPQ99QbEBL0dNY3s2t7Yyhfnz1unWDw49Jsp1w2G+9kpzcW8My
B8kLg8G09fKggiFViCP6R+uQrVSyRptrbEWYVAynVs/8q2IzGXS9u+8NMnGE+OB+Uw7/Y/NJFAYK
SFkte9s46XTk8q0TTw7UpZPJ4DEdFBICEe3Qim628ebXFSOjKQBCLhqlDeBiVKDjtY1OL9OFkV3i
my6/Ce6GPYuIaX1WGVIxsJzoumBBz21a8/pPX+lL6PfXbQxOexGePY0BrIKI/EfWAXw4fjBeGryK
gkHBcmfUGiIl3FGvR9cmzvzfGoXAhztXQ2BdHp83IcJgK1pejaLRguX6a9XBQAOritd0ZKTmalWn
GW9oXDWprFZ2iMZQF/16rgvkFmmoPOoP5fQwlqa7sBcaCw9ZskK/u4AsMYbuhzN/rZAMI7nkvWVz
+URSvAJ+4aIMWf35XuykD3be6kXLEjRZroQ/NhhFbwtz5qe2y5wZf/05MeaDcIwhsDj3b1ECagvC
S2jrkFZLtZK/Ix00oeEeC21xUi36eOY39J2HEImhVe4Cc/pVQBnlwGx80INsz/sZCxGTEzzHUXnr
m6DoLIEBJ0qvj/2BOcbb1HzWpUgIjHlF2t2Tj9REKmQeVk28bcyKzPbcZwaBAjZ5e/FbmUt/CCvl
Ryj/F+2atn9tt3rcf2d85Hkvo0zy69dIIQE8FdESWz3ol6MajP/epFbMnnyXtbh5+0gbBULlvR8u
jAtCaFEPWxGRx1jZr+Ynd6ErIjTVsHZHgcwcqWG43UpXTcQZdHwKoaeCNuj9ypwUcDhme/mf930O
ED6p1Lp6xj2GCJfxawBBkmwF7+LhAOghs+FhqjpdyvdxqB508BuOQm9ppVAgnntLs26yAfivWiw7
BSg8MqYZDgAm/SQw+IpAcrg+R70ppwu8Me2CQsntMShPfpVxosDiTNdSlEI3C83qlWU9qU4oilbQ
IfaaOzwJ5RLnxtWM+B68cERLFQk2sxqClMKc2FX42u2Uuti1TWDQ3udOQHB7r35cavucKlAQ3OIv
Cxix8dTqOPSN4FlP16XviKKUEm1iabaBuQl0igBm/5Wp+Q8n8XiwE0Ak/ljMfeEuiOZr+GhOStD0
t0Uqn+XS9uWCsl3poMWKq0ibCQA4ORDlTyOOD01K7M9ucuA1enScvtqtlNC46HCETKYCrk5JMNv1
IemWMNsW9KC4LtHQxVx1V6/CUV/6IKxs79u6gdJe95EduUWws+QDmHZ456SYPQmG+94z94QiKmI7
KT68y5h3I6xsnud1diYMXnJYDWTNnVnEaU11Ou3WI2rI74xvxe76ol4I9flQU7ImmF8mB6rdRtzZ
fTYS/UG7ENI6UWdt7iiPu4OLwtJJqb52qS0nudC2LbeXHY5jMqqrV+ZJ61ATVLI2FHES58XsJ6bl
ZsQ5Byg1FQ2m37NQ/g0ou9ZNmA9dqKVm/kKnTxvA2kV4uVup/S17ItCSmtmuErRFoW6krhfKVpZ1
uzzjvqkMD+HseCucDtsfaJROF5b2BFHlFMITNsTbjIRcpnNPQuaV4DxJLr8vCv8AZQhtY33Owcce
Qe2kGt3vz23Qkn4IaVRmDsyNzDHelapdK4ONWIXChMEXwqEw1/hXxrCadTET7UbUCvk0gMYC0M8b
l/NYW6Ng/QaVI4xyou/e742/vJz3nUqFNGOwP1QEEOEEwqHCJxsfw2MIYEKvnd9cbFKzOj39M5xq
o/4dApyVRtrYsLv/L6G4fqPy+w751d32foXOQfpvmufusb8gC+0ImO7TDeZO1RUV4ZBHpSqZrlt0
Cz+D3nsvkC72euiw8reyRKuxsvhoPZ+RwQcSh46iQJZ/GC7RHzc7YuT9DD+pccF41q3pSPHowanG
6nn/vNXkLA0fnh4MWPNSZY76+EhnrIuzEi86wzmNtmGAESGF1HyjOQdMVR/6CpTWBuONw8M4YZVf
YzB7MbaWMfdhBFyFEjH+rktlk1seuyL1rgkHZZw11cvkIB4Y2dnhHQtZ4ZvkCJenlz0z5K0KtUJ4
rAkSxclApYlTk0EWoF1QIfYgXc8Ac9A1im5Mxc4hkLpIW+MwwyyyP4+Q6NCJxaGrk97AqTsSTd8F
lCpPpEa48G4ZiT7Ks0IyKuD6WSlQypS5vDKETxVHwBlldLSDLc0f+K+skDt4agChhhWyhrSmqosO
lKbCxL8nMbRGuYERupZi1s3puREgbCNSbcJcncFyuUaHpPYk7RvW3bAxCZkE6cAxMxDUUl1VXsiJ
cuZf13XCoxnmWRdTSvJlXlrECDNlCgToFBnGU7mgeE7YzJXFNZHfAwK10Uq4Oe+eQtlA6EdOJjNa
x1Llt10N8AYuMko+0tzqvUlUiQkkWkiCEI1CzZaLKqrhk7lMnX286FZTGyjCXzLBMGVMQch2r+5j
dIeO5nnWBNBl7yNmlOh7ZVj6yi8Ou9Rro9poWvtH1TOuIFsYn8HxS5j6imRdYjw9B3BnFnNW7IHR
QdUo+rfesYmTPkgfl1HDnKv0rJ5iLywC0eitHhJaP5S85Tv02w1V2mJANH7N27+DuXHb+k4QPGec
gYbmIsLHtAhDdQBtZ3kEW3VdBbRz4UTgGBHa5vJbFtSaaF83U6QaiWGyCkwQh9Xu6YlBxRFnpqaT
MTypwuV+zj+AxEW0QitYTikwe84iPdqi6MrZGiwJ8u7SQxWwUim6EMUDd/VTFQYpVOGXRfQqX5lu
MtzbiZkb7/4HOsFSx2D2Ynfq4j9s5eTDd/JHX0T8IzaYSaufINXD4V7YCj2mND0/asUfefKzMYUj
YVZ6BWeZpJnLfzGhVcM1Cxw9S/QvqnV+3VWJW2NRurvScWvrwxYWieNnvWRX9i6VlJ8a+WdIXHJ6
MVyHosiPvVs7fMU1qAjpgnffZsEQIxPeDoA7kT+lLN+LepoCgEYspkyVjMFspuqmxoX14iTrHtSE
9tG7FFi84CEZ7RXYZhrP5wCBpKkUZ4T0WNFuf4JtkpqdL6hjYjwgOfVtQkJFzaCOaE69P8RJoxAq
gnwC4KQOVPi0HIn3WzqOw4YwCoVCA/q01c9Aw0aFgu6aw7ZNaVcp5UsUIrYH6TJ6/AYqX1wGQoK5
tClUIwc+3Jkt2Ake0WHXCLTCtUhI9NiRCzrX8ChRedXjmoBr+HuweigBcEsUcQ1kcenm5XiJzPXn
KALxT8os942myHl/1pSr24ommdu42HtRHiriZzA2uvobRMcoQ5mk7m6IcUXAoVP5BDqsv2KD4CEF
NaMDf3+oeDoY4bYL5EzoYcEmPmqY+j6U/WHCfuT+2C92Vc7C85qlRyLnK/wOd65uGpDrZSiP3Xar
4qC0zrY7qE+eqWv4rwIBE5OTEqq+P27FOQtmV0q2l5FYDRpw8G2vPbprYk3Ql/AjXfAwixo4gDtA
tXfSu8aqxe8CPL4760TPuVpWJ36TT2m9BNAgaoR2tTMFJFnDorIHyGzYUuOTZVRc52EiUKufPbCx
vFLbodYzCW2eRu/Q6sfYgwuTWmwWxQIKXTFvvvt55cfQL+mzPn8asHZvPEvM/pEvjfQENk0hGM/4
Re7J7vviBbiTuHNryLiPclllBLbU5sjGkkArGIF9UEP0pC1h4MO20QICY7GD3kzZcnv4UlNejPbK
X4jMjBXPGb017SK9t5ftv7OLgBqA/Yt2B2iS5WdL8jZbWYlBmWo3VBnuIBfUgZ3kFpuXibvLo3Yb
yLMJ29cyb7tbySalOyxZw1VQ9vqnPVyGFBLtu+WOWNF4sr84EtNr4krUvYuOCUgHXmSusFqKg9q3
JoXylJuKLyLCrz+8UdtateI+Z8lomffs028EeN+mdvcvWHF9/c/RVlhbotGhfqJNyo0D2rqD+S9e
mDSCNIQ5lsNl6zpwiO7WB1GtaKuZYV75fHqmkaHmC864WmvBbamQUtgnop7xZzAuagwIuKKA+SOY
TzDmcms/lfeDeSVWrIiPPm03ilkclZlLZRhSmlW9CA8BbeDEVIERrNaBIp304hlYccpj7SM0++M9
61vETwgH2C+XrRtzi0B5OkOvW46l9HzPgPyPqSEcPEtraWvXIMJH4AUsmh3lkfsjvezDhB+1Hk08
yUdjcqTDwz4XLkn6w04VWQQUrU6/5Ze/qf9ovp0gh1XD3sdZNLPQUby5kts8m8KdXrHQlo38r/LI
rojBhHj0mqm30qtJZga5IcZ5rGuDbr//5CjKmFr/sWyq/SHvGd25ZytXq1irBuXDrxr+Pq42kII3
XhRHzutzqPnj8zEqin3Ce9mt670oyBZ4MdhHKD+3Fm/qU1inEFkBTG+HSo0rPijWfBWCjRjPe2bN
CfQF7vb57RLg8vHZ9jGAcPxWvtX6bBHkrX4zUujdoPR1b3KUFFmIVdevqczzlpGf08zOUuXdRVsN
PRN0p99PcwgVKSDgrzo0RcKsnqMdclS/8PcbQLkTXx9OfVBdReV+Iw1bXoKVKVPKcOKPWlLfJSp4
C3rUhJ/lbXu7t033A7FdPuzt8DXj0ydy+FKmCg3Tz4r197PlTql6bPQxiftcZ4OyWkRqtRMmfokX
8JsMunBLZUxz9UQiVc9w+Oii/46a0KDkQYVScSfUgiuILJnbnJ0qEKxcGvhxqyGiVP+tLm5R99eA
V8dz46VDoXvSh4t5hNkQqqAlkJ20xTCwB0DAozknDCAqsZgct+IqRBFE2GqBXLArSCpbTqQXT5U2
dbF6aHMzhXhwOw/6bFAp2Zvg/USoEfiwyqNyyYdUkR7+8or9H1QAQoW3J7d++6oMi8rcbV3WXkaX
uLOTwXVR4iJOw5khC70X4wyZq1ZB6SEXMza/ymELkP7awdPJ4EoF/EDb1xNE+flxP2VLyIk1/R0D
DBTfqHlxhfUAXrh4HIFtQQeRe+rIkZN+2ndyEra24p+2/pvkWzgOcEs9LT7h/4qpsOaKZT9nFUXK
zy/DcRKgt5vQ5qlHFtmJmekDiwGMm8w6TO8ElWUAL9BJYCFaioDFutpKb/6x2o4ll5rmZSZgKU//
+ettZYEGEsaYgG1sCyzF/olmZ3Dywn7qn+gvxqMGa/npO2k1GCUB38x86RPWmi6nl78ACGVLLwSR
43/j6rt+RM4db9m4N3kAi2os17vgoIVGwq87pVuROlMkA1rBuFVq1TF4rv6VufbW1SKVdmpGpW0u
OgYq50aEa83UXkzesBKCEbxXoaUEU0JjMB4XmyMp3QwFPiW7xqWTVwE6oMvb8u7o9OKFn9PqPvx5
ZH0PaDM7MsQDl7F53YvdFHXuL6Q/VhlsH9rdC/5jvbl9Y+5je9Fm3Pbw/3teI70CC7IAquourn+3
Bl6a6POUpPkPccDO5Jc08WhnTJTZCL2eXaTLKmMdeILTnuRsCGd04LysqDj07fzVrdTvd4K5X8Qv
uxOrCUrtI6MwlLiGYSMw+oKuJUM1PYWKE4zbbTW87tgmpORbRF2M8J2j2pRJdBVq+aInorJVPtaa
AcKmtX6FRwez4lQiE3Bbi+uOlU/169z+ZuNo6Zc0fPhAbgXYG08yToLOXKtuIl7dPnOBgJCnZvuD
szurJhE6BsRTm/1EraOkK9MQjAwkVw5luigpovoILPMH2JVZ9cd40/mCJkUyAR1fqxRSSKaIA4QC
hQiFuVyt6/+o8MnLf0SEoxMMgGKkHW8X5N696oHkhiX56jOHqi6b4ImctiwqzOFzsxzUKfFx7hh7
xtrn2MQwHQnZ8tDLcIMJn1OsWzHwGnum4UHv9e+O1UQa5vnO4TGz0fPUoEwa03GpMdrTikoek5eH
aemanRyviVzDNvDa7B7oGfHOh02/CgEFiQToVKJAbGzIXsGkGN8063mMlaKkJE7WmntqLgNlrhd1
ulhcC2cPNC1r6VvMfUHeMgbH6Cp3KTQxPmACmobRx2U58tYh5LCl/WvxHWhy6PtxN+iCyHU2B7iq
YBu2gSi3qkuIokzPfCY6/8Qsdwy87CD3b4qSiSWqf53aHEd/Hfhp5LpUpP3RiLOECGI/eXI0q5Zx
oE47jldB+1dRrBSPtotHKDCj7NUq3gM6UZaXLL7u2J++4VgFquO0U4mW+KybSuUFNpGEU+oGSDYW
8Rlci6IWIe6ZMv4xP2A0OKP3VOLLqaJUDv5T+MGgMGkTtXIIV4AC71kOtfiqyQgTFCK7YiS5UgFT
yOyrVGyjoOcOzNHgBVN58ix8pFpfWweiamW2klya7tdNVGTwagcUmwY/5KgydagquTVI9CvzTvMH
HTpoAZBZNCwLlltSzt6Rd0LPTAY03739r9Xflq7tP0ktr9YyqkRKbz8wsR/udBlGZ76R9q+t7K0n
T7nIR8ZRmc/Sh2WkeoAeG+b9Ht328WAhli6hQNJIdSYO/c8q6NDPl+8j34Od9YtOE4A7dILIU27+
GEOhYcQoxP0q23RBze9Ro98lBQZinqhd2PX7lSxZWiMpnylHRdeJQOu2yvRJZIYum3i8yzHZSh7L
P6RigpByyDokt3L7fhoDhkqgpHG+4NoyXqeBrfN2f43gZfBJPQRgqQMkkzh3zyJyYNl4LP0txQsh
waQ/acXWi7dlTJniHj8OYNdyrGgX+tkkUX/CKMPdJIkBAX8T+++JZtPwyjKZ/bfn0wMsgz/OnarO
iWvO4TxFrgUV51ZU9lQ/4C4P7bP3DHqlvsRgJK1viGRxcmaGPay0pFt8PGwTAw8TsSz7Q9HE7zyp
aZLaBgvwY0GeaSUndiswF3P66z7VwoHosRupLAUZi9kGJvNK232NxIj04GnuqF11KbUZHqAq4EV2
diR8xldXARMPxTa7ugRUvLWWCi7qpnU67Otu3Y6kkUbNDXiIcbkV7gzZSAPAbE7xQw6JodqpFwWy
zFoyTiMso5EgoBq2urNKmsIa6hA9JZW85pAXxz18/lbZBkY29zZEbBksO7nHeK5grt0gfkTn4Yb0
iuE9lk7LxrQa7H1KTe9ZX59mZSPDgeur/OSqwYg+ao6l5mZkBAq7xUzC9TeH6qU2SO4pqszyc+lM
yxmfOqzPdi+CUeimqNuzg4IDkS4LynNJJpmDuDfxd554798Wu4OVzhoSXeRIf+rFeoDzMJ9S7dqg
i5ueW9gnCE2tVC1JMuMVUD/oIy18vVUV/Hw4JZM8jWht6sI80gR7Dvr32ZYJAwVa6LukFx+sFH67
DXreSsSMe+UrbFtSGRAoO+s7E/jau9LTBZ9HrTOAtVG1Xh0EFtluHS5qgezgtKVfGkZAuenY5rui
8TgNorLOS/1i5xTonbA+KGg2yp6I+N3rpD3qx4QxzCmSg+dRJNoaRWmBkzYQwbu01sXhbThJt4Yr
0WqIJoyN3YzMIS7nQR6E+MMdRZfnKdOWJ3tNRwK/OmE1Dp0VMsBhaHp9QxFPyKp9uhpxBph30Wty
zL0HvNTU40KtGQ9NRV/0Dslcwr5cOT9hiHtmHBhwEPulnLi34Td/Cm30DDgjyZKb4BsT/q75SzdM
xxv2Akp5S1E3eFPQ2opM6Sdi9Q7P/4IdbRyPI/3kckzDKIZNmu7vBUlKrdrFoaj1gSzFkgIljKMr
Nc/CEiVlIizGRecs96o/L6rfMUgxlPB5YCDBJ6/1rtbahRp+rpfNRBKHFW9axOcRzAhy5T/gikwF
9Q3ysWJJJpjvRiO0N4FpTe7EQXlSDF22lv8EyG+YAWt2KF8VBO5io9VdN7F7gNxqWDfVvaZJKqyf
X+3M/JZxQ9dNeWARLLRF6N5LWuSScIJIibCaf3S4DBlapA2Z38nWfQBWXVQZ73/UqNiPLqi+VpyL
mZvl8UKahV7y99ShATKf5x2rXOe71b6ydxVDDh+OFQGSIP6UqpPJNQB93z5EYZFh5GLvq35Qd0b/
GU+NOxdH3huQqFzHLdA/GcP1R1cgFBjUe3DEYccL+OVm/qhED3SJnybK+tMrWwou0PBhPLHM/9pH
Zxnva8Uyhd/6zld/mCU0T7FSr6BJUSUglqTqpMHxxfH1Pgr3tvyD0lK0PcOZG2Tpz7S+B4iQxWfD
YWmReSVYIdE4UjJnfX0s+HYeaGKinzPy8ntiD5DiwlUpO9ZOI1X0rwJ/7wUNLUX+CVvCDIkUitK7
9wXRsXnmz8CLzLlRHxiXH97ys66tOF6wVP7xvR6HYFkhIZ7v0P7QSoIq1G9td17GRwiR+59y30Gl
LzMyWeo9wvVil32ybdtTAHqfJlqHcAxiido3vu4FAq7dsgc0jFCoIZ49KDHBJNf1BqVRcpDagM6i
LlDoGtzE6M+0HyAhWIA0Dlc4Lfp61vjK9LbZGvWUGpUu6gcL4kyT1QOLlVLY1sv9ACJVQQSJ0bnq
xQpSQKeLBgTAYaJw3q10vu9iNLszdIF6qWH6oDNoaM8CQHQQHhevShL29TqXbqbSrlzheaXsQflv
E2/V8XOqrNqHb1UT/whVAGbVR8L1iTq+ARwUpYaAGfk10ioZ5eSTMvLdnxI9WRrzs+qGXxUvxIS9
A1bokZVaU+P1BSgn5lS1LBfEzhcS+ECfF5Sjp2OaezDI8ktavZqxYelX6wzvOqUuH2jLgAxsjyyx
mWJ0c9S1XsAm7o1sj2qa5Fw0e3d1xUGbfUP6KK8CiV9eLGo6HJORQFXBXCrWWqgflqACa/8pwAp6
+5MD+t+bbf3Fh0HOd5gDKuv7sqSqIMjyBvNZkjWfGCm735qCamhty8fuV+zw1NSgFYO3GvYRJ36W
MYqVs08t4o3o1A+/mKg6qpv9K5SuyuK5aMZzpL3VCRcfedvEmUEu5nuHaiwuSBopOZEI/XxmTt1O
+lQ/2akVbTE4iWuL6+lKmi1fDE/9ujg3iENkGkG6Xf29HVTAKn6kMGeZmnkr32q8f8p7h0BAmVuC
cpZihHNXGwPXknH9BWHOMUuS1Z9/D+iYiJ2E0QO1+JNwWNIKTPa48yaHUnLsoOR+xDcNfg6a3qwk
p01d7obuzzXeQko6X4hVgEGNYeliUNM5pEhbwr2g1+UTPURH3T8K6U60aI/6qC3pifOKvxRuzHHa
eYQSw1EbyVDt9N4KTsBbtYFT5WHZOeBJ+xZaXkRgQruVo2UHEzJACN4Mr54xNZFs6v68u3/ozQts
BrYzBmmWMXq0EDf7pMdQWCXnUhwcue/gbenAkm+mKIHXVzmVFVXet503SD2pkJjCfhRBFsP8Mc2o
lIKBFyMn0LrammiOox2k0i2MIG5PGLrpU+gtYYUH06V3VFyamCaRE8Sg3NS3HhapL8IzrdOQqNAu
drQw+J5oXZDQcgnn4WNGzyC8zR0swJFTMOS2clQPmsEvAXg13zGa3IXlt3n5PsWwlUnFpow/0KhL
piHqA7GteE0XfZaUqiDATaetnU9jhqmneMvcJGgMVA6W+Cxmj9JHGkySy70Mu64Nvs8LPJplseyJ
0yEnokqqCV9eS02bR/5g7Y6ZpupBjNiH+bjyXbd2bWD3aFyNVpp9ZEQ/YSbmWRvOem3XCSbCzfmE
noKFS9V64Y04a/25mBsWDBOWQkVfbY8x5limsawcYsEQx/dZkhSHhmhOC2yIf+r1DLbB3Snm3zIJ
V1oVBMwaVoUE32u5MOP7IFHqn/ONmm0mQubN3iq6h7SfpBmlpl3C5KyUsr38e0MOZVWuVQvbbE90
VuyzgIc5thoUr97shNW8myGS5q6l9PXJTPP9C2zYm06C21OaDBDOaOVku2A/zAhLHRNHv5mSknaz
aB2IS3lF9qY/v0QqGPv8TtoGZZrh4QdsMw0040+ESVCCkEyEzFC35vi3sakWWQ88EDbKf2UlmgW6
nBnOCQOPkSZg1xYj8FlQlP8TBeGfEDQa0KVXiEtEU8T1WDnzPzggKl+9W3ln6E9MC8Cul+GI4VN+
OM7mzjOuy8dvRKxKGP41RqRV+jytZf3PDEsM6R05zVmERjV7162xDEvT6/unN8QAFIsG65DFrGWc
rkKGSGt2PyEC/BdjW/A3WEH4TkEQAopVOZd+/Q4CCuKGHt6MARc1CA7evmuSIKPsZWi33eEARu60
X1jE63vPMDUnrPqXnzbkOiXH9Juf5vPqWTCOQlLYN2VBNZxIq6qwweW5staWaL0WxKmOmauy+Gps
U8cwmvtD15BZFS5j53NxWSlVQpx7NmGc/+E+RfBu6dEyQc1xvoZig0BsRvXHZHAqPet2S3RepNAH
BDre0vSMxWUvQmoIUF0dqvAwua5Kr+CAVChTLTGh20EijUDMnnI3oIIZfOHnCE25+SQbzAN6ESqw
u2Ama8bB36gFUisQvftzz0FZwX5UcjpZSTPuDZGM11e60i3DH3FBN0wv0w4gyMqrImQCMUrn++V+
ESi0ruk6mWf6fZ5QGImzy1IU8ZIgS9IH5lUEPxSUKLoCoVhvereGXMRwbzcqv2/9A+sOdRm6ggPM
nqpy6vJyjTHDaTI6AWUWsAXLI/ZMrIyWDCB1dZFOWlXWxaLAsNt6a4x8Dhgg34zjQy5MgPQ3mqQR
utUJXrPMaJY0MrbHIwydsR+lEfhJJSz4+O2f/hUebaDQJpPuZuMMgzLdhTj1bTHl3Y8ejC7pUNpj
t93iwJM04yoYoQ/5M8j0PBlqMViia2v1vhq1198nMY+kMGq15pHpKRJLaNsUz8YsZDPE7yyMCHQ6
Q4wnhREWPfOitvxc1dWLqHsKMHe67pq8L8N1R/6KoMNYh1yIJAgsCYUDtjnXoOKp0MMYRTy7U/xg
Hk013qbOxW6OplgAdVAxV579hC/uLy+e4ty+pcvYFjnsSev7HXO71yzzAanpFToNSk4KsNLqnNLZ
naAUsjsDTUhUhRKXErMS//9B636nZqKEv2cYZYNYbwmc3U3MfsXxNJJr3lw5z8W8g7HaVmphKoxt
6Nh9JDd63YWiR+/rgKvVV/tTk0FFHBfz13KHLG1HiHNDZoGmVcvzCEjNGHqTx6GPPRPvL7f722G4
0pM4wQwlzmEm/sL3f8Go7cMW5QdQ1Dkc3JIQM224gVRk5XBdj/dlywPhrmKRYsGHOzl2bYQciqop
D7tvDGw5Ztq7sxjIZXIfqbLDgyDnIdvmXYQT1GXdkOBew2haHh6WSXE8B53hxzDkyJ4gxYdh1RHQ
iJhblI8G9wo9g9KxTJetl7EdhVsvW7i87PN/IGm6kwgMd4Ekt8bob0ehZ6qITAhL6SdVpJXVxf5e
KuiaxtE8DmHVPvT/H6+X5YQLuxUqzWqeAHfEHZrxfuSS3WO0j2WZSzZzdxAJwjtgWyJRr5+JQrLI
r8X/EfDmYatBPVvi523y6fRJQCpGokUuFjonaQS4xHoofYz8Az0JgUk/JUhJhRrAWqYQ6Ksdj3d2
xFWvzMoDHKvChfC1obQBMPn6zVPCOWqg0gAOjXA4TdJ0V2F6/kXvJG+jeUe/J3v7rBkgf8jmjIMz
CcuXpUBxlu44D1XCmBqiFjIfkXUSKV31HbeDqdAI9X5nzzoLzMbtUaiETI82VNIOBvOtHvCxDdeu
ZsrwtIbw1zzgvU6UR2BB4GUkbHGMhP0v+FyJJZ8u5a88SnSMbLaK2M/PUpgTu+wEPTYYg1ez7nIe
wVLaphGPMu+/5SXbhIn9ux7cx8EpTq0riYd8a9f+DdKEB01rnFQ4mZdrphkWZohYxUQwJwKDa6Ec
M+jpTJNKUyOMRirUaPNeGHqbw1EVJzkd+QT090R6tZJFuP1wgCvXUS9w1sHaWP/CZKrnyuvsv1Q4
RnhRkWxG0wNW7GH1XmNhjHaCxEBQY26CZQad12d3FnuntHUpTYEmG6d2UW5r/wqvaFVi3dVRx7w9
mLY3NGkCy2BFupUgk0C4FrnBvDiEZhrcnnDd8OJWnAwzxi31CK7itaW4bZ3GDx7McnCW+LZ1K8hw
CaACUN2VF7X0R3r/YWAImYRFILybsmCyk4rB4VjEAfKo6kz1BCOTUgFYF0uZNcdh+jccbEXgzKC1
p2pQZal1Q1u7kwS2rM7u9ps/xSrtsh+8im8jy3b5agk+6uESignC2qPVRyBdhyeQw+sTU1B8cE7b
HEszvNo1BG0wMOiSM74XlNB0sKo1h5QIJmPYNLUrTeWlLXiuvDycLWCq5Y/fMPwLLGcuNVpjlMoA
edvXBPM3TIqExiM6aWzBzHYT+K3B7L5qXWiFCST5dgIa9Go5xagX68EKUyxrYZP4i3WMzKMRfr+1
+LLy92zwDcwMMddm/kpDmLjPkw7AQxmAdN1tlmdugIzCPSwd5PKcaEA5hGmgYtZCm3LfT88XyISg
Iw6eosuZprDT9mP9b8JnSuKmCFZgQc3r8j95zfQpI8SocHBr++U9mXvFAG9AzPo2AP495ctoDgLN
jurcHASuM1rdLB1CA1gqofAl3kCWeK/uh2A6NTTxjpVwleqIQ89XWUQE2OaR9lARZtD78aey5v45
frDdDQFHBHp++gaT9j1ULzWBisa2MMETiTweIhKn6vXH/Zrfy3uY5kykPbf8bVtnSyT+Kmg3XZMe
EQeK12Ie3/+qmLC6F3qMXxObF8bAivB39okzYPsAmAKFnkQolpKix5EMAJziFNMI6612yftdtr8W
9Rq8THAPtaciNZ6SGLbTMJNeoXKwgEkIDDf1QdwKXo9/DzDvScnikJfDvVMw2Nfihhv50/Lld+GO
+2ZUgAfv3Uk/hsUeVBE7tv68digPnTWR4xCfVAZSvQI4M8JLP2+pNm/0wfCkNs7uhkZ75eHS8Pdy
c025E7J9MBm18wk9D1OZWTIevhvd9TuiilQWVM8TDvUfSlmgZNIJL4MHXkgfUhixgrGJIw5pO8rw
e6rOP3g8qxZo9/g+gHbi0JM6kwtKUwJCkiRPw4mRkunG639cC3TQfhPu10bw71x6o97CtTt7ET6b
px0RKn4yoqJZ2e6oY5NX4WkJYyOVImTgKI25fBFFkxfrv1KhGekbYmYAg6I7saekhPSo+35FSZf9
z32LgxBtGfbRlYArqnp1c4xKQaTLWvGZnel04D+ZowTTURs9BUmC8jmteR/ws4zRQW3uw6hDefry
mdQI0hvj+6A02jhcOSs1bdQA4jIleVgnLxXN/K7p3dmkPnesCOvpcPCzj3dmYUcExkr++Xd0qhGA
gsOiWdNPmiBqFtI9BQAB7IVsw8NltHgcFzqeRLFwGQrO8SDiIfqS8f6iXv9ESLdPcgvTNIoHHKAk
UYMCN12Frg3DSdj6JYibos1dMAgmTmIN8cCt6HQIDwekZ6PbIMdRdOg9OQmYkKZzuT5Pi5n1h5mo
yNTipQ1X1diz0o/LU6Zg3ub/EErmvA8Igwn6P5217Fnhce6zXm2Ltx/fPHz0dWXj1+JJrmzFjPRz
3DE7LHVl12L/vue+ly+5Eu/m5wvmY1lNbE5OU8Cnmzae0781nUUKD4Hw1YBLZ7T8cgNQDL6Vzddc
ksDZgmGfFhcBi/KzvJPt6ZqGC+tpEHZV3mq4eFiw4LBKe2Sf33nEhAIZNC/OWQHN1y2EcC7DxgL7
DdaVmmoAkj4xlXRTkJGPcZgNLp9DNchfXYthYvkdgd7HKQ3e7LBdbTfAh881Vq0quibr2Syi7Pxm
zMkhPt7VbYu/tVziyOqXbEIS+ElF7bRsY9FcvFTat7BxOw5QBSpls7YDitJZ18pbuGiHXU+/Lqnt
8v+wm5LhK6wtUtM2penxPS1ZI1ThugZIOz6FsyZoEiJuONHxnNoQVIamQAZzj/pUYDjDwhnZ/XjO
gyszCkx26P6erUr6kAtnAcy7YeY3KkGZjpo1Evw1F62hmTmvQIp4R+hrFDxaV8Bp6PuJ6cTVherD
+qi5WXBbrUM7M7Jhj98F/fwTG2qXY0DMNgPPEtmjDyh1LjnI4q+S9jI0Kb304m6cicwfLCVzzEzp
1OzMu/Gmb9z6fv7zbSRkSj+sMi4fOdmebb+wJZTt2Hr7NLXJUSVwYJgb4r73ksC7zlr97ifNBgPM
mLt15YiJiOA9h8VQ/gBGg2dI2RxMBRRZdLIrfrp70BVhHSLioxK/FoNiaaEhbOAVMJKjIxNJnPrL
ETLkyeAtCbK5cmNSi7Nw019fG1Yep0qleZ1v7VPh8/1a6GYL0iZhrZf+n8WzUt01NEBnouM5e4OD
qykf1ozLjVsbRRbt2M9ZY/YteHtJP+xgnwsWsnnqj1mLqeV7SLVgBIho3DThvcw1JarIfxlgy7AR
y7O7tcAiXIYHZ4RlAQsuMQye8kNreUEw+F0j5UrddelhA+Z4YsxpNbUGBhOx2+V1QbhapM4qEj+L
txk3stUpMG2iQMqLsdR+p7S6himIrg8JMbaIoQf1GTvWJUCGE6rbQqit2mOM8uZAuAR+/ppXJSz8
Dj8eIYjLGCU1Y76hRm2AVJJ7KT/VyaGOqxtUKFdaAkpJKTXTohLiB3IuIPxbUVNpccT2PEJpZSeJ
8603Ds9wACGNUShFk4Vpk7LpK+J/7dtVjrV1AmCewvuYSH76YM7kY8yZZ41CBNwRpoNOtNGcf3B6
hTzuHgFk/6NGzX+6UwwJiT1zjDsg5gXZfS+3DB89ZY0QcQglmN/bSFvZnOBcJYU2gawRWkjpoHa9
wvhxh/vBX20jCV6aWBcDUtLQVP96PoaO8MC/L1Mv7y50cX6ygBz4KCh40iHO58lG0NrZlCdsQlnI
OhX0QTLhnXe8GgWPZ/I8OvAVsTMHr8PtEuKQvDwitBtLJoPd5bhE/GTTwgM/8AdK+JnZat9M3L4x
gDqyQvd9z+OP/MVSJLZylO+g+n4KOPBVgz4xw8wXRkSrjBGEZ7j7+2OoZ3iToZqcdr4fyJtKd1rr
2gzOYtp6UHMg27ek6KAFBV8rj/9U2v/Lj7KLKi7kpYStoBIo4FfXJQr7fbqT60rFJP4poKRWopsy
cSM6Iv2IOOGW4b1Dd1dyrjFk1P1NYHrAOKmYqKoPy6msbPtXaLoKgDq5KHguEiG7+ZdX8xThHjBY
QL3DM7UtTu+Ps1iloGIUizLQugBNBlUlG+Ek62/vLrVW2vclcOCHe9j7oGY9szLyXkDK08EJPhHn
/ig6pRsT9tn24fiVPDZ8uICgCxdKfDzr8XFpUiMhk1IBVw+obu7JJwvALJGOPPTvxUC+trUFm1FI
QwdOLEYQOzE7nuxGxihmJf2BMI0P3BsHzJpLs7qRg52MukeveUSUj59RTUyObCi8/1TuHqB8XM4O
mN4CSw7etyV2ho4QvpPCmhjxMCEWOteQ3COyHfqDej4qcUtkXA8MPJpFQ5t226aZ2d9E2B/c6QAC
BoAiC0uaDkfm8+NjA5BeFd+rlEZbrQZ9+WBzxHY0De+95Ip39C+QD3yQ4mFScDJr43HzGUTHTf/y
+aNbAU4DD2GubJwcibyIBFiLB6q9IrZLZ5N+A888LZNVpSapM6Y7pCwitFi9ycafXfJfkMkUkt7P
uf+Pn7cowvtf75Bs1m3yBbXYLAz+f0m7jenDu/RqGdC34hAmNMAbzlkM5NpPbRQzfqrVTB5S41l3
Mz+Gb8SY1AK4hPPtZNeBGqNbJNcTp3ufsjrwbCafncGBinX4tn/6e1JePzqtOWVhnQnbjgQ5vEAU
YU5OP6hd3VAmYqyUWqHGin3Er7i7J2pbNNVXtEjnWf2rhWXqSC2vUUPBrIFLJUpBDozkRtw4gm/p
76Zl/iryutOCqHt5GZzDZCdx91eStS69XImK0Jv+2JTPVAwP+6MvBLKrgLtg+rS1nndKfFuBvlky
duysAFFjj1loSSohBwQwZpuJqaJqWYz9WyDe+7O2Y0BvtPrrCEuGh8hkXK0EujII/JM5/mQPLNFC
6oXBBzBu21f7Skec2OQAEDexK/WkUEu+YaNfmlytEBOfV5R19qBSraEsNX96HMgWgD4W1NfHeh0Y
ZaJbjONW0tfYfv8wrJP1rGBInD3KYkqfZaMlqV5p0jlvXQx2lVLOXf3mpq9skgE1CE5Dkl9vn8r4
mDgRwXcv/dNdbMPxgysUSDizzf/OEzRKrJIhrOyLc8F5kH+myvPoU0qdzi/rEUTdVx5/RbnNJjOj
gA/Fum0PAa6vZ1X6j8ixqUCmQjsv2QhTynkT63hpHsA3SSSz8wixq4bDMj5tYpQd2Yg0mssaGb3Q
YrrTR7B8nrkYZzRq33mG1v1pOjHmpS+FexQMq6AZQohH+rjlIvVoSAubKkMLHUjLmfjaUZ48uL1P
jMCt5hlJlbACeYfZ84USYN9ZTdMNk5ElaJPBO71zLCtMA96P6wcBylQk/eGBo+Qeny+8wQ0HMPy6
WcB5KETyR3PVufdL8SxBLy/AoiwjZy2aogK4md0HKiTG7F3dunNriX4AGuqPRScl19SxLyYtVRl4
P1Z3rh/rVtUvrSV2bAVcCUJRo9oZ8Y6pfSn/9W2omMeG0+8qSaHifR86L0ygRrdxEaP76rx4rBay
/hOqk3gVpxPqi+xV4PRIt1LpWzkueYdlDDRTWhHoroKqcRVYgshmfc2e22DQ22H3jx1Vr4KCtiYq
srTMwI+Y1sEcClkdu8YsBZhcBbHbwhQ29SdHBxvayo/30xXfedWJuorcTdF6uv9noLXaWJGZQcWh
Nhb+f+ETpWVAMb20XdViy6ctJu1Ecy9eEn7lIoeOzCWuoTBKanD9Uxl4Hg5BpGvmlyO/qEVol++A
gYQAKI8w8kF2OHOGXO+S8hAeWcn0dgGArtDrX1F16Orj8WcU0wU1hHCKqLBTzV5aFHn1IE7TP/WP
8fnh22aoIEzAkeuem/P0H1Ksx3Navua6ak/2TglhRdg/HPSUCq3Gl1CoWm98qAvh+Ep1vp5lbhlB
xvbBaG4FLroJN3D0xzmHEgGSeeyX91QgzeDBfWJwVTDYqXd2BKBjx5QZzBu8SHeYPUsd+jM79D0d
IkMaO5Y3yhwxtO/A9oqg9TfgvBm68DjxKcZOGfkBFbphj4s+uUPXYosjipIyrkvRqYq2aox7VPP5
lWKvNcjSfwEe4jhcbr5D/mmlc7dFzm7mbOSxaaj/fCDsyZ6dhZFRYjo3ygyIBZ8PGJcZ5DXxndle
X+Oqx21Wco4aNuRWXCHXQ6LGjEOULxAk8oLowHvfgq7LcPkzpRH7eqg6cRhqppX3m8c5L5RUpF/8
LslpkiTz+i0V1vuHLy7TKQkrcWkX9BykglSMd+XusAf9oGR1sVmaYMV2LKNWbgxr9hh4zdyeAiqf
kDEBE76ISLgMrwiVJQtxm9KnYb9czHMvk74wCiMGVOynrzjiw9J1D7Dfmi5oHsYKO38hVygFnGAd
mKSaMo8r9JSEuF2Uu+QgWx/t9WSyww6PETEu22edN4cYYFc4FZnFkFfJAeHeP0e+vQB46JAhjJ0m
LtUiUiCnSZtLdgNRFKZnTQxUXArUjP+q/sYV4N/n9w79VGXz+9b7uZiRCj0SIKtqwils3iH33Ov8
NZTBHjStrLnON1ZlIwJLiwevpliA7CGSIUrQS67G/3I4wj842feY5xrlZBwMGNFLL5X/Av5wvmS7
4B0kw2sN2ap4XuIyLsCF0wrZjHGZezGwfe+U21h/+XxA3IWHAcXgIzOWF320DlZTCrBb/sDxq91h
1UiBqFTyTbnBtKTtOyxxVjt4R1PhQl3LlB3eiC+K5JX3YLTBIS9YwbsZYdp9qy3Y5M8VZquem+QB
bXja1ga/AtQ8WhMXKcFcqcyW9DsqyphSQc59C4UZvxSlMrl1vsCxh2QFINlDM3WMk2wPYBiUUU0L
So7lY3Ipz7C9TnktgEfWduIg3e5D+3cv84wRHDzO6qZHnpnPj+tIN+033lHu1IKiJfrHV+PI9dvI
OJmum95gpA2LfSiO40cVm/nLXSfpX2JAbXNGkFzpRScm2ZkDpsstjwkyIza1sbdOYOhuSXJgacUS
FXjdFsfGqXiJj4hWpqMVcqpVscdqzdH9EVHWn1RCTS8JEt01Zb+322EhIaFBDBCKqZoUvBSeSICD
nquA+a9c69KAwYAO8ahPaIirli2emcTzuGutdUWgrV8KmN8Ea+4H9UwRMH7JskNzqxzp7MKOyM5L
hk/DlKeAafRQ15vTKulm7qYpLV9oscWiPHVdF/t8CXf98fZ4QiI8NIyHxLdwaB2QXRaWgG2dvVpA
rqQOrRLgOJeTbsLvtLSkgkVCcFCk10ND5BOdTxHJzO450UsC+J4qcziuk6y9a9j1yrn/oLN0aLKu
Jb/SQfq4ZeOxAgYTMZRB1SAwnLNxw1j0Vi0KjLccUmUUf4Z5BLAM0CSd9q2qjZ/wfQMm6a3ImwJt
Z0aSPxThX5sLh2+Jn2SafQxqabP+31dxcSF9QeR6SrZO3A2o9Z5mLtFuJ3qAmpk1YsM+NuOcIlAR
Bmr3dMKbDeCvfxaYm3247meL3EJIiyrQpJnqeQkfVX7uXjV9dF+JH2i7QrcyoMUfoR+nRE8RJz8T
n2+tq6K6PHrkBR3DsNoDovJ0JxJDR0ZPZLw4dejAnQ9DQKmAiZlpxZ30I3oYrUlzMZVvUlXjXjcM
RirU1KWALG8Wst1i7pcuqBs1D76gzrJpt+iCnYeAgX7lQAukwhQUBueS2fDNmH2khhICvuXSy6XP
PwBQABhb2uBKYwa9J2bdeYiRmrTNNHQEvKlIuWIcyn5RurmBXSV24MrBfrOhquDhHvS34H3BJR0h
YiPLxw6aI5q2fJYkCDZlK7xg6cEbF8f66gKreTSqSDjtjkraUCxjyILU2daZHVT+yeGBQDIWOIYp
VPks1tQV2Ctdq3qGjs2aYqMbuySc0uiLqpk1umDOxWdBolG0iqGhmGvWkGBjKudWTBpV55VoY1BX
QX+Y7zJoGWmhJALJ6PjUgba1JNGC5bGwBUL+3MAefGMoRNXTD6EJ+RNj+CVXXmxSzzg6IXs5tSsc
s3htZebKEWtFe83d1jwwomVIFxWMYIQO+Vvt9IqXy+48DuNhJ8dzPKef4jXUlx+K+5ckyK0/JJ0V
Lu84jD/mSpQCJQfBJOvxes11QXk8o8iKOG4iquaWMUrGJW/82e+ZCkMHmBCbhUXgCjJcb2MPL5uG
ZcdRQGbE7o4cUb84cNnznfIowR+Pf2Cd1x4v8kM/gzih0Zf4BMQFJFmdjxQ7fDzyTLo/e/P4fJ/P
QjuRL57ol5r+DtCW17Nr5R8AUCDlGYaqvp3u8iLSBEEGMYbG9yKtq4aN7O8ZnO/f/UvpTmOhhnWD
6zAZQjFu0jn3RFp1yqS/89ANSRXGV0V5jJXJ9naTdss4PnMMi23SwFDU6nRRwb6N+pt5D62IDmw2
iPlXomTWkancRmiefDK/s74YPhRX974PkLr1dhgvbP7JcadehTj9SMdguKmT/+G8sErIntaHJf2Y
TLu1GpN5yL9H6p+eLj8Hxf35PxDhCRDYeRwZwirtiluimL7byFgYCPZpa7OvPdn1A82HMIUJfZXp
kxRJ8c/NaGHvQse6+l0UYTLqq2B1/QwNT1o5IlU84MNfj1Tanu6VWexMKMHmdMR9Tp3o9mqA9hYj
ZFF4ubiN8Lc3oMUnaH4zdu84PhtfeD0YKqBbIBvUQblRNAKgYQI5yuDq6j9Kpy5oqmyYVA8R2XO7
x4W3xvhlCptQPCd7CdqEUubrwwc94OtVB39gDHl9qaJK6sXiucCoulsOQ+PMmYFkP4yGdTCYu+Kc
laSA1DUJiBDCs6UQ72qNkYgGU3MAyTiT95aHAwz1inJfMqbnf3XW08Z6PCnuu4TORCGPVwD4O1fi
7hOkFg4d0i7zkchc3fr8fmYBfz5p1jkawf8i1oJOfBTD4Rz1gupvDjp5hC4n26/awsuDiAexr6ov
/8TK/EH27pKISe2Lgk2fm2kgOP6Fu0IGWaVgbv06DzNcgXlwH9pW7KOA07vKn0+8EIhGjEGUPj+1
TDFMnFYyF2/WwbFwjPfKUp+NQsxxKor/i2tTSC0aTaodxsGdIy1h7w57WLGyaddNvvpl9qc32o6Z
ULYB0lXjPZ0FtYY2T7bXloH/0B6m0Op0Wf6/VvncTjlc43Cy1GyudJEfWmyYsvpdIwbkxhDz+mHa
8MhZGj6fvAbwQ5EboObA/cf1roOrLo0rnBcCCvToPjp+z0Qr57bzd3ajL17zv6IFI7ehllcNF86M
OmijVO0F8idriw0B9gBeZuZpGoIbY4uMAy35mN6bbs8ilJJ02T4nrsiRVgZhR4wT0+7X3b0Vv9eR
+/XuMbiH/qt1xgmBCG51CBqb6shvDhS2ydGJPhs3Z23mIs1Fv+krnVrNMvL3Q8ttiM1V8lpvTOsK
VQYEajD4gp1Z9TUbQs/gCh3YbtmLVfu/qRmnXhG6DasCaolj2i3bcoutsCsDaHQCT41LElVjgn+T
Qg3MCh791bViKYAiQ3D35rO52/TmyyGksx0pX589pw266WDE0vokzaUDuPc8Hq6bV+Pw2YnkxZMR
d80Ic9C+AzhTpE1CvG/b8ZD0iQqhHIb48ilcWPOL5V8JXsckkf8twa69s7L1gjbFdCAY9UHoFkN0
NXgul7k61eJiklQvJ3REMK3A1U+i0nkdkwizDFZnldEnp2r78nqgE5j2sUB43nE16Sfa8NBmYoOT
eZsH+AG2OnHXIDwg9I3AudasZUruseJkSfia0566BSTdZPf2Ex7tljjAR/2xkyHBXGwgfFlOe3m3
zm1x6CI+pbzGLMEufUDClXHSvZbxV0YRMXw1aqVONcP2Mz5MwXN10d9V9LgRLO4LJZmC1kxmeZMh
sRestpmzksOa8xLoPDMRMYDqpMpQ2s7Zu1c+z/riiACftSbrIi+qxQvUttsF3ym0ZhpJCkgJRXG/
xYUpI8GANGQR5HWpLXgdUzmuZHzcZj4rnmOz7gYf3mzeIt0aX/Y2mdX55+GgdOGpnn39o/pXoPDd
44EWPlj6gNAm523RPgzsvwxdrvmd4lcya4WaniezzWZ9jxyIRI6Otp+yJ9Ma6IV4cZWPP0JbMpPi
n/b7dBhLUX6BigwLp5IujSg8wkBFAOJ3chZRQzst+rKEVa2YjPXX6UPfH+y8j1hT20jurRVMlV4e
r8/ItfeIoSPEe8SkJsM1rFcq0ck6gOLNbeA5gjtHKLhZsgUMPnwup/MyEjyk8Ef46U5By6xsnZfA
Ild4pcp0kepIUJ+8vFeDLYkT5xjR9Om7lSR+Tz8LBgR3De//abZQztc+gT/93F/6myC69ILNRXw1
E4AjjMx8GLMbDIyRvFZgyqEaCsLHOF04A/7Igw9EMcNYVeDKgng20ikgRqy2GqbVWUK1Y9U8pAGT
3VBGVJ3HBbQe+vYo9kD7sAsWynJBQ3g4zdoHgkRT0yr2+80/L5dFEPufmNZoPD5mnrXn614auqQm
LJ3z1DKk5/PzU7EhsS0IcRSIsirjmH+yAOUS7w5k/pXrOz3+UFDM6Qr5kxdFElwTlSBaio6fym0x
Xid4UvodkFiiVSAbl/zEoHi/vRV7pFnJN9uHO6TNDpXhkFRT2+eAkfcLhXKbxj7WG4TMy98wuXVk
awh/EmVl9HFw9nPJrDT9tLGV7SOiDd+EsFRa8pK24VwzNkuQZqJkyyj3umGIgdzh3OHNs8hEWFLN
RnTTvtFcon0sN8CR7Cepxx6diXKfX/sPUrfIBUjkyzc+GEoYj+mMCRb0IlNc7bcA1zrw2GlWe3IV
XPUnj/z66s6rTcLMD2dK4K3Ht6OWQT5RoZ2BWegEe9AX3vBFxf0kNfpBYii2rq5ndNwF0HxHCMCx
a0UJZ1jZl8fEHzYH+jV0kxy/yt9ZA8znYf9I5UD+ulxyRnyOoZ6/frdNWEoGAXxQRVX15YAJpgYH
0oC+GCdBO+MjZ5rkQuzVazNq5YK3/m8Al2osPL+Ww+Icj1DYfFdI8BnGgpTTxgKarfAXBlMouZOW
eSBOmx1axAZ6NJcHNx8ObV0ZRBRdxPZc140b93JSuTAoGw5Z/TlRL7BiIfLDysD4XDo/F//caiEC
Ddr1oQoeunv5tNmyggyw2sq1iolFEwTwyHU6PD6twy/xbZ7fyzaBceaNZEVhz+UKnKv4EDpX/Tl1
B1ILAoaBfGd5GGV8O+29194kY43DX7G/143S46unUIHkDiQCgdRsx2tuxumhFB/PWcpJWzvYPRwO
eZyrJh3Hcb5ebxJIWU6SOAyfZ0g9JuoX2aav6AOI+6bN6ATTQaLTeeoTQgrnudHdUUuuYX6YkwEw
9+7XGl6CvKrTCM/Tj7fGKoXYpzRApgcKKH9t2NShqza+C6/hm9/4OH472Y8ec0rKFwCWECnxS+Ip
3V3JdI+hm1cH1fRVZsUBVXuwRsv+5JyU6aQLX08YRyjZj1AksQR/35lW5QvQJZ8B/4YGW2WWQdUH
O6s1lHuTT4K5JlD/v3uw9p1NPhBn/PhDfSqVv6atEyABC48V+b275iROFf/1GycXOHXIu9nYvUty
Y3Rhmjc2tRkYRpl4VknBzWIuTioxcSsQZlNTElW6L9qm0C0sTCGIK8Es+1hbJenRVzc2oaRTbfsQ
OqTFeObCEVV60X1hVxHlwq0imvD33zSNXwAbZIIcdxnQqGXsuds2u20ia+yIXCZlPCTbhUj1hjJU
TK5KjaY5PXOzcq4owV4cZw1ZrOGXUfz+XDqE6akSx56x5t5yc2oItPsxlBIjkAJCp6PftDYyd6rO
CpZpMnur6iLIcpP5ezvAQMZ6ae4MAqhdQsjFMT4CQ7wXj6OEvGU3n9ZqN9Nl03r8vof10KLRmJtE
ZIKyZVkqhRa6F9y3bMGllEX0y4rieK5LlLe95cNBfEdOCs7lVbCSkYbyFQr2GHB2BPzpi+e7LFmC
hsO5zeI/JNldPSvjB5LqPurp+QokpoNYpcfWSd40Cdl0DBl53/4vbII0cifdqfc0tUc+iIPcVHBl
k4Sr/AiYIXpMDDjbRfXtNUM2FLYig3hKV2SQr/ngJ8FzlJVJuMxcF1aKlK8OXhZ6LbDxGZsHCCmC
/T8ApmcNe/mf5din9FoFLTyc4+ZaXv2T2qFlgbfCR3yb/xiA44YXQek5sV1V2ETvSf+Iqh2TnZGl
oeCkzrhclLGx8HdhhGHPhAOIvADlFFx4/QeR2ldQ+buruFAkVFi9DfsuyogbRaKIbt0C63MWl3Yd
XHwNhgd1vqT0bHYMlmaNdvjPrm2+TWwVhiAIglfTuAo2+WPeI0RsV2ETp7veeR8o9sBdssvM1PmC
8f6YGTiS4H7Y2NJe6U6GzofOMek/o5blA5uINpjZh9qV1Qeg3zYoP9ak9HAOaY0oruE3ORNKzzgo
WQCx2saSkrZxR6nA/34La2/6NcwTdXD8Bd7YjTAby5m4WXKMkcWgIvxyadgxmS5HLbHhL6qX3kcJ
kJgjCEdaQK5K7HqOxggT/gs44m2QQmWt+w0lp123FzZa1IJyLFn8NK/lFJcMWzOl/J+NkRVEHnr0
euLSbBcVTwrJdJRAwMx+vrRbytYi04Sh5zhnzQcr71FRsBgDLUU86OqeUrLK5JMcl8O1OL2c2pCs
p96iIxIfeLAjWSvG9LLz+03lNImIpUvvPy0rTNUYYoYPTHEY6VEBwaIW3yIwjhO+7CirNAb362AB
JbIc0WppmtpEQ4V+Zr/fjEUZgpcUHnFwOqJjWcMc2aGkIHegllz/BpgaaWWTbecmVdGfjXTyEs/q
1r62M9Q1E9QT3OhKMLsJ0E8EYBXsZVkyJ1lpKlwcbkQKnfGjokfcA9G3kz1lk3NI1y+Zst1G97iy
EyFcvHsqjrn+6b0qapoAiKsUkk+pjeEqcDeOj3v7f6sR4n6rlx9m1AyukGFvGsGEbs8bbcj3SWhv
TZdBpOVM+xvo2aExpPJZ8khFGf3Q1d+5sRbxszfXNdy0aSKt4I9juLI0UYEdbi1yCVuI3rXgpU1s
GS34FW30P5NqmrbIjOWVF8wXFgUHsxCcLNdvuJ0rcWoZtwBaL+N1czK/UF1jt8dfA5qd4wiUc8Mu
jpSX2ek6hfJtIf677O+vOU44eP5o+Bh71+b5/paUqjzHOckDPFWjTbff+9mr2n0LM2HMDXC+DUKg
4fFdEjaJ9OSBV0CRYynxbtFLLi2N4JRlLdpNZydDCBP+4Df4VPLZqGzKji3bIsvHzpgkPWOlBHpX
hBBgIRV0gjiKbwgrxuwzN0kig79q0FcU2dqBtD0Qfa04mA+pwG6TyUcQIgHT7Yn66VBh1icgc8in
4rNBQbwvq3kWA/HKo6DfZFr92RlAiLiPHoLDFnxsoehNuhYaznGV/d05WbZfqhlkarDS66lbg5sx
wLHLnMnmOOyeW/9E5J2kgJV0QM/zaeF518uu37Oi9uzg36+h+24TW9px0ZQ5lInMktKDu/NsiKhl
BHKsu+LZMQ7z1vgGQqFu/7cQYpEItr7DSUldKk9P0FyLj/27H4cOaor4BPFyZj5tP7eyeKhk172R
u/kDlhLmDvFhUIjjMCH9LLXANR2AUp9qQdCu9vmBoFt50XBA63LksEFLtOCaErb0CFuvZLzWERXa
W6PI5OE1kq1Dnv1MkgGFtI4GJ/yUG1d1KeNrwWQvqGKO7dqDeCKzLYPEFSVH7L+KTOl67rC1Qc/j
JsEFVaX6TDhupy7u9kdwky+hyZNTQn0ugmAh/NsgZeHU2gTTrJLZEbAhoUYyZ/WTIUpU3wY6oFXS
CchV22wSSXKYkEseMLt9KdjjhN+dzAyiYhjqsZUfZO5/nzCRwiQMFAcsGKRAp+slh0rlWORu8vHu
zZQ3KsuWutL4i/N8TbrAR38LRFxqn7lBRzrzdaUSj6khBnGPSBFyzRGQiUJV2ojSNgA0LuUbvp3X
wdx+aPTD5jOyfSyth2DbCAfXIO2aE0Vue6EFLJ+75LlGD9gIFGxuryUJX6qIDdTxBTHp9afBLO34
Lgv0rV7a2y5I3+FcOeq2Zqvg5mKdDqY5445mSquHr6nCr1WApwm6lUw/wU5BVHhu5Chcw+NIWw/y
gDiQsA9GDQNH2b0FrOgzmBwGYwMrT1AUscU28PIx/ivLtjRJLz0agOFeLVvG7ymgKXxYHYVNJ0tg
PWcmTltH/C39QfwKU/kmDAT1P9U5fE9f3V01DPgo8Lab42q4YnEm6WJhq7o9LZb4LNhhn7iwLUt+
PaR0r/KXVPxgMfe0UcjimylO0Seux37iRi7O+7kMKhzf0onxwqGeg6a0F+d0i81XaFrT+g1in8Pc
Q7MWY5XJpViVgXXFuyseN0YO4xvlp/qqALmwS6NcXOXzlL+v41do/+yI/rXXz0mDYQYn06ETnU9C
ATptM88iVjDiaIr9SWJDdGB6AD+LpfkgvHN+GjOnxT5yk9vxqDISS55rkKyVCrKASKVjJZohVuVp
bTvrW+kikzj04Sm/uQ9/llb2Ll3CVClxZd1p5OHrK74ksrw3FjceJW0sjJQYgoz5G0G/05T3nWB8
NVL8C/4kqDoiAb+SnC2OJdyoWjSGW+ZXY/J9Ox5b/pbspIX6Hjn/LKsEaNh2pUe2ZTGc93qtI5SG
Uy9oWpic0jRI9rs03uN0Q4AxEFsrAjG5LkyoZe1DRMfUW3RTOfU+42zycx1LY4aDFyJDtunUwkYf
sSs3axijFozAKjnKn5P3uWPbVOUHRZT1yjA2lpb5TmLFi9DGjOynf2lpiDT811Tl5xDUotw/vPQm
FqMhB6BZS+OFG3mrx+nlwT5meTyrlukcgIu7pXEy2smZqEVYY1Mc8AdS+b9D5XW4v1ijBBDZy4vy
dP65kQIOi3q7bzCuSYrKztWLd2SmhUt+3EuX0P0zxMycpmvTtUPfoxi55ixiZ1/6CFk2+d9fk9FI
/739OrhdnGipWdZMusWyFNuW/vzV+OrQEE4bSPCqjS5bNCwOSnb2JCC9XShTUozmPpOGrDFAZ10p
JcGDa1HaQVMzPgVAML7yeWK7oO9FL53qT5xGw5nlqriS4RhXQv7gnAwRNzO1075FKX4EbORKMbD2
h4zkcavdOIIfLxKjZJ+non0uSrHpb1mqjknyYLzBZozjcxVtpPSAW7eUgyyaxH8BNtlUrYKG5V3u
/+H9vws5kz8uQd4S34fOpwjsabGZiGXKaFxcgI4W1gtHJ208pI/xuBjhmRM3rSNaye6wiG2D0ELM
y1AsXS418QnptJhFGIDkQJEjKn4bADC3A7QIzeXshxjjSvwHpJkWlBmc2X3meEHwdYlPGioPEMXp
HOUhIzReyqrIfR/exTbIlBEDMf1z/wkXLPYfd+vKDO9ip2nZ4WrfmGazkln3vgLaELbU+2xxyBsq
6ybxqLIYz19IaeQDOCeHtQJ0LVKT0XUl+uH/cdJxcj5c/4qOAnrN4xs8Jjs9pv1W7D2y8NfsQP9I
nH0F/brt5woXRnJN+aJVf3QZdZlb14VkXA3ktDDA+nqAYOHOUHIMLzA5H+/adqUyavfzVZuEbDon
ZKC2UPjc3BnCZXYDkq2ZSKv9Q5Y+873pT6DKJ6iCOxAn+qpP4iGSZ63RqEMWN2uzOiYtbEmflLOP
KHzx0hxR+nI0ZI+Wgj3I7sxmKH13+6saM0YGTxvNV4wGssvZ9eTv3nRLHnOqe/9dwtPd4QDkcckE
bqpgW61MJ3yBmjjPWpy2HzHh9S7bNcmjCgsGlmHuOgPPAbgUPZwDQDuDre2g954WggyofuUC4r8e
cljWI/pKt5BH/31dutHKgqtDuBtW1rT2SCQBkRnNis2eml6b1ZsvaMiFuzJ/e22AXtnx5T5ERbhz
K2qgLdJE2QUE4+ccGOHavWuoTxkR0VZF5i1ctHA+RFb0GtB+uNOyJTycXvjM9YTcTjmYZgLa93b0
yQeSde9LQsziquE5ftmf3xCzI+0iWsfzBHGgYgywO/D4jzSePoc8bQXKpirm4Y3nzQsm9vKQStCp
St6Hq43/xhnrFev8Sd3RgLajsxL5DxyUBe9D6a+54KOCxNGB2EabQRY5nygGgoyazs5w+nFW1wPP
6MEUhHPsksIyVpwDsybS9qMB2GD30KpeYslTbE2OD9TKZpJOZHWzAdOW6Folaj8nq8PD6BrBNsPo
+JrWkb1wUntIwBwkEl/uyfP7bF43x12Ztglegv5p9coMXGzouL9s/zrVdKVYkpx+nG7LEJa9Uitf
7y7Zz68nYKVoxhrMpsygPcefnqSEe+G6dMXcA9CzRpAN/ILaPDD6MHivxu/u0MofJafrsdWJTW0M
Z/Lz/rgSOg6U8Krek9qX2815JeWMduWV96gggyYQg8cMoKigU75PykUiNY3k4P36dtRaOaalxCw+
mjdTok6g0LXD41h7hUt1p8uq09y6O9YWaWecfwgHGoRt5RQPDT8CdnCK38GVGwL8iZodF8Ee1xvU
kBINY+j22zzl2lLp3estvDmMTip5aOblFAL5KpVLSvVjh7mMFS0bXm4NwUDKVRpCaJv4uDk/KilM
/Et8MbOf4wIBcjbpf9mlXpZ4jq8e9LDWqUpjrnLyiNBUN876ptYHIps841hypeIMNN1dYlMG6Kji
3ZJ1wz7LOx1TFy5C8Utwc2tg2oeKO56l9MlzMV09lmC9V0VRX2zMSThjJG7XDVr4S57r/3/Ko9MY
InV77IKabB2JLDsGlYfkVMVF2E/JWc6RWF13A3XXVNBYjHtmPfZF/jklYGpqm853gD9+cVWFqcXG
yzuHifgnsu+QBf0pC9nHc7M6y2Flh4fNIJUEUIB2v9OSXCp73T8hWQn6ayvq8QhB8zMciSfJFu+s
2paWqakrtlDEtGYa4KytvpHhRtPm57dVjj1xnubDB/L4IKfir47CNIy56tWKK+gkR6ixkVejGUcU
hOZjtZWq39dwtPwVOnpFAtTEyRaRBEV6igOhMBXuxb5NWVpV0T4igUp7GYo/qzJ5v/GtEsJpGDyJ
Zm3rZ03X+KOqHeiFXtvrle5GdSYR1VzKQDqf3NFdyZGiMypRYmaj5NgXSkTd5r+BfRYfx9fZHN41
Sumnc6o+w0QUVd8iYgNYssppx0DWZac1LAljmf5Ro8dEf8oY3fkwod3SAAPixx+UM8YGoMicOG3o
1PT7QHEgVu2RVEo3nXfuEJN4jsZ3jXT0o/nqEtXLe3S0zKnEpdMpS2Y6dI1HdgKkDVj+VLNJCjxg
4t/LVDmfb++LCc/gOHAsb1jKfzkAta10i86gapYFhTwppZo2u8VGoPQFB7Yz+S24yzaHeiSr2nWs
zCQDdU7tg9OQ6SchPGIibkjUGpXyvwn6liW0oGB8UyBEriYf85LBjpy+oNRg3BtKd/F1x91XGLGl
zjSMyE2BNZGJ5UmnXi6pBfxo/Fd/yhiYHMk1T6002RDxUV9QWFLuObeqTULK46RD4fBhhOcdFjfK
rYJFc/tHPt4ScF49SooNxKaG+mxS+hGkV9n+KMGJ5AOcEbod/1cLsT5EMuYHxx4RhLzRvvu8j4Zp
6J+l3R3/e4VSlkFdnIyRA6uv3opHV2ZKWRLZwI48vTcXatONnFkgFBNt0XF/59ZY5RHySzDMmyvp
3ev84D19jcNlDa+2DguACR0bGGaI5fekfNgZq468CHaBqmSKUlq/tgprjo2BkPR0P/Nl66Rv4jPp
HbbQ7E7d0I3El3u5q0b77CX5ZpHuMEmg5WxXY5hmbQ337klaWo3EAsF1D2D0YOMHoibe30ZdxCBS
OyhFlxbclmbPEdN0sZTWhC0XptYjUHgOTDlT2kqdCCewFBzM5BOqEBFHPYFwsVI3Lb8SV2a1yQMw
xCrhm/BEwFAfnWtYwRpzkFGqWifbmBY6HHFTs01udhaZTE9tReBED62PrzmWTfhyh+DbISWQ8Ui5
6gbtfpd13CmCqIn5fAQc/DG+CoA6ZyeW//15VAZhlh4zBMCvw5AQteOBYF0KFwHOs/o260mwPHf6
3pj7+yDm7HiFsvkW06qFV+XpW2EOic0qBmTWmL+3GpT1QqNEADWEU3ODpwyU6kQjPALZg7g0UiuR
LNfqzM+HTCW7So5CHJ4m3kX/LVzvoOJhlubxm7PfT+B50p0+og8ULGesmfnjD0B5edOiCCscnJgI
s2BNQxSjr735oPYVju5H8HeoCY1Y2LeqADGoH5D8Zm6Vhf2G4WRQJFHmrQHVLl4d4w4Oq/1EtXOW
oqjh8esT/5EftCcrRpvrjK+elQVGehWjdPq0cEFu6tKoYh1QXZ4T16x8KvKmDmTXhV829Af51gbC
Wh+b1D3RgzfxHO0jDoIxlwMPpZ/4P+I2Ux+JgEso17OAvpJusPLQDcDiF+DXiUwunDbJS2oLnnL5
bVKZYwZ04NB+dWis2v9TeEH3yTgxEK40k9cPQDOQwz+K0aEl0B7NVDj1G5iNGvb3FOBvmwIbkMMM
eFPpWCoHaoR7LnY4hYXDpIEb2zp3D4hk5bs9oGODZTY/Ze5rZcyzMQgXFP4l/p6QlUynUeIZta2+
GcyPxM+XY/iQ7ve4tka2FwMNhjW0Y3lhnw5mFxQ14WtfbzRMXoGboXlcjXNHmSBevG/3+wVRINbU
ZhEjWXAJRDC4PAXCtq+4G0LXrQkuSZQNH7Rh8WhcEFjMSDrVYWLtIYjGB8z9AbxEDkRZG9vx90de
/EAJqxjAGG6l+1YfCh9FEElMS7Rx6h9SOwyvTbgUTPtdexEFHjwLLmJ9zOQOQO0wqXfDPjiCvzg1
LXOKx+g59DEGs6Zlk/DivP8Fgp28Qj66Tdo518b0ksK2InZHRcghZaGcnYOa9COLroiXWVBahW2F
ZUsN6gyMhtBBeOOfpvQ1grWOkSN+BpGZj4vEznXOTPksqgeY1P20S2aSMMPoWbRc7rt3EQ5HIP+k
W13nVgxtWx4B5JwxI/xXANT7F3GSRrxAIa0wLiEIUDY8JiYkSkS5q2/oV1Y0hMJwwWGz7hsuA4qr
BxcN5IXxrThpEIbtxLt8uXc0ukBZZFbLm+2hInkS7JwRdajJFX+98TbMfsn6Y6q5fYDSkGunx009
tHgfJ3QtSFhQTzrytCUFNtvBUoRCCSnHYMgOIBzTPwDXJCcEL0TeeHtn2lMS+Xiq/MNdD6tRaFaE
UcHQ2GL1u2slW87i0KhwhF3ATy5wDWmDd8kOI3OFlryTqzLmah9gC6tVQ1VRXLDQYvgKbfu5RRpE
fqZ0hYcShVLh1Z0mXhmrfTLXYSjWi0TUnuO4T8e9k8CTFCYpKnyXOZAmyoqjVdB5mgrjTqfJj2Ee
84OuAZWq6+EiqrqUqJH4y2wruOG3Ejs7GmKWz23wfCVnMjuZ8dBfAHhsUqPK3bevJWElzfoed4N4
u6iFsOK144EDFymeH6v9igR2J7USWtu5XqhSm6uKubBZuaS14mIrtijDW4xFYhaLeVpU2KFozMuI
FYNG9jLFPurLq8VvStufrVTMme/ULzgzY1Cr5hsXOrDz4z4P85SLTb974hFxHDxKKB1QnM8tqSxV
swDm8inJdrjKNeeXluKLOOzmmFbsI4/l65U1QNnx2NkcKDnaGhd+WXchk8zIiefr8AjU70FlQ6XJ
OSLc3mXk+mhsnlF1eF+pHEqMRI2tsrukY7qb6yHYp6FlYR5waaXApCrx75n+d5z22dpVgzgbHhEJ
NZBceuQOoHuJuL/zv3aQ6CboLlWll5TH7o33xXJrByOIB+FNf985LHR8cEsFkcVczoIGARMKIYfB
EJEi8132UYu5f+oomOc1L203czYKE8twpBrzyhxDSm1DGtBE9L8yaPw+Qr7AlpWkwbU25a9nRvIl
ldJnOAr5zBykYFBvCruSQuwBMwUlY1L1FOYw6ObQk//cgohLKgDJNY2LNLtJB/O5z5yI84h4KRBJ
YNHamiU8R+HA6QUxLm6dLSWz0Mc2RKNNhKNMoNtd1BCm9LYs4Um14A1vjM1oIFFFtgbu+GihBPAC
ut5KAi3qdU5JwVFRDd5QuWc2Pg3SkYzVUxeI9TZVTYcv7FZqF/DcidGMdojLrZp3ii/BQ7gzqXMd
nesOoqk+85198dND2WdCPdcb9AZTujRQuxrY5QHkIApmLH5yJNR7J48zh5ZzO9pHoH/3Gueg6ZcC
hEeAnYH2it2ZmVgPFdLarXEj8er8Zp9J3O7OnxlP7iZaG9IynymDF2lAaovx/Bnz3yMb4GtY6lEf
ftdTZd9oO/wjuEg0eXGv3FjdIW+Viy6iedQ/u7+8dlFa1+7POBBO48OIytUKSNzC4pB8jIagq0B2
qN2SfUz8ymFAyOXHKvY9jaiGCUe4/Cmy4HJW5xoUdH6qCotMTJd6EnjgQ9fCTK4VemaPyjNh9okG
C/SenrwcJzNe6ya/M9T7gv5fF3Sd2pZyWS2qs+bhk3aSmgLHJKCjpissEO7wChvG7WiVwkVybZql
TRA29m1STz/14NhhC8umvh6kA9OhFHimsw/f9jhSKPKNRQs57I2Ix1TOe04p+0GY5D3plJbtT99T
aTb2osO4lWPu82Z0oD5zAb53UlIgwG5BAEMoLaIguCCOGwU+kOjd54hQut5TyvWhQnwOe507Z3e6
EJlpTk0IDDRknLChu3/d04fCnjIcffKeudt9e5CTi66KD0fmRH5uiFfzU6JOTg1H5dXG83Gj3sUR
91u/yMx93wWO/7njiEo2ZuDVbBr/9bWlIRxI53ipQZW17PkZQf/dVBTygI7quQ0D3toDeAiUdQ9g
MjTi9M19r5iKWqt69CtlFWif23NiGw+fuqSwmGM0J+ty/juMHYUzu/OjPiguZlgL4NtjDqwFepwe
hN/Ohl7HzkGnNsvBZSYVigxlXIB7Qnihkxm/YoHnBTkbP1okg5JBk+c9VCsVmNwDtJy2lqkHxXrC
HpAizl2hovp5JlqZ3aD+qcz1GlUCXEPuyZC85neJW0YQ2Hs3j6FuKO+TyzHbCDiF7GytS4BGeHve
IMaZaQqPr+U8DtLFIwwjKuyhgM22QPSo29gNAx2TtCVJjjf1ypNBi1/myQwKPsl6PjPznqa+Or7T
KrmCuglN6ZNvYXb/f+7hB/onq2lHUV5qHLfnSHocNTdC+8iPlzsiCMRoPwetjoIWSSd+F4huMoAq
56Yt30E2FdQudUhobhWt8mlEfy1O3k5BoJV7khmnw++A6LZDeau+ptu83B8/FHvi31oxGbo6hafj
87VuNVWw9yyOGueyNxUV/PYmSxZEmeWADOYTSRLyjoM7/sDIaCc1h71tXdQ1EMlyL9Sh7DsLRfmC
MvhCZu1+zzaYs2ApZojAjKYmnuPwq79r2UhE7jD5t/1PIdIpvBwPuIGjXuAoWlZ+Nw6tDSW8wu1U
Lmysck6xm30o3HG+uCxUnDQU8DCYSjUZTnVjqwLYsovSKmE7wR22P1lCgDs4EnfImJb6qNNZiDOP
YfggGLv5XnRphfY9g5/fRXBVv7QMHoECWfimKIQMW9cPxb7CLJhS3w7K83GgDeHv0A+CWVWCjYQu
J/iJPJ0uiU6WtslgqTMnlsHfjBoTPTKW+++IKI5MJCqdO2pO1uKsxjmBu8owGfkO1xvFFbVQH7Uy
nL6dfKcZw9nL3M/d+WnANTnWCn3Ykhxv/YFUGZ6mrcoQ/rc7Eqxi1tZ8QOFUpR+LflZRpqbbq1dl
+VR43KDUctSLgbArNoT08Vxr5F6SNKOqs2iNHfOTlC7NUdJOwNKuDMpL8KNnUVpIh5Lyqp46yUzP
/OXRTQdziVZ8m1dgJNCgk7SMW9Dvbd8Dt4QAxkUI1wXB/cS7NyBErO1zWz8PvjXdPpbJ2Q88nFns
U1H7KTM3JDNIThDTvNaP89UYbfxUGGRbdPg4dBcIE6y8xEzmVO/HqbL6Zf+bB79HSGIp9h8lLrjk
gr1mLdtBt+5uOqsJLqafhP6aYFw/sXnTteh+RhTbIxnOYb8ys/qfV0OeaU24GHNoV0lpWsC1GiLw
biovscGr+sdeXTQhQpBFGP8v88AF96n4mMHvcuj1bcfP9eDgLuDYhyyJtPIio1KIcPRdFL5tZCcL
SfGVin1eVu2ayZW+jfMZ9l2/dlP2Vhl6nRTC8rMS2vKXE7vL1DLRDR/xTS5NVxI99mmgJXZPUiWz
c+Xcv7P/Oo0PRjavVjDdDalJJF30pMep3zIWdcbX1OSMXqd3f4mUglx0YXDog85CxX1qzY49ugOn
kV70MPs+/ahWdky8Em5JxlBCNMdAONvVL45URN8bR29CsHv+Z6EDpXtUfTBSD42/Bv7YMtgKhmjr
K7Sv1lsc0tfIcfxDWoH5w2qtZQ/U/neRbsRRReVJ6Ymw6FnWp8tv/bk34MGdPgDDNu74jBap9RbN
r00qOAKYPNXI0c4dDoswRJNnme9inTLwMVNJFKQCx9prZB3WXqP95ecGwwkdwYffxFcGZWCB4f34
jp4DjrbMor3TEmCYIENcNkZdngyQTVrTFRgQEb3TARW8bldia3YV/+IKW9FbmauemWrxyNbIu5H0
xHzFZ2DKr17YFB7YZb2FcLgq796HaycUdqbwcCDFg13q77GuywP80lkGdha2Lu1SsDxZBUj568yY
i9RVSfeRTi8VRwpXFR+lPQE8CDPkgoHazWVo75gO05g/vY8X6V0R/OdUV8uDVLzT3oCx7cBer9sy
TcreIqaglIMh1ZIdz04pTOX+kIu6B6AzmMPCWSYVADofXa0MIxyDPu+bR/7T0K3XoHUDeXRZhmRY
Lvtns3BFdRBLeE2hGvewQv2Y2Bf4BQbMfjxEOvazv9h0BQIKkZzEGUCHTx40InVKijL9+QsoxlnE
UptijMVyO3Yp/7E/Ttq4/62PrB4K6866wQCXqLF/CCl+5ecTJvkmYlXhHwAKW1lF8cmcNjhKadQD
Ktf8j4AxAStalzln1L7UGdWpA1z2xhTJ3/AJfBHzb+mRzS0vhp6VAkK5uy3a07yRR1HlFRvl4H0S
rdDXawRK8KVL6Bhrf6WHFM7zx4GdjuqZHbxo+DINK3W55l2s+NhBa7GGi86SFjOEoiQ1aidp0HJo
oRRyjp6k7e1P6YBG+oKtAbWuYhF9KyRegpkhF+Mquncc7imOYoxeP2jgrQIA7+xQVQcT+R+1+TLl
TdZXfGIm3NRDgWTzA2Ol6vGf42aJxtSSwNPPXSHxuGTWhpVkYrRKnuJr931ZwYTrfsHx+FKnwyOX
u3Nf76N2oFujadO2EZyW+itOzAaPW6Bn/sUDZxp9maStMAZtpyIfQUi9x6OAuk2WCTz7UkzdfDrW
WvXynJxOwiBU4GFQWat+y1FzjOVLGtJ3wdhqf2VcXqPDHa71LGa2cJvJ/Y6BqaEkwnU1cKd/jwTf
+Na11WtXczB5S+yywhrZtVAm+x37G6E7Y1vGEGuzk0tPQC9/dBXNHmCgKZyyXD0QRnMJ35SRB5Os
6ZqjxoU74bPPuO69B4nl0ZyZBejV2TiAQLgXDWXx6/0vLuvqPYfpUj8Nmg85f74e2zQQEtwmlWSI
doe0sVPUSoY38BVGGmAEqBNNsBQmHjxo5z2PeFScUbuP2KGyITT/dPx6724JYfbRHrZukPwgfPCE
f4zv8iFI3C8a/B8jXKIC3LCaAM47XmonjuKaLvn+bGrg4+mX+yK0f7qLWNn68myajtRhFaFQvDEe
peu63qZT6A2RIaAgWJwS9Fhx+2N0QgJ81mOHE5vcZkOTeqelVyz0Pzwab5bITj6QMgV5xirOHfZ4
w8HkQicMSsLhnUwK4oB0sOQUGZ6v1Ue27QWx5UQIzDBeZ/qFcFnO/+tnRhhsUOO7Gc4qAX0uEdKv
rDyq5VrEBhlYzOnWJBMAbzd/wFY4VAJMFFBtARwwcz2rFYCL5U2d5o3RXaNUbKR2ro+LE1eYlXM0
PVifJbOutsVb1Kj7SjC0Psd/GpFWfQfLpQvXQMxSe8DbcdBNzrmVH4EDcAz5389V2Ly9sTIzSACC
4OfsObeEsmn1+vIdNv0lX09rXMEA9gui/1ac4h2eAOE4achiSt69KAMRDNJrhkGcNm2MsiCRfIzC
CKhZbwg3qynTFjv8/cUh7/B40c5ZKSLaSovu48M0AIDbZLD8gBoLO1Mjl4/eHDBw6OW5+yKRDXkQ
5I61WMBCSko1ERCq7/AhlRG+W7F0xrifLZQbD1EvS5pMZxcjXJ+yHgtGljMb/nT1ItVqlznTIpgl
0O6gO2PG6K+gj4orYfjqC8yQX2XHbf9QPuo8JVrrXSYckAUEm/Rc4debNKslT5NH72jY8aDJBoBu
H6sju05AxwT18C7HpZpudWUxbHybQxHFwLV4dCKYmzHhZw1J0SmUrcNoSXBF5JndtpjPGU9eStea
5rrBTXJDseiW/Kb6/2aYKnfBteaDuLe7ICs9lg91M8q7u8OjGjCz4fgIU/TOHxC5XtGIS+giagmc
LFQbattmybGBu45T4hsQ4Szc5YTf6BH9XZKjvhwsxdy3wDq0yGSN48sXolBS5X8NSwy8lpXQYc/+
ECe0tEo4FODVy5KKx4iRU/ebCLb0gTY4is5H9ScvzbUoSSBNGVAyettRF0jhcPYkPjr2xeUEL12a
xTpepP2aWHOjlXVhbIFmGSS1duBjK4H+i9XBSL6IIQLvaB8li2TiRjFQOnORo1C+lX6U9CT48TTa
53/ghqR/2zEXfkCqXvmCBOd+tz4rSfd0HudmlFg135nBKFkqcF/x9ng9/tnIOjk8GL+NXr3bxh/D
S/ylYkdZ9kRKs5Ix0yUgo/vuk33Xc1+9zygzr3JXwQWJOtJ0WRShuA6etzHo0rfNPwyNDUR9UUgo
kVh+51f/cHgInjg0wBiaRfSmPjj9rr10cajiyXqmb8wzz+AbEigh5+q+iKkbI6T/fS1WmP4Pq6VB
VsQ3OQyEWJxHzyS78s2Mu/fulZ5QleDRXhtgvPfAjt5KPY9JELIEe3OCdn56yjesspVR9vuBTWZe
ZQsyjRb6ojSvhI6JUcEXh++iYOcMwe8wy4YrjeIl/eNk5Cb5l5pExDH81rR6ppbTnpd4w3smUk+0
aKAp6OlGDHyypDRq/4cdEAfgUgw5rCqV6Zai7qhKHaK3FOxXYd9X5YL6IHU+6Ujx8Cgr7aaRKQIY
xGjIC4SPFFDdJdke3QEg3+s+yuSCZKN1x7IpiuAoikBUY70ksn+w8e4syTAlKKqkcZk3H/abdSID
8HQ1xGjyyfHCkuxhkOmSnZKncr25Sy1H0stD1plIyoWd8xrQkA/ZXeGLt3anXq5ZoTki1ykGmg5+
ij7qmsat0o88+o88x+8Oeb932QfwKWUrUFO3N+VcFgyztUxp4yKTPIUPZ5zR8kLhuZpWWAYSIs/M
+X+gEkc2VOFDodSIqQiX/AZ55AfnDYzKYV7EJlRP709qQvl5IXfZzRuMcHs4qu87dj+hnwbDm86a
Pab/xA2Hdp4yGo7YDLBSYVNVEpQQGn6W078tXSlQ5IjzujAjzvnKNLxE0vEmJzAnupdMre/gU8b+
8g/USFnuROtp1EoZGbjVm98hrmnK0yUFCXzBr6UTbe71gwGLXmMXVy2tuqPFThw/y+Ot/UCfVm4a
PHVEXTqH5//T2mPTuK/V6RoWAQapgP7/1kUPMQzu2cXDcbEHSRhUsDwIjdmmL0cZMDl5VrLZjfKZ
7tKR1+hLLUKQ10uFZav1gHmjskfBIo8UMumqLpQq/pTRuU8wkssHThV28xceci8+2RcVeMDRAo3z
Ygng/UVK2zxLxzCrC1D2CthaBDHDwez3KQv/PKMWRtABpL32Q0MTfHyi8z/E0UpCOd30aHALqPRb
A0/6RRYun3Lez85QOtV/eUbXrgUIvRcEswN52SNJYjXqZft+U0iv1ZYLPqXsyfvIohI8Vp3I/VSk
V9T3F6iNpE70fc4DqSwk9/1bplGuNf+nlgZNcq5IhQfuWlVQPh2582PsMbwQWRCw52LgXQPt7alN
ZZZkWE3s8ZEt4uUB/X2Hy4aUfx6kzko/H9vZAzygH2GOt4gVhqPgYaleAfK7CUG4wm2FA7Obx7xx
0B/NqS+1ByU0ZsvdczkqFDtp2B6JD2Z46G1puYf3mfpExHawSJ6hOQi79g+B3OTftrG1f781x8zL
b3eW+cxonaR28kwv3XGxLYe3+ueFqVaFLfaz46EVGRcVxZDer5JxGonjuGznR6xV901hM5v5O3Gf
8y9agUT8zv2QMvV0e8RP7v4nK07elLi9iRAzqanwrQ+/H4RA9qnz+UMCXJ/nnryZHK/ao5KRVTRE
Sb6QuQVBZKBnAyKX1BlTxlrjFZyS74ktSOaMniM90AdxTn0iPGTFwEaFoaNP1h0di7wmX2NfXE1R
GpUR8oxdPY0Sv87cTdVWZi9lrTCcfGMyHje4xrJHvNxjQVFA9V7NYtbru2Z6kxJbGqAirHVOFiyj
zLKy1vy3lKSGKingZbJqMOY3B+RaeVdsXp3Je0SHM2koEoGFeGBya0Cc7YcxhkeTQlc0KWLgv1lQ
Q/ZJh/KMAP+sGQsW1kFTmo6SxG/oRYSji4Nl0Xe4PWYL+Ur1Um+azi8/U1aocvcShuj3eaU8Rjrj
E2cNCcqmXIYzU/2bIgLjzEvrH5QLYfxJBtRrR/ES81wgGySHL54ZKGxhpJtycG7hy/WYFu6oVx/o
yDo6yzor8DRDxakaSbCDu2caZyWYCVri3lV3+Nh7jaKuMTddJnZMii0l81LB7a5x/9lPyCXQmZ9W
Ts8C0r0lgy0gro0Bb4vwh5+CBY96/2H3DPDkwtxc0NbdGfV+Tox8tg3KmGl/eskqrkMjVb3kuYmC
LyyleFx1kElNf+bH3hSGLS8eXrCFTUmPFsCNuYM4nHtfPgWC7yFX4jjvoHCgTIAjbXT0b2TWPksd
Kf24PKSaLa6c0LMBdzxGjFns7e9PjLdHegjGt+fEB9W3awjPcJ5sKppReWRjZcHeYhVslXLzP1IS
rk0IGlK/MPD/g9ZXmt9/le6jlmTLqw8DpyCnBXAYjfh+VkBcBthR6Jw1zA4zkALRNC/JBQJ/AFIt
cJRlWoVWmMPL+YNSV6Es/NB6nSzvQWnVvj11Idzp1BCpstqvY4ClIuuwP9FEdUvi5hYtP1BMF6U6
+YBLhtk6MOb4UvzsigNpNr0T3xPA0dQQoFntLu6eOZoIc+XjZCQ98hbyi3tvWRXa3k96AsSp3O84
RR0rGFM6yodkvSuepUQOr6CqbRstmsQDl79cu1Iz2Mz434vbkfhkx2JclL9bTARCMGLabQ9xMTUu
EBGGZ+LgphxsGLPbtS65OLRSxuCbvQkPvoReQxNjap2G6RgeEiiuTlWJoF/6QBuSoDupQLFCiPwU
Jva5AW3UZyq9/zxB14/r2no4svfVJkE9v24H886AxPJUnI6VyD6Wu9gFVk+u7vv7eeYASvm/6+zN
gm4kD9saH9gIwgj6IZRJac+kqnHmRei8jl7IQ9QxrYm2FgAAhrXIQaiXhzkofynEeMMPSaCPIfXE
+12FGAFGpQBFO1/fx6/TICU99/PKrldum2l5IqtgYMJlvf69FnY1uTeDpCo/WaWN24FILtWIP53d
Y/q8RfYLoZ5ff+V3hs2E6ANZVwc/M6cBZSkhoaPnspitUrhx3ERSuPQjRuUlMw7o2JfP+xKX1Bps
oCNWuifq5WwFT/AlfyTuJ0SR6WU1AX3ziYsT008rj0YOXzy+qGA8MJb4aSULIBYdXTIme+SXbbD+
dUGoYLN3rayCtUFZc6iwvSoeCdR9wsmnz9EJzRgaLvFFT8Cair2RqQ+wkIchVtx34nGfvIgp+DkI
4hBpjXz3BYMrF4Nv0zfkVMLLJ2f3O25zWS2Ovb9pAYIT4yoAeiaFZun7gZFALBAJmTmfleApUey+
bgX0Am+F5wpo9ZHabbRVnBpQWPPr1RHdFL2RDFM00nVMJGAXFqLhrgPBq/cQodpqCn51D34Ubf18
4STxU9FkQEjD5tTMkYIigNER+AhYQqGmgOGwOb0mXECC7vF3M3RczXyXE2S7rB6Kq9TgMfo75Ssv
HiOw9Wcybcb3PuGzY5s4Bv5hVbEC+/BDEh1zcQhB1qz+fgx9ym/lOXtSMJoIUmdwrv/HB96Rxb29
oxyX+YBYyHRIupqonaPd5/6W7iFi/qyL9+DpPsslYZGndXOjGnbfhpO0UIYT64W+Ojd6o3p3JA3a
Sq1U1VoyeJMSaK+6lg6F0L4vtx7bXptsYZ+jNguqlhjbF7UnOJamY+jm7wRJeNX4ph2IjI6n9yC3
yAEhrSgRJG787upkuA5EMicqU8YQYB42N3ET6h1RjIC7lRJ+KLIhHDdbRGp47HAssa+i+o2yOISU
wnURwULvW6rZYio39uozaH3uIZ4yzdl2qTse15mpYH0ise3eLu+ms7eq7I5aXZi6fjZnvlHHftUA
ed7QOJijeswIeVMLsAOdBD1hgkRhe2eenkOVMubu/bLDcnUgP/vDSXIEgUUoNUNNsdJnnoSKrNG+
IVvGKBo0RuR5T4Dfk1RzAfFayp9XIBZ5uLp2JPEyDXx86o+3pYh4KS8oZOFeqRS0W1cajc+ifsRN
x0KxG+xp6FzFexg43cH5ECcfesvL5rq/rurhgQepneNYbRXLEtY4tn24I1nLeXScF4wgmctm8o2e
R1gEleuxxwBZqiVAGCfc/fGp66aXROcSVDer+lp1PtmKRrgeSyaU2QnSTnC2pimKVtbXGnw0Qn2s
GzpRlXfS6sPZZdo2AXIw7vQjzR/GgifAXlBjCclubKeCFL1XcGlr1Dt0+Vmu0+iXHs/V6VlwwAvK
apHmzPRVzxwG9b9PU6hSHLBg0609tHEor6wDdCJzEzDuvbEN2CxuoEF10GnU4X30cNLKBZEVlX+t
jd9BO/nQaUpMXiUDa3mLf4PahoYCXJR31RT3gWI4tQ5JS9Fgr0WP0kx+K3Agr8wIuN5yzWHkxnpD
deeK7AzZeUWFQLOsq0W+cpK8UmHBdquasbgpGYYa/EdLbXxbM44nYJLVz9L2UluROTqltZviKuou
RQaRIumatO5BIdoCRghJiDNJTmToG0iExkGZdI8kDx3BFJVMu8tRyn+8QDgKQ78HrIFLoGpjLa9j
picu1PhKfO9NMkdNT23Cy73uVb1OHOhvyKx1MjpSha+0c2TcDHx2+nG96l7BQy3W99aoq9EimbrY
46KYOce8oMzoZEmo1Ge161pvFpcvJGAm7YubmKE0aGwg2LVtrgntGQKByCX7hSoKX50iTdymWtlf
tdivmCYSZqTOx7cJSRNuhjz53Nky4PruV1KoA1VwzSm4WQTB4O/ucc5NRzdIs3xAm3TROyLw+mfS
A8NO1X0n04TYyYAbTNyPOpL7wzhujSR82tnLD0WCYbYme/V+NoJodvFy+t1GFgjWomTX4gM6TulH
V+QUWAwwRtopb9cQVcBsocNUnvBWKh/pxYod6QN4KjtPlx1LuXF87W6Hpxqv09O/15RNe4Wa2L+z
qaEXk10WYarHNlUizERKhLgF4Cn8yY1eZepkUfOwllN3eGBaPdcIRRtyxG1wiGTHFv9+ALBU7rPz
Yj3i13y4PyBVH24B9kULEVPuhNPrrRNKAXyiRijOJgmgvYyZsudttLPu43Dn7P42hfvUacaWq7je
h2vUfcQXh6hDxWFL8szIE/LxnNVfiEJtgdnZ9yUd4rGTE0xYiLNj9J+5XuWt1snhDta4B/h7tEov
bQO6FwGlfISvhSZNXgc+IUO57k4Xc0BtU2J2h+EAf8vleEHcP6vLV1jUzmDSjwzCPD8vWxBNb6GU
hjDX22Yj/iS60TlCA7y7C1Lr4+aAxa4dLcQHUmY1h4MCVEniedfm/rClXVujp0DWrbyV40WHsNWi
uyKME+3CIVP2AmK5sFQSGgIIkuYoJbnzXJRLPbQ0kp2rIPTH0cqw1H/9FchrkMmVGT26j8NdOk/h
vmBHvOROmqtAUXeOZUPbZ9pyNGtGhFFUbF4YhPSXpv2Km9Oui8yylSsCWo/tTCUOLz05P2dBIqBE
neHt0aYH6lboykSUhQ7QjVTsKcWDKxu7tw9EH0wPlxZhOkQC+D6K3sMl2zJ2xsOqsL5vBEh2xNs1
bdECq+9E3vjSV90vRl0OoEZ8mT1k8DVKzrFLzXY1qHIAqNMExdqXnvgvR0B7ntPrewa+HttfiISx
TTKA8sOORyWnLkM2IJxSq3I3cK67XfOp2atrtcg2zVPeXb4sL5cU6/m0hDYVj2SlbLPZKSe4YshV
9yS8kd9p3pMMLDBgDeGGhhnNPTJgfUuSuMmaG92fAwtYAbUKchCH0S1OWrInHgIuO19LsDQN9Ntw
I3Bh9G3xkIbVYOXiYqsSSWcOupI8eG4g4mwiGFxN1EJ4d+NPVezfpQcnfquImNUOii9NalWNGVy/
0E/P5HU2IQdYHB9Ec/oAxaDVwHwBqAlLm0wSKpIey+PTm1Y4lCP4G3j+SSInv8GoMlyFPVpxqrM3
REPlby7UmdxkSvn974eV3249wy39XTcehJF0L/vqpcCAJrslOEHKOQu+KDDhcCYye9ePPIVOaHNt
Avb3l80pHT50ZdSdulw9HAB7NNNIYCK7uuZFP/jLBZQKkgbd7ENwQa2ukXVLJNIBusj4XQaXAJ4O
57QXVYws/lTO9ZEin4Jqkl5TNGZ5Sn+5X64Tlu6qMH+B1iavonHv4XhiYkJKzqIh1uhOC9DBw9wm
J0J2zbcHVUCNM3G3upCz/ePxt2/2O7aP0JOGoETom9odXWJdUctrEPF4EV10Xmdk4CPy8Jqywgko
XaVQxWTjaGKufhAEgGRJf2Y/F25AQn5JlPP89qrHWnUZO83mAT7dn9ov5sbjGrSgDs7+XEIAx/3V
5z54vmbZGaFh1QcrPI9MfHml2N0MBt6W42jdjycyHvj1Vxg1aXe9+vChJJvASU5yWbHSk7kBzp68
8yMON61YyS/SqlWaBESsDOQuSpzwukHgiDTp6UPZUWyWeOEv464g7XLW71O66UogW2zOSSb84JGC
/DpsNSGWVj/Oh2CiixgAMRjm5J0mB/aSU7O6hikNSn1jpXowRb9bPBe/35hXwfsth/yumls/YiVw
FY4EKJnmjuW0q3HEfPPe6b8WUV7tHnDQL02hLWHqTu4DH3I+RKzoO7l4ALhtuJczxgy/isryDnOr
SOvRR0l40bDnznca5PeFzQXOGcaJwgv7akjrzHDtcILXBsH6CrFJQNYMSmdFjykIkxMYavZY+5ld
jTEhqlGNOLp5tqK6hEiorH6BaAOr4AkemZdgA6Vy20AlZ9+myf/7MldJEEc50uVEfOonmP21+aIm
K7tbJreyH6W9fvY4sgD9VdiXU0RzrXRqQBPsowPen5usnVXJtAmq//nBqNxq8YvRc7FBrvP4H7lz
rm8EKlZJQOpUdGlnxq9ITXIAlZzx56VtTK/YE3QlzE1xIAeurPjkMGy/MWCaJQUp6QqFPCmHlDnC
PiUM8ONk2+eMRCHtMkUrNONfJsNeBtKs4XoyjQnahn+N13JQ2kCVYENZCYhnL98Y708u4f08btnI
kNYYg72XRXwUWuRCxulQpkxR4HTE7OiHtuI/1fCGDnOG9nz2Ap7VBJiqD8mqA1plkznV7zNH4lXR
zts/0sfzKXIQIH1W5q6jiM/TYCDG6qPBjDzI3slGilzyTmja4MzvlP6TG7BerdyqlAqbSr4/aniS
utVCsjX71jW7LjnhiFlBtbm3R7aDYeU5VGTktOypYK/helzHPb5tmd+ZpHSJzmCVJsIvxv6w/X2C
VQP4SZSjg1JiOr+KkM4Wb571CI8v4QTmWPNSg9s4s1xubFqNtahBNM/ygIQ+cyHxu90c47OTGWO7
SOOjx0qfGKLB2pp8LIpt1+w8JgWCaT4avSKh+toT/PIo9WWV8ghYnFuWxnjtyMMgeSQLO5Mw20+e
Lvu1NDDz7/9u7mFm0rpfrFDtmG1ExuV6ThC3pgBZ7tGyC8py5O8CzKXEP/WYsWiHojECLeyhpNMG
jkGYB1DkaR+EDWj/CZCUPqWFkp0ggJTB0mpTz81cYeqgL1I3joZ32C6aNnWI3olK2o+6OgqHw6wT
BqpQHDVW8kWGg7RfFYHgQ9Stza1VjHGKdew3mQvvtlB+MAwpScGtMGGsZDwTEZcgkHCeSLirrg4w
5FVwV1QjA013TNbGmbrpGnsHf7HGC+zwAeCbB3E+qJRa815bAc/H/2ObF5aJ4Zg09gUqYm/DxD24
0JOb7ko6zgZRUTWHC0Owpq28RfWw75y5h5zj/v4scNeRpNl7Iwv+1THRgDic7pUceAVndT/2Lcjh
DKGxPoN1v193neb7zhL3MBIxoZ7LozYIgzqhJGL1nyD3OW9M9BVgaCrvlEm7Tb0No0sBmBvyQFWF
4SAf0aCa4AR80vCXliUnydo+xhbkl09jCEtQMSW8wetOCxboDbvTywzu21eiQYvNDfzBorRAztsG
sjsRftcsmOtlTQy0MwAwfEIHtW8gQxyk6hgFov5T4CWwKOJ6DGe/FDHHbr/6SsHPZK+Y3a2yOBp8
TG959MmiyL14IaVE43Tn+qrQp7pLi+ca42Ui4YvmJuUeF1GYK0eyxtf/pKZCQ4nr2LNr77ZoRkZV
JLpaNDlQ//muwJNev+i81fUfnbWu/BE4KASKtZooQHiAX654y4TkFxp8Ki4D10sqOh8fXxt0K/G7
ww+GbxUH+6bZnhaO7hMjCDsISfs2/tjo2WkvhOlyR/0E//7JF9Lj3LYS/vrBoK7s83PL3g5o/jfT
CnAMK2dCBzxH2Jr9yohWhLLbvjxJ2OjvQbpyCUQ1jALCYRp2xrC1WmYoeWiCnnXDJ5wdCfBwVgeO
XlJLVXZL/OAiBlmRB+SnE9GXOybViAwx+YAtgGkkrngaP4N407DkbME4YqjhtZknI2f76+aL5oZP
A1CvvcM5PORaA+i7wU53GPzRMXTBmQeJEEbH6JU9VEQvxc1y0CuPk8GiLPZVNgEj/gj0UV5sGhTV
86f2hzbCa7AuFV3hLYYNJKjAq6Wb7vJ8xNyWDHOyHOUU7sZn49kDPOOWKHumEG9NUKybp9Rtoo8b
1aNm3kfrQoPwUZmRglYiVxJ/oTbNx9+uqEc+uVO2sj5Md5AIYWm2zz+EZQXWa/Gso038n6HZsfKl
FkOetLnLROxUElQ9uTufGA7IElbPE+4n+rA8NpKQqkJxdUeE+EaRvxSV8CtGsYPv6CdA3xXcaoiE
oFVAdpbqmMyeriooyeTVXF1ii1gXA6biXPobawvwBGr9G5Yqt+dvz20qnvMAWV6n7GlbsYM7m27B
D5cjqE2KNfIgb5Xh63DbaJyJCtBAMorNQwY75fcu/IY9TYQxL6XogN3V90cvFPLSXxpo54EwLPyq
3gKlH4gWU8wjjsdOvtFPY8OaJGesYi78tlXN4mxwb1ha0o8XS1rVl6WxdQYtvF3r7g0xvrl0fOls
Z1MCtSlL/Q1U9bxIrtP7ltmT1W8kFzqqTYOjT/tTWDR7593MM3kHCBKQiFXIwTlI4cNPakwcdueE
z8JzmI4JTryzucjkIYYBVJwAEecNNaUhs2tbPpmgKsvlebXTUILEQyTKvNmhmArqhj2IFLetoimH
9RiUYdKRX0Wrmdx0t+k1U1pbw2O956o6n6YodYt1AlzC2/jXHKrlRtQuezJfzfzm/d2JEzilJn26
3FGfUjMpcXhftMk+U+LwhQsXKHz2h58qNbjtRI+0AlCt7ISun4iY/+VkfhBj1phfC4Ur2ZMx0Esx
Qy6G0cDSrepb12HpOvOQaAoq0HgUUrN788FYjmo2wLtRDvYdXeQAcuP8+kzpFJGTKDtQdYV9RPE5
kIofeP+YbMrYeg/zv/g8TePVGhXoa/d+hS0usasCHzh5k17o8xGD8DMEXcj0tuWXHT677UUHUhr/
0ql2F30oZfK2veI9zddSIrG4iKm+6f0fgKQz6DaemA/skmLgF8ZKDALh5cRehKFduQNSDFEANY9Q
Ln95ANrjk41Ot+zLBlVPKAp9PgHdmOtwHHfrTO7I2YCwKy9nFJbW67YsSTwzE9o4nLse/vQoqV+P
VjNsk6G8o7gzlO9eIsL57A8tEzK4VjMr9ZOR2B1PCRq95+NfOiorvhlLLQzR26vxHCINjNQSzkwz
mUX4/SFZO4wynPf8JiuRYgvU8KQ+kez1vGdKhVFRKOsJQJ0QylB9/aMpNLgy0/3S3o26XaPECcip
WhRyJ2UTqBbGWkTNbRT7aFTSyaUjXbjT0FqQA6vSWzmaLuXyh1WoJbzObXGI4JM29WGkMH0U7irD
zsmN/xVTtgXy00dP30BCC5pT3IikuCOSDGLHO4DvxZ5lImInn/fsRhevnkPcSXN2vBkkZWuTOyim
hDB8XB3me87eDgnnHIsVaKt8yrYt96mlxgLSsj/t5jWRpDPkYQccG9dUN+NUOiieVArTJgPscc0L
6UxzHiTv72ZiWvkhjltZa1siDIkCv85d9hKeV25xUXaVwY3nJwT9COlEc7HxxEMACJEXyujsWkUh
nYChmyI2aXrtGI5/ZVlMZexfYBTDADqFaYd+KaiTwdVUPB8uRombeDdYfSYxSTaCMC/rrVdkSw9P
mERsWB+IToFW6Pn3CLSlNQhbk5QYuvOo55tnF05FtUgmJx3UdtMMaS28raVvUUwtrIj+dRJb7gFa
ZIW6ecS1Dyh2E41CwU8WfuciNE2F5GZGD3dF88cYFHiQEwXY//cOAP5RGzg6qWkSUgBZGl9GW+H5
ALdPPuvuFJqaRGwtlj4JJuY7Pp7vTDFAJY2RPf/w5A+EcqQVU2BNEZDjgwBDwDWFSuqT3MnDiUT7
ig3cPFd7yUwgIx+9tqlCIyUMRbTWdDCWrcM0aOv5InaQABI63ckwjdBNPGFXCrQUy1LiuG2htM+t
c42jJqpnDN7S4iJJ25Mz739wPJlWVZftWzqtE7zV79bSNCiR0CMB9Y4yrnezuny+3jUVdXCYAmfa
6nkMXlnaESHIAXPHQ2lCSjScn0QBFDmMSjrZRCBECu794dJ8Z+D1qmWA2dqd/LRmZcVuuhxLg2Ik
029aXC7IRCL4yQd8G5Lbrs9HwJTkBLeCbfWxs7TLQl3VLejCNwD8GlXbuldVGrYogVfS9JK03BUY
lvBPHgSbLemWqXd7KjqyRg7igdo2BKhm+aBjiasYXm1I6Vv5K8sD8ovOd+S5j8A1MsysdINi1Hlu
7JfPslTeYJUkLbhO16AFM9eZfXo7wVmGT0V7DD6Dpmtm4F1fMpULdS0o7/H0TQKKKcFwyNgq14wB
ePVKjQqm7E9Kan97UUuw8YyhACTZKXPMj59IPo1h/pm1KZCTYJnE+sSet8DMYO6ciwVjf2J1OWCR
4zeD8Gap65sJQun3lrl8CiFQtHi9quiNCiy3vzZ+0pBt0/0UxGdXWIA2KDZEiM+7zXJcO0JqX635
P2eqjrT116kXpzfDvAGL3Y4MQ9qVZm3yTBMlIrvzAnMpeGoAji3cmLiZPVQhuZ1vR3vYItyRw0fr
aLfC1kBnbd072ETKN6RyZ0OrzdE9Z6azdEnahVr1QSSsXVedOObDAuCfSqngSPn0nF/q0aDkgctE
sgJ5WxkU4A4uHtDYUt8+Ldly/3JagP8EhQ77X+rNbGbFtF87YzD8BZx/4Mk51kaiC3JDLUrO1CUk
FF84PrgdEZ2gBaqF56/cZVfWmnHjhzd22UQ3RhlxsYmeI9FFM6LOwru3roexfkp5b76FLzoHdlEC
GkKdPFK0oHjeeszTK4BgEHWIJEJhR5L6n/j9oasW9nQI9s6g3JRjPD4aFkCXRmgOrxorA+AHVb4H
5JLCDxS1UIyxxfAqTYz67g4VecRXv+zMX9fx6cyxuqDWGjcam0jGQKs7YeuiJz9+y2uGn/YKIlfk
+qc+c2d/Gl3GqvP8gOfE4O0532l7VUs+HhJjKlpDiO9NnqB9utQ/T6kAcZS3OtqOsDdPFN/gH9wN
ia56FeQCB3svyDyjRHOmCStnCqHIrqyt9turIy6/iNyY+e5uRQnPL0F/myCNsTTXTjB/tDy+UzUR
+mNjMriWtrcSLdM7caOc74KN2SdBGIQGF9p0AMpmFEB+m7LZ5li9L+AKdcQd/heCOL6Rxfd6EbGp
POwBTo0rqro9/pAskkv0FipzuNs+41ubwC3HEdj5oa09H/B4GT1Jk1YdwMoWHFfBtOUb/Q3gzLfK
hi/s5fUMc7MJUQg9V7icWeftyf6Bw60d/OSc8K/J0nBB4sVg0l2vGzWR7PwjXXNAkSYtaBsnoTc7
DdMU97iFNtEwhUDgRLk5O5RLTJnurGxx19x+9h8kOpwZ+LwEArjzKhyN4bN1FSDnbI00gHcT3Y2G
QeQ3w5dpkxwNG6RgAePVU7IIoi+5sLm//IUrdI15s/LTewo3vtlm446FWt0rn6PZvS4g1mnPD4m7
c2FGDlElCuspE7OLIlV1i4jF+XXaBjiK7r4fqcldj1cgipM8ns9l8oiqXjHHCoB/FMqUfe9cJ/Fz
GKEczV/HKgwL8AhSzWqbF/1yTytRym0OjEuftgGcxD5WhfWCEh39L3ax/53B6FI21gW3rPyDp9FZ
V7rYkxB5RFQTSX/YyLf1uPH+5xu6O/ov4UKZLTmL20wgFwL1SAlUqIAqIa8lMXNGh+62fG+Eqx5w
EmADz2z6oWvTU9TILJWjLt5/vf/5TKSWr3CkSBAzFc++s2vSPLIDmaVmjq9uhTx2UN/EID28N6Ux
jS8aqOw0lPoD21CPgUOmIiPT3UoQCg0Iw92C1tBK9CsgTndxD8kwkI1TcK6gxJsj/VqfJHE9tK/i
z3QqNYmu2I4dGhaACnUpdVglyey8QtUjjGQkrg6hsXPqP61o5TTC22hQoKXmVFnCbIRS2DHEE8ju
U2mdh9oUXjibe7vXICRC8CTOUuXPxfiNYjpnyQuXiWYb1JGeHFQ/31v/YW16eTQ9MOGDaVP/Us3/
SydrMvjzW8EkZ7iarAJCn9Ge4gozme+eCN9igvZ2jFGxXnk4VxNaGHZgIzCh0w6lead+h/8oyhxj
3mfeKOBvL2JV1/w0OhlfloSu3IOusvmBhaoLzYiFHt0I100FJa/nGrVrFZg3qNi/XrpGd3vqyWdd
AhS3ELUE2dINJ/zsc9FhLOSGOPPVCUMwqWhuYZk+sNSs0v5ViBnkNF7/4B+EdKCzgOONfYd96RNJ
kCLXgBsL0awTwE2tYJxpaeM8dEuiAJn1lDzkNUjwAJ2peHKuigJaBgMFaFpT+fsntQHsXVS6RPUk
GT66GMX+p///lKs+qwDocVvjVVfQnhVEwlUZSoDZQzZeGe1T5RBCCpKwnzkLbMBesw4chUA9tviP
jZI6OELPiNZNpD7BPYhO/2XmPedxOT8gis08A5qZlhk/mwXBS0iqseWP6Y6wKhm+c98Ll3cdS+0G
wanQFeVOiL9Ww40a2o21wsM3j5zewMZgDZ+UHv5dxDAvVRZwq/5tZpxiFYNY+XLpHicljRcsCrHK
5wd7fB9qo5tGSGhpiAPpvhg6MQm34DrCQ05Cr1yQDFAwMsdw+4q5C25MRH6qp3KN2VJbx3H+cnUO
rGukMFZEAy/VjRSn4edIhL0rUD06b7SJZLuxsPIBuZX1L4/H58RZdUkhoh0C7F95ex3IjkVTKNqT
hTqLfVXPNyiXM/cT+J296jhtVigHFlalF3Tul41YVyZHUgg0JywLDI1+mtcPv+eE69GTb7XrkbPb
Jos6T0q3qpZrl0OpokIlea1YTJsx54vxhPzsOcb+6X19gPLjUVacPhD2wFkkyJTag/DxxuhXkpbx
OamzLB5K/yvHzmzaFL73bxWK0kw4FK+8PvVGOPsNPQsz5Zw8DtCJ2a5RkW4PAL65qKguyowq+juq
vp3ShfyHMMn8dDT7xBCgTw6frxqJhgz6qrLahqgexioUue6iwK/mN/jTjI+3s70+b2kG/UsX4zHZ
546/Y20viw6MthPeETrZIEyRQmUwwg3gnhfbjoZqitPuuh9jOzX8na0npC5i5lS0m3tLjtT+TrOX
L9SL3A5f7Nk8pnMdxtudSqfwz/VqFnA9SG24+Ws+JPTupPKDt8ZDKysjgq4fQYdqXMOAlQAJ0REx
lDS64a9f8CfiUeapVjDGRdC+5KAm7A+JjJPEpfnisZwpSNeQxsthNFAzi6/kGrf8Qe248MyCm8Dd
ph/MDRlsFOwMqG9/cexRqqSbfqn6WvIYfVZUKlFb7uEmB8xb9aYB9aXulkZL3bXmXJs9YAJ6FaR1
xnZojYYaPmkK+avXmrRWAEc9qGx2SNfmCJWdGacntntW82ziSw+Y1lF3/UjJJidEK/Mz260DReD2
9TAShaoem/7v8PkQrcNLj8ri7PxsIKlEiHunL9ZPT9dRgbX/d0P+zxIbJE3CCo987lHPHNlqU60y
hNaw1Q8vMKHv8EiAFfOEct70izeUqZewvVvchOz37hwPKfjOYvbnKMuDelhScAtatzVsAqw2xN71
/obTMfW9hoFYOMiDVFDxgadmC7XsU5Trr38bNCVgCim92woqFkMXEymxXxiIWZXyAlVk0zhMEEGL
6NTucCIZfp5l/LwldNXwBTTfZAbo4GfwhIAdsmPQaDxqLFLk/Kuez1Xc1kGLorypMOSy0hkiNLF4
6Ud/PDv0ZFhkFGRDUvZABWuj0LDzpl7nqaLFxtmDzIllVLS8ZCvdYVEFlCbR+XLHOEp4metumNir
u0ARCzd7EF3LF0A5Qb8IRSJG6q69JOcN42C599Yze2IxMoZEzqSZSZwOURetl/ryWhgxMrQhoFA0
JxQQPpgKfdd1f0i9aWnMQTfwt/dPVl8KLsBAedvf7bgAkYiaXEu0E+a5Q13XExFedcvCZrVfL0dx
V1PBOl2xgZzQELPmPJcIWRgddTAUQ42Ls8JwzZx28CNxRwFVNZqI1Dzcjk6CFjPgUy/OQiJZCFQO
Se0xv4aMv3qxuKm/14lfthOr6yAuK9DILKUuBQW5ztW/abZDyquBMdrQlYoepwRcnJqqnAgh5wx5
6eyBeYBjXCBzL6aU52DulraVPMw05kcX+uWUH7M5yDvbJvbarrrtFOcQZVsqN9RF+JJm7KyXLNf9
vlbhnvmGP0CvN8xfMbqH4WrYB3zPfQh0CoYT6K0Ll15mLOsDHYxltOv1wXjgicINbquPYd9+2o1H
enrhyikES5Zv5/WXZIwk/Gxn5UUNETmZZ+grnq0stdavGtTfW92/sOb3lLnxLAVEWmWyS0dCvflr
zsnPHf+RKSAuvB9Wc4IhXZSy5SvYkCh8M/3MS6OHQPo6hW0wdS2SO2B3DzfZ7NN0ZsBt9FFI6wkK
tuXXlXUxlReCEOODvcHfVL+3WXYqKyu1BWoA3fvFuyEaHIMmtOMghDTwhJ+6+yQery3X5+Ou/cI7
TYzjB8NH/FRFAkUnInKvLABj+JYDXhGsPY5lYQnUQM0vF0wHxd2qAcfjCskXc0n2+ZcYdDMsQjRq
9+zj/F8qRqL2kkeBwir/mbSQXb6kfFW3JG3aNHrb0QtA1c+334tAEwJFNAwaJd0tL+11T72Y32z7
4Ut875JoSisZHjDUmuPhvuGMZuMft9t+irTI+dDqozjyEvCDEj2NEIPERas8jHReCf8mOwFLd6ZJ
3Gf09/64ZxBlMaQCGqDDVd/gcdmOcAVEi0dgdrG60A/J8kS6MNRHK/sWim8y+GrEFFNeSQvC+OVD
lds9IUbKni646a+3/wE66jgw2erU/QqTQcDODF87slqNbGwU1g8H/Yx9BXrqX9E4XP5ICUkKIb7k
uDZmKrDnXY6BjtpaLKZeNXrOtEC345VA7ph3k7Z5MxwGueVFoUZ4fBvRClB/PSewiWY/eipccmyO
VLQrej2DnEGKm7p0LvG3J7YzBwJ7sslZdgRnsSVXFFwtlQOlLghig8qW3oYPelSBnLCHlrJrnekj
2QtpQ7fhWDGJU8SNNEbyvx50ZVfpG2zJ6zr6iMDA/IIs7UI4s5Vcl8/sg4QzjgHYmBNPtfbvmHDm
t0hggUddtxSztfuCZcZ4YBHL+601w8iVvJvdL/DyxwtpLcKJf57bORxcZAWem19lZT0O0H/SAfYV
67Ixs2FyvJQlTOQI6/ef583/Dyde88L3uEuYfjBPEZyFgQJAJ/ZLh/zjjqdlTrxKditfto5Rr5tr
AceCVSxy2mWpWYcO5nC2S4OFLyRwM0PL/GTkLu+efkKkQdmPVVyMQLne59A+8KlDHhTLuHVgd+i9
ehEclgJIWiiSwhGPwevc5nzkg3NmDtQ/iEqux/HmBfaUTYIZ9mhXrDNHbw2AbnLxnkyM5NpvxvPV
1rXMVW8PXyJn3vbjZ7mHt69F2wBozKgwIqcAH/e+4n7yME2bkNopv+MJgoYrnmDQ6prmMoqxPgCr
M58hT/Gfv3+z9Yk9lJuqmYfcEwGt0qexzdcIt5PZP3fRqnh7gcF7uHh0lntfB7JWxtMjdXGwOqKm
jKUs030SHzAd9TqeHIwotg0ZCpifcUQMVfqP/pgBG42ylxvB1fznRiZmrmVXL1SueMuRa8TBZlEa
UZgBKKzfzPl/AKh7HkJkXBlZ3FoUL8PjgnqodxaXtmTZqlz8JtVQzp+HdUPvk4vnZCrqrCphXVyd
h71OTqHxdGL7zV0jmDFe8Ssm2gBH2wCuqQN91OFTmhoaI7+4rB5Av8CW0E0lUEr075+1fpJnq5B7
VBSytJnQBb2x6CwAOGi+1v6otTn+y/NiA2I7BQoTCc3FHpx4DbOhjJ7M8YbzCokvGvb90EnNKQVG
+ODAveWpJ9npTT1u9EMslfFI9O+B1XryhsVDkwJXRRZZB4OVd9xx1nyicHbKh7Lhi8g/pERXm6C0
kyqMpswged5lVn56mFi6rTA+nkbjh4JCfb1jORwVYMYe6/IZVoYRafoB70OhdHQMouArF896Ck8E
VeY41+kfiIddc7GSH8D2LqFor42anqGtGWhOxEgRlbraeujBP04ptCog+DSLCDnrpQKkwbrWTSvt
CPjrnIuJJ0K3lcbJxl2RCScJDjOAPLjH7FMg79Ye02rc9ijfhG8KUS9LYLN9iS1AuKiC1lTtuOJ4
77L4YqGXonSNmSUun7xgGNtWndffvryvZwYdqK5qDaK/x+8L7/PdT6InV2lBIhk2L8DeMNnN+Yum
kIQVgbo83yXWImqKAHPa4N6dfENukRqe+JSa8vIddCzmAvKeThM4TMqu8TrQIF7PqMkuvkoojhVJ
l1iSTKGI4IjW2Q0dZDOjQ6XVb7/Cm5JdGgCbEzTCaQaGFXo97EwlZcKWMmoHd9Xf2CGGU7RfbB0C
Sr/FU11baaMS9vxUT/RQRAo4q2nhBEM0Xp0O7LQ2fNvFhX6rYHNbOOcsnnZA3Vns99R3pujRvd4S
tD6Bsmz3EFUji3Izn7zqHMHsL8JwnNZeiPBqlG4dghmBhM44IioHFDq/Rp9aCUT0TyIxagTN5+zZ
wEcwDBdburFzj2C8jSsIli103JdxofpGso46eFLNOhmpUOzGuK9yjicODQkzcZeyyF5cRckRchuC
HKq5ArsphRv6jUMrYu5saCez8DcOKWJCbuejsimCiekNyy5k4Y0fJcYfp4NKaHp7H32HhdkgC0vL
7XNzNYxMUFO3meAAMU0xBRRq55xyfp3wKl2Mg7WvCFY0+/9G8u/YFw/Pmh1PznwEcu59CX2j6Tk/
fT2D+cTciJNhrXoswoJxs4dKqpDr6v5zLP1ygZhEtkCLh4dadY/CYNnDEKddy8aXjiYpCbc83eJ2
qxKwuPwv+oBbf+DphVM/ZgPSRiijL8TBruxkmZCiun8dkV3Y8ooLvlZ4COiU/UNW4Rccrrznxkqb
5xIrAPxOQINCA1UE3fLlsCW0qjVItoCytwNLEeToWvLX/pfLuk9rzNEUVvAkXo7+AC/oP/DcJ8Vj
P7ixvz9khmhR5/y/ZeczFOZvidK1vDXieKxlBAXfIhpUXoPrz4P4yT3peTlE/Z8FPsYnqzZ0iCiC
AZP1jdv3popHEMN1rdjQfhYAbw+o0P011/iZuwjQdDc2vb1DllALnKPxDt3NHsyJ1jaWxBAg1UYf
OL9sNuhpqondjq5Oc2Kq2o+3Cek9SG8yZmrot7EsLif/2cy/48/smwgIwVOiFSXtAIF/HebGEbYI
cgsB1y95P1ioEdXh5CRoRymrrE+sF/nHGQiJ2yLZUt4fyQChAKy2w/RzRy/qXvAwrlV6nQG/FiyA
Lhiou+MCPLW5BnnXO3mq+zsQJjdEYQqyMg4lO40pJgnKzBJY4UPqn4zQPsTeAyG0LW5LVvksVzFA
0i3aMTuP1/D5WKz1wlYOLfYvnz5Fj7TdWZJJxSjehNhSaZ4uKJ62VCZWuM+7RRuJ1NdhTf0sKtIx
Ifw0JDBbV31+h16A0H2tLJciy396Rch6xirPpSCjalVwrnSizQgPg0olc+UuntS0r1qnvutiSNdP
Rp10kp33/cBLKWckbAz+JbgsFm5gH7eKSds/9jhI1IFOh1tfSQhYEWKX6jxYXLeJrIHBu2I+OHhb
c+KRchb2FC5foapgeUt9rrbgaiGI8L+nsAfZnwd1S8FZMq+DBsSERLibpyqaF43sX0qfMoeI21J2
D9ONfsPHGo891OMqDY5fE+9vqeh5RETN1UMfP8mnDPd8JY8s5zJa2v59tMIxGWS3ufD94mtOmkh4
WHTBtkiM9o/vzOtR/v5se1zpp+huZ87rg1AV37kJoA1uXpzi4pim0/xqPLbKXHCOjsreTGiEpTyK
UzwyyzjOIrMKQAPNnmAo8g1w5vsgXXugrdSVcHaLhj+dR0hk3l6+rt1mJRj409hR0o/GZ39GgcgQ
ElZFFPQGYg8jbXQ0xPZM1g5szH9UJMW22/HFcQe1zlPN6h3s4ZAXaKGOoB5NxPmEMvXo7RZGkJFk
ZRH86Io2o7mZ+IOS8sFt1MFBWH6hSc6ht+KvJe3hk6r2ZzRwio/AC5oi1zNvse1b7qyH1NfnnSYB
2vzNMS6SK+DhQA6YpOA9XvWwVMimhGOS0aUPYgsqS9KncfxKw8etPk6EUSXdyv9honkE0z4o4WIB
1ZmeaVnXVdc/l4tumAjcw+WEOyiMvYeK0oPLzHFmMdb3yT41bg8O8WlWN1JDGhdjX6EFtqNPbVbE
Tp7BJrLsSxz5ep5OgSttE+Qjm2T/H9NF266ybxDz6gMSKW8hZXg+ouW/L+V8jQCDhnjiSkh1HHr6
rZKJinT/cRPYzjJ3GwRSgYtuUh8LajwtbOfmcMtDcCRlPQ1PeZvsxukzb0LgeD3ugHvsv/ncb3Y7
oB21lmnzTzWDrfDUmgUMjr+FcyE7QlwND8pcPRBoiYbG8GWWFF6cCpFs1j7aiUXxE+ZN82zNj8IM
IYYFoNdFt/iugzfvYY2GS5C27oc43V2b5ORwvONKVQd6YFQ8zbVn6aNmDUOrAFYcepd9nQpX++Ae
mslV9eDuMxgh/KC2OnC4wM+QyxwgCAZ9G7taqLr6bhakA2GoJ+23CGF2AiqFU54bcTYLB1YBJGFO
D1u164c4OMcf4jlW8YSw51kpMAcKdr4jsmR60EuqN2jC3jvrwItRabdGWv+0RhcwEQbZ/r7V7REM
DhLJBv0z4VVsj2YvFwiH20FL/1peqT7GO56nMNrzRoBEe4nvVdY2eA/+pwwEXx/xaHx9pLDqKY7O
VUZm7Z09Zoowp7fOfr3DjOlAYGAmBEV7Q+WAkdaZWje/0n8nKOH6/2kM64dyUiNHSExhfZTSMB2m
kQ1AtNrQWemKXqWw79jATt9zbItLP00hAPGt+8ZAtEM9aDsS++m9WNgUVCEk6M9QHqzERpfUw1n9
MtB2dXvybPZeOMjwxsVoSxpqQTc9WtGQ64JAj3TIWY2GLgKzT8TlSjTdBSgwl85a9mH4fzomEIHJ
FM1S8/ucxL9xBC/JCvlWf9kvnm+LkRKsA8NmvocOchDMpLBJU7LeTVBnm6stQkikGInI1YfCWB4S
qLKO8bFJLy/zla8vxZAts6J1jdD1MLGnSlkfEMMs0x86D3Or7zgi5lT420w8cg8mI1dM/ep5uazh
fM8LYYd8m2ymn6H9eTVrA1zp0VnoMROATs4/c/TbHM70vDQAFIuYPbaR0h3IQg2PZiIEQ1mUCD2Y
OS8WGMB6XHCa2n+IOuXwXtDaec45CBPqVeJMBKHkUJkq9gcPsJ0r14A0J88G50ZQNeQYgtI77SPk
iwvwo/0im4Q1sHdCe5soUH/m7cO672Rd8np3705Z2MS8Xis7T1EC3OUF+katm27Q0p5f0Jkmcs5N
6592FfmokbVZv+R7DauSSui9j68/+aKDJM/OYxkNmad6uFiULGbLaorCfPVHSX/lsFUp2Kc4kjQy
wmA4AwmqmbAF/Lzn3amGA26FLdScMafqJ+PQgDA4e9fgSh4OHlMlAy8uS/BBiCvxnvjbz/6DGlRW
pJhXUEOTXeXv1H8TogvaT3NkBr+cakp/YmmJVM2urGof5j+1YNedU/iTvrXfYq+sl3Y/jfIhfsuq
veXa5QJaV2nKpMltdT+Zp+cC8i6ozKfTyvAPWK9i1bRd5GNSjezDFsRCtcmdpZvk0/6c5RqKbeBU
JsSb8Kaw5YnwqGGJ6zv64BlyC4N4dNC+1h7BguQ+GP12xuHJQ72dTW6K/0LzV45pY1YE/JE9HPY0
3EJ+u8dMdJcxVTQZ1/fxKCiHuv5ekfPMUv1V/IdMxRjDa5fXgtwPHXyf9VlZT2zda4v2tiQpHHwk
yR8Q1F4ithpQEbs8+e9553t9ti5x44X2PZ6/jg2giVsgB4n7SFOfWJ9i9Sddsa6R5N4HFQIsj89V
X88d5CVq9coHCceK+lgt/8w5txwvfEDC66I3VE8juzcxse7Sd/6VzkBN/a2l0umGWfUv/7EOX5Fn
TyMtlmZjOoXBNhU9zl8HHvKXiB/nylqY3gZPF6AXW/ezUR5YA52/7yrW/s0o0kBxy4bmu0zEfn8+
7W1Xwxv/enuyo+400cf5TiJchNFvYxaY48WZaYn+MSN11lkgBwGnk3CPdeNItuHzJwcLzOtoxQ+D
9BJ0QHKT0UvTcKpQnEJcog0l8kykjvBguuQCOkhNHRmdpnx/KzRrXCCRZQXdTNh7OPw9gRy5TJqJ
dV+/UqghkIdNIaWCbIW9I6ZYhB3+TDWC/dSqD+i0Y/57Cub5x05qUUOR+aGNZRkfAQq9OlvGQsnB
fiywV3ZNwAF3GvrMZS3SfbVGr12KyHrT5qJvHRc/bmaMfgbgFZgq2204iPRqYFNQPZVo3AEHctUW
62ncxlyhM8npA2GKvryTmQIOFZpKgb2btM8Nd81jFFk7BFhfnykWrt1Vhiu5KLHKOXyJiEdYb6MC
qYr3ldw+jfRUhq3R+pyksvvwfL/WC6A/n+lMwa06JPNPwp529mUXLJpY3BWvMQXct0K2FbT3R0sA
dWTF+TxQbtjFMLAcMX8EY5GE7j2YhFUTXeA15yPcqkszs2zbpeRd9lzAgjwr28tGMTgkwXvu3G74
yw5vCMrv/uYyYU1qPs9sIZ9yzkNILWRlUjXe4jbzNwCPOB2PVmHuxmWYM2EJdVT02r1z39jtXKip
gMQ56CG5Aav+vr+X7vz9gNpke3ZvsBl8FieQJD4KOSId/7drnjVQ8h4R9GLSwbqvVXe161eheLXU
qCh+SOfBKJR0fBs+n6Jky/vovCw/h51PwehrFyK1sySWHkRGfYoLX9PBSld1Gq8HjlFMIiv13viS
G7yCqCCfM77LDO1cycajj70Jkei7GKTvjxHQ9dGyYFU0KkoeAqBXclRvvAQRBlL2O9PLm3Vn8LrQ
q4C0BHNEDGI2wvgdd3H5aOjCa8VKZldGHJHQeiALcmonxskP0U+4WK4mMDhEJbM4ND7DrOb1vfcV
UGL4hTW0ZzB7OpqfzazEZU9gjz6i3PHD0yAdVGPHOVG73zAu24MlN4RDueyk070HezXxQoCXj0in
I7KwYrv6cmprk6vUck/VTzFGei1Onv+KlCJmwfnNUzj9LvnX/jzSOOKGbT4CipQW2OpOqAjiMCPm
aWX5ifJU4JIYZ63NQzCewU3fQcvsJFQNzuz/AzA4O/x1ZO9/6zjhOTpRNEyfnYGzAgqTM9M68Jg9
l2D4VbQgVHJe/UJo8CAx3i0sp7W4cj34XzMXAxI14Xim93Omo7dNYz5Udh0mKiw6rfqoc5vDU0c0
NLZwsNwMy7C4omdqExq7TaHbNWPhlUYaL1KLBFgHThGgMio0krI966iqKxRHX4A5wWdh9dDOgNAu
e9rcC7eQxO7D/ojos+Xwm1Ewz2YixyC7tAgZ0ymgmgBqulLQILKdtJVRQD0C8cU1iwJWb3eUdNKO
l/Oj6cr2JEgZqKtzxCeoo8ijQ5JELmk8cEMBE4U4Ee+a2QCqK8X9GDkVXQo/hItEb4FcGAFMukui
EGtKmRiJnG0/2C8DsLXRR7O5F0srWF+GQNd8CCXAU7eubNHaWUA7XCi7j3lN5OnmEnruaNEudFvA
VF1wR/7YOd3cBeT20qZ0aO6zbiP0htEiipdEUUafhZ8mIkcJWCksqprWgJyEQfVP7Qs5Z7vDb9bP
jopTnwJsZEEovsTT/dJ6AbRZEofS4s25ZD66hBer97EqplV8EGHALLBVzaQUjyYuQ37n/JnxZI6D
rPETLfw9UO4y/yzYVxk0j9I07b6enGEaMWxOBReUeYpP/vmm8Yu4JEFHhDkhIXsFNIqJogYDCpZQ
yWwoh7wQ/sBI9jO0UhrzKinSNihNZiEj47JsA0gjpyXK4KbFNczLLJtCuzK9gIbtGpTxYyQBvl1H
YBmcdglEn0m6wQuPdIBCtkxFn8pqBfHsU/y7rg0rUhLWfzKJ9EBAidB/8/Xed16kW1yfBul9cglq
QkJKu0xZg/x4lb8QXPWFU9ePgDC8LTl0TrDMj17/vKIAXpWO6sGY9F3AqT1N7+vZzi+8ExQzkOMd
mlQ3Znb4r+bMVjitZ51CWrRCnHZzLU5AhaW4rcA93g59KHn9LP4TbhI5dPGM5lN2N5cfEmcc5O0K
CpuA2bpCbu6IhGhwGj+oczg+yQMvIUnhG7bNNaoeQZSQZbJhzuPRMq1Rt1Ezj18yeo0GmNvMGDDh
aHjjgbLeXYi1hzUqRCd9Bjo+AgnuDQ9utEhOIYOwAwfTb3lZMKRtyPFLlrUnpAtxacn841ER3FYn
MYDV+jFqNiUmz6oswtcxUPkRuMoyBp3JQLikTTrei7FR+AmUXhFN6Kykzi48mhrRyzeGxBKnopPV
ZPnxPiK1K2U9nCspcIFvL9H2Bs6bnrNQjLbx2O7DWY3n8EvYTZ/4Hn276T0z+WLrsom1wLrmVkWx
AZT++N8TeO1VLKVGS7J7sVYa3QlGKtsb9kIQiZSohtXFumN2LrAnevC51MsYg2rX0LI02kNa77k0
NQtJSXegEnbpXQ2cz3DUPCBk7hBlT5Pkf85qslZe3elktjdqXvPrEZqJIRkICGuVZW2Eh46lYq24
Q9k/txycu6gfzQgGUk6uJ9WN1B8BLqsr45kii1s0LIRcFehsvik7QQPEP3CftUFwGO6v25QlQnt5
uEKjtHOpW49ThfvVAK5ZU60utaNNkC6FW0/LvgQtIDtLgYu6O9eDpJxWvPCdaSWe1St9Schd/3pa
XKuoJiAiT0t2S921JZizczZ+16uL1Boh4WdPvuAPGhpk9p7pftLU6x1wpQkwZ/CE8ZEz7kpuSR3v
qvsasNugOqQ6FRnenaVpb+A9ZgANbBMT2xRLK9YMwIgmhzcAhhnvoVbnH2QrAD0p+Dvgcojw6DXR
kXzrYYYTw45dNCLOAw1XVTSCYPumIKruwfJRVA4rdMabqm4s/P223uPVz/uNn1JL0Y9Vg1bJaFMG
eS/Shx9d5VzwSqWoJKnFUl0jaKzi6H2JpHgrXFgsZvUqZgLC/tno8GBPsPgydH/Gp1lk+84Cfxp9
IXQ4Q9h2RYcN3XiqbUIWwYk2Ed1PWAKJ2ZTdSyZih94qqE5KHestYIqKByHecFa+zoPEqYlwe2f+
CgcfNZu6DNuPa5I1Zmu2NYDU+sByUGCGozQuJNBkt5Sy9+tFIde9SNMbZED0HhsSHIya5C1/Tyxk
SZwUYWDhM4HhGNmO3mimlOPxqVvHm26VBWP3pTRrpuhVAHTzzoujlZrGS90FhAekDtkheyhwktAc
gETyaTq7SlwZRHj2qHqpoDoBVUayV/r+t+qaiQ5yA3myB4GicQxFO4px+i0sYzvUUyvaMxeMjpCm
BNaAe0ac4F8aNdA2ebDgYIzTMxxfQgZsZNY57Jy0jjf8W9uw1btochXdWnTcs+dvuOFjXp0EpoZm
3yZ0cK4re7ydmXehzVglSmNYi0ZoKGtCTki1C4SH9N1PkCCfpvOuk/Dl6dH37+1xIMMJaZ7NRgDN
h+1A3FbnqwMLkfzSWv7PnKhkXUcViIouSKBNnxS2cH0c0y3Nt2AOAxCbD9c6/a2uUhTWhhdLXLt3
keI0Sgl6c+yMyiBJ8Ko+AO38qLowTlahEmb0ls2nyITKtwNXhPhPol3QfDgbShrq+TahljyPabN5
x20Us+EK3PgGLZK/mwfsfNG/1r/NnduHk6b+++refDglervd3JGfM6SAX8Wt9Zib1vO8NwzWke3g
0h7P37HENcfqpA8CYBK+KplsQlj0k31xKDcKa+poI6mG6QI8xndy8cFPz7QR65c/XNv8g8VdH04x
lSArJGRsFvfU87SMjSS3daUWDmThjvc4psU1KmZ0t++gYezS1CCoMZxscjzuGwlsOmawNCjmQDOY
yfZj8cpaAFJaYu6sNTpw+M2LGh1i65qvlPEFeoiE/q7u/c605VAnf5jR7rCXsnYz+A6kaUp3y12l
vvtACJfMAUYsGmZCMq1XxMxyH1f4PJCzi4exXXkNYPTNyeQ69oskO/2kiIrXpM3QKMDeJ8LQor70
clGpzHN82jDFgLVtNLL3EsMrFh1nXSfDoT3zrn7nQ/9Z75Z+F55o2FRQ+XDRzvPgp4dIXnGF0wC5
pQFIom9lHsqAPQW1jc3pTQcjB4bXyJ2MaeMyKTafW1Y2RUJtgWXpC6Qi+4qpS6+jbE7QR//6p8n9
OrvktqXABMcxgo3ZU4YRUS+4avkgH+bFweEo408EIzPewbNUUyzE/tNxCveHz/lZC41drHGgyjym
8OJyCEfWKoxJJx2bKz9v5YFTQisqemu5uwXwjEQ0L8cqoMXFKalK2j1RaLKRzHd6cTcNym6bb6DE
gV6Rf0CyK8j3Jf6NjRnn2kOHa1hjToAXG3OktrBiNdXfQ+o15456oZyOxDKEH3KLOjfkN9FulEqB
3YfflgeVZkJvEQbkT6/2xJPbAQv93KEqv0Ajr8lcnR8NPdbXfGmmVCZ5ifjKthqT3SVEfHUm1rWq
aKPzvs2WY0pBMcNb1UK3PfIdURDa8A8zvEYkqRj9to4azZxJuO1opqkf0xwDJFVfRu1gdjUYldP+
GH3Jv8fon1jmzrCr2QbK7JweyYERFyPUuv0U5tw00NFkmjmGTdJ6rl1GMwzEBjdQ4GuH2M8JsqmS
tOtG0f88JN9dk9H1yC3MVOeH+UHKqLLlQJMJa/OL0M7yBCqwZbmIMR5pRnUNFht9wEEgq8Hplmy3
KF5+Iijmg3GWoTpRpA6/P9sHB7gIvAaj0LuWtGhRgbjxXlstlhhdb8XrRrjwOn6CtNJ2n4iirmU1
FWA7aqedG2la/CV0bYSD5NgvSKo0GILXnfDcKpYlKz46FwKXGUd4Pa3WVO+DZssqyXTk3LuXfylc
eDEH1j+7G9wXiIECKb+hicdjvg8UhpQIblR+0r6gRzbp35GdybVpzGu6fA+Mmbm/fnR/wCAQjrQU
2LcEElK9J8gqcPFJV046zBIEiLVv+lLm9+ALfpe8lS7e8pptg7bbAHNirXWXttPRdph63pxRZ4VI
DTtGxzQiYZdFAITfOq3Yyby8QLNQ1unrntw5dDCILMqjZDAmWa+AZl8tOno2sw/TXe3smc+8pROM
YuAjjBWMu9FpH828quBdjP0LMfwuOznXpULbM2INBa11Gwn4X9tQCt+cTDU1h39/+xs2qBKo4Shb
Ue4FptB37sJ3Ga+rLFO5lbR7B200JJXSAWhPB/QmLIEhH+pZBYnjoTZtEuu65h/RBDL1csXOqh8/
+Z5L/WLb3Td3S6gzgP5srgF96grMmtZ55m+vUPF5+m+84Z6L6D3HdsooCcUDsgez14MoQGt6rilP
/y431VRUt5v8wI9I6vb0JHGeid9SNqdUZWJYD1a6tgXu93bzjsrS6FT0ankacU/dFzuPMzKnTrKb
KbPJwCC7qdBzdkri6uvE19KBWfW7TR/tUV+yuOWL3lfFQEgKb6F5OOCyb59bK3Zv/LPGIVoLzLYb
t0X73IsnFOOIY+lUEVRZH1TRWYHILyyqCyWBzfla3SbBSvzqaA5J9jyOC5HZlckgve7jte8OLQsy
ZcbC1oaEWYoUqRDlT8ZYlkLh+b6uXEqSSlFqbGSOVl8M2OxwR1UEbiojx6BHtTbNBb/kfMU0VD/B
wV5EyiEdrzRDKDEmZpyCYGAnGRoQ1s8z6ibU34lp1QrQWCk8Dl2auoQFw59uU6zh88f+lWzuVCoe
mp7+14mS9SFmjvgLzoRubmwDabpwKaCRa+GJyHhAa9/zTsqYtT5BGe2nleBQJgbZ5WJEDzPW2ztx
jqFVsngodCeeAl4TBYne+4APndstGiad6iYvDD1kYASTCcYpYeEnfNjn82abiAavIfN7uRr/pt8a
SCTPfSLZWkPabc9YSCY1AtOdzw1JDqL/rn3v0Leha3SBpiGFcrbwnDWK+ZyTZLYdC/o/vXlKnbCF
00VC+rPC4CSjMOmdoU7Jlr1oB7t7aCVH5XR1ngFoi/0UKNizfDJepkL+MI0wDicQrvOezfI/VcSh
NigTRXqY0BSqF0Qrt7LEm9cuH+EN+qhoRd3YdP0tLn1dFhPe3/MbZ0qIuqfrMKCYafwDSNm7xKEr
nmznVlbOqdewrHOafdGr/fBaQHWDm/qDnzhPfjvtG7dNgQLv/eaO3fWmtlnMs7xzpp3ZGdzkl5vS
jcNSCJgPzX0m+hpUo87Kp5Az/Ku3S/S9qIIB/RypQcJu0UAoq5aF6E6oMtknd7wusMyNgvfLMK4+
1tXwiUT/m426oOBZ0GsJyUI0ReSrNH5SlEt8AAJQPgKR0PANuZmjYyYyTX6wYvcPN+wuTIovD5hS
/8xJ8EE/fI9i8ooqN7eOWW13LpIYVwcHjjtLm2OOgR+dQsj6C6aK6haxPqMhV3fE0fn2BCGCWEPP
bBhKwBgVxmXMf7AX/GXiSUPftMEnpWWLp7Q0hjJrKp8XE+0czEzSDn7DNP7EdZrocwdpfpVLY3Vm
2mnkShaH7Cr8B+JEw00H44BRsvr0piYiPsVscBM3BXJaUoO6OssJOUGcGnpYZoh6TEN/4WLgCHy+
WctUr/7RN+nnhIF1XOn6GSj4X0F8NsmxcpKAcR0rb51Bnh+ohGXqM4N6kgHLYqY9V87xa9kf+7E/
8E2IXTimXc4ksze+hGLmPgvt98Lp5snSUV1ECZeXE42WpZgUfBp/eDcdPNno5f6iQSHEf6UM9aC0
RhhwObCvkTVYQ+uCDjFQ4+RzAdrMT0bF42JC3qcFzR7C2kz4YHrIELkMiM9CDN/53aqopaJDDpE6
C0NARcOxJ7kK5lmz2z1iRwQrorw/am6oHINg2i3055esYwvROkylbcO5xZ55yzVw84wfEcvfwjdN
MXcagGH1D5jue88igF0bwAUyFGzVZn6FTmKc9YA4KeOCmSWCEls5hZX3NJkVKSuYfKx/Mvr31qWg
7A+mt9ad0D22wNsElf2DWsCOgDETE8+Eu588fN3M7g7SZYDu21p9n84hy3t1L+/NT3m2ioAWmrOW
RBaLkem0WQoOliDRQgFupq4uNcOoumSU5NRkLy+2ldR0RNYVo5KhgBRQbHvhQ7NaSkoT2MpJOhPC
e/kI5GnKPpBNuyw0s+kMx8ccW73dIiDWoqKc4JUz9F5f40WwMk0LaCXo9jo8Fhs8AUPXBqTCa6hP
BPz05E7EhIOapbxYGUwa/uPOtjnBnfsIBFoR5TLKCc/EfvjW8vcotRGLaGkLnjVO1nMJlAhNjzrf
UqKO75FRIxvkD9cKUCO+3Zqnw9hxCKTw/J6J9OKgrzWZ8yxdYIRkyxZOIFndXRNkrwXWRrmHn0T6
kPm5XZ/f1y/S1hbOZl9BD2UGjTmROYNZJG3lNFoD76M5Jia4rUADTuXlcacveqPq286Aq3bAyrvV
fbBjRRaCaKwyycYFVPQlMVuIF26ITHvwjFGSmTSRk9dQRetjNs+4rIupeYncfMwwmIbQSDM+5gPg
AaNIk0sqFbzsxsw8V4fIuBA1L3sBKEBdOBc4JuVPT1qGeaeXNpQCryCOCa9x1jlFeiG8xsIJsqJ/
wf6ZrROoNaW3R+Si5LqoWTR07+31aqEyxleGZOWu0YlyV1lNNhmnxXpE4p0XlLiToUi1AFBbIo4p
Rx+LSJ9y3/z+HUECb3GjM7EiKuuIDpCN1Rp2geod8CKz3rg39r3mQdMUcFNvLFsMUyKihgdkxfLo
rq/J4JJEPjun+H0eI7WNU68v/y022ohPyb4kFWUpMI9Kckbf859a/28oZ/yxsK40cIZusbo84Q6Y
iUdSz4LKmYtboOwRQ9D7VCcvYCMdl11oUYNywF+r1Dwkm5yZaUfroQtl+rfk6G7B7Y7nMVnHup6p
LsM+cdN9mAnfuVW+F+v62Bm6ZFiFGbRs0Iapzk+Ju/x3z9k8vAvePDWNh/LV5UeejvBwTUjNlzHv
i4LggjeSRk8Emi8vDO5rOWEobMSUvBMI3Dt55eE+AYp/A7U22ev2acflSbWTA8nkacp2By9MXm35
++W89mLmximclyLA1gbntn39uPQf52qMqrZ7MbY1cscXYmPS1fIf7OJGvL8qi4S+++FtYunLE6I9
5KJpzjXGFP/B+uSpvAGdr2zGJrriWVap8deAkPJQgvl9hMnbl47IG5qMrAZFqGVlIfmsl5iB7ZaF
QB64vQdEVtSB0GFlCIHIYqdNTEOn2IDsE/xSsk/HI4zhLIGxdnXtPoRz02J0gq0ZEQrDIK5eD1hL
YKjqq4QMP2Um9BpIfzoSoSaOJ3HHqW+Z1yDdYkIOvr0cBlwbJvXeICiW99fR3sKivx7dtFJbhuqs
obPJQITUcBUNTNiv746FJlbk2FLPMjQjwkzyVXg+aj6f/YVVLiRpUWz8lJI3Gz1hq3d74bXDtmom
m0oijGbk7CRwetB3YgCc/8lFVULZTKfKOyTTMu3Pox4cig3N1URRvlHySZ8dGKpQ1+UXJZjQIY8N
Exjocw3N5VViTZPWgC76jDpmgEZUEJHnTzLcsekLQ166OQ83QuZrIE8PcU5cRowlWqU2klnLIuOn
C9JQFJTFbtF4EMSmDGJ8IxSXriV2U30omzgOXV2vtuFOjx+702oFvDvmx1pBmsv6mMHx3nJdFsjX
76u0YDfgobJPz7jIRzAD3vi5Fh599hkmCKaHp4dic4nt385jZPGqKbySSB90YZ5iOVNHUvCLq23Z
RJ/Bv+8Xzneii79jRh2DWVmQEfWFgeNv/HxSMP6gXyAD527xITx29cg2kmZdVRqFnq8QQOxpD6pY
0jyIt0SMdLXfDDfjDYKM1ERPOfIuEh1CgKc6kQ3Th7Oog3ZY+4aRP5yrgKJ1XC4zGzFjJEEczYnf
dSH+AmY/laTSni7JBiFEoERAuw5hI3AaeXZ4zgJQNgVeeRHXblkxWd0B1HVE1/xrbKL2ON3WvyDJ
vPzeWaCi7O1purNv6a4SQxeBB3QEusgNNcPHO3de3z/vgetYoRKLa53/oFEYgCmNqZ2k3An71Qyn
B/pDvfTrjWunB2KEDbhk4Y6sKdV37aKpTspzkI35HMexSsMP2s7xmit4RW3X8IVjtCouY1GvnsOW
JbFM4s/MqKBCVtf19RZ/AUZWxiecidxpP36pxlsAsYjHpps9kzS/0Zxu1VS+PVh3mwt6UhVavPzZ
mvGDZeAFQsG50/cSW5h+vja6cKXQ498KIIYG+deM1wuXMl/fmTB3UlDJhzxGnEUnD5PIVec0lHEx
xqkNZrsePnCNsdjnX32wZrFKZhQe6+KaN0kN6c8x2FdBurbfUVf+BMPf7+099uE3jHq3HS3oIAfK
A3vLU28X/k9tEkHHVjrlAvmeMUpFnHt/t+qQdmlBsqjDunOCAW31OjagtrOgdd024Q1BhAKyO3u0
oTqqnFdvEILBguY2Kx0vyvAzbQo0WaYy44LN3L1Ppv25LbMR/7MOvBSB0KkH/Je2K4yFRFXSY5eW
b4cfDg6XezASiwvpapg74r1yJK0sAali/TkemiJXAQ4rLX5xp/GlqQRbe0WkAhCxo8pFqjBPdji+
lS7gLv2CAgGV9AC4FXuuaoMqSL02Pd6JPXe+PhMIVqqVVUuejpe2XEK3PqiyAkMDU/WJIiW8KKQ/
9hHKIeLdomvKBuP9PRVieqTDfeaFsAz3QWHIqOIIlv1og0UdvtTRoVNHDt5r8N7IgqgAxGfi1kWX
mrIBkuOme+rldGShUF+pV3H3osBYBHkGIaurdN+d1e9zSzRYiQiFQkVJToa/X0H/8To3vS1iZKRB
bHKv9dW+lxXpdNS0MGhv2Kb4EjSPB/Kg11iJNOg83xEo0nOgHn8HRPm1MToHySFRo0r1j9sNhhPu
1yd4eZMt/gWINQLtlZ9CgPJv/28iHabzcu4oKRErwYTQtnQq0lXG9KnOcWFTYPh+ulH6xMdOg7mG
AuoC4qKuaG/GCpSI77MNrSenWuI2O2NzorMzN59m3uCSxWUOgqn5TiVPfmTN6BSRXeQdTMWuI2zr
b2HMf0ojJ7uO8SbD9eBgrzrOBu59T9Hd3EQA0horJQByjiGw6G1OTKqeBKlZqHZ0nKf1AOH0zBhB
typ67rDZsEuBIIrXevM1c19sx88fHRZIks4JhbBEwzC/d4YOqp11QnLEFpWfViDV8ckEwSka6OnZ
sCG5eAUbXF4yckSV/kSK9he2g6xiR1D7XwT9XCKIbSJYIKJtUAoSb4tbqPQ3zheF5ylZM2G/eJyW
e1LG3qLMjpaVyJcHbz/1kpVS/bd5/6DTH0fZgTh6gim+3may/ceAVUKNQ1TwUsLjHkUxy1ADirsy
+KRkIVBH5dIOsVT3iND+MYfm1f/yav20JvS1XhoBxUZTHdcvUNF9nefbzRlKVz1H3o3OMpTi1FIX
gYRVXP5cscZzemGsdCXtmyro4FvgCdFb2/G0AdnYCSBMv9Tlrs2QOOst/piuuku4Qpqs7XNVMmF0
A9Zd/LVpA/wSSRb1KY73/x23G70wQO5Xl+BM5Y4LCehqKSLK5oUYfFVuIeoJplT5u60zHIQvpgSQ
GcnSrb4Zszoz0SwaQTPBybUrY8+4cSTpJ/DGmkFx+tFA3BkKq1jYWNCHkQQv/hHkTOXfMn7269X/
ipShfoeTvIq/sWcmAtUr3NaEzEDqDhAkUWZXtn4r4ARjd+mbLRcyPffIU5+OO5FR6WyQnx3xeSw1
Oj7EaXWgPwfRBNJGvl/wVs6uECnm2IPdDof6Y3Fa4mysgtDUvESwcO0pRFIoR3MV87X3aAcOyLRy
eLUzr2PbsClzMaoH7CVW59QEsBRRS3OXEkfTfoDcph2xTpouEvp+nnFnBykdCS/6DQsjmGmg3Bv0
stine3kawmDYWrErYWrLJkbb9gmH/ecbSP2tvQ1oE5/7KoXWyXUdfXWwK7tVMnG2lAX7+UzHSdwr
XC+C65pDxKDl4+sSh4yvuU91I35cYsyGoAZxDawBnUPuizaSpQiVm1CV+MrsrrAvXNfa9Ho8Zi8Q
2f3OJpT0EJKqrkdjWBWLHJFUu1dla+EAyxl9gcxt3Sn7dMuG7I6pKDlfO688xXlknNjEW4O/3QF2
+I6fcR5bt6cJ91sSCb1xT7x+HWT2HeqY7PE5bfJKP1AOPY3VuNCMiyEGoM3X7Ikr9qHcn2RTcCZc
SK3rOeT48q+f9bzC0KP4FGf6MrQG9htYGOX58scnpIfuhJTDWsG22Vl8QqyhI7LH03ioUBg+ShsE
c3CXEcwJSqRU8c8WlwsSFC9QOCxVTX0sVKf3grQKPWPmINSSdk586E8QvuyEKLKbxdrftGAtyXg6
pqt4O3GSKB6YTvGWeOnjkug1mNnKtW+34eM0Fx2IoZe0t2lbmy4j7COZ00Ng8ENf9TzJWrDQY3fa
ObEbUFMMqzj+L+4PONG3j+g73k2qy0fo/hd6CnJBk/t8hDjT159PQdD5eHVspWSUCTIJ6iYYocMU
yXT3/gWl/+NzeUV2QY26Kpx/oQYWx8c32AZcTcAFzk4XFyCB8A4eSESMkuIHg+mAx5qtaUJXUuTl
WgteT7sORbljGrV2/MctMGLO75ON43wQUFOAdaQMBSVvfZQN51sGbw5XDzl3hjFKCdbPAjaNSptf
HpfKMXZLKogFqcqmietEGgBa/zxwUK1QhYbpV54jLkeIM73CYbZs636UuiEptVoKHpgrkJ3aZOLn
9zl68b4iEVHVbMqg7Vs8AynXMp3xwS08BHktByRiLMciSKS44RMEdAOpVgW9HSCURKanIjc/BAbK
IFJjqhMk6h8PtmE8IoaNOkCh6T5tKRp0olyc6BRipZJq/ELfxnxU4I0mTiiPfiXZGfcba3J0kef2
hgURnreUkouY3zuDRq1J5CNMrhH4wFHShmi9Pr3xv2MkjDP7guk/9uK+Q+6K1DLS6IfqCjA01efI
OdJhpcmJ9daXeRq++z0DOk4h/8v0rq6B/5DuyVx2E+/anaGyNThWf59WA/olH4yDD8kybFXghWkg
KYThRm6xC9L2nB3tBMp1+1YKtQfbECAxmdeOKWFNq+6eDjx2pijsInrlPDcMhZ03X30jWO5ava9T
hIi+hXJHNU0zehpdwJWv9GB0D2ll0H5jBW6dIsIRjZsABhSUJicZbEnf9OpynnJubrW+CcWstrVF
75/Yb29bcAmIKXhHZxFKfKijj4O90K/NPD1EdVayn4dnU/sXECOb6+UAsP1zAssFuClbucgE+lzv
2EUUiVPzdqBPghjIQdFIu9d3Q76gdNydJ+7LkxGPgVAjMVdOYhJmQ8vf68L8lBl/tukp/1pFY6Ph
vr/0woNDjjHW8s+nhAho7hpIGY/rWr4jO0MvYutzNvSUfCz0D/7wquWztLN6DhSJXrtd35dcAZM2
YKbE8rRskkHWXDkZRVqkUdjoTQA3HZjlo5eyXyUsreKfV7IJfkTaj8qxfzPEfnh8ohu8mzKhERYR
n/WZnT1G0LnRc4Ko0HmJorGQg8x78rkP8hJoLR8hzZtZY2+Csexx5lB82SeLkXCzXgnQABLlLdQj
4KmtjlZUrIwjm4wKggcMUEwJhqMqQqO0AgeS69riuIGp3hDr6Ul2lHt9kHn2ULt0wR+PaymUlcEE
q3Wa+R7a7X1EKZYrIt4KjNAJigbKdljfbj6F8NoR43f74JQtQrvxrUz5FuYI0QRFqwH2aUnMAuHD
sA9GNyzgGjiDDIbQTIa1pxrfMwRTkOI33G5kiPoZl7Kb26m0uhgMIYkIVLyynHUaZxVETLqcvOwr
a2TuuTKX3BHu2XUEDCvOUsdRo4ZTTOSBeJ3LyOqcf1LkmT+GMxnU2wIhzRn4f7UnPfJlqbE4PIML
huYX5R9DdLp+HAo9anOifHT1guWVdz94He/K6rUbKtX8dTmrlDLIwULXtMoq8JgEdDHbDSzJ+O7U
o5vE0VbdJhmbp7sqhm17mhaM4nmaXxBf//qblw6TZZNT2HgriRWN8SNBvB9FZyG0xKP+zcc653s2
4XPmwq5BzDyDZGjgMgnXTKIUYnQYX2bb0M62QZvMorapf3NBuZKsEmPsJ52//31tUzsvA3yA1+Oc
Yd+WIhmCS9HcmX1ZFIIpOgEygdf/+D8lTX+ShqPb9fa42RTp2Q7DnnxEH5IXdCa8aYtCd4hHQkg6
ngRci2Qu2+fA4aZOwDOWB1u1iJLx6/CWbHT176eOnEYLHxmEpyMvKs1HIkFO1D0In2rQfIGGmR/R
O6zG6oxkNQci85unB16Y4DIYMiwbxoaRte6FQPhpT6eykiGxQ3td2j/dQG3QyA2Dwd1i+4QSCsZ9
wY+7UfWypMKuxGfBAdDOpk+eF5PaV9JBeL8GutYlTCb15Dx8vdw44tR7jd25ybu9cNwJVDWmFq1p
tnHzbpxXIZE9fpCViVPlzahsHkMBo+QOXctKXcHru8aufrZG///hM/izpFyzZQ6H82op95K2TRub
kffcmGfKUwnHcO8GD49xQHluffqxI4pdFWsthUKPZ0PzaxUGRdC4VQl6GiNEUZTaw+ePCoyuvGdg
+37jkH/amDrgFg2LUIcXSLE6+zLKSRRTLJ19tEJqfnKJQi6OdBcCzrS/4Zsmft5x6KJelqj2zM0H
S+uaGbWAfvdnPmgk3aEroLlW5ZAiv5MKriVBNNMmoPNTAtauCtNnDdHc5CQjJ9Uf6FiJ6ZSkabNX
NEEL1keTPWTN2l+tGsh8S6qDqQm9a/dEyxMy3IScRIOu6JnjGVp9QO5NOmr5HkdrEAo7CIhZ0knG
8hBy841XY3dS9e3j4V8CozF5R7iIjvbg08Aybi0ElPN0Pdk9ScYczMYYhJnB6EKFQN4J3yF064eO
LVMVoVaCBXYLPZmLC9dsmuHLTf0yHAoi80MAe1iAxvojJAzWxyANNKXfHbWehV+QPsWE+2/zc04H
HaLO2qyf/vNlhirloQHSb2I+1tmpsNzJBxJLsqFYiGUWAhY2gJbaZ3UyGHJ8TarE6UXtpTxKJztF
516VvPu5HrPgmlZDmmPDsl2H4hHEJ6Svn8n1ym9gBFgkhNY/MpG4vqtLcFspFyzV514bqmN/TCjX
fkjTv6kctvVS910s91OeP0oIaOWSYJfIh2TjJZFDD591Xq/eGfGmL4QWgZHokwV5YXz1QMelM2iH
OUDX1HtbpFBIHll4evxjO5pCZGXvbyS4aSY9WRj/BNoCGAjtTJuMQ5E7T2uYPPROqody8GQJEsNn
qxWbWtZJblv2HwG026+d4e3Fyrpj0X9XUvoo3+KQWPS1QCt+KfkZoYvjAUo+hyEW0SGF+PCefuCB
cLkJJkUbHOGyQ6OkXMTpnHpU+uxw5fF5ute0faZbbD9E1mXatFDLPOJTFZ7JNPQJgN+hCuq9fjSL
ZFtdeCe/tAZWf+XMoKPHvxMxQL5BchYfYylX1y/pCb0b4BAa28WCXE0P6eiuCmmCAHEjAJnDIw3g
X3+EsedSnv16i47byVdKPQwBZj9a+XIF1qunIpVI8uulRlrqDJ820J0usd96VT6pJZe7HefjBEbn
FTgAEHqKnNhye2yHPbOkElCgiL9TmBFI2oNhPW0uEeu3GEYmcb6ef0v2IeR7bkMaSnYbcxiL+11G
jGqedNo6KHwXqdHDGaF91itObfacr8Eu+skpVnSbX0neKdo1XISmkE/Z3pSKzFheJ3Eg/k1ZoY9K
cc5kWQ9VTzD1nBSthLcJZUbwuvBBNQsa1R2X7UESB9CoTBD6nUxR0fYVa3m5JM/uaxlC4KLaoyuC
u+MOeKYtLlrK6fMLbaGclX9pUnTw1q5eUggYxT8/7FC05JHuRx8VofhhSriByzlEtzpzlAql1Hql
3nzQa7+B5T+VsMPMgIiV7LN2gxvuCpdt/VCivPnXwMCOdwPGunVUn8amnA1Hu97yli7vAA6RL6hA
5G2wV7F4IjarJSdhlM09tR78OTD9617+eUjexQrqIg1Stlned6HUOpF2RxHOtU01eF6un3Q+S+Z2
gQxcHaRf+DjZcbjKXvlw/zmznVghf0ooFERjDIqMlHTcxe0uhJ/vsa2f5bGJz8s8y8YR59WDAEQm
LQTUIN4v+LaMmAHzoPsq+/fwjgeLUGAfBx/TTSpdZZVJ1gJ2T9tJsICddO7Miw/01xq2OdlLuGJP
5loYsUI2lKFB8+G6JWFbq3EUEoLH15eg2NQg0q6f54Zz8wgiH0neay8j5EIJz1u+hmz7bRltLGHm
KM7qN9/0xdVrydcsq+iadkAnZByLwILiLv1Lc5VnOgBF0zbyLg7z6OzMWXv9LQnir9NrOMTrhIIT
a15RbzmrOeoZ2YI216q6op+GEnfKJr8q43Rg6Dl9prLOB/UEKa18P70v6nX9L65B5RNgQsIpWZl9
gqBom5ESzJFukGcXsseH4lc3zsjI1ggb8khDhGdBBrjh9tyPNGC9PJjsYVEHCTIkrYXPJuzTzWnz
ScD+EgUx9nV8/2hIlGEXxE9ZtJtWS/E36Wkiqbln8WupakzcUW0D4Hv3B+3RzMqM2tgBTeFbLZBl
sfecEIkVpk6d5tPW7q8esCRT578GAUkHWVw5VVmk7HADbSQR8Z8bXVTiNVICjx2GK856M1J2/rpR
snIBTaC1MielTlhinyqg4ho4DAif7dtxvNoZkLPH7CtfYepYYKC697WLJcyZ7pwMIt+Yeu13hZrK
nsy5aOfQ4ijpELqYlmCFlYCJauxEzrbRaO6DUmTe5SAsU+cLahpgjxZ4I+yk0h1EDlOPgln9XxO5
MJp8hD9dTdaCF9b8WJQN9Mmwc6me8kWnLCgdjXpqHHtZdfNz6PdpvOOk2Mw9F0HRyqALQ6ZCgMZW
DUWN51dRNbrl6g9oMoS2R2PtFOz35CAOw9K2dIUi0pUOUnkUjfH2GhyHgi1uob97IxlWosVIv+jh
w577aJP0leuFA0/j9+dAOI9egeUuyCFryDH697EEa0mcbtHNGXv9g+W1HF+gU2mFtXo+0swB0ssq
1tFUJCkw1GJ3KQrXN4TjbhNbd7wQSAqzdX6iuaq7nS/WYX6KR+c/lTvY6ju9YXczrWwzcRK7qh8I
cAdyGaAIcGqtNLYeB4Po0Z0QkOHoKfzthF86nHVluImxy+Buye4jGZICWsOw2ozqlIf522V+eUSa
9DJR7LPDgKTdNf2sa8ZDhPoamrWZhD7zOZQakb7gwvXTFjxYVXDj50cj+ORats37L6yRIu6YI9gh
TMjoM0UXgJM4l8tWHgEV+Y9GSlxKSgM/NiHTTi+IvbBMjxqbz96lt0rf7uSxRcFjuNgUFnZUnl7B
Q7hw9l6aVRQeopVnZYDRONZTapbbAuGAuxYrjXqpA6mQlvE81B2iKy87qZZ/9RpvFBgIVfSyKcls
ol6JQRL7/i1pBuhZrMbdNsjPkEJ1XwvWuElx+8c3vSxy5NiqWwDOXf5uvPlIsOUfhO3Q66b8CT1Y
rC+KI+ckZrbkiIVTkmFQA7P/yFu60/tONN6E2BWXt8pPm183d2oNHzkTdy6lci/42n/ur7dy0NVF
MJWpEEH3EX0fGkP9LLExW9lZZksPFt1QJyOHIfkwuvYeGMLsfGabIKQngK6BpXQEiIGcb4e2Y2Ut
N1SbORArW5kOYXf4njI1P+ByKw3eDT5oQyvZmDtNgzpxOH8ieMjCUbuR1f6/xwn6sHmJB6duUQqS
j4GZNacGxPgDy9i5gHSa9fD8yf/HlKNGsKuWq+Cfi1yDkgl0E+UAMJrgTCDaUO3sl9LJbMhZKtIe
W0Shfmh+AH6OArRRAH+7LtUQzB0PUnJRaAylOlHrjOueZBpK41hohnzlZgwDVa51sB/OmDjJitFc
CDyhZWuGgbOUvtxrL5FQb97Igb8XTIVWAKoQwibVhvrsMz6whIJwZflo/c+z7G+M/MtSJ59oMrIi
39g3OnjDVuaFCu6/7+DLLTvaVpK6d0+SwXPJ2PdcvdStv/chi8ykaY5fyHBEqqw7FTTdSLW7QKNq
xpYZqUpA/MN+UzFVttLv6suwWOmixxF3X1ST9iWcO7PsGsjYG4ew2UY+zDJ8oLPeF9ANjzyAEL2d
0laxPquf2DF7lC26Oya3D7YCNWRUW/OQerzjPi2HBPL+WV9+VY2r0zru3dKcyPaNXqbbLVonNyIb
8fy6oxLYVoKSZ5cN51Xu97wOMMHKmYnTuz3DixHYFPivLTkrB2eWEp0HET43FO6tltJ2VxjqvEfy
c4f+GSRiQnaUMZnJjq5GEcmP/rmWzBaJM8M4uuO2BvN9jjD68rPq7TDfx1SzOnvv0D4Qu0wpbzKH
z8MJ4sCKZy9qaR74zX+g6bGkv93HrAYXSpmsc3YTM+BHfmqIEzp78GUvKX3A2CD3vMvcYX5oI/Y8
obIBv7JmUk8bNU/B7vVmNTaO+XWc1883FA1i4GxjRKrrU1kgzwX3tWUlMEbX9m6+JRf7pOojevpk
zE/ofPvSCZ8VDAoyG+Q0g4USZQJ1T1D927gzCwKtDJuw+HCOvMqUszXZVx/bm4etv84DJBGZy+wj
5Ok1TtlT66MOEnINHdd3u6Yy4+friGCHiRW+Dm1pW3u0jNNJNu1zpRBNiXHxNwiXFhvi+0bNG192
MiHSXaobC/q/K/dj+Vp4m7R/8pOoZL5tIBSpvkhkei5HsKJBHUheFGNX2j0nvm//iDxYyPOVfoW1
niBOiitPYUyid151u1gpXIg1qGgflb7dtoc3la2rkrI/tZ57HQ33S+VjpTT2jpc9fu5zYONH/4Be
qjGkTO9W7do8YBIKrJG6pKNgxceMyV+mm1CUDCUJH8Ha7oG7iIlrT+Ol4AyhLn5BfdLKbToPFDzT
sg81OCKHsVrwG2y4ft97AxQYraLoHgLDtqr8TNNjE17bZu9CXrRzPHKx8vGfo0cbmEYye1HAJjJy
CynHugQVZYgmJ/MOCgyNpSDak69ALGqYeLBMRPrMEPoYaOO4LkzZ2U6gyTli8CblQDcOcSjgXkDj
cwdn5cYZVNeygSGnvzyhNoSjjYOEnIKnKUX47AVSF1NVMWhe3IrHcM2biMaipsGe7PLYrL9k6+q4
U32KglwzCd6BLNFMQm3t1C7kDBzOfQw5l4lCerguw0WvvW1Rr6JGzN4eCAqlzIUZxBifVuLoHDJD
esB+y4p+g90o9Vv8Foi5Jkjgrxpuw1gTvGqvZpBlhxaDOAOtcezH12DmaH9qYcfsJurs2X1k9RTC
tsqn94kD8H+fp/ep8mjKBhAhLV/CfANfBVrOIzT9m7pq2tRmkQpBtq4kZ910wYZv6Z/ZSCyn+xGI
uh9fXzGpmyirNnxYwSvM0Jpb5YhhQ9b1avijP7dqrdDJN4IlRaqV4nlks7eK4FqyumTDxyXX8+S1
4cdEur9ikUNCCa5U+Z7TVqXy7ny3RZbu1NDPgzrxCnvsC4+LYCMseo4d9ro9YPpLyZE6Fn1p9DK3
ip8NfsZWoIlcNIG6gUMbgrI6fLMsqcnRKfbrGbp4UFPuz1tdLRUw/1cruhrBXGnVEvfxgoM/Oh3e
tB18Sfv7n3MwZn09a/bHkYLM5nH08FNiSnKunha/mfzDwp2Py4q9t7dNjxoNaCjWze1EkKPpErd7
ke0F1aGCHJzoRyuOxA+mG9KvgQiWp7rMzac5qCkTuAZLNeJKsL1lP+bxi4PVeFhcZkK7FIUezGK5
CwcEAoIQ8uGkoOnKpOqfXAvhpO/h0UmGEfgkwJCCashJRfvPYPHz05qdMTJEO+FhfJMVVqTTysaa
UAO9BGVngcPko9efUtaK+sjVqybygtCBz2VBJpU01pE/XKWJtoxqeaDiRxJjKDRHINWwGd8wKG7C
/DHOnEFnD46F/zOuD4AY5QLzmJq2ZFqEsSQJgcv5bCwYJZec8Iz541k2D7NeAyZft7lNDMwqTcW0
LCiKDOry9DU8Ile0URAZmWJ14PND6WMvZd01ljIbV1y3wsiIVShP4gvW8mNap3QOXtdt7XTWwgX4
sbWmaLhsILd3MLj8S+v2z/aPi1lrAT/YwQ8gX4nm6zgEAcWwORxGlP6zSK2WVc7P0HY6/6c17CK8
DrEUQ4jzDSQ/vQv45JIcPagQ2MpP6ueFZkZnVjvsZHS6OY9cnLWayAgCkOmbVACawcjeN6ta5IHC
oYBOfHOJuv0WMHU7bay4FTvF4N0MEauyFRZGcYsrbVAJNSDEj33FeeK+gRtsxVa37K2MIqCJJdFi
LGcL0NoB5qlbrgZLs8XtSVVEnv2+OQ+e4kpCEo6I3PZJcRwvv7t4APy54+PoyVJTL9sy0T4bRmui
psczgiEz74P+5gQifHf+LquRNTrgCvDP+th2uwtYL145rouZ5znKVOBN45SYPFhqb4Vz17wLFzxD
jwLpfzVPhA0zrGjCfajopuxsNhiPnvuAHTtFJHRxZcKjupqk0ZnmVy+Md5++V1tIcaboIG1ev9+y
9UlFoeZWRFOH5BwV/upfxUNaain3lpJwZaR8gu1aPcUCs/sPRYGMy8yvJJOR6seXAPbwzUlSgQYR
+/Liswl971qxkswunZJInqdLQCyTlkC6s85GUYEJUzvigIBPCcHIFkwKhcsWe7TJPF49JVyDO0XQ
ecnDwdVL7lzwDx5smjTjXnRgEBW4tb1Tkxym4BRRxJ72bXjULT5Ldv1G/2569zQvNsTnClHvQl0f
fKP5/v3jfz//yOGqFvbynYZ4Tl6jON4kRKDUYlKiUF5XGqIy0wOvIx53MhTodEk1GoQRR8ogRLWD
7PtzWCgStONMRJBlxFxbLmnwNyMwEMWDPLbDuKCaMxZ4OIGo3VQ6XUj6NMZzJ/uC4l+fbYP1HQEC
C5dLEEEeo7GXgKjWcP45BJ7ngrPNn2KJ1CSfFTs7VEPrWapxBWj49FbRx4ryJqWCKM2dHVDJc/3e
MdIaICFgDkxhq6eZRCJjmVRE0Mzmpjhjs5MYcP4ee14MI5/2i5WgSDZoNon0QtJXYKRvEmOspgrS
BzUC3HC+06a406TQeF9bgbxZhP/TOB8Xz7He+jt4z/2HAzfyctP0tgYhApiesFUcht3ddPhaEUci
u7u+hOkGX5iD9sgYNEkdkVKpfPyMb1DpjWBJbZL/FPvxNcGIT1pSxE6kHyeVsua6S6YKyM1c6RDl
o8eKhM+ByXZ1xZn8shYZwbEmSfT3nwDQF7fJi4jXrHveDadH5Juj5DEN259PqsbGC+TZQj/G5IG0
MwKzx4fS9d0CQo8PrN1QbngYktcgTFDMU5YvGpSkavfNj9m/+E6WxW26QbP1l29wagst+MsaghdR
w5CEXYMOSnhMOqmNTeqNyXr3lC1/31JkQ912wPpPMwnEuG2UhlQlSorYfp2gWYZ3QPzyaJ34Mwll
amdYX7Xa1yAyTD7IshIHTG2jGx6IT11MSTXduaHhql5ne4smaGQTLLv0GUdlZEcVplGR1kupA1Ry
8ZohTOxnBOYld7n6TVAUr6JXbX7wQCTzJ8P/UcNLnAbXCfav9SxWJN5XDOvqrv4Ffl4jm6Apyvie
zPEYerm+gYcd4LAWOGzPns/+ZF3G6C2fDwWyiEYqbJb4c5j90uHaSton0Vgqd7E23TAebhG8/c+e
NZZRb4sMq2rN0e+bGcDltwl6UXTHbmpk+ci/W1pkF/9vxQJD8DuOI0JU4lQxAYGy3zXAaTMvtvn0
TX6YVetXlKok2aB54cDeh4qT/FciuMMd20Ox7KY/I7jVCXLMJK4reCuotILAstyS72Ag5RN/XxHW
TLQcpMIPkeIL3dmqW5o87mo76sKIacLZs0sfvEtcpeGhNEtoQ3W4EFVfAP7Y77RJriw0ZEvW6Oon
sgfC33wPesmIjv3IZNiKGeM4yUOmH0i6V8rJAxoWAWUDJ3aUmOywl36RASlWIkQgrjyMPGq6WUOf
8Z0u4fG9UtuyXCOLTyBYxZPd6Mfzm0hD9EkdO5P1vqAIAEV5dfHlJA4jv+xuWjZL+hfauY1m1j0T
E/KOqZjMPWwBdTOD2UqmS9+de3cA7Q2KeWhspWpa4lDaMrK9hn8kkFdfZTdq5IayJr44PNNoy1XK
Q/fj5KqXkqm0lCBSLxjlDNfgJ3I1QdoW+Qz1kQJo/NhrAIdRbXcKMm+W8MKgn9lxzvhA/zZT2VV6
EoJBi0eLznyquAirMV1UhY197UTJ7mBc5QXl8/Af5qGI05YZC6we1oFZG4n+0Ol7ENXAiow8MCHg
G57bUIpMHaQqlIup/fNnegxCAX9b4pNHUGkysGMaiX3mvFi3rFcnSEflBg4gLFkE4k3gU0S9XHrU
WrnHs5xTxiJz5g7X3aoV9/GxJ1G9xa+bre64MtL6TkkbLmt+c2lJFMpTyDfnauq1VAvYNqMyvvIb
dkFk78nFaYfbadnjRhwpdFNthDeykEDmW+E0Pt7asXc+U0gIjwj8ATfER9aQ64IdQbJeqO7UA/6z
1+OFaUqbxZyozdort7Xe0y7cgapYNFiiJNk6r2MBavo5MZTDuzr5EyyTbsjaedRVTHFOVES/AUw7
S2/bmokSRMp3IrvcmsWhr6qOLDJwj6LclxQcUDLokK6eww+mOIjSXLvW0uzifg/Kp2XzxV1pmt0v
p6tLp6BjJaVfdOeixfRuAeQXgDzWom5SVeL49oq5lTbfESm3dFWkYq0Zieq6NcaiwwULQStf6ZN0
6Q4fnloVSPwpRxdbaGy+/o/lHHLfzGzOALnXeLcVLxMAc3Pu2esjOZUawLHG7EwMUhA/ig3GTyt4
pDVl2k8HLffmbka/YTqJYIxGlQZqcn5pXunglkkqGghdLguQGQCY49F5T4MoiHV2cY5iUPH7NNo1
Vec+lnzjB1kXYwmgRaYFk41OBTKq+VRJNbGjepJ3NPx7wEOva4JMzkusxao23D0qPZoOTeJuJiVh
qfg8pvzfpwl2J7BWks+91lE8s9b4FMkJai22odp00SkDCR6b+xM+gWcstdriIAkQHFQR3c9qfwlp
lIqhcirS8e8jqR8+dgdYk8hi/ROhd19gU3ToHomCasziDjF9R2tn+gJzL4m+Qm0o2GFC5ZuUa0iB
ahqL0dyAI7KnIQYFCTPutRO428ALd3EcfLAk2sjnyy6GrWFqkHBd+kxgZ3nxjMgycJg7Qpn/mgvf
CW8BN9GVrRByF+3aPKqX2gS0HJ39YP5favSlpnAroTrLMtY/Q9piJSj++8fJgYfY0Dqxb32TQN7y
5dFdxxNGMHKkudkMAQo8dE6eSn3Zr0CwbrWMUkPqo8dQMBZV01DFnrkPfZJSP6etLz8Jn2zK/rE9
19V8MPrbtjwrVmJKSsl8PluMmkyR6aApA55DyDKuY55xRWKtgUE24in+yK2xoeX6W0lPLEKIt+H2
5RxeUHfgaZcgxfsUv6aqZ7HHFHdpcNL4Cfq4dnNZlqiDpQ6v/H13nSnuD9YtMgCgwvakBzXQth2h
+iDUkYwZrRFcRMommHqEdspKA22D3eRU9sd6CQwFIpBJefb/tb3YV0laOXYq59SRJofLkK8J+G5i
vHS7KD0lEIcZKitTAgYU8mZ3WxYXTuC2FORmIWWpsKJrVHkFtOAI154OfUk4AjbKLYT3gAISSovO
LshELkCberderWJINW782x7lFl2mYutO5dSeEFpxM9D5lZIXWT/LAH1AbEjOJmEOhhx8ns1JmDEV
fp6kbBdSZRAsoSYdFULXRPUX8bh1IDcsWK0qDJ3od87AA4jvkqS8acOzhEdaZ5XygWSfl750Ca+H
ABL4XpMlbZlFa2Lm+LEETbV/b7flyoznQZirQXEWh/S2DxmX8z+nwq/kVkUnYXkt42XcodZ04S5c
NIjU86c0rQQvwod43ZLesx8BGO1tAkpL6a91b7LT2D/4ZI53VW5KLn31g79NSOeVWBc2mdG73vAW
ge2dpMvM/PSjWlGYXrhr/wqppILAOzix0mEyd8v2YS4F9kjh/7C/cicta4peZJzfi54GxLwePLae
neCcVv778STuAfvqCknjKo2i6CWnDXnlN/ZqMGVbWuiRL6B2cWOhSd/Y2K48ALKqRDRDWALNwot8
TVFLM9zniE26kGGtQd9iQBTTe6PLO4HxMUSrCeikXDUPwp9IWuafhkYGmWQ6r9NC0/n+pg4prgHu
wBlFM0t6gJ87/aegGWynvUF3SXr6jY/5G9AHMZlaFzYlLv+jSjyxnSzFdqsIPpNqCUYR8hioOlpm
xgG1Ikqg7D66s3mnGWPe60ncE/7E9adfsUUBOdZBnbcTc13M4VI5GilRw+9VYq5c6b6qRWdeRarX
rjNl899KvTCBOlRovsl1DlcVPShBRIpMdM39EL4wZ2X8Me1YrO4TQsNQJdWvezxtn++XLZ+viZb8
+e0+2cYYrZxgMf65qfVNRQZkT7xcKPeGeEOobATTTwUattFDFXbfSe+Z/hMZx8O7MZHJquhI6Gro
d7smOe9J7RjrUVTufy2hH4bTcFGzQQ1Eemm7d4fqmIu7rWlLOnfNcJH0Ej5C2gdg8jFtDfn3ALt4
xBEjRue28z1O+G/ESIDhrCvETMDWuK2kzFzBysTMwSxaKlv+7WYVyo91rIBBDVusiid/OSfq1kH9
6jRhj9JzY3Avr/o3Phnv9MyvZbm96/zg0NmcNOEiJnr1HWnbKYcsDPM7Z9vL+erdVu8u3ge+H/UI
OxnRE2m8FqqUIo1DPF8t7ra1TMySn4kTrIE2AVxLfm6DiLUWIMQqlZh+9ofHViQnx/L0AkETXkpv
tieL/MJHqlnjPY0lFLaZWjrnZs2kzHNON6ZRcgHtrd79O8OSOpC9ZOU9l6ihO7gRas8OrqewJJyV
T9dRCSiPaiqO3we2KlmHU0F/LF0ikdSNY+/Xbt2PGui8QgcImVHOFlOJLaI0DtPqwok8q0gA0VhA
dru+X/QMqqdBBVAcqxtOH5WtjLgGUf6R7urOOQc6+kVc5e97AEt/zAtLn1du5Hw/Q3c0J6JPYFzf
ctNDmQGtUbp3GaNpDhZI9mDyp3VxWuQ4HerdGjCoSqZoUqZH05mWfVwMRJ2ADGysSFOPEDFlAtA4
CTQQzzGX/6Mh2r4FvkkFi93hke4PwDtzqsHcnzLGZzOgMTCJpuDprpva5ibLoE4VvzwpNToRbSXe
KBnIpWR0qt132Srwe0v3hp84udas+33BLSisTaC+YUbXe3P5HMFcj2Q6LslGhXFqww008Y7pvh/X
u4W1GPmx2YaRq/Gach4j8AYyLSsqeh3DyTnx7i8v4rTmvwQ6QRkvwYe2Xz+jeDn2eSWxbUpqoNV1
7XElROWBesUJnXgCgOvs0ldj6Q+JCaqOB8tFiOj4PjFY+C1f+UIX60M88CUZ6ESYfzyIQJgk0aZy
nqTOcvFZH1yOr0WtmF2+UH4I0+lIq6GgrHSKjPB8PgAYMABspitD39N4k2PNWbDRCywsMATBnBLv
NgRzN86lGLnKs2q3eEi726kexIi5FWOna1H4xTvJIr72f+BwPkIL+MwZsEocLdWrCR0KhtARHPyy
SE17IXINkKcAhBc4f2NU+Igosd9Sz6AL9lfEIW2bnrnHAn9R4ABVV2tTh/6oKgLKRtJBPPda6WM1
DGaJ97yz5lOt1YEjblKZnZUrJhqTUCfjHzYILOv9Nffr/EnQQfGWn5yI3R99k9kvS9sN3nrG5jfH
qJ7MaV5ruCjoUBc5Z7u+aM9xYKroGfQdwQ11n7YuLQaax6LHY4uojZb71T4QzJb3TN5aN/5Q9YfC
+E3NkA1VRmAHxYD4oA7CsVc5GRK4zF2qPa6uPpwKT8FoeuDwU1Vrlsa2NYmuNKK+BaYIVytUwI29
yylfmsgnAcEFvGCNI6L0C6+/mpTZvZu875qYiI92sMLARpETV9gl5jNgVwsHO00xo/HwvOW2OUob
9SI5CuV0GhzQBx3QXybKno9fXkvKAinYXxqGA7pG1ks5tV0Q7N/Cz+hM/ISRGrhBxZqHvXd3H4C5
/MbESCC2A58FQJpuMOTqBSsYa4IfEMxDQh3/5bT9sywIkGj6pfpbnviH5JQcjUOUCelbVsjNgTS1
mvfH4z4O57kXtg7qRdA4/eRhe/6nMuS+ykWv0j2gMRyYKvMneCCF4/z+KZ26pvupcBpIyoiHsAC/
e9qskeojkIh76s5Wfm95itSookwQyW7CYUl/jJlS3MC1a06YxObwewK/mweHf9lgXYzJyR+o9IAH
flytCHKd5Uttne6MCX0WavLljmo0jHcsB/fkYvkZwlmtK0VUJtvdP7SkbJtKCpX9X1q2lEkV5iMe
r6KhOqsoUJ2CCoWv4aDS5fH7I9XojhqAH+MxhFq+9U50sa34HR9hptw8FHHzPUQKYwwt2rm8z5m4
C36nqoHrZ2+bXIad+95rVBPW+veab+qZt3j9qRL9f4M7N5y8ZCwA9/37vxuMBzO2EskEN4NAuu2n
vbMoRDJuQHYbdpCZm998gzMxF58cM7NKjJFIg6YLZZtlVlPxIZd5Mhhx/dw4vJCA8uGvq+JHjR2m
M+Rk1Ju1oGHbY47KdyJsnbo4iomMwDky8PRBfDdANJ4eSz/PuMn8235ZqdpQwvjkqFAu/N50jOYO
FF/K//CwDdhtn46lbAkmctVjextbCi+9D2qhPQzHtNlrLrYBeQVcjy04YJHUzCd0V8ZfU+i+f19L
PD2V7wS5FqO/7FvBhWltZg8xhSeRTs8AOzQsd2zLj1fJmiPondoFvrfB9Sg6dob4uGdI8sQi/6OD
fJ6rHTZ1t1JemDVvqyyh+qO40/jd75czQdwT8Va6/u2InR9SNaLoRAcefeYLUsK+4ARUYVMqvkpj
RBUo938WFkjDpn2SQNEFF5daCWQXE+2HH8tuWzxgprQkCwxbvb/QPm4uq2+A/ZoHOmA6cRdLZa3u
HnMZK62TSZjqLFtI07MN4RWxnGTq9SwNUdSqPOZDSPJmRZg3j/56tNTjxk57fqi+kybeSmczRvA3
2wRBhrigLvAuJQWO6QepSCTxeIFbY64zsr3kVZj2mvRiQuvbvAeOiUY3BPhe9rG0svwiKNEkWCEy
/gMRPgGaNf6/LABW5M0W/DrCdKuoz1yDDj56hJA+A59MF8Uez4efeU8uoAGkiavgyPYXQsYcOv1O
ZukW79Icm8szuoauKY2/kf/ESeySXyN8AwJjYQq9EAfXVjWob/Of6MgMdQ8JSSZ6+t2DjCYt/UZi
J6xVIDkLS2/mGy/B5f4kCXAd/cdqTNYWbQd/Z1iFHQo5lNuCNkvNSWw/7sjYFgXVmLi0IqEAzThe
CHP0fwRGBB+ny2nn2KooCNMjQdGJK658vmKK/8c7p6fbRKqQGAq7gL9NYr1r2F2Mib8j1LafVlzI
5a9u4jSGNNk28TV06pKDZLJk16NI+GqLhGzWPevl7a/uRTCiqSTUkskNY940DFGgyv9acZDazswh
rjRs5WRDPHBjahOyS0rOcn8roOb4Dj2EVdynsdwnX1X67MSwgF8QpmFfYddDU6WA/wKwXt9ovMvW
3jxYGgSyWf93CTwoTwatRXKW+mVduiQlYAHrBwcYCZF+33gA4/i+MmAJWh2nDzVjRlanc7V34A8B
THjqycvPd8qAhS9B/Kp+iHv0wjhkGltmtx0a9bf6qQp+Upnnk9DYzneq3sUVDOvFJV0nlJcVC669
+wzLZ4v0hx1fNHT72Jms0N7vCsmsg+R3oFyCWzP3EqCTu+N1shAyV97huUWa8GFKiH3U9CidYki3
ua6HFBKEXp5BkLrE5aMcA/URJTKuli4wtlDAlH3B6/aU9eZvy2r7TCMaghfPN83V3RI6WQ2ZW3Hu
R34lOZwM0uSmYCOE/IRveG7BPm3U5J72V2xImrjl3TRBLsw0QuIoBY3rlOd2mRK/md37DJaOnwO1
qZI3Q01uq/C+mVdwaqSZSn2+pr1FgHJ61eHRMTRJW3gywOUGpR0RJYh/JhHUNo6WFubeos+OIFBq
nwDWFqqQf1Jl3uNtWvnm3rdY7tDc9Zr8c+slc7BAADkxWhZIus/JIf9tG5U6mhO06oSoI0LKN8JQ
8mXSD7C35NqszYfzJfDTq6royrOQrqyTGpryq48MNJDYAr+EUe4JRYAJjaXOznx34DSogxTj/JxP
JPW2KrassGmaIIpQH1nA/O9LKgJNiSN4rqlebBrX8sHGT26L0Q5pubF3/L2xRKrMJXtn3uhO5uzC
mdIA+xZ8x1VMUVJN58eKpM3AHCMpaTTazOjAYrc9l3WThmh/bOt7GMENKuntWSGlBApsPZUOyfxm
wufk1QA7yh5Y61wcecPIAEkcw8rcHFItCDHbo1sxChC2ZDjTDkeiK0V423QeRe5ALhf2ImYz9MWc
J8Im8JR3rkt6jXRGJXDo8YuBVrca8utHOA6BNl5CQuLh8VCp+mtjWER0ulqXxDwFER3RRxRQGayd
Hp+5dnT8q6cjR2JM6hKtHXKMN3upJuz3MVptR3JJMX8C7JH6SoGhWgdccKqKDlFCtyzRM6NmBQm6
eG9VMD2rKMpOzwuM3RmqncDZI1xO+Lrl1dhMenscbS+6c+frL97RkJg18GEjXsStAZ/HLumLuI40
0LMC/WSyIrHT5Bz8q5AedqyPcGD+nCTy0Avt1fAGxYUR97VANgy/MD3rM0reFJ/n9Va9Tplfsg0S
eu1/1mbxdRNpbRiednZz4/VXlbcC4acaG7Y9lE9aHwwqcz2cnmjgXdis2C66kP2jq3s2rQlJZdEQ
55MYy3WGyfNQQ27/XP/Sw5lvhy/VpalzIcVgU/eu/65BvD6im26We3WyPab+sZGI2/L2veISgKeN
Rd9qzMVZ+NGw3bw6+w6GiB72lHwXms93m2BWTQFASVI6Ci7UVibDJ2cVq+9mc91QyTvNlvyT9Cw2
KbrRBpHZLl4GRjMRpk5BloXIjJ+jojNaPVMQmPhOH6/7PtiI66anhYQEut9LqEX5O9iYH1KSfB0d
RWmKtINkZmgg/gyDZK/wcx+fImEv3UJu8zoKlEK4TzC2ZhDihbEkwDWf+ZNx6mfdWF6CGOLffbok
Tx5nKmlpLkrYNE6DW/oTwJ6ZUpf1YFBC+a8FQLWJTNgFe3z6VCXUYVNVeZbN0o1JD3Gth626wFmq
n/MB02NU172zN8UiMStuqyXAujmdrGygCb133yk0RKzvbNSUhNb3LUQR8HQjH99jpv0DnuNpTT+o
guRLHI0X2E2N8rQfjDXLFIUQCVEyASaJRsWcLPxA3/6zXS6ysh9GDVFYYwFSYMzFN3xuxAcPZrBv
o1f7vCHkeSoo9XXsbWxs7bXeJFrEajKqtZSMCJrMVMM9LLFKkhLNkx6c92DzuB5Z15fKprlcUas1
HAqphrP1PLNHjJ6JV49napjK0PFSQRXEUwR0JfzypNtuRikanaMlmXlunnmDJzpEMrdyoCM7WPbq
Z8PEkwcy015bHBU86Zi1hHW77DJ6yA/itCZf1Thu3abizsWHx9s2fj93e6fHEEiegixilpgB0Atl
FVpkymarypqrqy8vBM/4uadnOf7UZ/gCUo/+nZk9w49zJ2EIFRdjMwgKoVCZ0EBMCLqkZG0rUjP3
8ywuMfkx5fUWrU1dOtV98mR10aE8ThCI4WaSlsT35LPZ3KJC+fjUo+GyMykvcg8myrD2zbK55GXL
h+oGO0xUJfjPmieZU6jKcq1F5rOfnLEiLrs39eycFqKqaLDx4PMLZjuXEQBSDpYwz8np6s/Ml5pi
YwGssqCcMa/lIxA7zyWnk4J5rRYgmWf8UtNfxhnyqWn5ZYHM2gn4OnFtBTFjHLuaPAGhLEOWCgXL
etyZuzpY1b3jS475lq3r7j22xXt8ri2Fq6OfS8cSCnnri6/KBwVyKMWvoqQnEJjkVqGHQSyY+K7T
0ezdItqZ8vYGccooJ1YJje7sEnzzzCBq75lOScIQUdcM7TH0YS+6Cn9OQB4Nm3HcBVXZ7XL9jHgQ
8VtgRMDM+4kXoVjb/lJVQIG3vmFnaRl5ACv2iDbJWuRUhAzcKpgsPWybe8J8se+8p+KCvQ9kU32i
iEcLloDCbLtJqtbFwfs4OqgN5/IzPapzblKH/0SVkcDFd0NVLlF1mmD8+8gNcK4IvEChJAh5+hnc
hVBKymabCvBJqnZXTTpvWeHCP4MmQam196OsSpOHYpwf9Evtqdq9SB7cUOZY2vgXTHvXwj5o2eYy
5QP+GEjwIJdU51u5wyfE7V8mBwyOmWBcx1cK/3tgWfucqd6kmjZeXvglPctMZAXF8SfL7caJbU60
oPtMShGegF57QUQF52OL0O84tioBMXab2mar6aQES9Laq7mEIk5ri4MSkFLuz8rKx5ys8RSKzvyz
b7jvBvjevPvwCFmigOKg2JAKtu/jekZs/1uSJ+JRRRpLaRPwSJz4EQZ7IWOeGWURff5Lhe6tx81Y
nzk64Vf9QhTYc4YqxvWRyZFyDWOBpe1epAODzIeRyye7URHgEk2/1YSJbOd3RFwJz/KWtzEBpwlD
R+nPL6SGavfo2M6hy0gXM28axtIwUfqWGAUepVEXDz7U3yqB8r/XbgF+Pub+HMqlH2j5p1+Q2OtT
JnzNRNr+2T9jSwbu1gjdmgm2rVMtJM0H6Tg2/jacb5SaBFY4Gc7kpFIaeETZ+I5g+KLQB0gKTcKS
2r9Uxd01f862qKv8rxYx5qSDn4KV+2ZaBAb51ExnDxo7bTkohO7UX8WH+4jraXXRqwdvVfd1vsRW
7+Vr2nsPOKyrqP5faoDmIQAN/QsgDqjgnl+WlKEYJuvpjHnInHF5W2zAOV0sst0/lRbyGZghatJk
TaKOjhzPdVIdLlrLOZ1fCfGWpnB40VOWo+Cx6iAnVT6qAuUn+YZ1ZawQTa+l/nnKWJagNCJhIv4Q
XbVf/3P+Y42McBheR6s6BUl8pz3qe8sDQQnNQGzmKn1Q+fcpH398vYs2dEMdILLNMqb5BT6VVEg5
UJbVS3pvV3qgfFtBkfvD3OXe6XhlnewQu66oY2ccl6oQJpvfVw/VnKODvQwr5MpW/yWnepSiDXjO
BqIHRI6Q4uWvY688XBkUT3EH8ZwAXUcEFOJAbxACN43yD9tqgkOFNtw+tTWLuUn/oI5pVa72wWS2
YpDCRaXs8aDRZ149ukhx5kf6hDm6+06mmGec7e8IUlUaHVfdlAd9AcKDvuVwKld5xnXhnrtOj8d+
/GjhoPvwbWIaikiMsVpKja75Osm9bBwphDywv0eKVktTjRq2akZidUBqU4Z5XBU/4upkx8KXJD6O
aC16LoAATPXWGaYJsgzr2i0BZaOcSNaXvlFI0IUKXLv5ku1xe+o2tacdHRLBRVRc0FpdzeDji89F
AP5ZNzxtWUsQ4E/ipp6xQp5q8oR0XnA4JMoVLs2qahElNB5RbYjuWsx6sEMnRQeVp/ye09m8Y1pe
O4NNwIAX34NJcgJmcsEt+NPUMzd0DRqYpyWMVyO/UJ9UeY07RnLcbvqMcooAgpxgUmPSLj/dpdEz
Glaf1PRBoHKa3TeJR8IjWCPi7PTtfZ7a9MEHWeKExWjFBghX7flIrw9h9tDushXNap4c6Dsauax6
D/MJzYoUJ+t9ZTQXZm1ia9xt4dftqgQcZ4FVu2OgryGYiRYvcFC+/lD7C5++3GuPJsIksfmosCpY
xWHTHuC06NcfJCuDVimHsOSW5p9IXly8DqaQv7KwhztIJ76z24dyyPY7oSLyYotZewNOsK5YuTR3
cbMgYS44C4WErlABgjg+d9Y7pq9u8ftsPUxYTdiQNfyyfasLfOTHD/qMWx31NqnK6KMY9pFhvaJh
isCUVYOYeo1MpQ+xzPZ35EgNYVY1dDzMnN3RZVlpXTieEtB4QRjZeOCvnI+TVOalQXaWdE27D+Yw
9Hpp35I8FVwtzO1QkPMAJNbEv+4B6lF8CY7G3B2O45mqNGUDq3qQi0qET+36nVf0Lx1e8JL5OFF/
8Zn1YcvkWgcmb6XdzbWEag+uLErRU99jfZUxSNp4kT9GMLqFK1DKrGdOJjcBsky+qbl7FLMX1LBQ
1DZEIqMtb+SrXiah4o0ZzKdCv7TppAfbnnY3QcDmFLkH82bl9WT462Oz1kv8e5JDjRm7P8/qQ7ye
Wfb2kPZpyKz4MQUAGja3XzCwkPb2iMCwktfYeE4ZFQhwoNe+wZnReFYi7s1mx9sjKziD63H/iDpa
XNB1pep/XltOhreb45D4AxluzjXtVJvZ7GEO0r7NQ7/mJ3dyrlm0+Gxyu2Xugxt3E/uvDKLg/pcO
hcML3L6I/EF4628iRQTCZENKjDN/jmHwN4Q9LYAtd3LobkYz4FAnsgs7KF3SCHN6tIhcQU5yci0T
1xvrnWVZBGr4I4alCAoLnJeBdW+XRSj1YeKPbKmI4fthf3wf4cG+RrF8OXd7QYcIoPkvAg9ncMjF
F7Ngun75nG0X4T0Zp/6ADAjlrh9mu2VtT4gIHoWqvYxJfoTYCuHMpBwDpQBFtFZ9hcJ7jIHVGlCQ
OMxrHqElT+9tVVpI+V4fY5mgVnRXWrftR+++qSECxz6+LfcjAAWnWhe5jTZYPn0ADceFTG575KOi
/J7RyrwrJcIMIdOdhD8EfxCbZmiO+EvurMePxZREJ+W9+kycg4TQkqZtxft0jxjcjSH+Gl2PpLLx
R42WLTxUozOA5aprPt2GW/zTTvkuGGPV7PXQYvcVTry23FEshe2cYk3qoQRJqr7AWKiffVpvdNdv
VpJ+1VUodC/nPTIcleKu9U0TPxfSRuNpSbTeuRVi9KvFKGKaZF6x37cuoqO+I3tD7u7+iUuZVzBu
Y8GPdyA9ksFxZ0xQTdmnTdxyJY0ZvCm96ahHzZY9Z/ToF7kNGFpm17Fu7YitI8kZnfGPZpnpADSU
iFKD0E5fBtX7RzrZHYyRNuIfFnAJmtEiT7kPvj4j9/WguXh8DFUeOcOSWDVRlaQp9B8XzSuoO6RF
VzrvuxoqXSL5bsrlsJaeAnt4IC6kt4k6ChUYaoU31QXX5aA0e1Db6UJQMHExweBR9vS8yWBgoRIW
1DWPjtmWxYaKicmldrUPpCchEWReg8bF7PdvLmOuFI/lVTxu4GCb2Jg/39+KnKclnUuO2Qc7JepT
Xzcir/o6nMTfFKXfFEKdoyGf3rO3BUqS58rEuTiwtIM6gLNKct2dyTicLZgIARmixU5dSg09MaVk
DBF9nwWOYm99OstDw4/stmbrjgP9xIZYKMzG93iOU0cGKQ31N10RsyQ3v5rdi+8Y2Eg8wl1hAGm4
IFZyKMDqcvpMj6IPdYShhkMz4DKDFRm85g0cVVpPD76eOiR4ZzqG/J58wCOsFyqnOw9lBJV3/N9C
kqSUPK41sloJkZ/cTHhJ28YG+jRV8QCA62RKlyoScuST4K+LokQ6bw1dxraAt+jvmNdkbHH4LL6S
TmDrItL3oLLUfcIoB6mYemFJ5dmLSxNHej3mtF1BB2jPXR/mbLMCo2J568EAKR2PZ8gBa469uwwr
J4LVBf3aV5KWuXvPJN9M2IW1DfnS50CHNf4/SOKAv3o4/abyu29N6Mhg0vJxa2dUcwrJe5rI36pL
59Miys3DTIyjoPspH/TxD9A8PQNShkc7DHkuCYGDfjEIo+CTaEaPAR+tkHuCQIyhsp/hg2u15GER
uPaZQLCnOC33Nl+glNtocLuwCk1CH2xqaXUo3ZYyvzswI3KUmYfrTvNvW8j5Cm6sbZSuvf0z1CKs
MUHb8Ga5TxBbY3w94xAKvwFt5ZvJbmMAwW/A9atoZF6hsx4YvKMuXNzNAfPTzpT8dpLRdDMfajg7
1qJdYFqLRnWORLuPPbaEtIJZT16rXoUEJT2XUuPf9oQXvEfJgnbX/YQAE39d8O0PqHIb4PUNbnho
I7Wo433vVSnaofH7c6Lee8IM5LSHJpTPCJyBPoBecqhd/km/FKJJzxQDU8AQYksiWlRLsTO0AG7w
PV9IIv7RCwuezb2onzs/KMlhGz88G2bM8yzQfoLuVYASm9UwYQWNBVDs5APBAwwQ49Lm828xW274
QnV5fDUYI+59ykycIAbplmB/2CTUJ1PRVHCwed2e26HogXSscKeXx2kiwbY6Yd91iPsCQPkYS/GI
3ZfmBiQ9CJuwmiZpPc9whH9JwDWthACJC+Itrb3vzhMHYXV3V/TyHwvrsc/hBRJIVz+tHqDcOSTo
+O7f9EaAKgqCN6b6qJO0duI7Vfa8WVFhU94e7Fm21yXpICTrNXFXyDa1V6xc0n8j6tyUbW4dcpKb
lH1+TDJU3c458ZiM/stMIHHulWS/ZH3GVzChA/8sfcglnk34Hpg6uE9I1Y7YwlQQAx8w0duuLcpo
HIndBlxBOE8SR5YTY/uXf4/Twh2c7rt1k4exDv2CohoLl89tuCfqLAf4Lv0azAstZpyg2yTwXFu1
HT/63Hw8pVC++6UaXn5z0JY0eyvQgmpN5w7MOU/IQUb9Cw+cwt8xCEJFHITQsuVHGse9IXcymZhw
BJMNe7RSaRvTM8xAxj/acBYsdagcTWNtK439Dsr/qLpykKB0/TdNrQFyEZrw9tTrsNY3AQNanYkQ
Y2Fgvl7PUiHmm5wunw62hhv2ZIlujbdwShXTOj27cD3SbHW8WhZ0DWWURekqD9GFa8my3qhKI6xp
6Ym6eoyUDijLKz1yUnC5AmKaBJb55eb8X65g0C42SbEQZWkvZjZo7Ndv8g5qSnkUMjAqMOo4vjZo
YunC17okFsqbC/V0z91iQbQFByAJAT8avXKGuU6sxl3AIJxODX0kCvoDQeNs4s0mXHMNt3P4Y0gn
+TeQS+T9+hU9VsebvF2LpjbA9Gzm2HJ1vWy4qm1cXdIQyuRMXCvIUwPus/n1VrtarxtSgP74ljgI
wP/208q83OYQvymQNXCIFosnWLbQj8Uc2j1nLMI/ngZTOkzAePKt1yNGYwQuw+VI0U4FVnjGgmoz
ZAJj0wWPVNhiR7jPL0WXComehbMb99J9acOrfZh+zEydkHYlFvt1Ww4pDnTtnDKdWO57F79wvbD9
lR+mjRf/BHj6S7IkhtYFDydM9wB8zYTAvHHYW2SkcjyrIeLZtDgRjVXVixa9yp2ofjGx8SPi/c6H
nhU6tHcDLJE9hc4a2qmcryIp7sgeq8cLhlFQ79ljTbpds8aEJL3XvEeJ7ZzI3Tse/xOoSMGqdjJx
f51gmbHMcJMvmcds99wxRapSthY8LmALJmffHgXFCFNj+BBh9aBnFF8OkeUcBVQr/aG/LoYJ4Xb1
9cZdP9fN+4Dzv0QanS2CvA99IU5u/TM67ub+jeix/cJZIyq0hchJG2DzOY+8GMpLzu4FID01E9+9
m19cxsRvZjqxDaJcCXD8zLD8v7i/nz2j/51ZnSRZ+xd/pz8UpX28DR/arY6yWiElNUgO91Ymm3C2
zDH6RyyxOpqz8MCn4spqMLFrfS5cz1U5wAzsrRW8qb53wHKkb1KDCd9/cM43T5oQVDkbRdUgIUvs
2jSsd4zbEHAHJlk4sFTaSgGSuuyhV/EQ1fw2PpQj0Og+FMBwRryyFsDXpfuABhoxg/axCOpep6wS
l2Ug0r5wm9g/8jkYgKSaQECq+kJ3dw9X6GrYMZtywVsvozKfLeEiQUKFCu2DayqRLSa3C3ZIr07F
yLLj7PP5PsuyK8CmViTZznLz44vJ6FZMZYxFuVIzjfMohoAvsTQEq2Mi331z9/n7xkmwQHznDJHE
GpxlZqMeNLbxQWmxmD3fUYGkauXG459osr4APEnZH9kpGYwS7AX1p34Fxopi8FOZryKDf4SRD+VD
58UDltcUio8e75/syy/Z4j9W7gfDdD+e0H0GaAlzZFfNJ/tlVlAo98qWub++GEPj7u1UQ1XkMcWJ
C+x31fEe5y/TQx+6gguOCO0h7J5aH0q/DnRzxQ1qsO2dkGJYqt3tWkD0wYIEToRyT4CU2kLLQ9Lx
OTHh3HzwP58vIxmOB82rK8lXOZlQqCnxsgVgd6PY5zWOgPIa1uYgcJk5N+0DrDWXVJsReBTogiTu
JasYiO3fCtd8dxAS5b3CTjTAsbUjGEaJCDyKFTNGo47mCbULsBE47EtSf3jI5bplTGaPXf/pbpqO
RDJooWliiNhPUZ29EW3eRc//ht45/PRBKXWHk1+ECECE1COzZkBGT5t2akAynspaeMXAqz9ZO67I
f+58JV9J8GRMJ2P7mH3DSrhig7opbiFFUbcgqIWR62PthXPKnT/llGM12AksZfTtXNzswzOrOAIG
e1waCPIi1lGtKxmyxbQk2TI09cI3cgVNIA4CIVXUjSp2zZwFrJHrx1h2231YQT5QAEIuKWamLwB7
T/qu52Iss4dBARMyixEubfykuw6ZA3gKHtQmxeL4QQHTJFT8h6WGGP8fnZdzCM2KL5bsBZN00XUZ
Iuzab0q+aCylmityu89p4RtOEbsWXs/q8Xg+nU4crrPRnglsKloRq2XcHww7T00hnpYjFU5acE64
GO89VN79mf/vGS7kccI2cpwy1ZkCIZv0LvA7eJ1WkeAHrpjdR1hFVpTib79JpQwrJbOw+7xU1jdK
zZaUTr8uNi8YqtkJmnlAafIBCax4VCxZRi7Ba+qG/tluP9yiO71HZ8hzmION+Efcm5R3c+HLi0q4
KPxEjii2TVdFifEZ/MMcckX786nMa49Nz+hrxbfjq4Q74qOAfL8Ufhqh+lOn3xzJzrVbIih0WWej
tixKiAe5L8+jkeyefdYg+nEhsKXvIG2WsPz+SSXtZdIJSieO+WzesDYu1Sa3gf6M0t2D1fhkLPxI
J3om2dj1BzEdusUZmELcinzbpBcm+uwVB8vNePdWypq5Sm5FoiA/7Xv2EObY4SHGK7xjyibfEuVt
5OaAOvsmt18tvB501ZiNbq4hPWywTuXnfiGYDgKS8B4K3SPUxoJz7K8eDdeADO6UdqJBBc/XEKqQ
0zlML93Lzaf3DvWt+UF1UAIvxl/GeF8+T4YKg1gKjhUvWX2LbuCwHr3R9DOHRJ5PYPFU4XC8Pr8p
KXEuVrOmbF0DlScC4i9q2W6Gx3gIh8xQRnVGaleTWIP1eCgKSG1PCz5Qf62A+aiILhThawvFSZKt
tZ1wZwHTiXhvKL5a8w4XSg2ludcXyaEl11Q1463Z+pmY83MhBcQ2jw1qrf54T6OboJ6NossaICTZ
Eu42Y40TGjcHPC3u3DXGePl9jGGKm4BgZiS0kM18dsnMFKxo4NPH1xm09i+RFHqv/YexEGfD25Nj
3yIJYG2tOfq25UqnQjlH8HyV38b/gdTSdDTJgRBC0Bffe3VkwMgUWceKtxWFTyjmsiu8HQ+XXxkS
CF05pvI5GWrzQ0ZHgdW7FQO8HuhLzCvb2Uo/+hLkXMvCPSyh8TOI08lweE52gvzo/1qlvkJ7E1gz
GK+BUL5kqVBFf8Cwe7brNX66NNRGuO6fUp0pB/JJn8+FJNZzF3pA6f4T1MB1uDH/UGGacndDktJU
UBwP9nYVGquwDJrObplj/OI5mNYJN2u8eXQJfKqQ/wW9GLVfo8ZDAjGbey6+1jQ06sqhQt+t6/Ul
cs4barLsOeKJ2ZYPswfr0x9Yt4FnvZ+Jzk3d63osIjkQWI2qtrbEac7cxvbbTettvJkiho1CVGPV
BLmfSy2GFU0tiJjS63bn1UgovpYKfSucldvmT8UwNXp99utj/fDP2oLzx4mC8/nGF5gD5KwpJkmv
eL8RggWH/ctmNuxY3PogEAvkH1m7bBlqBjhKxdGBB6BShLW4zpiNEkqw1+ixuBI+vcUZPW1UyzZv
RZwc4BExC5PLsBMD/SfsXkZqBQulr6cQsnLDd+PKLwEDScAeLd0Ab07KWmX5Rc6lcoKIxP0blKEV
rKN+njqi8yN7Jx/V0YwQGOiBIZNKYIr/YAxG/BnADuczI2fexXZ56j9YngyAu/zLNnmaymnaJrjx
1hKdTJkFmJvct5zo4DZIX7Td8Js2oj9fp4DeJXq/9kdiOexQnEuZsGoIpiqFmP5zNGKealilk3Iq
MbBW0MW+s65BLGlfHP/IBteMlDL63v+6ByInO1PHtlZUD+Ac0021dm0d+9AW8TIXLa9cb7WTeQjE
JdS/4XUVgJizVU7Lx7U6RFBcEGYbmV9z9K3vFY3ACOyt3IJ5vpEgBGl07mO6cvJSvcZojrhCQrHA
nJYLtxStNud1jppS7+pNypDIY0S0GvbtZtQ1ef0imirloNT8/eaDs5q1vWEwyz9YPJih0+XQM3Tt
PMfn7grKppV01V5m+Kca5G4wLmYxUNydqhyoJKNtNy+N2orSQxPQm/Wz2WWsGuf6YEpY9gXSKi9J
/K1cYkwcvuCF4RT3vyiMw6AzI5ywtSV7difHUgb6dbD/5fjZYSKWtwMe5/TEhtKwev7F4fTCeHci
r0JAJuyGq8JroCHkbrTIjSVLHkRqKjQAprZo1lc+KdyPZAhuvkMraRpkgfNkr+uOvLJuh+9WFLYc
9h3UuK86TxpS3bqK+ZtjFMZwaMxYi6TSrGp67Ri7apduW/OyzSfjiTKEd27yhKEewX8txegUo+ps
/D858rTDQJ3QQbTJmRSWJhXf8KLjUZsNLswsdk89f9CGNmVYleaU94aNHRCCWu5GXN+8JlXkfkoP
77xIk6MzdGSLJEHOyRauHUdClhG1Os13nCRDeYcgrHAcb5zABsGFTLX+hhSui1dGf2CWltmpc/sI
rQizQcxs0QSoyfZhXswXVbs8O8KA9kGYukUPck6197/KVIBUTjRw5zDDl5SNHZurGQILhlGwbuvU
xguw27+rInzClmcN/dO79hIA4lbNzQqBjCWE4XNoUtfycpIK63y5ijkY8Qdx9uNSiEnLaadcxo3J
4M+Q9vrFgmvVDV67pb9lEA2j5rQvW86cI5YR2KVUc0o4Xs0/EZqlpNToNK/s1OuN/qkHKkMEpZO6
lqvIfj0V4ZR+2gEjXxukfwIGhUg1RN/1+PHZjZynbTICbhQi00YyNLg872N790MiU6AiVVT6ytXZ
wpqy81cSY1gTYyfTRE0Pd9x9GavUxG8La/7+k3TjYmGF70qUcMvbClcHzbJ7HaXnVBgGaRsdX99m
WriCmCJNqu/KHoZ6eoXZFvO8cJX9+DrJ1kEM8GTMKWyi9lJ9gbA0aRfS9K9LiGX1FKag2DtHd4o/
dDHfId6EBSa8q2OzZduuMOyrYa1xZVIfh47CDm2BN5DiNNwPzjk/AyILTbPfGQITq9C5eeK8oSQ/
il7OYm6XlquTCAwQyfywv4NioK9Za2nLkQ7xg6vyLYvjnccuOP7EOkbHH5ZGO7o6Rb8vJzl+8vNS
2CaBGEAtYiwOtGOB+tvUlVUZKcDrEENw8WfMRD7Rar3VlEj/XpCqj27aat5oxZNdU2x02BFnoEV/
llFK3WMVaG7fEt+mwD4ypHR5pm2/9VdErOoSzyURh9gB41YfNraP6Fx+Pd0Nqo6w/fdS3QV16nlk
TOlD3GLzd9W+t+Hs0Ucru+Ke6FaFAz8pLfCEMSvAlnMHTbZBYH4eL4I77p74If+97zXGrnOVdos3
mRhMqAcwWhVtFyZLiWj1j9CB/L1dYTjvustVemj/XTJnjpNbGaVLCylnH5Jf+rLz7J2tSkCg7bLk
WMmBJRkXVpLSnGktU3DKkdwLoChv6T8nmwxV0W8XjrCvWsEl1j3hcHPjVEsQgalBxQGezgasbEyX
X56Qase+lEjrzHOqmkaGtCMMs5ByljTCFkxZ6kPXMpoDWVQ6gJRX9kHQgF2lUjzXlH/LomVRnTGi
z9UvN8ashF8Iurb9p/TvoJqUEF1J9EHWHacBD7XQfKdUU9q8Ea2Q/dxWyklRla3G6RCjDHVFtfy5
DAv70xm/djrg0BksrTFUnmqmfCC7jTqAEqTnZzE6K5bxm8WAM86zYQWZ/vle1zFqPz+RYk58iPug
A25q6O+1QCkyhG/Ubq0CA6GlEs/8Fv6yQSapGIkjc3ahGebKz4S1q5nBoUA/a5e15BfgtHSfdOrx
XWgMrETZGbwFqOqVTLUpixLUKRP/1G03O+eWqgvcJ//czOzvAPGiKq4kmlkniT2XKbBQ5HjVLFaG
ffWHo8rBsA21L5CtLmk3XH64uOtrMIORZgL58YCScTFP8ODd3ZOEQdIEhNvZ6UwpJBUku4TU8Pmy
LTc9hfqZTI63w5NUqy7X/j1bXJfj9cdFdrP8nKxCVxmLIWPQkP3McgnMOyFdD3g5pt5QbKvKqFB5
X0uiJrKv+L8WSf/Wcnl2J5Ce2zz4f1G1RQFdlRGY/Ke8tnu6nZ5WXDRFAPJU5Eudc7XZKxqAo25a
Vr+YtQyA5VMe6VVOzgBcWqBX8lU9VOdVxyos3rU2jB/gzdkrr2prB+EavAEAlj3WOAQO1LoOGQ5d
2bQz2nHG9q7DNmAT+xI5EXGgm2CZ9/tipDGhErVNteU1vrgoZeyJVH6w4jWtkjI/skIkln57y/Td
+jaA4VmU9DGrG0by+bKma/Ro9aMnYYMJ2mmEbzrs6q6DOis6Kc4XjzZbfjpzYVrBrpGlvotEvGl7
Hj8C7qSwOjoDHuOXl9uxDZSPQRMshQxWOUUoUwgQn6wHZ2LqeVd5Ph2a33wfAK7Fvcaj2sf6LSzE
LAp8KEI9CNrkZI4YkNY7k9f/gPjvqcluYmRAm7YUE8IuKXoMWJSYyFUE8vjaJQxLCcT+672Ubr5U
eTYbRyaTVVaT8xng+SOz5ixjbgy7FO7C1zmWKhEzAfFwnlHDFjD1EuQR5sola16yNp1cFayitqp6
ZojAZRnXK0p0mI5yRiM8D/rqERuVlU2VDt+ZGiEYZWza0hR/K6hoJIAlt+f3RJR/E8BsAW0S3G15
2wR1HIfzeBd9gQIg3gX85+0FLo1VsidvwuxP4tUppIzmoKfftNn4ZEFkSJZDI87n1wo70AbCiDfr
FGOS2E4ovP6OV1E1ho4lMZgvPnLrpkzjJ7YOgxG5L0TrqyCrAp67d08kgizoGurw6blyov71JOvJ
Frj2e3LaD29s88fwuDIUbGrg+JbUt/yAm1njj4pjGunPAiTCZKK6I3Esx8xKcp5cIZsD3crxZ7W4
RMLaUyIABwcUf3RR1S9hoMCn7U88b91Rf3If3abu+/sjI5raZvsxpCQHNlkIywIHV/jSZ8vjkrrq
8FfG4hDaxXpOn6VbnEE3lhfBSAwJkcz8AQxBXgdLCOM5IU0S0NJoxDutDkU3XT0jc1p1rMG2X+9m
9CXcw1b+MQn3KUc2NWGb4XMELavsSCOu9PawB+YIO2X+q01KVqjBDFEotRa/ZxhD7O/SWtin5BKI
2r9xJ4fdzaFG7AqyQoeGzfKNssXk5HUTLqHnh5eiIsVLDp//yesh8tOAe1AblOVlSXKvad/UVjms
diSYKbsD0/2hSCRpOsirMy9y89kGTRA6egqp6G9BeD4Fq4B8eTqaD3t60rnLpYFes6k8k+Is+cii
hFuiSX7z6dSU2DHwzE/EGbou3UTrZ64oHzD5/Rms1oF3o8bgXL0mv3AuvusgILJaiSKzsa122QGB
HAzEFok2f7xdHlbSTQFa9rq/Sq+r7pAX6+C4scRgdhApZ+J9ateDLZINGYswSjXdbPlKkk1F0a5E
0+Ua11Zx5QZNqEJ7u/OilBgjEYziqQTPju6JDcxsIVigBQr7qc/vM64wAr6siFxSg78T2O9W06gV
7VLcVmkV0IjwCXReqpAwV4wK8zjc97z3cOA4Qjy7Db2rnGGhppaXG3mbcxJx6nyg0i8i/0LLvUmu
EGFyZ3qUAxkbE+GCSNakkICstXT6QJh3ITsYh9ITX+OaNgnRgaUlnR0Td/JJvNOssSj9tfitpoGI
PSjoX/HWKGHPIMY3bjA0rmuBMFNGL/AYU4zPAQWAUkDlRfkQyjN4vepBK2DP3G0ApDzxmFpDYZve
lSwF9jcs6dz7WuBV3ZRZ8NwrVKQXGWUmxg3KUSTYS9ySNlkMcLsF3dIUGWMKETk7IkFlCPM4mC37
3mEIBfKvGdnfw1yRCadNtexn5SzFoOWSzDCvRM4f90sDtj/snnQgCJ3fbJK0dKgOMIkFrT985MUH
NZl8E7UNZn2CyXhYuwz78JMJiVtW6xgTSaVvc7J/mlfMeD7+iP0kxyH9pEdK726OFxTm7JBawjSX
CP1NpD0aG5R/pd8JQ17WF+EWv9cVcewxlW1bYV2ErKAUnPQbEan8eEetGQrX20TEBNjbW4yHisTj
UWAzi9jbEY13Kkzgh3ZvmeIc6uk+097GMY3F557IVWZTfFyEzImKY5pLqbEdNp5DWGCwKxOTRBgf
tohmQAd/LZzspO0m4KEk6+yyaaU11knPuqzpeDuvo6dF7ZvRgQzxJK9QIVQnqmIJZUtInrm6eLvJ
tXwKahHrrCvU66hcfdW+0Mnzl90ant+GeqC61hib68Qo+K/MAdFS1/0Vi/0EciVLN3nTR0TdA6Wj
gJ5SIlghz6fSs4oGFs326exgF7kBFU9izjK9brVm8FuBt5mCJ5fvYow0Vo/idtetNTVlqn9s8i+R
NOC1Xu479F95IvqBGJwq3+2RQAzmcaNFLami5DcPEORe8kd62a8NmekwdoGzO+A6WGoH0MSil2kb
VDJgUkg9USoeaHj3B9QyEMKEFvvnUNCfVoFLWVeKViqkOGBj7CFq7uldYnYkv/gSiSfikeCYWCoD
+1UqgL87BHMw4UEIbFzENY4GKdHu5IrT63x7DiGg6gv0NdBqUxicWHNi5pYWgWeU2xubrnOhWtlu
UFPBCOqVZ3eNkyZJneDIhKlv5kAIhrwxF0T0af/cDnLliIerG9X+u1fFvcTyjp7ak8nKU9K1zclq
r55hqplJf7OE/g6u52YgyFi8PrF5fR4dRStrUjdgeRsv22lMudsnsRjd2BhJCK3XJtQp+6uBlHxQ
Qr/47qbFKzxqG47nx8/UHzbwo+qgRNsymmpBXnJ8cXTBB/vVgcXf8WBJBRZWYFsSQjFAwpSoZbAS
Kt+pf12z98ccE+9AzfLW6O7/HvWPbGvTXa3ihIplUbZaKiqdwyBIjR9CElPHtkRzN0Mca7nJBaGK
E5N3qtnulfcAcD7UOVAamzfdo6uY5a3zGRnOCVKCCtNhIABRj593G7W2klTVuv9heGqhPTnQcyPP
LHA+tysPtoIDk25I2ew3XuZhbI2TFEGxk+qQNyl+HgwtNDA7/bXp7jatGk0K8ve44J1GpieWnAtP
fMhJXlsn0pNxdQIMaGtDYyMv18RMT0tYtGa4bJmn3olpKqOCbIa9xtfllYVqnKgORDEyAZat/9sD
WrHhhBYF6wxlqwse2g8moBqUwc5zZxfW7aQ2xkcxK2ZH+45Bs6bJjetFinlfNJ0CuOqLDIEcHLle
BYJ4TNO9x8ZTE0zQBgdsUEiYc2zNmpCbFHlF3iVcwLzaKd46vwBHNOb/tqs5h7t6TFD3ZYxgJCFm
emYy4CRvPVjr+5w8Mpsb99PM19XvLyjn30ddj8Mx+qFFO35C8lFF18jZ9/0iilwUItUFEgP2ujnK
8lwRzBih1MUr8TO40jskZP4cEwN9KJqtDbfDxC+Sa2eJDqt+rsYSw+5v8Dvas/vS/iTfxOF3s9XW
fSk7OUOLFjITZTCZifhJ5iOHzUyAml4hjyDYvNANxcJY/XgHm9+AWQiGkQbvHy71iGdUxf1MbXOf
D6S04C5PeAp3GRpXhT3ogxqtEOeXs1PCxdSVZpIVFht+wAJzBpBHoh1IIqbGB9IQnB3MBWI7lLeU
JjJaF59SgbEKqB2lCG9eiISer/v/lfh7WldppIlE+UWSMdCh2RvI+OJOxZNtB2qb+wZK6HcbUcfv
Ts1yE7i6/zBtxlNcYEi1/yeQ8VQ8OApbGXhOAarj/K1MeDWx7R65Brfossy0T+R3nr9zxZGvrc7W
rFMDJ2wUiceOheFr6zaEd2VGyiucBw34Sm9QWlqcJ79oz+XXy81aQb3xo0HT/Y3GSbawYv5q0Uh/
Y1rbenVta6E1m0ocsU2GTpy3CVKngxrM5FzkEIWz6Wk1kryl/6Ob1d05jJXhT8kMN9UoZGCslSiR
vH0a/DgSs5u8HHOVocEt8QFK+dRipGTw8KASKper1RYwZMUoQpXorOjU6oiybKO8+WPoXtxCwZN7
xYEIyECmSkuFWjr9g/RfBGqlCcl8OcCggWYhjzhDRAvHlfQ3VlrEMbsouTurS4U2RoVubt1uU7P6
XaX08KQLQ/w04qP98coRr3mguC3TxuXEtWUh6xltvCfISB5xePFqZzksT9oSoH7tjAdfHuNF5Hnq
YPKRMdvqKjamVsJslWv/zBX0bEz/3KHS+48kf58lAK6BkmtgDErR1kFSoOLRFPIiIcyXBLT3+8DE
Xo4+rXwqh9TVaTxgJjlGxTBP/tmmI4dXrJz92XegepnrECf+1VYvAaFxOD/I+ZrCRo9QrX7eQgDY
+SegAkuenU1mFdphgYd0PYMc12dnKVTR20JlNKJZnOABnVbnLCNHNKp4M9Ce0JLtN802GEWNLcQO
grJUqcis4Cdby2zhdd5Qps8eImRz4e5Fx1jvwuCNwaRB/7zNAXfwNJ8lVSQlpVX/Y8YrQhfPUrn+
LtKNOIdnjs8zV6ORrKLbbkvpvh8HfyD9GOVghdg0+a/5VJI/BKwounoXqiduZPMOpQ1gYPA60+Mr
o+Ydvz+zty4OC5erN6SNm7NhPj1M0t4FTiKysMNcK5crf0L/1Gzqm+SQ6QeJ46SSc7lukpZPAq0w
chab6+WKyuE66NizkqeL+hWHDFXxiiISM32W5TNNJ3ZTQdw+GUGO4RyN+HwM+M0lvj9K6R5wsL2G
5rBzH32LiXXW5jSyhlxDtYgeZ5K4wStgcFJ4lqzDX90KzQzfJaMJ9f3ym8eHA/NqAasRHfIuD1FZ
ZUQac3w89uyN7mxUBaqjwdNa3kgOtuc7i+Xpew3NfHcO/YrbxX7rIBFN/j3KJWUac/jQX4/o8qYL
omFCowQRZWO8RIJAiDzUxQ2Xb2mKPy5ZgUO4ok68FvSv4ur5aDW3CbkTZqrjZrHXDHA/q9qHEX5T
w6DQom3ojy4MbeLFiu6md/Sv4s4jxlEOUOuM9M88Fgubnx/VWcC/0nRlONiZhCg5qublPCFG8gR1
6dw4LuHEhWfK1rwWMVJtMp9NZBOIyK15FJkQ/YDRwSgDc0IccoHgfV/7fOqK0Q7qLwf7WzZYraqx
DwXhSJbEs9+ERLy1QQwdS+sAXk7A3jZpgTCDCA1M+it9wvKNdc0kVWQYCjhIfqdqwgDyaLmhm5Dg
03s+fNtWK+2uPxj9CkDGUvwrd5PO3qTy+qb3MiVsKscAbWVPpp7VJtLpalED+B9YsrRTe2QeI702
89LCFkPbZe2/QB92dKLD2h/HMOJ0opAv7r+u7gPFT+heeXhccFIOxaj/waV01nVMQHCscm/hXpOq
FjLnzEu4bT5iX32khAxEnfvRHljzhUk2rlL3KmikR8oPcUcpyPotUcaok/n49QhJQhGQ45V0/sD0
in2XLUhRP0YXqJqQoQbQiVlswdnYdRoosdaqvM6xxzk99D5LwYm/h9zgMNhPo8kwhx3A2UrPZ69b
wfW2DRKbwZhvyLtllv04IAMxm1sDNv+R0uAoNACZO+KJCYL7lHlc1Aa6K+rAGZ93W7RJvIGVWb10
4gNhVtlK0015MG0Xmhax4bzK1v30iMPos5Ju54Sd+Wz9J/DAZNHFZpErHdvEKENA8/c+YthJJMI4
CY9mL/YKMzMBnjtwxtEoAwUQK69+JcLS2yBtxtma2+9RqvPczIeo/zNweiZfHiit7ZfJBTi3YrPC
fV4yTA/x2dujKnoCKYiAI9aGjV+difF4fdALfR4Jee4e0ODrcX3HT3T+IdOewRqjffYzm6KlGrDu
h31wmcy4Fe2gmaT+jCVv1hN3Do/WGjLyikIGk1SPg0UyTYmN0zV2N3vq1q3N9+LWzH5j+bbdnM3h
fkpbzb1YNhynWOmGukV97bkDRxkp8LIoxsw1DOzFE83xfkXeL+VYOX3qeU4sKsQd74QGjppMMi0W
l+pKV9K4rsDMZRffV+Sd/fyTypRV2oRbdIiUkWT3Lhqwj8Js4Zwr6WP5/QJoaeuw7gnFCU2Hesu4
EWFnRxTBlqiRegi2zZGGAhk4jNpbv8z1l1uj6FEvSC47RXapRmiiMtJ6QMCm5ZChP+TJr3+0zP+v
048HPhK3IlaZaUWgO6OHuqxTT06HiAt8J0b1NcfohQB0W9Vc+azrWixVDm/Yumt10IV0B85B0sqi
7luA1IPrKQOqtEhcM4xZL6Y/ln4nnDAkeeGZlXNk98VmK5hUVsim2IYAELOZmZ0d0MwkqoGgWEAh
rNiXpN7mQMBYX9H1kBWn/rAydkEQflbnGf1+mdmg7fw6qzCoH+UJCmn79wK3LSBwvJG2m1cAGt1N
3JGHN2ZMDza3QP8Nq0zWELUjTYuUUysYr7T2sr0F0X7mLJENJrJfjoLAKUVe/FodBjV3P6Phl0vR
kgC/oMTYCO+TwEkaXfaM8K0Rj27LOP0n3mMp8oTSpKbpCuEhjvBMX5er0FR59KRRXwZEiBiwDQw5
Nmyygbd9Q4qwCwegFzCxhbcyiF1TqQ+aWS1J6vII4WYfGWYUU65l7Gm6w/Ahjq4PUa3PqGaY8cqW
Hth9/JF9YaZe+X5r/G9oI7ptnUog6KVURcLIe92zuiM/r9EUfd92I8NFNeTMD01XBcRjvslgRHal
+6LbUNtXyCu+IxGfKgoh3wvbSNHBKX8lZ1UJvsfTo3HlTSDQAOG8ME31JFTG03WU3u7wi1CvCu8+
2yUvFlFHjSkncvQezaCHmhlT4uIu5FEmYwfqsWDxmAMARfIZ0TYzzyg29UbpHEvfnXOq/Zrd7USp
WzXAs2yJ+om1WmRHDrNh2/oJvwqBkM06zJlVJTTQJW1YziKMBwXEQaz2IEqtMVXt0llGQQv4VS/0
M07fs050uP7UMPklx1KAce4pOQ0NI1P1H/oL2XZ5ONeIXDKCrYxMJwN8ZntvSf2y3+9CLca89d1S
IvXeVjO0ia2qQE/H+ccldb49fKSTNp68H4wfL46az8M1vKYnmCNr3bFSsPZnsCkYwLQb9YB1s+Mp
fIZx+UQWvb8vJzGwSLC0u3IYmUuTDb0sT99pD5NohbQZajTFrshmGRPBi9n8R/yJYfcQuYv3OUbT
NNHwfH2tWMMT/HUr9e5ob6iB60h+ud0sZ202t7gCNjrYHjPKlSa6EFnc00i2Rq94FYEYrkxhTe1N
ZQFZHLnvbktdkWedUPL7BhZdlNZL/JttP/ZljCtyafPt42OVgYdoPNcEc+LdailhSXLCfmJlaBbN
8WOCKfAGySeqT/WiaNTeute4fAQ//sNC7/FhN1XgMBr3AcHilmUSH+TH/7F63xB2wlZmu/wup6s7
V1zOpleoIMvuACbNHtvLRlCBWVUO9lMl6zbXCyz9BBsG4Yn8cELovg3MJMYuNrRl0dZ5eCi7bDVH
UQ8VJ/mLzWS5CrXn+eqPruAk3M2LTh5izSlKiDZGIod6kYqYtNuuVqnRsISKPWoQmxlR/LHd/AH/
o8oiJb3yr0zrZ25yMYr6WCroz/vNqA2NlBvNwY2RgerYjDNZbjh5CZ77X9/i0KMy5mX88vtosq3h
s16VQjpl5wLH8dW3jI1eM6oNpJ+Vnkg4DWdhVBI1jN4ZlqmMaCwuLvUrFa94Hisx3giBSKZcWpko
RKUGufXULjSJ8inc4PrlKBnFSiPa2rhzKHr8fsh5nrSuqg2tQrA5PsHiaeKPE27C5Bbemjf6vA4Z
Fl7jx/sJBWn9O4NID0hs295EvC/U36ReeREXqom3sm/M6P+D1kyhDz50Dydfvr8dl7Ebd/oi9obI
Z61iqL5MWGp6JDSwFwqFmebuKCuZfbKFuQdAr4lQtjYQD6ECSx3NgcTFWY6yXoCCIRiHhZoqoTlp
F39sVyZTWeUG+awJkvitePjAP0w1gutJHCT52GXFUfphYgdym4q0W2nbjXQyLaz9xmVnXuB50Dpd
mnKajqNEibj4Ytkc57vZmFEX/K+Vr0u6S8pYEbMYbA5vKCUwkDTdNNwovBJyPHHqHsX+f+0KGrcA
GewWvjWsjkFPQrChBe2/QHWulyPMcmeE85uO7vsObytni/ai9aR/4mkjwgfhPmkImaq57TUI21vJ
UMy+/CBzxoMny2SmH1u0IjpzDCQvWUXxeNJ3ziXW9wwJGITRbQv+fCyb6LSP4ZpwH8eSn0F//6Mt
nhV77nkLrNJnLCUowP2rwhb30uz8w/GnibMzMWBdDbi+cEt0DUOpFfiTVnj1fUFWzcqWTKuqZ1fl
wDyMaryO5RoomHI5Nzmfn6gO6YmAI7IPTv3fzoH3KnL9fGwaeBx9JbVWQW8Os9BHT+hwzOMR7ikk
7d78xbad+TrsoYrcLIjbfad0x9B+d9Hq+0QbQJjGOT/a5w+04plW2JZCqK/ZI2N0bn1DLpQmXNPE
s1eK6rAHgwPgLFho/E4fkZSUQYbsDdDb+N0erzL+69xmCPoL1RQ8gunvbUt7MfpjecB/C6SUayVV
GidfmyxH59lBCePX+rVL04F/lHvhWQ1ejchI1eRW/xe3mf20yPz6jO75eJxxn86xx3inm4ceAO2T
vOw9DMUk/DQol+TIRy8fjxA6cmnPUMBgYbNHcCDBLFdKvKih8Q3JfPlxs8Qo6CozqGDepVovUg9v
aG3Y9wM6jR6TI4Oy3SHUdkz/At7rMZlxCbpwaDFs6aTParkxTUapjcxqzyD9lwBe5LGr7dmpK5cl
FlnNzBp0cO/xFRmnsZ6SpUgxpinwbAl07BP7i0FQbKhHp/WJt9cf7waflyyYRE/BUH5QGVtz0zX1
KeJyhlKDC8SByys7SIQb/z4PkgAyiaAAs72Qiv3edn7uRBo95ulnUR3juFC4llaNwxoliPrelk19
0ZVYQc1UrzUifk7U0nMQWJ4VJMzpg3E1bA0+em+0Z2418tOv2lSAyclM0A78KzHpSHhxJjXOjEyg
S6lffpKwlyy6Tn03wUcRS+rmb+H47VuiKKMlojWAs6cGQC9i91/Kztu3VLevMhTOqJqAZQJeT4Ka
HOgbdGeV6KW2n1QoAem/wuq73RsupXLQT+9GMoeSKV9T4RQG+L3yqW2CuPIsrZYSZTp9axYuGv4D
tUYnY3WajM/P7gw6NWDf1v+zZCyHtd0Fe8Db3F9PHnd9xKUXEbjRcSVBmH3uWMwOoZASG8Zy2YSJ
B9mhlbhvEcBkGnDy5jY+e4YGxB52Sg5rcCZp7X75jwfKNO8EHBPADk/JyX0EH+Dz5cMAvsl1EyVb
2rvZ3eW4SbOgLomiYeQByDCi7F8HLH4e8R5SGNKiOZLHOuo3Q00b31mLxTkI6WkgGOATd16ww6gi
oxB2XN6p/tKvJb6jDIA9xwbb0iCQQwsbQ521EmyVbQ8Wbah4rLyfLXfdTh5K2BqOS3bsLxYLdesA
0tfQxbf7kp3P6DsbTMPXh09yCBm5djhHVA+K8TMQVCzG1MmrfOSpKiN3wq7YnzoZQ3vADR2ZTQWX
wY3GV7hb6ZAmamY2PZ6yTlB4LRHDccQXPGHeyXlmi2+CwCA2WtZbI9qIQPRcHykRd3Qpuz3d7LTs
ULEqsIU90Al5N9u0jZWRTu49hWKbY65EMrfWXgUEUEJ0TCY7PtGFK0keHFzbrONYCulXnuSbZZ6f
iBj7vgyCYqOxno7jAUDBJl6Rzz4wiMxa35dwBbnYMeyG8iekCkyMKW/Ho7cKQxOPNBHlA5rMSnK6
9Icu1R7axpUi2oQC6gOUujXyJ7iomNrVMC8Rw2+RVpDuiww7eSzlUk6woGlTpkjYfJsECPckPLGG
01X3WA5yRx4zSYeRHmqR9OD43PH5qiOsH+VtCyvuncFJ5sHwRtn8JJ9j9g84XHctzEEtz0W1Nq+a
smRPwQF6wvXeVC8bJ45XhKZsG+XP+Z8YxMBNjGjxzBWNyhuW8O6ImSrn5lvMumhNAgqbGriFRVLw
qwbfqGxtFOqUTN5V5FIG9CEJtvoaVzM6JFCoD5eS9O4i4rSbqvLsccmyU0ArGUs/e6PHT3La7vXK
ZLkHRMcMU+IxiM6ONBR4zQbi6OhQKDOCQZKgWi0tfoCcP2eKMgRwUtlTwxryYw+6CUaA0g/pi77w
5/bw0y30x4vy9D/XQRR09Sgb7QFUcUnK9OhorcGRPpy1cs2keM65847RwV4Idc+1pfLKCahYtuhm
EppXB/vomPfxNOOHBp99DCGus918+18KNNFc49LI+AHzmycVoSCcmltMGh7RRw5LaVHQN6HYhDdc
5lNVEdg53CzbIx/wpAGuBYRi1y/FBk947oQ6Ry3bGHn8IFqAvFxm5CCu7dDsbZsGH2Gp21LISEBM
2rH6AWOLBJubzpNCvSefT1dBJdWOp0GdcTXx78avC+1lfuIL9U2Yss2kVxqn/GkOQ7fxNho3gka0
DjEhyRDJEAc8ZCrAVdeSbvJ3B8hlPWrQoFc9y3J1Bkq00U/9VY/Tf+3b147XrD34uc4NllOH9FYO
HCzGgzJB9B5I2xn1s6svNaR5VB+/dv+e4gixdkyrFFrMDQZFqirdrOkcgHrHVSe/4w1JVPzfSd3S
HbscARB1n4Y0VtnQ2KeNY17aFx1j07fI9pEbjY0OUZAh/JHgATrrC2QifQqlQzMxfUgdQId+I0iL
u2T2nC6Qv0Ja5KkUNJnGdrm0zBIwxgs+fKnz2hWm3IuH2YS+4lppjdr3rP+jV39feNivLoPUxOK4
AUr+zMbraNQ2N4PH6LXmtg+dcBGsUvxJgt0xv+clIC2C8ypIlCFA5+xvnH+VVvxeSh4raHQNUtcB
396+mwdxp2O7zxVXdzlVbBZS8/Z1aCPh2F17R9TLrTKvx9Lcs+s6jMtjP+zCnIuFoMGCz7Uimin0
Ihl12qWOzYD2jGudYKZ0AjGg2Zmvkx0i1fP0v/4q7it/T7aVjHWuX1A5Nd/zbNFXUwRPP91jVYPv
mDc7hbES6ZfbGcSnbWXBgT492H34VWljim8IVvlt6jU2GgP1P/EPbwz55cAT8Jc+Ecf6xqwYBAPr
WcZ20RbD7ZMNDGQp0nh+0Ex2XidniQgD6oNDHIvovRqsL1Q1wiz7lw73Xd68Fqcm/mjvpSQdAuw/
bQqT/tYbER4O2mAYX0PbobrQ3vcJ09edrZt5sjg0TzXaM55JoGN0CnJx1KZeWLQL+JSQlx1U9VyH
e3oIagjhNXXkXbDof81mWt8uTwmvGad0HNT11zKxoHDLnNy0Lm+jHw31IghOw56O+6jByp5oAvZt
yXGaEJaWZL3XMBhGPSVhubD902j2dxoWGLdArT3nUD0KnOrvYrVKhsBFqCMgISzk/Ul/UtEWhe2V
YBgalF5XGQBWHXJqiDpCFPgdZ5DkNJnVRUxb+eAaaq4eGJ+56igbfGxIWO9JTs+aC/egeB8rMR1p
YxyAl3Fc8jtmuVYEkb9ih4P3P9iLN+pq6Xz5xN57VjGJAtsaAroYg8vK2NS5k8l0V2B+1uRYSiJe
FFrnF0K6+T7+mMn8rbSug560X1BuuMkc5tnIytX3qE81cFhBrioqKEVRE2+x/kKrCum4AJYDYPu+
TGcrRGsJTPrtQnkWoD4kr5q8ZjQh9T7lqf7/ZGOaCyk/gccG8lAVWorJgCA/pUNTROkwxDGC/1tk
I0/6BsI+eUr7q1ZbPl22ZTifqg1N/hR6GPXd895G75uyZcP49CJZGMjaUQdTCCk6iOj7Ib3ZiD33
4J7qnz96s8dEVFTbJ8ykSSNnrCRUfvIlHqKvbQHV1b4sWRS7rkKkRd0L7RSR7eDVrOLcgRLhvSN/
YNYTb3g4txfmeXMMmAfn4XGcd+9FgO4s/lbii/I8V7e5BgxVBYjZyqfLNgV/ap14vi/v+52lZJK/
wV8cvnn9rCmJfD/wloEXG1y0a/vGN8A1XW1HoWS9rQLPcLt94Dlrom9GGalQh1qTuuoTj8uPg9/P
3bNY19zhpKTS0s07dvuHLUfULREk9k0H+HYjgxhXU/v27jI5alSDHJFAZURnZ0Vpa6PIBNifkSpn
bSSm5onpjpME2Dy6sm/zTfkAojSv5aEFEiOxh01vAtEL8m8vQKFdsXBYd9w8wR65vWPWY6zAmUzi
OnFZD1DHdPwZ+t/LMuHrIbnnEIIFi0WkzLCdcVq6BGzjTZhkVp/V2mDDTa58wC1vvfnXT0vi/4wA
Awi66sLitvCRMdEB6tZzHLoe0NQGcIsT0ZEtHeftoOP0m9KjDRdyLYyg+xWrXM3p2pDp3xXWfpIE
p1mVug3dB6RX6Q0UjvSehjXgXBy8CtIrBbh/VffF+fUwXfaSKTj6CXRCJFUul/9KyASHu4S9BgyB
gWdQ0D5w8z5W2JqfQm9Oj2t7Livh5wwKV957nxkTevnMw78+pl/GZCyG4fr+A6lJ4Nf/ABA2MpvG
/pLVXpK6GIOu9kygj4+8S9203HJ9nY6Y6kArYzumEx794ohEwYpofhwAZevgQYcYHjMt/rinLSCN
aMyXK1/eodw9P42XqefIJPAKdEG9khG1CTFPSsEAr+qTFiLPDlAodYxKbLqsZqG0hRKaMafk+aDL
sWEtqoNlxJTbN5JeO+XxMyTD+0Qghqhv5bXAZl7J4J9hFnS50FdC6iGq6bPLpZPzqKBu4j2rX8Go
AD6h9xNKVEBJI9xeeOHreRHtblKe2qayor+fbwntlAxMD8uuE0Eo5N6QHzjHYwbIqrnJjcMzoMvJ
WlnodvucAr0vcg1VTvqzYw7XrNw3SRXSeDK8ABjoRrDXm7jRuFdt6cvRlNwoSA8SO1OfiJQHCUMG
sbzcGgJO4JdmFbNsKySRPBgirB0BREIbRGrv43gSshebsAAk9iUFK1tUw4IasONQCAgkw4hTd/H3
vE74FQanBRuM0XAX4AQEJoUUinmX9kzTq/LHdCdU1pQXUrerhkBk/wRij8hVPuuF5zKgZc0YltZc
DemVYxMaY9WN9z+e4SCNorAf8xKrijKau9BT40L5YTH8d46dAndoRZkQp+KCBT2AnP0guiQViYqA
cqkTXzsZf28WNPEGU02TTZsvFD80e7mMPaBKFPtmDpAnp0b5GEh/Dit/35NhJ8UGGQPgZtV7969k
bRoL4IuQZBgTiPPHE0E8Xda4McAzyjm2o+nepUEQcoqtpMf4s0FLQ1wrCYvTiaZj6yaVsut7kirJ
ZFGJ4HMHylGdEBvW1fkZFXTpoRnl6HCiyNh5EAlrH9rphJjBaS520trPUIxJ9GSgOhhnYGI9DHrp
LD6MfZu5f8coNXqseeqH+N3o/LtVqH7QTmlXfU82FMpZY1VdJOBuDivFiZfXMoOaCRPXx0oLPuuM
HhHWLUOjgU6B1LLqgZPQhX/55pGY/ifJi508Kp+GW0TH0y+tPRuaOps2nSeMD3a8ckksj7ufgBad
ORCUq3m+SKWLvUKn+QmSpDtu2zyr3Ae52MujQLl7pIW6keatuEnStKMvKWufwYHOIXto9QJTxAxx
9VGW7w326FH6Jee07Vt/5Quxri9Aln8jXXik+MqyC/qoNpzqgrqTSEtRWNGoynCnnyq/GcuhjhQr
CQmftqcPf7lZcjicoTit+UaXoOUp5Mmnp7cNFo8uNgLQPqMGJEJXVPB8et4IEXCfiUBcGbpGKvNC
xeBis8Gp98BtaCXx0j3maN0E8SOCS5/TN8kmdHL69pqSyzDE4NaHie0o124kSPkmfeB7A6K6Ar8Z
x5UMTYkovKIs7gQ4jomlhFTs/jKrGSmHNT1+MY3mTWan0X5z2CYkYQ9DEaZ/eHGGurjtXnBl8pfC
He6onVnaBUoUNabANzMFN7ApBIxidyummsZ7KcaxA+jlMnlXoMN/zuXkk6L/dwclgX6YaUkAA3xx
2TCpbOa4SZ72xYYx7iTGZklTf5A8qVvbjUwTFpbnyUKn4EyXsp8g8Pe6dkafr6Q/HW0dtewLo1Ad
9W+00b3UMhcnb+aUfq6QLDU7O0V35NIUrfQY+TNI4Q25lqc/HQU+tsonbqXuxkFBfAdXTSKSZwkM
4YLShNsna6e7dpHiP3FvX5Syz13F/TBVSiT0BvSmZmBmtN6Rxq62NVc2yXHyntF90WJctbDnKN6k
5xePdhvChUe8y3QbVN9BKvHwb1lqWjhil8D6M3men3GzKeseHTUyfWG/n3j4d8KZfTcThQEAakRK
GVVTnv4NrDZVyT3UdmUt3DxDxBcTPgbftG+/hiKsmuykZsMSkdsUzwAO1fBZ7iUbWTShLx+QmNMi
tP7vIBuj7nOrW38iO+XpiNvrR56eXfwUYlLabTTcWlSAYx59doJsCYT+vx4cUhuHD+QylGzIPE0z
NzsZmYD7MkTQYfab8oNllaf6TK041akW7Aja4Razuv2NEn5GeTNH4GhBofh8FXaWo+gouI154CFR
weRjnsOWbKhN3g3C0D+NqMK6dRX53TAqZs68Saul+lNdFvP3xwsHNu/ohij6h1biWOjsh0s6nLRn
uWrj8R0O/lquYHV5ydKjgs5bTPlnuIQnzEyDsHhOw2Pd3/9qUl6snZKw3JgYwNJoFBhabO2NSUbK
XR0iNJPcwPJNgVvsWXJIuY9SV76cpghU9BKAFbF2l01h7PK86r6ymBd38S3EK74Krvtm/Wtdveju
ENiwh6TWxztr60L6cBRv56EDFa2Bve4Vab4U9vPcnK7tpuktDJieY/QBWGyUAfJLAHaoYIRdcvZh
AQTHdzETv5VxF28FrKDZW8+9J8DFsJ1/17zYXKPVpsYv2pYpO5wE8KhXpuk53Bq3bN/SunNhCzDI
ZwPMCy+lKgXQ02fHl9PjPLV1v1pMxfCt3pj4ixu6NMTkkAzF5plav7xmML1VLW/1uK8LqqGQV/Ec
4d8/0YSfI7PonbhP8ftzRafWCkiYmsMmjBT6e3q1L0NwF+ec7dpVeyL5SsxJ/t7jH5NKOOG5/0L7
2xMvtMTSKzTB7fAcrAjlUOZ5BHOso4pnxdfOCfhB4l/SnsyUYOrE4Q6NDHzNuzVCpwMFo8bgxJ14
YdOTcj2dNlpRTpy4fvx6LQIw2XGRmMQNGS2Ta13ia/4PRw2XKxGCs7af7RpA5Fe96Mx829JdzEXk
aIMIC+RkJOpipD+0FqUReqz9u1ewMqmGXlhDFHcppK76w3/wgJbvY8emR/LYqEaWdEV1naDayWkm
2gcDSUECCnThfzRSBI5irteKIXHxSHozaSfUzP/0j5bSBr6fZbJcGdJzDzfooOR5mxnHBSKWrJzd
spmGfSyM5cnpJIzp1xLboHtoD/NlYJYxGyvq65DbEyQSfp0fXzWXmeNew6s3mXu1HXYlbZ2f1WOb
fw38edpyW25oJw/pbsqeFds72PnNxKrgfYhm6W9RT7hC9dbvGDz//0Lic6aNxzfBSPr7iq2MhYZj
R+pT7R4LeHji0ewsvCcqOAQd4UaFMabnyw0Egm6qoXWqE74pB+sfSde03OG2M/CIYari4S7pKKRQ
g4Zhvku9h10BIrTCaZNG5Hd54UqQFLN6pwAnAGMC4fJAUtsHWANk/RNDIwddHLz9WgB4AAU292XX
Jhwq8+ExwBTH2Az45oGFVEaOuk5gDsGhdQCaEKoF7n/hZoC3Tf+m285JCr8AnaFX9Ryc0dd61O4z
g3dv0oTtlNmksnOrgKq0P6S8GHGBCKCru2OPZk76RCRk15zshobn3FZgK4qym2fKvXKWcO2+oXxM
aus3KBGc7En5MEHNLuy4fYc3Qyvob3/NMgQfM/8cJeu517i9FOEbXWOAmJQU2L4VN3TJUKSIqyNk
DTujq0cqFZ8lmoEV24QyU3j8bHdCuVOXMxESYPR6siRIgfslh5Ux3ewF+v0PfhOBUYykGZ8nWWsq
n6Xh8Uh5k/5sKOHbCLneqJmOLCpe3+Phw1c3x3ASyHy30cY9xayckh89dPxBrPmS2sHVfbq+L893
n9V648fmk+NhJQcQqKGGggM5QRPIXgOHR6eWYYbg3EqjavLux+Ya8jNAk2S5DYIXCCmO3I4CpYi0
vFxfAnhKg4P3JTq1i9qTTOvNAQDEBJ/ZPyFPSv6KZVgKLqKI+vYTLSvemJae+ZVVSZV9ApOJorl5
H67s7nYnCZzJaJuQhwBZ4DMf4MWKiK9BUYqn1KYctNm3MaWjBUdJG26EFSjogIR+DEjFTUzwM9Ld
cEWljWmUeXuBIgLSFmMXW0pKbTAJdxjhg45XQpghGY7nKuOrZZRDotvPEVnGfH6ykGNIJRfKcV13
STqF2cRiNH3BJkGSyZ68oRj9ntZVzETCBAb8fVowUuLWtaz0IGcgF02Fn+XiG8WRQmFDw11e5CSz
Z/iokFsApc56QglEcGk0T3yIxONxdw8vdAMc1UUXNpxcJPilwU2TTu3EOzUTOBhr5NE7bMUSfBdh
zH90J907noQNsWn+NUEbXHyVpGpLEQW5IkdCQimiJiiwnVg1o5ryNXs8xyZ8yR/mbHs1rJtf1HCG
us87kF7jFG7hwewRySYe52Ept2hd+DRcbWNCshXs1irz3wj2+AbWvT9BcQ9n8t79lBT49bES4G+j
Pk7SAsMa5i/dya4cp4SlKS2IF8miwTmUFyy024Ob+5vZGjXO22fUgoJLzxyY31LqP/VzL2uCbmHl
4S8J+17XXzbIu9ZmSeBbtlK41g0Bf949ElyiT89uxCi6ZO0RLxPuTAjcmCvU8CyEIIiGSHwp8hVP
biGx2e54kHHtwwcHlH8uJU1wptSEgslXSfcRN7b/TPUAX8Z428vU9scBRGpnbl9N+dlcXO0Qoefe
Pk0YZ2R7mktavqdmpF5aEURgnSz6Kjkdlg831Zs9wHf2oAbtl71z3M5DlzoctjuhIQlT3g/U69sv
9EXzuQ9CkelTmtFmLP7VY3752xz6yU82C4gynIsqfvZBypCmOpCBlFwyKBNTvNwWDaTcBbblW6/0
vYH8yCSIHjIZth4kEg2Y3gMmLzKhSJj6olaM32M09MB7Wg1otHRjODbEtA9uAiqbp06RmZUhJBhl
34eBI4BvFeW8FJ7HvpQ2uDbk3TQGgBCWXv7CuMr5JBAdYVTzwT5KZzZK6xWKI5MvqfJVTZTlZdYk
RCJqMxUmzlTjBM8TCxhg13THc7jyRKgl6FynxL8am3vlZOpoRsne3fb6yJqvP/8+m99dWPdILRZ4
MM2zpmw9iQe7LLuPZoFdvy63VYdJMUMMyhLoF1+Z0kavvEqqQW3XFufxaRoT0XaR1dJwZ+/50E2q
bCuXh5XVYFVJ4Ex9ute634pzdoVmZq6pyvzMRH5bUdogY5vlB7WPdm4HZ+SFr3lS/UFXIr/aqqZb
QQ2hgNpongqW9242y9GIspXNHRxLOTLqARC1g5liUcQeYCg60Whmvlnxz4IHXyzlWrS5kP/4v2yN
Au6uSqaYi5rs6RJ9PIZ7iUr18mA7u3Tqa+RkdFAKGD4QzBXlFbgnv/eF3/ZIXjUHTVbW3q0zAbEP
jt1UxOCzjKnb9h3mr7J/nZNnrfLRPUErpM3yEawabL8chKS+gvxaeW5Z2qkZptTTBB/vIN6ZRsoE
rc7PoMOhS8Jm7bO2dqB3OwhAEf4e/Oz161pOKTMzv2fwADhxIjOt7ABeA4pBxKVVhiFyDeGHY0CL
u7koq6xmCM1oZ36PUXeFtQ1o2M+6rfk0iR1lZspDP1OsIKafLZ6GtRbD/LxYDicb8snwW3bzGa+z
1PLr1cAoAp0ORCKR4n1bs+KmA1kK67lW32hg5kR2Yt07U6CIreI8N5gpU1A1eq0pP7cIz1yqiFiG
6Cpym0mulfskGbUUgpDVHJf90ow/PjVXIJg5LZoMMzqk1Ac4lUZY+WMTPXNDfFQZeUHoYcHxra1o
UszsR/8OD029KYxdzu/STzDyS7k769VDsqOxwKUaAwmBQMTlP1bI6S499VUHSWOiryPuGscJYSxX
VlcgnrocNFBDF7lqr50pxqeNrd2YfbCfDuLjQ21sDDiZ60YUOqAPrjaYahWFmpUIl6EccKDvphYQ
lR6K55NZFTepM+Ror5vZcgdRaUJoV9NTbvIhGOmvsX4yFmLvhl0AnCqyZFLwtT9L/WdZGitvJ/Nn
kSrEQkMRytJb41o7vYo0l3OJBGJ+c1HOGPoMc4/0hBAvHpO9e4OI3tOH8O35PyzTvNsuJoPwRHo2
dwPN86g8rw//f4N42qO0HeiQzgMqMaBre1XxTzmPCN2qxyjGBtMQWWw62LnuB4hwEZmHSTMvqLa1
mEpbHX/hsSvBwyvEy2g7ypXtH3cSWUHHCiA5nDLBdYmhUL8AvnN1BcbWb2+GAjqEJFEQw/s5Fu+r
CmSeX987jzHieJuJfeOo2FdPhB/lJ+SInzgGt7sC/h2DakMuDkGtA87dscVc54cBF2t7lnmsmHWS
gLRFBNgarwjJsJq71t51XUobVrfQxl0nXA2vYvP6MalE8zWJKxJ96r9XHnd85yEJqglUGIxnpunj
PGi98zFm/7/Q6YsNgvqGWzQmjH5rBAifMmNBy3sl4ho+cBDy1DYqNaGPT2GeN/yghfZLy47JFs1d
dHdn2kG6DUtqqzo64G80LcyRGp/L3OuxM0TUMvrFD5MuvuukXhEhj5f2f+D/ffivMfrl3S0rND5w
yB3O9A2sQ9XOuXVlH1lOjGEGONmgvRzRkX17iZfpq70mBvCcYjp99V2KG07saQnjWoPdjHW3FNnm
MJSTq5R4eG9hkWl3x/qKm2PVqQn6iKlYYNBN7tQ4ecgvNnqi6Hqy1AlQhoECesPlRBJu81DyVXlz
7RUjZaduU/ZsZWbZ3Jd5oIFxHjWC592Ga3auPmAuN2b0Hg3phFu2pIcIBxnPfrYCo8ZTyjepBHb2
A//XZghzuGErvFY4uNTBJGhcxEnaeiqGOZ7hivWLYmYkdY71ZLeGnUnndApqBdXZplkJI9qrUw04
e6CkVjRDrYbcJKxXcXihTaaAXyWplO39HzK6HXuVIrSpSIaPSn+akcQDCzFYfEkhx8WGlNV3O8WN
44a5CDjT3BwScXdJEaB7LnQzCudIRJni74p7UidjA/tA1pE+84daJxv6a/l+y9+4cPkl/Kr6mguS
zkFMZ6XOjLTlY6EI+ehyxqz3lPNPAk1MRJ8NU6FBiUV/xE4A3uyGLH+AZx9t77M7+EQDq8ryN/62
z2bqvrMMSSWxzYbPCY+YK62UZ1QtFAdNJPuOPKBCKQGPo9NkcOl7BqZHSyQilCm44AQ9MJBF0vB7
HlfGVhOt8lhzuWVdosSYG6x78RUhVhbhbIy8tvRdxkNS+zdkvLt4Lfa67pWxawWwZ5jDrHf5lsVv
D1MX2E+/lVFC/IJ7pQw/nBvY1TBz36ttBBdF06BoHMg7uzNcMhy9VU+yaFfiIlQn8MNx+gWl9zMN
nFKJnREea4ZmGFeU7PTpmk+aUAAEHBYCzTZESiOsXhWymrW1vDPGMcM6gVTXm7vi4s2Aoge6oxiE
wySbRAaZ+VC5oVMQNUbbr+NGse72Br343K+QmZH2cLy0/jS7cWnIh0AtNxKApmqy8OlXvVzZNnCJ
HCs0gDEx2At891nHE4jbilwiqZ4MdROli9X2pvu3CstitkGSF5aEfpFDc2PHrCGjoNCluYRzWlwp
XJbmIE05T3cRVxMMiJ8oL0COuVVgc/swF0Rb8tGcoJLiuOG9+UglSa81oQedq1RGQ6k4nIqPwT7Y
OozL23kc5xmdG662FM6bdZqbTw7n/Z4zvO3EexM3K5mgW1R/GGG8FFNwznFaYHaFEQ6/JYo70amU
20cZ/v5IKNist4+TRP1JxGNkcIt6VqrKzCIfWM6wx9/myXg9bDLYj6CRCqmgy1U/Jqu6gvF2+/A5
aUpinoNKKLXl2Brq4rDfdkqMcta6uODIb4/IHyO8qqkZnCe7S4oO1JZ4hMN41AF3lQHr7x7PiH4k
NrppO76TS9sDmHjkaGis5QXGcUvRRj5YFZkWdwttxcI4DpAk4kvn48a3bnLoCS7P9aaCeThUDh8p
LxJZnY3edIAsmvDPdS4BUih5fla1IrA1RjqEfvTxsoXBNQ/zZzEUW0W61jZ8IT5iShhJ0LItoFbs
tThvmu48wwrKjpzRjpUV4jMN9ggbsOa1eIXc8tFpl7XU7SqZrFe2O8a60i80I+lPvkkPwa7ivtC8
4rH7bPee+JxVl3IgO4LrRVIO39a0ScF2BLyKxjdV/Zx0qk88U29OeV5uPt1WkDpZE2/fZbEM+xgf
ZDO2Ibqk4O7b7R52Dr+7pyqDnEjjG9a7GhDvxoMs6wxX5qNsojK3BAhy5AHk/Bsab06HR3H61paf
MOzxm+vV/PSg2FQ+WtAQYwIpYAPxQVJzPTOiKMFdXU+e4SmYWaAF+S+pLghu2Frx0CzQ+Hkozpom
xaz0xvMB9+rjX3T5AoXeEUGkZkZ9Oqz7YXuGuotdd9bzIWP2g5xudyQrd6Ssoum/9XTsqY/9u1u4
KA9f8zgIlAso16pgyyPnhIXE9Gzt0O1A8x7TA5LoxEO7WRZ2GjAdgeRB8Nj4EZiKcUrnMQN0DYjL
1n+/axNW6RkiMEIhgIHRpFMfgRYjoafdM7r64e7JQe4gd+MuQefkMe82ow+UsgCNbinHmZiMES61
pbfTa/IAOlxsr9ilL4tnQcMW4t+3FupjNCML+k6Sesjp8US8bTyr++Rv78yu1i90go5MY0BRmdv8
tGzN7R3M7YPIWnWlDl+YgC3aoc8f48mV9dpUyfbzKnr7U6Viulou4kgXkBuSiu/Mi6WF1XDP913S
ZyU0bT34IM/L7IolYHrMMTmg14oa18hemeg9UtYLoK3Gn5niBog7Sisk7SXy9oLs/MY5SibwEfwn
EJ1G2VG6lxnFAl23kFDxJq+FTfYGk4PA+noAfoNpcu7F3XMoroV4b2lUg4fT2SckD4ipTsqtC0Q1
009l7sTQ+TqouZBaOEP09aIGfySsIaV/ooeEsNSxZxeqM8y9BBbdt1JiSCMSehaBAYULoQGVSO8J
dmtZSSxYe4/e3qznx1Oz9p5Qmh0Ofk92wP7tJACvWt7j3/t+298++ELgjEvyLQrs7XRv3TjPOn9S
883xapd3Wr5PLbcRwOcXbAqM2AcKTMNRe7w4lYb4VrHgpSZWmnBxyEBFb8vLt9YBRlwj4atuOePM
Ed6isEO040K9vCm5nbB0xY59m6C0aMVWRmXt/dtEQXlbXinicmwLOT7wGQ/8ZX8h4kuTdWYCPyPr
shZyoKlRc47P1khriCqAgVDRPCkUlPWDtSVZlqS8jecjYkCZOAofRo0uSnVPQPasSXgpCgpq6drl
YnvbdKtwfhi3fEAViEzI+d7Ahe/lKQAxVfF2o4TMgdO47AESka+dyJwpobws1UY8AbMGAbADK/bB
Mrfh6q/a0ez+msPHBbrV7Hosy6DiSG5mSFZtIv25P/pXHLhlcei4fZFTjIfDez/WlinXdCdm4tVZ
ZndXklG4dZD/hQdV+oxlJapBfKJsFFTu59F8v3HQS6Ek4u5fub1Q/hmOm5RzZ0N4F/4kBPKWs6Ix
s4nHECOnt0ppc2y5v+JuRGKkz5YWFtA7Litx/9yZjj2CHZ9TcIGVBKKzm9dwsd5r6MdanxT8gKHB
sJ7UI/Uefvybd32U4TmaHCDKH5eW6vCLOCB91iFwdXGpfyAU5NKr2nGVI67mGqvo3EjxwAsH5miB
RkSqau+oJlmRGsEm/AcRdgqyvGSLqAEi+fQ1+dJlU8rM7aomXHwtx6VfagntCHeAjR2NJ/QN9ngl
UPVlPcb152ONZC4judhd/+matwau7wWT0R6dQQf52LM2BVVyHtB+7kRYTDLuGyBRop/9vsEpoKNA
mXnKkDA5gnVU6Vm5Lcyj5UZkIhM78218B1rh67cR09tuP7xePDtI2iGViGdP0BbiuVaKaMmKNSjt
B4JfywnB3hP5UxIgjfY6dWsCq7O75O5Vey/+jDdjP3N5jLbkBTkbOdOSfsFlBRBQclLYmwuFERGv
r3GpHBAj2WMKjVnU50Rxag9TjfVG4xABwMBUt9Gib3nG9RYY2DonCzct5cBDttIATFVmVQuIwVo9
DK/EV+WzXQWx6oRYlEXgzOfGr32ePx4fduig7S7yA8hW2jXFQzNJWXGOvapoGV/Ybo6ac9RyV9UG
Dd6iitApEvDZhd/a5YPkvpvZWrcVXot+jrOvwGnSyPCaNH7EMdQdPfeD2ebxJXI69R2OlEiovj6R
mSymtKeCXU07TYXftB8uC7ehs6lwEYSUs44WEY8lD3a6/0StkOXm8elidP//Vld1SWvcwD0GqLaF
rmq12OP7KGCMk0Fqg4JE/IgMu9VRPNqFXs4r6wswfjAmQrtZpddIGRhJSvpp+u2lwvl1+J1fwRgc
Dapl5w0QqeetrEvypZnebOXgYLOdcpWnEuKodHsNo71UZ32p5xTWo7AjrclKmsg2uk6Lfnioy8KL
AQwGiQe/yS+MnPSDhfuIfCzeCgsCan9kgcUYrIkGf0nU5NwP3IZo9K8rzoP7GRCr6NRlAA51bee1
oRl33nbAZwmVtkQN9eTCQQiphzJOky4kKNS5Ao4U6a2U43GhjymR6n0EjePJdiJTWeG8IPYH6c9i
ADFDUPO8TyjhSJC9SrqDUTRDzRTpa6ewRMaPZk7Nt9dr1HZ+T8MRaBMlzhEYy9MLrIn8chqjLbzQ
16FYuK5558lAYNrEuFR6B83Hn6lWu8uicNZmxlL63Y1dhxkboeiE++xDbxuEq6lR5Z0ZX6XWlDMU
r5Ejlq4/zCLAHlbfPofRYanbNYNE3Uyge/N4vm+LLR9FRs0f1hs+MFi1OF53+VxLM2717nnZnuiC
QEbDk0nX4MWMWex2cAYQjCYZFjYhJL6M9i6yqysgQ4Dpkblg5OIy2d3vqZnor9vOVMDhLk8zXAbE
/ub79uTEAujMgnR0VFReNphUuAlOJBgf9I+TUnAmb2QbdzuOvfocmQjh3bGjmAUjfGFkbeO1EHL6
UvIMVBc3rdlDBEcAYAuzwqtAOjea/xYDgErVBCbqUo96ZomNoKEKnDNbQwzj6+wlq46kr7mEa1/s
eZNQRmhnCy+sW/sD9ZTDJGsunFJRCYBStYEmiT0w6mXQHSxizvgMARIQl6ab3uds3ve6Qv37QRMg
BBl/h1Wmf+5RKQqCvtGbNZP/MtuDc9Gr4akLFEIiDyx4MV9opqFHZTGFvEnFxV7v1O1KLKBSqhc8
8VqfHDaAKCytWC1Ihe55foXK3TBdnaC7g64djo/nT1gYM0d2AQvkHvQpb83SHNzzVMlCqUJiItNC
jO4UtoOPDvy0mOrHjkk1zcBoADxTBvfSmY615CRTvwFdrCWfJb3NFMzYAbu5HIGDy6RWf3Eb2Al0
sfDAQBtkL+tVTftQdk0oFMB2XrMVLI3FaZTz93ppsP52ksoCFQ3PQ8kzfPFCJLaIXN+DVgCNalsJ
YRNxHjw/LC+1xlakk9Qf8+63YPnPm6hA2GKCCxh93JrseCPdf7j0vFCxIjgqi1YtQpwl1FMC+ajo
sWG+WrrL4nxsPsaDAULujOSss9xSKSbT8cMVYMr9ZdUcfx1F27pn1ma4OgNwUWHsJbYBZPMKtUDk
bXXE+uT0kEIKnTO5nrnloYdDWlbEsoS9m+qFDWBl+8hgmSSnwdHOimB+MgST+zmD7RyGUnnaqLcT
WIflGCJtKbtt0+7ZyKZRprN/WWm1GYzLI93PLdrlcy/807Qx7i9VYIxQ/S/cgkkSTgkcaGB2sKIt
htepzbG+zAuj6ZqriIxDcHwJqRHtqYnZjPHiypZtUURDWql3NtSySVp0HOqJOsPQF3rWDTDl6Ux1
dK6NI3kfFTjrY1yHcnPSNPTELqcpN+LSpcgSQjTqshBPFwLlE1/NNiHFR7bktPliNAKc0N2CqO46
VHyZmgf8FyqMayP36ECwAkKxfaoJ7fB2SfDtFLWNpwX02NDZ+FkFItxheD0CcT4SF9vXIEIXWcvO
837yPufwO2dgfjLxOevpg5oEXyfosv4OHNvn/SUDfuscaMWkij+4vkl2ihnzHQdpkvYbJA3nMFdc
6xQVkYy1HG8MY3wF057EoQhCT1vcdRbfeu3C3tRglUjSmk4UFdwLrFL8Wvt8AsicXy2HxkCXv2L3
yWrqlUfUdWA5WC77EUKXWq+6JG0Wae6fnxhAuFyGb4tKKHB0+QFSKE2+gBDj6O5bLsWGXPjVtVJT
c8szB3H6+XtenaX9IWHQpo8ANUKJz2XW4nipqLJUlAC89fdLuwwX1Ga0g6esl8Nkoz3Q8juKRO0h
JBMNkCG+uaIsxFknvtBF2kfLOvmdW+HrISh2Cgkebi7FkgGDzNDG4/fy7vPuZyn1fc7a2KFN3VaA
3NP9sUzcBDS8SlyIelBuNWQUHsJOSxsHyxbLSHz5L6XRIsTaw7bH6PFhr+szvtgOHq6cp48X+xqN
OqxtWH7RrDUm+BHCNWhKg52AVf/Ysihf85iHTrpVCQzXjDo/bQFow4xgNNSkqGDmjLQTD8CcBH5R
GdGAMsI9xRTgFFTvJOMEWY0gN2CDYP35luVHgXZXYCvXuRJBE7ntiFReVuIJF96oMP45a+H2tmiL
DM+2FE1vUlXv9Or7puXZio4h2L7BoRrHzT3kUElPcojnMMq7+Z+ly6B4DoY2GlfCo9UBHan5Dvqy
RulMvbQyVCqOyiS9TfQ/1JiiSA6pcNZTpzbV7mkaShYnw7BVV8mAKYqzcaW9/yBWnmchCG2a1cDp
RYCybp5aRriSG22XnUXmACeNvIo2OJxcxq5hZP/87yRcDXbKxFBiSlRN++yibKGg7BOWWFWnrRw+
O/3KYOIEwubsvIwRPYLj0SZZFIDjjs2QH3c1PB570N1v43XOrLdzCVf+MP6Uoe+fsvbW/btd06Fz
g1eaZJBXzDh4T5kqocGK0jcnFcnC0ELjeVya9n4AI7wajjT9TRm2fG9almtw8JTg7/fwEdL2X2ue
MOmhsf6wsMTk8CjR5xOtmQOufeIzQFs2Gy/G4ejQMmKe2WwM+piaA632zMR3byd5Z2GufBzOCzu8
nmXlfsxRnEyR5c1eAXl37ccPlATHBzjgKLjPLHWaXtJCLZgQJvcBQjwliCwUnMzSrb9ryZSNVd+U
0+BzcJGj4uHNtq7Gh7JbruX71IYs/SHiSvRrLgWfRljLwQgLX974B/qVps41cvTRhp3UV59xM2x9
FJQKDq/C1ngEabezO2grEvxWrx3JlYzhft2rFtsb0zdoEdCwMwBNoDF0wQs4ThwBzEdDITcPHcvp
BHHG7iCK9LL+VruMSoShFtDtNbNd1r/WBzD8iWCxZrhpIbOcv6uK/c9IvUdlVeErShk/BnGZ7oLY
Jqp5kWyH7NlAooUv1t7H2qF4w2shQygh8tgcLcZj7OuQ3M+/r6AUpCfzEAy+5SF45VrSUzA4q6MV
IpFpbikRCRvsbbBeQZZzZNr7aomwm+kj2C8x1I36f5DVAN/biGnuuhKw5xDPhCPGtRElEmlfzKJU
N1e9b+t2kOrv+1TiZoYDc2Q/G7v7rvBQ6Oziy7mqtrwqa3wnXISdP8Pb24T/RWZw9YfOnf7lItV1
djoqeBA2hC3MB8/eB6vV9FDkGlTmTZWS5h6+IX5Jl3ljjxeJ259oV5CxESmMI2GPUdJ0Qdl2L/Mb
DJAO7eZd457XTc/YnNS7kyREuXQ9QTr20wq4U9xbeRnSsKk6TFT2Om7pcXdJzO7rchkRywFS5LxY
F4Bmc5hlCyemtzZj5lQ21qLKnYPtp5ArRhTFdWkQ1JcFjlqDKFfhhrL6UWdPuNSqd0st19JzOr1I
tCJXSsbwb4jpH8wwl/VmRBw7mi9hrgUuo9zVja6U9pTX+d7KNY7dJdDGe3oHR9A2X6E3vwUP0G/3
yfeiWb6elB4Lm9n/tD5KocXsNVq7cEQkYGsCJBRPKjx2isVEKPHKCPHGfWOzGay5bkeyTIYV7a7d
IrTHg3hxFHdaHkwbacbSjSnF9j+YZVXSBsIrGZjB/DLLRFZR+K+LQCs3TTCvD/VUj7L5WEdHV4TR
FB0DXIBHp1psO61Z7M0Wq6OB1C/TZ9QBVlbnWWFpxHCDHfud5gtoanOMd9DPgr3gGV3CY0CNUyRT
EwF2Ln4Bno5F5epZb9EO+dT0MRcY4d3yqIaFVgONqMSacnwZ5yDi6xy6AypsyveUP40BdbyJgzVh
Z2Y8p/8gVUbJJizcHpe+tXHch9iGIHsbJZaDdmYs1bMjbkVuHstSHegBuo3kfd5hCn3wqzJu8vS5
XxVsIl0/cgcLNc7Rp8QdY9iwuWzpByui4mGTLSHXGFYk8C1KrVD1jqWJCSq8L40ESdu9cQECCiN3
y8u27mWfvtLdofurfE0lOi2ofslG/Pt7rFT6M+HTcjpbxPCPqdjDu6RpeazryIPEi1tv23aZ84ZD
98UPH7FqeWwuJyGxXFc5eQZ76mu76OjnCDWpYZm4EqKTLSUVXvoY/bsqweH+7tPNNIpA2nzFOqjm
jLYSuCPBchRq3VY60VguW0BORqYhIyrg6vdUs2ZDQYlmkYd5kOGv3cYaZ0LothUY/TDCZ7zqgfsU
ktLl/CIxs0YtKugExkQF5dybxltbJRbBHcABacrwDwQ6st0Qgg6fDUe1ht4I8GrFwcx+yo/7Dh6f
uSN5ZWsbuqzKx10DohNCvSzwKvPF9D24Jy75wo8SFRte60cI8kHcT/O/aRO3jztRIGbB0PW+BWmR
QUUwJ3aVQo5IXfGXqhClaeKKnSzzLqbL58fkXUJtN4XOpth0Qz55jn5cShjbjQIAo/CRNxl3gDqc
c0QHKALh0trVs8qGicq57eXs4DmUYTbJG9u8JICHbvmp9DH5fNfkE3d3ED9a7ij32e9pwuTgCj0c
PZE7vB6F6GzgK/s9D8MtEuSVyGxLiywt3lY8xWrAtYvgvbFuOTIUU655zIpvqYKvbo8MDWyLZpWf
u/7t5DYUFcD86qIDqm7orT2YlJvxCNt9kX9sDXLHibdP16CxmHAR1z4dtuhCDZXH69G1GGc0csg1
mX3/iz+m624c85I1QYesWoOfn/SXOqwiqc6aqSLIaA6+77Q3GtVgDyToJRfm1tgAahXOMcPf0cDf
fVKwu/HyWexnmXjspJ5gCD7hFNbaQvUPWkBvN3mGcaFhd3hGT3b3vQYgqZQKnTtPgjXWksoz/S9x
SaIuABhUdVj/mfCPkqUtySEZoOpWQNhX7FsjfTG4ZYbnyXel87TvXpgUmJXhyMJE1Idf1czCmcGc
1Qv2iAhGjfXZdVT854m40Yr+RWpDNI5jGKdh7e53pECTATR6Wq4KtLeO8mBq80U6jtuKTwVYnAwf
tumdR7nwFQl5egJsZO/N1bb1zs4aqumTk9sE5G55NLLlTMUoelx8KL52DDyHeRBUYus8ehTlb8M9
lrvWYXyS4EDCJw4BFs68D7sRKoUtGhASodNz/vl1BnkqWXLPV7SwXa6bquHc6Cehk/Z5R/bfvlti
nvo8SMoueDn4jNPLIgBx640iWKhBS1KmBqsRwTQ1EKLdeVacQuwV/fIuiYvzW2dMv4aW3JN+OHjU
u5G9Nnw7BqZFsjfp9YHU5L7JsH1PfM+9tQv4HYj5MgGggam0zDeDBlhpheIVhLv2R+g3Mwa6REHw
fz4vvcSB558mfV9CzFfKWW5Fko4iNqi0GaFMYDyxTGMcZ6mMO56ohEy8pSgzzlZdmXEyfA8o3N0e
J6SnlDRomqjLxFiBH0/osjI9HSmb83x9C3gG61BGFo5s8bY5F0pbttHGAH1u3+EFqob1OJW2Duyk
lA3zZFkkgN/8oiS/u9M0o6B1GGhISNAnoUIlhknpR+TZoZhen+2NW5uNnNDm/L/r8XpYPPEUZ+Cs
lxuqJLlLsxd8Usjv/55scEvXOzf5OGls4H0tHfPNVlD3r5HK6lU87H1zJi9NU0gaqnMljKZugowz
zBlyMDFexoyfXIIK7gXfaZEtyebeRqOQKWcls4z3XowJA7vLJovBlTwIM0YezjJ/u4r553XRMngN
stCYjcIsSFifxwuKXvHcBY/8vD7IRgJYyN3acVhaSpeU4uW4JDCgsSpuxoP5op4ysVzstfMIGAIf
JvxTcho4yqLdgvUSpnme4mgqGJK4UJC1ZPGdYNUXtPbB0Y5tD2Cfg96AXdd+XdfGWbY3AkxTm+Px
NqGNbcY2Xl9/pu22Uww73GB7aMBNYhi+n618Mj699KSo3M7ZY9stdEG7fVEolzogs4AdTAFiVO6X
4r5LW0LK9FVKsySElFVNfbqImlXKOiZG9ZEJvD39k1wSdu5XuRA2uHM22m8Jn94eHiD4s6bWWORF
d4tMW4nW1IG3F1Y71EkA02SYNEpLXNrPnwu3ZJncHdgEf0VDWp8NdjFWZxVVVN3ZTXUq5CuaMYxU
a6SHCdqhln7C5Lh5uwF0jFf+RP80jk1p4wL4cgxjLlXF6MvXur57nAWHfY4OuKAtQxTrMPbfxXrY
bAXZuAPdo9z748euSPW3HLRN37huKNzRMed47+L/ngxV8Vd7c8tbixWEiRztsFeNNbzLPJKwDB95
/ygTDN1h4bwFA4lVuvsQXBO6FN/11lpT1vcjjDh/n9Tr94dXghXeJ9Qfz6Pp4Aj6atDOJ5C9v05u
8KKrqJYJuOK8f4alP210x8KBQTa7qw2qHUOUYBFG+sEwlNLsLL0JBSzImsGKWQjvWLIMZ0IerX5h
a49WqtFDf2T9gbz/xpVH3cwpTCL6jkBvIDLrrqNOynaTWaSovqNdwK3Oa2zvInNflAmGZxzXyL7+
Rs6J8p3pbksHy7+nbzuyeTMMuigCVvd0b4cPrqYExhWlpCsS2TEdTkY53lC6AmS8GEwQg/29pISA
CW2tqWlIUdOtH5QByxynRJnsvAZdJgZH27eBDm8hVnSgL7n4JwqARvnt4tPtE0/YA+HQMVwoFF8S
9QfxXwE9KdDeaRQ6Rx/3FQ4Av64HHk825Sn/eih5xedO5rzyhqb35ooBTOmCGwl2HmudxBJAkIDH
K/flWSGKkbaOL9cUP0EhxKxtV9w6aCNWMkZiBSu+cCmB199WmruGCQEWzIRGchx4MzrvktueGMP3
RLXL61CDgQ1yshsAzRikaMS91NoK+7uuLUJ1voVmUibz310JrymGuf21KJh3XN6fF5cn5+9gFhY7
H/xDZbj3YoOQI1zjah1Foq0pf3jqiR0N7kAgxrECCwBLEvu5MSPFd4bQB5C4QkRL9EJHrSuKR/At
c7pyWYRG2fTHF8W7U4y6sMDZqmB7iYDU5hx8d48tO21lSIrlXLx/RKfuTnp6k+Ea95dovEIcq7Or
jk9YMOXWZntRRouDT66EPW+5JQYAqQtwgE3Ebtr3vfEj2/ghT4onBZ7ir08eS83rA+bB7CglJI/V
qPuLM9bav8lpBwBeCkdrT8NDln31bkU0igVQ/PidgCkNChQtHrm77UaT5ti3uo1qR5VkXF4afpZC
54uYIYSuel/wbDK9lwzkRJUZffyfkD8ikWOofJj1RPZ2IyF0Pd5gitAj+37iHC4jk4OVGof7exhL
wyEcYFZYPBpUr5ct+JpOXadw7ap2ypRMsbco3CRWt/8QuHLt7bYyhBP9vDWETuBzr/m33mBCVPi1
l3ZT5pdzsOWLEXQKKGLnBly6jpyAIbXURWY94+qshk0OM2Fp/sJZlROGGc9jM39Ifgyvruj54R0r
rksdO0aLqIGfG/DEMQ2A73T75F8PnqobnY9tWWjBze4f48tNvJwgJILzuZtS0EDeLLyHfsBLBZVh
L5crX9hod8awHThey4efjNXajLheJY/3u0TPWD87Jvy49u5qjwYwDDNATLZkK99jVFAzpm2NRDIG
UAVy2xQGGgm0MZKUAfVm5PDAB8RLKLSre2BAwlQkzuE8in8xUBj6KU8l0ekLXe2ksWijFH6Op41r
a842I5FBdLrHtL5f0tcNsU72SVy2Zu+p4MeAVRU8LW8wyA7IxVUZmkxriUgPRO/XaMwtTWQCDAs8
0OOs7js+zGrK0z1t2pB2eFKynIQFGdCcesGnBpVJqKAohhqt37gVi6qgS/hqin00ZCCNqkyAnBy4
xFqwUaLTiwGEXG3ALB2/oN5YUzlSWOkjOXLSRyhPA3v+y8U37/HEFYL3I2mH19F0aCjFZsVIUaU6
EJw54/ll7BmbjpGmf6XGh0mCOVHNWS7IuOhHE0/A8A1Cig30cW/31Y17p5IYnqoHZEuXYjwkA6pB
i0uRkNXDgldUx4qmfqXrjWqc1uSLcmoq1LuoJCRuKOFyMabo5fMyI5/EpGsr3nNX6Knn8SPPd9Su
Zp119xk57Yin2yGl3SwhRS6V7sf8ljqmRW3Y0okabK/qxtTBZcESFQ+WzY6qC+yPUIRrzDaSXO0Z
pv/LbiVLk5txRfwtmkcFt2iuegowkdGSH1umxYgw60BibjbWMgJeJXpGRLHVgDfturhDN82KJBBS
D7Hoa+PhVJs1H2Pw31+Sd5JQPZZ0oZwtIeMolR5k8ARN0M78Gq747wmnIhYAeQnAyf/PPImhx1Ro
C+V47YJqyIrsWCIzfq06cQ9a9YkvKAUuqEYsoIeSd7PHqwCm2Y5ouuIbBAmGXkf1BsjeM1cNToBp
GnLx6ksgknuPf/vm3pY2pQK0BAZiwxdWIeEGUFLpCXB67EFSTLajs2EmkrxlB0PHctZqMu5wAfTX
94GlFXVIWh03tMMCh3gkgqEYWwCxBerqLI0OCFt+NZQcqZqV9VDhR7Objq4LgRwXM8d7sLUDYYo8
EXoRDWA00FS4RxR6RkVqzpHEKPhiIjG95LhPDBRIg7lSifWHWD/LWnjnA9U7tgOc3RDy21RSe7ei
qiZECUZ1VtqFdvpLssrHyssjs/im3D5HjmK26hj2AW0XJheJPkqjmFdXmkJSi5aKBY8dCcMjkyn/
AVSRRVtCvBqD5ER+/RfrJIPTGMgKf7qjmEmKvoGy5I3WLbuye49e67Q62RGF72MEEdniWaVV0hVd
yp1fX4v3P2K3N/AK5waH1eHtVVO6+DUl4SYHaMcJnvcbHyeIsJYWNM8fjS05leepBrwQvOAEZnye
XCNTTQ8TO1Xk/eMpm5jTTrvqEsiErXDVBn+IqEI4UNZW5agjLzYw5Budl2YE7RUkOl6hx4DcITfR
xY/aQgjSUnWbLx1yq6kb2Zadg+rQXRcOxvImjibSvdZlhvopkWuGydFYSYIivu5M9IHzHUpK0nxi
0B0RLN0H+SNzPvtXmOIpQpHe/67dbseWQu6qf4DwGoLzIKhUjNulJ0Vg7UB15WLG22sJ+rMjIT1T
Yf2qdUbxZnPG5rSHd+M3ll8bCb/AbfTJE9+wEKQMD0MAeAzY6CKpYy+zwtKXblSG8oAM4mFo9FIz
oMsA8QjJWIihveOgf28U8jJOWwlUIlOL5fkgiLl6yEt5ejIogYoS1XF17aiHaTAxB88pZXyI8bXX
cw+SVK5frU6UeNi3Mx/gDbRUrtHWtHDs30Uc0y3bXEZRuJNWSDmlx3uTliYrp87O79tCCaRRwXVW
xsftKaTRMdP7rzNPWxHaR4e1CXnpx43nDD0gH5KTARoejQoHcc6j3CpRwTU1ZR5DLOFGpaN/cAHr
WnUwach/XaVHqORTOSKwexnAZr7b8kc1kx6DysqKrgrFykgQNwc2QStJw6k0WCl29nm9M0mPtZCA
AMcBVF8W98qTygFiRWitGZWJ8NwYldWrBApxPnAl3fjM8PYt/iey3m/7Zp2z0HjgQX5CRfj4MWX+
XxkPcGCRXlB41Kp/apgqWjtyi4I9gmjtacX7XSAAi7J1SSVEeP9Kk48V84JtsvV73kehdijUPqB5
EPJNMClC3prmN5Nt12/pO3jSJNnJb4g7Cl41dNg0sAN2CD7NO4TmisMSbTJeDfiYOuQ2eIntFrOE
W1ffdJfWDa6LfBrqH/yYRNAao93YFopmzcj5aJxk65LIGmrNXucY+fczochDo23qR5lyeqgcJU9s
DgWzlj3lgKBv/GDt8EDLCX1YvN24ejj4TVamGyRoAgrAXcbIDZmysba6h0Jk0GJUCNaeqatGcggB
YGDugzdiO/uA80/JYAzhcKp0+FFa8bv+UOqmrDaaLsN5WIpVf20Fi3p6sHluOTHSDt+k668hJchO
1I4RiV9LSxDsl+eoBXhw0yOlQcdwEsyOHJGqOBcGuoHVnsr/TdbWd6KXLmV0uGsoZZ/ywtuYuOHe
Yhiq3BIOdShZcSL55uVlCMaLUjYR3LGD74v5dXpgN8RBWolqWho1OIjDKuH+aMFfpj0g+5H+sX5f
+MNFvRYSaNApsuVaD7MndDlHzBnfptFMrGJBIyyrAi2wO9ooywNJ7ZgO5mqMvVUk4L1CrTY0kIpp
r3+k49weVla+6SEcAGeWinisr0uCrZ0CGOes0msQRxY3orjjgbvCI7Kj3+hyz4E4DcnEisfbZ+Lv
ObhbaKvYUpeLiLKUzjAd0u3BqFWBOheF/LJdlFWgmiOfnV/KzKaMtgZDikoLyO33UpB0aUF/Lt6s
uJSuPZ6PNeAM3gZBfOUeWoXbncnoafHQ8wy/+Pfr2wFf3g4L/uh2aoSuOYUJZou4MzT0CdRjBgfL
OKErktG9EHSunaPISnwsb7gnMB0wnBSJLW23dyhStkhKJ7BEzHCPxqTODi5pHfepZnUljwfHpyPw
VzfIVnN6LTcxkdd8vyoKedjqMOYOWRtFudtZEPCvT5oHuoGEjnZ32PrTZvKYbQpsR3odyGzMSKAC
gsq62H9dGojcZU4h+xlY7zyHYEprl+JxXKP+fTvYzL0tUGnbd1sthpLHFh9RznCf7WSBDAlv+O17
gsBfCjOozZqhUL9dVzHM/QqAC9rNlIalY90unar6qqejkz1xvGynVp0vK/d+JUKxOxsL+9kt/oMX
HbFNdBDm5jvR7Or6/plUZTHzhiAS5tMABvyIEolxOiJPOarFgASgyxwbt3yryrLmiezJu3lPLaY1
EO38wbntzS2T3LnkylmzyK9dWAWjh4XIbi9FqEBQj89lwKp6b8rsIDEfWJNVXrv6pEHlYKLrC08G
k3tV1Zq/oDA2jGJ1IXiSkPxp41qN5Xau0Fc9eQVhqpPpgF40HRoJVsKc2uG0raYuvw/OVL7RJbjp
NRqBBC4rOIOBNe9gfHnBBFk8yuxTtutlzUQL7y25rEuu1kJm3O4mf7FKHpb5g94FMiJvm18vIvby
Csd/xonyLLoD4O4R0Q15rTsqztwdaHJmkkH0wlEclXQ4QB5ZuraZwrNvwoPtzOfHKVrEYAIuRr6G
/8JdczR4QIK74ocXPmF/mT/vHM36aR0R/zXHuyusrxsH5VXDpXa5bvtYifnNk6mE3zmYqco7KEhW
OAdofboQ+bbutHX30DaANjgN9kufXaL2LxhtdHMWvEDM58yYgHznpgolzCZG0b/HqhxJoLL91Br3
nGW2Akv/f6XUVUB7ORnvm5EbMRQi/5EV5akuKeBMAp0MTV5QSPMaUfba6vERHysckDak7OvgOpK6
YFR29fl1bHYwCmma5+uCm/YGps5hb/mMObfYvlEk1H1j/ZSItVYnkpJurAWIRlV9hvDPELUGlR8s
09W2ePOIiaG0mDa5dQNGPGDg83w2i0gXsTVo4bAjg77DOllS9T2LQMDBRDSjSiiB5bvPqKky+E0A
vnOGJkg2QkqA916OpG6bSce6QIkAciN+pmuxJHiJKw0X4BO1H0aJrU6FofVT4SAuB0Oc1xNjVENl
OdE8+nkLqkgXLWxPVjXMPOkgKvgitpEzlKBzs0UMkVL5X5lVKCDfow/eDw6rS2CYjkpjiDRXGg2y
ubed63XRc/fknz5bsQVBBgX1ixEXcqGw87VC5aAW4qFK7zcvyOWV1Vx3CrycvhRmnfSkl2vUGjxa
dPTV+NErhPKibzm2BCWRvObJP+7qSMQKH41LD0BT7bDDKzJNG1RMhqYB4MkV8e5ryksbttyariz3
grOt8JJYPk9Izll8C/dapCHM44sj9QOX/HTqMduEKt3zPxKdDOYJHa22p1HyujAoyLl4OB0iMqNG
SnlfaJZ4f4YVfNx/f5KjqrmXpIzeORxxazLN65cHixtDuVDU0cBkRl3ebtCFsldFWdrGvjM9yqkc
d+AdMGqSQg+2q17cvbQ3qCL/opwhMCrGhu5MziZsFGofgJYV+PJa/WsdO205rN3agnnw4eulTC66
h/q5H5fz+lhp7lsMvnHLlKH4cbetE8wNfuoGKDL17bzrEYAAsb6/I3iF28pR/mMHIBBJYeCaxoVR
SzcBirfgDVXLmwqicXGhp+cx0U57XG4KZ25sbBONAcU75XvAJd8hHfVBlUmu1H6XCs18P0Xl4CVP
JXtDLIrkIPRzHJzBUvaVZmRXJudqg6QIK5oDM+YBqSRz89/tAGWd0XL5DDyyoiFfVHig9rSeFP5Y
AYNAWcAByOgItCPPvSsY3u3MuHs7vsaO83+RVPMjtp48opJsYXSHOOlkc1Ldu8QXQI0TdRwGCn8+
JSOFTgHY+jswAz7JmSljcJviBjPgXmW4xWVbEt7MQabpHYdYacAhlIdjmIPR/495OaCZhMs8LHcR
2jHM4U7EAOCu/AL/4tEX07gNaMbjXjtseZcePNrwwWV4ne0qiP+fP/eHTzBt3zNufCCPlxPt3g7b
yQ6xQoRK83fZ2aFnnm5SmGrIoWfcWB2JuRNQwb+6EBbUyIXK6BYTrImXmjGr1DNKwenMqGAkV1+s
NsUwXq5UQ49pe5HreF1+rwoG7J++94UZsJhEblxtbXXmv5cB+JKEqIeTe6kevYDjRY7CWUQThZ32
a8pGRqKKXoNIC7fKbW/SjKTrjXvxfN2435bjJnUJ6UchMtoi7oZEeJakSpHgAiB18p5vKnRWZvCa
qrjILUmtER855exfp+gI0jaHbUwvRc+N6IaMnB1Dm0kEUpA1jeAcuyZyODVgJ+njRVKZGpBOg2yg
nau1bQqfHhzcnSx6LTDCHiIjONLTYZXQfkaine6Hqu1GT6sMNUmNqFSurcOWWt1waXApC659yWAv
8chGZN+0Qp+n573cy4+QLAxCpMcurCVm/h5OvyHq+SdbB5ax1cpmGfoNtUBHZ+izc770b9S3L/Aq
BshBXxzjCFuo3vyd9wiw+ALEnYhDyl/mg87O141m46+JSM9712MAzvdi3Ry+tMiYwY31LsikxcXe
gt5Lc1QtaQInBeoUYjncfwcyonAo0jATClRCGWm0SHCl2XwPrLczS47uh1nJGawKlpkfsXY0r2dH
BsYcHPtriZ9SPH2ggiM1s2BWEKyvdm3Xr/y1Vyb80ObSHDYlwm1I8zsuVYP1fH03P7+OX2uU8ln4
CGSJIyJNM2R/TAO/ucr1580rIAJrRM30Mb9BX9soMdojRuLtYdXH+pNZdZgfbPLjdS9PI7o7ZqnQ
Y6Kcprcz0VFKuPA+9+ORjN20DoM0MCUcRA9Mo8sI9Fvbfd1xundayGiFSPwpAHcsd5PAns98VxtW
kO9k5is/AEYoaF4x/zsFaSO8JybSqHf7jMhnoRLEphraObJwTZVrDwME4BzDT0wqmi0JLpU1jsK4
FHuIo+rbIPUvuvFev0A2+by0CsrQhMdrr8G9gWFTeh0ra77d30by9EDi6gp3UIkZ20BQtTYj4B44
78cnq50k88VbuuqjWx0s0gXt9pH5YgyWB11+EJziyLBC9hXog/kAQvZsacmWavp3Hk+8Y1nTK32x
cwM75AxcIxN74gDup+BBU9JXd3QogL+UJOsQ3aiqypbxj6Hpw4QDNZMyuccX2DnRnvb80iUSQCCh
bDE7b0dxzSTkVNwDnwLDb5CdMW9dIUilz3Bn5cSzEIIvBClTnqBdvk14q2n2snuH32pDnBZRLcKx
4HJp3ZyLlZTueWv0yoE3+P2Mb0g/pSRvR92DDvP6RGHPChK1Jo1Q5d/z7rtsto31ko2kW+JO2y24
GFOvbHjBhYUKI/5I8PxJzFlaZ62k0xp8hL/OVpXoaIpcCWxHN8QDwAeCn8abmTzfSOFqH4R3anhp
qw5H/+CAY9COKGtmnI9psrQzSoRcMRQAyfukzP5m2rIyj8EHz0E2XLKAKwoXwnzMPxXlQpgrCq9r
ikC+TvV8SeqpVyX6iLzXOFevYFAx9fHU42owtLVH6K34A8InZ/WoEEFZwzS/xSCFHDtuyeVmSWt2
1SCQgAhD5MSgv3bdiqAALiNZ9B8f0StFVrVU9giSALefPricAkvMMvIr2tRNgHDokFaHQmFbGS4S
IwfhKtm/bwaMLMtI9nc6A97tz+0YvdqBJCYbTmyFY/6NYut+3GfOwvadvwlkw8odNQOAIDwY+Dhc
cvqGTrkU5lEtC08jaS3/eHTTlcx7Issiu2FCd5TR0qR8nCCLxk0lEJ1RN4RtOLqDDmtP1q49ERqC
mrzbUxM1TyMjqqpoUExLuILg9/qYkdpPribpjeconqYkuHxuFIZ4Cwz25cIv+hMLqV7zwDhS08Tx
WFmw+7d1hgOCv86YnXvmboxA0p1NBuARaoaWnVVyUcTJQHtJv1ocIkKPEN7DStJtMf+ReCvogQrv
N3Rj0TOzqFsAvsPMUNR4HYgEpO0rmYudMoo6z8ET8ZnGAzPkzU5ZKwrbI2/Wx7gJYrlXf8mBj2WU
ClQ1eZCa6uUO2Gc/Z4P8poFox2swRe5VQTYnXGXq/QZf1I52oa23UOm34S7IA07jWYgYhOiz0U1r
D9z9iexIpi+0NvXG9dlZrIo91Fh0UG75XtKkIGndADArEYWzmQ8nuJhbpnfWCoNbw9lJB4gmRE8r
mYt3gXe4mWV6GfEJidzzBf3vcxC1Edc5pvWwbksIRGDNB0GlIfl323eNqMFsu0HGFKohr6KjvTSr
UxveplR8gXUzynD8rRQ6VlJA/RmDmCmPgKKJySkvslRJexwJS0jCPiT0tIE8VDaLvNeeuJd0DOGn
Kqlb4lgRiPlGRDoThl/d50nfujYcdw8RG4MExPEIuMv6LqNTDl+MCmz09s6qW2LU+tomDvADPzjg
5QQs8QtuV/TW/uFycP3vmVAgTEkXxJhN8Tw1YNF2dT+Qvo/14nxqCXZbkpipY1M3hUEx3R72Wsjf
ajyLPY4aYRvGBwtRKLPTXd13tTRyVgqcnBeyTCO/6e8tO1t7mgoanBokvDtCLwAIJdcDpb/cEp6L
/DhRHwmM0sQK2RLl0jOl2u0IPKgDef/GomvXl9DLs/+R7PqZWpyijCXODW/R/hc0yoGml1qz1mrv
bd1ytGX/xN2cbWYiUIsItHGTYOp+ijieKwJ4p76HM+AwyCvWETprkw9aTAD2z4GVcuqX8WHFLVkR
H/Sf5xEef6YicbP11QDvvlKSwBkwnclXgJqX9OSC0yX09OsNwj6A91IqITVLCptu3KS7nkyr4mJW
fyo1YSKDjb6TL691pAzYyd8ahqk3cYrUW41M3MZ98z18md7Wsy9fxL04HJW6cdlfLFlOvbyzBh21
bT8kFt2YGuo0rWOP0D2sCJVEXnxlETg0JrfKKifSvgGnn6xIAJY1e427mzh1CtUMusEJGWp7w9AI
CHDf17AiVVW0wOsVgaIMOwxttvuhEfduKTc6XR63V362alrauwrvEClFcquO6QA8jSeNJgQekIdu
d3xteDc0TFq5cG0k37ToBVXLOHm2AgHxoSQ8JMAYUi9Qu7CSN0c/jRFsDcIDKisKkBCb5AHrf0an
9DaaiT31xJSVTHfnDoQKW5vj1uUhJpogAnZI7XTMylLvkm1hHQwQy0T75CtXikfd/tJ0TXwHMicv
Mbqk8GcJ1YN0f3GAK+7XgfZMTwUecuOKJ3EWyqRveL+R3olD68HbZDwn0D0/9XlsPjkTeZXnp9qk
JmyKff+yPZ+PeRB2uDGRw5GFBZYrniHd0IdvaqcCtE2mJa0CYnWtfa/tXJzqS8Vfh1fLf93yyMpw
Y/qHkeofI5CDjE71p6xQdeuuTwYF72R5oXbFrSYB8nCRqGRlmWR4wGY/MfTRWq3XmJ6LoZ0t/vgd
uLqAdhtIgmEQvDXDDz5f9QKz+vKmqWBpUH+EvCF1KM9HblG2ABE8roa8vYAniCSK6HGKT6EiP1nZ
o0Og0uooeJuWceMFLCozON2ZQFO3KhbgZOR+fstDR4GOIQHNZZj3x3nwywWCTpnjww969A/Acb+M
QKC+x1loczzRjzCc0erKe80zEXB4DJ1fJqUmjMAf3dXUmiiDKyjFSgbRTMbfkjUw0KIyoTr+D0df
EIv3Sovfvrf9coCwGMldFEyBHvcUJ4MaPeSJOlW4dgvyqhXFFTFaHw9CgnXZngBytW8eZXngfG88
zKAxRUIDCCHGqmfurGFLPOjLKgoBWaWLPt3kLVTfmjEjftrOramx/NcwFJup3qk4M+WlQz7joJAj
ghP/6EEk9rjVaCUSHb0iVqRm0QLUy7av+REpCU7GUJ/rmM479vvBgBD7NtFtwKmVUlI6m+O4NKE+
K0Ion+J5ra3dmdFTHY6qYP44bndDct7FdqTOk1ebtvMgqafcKcAnIxl0pZ2IzoZOm/PZ1ifbLWYt
VN2B/arAbAKMvRp7Lyk+hqjFxKgNSKTlyH0ioijwQGrcRZkoRHaEeKl7BeFo7un2uEpY4nQp4bDw
Hd6V56pi6rklhwIVU1J90WAI2aGxqvpxc/Xm87+gguU0moJU9hRrSjm8YVSFjTwcaJTABpKo6kcg
4I4rvIw07IKQLjlBfmKnwpRf8zfl5ZkvgYmKL3qn8D2jZe7EQKFj1XgSCylx2D1kFA82gbIsWSzK
7sIu/BJwdjfhm+RfPElHUzU2Q875L2x96lFkxgTuPp3sfga8x1tZUqoLttZMiD4deAEXP2ANE8Aa
wztSlFVVvHrn09CVeFAFg+tqH7IMHY5uCes19sYnrZ7Bg3hrufuzWSdZkXdA9odtJhH803p8g9Bq
ctY/cn8kRpxR3gesyrlOoIcsvDqjbtNGrZelJ5Qsn5+eKhGIKLFCAB5bcXY21K8ELzdU/5y4WrI7
2/YDMorFovAndoltCnX2RxVh6OhxfcL0Bk8AiDnGkoZHGecAQ+cwcLkpKnVRiE0YUpn3JKLZbx/5
oF4bozXaasv17xkEpTK/Lj7gWD+JybCT29BooWmRh46Te6yW20Yg4xlb7UeljVBpJqc61jf5uwC3
5RbsaDVBnRmTuAE3rmXJxUp51rWHcaiIPD9tN9Nuv64dWDRkr+XGh2ptvuZRFJpFaJFvCW/QzM4n
DU60ENa0ilgs5VDfTSBNYGZwou7PvwuAC3T27IFY7VxzmdmeQX4ZiSoepkp5suO9DGm1Hl1IBLBT
6Y6Uml4JCW7nxJvr1VIVy365O28Tm+yK4CJom7QfVQb1XQq9jTlnaf0XsGeAo4v7mrN3KEaPkulJ
YlEKgXAC4IK2M8P6kGfIjeetW5HdXhduhLbTwXxfFAygaEglX0LuiMhxqerP1cGwWiy7TdcHt6Bl
x/d3MbnFeNNwxgOTeGUjMcTTkQ/mgisBhlbrTd0uyqD37BQx5WPVi1hOaaydjesM1g98RgpyJpDI
VzVRo6QMsRc89ezQxdcB1neJ5LDux3sl21RDHrEC9poWKfRV/PKevhpu3a4WqYRwNWYDGoL5Gjx5
wAjusn5tXTncfD8zBffpzEt+neGQESKZeOjIBS/sJSW25v7O5USEWnXCuooNZvxrN8F/H6pC0rsp
XysVskdK+T1ZZVr191Hg8+c4SaXIKK14xVlmUJGVjKEVKKmzQidM3J4drZb+Bkmvqdq+nJJCsGlv
oCD8kpPiEiFyyk+Qw9xNXyuWbxoWwjFPHwXsOvSUih360mSNh1b6DhJaCA0NEVwvrYtlppjUwhr9
biuCcZ5MEc2WFj+8HZxG4YXAP7fKI8pdWXf2HEsdzu+tcS2toPsBVVWxfjEboJfZMerk8FsarnWb
i2KhQLIx1N5Q0pv6DMjwHT2Z0GLFM+G1PfN/x/77uwwshH0j1yA2ttBWV0wW3QYWz2+BcXshSZlT
PGHF4xza6HROlGeSYJQ5UL/QSqK19dPJ7UMXsKeLvqGbWS3UM1d3LT8qwvqz7Cxer/lGzqXd5kvl
AEvBxnJoA2ifaEMocbQdcijNcjeJTypgde923qarWcjB4mwDr+sVcsqAjsZCk+QmunoVGehCCIM9
GbufjrBuOtmqPrqD4gPqW4eeDxdbO/Wkyov2nh97Cm7GuhqVlR+V/7WmUk4KzrYkRGaQtVjA2lpu
YAgPANOsTUjakoExwrFQdY6beZdRrgxpjGFHnF3YHTM1Qr/pZ86TXMHcQfBdVvQwI+EawpIfWuzD
m+n+qoXoabmBbn3aQdaeWGan7qX1q77STm80FMrBwFAc03pFHyok4T+yfiFnSeWfu4v3MFDmnYmX
pgayNUw0FDhA50HUw+9H6jceT6/aksuKHxjFcoux4ZY+btTxUptlBpX8W9jTCSroZSTyEbF1gA1D
kMI83fjp1BvkigEeCRMaSdAVOJYk45B1ZMzb5qT7xcGMFL6uxvGnNsDZR7rm1R8/vF4Hb7iLmRfw
vzdyv/jrXTl6scDgp95SD+8DaC9FyYvRTpZxb8BTSD/bWbTr8YgaZdLFqtnsQAT8CWTjlogYgNZb
n86TbBcsNxK03EKIz3eOa47gIaHNHuyH54QBg9sjVx58ffDD31n+Rp64G0e39LPJWi0XvIwxovkY
v/yttiANeEbkIbglMbHMpm2bE6pWVgs0uGeaHMMnd3LKOMMKgVZc3UERUJZMyzsikXiPdYYyUflG
N9Jd1WSDTXHBsLYZv2u1+PyJnn0ozuRm3ND3eiX4YIZjVjYwBE3GS9aEEiVN4qsD6iM5v+9+aDFM
8DXYXYfYoMgcwvIRGFSpgIAAzi6RUDm/X0AGnpNl9GQnL/EsfvL+NMHO4T4FOqc0T/TL7dZtjhIZ
ow7AYP19E67/uS6Kl65LF+mo/MvYo2np2qUuzycoKullNX8kKXW4HnkQoKK7uURDY6eCtIyijV/B
RI1QjdBU04jRYvc85vMXH7Hyk7uNqqPif2iSx1kBaQJAKn+HBRfHfnNbXsSbytnqEAduJEOdsEpx
p2MRKMP62thJtJe9E5Y9tvFyuTr4JcNH6SsJt8bdKV7rmZq4a1sKBlFdUsvYCjTGE5fbX7CTwqY2
RR1BkLDlZzeGXAPz9oVb2l4aRIZO774iopxO/zhZ9J6cXJHVl0w97hwj5YCWvExT7+R8ZUYupW8M
85llQTBvlw1rDEFShAtZe9RjOIfR21GhV0LdV6P4rpeofKhiCBY+NqC8V8x31k+Mn47hQLEiAttI
6IRH7BIYl6pUyNpuKLgg+AgsQ7SjWUR9IIu8m2JYAIsj4dHNYLRR22V2hyZSAHPf5ZP6nBo9GKpo
B8RGiJLMqdWA3BKvhh1v8iZWSCB/wM759RkjuFjdPannCDpiqi54NUK3AgMC+Za+nE5j8RMvhX4Z
iL6DOgRSN8DhojWlokZfrs6IRfcko+Ug4NjaWZcpLKXApyrJiKz8AtX+H/pEbcwS/SwQDPGipI0w
oWWBcrD66/Nzt4FpIZ8aKBnLB9kWQiOe8Pdkwlg32wIi4x4BAu0+hg76QIjNr2BV+DmgtHcE5yRA
u8AxhHp6cIXXtEwvCVsWV378ZrpV2Zx2qJ9LylLm5/p5iT+E7OvCL7xKAjnMbCQs8FgzS3rPHE0L
kGHJONjbizwa1yt44PvJ55+vv2fotr8ugnvqoJi7I8EPBifRXblsNgde1R4JZAKLsm1OdJGs0LwH
RJR1WmhwbcmCV+Jt5uunSC0HstKs3Ai5DA/5m0LplinDtqCH1cqbIDn607RSZd2Gt9o7aLbSmzop
Et63k6gX7yqZ58IObLjSylEPpW4oiVfPbab1wbnv1/+3Pt2vLglePwy9JvM4ng0j5lv9XBqhWasB
5Msgc5jiBnZjemZ0xfjRgM+yS2kk0hja80w4pgoce+GQSlyXMEPQi3+XNh8ADrRvnsHCvS27yPVH
dmn2d12jMLz/Kpx54DLf8OQ1htSz6IIWEoiZDfH3ONUoCLT/rY4pBxJgvTQKkGrViRz/Sb9bZVUD
r+YiOvPH2dNTOxiQEQPyzmBiawAc6ACElTQ54FDUtP3fi/uhxV4gRv+F+pJsMzwxUvgEi76CNnwR
4q8Uyns5vK+DvcS7Ar1an//uxQvtWdDh+sSZc3jxZIFhHtTTj+B46eX7BWppWPv66iVcEfm/2T53
hQNnYyNWed153cOWHe8YAnmpT6Es+h3qr+u3Qvr3xeQhJfNYkxD4maLNRrNlcWr+uIiQmtkY7GTT
yPEhcKAi1dZPZ9o0NlTnsVEHa3OCrwGOHzgefX6VxCEhC+HwNgIYjWA5DNzGo/cDIKsktkivP3ou
ehRsoyPZzQOKSs8NSXlXkk1NVf2yE24qjcAxWe+aRzHWC2doC+s0zPBiQlnlIXLbwdseNRdZKRMZ
4gVukiJv8tv7p5DdKfJ/6szTUWnHbJCWKBUwcJIl8HAfDcwjIao9N5R9j4tveKt4BqGkC1Y+XY+1
NHjyz+BXJN/YodNOOkRvgUu//zxuN0VeafA/8TZMmM1U1l7et0PvlbcdX+IWW4vVqGp3NiQF8aVj
VBdvGx115CbTK4S1yAver75SCWJ99EYm8oFwtaXkwcMAUIupy5t7fKeNLAc5ithl7Hl2sdcD5EFw
7Jp4I6zQaRL3xPveWzU3fs8r9eSi9ULNByLfvWZL/Hpp5NG4Kr2G3RVdZ7h1e0JDMc3MKdlMSWOX
xsXMrso0IZ31/2zlOya7pqlpHh4HK2xdvUlQ3k/CcrIrf0hO8TTnBJjjI+YRdtVS1blC8TtEhqrr
fpmbByEOVu/7biq/o0T45pgC7a5lolMx4fyzYFAznktVi8f5MJnPZ7Rx2+r+mt5Wtxh3+jRuHvxm
RudMOPqt+uVnoYWkT/GhztyzksFOGig/3FHqd8NSkFwxKibgTOGq7g1PKZ+Q+oY8iDcMFVyhc+YW
8OjtBQCFBbLkgQhwkAxRG6d0vXOkeC99ve74xVeiLrwaHPPTDakmwjDXfjrpuhLnVTK0pX3F/Avq
mUXMITd7WcNY6mW9HmVkf103HLkFBKlgQuVsW/HEL8JrEVyszG59e+Xhio4l7pMovZSRPK5Vm/QZ
BXgAwSBDBTNrqpzPLcruO/pSinTwNWLhf36b0xLQ1VuicZFmkX1jtuH6hpP8yymdEYebk8FdBfWL
RuypqfSZcUgwvKm1QGjap/OvGli7LEhlpn6OkR+/R6hfUIlEPCXgl6BAvJPeKzu5XneMeHonKqtu
z1M0UjEfCEErTjp7y+siiJL6lSqCHZSdAsIld+lrA8isXDCWrzDbs+zSM/ByQ/QSrHNDBNkfaABe
u4U7AvMBkKuSXdWZpENW0ebgEoCCD8tTgGn7jAZQ/2/zSxgp/+xwg/rZbrUHY/JHGXOcKjouQGsg
hF/iLl3IjjG3uUem+adEUd9A7AA377WOHjfMyjb/XhJa1SadP5mB6YY/xBUP3n0lcbR2CE1qe4eT
YRQFpwzKpBd/9hwZp7PaCGsvJWAkzwAkSmi0G5cz8KYkeaOD286PZYQ5ei/bihbYBZlFFKJ3N3Dy
3mcf7+J6KBvPmkWDkitcQVaGWRUU8rif/nAH7vDwi5L5cEd54kq4rEdwxx/PCleHvfehBM2f3XFA
qd6O2EKoxhVJ7jUom3otXtdolGYGFAgZHbkmQXA+GgqIBl2eEaAhDyL3Py9fxE2QCcw82FgcgwXH
87ODbyWTFCmALB+VW+dWaHTGhGdvG/sozIyTWF4nunH9dDzyECT0Q60mfHxciLJmTShs0vM9Q+PS
iZ5xSBKdltWD+uJ2lbiGa07WSNDraqaQvdOD//zzrwgXfR6XuFgqJURNObagnPZixIESAVlPnfOj
CYbnNt+SKqf7MosUCVsVIyaN/ZjfZx46A/tvSgt+mm5LUqzEfyJnrS5CRGZwIAweUavxrlzN7QRo
oeiv7UC1nqXqJDCrcLegfkcO42kgDQIV+SmqtMJOHGsIf0u6tN/qTf8C/svDriPG59BMMax056lr
2u/7GtWuGhUjhxr7S6zE6SB7n3t9drRnHAixV0p4/sygqIGR43RhY/xsHoYXHigkfOxqXMEwgCxs
bE/5CQqq02MbrNP+4m2NUjWt0cNDac6/AiSuFK7ssh/LPAkQaCALad5M2xRZsnuS7bjEDp0RBBK9
npIsXEeqsYYz6g1l0pOa870NGMdWzGvYybafM+fBB9t/m65yqsTy2SC8OvGpzwPJDmV8kTfV1B1E
4jKrKojp9ORmH57fmvXvrMIcrtIAfhHi9hpdF9sPpd41lrCw5oLncv/bop9EUao5xSBwWkYaFUHK
PsYYqhI2DKGK07d9gxTzsE4+C+EC6mk2hIDO73F7tJdPDNLmle/0N0Pe6qOEdy5MXISaD2H5usSb
gzjSXPsRsuCXq6Kcqdf2+/fpU7Ae2qj9yP+hDSoQlUcpTXmvpodbmhqLGzE5sCYH0QfGSD8olzS4
+/kXHHWV0DwxyvayrS5yR0PvjS94MQIRq4C6fSN/buWIJ7t+3b7LghNboY8pmjTXcBSyRrG03PRA
N4bhlfsvLYtHSAla4W4iSZ7C8rPqktFm1yF4rB+/FbC8vhr82xlD/C7tRu9djRo6sQm4fDKODULB
AUtyrTaf2XaQl3nFMc7Ig8yj54pD2NrNfZTJME4DVtpVVx+yWcRKTvlJ5ffXpP6bUVIVJg1Syk2m
hwzZBEGTnWzfuBxT4fzqbrUAg85x5GTE8vhCf6yeJlv7ZjLBh3B8zFGp44JbiBOfIs/bnS+sCVcU
phqELmngcrQ/b/OgsSqrYjkJnBGoIgtCbFksp2JHz0C7Y2ci45efW6zzDG964+5MEd/rk9gNmobp
ay0maSDk+ypmbYwt6jpXjsCuHt1Q1XrPop/siSws1IECGymCOrkORsFIWaUYtxwfiNgKBLs8VKym
eygDXfTfM5gX3bnNTuRpQuzujAsV1N2MBukMtUOrXhqVoNxiDSiUqxcV9Khl+6HHcqNT6Tb6+AK8
tHAqWB53jR28VtCkzt5SAON+VsXHkgqn9LetCcnOYIItebQl4s1u0hMPjRkgur1NKJ9/Z/EEq94Z
aQHDFDjc1MvAilLMbx7A4fEUn3HpybDUgV+ZMBSera4H//G7Jd2MRGFWnDh2lMWAZeXw5Fp49cf3
YIxxCVsMmPCMpB2dEKMnOWpIM9NEQZVA5abarrYPyfTu6qFktSxKHD7hK/jyKs4xPJ+ANFECsimF
IjOVH/0kCBsqrZrQUGxq6XdVGJtsQ4FufuqVFOpcMIUd2fv7Oh9tR1x7tgBCdTNBEyKyhH9JzVvH
osOt7M0tiEcbRkyG9F1gO9gvH437V6klmlcXZyFwQ3GmYaiiGUI26dTOf1jrorFX/qUq+zqVhoOe
OXVXFPT5BAXQ6aRe6nTOQ+6u3ylvhHqEzukWjXK4ftgq2UTA5Gpu7lAeCMQaJazqAX5AChX2KG8a
SacaTAAELJdBPS3Mjor4l6ftEKqLcug53cHf4SYEbRTWCD+eofgS6h+S4nTlWGvsRQO78uckKMng
HVAAp7SgvapNIHtmEBs1UzHxcTf3OsGjP9gQZ5d3qcI9L/vuJiV9vvFvEFqjXW0aanzNeRGwZHyR
+iTjYWKdjw5PbqNOW4vBm9v1r2tRZuooW4466VNART6cDO0Z2BTnxf0sfdS6V28mEMQ+PLRq7A4d
1qnVE+ZXbzQwcHJMkMI25PkaiTjKQrPbSAVlCr3Lz1jNpZXr+Ze0XopGdoXi5aOrq0N26ce1iGGI
ZRmpOTd7RIRJ9C5hWz8vdPPyB5UWAFU+lbQIYVCEPPFRyuLuAre71b4IxFheqqtLfKQ2eDTZYO0m
nSWh+RAXQVCAmmAghDBd6e/y2BJsTntCY8yYkujfsCiqdYtIH9k+oPwljHyKhZx7mQfqAvbT8TV7
Gqle+v08rTihMo2Cx3jRLmFdH7e/WkbfHV6TOvvbkNTapMwfv+9lKngEmiaqXySTxbQejtluAxZF
4l3cK8qLcrEWKWVZroK2DzZEIx8V+G8czy4MYyTlzkOIwl3mDXG6PjrtDa7BR8nWFEPERpUu8oTr
P3hfPUwi6aPRR9m2pqzhjTPz/kDYOssAqK85NlBcJmlsB94O/sVE2EZZzFiWv/P5vNAbryn7BV3s
epXjCh0L0ie3PdlzMTa8JjYJHtxFQ01NS3RUnNHwXzKhAJtj7FfFL0sUip6YzfbmyxNMmI7JSUDM
ADXcYjfWJNIMA0cfyyrhThMrN7msBUl2XK0vkByQTeQVWGgpt8z6hAn3U7bn+8y60DXYzqb8iUPc
e8L9tHcX3+vYuOGXpTIiv4SMaExA691U5WeWTsFEde92ZBFzedsan8cMzgSe0yy/EEY6uBuSmh2J
ISawvFBjCFp31HrxK6r3URHR3/G3cPBfjP6LjDGpd7oORa9fKA2xwLqhOW6TsqlkVPJAy/QbSOR+
tkwg2Qx5T/ErkFnalmdf6i7a2zXTWjcQJTniO1bdDU8g7Y74oyAtsyRmMt45rH5zv7fAIjf4L+XZ
rf43bUmb1DU+/HSR9IiHYbxVaGBw9VixUMJ7WOLvTSOi5nM0xxJEuaHMmvqKUzOD5q7l7wGD37U3
aV9PNTXvtPpXLKvx3Ao+bPmKG++aymuxzxblpMaVr8ujSQF8ii/1FoVCyH54MP1T7UnfPA0r65HU
9ue07xFRzxqk3F4sAGUjoM/ZRnaRlJxQEcEFfsY6dW5LZIV+lBO3h5F7be4YMJpUX2f+CWqaR68f
2Z8EG770+ai42HucumqQQy/AJhNwQgH4DEbXEkTP7pE2tJEICXss3TZKcMO8pVfIokhXRIHBmDmg
urwuo0vHUDyWTnlpgu2UQTA+3xPeXYaRZkgVWUDNx7+nVg+FWRRWAgSQ1aL0mk2hoZyae2kZ0WOU
ZwDvP/rxQmWcXYXD/F1d3Be6js7Yx0BM24xvnymv0v4zO/3o6POysrLHFWeYttZDcqwDCI24uJnW
ge7UmpgAtgeBt/SZpIBY3bIkEPtx/eZRs6evW7H5Sg9GNanyBg14JSFp5WOR1diserLD3xfulUT1
g4G9iJtKsqUF56rQ11lfGuNQ1iksRk4+OalEsH+N05AD0CxsysoDdEjCD6PploBbxuqXXCIi1V8r
Xs5m1M/b8TYliXy3rg01D/lXX59j1RddU8e0KecoTea2uNQr1kgT9V/7GHbG1r4qMO5Kxe6l+ns6
HUD8tptxKIY8KWCIjv88T5cMuBf7nrZ1BnUYCGveOJpeuGMTZDfjidfeWbk+Wcwo2gprUHhmFP5L
CiINtEGPEkfMwv/jgNErTrrXe3sxTlpm1pZ8GCPo/EogLeUpMn2q9Ag02i8HU0wgCFIBtoMRyl6f
NwNGN/E/rD6tfSQeuhg/6ykdmFoZO9E1+PJ5+idFUY4Rb2mW/Ob8F+frBJWqKuOQul1/3JHZ5hgn
7Q26Nw/NEjCqRIa7NE7+sz6NUI2PnSoNzjZ3QBIgNCwomdwRK3B+9yksOh3Ge7eAd8lh87KPuxSm
yvZ/ptzQeCxrNh9yP4C11+UoWQ/5be+K22m588drsnLCFTIhP4N/U2AhkoYTql/ofBb3nj1sdKfi
BZJ8JU92zB1jx6LFZPTOKVYleOb4sO39JnzWnBomdbiqzOav6M8Y1WXkeJEVnRDn+/c6WH2CcxKT
/lPjco0Nm8DnvDGqev4M0XQjrxPZ1oJaA5v/hvqArSgGu+t0te0396hT2optBwn7329M+Eilii4r
kBsSNH9WsAzBm4kr+KJZ00fsOo6rZiGStGaC+GuzQ3eCkdN4QWa+4tMo8GvaWbDDlRQuoWlUouOk
uKy9tgMuIgGQI38mFjfQ7U4EXL6mTtxlBK+XROYAYvjbsrZnWqzZL3UWSxz78R1quqpV78WmkQlY
0OEhu6U3NhsH5p0iJPZCUUyG2yL3+6ZwgWZsLp+613/JnSvwSZ1Io7DfNm4vI0v6tsQkt13S2xeW
qYCeOcMj+E43/2jC2vWq2JXSpSdjeGSVlOX8NTqmknnP+MjZjpdVINqLy+IDkArc7eeTqBfZfhlJ
Pn+het2Kq2yBELD+1rXadws+oaCHX5+DofMRo4eF5CmvknxAYGxiLRxgPEX02oqcIN86BhMGp+gs
msdfm77WITKnsrczJKcLfskz22Xkiwp+XmQTlWNQ8euKIDhNUPtOWHsDSzCpkCDn99wjzRez1Y6X
k0bzZEU2J+ShB91XM+bXhxGey0zTMY6OnFQtH8ViQE9Bz8hi5p4ZGARhGW9zvMaGE6IvZFkwbwtD
H6aGP3a4CgKRf7Goxxd3CuhGsD/lEvEQ+Cy/jAwCCDUIEfFJ22XM6goKts4bOMZBKmunnfJtF98u
Yh9vBu52sJO6fgEP5RI8Xg6dnUXEmycuVMEiRi8fYbPyGesx3yJoTF8MVabyVyzuZah7ipg1q/Gd
7aKruqttw/Frq8rbOl71uxaOzK5ouEdoRFmjmKhRymGpONx8Hi0dLcm3bwFefnk7aWhUOTOlcmIp
Brbp6Fq5VxFg6ROqVw0Vj3ufwmIu9rL6uEFr7LwAJj3zaktt4Pc1vIemaR82qzdjSR/I507ZZfq9
XJZSSrewdcNqXkDR8UpWNxz9Ajh3SlZqBFz5z1PsDvBRey87y/2vbaIa849d5uBIUulX6oHrT/S4
3f3eqPvMlW3y3UmH49h+YBXpiTKQleZtpfQvPGYb++jSna1AKzUpwmEqzthStRY0w43tAtIPm6+N
uo3BtpHGF27QPNLLC85UJB9txGBEWRzAKKnf9PEfBquChjqbkFqTfuLu4OlhBnOoE09vPhcn2vab
WIR0UiJIgojotv2iF/KShgERJZ290vJ62wBtdxvAD0ksCJDcBq9JHKBSstC57HL1wEjKClhwechc
D06AlEVFbMIVTS+BzOVKiX88qfw71ORkUWLMnsaL1nvgTkiUfCWVnmsWfXhIeNuR2B1D3CoB4WBi
AG0pvqwXedU64Vrs2uSyyVUXN6q0k6JEJVbXUm0NX3478v0m+hlwQVHr+lwIigZngWCZ1gIM25Nk
RJPMRq9KcTAuweUvn7Yy1s2Q3JRoZyquWAcLD7No3AFb6H5dinIamfTiWsmkpR2EkYmUPmqLjoro
9iVgGR00X2KZyIlRNfWVqZb2x60pGrePXdEZJyf74uQPlCIPO2iSa8fCCv2i3Mkl+A7F5HSQufT+
GdvU0XhUcGxIQWTfSk77lxDm4KJRQaZQPT+UfJpvQ50nF8pj8VRQLfaZaAonkKVjt/5UW1P32tjb
MTl2nbSz+fsVZn+tB12n+3X9cV/IRwVEtgsC5ShdAvhxxkKN36n6pylmb2loZfgXTc+xxsujFaH1
6WghRUL7mCn5eROApfzJm95GWvvSMheFKwnKUSbttRSZLONlOK/xBvFmisIsolsZmN197JbyDh76
tFCGGAiaPOuKLFTz/wg6eULIDowZftJnlpoN7tBOCWutqaioIqqVBhSU+QnNw2kZNV+AhHYdqGt6
B8SgvQoTDcIA9wQfdGKHsbj+tH62ofB+zvEkVRo4pUI9PTUw6wSth1BHLJCib9RCSOXhJyKrNd2h
Nt+ifNssA0Kbaq5GHO3QP8DqX/QT+SPo7gLvPBw7zS/StnUM6JmSgOGIfHCLs1pJbH9JVjNHWIgg
mAp5GzuoqiGUysTeyei74fLUtWhw+nTS8Zst2S7atHbCa8ShvpcUDLP+LgGr+5H1UakOq4uENuj3
EsEPcYkumQ3TQJP+sIH9WoytolmilS2rvUdfYQ3USwITd551G8gS6KXs6PC2oO0LUdG2XXUTVovR
GcVGGBU7UcD0qqhJ/ZaKLqfP0LuCk8JtFjRhfeh/kyHCDPGJBI6UtWkYPeJ7A3NBJzcSgtfciOTJ
UQprgjxrB/8X/CbRtFU5fQOfk4k08azbVb2UHDlJ5v2A7p1Nc1reCTxy6WElI54hwWCjR1ZPRp+U
LcdgT+IZ9EEUJ1QTc6n1QfBf8iVDHtotH8qdDDyTRcEUZziOQf07auZndXehVDsvxEdj+CaLDpv/
+uXdM62xWUGmW30olOiOkchN7KdP8xC34/XdWRFc6Vmn70YmMkczDWzYvt4rwPCusZG28cdt4VGT
/xHWeWNE1YjLe88InQeQha6EOJa/J9TaL3kG4jBMASFRH3lIbZrAz5d/+LOBfYJfs6glDqGn4p/H
d0PooFtR0jTpe1cwlze4OQ9IfYb4hND+gjPxitWXM83XteHSfvKnr1QXPi5u8oPl1PKYdmFjokai
54n85jgewe8mgbhHKidddmQ/deAtd+fn6fmQNwAhC7YZHaTyQ32kze7vznqJTihSSvFnwc6K1G2+
FR99sDdyTn30S4mQR9t9YYQaJfGlf7yiycaAxc4JqH/F6yTUqf1KBkTx2n3h0n9jOZRIY1F8+mwz
Wa3ObnfvYFac5CJsCqU7yK6PW69wUqKJq5S88DtP7t6/+BI2uocbgM5q4MS0oC/wvNGSbMxgfVt5
aoURbaB9+oqs0yIImePyCi0Mrzk4+PQz99/LRURbpvy5dnpCEhneuka2nq8O76bOupZ6Kid3lUPs
Fwa1yXGyxgGdy74DZ4+Bm7q96+2fzrAwX5KlvG8vB+tcViDaRS2Ka6wYCedsqbd4E3zADzH9drJf
FDh5jk7gECxHaPG3TWZFDCp0ASNPqS2ay8p1hBJyY7JuhIdr1wfehj3n0/pP9i/dTT+MXPpADWw7
QKdjhHgKW/Hszc/EA0BxX0a7gqdI0zbrpe/Jg0sh05wRghFViR56ESfAZXdinaSFIwz7NZnX0dRN
JBOReK9lq4+r92VhdjoTm/S42oAbHE8Kc31krRsvjnq6WFzK+EvIviXDWe3jxbAW6iH50AFrJQDD
giagy4FJQJBgCKsf8rlhVaEAe8MCOMWbC7bfFvpvtcIsISKzjHhpUrgg7I/zc1Q6P3tvvUG6/dFs
WcKRo5nO+jcpulBEp+/2/u/U/kJGm5BwUCoMG2mODlo4ttNnX9AFZVB0uNSbiq0KJ3RX4bAm8Tb/
4yE9I0jLYWqGrByUR3N97Js6+pUEpn8SXv34J+DB+10XPpsaNGuqTegsUkoH8ZvBJcMyGS60Tosy
IyCkxZWCKcLWPPR+cJtA/JeJTymcO7niPIFYOROibFUfd5/qXqQiXTyp8l6XbjgA/gcEc8m9D0zO
XjcYI4ePg0AJePksp1Hy/rK8bifmhDeahNHA7HuG85AecqtXzXufXzr5PXoSuIS7rOsqyKJ4mrnN
PUvxqiy4/4WyFbRbPu9JGheFPhz2zLXVpJXA28NmgVbKO7JLfhimILE0lWyFp8Klh7t/5axeWoUv
nfbdLjzksTiOYAfMMBv541PifKlMfnP1XNt5T+dG/5aPsRAs7ZI8JtO1njH5S6hWzwd8mNeEZy/A
uWk7Ffim88vvf3llKytm8L7gW3sUFLXBJBAvqRwFekATschmKyresUj+QyQNEfZ3Ure1BKBLSH5n
/f9keBLfSzPjlxYSwaTYjALAktPM6gWmYG73wV9gQNaE2Yh7tAf0CYKct3oSKggtmZhpSdndC8ut
UjhJe4Aq/7IRKk9CAO/XpU3WIOifUNCMviZqycP3SW1or/vAuGDatC9L/0wTYqjcs1QSQLQtCniB
JbDhY1GLuOvD5c0h9xUV696AQNhARUOeCGVYfm4EjNARGqY/bfVD4Vyv7ydYmSYFYI3tqRBQFsaH
Y9PfTeGIkiIPT8teJ06H8ccfaWJskgeuhNxZ4LaBiPN6nGVIlrqjnFQN3geMSbD4ZFCNmJafuCHd
W0r4v2pvwBIzVC4R3CuGGWNHp02/SKRqhMZLDdPO4rddbbcec07mg5D0Bla/gtmaEpxRD0BolDA9
pt/OjQpuJA3qaVQjfSMRdnrUxHFMD8sfF7cWuY37fMKvmjqT1MYfYkylIjDHyp/tn129go9zNtzD
PVkldVuuWwaGFN+uPXWSUd7dQcjZBLEMjjreomxOYlqxEOWTuRkq9WIi0ffpni7eXp0GJNDHbjpZ
Yjtj/VXqeMgjyIm6jbCrKNB/vaxeP+zN6AUr1VHI8eWS2vHJJ+Jne/sCOOjMiuut2Dq9tW54DrjE
95VfoaK9aFWkj8RbwemueFuBeJWp1fo93aCxb4KBrJ8uXi7Jt57vFsE/lVDN6Oj8dGWLFZNI3UuV
wnmCHJqMebFadE4zjXYwmuHUtUyjBFOb3GNFGlr9+IfpguKhD5Pyp1H0+ip3JMGMz+YjieG+fw5P
a5SGGGZ4qdDsawdckYeMbei3nKaCU+h5gKu+DCEqqXan1OuVMmLrubcD7hfVmw8/BD5KOk/+u0/Q
9Z091lxBfiQ4cGTkDDGEZ89Viqkw00OjRIY3mGZGzyKp+Kqg02WFIZE8DLkHfM8C0TAfqebVuU5J
SyUueUEQyqKC/I4Fks4v14IkbqD0tEO6fMTFXiXhfDLiAd6NXUkLUXJ+/jW+ICrQIL1+bHJSuscR
hcvuBEAf+3rV5T880YuQKjUVBKQi3xCOu9kLu8uhqABURpn+8yBEmF9qjOfVDL+CuUc4irijm7iv
gTcQOsltPcekhD+bUuTJQNq1t3Co716b3P8cY94j8tVw4t1DaitA3GPvlaml3ITltvxlb1COLf5Q
UhSzvbNlxj0P8b1rB6xW2dE6kEAVMRPfLy9aIQRYgbQLp7HOzJzJXhvdbVifiyNzx5mN4jv5lWKs
9fG9JygbeNEhvQaHwD+HdE/JXPrJFEEhNfqeTJ7L+WBYUH8yUe5QJi/MY4nhzv6DmDjZmOolD8fj
5Qa2sXLji0wHJm5YB5KJjb2W8hH19ZiU0N/zAO3RE6v1US57Qp7fBcbhK5J2xbjClhLMaWQoN1Uq
Fb/gQk2NBqbJ6FDq9gaDJcorcJEJws0USm58NuLjCmyZYv6yjXch/kcsFAovTjPP/b2zJFlSgI7P
yvoxMAiujmDQg6qIXLQmg0ukAU7XeXxgbhd+bDKndwusRDPOxD8EgQDuRMRT9hrAi2Hptc9DTFi3
RW6x0+CnybEd/RFJMEteUwdKXDuVXcYizFiTocftBtPfJ2uwK+u2ZPt5jyljhEgKO9BQtmpJm6S8
6c7AOglKn/It11mNMXvkgkVvKLE3eZqk8VwKnbACuwDSwXhjJC6ieBFSUT1Zp7/dTHKKztLcwSnl
PJeYRFnC4hCnc/3kIE3gxUN/clwsNwcu8ulpmZnVLzNwoeBlXH590fqPHo3yRxt7QdOFND+mIMhV
6fRgbhbtecBn0QOGqKZorPqUCz8nlOIynRJQiI1nZFP33qG17r7lwvFQzHUtPKjCKI4YWOTHcPhz
DsI3L7lxCXRqAwm7YF9lSgtddImVf5YvNShH8zCHHBcjpqiRJ5wUKiQTSJTvebOY+UuNN6ra+Y7v
wutee5J11+qsm7SuBFc/4wABPMbg5wObpXg+IAeDE8c9kFua0EAtKZRQvgLwzpcwypyi2AbPi/NX
CZE1IipkRdO25TuWC80PA7RJU/jKa92lOACA16ljmLaSeO+Bm96bIrvVtTOTkEmhMK9n4Fw2AElv
xuQL6IdWi+tr52/wC4+Y0Lp+zhR2XyCZpoUXK6RfSSEshLaM8M04WKxDJ7kRgipB3GPBYG4pDBu5
CYA8wY6HB8Mkh9duCn2rj1GXE/eGyHild47EB0OFdd3C92T9T49IZju9Ky8mTbLTAjRZukWXZyqM
RvZhwi21kVrPtrMjG6y6VYQ8Ono6hH0s/UldX4pxEWC1QRMGNqVnU8k2gXc5uckCJs8tUXJWjvdB
3Yc7t3YGDHjMSJiqO6yrN/oOfsFUqQNCsKPJZ2qzt3yJ0uYgWTEIcPK+yQqjL7FHNScrio8aepW5
NbPYnDvJKQvFvseEomjOwshF05bG+fGLiehlx5pu6ekDh6zwP33t0lAhTRxILf4a9F4KTHsuohJL
o1AVyTV5FiMNfQmfKtPKftyPBYixskyRknEYnPXoYv7MjZUy8YyNwQUW9JyYcS1dMJgQ2DC8rlec
ipuiCLv2uVWPo0ezm8U7+i2/WmuHSBLxocXHcNqPeGHp1PCf+sXtYxvwtUScQV20195ujJR7FAAV
PjKbEfSYTRocGxgyk4R+8uUpXHVx5Kq04K7oVV7oz+2iiFCertrCBoCvDiE4DfOtAbx/AlOn06mk
7hlWmOvu+UipNPfFJBdn28FeYCqL6FXkahwN89Y/TdO954i9KZm0IIhAkLLpx/jb3tsgBw87nfkL
1KtOvxrAYrpDybbUpccK39hY6UQ/QpUBD7kgxbxPA61a7NZNqXJaptsCst+lkadzxPDWAen0fuah
w24T8NLS6KNmgRuxr6k/NJd1UTgBDZr1y2CLZH5R+2OWTSf7+knGXKJGETT/4XBIzYSLahvRFrez
Bx7aqRGUHZE/Vhxiwj//CCWubjs6P3fVq5weoZy+SptEUo+/Tm2pfhioj3iLQA6ntYRtplQzAKXh
GU+jOhPLTuXt4uPy22IWEj2m4UVjlQDDDMLbpj6KnqZ8M09rRihSgxgWJS6QLIuKWIH7FOzb28pL
DJxShFkr/PsEYGqXksJhubOLRz5Ic6zOL/7l2NcHjWQNRahsQvXFP7JWpvlyFQhAqvLTHExaPUlP
lSNbGgNlrzzczGDbhZuWqmhSFPgm3DPWfgYNc0S/eQs9vre6+aSEqLVBtvKSUbSRcL2X65/vBTCu
mAnPYp4QvdamLnsLGgzrTwoOTRv9nqpworsPVwPQO9oQtVFMDaKdQ6xsPuViLo+ck17gwasaXExw
6f1WdKRzzwy4BX06+9mM8hiDEakgKBUUshq5BSKUqgQWW2pma3TD0JKK0YJlxb6LRx6zWZO0F8m6
KwApwZy/KEU43Ki8N5EgNk026Hf8Z5JSC2BhsezE/QcJmJRVnrv0+XZ2om76f5fC6xg9NIyc3SVy
N16Z8uxiB9P0Ct+2SX1I9kru1qv5HzJ09DGlAYwlAA9f5El+C+8PQLSyogWFgXHQX8r8HQ69ZVbo
0qhPgfvX2Z1bAoMPDaEjo8u741D4ZjytJCeUjxHtcPvySbY/RHjyr9ZyWF0U9bmA25rFrpc+1kjT
L1+0XESebENoQoPCecwcQfaStM97xtc4DWqwDMj70x2atkbc+8URqIZ5kruUXCaMX79tLZi+d6ba
rLMwDBfbcmByuGYJBRgsHOesOsdv7YhHCUWWxvOoXesTrs2Cl8yy3gOVeKKTMXG8mKWbx75WK1gm
4xbz5uxEwKbts4XnXSt7dbGYLKhC7ossSvUsHFNblRwKfIUFhohcevZVoax/moq5fWQ38qCEBTwz
AHp/wvVfqhP35ZlqD23bbQYoeECa8b9I91BqVJN2AIfejakPFcekaNsO7DpANPKOLznwtFuBxpN4
geoOXPjbNfKMkK5F1f+LH2EKz0IwW8VPK3ew3alqk5Gs6sJM3VuRvMnHTBXUCU0T7wOlUXM4lxMU
8cLeAgUOPokHCxhAr/L1/hlPJhmCeprrt+ADnpahXS/kFHsQIj+vdYcPm1lxlVQxX1NCSl8cYjEc
wBay63SKnKiEGE/hMoQFrc3Z+gLbaqnodoJQdMIJD6yxUepQvtJfAXLfUf6KAUxnRek2mZ9ULnq/
EK6llQFWShjRu//C70W3yW3feG7Pa9K8ZJzyTo7sSb28aVhPXewYm3vDKamj3ngTfZw9jroZ0EMJ
/oVNZaqLTuau3e/U5fzbe5cBVxOFwYT/QoWkJ814o3WURc9kvkriJUmjK0LVYK1MHfbfaOd7jUf/
ZZAD5eaCppOkqQpqakZX0JV+fN6iaL2TdJuLZAG6vU73qwRjjHp9ogKaTYugH1OwQ9YjoKR8TPQz
oTKJofqOBohBykmeVBhR9dWJ54flFUnUy931GCBirogMIgxW/Unzy3rr5nxZ9S3R2pKQt9pFD64z
3kyCLCZDpggbeXju6LOdgSsffz3IJ/4wN+b7Ex9Q231lUWqPciyzjZix5agPeXzmRVcKXJRgJPQM
IJE+sgQ/Se55hoRrPZdox24Od5nYh/34bgzlrpG6snKX3VUTysv1WrRw60NLhy26MwwShKWv+4pg
KpcJMn4b6VvyGHxpY1X1P6T48QRkzDLWO16AC/rcxBaJwQj3CYtYQQvWc3vdJr0nFJi4WPpDMIsp
74oSPEp+QCnmBST/SEyV7AIrH9LoaoSbSw27p2IlOjM4n3OC6SZV1zNrIJe3XIfwNyogClSLoEhj
GJTY/sGeeoua+cK4P/bxBLKXYGH5Uok3ZyxXbmgpJtFygCrA9lQzhi/Nh6Lj42X0Pw8tGAOzZ/z0
6CyT20byOqnAX4GytXKPrR12Dj8PPpvdoUE5/EWVYACyD0QRxd4Sd7jUgUJ9/m73MH4GojhfQt9v
44+PdTu/TNM0HLcwDndR68O1txX+yGzlDP6WtVTzsCLAFjmoDiK5jUfAXFoVNvyEzRSgQGfUR+pV
9lmNEN2yaoL+ZgOVrdDlewsUbkM7EvLNAMUjPRpAnU4C3oIcyjqwkR4Bv3eP/xDF54NR6XImslwM
DiuxRS9y3Oh3C85gLKxZhSoajjfbM7QLnonot0torb/g0G1BcvrAd5aH6fjCY1eTHCOzJv2h+l14
Qs/jPYpWiwK6VVcddYcjRFp3ulCrGX95wQSBGqBfg5/t5ml9HvOBrrKDFBVC4bCIrXyOxedNrFG+
VUt/6nrB2wb2VoVfVkNCBNhbrT2sdQgJ3X7jmJjVM4+RBESUn/jOk5qygCaPx/ZxdcHH3khqesSR
9D9cnoO9Mwmr/ykNx6Hf76HjY37Ngis9cw2AoWSvnrPntkWtto86NQxY1jg8BfWocj4j8JgyKhHv
FBeMbp9kLADE/ZBr27gFC8ARVQ1ltiFXtPEzdJuDn4HENnUTtzXp8OswntBCBB5mST2g/3YRh/bJ
qGVM89b18fHV3h4z5BHZ29ltS36v/vWRRmTHaOS9TfEV0NbsL+L28aJn10mgegtzhHjqkWL+GaQG
XNjQ5fID/uHQVwmMVvNcOVjVSlz9ZIOgv3du+uA2yWkrXqHr3zRhFuXRGrk/MaeIhNGaca52mgvD
61Rwh3/n4xz6vUwQXp05vsakK3rt/Eih7028xXnWib8I5COvPT9Ou8+YTBgok8ezmkRrnj2vcR22
xB+yE8YYibWV+BlM3bKqASEd65usssrFcwQgcVzO8J5Oz2pRy/vb3TgjytaYtqPhB3d3SnP3/8x+
ed5DejCbgDIyba8WwcrBtguHb+3pqVxyvTsIQ+JWkzFQrG6SCjRchO6cSeS1g2qomyfA+jpOmE9G
u6GcxDRkyjGTLskRVJFeKF+JusOfGgTd9addhboay2reNj+226JWeM+Fm3/TcxrnZ7b6q7iQSX4f
ClLx5luYD/l6AU5bHMpgLCu2ILkGYoFljdb8sEFxPSqS6S0q6kci8NO9AKoofehX6gsVdBuuxMYv
JZk4kATFk/l5iM08PKvnyOqqxEDuAqV2GBfj5n709bShWYMvsDO0lrBlpPm57o0zzwK7PyCS7xxg
jy4vkCnYufn7GKTJ3vj8EdQD/4N4VtU+laTQs+DqWMmyNenCyb9OGyWnWLdUgoMFH+GgOTkVccC9
KxJ6XEHE3C+7pBg6Phjj38QBqtC5pMOyALw49DdfpC+qD1Y7tO4Jw48Ti1TWFqT/y6QtGDaNKj7Z
XNJZtUiE4kidJeGn0ewqH6WCex8pRiBQ3x+5/s4a+DX6NUU/d8ea4P3bJJ3+apgKH+zsmW6DK2HD
9MNtLsTsU/nx24pgxe+0QvaoeS7KVjF6S7izvP9WzIWOBrnEkC4Fx6PoVhTy2bVGTW9Rjmx4e3vg
tgnGq100aRzbctZ88tZYVx7IrMPkHVN74a4yXt07GGW/cJhT8xkiabSOT9GxaZlKphnpPDdM1ghC
XqOv5Mo1oazyNQgNJNBEKuIck0MdZEb0EBESQ2mstwFBdYYhCSDajPnGG+I/wO0nuh7iuvEvWPjV
WuNKBiH8zIokg5yaBje8UhDQtcckTQ9K7ls1vnCjyWsJ5wzSG/+TBoSVFsx0ZtiOEXdHr4QcNnko
amF+P5LHv15lHgkoTmXK5Yraq+7jgqN+/djdd9RgQvgR7b14kSh7rRSJagZLvOlIckYEq29VI3ME
AecATpn10ZGkfoz1m83uc7xQZMgbPFk+wHkt3ecFOZQbyBhvjKuArXr4nWKXcY5jHWjyDZsrrrD5
NoXhZTGCrCi63gMgfiGRV6qqGNBWMvauk8qU7rxjlqRz+KTtj+jpjj1oFCWuoQfnlKMSNV3Gj9RC
nBeX4wz4dtqwMzxQ/8tdLaq8vVUZtgqp4uihq7g2sPFfo5aiAN2JgcuLJiTHdXiiUyazdPscEmKj
KysNQ21qd2C/CiS4vNsEX0bAUG/mABPkp6X1aY4hWQ1c51Zn5W+Gb+c829lbGOqZYkqrtHkS1YIa
DaUtE56qXIIAix5PvFYi0fcN9+okIREl9HNwt2SiMHVabYHrOr2ekr5Q04j9Z/ugFeUtpiDqbviP
4MLe8RH56mArw/BDiOd91cZ0/obMpffI9EvTmK/DmgDq5HY3Adl7RFPnKf/tjyMrLgB6QJlEAKvz
V1OlAzRu9YoBlqmhERiMQobyHzyenB08GWX36hSVWydn6NcObNeRvu1TrFBa78A1edPpPDDvKGCw
BW06RzQvOsSQeNZFFh/3C6PA/fKRIAUrvVr6+STcicC/Ld/aWRICgfTb/pspAZpG89S8HrW7/ir2
CGtEIeUmbJ8/Q7lZvOfSHFBA5xb4XB/skG2jnI0tl4+Yhagunn05mtWy717P4m8onRCSZoEOxtDb
7FDCsgk62N2z4EKXw6qDXfIggcsQmSoDFpbKOlRVsuLt7yEEoEkdNvuDS4hXzRODozKwq8b5bsKF
JIkkkMRWJc+U6cnlW7B9eYs8bb2sN7OZJguwOnFW8V0Nb5tnAcXZT8K3fQMAAIVB48moa+qSKmyO
VOAweArTvYDIcV3vQC7J2STS6sTv169a3kC3TH1iTkvSrVQgrGNn1ltniMYul362WPSm1v4WKxpC
st9HxoZwJqxZC8/3zepFLz/FtoTQrFcm0YDFXwtws/FLM6OJANemkJYg6h+7RqHDdIFfNmZk4EqN
qTmN0Zntc6uRLtouBeTlp+u0Tt+QDlmmNIP/yX2Qsj77aO2zAZxvAkG90K6T+Hc3Xpq/ET5160tb
Gig72P2x8SqAmRedV94cQtWWJ8GaI+x9WwuuyvJVqPCT4qa7IPdRo9jcJMDSfcq7XVmYRZLf0AIN
wfmXCOpT6Ctt2EnRSP7e3eF+SqMgFmkPIOhAZsBENTqEyW6fSOxqMsDioB+uQyZUUdWLmsPNVY9+
/muQmTaUAD6d7UeZuD9U7ap7c3iXAr95e8e9mBnz+/2q6WsKe40unb6VmF4rZN96eflbrXxzfOvM
cXxFoLyhofSohgHSPriIyHuNd53RDrOdu2Wpm3j4LXrnJE0dJT7pFkmSmy/Uyhzfz7nxDVbaf0DF
SDof1Z50zcSfV7XwcUZtH3Qsczdql6aX5GLG2QRXX0AYSBVvG4u+wj7C73mMqakSlurxxYMHlK8l
jtH8m/JNG2Z2UQwqFDMld8VKapjZUjE5IkYuiYU0xDvX/VzaE0gAnlQLz6YWDaE35JJo9rqvgdQK
6uN5AdxJZSUzDM8eYP+tKNYt71Ujej6DNCjxp+x6cxfpSH1vKBLkO9F7jQ1C1t0ULSIkacOObs5x
gONZvyX7sm8Lq6pKPnVMoEthh4XtcA/ozIisjNCAze6cMSpWLP1mdZ+YvbJE4qtOipx1PoNVJ7lC
7tEqSSYtcT0wF9/F150aOvPGsoSA+lTXfKsAR6aBUYgzGLAh2vBgslvHHAgQ1fQJwaRvJCJKYu4G
mniKu+VelRKcTSMOfRzgwrfefaHJMOz/reSKwnqwqNiajLrACuIsCOeuQz4SqpJpKYqC3SpwnjD1
ZgHvlQKow9UJUK8QTR84wwRnBY+lXBMgg8qlPyHuOGGuocmoScJVM5B88yAqgsvGSmMjZk/ptkNV
pZG9Uk9+W/wzbB6LUz9gd99aGsXbacv/U07X9qhNtbfcOkQYz+ta82QCoN77eyNR+PpUREAyWG2T
LrtdrgduZO0vEtraviRD5TMSYuChwAqMnXNXy8QPSMY7X+7KSuEH4eWIRRTP+QjoQu2544ZQRouR
hA2wSmTA+e+b2MrmanyUet8KlTSqXdS6KoIY8mpFVuViKIdZtJgxNfJ5CO7LivOcrFzIuoPM8EIW
tSo03f95S0kH8b7OKGOlzRJX2eb6W3ZWUqnm+zLqrRqnGaQdt7vtDcVorZ4EZCkUdDxU8a+xxmcJ
7Y/ErqnrkrbVM8ZYOaVIEEKGVq7KYkGrG0sKKtDGZK65jrBEa5begBMhcW14ICFmMFEwhVybASnO
9zP0sugV8M8fLbNf7Rc+XMqJ0ZpHIi2B4PKCL0uy+Ts/+CkTyLLZeW4QEx4y2gKJ03DrKEC3jH3I
IIxtcBI302QhKvYiEFmyleXBW8nqghooeY8SkUy2Z4PM62vIrl1qTZct6b3bb1RR4Qjw5D03eWaN
+51mAE+E9UO9KbXTceLDLGbk78E1pM8jHfzGc7jBkfS+MDXrJpkiUB2E2n4VPC8/yLsJOSYDggKW
eIgHL6tw9kgdKopOTIRiQf42OrYPfdSosFpL8Dn1aR5d+jZU5ySh+x/MRZSCF9FulWaHQK4x644P
CanR/hCmSlhF2ZsIielESqfJS0Odcsm6hl0BOek1LUhUCRE++FNHm5QbctYuMiuhX3g9negyHCGG
Buz9z1O3wuaPjs8ETis9gHxKtXxDRuBHnFT02ZdjRE3uQt6QeDSq2CBjg7ETk4IggKY358VYuKSW
eFklw4R6yLNJon3y94R91LP75PRBxIAXOnfzTpoOKBO/8B+qbaPhys0oVyGfFDUvLZryZjF/ZhM+
adlAh04MI1gLziSot7VYNevOIG5LtH02sLM1qP3AkvpLlrM0yM5UceVvomWTVR7lX84YCpweo9Nc
paZBlFM2xHi7vnC/0dr5t0UoTKDKcOwlgOOc1uJLSO0i4hDJnxBJ7X5raBRtLnQUt7f3KGiZegX4
vLn4b7K0NZUAk5NFsueF/hmkEejhf0rmYmIZdQ2RditycKqzDL8ZMQXpYoKXwu/8LwuqrWaVRmzS
PUYFG46l5uBDe9au73JVeVmV0RuHECr8aIXTqYsuPDTNjbOsybFKf1MrNd5MEjjAWP6VErSy1OWA
DZfnk1ND22lVyL8uMvM8ZNX9UFbhXy00OS1WTCQsETlpeQYxoRDwmd9OBiNBEEVHSZ7NnUPN9Hjb
1NF4odmnQE0sExJxVvf+7dvA5uK+JPT1f2FKFju/rMPQhroUFH95tZ0srKrrdWgI28FrLQcx+7fg
eIb3xHikDcOLHVNBJURKG1Ux3wa5P8umgvmB19hiNpFbTO2/Mng3TwqD0d2pJ4SJuS5rFyXYS2zZ
U+4HOvRSmChGBqsmSDKQFr0w78PCFF/OvsXA/g8sXanBRRHyTT7RsieHfDQYRdFZShSkm3g++Jp5
O8I3L3KgwxxGo5ItyXBgP30BSksluWXPiJwrZfHSeMoPjsG2G0IFgxVYirwzWosRPJsi5FHu8tWw
NhutYJJ2I9jKspzYMdUSS48LZEh8GtcXC0TarS9O65VjsnzRpw3zS8f7833hT1WhRlYXC8CIcy6D
PagVtojSQBpcnaOINqyM5qxtFKDBo5LM03AeQQNvFhTRFIY4g7jRgqTtdFW9cLKsHkNjYk2ZEPOR
neLJPrqjzlRhazOMSLngueaR1G6HToA0/EV6guW7tnwiZtXE0MWnUobiQur2Rw43zX3Ygi+I97dd
8855G7ApLlOep9bLc/V+ji421kJYywTzYphlr/NmoxlNoT6boyw9s3xWcVKnr0kN7glGSYGX4y9a
ImV4oNyRNSGlvIIsO6Vks0VUdUh8gL0JTDNOH8pOZLDEuLOkhwD/j3/nh/q1gvWVdXQZMVqJ36HS
GZ1H6NUbfqQ6E5PhsVuFFH7VJGs+1dfrWZmUcPF7nH0HE6+3uGlITZ8aKqTVxPMtpm4KKzjKImnf
Zl0kk+Q71/bP0BzRGcMw72u2WQFWhYF3dZsH+JEXIZvuLacgYMO0ljme7LChLRw/kikpcACyjKl2
9Qm0MRhYvkn5xo4o0yGMldfVs3Y5gHoOU4nz4KVzwBfMUwmzWpT9mOLGJ5AzgVNUOtQEULAB/h6c
p5nA9KvKeaVBX3PnkUFkC7ALpZ+ryKvBVjSw3J8ePmZtfbKF6BpY6X0b0EZc14fvEHRsAzmK6Yqn
rHD8zR1PoWl9y2hJ21BOpoD2jmbpzGvVsuuBmChORvatCt36FLnbIwkUknwXtZ+87ITFlMNXo7gG
4H+F6yDZWSi2PgKzJCEdW1PHZXrQs78olU+XjvboCSkFg/az3Y+3ht1Ai/IiptBkCKK7CVUBLlAd
8MdiTRlVKN2IVaIP7WiJcRdjHBfMLDPvlpbufOZau2Cc/PVVhH3FGIP3gISLzUz7b0fv18+blbm3
76JL1uRtByX+qHTcpJS2x/mf3iiMTzNBa55c1NxGD9+dIrFDBdBnvMTZnmqZZS03H+9gV1qwJucw
TQOckEK3XyrWe/1I3+t8LSb8Q5pQwlNol+Fx6bLjFU4dc5JU3YxAAVUbsDHUFoO6i3WDxaJ9dWW1
2ykI6FEfjM/XpyC3D5BwbO3AffTbRx/Fu63DnHXjDEMhli68HfTKoXunoyibyyoFgpqxh1bwNKjA
UltpD/g73jXoG5WBVXANJs4XvDFS0jZJ+HYNUMsDQ32osUyxen9uzWyXKq9HYxMHjjOTu/SLbhCt
o5wVABleok/C/m8sN8pqj0Z7Mh5hGqfWryHV2AFufhtxF45AtEyJ40RUZtGpwUjUqxX7Xs1fHsRg
n61ExGESvOolqRw7dEOew6c3nn35Itn84SWB+jh2BmWDLFJOGErH8PfZa42cPfUN4R2bWrdY7OZP
ejJOPWQwRSSVH8KyboE7y79XyE2cLNCfOyCB5qxkIu6K5DycY7efS0ZUVyLn5F+P1b/72xUX1PpI
2d78lsRdlAfqN0THbmvuse3n4Pj5Y/53fj/HUwkYT0iZaw5pR4HbmPYa57Xs/s59VUzyTUMpWHSP
EFK7l8tt1hXmfZMccobXLPDT6AV+IiKsexqg09CP46rpt8Ssgsq1PmWqQqquefngjkze7/287ZRC
HNL5Hg0pVO6yvgugDhwUWogXPvCed8JXP0zyXexNqb6oijE6RJBZ9Sk0jdXgFmq/qlrU5p6lQRrs
XpTa1EdVR6t9uFz7e+nUd+NeFmRaUit77NFZgc0X0+KKPAwP9E04kovdBb0rvgbzXeLMvro+I+l3
gEWbbVgABhrDmSpjDHpPLS/DjNnG4ZxDAaINhscZPXMu5rxaspGWoImYxf0qL//Q7WyuvLmcXSHR
R9sAMkqYcZn0SteMT63+xp5LmsbhB15dam594dXCIzIhWnQ2jagQwZ0+m3o9g3jP/ZDrPy+pSdad
DvrNoFi5irJNzdVzg8Tk0dvj6RoR+T2dnAIJNqQsRQGBvpMaPo4oTwcs1FS8vHrb8MSpZRI1N3xY
ega9AG6rVa2hSIAMQLQWXg3HGLKGRiPPxi25U1j4CtHYefr/kRy6fgXRvfrXPGc51aU5N3oANSgp
bGABuhoHg2H++dgWoWQp4yGNwHiIxEJ+zX7K84KNsy8pXzJPD63FMAy85hyoiShtdMyxO0Hdbnkw
jIP3KZLQCX1j2utxnD6JbUei+4U5WAoA0jAydYZzl0Whgrg61zzrnsFK4l2yfH781tivLQ9N4Ht4
bNU6KAvTCSSIiVAT4bTqCIXic1+dPNx+Eyrx8qplXmB916f8uKmAzQlm11zf5AXneVAtTX2iNXE9
66SJa5OTqHpxJb8o5i4w0E56QcKS3xQFe4dOjOrIm/m/dqEHIewoZdgT66GGJ3Ueg0FjlRjdbs7L
uT1jvKYE1cVYadpgYGNgk1HS+pHxgPV8HNyeSi0iRBD6KIl1MyVNotjLps1Ylji3zi9MwCCMpShc
w5D7Otx162teZ/Gxpv+nxKd23FJdNZrILd1TxO/lwc3JHWTNavjumm0++obiEpkmOkqfKjGDL+0b
xc9EAUUcir96wUx7vgwzrkL8VtcOUDgIrj3Olhh8UVYgns6J0/+PJoTZP739D34y79o5lvnwDIgO
8j4lng9j2AoM3eyWl6pb9uYaRlcJLM/Jka4cAG7GjJK15sfeK4jTJWREBeeq/0Q+Q3//+UtQnQTV
HED2xyQIwRFFDJvLl5czYFHGa6tmDDT1SNCd+qblSpgTWITC2YhYj8M8Xi/LvDTqxQTC2105dC4T
4+xq1ovD5gexHVfCpVI3IhCYaKPsUi5SBWPEvATqipaa6pezQLns2Qq8Q5xuB4SXo+wcg3V4FFq/
C0EfSo1OafMsZWN42kgdtcJlajBXY17EJU9Dp4EJEC5wKVeAr6FSwzgs4e7abHKJpZdiRI9BW5/7
HSTy3jI+UZUDR94he0iqyx4QNElhyte0QLfNSjggYg8ib1RkjHxBO9p8Ruh3R5mp5FwE/d7rGPKe
Zg9VQFP4rkMn3HMDB5RNnbqB4MpnClLItxhYkBTf9GyMwbD2yU5JJY+yPCM3WoNt1UGyZDv2AnjW
FBvlccQ6eR5eO8bQJDLGiiTBPLGjQfr0kddHxixs/Y0Atx+KEATshgJsm7wDY4VTghUQCuYDZ4qZ
Mt1boHh3/eiC81WnjB4mXmDaSou3RvPlddBE1cAhqXaBTNCoP3TrW0G2Mj3iHPDsJA5UTqgcOzDm
6NFx0dViaVCGXHydz7t+BNf81qiio4UnXSBdDL8zzPmkB83pcYPcNMVk9beVTo5dnu4UGJnNiJ+1
goNeRIuQr/wGwDO1Wax8776LYgklUhE2vkQWRZt10j5/zci5Gyc74xImtY3U1rpgbfK6eFm+oIAG
mH23yZCqfOYIzjp+zxfZyXKZGziz/ZCQd866W7DbruvYxRObAEvSmcqrry7ojoHcn58+ON5hK+vO
UW9UJT8rufuzd0PZ1XSsd5kavjIvDcDEhNzGOY5atY9qEwEH4yF5mOS3HFzve4a18ESHjQ2hZsyJ
9EiNnM2y/M4nUPJaStph2mfJlbpoafT40pN4yoKMRG1l2O8IwqYaxE1uyVAIgZAJkwBiqzTdKh1k
2k6vAWCaz0cjQih2xFnR4t8VrOd7GHSW6kRtIqr0d831SMH6MoBb8AzSNuZkT0CRXdFHMDqpZV66
pVlcFnOYu8Ha86yHQWF559qJ0tCxM0V8rvoa7vVsi4n3l50qrczaFE9zP5oQtJe6X0+06agRNBRV
6+X9PTfhDeFBlvhjrrwBO9goPvy27EsPoEffUsugvPA1h2lgHI20FYRTFfyP4R6E3TcVGmPb93kA
gS4OYVRPJ+eUhlGy+lBcsN9okzD2iyeJFhCg9su9E2voxMuQrg2xB4H1tOpe5T9JWE7gRbeEvZT+
ccith2/E7cfJDLIfIMof8yf3ZYWWR8OSU+AkJXR+KD/0lwkDPQdvJ0YjHvyAlFvTQX0iPT5DrTQv
QyKYTZK828bAwHHPp8C2yeItyHNpCqDueufAFc81ZeNw0Ftg/b7cNPkTaAsQZ7M1Bp7ZgNGVX3w1
rPS0ZTveutS2NoHYK2h/guWimg7Bg6RCPclHmk0L8FQU67OlRXTq9iIxy4S8Mp7qYATLhjY6q/Vn
xYijjCa/DybJWwkUr6iTYlzBksuBf7joqDMjGwBeID8p4COY1wZILTvqY31Z4vyqaQPgBd9hnwKg
tGf6SmVXNFGGhciGCjzr6fAX141snOwrWK1r+P+p034BVtCIjzxpmotR1k4bKZM3qLNdWeWUSgjQ
Ly61m2sybxGPegIvMwYT2G/nl86TfddbVML+9QUYNw+tQZxT0bH97RitpCWjhKxoRaDFljmgwO9j
9rRpS01cvsXacBYdisdfcUrC/Mz/0xrA6auB3iQCZ5CeILWMlIQnmVAhxHx75UKpNnQUu2lwQweg
fon5fDyUTfbvRxHZcg0z+NSx8EfIN/vJSS4wzDiHNVCrhjN3NJ/J0mGz2EghbIsyWM1MeWN6NKHr
78WPniMZzDOczVDSgmpnI0nCen9R1ISYw01OSF1siSaJO2zn5xEyy99zoNt178prz1U13/iSS6nD
ixUt8ugivkZXabt8nzFOW4ZjWJi6low7BvegLGSFW+EHk9tniPRzCEo3b3Oi5m2giYqhECCgUXTm
gNvC39E9wsD9aE5YpSF9tKMIIYo/mY6T4YV3tQxkq2ZTdr7PBEeb8LbDnKmtqi1vvWupoXmyOwID
9slH+KMs0+2n+OFKDMYUSfAUExJCEz+rcl8HhvnNzRzOdkf/KbIPOF7C7eBW4hW6B5qkceEpQBHL
3rjz38rwQ66F6YWzpiBqgo15E3fF15pJvsogNojG3UCX+dSn3rzvt9BTtPsKvz5MqDOGurjJ62EY
Fz1g8acUprNnwAEM1vfXWGfyXivELbYqa811snXNApksGGwG2VjW4nIFvgD44tyuDIH/4JXRi3x1
mkYrfylJRtnA6o0QKqO3rgat5SYCT9B7g7yk88s2qVf6/QhLfUBgyFZFd5+UDbezRSCjI0x4MDZt
1WLyO25c2s1K8d6K10WiTYGO5dI7GB5q7jsBNdTY01pHSdCMb8J4PycYknuX+jVFhrhOkOyyLnPR
izS809IRowZM3B5pDCvF9/2J6SgsUkJZhwlHwCuqGb0AweIYM9//5eAjNs/znhXxOSLG89oGVczk
b7l+bLDmmDo0ychLuLIwLLky+p7yvkGiFa7gZKt+IL8WcC6daRKgqlCV3rxQxsWzDvvAXEcdqWOn
h6z3dwiluWFZvUvJGOibe5SJjo2sUFc+4stoeGF8q881sFzKcpQL1nBryh/BoUWaFkzWgmnNbHLh
gKmZYHPhPxPR2t8G1gvp8bg2FbpEfZ5UTAeQ2jUgagX1EQ7etZPvv3bF5YXxIAt5gYNI7o5KI1Pr
jhKYqTz0zaVmAPcnTFMRpMVJEqSfI49HjnBUZ1w58q+SDyNP8/1WQ+EczoTq46AjL6KJuv3i1VLB
FpmX7GW7NPZLrE+yrLJ8tRCMP9c8u6E1SmUOI1GhwqnktZt29dNUseSxv66KZctgkxuY1LQJAeCB
scA/Xr+XeapZ969oFqRphKQ6bBJb+wkxN65BCHWGGeRijhK3HvnQcnLpiWHAEJzSPvsmroSObjW8
4riBs9ldOCh7U3c7QmyrOr5zHq/pMWwUX4MyzlN4Rd/g+YzCoVqJNYW4ftuSe0DktZ6Klgrk3HIa
IsroQFWvVW9rUF1N57ikDzR2ElFUA+4/+p2fOM6HKp2XRRnf/PQqwcoXpqKVzjMTDxJjwWfcbhsT
h+PrgU7OS9JrBbHG0tQtJJ5owIYRu1NG4ERgJbx2phuA8up21mEg+FQnePahUOQo0ED5hV4JK0ZL
DwcSs2Pwd7yXZF4KCKp+im3SN+zdF6oSjA+G0lt90X6BIPM2lnwP1FPQBDKfRZpI1UgUF3e/PJZW
d2KJ98YCQPrdKQA8FRnSXPt6V9ho4G3/jWn9bYrUfGR5SanP3HKNylXvNVVN68E7ZkBvLqxiDFUQ
Q+VYFFnzoXsH8InIkZhw/MhNPoT18BRK1wST+FukZwqPwPhTcKHZEG0CjgzSGs7UailGTZ46PhsS
4f1eXmdFEDdxcB+RJ8k13LrML5GaADw4WjU+/S6EGQngIKCiS0Rndw18d6N6E/NQaC+GvaG8E2gH
CQqFHGAQH2tfzELtGCESY37jIfEGxy+O9zh/GvyyeHdU2X4cyPt+8zg+mfPQQ/Z2ZIgfcqzPoTEy
jc6WywlgFDQn9Li6efVl0gRLVVT1/4GXHbSAuSmgqkHvolvRU9qKcelbMbfXJjke+2jPPqNwGgNA
su8Nm+LiZ2vRqjuhL61we1kjxc5vo1FnDF43UFBU/jkulwDr2j02xh7r5hOkvNbcWvkvLjw6+TYu
4d9/88ymPHWBXObdNXdS9C3Ieeurjl4TPraNI4Vg6Bl5iEAHt0Es6HSbAoraW1iE8o8YwtGJP5Hs
uCIrNyCrYXlHGf99OesBvLN2+uGWsl/l9ZZddsRDDyQrTT6w+R2sqZi0b7r5oBBO5Gx2qM2EfUR5
/4XBiKomjFRD1GDyAMwTnkVk7OraCCclL3M+dmkBi+pz8ofPCMBr1FCgDO87jHp4OphtmOtGyRA9
49eE6C8zhDfyb6jhleViyHkOoh+knOe/4fC2SJMp1V0b7GSbQ2wOU+cI5MufiXCZzHUnixiRvraT
F6YE6KniGD0XD4UFG9IevolkH9IubdzRPdfy/38X11LJzK2DZIxZWf7ip8n79sq8lNb7YX05+Rwe
wDh/JxJzdCnZAINAorNm3JthmzKqlq1gXHnzI1xNRRa+KJiENP5vn/r6S+t4Yc/AFN7WAepBym1r
kHEHVuSjiXjcjHwCKFSzkAyasW2OUC/ydQuOcUbzd16WTKiCH0gEVsNZMq2mvo/7HlPpOr/a6Dmd
4XRA321cY9O27JJWd9VFmux75chCPKL2nP5FJr7m9ESuRxDJq3Oiq0koDkShr1xIHcsaAkCoZVUy
ux2g/PItZBvluXG0N8dumXLpmMV8rFO5HWnDqGk59Aw0IfTDVg8deXl1x4N9S2R9jetosU5FSPvG
H+mH5OLRPr5k29wo9Q6EMqnkxnLG8dQ7B1kXDgpCi7rERcczHDAqNx84qPMp61mO315Yb0N32XN7
Kfe2gJiEW0jRyQOTTYl4wzF6iIXg+omkJreKvnnsHNlCPi45X5tNInnrxD6V0hX3V0uruOmhSS/6
58zOSOYeLjaj95p5prI3mhCX8TgH/ySd9U73f5Ao0QxZl6XWUPLNG8RKxEg9CM0F6OW4eDQpeYey
LKzCYztSoJFsexzJEdUn+IKWbEHF2gUrrFPr7243PmUxGC/PhHj5aLABZKZwOikzTwPozf/BvZIT
kuvbxicryLk75jCEQkygjJrrccr83kWv3zJH0D+Su/cTwnjkTcPmEo6i+YDdcW/KYYfdUpHIdx7r
skWphfb44bpZF0h7tm3VOTrbLBo1Wm8+NgMgk7nQKZ10ryOrIKxbosqiuIA0+Q49dwd6VHpGAMet
iCyuRrgRv2zyHsi0WqtQopGu4TDTjp0rE0H1bkPe5O6qHJ3PcySGBv69Lb0H1hLsGg6obNsaVxXZ
ORBO+A7oOA/NOUp0gqyFHr34NwiZ+2nHyOOe7lRl7IOKCGeoiCdRQ7jOuO9MLVP9uJKnmKdPO7eX
Tdob4yzgREofcvaRvjE8OQWGjjKVfjYfHPfvJboRF8gtoyzKzHKu/Zwtj0j9oJTLgdHKDZYMeO2p
+1Fk3l9kSqC+sJBYU/wdt3T6mtGWybAy2pgURI//azupeLevrYZWkbEIklCE4TI97ih3xqyrx+fh
9sXNb1lwmnHl3ghOiPiHx63Ai8vxbVHyhUbOPlYLAeTkK+kScWajtOxPh9lc6kcCGHxTOo+dxhmX
W/4iOtKecFTW7zoMj5EvLN1z/SyJRXt92ttinsRQtp7qQqHYOnkFSX9oRLOoUTWofBR+dHmxs5j7
LZ8nwNc9iPv59vOuoYvCWgsa5p0Yfq1765keGzFIgm7yHtOkcWvPz5robtZelcx5Zuop8JIqVM6Y
Et8iE+E4frmsg0wLK7XoLpiWQ8CLagYPfRqPlQRodH16++6Fqm0+UciDrPGWk5QHqN7d0Lm1sGV9
1dC7UG6Jz3t5G4YU/AE+AzFVLd8StVSv45EsKB4jxQ+ZS95wDLEnPk6gCoAg4h2SQzNHOAOlWR4F
0GDY+cQGq9gv6XMWtVVLupmMKqPRMTmDPx6UyxO3LGpGMxaBx665Wy6pIiOzxr2ektgxdbCYtB7T
RcjTiKeUCRWH2F2n2Uw3bdDlW20NF8paOeMamAatJdp/EqBMHOqtCyvV5+ZNL+bkDpDsG2BPPF9G
0Pqv9oCJkr9Vf3kyD/7K7BtGXY5XDD3oiGEa5V1AWUwr+/8AHocShasdpwKC0WAXfGX5OHY0+jJF
8ra61ECsUnlX0+1XfavZlYd8xDbtGgoFRXZKE+uigd/An326OI4ZxG71lLyU6nTZeD6JKrZUseAM
QjO4kWS8P4iETO5RUIGUycfCJM+ZONeYy2ddLH/fcnkpe65rKMBsS6yUg5Aay3oi2ZV+ClHTdYCx
StPDg3+u15Fvjrlfy2JHTZvYeEykB/ImolOhktTZi+oacjofYM3YemZdHe/hW2BbT3OGCup4iQ/Y
czrl16kKz/hnan0Qxnxa4Dq1phSqB0xFqDBab9BFAMHNPpeUoop8QpXVCaoJbuWJ15N1/1pE1Nyb
a8uelq3YEvzb/eXRA0s9MleBo4hknUAoR58S9qDC686JZDkJpt0m0rDZWIZ6vp02Rsc5ItLM1ViR
vz1y+dN+4TcpK8OuGylNW9G5VlxtGUrGX47IW1tcKfM+nH/1LcI3gW/RS95RdD5LXeNTyJlTT31e
7RLOZ4mPpkngEPg+Ya0Mp+ewWY63rCLPtXRFLfrgrVDjcKehHl8OnqkSJYGgOQaCzPrgTghyC24h
eAG6hfwQYDrMVHjtO9Z+TOXcPFFsztHCFqwpMfwGs/HmTNCJhCrPa7FeOp0N5L0KEDPVVg0Anpq7
uwemnGJOkaV7u4hj/9VFiHEvIz/GkwNrHrgcg2KM56ZdvRk2GYtc2CbbOEW7dikzNUpM4zvwy2fi
k6vfSdskB8ol0fw5aEmUI76lxgQKbU/O2H0938ZCQrhM0AUmBpuSZyvV6UZm/EzB/Gh1a/B+ddrD
/Cq9Yzl1TLFSm/pkg+HFzKZiF9NDakm/98BPifVUO3lDsRGx+iNvyHtXESHYkYHCQRcmoi/Y2Nt/
bhp+0lBkS2rpmBPybYOHuTVoJHZkfnD27VTyngfkjBrWA2dmgxZRRupdXTxas4bJPCPBPIPguC7+
6x+OuejYyve+SSsWd2KWBOuJE1XgblqwItJ7H83xkClpsosLsPNrVlbbTeiHKYYavnJAiKD4y6GJ
oqayEJ82ZvMHauADRPNMa+eNrbJ8x4ybsHCWxjG5qcbJF0bhh/acBccru3s5AI20JRSdVGGqJPQ2
zD//N0dShQoJu0nVaJbPoNQc2WwKWkRpKRxl7VdsHwU3AcobuVUsV4ITlWIinxkjrx4oAVz01OvG
g/JxE0Ny5IC4xwyOPrSaES+4QW4uVzCTLpRNXdeZ/u+YTu1FcmxTyuBwWSr/X4qv2VUe6xRIrwRX
v+bKky9zu08retB3k6Ks/7zrel5n7EKeZSbc0j8Ct2gSf2udr75cXv9TvpAVG83oGsRBr9An91Qe
OybSQCqAFUyCoLxDdaAJbDoBT74JTO4GoX7NOsd0uJkVZ4mLWDS/2zCMCui89Q662+VOSAyJ25EJ
V81r32LPSnzT27pPicJeN9Y/MZRDttV/wPaAxVp2iQH8Xw0KKWNQlEUNb416efpBagMG3c8YRJH6
7ESwzlCarY/gwEEFDJW5kROjpATi1qnF1lLt+4SRa+3R7vwpUdgXi+3aKxJlqxYKtcCFOsPb8qYu
+oF6zhgBaVbUj8B7dI9hVm8HTDIn8pYCbCJPyY3yts9FFrZ0kg2mAYUmaFLn99F4FljtcjHFO+XC
4FGJVCPjjAANPlloChjN3xOPQkEteofRhIgSzQCciPfbuy0um8vlZTu8xDTc+wVBa0i+QksD5pjm
AzB3odmLa80C+Zeeg0RmYbrhwbeySUWpz2HhwZoVv9JrJmdpn3aysti12j0SzRZX4oaS8YWIlhFs
ThbD590oAFOWt9s7JE8JZDun+iR1xuAKaArrtTq9PEh6kIJO/twModkrwpdf+zG0EcH9CH/AY8ns
CAs+y5U1N68fbC1sg0D0KeR7gSx1+lBhKhWIBSPK5HqvQqQ09/cce9gvKFElWLvsu9ML/Z1Gh0FO
RBT2e+ixYSS/sTgIo1eIacskUXD53uI83WTTx0VwHME6BkyDuuDu9RhMERgjoneiWX80UoZ9QGrg
xDde8xGqgBT4MckOi9vFChlZjx7Z+pzRB0SI00E9kOv2Hx18FnbMOC+QVli0wfd/1Y/F/XnToNZc
MFJ6RwJd6RrEPVcQyCT6kj4mbLYnwaSphOAJ8rOG0XEvfhJTkPwpfHrLJLLhsNgpLk0vWw73C+SA
iS5opE1uCfrF+ZCmWgDIcsI5nVvb3IE8mb4F1aUaScGZZk7h/r+Mk97hOwxxrkmllUFpvk8Rc29v
dtAUd2CqqUZ3siuXz5c9v/o4TafiITPD27hu1CDwcFfqU9b1joPrnZ/90VqW6mVtn3+gk8Bt/FZk
ZsqLRt9NK+i2DRLsXLljOdMORHnDhSL2BiCxQNC0qWWjlQ28/0QY6AyM63xNpamaNaocFrpqzvj5
FjXmXALQOQEfXKE9OerXwKzD+dk6TnhJH/iBL3TZcOvfd2JQ3UvbW4hXloe5lV1krpCvw8+3WTxp
TbCIdK3pioGaQ56dduEKhhB7GcF6pKeVUN1HoCGe+df0ENoZT1cx/j3Sq+8EFV/y47vvKq3OT9vv
sZ9Pp+8fFK2UJaI3vS7y8Grb8tTGjJ6hf7hPFu/lR3Dcs3fjvNc3E/xAuy2ADwbPGHDNRaHUvMGf
Z/azqrLYoe6C0IPI47suMA55d5H4oAQxXwy/6MY9n1yyPM7yfdCEHmAC/EvwFITJzIdcsh2XJPrq
gXDranhw2/jYiKXHkkbQ1dTZtlaxHjAnN9UJ1aHlPzQgcyDcghOzQ9EfdZZh6B8Mxn/htJGxNFYk
D/Y/1XWdAGcApKz8m/aBSsDwxtWBcSCeprkTW816BpUWpvvx7y54yY7pU844Zmgj+DnRsPKkj9mZ
gRK7xGUOXiSMRQCi+ff/RGFEahsUlp6bUlGJ9USwQfNn33O8FwSGM1zoSQVyokEgXI5RThGq5rDW
bLepyT7drfjYXpzJlVcKZTothJ92SanDf2AQK7CdkxEtbpv9+Q6M1Y232Hojypb9O3YSaum3vhP1
YmYim5T86iJr6a3YdcCnw028yNOKZMW2qjYVp5PUGblFiLXoQedAcDUMoRvAFUikSW6OVOKOA/4k
XLAs+kAEdzPUwXPBvy2FOMz4iApjXFZnxCRk3GTXcK1BNyTh7z3DqqUfn4u0Wk9g5CsTmte6s37Y
uOiHUILfAg/K083qvwuhDRk6F5FdOXJbcustDHjds7pz1mSkgw55hcODpXxi+nqPdhxYH9sAEqYU
AfpuvOAZC8BNXGuugluNaTPNNotl+wemU4K7PqAdxP9NiF50F+DxsL+bAiTHP3qjXRsdm+j72DKP
t8ilIL4KHK6BM7td0ogjIlkiY2EwW6fRS4SvFHuN9e/MWZbjnPpg1K6TzmTCuRJeQJsdl7N4WaSb
++r6Slo2OPn03de+wHs5WWz74AG21SisizEo46vffsVm5kI8UtNbrHBK/NPmRMg2sK6FTtkD7LrZ
hn11rRTRil1wQIu5DMotwG7slpgfF+GDR5bR1huIp837jRHf8VrM8sBuhi9XqgSz7E/js9oy5ls+
9QECjzjVqfLyqiOmz6oia3awk0agbNyqzEFz53P/wNNT938BrkYJ4ACVxg6p0+Q/ZTRlb+1TO9gb
3/rPH4quwXTqlT46ifFuVLepanroVivo+qgBnB4WGEZE5+JCwXGUwEQ8sJsJdL17KRJtUSra/rd4
CmbRW6pvV1OM+NSzOQrus40iZ0TDQIhvUyjSBFcDYXM1EsL6BH4wgE6TNS+HNqnQyziZPIsQe5HQ
1f9go9H3o0oHL2K6/e4GME1QXSOxB5B9VpPRh49iD2Z0jvGMTOScO0VC+/XOOlWeeEMAvY2mTujr
TzPuDomg4bO5aAcVZUSTa+QlruzGpYh5OlI3x8Eg8oYsBSpzHDpowrrit1akCQtJuItfW6aYaJzZ
vpMf5nCBbN/o3fkFid4yUJGtgJUyjkUkMSVGM6HJY+N6uUxL2IMJo1L9MXB+UJPHbImtZrgAmOjb
UFEExBd/UjtmBGHso5ohAor30dwZ/nl4wO6yz7NrWIZn1XPXbSV6Bh2E2rB1nR8cgZY4wLmNVIwU
x4k25DFKnARB7azLjxzKGx+9NKQiXH2iuUSrAAMJ2+lISe4KGr+K/9eA2fL0K44pue8pKnJLsq1X
Ih/pnrDBk9SwJm1C8jfwSnuiEO96aHzruGnD9bS8nGsNxTDiEqN/aifCxBCo2bkRqq0OrEWCrNWh
08aibuuQ1Dp7wsOpuSXyhi77dxPo/gavAGZF8lXbdC22P27MO/RKoSRwprjV+Ea30qumaxtuTuXc
xlryhsl8S8/TC79n//Y1/J4AmFcNZt+iDq2V0AyJCs8dYWFH8UUrm9rWKA1auvgkKdE9MV3l/mJf
ZuDl+x3Mc0nuQVvXIM0IUkonMZS8kqQg2dPtYI4aFbZzl6es9k7+5ubX3pKWjpMw2HX1gLAVyFy4
Du4m4psOxoqrEfTANxD4AM0Kq0Zeejf6pRF+2TkEu6wjZHd9WQ6T45bAnLMwpTTHe9VSad2KjKB+
/Nnh5A1xyyw2HeRac8V0ibB2qVHqK3UjBW7t1cLa+E5bULI693BumMrgkPJLt+M5hqynfxZOd3BG
WoqBYdza4n4xfn4nC3T7LsJNz5zlB0pAfTK82RqoIpFn0D7AAfGa7eTaut626bq5x0Ra+HiQt6IZ
jhEMMrcHUtk7M6UdNgTS/cHaxBfccJvHLphsycbtT/YzguhrJgn6aJP1zXr0/DRNhBMSMeP3vO5S
9ugCn0hZXcxLXPmXXNXmMgU9EfLeChbW2OEAFxdKRhR2ufjf7x2ROOm/5CJ4TmHoUvr5WucsPAze
KGHRZAfS9vAHtf4AfwHr2qU/HT3sqc5fwjxyHMuU1HxPHVHG+iKkDhpqgFDdUDpStmzXF3/p7OE2
lMpekkd+zGBUiWFaqsNfnlK41367MTF/CjQo0eYE5YUXUA0kWC9g39E2j1WcwgnkAanfwYyMi5cb
C+6wS+f9d43mPEkfGOnGCH7MxViGF2hw6hTDcnIPOPUQzwixN2EW3pJyicEowCqsbFETohOxU0u9
9jlK7Mv+uf0wT6q1R0bnSbHMHK8QyfNGkVkuEoEnXsMDMfgc6ZhuMTgWc152RsWlqX4Gfv3ru0zH
qpFn8+SaNNg5pfFoEDMqFvq4KLGsFkzWZs2xNTF2+m/a2k9KwafT6qQg01hkcanuJ88FMSuKYTCy
ZJPZJUOHt9hj/yqjZJJs/PTp42F8HN6qNTwyNj3zxuhaHdI9VsF+ck7nMMsFY3ttyXhxNPgA7qEi
MBZaFmim3v2qGUT67OaF4kemzYiI9njg8bciu/H4ePiExK16/mDWNtTHHpJTx3w51xZtSIMb94Td
+TbI90Jwga9ZoGd/TB6YIzQ6Qd9NmrZ8lcCNo45i6aw/NyYxFVcPjrA/wOKlTHXC9jJaqQkgSl94
u+pwWoZuhKoLnBPib2miLdgsouZfVjv40EHlT/A5aUQLhh77Xv1U/Z4IAPm7aCJH4GchrDfIKCa2
Jhvvn0rkelyw1LfHeWGjc/0+/C7+bWxwFaIl21gvmaCBwWSkfTSyqkL5DnHmZ6bFIU8eZ2n144Aj
dkLlDWiDctelFlfvFK1NYwJOHb7pEySQGtVsBNS9cNYEZ9Abfr7/R7tgmDTPeXNNsHRNnV0ktH56
hrRtpsTfthJNFxJMPrfBtgx9xXlB1IY/oSvFM7ri0gE66yxTPRhlBCIDxiCeVMi6rdLeCXlpLvF6
ZS495nV7IMau/zO8VXoCH5+jf/QLjpWu3m8JohMEe+OJkxUNUpNR8QbMSr+3nW4VYNQupe0IQYDe
WL5Jrt3jujHmvvS6j1Nl2eCjBXFWZv9PJT32Uo4cutNGooTZTeqHivqtwee9KRJEeChLq1HfnSfa
3x4wpajCa70sRDRRFQEVpp/G3W+QC048SA1EVzVzZbiv71DcpYbjEsx3ZXzds/QhBSZDUU5G7oSv
itS0WZkBV64yq9FnVbayD+cC+6hnl7EGfxI95MiMl7NvdQ7ZsPPJeYooMJblbeP3s4okeY1L9jGH
R53Njaf+RBEEQx3rmmuLpfMnAiKx1/l+vEDHSEVYvhdlCoEaGeSJrAfK50fXdFQb5Asraa3CcglM
rIXNqAluEIjcbPkpSN0yiEeazf5zEEso9HMJa5tcFiGchKzRUs7FH9uVE42frwM1AwhKGZxIri3p
CyheGrZ8Eo4Grg7PvO89FlBo7qDWwuCitfjZb6RD7XPhSNAF7OvTnwZpX16PMiANfOhP3hpSzP09
5yCqQ4SYNve6vpYyQWKhznKqFqPyPu1rDfJYFwCBto9mvx0t3lRzO3Qs0bl3wEGofnJtmlNn63F+
WDHU4c1LNHtrVNyAZf47MsohH44gIt8X0mNPzYF2V+xLM8k4OGSX5CxKQiZou6pBqiPUvjmzEplT
K55k5yelZazHIbrmMRnoxMRYtjTGblUN/M3zsTF1YmNMtD+g3LXQu6nS6W3EjjuKIxb9BOGPCv28
+2vkCFOWKP3uqJNT9LD8US1ilNJbUGYC3ypb+Y2hbEcPzlvISwDQxs3NbQ/eMMf4cDDM/gFH136y
0DStq+AyT1Ho4GHhWMOkciUCxrk4ukc9LQsy/P+wjUcoM7HX2Aya0nPrI36U1+Ca3kMrwbgAO6nI
g/OdEgrERh5+rZE4PwCH+Rv2mcQI0X0RC1mhaXc5X6FABhaQTySVfhfKxf0AXHVKTAy/51NWnVjG
DMr1ykUUyOBKLgcLEconpM99YT2DxmUbbIQlPWETGEXT4FX0/4dn03LXyErvPWkrk18w++GQC6q7
wTryQvTS1qLiNd1GxwsCfUKBukgtuJZ/ihYUk2l6syuhhV6XebX5KVpr2p2KRbKTi6vwlxXSTQwK
tYGY7jKxcE8QQBsl6htck6/wv3g3kpK8mYSpDHZ32n42bMdUSYosepLikqT+GAA9nz8OlpTAK52g
iFJjQGXSzLj1zQ1sHdz633pAyIdt4dpvuJz+20lp3sWiUrF6B2JsHy/TuClM94iFoz06WePAxQzB
Dl+15+QX4DsTE0PN/MSfqDkmZnOU3eQwpVGPzHPg/4VSUpzKKyAyH5/KOZdSaYRbPw6eNXf28dVL
nJI/Swak8/7FqqHZOHZMFB1rP/CHxexM8piHDufRtCFQyMa5BxMbj82etwglBrfvqrteo1lrunON
Si//gPdH2e7pevgoFnZGuSRA4ihcXXOUgTUhFBlIMuBIM6XvGKh04FpvvNhp3rIUZvL9ZCd7c+h6
8a1GA1c5e8xtor/L9eRPC/6akLQ4QVQZeZENYE9KdQQTTRsmN1LzzcJx+uzNWh1gfgfV3c9zKIA1
eqIjCyC50RjYTN1nsHi7b/iEEIsU9/x3EiaOFl0oHXkQtVPRt0RI0fZdxexHmAT4M9H1bwOKlMAR
4E/+IbWuLY9IEPJacncZHyByfrckyIdZWUJmPLKubeXWwQDZJaMLUnugPlI1gnHhwG+XQdvYgbYR
M7iNhzZOLIqoLuJ1jjhPPheqPpmbD8ZCGv0D5sg+y0TI6lQpM08anVRjJQJWQAzYhWXjh3jiLbmN
P8G/D4lPlnLD6M93wY8HmXo/xs/okF2ZXPVvRubDBGbZK0UZ+fLNAkCZhBUrgYF/Vw1phIa4lRKq
VPzYABlTNTHN9JXJRN/gglgj0PDb43nuO/1xAF2SBhCUwArJYSr9TUSN4d1O38mjc/C2c0e/8R1C
e/gmn4WHysvf7uyQ4kunQKw+Fg7qR/Z8NSMTd/TUktIuYN8hNF1/dAibMRupCSUKDRsZsb4Ng/3Z
RmewWV7Vz0voLOtOPBNnYTPM14jFD/KFBhvsRsE+9y2C3es5OmsuG3BTrqq9XZGJbKkF68JafE9B
be0No9OY1AXVq9xxiGvYrcI/xKF2uqJFiEGE7ThY6IlLoAwMHQLJelRr+90mlptoJnDNgnyI6zpl
njey1OMNNB0UiQeqeXj68zwupi4CwzidnBuRWtbqFsOR+MzVaoMIW5NaV5PogekGAULlBFSz8VZQ
QO85ySX30Kwnm5v1Yvoy9RWYsej4kpRCX7MmpBxqH0B90z64xixbHG1bOPe3n/kBEAONt2AAIq1D
uxFaMloRVVfez54K1Dr2O8zhrnWyksEN+cDaz5NUFCeQODo9YlQ7nXEDYxRPRbZGkqtFbB8i6twQ
UBrwsHibDURRHHUBVxpIUM9Rmvq+TAPaMacvbCYDV+qznn4SvaYdGJyD7kReJD4gl81zagJshPvO
dQyyAFkXSXF6FAFzQt9zygF+K1l35zVGkgT79WI43UJ6H/NX4FQEteP7hW0e8KsQe5xZrVkZ1wI5
RGBqF3M8xta3Wyh0EguChgyaWfzMpXo+Rw8gjFJiQIlUwfcJNNHsFOU0CwI5Qs73X3CJdXIroSnI
u2fLp2Dv5ml44d2/j0/FKjBG9m+ghephH+H+nVCbM+9GykxletYHtpr94Bqp2dvYWMX5o3A+aBEL
wwt9MY23Y4XF1W02qO8urr28GkqgIBfTynQix/QYZF+O6r9ro483u/LaW4CuqIXI+gZ7vVPD/v4+
JLFDX5ssi8KGCm9syaf9FiTEo3xwvjIpZYy8EPmErOntGYRESmWLmZVQKhXxDiWa43Tvdl57Rmaj
OJRGlbIQNcvHgRUn0HzD2oVesvMeFGmAMh8XNUc/cKbOJi6EQ2tM3RU9uQW3PB+A4nYjZUVnKFi/
Grda4k8wyb/RWRB3SAxPggqpWMHoj+OP3mrCi3BvLxeTQkuCddryJ5m7OXoZh9f/xe9jH+gCoItt
ANmjz25SU20LfjLco1FWSH2Ndr2jvY6WCnLJI4ON8ubvyhNgxi02xmHphLF09S/sKCmTXPtX0YJs
CvjXrQ7vzeuTtAr5+KVd1iVAUYwJKGs0/I7klBOLxG6Hr4B5J+EvOrPJ0Z/jM7XuTFN9/4kgdHdO
sHShNHdhitW03z2z6Ok+iVDZMBsv0if8l+bulKMA1puq1rxKYZ088VkT+ApwOM132q97cOjiSKZA
M+D6YA6bsnYBrrDHp2QLGe3x/loZwClP1DuB8T03AN8KePI+oTsqLC1N50wpk5TFWZkMmkwl5HVt
PxR+jjnX9SdlRng3PVY7CPpANANaXtc+hmQDPSa+iKRXxPZK0vp9MreT0A+R/MEBhQuSsJcImS/4
q0BrpXSpACo2kTYZdDTdfPpXbw9NswRviuZT4+64bGeSaTCuIPwMXGkk2cKoTB/otS4S/R6PvBfe
8PhMAQkFX7pof78YzZaB/OgehTcTpHqdjvY3PWwqJfHU95pQJZ744ZQeP5enIBQqROJox6Z260VK
29d7wVyOdFGKC3NDbw8ySNGcO8U9uKQ71ZcKkuItrQ3Pl3CsMKsMAfHe93Is8ZDmzC9vJEGaK1sR
ZVTTgBdVOBBfAxYdi/WK5dQOD95hUe0g9HehmsUGksZ6X9aK6vOuyXaRg24qJmkIUt7r7NbjVNIy
5F9rMVeJq8qHNhRhImyG0x/nDqpZhpuHcAYMChs5lFcqZWgV13bWVV1QvSYwVqxA1opwlz3Dgm15
sahIC/FQi6jeoRzhg67JPfNcu8ErR5o3HAiP2PUuD99pO8CSW7Ot91g1YNEWvIpbcxnxnByDxW7P
aXROoUpkMnk+uOypWN2jE9YYqTWG66MuH3LkRdFaL2QbLO+3/oijCq7+4Ejpih8i9P2AI3Pr27J3
/LvrTAALzHnTiTK3paAv9TCU9OKeWuE5aCRDKaLXW4Qh1OALrM5OhH4XYu4EkRntarq0N/we/GXo
tD5uol0idDBKYco+KPKZXdcStHBR3A6DBQEsUgcVC2GoRFWPg2iwYFuqkdvuuV38IEBQ5ypdIpci
UXwIrQrq456LKPX99Mw5AEB+kadf1//7QQRx5N5nXf5MSI60uO7+dExMqss99UzPDTbIEnlNrkuo
gJIZALJHRvAnFfBvtP2/zx/qUJOvQOlObVw4iTVn/hi3MffhS8N0jQ10NPKJfdCott9YNMrYC5I/
NiFF1w4rVz5wx4WUbocBTFvf1ApPARRCsKie+5XnWYyQEw0Tr0qIbwdBiNOgcj8qPI2hQ8sFxg/b
ZmOJf7zLC6pfVXEBsMz8/fsbIY5DZdeTmgUCHg1wgSE8wLXK7UqF3uF41C64ew+JnrdkgTsmQOin
rr0Ng5JBjBJTv4xwpT8rYnKiKgg63kasqEeJyNAKucXhS2Skqx5FE6sPkgCNHedeaZHIC0s1szBG
hfki9ErS9oRzX2SW5N9TikYMyVqofHNJrIVgeh6bBZrYoDzAZgX/u6HW+8TdsybiZIPTPJywvxfs
rtinwQR5yIdqzk05JiaJLMiVuq3l9DAVNgJX4chwtQg61ywP8JY8jpcY1lcURe915M/3MmYDd0Q8
SZNAtvbnrxmyMEAr4HBaEC/7h6p++HCQs76zL54MFeCXf05T3ESH8l5VrxH1K6xELHb4uh02ms2N
UEeWtxxvIM9/8H/GlzjJ4IjrTaaDSF+i4e4Xqm3v03ytsJ3aaCPZyDv22mrTPbBnjb5b8vS5j3nx
lGcbqh5qjpZoBbKGK11ubpo7sX7dAPNnCq9ctxuygn6Z6CvY03N4J0gHQre44RDDZKIxkJCWiXxm
qwAVcolxoKldW9Zq9bmNaOcUXddwZL74ZPs9IqonYwu8/UzyIpU9Zl/9uMLnAZLVhKQEFupDyMF1
lLnuGG+PhoPl0t2i09krm7M4YRi4j4yH+wGdx57SxuwKdA6lqMB7wpowe7vDiLPNkFYSqKJjCoj5
yNkKuN10ELUx39nqk6QjTp785hAbTrYpbn5ycHDQENIp5zFNqBoJ1oSA3oBvYE3v4JyWQdTwx3eW
Q/qLQP25ZkdPjq8r3liG+MfhdGjZjijEhe5j87xKXkKuEKgTBqIUFMQD/mgmJgDfuPZsgo6F+uW7
m3DIsDNxkF6OPokH4rS8rfF7LB0fzFVSdAF24p3NozBjFYKSpAhL0vCtwtiZm01SQw0epaPXGPNu
tBdbRJJYvpQ9mjpCeJAJK8+PLKxCMy+B/BD+7bKvtrmy+fCC225c4P+DUbmcZIXKsOWGCMAZkpc5
7krPEogU2qYBbG321Gk9WJfNjWO1LPjmB0Uz41hMd15YVBQPFNE22Q29vghR8VttrweaHvnxv9iN
/RC3h1e0FRVWRKJeybE49tEUFCgXeVMNgHOT51TORpTeKqGjRuH6cqrYBSGfHw2mI4uCrNHix5EW
g/ekHom70t1EOiucLpd2A68TaFfGmXvOwEAGeTMfgbDxUsiL8yzLOXAFU30HBiywIyFCCDynUNKD
4V2Bv+VLv/7zh9qmh5tzwZKtG3BB4JnlhDzP3X3enAh0aNJqYqgecMS/DXBfqy6XDA5mi8Gb/LGj
yAnvFXbqO2qZfuCP73OCs4FFvuaMsjjLaLTE0HP+PAz4aiBD8pVqT58cmGM+w3Fxkjbsvg/aGZKi
Z2QsWy1O9enb1jQSu/jVDH8zHv90JGrwjRHVuBZKRxaE7tRyHx6XPg+KF5QGHCKJmqziubmEdcf1
ps647z/7XIBY6aj2CRaMYL4DkQ5kjeSSxKUSUlvWo9mxUjfwkpOzFLfrRyRHwRbDDR9WWzc1dOzt
RjuOI7WidpYLtiEGjkad7VvCM6m28DkQ+lV258MMq3S3mY6BGNkwPjJq/6kUUI/fgWTQtDFiATv0
b6c50rPc0UQox1enf4fLAsj0gQGb2nMp9zeL7Bedk4eJQfFc4LDs2BeveOV6rjK4CZ1SP8S7GvNQ
SdDAUam9xBZXgC/AhF0S6jwFuR7zRwA+rn852Mw5XIv3uDyT2nhmvh+5bDWIxR7u4da+1JmJjwUh
KDE1lnwEpYE9ns/lYobor0X8lDYuWJhaL9qTBqxD3Cf/2WIGAp9Z3rkr8i//CKGDrMYzMGjByflk
XFjE/waAZqZttC3c3wBMhTyYF6owtfkUADKr2zju4Sx3EaAetl768ozkBONdEDfpQ9F/KsBQQvma
/kJgl5h74oFulrURRhZKtbE27DyExcyOufUT7otOiyO1bDdvH928fqoXe0mGy6VsiI0QqjWwJBtY
7Kbii6nQMoJUjnU2IpxvmgZMBsWci9+6/zdEOygLtA9ovZ4RCLWu3P1VXeLG884LoMCL0GVmLg5L
nMkvKnJOu97i++6fiX/k0h6vW6BfNTMtBmh/s/fDEvT+tlmD5WTtxNmOt+CwkM0p8+XZ8sUhVBH1
PfSjRpcUdyYbulSJdhkdfRLKTKX3JRa4/YEpGeZpq1/Fuwoh4wc/R20U2DyeFkbuGXoAB/oG6L5K
tJq/QpXzR3Mr1QVshMt2gG0Owu2ocpa31OdALkpw6zmz6rBSSCZXQBz4Ld1pBohgQyczdyvI2VlE
qbP2lgHJK5RAcwfo/JPskDlFzpbKgaA9uBz4puiYqXbD5HOeRWbMw17K6x3YOSC+7qzWREPAayYG
ob+JWpmlQL/s+ma4XkHeI+B/CFs93X07cs4Zun7sXhIrIMSWmzu8f/yehsaU5BLkIQvNX0lbFS6S
z8KO+LPeVtC2yCe56ixayu3M4QKIReXnmZxQHDecFVBi0NMov35SSykDSUR/Ltyoa7whz2HinrP+
+pmV9LjE8SKOaosohRzR2cSVU7fIddY8yBNJrRRoBoS13yox+hdUG3LOsbjCA5YAzu4Jg7e80PFF
I+21j+eUH951hS3n8dxZpUVx6EqMM3VjERTBleey/Sh6CaWuVujdqoGmABbqAMv+Q6+ft4B6MSap
NIWeRy4/gdDpeU51wSJJUkM2ZXbCHFrrrGHMIGX0AiAMQx1LrSFW41WGsypUFrP+G8PQVHcRgYVN
ZVqFzrqe3bTcqeeagmVq+9Ueou9bKIbGLSt1Gn1bgwmmKDmGi0fPV19EtnpHC61ZzmWCwY8x3Bm8
BUkv8dkwZ498vMxhWB4KPtDCG3ghq+SU/pUzfSxovVVQnu6bjdLI9YcTieDBo0qA/FhvArVwU2a/
ckh5F3G5BmT0U1n9I0sz/1gGX3L9Oq/epaXQvvIObCWFwhzFla8C9+QEIvPaP9aZLoipBQv8ypvk
ocMcelcm7OFbN6U2lSsVTeQGWZdBBNlSBpA3eHlaKRiaQDo9le88mDtaGY+sATQ6ThElIBLCXcLs
UgiPZrV7l+0JNxBv/z1Ht0QwAPFpGepib6w1I/eLfWdY4zlvd6J6oUgjyO14FLRtxgUdveVXuSUK
4OLLqgmmZ7Oomav8m56tKL574AoFdECwjv4jgF4uOjHVafllXkepx6ooTkkoDVDTF1gqD1WTpnQc
garymQK0l0KWMHbqEBmrjk6620z1Vn4mNTYSRDxvkGa33bCg56azb08VfwmMIN66h9LJBSMVPlFO
/JjTYCLWcfXZ7erDIgXgcDO8SufHTraDWFHOfAvuqBU+iiHHn90uNf3nW038Dv287L63ENWOm2Xx
lJgrhbmh/M4WeQlaBhfLjma3ANcf7lEYIBokMsmJd0dAXyrCwtZLDN0dLUzlv6RwzG61bGHG0KhB
vTDgOEYL8CqOdEXR2+9UhDPnNilkJIcGm7cJxv5+Ny3UsYg2BWMeENlK4J+Q3jn4T2ptIktkIBHL
h4dYEcAWYH/Lt5G2HNc4RRtQ9HjJzETiHEidG1nfH0BJ9NB78b6upkO7Rj9LViODeaNdEXEJwisN
Oa7rpJAQk54CyzTl41/7FcV2SlZ8z4LSfsXBcO09hMBHAkjDEDDTeqScYp/juvvNTVgOV3ZiXZvJ
Yh1+aOEXLylg2b0cxgpDqXY+lpZCzY21JDibk1Mp01nReCuKlC7TMCqFV6OnQ9RKcgXEdhAykSBV
A9pddbg1TTg2PM90LWNQ23zwq8lTsTe/VceJ7R00ehrv/uQSfPnTLCtRF/u4HO1PNm1Id0fYXzIz
wMc0HBxiitrKu6pl+j/6RHMBBO4Mr4XOCYRedJHbGOfIyNoSAPVcHd6WAAGqqDvpKSmd2wjb2T3s
XryVkFJ66XQWphablO9pkAkvXtBSD1m+zUww8qC8hHotdvFFhuDX6JNaONVPR+jpL9jdADubeZXW
UrYQzHLlOGSqezSe0iu5bt+ThCUnoijz4u1VR3S0uaE4iVSIrGUjmLE1NuhkqcCjcvZmAYG7jqVc
GvW3rPtj0T6BNQU1r+HndBcXBWKBGFO2Nfa0ksU4dWutgvcPFzrpxjbCdCfcNWf3Fp7FZTVvakIq
U+Y7QNIVWTLsu1rGcs9bOUktfs9Fv9wZ8edr7w1B+prbg8CkWTTar9CstUXlj3SyEiGIMebW1DA8
Q/lBe2wvNiKQJPD27uISYNPSjPQq7LpReeiY2aDVsdxBiiYgFvWFCcGwzIMbuvTBkhd1LJngn73L
Pa8IOAInrngov5miFM42loY0gGNP78K/p9s06d1bKK5/ms5Fx7WBvvTDj6uU4MOBDSQa8LuBljf5
/ZNmlA0G4kvY3BSLMt9tPRggqm1yfotwZX5XfcTn/8nabBCSvVtqqDdc+o/CBSNG6REJaJgzIgU8
4cutr4R1Vy3/ax373xRIpNJigk0nOTONunCe+36/QjeAQlV00u30K0hwNfGUkHGm1ZnqJ6JzsrbH
ucvgZ0tALMdqX3A9Hq35fEsAdRanYto7Pa1BziA+mqs1mlv2FOiebi9VxV2BLkRe74+ytP2iHFWR
Gy9Y/0WN0G7X+vhwgZrGuD0x0mLyW7IlGVwcHhGCzSXFgRqV7ohobHWwbtwAuiMrONJdewYIPaiH
CAcwv95gNAgr1qmLIuxZklzryYW664COMlTZdOLkROtLDUvoNnpgGR5f+1PV5fdEcZcwCG6yO8+N
5jN1NWCiNPvX7ci2EwnUt3Iqi12fDDM39rU0JwQHVUUrJC8PnMLsvIRE2fAVRGXRjwUcRUxAskBt
gG47IPf725+DnBLpl34IduLLABGQ0hf9EqGsZs+AHo3Z/bzw2jLikZa6tX0xy0m2qRUjq783rG6p
Cjj9ZWHhycdNn/bZMcfTYsgiM+kxo/l77XDxS96oknaZ95HjFfy9E3AadE1R4CIZU0SnSl/VpSql
6tqfyqqkBwBBujeMBTQkY1eiPXXMJdiBccVTRkNbsU0YaiLA89ium2DZdwvJmS5eWAGNDUCT4yQU
bPp7c94SxDIBpfSIKAjNdemOzjxtDLSHw5/tUlXWMgCmylO3HslUbeQDNyTNjkwRCNkGbS+MvXkn
3TUQKE3mMFy7ilWAuj+IVYRPVwsjBwG0uPGxcogbjmun4voVCXap6PyGa0Y1Zs3KF+z51Zf8GaO3
jlg+sBsEPIU0l9AJtyVGg+l445fJSsTZAhF2YB1B9RkdJ9YawApRYrcEFE5gGgt3ghg+TCgW2NOX
TjzGxVMm9+gZ+sDSaSu+B5bYOdRq0vUljGfedZWlnpKvAoWcq77jahoCeSBpCUqfppesmEB/0SMx
I6fh43rxNxgFsZG6rlCoHaoEueynhanbKjHQ4AVN0ICDdXKX5sdx4Wuc9vGvy5AJCPFTzRE65GCG
QPv0hgsJ0DUInikSkFXlb1QZuCe6b2yeF7TZQyo52gC5mg8a4vZWTEQT4e8Z+D/mUCbrg51pndXn
LFUTFB3SPHCl/fZb5XY2d+bRh2ty8WIlJMYlCnO3mVmhzrtnuAQcRnHSeeP37bhwVIfhlV+mgyQt
61OcrueJE8omhv/84MO8mv1L6vKvj2EuPUY/SLgU5cGSfnZCPUqSUHaeNhVNOc/laqoL6vKgoDEc
6jNJmoQPNoHwz+c4ZFccQEn20cy1Jw0ATf32PWPW9WOF1Y5OZeDUBiEpLGjDXdULN3Ubjq33vXic
E8kzCbJbJVO7je0LvWZ+l9SI+DYXXVicowCzOd7xdRG0zQvT1K4und7DJdvRwH3HabHaN2v10nP1
gKTjJjuy9iNTyR1rYIa2zNB7Gnkmhk1HE9nKXo3vOpwHNgBXvZiQaGH+IVMn3cgyLU927HhsgrO8
QJ7JNYfQNamoVCQJLH6elu1qK3JONt17V7xstZcRb0IwSaBhEmQ5qPJsXRTp+I9i4tWP4RIN2tud
4qnVZ/R9p9+bJ76I1aoEC7fC+hcRPJFwTI3yifNEyu9ssc92ink6sw6b6+GK6IKJHDaIoYr0HAr9
XOX+ak6uatAW/3oVJcQvgUUO21Mefu8hoId7W/VnZJTOzN9y+IbTWm6khmDKjxyB3mxf9av9yezb
tVbQbTwb5Te0szzLJgasrLFWGuBBBQ3bGhNRuFAXsAhsi9toVJ/ZnhAB6BVDbKTmTGh3jAF37unY
uzedrUk1X+kcTad/PHNTiOs/anI6MoG9Jbr4TIuC3qveIfwvZJRjk8djNXeLwLVKLAZesH749phr
cMBOyUr7ADFl1gDNJi+uK3U3//hYJLjV8smDRyDK7JSBYRAJ7MqcHFQQxHaYNhoT5jca9HgbVvqa
WlIg7+1CLV1twrLfLp2d7JXPvQEf+8z1VwQgMHHFds+qhKow3pYJZrm/XezzZexS2UlrJ2O3CLhV
lHVQtjV7OM8J5s0ZQ2RrcFK319dQKjlX2+90qdP5IRqSiqzqIfKVLvrBMChf3NwPVSwcOHtJn9vi
sFkVjT5IeoFrbxL4/3g5LKTAbf8yQIxP01Wj/6hDzbaYQnlyMDTbyHvLdDTbOc4YLTkpFEgVHHE9
uc5f35DlO2yxzShnyYNpkgYmz+6WUJWU+fV8ESaGnZ5xYTbXmDObww6cSTUGoOfNyvOPYRHx3ZzK
wjPpDzKKq4QsJli1FlGrOG5XpGGy7LeYxMcCfbnXDi3LxcqVwworcH+YpJu6dthHm7B6rsLdv4kY
8QjhA0Q8LlUenFAoixQryFuJyyWXbllCE+drRyX82ehP0zPBdh1mHLpPOTAGqoKG48O8keq9pnU2
2n1SBuvAPc24fplRpwmz6D0Y8+nyf/DXireDRHgb/dncPguf0yvD15Cz7scwoGZ01mgkRIVTuWiF
Nz2CELlxKDyh4EhuGU1k7KDaESiE9Lo8UMQnMe8fWELVNFhi93+47ljhVHuKjHnoBVpxkoB4ZNu6
OZr1u0eYqZBCg4x4mcNcxiwRSVIep69ssOMK6Vfko4PSMZQNwQMb12rc2bXZ6YTQTvrKmgHCQ2fo
Tsr4E6yiaecCHMlsAR/2XjAjdQg3Hejipo2bjkHsw8INc1i8/YU557hFRu00YncudFg1mhgNokxw
88iQfoZ0srNGKKS3nD1LF7YqOqZiU4Vq7sP86hL5I0W+jIOPXYu6v9o9Z20cVCBY8hg03YcaCaUH
dfLhe/+9GqHhDJt0JmZm455detELPWd3mRCSKloeOwQRFTyho1OVs+OC3+mwD6hzLgptjXTZeU/g
UhvD7itvv8Io9Q7oykuI60GSayNz/EREN+Vh++3WCDlis7gQO0kY9OVBmw/fKFctOI9IU4ytNUYP
oYkNr3Jgzl5PnBlmEK3HwjJ0nFcbT7qQEjw4C04ZLwLjAiZpjVZHCB4BxuhZXjvTl3tlQeL4Uk2K
8mxC57rnkMBmy7s/N3jTR3aNyP7ZK4cYRXESWYHF4w7+J6YrVP+ibFLD7h8icNfkWcEzA9qxMCU4
BGuzwbyORP5yT+8XBkCyAvP8BvNByKJ2hzk7DhVHB7xeVhY1et5rFZGUPSf5fhExmkeq8TCoUPqx
BZ/K8JFY6tqb/AYbubWHCqDYDvZQ277+OiHgbBHMKTG64wE6R45BH6eR7qNcUkP8sx3duvEN3rNo
aHLKQrvjrxbilw3D4QVx3zOMzlXZt5sQ2AbtWA5XMgcrFnoPcFoIpwTbhfFRmeQ/OhaWtqhuj+Go
qDQgxsNMWfnIWxumIkvmLe5PlRnpanZ6PNsZn33OPM4i/t7rt2QXM3KTScTnSYkx7pNRxwI9DNFt
MQTCPDypbp1frmkev2gWBVjJCCm8pzA5XiKMWtNwU8JsqkXNVxdpXeI4fGba9y5HXnexL5QoTI0x
dOUYlAl1Kg+nf0QLXmH18qzfvcDGipGRsvB60lyrhHDU/2j/WY3vm0M48icuamdD0IUsuG6OGwdj
GAyQN+Ce0AfL+QpBVARDE2UZ45OzIYWy98CIBk/RBTUffbL4ZgF9JC0s3cJxpn07K1dUJYic90wO
FZkCCb6qETarsOrg8vNIFbvuyyweoOps7JpqHgdF17bZUOAE0HCfSDH4A35b9V3bIYZW44g6P+P5
brM/3bZ+eUoP2kIvjRTXGTSOiIyZMRrx+HStcm3wsWbuqhNzAFQVuGHMdTUSvZC9U0ExcrF7izff
pyg/4WUQlHATgSHuJzfuWj1GDltpJfNFEUvKmvYwNyzVgiMWexOHjYjQP9t4UF/5yj6aGcTysaJD
Mer3cbb5GejsyeyrpkKr1KsT1DWa1nNjKXXguihpVyG4cS57tqOc0fqdUdrnw7/pWrSH8S5k7U1w
JT5Cc4Xzr+4Otxp0kJbZAxI0ELlP5MptoWG+mYK51j6CvuGoB6PUgnlDXgmB9vZ6AEp550qV0Mxc
cBpYIPnlch1wgUZ3bfoTtS/Kr/JMXiiIE0pp+X4taGtBMjxVbC17dSXvrdXQhsFvGm9A+plGN+ts
g3RzP5k7k08N01VUbuPfDHeLW2qDEf2oY2oW1UcNyjPm3qulYVdDhwyU7257Wedi9nxHSpH3qLN8
NKXgNOyieBJH80FMmdExwLMtfubDGa6cS9u6CF5mPP56vSiqsnkEprlSoQ7Hwx/Vw6N5s6fEAYU/
uhbuIZLe6W9EuF74vds2qz/ru5Dx1z9QdQgBtRwi1VrlgXk9uyam/pSIMLlwJ+FBST+nEi4IPFEs
eSlHOD69a0tOG/HMi16B9QIe0FB/SoEIuIN0ESWGpZEvUgCyHmlieY/i9v16dbFQQ0Xpnlv+g+d8
y8MkDc2Mkyfhtf0tFc6oAT6J45r++oZYxzTFNvjxGTpsiY7rFDdz9Hlpp+raAOwCHAYRQ54mqNAB
ubVEQQs9NeKVCbMR6naUaBV9u2y4CcoRclugI9+GrxSFygzoEiXXQuA4PBErS/ePlTtBjYtzQAsV
oxYtdhJdniWIou8WHZSYFdtbxZB8ccR3DwuYbVHWxTBv8nNBpE4lSr4oHgVn0XDj0i89qHIzov6z
V/9eRJUeGXaPXmIRNB+hA4i6588/iRMjPD5g6c+aAr8OUSZVr9g8cUNtuXcvSB/ds9nOKL2FN9ca
5HY09zyeFPvGKs2Xuqpt2mnWRALpnAiP1SNp8ZTbtEbx2l9cJIoOLPZP6AQLtX/DWRy48bqYaOnm
g7LFe8UW0gJRDy+9j14il+nOZPdclGBcrxAgKNN0u8UAtZN/ejcoSGy+mATsiiUtRp21IqHbhy5i
WbvtSTDLiAy+fP6Fo2bwsMUZDn6kenI51q6+Gd/TH9Hl6Mv7HA4wyev0g70WnBs8mrJghfMidjB8
XsBZETS4lJLaL9oWWVoNM3JYYMydrF+IjQPzKAjhTRSjucJPftiBaxrbQ8Yao+n4UWEype6dCw21
l7EuBYkt28vJlC9V4Kde04bBViTPKZTHizfzy2AQUMuyaKvO9y7kgNLv/zKRwytnUVwHl/sSVyVx
MdPi4F8VIaRXQn+EZX4WGWRWxBgroOxcGhPeUiNEEnVY6WBZLybERlSI7p+Sg9zCdVz2VWENE1XM
CL9qKChoTAbDJ8dVBxmmYrw/hZ61dKZtkd66SJnrjoxlijadzHLGm4S3KnEF+Nf4TlKJMk/3UidG
heb5UfExji3EUQnm9BLFB+uSuSraQ7xpW9/ZWGj8QU9Bkh406/S6BMrZ9mCpOGRytTO7pCNEKnDl
qr15eFXew0PSJNkHE44bvcePqxGMHfJDK5NHXJnHe9+swF4erlDuJ0ejiBpLfJi5zdJh+PJ48uYF
WJz4w3qpwkVtRs2oLcbbrzCKjRyMV89a02gf1hFqnGkTLVCViUtOd93G+IcLj8Ewh0tTSQIaiTJ5
EctvqxTvp2soFr39l5qU2SAQ6j2g2UOJ6+h355opCOC0OQ9RlLAkQMr1aBy5TKkZHrSbDUDkOf9p
qN9vkNQ+IjdZLL7pKTmL7i+FfmqlvMLx2HfSU5PqgMAr0EFv4D3uXIUWcGFrM9RXMuT2kMkalM1W
XTg1t2k7K7PRfBSznqsdwslW83MorW0zFaX9S0qI9anXksuvW5tEGNLDL4dkdv7f0rlpJzigSn06
mCCkStOlUPnxcm9cKrqTSrr8IKamM14S8UNuYqpXUtkVk2+T7HDI+b01cvvvJ46cJCVGON0jVsNi
i5+jSIAFeMo2G7WdBBZNH1IkHJdGfxO6IQ2vwD/o++20Fpnh7H0c6KPgf9mbYnBLbfVnhz06W9CZ
Tgb3hbK4YTOOmNDQABzODvh/pkVYxPC0u0NNTU+1RWqbXjuqZSUvkqfjhL6ufHynKa89tf3gf9Te
LnV1zvCpInvAPelVLkir81eLyMvCoY3vsHC6zc+jsXF0xxNU0Ll5bbvKhpQ0J344GAi23hC1aEoo
w19EJ0F4Oq2zIvp3Hm5IzQYGhWwHXEXwxbQ6rHO8lS+xHFAHhIgRFU00PNG35NBp912IIwZ2d8/w
jAWaQiiWKn0/BX5vwVYflYHr53MtAmqs5L700q4MJjgIALFk7KyW1iDympqaJIQ7lj892oje5HWT
gmG2oV6qiQNX5EymnC0Gbz8NU01v++p7Q26lJJxfvv/P4StN+OzxcO8h6VI52eiAz+gRyFvMhQ9P
7l2c1/ja3B8uD9eKXrQORqZMIr6AavUfTYjEcjaNaw5QsSBth9FnSV1sL0DyT9AJAcVdaxa0Y2pE
SoyB8083IRnhp4kzbcrjFBLbV9SeL/NXqNwum/GYvetWTvtn6W94dO9ssF433MkGQmaHgHckimpZ
DvWI8oVQjP7LIXhA/9zj1pMoXo7rG88DdGQuciF1e7/iLTBL09MZwkFqfm9xX9IEOPei0JdzownL
Gd0kdFcS8W0TdA9zbb24zQ5WRkBJwnKo6Gmy/P0PG4nX/G9+6U5/s1bOw1iReSC8BJX6cBSumK6z
9+yrdTmvDxbIp8OiG+WSwAW9ewgFlMLLAM7tZMQ8ZMjyj+YuRaIhIYlKKxEVsIJpAQt9207YMo6b
LnxZ+i0U4U0YTwSAxetKlCkucECukAmsUwxMOQpFyB81R8vTPCJoIPqnLS8Ok0mwDi2rJdToYkuE
R15pwlEdPTdR2pBBEH8lQP7lELO+MaoCVwVpaL3qWSGiYgJFqv0gFdUCwayX24oUjhnszz68TSkb
Qtgux5o/NEc5JXkKbJg31pQKFucFg7tzj8iWQKHtHnuNGuyDAoKylO0nWicwXgmcmeCU5LqKdrIw
/EpPWCitfSYWezFy9Y5efKhdJ7Zfr0katAMx5XTMPYZe939gIFoNV1ofbke/qwaOulDNoE+ckjq2
ytUJjWHZJ4P+d552duH9pXtbV251wlc8nQ0qJzqAsQH1rT7N3WCjq8i0BPwbL4uYntHFoS73i89l
xBiuBN7Pyx61shctdGBGBuHGx7/d7HBU7omyerE51mv5brsGGGeH3SEhCg9M6VqS7Xl3KAaibYRb
yiU8gS25gWu4pRvBg66i5j1EJ4/lfgvA/a07b7BnTDT++QlF7KfP/1NxgZcqL5pYo3kCVL/79aKj
0QInu+Ncq9StSYEgHGj7oAUp3dfKVZLUAw9iVmjHad2EpMIVI5vyI4tHHIPfy+3cUphpXzwA9Htd
HfZE65Dt9ymHz/fgvE51deXNdeDJcXJQGQu0gBXx4UDTg3v1d6TUS55eLS8GHXoDoYxnSvausnAw
buGsS0fXJ/ES0tldfQa0TAoYNWK6tBkG3TuGPP8aAClTcMiWkkoaVwweRKzOdFug4EoI1c3WBCfg
hVzwFpC8hyuiMpLoRIT6vwh9u0FaYG5JxZKp1/CDXXMRUEV2UQJN+kQTonRT2bfLp/AyTNgZwxbe
ked8kxmPkkmRT3lZMcsOHlYlnusv8w5PvCy2Sxdgtq8Egya3Vq13+X2kpxpZrs2Luo51bVD4cHr0
BadSsN0ZXFkwbps3Qxxl3Z5QbgpvQzkoWl6lubAopCwKsNw2SRm3y4DZxA1DJOi5ta2z6WS6vUqa
YK6X3wWWD7m4t5tIGmiB1/GcWm7AUPHdYBDUK5qCG41jwwaLSjIFX88AFziKjaL9ln/CKgWB+G0d
TtlYyiS1zXOm6E//woLdwSh1+JAlT9CMhrK6/KJ9vWcQsoXkeTmG3vPUFdv3FqWRY8xcekK1VzBk
MyhrKlDcMD4czsqd4giinlkIb6d0C3pHplwEDLARZ4F4PQAqSxauUc2foUKAqWI8pEKPFnAwjsqK
NmB6Ejx9cNz5rnVCwslyBTJOVrVB55MZAhZb5Dvx3GGCee4qCByleYRTbi1vC9voTmcrG9xG8ZuU
fKOKVNyvBFigluNuSzUEMTUJwVJ/iOVmyXZr3lREarXrFbDELmzIhZ5kpvYzNRs64xS/NJ3IwzQl
nemcuw1l7K/+YuQz9AjuTFthPb3uptwf21f3Lvg+EIhM3T7eMS4jTVVE7m9EwqCUM3pYn+aMKxKy
0qw9yxkjBxIru5GS4s9ebysM0I3ePt7IurqRaLN21am0FzAMK/39L85lr8OA6V0L1az6+mHikae2
1hdRNFd5sQ7hQMdrIT6ijIdGjBlxB8+2lUqT7h4xqGw0lAQ+YwqoijVQ4GJ7kNXu2LRzmcmuzFEo
F3edHh15RHjvy3xHfT/D+Wr5gs3uVQanyNBDSJTd7saTcoAzc9wBAL9lbS22H6F8MfQdy8m9j9Mg
Dwx/SuvlLhONvvJdfnxJfSM3yO/TTv5Oh6dSdvzxi0kzH75hZMOxDxPtoI+7duPHIkSQ3ZheBPQs
CHA4vGcRXEbG/7ovs9o2jSNKW9Bl8M8jDwhen7xUIZqh1vcfOa1plcrAneve8Q2sMHvxMZcGgpys
rUDga7PPwoBNED/miGrFXSmpR91prSoB+GIjCXgVbli/Y0p05G0RiqjzgYWtVN5S7Dzqb5ggpVLu
hcfC51VqODeOCPyfWsm3sBTiLWfevfnwlgbK7cTf5+2TUYv5Y6D89smfKw3q6NKWisE9QQwNLrNx
n21Ry6XYnkMxwPr0HE54zZkzwSR665MxyOz51OKmsu1CwFjcQRyCw6Y5u0XZCTjNY1mPX4oRwg7N
ccZJzghJskSyhVxNGVDdyMjUXdESisfqyHxa6XfP3+NSDNIWTA8MhTQ5R8/elqx5T7Vmj3Jvpp2m
DX0s7ojbS0klXgmiZVpCCuND++sVQ74Sy03q+O1abBQ9Vk+VD1j/OKwRYRby49KFxQevsMN7TkQ4
ht4i6fcQM6nJTlz8+vaqxlNBebnSnufgeSKScgnUxi8qrhBl2fLmKLfYvgzL/gV5bK5oUx5JK4/I
+pKgpU7Be9fl7VUUfwPBT7KXlVWeYCHyxg96hy17tnZkxFEBgdIc8tg7oR22EJ8lLabBx+AwayGz
TegTPLOgRZOWBozjchW0u0D0yL9KYhzpLHzofknVqYsZP/LiB8PIg8h3uzJcr9XwJn+ReWZIY76d
PU6vL/sCDH7S75Vlu0lrirDh1FHuvMFCyGBoEEjmK5U7uvVN1+i17nycaj4ou6JoDLk1f8OoDk/L
FtkcxiwaaLZJH1/p94O0fTyUHsN9TRHnfDuyJX6qcfJoRumM10255jyr78NmebrSMX5nhsL9SuzK
faArkUpyKpU6FSFk2OvSGlsigqQRi54qR5fkLjZBqY8HRHt8LgwzqMuZFuk5bvw+cIdjHuugWP5k
raNnSZiYDNgnkA090sQKcjHyGDoZAWNKWYg8wf78qeKvGL/TXdBcU5ZveBGb8wSwHGtFx+ZWegSR
utp4XKB30bXQBEU4Bvu22FMqFD8+zVGMnVYJ07UHkOXntA36NaztDWPWIo/142r8+e1qUZB5M8Ma
ARcZ85gimAz5geSEtfB5/kVTDh4eTViYkhlzdLNzqlGF7530HrtF73n+tCdiP1upMRUHaP385874
wmdfPLFLLfZ54Cgsx0wepcfda1t9MNI4KDHXITkiMLJ1z2ZEwEzG2AcYiKWopzH/OyJ+HTQEgZLw
uI8tHFjFdx6SIgFnNCJDQZIckGGJJayQ934uYCWktKjwhLANDkhkoeESfY6YMxRF3hTM19MP9CKJ
hZKkMiiavuX1IbSecbIM2fijSc2NimUTk2MOvB0BQYoSsx/AeXTGOKGdrtW0NdRGrv9SIVGbnnGp
FdfNzvEpamr0yDDf9t0SvOasQBtfWZsRyppaL4OjmyQ0qi8+iQTTd81kA8gFn9EJfpruG/bR5sus
XdophN6fGLJpro2O6bmGx9LzFPJAidD34bjtH+f9GQnWzoirZElvcM6mBlUROhGFh8BIJAy6sORW
BosZxaQQPEieRDDgG0Gjz7neKpsW+s9yPXZLxltR3DjWQMEk21WRm56njoVYNX6sQKq1DT6CphJV
InaTL1b/6NJphvp+2HHOlLgueJoX8DjQg280j8ybvkQLFG7IWrUADvP0TXVpnH6BPJOqCEgi7gtT
psiMNtG+Q+Xor9wdtq/ur+VEdiqp79p46i3/GRyt6jOMXOjAUIwhBMITbeEC87CssBvh5Mqnfu0J
klgfn/6Zn5mx7WWO0hKW5aGFZFKav+kkz2AmcKVV1M9gmOSmCh7FlW5bjLQFfnplaPKVsGmFlYFu
VpBGuCHoF4tC+tEuFI7uLjDe9rcRKaEk/69HHNS1S0Tuyta1FucQ0eHzJom+UmzvVgWMJ7pMl2a0
CSXCyF8SLkLH249yte3ZF/1UTk/DFUbqPzuwhn1Vxu2SrGlYSvG5+YX8Ttb+fWGcVHDJqnxF+oMZ
aGQHbTegH2wac9DjZyBmzjY15dUf6j6Q3PKM3ipAPBnAdaZU7trneGKpP20S3H0wTRIrof7z81/O
9Yx6KgUuSqXI7eo9vCi/kfsfyTmkBbY/HBoELIxJA/STSPXQYx84187yBmejmQ7HsC1JI23g87/K
4MNFTtb9oYrA/7qqNrwhLlDmfm78PBFAmZe5RfkuYsYXExyBUBmg7vcfZKtrPkvBrZz3uMoklxra
ksqUwODs2CRerLsiHaQEeeYFpkmbv8Wml72pIT3wh46p7sSoJcKrH/hrTh08MANQ0d2gXatkuiC0
hecD0+jLUB/0bMFK96ApKCYdp59tpU0gBR8ers5dT785/4QEYyBqIGIfWVcCBzosEMjORK23x5er
xXG8EvP4ZLSRe/E4UR0gLLMu0vTw1dv4RRSPaZuDBi0vJ8IFecn9qSLL7Dndo/ZV5aFs7jE5h8Q6
dukDXEpQMUbIxZRQzwmf2IbozILu+FXBbdqskGRIAQR81LgwGj4xNQCz6EPNOWUfe9GAX4LTNdS4
dA4ert9Avv2IXY25Z+Y64pNNdN9KV5loMuo/gaTh/TfkjH8Ywl/Mc0CfQohFl8inv2G80uOTaex6
PHktW306UoiOyDGTgDOsuIAFX7eNzbidF4z/xdyyI+ziI0HsmxSpyvH/zKrtJQL7b5gbf02Z8g1b
DuorRRZc9nGZyB4t0ezrr4igpBrTS2dz63b9zSXHBAMEgCSfr/QQVLzUTfR8OFI0XO25Hd2Vk7XC
Zl3OHCZhz6NsmdKtnBHLjS25nfs496lzEkQqcG9MZz9SUHIQ3jUXdcJ08zwqWZ88t47G8SaXTFeY
y/5sa1tyXqHus7DrOzXdv0DSLjGLdJpHryTXNLCkVfFv7paZ3XBk++29+TAO4c9JEAtCTUZw7gLN
oXvkjW3fYhKGaz4erWdtd2lkcu7GkRcKLf7G/plKtlaegda9osB50dGz4t9cOaWI2Vei44WuYfzd
aAi5kVZhe/aNTpFIZT0Tb3Rh4tgwBw6Cpa1RxOrX/6TWzC0VZJks3VlhAJciJEudX7pRTb/DWMJU
9+C/UDvjRzfxf2Vi/Di4ULGxpLFJk2aqKHlJqDitv50R7S5+T6cDWamtIe93SPeafS1frdtAgepy
OJgFg3hilnR6bKZL/OIgXdDsVdb6Vh0tTmL4VSCpdYzhLOFM/+sAFIoQ7ozJzru8DFLG9eEX7b2L
7R0qRMjrXSH5JdCYcGeoFZ4k2aA3m2g5f/REsm3a48/EmM4EZyvZVV8Dh0z9hgaZdlaDaFgQIB0d
UgWuywhFdU/EGOebJ8rPGGHEamYVi+VaSKERMyK7Ib/HKazLxya3Atqcwp56/lDxlHS5Zl7FwZcL
EXVZTh4G4CCa3VZlay7l20lRbaJ+q/eDYrZxvrjQK4LNo/0XrQ3ucPUoZK+X/ZI01LWQjR65bZtm
NIfBZlKcXtp38xCpa+hmO+y6mZ2kugme3beml8jSrv+jaZZzexZLeiI7mOzZBblw/18EaOQND4bo
dWGmDWx9jswBsfKvA6AqpGDcDFdmaIIl015YDV8s4EkAHfH3iXBlPfZ9Vya1rDHn/AqMyJGn6IM6
X0upbA+I0bv1g+EhEyZp+4Rv2vbsZoS/Q84kFAUg83x/wYTkk8Z952ZJXGh3951k5dGEsUDMYJEV
6YQDttC8zESLx3oSKUWTrOifYt831lvaGxbtDBK80jnTY9bcAonJJsPbO4QeRTKPh6kNu/mYbHye
Cd5NPdgJ2WLkblz4bxzLG7v+UyYVMOrkDCkG9ATWVz3G+BSUPiXFeEF9RTBQwiNkNLpwT1pqw2bh
ghFqnjgkWl/SpAwxQLeVFSADm7F408cw+/eahIBu7QYTZaxPq4wk9IrOyq11U2RRJRn0MMGmI2A3
xl86Lh/wNOUQ4sfORPQlfcFbDXWFcWxuCUBL8/kwVnK0xY0fcu0u/ThQxi2QkhUnliUDFSzbBw/N
8kFbmnG2GjCd6XT7y9avZJcJuWN1zjGyqE5Zc6XnDSIXqm2i6FQVo4xkfFs24/RLZ6a8zc77jeof
Io26yKPfet/UYX4vaY486tVOzoA3IJI6WqhkBnb1w23BeN/0vPpfcbE6dSGUSou3v95JFKM3QI1s
k/v71yhNuoH/02RNo8TkVVR2TZN3KUD/aC77VDUgyDTcrQg640VjcofIJDpK0z4yAgK0zDX0/y4o
2yeiBgO7h4jDHlgPYeYROi2oPDsyAINIARJQljwkc7cnlVQi+qAI5t0CI/mdIFogSMUQCNv2UjWG
szo1gg0u6rqekX8GJimnwpNOjtWtHczLTHb6hISGD90ViY0UDF6+6SbljxXY9hG7cYKzXSmZ91DK
Nd86Vf7aBowfVoUbKct188eze9Y7JgEj8S4/O+Bz8Ju+dUZaizTZFX6oqkyvuwCRtJmRqiyShZAU
GQjCT4Zmx1Y78NZ3dHyoUbiNFC4x2q64x4mjCNxhzQ8mM/m3b70cuzSHWnwAnXbI7QwsFohR2YsX
yBmmt/D9OtpmoOiD9TkS6PQzUlDmUcAg1FA/4+/6sMz2mNRgAn8dzLMZzEdnPIUhSNZJle3ZN/H1
Ighk65lZSZiuKk00KyKTsLnsSX243fahmGj7dSJj5GeKKj7sVd2P/hY/4xt7R7oX+77aYkMur3bX
niLPdPA9wkYApxmHq71CqG6Hpg29ZYYKurGdfTg9zFAK1Dy9TZAIs/Gw+HNXVQSOqgiftV2tySSu
1Szdia96HMOfZYLpHArcOXju/5VfpJzBprG6dD/dZrtq/d2fG1j8+uHvvXxiAiHnKNxQtGUUMLPI
FHIXAxTB3cMVlhFZ7fUYabkEUTm+rgG/tFt9hN9MF5UKrFaBchkI6zibSIXyowvLknWOt9XsAprW
NM5gKYtiR3lgKpVIdENn2EN67ZrlAHwwxJSOXzeH77Qf82rAHQuxXVitvwcUousnB5Sag/OSOS05
9dGBhLyETk/g150J33TVj7r25ay6sxiCKWsUspKkoxREdFyi3Lv9dns68SoFgwzDYgIQ0OVq6lL3
+xs2EJtHYCU9Wnwhji4/M+mgmxY9uCGTsGXgj+BKxXRvitbLNki8a4ndLlyNAoPLEvY0JkBBt9FD
I40yv7RsUfJVT2X40ZRwWfu51zFmzv1lamiT9gO7aR21zOessDKNvKC+FmgRpq3/gV51UTefLhxz
F94385dSJwhrst8QQifRi+Xj1+IOVOu2Z8jx25LctFjX1f8BOXeRupjxSNNYVWgkqtSeCeajpjy2
QgqB/ydfh4IvJIMPKfMj3vWlG8Y3q1xj86oaMxKV4kXosbptMHFDKtywSFCvd99NL6EMVNVLomN5
z/4AXrZ+LZPjuJL3fm5EC6rKB45LAB1GcMz8fvSNtzG0Nhak7nhXdAMO8F0SsuIt6d0F6mcE/5cU
RNVdpHXoEn8Asub37SRE/VPFfzxz4hzQ3DxuCDKer2vX8/RoKY7qc0HgxwTXJkC7ihWkPp1RFjNc
7+YIfwh0ciie4OskKNhrkOVhwBLAc1/pb4oIRRMnueKHW4pRSz6SvNkkpt5fzEGwH4l3N6Y+fD8a
JK3/v79D2Z/OSrWjNj005YvjvRo4BobMNF22VmDrTZzlqYP0pVFWBUFIDeBw5BmMDJkJLSm+VSts
A5P2tQedYi2e4Ct51NyYlyWiCOSDKXlUFBu0BzxE1hlF+C2/rVFKq75YyFw1o9LMrqfLSQS5laFO
q6hu4kg/brw43OqQT+nUPNWB6GErjmQb2wItQFAZVe7HFgt4mhUrzSFARSbIr83pSQwQvoPxyIXD
zSto1Fx0BeKranv2ea44KTouRo778j38MDmqLOCanqbHaOCizfyDVOH3EQGzFK0wg37P+8+b8LeD
uuy0JtohwopR+2J2R7y4eKPv9uGI+Fqc3MXGIKP03FqemAHsUAgKAes2ZnX72yvtK/i327XE4if4
3PJ8PVlnf3+AlS3TrN2VoXLdH6NJMAV6bRch+j1f/GGZzH8t28+7iN03/HTe6vy260Loy8m3V0vd
T6Sz8ryzA/3iFwnQf7ONJyrNmKX15h0Ni5X6bvLsiZUXTwoE9KYkAluG2BawXN5RCTkW7Y1Ed8kG
Uxfro6yFw26H3EHilWr7okARi8WlbL7Yzu6Ej8WWVTXgiwQ82YCq8LeB6Rn+l4gUfmfn99yZY95t
bJsebXPpg2acD9CQF82y3SIPfYOtJA8ZQlf+Yn/E61KICUA2I01ej2RPWDJpRn68l2PaNm82iqMf
DjtRJWZftUmOtBY6JP7GA1wvkGQheFsBMtr37Ryi8pdELP+7ipGkhm48hidPqWbbQDsP1HmRc45m
TeweMn2zz66i92/26B9bGyuUoszmZWPPhu2xP7ruSzM7KXC9HEJHr6UloHzdvUP08B2friwlIz8/
/OxktxXz4638pBYuPIDsWcEdpN0JDh9Iu+9x4OpLTXUzT022W6UNi3NDW33Sl3clZZbSAWrP3T88
RxREgB9yv6VeUsQxy5cnUly+Vx8IunHtH3MqqaNVtQHRO6VULnDT/svsY1V0zLL9tfA5iU3NDpxJ
e420fMN9eu7ylBj3pgqoON+uqYgdnx69cODsxtIrREKeGu6dV0eNd4zVe1zUvjU+pWTeE51To0Mn
nCm/pE5geWaK5v5e0PD+Je6IxCXA9zSSK6R/AwhOc4umldJoAYGjjvsiW0jYlDoldXQ6WmiwP0xh
3umIb0V/cXrENi8nfhEHK1IC4H+EkwJmBP3+km3+NfPw2MLcUrmYCpQ50FA4SzZOn2lEIl91rzYL
ATMaVZ8RvJWsqstaDamr0pbD6OS3iYJDAbPh8XfllCIC75CZg+o8R4+QLKzgrW6MpAqtBrLSSzwY
czOyPaJBR87MoNOr5X5FCiEuDsi1MT2Uj/YsyjVI8+KeX24gIX3o8aHouy8qETcxtGWfM8Z3zB1R
eZZTVTwrjWSJA3ZUSaC5FrqAOYQi3ZVI2fvmAA7tvqGieSzptJpnqn1c77v8A7dVfBjCUHZbn0F7
h+Y1rCI7G1DaaEfH04nmwW+q6YcgYHPgd0r8SiqmGw+xGvctMc/+amrbzSmhASQKPvXW+US17qLH
q19/AZaqq9HybDboYiB6t8bsWeGfhRHLuE6l9mzGa23FZvoJeBvEDjbi1qdKm1f0buo1MgIFFLFJ
WaOiKvxo6f4KiiijlghuBj5z9WL70GAcN5VD9U2TnVslaPUnBt25JOQJfJf17M7hn+v4Apd/kCes
Tomah5rx2buA+aZ7KjIGCeg3XS51cY27YnBK0sFa3Y5X1z7ME+41/a2QYPAvB/pcU6R8I/HW0JqV
1AgH7qUOdHR4mHVnk+q3GmHgHlAtZOkOtjlvjsVLyqAP6hzSCrQNxyd6vfdq+CrG82N1DOgHenF3
ZhyKZUr7AgIzlUfoZwZacduogXh1w4QKoF/AsjcCZm/Siie2Mh2bqnQAKUn77ch81rvKZ+wNyomv
MPkb33JZQKcDqHf69dH3BH4pwWtgSqcEIjA7CkrkpErUhZhn4ctEr1IMtb5HcpFihhSauCXlLK5f
voKS9vwyCmso67GixF+CaWHrFyyilMNtlJe+IKvs9Mx/oIoaDAV6ZFPorZ98u1xprYqPuwH40Fi4
+gDSYHqYuTpr8ctK6J0OBUwfxlH2H+BWuGXu+UtuIq71k8l4sKfyRJChfsgPvc7H3f3gjCrsxjyn
KpsU69qBleC00eKDkhmYKi/6SBzEPHs51RvNU0DtV2qX43OB1aWQ+vvaKKUB++QtRVmjrra/6RNb
VYuLfOI9kVONapRHzHPvRgxxZQmNGxm1uQwi7RvC5cAWygRbVys6TOxjGj1PAq6ZtCRPQMaHmbhU
CMSLtVwfUDuabwXG2DzriuHZfTLqGCUsld32ti2wE+V6LEDpHlGlt+EE8bb6hYi8uEIZKUtqhe6V
CSUqEGdN6poAToOFbYZCayihiWbZSUoBkLFTRm8s/j0I7d+62ay2AjQz6RShMVINNiWThIXQw3+b
O10mParsTLAzuzuLVEKOeeieofSU9CEyCq1bsMGVrh12t3GFE04Xwy1p/7AxUSJrabAxvvuNO7ao
rrfvYd2BN/kQRkEN/mokSq2e6ips9EG4gGWj6IlEWKdH02lOEt6o/YJ21l+I1613kPqA0drl+HiM
daIzJsL0ULBoxaDLoir7aUu8uwhXuAhoqx9l3okFKFFQxsOMxh3C8J7KlFyliYtQcehsYn8G494T
VfrzN5+CbkluEygfIkBEyD71rF2OXPQZQk6rJEFQ5O2zpDXke+DMjOebITlHGqJpVaA75xjkcHpD
pt7Z1l3HYrrtga9yL80TLaPrs6J8DY/UJyyf0KFvnmP4o313QpJKTni7iAXKf0kRmTj6iBmW3MV+
wqagEJM57rsTmTO1RGxCsR7Sk74pE686MQ9RCNX3qN54ImPPRzR6gdoLxYQkjTfvzz7oedIiF/uf
5DJh/J0vdQ6c2qtEkD70e5N87p0Oa64omTvvOvyAt+jzHAmso3x+e1o6mBFoFRHhtv2bvYw7CEfw
ucO5Zg4PGXBUkLt2GZMFBw6o0L/wp59C1N8HHRJoAliIL/yYm38N1K3gWF+Op9gBMcyveScKA1WQ
H53YDb8LQeNPARCsePoXADyQwXMSOisa9qnL7y7nLh2/3iW61eGRT46EOnPa9ZSp8ajyYFXKWfES
i1Gw2mWOtNv+cLBslNeLE1smhhpGrZFP6AsK+Q1CgJSWW8Pn10BLLMscZpWCVJwnqdU4yCn5uNNg
ET9TCykAiLFdtSwBvZ3l/MX4Y4xAro0ipx9F+jfsWnnW2K2a0H1ESxcwBWeIrLQWS+CC0dLK1vT2
9TS5l4JQFRGsimi1RI2E3hJVfXjmq5Z4olnKn2wQyWx83ewCaruubLGiLbjkr8EGvckBdkGLbGaz
TIdUrRN5WI/cCn+IzvqutOb43uHo+NHvj770zoSemDoL6IHBsY+Vs17u4FV8dxJSL1LZlcY8gZXP
U59yA53oFb1q1z1F//T6uaVhZMYQa0H0kmXnXuXS7L6UdVvcANg6mZTYXKuRNOfGQU8JZB+UnjL5
6xQFvxz3TN3gcOt6xW+xJpRjehC8Tt0+YdcgUpFyal0rYXZF9fI+oWfhGQHsrCDM+l/IhOu1OaFH
OHF+zbZjWf/0TfOWAltE4zB1ukWb8Yj1Knk4Y7sVYSMUNQ1FGI8QPeC3GJFeHKnkwQpMeyLjCnq7
lyP+mknpiq02UEV/nzgq1mJDS/ZNUwgJO1ilq49hMKTNMnRP3FPlf8CR6+Fphwjt4AQ9laR6ksmq
N0j+LJV0jkGm8Om9o6RllfJIK5Vbsl18NExtd6nJP2dDoON16phgijnRdnwhSC66CkYMBh2cpaSc
DN1KE08wg/kKPVZdNGWOYyWyTs0/AAd+qh1Ho0vNflzm5KWm5I4ZSwruwLgwqJ46IYcXHDY/G7YG
wowL9RkwFWBlqRbTksqCi0+sbG8F4YRpvQVxIEsxgECp6neJA3LBEy59rXZiJ0iB79E2EooD3YUf
fhvkywwI8iVM1hAC5UevNmPHJoMX/R391iiSq9dIvF1gu+GZnS7vZSFdZUZXQEgOeNtbdvvz7TTd
wPB3EhUIBaLA+pkuKz88AP4mgd6bqqNATjlYE31Acj2XFIpaSVFLU2Z+AOixcfcD18fb1Ige37Hu
pMPIhA6qRec3un7HZs85g9U5kRnVZgkUa++E/ePaOxdR6x1k3mUH24NdMDwcT8HdX1q6OAwNBb1B
eS1xb6gviuYaaSlIveBh1LVWhOwC7G7EuOnlZAO8vti5qBTlLTztfhJg4PcagT/ot605yncMqIVd
PMudNKaca3R3e5Z1YNuRepzS+2Tg+99YcfMlpfP2NcNPEigpbsnuf6RdjJe2wvmaw8iLZtXtl0Va
kH0R4HUtW36C8Oddk/E9KTuMBwrygNhguGxuKEMU4/wyHY6DOCu6J2/pDn4TMstzvg1SzfQkLerN
h08gIkBCJ99UokBAg6KIsIs2/P9AZSuvjNlhQgaS6wpYQf/JQ/mWyo7OXp+TxU2nKrYAyOQANhMs
l9+mLx36dFqyPrhi441rVjg5AANmnEjQ/cj1MGlzrGns8oWB7P7fiOIc0O18mHeMdID0QwHGg1xb
cPsCea/jurUP1hC8ecgY6SyHKGP62jkvBJHsxAIMz6XPv9limXMYJA69hRlRV/Pu8rZQ7Dk0hUdx
3POcJzbJoQnLmf+2n4gVtF1x0fG1IxIkUJOsrLO+Pwmx879HVs+JCwpgAtww8XBAiq7OZfuzL7xf
YxrOzCSaO+QEElS5vLAS/75IZSbdayhmPZC2lYLEgYsAhQjnBfUfREhM58kjTjrFinm3bCVGkJy8
CPKjQb20VIAGAjUyEsV5xFCE1PJDROs8h+GOAeTUOwsBFafyDH/eXGzoqYNvRyL5ipK69RgMm28E
MOkCuYTFrCG9IstDUt+/LpPeYzBw04ETXQuYYuYQJ2hQ676sicAZ59tqcrK3NEe09opjZVSJ6RWf
3gMBIXV5h7wtvCndJTKqQKUpOTUxFt8T4wg6GMhpt3z14JhHOkJoHF/qKgQoY9NGb6L60LxOuj+W
FgzWrz5i5J5DACFnFsJRohfk8RxVCjoKcEJBAMDh+uii8pFHFJqfZKn61zdGTCJOCz3Qok3grwfd
J6+7k5PYdZpk783ZkoBTHwMCsUgwNji8BXSALjpjBduFD/YJECRul9WucbtFzA2gkur+Z6i/gbPq
Ey9V8gb2YzbC8rzIzAjP9JftEIZJ43NJiqEfExLMjLE1OkaTEEvHxvgwnxVywrEU0qNjX5H7JN5S
YnYyUAqWpAMDb+w8t7kKzk67B794KyDJECT4ud2WUyU43jjJ8yfHaXzQRWK/QWEn9GPs6F6zLVPy
8eKG9iGWsHizozSLDjgXx83RZeotT6ZAQrjhJ5/QdIeq7Dix7FpvKnbECAX0RoRH9wqMqRn27Ym4
oXd+jY6PUb11Zk+XOr0/mcyYcBjYu+lEh9VCwDgs7nQz5iW6LwtU7J1s5lbP5uSa9SmBENKZeHvY
jeMIzV3lu4WAnVxUNTFSXso2JQ9pfufYM15i1wA5wNZr/pbcZYjwNWU75WzxWmG0e23FnqNuxgkV
8JH++7jChcKT2IUtaRsJqrFVm4UTrB1CkHRtiLYTt9VIV3lsgam6qaXtM9umoeZvc7expsfSTVx4
noIKQqAnJ4D5Vb4cQHBD9i2Lp2OkbWHJD4Jbp0BzeoaaOb0Qiw9VAL+IPQFIv4WFzJWSrczwesFe
5L6sxiAC6DaIaMRRj5GsTdcL3yqzxG4Ls41Fc/Q6qTuwv3VXfNnlDk98DAxZ6tjY6zQ/C6ptP8BS
aVXT5khUgcbXQBKQ6M5CzRLoalMaUNRcpmdECzBqp1FBhtiz1fafyzg2rJtRzRtQmGbD3/c9wkn1
Zq8c3obyAYoFvnmS3qvAClHGlXeAR+BQzBIOWfTiOL8le7w3zyI3aLu2dcAVYrRccBXNmmTGXJSU
dAzhTjPi//6aHquT/yTIFzy7WF52bIDEg+VjGekIo70ApqR9xN0+JkkxuYpjKib8VPMIyisXQlud
eweeu4gN2n46Fcc97XIgnW+j3btYW2PlkoOeqiN0DWpZ+nB2gpyYaBghMXcW3eWRbCZtUJX3x4tZ
RdjRe3RfJ8FJCAq4ZI4ZlarMBIURviUeu08vSBE02USgMWMqgdjkGI7lqImPv1pLnp2BAc2srClq
iuW2zYpAFc4hzwLTLuqSvlegNrZnhZFQdUIqL7E8guvr7thQUxq+FvtwX8swg39smoCH+v/97bBV
tcBJ2Cx45LK7WlcJEBUdrWzqKshuSPEdDao4QUha8pYwGxYY2M7a4XDhKTKgce3ZKowPafkxVbI3
Qryy8bS+wv3s8k6p5wn4xEEImbHTvaRtM8uaC1LPcomsGtvcsAkMZ7efz2kdGsDHYHE+zMPX1ynu
rTtrTZCO31Z8Ma0/W5udy7uF2WIdZVQkHygzB3sYsoYo0D+6PZ9J5P00R/ZK1CTxIyiMIPtQ0F3I
JCnRAz1Lw8kMH5MMoHPAZg66h4IF3FjoAe9aJQRGFEf31T7x6Aifg6mXOlbstqX9OviZ4TGwrUZc
BalEJwA1FoLHZJClzBJBw6K44g1EcsvgGMFWGYeDLSAA7+HjAEImn91mWoRoriWOUk7Phoi5Z3kz
62KTWGqtqMQdu5+L/mqX0KsI1IvG7myKhX+224Ed2g7DvLynFXlJ7tErMCvNxKc4b+8iBKkEjv3f
geFfJckrBq9jStx5Zkdmr4BOtjgj0hGX6XgiLU/HunWwfFLZZ9UI+Cv0iAm6+ytqOw5Zv2GBTpJa
q/dGBkwbtvavQ6SNcAQ6lXIEfJ6y7GXV2LnjzRAMLCkVt0qJ0fEE0fovNLAWN05RwI4w/UELtnWZ
BKv/NGtQDUJuczrfUB2Vgoq6vmuvPjZ/POt1RjNhRuEJiP9885aNi1rKoXm6BenLAkeS0YcFQS+v
MyQ1AUF1fy6rxMbgdaGa/tdKhnPLr0a8HihfIPugYjcS0YB6vTq5K3APncNnD85l1hSvS0I51eDL
kIeGcxwYGFTDkBIgVLEoF67W4NgNs1ehMOKKVG5pilPmWrWz8I6k6lStNNpj8xMdviolYJf6anG4
mnqHMBOPzPL2TcHSe+bZohrRy7cDCpSDdSr5uRB1HoWjjwlYRFlk6Ck54iELtv5doowpm2vJpODP
RXYCC3ywsKOJVxg4i2EQffTOxRgfK9FhIKiVOIz20RqDTwfMu8aL8QRxeGKFykSbtNCaeFcS61Gm
KstVIV8vfu5BkndF/0pQbRw7brhMO7KMgm2XPBPqeypbHl03xVlOXwDr8IJNKb5B6/0YvccK/vqV
+s22xN4wusUZ/FAUHZG9/NCoJkkCY9SB6u9/zuGJtTcM4OrSrmgv/U/ryU8FK1ingsHmHuRBo3cY
qkRWaTwOb8/67FvvMtXwSdhhOMMjgS0S0PCtZjfJUQIhk1idf7Q+Lx+t8upQ3MfFsOtS4KCb3uOo
VdiswkWQQ+GQWqyZfWY8oZhPgST4uya4PVfcr8zaxkb/rr2Vw24nWdgpcr/1FxmvEb9tDNyweecY
zZNDowgufoHxUIG8fxezjWAtvYh7UPacVbWPZw31ObxACEErix7gBv6Las1TI5qprpK+S2FY1rFw
WyDH5aJSsbK6wod+X//eg8PXtN4or16meBBuK8YdHGdYpCy6VbwAEpltGBCH+++Yr5e+xsgvBjxe
VsxF9jR2BaKCYlIFJgTrF7orKKN9s7ypaaIc4YWVsZ2AvEoR+SnGEztq18xoqK6ju9gU+Gp9fOQD
0FkfvZRZrAlaP/Des2mGEg22Qe/BbpWozhOm7pcv10bnuR4uy9KR7f24LjE16EKkCPN07BgFhdji
WVP2trlYdjwSNs2wTgWvQT6e8ySyDl742vO2yNlVMbIJtXwUTv1Q7qhwpIxBirvfYvBhuApdHZ0j
2NBmbEoj8V6OqBcWsOTMeiYM0UE1AC35mdfTkLI3r8KNOmQEoPHTI0l78jfX4RugcbDTbnFfZE3M
Rg1RNYQyimie7fKRYmPlyPBCkeRC0Y5nuZsa80viuXkVkXpTbA3vLk0p7v5XZtj60D7/z9Ey9dB7
skYZurNr1c/xCa0MwkFHaOdil4FjyhlTM1lXrMQJB1Ogco04gD307+MNiX5jHJM4my7XnowsqXat
EYbxRV0t2TxFTZRvgWZlpIZE5tRosgUuigL5cHJ02FbQcwY3Ty6AnebWy1Ok7dw7Q7jMbuuVBjxp
2kgA9AYWOAp0T78YNCChroHF20h4g0kWR2lbG1mrsC4emT5RZktRsuIah6bbL37d41pI0oUOuxMJ
HVN2L7u+xJpAer4FO7K+TUOHbPVUn7dPG3v3mz/hdZHPdlyoxjh1F5ooreNusAYf6HYjQlNJuM2+
E+YFJUMCahntQ+zXeWBvB0ceAqKae7xZ8OZd3M9EDLPytHKrm8yVaC8B1RVXBEN6duxGg1N3t1UU
ngCuNHhpZdd7yx1XolXgfTknxxBgZuJ/ORKQsvV6wKo1kZRJTSocg0zqrZyc5r/5R9de/0cB3fU3
9SVyxvN4SvjMuxesJEHqFvNZBI1eI+bW3L7IoT6gO4zyOpj65e9O4fqWsklG9F0a9I7VeDKidVqT
Y56M8t4cfS5c5PMBaARUTHw/qDjgGZB4nTf3MbU6lo4AtEdipdjjNlTiS9dMgCfLHbUQzpHTD76v
l7LtoLhrnay/b4++y+OhrHlA2snsnyfFMQh/OxRjYGR3Ne0no98EIvs2cUOPMWsEYo0qtHdeT3lq
ZELf+s/5DVqyW02xAgMW72ALiuK3kJi4pWN5Lo/kKb/H16iqdxXxpky+D18tvLwl92vAKfEsU4hN
qyeEDPRB2H7mZrcDWqWZ3chKbcP8cH4eeKIHyMh0G3hg7PnKA2Nw628GTvlnFK/sS9LaGizBq/Wm
yU01aw4b1D+Y8GD/EDgBYOW9xS/AYs9LWKX/eMxMVGAEilr8zBYIkQ5adBp1NlsJ2fsBrmtQblu7
zp56d2nhvxdxT6CuAorC3IJloFTihYxCTL32G207VYv69qVAaFg9JD7S8ZFuMJfm0K1TkKyQANZC
HNFj3N81yWta/D3Ja7U9kxFOQf+eDXf+ngsnXTNdxHgAFoAoqgk7nHVGr5yRfEzdbmiE+8e8zmLh
5WnrKd5FTg4adtb6Dihuk3Ph3v1e20If9OdYI47b/jjnk/nt+RNNiM4dw5QZ4IFmeZZ/3626IM0f
qL+iLsLDpnXlwKOugLYyZartft7446R4wy9ODNaozfujbK8Doly8wZsN8mmnPtfeZZMstOAPGsvA
X58k8Fwt9q9kQ+aRl70zhrUHPtJBk2N8Rg2k5dS2CIqhFZrD2kS6mivf6ptG59CJ45e2ZPRcWJI8
rXYj9bAvXK9OOotGEPByYxFwuT6MVGhc6EBXTnylhuB029Cdc5jaZ951MqXQ4690tbUhgMgkq2Y7
fqS6yUdC15LSe1rq1o3bXg9I+FVGPGCD6v2u/9BN1QIrBf5HE5V2W5V1JclDu+xKKu/yQCtqJPXh
qza+drSqwvo8gN286tAIpWMHTfe1+JzOH4usybi78sU/tCEgzTYOiQ1evzWEa3ukpX3X0jBY0WOv
Z2sZRnNSmJ02uCSK8rWj/21xqK778mNH6sbweuvTUAjU52E5ANnu6Tb4WrfrjbpX8TEYrCAxJvf2
ZA475SoMXz6UFUgkMsa1qR//PRewpV3xmb3mgA9wK2gXpIahPZmSoAdG4AjmAmvT6Q1dFVpoosYs
Pwc59Pifm3+0Q6cNUD4McotL4ZskWJiiwgm/1JeX7B1IJt2A9hNU0BQ2I8hcmPSBk6clMCpblzXY
F9HEbhWVQcoIbWkWdY1e+jRf0vNxnEPTaMOqr7s7HNAj2nZj3KXXFaUNlAy8R/xXdKmsr3/bggPZ
Gne3LJAzcmihQFv22yJ+ys4yBwEUrMbNp2HNXBMAo7psqrvXXPB5eObPFfep0pb/fKWElSIy/8k2
HZB1sDJOclVUcDwwI64yuAlNRCVitCeA08gZq1bJCs7gwL5/ozUFFtttyih/jlezRgtpBy7oXAEd
pJoRJjTyzzr6KkkbBK7y9diI4EkCfyfjCBiW4rMibZLVDGvA8k5tXz9on1y2eOjuFWftj2sfShMl
msmgtjeuMkXrtrpdRxyJ7jYd/B/QoRQFhegGzlP2Usec7wGQHpZbIgUl5sFyKd43/oGjeWrj7L5l
0YgHjDwGrZf9iQF2d5jWgTpense/bOO5iDyXL/C0rOqAdQCSLtEALALlcijP6hVJFlk9HLaXG9Xs
tRoWBlDf8IAfCq51QbrGOnVi1N5mfdLcaZi8tZHPlFyl5SXvYA8LSlYwTyygSg/gR5o9W2Y9/GeA
9aeV25ZktQ/wSweG6PX03U+zNnIRhbMu0NaCepDTvFrQYxCSnnHhpRy1YF8Ci8kl6XprI4rlRMhC
rz0gJiTI82XsGPEpP9kNHkhRnsuLeHKDDux46pMQ/YipGHx6eLiP48EVeKO4c/0HjmK/aSWIgNjw
5CNhY5sjqkeUnTWqo7fAAD3xEHrjAYXYUh+a2K4V17Y4HYIRakYABQZz8v13GNkZiLGnIB4mNZpK
OgFHVhtpg0OGaVll36TG1ibJALryJvM7VZ8gep3by3IWgzB/tm3/QfLLpycIwyT70Z5O66dDCI1O
XDg5ZedUTuRAcXSObBa0CuhXH5mcq3dbKNv+kZCAIKl+zcNJZWKwDkjvvYEL8Rw6InKB17EG6+eM
Zbj/LYItHMM2q/r9ownSUOm4eyy3VtqgYwTawnpYxJbTglSrzvL2AQTGPEGIZAm3oslw3kxhjdJ8
Lzmv5NsBzbYkUx2iESohvzn5uiO5i4XQ5QZMJuMxCcozKS9lK3PDmcdZjD+F56Cn56raqvvjF6P3
Qm+D/mwQoblUUIkK1nW1uu+BKVg0Z9DHUyhaYqGHCzBL0aJGa4BtTmK+uieWgDyNb+AzTV5ezyFx
HEcBVG4tYK6pakWqkUgrNpEO5NSqKSG0CdJK92HcmO8kB88Ex8b4nMFRjeZMp77kcWA6iFU71a+s
Wm6cU+Zj/pWd7DYTe1KMLrOHBrojXErR0GJyIkkgN3EdIYghQDh8EAouscJ4JpTqVHd8ahtnh6tX
+BceEaSdMAlRilwf+hsazlRExi2Kiyvmr0afqLs2sFq1XXqJZuiYBenWOJ+U9YxtLJeI7BYc77F6
mlA7Uo5NDC1wEtq7hPh4w0vp8vtxG+msmxxPZ3aXN7wrNjFktTgEQ+eOaUxrzwbZi1Y/s4VgwzI0
JsWSMc7EBNnOJ3+0S6NDQU+/AsX5HyCth0qRHhYFjtFjRLAnjWtHRaCjmEU+eSRME39rhGJWQhRP
C/s+zp8uC8RTgyissvVJNayfC9nLSVvlZ0SCCcUpVMuzMGfx2AIKAoP+qxVqjkIDQXZcoxM/d1hu
D8AQcZlp3fgZ+7cwrsJBLrvcewnLA6vOk8+guREhvEuwwZf/dzjVw/mR1LYnqwTGBcJ8YEWBbdze
3bgw3QvcAEW2YmG4Imw1rQ9PzTDY6uWN2LukYcAFFsIv3QfV12zYU1DbRrZcRz8AGEMpwjNkFfwA
Cw5Qu/rMhiH67aC99KkRYs8i+qYBYMLBP7SEbncxle7GOwYcDNHZl/d24VSJKdsBuBC4aGWSaN3R
6WNFDv/vbxyZp0524Zjh3tlP9j93+pLglo5TTCgEYsJhbMjyoeFxdqUogqOpyT1FryreDKTz6BJw
FAwfAQFNbSJ0KX+qpwX5ZzMZ74Miz6XHA5VAgudOMqcK7AOirGNtZ387qrJpQaSb+ohk+27M8pMb
+s+6vg84kqfC/BsSZwe9IRFAB/MU131KLhPuPuRijlcfNjzZsMM2CaPfgzz45Gh0mkCxWOiDeaBa
sisUV6uujZlaoYCK8afdW3f/3pl8LAFcFH7t3EmimF0M6/wMi1KcUA80NJ8Cyb14/P6RRWsUg3D+
8MlLvu7ApB4YCbbV8MgpSTq/yJxaPluZXYhEhfSrogGp1w+wZMmJnIY+taHvTedSh3qP177vcUfH
C3lONi+Z/ihIt0kRH67zMU2ukEotCJMwtqC2qSczzgELhlRJIvpytqevHKW5VucBWy2dFmBw9218
a8iSxPxPTl+ScptBlyJfzCWOJfg6dDyrW/tjdyB3wyYAVD6rM5Cc195tFUeKzbHuQ3Lug907u4ME
6J6xRVWpDIudSm97rNo5ca46cg5UYJadojIPwddE0f/YaxKtYa1O2LttSp8KnlEGgj76gwsEd8AV
D3Lv/cT2gfZRVo3HuDEtfscxiGxNTMXJZDPzRKJdtXtw3g4HSMYf9sF6Cqr845gEqOph+QA8EiKY
DE0vEmXQI3WWGBptkqEC0My9XiQzmPEEM4oQtvmNI9q90O+pfBzI40ueZuYt8K+ndHIdMFi4wnTs
xUvp7QVC//WrKQRuI0tuvPNsfDCTy1ITuvqCISYzpibOATY9wG61gRTFaPSctXqu9FQ5CMlRnMlU
NyJ8wpfNjXJkosURG3JLoF9gpSJ+Xw7rVkq8zD27M9juGgzRM09UcDPDrGDTvb7wyE84wS+xBw4t
biLlXUwczcKsxJgt+v8aBQ4/ZVJsEmk1OJW73Uf9qQB95K8gs1LHjV1idLDh1+0eIEd0wN2hevi0
/SFcIz+aHU63Yiqcn6NaYHaL+ml7wJIwjD3D7ijfKcdUsDe/K8dK5U5F+ItWQkMVywgvLOM+naa9
8XBJWLsXfWfSjl6bYV8j8Qe2IYt5Z+EjPiEjH/ycC1notCPaAd/iaXYhJqrrqYCdsZZ3p/N+6+Q2
+Bbdj2DKxg+cmI6kr353ACSml1xfrx3uA6EOleiTRtl1SZdK4TWpZsLaat3Gmhycd5Oafs2LXMyR
/s7gKjPn0l2PR+/Iq0n7tzh8yKpMaQF2diNSE4XflRaky8TUd9yqBriQvtMK/QjEhZpzitt2Za3n
BjXAkN4321KT2GLCtMd9O1yVarmcomBIA67qdNbh/A1V3gmAFjkwFsnjJD777WHMhFwMEH13UYo1
kWxxv5GMHiCvEQ3BloVRlsIE+po9KNIOpKplqINRPoJsqliGtSyzjlXs+C11zKwhaZ8rtHV7LCBN
CnJuEO8zOJvbbQPVLX1916WTXKplfQM0HoO0jStMPGLtyOwXPUvf6iZ7wcCN2tgUtcf0YuljMV4z
Z58LZTp5zidfpq62VMXtKMlHieHgIas0UJTK4sfBiuTzLz0pCu0PxzVkGiutLPHiIeYxYDR8/9fy
dlGP4ffhdwGFyNexfUw522sst9gqlC1j3sbBr8E+2/kuGlHDY8GsuyMbVrpcMwpDduOztYSJvo2x
ZmjfgtuNb6dwE0l8O9vsSeC47G9rLIIs3gO9zlO1HJjNn4lF9zJ5v35eInexrJF252I1oNaAvPjE
e46HRxJsGc25KXs4Dxd+98Atytyy6Im6NTfgk9fBgFk4Z/L0/9zM3xBSpsjpK2i8bsMlKtoPTQbx
1na4ne9oT1yo+lvrFPCFTqVDs5ZJgmIzgRjVYDE8XgU81RpNJKwJevqQ+vuwYnf4ufT+67y6/lyu
k7jar1zL5tDErOX65BWy4xpE/XrPkQRbeiYpLIhMmrvnl4LOD9PUCVSZZ4/22xguI0pwtTS9zHyu
AASe7nbCeHI2l4uQcTTSMgQROKZi5zYL3CTjQ84alOU2G0LOhNcwIsoucN9zVLRWV5NP/JydN18c
fI7wzLXgbLKTWtfv0Sa43Tptp6vnnMhfQX1UNLo3YiIZQq8HnTIqM75tIaUaokA5odz0SnxPe9RC
W58/8zvX9xcebppWz88iFwlaY84mBSx+bCEwQynJVEaoglqaN/1+2r+4aL1zXcLljysJug2msg5c
bkeSJCm9nL0bo//SnemqdDC+UYUzpsiebpevc5hv4Jkkh9D2kLe6LrtnQVKhOKP1M+e3+TBR4Zw/
0nUg5xysIJiquAKPo3kcr2FOXwf0dmu4UYLbQDLGHrDrGwmjm98k+THguYzXenyGV3a3TDiIWO8S
j3IO0qndSGbtPVMexSSaRJEhZ8QkuMPQMqSnJjHSuwXl8Vi5aeev6njsJgf+2TsEpJ5GGz6IFCv9
45cgVNYYX9bopfkR2ZteNeb6wCWgxMU7lhX1SmyKzTk1UwwNzd27i127ZZ2gGcWC6IcVi8KwqiMA
2kuAIUE4PzuAdlUQairkHsMkA9UjatCsd8LDzoSCPRNhKec3apd/GDGxFcy8sXHzrpCZI873zViC
+59shQrdfGHUPd4T3B9tNJCL27oFWLZ6fwxd6kmuTnIxLL7tZmL8Qejj6DeVbBrwPcmcByE1bvRB
i3gWPV+YOcEhVJRSPaVb0uhuESmQIpbCYEFSl9MKfd4dw0fwCJk/7tUAbnQbCRhba8ZXLxikEaC9
F4e2LZ2dQvjvlJ17qCdUrprNHY8rzoPWoA6gYPsCi3C88zjE8v3rvL7WMwaAypEyU8H06hVYp+Xh
/s6vSD5Xzrj7ToxfsI0Mx27S0Wn6pYedyWxgLGT8A5RtQisUENQZV4fFrO10tALAak8DLYtbPs+a
ikCcDlNo23FRoMUhIG2hckdRgR25pkasSLjJDmz/mP6EsJdMLtM7TeGxwPEuENdTCcKifeMn9tEf
eKeMOpkT0KmppJK6OTMDR4g2qN+sLKggRoD+7pZBpRYmGLqscfmDEbWAi+/KzofGtdrMUWxmIooX
4oW0VkSviyna1IHuSSF8gxc0ZAy8KLlH71wz2ZG1VkuV1n7yNA4Upy8H9eQEvAyaSVcNTkCR9/bU
3IdqaFYRST/ZtMqP+eQwxKjebT7jzQsEAjAel86GOk0zdnRe+7fkDB0W09o7gs2ob4gveodVAK6K
Fxp8DmQNTEiJpAOCw3QBdstPO2IRy7y2ZLOSzT3jDgcy/8JRbyXx0Ruv+i/WaWZcxE/fXJBMLOu/
+9R/HZaWlvo7lzqrbejR8OCcv+0Gc3bScMxbgx1o39wUcdUW6uUG48gyIlPfP9WgwaqEK9+BEVzj
vhVwKKyDCtE9+RUxtBfT6Nmsyww0hMHz5JxEz6mniQFO3qpqje75O+Y1DOvNNwzgtwisBYiBsoDC
v8hACaJh5cwAadCbanupBtK0Oi8pvMHkzE0B0Pf/qm2GoaXUFqXDAHZNYwp69HL0d1ZIphOObu/g
n2e6l0p4n/kNJXNZ3nXyaVffolZfN2M0LB5prkS8M4+qmRswPCwWne+SwXuyTwLhAQnnjljvTzm7
N/SWJMguGGSIKBHaJ1wdIgS6Hhz3gEpJsIGlWiJYMbIcWpTYDE/sA3zMv0BqfegvFZDcmDgDRX8d
7ckBJMvV3io7xCBaSN6QmLdUID3gAArYHpeNCVJwvgXeQM8oEZdk2kkNEDltYI63GMluCF91I6HT
42RCE7iyxL5FWE6KPvgsp2nCdqNdnUdmRhr3QV8g6xuFeRD3WtLboOJRNX8lxN4K+42rsUgJxgGl
C7FY7N6pY94oEJD10mAbxt3QpPEy1PQNjL0KYriFoDyg/nSQcBszzh0SYmQBcF7KjeyH1i3OJBJo
+bfHjzr6d/CLjX89YJMPEhUzvo7ZQiunoIBF7NYMmsbJoxO/mYL5V7zeOyRezoKOKb/EtjfGhrIO
RqUV3e1I+PZDlDAolOvRq+YtOPwwHV2fRCA9bz67frxrOIbpXRixNbus3jIyPxVcZPK53S4md4Fr
fLU//fb2m2s9wAmvWH6cwVxnfTl7qWzhL2poS8zUE6eSl4h0wKdsWObeRG7Obfyv67mrsjktZE9a
SV8Eh19d9YqfTr6UEsALg0PxZ60GOW6/r6EcidbkJb4O8hUzU9c+aT9/Rxh5VsL39yvnSdKWQGjV
hv5AVqbucTf9nO6NEINItAJlfgPlwQXHdVte4GgRWoFGssRCpkPiUs5K8/YpH86EMM6YOVifx0C/
45r4cxG5GZrBq1lgsYTxJooGoC495yHnsMcYFwscpdtRy081ndJhP5biP6UCXqMDGIuJUSbz6fdf
AE1OSA0+zlIPwV0hEsXWJO58Z/aXGzptmZgul1ofu9HTvnUzHH2/2XDWQbRRGMb1f9KE30n/6tBT
5H9zvZrwsHbVf1ce6oIPxW4Zp3x5pqvVcYPhBe8G7CHA8w0PAby2Y+D/cwqZl4FwPsRMODt04Y7K
uzTXgJeO7PjuU9m5jxVllef2FLi3b42d5q3jC2AsXk2fPtAHVS4I1W6FTc4CK7qVncYNrM1EKHHJ
PnQLZGUT7kyo+jG8hJwJnjIJSVzEA8glFmPnUVHTzw38/MgOhBZpTWSf7Lu9NH60UlFcxEEUM0yG
z1yes36td6LCZBtg44+mGXlYjuX6V50yBaEEj9RBn4XXv3QIo1jzsadjtJY/qcO6QrHsIcyUJEML
IzNzmtBC/CoF+wTuCnLgOuStRKreQfJiGUs3xzX3o14UL76qyYhQ8uYHkMHjPBnTPAruvN6hGkFK
l1ExStCad7e6Ze1dqm6ShiFb4pQjYACvZJgBF36P8CDK5YuXoeM7jwONcHHFKU00rU89n2E+PZ9U
gnaDHd36DDE+bjvJhNSd+1rGxqw3QwDx2l/npP9GBnmzmIxCGATPQ3qqorSV3wQJGybz7cFVRrUv
Il4IuAzVg5bvF/J/yBRjIqaLsvqIwEBjA3CxXhjU1LfWZIv1q6y5rxO5zb93AxPnw+egdO14DWE2
94qjX93i1QvOg4oVJTYy6qt/Qg1UX99lv8ZPU5kZGSlXz245kcAfQIY9nrs7Cuo0eXFVjlsyI/XY
S9ncDu1LobImW41WRjhQ+nrnK1cl+Gp0oOzBF8sCxi0aEY9t9Fkg4lRUxafOcupsDJ1StEoWx0o7
yFdNRSq9CENnc38+z1aoFQzeBJuZrEgJ9TlFmqm5acEmrp6IsFH4gmTZUxLonurbQXOoI3WfCYRq
nQO7Dv6QnMrtH/CbErnRrSbP/gEF11IEaxFXSawvnBdzATqjdaI/a+B519nEQ133QtYfRoN81S2E
YK+KKNS9DCFbic8M1vc4T934eXFKHhmv0svSvHQ0dmupz73VvfiaS2FPcnkjfED8qn5RtykOx1oV
70Z+7v8Q23XXL1BmPFHOwuXixXb/q1cryhLiC6oWTnScKPcPpgpGiWj+cHV46WhNSXu3UmGIlarc
o6VJxN2Ub5FRrV6HguSyKfAU1hA1VgYjbOYXaM1i4vHs5KhgqXwOV01xoC48Hgpx/NDs78K9v4o3
Wzs1Nf7ut8kbbPBF5Gyx+nhmcc7C8oeAHQbbK2vTx9aDQL5NfhT2DjSi1y9KWkFRW0XgpCXmmjYd
kgbEG/2/w5v002JFz6J2Mq5dujwsBBn9AKOR4RUm0U8ZN6rYAf5c0KRzY4N/xX1ZYdU3s33ohL/K
96/yuJWVDZB6L/QQpwNOjdg1Jo4UuigQRvmsrIIo8kOGswADMjytvz31k73U8td+0+8E6a5VpsnC
e98KmVIi3YOEg3XSF/cXCYQQRqg/rzTu5kWFCcj53AS/qyHus0Fx9HlUceeG+iuCVyNWcn5GeeDF
knqrvCnb1iGPVLWROYdUpMj9VNfHl/lT3bovse59Kzm70E3Cgwo9iVT6Vi1xYp+KNrnq4sp4E5r/
cZn3lynITHtWdMT6thv9qaMzp60lMCp6g3fXpEJ8KiCCcEzSFdAvWNBKCLmut96e4G/qbWeGedj7
I6RrA5cmyxbAuD3gzjaunexlhsg5vquabe8AgIPaBD/UbX3AP2w0AvnmN88sPM5XRunu68qducIh
VU89elCYAHRNMNiejQVKt1Nfe9tkdSZWRagzKO1FwopfNL1mgNwobf1TU3q7Kg5eJ7lbzmhYWNk5
zXFRM041CH6jDFRHWIsjrF+9d0IMrpczpVmG8WOc10/ecxeiAB9tL31w0I5yKfoxMPFhQlI7KZAW
lLRmJH7qi+i952V2wW357MMJYtZYGQa6XwGhjR2Wa7Y0RPaFPm7lnkhFNaIdPzDDrvDkmfamL1ZR
93+CZlwL7Zsnjgserp0Q0kcwlRirQgmRzqDlN4JXLG4aw8E+PWlDSlVbdPFQQ/It6UcSiyyV1+2b
h0OrIf4d0+krtA1aYNrxxVUTUejC1UTUa392iOP8uT7F9u6TTNIcbSxONfZJNkKDbhOgsMV/fx/b
MdCx3vOJbTCeCDrQ5qMd/F7iY4o6GleQP85XvJx8cro3R9JDc3bh1BrQ+QrqFfBVPKDFk5MJ0vEk
mcIBZjIgS5rc7i03NgewAGCIbepzWDqoDL5bNIEZjmhFscSMTzVANs7VTZOsX91q6alNWWiVQGYX
bTRyXJ+SeMW+ZKDt269j5ZWnziEyVDaBfu6Y3/7cj85YjNXV/oz7lbUrLI/XuFf0EY/ydqO99xZI
UKwBmKjZJthEZxm9nbaTxC786aZuG2NJlrnilioIqR7cYBFPxHEPOSDldwNt2PaBa1KFHk9j3dom
l1Nqh2b/Kq6KHR+JgbpJKvUqi5LekEYxAbflYd7+iz3ua8mPklFl0r04/i6A+Zu+rYjMxIAnkOSV
R0gkdS79yojZjd03YwBGETAKINEMjBktZNp/LPeB1sLBnh6afK9F9WXvANB6UCa987H/J8NoCTBj
T6qljKwHSOk+1AkgIKAgw0OLY5eqROhgaKsSSVMbhZnueMTzOZ4NtuaA9L43pIEcIh18fl9/m30v
5sE2/+LH73mnamQfQXc3h2axeQSYC3jj6E9EqogycXhc27TLDXiL4g18pTyZAeTEW4ElHBGRLwNz
/2DmqX54W6K+zOn2JFCIfo4DVwjCfa9/xjgGUEazsr+TOcGcAfGsCLAsDeCttGYOODKuxWp8k2tr
b6/6KXhj+nxbr/1oAIgaBhMV1/HHpdil7qUVk7hgt8wA6cjkf6Ehe/hysAdWvx1Il/TO7HCJXC9I
V9elvkpDFAWtQjzb4j0uOuYcz/rUX9ULbd9o5Oyl1QvkNg2iOiikYA5WCrSQwRIcODJpDxwVhfjY
L7yb1aOhMgzT341bbmvoRVDatw2bkGhbhL/o74cIjvjBGvMftwIA1z/TvcaWPpFFaQjjNcmUPA6+
vIKq9FuxzLXZktkK/h3d4c7qXZK+QaSj/U7E4yOzuEh7ZkpHgGggrdOfVGxmQaNETKL2PJiYG3he
2+3xcRHmqtdMkFYzod4XMueXZPcYFCxlXa+t95HOz/UCnimkmWMR0I6rElpGXTDxDVK13jYM3fDR
z+RacRc4SeaptKOsw4yHI2jWxOBfmpptd0jr0LEw8ljAP9h0WhX0UCdZj7S/CS9+h318N110tIGm
59irG+iMIgTKP4ESx8L4da5VljKk4CN/6hCCMks4J2CYj4xHqeRR/837Rg2nL88FC08VnmvbqGoz
SKCSlVdP7jhvrUW3R84IShPLirv3/CQEksxyRVISCd5H2Hn6iAeH1aHqiRoK3HWx37J4zdkeMHau
j54gIqfru5dLpjm4PFP+dKVLwWdqPgF9QWkbw29u9Zs1JzV+gLoQ+8YkvHZHeM/WDe+fS3HSISzP
Dl7nkOubJSpv9W+VSZapQGDlFXmKxulpdWZUMzxtx7fKelSIwv/j+jtyyZxEAeesyHRY4AHVneu6
khesTxIGeR1D+mo3Iyl77xITvgdQzTBvnYGFnk6oqZmu7LbJgIXtOxCbswKG+rIU5kS4mKjwo8yx
OqZoJgbRydj7O1+XUYFCLO2CBUsVqoIzWtibgjrmAhW54bSQMDzRH1Y0QiPOPFc7d+WMCPthiJVS
/5ni5jvCzmm5YonmQE36BD1L3AcIGKJNe4FPtmceLMQnmTFha4l7jPWZAnlVZ0Q5dsW24jjKsSph
OHLTJB30qJqg1Zw1hL89u5xgR4GeRa7L02NhaujwX7VV7dd10QSBY48MTgyi1El45uTMqPsXEadl
04kAH5PREff80KfB9t5WR2g/ZQscsrjql5aSxKP4eFF8G+72mYd3xMMVx8G08f609J9YvuBjOvgn
4NCCZ3dbVgPCGWf1Ngg5KjlVBnIGPPAri+hGdcjCYM0IXV76CTjI1QBl4oAst8200srefcQHVVFz
rx+ifVUlguzdMpGg4nI99S49dEFTQ3a/nSrtehkqD9WrNXSEkRI7c1Tti9VX3t9CMMVgZbDxhP+o
RR7347qMcQ+WUTLf4v/tuBu1MA1xGoN07pOP7Rk9LZI3kyzH/e9O+a/LN1R8GJIIcW7L132gsQjP
BvTMCck9GNCYtAemtvrX4vbo0HFGWwC4uKhM8EErESrjB9JwbPT9im/ERetgVhI7n04hivOMq/bs
LQ/dYChCsv1q96keAxWyJCxDlaOFlBbsouDvyfW9pY+eCWtzIDsNV+me+KkzEyGJ5K70boJXl7rv
skycUNAOpaf2us0GoWQ5bpl3ikv5vJc+88RQcqwjP7aaGZHnuc4C9gvd9jkRs65U0MB9RvZWyz1S
7zQ/9xioOfuTVBE+CuduAmzdKaNiYLr2ddpAmwKwjCy6GGCuUFHoBNNabawverru+y2YEdH6VBfa
En45VZR4GYpn+14DzjdULLhn6wVNdgiNVpkOU7oJg6FTwTeIoD9V3cY/s09FtfrOzPTbXVC+ONWY
hPeQuRVvVPaXOzYJX3NAs/7Si451HRgdFnjP8GkHxQThHUogvSpdAuegOgOcwxjp0jMFlnXu91Uj
oE/qDep7JN5ZqJx38ZsFLSGHpK+7mglxxtkVEovxC/sQH/gRmJts8V3x+d1gajeu+2cKCWDhWAKV
CyqqU6JopGm77u+xyV9Ly5NVx7Gf5N7jHUqQtp/SZjNZoBjBSohLM7HSk2gYgPWJqeSwD+0jvCp1
sug1s7psvQOzrJkYtN1ylw+dk18fa+VS6L1kDGIM23GIgOBrmSWlK2p0lfrwGu8SIAnJM5AwchXN
ospfpcgHm4JZnSu0PclMUH7XLwEaOVIz+lZ4iDXpJdskM/f2LoIXY/JF0xRs4b+YAM/xQpGEGr5e
7kUPUxSR/X2rQc33JZz4ubyDrp1QcEfYEK9ZzQbdS++bcpjNIcfD4KRPV4RpTM/s8rubL6U9Z3KQ
TiTsNfjp4O9952+n/tdNis21PwQYuc2Nc8Q2D5IN113KidBQv9VtYml5fGGM0RrFFtU5fx6zj00i
8VQm/+i8Jt8OEW52YrZaDcxndze1n3GbZDUECPtVOuuoBOzARaBPgYpJySrs2FDP+qruW1RsTLv2
uaFLbrFK5ABcjw63+fSEhXpztB+BSCcCdgimcyOJXiVR8TI7oQT8eOIqpuGeoNCdeWeAeh9v0yoL
4lsaEdaT+FdXbLpLYuVtEAXUMwSSvdOYqdkzLgqHrGqAbiU5TPFJySCv64VH256faVOukvnv9HZj
yoVLmqQsYFwcMjHgAPi2WsDUI96GtcPbISBNZ/UwJ8P6W9xaprJ9AfNmwBWw72ECHGln8By329pP
1WiTJpHhdWRPtO7yjlMwqteXZjzjyPe85SMf/B1k3as2LqWQyiGxJAS6szrdg2H4c8MUZgCi7YrW
6WWuEuNuTLfZ2PSNPef7jUX5oGUm/zWCr7OHpTL40YfxTYuVdvWY1uYH7akiORUrh5+UOB8jw+aF
VW5OW82RUVLyG1mZGzpCN1KuiyZ2MMcc2Rr20H81G0kkFzPYefuAIjFcSKDBBEyn6mT7ikvErnVO
RpGVdLANfyfCbZyYN4FLjzG+Ca+hwcjhsQnb6fKKf/RvT9I4GP1bqojzgbLiyI8td5wEH2tQCX3C
9/vCCZGxyiSGbqgqAQ0EYqThJTc2U8hjdRqkHgn6dZPmZE+IBuaYBdeFFh3E4tQ7riJFpEzqD+4P
mKax4egZb88iOQdDhMWHImX6HRxd3dCj+LLyj23CO2n+bW8RXWvC2pgPOoPVYJ1escx8/HlgaMm/
XBXlpADPKuzHhwacilkDzTowCKpmSsTVqQPDCGAMddxx9WpMdK5RFn/ItVYepyqX/wA/ulADPGpY
zR5cYLEJKgNbX4gCC4gf2TpZI9ORJofEtW58eLmlbMXrzc9PZpZwEQ2YGS2tZFHye753ZlcFbvnA
20/c9H4D1Ebv06cLsNjwJavCEzTiBWCPQU7C8oqRuoc7nKy32MzEDAu06jEsbQm31NGcPEjhFso/
xi8q+UIZDUpE/yyud7PmpSeF30ICxFZ5kqdchUwmrGN9WwLcSS0sL32xqFtiqT6sjsYam0gnH36z
URy7x2xDhK02gqJjAYg+x54FiEVJh3GJouox4CL53spSrHgNDeEbosMwDoohBk4Bc3zj9oAOmbHo
ZQvW5Dq4IdR5hcpwcYXJcKuST8ZW1B7+9S5ooSvidEKkvQyDgNgIcegdszapuJB99SmthvYb69ge
3YA530iq8rb6Ly/coxIGbEwndqDM4vJFw+yFgQLgwogsUnJg9fP8PNl67zEUe2wle/LAQsmp3UFt
YmPR/Fw4ce4oI54usHHCJokEpTscPviUeTHcU3vUDEWZ6j8CAfz2a3os9H1D7Mrn2C6oWaMTnL8V
6UIlzdJhsThXqOCDNQrvhmS8+PTW5jx3ziKLseOXOkSt7lU4XWPAiySm5p3trBpYvwLTdRY7lMZI
xfAzLuOD21C1XEZOHo4SZFDQu6b2pxFcbsf+Aa6i237tZ38CTTje2tvJab/XqdJo4gP9TbY1V25F
BNSWiCY+jVVvV9JFQ+m33daiyrkR+AdlGfr0dRZQjOHEFEzDEagCdz6Cxjh8m6OgJPX6X21kxpdI
yby0qSEIYmfGKzIL53Pku/opnhEaxVVR1ClS4Eao5HHZ7XICWws0i+od3uE+L1CJydJzt5aqPMn/
6dCQPuFk1fTcqUIt8Vvx9Co0Amvheo74i0Ex17eW4hBx3dPNxhWaxgCylX4rzDoWXyp7zBiVHC2R
JodLvmOSMfhI6bPGUwihoWPLaORqRDtYrEZhKyKqt+X3ygdU25zCs1dTlOS9tWSfh+mLYB1qvLrs
dZjmVKhiF98LAhHAGCdM++Ozuz+VdeOMVZ+FxHvVPC44YHno9o8WSc5khzj1PaRUBn6KbQDM+Vtg
WvO3rrT2sNwyRKdQnlHhUf+WzSxV+2igG0vN5yJTa2HXGtpfRTCIiSAYNMPhFRpq1Z9sgeKy21J9
hbJw7a5djH2lFK4n9zL1fF4jpfGkW+EF87rbPwbwR+p8teWRloNG68Va0V2p6P+ZW0ZIW/5as8gE
Ez6Iwx4FL1h+eS0P8L9OxTFvArFxCJAeogRSVTWiOeKSGnSPtbAqRXw8f4UNHkDAflIkLLZMMxDy
CULyP0NvK+lch2Wv12raM4bHOyJYo4KtLjIyN2CpJVNfdMNZz0YUneJUWRn181PaMeYM6e7Wyc6V
5WlJOH4QuqcbPKQUV5IRBpAir69IS6Kgr2P9ocwpM8mETQ9556gLPzwFzArm/74oDKUZkoOsksVq
yX+ReAAztcZkl5IJRSZzQz4x7YoXyojRMQ7xKzYM2XRJz0hguGCeLLpRfsrxzkiAj18nFt2GEdgr
F3hQkdhuv52YYMRyjJWgqCWk/PzeZ3oJgaIchWgVIC1gawQ+u4CpCzodd7Tu14x3RXztvE9gqDqm
irkfxdKdL0YYF2XiixbQwlsbzlkFFZecfa2RdG/TPy0XYYhxc8npyK2HNywdyxK/SL7uNlbhAVFE
tVPs185GBMspZnv9wRvzJtncPdITrgYiGFmOzGRDi0RMGklKRVBnfUpXPa0ZuXmS1N63mB+HQYzj
24vW7yQkERLhkIp8/3pZoPj6BQiJuGaFqpc7D4IFm3USE7HDCaegzIf3NdrKQZNAgqeYt+3LQkN0
PkUsvVrQ4FSbC24pRXNJkLGyPFjEJVlXSkKZigMo9BbEcPQO6ymSzPRWtxSRbk1JtwiYHeaopXuI
EL8pVxrXQL86+XguIPDGtStGPjU49zryG7w53IDpCKHGA4lAvaDpc7x7M+AX1BSkIrIqUq8TNU2R
Y+9tkM4t9hW6jGoWxxboJQrq/cSrlui3P2BN+rImLmrzHSsyrBne9tsxw4iXTf+kulP/2Lh8E0dq
SSE9XpaXk10ByC2zelYpsGdDWdmAgKpw0ymDSQxT0E62fR/Wim1dqobJhvFKxKefU6KMuuaQmXfs
TmH97+RFKk8RWlPasgtB924ytkB/mejr6EYg3jUGoup7Q0N1xmJ2I/E8C/GHGlM14llKXLfKMrR3
MPNDFyG4XJEL7QgsWmsBd/RvM/kvFdWf8aYmJ1ZN4Ex9uMOS/wNI1TE4Yo6RMix2P+wBuOVQq2MW
O2GGAxLRHS/x8S9+k/w5CehFzYb3w7IOToFY4itaR1NaMVw69XjJgws+qbOYDBmAVV0RWlf7ncNd
QD+/KWnzlAYtF0VzzD57z9B7jAmtLUxY+VWVfIi4x3Bt2ZflN3+Uz+5QlWJXE82MsJGDJRUHDY0r
b1KmR1bS1jd1aiencpF7Quph8vAwBR0MzAy9Tk477Rge4qihuMyoE6uUtCuXmKBRWqQuIsj2V9CZ
lFraKVoVUgSj8f70e5beBTs7cYZ8V5UzE3Q0DgkyydlRZBrz1wN4udm9J+r4LwhU5ydAHpqmPM0r
oEc6NIFkvjNAzGAQ9MKpcxDvW2bKcWLClz5cYZbyILkrYEAnSv06y0MTIZeNwCzRyXpGW9lxqUfu
PODtC1GQ79WXZh1/zDtkFAaqwcLv23N0HM+uvrVJevMi/QxOYbjPCiSYoHWJjUt97BxFZ5kG/Oxn
gJRkdoP2s5YaDBgBCD/UPAlNacPW5p0tpr6mjs+L3NGAHSxCtXd/qlvJtpYcMVAYhlcEpgp6oAOo
urgnewCmnbGFsmZSGtQYyIioi7w27PgIhXqqrUzeExufIyWgMRUr4aLxriVEay7Fj/z9QXLNipFt
0al6mkmkdyRFL18BMprkqEb+rVDgQbmpUf/pIp+vLgJx5+O0BNPUsPTa5vyaTyiZvhXhhuMD0Vy0
lgF/CTaMJljtlaUYDgyiPnWegreZtc53XQR0Tfhe7f/dM7DQDG+aTyaAujfeq5z7JYJ6IIJVuhr4
24+stE64G6ACP7/c9RQmd4IxsKO2sV1sboz6QLSQEwQk+hZoAK0ZMiPSEQwA+8B8NUVD6dLB/hWJ
R3E/hSyk1J8h+ZK5Kaq8Yf3GEuHu8Tp65jrlc2eqtl/t2C9FYRPmu6GZNzdB7Pq002etdiFsckGM
NCV6ADLiIjprkH9VByRkyHZx9ALmQbS1HPFfX6htHgd4ftDg29g6whS+/PBHye/Q6U/a8p5GQ207
9hDoHCCyeoOsOb58JEQ31ajKcTXPtjlQsNQHlO9lDb8JdLRR75yuSbzflZvBqTwPCkQXxU5qf9YC
SuHqdd/FywnHeYb0uFy/vP5DdcytMTaKY9g53d1e2XW1bh0ztTQHYORmrUV4kqgUfdaMDELfl5Kx
cbKtL0vAgijgNAmYJktFSVYHYPG32Li27YwZaPRAhuABPd3bMtuBk7uootHV7R0Y/DI9iCSaDrcI
QphFMnAF8sjuzRZ19oZodjH0LG+EiQt3q4dAE0S4uLFqCFR8Q/NrQ0K43DQ5JlqCiQb5gZeaaalX
6jF5vAc2YojpUXem9NP298h20JNZUf3zSWsdJtFcfiHfTOHQH7xDZOYnZyEZtILOEVLISvYt/Dy8
R0TCTFzeV8n6FsDmbvKpec3RuyebWMr7XMDZ25OvVJ0g7vpS3PV0BNZSCp348BuL+/DsH0y+4+gI
3ySR8LwuSc4jAtgi/IItA4zNbbMKdru0BkfQlKyAuxNFMeOCkyvOhLGe3uWZIDlz5iIrj4zN8HIl
FwntamkgOKK1xUraKlHGe78SYNQaotTk9jeTsZlHXLxNKf4LeLROCEMmN9B7lM73fanDEiP1MJ88
NjCNZstbrdgzGk3HhPmhZ6y3smKyHJx1stTlQ5MfnCH4zI6iYxzxE9TKZRk3rw/ETJXKc0ylbwJp
X1SbffmEWsF/0OZoV1+NzhVfwrwJifPQytUYqitm+KCokcIYVC6KOvLvVhlD6gFtWxNpCQKpbWnv
hIdJCNoWHdW4aw7rDBRhRp2Xd3JmAv43/i23Yetde5+JzxSx5NhTKzUScmgCl5nXJ9GbUeqAuGx3
lTLIT3RVAO3EhtfhWCvoqupL0+UKeSluGos73DQEQOGslwTAfz8X03Yiic8udxrVB0wJBr2x552x
Tca4Ptdq6vG/MJ9u0PzEWIFvDgMssCsy2KFvlCw+iFARMASquVgOLC+AXCs7EbJwBR6ZLXixQSk6
s93LvmwsHCRG5aMMMrhT5pXdcP9tCrKjeakA4qn3oeFwDzfgWCnZsKeXLDLKnpmJjU0XFA2Dn4j9
KpQdCYL8Y5U9iGZ+05wxsvdqsS/7C4T6RuKR01OWizjz4p+0eEdU74z604jAwHCW6rc4AfP3/R9a
f+bNX0pD8jiqoJcEPi1BB+MxUhH5uQ0A8amliUzC2GkQwkg/pPw3HuSrV/iN/6Kg3nnFm47sU7+l
wzVR0y3/sz2SICy2ESP3tzgIJH1dvAnIR37lbBMgXYs1HgGWo6SsaRAegsyrpQY8EyI/0TRZL2qB
CVo0l1vVfZbJuV++kCzzgjKRmK9waiyQbiHfzlPfIJlvAgsLrfpkqtofWQlvWpMctq60d+UGgFGo
ZeZbU0/xi3L5hSugstqZ1wSpuTgeAdiNyxxP/+sw20JJe82Rr5956nQB1m6oJYHdcMvyPPjo2Us3
jqngrpGjWmjEo4BslNiT3VSsj4J31gyyiUOMh6MLf4MmTcf86RKKWa3LwAJcE+IuLGq8zU2C1MxM
z8MEHPi2EpZ3rKGFlXiEo1JtEUMHZM2xZGFr4l9xdUHiSuYuvG1WSzyYsVdJHyVJ4NavxjMAXAnz
HM+uNW8quJWgANRLCW7Wjr8VFR/wJD+A9oQAYRN2S2XqkunYjac/WHwxZN1EY1ZHJxeYZJcUrjKK
Za9QcUEoDP+wZJma+iPw6dp5X+tBkOg0VYibXZnzAi5h8tznI21eTVc7wB/bs2oxqIUa8VepLqiC
8zJEoURsWOrhxKizfqXrFrtJnaFX24plFxnMQ5DLqQyTvjMzOIaZweVWlVtFwfpSqItfpmjhUgSW
9hgBwD3nt17WaSP413zhdwTGu1711gahBSkJIrCrg2P3FTsMYnnwUMvZHrQ0HkplZCt6FhQIch9z
n7JkjeklVM0jFh0DGgEnduMis6p3QT1E8FNZ1Vjw8e9mqr3aXO5P4r7e3kDzsdmX6foTKr8/W9ql
XkO4Sy00r5IrT+ux3IJ+1FCE1icGymarrbEy8ZMpvCO0cNzYJVR2aUCBmZQtCYE13KnO2bKdpP7/
1zpLRbR12Dt++Tx+L3iEd/Uphn4MdVILDDsG4kM+8zl5HIVQ+NF89jLRg7KcJ76OPjOO42GTwwLh
H2UFH4HU/PLenHq59z2sv84yGBKzYgutueyjUxR+L3qsEk7O9cl2faIsAjODd2mUTx7UgUNACJWb
WUoqqW700KKr610cNm9YkP9P1Gc1a6us5o7DdkNTBQH1L3aGSXW0sAtVi9XNMuSKkDhPP+WHfw7V
bc2oICJ184jKhRDE5nIgbPsrC/PuxtvkRfyu3jAPdUS+1o2vHfIh6vWGYzGTW527aNHiAbdNI7Dv
dL+rFc0uUYTUYUnniFsElaGtHm3NJOaYS11IVw3iRCOw6GbmjXKfrJG0inoPIKQXj9EmCwo8nYb7
VBvI8LvKqBr8rl7CIkwR9j3LjiT/ti5p7HQHeeX4JGhebEZ536QT3FP9e1nIPNCxa4v4c+L6gfXP
kmJ8vmjDJMO2dIyIdjVX2nxO9NAzjdrSQ0St6WpXoZ8kGxI7pDDa7gBx+vwr12y3jkM1xWp/xY6F
iogbPQy2eg5YdRZKCg4qZjVrcER4ZODPrGuNGZ0H03kD4yzIIthU93GdseJf0ilbWq4L/wA1/0Hs
XsRPIQThn4CRF64aDduoOGArgzZxFWTAI4pewVNfbdrU9XoKM7s6ECi1Kj/6jVUp7Aq/GnIfab/N
VyCvkwOZ8+GEWmkRMAcK4xM64Dpb5ggvm3lHqdPBIbnGPA+F/o3JIeTR0fdxqZPwxL/kPGSF5PZS
XQKiCB6OTebOLT+WDfAPyrAqkroe5zLX8r25cpQ69Hh5c2ZDGsONZcwOm5c9PBiIfhgmuZTFBfl8
Smu5i8Xt08e6z2K+H4WGBo2xyuMzblDHARxiniz/WqfRwVDR+3DqRpwkfNzFUiC05ltsn3fNhEx5
dloiUw4bKaC5C5b0u+0yBixhoJfPdzR+000PwVlyIf9mLL7+RzMeyhtRDXUPd4dlIvrct+hw9RPp
AXTLHJO9OHF97qBRhz3gXLbJQLsY83gbokAJc2ecu4JAaxMh4460O55SeCS7XpCdKCLu//E3uZte
b45mKd3OQme516r09ckqGEc6C7BQC2eOrN9g3jOmAVVENaH2nerr2XMMSERst/IqNdfvQxZbFfAF
uJZZL1GvuHNdzNlKYABSRze5XagR5cqOVgSgqY8/B9kWTBiNG+jJP3ASJkO91drKxkp8JT/+lXjg
FKuIBiuwtIMQAhQfl5RUyzt+l89YnFNFhmJtAwZV0K8hDIKiItxRCLxd1TdyvKjkp7z+MeaQL9nL
7BGOkD0EfQt1HT1pnu3C3NTcF/zPFQSbvabsLpRisT8XwA9qgJcAlyslC1D74cY4ChX6Y/FoELSs
jGPbefMxN4RqUNjA3hJ7QKYJjgy0v7VZp/uaOPa31OEXVRfnT+gvtNJlTX9OnVBul8UbnTNn45fK
zpZFzi+e+GANreDesITQPVIJgDL8ySVc74dmUNe2XXk19jtGcKaRrV2xEeCsTEUuw9OY3UJF9PDk
XRCBqYpkrg3gau6W+Irz/mW5dSJnVeR3uzSR0pOPKAzqQkzL56zPXrzrzo6YakWbq25F+UyzE5xF
9aFPvFIOATeQQLep40jZ+IEM4Q1Vy7bk01XhpQe5SwrDSthQ43MQrSZPga1VfofFq9bMpI566UFm
PYoJvzOeASImCqvfSGbifZ33XjnHDhmQ92kSZVtW6JjWyVmLmsGAKzSlHTWsNZA4Q8LOxRmL4rHF
iLb0fs7Ms51a4WzVuVmfaPm11RR+T7amk3cV/8K5r16gV8NQ8aUkjYZsu3A2jydYyBFq2JMEbfVz
5l8tvXACl3GzGuGBvWuEGxok8Im3wc2nLOE3hBpZhS+4i5zeT12t4MCK3eQV9hKXppkE1UwmoKOD
/k6EJ5x5DASIGg6YyZVZ0gzqLaLb0mRCCiYl8cBX5CDwsPwe1JISt+vxpsWOLHe0e+TYSlBSBK0X
avYBj8CEUqUaOIdC1Yo6kJsJk6j1ToABMbmVtO0bVU1OPHidbvSDANnu2OpG1pcSDOr9Zv+3195G
uhonNOq4AOgYSOxaXMIDzjf9pJLjN1T4MMuzABx9WtfWLQY8GGSzKeM+zEBYKSFowtnoLMS80+Q7
I4xBdXmCe3U7Xe1t+tA0eLhpe26+3fYQbsBnAaiPQmtAdJ9MBX99RnetjGHC65F/NzYiPWmh6onq
/3U7S7OiB5L1xnEbJfRw8jlScsU3LVpRH5Y3YmZ6kV0CUZ7FKPLWbj4xcrONbUGUDKzvvjhl+Htk
OV3bw8c8zXBkd1Sb7UfuFdXsLdFwH/TCh4lqodd6KByuCBye+//55qfnlc8AOIBLSiUEnyjFWNk5
Q2Y2RUXhjuN0/kxDBFjzsBYKaRmVUrA5eH8Ng7qMexAOWxx7jbt7isZ26LcEu+mVljRPlA3ik0pO
ncvtHOrbuGyEZPFEVbXQPMG/e16PzOFKw0WkOU8UoKIljb+xQ7HJGBswZgyjVXEPao1okxAkuaet
f+LmO+5BAtiCWAckgXP0f7qGsXBnhCOHGPWYADkBu9JnvOK7KB40E4waIg1hMmIcs1cjtgRzXGUM
OKTUa+dR7EGKZ26NnkkqqdHPl2SymJp+gzgTfI63wv1a+YU1OfXk2SOZIb6lInzvLJfLLNX+Rqrx
xuMgNXnqQBqojj8QxGDsPdaURerB5DrEi9qM6HhgycwnOFab1w6I+TXvKS3fjANWEWIVTENYk7O8
X+kRzdliKcKvITjmtirNCwkv17YaIQQLGn9JQf/YpwoODKjW+TNjqLP6XKoRk6chkdT8SXVatkTA
twg0cbMW2XhvojNNT8D+NBM6DughmN22vay5tP0deFbrfaa4tChno+mmJ9IJgE+ytId1AvhVgDtO
1N954cqq72EKAnblh2+V6zly6txj+agKR99vVJ+plvTCFwlnsK9RJ1E9hVyyqSaKiBF3tVDI0HmE
ufawrRxn6JX9K67J9gzRBehz3gwqzKGYIXjlivZwp6FpWvak8q2wyAA/XJm99J9JTw7YALBSI8No
WO9O0xiWDaiOSc+2v9PmmG0goP0Olr4tYDEKSRMT7eWEcA8Pmp4isYBBbVKup/u/Rj1DQhqQBw9N
HDcsLRpSUEA5N9U9F+hE9xUi1+6PcAhF7FVnugUvm8lz6zNRK0mCEgHHH6EKjqwyqCRK6IDK9U7X
5fyMfqlaVkBEq7EuzTtanUWC9S18rK2HQLex7450tpCCYQ+gqfEdtVKght02euPoSqsoMg3tt0p6
Ln1qf+oef/i7MlbUbtdUS+slItW39LHP+BhgMjO+dEItaf9igFMoyX5shVVnL7I5uMym+lfGOHpt
+32cTAe78yC/KzXpB8NeP28JaaWGRKQs9Cd7lU5582P0Eo9I+Q+33rVm1ZOvOCR/cg6X489Cw9h0
4z/gpR2tmEFTgLEPJLhBtpgdSU0Nwf6kHlneGTq8SX5nkwzxeLWcy7OJEwGS93ZTlVnZUnO4KgWw
j9NrC+uCQHS9RJm6b7hzo5qsS7HmEX31XJ8/Z8Kw5BB+g9yZ6/DDgcxW+YHQfldqcsKU+nJAEWMD
tB/Yz+wtoNobImaCTYshMTAqoWQduuBREmapZhsfthR53LELP/cWOsW98i3n3eChCelf6L3VUXUy
J3TJYXm608gfBZOwUP8LA9eulj0OHdjo9gevWIKESdGXmYlSM+EdcNwFeTpeto+h6pvybxY1fUA7
a+rm646ttad6V4B4XplwxeE62dG4U5AWkhaKhzZ5vce4qY7j+bzljHlf5A1FjfsxGKUYLjT0UvhW
LiAUbpmP7n2pS0n6+0TXEWA2ubLuBDoVFFCP+hL66e9PhvDPV/NjO4sD0UwhSmdjg1K80S1V/b/a
dWCLWY1+vzuKDxOMopiRCZmWK8hUyeBbPc03PVZmZntqxd732jCbTSH3d24vDG+a2tS4E46hkWTl
Vb2Pve/q2P7n7YOmXNNO20sR17xnDr/6ZHFjC49KVyVbzKeUr9RZ4kN61F0runVDrusOcoBp+thj
ErV+2fNjFwg1ldJXMESHUCIQ8mY5rj+ShhPa7VUX49qnY5aTJtATgR3IiUt+6VHKRT7UtrDWAVtt
2tBPRmrs9xqLiz3HQuGsahIV8NhaYQfPrBrnWkwOa5FzgSBv2FM+Vb+YIC5twV/M1+UZFwXpMv0N
QqOWGxHpbcv18s840QuZ3NSoFVG0wWdIvx4H2Y71WUzRQ/jB2Xw6TRvU7F0jg9ULLh8jp7ZVdjld
mV7SSxpbBq399Jzl0oJ5ePjZH03dR4v7LvAixfrsPJuGF17d336j6RzUsZ4W2wODHu0TdKbcw5HQ
dyMrFDIpYaqsfWDQqQAo6tkyasb9ySPENPT3SkvyiC5rpPply80zfJbyfSjU8r02LejsC3NF6huL
iehpBufGNB0xx8QIXxv/Ykr2fvF2n4cmeJaQPJP5g633Ox39ycD3TpKFSnaPP5kRBTsQSQnYrxpf
QorhcQR9LfTrAiWuWdhdIklMm0GnrL1kB8TZODCeUqP9hoCx/akZm8DY2Yg8vLGJloRH5Z2eivkJ
liaM3tHAV8uWkXFK62+zDZRhPPL1kcKVNQ4fvPB3hMKRKkXrd5T2o1mrgXFe39/Doi0+sy2FJDWJ
Se6Vi6N0x9VcWzrVL6flCYEngYBw/Z5nb1qjfqc44ZYyMQ2DimbgIqHcQxNO6O+cArQMVpqcTXG5
TucJug1zoOBaq/pKKuK/ob16a/eEmjLxXUBzKCKNdAsLL1WClNou5frgmoDWERq5enW1aDBMcPtx
UNGELFV3YuH9qqIqXYY96Zc3xRa77Sr8wz8A4HGINBxavOLaPFTesVKrf4EzDna+cOMrXYwneOsc
VebViXx7BpWZwxHlGE2K+xYuwQ6NXqLhwxjndERFdVoSvFiVcSq5NFHL0IXwTcoAcgNbF8bDVDZ1
v3T9pJ8eYHCJd508lHvtBgmyuJl3+Jxq37SJALartcSv4r/Ynlkw60d6Zo9ettt2PF2+LWMPb845
MfowT1p982wntcIyjhkhGg4Vnc0pN9SZwPGHOIBMzKff99ZxuXhqsC33cBvAaBeaZn28JL8iSjdM
QMmoGxllST1Ans80+4n+AN7wsG2xaYhj4PxvdvqX+mgbIr1Ep5eKSCi62f8tpJjhvkH/KbFHfF9k
ovOkBqVE5upASDV43AI6J0ya5XsgDzudDjr/3uxjpJhzPWG7hdg6/MSq2ZcRef740MB0bOd7B0fl
L+Ml6Mu2hpKGbWCAWAaN7R/jvHSMiQ7zSOSaPialzYJKZFe+a/ncmXKfzaVVEr2Q22SlAwUhB8LU
P8sqAtvtrfWxYhJfoFFxCnf0IApbzDWrcIGgZYFdqCy1sapvPBz3UOgJPqRbq+HF2pewSHgV2ln1
S5ExnHX6gyGST52owWW2Dk8ai6gWaX8Mv4Pf7j7hgl8wrcXyTuzHhY2DF/2X7PMtrBlU8xDinm2x
v+/LlfqmCJalqW/WdQ1aSq/2+1bDHkDpwJS7GnECWP8b0GJGzDXjSfsdDeP0SeYp7KaKGrv3gT8S
SMwrfCpDDvaLMdepLoiO5tIR+4Kob8MbK+0d0EbWsGxzkFw3K0POX1IcBhpQnspWXowQLmcQXUgo
WZlRQLh79/UAz85H1RFDY0gPIUwPvrjmCuhaHX4hJizFLDw061CMnbatA3Sjrz9EfdmGCWxmhkaH
cDc38z1c42hrsZIoqYmIpCNTw0eK+/skFl/wDze42Ku0Mq5hTvHom7JykOSSPCXG8KiSO5JzwQB6
oU9mEKz2JC1axaRlhsCsW3wTQdQ48EckjTYCrQRKLIMOHnkK9jk4hi0Gzy5C9537RQdcjvqCu0Gg
+s0oUgHgVcFaHx9tOJIFSTDa3gLXksTnz+dLlUzGg+wUZEdo5UTsvjpR2QSDl6gdjiXhnms2ucwB
Em7z17a182D1ZHYUy3FIbOowo3v47u/F+ly1GrMVyIyId0AFXwv26DbYHxw42OQ/Kktz9xrjL4G4
1BYF9xpZQcXUMpzk21RmAZ3IPvF29XtW2gn7rvaRfSI5AFmufihr3iRGHLGN3Lkwy7sTPCYvEbup
ss83EQwqmmo4UAh3/ZesYXTKZhtCeA+0fHACakxkCj3R8lwwgrN7xNSeS74ey2v4pUvU/8OUR0eg
DNeL6YvvvqishfyWENPKiGZdM4KDqct1rH+Qyz18CIc1g7uyn6HWfQXdsLiQXIudVE9b56HrZlKt
IU5Wk1/TkE44S4Vy4vuM9JluuN1sGg9xGi6UTalCylBSaYjQSym26kqHjMQB7nHa+BBNCy3Z+SfP
umcVBSNIZPl8rAdOTpo2oAElhnmXhMhbyQ1wgUtNMuAJFB+rdDuW/BBrLZeOjaZkK0wQCWkMlnkc
ZogUwALq9nbHi67Z8ex2mrRvyfYyV9PJtTy+D9oP2HWHl9/6LXtYOaOcHhE/nb8QI/byhQoR3+XM
oyRo1e2LYubw6c4OE/HGnBgX04T58+StuGYebYfL5EHKruIJjW/BjhYxy+DqQc2aK8aZ/U99jmbX
6N61PEM9wAwU8dIXVV3yrUTT42657v8pE6X7ZBcIML8kXWh4eGMELPrUbQFBNm0mN8gY7zhobRXd
7vxL83KYK2ysHWQzSp5CGOMOnEZSNJtQ0YdstIRe+OfTzYMCLbxtJYVj26pD5r7wKQ3KOf4iBFEw
MDqR0N39iJ80gGWepnWf5Ub+unZGCrbKXtBzPFx0ikS17pDzVBfTBU5/WkDOM7qU6L6cbY6By353
Sq19HMKQ29d4hvG2Z+NAXVyvVHdCA/2ZZDi1ghy1N3JPFWOoz1u6lDurGRHNN8r8HKwJTq6IwzGx
QC6AxSOla4XjjKCW1XmJen1KUX7zwOOvqKIvx2X5GsLV7YLqHkZYU4I2sQCdE9YPMOi5M4/ESHsV
QOB8PCM02UT9gPYEvqO3/0MBXCD/kpdELSwE7ql+ctyrWIhKMCM+aW9pSzzbZo0Afp/1SLpC0blS
kJgfRAE4M7rwRsvbUwdrLgrP8I3PcBTsYFmW19x2h4CftWwspAKHDme1X2vkWx5dfCANhO0sz2xr
Mxjy96h78a+8TVP1UTIoteromR7mp3TdnGAwo2dIfLpqsmf2LaBm4LAwqDcd8hjHBEGUZtOSJAEt
/8Kxa3jBfRSG1snVVjWDVN+8T2nQnWhX5ltGf680fxyJcfI9haPBOqzfC/SOIeeFqH338i30zOV5
8nVcnhNIaQnwgNeCK4/lASAn0rKI9YQ998cPc9AY8ueNTgaJd+BfSYXKb0JzrQbZKUp5LNNq5boO
UPZXmca8r7YtcA4Wge4B9Hf/tE2EB+Xu8fKeiogbPsk2S7vIkF8sf4fdNh3N+MGaI7MB+h7QVEC+
EYuVGLIKu6hi+RU9CV+R+aSf7CC9a3krthP0tI0sNwlc6hpFNhhpiXxikTuQAMQ5jquoYL/Ri1Or
Ie64JdQl5klYeg+FJMLSe9tsFWoGcjiu/d1BHS8EcemeNCbUKqkqshp2va8fIeiK6dB/8GGMP6OU
SeQrXCH7XxY2mDoh6wHIp6El8urb54N3AT//SO9zEmVtSwITql64HSeqINIjOuPttWDBUperjGzP
hG2RvXwiyxfVbLLN+iLuZdEBZkKq4GS8p6Y+4wGvqzXKqkAZvj07DLLPUhlUitdvQC2IhTRbu0I6
XJhLZP6iuDK9P2AoAJLVLyOZY8d14gkXZkxVj1lBZ0oNv1zNLsocQzkOstxlb5xbeK7a9xe7C1Jf
lWv2/blr0gbXFpKgtMzDL8JYrW3BRLgWqmYxYJANGXHN2JHKM6+KN3U253IcvSHK/Z8Azg0XHeLS
HVIfCFtAfdIKf0+4CMVaOjoeGwPBNcNP2qIBbl2jyvmJmCPMtJoNBXAXX+WxeFv4eiBwdEhN/k1D
ozkHzyIClc5PL8i+r8/4TAi0Oyu8QJk8TVh7uC9oG8WnCW9WGdSlbmwWGvDHVORBOWqx8tQRgXMQ
wgegJgQDcRIABO8d3+ysOsOlvYP3vuNjZEnVnMTLZYLWyRhF/PmsEZZ0rVW3ncatM/CoUL2pBVv3
d79xZV+k5QPhcETvgUG3sukfzkHz4VkWLryza+gQnTUjDYUrCEWphL4itC28fYerbkQO9JXljYmO
KIniPLiDYaKwMlM/fW5xshSwLVCCYhiaSeRb25B2DG/Y0BbjRUmqdgfNsLbgdvf3BRWEd70q5hWb
B+VdMcbgibvscLOh3rOWZED3lvclEbRKxxh8IFIXMJjzDdo+LtIishJqOlMA5ULZrshltnUpVEay
TUnwCVyZcYTNOve+a7L9Ytj9MjgbyIjiGhJk+UwVcqsj8SQzOLBAKaw9rknV+HWWjEouWSpcVGJt
I7mgcX0vWzq7sMgFcKNDXXXqJrundVI5I1Kh3j87PR+ty2/3E9FdhY1G1pfaxFoYYQ7volAV+fZR
wFnJ1BE+Rirud/6CEi1JmINWpQegtjmbyySbWhKa7F8Vx2rxatw+OHJ13ZgMN5xZBsVVPgBnL6Lx
8/Hh/jdT1YcdLbzRthr/JJ7F0YDtikuvNrJHfkenHEpn9JDnNGHsdiqSqWGV0AT3VZkHoiP+hfBs
j+/k8ljWBvaV6Rqk9Y6V9ZN6yHlz96SNAS9oJzjemtFohLfPYQZPasBP9fcUGXBWw9k5L0glPU/c
riVXO1BA7r1t96dujwevJ7842eF10Jt6hex5iSa7oWzNavaG2y4RucfB6Zcj9WNeRdmY+61xHFcK
Y5yiX55WijrJWLtxBT3ql4hLiV8T+bh45NqmybIud5p/GcgNPNrAdhJclMZstWlqNUBUuBEhj0dO
5+IwdYMY07PPmd8tMa8eABI92gJEKpS1gaVycPyH0CEWwG6EoukFtn73SWyxjYR4eN7Ap3wkexWQ
rrP2zeH0eCuNhRGwbitB+pw7V+NxH4Vd5BUr68hySYF+7tTydHp96c5fHA9hKTwaPu1DhsZCqp2i
nBuhXxweUYJJ29OtOHY/v/oqzW4wZHn2BgRd/2c7fEbYOk9/mch6cU5kJexminfzxXjivgE6jQg/
b+JBrXAt1RE4XgNHlCuIn/iWlrkXZe0SG7m+5vSRNcRQo/I8J45JcFTmlyn2Y7LrVC1BzFj09S4z
uz5bVB67p3zex8XNS8RKjh5xhtVlhX/WVxcnzpPiq1lqrGG3s1NjD+cASACSa4phb5RuDBZBIM7V
LctDeBHuROAHUkWREO1Mwpew+JgX+bYEEVxawsQaq79GGIlXqPcEVd6MIs9x5U1n7p6rujeyxdEL
t7dnIwzVKQ2yL3t185VimdQ3FtxkKnTu9xjt6uWFbELGnPHczaet/AiCczOfHaC/f7oCRiz6yeR2
waYY0cXqfPs+vgJ9vOkevrfSiZoDPfsVnnmkQCKO9XEsr3lwo9pXHErPpnL7x2iC4SELGF3YNkES
Xq3c9d8uYeT9Vo9wJedDcnb2dsonid3tk/zeimnzAWjI/UuUlerGqRigKo+FkgJP1qPJNp9FehRm
bxt5kfdh8fDsJYqOGtqV0/YmX1Qimvrx+ZQ27SzsT6GLnjvLG+fYJahqm7E3kIOC0k6ArYQ1aHNI
LUppupOr035D7PqRbHOl+u3HEvhK9Zz6eb7tEgWh7NhyX4pX6LpKwwNI9IdxZRahx6QqSxjokEOj
VaizSHEzPuTXzAhqEtSxTOQM2/2ojfwW5AYKn/Ej7/LSYYvr6L+yL93slnOZAFKTK4r2uUgIXmkV
hixwgfufBb4p3HWyA44LvEsefJ6dk/+g6qXk+qDB3rVnijdK7Yl2eGU/FfSl8eJu1+Ekyy20C2Y2
Bb0aUdaUreJG8V8DI70SM81501TUQ7b7CYP70z8OsNrulk1a+4cypBjA7QIz1pT4o1SNyfd9HaQO
Mty9Y3ITtYl4XjqPjsPZFHtsR3A2X3M5ogO3njx+lG9AeSY564kjKVWARqsDYIUi9XCbO1Sv7mm/
QVD8fhBvYfy3JhtvwPY9pkv+/Alk0B5fO4vgrqGzYdiRv3MQoVLjxOb9gVdxMMYHYfoEFH+e5iMZ
MaxGUxQs9I4lYZIYejBW8oTIyfqYZy2E7ISsZS7V/0/UKwSZ4vw683N3RC6UxJHuS3eyuZCnL+U+
t1CS5yMpY9EoFUX2i3iScwqkc8LJ6afO33x5JTwOQmVu036KDrFIvZpGGrqCj1BCWhZKSMrOH7Mi
tbq0CSLAdXs3zKcptUfnockTEHrK/pM1QDXEd2Wi+xAuUT5Wn98TUdJqqsyrnDLQuN0as+2cyo2Z
fq+038cJ+j+TptH7fnpfqF50BX1mnaUimZ7jmWsjfpc22jncG1D8Tg9OrgpOEKw7NXV/qU1N0Uz7
Hhuau0dtEufP2kzXgdOgUIZ665vJOvYNM4j74aPP68/5XfwtSoFaqZIPlT/HQ6MnY3WjPeGdL3SL
Pg3gDCVfZohgZ9tHMaXTSyZ7OKDHnOBAMlSQwiAwR5TNlHH7oHak9YLz6k5bzS0/xSg6ciods+/H
KShwktbMXPKRce6IFr1sO/na1PIsoVvjQooXElv6L5Mmc45F1Exh9P78gYCnr07ChDjW31UXeAkN
Jq5CheAkMqJokUtAuak0tYnXTvsYRdIbiGeNAaugOMCRdhebv7eQ6irdQwY7K0djAIvzH5EQjITZ
sBGwH3Nnckpz6w6CSdL7EUjg7igOd8iRx52T7JADCp4FdDtFBvQ43jLPJZIuP2yzpGoItQFpfCqH
U0QqyvKxCUiuQKL6tA3ygbGnqqbRLlu47nZ71IoqztkZi4N7QYrWu3ZVr1HwEd/1iljYsqa0ouQZ
V8Ifn7N/mbXzbO4Lwd39+V5wa6AFgdeNnIbuwlSWe9+gKBOIZEX9gM+D8oF+gDIx2YGlGtaweI3d
+wv1t5WLtRwtjr0aS92mOlDqSAyi/85Poy7/L5cO6rgwoPYBT+SDG2ZsHUMICxdmQYSTB8FG8iiO
jw72gB8Igm2kKHWT+Y/bF19DNrz/oonqsUM+IQQl8/NldXqLaLPaDfgxM+Y4YOsWRlAGJRF6rlN1
JCXPMS2mdSQcQSSB/vsSqvN5BmVQyJ1dQ71CnqZBxRNcgKJ2mHYE8KVN1XVKdrDUoFM6xEOMtR3Y
SnCGhoCuK/cXREY31+5wp3zytTExafV9IQXd2+EoQNa5aFaJd1jcDK9+Xwh1S265xnmU8B0QeC1w
wUl/3sb3xw5ir1McJPFRhLRfXNgPiSHARsjpGZRmHsf0cKw15nEFNJBcw/nIwbYbubE1NvKAsLlN
4SZY4BSbsQ/xUTQAkNFyQ5U1dDuw4wBYzr0nksD59HqGTG6RPvb14teqYOTWyMMMRUvMRGLSOE6o
OuOKk0Z9V1SlT/NE8m7FrkZk1YjlYuf0Odi4c9n2K0jnMzUE2cqLuPHnEDvvO1eF++MEpyuGbB5J
/48vvY94WUwk6F1Z2VCl08dswhuwNLWRFffSecaaw+Ba6FHezd0LsMDmoc/PugXx8Bdu0Oyce1ST
UgrUJ4Dz+G/3/w/d2ycnrsux7KsIMaMbh9CvBZW+vfqSJXdihbZHFHQE8jmylmGVqSM2ToKTULwM
vAFLgj1YXXvSeQkPalyB9fLCxvc7ULaKaWiCWZGMjN4U4j/VYr1q6pTfEMFjosCIKfG800e88Gpv
BNfGiAijKDInGNJYZwxwrsY4FDj/SkOB3qRHxHLT5EJMIHwWCxaThWpllFoVHZ/DRYhkjjQAky8n
77MsVX/2Vhk5VHMeSP95pynZjbqJXfm2pyA/F4cZHGv/GhQb+hzi+cUoOSHWNUbleityjsGSDICY
HlxwDRp5supW8J0vscUfv87lAz2/lmLWRg7mdE1woIIw5iok8va3wR/LerJIG7/oYXBIsp1tEr04
Yb3J+EvzcadyJOBYA1bofiaDe3xV5jt4UlMJndeNQhBFUcKZbZOHCDbIfhEkcO7NjrEauth03zxo
a3oN8rc6CEajQlL3JeAOay7jwCovoIri7Gynds1rGqQQBWNHwJodqqYefObcchoS/CgB6uB/D3Dj
gGv5CY7YwXQRA+9n6TyACevCKZRAyV44RerV5PZoWokFEHFN96pR4QM5V1SKoi8X+opHDTAPK15M
koiMCaUYK65n7NXLXhw+XgXPT6VYeGq/gEYDNL8IYxY3cM5y4xnBK6Kc+UiYmgG/jf1ZVlTgJu04
qpE0vs6jhuC2kag3lMP9WnaRhyInOUJ5+gTikYMYfph9M+9cKxnpFj675II82z6k/jhVakYzwuij
g+FZKliFHBepOif6zhrEgpeezQuCFDFtDyPeANtLUkNpxT2/R1dUCB8pWIBHT0+vG/PX0N29xvVk
hKCMdhfgx1gjsuWFN2YRUeCUNyKORZBsfsJTUsw0VtB6cDLssz+Da5SK/26TCpvSu6s1kC1m3EBt
Ef4CZgoa+NprOidLE3Qe2FJX0vEhAaS3F8Gf3Uye+XLqoPLQ14L1jfvaTukUeT2DvtnYRxyG/6kV
c24c58V2FF+iP3/+JUcwa90DE7ZYaMRyt1GK2fXtEZ0coqNwtJMhUClVwsTfYcblOn3RIqu32Yo9
XsyZGgEUccltCda3oa1I1TNuWfpExBRI2tak4lpakBktkp9GB87zhLaOV4Kx+Ko7Fwgs4cKa4GhX
9CPQcyianFIkfwY1hzgIfVrPcVOJM+KkDMwwCSNU6ZJYhpH4mRjZVIs4E5Ux5k+lbqzgvsl3cHe9
AGdStOKQrtxerX0HvHawJ0JLWuAhxrRSiE1sB2kdqV0V9rPiQ+cYYp6uM3LlSo1e2tKB2toqIBbn
O+4DFTR89CMRBP7vBygVq2sFW4H0XsjD66btVu8wY5heR7yEP1IpLiiYc7RBI8c3pON0I3db+l4z
gKrU18tMRyAi6mmvuiG0Y5gYe3y9HWNOucSugVxviEx5g0O94BTEmeQY85sa92KKZPUzXrWHomvz
VvYBWcedh+AyDKZ6VmBCMIrhOEnlMhVm/e0Hs35MyghKoh7XO6ECzTmVay0paP+0eA3bUeW9yB3A
1HHyjz5mnJEfabHTDBIQDzZR+YradugwufcBv0MyRZ2Dzyla9Ks9amCLVTisC6lE3uBivB8g9ir2
UpfQ9vU4qOUt0sz3egWUxw28IySRI7ycv+fB6zi+jlMIHwK9HB6NEkDy80cq89bLsiLxTRA4uYI4
Xekkycc9Dm/n856y5F/NzoraxbfK/cRsPt8ycIcdM46aCb9EQL/d1f2Clo4LEhdJLYIGHY+x5dGO
U43YOOIYT4hYWZhvcRyHJW+KoU3a4EMrQf+z26vHSkk7lDGoLOs8Xthas/RWVOxvYeOFdx0F3mEa
buw2LVaerTbg2Roxw5zC80oGt5VyDhCu3dAwowiYLP5VZqQKmg8GzGa+gdsxhzl1n0aUDWwm3JSR
OuXMBSG5Xv0rOaAj3+7Va8B0xbiUsc8DcLeTTxKebwB7LvPzE/F7tsthsGSWlrRFnTbPKBXHGKjj
Bq+7Mx0DfHWcJU342TL9jP8/ol7mENYz7OdS1gq7iajZooy40uu92UXPBQCsSMFa1VjM57Ie8Ljb
ea/tbQntvEPdsnqfITn7d8JkUYkJkFc0bu5TOjsZHIjDK+WO/EmHyaf9rF2iRr072D/bK53XuVJS
agSguymXsmzGviu+HYSZDm1+qy0yeua1pAva7P4eduxJenv7/1qpIF4Y3GC9R9WLAOcnLMQQYZGZ
4FPfwfVSQUb3tl0c9e8rAfRbzRJG5DVLvb+yQ94AL+eqP9EWODo9/FJFlLKYK25eKUdxXcDQ9Kwe
2MjlQUhahaAcmS5+FFwvSv3uUaRhe5DhXrJmUosHZP/ipPdC0AYUdPAYBlXG6vrEl8YSpWAOe3Ay
LMALN81vdGo9HZvR5ubfTw51vJVggWF5ZCjfy26FZ73GEqB7jYK6bhHD8XIjS/3U9VoqEmJylux0
BjhzsSbVgT5N718pDi7lW+wLA79FmQrrxIHs1NEhk1XqzFMv9YGBI9l72KtD297jsVI02c+w+vmF
XppoLepqXnnU+RcBv8dNaZtNLU+wnL6ArJtUCZR9hrirwAf+dNJjjTIUXHvooTmaH32zlFR4vuJV
2vz4e96Z195+zCTRZm3mDUx9M5ORPgwdWRQnXdNHnuJxHo3j65K/UVmIxEmLG/oMeE197DbaUTB/
fU9GkT9A16qF+Ocrtxj+9HFZXQQ4SN4w703sGz9gQGCOHQ8WCLdxQuEJZgaOvKpWiD7PNzqmXpcS
CWF8pphrEznZR9JtnJfIYnXs0jzjiZQOGbjmIlJOzx8Elnq23mWYC3zo3/GGFzkACDbM1SgszqTe
o2R8bFKSfJmQhUBWgKHxvT8K8XdFsy9R9mgSPIVyqvrv7rKgb0Uk9zMUoawlRKg2W8nXid8aqLn9
CpCSXMP8mP5h7G8SXFoVH+BDQIJI7tlAbG5ZHAy/0McmZXDmXw1bS3+RToeNz8Be2NwGEuHYbg0N
/1heKpTwqxpfuUMZMzbclNRn1ir5/hTCsT0lyUgcFu6dcvhAeQv7SIQcab0TrkI6Fd+hHENNt5k4
6kQPJggdyRCYZTj40bVPvU3f/p9cTglCVUU+WyOTgu6f5QyNkrm4fUscNCUjAr1xTdIV0sMCMbU4
jmVDY6urfy1EfCS2nWd+baGFSwUbs4jqmLDxbAQGeoPsLlGLDcnGb5wqXYhgUSEex9eI0vN2Jl7V
tuw/Q9eAhWG+lY1ssh9j8lnhiyYB/5TajtrciVTuPKg2SG6P3xsyXoESqvDYVcjyZJ3touYHz0PE
URmAxXrt3TVTfepMh0+aCVADZNxfGzzblTA7LWHal/3R97ahg/NO+AlPgVbqoSBmayhIXZed+NBu
CGaM1ip6Th2S/WQmxQF/vtSlTEe2UUI3lkAIpN7czAsx/hWrld4cMhfOJNgVPaZo9Fq91SUdhT/k
bBt0k4MBIgqffF8AparbMuNY6H69TyYW84tRtpygTEFLLwa+ESK7B+AMGXrH5cfcnegnzImPSwF4
1Vrf7mQpWFI1UbCoTgcwyh06dyriTZ2k5OzGeTm3rIxUq2GEEXZWW1JrpHWthVnq7hVxdyNjaZ1A
GSqJdlDNTpq+ACeSGQMaTWCbMHBDY/kYMX/izyVXqBqxb4DXP9M5j0hgI8sjZR3vnPLGo+yawcjl
OYNF6UZboRPakDzIhtdMxawSE/sWiq61OjLN+SqCSOd3Pfgvd6noTL+U52UGw6FQuJt/m1M6MfVt
YG+EVn3a5yQfbmHKB10aq/gubM0eu7wMWEXbM+OM/W/YWso+7ryL6djqniXwHDjXxd50iFib3nNv
1h1W8/OEq1Odbj34gCcvAtKx6p7LUG0LmsADrV81t9D4tKK0p/nzEJajOHZS7CvSG1gTU7sZITls
qKEEtWqzb4HvaCMLtdo0MNgluLo9tez9v83wVAiNLGEohl1VGZFoaNzmuILrDtPqCpocf9xic+2A
I4SUonaS/stTS6a0uyl239T5SoSZ2ALebOM1CEd1O094igd5ToZZ6+jsOuP0Qrlrs1jlskY88RhK
gM+sNYpkBGw/3W8PCM3jqJIHvfNL5DcuGD96R3iqYnzoURhjdYbFAO82vUZHpOibk52hCxlfs6PJ
EfS0dhsylWkozRU4axH+TnZq64lq0xgViTR1EaPU/RBY3bNcUff38+KLITSsZC673SG946ft5Uar
B2qtgiA8r4zYn3O7xwNHpbFY9DtU+/XYhTF01IzUr/1YKHLyae8m4+5riwWga+6RMIH8dBMdevrJ
CQsewwIs5Biq7PVR2rM6Ns2/MZn2E46P4zmsk3cWyh5SzZvW3SZlg6kyhaQaDXlM6byJKwVJdJxe
y8fluC8f6BqXXbzsiMX63A9FNwBpcw0yJ8nYeOS8rTbQyEmRvsfi28bWNhPSRVq3ALJYlOk3D2OT
ejk692afpc703RGjUCqmkszAIxBPnYXa3ozBKQ9mpYYqPWtzFdMfthSjPMOFcpeyENIaJx71x0L4
CLM2MpeTpxIwosX96NLMXqjOUCbGw4WUdOMl940FIChkagkst8HTUPUl3r84c6kwuWjHfdAOmLqM
BBAhOOotEAcb17DsVtXqdxMIDbBEftPHKXNNbAOt9QV/ybzH0wcJj9ygJ5v9KXoqcHEOYYkR0p0O
Rc0Q62OCHi6xOreAeW3ahH0HEjDU9DYlZHuo3iFlC0kUh40pYkfyctahES1DrfSUs+F6FsMWZ60Z
iujrLJrZA67vi+xanqK4wDr50K6iKzw1tSf9vtqRQJEWWN2Qxu/auZzPa+oejkXiG+/JsY0U5fpy
F48Mal60A6pGd9oeUuId4QI3YAJ9swhsHzDYaNFNAUOvtRowtJkRmcJmkF3F9sNQOzrZ1vPZO3Oq
Po1z7rkdKuCq9tc31Fx5dtlb8jwORLIumm7F7abKZqyZUimdq9WZXdcOInORNq3S8Yvqb3YxqeI+
T6nE6drRcMmvROFGR8UjCNv9GVGhUB0JtilEsGCqo7OLIweUIxhMAaS25yPWlLkG866K0YbyxfEm
VI8RQJa5Sjr7JGxEHuhUvAcuwohY8IpF92HSp/3WzDTmP05q33V5XmeKGbD6LMQBAtJ0zxPZlKUv
8EL9AI3SJqkQzGYoIzeJuFsThG4UHDSUK1l9IoxcTZf8dLOPG+x/cizMoF4XuXiinvSNPBMOfk+v
EM3NMH8FwhuGvir2+BUG7bunRdsA7zXL1ol4G0kIhyBNqfdpi6n1Ygog9bpu0GJuFzrPU0ppbFmH
+1Yfl0EFi55APLny6mACW/G1I+NDl1dpWw6wf5rmw1L0PXTrXDMa625jfqz7pyJsVEIQY6+54IQV
aFtnECZ9OMMNF8wFkzr751ptlZxu7ImvvbFrzugNTND4qcwOPYESVesAFGMhPWkmhC5vbdM/4YPE
iUwWbTELo7hDVn0x/YedlQzA5ef5Ty43PiVvNnRLyIPzA3/B9WzQXtmtS4wIezU+LT4tF5vd6Y33
Qs0o6n5iCozYzOFy6h4D+ej6vQzn0YHNJHydM53+V7+SbX3f8tuLdacKvRvsZxlp9jVYgrrGy1Az
pcUnXaEshbFQvrWiS5Qeb1Fdf7jdu9Xakd8Q6saWlkYvyNE+615D4o3hvIMY5eD5FENcCdZdy4W4
WRkjLItE2br0y6Xdhd2RLu7S8GWnXZjVaMKBt1iAYMI/nQFn7t6QQ91ANo0toW3Uo2O2ykXV0BNS
A2CwJl7Umc++/q+wMAxDWqqOdMPRuIKV6o/yEgnXpnt5R9+PKFCJXn2comnwcldXUeYZYO0651PZ
OPZcwiJG3hx9V20mkDV3azKQ6rXWZ+UvoJRPhw8CfC+ryw61joUILtpRVhDYiY4HW4QjY3HO3ku3
nZJhw/AeL+BiETQz8An0Zo+iN7jYh22VtzjyFe2yEA5axMllZraE11cKv+UiaRThDZVaPD/tcCx7
RbLg+JoZ8LD8Zij8EwY8JKYVkG/+usCLiNqrMd3UfbpO1EVosR4oqkwfioViWoS29wIhNVLftQxm
IYLacPDmmD0PXl1mNT8s4bukiq1h6bVj2KscCN8rDMAauoAUTURke8zdbSgbEQcWx9DBa9UH4IAd
yyeSb0CvRKbuGtyKJ5kRjvmedvqLGblwPZ6wKyxdksQrQEXDkdTUOmAjADIwLqDzDRtD8SqBiYjK
JAYwsZf2L/vyMY9qSkF9pFiBQd+IHSvfdAPKbpdOfczPm1bqVfmCNXgjzVDjNFsm9m0DiBDbnmFE
njQ2YeBjTyfj9Me5bPaN2p/1Lgz9Xc6x5d3XmcgDVe5Qab1s6gXUxxpr4bekKp9p70ihd+Hu0LQU
lBSnxZt3C0zbeUuJhCNyqLqm0/EBPcQPvTi5aTp++BwLyNtGW7IsZV1osnT+i3g11X4KgpQGR7HY
CyDTbMTs+IsuW8R9JEl94jt/Qy4emSurjgfeYLk2OiWxQIgJwSQkw6Zwen5ZjHtgv2GiMwVPQCOU
jydi6fUBDyWMynScMAUuNST+K/SLYWf/YetsAFWfHIomJs13fUTblQNluHgNO2pF3J3bsqZsAZMR
os085B4YraX/rsyCRYWxH/6wUhYrMVFdJ7GYz+76i/A1+RC9Q9r9PiGwrwIUYEXidNIsKvAyLnbY
QGZUwxUL3zMt9Mb4yHhQ14rq01BATkTt/F2P8ZHeF/KRQxJsFf1Y30Dm4oO7rIizTr+wCo8ofQqa
2aPrvn5jRjuX62mfArr7X8UaPBscakpK+7Mp13et4vfzNexjrkyL6+dEu7xZypcs0OkyxeKDOjNY
0uIodHOYkM3wchYE1Z2ZcLaKhKJfZSpJMWvQYYE8wyPVV5KTrIoTQM+BwHC6VCrXxgjq5ORKBlZA
mlUH/aqwmfm3O9B9SDMRnvsjNrd4TsJl7UAuZfK1St241ASm6PHYebtfwyPSNRzbGSTVVi6+ORjF
N72muGShUkdReqdlOS1CLI7Herhp6zK/e80ff2ntwmlcO36grjz0dda4c0bs9xcr3ooSCnjUo5XY
dkGNvT6rq30UAKkYCWxIvbQqAeokceq/HR5TQ9gBFLj2n5ZZJcLMYZwtN9ncjwdRDzaynPWz1O7n
onSgFq8C8ZsBQCllQAvq50VH5eMso0/3sDM5wv7eiKh89yYomWiAmyP+WTcbakY+EUYIAbbFH1Zg
wmyU9S0u/MaadugL5XJW3a88Y5Q0EEFB0LAp1ZG9FCH9RXOfC5bCzOeG8nGusTFKHqFAvAU2wyMz
WWqt/JlS4QLyjHUuUu1rMDQKgnbXLY893Xf7Z/aAMTvMJLEGBB2NrcRqGI0Ye/vkrALcouFBczJj
IzadiZv7bEOLkAg+kacpNTBBC5lSZu4R6HEuJgfa8fxE1VTANbPSRXhRbTGMRo91GSzMfjvD1oNa
PAkcXsdAv7Yy3RzzzUl3fSSwI7lVpY+Q7yC7Jf8QdbfQw/EfUH9tgWP2vna9IatEbdjJIL9Ntg9+
FRvd7jYBf/sIscD2+xOi0KiiRcxkw5bHSXpWaIogwIS4a3PKc43wY/RTkFWh0DBCWoU/LCiYWrca
60DfjD/Q0ZRQid+AzAHPGzpIEKiFdZMihCI1+aYUW1zGIELH/FTaIvjhWDOmH+iePGhIyYgD/L1L
o4Pvcd4SAWVXi4PD9VVZwWhoc2+O5mZjMPg6+nvjFlzKTOwzLfb5Yil9GgmubSD400G4zLdydE64
xlDuFVRSjXpigJdQ01aaA3dpXusKt32FRYLFXWZ+v3sKQgqajrD/lQJIhT+ugIDPysgnQBmix2BH
W8ngUhC4jA3hBMcNLFOPUgg2ZXNhabcvuz8Oy4yuzCcT4tYfIINDuKRK92Rv8+7P2okU4vGY2RL8
ElMHVP3nj8rgw2kajjLSBc0NdZyfbqoBFO6Rsf5RS7V8dQ5C9/7fCUtHX5ZDZKlyoDaD/MB66gBx
JxXGBuiFwyyz+zWpLgZae9pNeBHcZjdVK2h8D6d4bkr2pKJQj/Nl0QiOwZ7xN00ot0tttWymUqhs
viykv5/C4WxP8aIFGvwmidZ2gelijGvEfrWtMuRYdYT8E2lCn5gh6FKtruLFI8qy9MtHyBsJWCl5
ictaH0JXwF6hrovaZTyxuHVwuIbp073HNG95TdVAkdxN7js55Zohj5Bg/JfYe3HepC2bw0PPZIOu
9uepuLxvHEl/y+KmjkNa980g1WxsBbcN0CI553BNYr4fPfJLsV76lKVxz+s3tk80GPP/PDKoCYIP
Y8rPkE7yxX64VuseNo+4FhmLnaTffgIem3x1m8loLBpOHkZP2KL0xI8C2TEEyvL6lMD13C0PbPUf
XRjuTuG9CQtcy2u9pv98FKyJ/Qf3520f1mBbGZLdX0SLY7AtreI05BPNBF6oxyQ8yhvRufWElewQ
QnAVYetYUr3+AdndmWi6zmNO219gBnI3DSbBOKeNJlRYVOpiZDObN4qrRtBESeAmHNR8D6Hsdyxq
3BOCVhAoM9NnSR+3t6azAJQqabNyQyNl/wmV2Qua1mKnIdOiwOyhTe8tQM/bABg2D5mFcKz5QvPv
CZlhy5XbRmomAeAcyCnzpcGrL/MMtBcXeaYaaBdZXb9lGj88lpoPP/+pcsNCDrwbMpbfJIByBGFw
fL/EpOG21uTtPHBdf17iSiz+jHklOcy5CzbX95SBp57xBtMzUwEw1dNxOnpq3AYkoazRfQvWz+QR
15l9vsZP2X+Nm1TejZ3KzFc/oakvSdb7aSaMvrOUGJuhT4J6vE486d7KYue0/Phpm497ftv7YGzv
u30OL3fbENbIP7jsYZ/e9ezlB29MvHF28VU5R7Lw2ymS0C6GUdRlnfNvbfnHbKwzIvYcDCpaMtDq
kfOsf/l5uMkmtBW6cKweOZxUBWI7998PphZmGbNRfzcP3Bx7gQVgCX/M2BUGa7iOvT6cPNkhQtT8
8Jw/UCjdffEw8DoZywfSfsfxPyWu7Sf7nsD2XReMDTEMqggn6soAVRXXadIrpiSq6IyaMIj5duoi
jLyTkMga1FRzdQv/khUk7S2oqYRGqmaLIYsHtQ9puXKgr3/5RotMI4LQr0MVzxAPBag86V7G6jfg
7A+pBQnT2gQdLGiRiIwfeYwYQoseF4uc/oRtyMjVnFPAseNZMaTVKM3AyJBI80FWsAb3F5dlW3wx
1wb+0zHKzqeOEEUcR/7DnxVzbhhQ98FA8zRmfLf4DGhLJWqEtgVHrH9MMLcP4V/+4Zw1vEUoqWKX
Ceww389iBjJHl3FK1vOrvL8Vnrn1/IYVDBVKMqoq5PtM3EHfx4nFoKEEI0MeGPj1U8cMinLJsjwT
HK4ihTf7MxYTlkdUPFfYHHTZiOhD2oyG5vwGiimaZCSjRpCVThTlvXVn1HtVvPLUA007kA2U/KMB
9i4cUyYJaU3aUqyUf7NRjtth7rbLnqzeNuV/P5gln3RlrJ/fBe3k98xAlP78PKixq+9/mJaK25Vt
8bOg86iXvcTc7OZ45xlXv2U2/ZQ7Nw+l+cmmXhB1uqbtS5q6egm5b34WnVafgEUI57vjwqlmGCYe
D9rLRHHL7IxN6NwEL5Z+NifqJQz/wj8IdxXISIoL+HVal/xpmGbB0wWJVmr7W+j9yPDmaXfCf9dJ
cymD+Z6yRGUoi/d2D5tkoeYfQMmYtcqqfO/+KpbdL0Lngkr9riVFfyNMz23Pg0/vLHsgPegs2YmS
UZp6rk56C6ZsmRC6t8wuC3lSzoR2NCObi2V/BkQ41nbsUwr42Vi9fUyndIElxnSNjS2YqGy0vlZj
lwRxv6m3vtHbms9cmo0iUZS2yTCd3Tf2z6zd+hG4Z/H1bGC9Zu/XRVSUY6s1dKAmmuvjzPMOmkMp
9a5FJE6MxUAUbKCc8hh+dq2inXyv33dV8s4hpLT66hOpatgREV6RtuG9i0K68FDRu+yoRBA1Ck3C
t1DRxWH/4p+2uYAdSQxdu+/dOgYIqwdP18mOkVDp8mttixT7/YmdJADaoGZyzA2GqPp8fydLPlDT
jf5kxGAzVlaP4uID6EO+k/c+mIX0lRBEmFUzkr0fJ13WouxtCKhF6LwiVlDNqr2C4JHhNEuSH3ik
tOKw+7+qutuFZvnWq5UixbqvNV3cdoa281HJUu/3dFxIgRHsGbAOAm0sOf0iABEe4y4ZTraKzjcS
m0tMRUchB9HXcWKGcwiHYERJ5D4WOH3Nf6NRqcFM4CNnjGKl8GhBxL9a76ogn6RkWbUgV7d+VSAm
drna+SFMnkWT3SqY55vddtsmoz1+anbIlSpDaaIbRYFtLD2OwgwL1BldulqdbmlL7ZsIptTqwPDH
T6ZbMqr+VXQG5ugsKLxuXZnXg+38y81PvPWaZfaBlgeLPwScg9Bur277bqsJgYx+q3JrqwJiwK1G
IpVrAQpAx43R/65d73ZzArhAimN8R2JvtdQsL++AY8hTeBkmbd5HQevkky25ZoAYY2rXem96TJpk
yWlgZYjHHqorL0kphTSyGKFeIq3G/xXT7VLab0LjOggSC8yCH0IpfeYsL3UtBnlDXILbaKoM/4Zd
f1UsD5KyE6oHvKSpPSpKLEB5gzK311erf7CWJB8jnhifG1ifmeYJcYS2YBs85ARM4Olp15JGTNVt
Q+XLONj3Y0Mb3pN0CWjR2bXu1qsRjnR6SPvBpf/8ehhpTb860iGeu87kj9XHV9sBCM0mKM0cq8Nc
Xl92H+m4hAhX7TEA7em22xH4MmdY0BsVd9fv/zKP9SsvALiRw/PrgmQzftpc+U2LzxMG04ljWafz
R2Ese3evRf7fwURYeMEaY6FhbDsrSbvLxOyQFqLWBpc8L774ds84CFFTWAPsqYV1DvW9afMh7h6/
+qIfis3AFv2mPbKQItc5thvHB5ozzP7zf1Ze52Fz7zjMtt76j9hjwzIovhBDcLdHcsycvvVTJwPB
IMHaL7Nsx5/P/Qu6tqL1w4k7xbpu3CCRyhosW4DnkINdCHgt6bj7sxGz7Iyt41oyDMrRyr+5zocN
gdz8n1WIA5zczhqtZ526TvsKIBNrRQP8V+Klh4sFcV+igtMWvPLmmKFQ5jRbdenbXCITKUHrbVsR
jD+4BpHOMjTWoXd8+Afu4pG7NjbjbaymGB/OPY9bCeNls3DQAE3j+nWJfYRuKj52MquCrSCRP2DV
eGq7ssJLVxhi0l5r2b0AljIVcRwWSuWvmQxf5r6rPQpZaA+gGbqJlz/u9dzBehApah9eCkPIGYL6
DuCLZIBn0J0V5R0vbwtEet7jq0ow3PmhoO7hiMvMv/FZgQGTLC+LnrsYqwM1KnTgHB8EYNTYH+vB
mRjn5/A+IC/KvYnC7BjvyRjwtmqRZBZGdjmhDw50JR2kTeLDu8PZ49WXcKWz2YUAndTBsuCmuyXf
bYUFHswPu5goZLob244E1sU44G7SqtJ06+vzRGpoJF76FVBPQ5J7xWkCtaN5Dvz0C4S23DWX123G
gQ1DWk68GdwSKnngY5ROBBolDJR4N44nsMBGB04pdvjguczaJOhisn6rKdJaCjdSV+WnUFur7S0D
VDA1Z+z+igM8FHIKaBviGwOIBx0GhU0Sj6x3Wsg90sWK681o51tPBQ8NnBK/y2NzAhA8xeYyWjxZ
vTintTeFLl6ITFBWxDxAudWYpGJ7tqhONxXg6njZfnN4HTT1hzk8j89n14Whp3iTNcsjq0Nj843n
BIz5QcZblfIJAabxNGyuxiojSzqpfuNRYcc5dguUCl+2jgdomL0KWmoIKM2nrDP6aAkWYujMllrP
tOnWrnK8fOKYGusILqMXQYHrwiQcq3iweIp7zLzTP0/WGqg0WWYe+jmN4+G+AxzrSRkoKKMTCWKv
irGOryakTImr86LKBgml2x1aI57s645iZCXJOPG5mTiyFYYpMH3tVxgESLOPTzxeXGaqMfUZcT8J
2h5F8qnQxfUXZ8YksWXMHwdXhevwhRQ8+hEEXcjkpxGKFrBzG1J43/RosJ4b/AeyDQEW2MqHWIef
GKbzDwCJihz9wPq7LtG+LwOLy7JAcW8HjggipAvxa4Pjw8yI8q7Qgx0Ic3bxqtIkDywuCBZ8sOnO
+V0QmVAJCvNHsgFBuEDo5BexH9acQAzI8tcehjKf2bkiVXmHUVZRQDDSWcXO4N1woFHKK8A5h2Wx
i8BSX4aM3q+fz0adpVEnxPbIKBZH3QaTuXbENTyLo7Zb7Tj9PDGWYaGFUcNSlX5DEZie5klbUz6G
itlpaIuynPftYTujbL/uQKa2SAEcbefVKM536peV9B8Yf66HHpnZbKkS7T6MHEvk7x5n9AyxHewM
HpVCWIeH7ZGU6ZHEDqsC/QXb05Rzb1aXZEptBlVQXPsIr2PfFwK1xTeLbGCtNrGoyECJcVFF2c9G
qz+F5VljizwB4WKJTP/dPd+hWjsoAeMW/4ZPo0uqNIOXZO4OoMoEtSWyiI3LndXnJIlNqiU8Ka5N
B0uP1DUPDNRBKxbY+KEQZ7e8tNGNzo3Ej+HchNfkV0mjPeu7WwSPkRNkqRz8lxjq/RsuQwru2gTY
SG/1u7Y/02uKo6Ait5K7dw3bKLIzYbk+u4KPBygeT7VqJ5okhBygkpAWaKMcRIoaMoGUSNJMa0qk
gjVUzihU4ieszbaNprGL3vujQ8lYRIaJL1fz8grxtlVj0zGDSdYTh2f+ad6DJG2Tj/qRCFvRqDR7
2QL+pesSjLEJfU1xLmT5A3cT2BtCwdRmUry4gqMi9WQp7Z7g4uM27MtCdZxd3ykmxKSjKJf6EI6k
WQHZxkfuPt9nZpB45J2X62lH/b2La44NB9eU2uQmi060xtXUK9LOkeO3XYHV3ER9hl2ns3n76US3
ba8ii1mmwnYYxE+K/JsVafoJ2RzC/4CHvQJQRQXY6XhvkLPzz77wQ9es299AI4u8pv0tEj0FQ0iq
Msq955Bbi9eo+F8bZRTFzn4p5ip+UTnvCQ5bUWbUqLcHFtO9SKSb1vzqLYrsIkg+uDGcKstLPL+9
XjCNcC9sp8GdqjTu3mxg3cEQVNwbFDXgBYdBT1T86VzYA2sgjtu79t39v7Nk67TI3Wqd9kIWRums
MgxCJVb54hqyeQ8MEqrJV3P8bkbsTnrtPOcA5OJ/syDbelwJC9bLbWo3F+69A6kI/MEQw9hwYelD
6hXub9SBlexLHIJ90RqUI39fT2JS/iZAZ/XiMDBETt0xTt6Cc+lljQ8pYXVzfVeh9flg1XUhYtHn
4R/kuwN92vT8N1XtdTa6uJgzsHOWNBwCdCuGZnfTG7Od+xu17CT+iGpsHvtXqk3m8ChOAQTwzY8a
kAuf3E/jPTNrQ3ni8j/O4khdNZnAVy501XjeyQpk+djatEMmd53Kij5hdCZQFg1mkrMyYcMDFmcT
kcAGkaC6Ujhah5mBEeKDPxJRk3Pstb0cAvEz+2cUOYf4D697hwlrPm4I+X8PuePSBKkjoDqf6+85
fJBBxSShMN/w2gZRv8Ru1bM7Eo1b6Po487uNSH562N3QEoVlw13uEQw/Q5DoS0QXOSvld1lbOr3U
DIF/PyLHSQYQ7mP90pDownV70FtK6+k6Hc7iWUIutnWuozwhkSdUHCFRL+e1BpDzpRznSwTs3Qtn
yxX62S7cchfRkMzCnQhGGXtv071eByZaLyWImS5HWNLpfy9Ic1hmqM2o6l+EbSUddhoM4VLoYEeH
elujHtrAu1bGiwdQiK6lV3i3BbGC6ZBmlKzl17TPzSoY/c1x2OKVHUNRnIOcSpQ7HcIpPt/LzhP5
vI7vZQatMZf1wuoq4shFxcgVLKzzejHMipKyX6AlRCp7wi3fUOoDd5kTNMSpRzt/W+MX5q55X8tI
4HqDpwbWf4tdhtMRfoiKp3xaWHuABnyvvSCfBP1k2Kvwtquo5U7zXii1fwHfYQst7Bpi4YK/jcIU
e/BRSqLWDUIsg/VFA/Hqr17/UwGcv+xuzjwNHEtWorvRLoZb+5Bp2J27QbS3sS9qIDlqrt0rjF1L
OGMekn+4PuKeXx4CiHI5GcP/ytDJGf0/w/P+U9ujoi+3HHkAHvXNQHkcLYr4pkl9SDeui90D4ixb
cHvc4ViyXFdhLBEbHdhOg2hHjRKoXJmiJEqzKx6ri8dJ6iJoI2jmqXY9/P61SbIMP/Bw/8RjA4yR
ykBozJ//Fe9UNn+GP6mvntQ8CXfwQz/sC1W6qXsrIzixtz6AFrJhUu9Bwvy+taAr2CafDVBfGev4
6KFNc4EnXVH6zkE1T2hHxw6MWb9jiVGvLHdWrYL7ujbHWendPLm2OV3u+vE+DuHOQrxUSAnqH8YZ
c2nftBV0cJpFuiIk1PXb6quL4zc3t6xNNdRiLOhf/hMzeFisqp8yU65EdRYZEwiVc6QrqHBbpnyl
wcNBbxJCiDnvOAEfhkFLteJo12DVSOqG3/vwSlLdwkAxHqBCuVOQbi9gnYplNiK2tRAfPS1x+MTs
pTYSEfVaT4CB190NyFoU6CWJ2UxyNda6YnwEm0kVwng9iF/690bSDsFZm3BnHST+RQ9pW8W8xmXh
XAbHKUgTk9JxapG+ntsTmoS19LV/QtxcpijwsvwnsF838XZlXmaMciDUYBQZutc9jbtg7tEi/Vqz
QCAeZB8JHpoFna+8NlS2NcrqJc6+d9SZsKWkaU1N2PDn0WlIYB0CsALFGnmnZDo61X0dypfeNRvy
16ETJBLCNRUahAWxwPc2bFjdMNWPZ/vQJ/8uLhxYoIfZcJT1+YafoqgzV9UYwRowzIaDeojTROpV
DlSbPyKezCXC9FsnX2boEL8GyLzP6hUoLe87yQDe4ZDjlQ6NQLtHd5TuD2tooDz1b3HvBZkYYFZG
k53IlMlQzYcCfXBfbkx3aZQuhMi8bbulS0uczICSeLvK9Xp5XC8wGzYdzY7O7LPNPvh7wyOKWsfy
Hzqhs1dwfK245/DlaS9fAaGtdWFlAGXblnCQxle8B5K2QfQFyvfL5k1v3GxsdPz1yRQ4h/MIoUOQ
O1DO3xNPkQwrbth38vPmgC5aXc/k5qnRMeMFvIjLbm5Ld66L0jFXOBIwDYYZLD+qjJJIIIp26+v/
YjwjLIfUrrzQIwopqHTdAKcCNam/YCf+t3mXxgZYmB/ORWZrZzbYCTAXc4PCZL6fF23EOuW8r2Uh
9TwD/Y4dmPH1OmZBPHHnEa++TpzYwLiHD+fXXn/Jey8+9JvGTyfMc21q7sxzFJTYjHkPoNmcw6+A
GGxodAGamEIienZP74Rq+GahYJhwEpHlVrOX5tzpPWxpqU7iM7e3f6Rxvsu+/cs6sX37V4QnfdCB
TGSYpHkmCOsZHoMJ103qI/J5iMawcMF6QX29b94yI00Dn+CgHQYlg9i288+hrrjewQltry8yjxf9
6vzBuNenqyqOSp5CLj2mHM4nre3yfcpQFiFbOhl5atLVfkfau19cQ5QDRsbqrusZV8BXP72BG+zP
fElRq7WVkXEznFW657l5F5tpKptE+r5k5/mwi1KC8RgDi8gWY0Vium3DukaHDbNRhmTYSiaXIGMl
wQJ/CVI4i1U1HLiukKhIMtdWxi2QJIffSartNMeAtmFvqFHSSb1RK+S3OkL+0n+MqKoFF6D/WOtS
Q7EHHtWLR39CYHnM+tRrScolauMWenziQfNXb5GAAGKe+gmqq6t+YJVChmjkH7Qxo9Skwll4Z1I8
F/FNLH/jdVlH7dENWshtGfYGbBfmPr3eYXz1E69eHdZGCEZFELFQq725gflHBQn9ja/9rxm2/Y87
yRobvDlilbSu1Ygg8LWgcXtzLQslQ1SJjGC6gR32EzMxVikKfJeXQPuOvyDRSYgzzZZK5MIVch7D
gK8iipsN+8PeT0qsdTM92ZGDufGG1Dy0aa+/Y0wjBELxTR8T9U9zZsYiQ1vyHNClecWOb2n1IyTE
2yhLJIcraIwmBYPqA7N+cnCq8aVeCkOXy6t9XVuBtrO+LDWS5VuPpSUXkos8eXERhGTEBc3WzoeA
+fPTVz7kgOMXX3KDONKRBgIns/5lCBjDx/ZLYmPMQksYLCvfPdl+fnqwdflEbKGocBiqYxwmsd/+
w+5Nx1B38RWC0NAVh60IG7yZeiJn22Xzf6prxoyAVYHgoIFXF5stN0PQ5JuZC7iopfaztWEaMPLG
7a46Jj4ax/o8dmk46O4wtXUNPRVZPyvbHN9btFr4+wxjiMtwfF8J+Y8DuwecI0PnbOeXUQWSOlfu
6OU3IW6teog16hqm3kbBgLB0GXX26zGbwaKu16feogwHaTBNGg+n97N1LJqtUzrrbeOe92niyfht
4ibLvuluVt62S2PGF8PuDik3Jbvg+bE27x/4kZgMpaP45k+Xccdx4w2Kfd0HV/+M6vFk2nbFj8Zg
7FuMO7pNlnGCueCFotjMr8b6xfVSolP4Hl+c8DPYerxW3sGiqW9GYOTJSxwa9mJFyNYKINFocB5N
yltUOvstxSp2xMNdqBTBEQfeSweTvEzaIrd93rTDYpzgZc5DdrgPOUvl/uoTm3w0E/HxiRxzBzvi
6eYEbHDbBxXP8Pnpr16f0+OBNZUQieincMIQVfoaOfLYVEyuHB1bgF3mz5rHsa8YJ9v/6EKiAVkZ
T3UODPT785eBgTQwx2VHzJViYxOMvq8dz4X7w7A3BdLrg2hM1T1pmGNgO8MugbRO4szZMJCeBCXl
LZjYBI6Iex5avSf8J7QT3iFnsiBDmupbWshBoG9f4uqlSJTUmOotgWiepgWsyUv4QdeSub5uuEEF
utydP7qOuEky8M3VQAzco2Y+WO0Qwbam9gSOEt2QiElP+5qXp1xAvQfJvQKb9Qm0UgLETbcikFt6
LnUH3XQEch10mnlUMiCia5TgkDLgAKIgpy84pnY3+1izz95SXyCO9qbki4gfHrHE5cgud14hiGA+
honBgtAYGWI2iHrrePEL/wpo4JzW+aqvcGtmH/6w5989ICYKCfuDErV5pA8k5fYumiL5I3+VoaGV
hCTAGJHZWgSq78oW/4C4WznNhNSNqwphvb3sGl5s/aotHW6xyM3PDdRkcs6+hKGfuNJ6EqyeSZtX
B0vNb7UmkKWIsttCYZELxHQkKMgwbSoregQiLsR3lD6b7dFpmwLcJhiKeh04mvGGx1ieIqWEYPM+
j1WMFa/PvRrgLKjr8zuwGNDbBOoT8StcyVOBMAARyz/ksked8VC8di6vvhwnbDjPsMiF1xxlrV0v
4k8ZRzPc4MLJrYivBWnUWQsL92YDZh09gXYOJAblownPgdiWp1BWgxGRvxDedUYrCcfCCy03DjjV
HSry+LSc4ct/j5kgrOJJM0x90dsAxImklBJzKRzuIwjwqyZvw14gfVL6vLtKIRqU4hoZKA0JiDS4
lk8VQis8feq9SLjzGsa+FkLUfjROQfBokUmFW+k8VyeH8LE/ZQsM7gcQZfuwhD3Ds2zt3PPpwtYd
awbZadP2kNURLK+vtBnKF3BLqopErF2NTYKx/I2LM3JT15kyJD7TKVWyeNgsYr7VARYH/QABloSq
w9qfpuBCdbib8wXbRgJtGKenOsf95BoyFsOqM0UNq7xczMpe6INCo8fluixlhIhAd+I404Whf7zt
fX8rDf9a5hNHdENqJvIlFPclEiKXIJrr4k/up47w53mo4f0sW/f1roW3VszQnM9HAU98mrkqiQJH
DY9WlEMqcyE7TWJdqt88GYoKIDKHRY18dwUJOQbchTs5tUzd+3ZFWrMYPpknMgFnEEkOUrt5uYUj
gVnOFm6ROZC1fesNNZLzp/OxmAs66KYnAZCeHidDftaJSkGtLm9/C5gpDCN1/Bu7lDbkMyMItTx3
AX8Zt2HMdN9zwDPbcOIFNP1ti1E1lLSheFofgbSibvpFxtoeFXuPexnmhesLqPqFWYRMSXtKWUjX
H62XF6aLQbvnlbbiiLKnlM3WteIUOuXWrJzO4JCYuhV/BRRfHJyMBGRseXJ+IJQJQfvgaxGHlP2u
A+iusgsIGg6mXaqFIK/D4mdjnXyFpiwKPLuGH4uFoHhfOb2xuGT/5BEZSenAcG1AxvOcnnfKjKZi
zaw0G18kwBXUMcA97WEFgaWNxJWMtLy4TP1GB03Rlp+WvJatQRiXuasvlbEt9RIztBG0VcAEcw9z
D8iXOrEgC8JR7DanKzCH0UM64yxr49IzUFR+UpHJxrjb8LWvRbF6mFas9LRfPCgGcYlmAZF8dGXP
3ZlMZJ24eb544dwgr4y9LzJV8vQAy9UC7eeJd2mWZn7/jxTQxXPwd9DjyccbL3hhV/Td1KsnwCTW
t4cMA6dxdEbYtODJjeTVZMobuqNGk+DlChdAQ2SzjAaMMjX4GevtZ1waZwUPGWb7eMH+IRRggzRj
rX3iSpCdIApRG3PFqLCcz22gtuCzxSV9Q9nhjNx7JIQ9jUmMa383J+4W07kX3QqcXaNek+vqkhFR
IBJuSAx8Ac+NNOoST+xsifQ4WEoX9H7jkF6IZF+EzqRvlisRHUQFJ9QtuiqDsfOWE8aHC5W6qG/A
wuPfhy8eGh9yaE5NsBH3oB+a0aWmNwpz412pE1OwQfb96Zk54+GWjyro4ilG5lX8x3wutV20CR7p
EOJoZH9bz0Mx2ZcED3ym5LmB0WA6DYeCbEt4ccIw2Bas7N0Peim8nIhYrmTyJK1U2sEG82l/wSXG
6+lbY/FSWfOOhP6FdjECG/3RlKCVPynYOZ0TnxhZAAW59hCxqgQnLcjjL1BotxQFU571znC5OaVj
4jMc8fGvshAs1Hqu5zVvRPYgtafngk6A9LDXYuwb0/CP43zsCZndwOJLNldGv4CvtHhb0AGfm6yT
zU932QEaWvGUe6wsCOgm5ucuUDJHbdjrbgyXrbG0OdvqM+KwgOtKIOf+VjkIeZCPFleSjIvYKRax
MeINA7BiPcZI3ZvqyV3uR4OON1MIXyiV/jW0nBAUzPLg6I2GgyaW+0r7VnSE4cq+hYjXe3vW5/cK
SjnhmVpoXchMO2BALydzK83wAvzDqyW1VpTh6iDftC5naseVLGoy2kkkL4d6D72CnDzPlb6t8+Or
OaZCJ0nJ2fiN5RcSFXj08gxBFelN5x5ZZ7QC+gr3dNalSDEhQ9H6r0jCQKFUCz6mErLyPM8EBRxh
cHCw9MFkDcOxleo1dDVlp4tEdm/xFYcyj8NjrLULP36aSSrlX4cLkHvR7jNAI24pMOU+e0+GGo2n
AOblX5XYd86x8OurQgOZKtYYPL4APA722hNjI3+7yaRRAsgQw0rroyawgvQQ+pwphjBv9FWHkkDf
y/cuxxBJaTlMZ/SK/wO4MSxG1lBOK22R5zOhzKjSmrpvCMYeTBa8ANiZRh5qpWAF/2RhFF9LK1gJ
1p2isUfvWEB0Rm3IPM4fjy3GaQ0tr8c8bLjmLiXDo4HVMaDxewv+3SDYMXcEt8sTRDBzUgsAkLh1
1ECCmDPtux8tXMFvywWde4mRIBt6a7DKs5j+comPlvu3EtuQFjWLvSbO1pKJ90a8bDTr/PK0h2Px
jUNrQksAyJqpRsdklgWKDTXuBpaT0+ib2CUoEWB+KV+NJu6OWtZ0ewpivPfjvm+t/a+SNQUjFOjR
Qdt3sWwqroo4FFWUz0iVPaYcuTMfwJax8s3Dj1ee1oyMkJqQLmBSCKHuQIQRAkQQK+G/dYSigDRV
eHCQtoqWunk2ZwHFqT0flEUurCQ0lN4UGyqXZzZZAawn+/6tSr08yFvCD17CtTYcENPHPIHfs9VR
xCPa6LTbUgKBWvB4fwQx8YaMaykRCxE0nJg+3a/jzLrlbkbF85kAB5/m4pzMGDVm0cJLZQniIZOZ
v9i7ZyoW3Pz5u3UeOSmu3S0TFrFD73GqcKT8GgnCr0ehOQYF47g5cWLMsALXPG42ZefHlSR3Vwo4
lw9PaAjp9eYG5qVLb1MxLa05CiiqHUuZBd3ZR5w/BmxAQqyZQzn7GQFVDHDDb21RUbhn9SPDZLu3
XmT7ciVkzNIQ6jLP3UxSUtmEKnraclIMzo/bYXxQLoX3rvK99JdNMOXTLfY/TkDQVCqPTmIxenD6
hmraBKhS7QtJPLxUZuWW9HFBBcCRk508KRBQcFgTKvfGOVaJIdMyJTE3fMhhAJhpDfkzmmZ7d/Qa
VGphiPt282t5vo/7d6Ub/KOHc5CQT9QVjUjL4woCjYWGPunq8HM7P2Z83mrDYOXyxEhKEhyBu5Aq
/e6rPpySMPNuVNAImOSUrmy3+ic5gjTN0eaYFgPpU9ZGHuaVD1ppVc5eJX3TIhTnvQ15j24++e4T
zVWHTbVXpNNtE8XE+dVtDP1AO9ibuqGjw2AVmVx0UqUoDNcZytLtuY9t8A1hWAdqYFQajv10lMDF
YbaF+u2dW2RZNGzoTImOMpBud86ncePDSrb4IKtR4sCgsmKx0Ffz01QdN4CICuP5sTm6bk0MoUM/
FOt6epiT2tQfYsTt6pLDTHz9e3jTMpjKr7hsBOpxETm/HBFsw6VmJfsWQmkUaDEmz3hExPy5DzCm
WH3sbsyKoxW7z0L4BXgVS1aKftKwM/5Qn2v6+rIziaxtF6iJC/UwMpPSmd61D2UkasCdDZWrmT8p
2oLQjZnDqYPbwjRNix4utqsacqspZbou3o48k8Bf6n/IcDeh3HDhRmoiDgU+K3w5/OzbaDZ1wENN
ysmX2DGZnRzAaGh9q6YjG8PlM7nBqRxPA+j42hCpNSLcOUfk5yxfhl6XVO/3RLJ4XKw/wOoAmzMm
YI3ticYZlK18OXmjWc5YvlWARPBBRLC4OxygsqeDwz8s5HelxHFKTQ9nwiOeaC+wTG0RIRX0+lX3
eGc+Nktee10C5Xl0qBH/kfgUoLFi75Z0u65EPW9z2ZKZKECkmH+g/dDm6yPqAm2XzyEeJjdqBlBQ
BMk7VXTbMUXbxBgiTXohdHGHzm8LSdOMg8r8CtNgbUU/ob4l0WH5Ii96P2LVfnztpUBJ1OZGceOz
PSbwatrvyM4HpiBrxy2uZ568OeC+UNO7KuT+lXqEhPFEnjEzYeVAdb/x8ylCknQHYZ/ME/+5BbXs
3/12Vx1/qbOH3lc4k5uV17kcxVojRY1T5dUH/sCZdXPyXjtVZC2mzrnjSleI4N8y72iLdrRC3XW4
h+oTrKoF3pGpZ29ksyLo1j2dIx5k1il46tITp6lAXu+08J2C2DnXI5Z71WCe/ipdVKclnHEIJzKW
1H5Yt8N3q5V3NRl4UBMZPqOlkeF8gH8yXT145Mrys7WyWsLP7NBtEuxd0FqNc+P38/D1jz3UqVIw
NclACELzjdQY3XG7WOga3YLGEygna8b60e/HZdtWcBNKLB9WjUueZBb+F2Vuo2laub7y7oY2zMbt
UnvEcPNX4xIErmQ1FROQguG1N3E6/W+GmiEVQhsVDUVnJirwOWKrs7prLyQKO2bJ0lzsI15FtKZp
uR3aAy3anxCpeLfmBNZF/sEUtwF3alwxMvcNU3hv1zVxdN6nGx2p1Xgr8mB3Lp4TQY8xtjQ8T2yN
ydZE1IXRNjZvIzPF1pD9pESKD/0A58VCCj5O+PYkGPKmJxm0C+M9/DD6mOIbTdgN8pDh6ayoHknR
e/UirCQ7jxGe3YzEWZVeTrumu56YtG9quwVQPDlOXFVfta/FwpLvvJ0CRIZ2c1CXLuWz0g+yNCri
If3qdJ1hyF5Nlcu6vh6FBVL0rDi9DABskG8mXYinbxKmHowv0AiMRQPgaCLbyenVnXdw6iq1dRgR
2NU6blJ06S4aZKI5J3jZcqE1Czwtb4iNLVSfNTgpTd+EMrW1fDCV3w2fb5hpLfegaruEC8MHNuHX
dpkOXpB1p1fGkT8ywx1IUo6PfTiUcHSe53cd68ZA2y7Fz5oOX4JcgpIuKpHe2OVZMXvaONQ684h/
9qYyFctpQGjbWTm9AXe+WAaEmEhL/gSx9GMd3J37y4OoR6zayaQ9IYZ38ZZAj34/u5mV41WALMdL
zFSR1XnH2OaJMBBnYR4oVWEpd1mllzh++VmCq3DvNst0OHvPb3IFOMDmX+HLFPg6VVhJw2p4ul51
K6Bna401PJOpdtlvUYsA9o9mjoEsx6o2RhV/WyN2+fagsbAdhSwCkKCIBjYG/rXi5zuCncuUrHvU
DaMuH+/pjv0rdRcpSxgsQmgkgIskGQXU+b3MJQReJGojwHQ9KXSEUeZ2NYRFYfEFJFZcK22W5mxQ
rBM8oI/lPv6jddcjRzoRZ+GlkufGjDIQee2AaXAbB40J3akXZhRH065RJkTxoCmcI0o+Dn5sOVGi
F+7is9UjdM8Ek9exYV+2FUEIWy3JJEIhPuaLujhTnnktJpQzXfNNWAnqm3JCtPHEfOVZLNXOE7rW
ScRmZ3CBrv2ee6jawSU2NG43wzvT8Edr5La6xh+kvZHL25RBNGJaHyCF8h/nhv0JEw11f+qmoLf0
7eeajX2dQkbw00OVkTsztE74noCb9dCV8MpSPZ4VgFfZXrfRTHzhlVpGHjovE4yYt1rBdPicCg50
I6AFHGT1Lh205tNR86OInHuNcgZdK4tlgj4nUTSNXEaU8/E2uLBQDDg3U5C7VLNooYWHFJu17cWm
MiRz5xWwSCXwcFWP6+/12OzIkqodwqUxfam1qTTkv7x2FmQDvyTvDkNf79RF9/rJIyTD6Yq6R/MG
MqrYSf9HXYuOY9bJUNitlioEaE4A9RwWAEj0zAQNeA+wsA3QzG2g5qbu+d08u00XRoALTk8Ha8CD
V3R2jhJiR6SVzWKagXM9Z3XPwn7oTCz3KKRmDdAA82j3TXIj9e1GrSAIOXGc2dBGs7CGKgW71Rhv
S+ILymRqsB2U2EvbYIrfjJNMTU6kUNeIMw6VSWmJC0XhwqhKeSHzxl9wLYekdV23AMBRMoOkEOIV
TCrActWFXtQ+g4XoBZ/2xoN2y1/bzbA7NIEZGl60XJYSehalDg3YQRr/ILydosoexwO694RKqvLG
0Um7zs744g3TcABaBnMwpDProI9x3fOgML78Ha3Lbcp6oZgl/bLRAFnUH19b1ZHP3UVzn13x4x93
ZvyuQWVjgzL1wTpfofPs/7HeYAz5QhbF/KVR4zF5ilqIfPpmczHM7G5b5WjenXLqF1NzBXEmW5/A
5lRjLznVt6J5WCYnJ7IhscJTdeATXyhW+BNtAu0Ti7KJeRHPHA70pKsr52hd+pQ+jfZ3wtgaBoWS
YHxB2nvlbfryB4liRScDiq4YcCmH4YSsQ/3GGFRtTB51Vt5r3OBvZqsqV35ECDGQsRRwYVW8zz5u
FzkUc14OjGOsSvrmF0aJJT/v0kIo2EihQAjANK3mWBVUmymQ+E9doaJi65ws1vRQ46RKWROJVSUR
8f3RDhxXpPAvyMvWPmI1iTs/QD3U3GyQSLpkt0I2Du+ut0nnNrqkeCOsqlj01ABe4SoED6AGSNH/
SUZTWfQEGVJxcUOqOKw8vT3+AHL7hyOGTovEv4vSFil+7SQpgTnifR1H60HLu7RILt9cASx6JRxO
YyS4dSCZJR6V/7Zjt2PtAHJ0XozMAoFfnxv/aQtiOjbO9yquTVkbAkjC/BdANdgpZAWb7lrt5QoW
TYFzHp14LkZra2i8UFH9Im3NOKLtz+Lw6vrjgWWVer1GWDXgnsiuXfN7zWEHsHRYSy/irFO/AgIl
SGWzYUsV0Y1QH1AJCRUqtjq7moGb9L6Vkh+StuVaSTXP8aFF9xJ9TY5/OtwDNsqEt5L3SXQUwWeV
l4lktPFA8C7w3L/wIg1Y06QGA0w2eUQmV6e0YhSRwjSAl+RneEOjBsQArXUVFwa5z1seOx9aHGNF
I9qxQXwzhAyZzQoCz1Xit6KAmoOuc9E3MTr2AXKw7XPb0Fa3DcRDbabXFmoor64THQfNcvBxgQ83
Z3gK14837C6CAs1UeH6xSdB/NsxKTeGolur+QN+twaXj81frEf4QtDfw+Wpl6n+JDjFtRx+SOdmV
XbMaip3Qzk3aIjT6wlGtGSazfoBD3h9STbv3ePKoUFqzz4CrILls6sqDzHgkkvJSt0DgqSqk62DC
LjobFzofCGpYDFeAS8FwoFrzcIy4s9dDcbUpZvv7SsXBLH0PCvOMn7RPg0Ow5qMytPJGCgzG4JZ6
McROjTbSe9yaxQzWlXlBsqvLohrTgcYFEpnQCOO+YpUBz1KqJqWsm9AUEs0+Ye1JNsSwYH58+EXF
Yt25T1NzV7JvNw0UifI+xpopOkkDTEeDflNeovdri6SUTtlZfQ8nZe4AbxRUaQZu96J+CmNRyK/9
fcmdE82+tkQiOAfvSapfH80UTXbDkoORk+YFKl61WwvdoIU7Mgsh+78bReW2+RNJvVNzgLF0w0+3
9sQZITzCYlK90koT3YRI64Fn9eXXV+iGXOuymqK5GxqyDP/CllVSFAromjCkpAFn+ecpqZaR/WxN
TO3vwtvjWR1vhgIEZB/l3fOoNHhGdZ6bh61R1sQOXjUV5iIPhSsBXY38XV+JwYdCmSot7OA6ip+f
GmweRG/Bs32stJ6rRotffrAR+5/kgYpseceQivevQ+UBNJ1AULL39kACQZZuBrjXwBsDybubc+VF
eBdhSd+fK1xLsMUBrPAm2zLcQOTozDwP46+MGn2Mzd/oTnY4hDQ9GB0TqdUsyyGz/bTm9b/Zkug6
SeQLghQYF7InF67aKK005N8MUh/XR0y2UwGaG8mjGiIkkKfr3nOJ8om9nd/ZnlSaxArEgsAjNfGW
zMl8crQxnE9dob8OQVLmfk/Uya4QmPidPpUaoDxpm3ZdxzEZphMjvfah5raI0e95HKs90VjMBaAv
Att3WTtJqx0FKun1AEK/BxVkt69BXIeBmbESlB+He6Xen13kzPdnn+w1ZpLowW9XsqjyrW4hyqTn
2a733TTbyqZOgGaOjxgD4yYYbTFZsWgDUWn2iA26NOAVNL/C1kKybO21jhEyRaJJhm4cc0hD4+wn
yZdx0Gkg0yhnHtCr6byZVvuXUbsWaApGjx/9tRv3d8UgpMbVoNEdidcH0AoOTV5F/kQNFNP3RqJV
Upn15RVHjyNtRqcZeWGFZKsi+TmDYLAMJ//7rSUzd2mifxhXADJlr6vxUQViGZ/WT9CPnJ4q3q+c
UJnYyp9Et+9u2xnbPQVdWbFUwdZmzMIo1I11izJWgHMNrfwCAsSDJYtILbMgDkS6vk8z+Yr2mFd0
I+8gJfwbhAjUzFVUMeUaXzDcV4RKEwROR7ErFWEWeRE6rDGHlbH+lRxwKtLxrkKpCK+WNnp6jAQ4
7qfO7jTkbYYSLdE3LlaUJVoZp49kOx8ka/9UJEzTBlWjnTzA5eBwbnKWm7VrHJCC10WDvYNgMJ/L
OBKbRZrYimvs+XIKPPKF3Lj4uQquTvRrrq52NrkoxoJUjyNhF4kqmGQdYJsaY7GoX7/YnXF2DKoc
xOUE4bARKtIX9kaTNnh+/hdDYFtjMSMrD5DtwD/kFbWABxe7gOUsxgdMIWHLQvdyIPP78qrggf68
dk//UcfGC2e1DV5Atx/rM1L6P2AIa8uAgkzKlh5weGGOAwHwISmTdKQJRWjB0Zgi6pOARmicx5qL
2ymrnfEkZ8gU8HsGzoZWwJR6hwwfViJTzJJ6H7UDwaZWjwjwnZ67XPSDBwFV9NzfFFa6rGeAiJb0
KZhHyCJumS14l28VOTMBj7LDfa/83Lobw0wDcHf7vRjtCA5cvZRXqoN2Cg07bBVka6foO2hRmT45
nrVScZTAfNDfD+3xObWko9V8CH0vsJLH9wkRWKvtE6gzY2LojCnYdxMealEWJZ/rPJrJs8w1xlZu
JnPjvLo3ldQn6jkKpxiDO8IZcQ6RWJ1ip4hMRFLossUXdcY5Hy/NBbA5b/omkaeczNdxKaH4FBls
bqgK32a6yWsfta7/a/tgAWjKvk7B1Y4IPUSX6NyZ42sz+/g1cDL8A/3p+RZcsOT8Yjq5sImpJLDU
Q4XWVg84cAXyiqukWWdze3zSPc2BAPxgz2tv16occXIt5MVi/8x1ZSEskv98VJDZhlm97ftCjlKm
ykPEUeTSXzujzvdu7y+ofZ4edXgskbEMw1/Mk1qBa1OpjJsCGwxmN0N2ZGLr4rzNQUhy5ADgGPBD
I1PWZtZX2gAo4t01JYoMkT9YSL4geJf1fN9MledJJouYiw9MosLnf4M3xKtrMW/oc8tWU7sE5tFF
m/qNzC/CyrQyJROZBdT6wZWvocnlv4YmnBHegy6L8+4k5qbekI8f+z5aKrNYpfvkBM31wVIjljn6
tyytsP49u4LmXydGBHXEQkY9GmsxDl+CKs8nB0ccXJAKF1pRx29gA7FF7PBB7+UOy9LZ5OHZkTFy
QslZN1zyoqLCNmP9EyQVFoLoeUyEPxUSX9k/7mS+uGgJ8/kuWDhYHeZbnXkxkf08lo1PsB982X/P
gRuNvICCGgFfVTrCIxOhFsSqJ1HOGVTFOQNl+ELHq0egGEQ+EyGYad7/B1WoaPCBLVI7iW3sbpEj
9QWMRipXfMoH3rw2CZV4JUMkIcU7IrualHkrHkBefGzrH1+vhiAoHQydYLQRzTCQqSSrgrccbrJg
qv53gWapzAhHj/s9SGU2kLL7FimEELcPNe6H5GCEwZ0R0Qjcq6d/se0nBIw/bvkt7Ru5P3QwitN6
Alroep+VYlqNycyKS6EWMGrfn6KE4lJBwtNQT2LSXLs+g9HvRnmt3FR5BXud3LE6hDgAzq8E1q82
BtgFgEMjkD316MOf9Fhv6zfGJRbl9hn3nOl4rB1/kZZkIZU+bNQNlTnt9TCbv4drIAQGDW6TR2Uw
TSGOoejCXZC7H0BGtl0qvFUxUfGCP9zwCWbpq0JEkeSz2tB2/LPQahZE4Tl1xcu4E5FHuoTZrd17
4Wuy9B6dt5AvW3T7U4XKfCgzY3g1hlrwhZonFrn/5iqkPIIgMGLgYQ3gW9qbA9SotnFlNpag/XvB
av/IaIhTvrdCZeURQ26gvgFlfyb8eX4cZrY3o8fSE2ls4mHCPfqAlt+GEMiHXT9+/3a3s4fvRQne
s7qmodyVaDy3YOuWGfmsvvD+73lj9Og+TlWcRLUZnfZtn86Y1Xi8NNTu3cU5HzJxFfe+heowsYv0
pkeHxW1urwmWiunldg+jSJzZeui5iOZMiw+KO5+7dMjBAk1qXcvgW3/p2jniahDQaZhLQFtD7sLo
y5BNpNMMzYlRLoqDBzmzBlpYnTPMAs566lq1u4mOi/qjpOVVcML0fbgC+Dqk+IWe8/3YRH8cZbEz
rD83FfPPCvYIJFCaajEi28t94pOEvUyHtO9ruUS+jlYgdCD+nZvMtKk+c7uHGC4h8u7wsQ1Nf03Z
YNDAp+FIF2dngaq721XFjCrcjeZD+vfHLYM7FC3I2xWkdZTCsenE/gZhs+8h9XwLsyKNkYnzvjq+
fasJVA/tjnzeu/YOUTiBe+gI3n6ILwxP+DFE+E2By3jr99gK4a9PzUjWnwEpdG+SEcf+iW5o0h1j
RNVxBCM77Fqi9pbsBo0XMhh5FCNLqV1YEyOOjdxRGi0Wbd+GAeQyYl9QmeJXHiZFOsd9anJSM/ZQ
9BVvrYPnWGYCXNANhmhpEq+FP2mM9GRVcbipQ1H2snSiyOKS7Z5JnAYUvTIzYq228xvzD9KXDChQ
/lbH8TF7r4ubpIz3gM9oVVxaFv7ElDkuI+dwrhGLIekhKiDeyDVqpi5yvR9lmdfXPeZQXBTBresj
QsTSsDfSGf0NSdhWD7tlLTn8bgWM9Rc49L1Tl+gkUQU+jHaHQn3Q7WkKbp2ggn1jVh8k9MPvPrmS
PHOu328I1PWnoKF4MXWHCjrrgpKtG2q1o2mP2YhuSSGvGYXyec1G2hN5wRfMm8h91pNks7rjYsPA
vpGUWTxcuo5H/79vMCyBSwgmxhjXzkRU91rVz3ejq/DNlHohika5eJfx7YIaWBkmrnrSygAHEOzA
54mjGRKpZF0/W7GpWsEZrpdrnFdRPP+fin8dFys/XCRDw5DexvU2Ul1BZP8rB5Yn540mh2IPloUa
pCWISDJpIO1N8tZ/Z5f96nzg5xHi6eD83h/GYjnuHYn3exJSx5Xs2MLogjqfbewyY+nAgR2KiYir
JOdrfzKAugIyeGZuzzEC6M8Rk3vP+rNdyx4HRxXpPxQQmpPXKRgsjkgtWMVPzW/0BdOsONCUhXQg
7YPkVYIf3u7GDPe3dR1EESsfpx0ikpqod+qVF8kVglT3yWXeolMCLOJTMSmDsQV1Emx+hK1Bmk+8
nBI1o+jwbezQ95t1/CBbB+cJd/XIKB2Zp0MOJHDh+/VPjkWz4CasZiYUPye15YiiHufDhdQpoD2J
BUANbTO/GEdGkxWpbKEV2i4887tfy7uqKvFKcjBBXeH/yo3MSsGRcXqL/V6luDkHOYmlUDJbtwbd
r3vI0X+1XElS8+ItNPcJ7PpdFXkKgm07umTAE6QasirAcW2Nsp8NDJPLRYA6laEb44xV2V9B/EeB
VqpkGJWfpKhcAOeSI9pGcp1t9EsTSv4cX+3CfOetuU2E65dTiwMD2Y+YZMSYlMsc76lg+fQ4HOLG
6V4mfk0AO8FcBKPZbM5TcG/OIva/LiAKxyAhKxOUW56Ac2Ed0G3ZS21vsW/EUDEomCUSdJ455XK4
/sJkQO5VVz/rBC6I4dQlRJcpQZNRvu3HbSsKzryaPFShmQnZdPpC/Is5PltuCW2QI/YIPDWyV3iU
w8tXwulA+GakbxsyQC3xUorCM8nN0xFOlJM77FExOmBpLL1ViZuoxAmSFfUr2N90RMFERDKV2AT8
lJWkRBFKx0z3GeqGMlpfeuq98a52m0ie7be9WcUbb04yvRofdR1dVVPwPz7QdDomz5SNJ+OlDXeM
8kjbpKY3O90Kl81j33FruoTCwa1+gxMno3p5Wk1u/EIpNaaemBSp+1BdJkt4696YsTQvmcrRyiif
tZ0/eaJQ/a4Am5is6X9mXe6fZTar5VhCO8iXVZH2IZKfmzF+9kBQBH53V4mHDWbCO08QFIsVRRAO
B/b3wBXKT7g1yEvjtTcRt58m8qL4+PX7lpOYc0Awh6PyUr1nhRNvFN/nessyi36xVZTT0nQtBnql
+LHewJ+CdiAA9z0OYKToFKUkwNc72YNPMRAOgK6q5nKFIQ3fGn8Yz1CRw7CgCE1TiX31IY2ELCSt
yM5ENyQdhReQVm+pSYNJv9sc4h4p+2rCsMx/cF/roPFAYMuNc7rY/x2egGWhmfwOalVoQzPwyJs4
qTgnChZIJRMpQUnsoToYDLooiSehTZeIEC5BOMB48ZWx0jIuUDBXd/r9CnKawmS5xYAUEyQ2tE6/
1o2cKjLm8t1zPLSGMFk7+ZslAKfDsefcOiDOWEv0iA0i6JcpF2MoEIBxH36xQ026sbBS061t39Xy
oYIagAATy0/a/45xKipEXKndUltETpsb5zOb/qzT4se2TJkCMh+Lqkfs2tA9b+196SxoXpQbVZlb
KipPCWAmTMi/OrRaQrtRsALKZiC5v3QK5PIV5b1CtxaG+2a0pL60KtkNzbXRWhBQi/5P8n/G+u4x
ielBCNWCfxz9Zoytierc9FbJmZ6EkMT5bRhu0QgG/IDeR7SJoycdGpKJm3nkfEqc0ONuARVEvLbW
Mw6kBXq/yBCbCcP6bu6qDhhSQEzS9Ec+Qo88MBaKr+p19KKfQ+PnE0/CLHBEuHIKcBvGT4CopgPF
zhO94Q87/ILmmdZB0uAhA+gAv9Gw5ofeI6m24mEKEfCLTWZUjzP1trayfOV0pf6ft4oNDEq7N+Dg
UAtPEraQQR5DfKhDDsrT9hlO6uSG5hRJlqi8/3+RRsnknxzEI0YQqmSooTmPCLH2DhR3NvYPDzSO
WlknFc8zj8j/ISzCo+JpWiPdV8cJE9+j1p9c9lvICW5on9NejgVlaGXI4vmLDAMhZWCDKmxUlHCz
oigpQdZu6WQ/HpgZi4Lx6xeX1C7c9misS1DhpOr0jt03O8ZJNGcql9Juz6HMNqMF/K9pzC9snqlq
pbxm/8RDfOEwmxx6G4BU2h/iniFRK4TnZzmJLmCd/+dAFTcyLqFWJRwaGCYqzW63LisuqiM8a7QC
qwrZiwj9zlZvhGlC9bs+fXRnS2ReaUJXqp2VNggdMqLiV6dJFiTHMLnenvp/MwpHwlUGnzhU5s7H
RtjU+wIdsItgFckdCkQnTgX8eC+/OU2RthriH9TjACdco30k83s7tI0NgpZ46nQ2Sa/p6161pEyY
baIeWvD4CcN83bNzvxGAoMBN8pQMLzqhU7jX65dLMLoXAxOP7+nVHiGmdA8cVb7Iwy/VPqvUa17B
hgcDRIx2jGmqb0RAmjfToYkSoD8ovjH/xqIhXS7ZbGLx35K3K4Ipnji9EAVDrN6unc+HzOIGswzD
5V7czm6CUi3B2+48QrIZ66TU0GWer8vtVIqCV303B2n72L1bYCqda4xAq06Bbun4ILg5tSpKgpzN
fIE6uTKznmGHDoI/FN8X8gHZ7HCb5H/7o1Q9xz8MCPr0hTIpVX2eDFMF+4pPxDG8AAPcX3en6Wg9
TqdkfNTheUYjW16Lts6DsBimnUpx5Ypoq6lemCjt0TYnwBG1Fb3odgUzbCWVTW4uNUYYTJgTJCkC
AoZIYjiXvXBCTWYHhzO06NVCBz12oG2Rzy4l2hyetYjqwUrK9bpkWfwCoTACq4cQpYjJirmEZiKp
/zQrEtaTxNo9WtnWaHxceFBaWch2jUuC3Y3ADH46H8g6IlwW1GlE8yTibmER4cxtKuQV1mMc34Oq
uXvkApCoMcIpGfv0dYlP20qxQYsgNSUjkEuV51GxN1R/7JBnz0Q1eIffC3yQSIvaJwMTJdtpzw0K
TKNa07wOT4mkbU955BU/3f+P7dRwHdzta4QvLpj/hKuNCKstg/J5cJaxxtgiO7EznsfgKj2KyNBA
L1KGYXfqS0tFHQqhmMK8kxtjub8CdFSIhsgsDFAwMTlm63fJSCcYk+PkZd6SIYc3hVFj5p+7pEli
9f/PM7CEbKveQMlbg4LTAnZvN9my/End07gg0S2qnbkg05RJdcUho3vC3aTtyE/A3MeOewC9X3PJ
vCwnzUYkwKgR6qdwT7GVP43ViHpTjDfJAq2bK0Xm9D2TmQ8QaXJQlRGZxc1LcRnPUNsfkV+LC77V
2jjU+VcP5MJJC2GJZuxJtQZc7ueGJQFutnfXLpp2suxWSZK3F4HgeQ4uGxAbLYU1SIbr8rbEnW3x
PCMrppBJtWlk/a8zlbh2WIgFynjNUUyc6H7ix+hBU+FHLghgEfohZic5X0ZJ68BYdjzhaUqBMD8c
9Nsrc5Xb/OOWnDCWSarOthNI8pbhdh9BY7niqrae3psDrjIz63MaeHrhWtS+KX4yUrqV9ngr0366
5s4DTWGOKzAbbP8IycEtDyBbTiBJR4+W4848vliKOixIkWGSqWubRvF5VmTg3BVnjxkJ9rtlDPVk
2KMTruNZ9gZJ6Sb+rvmbsGki+AuO5BTwEG7RL8cJZ9iFkAaGmDqvvXwGzRHqTHrsrX42FCA+QkDo
c3NVv4an8EVUXxtj4shXEpLLpVQfx0nBpULUqNHLX2wsBOzCK1ACW6RTO7txx6XHZhQ1rm2k9DGH
r7uN5rTRQ9enZcX57iiC3xGv25OMlmH9eQRHi58motpjl7OShiaDKDEkZdQ6S6Thpk07LL7G5OPQ
rWNfDZ7AJVR9U7o160B+PxY5/qRGG4s8RLiHT5R8QHONydWuLtAUx1iwo1gwJwrBeV28RHHypkro
Ci8VEZ8q+DHFBlCK1+pqBF2uKmLTiHrd7mQEGtwhuIpIydivqH/zTwHBkMDA14eEFPdfTsHOeaiQ
OwjAuK67aVdMxaI56i+1ITU8upgLusrBrz84bg+HReLTSJaJk926cCbiboyOMvmWpDFnowdHmpVY
bnpj1x8BnK1nQog5bDyUc0byF/Iy+zu+8TBaI2H56jlkAumfWyMsOKPrbssr+4eyyhmo8sV8h60/
yL0liwA0VQgLj3cmJNqww5TkSnAxkwBVSQFyNmgdl02VPbmuhfc1jcJzeJQA5bKY8YMgiXSoyznG
AFofYH2/zKCxyJd2MM5LLWK6oPPDXVcemfoHFA17Sjc6k9sPkbN9chO+nFi+YZ36AjBnnigY02KE
B4PDYrIH0qB3vFTRanCC/F/pREvHxS2NvMi9WjO6oK2JZ+jfEND+eo5277Lu5mo/Avkj2gnfqGFZ
/+sUxt6Cj2HV6D6ubokIvHx7QwGf/nyneRfDd05Of1f76YvyetaeSH4NtmUQle4hSjm14ALlCOmH
Xfxzr7GnLicQGACVj5PeEZ5yKn9TmH7VIqEKVRCu8+sR10tagrNcrEo5CTYh+Dul4fa4iCRTCllS
drPcbraclLNDHzsFMRRNRWpOsmwCyfsrJq3l0Jwsmff92rVYUOetnLev3IOCZOiROcbkmgZHrS2+
8z7Y5+e5uZPFBGR+apBaXguCB8FblMi94E1UYE3eZtBFVUtGuXZ0oPFNMFkbI0qAedfFYspfSmcW
dgUGm4eBOtHYIaa8OTB37avPab2tT4k/25uIP0AdDgfaeLlxhzk+dVDzXDecnVITBNsOqeKHsoj6
joI2Ow5TmocxVzUvN/stZLqGQfgbN3swEeDbYDvUObdU+yZGJesdqGrCdKIGs5bLwlIq8forCR1k
Oa3RtRmjg4akqQzDHmw9y+3blobeO/p5dolHrA/0/xacFlt875RVE2fNnQJD+mW0GerfqfRwAUMm
XHV1dHyGdEQppyKGwMP+E4TkngRqVcaYD8Rv3B6cf0duVgM4LHLgtiVpocKWxgYTT+HNF5FWzeS0
yv8uXT4s5ruCcowobk6t7VbDUFvwHDI4F1V5N8IRiSJgYndw/vmX0qhD4LDSFd0PUdixNGm0HTaC
4wkWWvWJS9EIBC4is6QPnQ8c54Eun20Wqj+r0zK0DmgmGrJXNfYmqRSlSeTu2vAfJStkBCR8uIf5
1fWLtNFXranbRPIsPLH3IHkKkRb19Db6hz7EZqJZJwSz4VCKrR19h0WoY3VwrVVUDoviORHtnJZR
zSL9w7I0CSILIsEIJydecQwMurS2UF0YflwWLbBoNeqwFkTkbe3Pqk/qIwYylpnJhn4zV1fZya0X
YOWL6h6lnwuPFP6xYxd5Ucpk0kIUziqBGHZUVBN/j6JiZF1MGj0lSwTKJ/CQPjXoozbJtQ/NJ7RU
tAnpnIgNFp2aT7iRxjhVJ9ENB2ObleH3v1Ho02/v8rtE6zCg1IJt6IYNg6lf+Gf0uOwFUrkb7DC4
AQ/uVVtf3HbRT7x59EGS3x8CAekR6sGzp1IfzZdOC75jJch2BaWx2Hkv47nJQK/mRwFNXSdqRO+b
rpbrkbTDN6tvKjaCe3Eol9AsQf/7pF/UoWa/uq5qGPV7L2/UNKYf2tTpNciJjvufEms0/yIPIqK/
/PRcTX7u94xrR07u7/UAR46nFIDoh7RqjmzPNW6ggkuQ8AnqNkJhJwakB4IKZ1ZyCixjQA7ql/d6
/JSrk4HlW/irqHmRUkwVYRVueTcRUkxU+bDv2DKdtdxFKb53KOts1DH2xoI13hNNqzeboxm/X/8v
cb0m/639TXCU1OeglsEwXTeis4y3BmhURWTrt+rru56CggCChaKofxJqMFsRB1z3b2WEM7N/f5G+
mQGyx8ckns9z1w+uG0S63HyvDDWUeen0JdR6nk9iJyMV3+wJI+wvvtHWHJqvDJHsmKyd5T2r2xc9
aFMZDWzkuKcqWQeNg+k9rm1hGv3wG5phg+7ylyTRsjznnvqHPbpJbumuhSrK8dN0rBTsFjjvv2rc
vXyVnsj6d02BcdtaA2S5DG4nnrIfkeHXy9h6mECceRlXqoM7QpYfDmhtnZn9eCSA6SxvuL9W5Pqw
kTp+CTHdd3IYJRW6mRwJGsihaDqZr24gh7OsWopaAfAFtvFWzQQHI7PErIVvSOs3AreyTh16T8pV
imiXY1ByWvk8Ke0N589gV2bCxO24+sQv5JahgAWBCUmQ5ibmcYMRZpCvPyu6x1mafjtUqVPT/oC1
yTipa+VGHwkGD7P19QmJl+fo5Pzn9WQ6/7ToQbuXm0S2NA1PETnZV+HjHwYrNdgwNwgeeN+tHbnc
PUSOGiMPLMVmSbnvyZuvoAUWtcHMN1P2WS66MUyp8PFxlRH4vgsQIsk3DH08g9qTTozBrfcyY/hQ
lQhhQhOiGEVos8Gm8yapiO3Nq9+l7EVQ08eX91L38NbvMy2RA6+B6KcFhBNBQ2TWyUz2DQJYO7h4
bS5CaZhJ8Mb1h25CHIwz3/qC0y3tV9s6wptVbA0qyhRl+LJ7bhNA8QfKjrcCLVOhoLaG2Sj2Foh7
aZFZQlCy0Yr1hYox4efrgPfKasPTsDmNc90hH0iYjA1SikpzwHCTtYrM4UaBukOMEz9YQvN9jDW8
S+iuy5bLoXaUB5XJyFpuVlLRo22Mj2GvaZHdZhvEBhhWMbspC2ZaHDq146nZ6gOcRgHjX9gsGYqd
gd7JWtTq0L6eYF+nCGb4NEZhLl/u+De9KHrn4kJdqYZqvhdIjFLNKOyN8Shyr9DZAK2ybNiITg7K
pGzv/Kabi4P0kriPBgYgEI/VUepoVNFcXsnQKsa0dWw7lMU3pln0zYG944omLgcfj+oBgWAKI7vV
pMDK4kg4g5V75eWrKcCWc3S7xK8b9b/ZmleU9QGiF/fmhoo42tGpW09xDOKe69xsrPJzwPH9gJOw
s0fgzBYqzinPc2GKdawUhLDEPZlJyM1bLQl51Rv3DGlSrqWRJyCr17Q36fz3AgUY/objioYeqDWJ
tPnYWxvGllLdK+Rbkie0LB+L3YZyEPtys/mDtPng8iR7nJS4kwneG7oVgojNpG0gzAzMWx0KL3gT
NB0EDP3kThGUQuwsp2MYKQa/4X822ox9BIr3vDpShfUbVWhW4IvgWGa4bMkKLAEjGL6v2CobGvjt
6Ui8I7Tr2ZRhv1K3+LsIYQrCqlGPDR0BaY60+x4RIhsjhbg/Lrz/PSfaduFPprpbCoVj+wSjr6Vh
lJN31mgra9UEam1IZYVuzyI13gF1SPhv959TMUAClDLcy8gwuAJoPKRYBdX2ixsdcXShl2FAcuyX
pILAaCsEHKUudn5ZP2KVFJZOYPIvJ4e0eV8vsZ5ex+Px9PjZqSvJ8vOJuZhYxM47RLELU0a6nzo2
o7swXaQHQEoQGtU4oI68DdSIKEbXvX4lrhCxh4R0EW0E5gEelZM3oHC+LSkSTdVKPrVPXShLFXpn
VqFATEj//t7Ei72xfKsqqLpMvxYyw5Ndo8AB5nCUGqgzGed2wn685Griyy+get3XL113b5d4KhIW
QDuerPlKwy9ocRDCb8lnXautAgsPHcWAd1LtSHUPJoo3CGj9bOyKfC5XIhu6kwrWyQqrQA/7gmWw
WihD/s0ddRGVVu8snjo4qVkfgz3ZXIBmC7wAu/e5KlkbrQTjwZtlhav1hcoaVW8nKjV9lminnmUM
4If7dtLYa+hb/N/xOC9LjpR+PO+v90qn25XT0xkdUt+MK4ShDp2qN14AJEzVjgT/mAe9q12X5tk6
JBnfAbLIYskH2Z0RRqBDwK9hCsSm2O0f6vxtzmTIFInziVcS4043Wkd3T3a2vstt5bPuTxzpDk7D
HND+xy2irmrgXagwCtWCcYHiqpxFieL6AKSmlpKvXucl3kK2T8aaFGVf/yDdSJnWoHxbdWBa+Lt/
P8VL7K3dRC41zO4R/3vdePMV6zRccaHwsDznAM8BcPV4rdhPuCRQ6B7y86JcnfFMII99IEYA6PBU
JsNGDBxCCHlmFe0QwHwoS5+Wm1w9lA10w3+KwJ0Vx92DtWlasJJFjXXLbzErRrDA9u00bIZ52tqs
30ZqIp4S9R6yZpf1nEeYqjbLI3k69ejpVMjfapGnern74XYP4BxXMRGQS6lXocyz03NUpokBx1qh
ddo9TxXKeVGCGUDMV55EkK9q93OOivRWNNKTvz6bJY+LBwY8q9jNhaPHCgOomSD5R9xxsUiFkB1i
X4MnJdTIeFIbDk8Kth6zxsQXbmUhQFWg8uRa7FuHANYsP02AFRS+sxXHxGKcQe1z0UrLOOVr7nGf
vaq1bAh41Q2uB7mnAuaTY6xnov985xj7FGegVDHHIkOj+GCzrl5mlXVGJ18/ScwCSVJZeS+3FfC6
UMDMjmLLj4C48WFgN5l69ufnAKvAevArC5r0V39IuUT486xdMn+xBtWdvMZsmJUylQwFXv6QF6QJ
NWzn5c77TPT/0i2shfeeS2dWshRsmKzwFU/vEQys+Y89+3mXK1jFDD7EryGoDQX7tRng/3WwdWSE
q8QVLkWoPm9c4H/SlNrrUINcGhu8ZcntKubBkkMnHzFwarVeBqSBjN8s0tZhD+V7g+SSWciD8cOF
GAOu+Z2JOyH4SOpYfx2K1K9Ibht9j7/LHiWsTa5Eawh39CUoa1I3s8Rhi3PH/UpqDr5IsBnkG6l+
5Vc5rhvnT5hRm9Apl69ZU5eeEwZR49qTvwPEQ8MIJUYZmdyb+8AJ9LQFWrVVdoo2/0FbnvSR76G8
1BfX+pA86rVXLUTXJZZdm7lc6FbLOvvB5CYJWgwlcq576iPIe42XZAiiZjJm+qPzRm58rXzjtQbW
bSaP50Z7jV8XeOw/iM9PSChyvMrVOio+6Bv85dkA/U11EJwbMJklCFUtM4N1DgfQ4S++pGr69baE
vZwaPiu3a9Pu7RM9O9gWJdMMJD1FL+hVJpcziqfeW2YXQnKUJ1VpG0Nu7BMzHSepLOwWWe2pbkBz
TrC6CD6t8uAOUbFYAMrRu5sUgXrO21/9rEUh2/bRnZsKfIwtZrSaX98BWb35hwtY6qTJI4srdRpA
IV3AgdIGyEOBJE+I3J1mo5yd4xGq/67TyFHWjHZCDMAN8tvw1OsBe+AfY38lVKj6kM9f0dIh9Tjx
ESDq85WM14x71Id3BDc927X8C8tHNmlkjvgy04KoBRl4CXoipLEdFtE+/qtQ3/AcIOA8X2YGExMp
x3B78NaWKR+N8K1la8fkcxeJPGPh+uNwBwQurnQLM9brKb+stHhZOfzRdIWuNlfeTtfRVRvaDbkX
l0Zz9x7QDdtVirDd4/8a7v9ItMeFJWgIyCzbPqRMmqtT3QQs4aBVBNF0QvlyDQBIlpXAbhh62i7d
R8pSPDWDoIo4wjxDzrZRkl3K5+/hi59WbFEOL30s/yEWeCJLKhZUGcQkyD4wD3nVF51Y8NBRNqwa
37fBmz5/Y+8gCOsXjYTD3iQyv7tFEJcp8eMpWoBW6YoybzuKg7oVtoYHpmTwvJvgiDW7kPIEEhHB
5PPIR/mik0tPjWqz5/w+dcRTGjDacWBAFzYwLC6aeN2xNjnfWmaXQNRX0nQLoV968cYqZ52g7VJy
ofXxYkC3acx7z62ZAWvOlpp+zwKb4iZDiISjYwEGKusbbru9Z7zrmHZk9dG9raO0AQIRUhu5g+1/
qF+HMQNcHyHlqYSk8JdUe0yvWFkrRyQ72zEMbAFRbiiJXC5rpvAQFoq2FNta21YYsUtPQAad0Jb+
hS8o1W/w5M0k/obZzcI3nxuDGB8zsEx8PsZFBfcK2G8a6SblwKOCZtZ3kUpuN84An9T4SYtW0A6m
uyJ9zxvm9FsgkiUcoprVbiYNuH19sn5ucVa6TxrEQNH/wajNHxWJA2W/Cz0YylhuXKVdOgFwAs23
sB3G2j8yOwNRiTe+lMCrnmdq4j5n6BxBHkJUl+VPcDJVHoRP23dnWMYWCwKqQ6efhAuE4pvvwaqf
VP4kyWAcV7cga1A7HM/8CeUINMtQSlci65n8Ae9N+Cx6oxlVoCz4rAsquuRqm2F+IKEESkPeV+eG
uSqo5NqA5H2szNDBIvTqEAHZUY5K+M6AOpWH/YHpfOacM/pw+zLDuBiRtIPrg/pvoa6buutjju1C
65tsTOfNDH+T7XwtCXA4bYGe2SiYMrQBevxRDarvdHVFnjxsggxbgwq/oVz1FeJgLAAV1EqexwkW
tUDGwrnVwSfLMMBJKejBF4AXO0YOLnQJS3OSyttxYbgrdHmbHkXQjGwlV3/6BbkvzIyOnxCpkL+K
6mZV/8Q+U9scy1Ow+GZtcItkZ3T1IkEADMjWYBWQcc9XttojQHmanbu4Pknyb+1EkZkHtR4GpZgT
pq/yjULOS/4WMU6UEpQdcgi0jWZRmo/SfVsGeS1kBC5la/aLxVnnnOwW1SoGc+tPln+nT+zf42Wq
xUVkoQMUP9ik5qVvjIbkfaUy15vc90gq5UrKRPquWtTuCWr7V8IONLI/7S9j6aclgc7WKJ7yQU7O
8enwjdFn+60C53gzSgVFKSg4J26dQ7/LoAzNRPm9lINKQGI6Gcetao3QzsTjx7W+OWu+SwHfozwQ
eo9SZKYNzK1IHpVxtJ4jmPYOUMVvdq05YRXsv6iyatfQhaAWJYHHhLLKtuRWSXNhRL841vamC0Kp
9YoyVYSggPuIvp1tbBcBW+WhjXY9YRLsVX6dm2AGbV27lK9ZkG2cTcATy15z5RmzKsJ44W49jXcA
ibEGcKuWHSPORFuHrz/TU4GCpwRynRt1hQUpEbjU1iscFMdIzyVvbdd3DWGhJKfNeJ+1TfTnKcR1
gWiqkqGU0mwPhUn0xoUActBgtmZeBxkwZqA5jfPR159eGRCaxEBN2qVaubN2T/MBw4dGsQpVg2OF
RKQ+DpI5MHrU3sxEnlHXasBangENPFHyVd2AfPHnCX4P/nEKMiJ4BG8LUixk+M8zBbHrz4IalWjP
GRG0B8i+Ux/oaFp6NC/lZxnHgJjutCWHRG0gqTVxtdlL9gYZF35v2+UiwyOKLyo752gjH7Aqmikl
MDrLys2DkdkYW6CPuEOca+GfJJgj5zXze0QRPwcMm40whj1n+Ji4EziKTQ19BfiTBJ2pKEkEfNFD
gsBDtb9HyQOOaM8zukmlvOIYOJASuYM8eoaMlJv2DcOloaeRlkMTz4vUaTXZqrDpzStX43Ja4MMV
9acWXZeXy4zuQV6AXNmEeShRzYBmMSgne78rJmq2yWya3ZEqez4bHn8E9jrH6I/lkIm4PW08sI3U
GQxcIYgjgnEpNJHvKM8HaCnrIUwQOYntrqwTsQMuwhPs7rlcSMw8NwjqITGqKOjXQDNHuZt951JH
qaq4+z/ejZOvrxAeUyIU8srwixrJMu1uB1LNz0pw/dvEzQmY2lIr/BQFaVRE36SXqYH9utb3w/6f
4V0P75RjBpZV/QSKY7pPgrBwemruu5n1xVMku+9C0cbWAytHMH8+77olcuntzqTtsBpsIysX1hKd
dTRezmB57SYZHBZcpP0EvHrwCuzMtAMVTM4XtID7SaMB8/Jv4LsqxtptFELrLcycrAG8Rh9o5Gpv
FdYpKtVGWTItAOEf4e/zeuf2DBIz2AavSEfTvH4Viw2borrFld2pwjpJYCLoPURxbKBdMigg1lEl
oRn2vOQcstZVqpSpIU7kUABPZ63scI7Xclja+nborvdCfEh+JW5IlskdB3XHsf+4x+8MZ+HlATTk
MMwpuJ1c+Rq9RMMpgnJyRxuFMWCabvs59QBY6HLTRS7uB9hYrV8bAqMvqOw5+69AqMpmgzY+dkqT
t0v85uqY8xeSRSS46SlXp8qpRIpiT2oetr/9WpVSD2w6QH2IpeimkEdM7+0avkwtYXBZeNYw1zVi
MC4eF8MelyW+X6YpiAYhoTR/ypmZao5ko+dbfMOT67YUz7GTiSA4je2B4qtu7/rEyYpnuViZZL/9
X90PI6cQTR/kZSY/iwGUzGzxdXC/3/tg0V4KXxQPQauor/56j70yMj8hiG2yEsYk4iy+2Cvw/4sF
DCwUVfLf2u5qnA5HIfWuEu0G3NVddr1EADSloeEBvqZwx2K2K8oUDQpRl04xY68fwPNM2djSeYzF
lFPnG0wwsZco5SH/Gm7jp3CnNVdGqr5IDYnyO9T2DEyw03c8YSdqtexVQwHn9UIIYKQT8Nl7MdcA
2pKuvSw/FVtGs2FrW4aIzA8uKl025kLmwY5+bb9AXFM+TAD/RZgFkT9benxGqHMLZypn3dT2u1I/
3oIZ/HjnEJNQLUTqLTs/oBxwV+yIvKYkyG6Vr9zBzXrqTcGI0tK3DKbjI8/oOxIMnLBs7vz10aFA
kqHt+sUubLObq73ZHpf+u1Z+eJ0StgJv/7puH6YQEUmZslmXA00/6x1uYFASuGE5MUHm4VJHIXed
BM8Y7OzS8EFyGAjPtbvq3SmLVbqCYUKme1diwF+wtjqB0XfLfl9gfzqzJLrkjvJnc+NtaMm+X9yO
trZE78RlwI/oF3W7oPHHpDpjmysiCvDL0MI5k45d4nMUd1CqF95LH4lOlwUooidYmZY5E8OQH0I1
idyV+Ezt8tLoATZUcdqEvkZiDuyeqhVNCqGXxZFbWRwv+eKCuaTSjKAoaikobelEXKFfc1O75JzM
4jjItgbFO6fK1KG/nkGYz2Hfwrh82lI88ZcURFF+ooTqp933TsJ0qhv+XqAiWSAnEVtZTmYqGVra
sHhJb2cJH/BJe0sA1Azem/maFhwxRRcLN1v9KlegCdRNsX+FAYpyPVFdAzeXQwGBbGDJOeuxy6bE
ink8HTmxaIaWiZpgTxiUq5gJTWDxjysfVY4Ir3glpPhqLOdVrbfqoe3IqZLTxXQp+MFu/yDRd6Vd
3FkbRaF4te72TcTRqlm25xgwazFBCIVZmq23TeEFFHHc8LehqaxHsyKtlX+2n68ZXEVj/PQBoBeD
Qle5dBKIsbpF7RZapnJJ3Rp4LI9fjk6/grSgDR9np16lc2Z5d1DhbiAi3e2oanjXtTcKr06bvxzB
W31geb20Inm5MiMP1YTxlFaH5MrTFGEac8+J3y0mRE9pttXNmn4JxYS2IUljQjpC2UNtzrG0CqzG
YP2t75lfIpNfxADLnyT1TNQDlmXFYiZgAMkF8pAs8arg0LrDdNbjjhzTjQZijf/OduR8pHHNkojB
Smrs1UQX4k9nmGw5JVDzPHD3w6/ZgLTsb2WXFreK0Kv7Of6o7voOjG21XhetoHto9t1Bi+Xue7JB
lvIHrMXOj/eUeHzEc7D6Yz8zNUq96qqVbpvK41SZPcs6Gm+1oEg0Hx50zZaLoC9cjnYs2LBBnKBY
QGMoipA/pw+XnQ/bxXjFIvH8s+JcQ5Zp18tn7zZg/rjG/KfhXuVuYM6i/yhNQlCN75UQP8uLQqi0
sTxLTXqUXbbtmj1epkeDhGTogLVS7L515GjcBal38AyWJMqRWQvRk/blvRI45AZ3iWis4BFAYJvb
8LoTQ9sjfu1Is9V0PbXrasqrCALkOnsp33KG958mv6Twf+57zWHovurrtKlYTZZr7lhbIJCmuD2R
Topqwpzv5Ayy3UDgUuV/cwYYQT8lcfKwJNC5yX2Otgs26oU3OYxrR33paVmzzlobsgwHHGOdBKmx
hPVZplKJWIAfOxdXDNT4+cckw3swmBpC+FUQI3nKm/rpaz8l+rJdBDHXXe5HMMCCfPjd6SvU45PJ
oDs36oAFhGfhQ9FqmOGHkQRpRz2/64ZtfGRHpoBDQTqIhd/slVM7qruBD9LtiXGCTaois26cINuj
jcWSB7MfIE7nz405Wcak1GmcTlyA6gDzmoMLLXMMJlS9RK1zNxd7pnvib+JAeMG2OpIXppHAhPSw
7pira8ns8zwfUJ43gXNKMiDv/l3GdJhZAbySBuTNtjrBHdggzRiLPbVzZC69xxgzxO1W+BtmdczS
i0nFOCDTkZNjdgWzg9gBoStsuUGHA2Urru49HCBGRRQQP7+vcHx9e/0D7kZ81LTHSzd98/sgbYn7
v5PVTebm/btzXhyeyysLPuE6Nh8lEhxznTgqQTxB1RRM4tHoZZwmnX3qFfgp9Dsp/Pn8T+ngzO4Q
DsqamC20LGMlN48/0T4b2x1qkDr7cm8+Hu7u/Is1GGz6WmEtFi1lm10tX/X/miXkZPZsqjsToMX2
fgz8R05cR4+jrf44n2Pml7XQSziN3qMVXpk5uHIqRFwkH1AuiGvILFbkS7Nwf0l5IVSUmPTL1vfQ
EwtvMCCVaZDn2EQ2i2jvZHnAxuTJA2FpNwDClAhSx404OJ5TJSkJVM8bzkk7Oy0OCKZjSPL6GiXN
zy3US3pHG3N6E2g19lJQ4lwls7cy/k9Krw7qnGQ9deVeaJH00VaQlAPH5EGwOeJJmlIvDcDnzEw9
ZfFwRUrY+u2bBkbxvt+qnlb3YMSTtnwWy0JcbgZKgEt4pLIsxtZrKXlmPBejAg+AuDf+JfCpk2Jy
i+dX2yKEYTgwNhqmsIJ86nkhHa0DM7c9zh7gpQ00sMpyf7u24UqYygqHfMSnvGHQ2dGsfs1iQcy0
Rj7wrSCclWH6GkO3haEkloP6WV8FiF5bjSO3cgwkaL23DCakQUA6tY6PLZQAC5oaUeYtvS5kjKKY
8cMb0y7K7tmze8NAtTaFNdVi4dv3pdexrzvaYlcIdyR/tTGTtJ7d11+C4Lid14qSD7KMsVbU+zZ6
dcHvRjibMnoqcYKTPt6il9HIqMD9WLfFb9fXjG1FVX5JIXIq99dmaB1bJdZhqdLymV6eMXdSvNDc
w2HJLG5wMelpWeA05NMm/Fx+k6WcQNyHrQCqYPFyp/KD4dKjDZoUd3XnGc0pODtcONwo+xlG5F9D
ItX7H2MHpUrohv7CPTXuDMtnkJzALAQKmhNjfysgX4t2rev4lhuM4MzeUnUTJ5BU6b12brT9IjjG
FOCT0nIk5hsbDeVchFwbw/KI4LPt927RHCYSeY7ea0esAgjHnkhHTt9PqQWNvb5DifJ2UMxqnGSZ
7YoxTHVjF9f1dUUk32HgWs2dAkGT22pULkaulGbzzArSPkxa19MaGqKbOJ8mu0NPsueafpOiwTVc
xzInoREMyyjjyMaEHchlQGA9HBo2fn0KQMv4Mm9XD/TBx3LJjtHbr2edxHlSLtMs6pry+9DqXlZR
9+SZt24ahErIBjo5D7407UTkAseYu5C/c9ZOMhZB9RLuOAB7JFCFn5iXtlC6xpJceibZDfsIavgs
o2K37LtD//iTKbttbYLw67no2WqRQnsax6Ctu5OpgX2t5NpX8QXyEOeY+9mRRcoXEGkm2DQ0Vu1M
FtT2eG+d+wsJe3rC/dxOOgf/dX09DXYlLHiLQ/ogrxSMC9JcqWSY7ihzbd8GtTsR5TiIP4YTG1sU
5h3KPN0NHIj2Pw88iqsvlh2VJ16JAPN1tRordHH5yoVEWLZU70AOqLqvS8SJgz8azi8PZY0T0INQ
Y4Um3lUHIamlN1FSRrBzmPcGjIfcclxT+/TujtNBOHdzXDG8zmQK/+YYuhtNlpnOg44gyZwbPJuO
LehRbiluqV0/yOWJ1ub/zkPspT3ZrBbQx9JEZVL9NfbAfr/nmmLVxQcB7onQE/oTKBNwNkg2klA/
kOaaSyn5OVtU44P5UitO3gMZspjlEU9dtmXVpcH1JEm8IcWb9DvnK+pV1uo24J+k+LglEMjikwzq
zE8zu0Jnjkwtc8So/3I378qS4CXiGMlJRWdSgwol4OUtm1QGnq2969VvL3JhzLBDXXKvlabI/RaC
aO4pESz6/h+ocgX6CGMOWTFc+Oj6IXzOvKl6poWqBCcbok3D3cWQUx8l0Ii16/SSa+xQrsPIgNe7
utFJLo3/4cKB3vDYshK7EezIfeMonzbz/Ou1nd11JvcQ+Qu4RU2t+WCpNCR1oqXvDz6wQHv58Ky1
jAiU+fA8Q1Er+Adj4tIAUowt4tqjp9OkO+RG2CYyyYJz1ZjmfvJ18P+qqgcT/dJawrnlrQAsSbAr
Hll4y30lzW104WocMNRdW3fsrEcLY6+rtkPNes9kLVoVaPUZr762lRthRbeSgky+CJLRezlCgzgx
QsD0+y51AfzZvGPdosnGNxpTDR5NmBA4qbqywOqvejykUNyVaU1+HhMa8YK0yDvPmzZVbJ/mq3oS
RlRcgF2KT8jDeQV1ZwmyudfJHrV7d5tdtJFqICPGat8B08+eJ3blW+RldNRrDiFIxa9kYo1nqXo7
Zn/q3gF28S7P8n4beT/lV0C1CinfhUu//MFsOir2szBiOCZNnw8doZ94GNf3IlE1PLJxOW+O00EN
500b3ly20aw/Y0srWbQjTZeXaOWjQ7CUL+gVokiQIAnNQUeA/U6oLi/xD85LhdIb6fAMZGTDaZbp
X13XMknsWxNX9k+DJGLlU2NurYtVr1cn7hFMkusvlp6ULF+Cn48L2RxMzZ81ANWE35Ch6OIuQG+q
u6XzVmcnFlBnLFSs75jYToW2ljWFBc45ARmdlOCPQU8nXRu4PIAtZyP9nIvAoJY+FaziS4ibc7C1
8CbW2VvgJpL4rLiRQurYfAy5HRsteTxEAWvgQB7ExQZGRqdMMd1BDQAZ2jmQyVyI4csyPCb+tAY+
Q7T7R22fqnasCiHNtmbaCGcVKIcAoTSq0aUOXZIP1yTJcZdCglqqxrPfmykuAFNDloAIAnj6PejS
k3kFeIMS+Xii9DClqzc7Dc6mIVov63f2jFmKCyZCeCaLZQcWRMC4UOHBTm5OnT1wYrvlC6TF6EKf
lmPIwZGqvjFzXiqfD/CptB1OiabkuSDPwx7B6zZbWvVr6CnTTy2Iw/gojn2sx+vHqV0CwM+iXjHm
vsinVMYXqLfVOhWqX1+zN+dfYm0y2ehjGap/JnzzCWCyi45qOPOs1AF6My1207y1CRwH1pMyxbh3
uwR8t/V0EXIgClnMwTI63LemafrT+iCCqHrP2g18rt/4dUq73JHA20iNzqzNbwhraki+uB6XVE7C
Fb8z8IjAv5zvFwxoWM+VUl0QeFGZrZyOB0ajIAIh3+ZDd2juHigcpdgpdGOxElEEPYEDnXcp12WU
rSNJqVRK2VCATCvxn9zohcmDhxR0XWKpngyQ9BJDEafyJIs2eQ+0+iQ+YaF0QgCCC6xlWXtvTM2r
1lyJbRWRaGxgcnK805CaVDGARrT9zeeqBghaww8MocKiFxAg1xIQ6y+MoEqUyz2/gL3w1wkHvGo5
q1HU8O2NO2Fl+dA7G6GKHt2POOBWF8415RlLcP9B/ZtEW5JkzrNxdOKKAAcFqvvZCCpIeyQKDYHy
ZYi5LSMZM1FzXpCIffcwqBo45GVT1deDmhAI3x+x6WTG2uMjfxHO5Gne1RJCmKNNFg7GwHUz4Z9t
NgzAuNmHGSiC0viH95dm3GOwpoA7U1dqEl8HpnW/2KOV1mWiT1+0bEFLO/OxAYIRwHJItoxtzBsX
AQDYc3wkC2bVQwxBO49gsbBvYZNad2nCSQLwNeMhk2b9D6vUEFrsPmbZ1iq6Gjr3RHjkec6ujvft
biM5cfURdzhdvBydY9H4oNBU1ZOVlvdhVKYLRsdSQLYsGU0i+spUrYWcR9uhtSJ8Aiq2BuloauNl
dLt1jkIVTMVt+VS9yNrcmxZSKgLe2OgacwRMkT51fKhm5TviATeRISAH6HQYgxp1+2/NCm7QoCte
aviRR5LLu2nwbNp/dvHzxJrBpCl1sSeSsP+Kti0R+ZraLfa/+FrhVDa6ZtfsVO6Yb1E0myBF4Z6r
EIaA5CVFGlhjwNkAYEZamKqSs9yh9TTRJOL0y/7twtuGtGX2W8Ss5bdGbtFlkUYOufx4As6tDZPW
OsqiWX8Q3kn3BaKbsHz6rQZpkCcj0yHhCay60aAevZZXxYhItWko9w2bxrD/R7Mv+aqs+7ITsp9J
nCHVYHK/c4YEnukIVIycoep/6ZjOZeSGtrC5fEPMXPmmW05Pdxbe3tU9U6qp0KLrO8ULW4NDTe2X
et7zY9HbC9sU/aBT8mrKqgn/q6mnP2Fj6HgW5VRsQEaML44vrW7olmbH6T7SI4HT/8LfRSMlVv09
fzES9RKk3pk8LvdnBzyl1hKuqI4xI+klq1DNZBx6abF/UYZy1HReIkLcVu0aeJ2qxTUrphVW7B2S
zP4ARYnD5gbRvLC/R+CX8CRMHjUgrMAtBkMCXBJrj7kO4HgfrSv/yiMonq8ifeSEVIb5RiPFeAnf
sT5lF/BSXQ9CQPSRFCCC5DA/juLqp0RuI+r6m2MyKCzf+Tb2WFlaPUpDRU8dkSyLXZFVXLgoP0sZ
u151ZgZn3IJXwDuxaQqirGd1S+7BwEqtxlGJVhGx6p6s1HiiFOrWb4Cl1GisUfk/Z+Gej1pSqepb
uM4MhsdY8FNRM6n/gxAqLqEnnM5NrhfI3YRqtS7BdfHULYIHxXrNU8fTJ4aDIkYH6cMYUebKjrLH
t0fmzRBINyfTq0K515l17MyoG2N+F7wwKveEJujfggIXKooobZWDOb8+AWq4rxg2qMiQK6eb5c7x
QJf6ksVHnrInbp6yClbk84xFZC7leUO7cNzeYUOKpXlU8SI177fT2B1m03X+55KgfSyYkmp2/Df4
fR3ormkLLu9faJ6MFsfHTL2Y80f0eoEGVJXIHTZg/Kf0DT4IZi3ePEAqKyMIbhgS6oyVBucdaQfy
ndp6ZbqsMjxzh2fScISbx4DWbuV2vLqmO6oDQesLtTfwFT5+kj4aLq26eJnK+hIDqyw66O85dCqE
xNNof87Cz1j2Z7CS/2zVuwKbVUMHoqMqR8fmokQVXlpXpWweBCaJrnCc0n0iPkDV2+dHemtx5FJ+
HmeaIsIZzvUbahaD/IiKz1au1LYcyMU2M2nG2hjWTw5wlyIQvnTveGzQOK/b7OvvkucpBhWnXWMA
64S6k9+WvUzso/q1AnvUyZs9IjcG06limKAB71QZjJqh9HQVHd5Elc3OZitGQi4dQB/eYUHVN3X9
ZvSiqvmcsaNtuoqHodhAUH91grxPZW8xGvp9mBbLYPhtun3obxquRJBi05JvdSB/oO6GNefY/jdV
YPGKz+kW0oFbl2jZOse9p9VDWEJiglaPTyvM/BFcJogvUk/QUecUKYoKQRgcvrSEQC73ZiwUHmBs
/Vmi89PSbjpXzdhIFSwBFhvHCES8e+OWHtjdgXTNR+hSCBjt34BQfEglUkWMCEe+h+qsk/+54Qtv
vSlK2OU5vaZIf1w8/InwWKr4GPibDLytnp/vs3kz8Yp2d4BWlKbrwAi+7RNJwbwo6jLqCPjl+5SG
yivmsUH92U08ChtxNRK7A247YxGArJy/NZl+QtN+jmi/GQP6A1Zdg2HRS307y8YZEVewCuyjyWuU
YangPQVcPwxoQWoDiK0SCBuprUmny0Sv1eXnYzHzzecvHmloV53eBndPeUl4CHmmIDOupqI43aTE
GFC4mqrLtZcIfN+ucRdzHwGstbmxGd4zqeQsXqgScfDnwSTWklxm75KHh8c7u6jA7zFIYH5v1UoE
nWCO5MT8Tta9gpihEqpVkH2FanBbMtXMsNvsE8HsaeBx5gtI0z0g8uojJJyiwISwC+e1/Jw7KQoh
1vjIc9FnVuHCsDyowsr+IMZH7Ju24/q+Ym0jvHWn1UlkcaPHJLewctsit9zB3sjuinGBeEIV99Dj
2b9Y8/3IDqY2OMFshZhZv6yUIcB8rBqZJ2YYZN1ZnME553zw0ATYieHEqlyzBUwdn6d+2k8a0Is0
4bx+vRcDhbedFuFrhsw2FQ27ZyEq8cdzrAftrO8+3bF8zElJ1jV2RZYNFYUDLDvY4vPT3qtFMeyi
fzmrPwDywciNq0QMC3eKPxRILZr7C016Z2u2RxBss4qahYIWOgh0yaSr1qrM1N/AA/URS0fbLlN1
f8tfaBoNdeHcdLQ5QTvPPh88CkvplR9ETLTyJgEtucLkyy77TW82f21P18A0E+cMvBgfSAI1yRHs
j3GeALILDB4gBTcnLtv93oLYJP2Z/MXiprJ4TfBjtovms5NRvwQnmei8CYx+K6QudMAeMOaoC+ay
yfY4/J9LLZP/xOcrYyW9yxiczFd1vzMZFotMtkkzER0YFqvXJlLfeZPxP22ZFukURAIywPnmgVff
8e7sAhk2L6JnqCyNnIRDZOF0hlBOl4ex5DSJzZh0m7nFpX3etidF4AUfEzciM9pfJP8EURH4YEdo
lWekXgYKJj59YVeVv2bv5bqGdumCY6kLwfL6dE1VUXOs7XFaeB10G1Rr7rSngdcXBrqfp5ZoXod4
0bJrBcibGnn2YxSLbyinARVaiLucgHDlqfU7TGH0Z02Xu3z77f+D9CN1bIDf83Nnru5nKmy77hdW
K+jAR9QBz+p7n03r4nPXITdjP4FzXv5Da5qSn7UKOhG3ArxhC32SeAwlZsXaUAHWVTgb1e6RuRyU
gFSsttJugUJJ2i9mo47SIjL4wIg0pDgTSa7+pEHXbFQICOwopJVcUEmDTgQY69FksgC5nZIygj9g
LDVL2FIkLbGLXrCk+1cW0+H22bUx/L4ePMex6koScyk6J2x2TlDa9Ul4aOrgyxP4IwCBcG1/puUl
VykuGQObg87U/8Li76L8lsVJEr0W2mkcI1+X0UBQPDgF867CeISTpNcdzz5bTNOGxGtxTWEXFrYS
qxYCJQ+huAKopcju2oBbJGfdzwrthE0Cyr1Ku9DHt/vIaWj/SgbwtWkefzNKynUT0tp2utsai3My
2yN02HG7/Kf42bMHGsgoGZDVRTTtuO8Bxnd7wFTrV2xEQb3oBIZGe3AFPKZKq3yfaOMxIxJcuhRl
4B+X6HnxTuUIfi1qmc53tRnX/Ip0kA0Bb/YhUoHdAt2/h0h+e3/WenPt5dZq/ki2L8Hhu7NZ4NCX
5BVhGsiPFkksfexOTEydnVOLTylu98mzc/dvWvuqu2xZP+x3s8JmrVX+vUcjj9i9Pn++LDnXbGEr
PILQ9T1GDm/pOH+sFHJgUrvSv0lZrusU+qssV34htr/WkqdCslhwY5q1Kh7gmEtbZfLtqsaU83ee
i3ilVz1IeuUpTJddHFJ9GFFftio6WzUnVz+0uEOO75uol5s26UgWNnRb+nRNLdfFnmfFAhWGWf3P
L6vP1Rm+ovhmqGFMLvrGIKvBu9u+F/qOhpQHOClK+0Ivt6N1Mhj7XNDZYnlm2wLxkxlzaKXRYleL
HISyA1trq7uuVIXd4za87rhxB7I+MdCYUEtYE8y0/RbcgIGDKv0JxSWYHcKTHoZFuBBbHFtqgxdz
ZNCdeVnWCqSPvp86RPB4/pQKMSr9OoSZvjLuAex7RFz3h0pumGqdQpi2MH6T+JbByXisoqCt0wzL
dkXjdpBbJemBkTXRaWsZ+n4uyZK0lbzp/n0X1ci+mysA8KlWeV0RiFZ5tTcjU3tHOWwTWF5hHcQW
cAV3ZTYoGUV1FIbgYFVQXWdWHlebr8PXLZ2GrmPiXromFjJHL9sKIgIDcXGuyDwdb47LGjcA2Btv
k/rD2pUhYF5K+LjzKzhZ76ALCfMnipavFAtF8RgdJJuRvymlEuGPrGGfqv/b/pSQ4tV9DBJo4R2m
+xcqI37W2jwZ87nRYbgzngBTfFxLdQI0V45naPSjqWTJKjGwxn5dKY3bC2p6zVhEvfZVjkqrfc3+
hPML6X/2Qja1tLZA+y912nK0DHFZT/VjRMjDcuD2OcdpLD0WlFBHeiakSl6Zw15IARApCbndrxMD
oivAxirwXHrM28Nziq33IyhYgmR7kvQ0kmZpkWBfRXTU3H4vQB5Gdp44RL66p839b9NpT30hsKV2
gi27xS7aR1aj/K9AOD4yKJiSt+SpVlr9EvY8rJic78PuOuHvV0ns8PXkZxsUuoQkecCpXmYgepbM
oNxCWYQ2zLwza9W+k/3ZM/23TpPczQ+kCBlhHVfTYoIlkpA1oCEReXgxbvibUQb8Y0Jrgc9CtIr3
bXALSVmcZCcG0ggWSXXP4GAmW0ND2kswlNFliJl0LaXGgxDH5pFq8CYujig62eWRlMu8BMwMtMjC
s2sSksbF9TsSZCAVEiX0EpQPkPu8CG/CEhHV9+kqMpNYsbSliWsRyqlGFvz4ziNiRwHx1i8x7MJe
tuIxkKBbC25r/Pe2C5OMG6c1HTq/gYuKQ6cRqyBsV8MX8KlC2zGnKjhwQ4MpOWqb84JDqeP0d8fp
C4SGIl0YcYiImdn1DO9/fZrfQyBYW97FXGC8JFTDIfUSCbmiiIHv6m4HBKo+eZOTCfv1BAAuN8Jx
trGbmG1bx/zxXU2HDTP8St+i3e5GPrnts5lW/abNsxTofpzp8cnZe/yD/SNzJLE2oRuloEOkrIIp
2FbOKBoEwOGBaYNiab82xLIAK2v4pM6MuEYQ5jSg94HvMCsQ/v78j2pVpnkKFk/85kEjX+myzoLB
c3i/hc6jxdG8JPbKkmCf/QbH/U6cNjg4PG2P3Jn4X1X4AvsYGfcNO+MK+bIBHImcaZ62Ic6e7csm
GCpY4RrGwg7EhI5iMk2OstjvUXX9yP/4vDTcHsDL3Wxg5iO4dq1bnKXJQKU/6/MLJGi0HINqT7WQ
kCSeGNRYy8CK2V2F/gr6gtc/diFregCy1WzIEkWa9p04ZDkF+RMhfsWRtZy4Y9CpkUnlD3b5CKyb
HAFQ7RCgFq/Dbn6F7iVDYHFuAzVKOODhAmkCcv4TYz5WagM0yNN7W0GBbxL+/KaEFgGcXsOnDl8j
+hg80gLgVQNtl879EV0p9FbscYK74sWu3RtS1oCwuKk1fvx2MD2VwtSB00ODamgPvda+8syCowhD
M2POgasxkYs69ov5lMuo8oCifM90qyKokHL58lEOu8KDCmXL80vv+vz3kext8bZHfcpNzHu7Oqvc
UebYfvRQvLbGmQalxQu9/DR3X9byfkDsKtFRtux+wSh2P92B7t7w7cHhGlvsPC2Q80wTAX2gpK9w
lGXLaS8Hsu32svmdXtNqYZRd2TR3GCqZ4w/T0rnWhN2vZonmOagwZ9Yq8hXBjCa6p22iG6o+GCsG
itH4RwJL4FBqzftFgJoMXfOaTlO/eoVSy87YAeiwAJeuXjGSVoNYrY4r6XlyAndnHnyJM6/VI0Pm
yXmN7BV5Jd085l9UjJ7aLPvQwNDWGxxJD0x7LUpsGie49vTzY5itEbmU0l9eOUjwb1AW/21IOd72
/8it5HzEzLGhN0SH6BClxStGdOAxN1HopkMYcnX7iSxJDMSOKEslC7EZyexbj3LYttAmbk6MEfzc
0CYQA08DwPvzkw1XVKS6d419ONrcmWd4ZemPY5+bL9zwKSdH3BaqyiiVGr8V9a7EWCPhU0HLnE+x
V0Kcmxl2Id6AACu2YeW/yTnMDFfXMEhdJJ+FdDa+aTJ3JloHqpkQJnoQDfFCSzhkcb2GgBgsTtA3
A86tfqNGmehTXygOLG0PGWdtJ5Pf6JrdCx0LIiCAg/phRHMlzrgFs5IB68qU+/GUru5aToKmM9n1
z3nUwJoMooJlA6nQPHqaTH+iHQVBa0nPCI9U+9Kd34/lp05KegS61LX8C9es9sJRy52caNdy9ZYg
lZL1IMav2nLmDYqY6diKwNky/Uy3l+6wCwSuz1vgALBve9HEjYJHgYGi9hJ+tCZek3S9cC8+/L+C
B+FAj19WS4yM6Om7+oHrKaITjSzUhVP7mYMjMKah7O7BycDTdWjPvCTN6zz9B0lgex+flTnx8fJf
xNgtxAavIELTuR1hS92EONA6QH2oHjVdKFvyBN4y9HnI3DC0pDmXwLA+s0qa/PEeJCgcWlW5hsGd
pqEkQWuGZAaMtg5wSyETvLEtC+jaMTsaZD3BWrQE0YoxB7sX0IFLtknGjg0h8Fa/qf4XUy17SWwz
ojc8GX4qIBRKCtUS5xfrvjyfCbjvvj+eGRv1r0Zb+hthiCGgZJ9pZQKpRjUNDJg7hOdWvr06gVE1
+Tw6VoyLaLfF+X1SP6WYo8tgthKBxox8cjFhTtgB7CUE/cbKygyfGy7TbMVL8PDl8c1So/DGkIw3
tLt7nWjoKLYv9P+4M/ZT5Is/wXplQpsM1/SLz+EUdFylyj2X5vSP4f8mrOtmJxewoGWAZLlvxM6C
r8v2BbFYOf866XN7g9MbtKPu8HSs+DvHsQAtxDeg0ozFHJ8CGMQFkW99vX0gtZtfeOCPaAsrhNhc
QTvDVHHOf/bI03PBe9y1vKebDGtgdFtlbRnwVUdPngWtPIi1nQZHj7tLmXYMxmHXL032SRmPPvhg
7T7w20puJ/77jk1zBFDswpSKyFapoiSiYq+IMxMHsExTFWsKnuKk+Nhf0rNf3ln0HBRpu5uz59fz
HFaOjVT5Xha2ITuKqThWmj/kgTEmTVNXYqN7zWJZ1lVmF2FIEwj02GpDfZBvueh975AM4eHWXV9a
GABWCGOX0E5a1akK8UfKXr7sFfTSIvpJCWuSjueiOBLKKYtsIBqe2xfwf4ewfv0mOOY0SZ+Lx/4n
wL3BMgslP8upVeSuDdtGLW7PryghLeGEjfWvMFzd/yzrWY9G/LxA9P3M/3xke4knpyPhhrlg5fpt
RzoyRHBaCOgqenuiFjx6Gq/VdGFGKgplUKa3Mw2Dzf5XPf7hqa3xyQPLTxbmxSXsdTslllePbLnd
68H5v5uqVh8PBUVVizqiC/KgHhVf/XFQGR/5ceJaz36q8SOmiFNcunX9B7T1KUKrEBdlJemOVebN
mX9wuFKDZmS/Dpupad7ePxl1W1BZPXvlVlsWL5Z5HVI6TZXn6CGrEgc6DylNiyjsVIfRaqqrGYLy
fQ3rA+C8cStR77PlHc4mspMZ0xemc1P11pHbJnLcrX5JQny+QVRqbyYWxz8qZm/9vlRCqQJa7yPi
hEKWOvKhSiKIc9W96K8D3ad9xW/YmP/0dmTR8yLRJHyXZ9cvG03qsRRKbXXRT5/w0zNUzDyjMR1G
j7TIQq06Ax2A31+GaLGR+1BXq+v5HJJHlp9f0h08hpO1V5A70mu1Bfbv6e80M/RNZsgYhEALpAjl
Wm5yTLMKM9H0B6xmfUYyxXf+Lw26CUWrIzZIKJqk7fGbAlIH6BY6ITSYdeZ754lxvnf6/QdZdMO7
Bol3WDM98rjxhfYJtFkgmnwzQbQu95jALDDVagHLy/hodYiKtqhwCJGPtuwJ/k4p3oypfDCgBQcj
djFScoqu4s4agOa7GD6Rf6jDt/N/lXbOIfqMmNYJsi7RTlSVXRK8gdlIpsFJZu0E48DlA+rHF+k7
XR+nMS2AjVkATI879hvKphl9NsJjSOrN3ebaDCfR7nnFkkxJG/jOmK/0Hxtoz4L8Ob7oDxvG6cXR
9XoiTun8kCeGzO3v3Ir9mGS91h+cysCid69Dpxwiqs4vAkuLadOYJSzIhdKuzX88xSRatefds6NQ
n35UbCCdidT7sfTcEYoS9xQ6BdEys+tayINonjqYNZVBJ7KQYVi5w8E8boy6u9gaJR9MGmha7JvK
B+Y+4ftxN+5XATAK9o/QgdPl9zvjytfjci3lePGTxWApma3DpyIU+psL6WkrA+bRuaNyn8BFz4B2
VgMggPPInzCSjk7zj4JJB7uVrfv8wstARXB5emQ6ZCu/zlrIj53fchOCF6ibcGa50mVdL0gF/nM2
OxGR2K6E8i3T8tXy3aD3zXHhqYKesthzRaHCVtkPSdtg9p9y5mQAOf4esnD0r1nEPRF4lt3L4mfb
EUN9EqdvCUiy7M2s0LsbZ8XgK+bmI8qBtrOR2lZ3/s40bWJmsFOBJ+MEnveB1TPgcR6D7xKVPTJH
RkT96cXv7HmYIYIsQ6NmwJJuFRbXVmxKO1TYgztU2D2YJW/0aaYjg6loxcfGtA9yPwTOVGXiUkg6
KxjzXABowZ5ANUwasU5W3t4vYoMHoY4TlQA/u+PjtfroIPqhoBZc9L39cpbZKNf2mAk38Tx+SR8S
uPzvrgn4ZCgVEEBApgdvmi3mfopzwzkUqPUk6SGmA7SmjnHyCPIQf51N1PKyc0lE5S8KaGe26kKn
7aJcSzvAkC9iBbO0ZHydk/6VEuTEKh+TrpD/0Zmb/LCH+fM5c3PckU3x4yiXZ3niFMv6T3KBHjOS
rorW2uB2uANoUhiGDqFMIsrOJOrtXEZFb0T1DBRNVFzlWs52JZHY1D1RWkg79Vhf3k+sjy4j+j0p
mqrA//rk1Uj+CGJItv68dHtVaM3l2Etq/dwfqulUnYJjdezkWDTAI+svyzKomhAA/Ash+SvJ/npF
uPBV/f66TlvlZ8SmDnN9de4i0NH7VfjaNo4xL+QqXgnmc/P162ObLKmBVYGEvCVbsJYCKI3yJ0Xo
FdrniNXTUoTOLX0A36PI8HTCBAjWDdYPYRwACPUfoew7NxXXpC3ST4IkdLd6ma1E//moRa6Q65eB
0niPAzzX4sRxbjaJaTSK9i9AyRdsFpR/bnXqTSNZiZ7J+8ViMcIe/1m//V/UxvxEsOVYCASIF9Qt
yJeM9Wk6z/jR8DIrxyEdDGF30h/fb05X60H0Cmxr6Q1oJloxniLgL5nzLhE2vKQ7ANFh/T1FLYHm
R7lkLt4vmx7+Jswr1fT2qYSYM98C9oubmKY4+3s25klkq2AAeuTnGvXHmTnZObp6/6uieUEhdhcv
9rOG8RfInUOyhYMWXQmlpYahQJbGzc7fxyjRnxhK3ZmMN+JWBl7BDE0EyktHq8u2JF8XwVEagQG0
qfzsCZpSQRyrvgCNyX8ukdcyT0h+uonZlvW3WQsrbDy+x2KOmDcdvA9rdzc2JMPsFyYOeIcUrHH5
8bDy/tIDSN2BYhRu65suDASkCi2rC+iPJ8kHm//bpOE3KlySNzr4QlzPl2KyDazMeAkmsO+m1F8r
hYegcDS8224jpuQEiSOqeVonc1SZPe/o8Cp8PhwaBzm2q/q2KB5fRevFHclIIpSXRjwHkd971fDm
TgUn8FPbCAmzjtRmsxhoD61TugHoPNCd4rkmFFpX1mNYe78UD6x2jz1roGVymw0zAHx3Ba7CK0p8
X2TweMdE0bEti4CSHDI4zbSS8SK7OdjfXzq6zO+SuurC4a9VYSYsqhaBb8gwFxNYxckc+M+h8vkC
lMfeObfRd8ffI+s/XyBXrysiRIQ9Flw6O5O6i8K2NYZ2wC2w445ch81JTckwDOfYhE+Ij4yY/al3
oohzCP2OYBZqPfdQUzUXyI3ys34fN831pY7rKZ7odEa/GNPz1yAdeMJGuh/2Vtpy4lKqW2IHZe76
jYcUmMPZ03kDQ5AAKORpFCABo85ASqS6qAXpxm3VZoTFnaK0EeQjEhfncGLIKfSvArHo3jmb7an7
Br2gFX6XwbSNKjFfvbooK3r56RsWBOAQPfsr/uT4ISK7TDiOH6oe/bsM9UgaFt79llJAP/Zi+g1s
pyXSBGY+55EDHXTlXLeNhDZvwbgfJVdmlAyf0tm0R7WEJlO6T9d9VAwqOs/l+ZmVbnk+J3AHq7Gi
B/Sx/ZaFEZuOZzgQP/mZkS6wWJpViIVqgIVCWiAQ2TQTSK2n+5dQY3BSJH/vYHqmi+/oZPe/XQaN
t/YUMPEv1YGHMtQ9YDgxYFqpJF6lKxS4R6O8vL8TdesIKrJJNUlqqL7lv5JmKH3JcK04FWrOBY0O
0MmPFh3H7+aMVKIy9dlYa3aA+gbQoIlwe6QJfSGuIYp7xTLvodIwaIrYEnUp0cEA9rZF4IA9c8fL
ZGAwSvb0MgFsBQavsF7nl9qRLYZFDrE30dZyPdvXZwz0JQx3X4Pnie8HGR0NvdmEpYpkmnwYMIBg
HcqL8lC9mnDQWtV7YX4ZkbC5sxPa+q1KUjjA5A+lMxmhAShpYVJMHuPt0b7imIwJSoQVLxp7P7ti
a9YIyvbRFhV2jk//8TVlK2oxZNDoCSRs0jHEv1QZyGiFEqrgr9Bpn80tO4A/2e5TjP81Q9y/8Xfk
Lhrif9Hf3ucQ7M1j+FKL6nupneBhZWjWJkq5hWZ6F19PdZ8b93x6VOKdyAlBhIrhpEtgDByT/TRr
N1ZPXS34CY97XORvfifo6M0+lH6ECzo05G6NbQIBz2Se+6/XbWpcLieKw6VpaiwpXYXpHSxnpZSL
qY8DNBJAxxn3LO1QI9HlLjmdx7njU57G3k2oyrgytL4bU+dkJ6zO4J3ssKSpw+jhN0d6495I0l76
feqHKw7bBNMIaypwP2QMpo98GSyoZqMiI3WsAoXGZtf7XlO8n7bLbRuG/7EcGmuOdECSf99IhQYg
Ts49qvqjfjoMLHk2m+8zT4IJqYQw4IpZ9dbf5xH7qgVGsBEH46HZi/YyRyReTqtuy/FWgpTgbnTj
2cwOECP4HLc0ItP9TWyAHjqUVi9cL5tc7RNIRCZescp9l3yCagpPqMlt8co4FkGF5ouNqtwGbNy2
W1Mx6L7z8TQoQ68KPHcjAx6Pz2EstSB13fZwtYV3NfchptMrRYS7x+RnpPfbPfWrlsqK3SMwV51r
cQPUl00vs/jZqI9E1bZSLUqPihGPEPuKYo/9hxCPpxjAcpnYYm9zu89h39A240UBcNSy/Dk8ntV2
oOjraEaLeePo9NEIy0qmwIlrVdU62BC6HwzgN5fSKmN1eVV/NQPXoysURFPqdaBXHTgzuOH+2GMB
l1fzWL+9QXoS7nkfLPrO7dC4XkZHczFoV1G5wfahgkA6AMwuSbzzX+5f8OaN5NrZ4lTXuQdRExHi
d8kY1qrJkqJDAXWyMr/xmFH6hP3K3RIa2DMjIb6FoyDUa333sNUTfg0PynGHh77U8p3l9WPV1rK4
h1qUHhCJTeqf3tNfx2Yq8sWzhJ/CD2nHd6YyiEinZlKUvWp4ZKE0xfAMJYePmaPDJCdBUhvsisYT
HC3VR2fTouIWB2ei5318o/5UMp8gfdzAqLhM0R4AAeF1EmlpEz9yy3XkF6sZJ2zPzFU3bgQ1M1SO
An+FT+QbelF+d+5tN+kCOxJiyJqKPrr4w9KAQpB33H+AOY8kU5+B8ORaK2zOU+sVzqG4kOO/c905
Nw7stlY9XVNtp5anqb9xXCvf6y/7Tcyn2ceaDbCxEA5s5cIA7jpocXzrmZdQ6fDEpQfEixoVUQxn
lGOPyU2lmrR8r7Rl+/WTVREzJYwG57rhf0zfkBkswHVwH1UUVLhg6kqqVpArFlVBM7gDFy6E3n6T
GmOV9VSacYLr9PnEmzPdgRCuULfo6APslYWPWo9EcBxIISxcujlfo2uef3XwMFZVYK1RgSNx021c
D81c7gIhvGYRxRANL23l5LNor9ZWwcuwQ/ywrigkq+NQ4Gkd+Kmqnrjv5GPNVENhXQJ7RI3aFBTo
d7kp9FZjmAtR0SDgL42+dJMlajeeqfGZneUe2XoOjq4GKV56W2H/rP2FnGn2tFkF1si3OyLaSvPJ
eadaDIONOSgrcUZcK2pHmSfg10FwOJsIEKE93wxocDMFA2zLRm3/NzZd8I72+PoK2LVXiSpqKB8e
71kLNiAo5ChMP7Ac24CNyYvy/HMjUTcGhUX2vmko9fMT7xKceAKGK975ctdW4MAaK/hhE66Tn1/t
zAuvnHlWYubTEfXW2q5wsa0Aw5viQ29q/abilAFycldiLwSjWi9DevKyjl9kbM5Y8R7nhsCIwnOe
WEPDe2gHR7XNUHiWa3WkcRJGyfNwnEdJA3d/jq7UNv6yDx3fOcM/zic4HWHbGCBsQTMjLFvqykxo
3qiYLPvPIiB7iomz7zF0IrouAQZXAIxoHSCrjb/FptwUC8Kju8GGNpnUCcZi47SGE+KpX9X0UAGO
3owDpbnYWZ6johe90ftXd1CktgixZUEMZKW1Uy+kjIUZKQ8s2CKynndeBSZLG/EnhaiabQbZmI/e
5lPz3qM52mQScmD6FKsskcr+F59BlLI9afE4o872i3/dFT+b3edIZcrZyJfkxgzg8Kuafs3kc8TH
qbcAr5alAsKY0Nabt8EuqHhNhSm2SchgqS6CfohIurxsMZSLEWlxNs+733Gmd8KtO4J1R2BaPPdW
FttNkLJx4FRxGz1JULSISdHzBaol0lvuuoBcG2HoYBtqYQLa3dIILYZ78U/FvHdtBgrRTe5y/tHC
gUID0/lTP8nML4cjMJy7iMgUnEDBBewF5rLh6LZtDbjhWqx2YfxkPMZ+yhuuVmgjAZuJUXLhAUS2
9OOjtWD4UTOdYw2dqff9ofFm/YnoC9t+xPkrT89JCKl95t5btmAJjUkYOCfiMxkwnxPdkBZm9kpG
nxNsIW4IL9lSPhOEHBTYuLTcgn15yEIcneUx06ctPrezRB08ynCGt0IId1Zri1jZj5oSEfPkynnv
pLQgVNPva477xIbPvkXQQ3aVuBAIXK3uu9dbFJ737lu5UWWCXJsuPt1b/1L4kM/Hfzug+W5fT0Nt
SNBgfQWO4SmipDEUNKoV6clPdo1gb0/+3a7biKaQA5gW/CBwrcb15+3yuuC3214gM8RHAqCKuCTj
wTPROMkdFbjkSQKu6X5wVdwq2QlSIfhr3VMVKBmCDzncXcc5mjXuTEhh2JoJlC7OGyt3V386EWu/
xDKuhJLuZQ9D9SZNy2EuKUTfjNMWa2aPGLrOIq09eHFBUsnGVTuAdvcUHllh98P9hCmnm+cOpfBp
sdh70JS5vf5sn1eWriiPHwqEh+yzEu3h1GdSzQ9iFHdf9CpkLoh0rK/b8xP91cwPawKDfrZRMWpf
vST74qDWyVh4XflmRK1VTywaf5MZwO8d+CGb42AG+15zo4upcgGoMZwdd0g0g8xQS4HtYoDiXCqO
ZTqxDylO4kmkZ8cGf8giJtVBPeBOZbLDeoImBHCAtl3VLmdI+gDPCMNBBaVcCupnlH3lfqmcKsaG
hekh+D9AWNz19x0VqwJUwFJFEtU+Ylv0Wh+o8MmTmQFTa25d+nTgmULgUPRd2em2m2i0bRWLViPB
pQDWzyxFax60QZCd0vP6pwTrDUmmdM+U9i0B8++O73ziny9s7nQzZtHfl8gU4kBJuFQFzwhWca57
lVYP8AUjFX9qmP5r9236xaxMK1kuAAriAABsFUbUeE+uB/5BqVn1VpYGoLL/AJvG3oKW5hRBVIhp
ZctwHSl8/291eFiGIPiPwURnAjPTPl5eohs7P0/NquNnjyCYdQiHqqnBfTMPzgOK1pufJ3J+Su9z
zoRnM/PHOZ7dnSNN5mSNsbUONCDOHC6ryoKs3bs0Rm2RtlOQ0BO221q5z9FzPq7Xdu1R/UWlZDOp
amRAwnTkJ4EFIZOaGqNguA/SdJu9xzhPc51u+h4v0x6WvfAiJLzQb2ygMfB2k0JkbtnTC6jbt/V1
0TbKIaYq+J6UJNXzzOlGbALqecx7LwLdbuvTZO8pIbGVN6WTk+BmryjWZW5g2TtjeBlkZ8ba37o8
s75PQosvEbc39CIrbmRc0fYzE/haM11MwQ73P2PMY2DC3vk3V2PxqLHE9L5PE0QalxV0RzKtFLuL
kN3yldscOLIhO5RUsKGvLIzt9kqgJiPrg40GR4g69O2CgydlcryTHfEAr0tB+DIY+CTfSnI/vU+D
lbwAmzstET6ucKBUJklb6GsNZLq3yMvJrkM+EAaeS4KlDYUmc7TaG4cAyrTleEIbH5uxyU4US9ky
QXjAjpgM4HMB51icRdy0H1E6rYNRzgGrpMDA7STihaw2jlZN0Om92QlNzpGeV4/Yxfq+ECvQDnAp
jUizrPTE/RvLm9ti38qHcCxa0o5pPkCOnnr0gtNbzGfr+VIjg+A6sYgGWl05ycNtkdHt94AgPSi4
M89hADn2yhy7ItGJOGG2j0smeMEc8gWNMKxAPdqi6ZnJsZifp/TQWYwN66YNChGkoCc+PdEIzdSW
XfFAsBYsseZG5kWFL4ZWT2ozjZx3sZwvNHHV+mxObzGCI05g+8tmC4j93bQ5x5XkNytVuSXFD/4F
zFNt9LAV++VAvtqKra4ELMnTvbafO7ICnwOL5T5nMBuAQoikWR5Kz1EdnTodQ1nZ654DqvrIaH9S
hp05e/K2pgdp71xE/kBNv1WbEUshC3dytf7ajmgOIcQG6bbr7xtEI+m+lH8+Fb67F6jifdmUihjd
1nBu9oe7dXRMnrKQZMbn7Ox1RyIRXDDwgTsDJv76vXMiwrBhaZ368xQdJwNQ7UVijpQztKWSZReR
vx6ZX5IrQ9SqGZdVuqfpDD4rmMngd7Qde8zjy2p+K3+EfRmlVwPQrjcOKtF/Cbxa5ylCAukMypV2
H17iRAXDLs2WjIBITdrBAIsn5KyxCDUpyxxq3SdPINz5oLaXf/579MkASxcm4O0y1jgbRWUTAK4u
3RMxqFbppW7ehUKK1bgpOF3FnpgU5FnjGmQwX8k/69GzXBcGaCCASDmy+63eyZIx75FNdZBrsi5r
HkyGvDt24Au5+piATZw4lUBiFYnqiE/3/oKW5eX4WgWCa1syibe1PZ0UBt7eABcCWQVJ7d7IppeS
TrjaYx9iYXwPHnUpqhuuQXxUDB4JeaBcajLoU8TVlNyDzA2AZ6E3S6Rgvwz2TJ9r0C5L8G4/Yfrl
cz0NQfJ7fYtAVGB+P+G0yUaa4mmmMEer0NwjRbDhGXuQ6KpBkB+5iqxBb0hheQgz/LnDKu0a2EKB
UQjknthc0cN+oJOfTqN4wfzRT9I1OZEC4v1+Ky7k9V4J984ptf5NMe/jQ4dttqHImKzZPIxLrkHb
UR49jRw6Lxnk/Ys79ICzIvQlXEVf8QtlS4H9eI4uHC3CjhlFoquSu7JvK7K8Vjh0+YzyZ8wVpbnz
LnnmSuXyZaql1wrKiXXKl+FnkQk6CpvwGiTXsGwjQtOv3sPrykear9zFeH71jOKJeWDQnUx7OuwY
xGk9sc3XDlzc4hobp/CHQwaNy+gpRLzPFg8AQsra7I7jyAtrhJRxZGnWjZPTf8mLc8gpqoHGfHEs
ZBe7S68HrcltjARQT97cyiPwCRQ/8+/xDlLuMWwgZFJ78Ti84U1GeGpdB+em/1LjDTGOyuFcFwsF
pIaLv/vhURCqNY2eaXLPwztz5fIcQUK2HLbbHzzD/sF6QilqQ4TvQIGD3paq/9BBolng0rwby+58
HMlczEOsVS/9LRog/bKUqAIDFhFS/3JbZTBmks3iA5kSckr/zBSab9XjJ+wom4mlybnvti4yCt/n
QHFFcrFy/Ae3Bpu/2gHud+yh5eR9/ZeLLKD/bGWmq9epuf0hjyQjQ/lPTraN3hwR1olkUJ3aTJLS
t8gclyICn7eIAQmW44B03vVcRCbnfvMyB7O5l8+HtSh8ucI7A+2KSates+KtlUvejjZxFBc4sFUI
5Gu3XHsNMyTJGZLul+xu+Y4EbDjY+kNZsbOOLpUiR7/FQwPs18nLjy2TW6Fdu7QKakvWMBCZ7Vrq
guwI4CaASJAMbLy2k6tN6a6O6ZXseFD2kLJWAtRXeLjvEA1rG4zQDvjW5T9dHUMkqsZ3dWdJ+fOm
TrTGACe/sFvuUVTWEQW00KpX03bUqzzVQTipa3SFM1iGPFeC9H+ZVXF+9/gAYcBEN6ZtTJ8A8pSR
XdY2Gt5l2CxIqhMgKzL91RzJfgGdkpkNYXZ0fkevWsZ6rm72Pv1KEwzf+GrR3WWKM5H/oQCSVBYg
Jp5c32UvUiwrjt65ggD86uTHHydkfrEaKWkWltEXV06OQRGb5TDKiVhX8X4JSEyyYDg6hAETHpHC
cbcN4QO1tHIdCnmy9Qllpew7kqnof07/iRTiaknJY+PNWMNSfz+QIE4VAmD2VN1/SZzWSRgXH2ui
RqgTupSArNDqv4rrDZhfj8EfuUhp5BwqXzOLB1QtwkQI8BpX16KDKlWUTXYgJjm6PSf40YFrKP2k
6yZ8YqrKWCaaYCrRELP7RZeCe19pMNjCxqukxFYsmUb1RRiZ6h7Ceb/zDKfX/t0ASeT9/tWHBkah
GtgLQ2zPPZpVgn40sgkAIzM4kQDkrcO+PuZWDO6FteRpfPa2XQPIDt4f5iazX40V7hMmuEIHFLcg
Ac14aIM4UXtYOj1eMtGagOlGUWsPJPSufvYDYu4KVUS6XJAN9SIbL7n26boNldtyMSREXrUOl768
TewjU+aFePyyloXNGH41IIHBQw5M6t1rhzBwGShiH2p3Gwai55i4tHVtPwkIwaShU+gihImj3MiT
/y1tYDeYLoNl08w6we+9Uq35e0qm0i+kGZDZrO5sv7okIRDwk1LUHjXdzOs+zCp+2klvQUWk/hkR
4uhdy1C7Vqyzg1pG34JDKegZ2n2mnZ4YR9yMbp2IBCJm3ud2UPDq7avlnw5oasp89qQv4eTPCfcO
Epa7ctr3htHH7NWZNM73imxLFXrUq13ma9zJSpcto3ws0ff3fcyNycMsh5UV6AKlXh8VqUlJFquV
RW2dPGxIvvAGDDTQ3oPIzhgA4rnXiua5zD3ewx/YMNdppLRx90erIIDrJPkSeLZtxu+kLI6rZcU7
6zOkZWvznVO9auW1wsWCCugyeRPbnLsb9v2KYhvzHzcKJNGFQh8pRYy2vzzVW32vhdbyEvYKH5xB
GJch7Z0BjPcIPM9BfWPcGW4O++wkgD/73WdWWhrui95CP9QFs+iH5frBH7UzLNzyswQZsY98IcjS
Tx2mtMYfPTc/E9HMD6Jp5LvUYWLR/e7ARInRvwPMM/2FcCeUwDoEy8zI1LjRZT6icstZdDDMuhyi
ZFAAxq0MhA4DXrzJkaPEaPwwMmUHE88ZcJ8dqeNKH2dNAR4Zby6p5451KMTwOmO6CEmxxBBUO5w1
oL9fNfr6IwC0Of2A8PPdTmwqtx5aHxXgAoBJoBq6Ev/WrXEG2GW0P30vUpCmoYxid6eLFr44gjsF
OqpB2E3Dnluiq+aU5bucTuhvlm6W7o3/BL62URSp5qB6V15e8tMxZOkLeWwN6romoz62T5OQschl
gLI5gE+Tb0jwHPZyfSArXdRDmPQulGeZr+G9OwfC5JKKm4r7yyFbL8H5Bxh3VQ3NXJXjUzkKYkzd
iEUUZN6nwejjYb/5KnbXPOVwmWM/xpPzNHssu++mk7K+z2lStmB9VUyukLAwadW7Dmu9W9itGLLl
DUalS3tK4+Pdvvb6qkv/EJuDkqBIrXCHAxmD3hCqBObGX0DJhaXYjtGQv5Fp/4IHeu9T793t+W+v
C00R9NuV3Rw6qeiBY3rxzMmEiu8XsMWzpY18KaJbiyTEhYRnn5fxpZNGYiWazgYQ3ZNsq/JeT+iq
4Cc6ISEtB2WTkiBjmxDXiZBje9tGYTGE5Ub7be2nRDN2Hthiaf4pIZ6VI+Jo9aaeuokI7GLzqI6v
2JPo300Ec4n6OoBGBJTkwqsShHn1O5x8Nopi0U9mDUQs4x9aijFHJJlqcjRx53EAAhj3IbOMWtfD
BlmgM6vAlT80q4PxFQo8DUVL/HPEdcBEXOJSLDpRw2FtMSxJTUXUTzUdKo/Y070Qi3pvxCBdBRqd
r0aQXpFJXK0PBEqfbP+78sc84wYCr4bYLhuon7n2kMHUgeLPpEHapDWNwRKcE/H6kJ9N8Z0Eg+ov
zLM3IMFhEfdjwsbkdBHll5+VmSsCwGiJv8t43bMgzQ0PDHZmlgQd1aLepD8bl8qnGVGuR0JEIMMY
bLdo//GriQLzTza8L9OzujZp5CFPhs/FPbB3oriXvf5aMOu3XM9kEwoIy7+HD/UdU4qLBlRN5aRb
JzAHHn5svylZTcR237/3KbVD9a1YMqs/L60clR7rlGKlIfpDZflHmc+sEHy7O0rOi77skdaR8N7t
LUq0QdDJNdTAgzdgLk/Kj4JoX9p5qmlBEP3gIFEvwpnvl578ccoTE525ocOsVJqMU/pc8cLj2Uq+
/OHcmpGb+ClIZIAmKCYXSyDaDEbC3YnXwWAU1viSHWsRWkUzss3m2KSBcsc5V9cIJwTwTVIxPwWh
+H5bfUK0cGXAlLkExTT8bLE746IyNm3Vz19bTuWC2XkJWmrBcy74ZW5xsbo6KyawdWy0kGcHJrW7
knC89uA0mqesCn8enWDcwhkzOvV041dKbq9wZDET4ez3Bg2P6v8UfweV6K7YcZpikNRL7pFgQrRC
MZbMdalyLWKM4nAt4AMRwNM9WbPr/JMt7GxLSPfa7p/0arIxF2SwM47UTu8Xik4Qj6ObcS4CuR66
nv84xT2bT6mh9Z/JxUJ5a8LdEncr0OOk7mzq3EfCdMFY12A1ReXkvHDnCL97jDLXTT50jfaWLX+Z
HYELtWZ5/4DlCPFRNr3lfOz55G+AcmHVzl2HsyF5X9DkTa2cU6HzPyfiVjbqHKkvArExSivLE7hU
BwW+ETGE7qY4i5s3Ex2TyOUOwRpfwJpaJrc8ekzPngaJLEpfH5v/IkEBP7bngfCo4loeI6nNTFJ8
OjxpjhMtOolKc5jLnj4+CnfwuWi8vti+qVqRlvW0i5zB8pUAqQ8o9ot+XCoLiwmcL+h6VrObtrNq
ublyLAerCO54O7qwe2rHyR5oHI9fAzMqLMT8LPOXoE9rg2VttM6whukcci1WoXtuNF/qREC9jGgE
qldQ+C52hnsuXxFE+jizuMD9zLWslJBiTXn4hDuhD6n8HsmCtyrrFxw6j/zyOxfCOdDDwMq+/FQI
wThUdKweU/8BgwDCyDvsiuIvDfJzlM6QrpwPBv9a+9u5R+RIR5g6MDtUV1KD3fu4Qz9KRAaGnSc6
xrEeB/ZiKcJkwgo+s+Hq1TvwCM6FerBYNcJkF6rw2GkTdG6rUzd5KhXfaVsu029K7N402h/PLSZd
oPS1Vo4D9HVEXVW755wW9xlVokAR/chH2Qvql92FgWWzAFeS4yndgxhAwdDBEQ4aitQa4oD94Et8
ZIbvOUSBZOUwoFt6EtbT6ucrSraC4BR39/R58uOyYDeeY+NEeGiUwFANd3ZHsd6wSsWHf19tAGy6
AyWgGIRa9L9BVE+zPZ8f7fWYT2Ie/+TEP9u0MwTMsA0YN2ArrUNk1VRV0eaSBdYzWhQEzWPKxqwe
qfp6mbeP3ujfeHpbBZ/ZRkmQPni1tC7ZCi037lGBssWqaRDloXOJJ0gm580WXEp0qzjOkya9mmTI
AEoYw1H8hpv8kCY7BajxuWmwvsV24MVNmh5zYA0MignrqozXjGFazoJRIxppWBkUOv1JqO5e7W3C
neS6q0WarftuKrJYUUAAQ5ezKQlKN1yXTafKkYL5eerDRVInN6QdAI24ruw8WQuV/S8F2UcoDBUc
0fu6QfXRlVSWZH2euGPMJ/1+YdrnrXHp+rw/tv/Ng9L8WPt2oyZnJ7Bjf9mDqqG0LVPWyWvHcTUQ
YBtdBSHqTMd7Qp3hKKcp23p2eTnmTJjy9SnWylaeBzuQqzYrannd9sTlJvmN/u8Scl+yiDnaKM/0
gyWZcTeAq53ZqDSNIx32rqb8Vld8xGbaiEzSyacllQAJfK1B9V1BiQdPVI6FCTBCfAyz+enG0V6i
OwKW5qsUpc7qrswYFejb0pHHUEXT14F4gTqCEmVG5HtmrtLv7vEC3Pe9x9sG5UCtoBJjyf3Uu+NM
12B1cdygLMhP5nOY7Fi8/IPtuss/C3NmvscAUZZaUK32yNazLa4Mw8K+6TxJ42TLjXXEkpg8SfeZ
llT0bWs1MVfY6epxOIKx4C8qHvw3lqQR6hqbhCN1jHlHYbcg4/Z6cCl3Vz3GJ7ouHNhHCUc00z3L
OMJt3N58KpF6LLEkMV6OAMaLtHXzS4+24C8PtZAKkc+95yrbwChL4RKlq3l4YNvCBZVjHxF5G4M2
71YLiuwucwUJPX60vS0e7kveVQnCq2UZxrlKbj69KJbUmZjxl6OKhh7Nr0hp2v4Ss6A49AsrOawU
3zMFuP2Zq2BMZum992VyTNqnwCk40qXdlLZt8mh8iCaPt7yqPhiXo2K5K5PhbTHsO6fsnjYGGd1t
MxJgBMp7sisHPv8KrHgNJVMKjN58s3NlW/90U0cY+N5B0Y0shoZgk1epe6xHi0eWXxOX/vOPzUtd
RU8uiBYKDQ8dKcUzfHmk6v8XvCooRDkdo7OKCc/bsazpfdbsavS6lJsvQsh+TTot3KEH7xEh5Bhb
3cRaKE69BQ/Obiua5tEjeRYkCsovHzVbSJAdZ1bB5rt3bd5JPOyfwZfmu7c5BE/JgI0nDJM9DF9C
KnxbcIkKMofXHEKG/Sfq3l+ppiXoyAeAlinDHAYKWhHvUGicwTR0i7e+0pDy9V2RQY047mExiiZ1
Cu2t5/DY3QISAreX4wP7egVFpgROFBbGBKDq7pMdyJE9wgi5m2O9VhG7Q5LK8QawtuiciCCT2as1
ts8WLnGVlJNjwGlrM2M6QUFyAXpptJcPNKYFK41M7UKULLymO6qYtOnmooPGKktyHQIlSc2w5GZy
NokrUsvzgP77lx2gSJGlpuwYDnoVGvjnXbYUXQ23/XkytJksuY9uLJTh2VAAy1re/P3UNAAncLps
pF1m9sLIbzP18OLWLEQCPRtWQ090qMwegqOn7WZaP8h/6jSDHlGX7POS/eGdZkGpYDMGd04U0XVC
hb/+co6+julk1DsHNafvl0UMzNdCSZFcABkmvyDXIpUVfPIoCjGixUpFk4FtP/Bv6SqgTU6petYf
0qJ8isa0ZvdFWD4+nOELBbwknD+PvOPnv85bPixuMgnHoM0cCxDgOWOEvccZ2L88LP7kyIVzfJCl
KyLxtI+6qgstN3Zl/fI23ZzxbYNdM3N7UG3tzvF5B4QHz0h6V58ut+ZRpBZ2tN7Y9jaAAcNR86iv
2hfwQqpMVee0u12ZDUfHGiTpzQC+iYJkyB7sf7jsjFMI5wOqk7uzqPLbK8rv9CZV8efBwrcRKL4h
APL9esANhZvIjXVdgIkRM4xbim2itxBIaduJoq0TqBtaB7u81RpD+uqAGEZtBa/J2qkOjSN63Rmj
UoHV/oXcP8ah09n4gAgCXtkKD23s1TaszIfigoNMbynmDX1d3QjMLNacIDdKPj+Q/IK6pkW+zDsN
tFecDDGbMvXuGy598dLAhtHr4BSK2kUhc38RfPUFiODji+mM7/tK4ucFN+OydNnVNgQeSmu4SN8X
g+xGoo6wBIBuSLCs0d2i426IlCDppfNd8Qp2saNqhNWY+w1NTNIqYcIPKJpcFk6UOJV8uV7wgY1M
Eu/T0vhw4QUCoG+TwvTvARDn6QRZdp3ZP+M1InVYvyft8ordJ1zxvzmDSkxeLvBrqjXlyuw1Z8r/
9EhSmaYYyiPBEJB/esUcHTc8AuL6xbZSC8pkDYYlmoa0EXct7J9IHm9vtE3NEVrp9w206UUIa9Zn
6GAGD5Gw1GvUemnRLNkAeZQWH2FCqERMk4o6voZGskgsJoiWymgFMn50R6w0o176PW0sikobWQOx
T//2dNtxY6q/oOBZyMzkFpwdDznJGW4zc/gAUErEC2H3tAtlQekSKC8kaPJ4vctDlxqn6srhESum
E30bImC1hfOt0RJKW3lWvZyqgRb2aoJm8kZmAL9AwQkQmGaiG5KZPJhhYr5u82mMjW7AxaA9lXkY
goYrKlAg5TciZ8bJ+cMI/Qh/T4NE073bJ5vsPVvyrjb42nVFNeizzwJ43zHNgbiSiZ5llk0Vozgk
JWrOs+3JTxFc3KAcmGCSkdl6uXP1p7O5extjQj9HZcucq0ja41EUOorXj1oVNxW1U7o4zg9u+d43
d1cZ9t6evt0HxUBCZBtYlVjfb6f+gTQSWkc0hWYtkr61eFRBNYfLE5kcsLu1S0ioBG6+SOq6iU68
r6cbNQTih1/dYA4AEoMGbvewYjS3uVFLurf/YsWr0USXdZFEhxq2rHKeeXq5ONQnf5i0mY12rzet
KPoRKyg/lV/w9mE1qSAk2mY+2aNFz/QMoeMLIiyU24rpgaYNpJHW68+qcAZ5uKhzsKOrZCog8z3F
Y4Qha02O+SRUfclEzHQsiejRuMrFoLVEuYcF842Gz1Fa59pE5vKIa6iRUlp4aj1twrvvlTqb4AU7
a8I5OZJipMQe+Jwt2eWSYcWoWMnPB8VNseKC/eE8MChGCkno2X54IsSj6igWQE9wv8qQp2yzCw73
G7UT8kk2UWnh9rtuq+6mUNa7sLBee7VXFI8yt7/2KJztgDynu9Jaj4UnQ1srpf7xWbScjh0coyyU
GvdnsIAcOYDmipMidjvM0X+vMduVNe7NMpIoROix/5i3Uf/SiBsKO4mNFP35Bry8zuhWg4UkHzcr
s2N7e8aBWdDXk8n7SSaVZltxmp2dEZDtANxJeSWLQB9FSoKc+TcLd2VWTUT36eZcGKkD4joaexio
txfnitflIRETOVp452DJpHvyTbDFpeNYIQ52mcZIeF6mIdlT+86TOGpiYfjtBk8GdsTYSchch+SO
XhQUjGlYalzXSXihwCe8hqCyx/hqEK+BG57OTcpQShTFqmyRe5F8FCIORPaGpbcssfTFPbMAkKpN
297wg8BMF0CpZU8aAGITAM88AytAKUAZaw7xIIh4CuZTYEYVg6JmzHTU1Jw0hszrqlc78/ENn/Gu
reNKKC+GCrDZz6IzEEmGM1zFpZJN3X5kNCoefFWnEiX34tMWvlG11g+ZvTZyqr8cWCxslOxWPq79
8qVEcKbwydD1b3PBXp4vjKgZuY3FEfLlF0+Aub7nDOfJD3+CnSuX6kpC+2s3mZ9qCZgaQoWheQAe
9y6J3DfNdBaukUwNtOulSBfHF6x7ko5tmzLWap+EkHPFvToTnOmdVl4IxUEwoiklVx0zWSbvRLhL
BgtdzU45AbuBdnp+4L2s/mgZgjEwW0hZXXgr8ONWtzmg80dYzrC8Bcjssr5faFC+Sz0f3bVdknXU
lIBavEzxtCW3BCXhVPjKzia4GunSLLutwQ8I58nWQ2AHGzUG9aKHPpIXMnZRdXywnH35zVIEjNCz
Nc+SYlQzL5fn2Cm/f+PJeb5n6vW5N3fyKAdyCfNSw/85whZLAzEzQL4EHWTf94+R7T1rzF4mOvhp
GGsL/KsUK00C8RJLxnpI5j6/Lp4oF0aBrH+xTFifqLkkU4NHI9TBdJa9XAJqNwypeCu7mLhR504S
KCV3OGQNBNdCGxOm78Xq/lQFpJtPM7w3lS+/yu4CsnqzFDBsWzOjD9qKxP5eAIZuUqYqUp4sx74C
UzUui9tfQQlxqczlCPeN3E6fMrpH9vtOB0x1AOTGbS4E8rgnL0RFZWk2ljm1lrWU0GNPZYlLZHYL
pz+Gth2DjuW1ioF+ceZFCeQ8mIO1/bLtndDZFc2rRn09wZnuayxBjZVXhU5axj3eSTGP/XIKQPBl
FyvTeKZS44wAZpbKi9PqId1LXiUPFzC3UbZnyt0eBdeIlSEsngliJ5fEHoqkJelXfH+1Cmit3tGQ
mtt6bG/1SyObcmopbcJNDLOj3uL/d92RlL7uhF6uQxBZVIOhvbAJTjDaKd7FnTzx4Kq3LneXTHgT
QAhIZ0ETH9qguQh9gTCOPuc+fQet4ivLgJ1qXF+3ghShFFzRsNzdTXsx2Bi5fdxjaK52HSg18Y8u
oWJT8NAuIj1pkxl2/Aa/ynKH1p3bKazTzsCGydUry//9Bw2ADM/MIBZgPTahnAQXReWp7RkBEKkg
pkEhETmJ4kvuf/X9XQJPClBsAtx/zPVkPBDe0+SuMJdOvGXWGkuzW7bK5IQH7hexcUZZUvUmBqbk
EtO/ZD5UFbb7Pk2k21WXYNg9ZIEZaigqQTBCnwdgIy6YVZqvJgPkNWJjfUBg9jU+KKiNeytHi6hY
0+9MSF9GetY5DFoDq8DmGqvdB7vxjlZ3qBq761ln9VlVJ1G+xzCZNMjHhL3q5cOo2bxdmxFT3ZhZ
h9x3AAbcdk/U1Rq/rn2fpunQ337WsnwSA+8AwIlffwOF/45DwsEHILH0CPYSv0eW+cKkAWrxYtmp
3JP37TRqPr9NwKL+NW+MFj44kcMeBlytelzmYWknI2Kg4N9IqAsXvliSFA8l0oiApFwI2sS9RI0L
OaRi59F7KPag1wgI8rPy/AXMilutmCIUeFnrVhnGRY2dnCkPVUQNZ8dqPTL2McUHuNDPBy9P17Yd
5uL1vLVAKWT49ClTHbAsJEfzuiXMjyNjrWd0OReI9mCC0i4aRo7aJ5aHSeQkoJzCLWha1zm7D53L
rhtLKhiJOkaRukIxqQSlf68kjpIaKJK5t21O9RrReISb5aHQzR/UrcRsCQhYeXFaOXfINF4/GSLC
c5B5NPcfrdshWlkGk8dER2Q/HKZN8eLkJAeeK2mPRy1emGGZqcDGIPrXO4CicLLW76XtTNPPZsMK
Jz1rR4LZsic4Q5nsVzQBM3xZKEP2zHZEsmYiFIyJShQa4CfKFITeE5EplMn9SL0gIepQL5PB0RnL
3kjYh8x/eGvh1GFzdMhV7EDxxpiYVduUxlVrLNJPlG0CawaRd7lygXN16nT1UnwVlU06TMHgg7h/
3PLvZWWeTlGvTlXXhkcmDQ3CqYbj/Z/4hD2kBgj+89xLMtGbU0XO1U0U4S69A9yiyv6+V8mcfDCT
zU8XiRYu1kyOFuYd6qwbJKi/Df7JFJBP28oq4EvjU57wJ2EtDP65n1HN9i/ydKDG+4IbQUIH0S5c
Ke3oOS9OXvT5NQPQj3PtMHYYsYI/aMh+mi1FpLpgVogSjxUg1D22bM2bUdWLkdqc11gzsXae9oxH
HSkIOLHXfJmyPnGNUyxqhjvJ3N4wnbIqh9rImL4TFSDlo/darwsT76y1u6OMiX91asvDM1l5zf7H
06OTq0XhyTzOBOfWo/U0YDp30Ah/ySK9/comZRB8JpVoECEouwtDkPy6bTCc8FFscYmg6/d8RpD4
qKYhYng7gsbwXWJvatH2DrHfMxr/INRNLRlrTnjXi8gzZohzHKiK3bqYt8KLSHrsNRtoBnpi4gaH
loK+X+1YMiIYf1oHZApqGjsMQ8SajYkMcmWy9UJ4SvwrrlfJlqm+hcS6/R7ED4deKkH+3iSA+faP
eEphNEzjkzZmTKsRLn3m2fPR+EtIU2Wjua32hh8qygWetKHbQmoqWNYRLzDzafP7KLLX8pggHWln
LV7dRO7jwGlQ3W6tYge4i8tcNuMw4xC+4BE86qYtBVokM0EjkN7QL5ymsVctpW4zLPehxDYfI6E9
fCbwfb2SEYV7gHYD+x+j/bBkJnPmb/ERip9HJjdGsP925qG1vZ+bWH8DdpcDunyzGxnu5itUoxZZ
GdmQdtPofUGdqPv0CCwFU1Hts4/mxf6XR1BIxzuqHXoMIbnpZJmRWYPUYFZRUqm6ddHxKZ+h6eAu
+yUoBnfruaMWZ30d0KfVg66r18uqlLLfUEVW5Q9zFwspdJXcBIB85Wz1ZteHSSKidzZYNK5HRr6n
d6cImFv7eKGvXVc4i3zIVLxQizDadH+rGkBhV/fWT2UFoy4Bsjq4Bx0zYnpHSSPi5NUq9TCxusTq
5Z51wzzef8liBsvLf7Ai+jpwT9J7FBt31MVoqGqRzD45KXF0KagfLJRYYpcklVblovClnD+vPjq7
wu5CwC89tRTK31VNIgVStPz4Iu2Svrn4lX/NdIxA3wPlVTnQalMirwHWk7yizt1UmUMFlIu9fwgD
5ER8z+JbKEK85H8EqiesHAHEbxcESXucYwAWaJjx97W1KF+aQtqwAIpmgD2Ot2Xf5n7ttUk+sWQd
i+fDiZOg3a6RMk4rgOfdwFdBZ+578UfUryBKYWxBrUvfmtgB98JLtYRyabjJwS63P/E6ejqUV5Mf
PS2GN6z4vC94tfNgWrLJ7zVzfbJRd7LIO/ayGgMJTQjyE6NVMTWlrrb534arfM1dImG6jjC2Yt6N
wXY2kL4W/Sn3B79MT0ZZ0RxI8PBQaica5o9WlcOHhyXupRfIZR5O1wZfDGQard2XCaIcSxFblpTo
xqgGj/7gQOP1JVIDMaHFJ23EmSdHwsatEUIaaCQTASdK9SuYGByvSFC8VArqho0e3btruyWHkGf2
rD8nApY0+SPvBbNIUbacoZZedDHdMmmwEV2FQfdO+JajWx8iA1hlmEaxUk1r+iXlEUp6BQMH/m9U
VJMWLbWxfnY8oWYMGd7ogSdpYK+YIFjoaMxHuy7CAVHRjuI8zCrCuMjdu4FMRZ8FEnDyVXRkLtyF
GeQqT5suYcXUzSHU6ObYeaVEeOEzXbrluhIEofbojtcTOHpGxBLbqPyVyaCvd2an2rQ2nAH1TMNo
o/mvmHs++Ug/bkhic/f+aOYOtR6CIoUHYxjZjfGSWuDP7lJ+i4PIt7YUdN9rfZnXJaER09FB/3w4
a1jNBrr8WHgtp1K1Shxcbxs8tmxoFmKxkYSg4b0yGZSHnrGkMKN//qnzo11Aia6aBAV9udCug2XJ
wW3oDr0UdFsioAMwGEOCetWXAeEG3MtOTR6aS6U+TrHKt6NvzyVlpQe4st9PGs6brZ5xbNO+2DE+
8KozQQEU2mg78kBh2Kgun0y0pqN0apcmNJyySt+AZvOVN/EL7UJS5nDLLmj+D9ED3zvKLuaLvjNw
sW2kAi/Lsj2g3WyPig9jAGWtHhfkw6/iwnQJgs/89fKru2OyXsyBh5OfPhQEH96SwW+ws+kTVypb
/fDXDigjDtDwWTBB2cJp9N5MswxXVdqkgqpzBfdbaLv8Zf4KNjgtOodl7bSIUdl1vtw2puy9Xc39
+Q0tKRF2GHBnmauXqLvey9sowkZ46erskxVT8Z5W8EWLPU7hVwxqhWrFPNP5PE/zzptQtdyOhCKM
z5TO8l6dEX0mIDtnGYjuNPWbau9K0msbnOdsDEVZPhcYgGsTFZLwuMUcRNGrznC3HrZHfAPiuSNz
Mgtf/HNuXmx6PvFbkZ7YLnG884Ml66KcO+5XoU/CfWdUHOdUri3YX3ihr0YcFnGBLoUM04rLIjNo
soBmhGZDi15PRz3xH7CECLHU811Ii5KevltrsItbngVXfmzgp2k2arfDk+GlCZbymMYRjUmJ4vO/
l18uTmbrFH5s4IZkoOs7tLF5Ep++WDwTpDiMqX1S0lZww8va8FNuSvo5qk2g5AnplHZIzZ/bveRX
pRciSJ2RAP7N7D/Dof4b98V9zoHQzjBSNC3BsscgEBMeWXi4IBMNDpKEUy/jt87AOqC9jhEYZc+O
ChErZyNQDmAxlyQo0BCtDH7tfQDYm9ns7MM7Pj/zbDB5pNmaJ+7nCsLI+/Cb/smAfjTdFEq6Stnn
xgm5oj1q2LEkK7F7eC6w1DqWazCDPpTj/4GTAH1HCFq74+uDsJd682kN1X/ftOh4MgJRLAg+xitL
V8Y3nFCnHKDQ2mnMd/Feroe7UiZFBeuCJsWqob/LHtX9XAYZ8kS7FzHaylq2TshRvKJxkRA0mtlG
3wNM9eaEYUI0D9YatiJ8aHq6Mn/bBZRWBckwqOsulvQAao9u0S3Wenz5T++nDDT+h0Q16P74ZiMH
WdJlM8sHu4NB2rNNKmTn0zQcmABY5EnLNH3bUcqPL7+ULKmphnaaAdA2Ovf/LPLuKeWtNV57830b
6fNgutf00qEq4OppAhBe/GMXqB2ta+adX8KLZOtvaxaKIQ1wCH0HUWSjdeFjJ3Ml06KhPARqJH20
QGq81z+dbCiki14YzayV8W/uklI8Auptta6lmYCpkBvzHeK23oM/UYYSmsQBSEHpJW0t3YnkFHZE
4YvCXomSBWIdkVpXYwr1f8cjZDOoZCtI3+hTuO499qeXR2PnoGuBN8Ll8uGi4d3DhtDQTbkEo2/s
+8OCN5Gb9hah+1f4KsIS2GNtTmE0aBR0yycJ5coezAfSvFwA2zM4hwqab0Qtn/ZVnltlcLsaWxPj
P+SIAI/gbzo8VmFBXLS/vgxEHKRZW3lh6I9x4BFtXRQvrrjyer3RtbWuf+Bny0PRywQlj3+bGeVv
Kr6ssfNSZ4lXLxIRfoxZbBsNtb5LyzitJwbg5tXxiwxpcGC81UkiXjfpia3w0t9mOo2ipHu2JJeZ
ppC++H8vV4fLJAqPHbejMLmHIXitwgT0zdFVAgqaNdKnGEOeYv9337Hf1gVJVpbk7POt1mmWLOlq
UoLiy46bOHaq8+YCucOf+padEJ1FX8pfz7dh0HVl8z4KM+A23E3/LH+Z+T9lEsHsloP8iC0iYNEy
R40LHOIOA0Zz9MMMMRC2j5xHL9BDYx3SDfnh4EzsXiHU3gslKoSWROxjsWS8kOCTi9Yb2WlOuxlO
vneBEqOtl22jVO5NNas+JVXJw/6EztKvNuVU2ZLn4wUBX89yb49aOsFDaWpqjLYANtmc/0+gttxB
S1gsN1krQpbkw1Zcj38VgkzMSyTMW0wfF2Zfc6COUtLV5Fus0rKKwQzB3jYov3+l1SdAF30WCAZ6
GRjQi/sdfJrhlLQFD7A2xvfEo8yrkH6gAtSL8VlY+m9D9voC/4RkRYsAn0AvITeE0dM7pJ5Vx4pl
EmHznQ+/oLbAW/82CqrYNU38qjooikDhe9c7V+r2KOv0Al8Nlf/JgbD0q6vm0Rq0OXHrtD9T2PZW
R/N9+jgnjl00nmuurcksz4r8jRi1cDqz0gbrShiBfX3SRij/OVq9g8esvbnMMOvtFaeK0dX/fAvy
lhuswf7cmITZ0VHR+E8ahLKmjQEoSkYMjst9Uyzuy7HPDsy41wfI6+Puom1OEjRAaYvm3TJNK2Z7
Bca0i8Ssys0iNqgiXMEEMgpAU2VWCwW7iwSDB1AdtLJu77Twhqp/BfA5VuRecZJ1JeFEzV4OPZao
R+PNNa94Dupxzl9fB062N6tZ36ZQxPnktvtEqxc8NWhq/E5U1M/nsBXj0h5Xg1XC93OjwV0paBkC
j53LSiGMZ0Gkipu4YC/dw2glq0c9fS33RbaGDNgf07ofnwLyw388mOMjzn4TVs9+tro8/QZVjsb8
Vkq/aKjan/RADldi96jb4xjT97WSBPOa1X9K6YMsNeLHr2qEmkhOAs1qSxW2weOT/KKeNYMbIpUq
NgWOkyB5mFxH7q5/QW+zyjIzUBq+OkUZKHuEidUP5WpkQxv0dINU1yd6UiihnO5X0PygThcBrTDA
WttIdYLFwk+nP3AS4NkbhFtSMJR8XxPBGJTZbH3oHklWgVcNnO8OCQYLXlxJwPwc2TpuUeNT4p+2
d7iloA+r2JLG+G5Tx18wP9sbqk1XwjbBY2ERnIajU0y5R4lwLpPs3fnJPnaDZBAYzUWa9HzT9jWg
mt4pk90IoQD98cP9SaI3gLQjB1YbU+Lh1XG2recE5aQ3P2m7hPPrwYDVFXuL6EkZhUOWPDwQ5gLj
ZMC4sljY2qSmu+lDte3U8cAqRj4NmB9wD7ho2uNIHD9JzPw1y43sk+IXLxs0QKuiGmBolAmM6UXw
igB/uX0yl1n8SKz90Iqlk1SdQ3JLN1lK28gsqSAqgWu532GFVmn4+snT1jhei/6Dmje9TVYP9Pdo
H643rJ7TI432tORh5mHo+hOUlH6Iq4vILJ8+GRm/ISLzDLcvrW6rQ66CzLB1ClfD7Tqk/ZwLwqZJ
8xTjXdYSiOKp0FXWbSdg58DGYcxbu3kBAlc62jy66ADuklkuEq7vpsMSjZxZo9+m+r6AnzT4hGxw
E9gZQ4aBrb1cGpj2yd9GXPr15cHkZ+NpgrFo3tQwMMnjbmCKosRm8mkiSw2AqcglW2Eiow0EklmT
Su09j+Knw6fwRnbdTF4O0cAMVe2wQQMnHLKGBs/y4p70xxTpYKCPB/AIr8xPS/GheA1dex2WCkh5
m2M723aG5s+LXoga3USi1ijHXKISV/tPvQsFn6FN1WUUbN7AApbXnLq4JbukPy0ZScRbMT9uE+5r
ZQlXD+2Ww/dvIviaji9Rl0K37fYeSfjsIt5/PA+Hh2PYXSwuvBO7u91We8T2ar4Ep/oFuJ7Yj1rT
zWjMCfh99Z1ENFYnVaxjr3HdkGZ96L757Wq43nM63mik1WlpMngpnSbGd2m2MIUwGmHzGC8p5A0p
sx/PHLceZo7O5daD9M4hc3NP2AUaP3HAN3u/E0xqQqfZuMoISjNwd562WSm2iR6XD18aZLBI0GSe
qyWEHAhFLHGHo+gQo4B2O5JZKzlLtoDIP8lkPpXXHOOoXqXx+kkogYKjKkYrw086RiZgySwVnYNp
P7bKK+rE/4I9pKOXM2B9pXzyXMrOWMH6dVRWl8Bn8BZBSRcyWb4MRyB/pAL175RDBN+1lp3znzb4
/mwk1yDz97Ija+r3FMsHNn1RlRxAQSd7XPxw1Ai3dSpmiPyjrCX5mTSfzMKJTwFCzzRRDCa5GDyq
VALAt81MTu1M3PghxzHVPtieeTDisxtHcFGVrplCi8/IIm7VQx8/TUBK3eAygxAhDacl+e/nLAMh
S/M9/rW1PDg/IhReKTASe7NamSgqI/debGKAjOg9xdscc4zQB7+ls/UN5UyulVUZdHcV3Ye+oNF4
jXBRn4EEDxqy3i0wrd/8Y3+Gq+ZywmjlHxS221JgJg+YIvXqovJC25bo1b3qr/96tiagRgV9Hm+O
JuSZavd+vtioKT1NwY4pJs93fQmyMADJCLnLdE2cOyVHFXFJZkNfUiSDLzWaGOg5c3Bf6KFoUJgP
t7oBpoI0gvnxVXszXJpe8d9Voi6Ag1gf8eEMuIbAthwv93GTe45WSpZcX1kks6u9+td5UW8YTvcL
qKCICsI1W+PgdVZjISRdvQy5vXF4GUDgJO2f0NxQDFea3GtpTb1M+VsTW2Ts6Yh6eTtajeg6Zy3E
ikYyaVsNFPC2Z4NNKuxANohcTQdz8w9VVQDl+0TXwWl4RQ1x8L5jrJqimaESTV2a8XJb+mBiYvjJ
Zcr8X3fhNM1XOIzRtjiC0dJ0VmZsV8GwXNdGo1YibEB6/vVL44k5xPjF5RAjzvwKga5BqdGvvVSO
SxfmAnHQUtFSMf/6dCyc91vkAqFcNEeJScR7aygixNYigmuZTz7pGJj5iU0kKIPyF5DpufkzPJh4
djC5M8l/HhS1EFHxjO5iTBURmLE9YMROwyGcfpGPsC9sWhZz8t302hUVpYuHeLgi9Yhe3a5yOh5s
2mKpAXOimtAImXsjaaGlT8Bv+CVRBEETmKCizMW7gx4eHgwXZ2VxcSDQTaPkE4p8CD64xPfabTpa
4V1hYEPK0H8A2ZjEpLZEPq2uweZ85Um/ecn+9rrC10Lt3LuXa0slJDUmDtELmnrGWnimw+Y0icFO
WoSoGr6xmYZ0p7PTd/5NMkWa9Qb/ZOf9plJqUlu2348DQwJHqTQXEtYKLzxtBeYHnZZK7WNFt1Iu
ACcsGBv1sF9lEJl0j9TBbDkABEvWflJmMYA8sWLryqJmnx7Dp8+phGZFYHaCOJCzHd3Cb/8rpiuz
2fzVdMicxt+TN+1lfh4zDtlxc2jC4vgZj7U660UhnpMtDW930PeM/4rgBnmmDzcgBN7CbgPQ9BIx
Ob1pgacYIrGCcbmKMEdVlBd/6EmuL3VPrtQ7WAeGDseZHoEhU9gm645Ll4lKblAGYKfOTesNuuQd
PfxeQd3E9/49A9K+PhrqL5mi0FkgfYD1kmOqPEC7KULgTlMX1oY3YMFtXJlkJyZbXt5lEqY1foc6
ZUm+KHXIJsKWqdFFy6AbM4kKXiYAV8TLXrjFehIBgkyytwLgAckdqHXAuJtkyrjF1hAQQKryWiOZ
/MCZqm49KnpFbZZmgW4zONXw9iDtvPqM7x0si2ctE3QOnp3wNaz/pdaHTbPp7rxslgewjwOrnFHH
fiUSjK+PVLwPz5kQhQvc7PMLgrE7jIEz22WUZSS8pGcnpgBKK8m9HL5yyZIp4q/qzB7J7xZUR94d
koV2hozWGvH+YvkMKZG1K5Cjuqk5hTw/NBGzdswQyW/Ok6cZGVUJr70od6GgWy57yyIio3c31I0P
BWFEs96fwS/2jEuYbpj1W7XSYTKP/0+qO3u5SnEq5F4dp5M0LvcMMmJ8a3KJ/aMoQdKfx5mqtX3p
b79m2GdAx3/c78Mak7+xygLioMsQG3XCwKX4G2CkztcStR75CPCuJdDGnjmMvBDP9Kvb1W6E35wX
+WDuEGp5IaSttKrFgxjq6JLGzBAVaFupGKKUPrAaiHCwQxhDr3j+qdkxDF5Bxc+ezZnoIthf9o96
sm+11IohOcS4gCTO3yulBzRR5b3Xxym0JXMrmXIf+uqirWarfoS+UF8WKjrr2MIt6/2d0Z+1P3PQ
llV7woRFuTlhrc3IDfIxsvx69Ajpr1d/Nh+lBQKDxA0FUI1JPOCF19hEb8IU/6bXdOQGZFzrGUvD
XWxw9Gkncw/kGEGOIE9KipjN0msqXBbE6BP9A5civcRd7aFczJaPivaHPCEa4iBJ9xVd4v9big2Z
gWnuETXOkz1QF6rpfUYMgTyjo9+ekju54+VaE+WkuJDV15cXf4XreUdjB7MTNc5G3OXlu4kA/AnM
tNnD8/TBO89yx0m+IJY/ITbY1TifIaAkg05/d4GitjpmkJ47v777pRAjUKHnsJunfg4+6kXd/CCS
2T0leMA2BWjFykCQy27SVuPYDemIFRJYLmXjNXYGk0frSj716Dcj8uITPqOAfj+1HFlgqdzR3xfb
AetXtakPhRIlM2jnxsSfUTNh9YwMLHTtpXhjRW38rXBdXsX7Io1rZX9Jeusozr0cSVApGGvgos6R
g0JaTF9VMyDsyj5P0ah0TW8G2Q2q8Mjm+xSrCo1Jm/HwhYXCE56zbSwXJrhaDyk48Cy/rzQgoxid
AkYWoAdEyxKgV1Farbpf6W5xsVG1cXAiSMI1rybgO60sD8XZE3/ruzvSW9fyXuQzugIGxjzyJR2k
1HK9U1WMvC2QoV24PMN0CGSFzqS/rmtAZ51HbA3f7bJfF/k5pxyBBtoyPy66rhAhJFwp2hgPh1dO
9mNct8TO/81DQYhajitFgR8DvcFdOb1cmaDU+36SZlbz84lHHdkgXyd0ETRYO/5SbQpgh/O4FNak
aOO2GaiHJjxaXwiYzKsHFLmEy2gZJ0Cknmr7uJTtEMCpMn9wlMEQKKZKxG5nIjMl6O47esYXvsNR
Oil/eBsGt8/wuNkwM5HMDH7OpS1oEuEbzMurxIUIxTJJQQmE8xKTsFEgjEEET/Ot+6ayWcM3Z7/w
HJRwdJLDFTuSbg5gtcCCOtMMXCC9hZgnK3ztgzm9pjjKsb9uJADmTiVgFLSryC+IbE9DqA6x5wCp
usuDEfaluVLzUh6RgAdhWJkRQBebCdAzLOrCVA6uWNhgsmiY0yWRfkjn1HecJ42hwTd2V48vBoIK
JIPBefDhAhVf1Kqs3WliNYu2O2AYLdYmtJgBnWciSPWeBKcRVRxsT3jpPOCF+xpLcAVWvWbN2Dab
JsZaYbDulsKoyrBW01tbqhGgqkhl+BQNAKYG5T1ubcZYztmIdGRx19gXADOaI1cRntJ5ZrktK/Gt
2qRjn94ZVWI6APqec/aOgJbUIlyEwfWx87sQRgkfIePm8G6uuvsV7nhl2JBglfU9BY4olNCQgSzL
LCuMOWm9Gx+UnERddCPdO8p+DHNrRexWPezO9o4dzSKMWMp+6PmAXmYTOHYx7HinffGUgP7woFTe
pM/TcfbEGqjUUJJLIMf6eAR6RcjHY9RHvRvmbjJuKqjGsFMyF3RnEw1m8XGv4oaec3tpRlFnNpDp
nlKz26U5CbRXj9IL05Tf9hfojIaV8hIDD6lZ9svGgM7Ygpx0HgVC17rcrpEPTrP55m8q2X1bNnmo
JXmXWfPA/hG8CwBcthqh7yEVGAWBYVWKkUWyZUNHY3j7EXxcy6meXnYc++q67RfB8YNQ8OyJVkOk
+H6WfkOk4xVqNDjLOYCJ0aY+u/jiDi4dQUJDHgpDlvx81ybpCN5MwKF6Nc214lLydsccWnHlZtlb
jjImYqv6WbOQAJT3mHCUNsx5KuOoHqAXCN/2m+rCJA+1ygxMiWuAj3oLs2GYatcOhrWTMLV6gevC
esxkfh0Nmoc9k0ypoyBWN9IAnR94VyjlYvprl/D5T/iyF9MtOmqKGLH2ma2f81I072MKMuHegbwn
chIK7RFvvBfnmbEzkh9nATbr1+iYnh3eQiWqsi/Z6nhVxlQkQNoPxYudH4aN7dVw/4x1/c3hg0ad
mqKzeYbZTVWjJuk71F9n/Ssmg38dHt7wBN6eWuNSpwiaGZut+1UzJiEaMDJhkU0SoPKwTZHmMaBP
6wlDmv0IidTld2gFZG6YrUXORN6pGTGCPQ3MRWtA7Rb9zU4JctsCu+ItHlKaGKI79jneqCSJpCGI
uMseqhAa9aCDZCI2WBi2V1O4Dx0C/QVgG4uCSjd4RJzKBBr8Hxz/pw/Q/wadyY7nTonVcsTaVAzz
IZ4+uCGMc2fsgkRYoGvSApwfyQyGYoNVWn32jZ3SH8txmrHqjlm9alL5gVHtW1WdCgAdoAK9sxP1
Vx3UjLFk1QSZsOpSThzCjATK2zsHVOXkzrYI0WuG25kb38JSK42jOTYTJcKhFe+lQelGAYHi3kHf
XbDNEiX73vsgGNwJqsCsiRv1Wmh6cWV/pYD166eNluojv3F3Ohd4hXPVAMte6cdeeiGBU5+swkvf
DLCENEeQMZkGFaLZ+WcvLLPQsmVaVFcol45t4srtnltqib+AAnqgXWnzjgViPguFUN/UzDdtX11X
IPlPpuOAXl98meyBmWC/h/BLRetMBTNWV6/ZCxTL4usFMs6JayPS7/OXxdL3ixW81WswnQeu96CR
Bj4ihwVSUFTm7Hv7l1mRf2CMdVcvs2UqZjeid7tybDYS+X2NqpVxP0MFATQ0dcb2HGRfrOVrmw+H
L1APjgw6yPEOyxEaMF3OPJ/XjoTTw3ef7ZVP3K0cUqvnfscvWvnClcvoDVvBJfbj/R+3KTC+/oIB
G6xO4xOIQYwvbZCFEbTTJTjDcgLIXRbZ3w2w/rK6+sD9kjVe8tmjqpcUiLuA4a/tJ7ZcG95Sypns
P38WLH+Cdm6Fhw8gGhrOaNTE5Bbq4cLaYmqAoO6CVVZoWKKvDBux0OOyMKd3v/oeROXgMOBBxgoF
w0SU72GPmOf9hX9zVVB0liTb1EkEfd9YxujzMtyIIN7914k96LaTQkPaOI1N4/UvrhJ8hPNHeGuI
xzlQl5YuWZ3lIgkNL+TbEBZtJ89xNzvRJ1fgORnIo5kKYCw7ZA6miRr/aNB+bfrSoVmK/HO4NJmU
NQE1AHnmO1wRDJ5iKUbT9L3lhQznVftR/P93rV9XYSVleP8eve1hpnMboA0N5aSMH+d4+WwF4vAJ
5JRHv0JAPN9rH4tEN3ymFsDwQRvV16XLH49jxjAETreZ46Meoi3l44lU5r9ga003DOvbjTwnZpFq
jFgYAfWxzYoWf22Cd3mpfD20e2qWUGoJuhaisXiGZml4IwUzqd6w+IzaphoSZnU6r5jUSCblIRof
8a86izmXG2d4b53UE+eR1SofcIs/24L25Ep4epQ9tAmsQuc3FEV+HWvBDdPTT0tHLPAGbLCBdRGH
Fjft/eSBNALUSFTYECWStcMRyFLB6mGLUufWlXHvu/HJFNzlQwPasRsX0xRbCkrjbPT4iiumV8wF
5OxD9K/SOYJHgU31zbMzo0y80qVjGNwDS+wDIZnuF2qzmYJTRckfGAF8D5fPAiFmMK+8gFWcCFW8
/hwez0iWgZUkKz5RfB9omOYrTNEgPEZW0ZQVTbzrEvUnbly4TvN8r5rDYiK62sfh6EWF6WW7A2CB
yIbR35GcsYOXnBmTttCq/GXT6wQpn4YR+rqJlWxgc4tTYtDpV5aGwp0GVoPccaVMJxu4cNnUOaVn
Jn6VVev4dOqR1Kfcek/uzjm698kVjNQIisXbk2aTUyVyHiZyFxd2DR+9RjqXEKtolvi4YOqEDvIE
fnq5ve8+6U3WdXT9ThccE5wkBDgOLN/P4mafxf/SfailoJIgKXFCHa9yNCCCWM8qvs5GaR5D9cca
yFoIc0YDQT1Sc+9GWZ9BgHSXOF3eNvH63yKeZ0j4Cjv/4fJy2Og+1U2o9CpywpbhN+YOpmk6AfMg
+6KtGCv079zcAjDQ1RbrBC1xnkpjMbCUyioZg2GR3Jtaf/+ippG+uaCj8h3tRwZG8Tw++Iusj8mV
sW6a8i+n6ZiCTnRm4+g2hdpqEv02J5m/1W3wKrM0eNfj5EmeKoJ9k/pibJmzBkEjPY89VMs2ZfkI
oZKrDOaVuHwoHErzKwwtbgEW1fR9kAxVw8NNO6ViezwINvB7it9d00pI4weRtn0EQMhgg8EAcGs1
K1CAv00LcXuye2KdmWnOim1QHtR+bhwMB3AvqkyK9i3QnLI5xNWeheFxbsKibwGyLDQZ0b4yJQpA
ujeh8FW5HDhTmnSlvQMmy+ldATbTB4V8BiswqfUgYc56LPRMoDKZSVXdkVpGYLfPlqix0gCRpEtH
AAEJuG+LgMuEnyrOeVjfSv9NIqMTpWp2pngpc34/k9eEkYn9D4+1xXCYxuiWkJ355DW5FYZ4MDCP
Evix5tnvs+/d90Rej/bBeW9wGdHOArXlMJy/jk2r8aARzEgeJzCNAutkDHQ8Vl39g42od+FkongJ
nMsb2pgCeadIEvQA6HIyIs8Z1b3dpscnQ0mFXorsmGDvQonNrezj5Z5Vt2qVOhbS+UGldmTphQSQ
JOpnLaal6iqeB/rtZFx4AXKJUW6D3mLwmFH4f1/AE5BsvF7qoDGReHyhr78I29bflcBrSAvoZBId
6zyIsufIa3gyCZ/GoiXxpMnW+BnRfrP/A8NIMKMkGn2/3q6ERtlRexnsSCRFzubbxIp0ZcXbiCjm
6LEHPO+fiZejnERq5R8kkClm2ygjrTYfmfUq67CbproS4VHCSUk+uOTBPXYcLqZd5drxJJuizNow
qRi7+rEytwAztHp9/4I5OkPzuKN/UaK22LgCul+l3jSA+I4Z6zzgZ1lS8sPy3MG9PBujIpzINHqA
TBjf9xPnFes5zHfUfzdCBH37e4EWbFPQhPZExML8zAWqAdcVq6KBQ5bDw69Ha90ed+9iCIKuhmUM
kIMlqPMTOuQRpZ5xOZ7P2Itrs5bNfhnwWX2f6lkaGAEB94gkvOnLSIHQnFj6zKfAJGf/LMhotz+l
dqGrCpaWuEYMKX7+Sw4K3zpaf1R7UxUx0ZwhmVu6bIBJC2TjYY9ztNssOkMXkryjLcj0wcmsCYrx
vTeMN9vIFwKwFKl21YlqffcIF6H4e8HCpjlGx6EF2bcV0pzfx/Ap2TUBniYApIBPe7ZXtH2eswR5
BaqA0BQrt1ARSrrJ1Th5Zkp5hUvvx/a0KgI56q0fIFeXgyQ6R5w7H9Xe+LRySqtIQB9DZ9QnTTgH
Lpe3EyolUPWIgFbYCT5GtiIyz6ktGD7m7Nx5HPhu9TuZ0J8F0tBRCNNU/zL4K3srm1yYjOsaCdN4
N25dc/l3KHvSADnuJ21KyATTAV4gZ32FTDOU8bjTFherwe9RNPB9UIctW2qT/91MkYE086ue4diu
27M/UU9XtCBJfAn3eWWATGAdAttjt8sYCql0TyMRrR1f1IBVoC60SInE89fb9B5QKBmmbc2tbnlQ
QVC1fhUVjDfkd6xOU2v3ABeAksLfQWKv7ljCsX3cyW3lB/C4crGgdznkRdP16mvL8DdCuViUEK8F
HP7JYDnbv8YE8zjrE/ZhifVQc8b0Nml35bWsNx0DOiAF4nO5WIWa80+yaVeQz9tGBYLhARLc4gf1
WRaIANvELI8C0zmBilMfSoTNsDs66TX1qHjjbdM/MQ1lkYjiRhHAeoT4+P5ipwpBe+Ie30zOQqjM
gtaHlf06DwBdJom+CE0s1fUjhkX2CmeOf/b5v12vKkcw1Azs24q3LEiuvqdgPtJLh9PyL2PNgnwM
VNt2wc0sNXN1S4Wn6mfrlD7wCx/XbOXVWc0GRSCNAVQ3E4xGK8ub/LqCNSQoC1TH//WkxoE9VYBN
4AjlHidwNSaDSH9kpKyP+Y3Xr0DRzS7wfhU8Ns3XdTMmy6I8V/7A48K0/yCSnLJbAKtH64Uw1aaj
5Kj1I+RB57Rzjz8HlUS1cSNcyNP2xMyzU4aa1Aav1z5mrX8cOD/rQwIAcXLWITMz8MQyfdTipMx5
xbq38QnM/i4RbSmVGiSyHftOuCkZmj8ETgrkpdjmD93/k8do08r0kMoAugLkiaiaaJX1ZHRfZKP5
xIbhE0jYuh6kgbW9wuTj0frOXipfDjc1c4K4QxXB+MitPQTkSQCk4gcLmGmBT5+2xMzYPyiNAzIL
8lK7US2Qm0pvuwYYi2DRkwdANMuIqK+JJ0YgZ4oEvD/WeUlUDOiw1HpOhp+la5QorDYVU/Ryt+5h
aoSQk/S5vzzrqadBUEVEdJaOZXddc/a4IqxkQs7qFAsvWp/zqYHMOtgDqgKUjFts6pYyhGGy6qBx
sv/OBZcFWZqDGsnucnZMziKB6/pmaResyIssR81YN/FubGy7ICJ8ZgWfA9qo2DO3W8vyS0Qo0Gyi
gYSgw4IuRAnM1BYcUVNSqQGz3MUWbVW53N4eQpkY80luxr3xcR3v9I+zPKWQ4rKGyGzyRIlagdEf
hLUf5g4WqoTy1Oi3irowtay00zieOB83yFn8n+VgHO1mtKb3g1GFpHCOwl5XX/Ft0akkYTIGxPtV
WKAShEm1uizWWZcOIAXnVdb34K/QYvk1Hy4k+7Oecf9w0iFBhrqYx2HY7g2mn8VeuhYoSsqTd6SF
KnF8zMZP+9LGaB9iG+XvK0UJAUq1c0WYq/09I4G6UQ97UvLI1bfjG1fbEB/OjH3cYDwuxlhwPwj+
wvHTgKtpOk/tmNxl4CpWMhjf2eLLAlBEpQfdXQUMefO9hmxPyU0jRvWOhf95/JSJb590dNR/U/vl
Gz5dReM5GNFnzPDkR43tT5aSdPgpH+hhjecCTurDUPVzzUYWlH1UG6hQvsi93EA3L/JKG3pfrkju
5dgBBGwu/tJc3a11Fdu/TLzpDIeYf6InOacWZm9C+TgXT6sK6BhUascHGOsbUqzf/QqIWkuSF/R/
3qPQxMsAi5WhWCyPV22ZZqnDIjpqc5PHEsAv9hAbc6EcyU19fwLWDjv0Q3pw1p3HsZo9EC6yeXe9
IH1RqoFdselLj6icthjIbguPdeiZracXbxFhTAuECTjqSjkirebC/pxEP4RIcpYWJbBuVQVnYEBI
FajCu4P2NdmrHkUT2V+tYJMLgkDlcBjFY+JDrbrbwYXUbO7vHh1GUEjO1FfWNX/lbypdZpvu2bpC
mO+3wPkHZoHZUZVQQXI1BpeY61hHEUCY6d188v4nMhX6mH5nfu1SSj1yUoCjHyvkUCri6jkbx/zZ
onvZW7NIuSA3M/0yUL9U3j828dbdIVGMdg9GmP5bxvtJqnEFBMqvSL6g24lEOzZRtZe2A2pw4yZs
Zx3K9gOTNQEbID4cRuq7co7lk7ZdpFjH8fxK8DAVJbrP7D235SQ/aZNYaZ7B1yJGzgVjdkzNGRyz
225MZ0fnANrAtbQ1jC4APjaliaiyWnaebmL8P0fdoQKrof3Gxf30DNYaG9uOpWBf9DRBBoNSBO0k
hDFvBpYt41I52b+WoSIs9SF5KkU+wWLM+CvEfIuM+F5R+mLSZSj5LCq04ctbGalok416z4v2a43X
M1JH96YD3icWdtuPE4vRmcH4gF6Zt5qPjPh1HbfruM1oP1YKj09hVE9QcJyrxuHV6wVttRB/2Lra
VgErfvhBJ8jRKNPsWfOGdmz4vG5uVW8H8DXupKVznwmCVXgqyl69jOc32KUm146fqM/In7Gn3WCL
Gq0lOIGaRpL8Op9iZ8kblN/M+SPAFsUe8AGreCqwpjiEPouz8YhajZcihoA6Znwi46d1bkGVfCkC
LGCABXHgWY6Mr+AvxBh+kHfF3xU2L1LkIRwZYLLeAdpO6M75ApSONc17aHaHu5LR7UdDZQ/mbAGr
Pj5n0cAcs/u9oGKmYusQMHfzNUNhajhtYJNu1jYDa1OHaP9BYw+6wjDETQnh7icdtEuCHs55SyEM
pd0oX4Ejbf5wUyUi7A3W68PR5ujXXnJ9d1cgKomdJSDA8Y6isXfEkVXSWhW6wOu68MP5uD3ri9MD
CD36XRAP0zFj1v4bt1bjxQDtBVPT+c7WJ//xyprViZrkwjUvWyhB0j4tjiwn7SyFw3tki4Kcntw6
lS2uPRPZvH8+9TahefoY+EB5uH66sxJquf7henzS7rx43YPTkrfqMdy5ARrzlYEJYEbM8sn0+wED
lYExHr7rgIwIcsGHEWSXSpsTbqpuAn+amLI6XHfQWwKVGRcDJ3bDzTqjyhcJfjn1EHv1J5s8yL/g
CnGHelT2Qs9+Dv46A/CY3qizgX70M8CvZu+Jg6nwu138P2GmhEMcF9FQkhk1vVSJ+n5n+FXAjlAZ
iopqYLI4BrZS1l/2ljmCouaW8nFIEIaCAD5/YPvmXYPKukK6iAaSOJH0G7ToZnarOJ6ChC7Ykw/P
FYHNO2QiHQCwwvzuyJgX4DmZfaA75hxwtnvDxikBZrZ+Ynr0foNtk318lkylT+FlZX+bzMaHMwFV
bHXC7UCKq9EBNdEpP75qrShGXivs+XEN95etrlhYrp8am1v2gZglF5wsn0jirgTCCmoyrVDvxQHd
UFszWh/Lv5yaWgmhj99fuaL+eQUDFoCsvUWzBxLL6EnjQ00enRkwUE3ESlmUBx9an/1ZzQylxq21
ld+3bDlgUDORr+N80Yw6gWC1ZdeR+fJ9yqIfaKaNB6b617TW5JCoXeLLqTRWQ31InoveXOJ8anp4
jMGNcd+QBcPe6VqnVRWq57Q5tXQtJmnR3zHLUsPPnNme9UNwl2KG41auvNzniejbLPpVe+jNbqDe
UUdziCv0IuRtDMz61FP8vWTZw6Zm+hyFaNnqIugShFOJ4IW48gryYZCvfZOr9qtWLsR2+oy4XwOt
vinMLWOnmjNa+S/jmGl03kIXRtQ/vxrCkTCERJ+LjyYsLEh6DpWHTXzcfxDXuYesu0fPG5qRy2Pk
XPa6zuW3a7qo+Z53cp4fimGvifUL9xSTn1tYA/9vIlQV7INuHDRgAEioK+melMnVq34bBAYT0hsX
cK5uNB1iE9xdsSplgKW9DDp+WScNuevD14KsVh43NxF4jo99sS5n7Rj+pLnDW+PuHtdgB+GtzOba
11sqJ9xTu1QLMHs9WtYG19gZWlSvTD2ChOxU3NKZOtD9st5BsSLG3enojTEiW2MJr0uuMiz11lfP
ssnG0/btWttMN6KzsWlEmaj/xq8prGP5+iZfDBPf+AEG31uNi/kfv6y+UDl3b17oUxZO0pc7C1+f
b6CiNe9Q7Q+sCnuA1yb6z2bwIpaPSu02hT++J4uePts1NRExfzgl7WDuIFbO2PBvuIzD9A8LiyST
mVc8bB4qplu/bCZVuTQxK1D6Cz4/9b2oiCP+3F7LZDOaCQGLXC0xNZL7gw6i7h/xpdm7uRSZzXtc
NSUWALC0Kowv06RcMNnyn8k/WYwJoQj4wuq1jIU90CLCbQLJbGrHaIkMw71Cv7PcJsZeFT2e0rSj
IWv8sRi4i9Kg5Ygi6WHFeW4eqVuFojulRdX55zMhJ3ahh8hFOZJY3NT4ccAzvCP/cAYGS23WQ5Da
1h2+VCbtlFiuHAEfd4YYq8UQSYhbLPH4hACHlgkRhm0ZVJGmxOq75alygbdFG2tpRfhLmPX3S59t
hxEZFH9s1PJ6crUH4zhOd+QG9dlcY/RKQmaF8Hi7YDRzmhQWSecNYKTy7cdc/Kn9rXtEEbrlcY0d
6NEvMbK/CmNduqWYAOfEJ2AoS6ckOZ2UDuc274DcbBddKWGSHZInvIaWnHR5mZeoUSJqf7486YFB
YsgcXP1bJmuiF4wYGhegtCzGpWANCc9xjyTyS1wADuDFRuDDUHxB4yJWr6JIhUr8ZkDQ+9H3w/k1
sbfZziHKIXb0Q+ehyS5eFN2nb/IfVS1iQazdKKoraIVKhciWv+mtHjWsa9Er87S8QSxGyJPA6xg3
otVhXwHDl0OppqHJMVLUq2AoOKEbicDLiGR8o233B1udAxxOTyCDV8cJFvC0aDQz34JFBwzO6O9p
s03SDti7WqZ6znfToBPZrEk3S+11xiupE6MdCoIoJtvg2ff6G5qFJvX+fNeDRw3D7q9vbrIdFKlG
MIP1Zjk9z2cbZm3sG5/TeBxY741CvyaAY1PAUOtqmAm/0oyaNOUqjtAknBWieP5MPAZFv1COoKFg
frTYAG9J9UcQmQfS0RNrPzfMw72hL2YneJCCOP7nvoMvqY3rnhMrpY1l5HJ+y24mOXQyRel2ctLd
KHkYhwQ2kzx+WzMhhPps/O84Kej+Ph9zuAAp4UUdouSbRJ2t7mai2ySmcPc0D0EuzGl5mekskwSk
f2OyLRiRSBRzf97OkNL56oun6NkUid6xhFwGloOZw0fwq76sUz/YpBRK1IwAtQJ1495SBDma3M0T
ifDP8+NwrH/+vjnVSPtHPGWFWNWZiroTImVT/8SteOlEXKPEnlJBD7x1/CjWuOIyrXzI+G8cpvgo
yVffL4bO1UXgY+N8HlDsdnzUNoVFosNsAodMSSy5S82gccKPW2ZDCJQf/W/75prL/WzlY/FWf8/f
tMnIHJEGX5pWYeqTdt+XdVSdURyOqIwhsYn4auzUmVBtx2Jfo6iHVibfB9KRYJ/kGy2S9/Ck8mxs
sKcKPWXgQ+k0246DfsTprT7eipucUPEtUwkSQU9cigDUJ+6C5vXY6QdZA0Izp7VCu6VSKz3YE5J3
FRcA4xgJpMAxFGbpttVQdoHRKYqUBol91GTQCQmDt5GxcKwEi5FqS+Vekxdmb9kAbQURBGLSY0/h
R1Pii/yBo0sRGD8Aa/GeZjaZ4uICxQeT9I5oqKrT53YByHfPP8Yzm48+CXR1xyRGpxIsWH+N/Lxi
1f5z+X/qFryQxibjMBgttePfuklIGpjEXRszQASm33O8Ro49+aORlUtkhUAo5K9yIF0kF2jZqNt+
NVbysjPS/nonehScnkf28YA9ZL0BH4uoyyMES2sYJQpwffsdwv+DqZlUaBEhppgMSCm9cUJpz/gH
+PvLNx4lqfx/ThbKf+MPop+SZdRb8iMwUDCLvqBNroJoIS91UAIDbtqcBoAbcb0ViusIa8xANHRe
fv2AaRR58Uu6UiGaKN7XqT46eU52p5Co9qT8jBOh8jCCmscKQSPPKL9GQiqQiA6Tlt+QjccdnLAc
1VeYhXMfrR/Pq3wXstjZyi4Vl2y+qSzLvqCMjW7S1ale5X51MVN1c4dy8Jm+9oHag1QvDPXZTGS8
BO4fA+SvvbDrFDA2zlgh1/ffNelFGO2h4uY9oS7lTClkT83P2fcYuTk/43I5bfx3WA0m9sF+ebiU
kcabRCBLHBXbejTljsMoC75g8Dq8ES0Sf7Umxyle/W2mjJ2TbppEhvGezW1TCzOyQ60G0PzX91YX
YISXlr53TAWE6XHPP+s9oPo7Q/ncbm2U+OJY/LGsHLdVEO/X1yDbYRS1JYJ52Usy58bhp4RyA8WJ
fbgwq9S24BO+ABxSadXt8HGRwbtkp/2fe5u9+ay79z5zOBctC5CD+riSyE/aJm+tyA2nAeALufgV
ByUNyfj/ys5XzSg3t/HJJgyz4/D7XCwerMcVio1fh7ryuliMkoYEcMCkfw19ZrmRBOXQ0IXxc80L
7fxVkUYXxn9k9KzGD0q5czcZGXoGi4taGn2GZYdDnTb6141S9AJj1aANU35AwHBp48MU/kUluluW
ILuVUnPTwbZy9oc8QzzpNftDXgQQLlWtJIEzCrkoie9gRZjJOIWgZ9LumdsU4OUKbTQ7iuvQxtKc
95FmZlWwBts4zwBm83l9EZ4d1CPhWBV67XPvkpecio9a9exywtAtILf5FyueS8Q+XpEk8lA226eZ
POAKArSHggXegHHt2wb5hFQpFCU+8gTnQ0vaNiviXeAtNF+AX2sZqfM3iqzVJYqUJaXpUkoncY00
A1y3rLRTu1jtTexW/EB4b+kI9fFKnJ9zJRchhnJ7vlUqvuTwc1RtlQ9ceErlmqK20KfBgfKWxhaG
HKwRCUOm4RgpqjCuzNg3jmO4MWC6ewKlUIDcbARQ461sV2ibbidFj82Nc4SdPg3Np4WbZPnYKo44
xhUdkJFVWJGmUaU1vNgj5hCWbwRMXKHTUxlJlth0fh4gfLm5XQuzCI9YmNG3gwOpiBgm6cP++pui
1hazB/V2ohaoGLPSjLKifeN4lTVK+DgvSJItnsbWCJtbACDq26xGXZmXKB4Qob+eSzDjaTKMSiA4
0chL1fSOEFv5EGeACIgpIKYNC+0UO9se+exSaCvUFuaGLdOrOn1MdftTXX9iI0y+amZ+41uVR0kK
/l+/HdoSrrBPdLYNg0s+lHEEEptcE55ivTmjaoGtd0PMlGwGfANsjC2KQG480SUTb53G1bbwSrI6
BcCkj0/pj6lbcEMl/iGj0zYnToMsyXA9MeBXwUsKmRcy87ar94+i4HbPW1IA/PeTBPVEG3LSLO8O
U9eLfUFmdiwBGJ5E07q66U3/fUnafLJOAIzFELjmQrMyvousz+9F/FGxjoO0dSWf97CvJ9BNPq5i
e101w7jjJ6ZIgcETMuDmnlUHFxd+slBydxpGcPeQhhcUV1sjXzHmwGxybywiHNpCy3Am1SD6R4zR
UOrpQQlxTKYcYlIxacOmgFOJSRILpGnHKjGuqn0ubKb2T3vim6JdZdahFV2mrFMu6rIZgjb4aEWD
wVwT1H4/K7HbCsV8hvZRla0E1H/DXEvI1qia+wy1JKUU8VT/0WoQc1eYeBw/kMwyMGk742iKxe12
hHmQwIuHP9apoIwPgpeQ8xtbCDrUmU4mayHwPgP9MdbO+CQobp75hnz4HS/grdLJgatFO2UcKtF0
n5tzL5Zglg15xeHSmfhExHRI+j4wUy9caqtUFupiv7wRh+CkqHP0M/AWLlQ0Kw45Pt8j4oZZQ9+b
SNYbfxH1Wb+udfLinu//2hkFo15zGWJKvo+nnkc641oFRYR8oghZT+kJsDh1Xq9DyUgLkCqMophI
D7JdhGwgaWmOfCJKXSGtP5HdHuGTjYT376b2klUeRZXMljBnu5BmJV6r1gmdM16vT695KQaI1kcs
dwGQLene9ROU1ROhHKvdO90wpvSB+7Z7XONdsB7KjFFo+bn3JHBEtPSUEYAxigq4iV1mLP+VIm84
+E11A3f+ch17fdqQ1jPrZT7ugtHDgiT3tH9wJaWbPy0XgD5CN7yUaCsPHBAdTTFKOYhW4fkeYGMx
x4oRkLrRdk3tQ21EbhYoZBcSMLQTb3Ei3UwkLTMLOLeNcqYkIuiixTQGZlXAYR4AT2KW3az3VT5Q
kie+cGZkUBBCRCgDIjkOfBbSIh++IjUsm/W4pvx1QlTZJyj56W+oiwDjEFrvJZUteoIBaPurgjSZ
5LGTPxmzbw1rn8viWFvNCGIky38Hp7LxxIeJuRJpD4qY9uVHntu4NjLwN3/lzD0BcpDM4oRCCgN7
KfqB3idG76ntqBVgJzRvLNyyAWu147SJd2+l9hDPaDPvfPLmlOJbrMuN+HInSh2W+k22Bc0GIDuA
spFo3FrvEqS3UWv5AOpY5Ke7A4hnUgur6ulhZ+5AlsHzWfEjF3uCjNqzn/0QB/PdloFj4UF4djZ3
tnYUDDm9KUbVVFuvAlvzwjAhX+6W/RlA1o9e5roZG5brQV4fzyCklpPZuIaY6Fbjd3VGS+lmLOvZ
3ZwVNxxxB52B0yqz4mT8DrpcGcm2mqmyoRQCZqIEiyy9YIVhF4vUh91Hhs12xP59syrKEIEGxQQY
IN2dYJHdwEsCL0ke82EIr2fkq1CfpgrNcAekg40BmX5L1KoSo116f1Tt9yMilNRfWxHGlUk6uMGX
KLlSPHonxRMUOAXw8vT5/sCEJ31cyc8VaurphE1QhDVkO6cbEq7pl3ehU1+cv67VsE549kAIWB1I
F65vzXagXZtUlDWuHUwqVexmkvidKSZLFoAzWu4og4OEKzND2aqHRrKMOFQ2meyZXMqrXPHyfPN7
y2Yofs66nxGT+cZArmLD8cjx1Rl4J+Fohu7lKby+D6uT8w9PUVerd4+g4n20+1qCBApibJLepApZ
qdxJs0zCzqQox2SEcjUDdNV7LZenOWkLhVaneiXhDUUgUsFC5OfMtMhkbDiRIQNXETsKfFtU+TbK
v/KvOLtuzKqf9XoFi2hbVa9YGVoKnBQ7vB5JFcHAUT93xU/8vsUVfRL8CSbQFQusU8C7NcMnhcAl
TnFW0SKXm2TEKixuAtRG6GO2Au4mGhbL4HxhPlzKcM34Jd5tfDA+Gd2nfjUYaGmho/+ca89JoAmx
KiCeGw9Uem4CtX94LIiW2hq1HNvfJopIfGwmGZS4rpYUB8JWtiLWvyzcZGcGToDWufsd+GRCK5xv
ZQKKIXtY/t2S1TPX0s92qJuAXNrhrA2UdLqOWkDQajWOK+L9IIrXMgAMIvU6QauGma2JP06F6EoQ
yuBYjgyBENW9v4Dd2OZJRYz+/CoprwE0r9MVCo63XafGOeKqd/Ub5C+JanWeX/zkRAPx23LyNCD/
f2kZm2u4OJK/aBB2PjVDRUWRrtoOq/bJHyQWEfl8rBDEUyN0fl7VNb1jqnUbShFW2o2yU9oCEthv
9nUb/KHGFDUsUfPJyjwvKBPScOc6XlfXCOVKNmrpAQzGzDB4ZZ8irCYADAEK1+btMEjQGoNYJFmP
ZXgBKbinVTe35J8w9eNvX+Udtu5BdyguV2RqVWnhGQbx8U+vqKta277tgHQz8xbHbB6ajKj2NiSk
DrdRzIgZRza1dxrmWTRj28vKOiWf48k9aMx7xCAevTmjjQrmDjY7/w7qfhUiN4QXp5N1ItivJB2/
m0s1AjzieSnGhcGV2NCx2MDc9FDsaj3FQbOriSCOSySEnbFJb39sKphTtaInS1jKlzTTetTLD2+k
7Q1IfpUr4lpvTCrHUVosJCgrerTHL+BAm20sNAQEOiUTgaLH/lhXwW5R3JLjim9ZPs0TDhkk9Vxf
F1V4/FPPEAjf8ZAz3sczoxHdU3L19p+ea2ynEWAnffo2QAwOkDeK/isTYEXdPlkkBjK8pPj2LD3e
ck87pP3casoVj0kbzeGlX/Wn0mZrmYOQ/4iAoW0H+hDq5JTu1n/t5QZQOPAMP8Z49QLUl+U0GkgG
YtBE+1LjKsZqOxk8Jo37ZsnHrjc8/rHAgNZPDebExqEpn0oJ/PQcLxUOD2mLY1r/A7dL2W6nJKuu
wp4EUuTuNJz4gsHgK85bD9BEu8nxCS7aUSIL2sogWORSKcdfpBXdac+lVTA2tFQfiP7Pd7PxZwYg
7A9Us1n+1GMqNVvwFT4UKGiCYbKhvIGC8GS0W7sIB+UhoiLsBuUX7pTpJEhCSVUQkGqz03L5xTid
eVg90HYb296lcQN5VlfpHnlRvKzmkIoQBGGlcyerLWA+lOUUhD0SQPfHcawR2NFPPU9dxLF1RJnN
C+ERWd5pq3o4cm7vF9jYEbLfH2xJCBbbQMBGu6nxXQzoSl3sVYD1KhF2S6B+ytliWePSaT1oMl02
S8n9zA+Q+Y68BlV5iE1WqMlRZA29Pujcf7WrvIAcUVhgNijqBMVstFxYF6NGVgyhbOFepZkj1X9d
5XXkcIor87TFTPxH/weZzNbwlQkItklf6y8jRtJZ71eCCKIqRKLIVs1VIQJ+xI2AB/LUZWnBQrDr
AhSz8TGpOE1Ufng6fKb9zq5NFyS2nSDP2S5x1WgNqwwnvxMRXlhl1sMfVm16palEoMmZfpk4QcjS
Gt040McVnYLF+rnHGaM9Gea5VPAxnTIEOG41vhNlBEsXf3ZSwiRZOq/+iFtuXQQmYTGuj+IxOM6W
x3p99bLiVvCGy7q/lPS2lJVyNhaiLvBWj/r4no4xmcbIwVXTu96Ult5/IGbpSnO68+tt91Fz3F4K
X3etHVAjWO29NT+rTBx2LQBbRh8RANXQVPkUn8o37bfGWR8/Cwcqv4M7cs7yKl08jaF1r2vXXGiF
DmpQtZP/Q4C14NACR28GbWTpC9btza+Umrn2B4N4lADhlbODaMmnBsg4xV7sKjfX7o/OkDlKCX/d
/M9rDDMHTdhyTTA+8UcDjwI+luN55PaufwyzCIHxDubMJiJw87YwpwPb07iItsnNr5h6mlPdkPnH
S9O8BvVv2hL1Ls77t6cowvbLrDuKHYgvwpRNk+1p9U6RSpbFsbqfcKT2p9jCsvIx3dG9Eq/lHuBa
cB0WURU2FalGhLEwwTwrRlvdUbMDoTQc3KJL8gFqrnmPKgRrJFEXegdtJe7LD968qSZeAh0OW7LQ
n01awlUBjojkbZjMCcGUx4Xahp4HkKeoHP1ZnW+Yl8uyrBG/rqEW0RLf7+sk6LnGw4zwDlVcVws/
oiXwz52LCeLNI+0aP/wUaVgTwncKIgr4hyvhgcBdtsZ0IYdmuOPfWqH8Gnm08oThcy/eLsJ0t6Bo
HknPbnx0Yhj+QLPF3UE/F4Pcl04dE46tHMn0WJ3FgjvCnnfJTfFrqkjTm2726BOZmmumLsj1tY96
RRA7SUTmB3MwDKwGuLGDoLhWTIHOHA+GS3c2l7RJcFxEVfNuGmZx14D6OXqDtJKMs5q7pCcIrsmJ
fBrt0JbQOCqwEBNaFSVl+FxL2yumRuLNUfq/FrqIUsJ0lg4WybUkRjBRzX2nUgm4kmXAM97bw8yc
YivvyffsLpIC5ZsZXiB5a22h3eGdVVb/EzpngNHVPgqWYko82mGqW7zu7QZZ6G+mcTyidZJheJ5x
lqbE04SKzMfB/OvH4EULi/btTweOahkmnuMdLrn5cPOmMdVy/Qwslsr4GDVaUzqkNtc8M1ROBbwA
BQzap1efIluVA9oy9odGtzL1vooxVs8CvIgj9jfV0ZhJ/gfK1hc3NS3a4pwcdT7iVKAvbCISd2RR
r+IM6yAZ7rLXxWXHK03gFJ8YX3QxlXehYYc3VnjFBZUkw483bK45bdwXflThBWvGNUbdAkpD95hG
8i8RuyKxdGtF48X548Xsru7SyMZ4990Cg3tLVdA0qvha/Id+928K6uOHyCG/lI5WTyVn5iT2hLeB
y2cdmKrN/23ZXbaqAuaUKB7Ht8xwqzx0N8JMjIt/alNneKLL3THKvPoZcbxbGt5O9YslktIk66o4
nuJK8tyL3jXy2YrVXUJZUjd5Tmxev2oUVhaHSTLApwkE73s0Xw9MMVeQJcBP11QtzTIXoj6k+rwS
agJ03+tkVwZsDLquV1eG/2Iqeskzy5VwdOqGNVbn59GnHH6HNhpecZPkEICTZ7HwKGDikRKDnoIw
r/2NqThmrojecWegitN1Xd9mqpHWdbbkh7vaINNu5G6HVKyUMv/Su+Ao58gnce8HzpPwj6XvXe3/
GNvu53F96Bau4wJq436kyiBEQr8su+3T1eK68KTpvsqfPrsWQLllsY6u+ZgMKC+NQrRxNmT/ampl
fprybv+nGIMlq0syViFFS8QhK9m+bPG4Y+GsI9GU+kCFDhqxjR35pnkVVh9Da6kSaBy60efT1HJ9
nePxgOfeH6BGEtwnC1M38z+3AOjkDDKicVALPb5jIfiWtdDbNHCPsfcW7gDDCIjh65/8gI/a6lud
cMPhmOfAG7QfS6so1zzTAs9yb/P/3Cq+0EmPEVJxNEhLKGMUMKd2I4tAvllEitPZTVgFV+TrgTzm
t+8YVL6Yae9+1DzzutNf/Yq6NG8AC4fawkINnjZ5VJQQGoIlb2flpRrE8KYz8k0iOaQh7OfdXO98
whdapZpClbefygRkqisw247hoPlynXqXV59Ky+6uDQw9O84/Q/dlVFuV/jjBH1nEHWpW89hQzK4t
U+NCTzhqAjEq0hvOR26+3TftfZnayX+ud4eo+96f5wSmNBB0UBNme1QHnogu6lFayzKjNOaoQRcG
uP6sRSEVaQK6DmG7FEHT8Rg2wtigRjVoTwLMxOXkMo5w2agcSj4Sddwc4Slb4CkhPX+J8BgXFBRf
btx7rDz40oDN5kKj9RQQSQTh6eKzpfsm14x8QmD1uOLdAxGCISmqVY6GcMnDBdSHFUFKgqdABbq+
CdpdyQ4CFSUoJTYs5dumFnQH3iN7cs7QleV5DMUbP4R2Yy1FLrzjFdPkhpSWtVS+dHC9Nz9ZNM16
28Kvhspw8aOkKZ/9MWUwo26YtNwpfgTBYucH80gk90vuDoCZSe3rvTeH2ZoXuzqELtohmzv3d34h
XPl/AzD3Uqm6qGkuS6/B/JWR07Heo6AdWFLaZr8tfKGSCOS7uT3qeJ19CVFVdN/bEuhrfGCeu/pU
hZzRJzgowkSznXom2Eu1/YALp3/+R+I4GryRhZTOXKV3Gv3Sj0F5M+uX5w2HUdAEzIzSknm8DZOO
6harQWlUbBKXj/QCw9dMyYru0WX3EdCOB3xLUHATPDlXdtksYZT0MaIdBwyzQen0JS0L8PCqsVlL
Vs1KCX+McPkXyVAmQzytz1GFPTFUaHhfDYeOypNe9VZlKoABUNcJN56XvE4PSM2Vs0K1+QjfMa9V
MgSXmCQUIXNzwUdrrjN6zw87BmzQq+TzkDKHD9cT3lp4P5ekAzi6PwyiWUzOXHzrThzlaIYW09/9
RJEKmGzt1E2xF+UqhGn90f494MPv9a6B5/BIpjJ2oNSaC5cMTS92guTUXmpZcCtoHYnrQa945FJr
wMHLf2qjptQSNhoJsZhtO+cnBEaT14KPZHd28BEoRHOREkrQm3fu72SGZub3/flTqEeArIj5g/uV
EkIPcYm4Nesf/PLfiUX7OgvLtiNaw3RFheRdr/ilXrchqeFio4D8v1Q/lrWEILka5lyZm9PQfzE4
pI73IEnlV9qf+pvsGQbJW3Jz0ZaBS2XDPAjO1zIUaZR5UJsR4UC6fnMRWciduyWDHNlHeT0WW6J8
sOMsV49S0Ve90SdM/I5YoJa/yKDSt34V4MlQxxBJNvUZ9rl5iYPIBgux7+xfILenteVSUWDH+hh7
1Ct9L7rpl+OZiIm2rTpQXyXIX5dNJIvBZslSMGfDCK2ALLJoRXI0WHp8n/C2mCN2NFK2DnhDjyNm
zo7BqU6eHUbU4eR3ETpSXMR3hRBM3YUkscy3U8amxRcwKe/yUj3TcVion7jWYcmlXON6+gInBcqQ
RTKWldTLZf1VyFBSGmNagO0UwWTvc81T9uPFQMxZ7An6aYpX6p9jgXr/68vWFQnAz8HxJwCFTw+t
e7sUkYOOOJS8CG7JPdo2NYRzipejmMcgB6kRbylWBqM1Lu/3YElogjCBPuCSjxCA5kY20SPdF4kQ
fANjB430aaKoy91RpyiRqJlH751vhMNH+sU7lnKANnJbOAq0xAh/0s98LUrnkSa489BCmZDKmhdd
W4sC0XbqqiPiZOeJWzOVd86qpXCCQ+U+RlB/o59mQ1zVY85lvBEeBA/dc53gFVF9aE5palueh58K
EiedD+rEyGtA/1SbTzeVOvhZ/YcG/VctXXXKB5l0J8PPrHfnEbgkTh2XyM2F4nz1yuEYubbvAahr
FfIFR8N/aQt7Zn2UrIe+PJ094N1C5nbXKT6gDQbqJP6P65lZa6RKUJqF5UetDrkn10C6d8VVQiQH
JnDiJ3y6Qr/rwQdNjlO8RE5PTp5GJCsftXNVInDXnclVEsZN1FYgCdPTUDsrxMAxTG+uGnE/LxDN
MdHbEER1x7i87x2ME9RWe3R+SLOurCNqPqI3Tqg/FxrYlxx6AbpEfgNr3Htku6wvHcBllVM27t7O
elytCaDSbaMfk0Q4V0z76Hbo4jA4XJXkeMs9FusSGtN5FxSgGoMG+g5IFKl9SkSCPYVVAwsuYu7W
vt9y5eSfceNBAkZxdIBIUCvEvTpMr0qjuGiYGUCZ1j+Zss8SzpC3X1/wimSfFzYKPqLfDuxQ4b19
ZYNAiASLnss1e7XzVMpJ6I1n9oMaaKounolnPWkGo5QKXPgMNy8NHeSJjLIOw0Fao6eACLMReZxC
65EslQNwzRnJPWFfrwAcK3Kp0W9IDEmIvvTQp9nVJ/9xmMwGp8wx0ecgSUW5/t1pX540NoNUUe9z
Q+cqZ3UOqRLtbIzSOQOZCrrV9ZZ3kWBckeqAWcJDGpAxAlcwvIkLbATqyvO79utr2IJ0bSoJG2BX
M9/Hevwmpg18YZO1Y8HxG6C9X6jrtHgjLOT8f3/u9AKrs9GZny3kUY9zfBfCOPTVKpaU20YXzaMA
muxllGx2fatNppy5Pj2dSOrY0RKHIlKhg59LnVUUahY9dYMdPW1Zqe0YULFgnKy/EnhT8huDU1x4
xcqj/s87gkeUzYW4luPrCoGm8knNk7ncWK9jCIvIKpv/N69f9+0RrboNlqB9I1TfZNVzAePd1cFs
0SE6XqY7Oe2rQfxrExcyyWTb6zK/SPwVrripZRQUvK5nEQq9+4OaU25sGfgTV+QqU3xbU1mhb7k9
2C5nFWi8QDcN7oq9fDF40/OtMVbe1h3zVPS6feiz04/2uzdtaw01t30bbZRl3xvaqzUVlq7+UN5t
LJsE373dYIyAcDkG+aT0PsACzl5xmK8UJ5k46Cqu+BnurQsPF8Hb+6prDjcPUc6nm7mcqTNmM78g
FhMoP2m0kcGIVhHmIecr+EX6H/ptoRvKKxMXUUHFbN+Gbz3ezofNYpV/UDUHabkU0ViKYkuKH9Qv
1VMirRe2C7l2OICWSI4JlxCPfcXrWRvKlHLdnagbQDeR9NfeStb96kU12zX1amvDzp43QYy6nMbF
I498dNGgaVtKnH1TaLlnsG+0IurrJjxGDc7A8SVQVM5Of7R03urdXlCbpAxrib+6GcTtXrjm0g8l
d7aNfRZ8lHFC3JapJQ03g4mTgbRw5aQspTyXo50yLTf3sFlgTNfLwH9/fmNdtpUW8S2zvG+EyfpR
qUA73pza8u7RNQfMew9Si6v0kF+yC7Cq487lYnMQElbLqd/nLI1aBN10OCjCKkY6J9QscwmFLSC8
cHFqTKGdymj31Q0kajcFEPU0N2Tw5wKnT7aaLLLJAD5z491/1BiDnPN8mL++hoI1f1hLbZ4hmfUN
+M0nRscRlucsJ+5jVgQSK8QBbCwYSuLSWaunaj0iWUJ6VngBLH5EyxXvDD0aaQ/JJglANGv3f96L
YpNKSKsCwsb1mgA+VyKXdw/B+dN/i+U253PV3KkEo+ixa9Fiz8d0h5sF1V+QevAUEjpeNEuEGMNr
kABqaaQPGOJWcSEgsNe90i0i+vEe7sR6f79Ocko5QYrHiAZHWg/JkG7oPAXOxCX1DjoXtrykPYJa
gn1x1zTn1rX0aVPoZgifbw7Ioyom3cMO2UAbdgaOnXRzcqykEtE6BBEu27lslbUOTI7Q6uO1ec29
MTHJxSqkDQ5EAe8+U8xmipcNVVIRPzUgqKh0NpbPwXy0SYbyogjgbHhGcmvDlHx0lDDWt2P+82V0
Imik/34Ag+jckMhGvrjyY9zqJDcAGW9W6oLnXYrKfKYiX7Gmtc7POqcBwiMYhz59o0Q1Ruh8YFEc
c7zd7VPwo8IEy0xubzm8zCAH91vmHdURV/BeVY5PIIk4CRK06FP/uvMBCOYzu415yCANn+AFtaJV
Mavbv53PMMdkA10vxlOHHPVbkk2oPSlmI1jXE+jTGZ/15CSCF8oIV79HPi4+ZWjfnaEYF2shYiRJ
kokZxVGZK3lDO+KDixpFsxz6KqpK8W4DGFOR3JagLg6BzVHpGi/vl0HQ9LMBLb4XpaukH+bYfzOy
1BCSGlJENVDrQIh2ZmNBBcHrYrZrorYn0bS87ir+8/DuUrlbr9ayKU4WwHWTADB1t8MGBEBkXvW0
RIyCw1tljgcCVzcHlT1N6Rjity4sre1GTe6gO7Xg5G7u48Tjm0gJDUemn24cVhu1Ou2naSNMDQmK
LAxa2Q3Qk/uFORoFk+9aYi4KB/NepgJCZlwylj782KqAgVGrPnC17qdeEDpQEM1OroWuBLAX9MSO
BjD7jShNKz159TTDuFY9x2id05F6WOlgdobs5N+9zYCD7TggRCEpiAeri3UdvBRGuEjBW13NVYkU
29d6VYEmEAvhj/K26r1p6T0WmAhotJEu4uVz5jD6rF+eaNrSO4k1jYtRdRHFoDRZhmTKvqnhXgkL
AP/kpHCrSr6iJ3zzNWdXlcrLxxm+gVuSDgnqEinrVpWw0bd0IkAhujn7DWpJkp8AUwr1P6xQQLwp
0ZzISymlYmAvnac2GTG9NZBwEg+umuChwST8GcdQzDhwaRvObe1sXttiXMkzZM1RNoOZAEuQ31EM
3ygHphZzUZASvbhz6xCSJhqXdMECS1edCVA4ifJec+8oG2/27aNftIz3wqpyHp+K+Ks38FsuCz+5
TPVj2Nuc3YbENHReqB8Lcs7TUoOMHXeSuXmwh+1wT2MXczl5WY1O39zUH2ZT7P8x/bg+nYWrxpmQ
UM+w8nMOMdr0fzxGO/q7QW+qp10q3CKgD0RATJSD/JSGyw0BAxaqd7Uv2z9zhFDOjGwLCaODe73y
HsSxsf3qzDWHRiXx4xqo2ECBb6VTUzVY9ECSlbd1Xep80rzSVe2RSUPdIZ2bb7h5WbMuHFwD26io
AzMFQMbwLS74ZogSa/rmD2kaLEeUgMqz/vbNy6MogKhsMwod4xBx8wxY8QotbRd83fsfq358z9tg
DyEtld3N4VtIZ1dfZhtkvnJFy8XF8fE1y8O33MtO02703gFH3n/SlPHGt+f9JuO+co2YhOmftuVD
wpu/bFSrHeApUaIxJY7TLIqtVe8TDmyA8QMYE5sfV5hrA9qITVb3YcOmY0mTDnAyfvYva0ct6Jnb
tzbE2rX0lUkm1VsEX7fhNrahyID2yGdqAw5ezuQn6U2gTAoPiqGStJMcDIlYJTgqwNdY+h7McpOb
LQwfN0Xt7e1vBnG0J3nAzVRw8Kq7A0JGJRyPMkLNWQ6AxpbIUfNV/2I9TQRR0qgmE7Z0TF1lmMHk
ds+gwGzAQ6fmkI5R+mQH8ZzVHkzRY3y6rfyfFdu8n3hBhcZczAlZGUYyZxG6v+9EPV5O6g+gxexc
PP7i9PAXyUJjkjv6VzQZNjt73FSMYowtzA/32SshmJoGwqrkDmGriFsiBiikm7HnJhJ0unDr7wk8
BNXtd1lWtAjwMUVduEX8ynCUk6iOvs3k/9VkqN78Z7nrCAyHIWKccPEV+dF3fpjp4QlSOdKcAg0Q
GF6zo5QbP62vjbWgMT7Ga7WhkIxtmvK5m9X0tCDGSCxEpCdSxav0dy06SlpE40R4i70v2OlxMKC7
l0HhNQku9v05N6vXAwe7YZud6gouPOK/pDyi96fSiTaLR+ZeeaiQq9ts37TxDJPs65sqlbp+0vhR
TnCyfDlJ/z725gu5HEcBBwmDmafBZ3sz1JTwbU0xvG7K7dWvrYCbHyZ1gLvmmUJoNW3BrTOOj0Ba
R6E95HHMiw123Ab2/12Nu6z+NN1y+Yt4zIApi+V/uRu16YlSiukkn1jNZOnx5afMSTYLz01qIOHL
ntt08viesR5JORNjX8uyO1BcDdHg7VhV94xN9KcrituJs3JIJXaroH9Gz0nKodcVaxzR/8nIA8Dw
ov0EkJn1y5UoXRKaKRipmh+UPthH/Ui8jl/LW27+QRezIMs3yfYr2zTPHxRJxa1wcufpqNM44mjW
vkr9cRSueBtlVxrKorJjrz+fLREiF3PERbZlsBU1KEIH1p4RX1xlK8PE344uLDIi/Aafc/FizJ0m
9JSHOeBFEo8XgvbQviA39mEOf1tcE2V9NkSlMMeg22fVRDb+588YXSbHLS78LLfh12vS8zdLcn67
mC7ueJZ+5P6XKSCTICO3Kc4DYsGyENWZQctckFpuzsEyS1ohnBABMdqQoyDLJc6O2tuDmCWeujfq
4te64nyt+C3o5dpmirKU7iUou+DqJwivt1lv2fILiT6ji+qf3kJe105ttkHras6QSK3RXLVNac99
Iav+Q7yza2HTiDd2vZCzY+4JjIY6Z/pmRsci26+0B/xMgwH+1cOKQfUVC0u56UUqU5OYTWEcXCAC
GHJsVNAy4FjMXjdnzZq2B93AJ+w1thCBD4rCzWS9KDX4JrBaDWvw0YImbKqiZXN01WbYAZ0fI5HD
IpHjKgxQSZKWIIjM7KziwvHUYpCkbISoZoUeYwmYtf+6DgJ1sQuhZg+Pzep1bnNOfuK07AD1ZR2C
YRojOztY1ODhreROb+6CXSNaxH/2sZxmQFadMy+K5EpMqZD/vmKlJzdeHBLOCCrItB0589jEdrtL
ysByBSDI/RDz9GBEM08Q6uiviJIiNrS7ykwqh6+NS+Yhf9rjVtLdb4W+0YyDpaj7B4Lpm4UPMT4Z
bg9Q/ui6VMsDZvfDrFXZvM1BYp8y/Mi+haUTrgY3xqKNckDagHsixtIY2IuaEITuiO1ww+yDqQRq
mjgbDkjKUMv0x7WgFSTtdpY7bE0x+ObWZ7fAA59HlCrrtciHbQzOzx5GIz9Wh5G72XVYApnfs1+k
FtFk8Yh+8SrtJxQ0+1GFNjk/4R9a30MYLjgUKqg7/xp5op3X3zknfcQiat47o3JqUK2hRum7h2ND
IaUVOOJ2mfMV03SErm3fJvpedcxdgP5/+KcrtnFE8c3M5so/UBtUJcCMtd6BUlKg+dog+esdKRyZ
+z1vp6ThVXQppeP3tKwapbNoG+PNc/sr8EIbIeOW9MAZZnlxIH2ma7YLe/lK5xyzN1HMS3jpYNig
rsJ0IjSaLMBmiGxEFHMw6jPxICa1nZKyjV/7BcS5YogqfSnSCAYWdDo++kbvjYeFGOBw6LuN/GUy
2Aio3zSCfRcQneH//JoxHzotvluX/glBfv/0/iEfXejc90daaj5sTypnw01BqG/29vzCo/TOdkuG
a3/WbDScIRmMKpg2dJ9o4dNYKU29LF9T8ObE2mD/oG+s1YfHxqHyXddO41ZC0CiSW8A4B3iPRU0F
mwvjjzZSuVbSvYiNAr4RJ2hFT7LhI5noejJOQ21u8vezXPJVgNvrsa+hkPJGcD9qM2zpKh01nvPU
h4+ZlsBdp7aHBNlabyROBaSF7WYY+yzZdFMU+kVs8UWSZTUfndForjRIYBolRzIb1p/0wosfX2fY
A5s0PTUm/sG6o2l5UEgI4uUmChJyE63vvVExwfeQPfpvZRtka81PUWI23b60ebvnkQ/Dzcu8q1W9
bXhSpRn9+o6TnXzTYZVi4YllJEkYe/UoCuk9f72FX3K5wuW1Ub49rswKoFDbIXKGEJn2aHLe+xGj
R22js/jPQLzzrr7MKyJ/i+8kVON2qyTtXe/X5SxZ73OETunWvZ0KJT1us81wJccBCXfp+nidESbe
IkTKxBg6AgUeua6dgF1J65LuYFkOA/ligDdrFYXFlECYVTVw9IfzdRiYofpaxc6KZyDvKs3lPOPv
DjxPeSOO6wwLIMCtmd4qBXl/Zc64X07Ym/CAkPJFcGH37GAd3P2FTwDzC6lgZKxLng4DeHImWkxv
zQ26u5y4wJ9rNKoaZc6uAASLRktJn5OFaVlIIJezdytP+vGRTIgSNi907pbYv681phab5mH2pgdC
A/ULnhA8zQfaWhWs1ixJu4JkiWkw7IPjnAUdkkNT3O0h0JMkv5TexS+liCzyppE6pKtdHYXsDYed
KHJWNExLvAnMlnFC1c3FAIOI9VD06wCQz+JlnGa+CGMrier47ar1WvkXdUg0DMkTJMTZwY63WkIw
bWpdcRTcqINry9vlbGXdMnM+tilfVCIBsX36ck0MdFJLNZw7R2LQMUb+fhHa7sPLirLNj8B8t6q+
Y3X3EYTYUUESYYbi2M/st5tVp0MKWl36qjp1bfxh0EfH7/Ck8QVP6ndJ3/VvsFetl1AdEn0GkBKb
kvbBrDvGa0nNhXs2OHgaL2LdI8KmjVKPafEzeFR9F3PL7Nz9yoQcjM1HDH9QNsqjeOMQ4eJ7hMwn
2FSoSu607ackCOMqqal8Wc7BUu8cABg1cgFZt0K13j6npwPz8ZPAKSX3gcdKtUt/sUReQgkD6qLk
I8Slu7y6LcT/+eair3eB6GsMCTVtc3pKwPt122miAvtlby0vQIa3D0w6cRwjWFRza0ml85sxg9MH
+iDU0ZYjRO1Dfx4PtbObjcGtRLGQpszh+Mipwd5bestWaTVscOqRGCb1QAgstJVA3D+yd8E5YpD1
MZLvMHyfNgLT/pekP0glUOAJflpGgf3Dk8bjos7/AHoONy7opiFq6zYc2pQ3vn4GZcNTXwK3NMfY
pwMos9pj2LG75XX833aTWcn1yl0lSOokkPFlNlsPR+1bAjuJ/wJ0PnsCmlCTUmVW+n4dHs9ZOnps
LMBXp6e7izYFKzBpFFJ8QGy/wNtYaAACP5+SZj+DkIkOEFkZhU6d5FjljlAlRdL4f6xvB1rO632I
J3bkv6E42vX9Q4uxhbKfPQiERKKRkS3AYPnseU7op3hmfoh5G6zMVoypYrjsFJhYw3vNJtu5c3v5
wlNSE8zh4nDmedQjbagELW0E/gd4DqfOKUY6N0BtgtLWJVijWFkXNMonppFYxTZmmGCWvJz42r2T
11Ept7YQvnb6EoXiKsSyW6K2netCv09j4uMU457ISWeVy/d3lM3eajp+KG7kCzROCD4P6w0UD/+g
cU5NMVpZhFn8A4o45TcBJu9RTcD9es5rdeL94TdtBG/vW18vRbBqdy14VFu/wtG2orxO6rCgbbcw
9Dt+rChCJQYjdoWwRKDyMAhzet8jn84yJrTDlajoE4/0t+lSljNd9klktiShXVLGIyV6Rdpp7adL
yZgKVfuRGKKnmb/6UKZxFVo+bu5mdioK0HAwxZ1xb0vUmswrgTcHNQ+6NQOHCjopDmW0iqTjGsBC
lu4FAX0+SKaFW05xJNVzi6Ck6ZfM8P0cI5UtLI4MRd05wwBLQoFtiNibwwvCg98NmGUE+cQHTUks
LtIQMvI98WRYbTy7dsUXoNWtufEUOjWk9OoT7YUl4r9ySftevEEwLbuwY7rAi2ZVvY18bseDTw5l
x/AD6NOlcd8jCDboWtKh5OchDc6oX+dumyU4ZkKSnpQXiIH11UKpIeNePsqh4a0NyMCpb1jjnwK1
NMWdyEVXAJ9TtpOLiMaTz7sk0JbPIzoNFPJv0fz3Mm65313ANtKiFy9F0P849pF2zoTANsv1gyCe
3J4zBaYKowY8OI15kEbQnIaVbKO2+Gdm04Xyp1qe13LCp9njp2LqM9s8JDK+6JhXiS1jhucqhjz0
zn1IqVYqwmRe+UTtAOzcwZITvk7o1EvBUJVorMhw9EiNEXbLPnCiB5g28K5C2MkGphjP9vrJadEJ
MmkbL8CHGbZO9EHx0N/4hIozLvkc0fX8SBrNsgOliXU6d7PROqC1EtL7hERSvZZaQmbJS/CtoSrM
4aczT53NqOR76TgJJAkwK8F88NICJUgsAC6ABVzLVrXFOd77f74VYJgQoITtisU3998q2RBhYBji
962vJ2eQN1uoFUStRlQoB0p6Y1dW4XVhI+ixGx96D5lDGCYK2pfMnvobQmgy+8XTqOMSnCYA1omG
CZ46GCpV7mXng1yb48dAUReYXIDTbVyW8SMyT7ILhB+eZJWwIt0ALLhk/el/HLWE4rDCfsq3wnUa
DY2/3WFSZM2FlbGLEK/F1AZ83GAZqkuciqKi5FTmuDUsiwZH4/E/1aA+wySBS2Vrpdhn7K+cvD07
4aYRoGp/AJ9QTVI4zPPs1oGHtJ0O5Moa3sVD6D3P0gNZTot3cXZ/+1V6xagm8DssNy/5pkdYuPf8
XUKGi7KgDVvTdCrw3A1R9hX4xTEMQyQATGlSOQWyxY3uQ0lAnr70V7c3jH8hWUKZ9qAqw3zuqmgG
EjsbH04TF3P7rLAxGCbJP4dE193Nv3QzmKYFkhxJPRjZHQPjP0lIjvK6GJQ1IojE5Kk4I6rLxQCw
FXrBIVgoVTMJaBlW4rXwj8e6pw7Snb29Qtr3JIcjXujbm3XGNnnsypAGPOMG/z4FJ4MEitqADXdM
0ss5TuesL6/ZpAvCwjabMXuLal/k98TaUvZzxnEtmat6G2yaXHlogbUbfxt6kj7Z/ViYni4TYo8t
5awrXpJkpVn1n4erxLUacv4409RRtrRUmAp8EGESTSrNP4thKaaIf6QtEY1vyV8QlsyHEnvHPaGy
qc1BSkunFtkrF4mHPXCCviE5NZ3/eX9/dr4iYFb0vn8swjMaSSZf4hqdEt4ZiDL075pZSHwmr1aT
qQX5aPn3Xz+8WNztrQ20g+SlxxPjLH1/GuUZtQ+YPFnfwc34abatQOR7Ty6NQQPtON4sHPg7DzUq
OT/9WT3fcGf+46ZPZXKldFzOZvfPS+bb/NnxmlGO2MOlqlOT8NPh2n5o0DKYA15nw4bpeVh2SniQ
fkN49Q4ALmalkmDVmKKJq+pNDK5n1GyNDg714Hi+CnzSkZwzNtNWR9uM59gjF1TSqczzTdoammEV
NJ3O1JOxo0+lZJu78fV6YdZz0c8lV8NJF5xHJDZtvZYD2uBxSMwCv6GnIWn0eZr5zkyvAyvr7dJR
RRzJ3h9RxmVdV7T7jyXjaAgxWAxVerznsKQVyh8SSFwfUQ3kLDeCLUtPO7EaT3al6ASJwSpQj9wA
nyRarPUjCJ/uIJfJUM0+bT+Xo9xfs18OfZkIpRLCZNxof4rBKgbupn1j0+3A0NumySS0uKo7HG0y
tIXMSF9ZGfiyyBWeET6McU17Ujv7QVS3173jXSjsE9kzZT2bc/xcED1r/ZSvbwe+hLxJLqHHtjZp
29ljQLkzbfIhYX6TGcDH6MnxjMjKPa7Wbm4uoCm/iluKYgJqyghcsVEJm1qYNaHVrx2u4DSxFLK+
IOcoaKfVbXit4pH7K9d338AB4r6usyK4oJgAuF43ziyCQXflCwDGow1MBnVuxn/HMsdaTgiGelpG
kES+hCa+mJy0rFRsZzkeMjU6QBiWOikf7tgoe6ukKS5u+Qckv8aYcBb8cyhfKvRZ54P2uGN73IWe
LCyO4WymcVTFzrc0MfIMzBEKZOl/s8O7dLgbLO0IqzXm3QVDEps+kjBizP9SHTKF4fxxXctyLHg7
MsKrbLp1hCK19rEWSrtNhV4g/MvggJqq/M4XMlzbasYZgxhk9Hw+VwN2FVcjlyAP3ydJt7LcOxVq
USIokf94UD6lfrHnOgNhc8ULJ+XfwqbY1Uj4M1ziYAEQHEdifPhNJV1zZF+eZNZ1IjxMKSKcgm5m
J/5vOZnL7NqiYt8cH3s6jeRUMdqRcDSWe728k9rRyqDuYCkMpWRjfmTyS7ydQapLMBLGOvUjuG0q
wNZQXFI55mGo+ijnh1GsSL6rqPNp6kzs8XZFyt1ZpAdviDYbyggtR/0uQfFnO1qcInTvGBBj7san
HsG6JfVLqklN7C36N/t6X99YPxCKSzXia3AoMW9hE53vPN9L1bZ4B4Wq5QCLi7j0ItjyNCNLr98r
lEgLyfFRB03V7fhn9+CbsCN1FEzzhO+d+4K5+792dcvcfc2G3hTcY22yd2jzV1G93JNitgW8oPbH
XpEaXdTnRluYLpwae+PUnF48giiuC4j3/KUE7kcOu0xNM+PIjGeYXj94hRVhAKYiTIWikQDXF748
Kpby27vlBIl/SLUhmbsB+Cnh3onNBcHPt04GvcAmt9CBIJES74hRjfRGZTjbhSY1fG4ariFtksLR
/GsAGxg2VDilpj5q00NNqqMJlmNeWp2bh/tgvtnGuDcDd52E0WQot41FzzgeOcft4wMABQDfTK+V
Yj9S/gRsKmWoSK1s0JRKu63u/zSRMM149pnmXCV3mmlMz+k88lkuKlmguZgQrb+VDvIbbNUrpnvZ
x/sGEbAdfMDfH1Pd2fgHC29DZvmM1Wzi6EmxuuX4b6u42En6gnPgeNUGnfU7z2OvqWKFOjSfdEA9
oDYoDBU8K8Msb/XwmQWRRxEU0ieH9x3GPRCtBlgxNU7peChJM8J3hiJP7N1gchEX776Q/nYRBhys
bcCSUWHC9vobEIVq5qumRBBS+2Au6SUBVn/mTJLX2lWLqXd/z1RbwnYWs1DXdauhOMP5gWgIAN22
J4+giaUKP9RZzU9znrqYVfkQiseHrhw+fUOEl+Qg2iQX3+MM9DB3G8Gr0OJnpjtrMy1VMx7Tt6lw
pBA6j4ue1oCESlFXanoUSNE0JxGJBwu/LU60oQwYGy8u7peu/XegAmNZRZszSKNKU0xAtAZ9K9As
6HbtImh6nN35+Gzw6ONej2C2oYo/RY8FJkmlZgBZU6celpUJqsedC89eYYn5jeglHqjipavoVibj
VL85OjYqp9En3VqHnafQbMfF0vx+eV5b2fKYLXlUnbcPXo2VY7ETpT7SGOBac0kCuklBh8JiRjXR
t/5gqLd9NrmkjFiI0XEjUEczZI+2K/8o2edjggstCi42KQbjUl8VD6GbdIAfV57z4IlI4VmUTWdx
Fv/othhFqzXv722L1M3vw31wTei4UkB+8kkAIwxxDTJLQGSMwy2dLxsA7z43tB1SqCmLpRbvsCxT
yx+kya1e8ucf9DXS5wGiTWs8syaox96O2OwT2F/YwOKmQgo7KBWQEhiL+eZFG+TYLH2MIDt8SoWe
hhV/xuVGXE/numhPeJbQUSddxBm5KWfMXylfbirBZvJAIC18lcXKNvxwYHEIDXKtYhXrZFgpIsvu
OF79eWj7FR0qmM/O57RmEZFYDB4zehSh/6WRLNnGMlF/A3VK7QYRS5XaBFtMjvJrqqk/ZT+f4b5m
3UaYl7HSE69fPVFiMg2NQkLY9dq7k0qHOTsFGCqThyouHOgDk6eGo22brMwqAN3qv+C+szY+Z904
q1xxroLvcMqCS7jmWEWV8nDhbp8AhbXekzP5g6EKsba0RBqK8t49laU29fYZpKmWjpvqgvpa1H4/
EVWwF+0y0sjIsflMarsvuY3tKNVu6kvAShe59EmJtCZjTCjSJ+i7u5bz3GueGI/jtVWRi71e0VqZ
G63kkQGgJ6e8BzR1NHJCCt//3kn/xlI2JAtqO58d7R7bJz4+v6d5wGgp1a9hPq0QY8ZJi4VVEM+x
K0wthuMon8u6tl3pHZlolcS3SUUKE/+DWn8/pO5/WJ42ZMml5BZcoQGAwPAgV6XKeoO8N7JPW7Qi
7PxTP2OlDmszvOJwRAxCnC3VlAdy0MF5R9J/xaRR3MOn0Q9rmkD40nokOyEn46+TKY3rfRpRI4tD
Ek2eh7RShsZowemJrld317PiPO7LCNenV251AQsbxG+3tbsnDUU3ZKOPGp5pfn4okKgcXL6mg3h8
c50WmloFpjqDLF8EwDllZCzysAPxS28BChQTQkzwSW2STcWasjceUeFzHoI3XU9s/BZl71fGl3eu
BvThsOJYnA3cggoez9QjV9maPF8YYB0BXIS23wAvbBOaJQYMQ4gzpNeFn545HKgoGZy+53EwvmVP
EqJdIYw7W/PqPeEl74FVKh7rNodqWtsuTtSuqFw5RioSw/q5dC7T6OUTFzGEKstYZkmWyBGGq4Me
urV4Ipk4yjGCbSFeo5JmLc4tjODvlBy9ZE7EUsb9XrxmWFIvxGQDBj8tL4zbg3SKhPN8OANywHuR
WJ3dtGKVFHhXm0uY1sHW83v64YdY2iiOJaCOjpurg/hvmTKuDfElWo8Wp4RXMmmUbHTifJsbVuOS
FVbKZsg1IdZxEZSeBnJVEU2Z/4yC0iEBQscr8K8T2A24sJDP59j43AOkgYXobwbW1/9y3KcWqE9p
5xV8/8ewLfFuj4ejl0jGBnvpEYlG8i3pbMKdx9JwqUJ2x4PDv3N5jPTln420daqfwYzDiv9fEe+P
hetF1nBdKr5Yzue4CYXRsuPki4JDO7v34kb9wHwFeKGBidvDB+sfJpHG5XBMs8WVXFxri3W01TIL
yCdTxCaGrlgmxNSipDKyxfVQMMg5UF91djOoNuVbeCXVxmAmWGyJum549Db8nPCNOXT2W/1dHUNR
pu3WpTJYlriDxayXbmnIOMSnsl6t9A5wCC3yegWNKcDF39jxku6InnVjiZzMluntzEoeTOgzbhAw
FLXLjEErdoXdeC9oAmCtmPxGhI6TRM7pmqlDRbdkAumc1FdUKLKKkKL3NoMDwn+GdNj1nXxwy+ET
hJGT+S5tZ1sWq0LYDJod+lSZWcxmLw37MPN+DSHpgx5NDF7SMrHR6M5IrjaXHu/gDCIfLyWVVf8m
dmqA9QfDaU4MXoNADKZjf3RcPVYLnro17wytcLSK91cYMOhJBsgyP6jVhWluhzLzM0Grs0yrKmNb
QV9I6xEh1DzpWSqLmPafujvSusbwtHx8jdjZXwLO3exCSlutNZKlUN5WpD7BwuCep5/Zv49R1EmR
4I0BG2pBVxSg1tcIOx0JX1NR5q3nbFXiEqN8omuupzdCJa69sHcxkEVslhxR7O+cOF8O4FhEWP8N
gLxhDXlXUMNp3J1F5gZwAfXdMqjBXP/yM//TBdStYhKNoQhwEWQZMatfYhzsVbfB0IcbpVXshaWG
9V/vmoGP7QCz+BUksZXUdA/dGZ77naicrn6DvssDFpNj+WchXMF4C8DYOD1iobr7S1qYGM++KRDP
/f2Ma6RIgh4iUKI6KBYinS1LsZKAI4VEzMcENkdDTf5jJTOCLs1IoiqKgzVNh4jAIpRTPQ0QwnYA
fsBpW4qBvJWaWazznwrlqWEBKClicBrjITJY43z1I6QJo6WM8LkYoPoMe4X/j0Dxv9FtCK0RisDa
kNqCqM3LWBrntww+KoWHV85NPC+gxLbwx0+BdabZq2LLQDYlwAT0RKAavqxXcoJ0ujyZBwW3btIl
NUzQdx1kSj2u/S1Oa7jKFkHWDn/i70adXFABi4whvhRPlQy1Srb/AW5BvR4Q1kWXs4AdQRMT3v7Q
h+gxMHOUCAUhMRJT5ejhgPa3B+xxVw+4HPmnXpbZogZPCFhpqeaTiyO5BJYr2rNPz3d8f7WJD6nW
P7YQzyLsnEWjBYPrH+ehyUqr9VtD1g+7NV6guF7uqS1H4PBYI2OyQPZlT1ddibc6fxHoBzyYtn6j
niPD/G1Qs8WwAOvpET5IT1XAFnLtC+59FTSbfsV1Q2B97IJlVQYXJEgtMRTrPZd6uKdgjS1gJpOy
HCa1y+HjfNO+1HrwUbyKrCV5Z7hCsEbptqHRTsO3o/hHCBwuqgmCEJQBZ2XUMCHLWUjFTddwGy1n
x0Swu3PVh5gXWn01Q8Ak/rbANv718yhSvjxg4js9DnzoetJBQ1Ldrkv5gSA3ya2FCx0pBlj1uXOS
J6Njd1+FCKw4F4LclFamMfD23hz9Fq1m/T/zIUo9+8tkDSlFs38kiVSG+Hj7jUV2ldIAtwua1UAX
LziumRPOs/wQbAPslnDcStM1hxBCZyyyJUrVvqKRezl/LOAHEknSOlnLu7IfoCPXMCV32TrlZYH9
BoZRRnHlwI1hRZaPvQpU5Njy1ZSKX/r1W23L4k2iH7askX66cOelSa5Eqszzql4e+fSyLbN0bqcn
Ssu1rYl7y3u2poRLlhgoka6kNN2uTEDJLN2gxrhk4AInPZz7YB3cLUVEu/mmYLW78GzPBmzlFmOw
OFLmG8/P0RTweQxKL/gWEiWfHzwmFw+hm01lo/mjPfHf4tryERNCCpaCndjBDb09YoRhhTlzlaxv
VDnJtLYD+UE/FYO+EpCZzdgGL40kMjAaZ1r6vfYHT+A8Ksh3DkRquM4pWfYzqqVtFSPKHjua1ooq
UW10I1LqwJ0yb2vzLu41dAXahrUf8gznYcpW4t7O/fyLv9NHdjbrQXspOLkK+ZT8BT8yU5SRhmUT
b2lFHxgPkPMZFVXxDEpOlr8roBLB8/X8NZx+OnUL7VGTkM+VzMMURnGHy2DlIByD9YOApZ9803ye
INJw851VSTj+iAiULfF0+tf1Z5jTbx1YhSmOayMT/5aeTxWb4R/6URfUlQBMNQT8bjnKL9u4sIxN
4oSK7035VXrmfM3iC9t4BfIOTAKmxnGY1aqU5qR2aSVhQt1eni3KZAKwhZGLf6/VvM5O9aQ40ngj
G/VSyEIi8Tt/mnCA/dIgYCY+dsT4C7HS4R2OCT/gDgs+TxWu+dvunbMEtn79y4sK+m7MToGqW6IP
5Wz3jnWPamoRXxXQvQV5LKW8EyKBvWP6YlUlCXk1oGvd04AQIfnxsvGF+E8+6iuiQxQ9FsHq293Z
eljFG2egCNe3XofoaeTw54zGDFwsCl7/gIed09/jbgnZoS6ixss+QMuQNSRHP64RJTydeq7r0Ovc
AoymnJBH6LBEItA7LK2zvw4XqsdFIOGPJskIyW1AFJuGd6s6Jqht4OITjpGEpGmYM1fI2sbBd3UJ
1Oo1hS1PegmEMSKaYtIT0/wjw7Njy7mi8H7PlAYRFcQUHHMygAPcOhOD8O2LAlBa0zRxUweB4p4n
gYGq4EWRoHLwMV+d3Nb2YBAmVtezH/zP3Vqa1OCzubfAnAmYzSkmgxTSiOf+XwSmEZ31RMRWBONH
MXQscevyniRP1dNEKWO5uoCKZ3zoSO6ZtLTbkhw3ucXi3MHHhtCi8X4jz9hiKpLKrYjizR+W+tvd
bmtSv/5CblloqYqI6cEnJGIjUw7T1raRTumvF7VLy3CRL6EiH5uj2GMNSb8yCG3Yu35B4ZzZBC3/
Z/MPerCYRl9cbDqwI7BFBwuKUnhZe7Amf0uu6T4u+WBi1Hry3FpOtDBxM2j7JkAixl0myFWLunWp
ntl30Asmxbq+BumipnhNx/HNDcnOUsfqStG0K2gJwSOeidM0RQsyj9xXK4kKE40C4+klzOulIv2K
9aEzTon0ogNQkqS1iLGDm7dS+ffOTe5a7HAJW+kEWFM/yzXGR1fZajDxop7uKOEpWAV6DvxUa/Af
Kw5LXn3rYrscHTSyO8S4zXsPI9Vf8lNcPsbhGrRtR3x67JzaUG0qlBr5maHTTKEjdpdM4tnhS+Nk
RHtNggUim2gnslV4Le9kSgzxbIhkgUjY20O7ngd0grAz7kmUONojUZhNBHFlEz+X+kocK059vrKM
qICLjZOADf9NasS4XzKaZDj4RxozgcbkctQ7XOVMLLgR+JRpB3Kpto/g1bYcjuURU4BWLatQW3fl
su38/bajHk9jjcOyx59J1m5R9UUP79BN7TTrBps1R3gAvtvg//sdx6xyEMFDKuf98GIHElDdLDTf
4QRgPbb61vQzz/1Xozz7F/7eG5lzs9f08VOmVTV0O/0mv2wlsIgYBXrbixIIdGqTdO5Q62OjGaLc
dFx/GJP5bwshxchQpWSZhQ+SSI9i1RcZDJBobmL/0MftTmgu8h/p4M8po8nSmGGGy2BYB+9s6CJb
McZCmY3QYfgvPQrxhE2Jm4QABkVOkOz93sTRNLe22TJdIMJ99/d5K2P6vsqytBsQMN+vJce/D39f
oqmsVq8yml+/pMOnWd1qWRYTwDKnxFxCXyWy9SGmzOGBqFMV/u29+h0IFkaE1er/m8CbpLtUjGnD
wA7aknx9Su4gwMpIH3Q1p7GAXK7QrydnUckR7jY932myk6/alAIJ4sSygt7gusObJQqyFUqHfXWM
BPRcsGZdC6xz/EieDZ/+rFt0wv2iL4O63Rt1X7Czbvqzzhn80IWE3k4f2PL9Sf5M//D95fef1sJF
Jvk0N7KTvsGf5Vj3TtRnvObbIE1Oxb5JcIl8eKNZIvNyHPzyAoCnEsmXH5XN2lgi4av9B5cPBvwe
eoCtolsIhHer5rvnBbHrjquKmVrktlZ58CFBQIr6+MiaLNggiLvBK1gsT9V2dYeKNUyIyHuIL296
rge8M3fHBpGtKCM5kPSQm/1JO8PCJ9YVvrRvuAf4JBUcvUSjsI+colhDMzYIWuqATTPx56/j6ajE
fpcppZpDt9dy+mAwiwQukEESJz2sZ6D4GfFX4b9mOxasEFGNgifKN8AQkDmVgFg5aAVVMdKSt/0J
/SCuVedutod+sb5IZPHbN1LuEwvQMfJAIJJYt0zbGQ3ZFdsoINY+QdZ3liiMjiZg/QcVr6ieMSQR
xGoj9GKttt5WOiUaFIqPW977k2LgrkBe/j/i+KxKodIsubUgt0ukfTqXEf6u0y6US2NF3qogit2a
7b10Uxh+pfug4X+0TGTNiQ0o2Q+upe+IHrzahuudlfJrGkS1r1bBFpzqnRzsFS8SfZi+bCxin4fB
cNqIbxHaL9gqBCk9yeaow4PCmpjeY8nN2B9DDVgHj4nEOgPpCtp1S8ikZecVfVRr54tgVw0LQZT2
6Am673MjFuNLGVvDUK+GIq6plRQchESi0Xnj0tz6bYGy6GIPDKMvOYzaHE9OwN8s5zqR09U3SEnK
0GFgIg0XmXhmfJVWWiAkZgN2G7PwMZqvNYfacgkZO4Pj4V9hPyWX7WqP7sTWid6P+GdEto66fr9b
4cxCo/k0+1Wz80A03UiBIsg0bvnaLIYEAn1pzIIQBAR70ubpDViyejBF0jHuLvqHvUaNO+gWzoeN
NHguGYq7+9K1dKvxxf011zqwfAa6FBFIT47EYnpb6E/3AEuzcv6UFISWszwPNFs2gwMuG9eEoSXf
3ccnyqg2v9KFgHgduSb0fwq/SsX+zX3FK8F0dNVOg9wLXYxYXNtcXMNcJzP/Ll0q9vr+PVCuZt1E
qhZuNeCx0DrPFiK+HA0VDrYHZ18HBex1GjtIaS9KP7fv7W96X7Kcr467LgQGExZySUbQ0kOcwj/Q
L7ObTbC8WxJEBZiDkVqB955i4W8BP1W/y899W9UqN3flaX60WPVH+X/TLwxxzM1iN13EKbhMxGEP
Kno5TcXo0r4ds3Q/81s05XOKZVgt0CYIW0Pw+iXXvU5wlINpaUvNEwUKoeFLQr6tjpwESOpHMwn7
ZMBfdrmhDdbqUKmTh0rj2ARc5mYdLU1KRAoo2rY47I6E3pwlB2Mw7C7KkCXKfHIDs6Dl8f8WG1pa
DGUN0zKmiHj+9RUchTdJtdes9qRYwgaP3kXXJdTT4lWF73Q/+hhh8yvQ68eTQEwFvG5Z9jMn4Xa7
VheaFJFEP9li1MKNrQwXJWTJEn7uagYLckytUo4FFIy9z0o5qgVXoKkmdCqtTZs2hX9wO55/7ODn
pqddwW0M4L8ffG7iEDBmHg2V7GaYuHJFL/DODLPswH7yzo6s8jYHjEuFLEOPSRIAAvit+UrElWlD
3PTy1nAwy0gywIjR1N29Nv85F/bacsEUfBRlc42HVC/NGvQC5iZZq8RtG5Ty8OZP+gSuK5NYDN/6
B4fmh38KwyRO4IohtiNgqfdVpyXY3jfJJVfBGkR+b0IgBP/96c7XCsTYWT2sBUGAeTli6E1UYR/j
76yA445yHpmu6tGvAvPR9cc6izLmCfCPPzF8YYHsTLTUskyOP7xvR8PUrswTOw+EQh5VcuXMy83g
cF+Q/Tl05n0KxqtUcI2nvcpieNYvonQCKLbubtc6TpcYKZTN7HNkka2xHGkkOmCgiRZuWJ2Pke9j
PoI7IAED29BFgJHAUtboRzRCUAv2S8SyNKV6tkmshknzh1HLfzsaiCRoxtOm5G5K6wai9P+p5K/Z
zCqB3UHy0fujtaxHphgtxUMDzZWcaa1X7FdyN43HQAro0zqd/ie6+Kce3WhAtMb96/aXifQo4A4b
Pk+IpbErEbrx2fz4XC5ien1dMo479RoiFVMqRCwooL3clW9pxQgiy0zECCt3HM4ZNTtt/k+AsVBh
3Jwbw4jA/1L2PFnfVpo+A5Pw5a28E5lUHQzdXyxWdoQRYwXYBqRqmq0X3ChhTIO0Nm9gNUE9tznh
JhzITKNjPcgnjN1kkv+FuurtaIrFdD/Ji296RBUalMwa9SnorKSB+X+98TOveRX6p6eT95jo6b8W
sviawmyeuGT77QeYukoUUeXY7ynbS2Z/+9vYsVA+0qj1dmBC9Npx03wiCcr99Ebd3LeT+cMh4/6f
XLRhI8mOcBmcHU27ycuCcoZThygkDqOSGtPq0/E/lRiEEQvFPLRP4chhFXxmRzZkLfeSP+Ic6ysT
bOlxK92AFtsKdAFCHCvDZ0AXrG5lcIAeJnpwcH5wSb31tVlwb+Ziwlq0PmokWys6viZJls6JwqUF
+lsugyqCUexOuY8j5YrTRztDgrS1g9kT9JpsjwcbmHReLxLpmggf9lWLYgJuKkqIrggVy+Bx+j3S
q0fmjxFwWkh9XXWNxjQ5OLAswPVZa6cibowKi8l94J7kTgnzv6UFtbf8NxfTN2+vuiYZS/OTE9Jb
0ZyFzXS4rr4ab5BFDmvwIj3jssCWadbWuEeRmgyH0d19qHx10af0i3TMvEVGzB30cyEf69qmRbXo
l2RteH55WmI7VES01rG0YFkqgIJQ+X6y5A8O5X4s5gN+P8ydVh+tTUhtu+38EmNMqrN2GTXHOI0h
ZPKHYFT6PBMxLdMAyLef7qJHfMMOgfS4tm5Rz68uipBo13Jy/TKQXa5mqvSX/dZQigF5AEJt/g/K
otMpxb4v8wi4lrFq1HTZLke6sCcMCZ/2AjTr+u1ySpObHKjmbbIV8qA4NwOAPhGNNDey0KMxfQyU
LlQMOzoWSAGcGz2l0SAg95tjTOrzl8IvzKNmHg05M0XibdyFRhMY5DqttL4X2FEDypWkKp9McN50
xiymNU9Pixk874OrrQ7YBw4/SmO2hp0Y/ALfTvYcAun//ixhNgn8jxLfhKkhx9xk4XJFgT6k2xON
000cPIagtrpBAvsO25SbbF/9/ucZVexiui47jDJGBILhjYTU+r2f96B3XHVkyXRq32qOQbCnGqSG
EtjsIEyjLMV0q//IeORff+d5OIM9oq2bT8krDqQ0aNHGosxqNwVVWeOpIr7fUs5GtDBqAcqNavjz
gAV429jpTRQCSH75AtrF1dXEmRZnF6D3exIho4PgbNYEUvq2r94ole5ymqoIDryvV8boQvOukeVZ
iUWDVTJ+1NbkwFFcZhLjQEnNoNZ8BZg/ZMY8A5H1+i5BCwsbas6zBOl7gh5o2yxwMnzVs3EwAMyT
W2AhopFt6bPPY3Tgd1jU0MEfUwlYjIlkMyvYzMToCWu3AGG307nqkO91lTxwxenuh1JTndxirpjM
XB/Oo/Lw9tGy7hqg6/JUsodZnLKod8oNnxTIoSYQbppkZ3oBJjOMwQhdJJaVBOAFhMU91ofq7I+N
+sT+ob5CkxBNYZjEa6AZylD+jwkYPgTXmg7KEvipQ3WIA9EbQl3z/nURTEBUhDDjR+06bVrGsu5A
uezZjoxNr4G9j8TWoLGl0gVpE7BvG5oTxfQksch343AT190jU2Cmu7hHu0H0zDnho3Fcty+dqRbo
1a72iY/u0EM5rukZj1ZFMDBt+xzIPlgb9FFB9fUsjFs8rsFGnIOef3JODqijW0io8VK6PXc64bpB
eqpLWnkBewDAOCphsWEsA8/2eDAn98Irn6LwxbH0pGxYaV3hp1wH+NcPLc2onYGcRTnhxAp/yE9a
c2qJJpoTM6/4NUYdEYcIvFNVqOItp5grkcMNrYYxIXZoUYP7qJBmjaLxVCCmtDA/kWkJU6smIh76
ovy8tVi65OpM9M7XoBj6B3B70lKl31VZ9Kr9jLalYGVPUxQNZ+AltapZg5qSf7NXJaqDPeYuwkiW
fSfjIT5CbbVX9Ji19NVQTHsF8GB6PZautbNl/v6aHlHyRSWRMssafkDSeKuzuVbIqM9aDPvRVqNd
ZHssfc6eIJOTqMwk8KwkFXUIOzgmo1xrh58ycn0bvLGDG8Pjfd/IY07iG4FHQCXcAsLVP7uLsB8i
to79bFhUu5bv8GrxC6VqmO/yWYBRutVoG0OPrV84EETA6wQzA9DAx/fq52QcKbRU5J0OD+g7ko9w
KNtSOs7UqiLaOvYyGnk4u8ETDxmtwM9Qwj/whk+kMpU4oAtXMIY8KRxPkTEn/7Piyg1UVvC436XD
RwZxI25oSEufCorQiJPjBqqxH97lmPwC5Ce6sZuWEnwX9CSAx2VmVnVD54PwBs898dPerl0DAfmp
XumDLv44jTJOQtT/pSAGQTA09Zx430Vc33Z8yReb+sJnrMPTxOS6tgmZan94zpIdmw24XANZhR5K
A20880Smoubfn3OfHLezhia3F0QHfDCrQQOzrknJhts1TY5sL7qv4d1wh9Gob/Iy2lWheAfiQ3T5
nhZFsz73pUqnJBPIjwkXfbVcBQ0G29H5AyNgnYVvQ923Fc4lHgqZwkurFZ2DPr6l7kOo5jLQsFjC
Z2HexrrhEDbJhZGXhhXJNZGEPRj7qt7VGCqzgAZrfYxgrMDElpzqzHHIDMr0aar0GpCqnSQxXmEM
hla/1M51LVExABr5EB84+aNvsxjmEBdQsDeOvtzz/7zxr9pq6DOa5XQwABG48KQlmsm2Xc9MKR83
6tApKOpOYdHebuZhnyQkb26d9ECldaHRg61RlSwoDEQMWS+YuHjAlrzVTJJFIUvmPeBYYWqHvLHs
ZZsdayOcq4ilHRPg82XOistUP2Xz29E031996DNrtLUrQCukRKSzcSi79EPT5TagcyOqvHTbjNml
FRrcI1MrkopmjNavElRGzpEE0KofW0jDAXKFh2NQ7K8UIkh7Zbu3TjzFqXxcfOKPDksSAerf+8C9
PN5b3DVkdUdVvA6V/8AmSjYLGCH5S2t4Fv9fnNAFkCVFjR5EnVxhThyZpwGmRt+QmPMr/XqZyFOd
0jc2ZLRBSMhYINYum8mnDFYeva9mq+XxkVnWIxE1unwn2OEPpp1TMLCv/9k2yz5rsqcGOUkKmneB
93wPhcK0bXSH5+RhjGSV5WgiltnEYh6gNY/lAipmQ7eRrl240h4z+MjIjrBx6+ZC6o78xicg0XA7
dALAsr25MewPgzDwwty0bau4I6WvunyeJs3KT95meIShrDHTPzdgaPKYZ4V8ol0qlkwX18gLC/Pk
51WHb+dIh1+YDU2l0fiC3iLFlya2HYqVWR9QyGby9DaIkrFsueuLPt2jTI+DmErRTKU2GpjWkQ3H
7EEp7DCse6ojZcE+BvRiuckDxC/rS5pokX5dYCqwLQZvTjvVjAlwXO6RpPBeW4xtH+i9PDPLppol
QkZp0/QKu9Edqudu6yRgdDEZwtCF53ZW2f2pDUf+HjvknGw0Wp4h8crpJAcVZsf4y2IZIjUQfkgF
fna6AYuUC+j2UdcdbOxMwSHXafJfMdF7ZinrKM1+sqY/HViSS8qcX6KJiE1Ye/V+f6ViCv+lrAPh
tbWexWX8ORxP67aZU5ZPq041OX6GPFMt9Np5fA1YM6qSb900ZS2flHWInWgTxfiJuz3A8CS6v2yt
TNxQXpFDHiuT9UBFYjm771Fw3HnNziwcmVoJ5phihlU6BmST9tQDHN9RenSyTHu584Dx1Gg1OCVq
rGl8OQbZ3cpHKjEjjBb5qxOASRaeYKsGjTIRbbfK6H9W1H17flgBRKPJ9J6SQ8aFG2c8z9G8/PC6
EMUuaDv0sKeTKegfUUAS7eE+y4vbPH0oXxmIVaebCILB9mu3sIrmSV6ektPqmGm2X/B5zgljcbX5
rWIEZ6W/W7e0RCWms/VRaRk0slUGN4UpV1X2GaWixClhy9+oNamAa3S7I2XMuolwb0Uc9mfixsVe
0IfZxliXLscAs3/624Tcu9nn7rYGL9HAghXnCz3yPeq+IhRvk5ZcK3CcQWCRrMs0uusFf1b3FEU6
UYVmBMu6gt1ZRPeOujLTM5fcFNsN2tl0sC6V4/R0sXhViEpH/FOaYQOe/o4lvMygWdDJZJruJUPl
CuLky3YZUf5ZsQmfn8vY7PqV53O48Y+45z471WN+wcAXqQVO12RlkNk05cqiwXN1ZM9mbLXh6bLG
FxW8rn1AauPLMy17C08MipQuc5f2Nwbh5cHt0fS/hT+VgCrRtIQmoSCzKdanS8MP03Z/qg6YvobE
6GF2i4Ik9jZXxqbpir26IJoQs1gsd5kPPcpmhvx8TGnjU/0lAFxFbWcwtcGHb2YOEICSSYnlVDLO
c5J6drY7ZUeb/kMgtR6VJqtUeDxR4QYXn9tIc7HRDx8kAJqcyWMFzS7PSMFT7BshgvdCKzl34u2T
c8U61DqF68klEd2uoN8m0ZqsL2kwB/hnbDFNoKyfEj+t/ZHtcAY0/lEbQNw2qafNzFxt2nYE1DWR
nIlUFLkD3Guy8mwZBqeu/MTU3pYdKKnS4n1+A12dnb3KQEMqu0xVZehwkJMZC64M3ow53xb74yGL
2lCJCERTIz8MCAGwBeHmYY1az1KbqMesgZzMCeGO0kS75JlrasviCk82Gc053PzwMb2Nup/qJ7Yr
7Cj4EdtJeqqw+rbdS81XWVPThNQYi1T+wUv/AgGMsynLCS8XRdEM8gotae1exSxMmLUz5lmgEBsZ
yfLXYqxv9aL6zMvPHR4uC9Ky59bdRc7EOAZ4qagIHPJs6oKfpYk0o6NalxPqxZDwDnZ2uI1NMbjD
LGylQUa7wBFOFPTiqlF3a8XMgmoKQuWHXGpCLFxfIknyJDQS9vf2AV2Q7qUhoHr/B1b5HgKvp7GS
Sll8P9iPhu02SIkqQKj6dQYpcBsMyB3vzzosViTY4XDY4WTwAwxEu/kGawVFkSoabT2Rb/llnPG4
Y46dgsA3I+CArid8H4a5kacLNUKZ93ysLAjHQnCbBdYyrE9HMTcW5n8Dwqa91ibZjUcUoDicrNw9
Sfv97lMRooKkeCC0LWUXIcGAjN73xo9RrlVW9tvU9JiD2BSfoJqqvpvGSSUETg93iVA7N3cv2jFh
dNbwJykT0kzSgb2O7jt/rMwiS+sjLfdzaIGYl9ewyw45A+CiMh+jpajft9VKfcrbKhsl1O6NyMWV
kG+3kHu0J+oYPzPROjn51zXNtDoWaJ+eIZoWhsV3kBaSfNt8tupebzvzWXKSqLoPRMHFo1npib/4
+4Rd4pC88Ue1xIBWWh00+d0tHoxm2OuChPysoivjO4wG3YK8/2A2g0qB2N4y5fr+vDbhxRsTOF4R
eHd98gZhJa2W1AktVkB/oQ5ExleJyLniEuxuOwhA7LCv+s+rCGVKYGAwy6EOUk/ORbd9PTXjrtqg
+ckZwmqg7FQKz13fKiz6fJft8nBdJ6IAWAJkwJTgzXgsIygmu+SAuqI55jHx9rlDiUhsokgwDCPE
lXMLVFZyPjB51a5btYvqKcpLA9sCQORScvwhxcmtbb8OWXtKEH7nngBjN4lUEeVRw8aM27nWPdGe
jy1VCoBFCkQRC90kQ7AeTkNbyoJKnfMlMWSzpAa31jd5APBKemo0LGRsAv5sQGasUNdxMZwwZ/GT
DSt8cJemsaVT1MED6E7CYM1wPM2ERWWkwNfFN7jlvGSdYo3l1TmdtnQGoElcYLt+NYRbKDZerzjC
oJm0PO+jvZ3GMD/yIXlqRNzyikxNoz51ZXvdkqT+wDcUwm6UT3TRO+y3orX6NdHkbQuj3aOrNILt
Wd6oOCrCu+g4QHsgJOUpXzo2EWyWvhJiY5GAFg+8dMLaT7ORmygnFAUP2w5DB33YADqq2++fyAGQ
JIaD/aiTgqpbsGqcv6UNlCDgzuoWKlmCveJK75mCEDHszZXXYK9TFGcOtMhVR0XYNGnJYhlZl4oy
h1Un3IoRMcyjXQC/qUPDC+FFwUWvNIFrfCpUeYdjoo5r2PYJGFm4e5KhJX6gDGfZrwiTIDmuKnY7
Bhk3z0KCl+opt/Wq1gfaxnMBuG16QYStorAAse2YybPFb/bxGnLQl06oBpoAPBU/S2LtW0PItCjb
XSue7mn7nVkmc5Igg9JEWHKZVwI/HPqebf+qNrVv+4+1kIAP/rcJwwl1qlGjpKuHC+KYPWN3Go2c
v42xDI86puRc6lk9yBC6QKAQjOliBp8aSgqwmZxAktoYcb8dPCRiHzA3L0+i1YYHTfvrj9LbBVxE
+pA/8ufzO0LAlyrXAF2kXz6gGKA7P8OZa36Cn2cY9B2BOs989nk9uCKOjm/+/uWq8iS5yAhKlX2b
sVICyBiqMNj4UQsIdq/loXa6UD1g+hfoVRpxkO2oc3sUzhPYk/RK85S4sckIZ74kETV3s7uFRLoe
u5qhaxZbb1n3XLoariFK9mnysoazGa8c5WLzpla/RjeYlOqJn3ICYqYmel96ptHEkNfcG2be8Kvm
LX1oW0yZ42QvUpbR/F7Z69s/U0ovcuTLD17hKLpyF5FIk0NOs3ELaG11Qk0Vaa28AFWCEcCWkQNq
z33r8XRn5DQtdGG+7q83lcmFPF8PNrngP+B+4U7IdFMwVxMcn8Gkb+ldkY7rgpHf7tZefcw0iKmQ
mN4N8xzFaGo5DVpUl5G3U2ybkmmmgdqk2jFuvUt1dXgUltcH9AFy5KyqwhsN3k1GZRpXMjUqwwvQ
AypxT3X4C/ECk88I2J252yw2qdc5KGZ/HkwIwAxhMQXYfVtfEzOlnMdW7YOKpYOiADIkXsn6hM/F
buEGuelLWfqNarP4jl8rqHxuYNj2GwOOAOWBuSQBWto+733Me7FjNGSHdx1D5T39zMwbW5eGafV6
kgA2jJ+AZHYibnBm4vF4Uoa4T3Ny/1/MDcR9V026ZdQcWTua3D33lSeqIczNhILE7wEKaYQIGm9M
+V0sLXNjVD7iF/1S60xUYw30kPIKWxzD5ODDn7nGiPA1Ny8KIo7Xvq338OSCPH6hEj7WHovnRnDG
SGOFjS3eS2b0H3VGLcJ6tkT/YrBGowtBmITn9vyALkcCUsBpN/UYDkA+9NPLkBnIOqx/7WPrGpcg
llvUTsYc2pFdPnSLdovwnGfWodWfORg6BP0XjUpwrDMhMoUqPwKg2+SebZ8EYUQsjrjpr4hWirWg
AmwQJ7sBDJwWA2sqQR6ilAjqD6ARuJ7o3/UQ/N7HcV5NZ322WUiSVshQa7nMIYeyn4/aL3xLJyuX
bZn93SrGNbJ2qJfLE5RlLLYVSsDwMCiGQMhXurIgrA/UUuMTPBWy8zIptZi9NMkcH4EqI8QK/11W
GLcf5tDs6F1OTbOvu4oV8te+nEp99bKrmhcZQpld/KBXHFNE5Z9FWwT+Ys91XjDnGiTAMoXpONDo
9DnhLfZYj968gcVJDxElRXbzjonUu2qtaQkFlIIskjtGWdn5ih2HF/f1MY4h8tOxuZcgmMmjgfnR
eWOsrTMPT4hPPA6+MqUJR2FaTcEC1WwsiFU7A8lSbXw2Mnd7VuoPa9DDPsgzYelKg5+ZtBA5nRC1
XL8RGjNn+ze3hNPjDFhX8Z0XNS7Ecv45gLXTlpqf7gdU8Lr/K7WeeG1FQx2+e8Ps0B6D2POgiG4t
9LfSCXlxK5SZvGjxfp/AEECWJ84900OsNc8O9gtBH4JiKbpiGTl8VEg7taBEIAusHgqZzij4W4ZM
qLK/WDvAGOQUeFrah8hR4/iUvIm8S1AXPl7Qsm8Ebqfj3VEgVD73Rouw2UEnR2uTVEnCAQliEvG3
84To21zxCWo1VT/hAw94OMaM1Es8g/uNNjrXjPlgN0P4H5FYpdwTqI/k9gaQhYS+zxQEn+NIOCpM
IanJ5pEZ+I/jHrvfbdhGaZMqYLmMNhBcOIRjrv4HU00OJ971TBUu0BfOiPb3k4SFqVyTcReG73gz
E9nDLVASvV7j10C1gRHwEGx291OIQeQZ0euShljhZvum5vAkgqKWqEk/tP8P8ObCCOFWXfInqSQn
SewAf7XkNjtUZhY80AoEpvXmtFN8SikLbPTndd4G/T71p9WgRQCdpQxNqKretZauQNiOUeH/0rba
mZOmlVn8WZ8kdJh6gbzo3ZcmB9xfU0jK5YC6dAto50TlrfjGNnKEhNI5++NwxgG5jTzgxxicvifD
2zCAH+B5sPxVSlF/1U876gurI0sY+RDq5tpRHjawG+2LxKycAECKAlPBSlyomZ+eW+BC4uFuSsFX
gX6H5AGWIfZN7GBBLljMB6TzBUGlwRnbBazZ7TltKIF3mNQQPSAXMBBPsUdyBllsQUps2OFSwbUx
prkYkLINV+Nu7s44Ma47slfNLHv5vvlLip6WmHE5W0f/T957wIVu76tJKRsxlq9/6iwybc6Uxbnj
Pd5VXKSooeVSWo8aGbR9nKvOWrh2328j5UuQ0idXu2t7MxT33VoswuXu2mZ4849U9Q7xIgwUPSa4
39Mp5+u/La8s2H1yBd7J+YGnRsyLWCOuPpL3p5DDb0U1/2q1RkwhTamncs5thrlHZMn1vUuGpaGk
mRVEl+gEV8AYdmDBJBOAgeCGfjodjJAcCdH5FLjh1vX6gUdtj7cyqd8WGYVHjQIZWf4WqxsuLuwN
NH4e/7azwftEOs8xU/VaGTzWEa8+aq/s+JFOTm2quS4tSVND9X39LcHNDtS0Am3wO0wjFh6rm0WR
QC8zj0RlwADyt39gooUjpHWHEgO6zbQSXulyJBL5aaNpWRu0f5yhbiwyA0lTADmPP9JpI78+w+sI
CwQzVDJcEN/YUyJlxvic6t6NrHR1nNdNkjGwhC9Xni7Q/ybRwhciwenRAeZk5+gUnbs6DRk+IviY
Wnu/h7cuODhUeErP8EsBfBd5OjjfBdJDZ03O8Hy6+lJYV67JNf7L0iPNpUnREKdV+FIeJcfYbddH
pf/eS0i5yXFpoUKG3/732KTgNZfAub8c/VTgqMVE5awKU3MC6Pw6vOYfwbUrshLD68lRwJgJJAyJ
OjsdgHtw+BQLd+58j+lNlnvxzs4Rr7mULWWQEsgV+EG2FFZNJJIfwU8MS9lEfsdd5vsVJW8nmaEJ
BKB+u01KrRDJ8hIb5autly+0ypAdvsXq5HY2eD3CVa1yI8oiqL9OkNB/gmTY3al7cmHCJlnY5DZr
ay5VY7GfOui5OIW+GW0qht9/eJhNPJWahTa4SXlcs3CXykMpZZHrY2vrg9dm144D/WgLeVU9Z/v5
/R4XPo7zJPNeR2Vp3y2yQD/hPxIhdKr8OWID0HGNgEBPbmlrZfjK0apEBwTf05yH7RIuvi99/URn
KXpdn1LJ5bd0Dgc5a7Uk4ZCcmLxAegBraF603LUDmvPjJnO/YZ704MrS7gw9u/wvVqQ9SEhxmlw7
VM3Ys1Io7tcppexFMqOgTiMkXn2T8vdtq/8zo4dBs3H6fyvMxhB4qOeofIK4cfKzvmu4Df/E3+6l
/Tp/j0hujGyxO2VALje4gHFkp/ae/b/AKYbQ07FKfrprE4nShidsXypCZ5sSy38ZAZoTUfGXnX7t
bLJ/Z77THih37unBm6e764jQgW8XwQjLvhWgvfP6e5G/WAPmu/0R6RGqN4XQekbJ8sv+KWs1h7KB
4Is3XVXtghKtjezlWatYRYB0q+/aECTD9iubAAJv3rs5a40eihOG5aNdXSAaQGB0TY1dS6AO19o5
ALgfZVxxIYy3kfAE7W8bmBFud8xS8v+qNujn0xpX1BqSYNjtOM/GpZnEK3nrNo9Hn5sWIDJhv/uN
af1/ulDGmegOfs4/122o/xigLA5Erclm+mnqeNQzk0n/UxQiVi0sLAzygrKDGI8KyFZrhMh1mUsP
BueCpfUwOncJAwhlQKCCz6LVjR1qeG9uwS5Spu7mwy0tfNHTi4dvwQMTh4Yp7V6J4fsCcizVDX59
aOI3Uj4uJt2COPvLuqisqIZISCY8k2RUVyAKhnjVNjJraUGejBCHMmvvL4a8zbpJBWXD2zgkbBkL
Oatn72KrxmJBiWqXT6HQwrd9XqYK6mVLhoCntqsS94SmG8jyU+Sey5MJ+llkv9CtHnh4ZS77H0Zy
u08YufvG0TsPt3+0QyA6oh7m8DQE1/ug6B9oBm7kEbjhVSMlRsZeLV3guDN29tD2HMoseMlKJodb
jlEuCrxi8lpy1+T7XCh8Qjv9/DHzAQPR+AGLmhrLbHky1ZUznG2wLg5OsEtBfASMBDNJdvyTYw1Z
DqKp9sMnRcpAAkNrzOMGwcb5oowS6ETCE4wqTQ2S/Xzz0oTc9pNrwrXjPD0K7Svw6JRdTPJ0P/v6
50GhKCCK6oaQ071yGxGIhF3dxBWXjzE25wetWhthmPtJ4wWdJ2DYwCw6vlV9oCkIu5/J3hjgqABR
MGtEVe1sc7wfz9thC89WIOZ05nwer6Eg9treQWp0eQyVeBM4XltNEst3VXi6LFhvb9Cb8Bynm+wq
qMuD3zG+nIhHgPwF/BVHQy85YTaqMuEK7vcSiLQUNTuk/RmN6NbouyLFGyd6LXs+4KXTVktdn+Cu
qvVm4R28r5OyJ3/NkdW3gaw1CcOpL5Msx0u36iO3pQTk57QoBjoEFUNlUYlIeWlTlV1PFhhbxJS8
BF2IvgmQsIweuGYxY9Molfw0FlBiGXEOcL9NUKsZYPgFxspqGvFZegS3F1YwRC0H+bPUrSW+0YKb
PWthb4YQ9tBeH5dI7BJiNHmFJLzV5ZqSnusO6RZZTEGf+hniVIhVDo/2H9zrRyfjda8/i4un5Yjf
pAKpyGD2ZJhk38/+7gXj+DPa7fVlphMusY7PQFp0nZ9AHOh5Ykk1ERNl9ye1fDTE5x3Je/SDdjiA
I4o+51pEH8RY/zR5yxjgO43kcRanjznUMpKRh5fEgwrSm3lXBdyMMl52eEGpT9uEnTDF0vMbtPTK
XqS+GdzGjgaZT0uQ8iJDJw6MiXlU90/n4lM7pSa33stdrGyeSpRU4QTgylC9bfVWEMbe7Qn7s8aQ
9KeP2B4cjQ+fVJEXhgEqsPanrU0Ung/+SU0yyuUIqGrPymdFYJghqJHjn2/RpTupvU5D710ixEt2
ETUCcTi7SBRNdWInMO6k/z3tHwiTmCoC9vOQFmZfCnd19AcsaWc4td/H7s8Ht07ohYjBiKNIffcE
vcqSloVTJWGh/Cxw09E2wwU6DdCyTuuPRUuwD8utdDWaMLqqDA51PDO4SjWWhCT547BuOlNR5W9U
CVaemazUxpGnc2/TeilAemsps0ZYf6Y09DnRgrNC6ajinbrhO0/CtNCUuWYvIydLcmst3fE+RBNl
rf2x6RfS0VNE3PXI7UiBBPFBzxemom+g+aFfGWmi1aw3+rrwVP1bo7T/Tsmt7xt8Otq+ASBrPREL
xxbUHkURERbHyBicss9y48/0RsySVDgwWjbqSiZQEGHXs7mbwHS9An1MKH3pjMPWY+yGYa3KNNkn
+L/x4B4H+D1CmylexhwVBYTo7PRyTNEZnOciAO8K0Ui1WPRNVJX90JPxt+u4Ba8R69xpuLdWodhp
hVQot7wVFEStr5XIuc/plQNXIVRCvBdo94069fLJZAlr09J83LsCe4qnJgMgl1sAJwLWfBg4iSda
tVqYQ1Jp7RLdOab7SgC8AafPyNTKcMEoMm90shBhiQ4fH+PylPFOLzB1yhWOKqy56RLkXK04Yteg
JOdaPn5YMU36nPZFPJIRS6o+hzkf+UrlnPOmXXnRFygm/Bwy9NEPYwdbyaNFb4PzXI0+9nVEPt8e
XDlroglSbbnUEZWUfdhmrCgn+lZkZH54yGvWAEP0TctUeJnf/x94nNbAzZ0+Nj9FokS3hDfuTr4R
km0vicVO4F1HGfPCMBIdD3m1BPEC5UDKfMomIja1ju+YHwygpHWDsz6xSz9tUsq2rj58XjCLoM3d
xa3lAtFjvi2/4TU8JyaSoTKOssKlPEJiKj6hm3rC06Y6yehpwtWTmCvypzVJHxksMBVJmRubVEJt
+p1YabemjumPvU7OrgArTar9YdFBAjtDj4lR2DI1re2rChjPKUnf1k/1shgpwxc9W8+D9b5i0Arx
dKgx473ZRrkHlmdq//UgzwUs5lYLmOciRLpBwg74kBPjOoJy6SY0NzWoNkxZUh5jehOIfsF14az7
fhKNFXnMuNzyeZc+MRHjnyhPrp/pDuI+MkYynbw3z7wYp5Mx8MjKExgA/wG3waoWY8A0x7bGX72p
f7mR6RN6zVilQ64bciW2pCtj49X1eI/BCb0ZFpl+lYaKdf6EPbROdmKAyTqmVCItdBq3L/cigK0k
aoiGRzLZoKUN5mgEIl+qEtCjoQPfw9T548Rrmatj49ajGrx6v0DTWg2MBDkH6uz0kBbZSyctc7Yf
eYD9jiLW3tcIQy0YnbQwYMcaJ+aHUb/jhSv3FMy7MmsTsd+Nd8Ekzi7kf4bSIysjYXhbcyBoS5HR
545yH6kCijorRnF3SwzqT/tPpI7b4Kz3KvYYhmWD1i8bdVJRuTF52M73poCtLI58021iUlqSCSqA
6CtI82vXse5jQg5rN+wETJpTdk9gwMu8zqKbudBiErKpXgedM3c5IkifIJ21L1wjvo+fxhfd9AEB
q/6lEC9fxP0g6C/wFcunMLfSgE+Ve+m5A3pxsS1jNT6Nemnc/+oBcK7yiCmyEEnsZSXk9AibPYgQ
TacJ1KezuhEOo3rnxQp/KTGzgPkfQv8p5XFYrbC4A6mYgPzm26bKtDZ4IB3l8zmlt2bBUsQaZwpn
LnuqKURjyBv5xZ1UdtiG+aS9ysj7qIf9NPqbMD6wPwDtd32lcXXSyPFctSEyD4OGCSdVMCdBukR8
/z/i6qvKise2o8gvM+7pNVyhNNpHIJir97edo4WppvDWGKRdhRzJh4JEO9pr1K0RztDlf9cjRFq2
QYOuENlTLZpyeulJZFvdWReiOly+QOxqpFxt2meCs3nmufTQodeEtcdGehehVlHDP7bzyX5HmXmu
41KHPAfkdw1XVt2WgUDsrTScRk9BWL3SuxQob+gJn3GMoBs5UBf12Kbb6V1bO3GuyAYRmDydtzEm
pUB3VdYoxQgIZWOR0M/L6e6ZfRRJaplzVR18Cu0cugRJdLqUaq7xSO/iKH8hnaNIP6/N+r+NUWOS
dkIC7mmhKjIGxTqfsv5wADuEJ1M+2auuAq5ahDpDXefYftTE8Q8AEie1vc9r92txOY+44LjsdMKr
f/ZBGhk+8qaGwJ1CeTUQO4eZ2np3rCA5tJA/GDRJMWR2nCKnEEGfPO+ik/ceCY+wgwazTDPfr+lG
BFvEVyenWEglKrrTfO0wF4JS98cb6Y2C+7FkbBMFrpGtOufhUiQSeMz5Mi6/3O4690bypy9JxMXv
/8k13CGvZywGF0SBzGziSJMmEUbtufQpZzh02vFyB9HFad+GtV6loZHPa8ZAShtjjUqJA/zFxGpn
HEV8Kn3o6ufAptdJ8jxEYg6ppc1ATUlxab9NLjD33AMAQLY1JsAjVIEba3ZkTvxC6lCTgR8gW16t
syftuPT9Z79MhHd4qt6suy06WtOhhI5+93bI5d8UVLp2Q2l0g2vlpoZlVYXeHeHiPZAMoUaqXi8v
V8P2Lz8EmLxLWbM7BE+m8A2foFp1ewwv1MqNR0QhCvFq0BrQPs16YUCcBHu8nmK5SF7rQZVKssJz
qppBX6iavpttQBMf79lelyxVOuN8H4Ac5DbfiPzA5dANyAsTbLlqPPVWS5rok16ThpCj5jTYm429
NPxKXY7iz+H7tPTPwf018QbJF+CLpIohRDsSDm17+khPeuQ2AIjLD20tvqH/h3wN6GAc4b9s8rmK
Ux9Dn6SSfNtnXDhvQAA1bIFT3H5/XutspARDzVFf5fWhJ5JoC4R6NppxBPTWcBWGfdxwUWZ9S5HV
jjTDnfb+ULTzRCp7JdZu4uknDG2QcYaLBW8t2EHBzELMiBcL4NS5FmjxydgDKWbcbjpiHmBO08jK
ML5NzXAol7X5nbo5jXd93nj94YmmJU2v2CNvK3TEq9o4NdXxLgAKi5kFl88Z2dpWnw9H76YnSPjP
PFNrgiTZp6vt4pV1ogOZnGFPTvnW5ehL0EXUWlxdfpAY0CHQPuo/21E4n6P6TBlyMejq0F8nbe2F
e8cpJDNDU/kcAqJfLNH1MoPVZ98XdEMyvLvUl7jEEfplBv0vLdOyCYnNXvF5p6r1rB6qIiNQSzyr
Ksdu6iLZiYLxxAW1q65CLNpi0bwmpga6jzV9CaB/8KHvLo0YakZNExMab/ILhPIlfaC6AtLZykx+
Wv91BDO/OogsTH7hOzGyc9HbRMaTpnGssq4tNUAT06V2mwQ3PF9k98rgvZugqYJcR/nQC1mCfu+Z
+HPLENPPWm+GqySjkRd/6Yj7X0ee/43LVZcfWl1xLoMW66pIepRy/pY0veP150FJMLuCyeoIXUy6
/ePsMCahGol3dbB1EtsHwUlZ1M7NmZdzJAiDRYex+xgRimGen9OC02EWp41ugHqN7z2S8Bx4W5bK
g1Xz3K2RjbuiO/jnKbiIl0aAh0Y3HJ56SGIeOOH2qCcWrr53A6OFdhbq/g5JgZbKcSmEfRi0C4p9
5tnbDkQiHUqwCXnd+nMN2R5hIQmi4Y10SEx3ae/hUTYvocR4tabxvnSlYaGJq8R+LARrrln6jFd8
jUnGwQQPtDgazDoVox1wKVyECTuOvUOvU/DOT8f74s5a1B7vwpbsSpSP+3JrgD62vqvAx9KJta6s
CoGpHDKXzkgaClxV4756YzXuP/0CAIQBr9i8RqK7R+fY0xE0BD7KjEc5QwsDqSBX0K3BKYFjhoMp
J+AI/ncZHMwAF1Y+Oj44vcJmpvsRNG15eKGO7WlwwckAAreL3pT1601sSIxMdUqdyRARaMuNZKJB
iXd4JFA8fw66uZPk6bFhkccDgR53L0sPjIF3144Ka2XasVL45nuS0JHjV93NCS8a8Q/uG/ckUckd
ZMUbBquxFXP/FQCXmiYtIVRQPbPHEgFtZp9hcInkHf7u6PFj67be0+kjh/O9r9PWAq6iKxEHWL1l
Li4c+Np8E2MWsIKe/gmdDripn2Odrk19Jd70YOSvCI9fMd1yE9HW0UnjoXYayJrpnJCX+Ym/6rbU
5I1bc6diFfrjWUlT311q8/4syspf2Uo9t6HaA7joPRkunNpyzrJynK8+hsj3Y5tSaTD3rNDQn0FY
nHy1+yvEIuHzEhnchAmjoqwT9Ur0Gt3xKPPqlZYxO/D9RhVHG5GteRJOKU/GLwOYKYkzGmVcaMrg
9ltAlErTU8gKHCd6djW396eDcI4H/Ghb0GvImNcM85zkTuDBIHu2VWTP0xvTmobBuUrVil2HMmLi
diCEGoATIvIrCvRwFSHXjFd0fjLT1ozDDzYg3vTe4zMA88nvY7g0lRiGZxjSlMdPr1b7/e2lBEvK
kfJBTfG+6YxHc1qb6HC3GpOX8+epQQT+dkOf2DUu5jnXZIpgl24Chntrw2nFJiEDCDrdRefka/EH
N3eRTJnkWxO0J0t6ZSUy50zeux6s+bFqKqSht+WMo5V5bwF7PmZCOrlMl//GmFplDT5L7ShOb6Ze
dIpDBmydkn6A3vcKYnRc1Vq/PYZykuzhmh4NTnaytBFjA7ds6k5RvrJJcr+Mu0n6OyJk7rDx9SeV
HcXsgEW3ZznQGbNJm8K+aUMMGqkiQTLydBk9Qs3XEJg8VD7umYJzkGdK7BdTMry9Mfvgzywmt9gR
QewRRHzV9ieSwyMtdAEgIkS267r3HIpQhOVuAyhcxmD7OyXTgKTk80aUamrtknLZj3vq7RPMvdLR
fFEc/Yke8UduCIPqSS9JKX7TKfpOLJug8GpFRBMvaLvpYP3Wd5rFNcyXFM0JG3z5hWehvtLKyBVz
qH3rPkjuVglaViG1GJdjhUtUtXyYyUlOwOAAp2fmi1mm59R4o5MBiXVczkWjf/4PpTKCP4FKtUld
YvKIJMqLgKRc2GtIGO2UtKXAirEsd7S1imAUt5leGd4ukMXIn/Qxuf3v27L1JhxjdoT/zPqTNFIk
FhdqwJ6Qczfc8tJubxqbCSuy3ALxT6/Jf5PR56ER6YeAfW/43sknVaq/a5lp0XL4CxLDYXtmdPiA
79zs3WPi+AbLHVjNquht801vgG+pUwz5w54cWka8ubhj7fWDlx4kxC311hcATip724S7O/CevU46
/EE9iy5q/eF2eUBp+38L4DBw/rasJ/K6OyhS1Kjm7xP5kqA0B9W3JiiZF9/7goV5LodEm5umfla6
/ZDOvQ8wJbsD723hAOSDJ/Y6/rcVofuAsWvImwtcgdti4lo6Lpd/DjbaFakTZr1AoZmhKQqTmWD7
NRnWHNEVhXnGxK8kXshHpLtuMicfG+R90nXtb+rDN0cIvaJsTR8TbWdHkhhQDFHloONzOiR11w5z
08bVTrJ1gMxFbJdBl4UzwQxRzycF8cjhSEdcQ92meOyLjaFdID5zD1HEMRTxnwh+wMd/qOGqHynK
blcsGEdduI5Fno02fQqqWeK1zlgzjQMCx9fXRSRwym6dfBylYKYfoR17xcBy7GfNmFYNwRDSEY+u
QuRBleBeSpSqg8SJ35Wnu5uEjAQ/L4Pca081ThFx2y+VHxfJq2cgwuuVweijoLCaGyDA7OEA/7vk
fCzVdmhSioC+DNTvZoXq5P/52c6gTE+ZW24VXJUqg2QUi3shRZqgWi/YZCFXpcQ/cb5xApAAXXok
uoBRcCY4wMuf+/0Rz531m2Frl0vlbgEcOawBJfHqm9qofdvVZx8ZDRxM9Z0IEapMNnJrsRw8YvVD
uJgtAbEV8j8/4RzWsHsbwR71Wu4BXSKzuEdUV4nS4QdBGno2mvSK8tA0MpIb1EZmWmS7/rXoNKLl
dYiHNLaVmEx1yhR0AuUv/eeFb3wZET4lVe1+DGjEUfHzqHtEXQ/iLaQjW0B4cOsU9bwPuIHrKYL5
CXmiZGjN1HoveACctw86XTANXPLZ9KLtXjqQU/+QYocZRRxqDC6cJSsJ7o2bbd8ca85fkzCHyVPc
f/AVhImBaNxlrHq4erXuRuFDYERN0Tkq2KmylGoZdDN6UxNy+3B8jy8i78FWQoL8YsMbZgtEOhVb
f8ACka8uAWZoQEdNiFsh9BWy3+qNB/0npiysbyIEBch7FtBHB/4gQP4Q0TnnHZepQVdaYT+QuDLo
E4u25pG5HoW6qjvBe3kE3lDuA5lXvK/LENUanWMuvluBMx2ixE3CBgB2+t2daDKMCwiAvWLOxT96
sjbFg/BqJUkG0POhI+mc+N6XFeYmbS9vd9mLPyIWZkd1pdeOrrQGY9NHBowtoQRs5+3UVzKPULvl
8aNtmZXCFf0mc4x2oCcDnxWA/dWD2gsDsMfnuDo/XZSH+CPZg0wsd958uMrVoL5JjmsYPxHHJe+t
q66GEVPT1D+7OONX19y9GNnf5iBxcUM4lYtUmJIFvqLFXekwdJThkonXl7DnMCxtLj8IxdQ5hJgl
6PD6TihAy+RtHwC5Z6+nX9GyXZJhDfgktmBrJbWtmQ0T+NVmlktskmCEs2xPpDdv57fZdAV95KBW
GNFmxsdGaoyZ11oi8n2f6nBReca1P+OlPVTQMLi5KbeBfIH80HYTrzS83C0bzx49i5D7vwq2N1if
C/To3VxJ2gq92KdnejrerDPHmns3Vh30dtjKtYOwUxEewfO6ngH/adsaWIWK/celx0mBFZHLUHS+
pR0FwfHvf4niz6a1U9EFinPpqgsWy0+OozhuZv21+MFE2JZG4s2kf+eDQWUEMKuVK/fRFVfnFHlq
lhASyGmVqi0ku0ql24aS7qKMfkcEHHy3edwZVG1fZUJJjM2tHsO3McYb0X0iMir7D5ACGXI2UJP2
Fsu7vWVG3p7s6jbK+aSM0NDFwY9yJAiPczPProUEtVcUUAOQztA8HrK/mt1XBFzCu0wAHKFrXbgx
uBBgeN35RXqwVUbC3fjrk3dQnN/iZnThYld+AmO1yAO6zaCOlpM1n7QaQzCL+3dsT5zeb/CbZPEp
cXWW6Q4HtofUT0wEDn9y22nX3mGNYx848hU4ZksTZ/gUcrzOdi4MEjmrx0BrRHYT33MUqYOWeOnI
5G/JzF4QztmsOosJnxOKWt9hZVZQ6JLbzLGIBjXx63SD08EDpHXwo/KZZhUQ6J1Sb2suZEtnhdlY
Bj3+q/gZqiJrgNWG3bA33bBgDFD6LfDNZ2c8+GcMK2Q5EORcZaklRj6wWZ3UZDWOavlUa7PaNet8
huf9cfeALlAJ4UpzSeVgPk/as2/IbKtDwBf2ujpZaG633vA1KYZX3ML4qeTIvqiHqAKsCmA+rs1a
C26xASKAnrG7fXhEdm5OguZ+miyhuSqrjfRqrtdRqy73jUBng8m52YORv0IvV53S7UC2ugnS/r8z
R+arxkKsWilwDyTZ0GmnqTTPBbcnju6OwyBSLcIQ4K7KIkVshDZUHCIoPZBzJNyNWU12Lnpg7w/h
X/N7oFKfUJf+lPGvvyT3Ej23jISJbwOEU7y8qWirh2FOmXJ7g7glXu+8d0TjfaWH8zAcCY85c49M
H0H33v/UC8E76gIBXEDrA3FIn6+6Aoid+QnqaV32ZfIOCqDpCB7mEWm3entHpjl+2pTuvjkjoyP+
X3d0iOnMDKYmHUmz96PjwQti1yiyxZjzyMU6VJm+q3RkBLFtI1wO0G04HzhtDTCfIuE2G/GlFFSB
xuFYejCIVLqT2W4qH7/pGoOFdBuZtBGpAHvbQEDiXGsf9xbKTi44VegTK6G6u0ARAH02ZgzD+t8L
AQqYwA0LzWif04mZ7RqwYdZCQkQxwYGeuPSkJ41BYLL6UporHbZiC6Ao78VriFtn2pnjSExsLZyC
KcYrVqQpOsYpJG44uoTlS0tCqqd2CWdTBa4ivwxxIuiRRYhhdrcqS+MTYNGt/tin0BtSI+IRvrtT
RnYz2MZ3gXyGkecwAIE8YJI/i10KZbK5H3Sz6FX2Hn/uDXOE5iAHnJANZsanVVWwtjQKtmB2TKvV
PwLCJtaJ/3+KBnYoQZ9+Ocb53o6JUZWbo3mTZ9HH7idbsha46wImcTs2SgL6XVyef4x1hCSsCFbc
uwgJ6848B52afDNFUzkGIV0DXnBWjGPJleYv28oumZI3s5y0ialcXL4f0VZSysnV/DwFGIlK722/
akonViVJsDmorC1gnIjKoUFjMmsjwvoCmUsTZXQI6W1fMfNX3DloCKUvbZI3DiCcquydK+qTqgKR
5kt55glCWTvdN68AGy3XBW/ti8y1U+68kvETJRsSCuItRQynkeOPj1z243KOttfRqbOoHNzBZijm
mzIbc/nwXNhtwJvrY9XQ5xNdHcN5b0PIe/dQgP6gY9EfJSRYOeZQ7HrQ//DXpYB2wMmJQc/WWEhF
ZYDDi/KQ8jom+cN1kMMdCpXwtrPimrGD9xTxIHiUji5ODwIAqxomjADHI/N6eH6KXVCWPWavKJTY
5POtMjuTZ1UwbakMmYAviTRDFf8ft+dcn2lCP5jjENB2L7dmh2umZYh1m0fab8sSsBaCCwfKJZ/4
IkI8jXSUinoZqWrY1K4IvK5rzhFN9d/2Oxr17I3/ITlR0fVFZQSXcDdT+kEh4bOZUfzV5fycGEcH
6eOtze6/zmMubFF7Xjq+WedWKR01xe2521YrtZa508oZwS7eHtoeIkaIrSuraXPr7UrlcVJICuYE
pjkoR5OoD69Bkc88Ca7M+KYOvkZ7KyNE/f31q0P4PIY7JiIYof+QgOtj7mSwQdeDoQoKjZbUWUoM
pdTRVZqocOMnN5/l9g+MoAglBacpM7yy5VGh1APSz07eug9X9+rLqx+S74uLG0F1ouOVuJ32Nqeg
ur3tMQ6d8YNph6pCxnyOX7PvQ4mDv983+ViPYVkzsF2DSnLE8YbBmxp0dY1D9A1UkhnjcNBLx1Ck
9QuoUEdQI8BSnwewZYPBcijFX9lwoLubSwurCACUfNXGxzl3KaTYSeRbFkEee1hcXr6WqeC1Y2Xl
eTCF79bNxz9/3y9Zb51nXbEWfs3VucRY0ycVwQMTBPx17TeuczsLL3pVyjer+j1NgI07/x4qLm6d
moBfMYrRpzRs65PwcSuOfGc6eLYE0D0LqJfThD0sPb4Cs09A12E8qCggQ28ypH+jY2K+HNvyfR61
xx+oduoSA6o1yn+FyydyU0/cuIcgbDfy4i4vc61JFd1Ypmp+12DATigiClnXaMbc40eQ3i2Ema0E
0Y+ksqIl7l2lTE2mazjnoeDT65S0eQU+ARY5Ia19NKTkZxgkJqpNFEPCKKpnCnGBqTKpjGCt4+dC
RNza2XR/NdCqzbXoUMudvaYfCPefnDwgp2WT55wD0i8FyAjQ7o1qVwAxcjoUueeDnBquI+oVrbcz
/4P8UozMijalWLFgataWMbEyX11igMhVW+SQNEtmO4NBSJz2tfnPJDU3bcDBwFOdBrCd6y5pKhC0
klEL5PJYilsczKxzHLdobz3AuctNWa2LSqSWf5nkpCwRwDwV9E+RISPO0sVG1VqHYcvO+c4ovlB3
5jeW+E84SaAX7OXDmG9JZPmoFY6Qy5G66tryGATWLJK9LioIPEij576w1AVjZKUHKFjqi0SY+KmJ
+Pp/WbzAAqsbB19CoKs8Hz6SdHU3UPgoTozSWpNik/NuslaSnBDSfPL386f1+274lgYl5v3egQOE
Y+EEJb+0ZjhpU9mbEip3rRlVj67IhbRKdzhYCTTkqw6+6rE6Nd1O6AzNaaoP/e43pBl1FyXzrqfw
aUr+zSEZIXlqFDQbQB6IYxzxWqGN0n7Y7LRIIoMc3fadxu2nGH8PwwCzkjd4Vr8H362zk9voIMUj
Ea/PpfmtgwSF3IaKlxsMFC/wJTuV5xI2ihzM0zXT47BFeGsvmcgEZi66EiA4sxTCS7fPHCz8FUff
UH2gTdlEF06Z2HiK9JZnQWeUVnUDvDHf0xFce6yhpsPvFZ17/QnAzFmQwqsGgTKTvEfDlp/KREia
DR6iAPnd+Jm0oE2tsxepSeT2x3O4oAFtjzNu++MtoBWrZj7GqYEzI0YxGhiTmNgljrMqdxKFGKCu
Mv8E+epvT0fPujirv7YqR4/FXMNZybEFlaHO8fMPKoAomZhbY2N9xB4ncaE8a56Wtg2ACEc6OkYi
8335CXU/fC9ZYO+wLWJel293D8A4qj7EbMiP92TvhsqtmKEwXB/p5yuDCYR5Ph/cgUZ6Zv1TlPXa
V4FhxSDh0q9/Xry17Mlvilmkhwd0fLR0dM5IgTfPIf0TfPMX4l2HIjvsjYwEpP1GWtY2g+G93+Br
rChoa3hRpOLROvEGlSH21bWqv41QI2e5pkWTgp852KnA0Uc4GzVdnlHjk6dCNHwgHj/WMb8N54vJ
X8jx2FwusJ4R3TZ1VNKjoRI20S5/dAdo/pdP4rr269JHEGXOaaJoMiG/NtaUrdw5xF9+IVnjaxcT
V2zF0baecC7ZNXeg4E2m4qVuJt7ZiXHdfR7vf4/MXujkaCkqgDG4Pglf8jsnq5qZ9jNcikVxbdjI
ZRi2ga5kzjeTgNXQYGIqKu5w0OdMfA4yWTmP90N1G/4uNPVT+u1RNrbiBbQ2TtuAevVQ3InllZCr
7R3n8Xx5mCyUX6fR29br0ZCK8d9ZaiFzexVy4eG63/yJImRpA7ND7JfSaVzJ8WSAX4llRCkKcAtq
HjnBP4yTJokHy4xFEjlY3O79ELRS+Zc8bw0HpNXi+gBNDKAdqbe5gVYAk/cE63NNlrHcVN/R15aW
G0IG778pYjwgbqtPkDlcu/mv5emheh6UpenHCPC6yVhnLAPHAQZtuL0WoBOK6EJnChymMGp6DbVL
fjuB3DlUIe3opNJjRCVmvsK9Yiy9mc96FV3P2YRAgvzXU67KQoc2s/70qfSwXL4IgPLPBRn1L6Pk
fzruPDvUOwygnBf6Ma2VWUG5TqqWICH3xCEERBd/8F7CJEl8EFFa+Znxzgt7bOmFRZjHuRnxlg2V
ZDlyP+cpshZBsvmx9GR7JpMDO1iTM4M7UsPF8zpNJMrfNa7QB7WLmAw+pNsZ25n3Wc+NBj39VKoY
nuxNwmgVNS55RJ0UiizzPckZDZoOfsSsisiYjqx7mBf+kIelVrOxJJcBWGCeWYoHI8C6ptjAsb0a
s+q1R9gF15iwhkWLGAqgp7bQANWzAI75zcMurL7O8LNKR1khF6Yh1XO0tXunAbg9G3WXlTVEzj+I
UOve4C7wbVfoByHhUTcENX+bnHzadcMTJXj8CRaUYejB8lDXgT06+SpSmhP/D88uWTXT0iSVZsUf
A4j/kZ6LiFuCTLG8XYBWVUB2khbK9U6LtLvMyZMddcn1CciFRUyCaOW+V8d1ORCLfpaiCTrhVGA9
cSRzR/hP7+EMRthv6fscLBjrMrhtmgbeMzO0rc/nNgBAaA9ViMXm6tXv65rUIULITy/pR3pgM7d9
TGex52BWk/sPLyyMNYYCaPBlmtR7U1J0/sGRO6/hHyFv5twPtJTmDJkdszHY/WOiAZPNqOki079V
qedLp3ynZZl9EM/Qw/3Kqqy+509Vi4Y1fkmWFpQT6kiJNje7bi3YEjH3tvvq+sMJOEu28+d0ECA1
DrleQpoZ7gcMxktkRM9dy6G60NtL3slXbQTe5f8NShyig9+mq1xbY2hsrO3cMnXP++hSmO/ETxaW
Bh/cPc4AQGYng6lTNslBAAHhmCppzX8DRiRTsuT2JQht5+5OFj6eW4cdckQZ3JFue0ibrO/mx0uf
ups/Gyb9dxDOmLV1LhvbbCb4srHeiT0hPjepNBjrLmz04X/0exO+PPYTLieZai7OXhMIC+SNdmZY
j77eI4FkivdYzXCe7Rnw7h9EYnynkC2kzsj0lXi6SvAuwnEQTMxPlQm740Liuw1d7QowQ/eHB8Bu
EWIvLab3Ulf9C7pTziCI5bl1xyUO0noIXsg6jtL5aiZ2ZHgRd9fIcjc8HJb3OV864iwsVUnvN5uX
QmOwUCP4xGf2+UbNSRrJib/QUQB04/ctcCZcPF/c/WRtmyq2I8HYL5JBuMQ05fQV2Cvx/O9moPhX
FusJnPafx0AbYO8NYdc8ZPylG83IvpJjhGm/vtgQ/s4dHc39OSfOSIyRqkw8MJwlbhk5A2cC52os
rnZWJgp0dUe0v0toIrQdAVVJbAwpDTZihajVsjqJE4qazYjentQHNOJcxlhWgI1Iu5ss4bqSh6Dk
6Gf5B51tSbvA0aumL53+D9zDsMj08hf+0UITjRgAU16v+GU1PWZtpV6NNm94GTZMn+c0cQ6bPB8p
WK611sbhLyL1jWhHHSXOC4u1NVSUxvvs6LgKZb+EMkMDVOeMLY4x5njTod0drvDaEkl+9TP+ezdY
efXHizZx4l5/Aj667Q0EAlKjiis1cSBgwF9RVHY8GKeJmeNf/R8Z6qSgFKbXD3e3DeeyD0ZVlR3y
cvLrolhzYouXGJmZ7BlUktmo3c8M6MCV2rdmmrqk69RrwDLBuimGJy2t6mjxw/2kVsChhSAlFNmu
6/1u9uWKaOlTRHV7oDPLzVzxtOv1LbDuFec4FYeaQthUHDypeKGTYR5dmKtFEvGLlu75FE37+wHY
WxbxAidppswYlO7nguTR3xOlkoiTfwqefeG9Pz3QBlzk37GvjPSFdtezhcsxrRCwezPdMw+Dagd8
InPE6qoHqsX8i/0Xs0cesnAyWDTDegFqs6kWZAxtwse5uxkGHpWBhxTtASoFJ+KsxSan4BVEsnnt
E3hKxck3PXUSWNYWDOLKMDrlu5ROfu+xZd8K22aofscoBaX2o9/vhMKZeEig5leqOVp7+Sf7vpN9
mz38LhjbJZ/57Im2YHREANnGyrAlEkuUacziSMu1CipPvJPeO15Sbj7JpCowY7aGgwixH2P3Dynv
KQZSJEgN9gbQodzQhIW7/7pBkgBY6GAdUFG74ld/OBXwitVYmS40cCrSwfXcZi2dAxsGR/ZPLffC
psALYxt/0iSOGpt2WOh0fRWdEOfL/Yq//OW/5hsMP/rd1o3SithEI8vcj/qaN29QeWrGVAVFtjhV
87IVVt2bhlrdBIDIM3wzUVnyyfZHhBS87oCsSm+ZIVqJfbwg6DqnGu7NV/EwQ3jUTYSLffkLkmCF
I75PrXUB88zZNIZ4D1bB9x8OBXgRNI5QYJtWqCapQhNBTAir6tpyiAvOmWTzAokwiWE8u1dhktFb
pp9zgZlcVx7tVWlnQM62dx/sY4QPcFAkLvjeKUqdA1l3Cj9jYBDeNvbfAIKogKl3NyRV/XY0Mpxa
kMK9im4xbvrzX81j1xaueN11uPK7LYWKNwmgCpOEUZi9swB2f0wVZI9zkJ7FHmMwvBfE7F7zhyec
VXFdrGi6mTt1dD7PeSezpPlo0NOhwx20oQ6BBY/UKA1hF+TvGInNUwLla+/oLFoSSLEdPqg8JSlD
J/w3FCralZ/wIqNa2XZZpxCCXHuYgZ24XaVjPNOhybd971Md0s8VmNJkvNyYP7lfzq6+2gJ1Yn+9
jySsJDbLtvvmG5vPOorOiZH+/ubyXgFP4EkuGBKOyD1ktZNMOWzUG3DoWLCnBo9Jec4+FCdcDQFQ
CAMxZ/8Kl6+n07gI7LdC5Xz3Qzr5iq9cC8wIjbuTkgYoGH4IjG+ohI5yNOrwAngXpk7gWDuO+65K
vZeYe1kuw1Yqqwbx8cvnBqJVR8cxkhUmlIQe8Lmcx1a+xl+nzNWHw7gjRdrq2tCsfQhUTv/MGy7E
55YXev9V1GKaZyKMS6MMR3GlFu7TBR7F4t9I+L6l5UmH+0aSAIZgHwU0dRtna1F7WhFVD5wGUkuW
vPgNdhWVPnA7v/zlKAS55T8OgKrdZxdGeTBlko6IPM+/tHt0rwe5dqSYvylhTqcQW+kTMZrJoWz/
MpgoeW7DVjx1AFBR8mLNB9nGNIDJFcQlW3iM5R6fB0uBtWEVXTRbghzCHEe5lt05HoRsckubqjGa
aYNWzpHY0eCD29o8aXo4p5M+SX38izy9sVcXz2gP9/q7eaauFxUp887orc92j7mtrczwVvNvLsuP
HeDSAb9RWt0GS6mjUa5f1EGE2IYVGG6e9OwF15bUbPZwnOvJsmEoQhVjSMU0ydZuGGDuc57jzSRt
jwY+xnWiksercNCVTC7QIFlxwv4cJPs8OzjgMsZJ4MnuSY/bLoy2KCThTNpxGHgK7XJ4yNZnl7mN
uKExIZtyZ++G4qZPYjq0aFjR9TCiTVYqkMozZQH53a/KJ0TfRHyxR/cVLzAYnMkBgAtE+9PpFM0o
7+LgDxHNm/orBI4g2m1F7FYPlrsTUJvvZMv/BFzuDzkblF+yn6a0tQVCXNEoLDk9/VuXEELtcfuX
OLCDYQMbGJUVIZRF7t2vE8MHc50rWgdNNsRrrpL8DCG6Kh5w+k/mtTwlkv83scw9FsuV/FdJhWnG
ByRkMC0qlEX6tZgiYTjLCoQEB5uXxeST9kNlfKF7/TujTUA5ReALc+l8V39hEogbf3EuKnXAvMLL
8olqKvXP6UD6z7xKGA9xIIYa7FTg8TyM7iEUb/HhdRuYWCz8W2uNusy4oGk0EuZHcGvkqSvebOON
IbJrA279MITh9x+oJafD+BGb32gELQEyf8a45j/mmMvpeYStNhV+utaSWIbCdCFNlI7Xx6Sc6cOi
Ol72jwQNwpzRSIvP/d9lQT+i3VU+CCvpDuMQGO4gw6JBb/Ib5MlAm1r8DppVqT64QA0O+BafTFkN
2c8NTgXsKnThnMTJM+vqndwhK651bf2tIfuPW4k5mxKfFV1fuE3i3IOu8wbJ5INSS/588jYoKtCN
dbXfXcYU4M6SNVIqUtuZesImzHQ0Y4ljvGToM9LhLvRHRSDACkWCFyehA/9cm7kakMI+C2BoQRoo
V48kmtFJvStSAiI1vYm6Ij9HTxCHK3bWOifeWSG9IlSF0ASUK9uuh65GomxMGtLUDbW6IJ99gOin
T1y193CHtCDdqhpK8S19cBvi8Dk8k4imrAesf/0Xgt9RsKAnpcixe519Q/31fWVo+zmmnPG8AplP
TMlFiY2NCR+jIFvTLI588pGnO18PF1Vat/t8Rr0Q78vNJ6G5QIxsejV5yIx59skozQMTNCozAONx
yAsrCqPBZg+jKQ7mX3Y/QHGLE5qZVLUYwCtR7HHaxv1LjM6xuzPuIwhbe6VcpkkVmBPLMpC3PK6a
plJy44Z6/WX5TuSEV6nst2+POmYgtbhd4g4Gkp2N5dTsllFDuR1rsvwnIjfXpHvVua8T+I30uCC7
dQateEo6YWPUrpACqXXf1PWTplge9U7erXznKSeSx6KZ3T9JVCEqIvkAx1ornQEnkZ6EKvxJiQij
2XbjeDwmWBWFTNeMKHzUJBgUc8AcxVRiHiJdeCJjKNxEig6ByO+BpUCkPv+3KLodXfB1DbONCsQn
W3qp7JYSbSIEe5jZhciVxr4hXbGJuAuEY/Rd/fX2AFNsi/ZmyqbzXgA/LkIgzZFJdA0TheO/pDwi
PhZov4BlLugX4ImvyrvGHb7b89xlTnqoJNBwFHfKTgYCVbTiOz382l+262oCU/9FVeS6SO0GQAPp
P/V+eQ29EAkj05ZaQICj9USZJer6MsXFgbi5ZT/3A8CpqCHoHaS2ilDDPjXLcQnHTy0WFPGa3fPA
QDdca+GbUYMaNXrJ8vnN14Yg79ZQwSr2HVJ9nL6zT+62VtFGJmnudq6zExt5gJRTIW0T/gkrNye7
XRa8NSWrfXjdGFS03qSQLQak4ggK667/U1dt0QLg0zVwIzGLR8dRrVCErFTViZL6wg5TX+cmd/SU
ucYMG5/BqW+n0QO16z3JPoXr1gAp16VaZ7PKW3P5ksgpvhv59wj+2lY4Zv7o6GF1bVSy5jbeNjed
DTZ4h9a4c8fdxbsiDpiTTht6W3nYDDrBina0q3IY1KEUTAaUUUXs6uGGDRKNw8BnvXm7NUMnhBfx
wwkSyKGjRGOh9RacfyOVu6BUegbjeK79+tzS2x9CM64Bv0ytfEDdiEOjY5Z87WUW0xXjID14FwKG
XW9MTtYFKQvkH1Egek9qjY0djuqhyS6JF3VG1IAjzgXHtnIQZN7Bdnj7aMIwbovRB/OyveLwxsvj
CTu5OzquMEoR/Fa124DtnWEzYk52YmznvPTsr+PUbnsK8EwLs8fScEH1AJMn2TQAWdgwZC8opx01
tFHtaf4Feky4qm2PveGPS3971jOn+g/bSgg3u3b06ilbqsb4ERIXBDOi0qsC2M6X/Z7HmeXMtU+f
h0t71aH4QfsRDX7UhcbsesdAjjSAXp30Z8vmtHUPt1ZanRHMMS6dK8BNkCwgpI5Nc6rsPi4uE0SE
R+nu6tMK5YZxpjjAwACWAD48MAeORGuypIRvfbtl3GDUjBO+/qB79XQjzOakkj7hDVAm/j/JbdS+
3RxAiRfal4l+MMM7U4eZ+SXo2geKSmZY/j1zXVSdL4Tog6gSXbAv/pU3Vss9ae14l2NEqUpWg4Ig
+jw/FJzRBsv2nFp4GvjRSBqIo4fAofVowSxffK2LztR8dt0HWF7L/vU5V3gFlbfzCvhzevF8bNlt
4HstJCfUWektNxAZmfDCcf/6Fb5TK7tVz3A5I53Xr8PIvqh+BfhvRrvyE988Tw3BEgQZtzRMBzUs
OHqeCco+wmBDBIwESriogH7AJZ6if6EZmP3dTVnPcYVYbr6pViUKhU0xuA0Nn3L5LdBzf8gQVf/o
uFbnwEnejt/YcqvUcKn3Fm7wlAx5PV75jG47ZWtKVYmc8r6sCENpqYNVDs2SiPk5E1/tRXgl5/eO
ukoi+N9H8fFeYROfNDo3yD8wPIlr/oQCuUleRjwFq29H084G/nXgHV6FSoWVNJIqG5YG1FxIrU9l
sd3YDj8UrEhuhfMatMAx/ayT8a9w2bnBSz+s6DXA/rHPZtcjNw/vktGROJ7/xAkUAfG2X2Bp2HYx
8oGE9yO9Ckb4Taz6FLts0J99S1m3XUaNB5HcVlVVqPga2iyRLnL1n3eOLRfsd03wA/KWWQl1TWX0
Yuts6sOVDAvpFhNFtOJegz9WlUbphqycrM+LxUUSdMW+YRuRlqVQrdI3UfqID9dmZlpciJf4I3PU
/41vqr2yzugRTkiCT0T7H66QEFtOpi5Ivh8YDWfUOotKiHj7f88PRjWWnmHDCkRX8C3gTRKTffTA
Z9r0x1WwNBCU9w67aTYy14iDO5J+xF3A61rDUcUjtXSVMtbLQ8Ex7V3NchcbsGfGqfDskXYFWMHB
NN1lP+TviBcaPzzV4uoGJZGqQ7YGOILuIiKN5WBsfyoiozOotVVACFfNKtY/QZV3q2G7x+mrwJ5l
IdtxyH/qJxz6UPrl6kkf5vJ+VnuZJfaP99zvEdV2Kxbt5YwxZEk/wFR0XeM3F5QOFk60JKw+Q6aB
pLrqTFHS3NehL0OYv+mGEgGOleeRTTlkUX3aYb/T+dMex6X/SxUkuYqhws0N1rR1lUhdn9JjO529
bTDtp4Fvz1RsS5V9PLZxOOuYBBPBh5xxOhkaJu5w0PRKj/clwF5Wsh6ecURXLk/vZdR7MqufoC90
OP1n2/ckZmgxNv3NK5TdFbTr5RoZbsnXRHgyCB2F7z0s18hD0TBFf0zUV+/BvfXwo5c2yKbgEIBg
9xdi8Fn46X271afG7V/3rp1EdCRlC3ScvyDevEA0+0rz1hIGIgVMiItnqZNEJs1gXzf2TwF9wajo
7H55mnxWYztoRDXaVKHbFRCPxyI8D1Boq8otmZwdHV5XO96BsWyOtDgxW2/47xWUdMxUuTTk8xjB
56S33oDHWPmQRtqngqzjIVEW+XWIctimFVNglTgIzSfsaPf6tAkPQLyErqedpczp2O9AV7Z7Fgt+
pYQN8mx9pBDgFubiztYj5H4q8/3m23LK4uO8m1nZ7lRYFlwzVDM3lsDoctO+LQxulIRGNcno4vZJ
nD89V7xY8CNPByVkYAro9xUI6F9ZbmU9GykMLc+/GWITUjxbeE0ViMmLEoeQawfgvbBVcx7AAqtG
6DeWXgMrz7li2ye49J4KoU0nfPQg0EDV9FG4J4xKbP55XJlaA9PdPYjj4jLQtUdeR4mSQxZn/iBc
jd2K6uTWh9NWnhsCrRDtq11SWG2TPT5Ab2UVwFdT61xNjYk7xLpyh1Cyj5mUqsQP0bwKw9Nj2uY3
xV+dU+cpKLdRn7PycvlcYNK5BptTTcjAUwMWxiD9+OlorwNXsHzKXQYhVhA/9p3753BvXYPk/g/C
pjSb1g9yC5Is1rYzvy0u4li2Xj+9zSO6NkL1mClTBy+/ra8Coua4MG6o+n8rx9zuANlhvJgbXxBp
YU0QKHpoH7TJJ1cqy3ei1Ftffus1q19qsAONvH8GmE4V8VtEV1UCzMS1r0fyBvdvJ/2gJHtmTuX6
81GcYzHXirIrLWX37DzfvH4yEjjBq8MIjLaEB0bkYn1ZQsUXYY8FDqJdReJzeJDCBgBG5UgV+CAP
q1eOkRJ8Js68og+TRzIJCzNlHIT9KR+2F4FJQ+vqy7jW5iPsb+0Q2RAsnHx6aRNSHgL3sEuHCXvC
BLV/lRehdeWjpSRcsIvrxnicEfSklysVZrdpCtOHEDlXPkp4eOzFdggEwQ+GxAM5xh839vruWuzQ
CHia1k20S0cJIf14r+ZyFpsLWqDumX9sG9ncoD7JRZsG+j647FHUNQflEr3Gx5NA5c7YF2FYUf90
u5KjeHGUlaROXYHFzM5xFNDaFqElUVz1nnmNfgyO5opryjX8E1v4O7O4byN5q2FNwzpQh3dhhMZg
dGrBQckQ78LeFnxw8GuHxJm2eiKYuHVHlh3icYhliz4Vpgp+vIdkkFLw+YfHXZ/jbvD88UTtETM0
MnYUptdlB0fbct+ua1xEe4MyIAhwhrZM9z4dzLhEfNA0mPuxaHXqCyjdBFZv02VQPECQXWCGiX3o
Aaes5mCR0iK8Q+K1s5gvIZNJwDI5ai0D45gm6uWXXzV6j+3Lgh5esFnUSka8qtqLGumPwVBlx5ra
2Hxr4qSuiculeqR7kYjyApS4qu6XZLheQwr5WVaDJMsKpDC7FJ9wbxdOAxOJzoSfBS4E37YfxPSy
q4yFcMxN2mhrKYQChFtzVLrfpm0hRT46+ixM3XANKSfAWpAqbXE0l2fdXRvczIRgZJVrepFyH4Fy
q9mG7ILvb3wNIrCDvaizZuYOJquiZj6b2CPIJQ20xYm3FrxHPirWXUZ86EvxQZUJe6FVoq+8qOe4
Exbt7mSbSdAoYTl1px3gu4eiRVkuNLpNDrosEWlqBw4S+20Q6tP6MaPoHzKbI6K3mUzK+vwP3Kew
oFLBTW+P4AwguKJUPCDHFP/x/y3Q74A/NNEDQ+Z/BsU4jQmL2Trz9mdWXiXp9JSXtJKv9GduItgg
yW2j31Ny9OAAsJ8LHaG40J15i1Oo+yHbEZ2crOxHROdCoWlnhv6+6Zx5LGWxlloAjXiwSRqb0Ti1
H1S0Lvyh9hwcv4Al+WYfXF1xHC+TyWptJ+5LtZypo+LYKS2JLpkivoUvWX+BZeNxDcydClasn49A
sEU92PDUY4qhX+6V7NtajkglAY9BDT7WByvKv+zAh8Qc0Ed4XKZqewrt3hl/StjnR8Tx40uIs7YP
iJ56vt8rZrMq56+bI0km95V4Xv6ArnmxyUqSm/qqyCn3EhSSt1j948EmV4zsv5HOPHOTdayI3nlq
tzpcKnl/HMEXZfeNddhvaSc4fGT2XUOS31geuBgx46S3QkoLTbaOdZE6htEUXczznkxfkAVKAEgc
Sxc05tw8Xrx5b5xE6VeaYH0GlMvWcvGgRCSWeQQTBhGkF3O94mktkZ71mXpUijZgWz3AdvHxMcWR
YccY/L8iFRZi2zbgo2OBBl1f7UB/1QiMhad/mO13rGLtD7t9p7UzB2NZ4GMXykUHhXT4YxHdYNmf
RXPaisQCo3+Lisgi3D8E1W+W2eQp6UiXTh+Q6WmMOcH9+AeHUKz7Z1YIKKt9/pqGYs8zL5oTJ7Bd
O6/36qPfDILDmekAtZZ483KHIJl0pLnt9LYpqZwPPU23y+6cbuxXcH467NMODR5jaogUV5TYnxM7
tiVWWtytIW8G6hqEvntexm3aMKKDDmKTo80qm3Uqa1lUmaT0rKgQb0iUSs2SSyjYQ5YkR5wPHsQS
j65xN+HPIkGrfjVlXdFZlo3M4q7Gna3GShOlPLEuewMuo777ZQqaftMT2AoLGvAY9yW81XeGmfKf
N+IqckskJV1RmEIpaJAqFrbtzs84GysI/r5wXgEA3t+URkxGzy8vKEYZgH8DcoU3vAHNK4qT/sZ8
tm6earboyoWaziVBheOLcchD9Nnsv9HVrgaasybvDue+Jivd72CvlgUl3LHpjjkBYs89oGgw06Uy
Pw6W5WGV/0lOsvgLFSvHZ1StBTRVHul4xjR9O7+cb8tmvMMa7d24astadUwdSiWq6aNXXB7/EM8E
W0O4iG+sVL2cByAL0xdZqZdQbsxM4lzjCpDGmcHbHH/5GIbjmd2JTxfxT9+JUcBTxBGFDCIWRjJM
dQxmKX5986zPbeb7uYYWNwi4ogaOumJhCOjlcgxVk5hSO87blEU3lqcCKDqX+PEMAe/3Kox3mFpu
WWSAOrSU0a0FcJuzSEMLaS0CJDuKutwKWtEQOmjapzYBybgryQE7aNNabTelFPVFgJYU9Qvor85T
jYbKoF3sy7bZc82TxryPf9BS8p+C2d0i1S+DLzr52htwtSI9VzfLFaMDncCil2OhBI5Ffg5E2M+t
SFLgD6pSQBdafIZCeyr7OZHBCwJSNGpkopRVlYImdfshUGOw7KyWG6p6wwaf7pY8YcL/8B1MZ7OL
upyvA+cC1vQpt/YF9LLoqF9N4ykzZMd+zBxnoIiTFN1ARwqicZWkWC1o6ypcXvi0tTC95VGw+i0a
krclvdOxGFBT0EjOlp/7kIEHcX7FmCOQ719ibyPF5JxORP2WLbnqXTVyRICOUurvdSkfEqCq2qRG
tg3tDZ9NgQOMObApMHvcRY5ILBAI9OZpQbcKoteUP44LZE4Yt3/C1QaEXcIS2Lb8hGmwl9Kbsi2j
vsWKKqQo1tpxyu5z61eRkXRW1TNjdakfGU360m5OfZbUSBGyunLt5qAAZ9Roh9Y12JxqQG1xVTja
RB89XWr9dd3RkesLnI/paa2iKM9qbKfzHRvIe5Pk/DXwJsoNOyxmoC+5qjW4eC0l/zb2t9XnQbvi
bO92ofOtxoyceWjg+CsXo/iv50/afJI/SI+rBSErdxynzIf4/heF9ZtILovn9ovCtyX5pJw8WteS
0sKHLuqjgjM0jL+NV2NTd+o3QU+Z8bXeSgzHeXRaXn9PqBtr9M9TMJfpZBvHkeKhmhdm7sU3UV9W
VgkZSOmNWmz/nQrrQSTGZqzuzUlDD9pQyA/eOiXZ4h0PfemBx7RgtuaOAYDNZNIY73LLCIygsjdk
Os5xRGNpH5moQlGqFlfZRCNhC+5JL8V5IiXrH0gQF4nstEWXRPQKrnvB0SdEbxkok68GAydHxG7p
42U9W9rHsaL6bvttm97ew+nhE77UhkQeG9/WzQ5pJ/AxKjhG1xeJsKzSNDDkM9HXUU/k9A+LL0hM
ZN97hP62y3CDmkJsiYBMVpr1tZYU91c16JZqyF0JzsWktJcLo9LazUHcY8u+e+VbqfksSq7XBbxs
oRtKOvmX/tnFVU9GX3fFz5zxP7S1ebvIqsZSiONV1sn7IHbj9itEVd8IAVmh5nGn2FntZIfOOaqu
kXKeX2EFaEUx4RA+K6uoqp+v6gVHGRhMsP5JYoOkIHA8TNIFGH8jXXJXeUlDAc1OAVduVt3iTefY
at3YhNjHsHNy2btuIEINFwzMkw6W0h1uV0tsxXiYKT8VOX2on+yOiN8x1quoq0JBt/f86gGLSjP2
SA5vBLIzzfSr2ofyX2zfykfUcw6HvYEZYddAoLez5YpsNscDzChPuTuAn5Wyxo5IQGNO6MaiB0ft
XMctYD8ALZRv5tWHBuFFtkvtkQ0eRW0fEqm0+8ovCr/qcQ95IvC7bbX8Oulu8qLmC4gACwrh2L1n
L686wpo8ObzmPpcLrFmD3/6mSeCE7oKPpGnW9JA/K/rVzpr1SbJb/UciejanvhCw1M4puQFqQf2q
VdAMfhuhOaJOCMvPBF/BRxHk4iKQOODLpCDK8GhsoDcaqx4A62R0avdkM1B1lOKlOhQEB2Z+7RZt
02rjZpIf1yZCysnx2u72iCnHmfwOadyChkqjW20RNxfBBrtvMB2bP+fn0HRRMtx8WrLDXi3a+XFe
+QzdV8ioQXhdbvpiiIPK1xIjLMv9Dakz9Xa5Njv5A5vW30hc35AmHxwTJJUpK0vwDGLZ6wOZ+yr+
lyWNjgv+q0bwbp418eqOVrtg3+b+Qxqd3K/a8PwLEWF3AzcsZbYb0sLSwvHDIAS+5m7ZmYQ6jyzg
wPNR431y/rqsi2jAF26koNhYh2I1S/gccBOdScHDj3l/BmIQWHMj0pGMgrhRNg9NU4sqSsVUJb8Q
6KLPnXOfMqYm8C6h4rf1/rYz3ywbcLTWcXaPaMu2tHiK9EIFcYZ7sDm6TcXC9sqAdNGuFMg6wgZF
WjHYhhESYzhUeUgqn7I2wEaZWJrJSr7paQ9SRY+ce9+XqG5AsbEs2VjVA1mM6H3SAjUFvc1P27lu
pfhrDypQvdoU/jDgd+fOS217SPC8pIivA6W9CWBPqrT/zLQiV8tQijonmEn7b0k7ccGGmQovaMHa
WUpGSPDuhxCvu0sTcS+TXgfJmGbX8Y/M/qBno66B/NftEjISVBAlQGOp6Yh0fRcxFd3Frlv1uhNu
OU/j/oKxhdAAa92uXi/KDHkp1pwH5E1hT5fq9znZ6O0w45vrXQ2MyjwAgScS78kJuYDYnBsUZU9c
MgsmtfuEHNz/IlgjTxbsClby4d/e389NrGZC47huoyhx/hBOPJ22ORaJAaZeT+eON4RhEab0Fl9i
bmyAX6T8jjiwYBFLsLZ1k8hvdnmyOHX2MZRT8uPVXcCNKgvRuMhQ6y8EPNQ1cM2r9o471JPI44Q8
SRBE+IQ4QUNlhh/TOsy1JGf++Kcw83XB5i6gqeSnjwTdzIUR8DF5snvvXffQF6yLUynxdIXCnZO6
Q+1SeciG1Tlg8umcJ7K9xTz9mT1INAC116NQBdIQIupavGPjVHfgCcGO+t7Ze++tCFZ1GiJ6s8Vu
634A2/D9Qd91vnudrODnG6pMLk4Dxn1sQW60WTMRTvAhCStqRFUXRV903i+5cT5FYRK7S/MHv01t
Nyrh8H0dO79s9zvaK0mDEpvNdjIAqDs5R1r80MCURMUMl6x85EH+8LQYdnR8qSCWUcEpMcSJMDQ/
lJii7ZvZ9S1SRE5zWoXUU4kt3PmaFzvZODyTMLOMWX5Y1EhFQR0s17jWyPNTMe44wcQg89xvqYfE
0TEkcg/WQILImhfTY/f4nhoD784LyZBlXObYjMLhbdP9cnNnyH/1XKWwshZweUWvoLCDQycrGoOu
8cfArdkXenDPZv6JQZ9mX/7A6q+kFvFQUtB0Sms98gK3FuatU+Yt/StmNgAX1osKdzwrjQEHBwI9
u0UZTDdPYmqF6TqTY5UdYFQDVF+IiWth+Cc+FFEKIFvb9W8XwtUrtxwyE6P3nAiwO6sPN3FBLWAk
/932WYOXNQhOQ0LDvt+EkkDIgseOj0ga5bb78hWwzDH8AsVeYGriZWU2Z3wECpU0aqYtzC86NomR
CVzJsn+0YhSTxklHLTEFIzdqIBA1KfNKz8azSQtlETRsdg/jb/rvMMU0mIWtLZfPzjjkGW5n2kjc
j25nO0NfmeZakr+3M0oN+CORpwz9KotcGCXajRfGDknhzr/34Ww6nf+n4rpq++QOlxHAzBvP/x+x
TALxRp8Svhm2i5moAURKyrYQYK4OtsmX5jqBXGBO9tB72LpxVvXyYSu099ogCSQDY7mTJYmNo5t7
3xsoxgvG9+KkLwbljVcL4UAmmK2byNQDh/Cx2oOE7/LPlz80bRkK1p2V1RlTIAzLTeQDkUhoMMTB
hzdGD9f1IEBWHcecSDOeu6zSCeOnIbCEpCCFxzuXXiH3ggteZLzufY26YngTH0w0I6F3wHCNe+kP
DcIv2b7it6xVMYT0mo44RSefSbxC8KZrjfKtPuxk3AquKq8EEGO1sVGaj/RfeG7mGNsF5MKM/W8q
C5HbwmEShZiBJUfHEQUYjWvB7808Zv5k0SUTNso0sZ6pE6lm2kZ12AAgsYts89mo6lsCvhHEH/eu
BRt+S4ixdoB/0JWYT2Mtkd7sRxYiMxNNL398WgPh6xEVJOS3BuZxFaOIX5LbcMNd1FVn6XTJq8LN
tw3lpI58UuUSbHYaa79SJWBb1IaPLvIOLtG1ucuHcUL/aBUHnYHaE3S9w80U2O0JlRgJ6lsW4Xp9
TXzJldZaqOirr+nCUjaMNtLs2/NSxwWTanDmNtE8UYJWH5+zRDbur3mMUssNWAApOEr5QdtGIlfW
NBkottjPQbC8pRjl4MTO+bU2tsA5bW6taMqFm/3L4wfAHPobK9Ft0j/E+rPBOLVDwR/fxA0C95RL
kN8plfQT/T+SHMJSOdw6rQZEuLtDhS19wDvTeqDTmT+XQwPdDnT09aAjQK5B5/OnQA/TQNfU62lg
/8uFTTeaqIug3mdqqnBB5muEHLBVXf3YfFLYgfXOgAviJxN6JzAISyignc8t8NkG/8aVzGsifYSE
ZItsjygNKhio2863WTSn3mQ0/lKqku+Pm1QN0DpQURSIKeijwEbHFY0hseRII5b+ANhNCZU6wcnA
In7YQTXtNM08ytw0TZpV8wmbTE0kBN5DkYKAfzUYVc4AZzj28qXepb0JU0B9nPsXlX+K3zPr8rbt
Dy/oHlfEP7sfa5WtAaMXlpidAvB87rjCALOTvTLLM6DaBvZhE08lOgb8abzKJR/LFi4M6EZ3DBGx
PDosAJs7B5TSW6WbPVebmxYD4UvpCRusc4g4P7Qr9tpWSgyRTZPB2cUc9RK/BG2ZgDt7w2cwaO97
C3ivSHvwXye3b1itfcYlBll+8ZG9//3dBt3bHPMIuJtZZkyeDAqOTyoQwUkSaSpWiUfpFS41R0nq
PT9qJdmfCYiBvO8nZBgUGwhwESDjK74sIlQGIqB58CTXnOiigXCH71B76d9YmT+IvYMstt+Q92Xx
Oi7ltWTPdKbzUQEqTDCUA/vAI+9cm+L5Duew4nk7NoLLFhRiq5RMIStq9t3WklktyGj9oYwi3JDu
feCj2qXyPhjyQOscXWO23ac6P4DEv3u3mlEG4D8vbmqWbLb6svZlFOSkBM/CfjqbX7s8nn3gCK/G
aF4+LKD2SsjEIRG11KHS5mRg/D+KSBOOyjT4YC2ClREw/CvXbPGnBztn/Pt2F/8ghVzi/v9lZwBe
Vqcvots0DHpyDdBcIsZdM5eFDcbhJxTVYvwDApJUBXQF9ahk/2Z/EtVntImzxnJbGAkU8KWlwrOD
cAEmiDjQbXeZuR8sOr1aF7jrf6jpLf72bpG+bE/A3Ump5Btw20caVVD0+Pl4R5fQ4l7rPH9uqJ8g
iYWiGwUU24pvVrbSDv8Xn8OqIHLYIYmOChYgTr6PLFLVG4X1MOeqBUkjofvIFF0rlWcVy6DF0Qgs
rfkGOYQVAt2T65y8PrfAlmtVu4ZmUzhzYM3ylCauMIXAdKzlh+B4bmaL4X2dy5jyqLQtXo+NBG3g
qfK4AMZyJ2+JukO3ZaBGxoGvZ9WLZg/RYZS2nG4G30CGZTolX4jjkTyvk6xwSElLZp/89fxrghAo
wGcfrw72kdPLRA2sLNVSwDvsSn1/M+1AN8czXFqpQUvIPGpQ/+55bzj1hydJcyQyTul7sdUGDcRw
GRNgZwVWq63p1SIV43jXwFEvI0WzBJVxP0nQ+cCBZUzXw8D/+1v5YyrBOZwqASAQN3O0SrTDQIZY
UGORgG1aGblU/LmcfSnC0ofCQ/cla+iR8oenev4PO5MYqfj1KQ3I9vGIlR845EyeV1GG+LWrPslo
1Rvp46M9OVo6i6ruNS//cRHSSSeYXLVUeRgBOkRfky/3Nh5d2Pe9FUFEMiItt5D748poxQnYTy6l
M8NRWey9npPk4MwzkPocyP2SIV3jN7S/zC3B3XpsTa+slJBId00WABqea0x3DsGayYifp6d3kaGo
7xkamFdDdkAf41e6z/LveEW0MazBQGyLR7qVWFec3JRzAphC+v3SKKnsA7HvjNt5/y4r9pG7s0Or
qfa1qlRS+kSR0EbdASlOsronMP5CtjyN/cR4a1tyX/Hqm3BsDyUjLG987ESNG5dfpwr2lCacb9md
iDeHgL+f7Ab/gTvLCR2+9Ndv+/y7EbTGITQacQEMXjasTF/wvkuCSnqMyXcCRVOeX30Bl3vuBcgL
62070J+iB9Ev605ABkhQAMV3utw0QfKKvTkqPou19lr4E8YK6d6ruHPnKGL9bA3NA9XHZVKnqERr
BKoh92+tUtohkppvkq65tGFqYMCsDI0CdwonLA0diDT8v/ttBDnp/kJeMBh5pTsBSIbb+4cTqq0g
/v0wpoplOE+/gLWoSnbrMqgrtsvnmR8jh4DG7OUt/3Gu83//+cUYJH6hZ5KZKVOpXRzP4dIiEhKp
3SGTx9LpJPlsmWOOLnjWdyfVo2iGdoVzPbq+J3cX4NvhBYp4DTWYgttPotDpPkf03/IfMnqRAcIi
vqROQksWQbLJ4GYa/qdJ2wpYabQ/bE7qMTNQ8zOk7OH1sx6q3R1vGUB2kcaI/RAy/F5BMFOpgF7a
9w2EyUTNeDT6Zuamlma17ER+xXXGzVHuCiBzzoBfFGCXXcKys9I6L18qgDpVkvLbJH1+zhD4enju
LDYlEmzlqrCPEvf4KVyoGtBkMdfvKreVHUUhoWYhkSVMt8rfRobN2JDLdxtIJxOrGo0PyQc87I+z
KKTkFvLGipdvCgixxHzpALsYs2DQLVGXucaCdDGnHSvagR2VmTn/+b1+cDTQXm8qMlQZNPq4qzT5
YJLNaGCtm5uz0lGsA6ptALQIjroeJVdR4YHhXMt1mjoJqyjJGRbKjrVowCBYJeC1iCSGFvZNu56F
w5t37lKMXp1bC/oR8LvyfThdL6+JAV6kUGFSbDIDazIbt1L4rXENGi21dIjJSoRGi6qZ4n7Zv9O0
6GRqfrt6vzU8GWYbb56Ten0hQkzZUDa5qgOeMPQPaOC5VJ3AHoIr1pCJGnlm0je7i96mmxlFv46s
TafROZAcy7853AdgnVRgt0j3mkwkwP7WchAp0UYbvi5V1s2U57T8IN3eCDsHzPZLeTXsi4ePmCq3
wtV76pH2sJWWuMzP/O3jb5ghE4+Xx7HYutei9sodfapTa53WHQZB+lp72H56OrQSzHRjHH+Ce+D9
93HF0c5MTrTfuSCPbWEd2p9hw6K90zmZcJ2uh3bGYt6pDHq+yShT+IjA6FfC5auy+A0hTSFMVCvx
OAabcyaHmBY+YjHxpukVITBgZ8iTbWEPbD9nc6bAggGMIjouF48x6V0keYVjcvG5TCjnCduq45tC
tXYRYztCDoVx9iATravKQYYEec3uVNPyWvGbl9Mfa0YgF7XIBhNTPqI4pgEHZvKzB20O14TFGbmq
rkAuLKGnWzHUDtzM8537bq6W/2phEVRX8CXNh5akaRWyViLG81UHCXKuzwOYk7UfnpfV28Pq36lk
SfSM6NEGYdlRkt8V7MEa7ZBkCEiHFHQg35YmFPCr6aMDXMi8QMxtTXlj7MbMyotpa8e4mQ0dT2WG
FuKc0n0YlWs8PNzF0+eYawgi8klfR1xiQCT0EUpoZouZUqfxaCGv92MbE7QcRqw9KFvnJNm0czJd
0QyTgjFVvMxNn2nmVSqnEHoTmbfb+CVgCiM+YIeSwz/v+kjg0rirXNubwCYAUVGBs6Baply2gsXU
Ftw5jUJvDvuYlgbr+DQV87Zozp87K+QypHRhWCw/V7FHDdatbLJUJXPqtrkYK1T0IQuH1HQzngAO
VK0EWyxRKy6gcMO+OLRTkU5rivSw+n/eTSD1i4PiN3SVzUnkm9fsdk9OwPQ7ikc3vT6ZzbEeHODU
CgwIdvjdNZstEVg3G+MJmZuE4vF6JGSVUjIWGGuODttkOtXkU94LLa67FZLwiQSJijszMV8/Cq9Q
u+7vD3wcm1MkJYtXg44zbB5k5AcUxlsMSefpGIHgus6fak6NBZFruhzM1FBZGkn6ZM2fbhc1wrBt
klcaYUlggRBBVhqTb/K5Ug1s0rcbgw5ur2ZPmwRhJbGupoG7X0qtsmohXqa5GDXUsbFlcQWRevll
8SLa5ReZvsns1Lsv3L2XN5gWbgaYnhKChNH33IBLmEJPfT/plqpVePVO0897AjUWSapoF+iEJDis
jjyqozxvH/hzS8epCIbJoKHZK6bdZXLE9rzKPLXKDqrMg9f0DYkWeRBeyEslePGOOJNoNxa79Wz1
P6yj60cvpELmddTG+ru2ARUsieiWYjw2VYqB07r0YAHQ9nk62HFbgGCNbgQSnfXbn8AqNztB/C+8
tmvL06nrcRdKMvETOilojXV6OVQyOVls86cpbxMNhvPPNpPLE7hohV0/8JzVSTpfTwz7000j5ntj
B0o5KlzHTsTCWmgIdiWSTQ6oWreCzJ6BqZbrYcwufGr6BOuPFntDhzKvjb3K+P3ITaKedw6cluZz
s7AAahosSXeg5BDCo4STWu4r8tR6VXNcTjxBWnqWenYwCaRbE/wHlj2myFx4SDHEu7wgMaEAG6rO
GJnCsVLu5MmAfH64CF3lGWPDrfjOIB9KZ5prezMCkq5Fpex0xu51rXbE4cBkxlnhU715WcPehIP9
6HVJ9Uhy+9T3AreiY86Jcb/eD7BOP+xCruhu8Bejm6ACCy0uSQk7mmJ3uWNbkbi7tBfA/tYflmpU
l+zP72hcg8ospL45XohTA4F0jDngeBbXsGEsvTVEG/nXb3KhnJtFvzXWfuhThHRy5v1rGJXqRHTt
eJPGS31e4wNqgwnFkJiwSGDlaLmuYZ8auYv7mBn8e+8wfpG0iQrD8X6oVY1ii9dOkFpz0h1l4pPf
zPJR9F1f9ab1jrPLvD5hFKGTDIdCxDdi5nT4YQm6IuUCxbJu1tCkNHcfctdvwMcwCF7yZ2ao8yk9
qwxXAO0H9Ql5WW5++8zBYJskcNewPd8k5OP7VKCUMknSK1Ll8m9RX5ftTTax9ox3n1vAMYkhz0mr
+4e9WFtnagnFYOO9CI/JAiffvaJ5u9t3SSmWPDz1tdlaAC+rIsYUIje+8E0Z5sO66v9u7uhmM7do
mawxVRilrHP+6nCStws2zBmhsWMduCT66SHHkdzbY95I/lwmoJ48UpAV2jvqSzPAmWlYY6u4fodB
UJulcCQDaHde2rncEOQ3yk8ayJebcEF5ADgINc4xdhMqRS8Kbi/030qb5tBn/9eZUB3StSiIaUgh
F6xUmhGVHyonFzuza5dm3MgsYN68vSexRnBPGOWCGu54/3F26mQNBtqAvPoZ68MTjatt6/HImvsT
PTaZnfcLfwjcQYK0yYvExvebQ5+kZ1NmoEq/TOpMhvckNzy5I5KSfEU2/W/VpoDmOtxjwRecVNE8
40+YziIYoTUqd6fPULHFGzZgtpuKTdyU87imaO5Fkz5lVeYvt/Wkk+BJ7+0z2TmbjewCJxjjbOro
bO/cDut26vTyVEfbwv9wHsJnDPlJTWhYmUwmfVAQK1tG8L/keoVS+Mo+gwaLj0Cd45pFqsdbf04t
WLcUwIKpg0zVoZfvNYoiFeOcYJM6s95jc2j1yNqc1/io6Qxb36WpugpKAAwgrQ95IwSfAR1k7+mF
Et4zCFYdFCAKEUczEFYplGklnRcDQQxrhpx9P29975K2nAgpbXwH2WMAg2821xUXkyFSaSOVGGI+
kSxN819c9cYuNVeIcO6DlmpmSXVBj6ufKli9ZgsDL8lXqBW9fGTi4AwjO7faUprTA3C7IaFDF9Qn
Va5yf778X9aHDvTyYPI/HYfs7zcltXx5zD0xLzdtNkxV44pcpNYghTrSETjmezXTLtOPS2F2q0Za
8ilo3MPFP7GvW3CfXG/Ucq4L/b6FJm4or3AvL3n2nvrwQCf9zW42akaRdo4x2PznzG+GRwxNxAA9
/fzSxHE27Tou7eMXhMmiw0aBLsOK4CV8uMlSDX8xs6vfVDjQ3/VD40h9z92Ikh/djdE+UBRNbrGT
hSGXI3cB3ioC0KMVU+MSxrYWEYSb8MCLOthDVrhVp1BtO0fSTsMpE8Dz42pmlzDLxooUa4QKqq6B
avUgrGknRI+3/IhyCmpkKsdBnP56PDZ5HIfsu96iZJi6lrQxhxZbkeZ0ZoCwr/okgAF+i36Whbck
RgkGDxorb5FPnBhi+jhyfSkPbDdBfFhoGHOobm6wqDn2v07RIB2y0AyNJJQaYAEoA56CWYOzgfYF
qJ/HYbrHaKv3ikCOIQJQ72/UzIublyK5jL1fY4QMpLEFJnyysRb2xL0V3ZqxbxZY0uggjSSZctxq
bFX2Dp0IGoHi4a1qfaaeRbmNGnSNG69DYDb7k2UwADM1yhEk/5Y8kLeFmCtCuiVcshZDGgkVZ/Us
lWD5EQpUwdXobEwDCHZvtkLsF7Ij15Hrqxq/HqssbBo+UTojeVmPbi3mL6bgWW6jtui04Uh85LUD
WATty0r8HeewfRr6eD80ElN8GSkUdNEJ03ANdDZaen99/HdCw29fpq1KS+Op2rsMnUT+QLbWt6BT
4fTu+TU7ofp0G1JVu8cL6QCWVWCZ2nGLZVFzLJgrMYWDyONEw1gg+Uwo3OjpI7QIuQpWbwIoVLUz
fa2JK1C2g+AmgQPKYKQ3XyGxQ5xryfK7dx8axpeWqkwa6oc+yQ8yiEdkx6zr7RCIbseohae7rWP2
cOyA23+TS+cjCjBr2eZQp9MEi+6mOGqSKQGWogqoPCKfu/VrShn/uTwLkNwsunlJForIrIIpD1qX
8rN1Oe0gQoUir3OI4jT9UMyI4wnyd83PQuqLWFzGtyiLXBat0UVyaX6XcLta4cWNkrP464q0EG/g
FMBrvrV6crEce6gz4aIijdjF/bzKe+WhgYku/G///vMPhqZdeDO8l6qmixkWaHFmvdGeITnfTFJJ
siEO9fQzENpAnJpr2RGmFRcNMKZ+QXCMdbtbdR5aufWnPNR1D0/M0lNWzAaI3p1sYAj4jpXwOJgH
NNYJFe9LzcmiWp0T1m7MRuSJhil0pmvX1SQbPx/Kn3N69tJlUjqjU11tr+yX3xkVO7qWXjckdkph
yhVrJNzcsTrc48sE475SS5E12SqkLL6EjAiyNHjsaGrpm5FyL7blUcSet7sXTnuUTql2le6lOlKv
xTq3Mlpxs8MxtIpIog9AwAVgBCI0lUwMtjD49gw27++1D8vLhOZ01qLmWf9gFujq6qv0aKZBquok
ryc/ZE8zTC6puHqTye5rO2Y92FR1dYoaaekMcrtTD3ley4jGiGARgKjmBaFtj9HEy/K1NPXIlwjf
9+4AqcW1hGFPKXB60ZTdMCzI2rJDtLHbSZXHGp8YR0pUZRj67HXZH3R1hPPOJUsQMXgHywd/DaoJ
xXD1OlGSGZahrveeHp59tpHaml5FaDCrDOGP5jO/Uz5fcv+O2u/6s7e126fjPtAwwgOJ+TXTQqiW
4RaKYCe4mWAVKdRR8Xh19BalEiDKF/DEJO8R3IZhE6tOZVQQrifj7JMcjkmxmeyNYH84dOm2FfJN
XoUNXHYoFBkNPyW7RkXKl3IdU+chzZG891Tegl40l347X6z6efnKiveeBM0JUlgF/Fwco//V6Y4M
M0091gLSHfSrY5pMfxLabPzZECE1ik8cBK10JaXVAn2HNx1VD1r5Thukif4SaYUPTqMIsHW0/e4n
+Di9wK47+Vs05C4kNRVsCNab/X+ZwGq4OkYbeRyNbGS9DmPk38x5wT5WkGW71jXePl688Zqx0wFq
RISOXLwG7IgQUzZwipWdknKOOPmBcDnJ8KKxHapjOWCa29JwXRdW5W4jHy6GVpBxVyOxBOVuONGw
KOIDeioUOfPg8BNsGmK12K8ioCFpr+cLx6qM+xF4NYIuGriJacWASvf6iptci0abJ5PqCGHiI+sd
a7XXeWlzZO9hexBDXYqKL1p8aOiCLURLhh8kNlrCYEovCzMSQZGyMNPM9VycLgSogL1MNQk7VVGV
wbleqCEEmshkOTs20xeZyjRojJoX+uL7qZJhWTVn0bE5x0GyiZW9qyM5kE7mxlEld/CpSixX9XKu
WrmybW3gUzdu5K9pZJgS8uKhJOEXrVeuhxqaXRB22rSYlp2woeoDarWiHvaZfWZgyrsAmwkBCGjW
p3aUx4IsYsd+SLGDEO45xuf5BQUevpzcImrTClV3Q8CHR/8/8McbxSMRiut9aidTNF1j81gNqZFf
VTuMmPLJHDk9jATcfXqkaax6jJSa73tNXpA3HeMyyebD8VN6uYciGwArS/Q0lFEPNvSQrHqy2Jc8
wmMdiChkNWD4EcC8Niip0tU79/+oIh8aFfHgu0eNd2JNoHmvgnTRurbNRtpqmdQk++3bvYIu49Rb
27233YefCVfhhHAoe56Bmqyl9ydXJdjMOVp3Pa0jVo31aftGu47e3sIyyU2R8v4cyjc8MVFfPyvB
NhQ/pYAyWPaH1BqHFOM7f87+9vI+5QxLF8ff4FotXTfKW2Fu035GwZbdKRqRs/ZtnrS9UqePYuET
DOxKFJcDVIW8sEgg1txt8ZpO3vvJ2KwFCBlrN57S4CGhE3kENr5e8tdPXo0rzKEvxNpIi7ukr/uS
Tmxku9x4gk+TuaTXe79E5dajoAwjiwkRUz4k5Ju+fCmjars7Gf0PfJdXtPeUbAPKzeQsbkuj01au
3OsFQqYNOWamvnhw2tsXPGZ3fyQWfwDSo6rx+SKO21n1JbGf2z4IaDLjNOFgEVKN8LTXgQBUfBUV
L93ZOUU/wVrC9s4yvlTfZySnvoOoIOYuOLTkHs8C5HkexQaARLDQIn21HZ75CRzXWHnbR+lZND6X
YLRZ4Dme3B+8+9QpOMinwKqlZPsujsFFPGV0dCmvdV01AvlPlqFtOPVFtfhuJCGlZ+6lHbgeBWOx
RdENE61XpPgemzEU8nbV4UqkL9nqWz8a2/Asst8svxiUn52PtIICajCckZ43+15GjuGu1xgBo3T8
hB16Bnh9Bib0L8Qj0GncDERZKyff8XBcQPLtlMda3SrBg8oO0Ovrp1ZHig8LEnkgYqOo/HeDVktf
+igKk8RdkCm19h+e0agvurwBdPQXL5e7Zs2AGbpHNSCj43NKmtBP8a48YrpZBPlH5K5gD45vKAJP
LdNra3OVGSzTnLAtdw0gOJnY6usRBz7hyizu2yryR5j1ByzaPJvu6IQmodnl1tPPWlG5lJ31Mhe5
U6rHGWialj0YXhD+IZWVSkcHZuOAeddqsMdtcex21M3WTxJzKnUTxPWzONoDI0sMEyNDKNlTYZaY
2UfA2bZeYO7jXkKh1RJE0xo/wP9zxir9Jw1O0q3XRncw/s8y7CR0gtxJSrN3xrs5zGS3zHeRUq/9
UXZXa6FB+ZPZ+3koeU+gl/nSheLTjo8d4m7CUJZ9KU8Lh9mjvku4bDdPvrZuSLEOrhaPyMsVsa9G
KDj/20vSwY+hWt906db3UdGfHUs3GRwSGXR5fJhtANQNtcIs6vDWyiBK0hdQafbLdPBTTVRM4NEN
Ky80rqrN8AKOrB8YvIv6sSkdB57VgtZQiDrsjsSyvoAQumie37o33cz2PpdwPsjwJ2aboGy4+rYw
RcoxcQVJPQbKGSvvlk8iRYDnouuFkn4SQa24um9IQHCJsQKjRca3QUKVrmhviCdZBEmPy2gJ3sgO
zrUf8UPkxswd4I4wUCEKrV0SZYM1+Kth8fXvIr/MS5HJOpwSVW1iDR608iHxx4/cBQ7F7Iggt3R0
NLAY2Or1/XJXmnssFs1e0EgWGAw847oM+F7Azl7JGmxlXbxTNWwfMEWDF2svi435YDQEk7e+tP+T
vnOoHA8NaIXS46MAL4zRSAHz4KL0YALEIx1HPOKfwc03uV8Wtph+ONcuvSGNUHhFXyEys/H/qpFq
VQtAZrexvgZfdUoyS4WhWw9x0L5Vco463KtbmwgLwKjOPrLb3DBgK9C/qgPRnM+crr1wNEzis9ef
oLutShUgJf6t4mvE775g6BGmqoUVMys6FYoLFUGIkoR8tmYTKVZU9KoeoOUXkdhIBRIdAl4oR6AK
IFLUVR2XXSGTBLvYjHIzhmGYmH/RqVUpddUwPjzx/0MSMWP4X4hWx/3xK1xw3rMg1ZeqrtkHZJtn
cHViIYirN533EkKjIAHXfd+8VBIxK9PwJKEkyHGrIdyaF5+077tivWtBtC/WTQVRPLo0qNPGWZX9
PU7d8Ief3z5ZjqkTcNL2yhkftv4MQXjL29bVtuOfEVTMx1K1hYhXpfuK17FOrR5qpRzFnF+k/3dA
zLvYwC8558zmso7Q+Iln0UMPXQXxr2SGrn2czIbDgsugLHB1omR7JWUb+H7A3YNA3X0o4VGkpRYU
BlOPcmy/M9O4qnZImBtkzIAbAvOZcrF3gQ4XTrcO2YZD4UwN0cLgv4klPmgJaCQ5297mE723IMWX
hyFHpQRZrrVJOsIpLJ6KcY9+Ly3YpP4Igw58JLNnUvINZFXtBdasgUKYe9OJXxECfdKMG4n2qZ9z
g67GlMZjXpvVSHYMsnjRpQswHPOiIVVxZ93Ev70ez1ZMbRhL0TOoeFT8Fo6qCBBbaQ8rskTa1s3U
+ta30ZmP+JTJFyfiFuGnKpaAu71f8WB5a3GamEi2OJ6E+VhuAyP/SDshBV28N6/Fkr1lhmVqLagf
0zPcP4vngkKrcgXPurk3nPa+83OpMbyM1et7uPwQRTurRVQEiNx2Pn0ZbJzdAdzloM2B7qyoBezF
2SCnb8HcCSpo0VzBbA5Fp+uaqaM/M+xLxeH3bfLHL/BVdnNtWEZTYq8o9QQjGqFJwenOtYWHyEPp
gGVVvLM1cTnv6tifN1BYRVWPngtVTnBIoXV4riGnDWBA//XSngkamZ7FAmhRf+zLcAbtpuTFTp4l
k6lSmj3xEmBnr7a788TXM2E+b3+vObVj3uPyTDOhqWtdj2bcLL8OgqNRr7ww1RgPftDuhp1JUgOa
f6CyJcu6edQArepufjUpntWrhKKtH9WQqefK5eXDOSyorKrFQ++dQ9SCfGOOo6zHA+6uRuS4nZEA
8TEgOdzNnZVaDCbGBnUn+0A4ye9P8JsFKa8D1/6QDxIf1A3p0YJjGbFr9RMhntZ3GJAD0Y5edy6J
T8dTMbdFx7k5fDpRDw01vGQ33WZnGK4X5eYVnm45UYPZBEoMj551qazQFXnySVny9D8kuiiAwy4q
ME30pSzafcRK+FQwMO1SrlcBmsXtg17x0K9sOCHPLYLTuj3iIHjy0ylLAlgkW7sOk1rxLCh2l4nY
8I0PkWe+daBeHiAnA4JIWWjS6ozOtUfY09o4/2tDWt7RimbEuhNYNfzttz/mcXEK7Sat3RWSUvPz
YlMr45CBC3gmxfQT1rygoLZSWGTLWzr3UzIzIZMOdK7PHRVd3OKLVsZvQtkV2Bh6Z/Ifkhg237yb
TMqbfjSZAyqj+M2gggDRQDOZS6P7kQYZgdAzedZsF/CVxpyzWaunJXsKmCC8QFAuXLRsBZ4sWBMe
9DHbC1Y8xQXXtUHTlMqVlzwd8GTdK+++HOcysu3dfk26l+qCzauFGg+gziEotEB/IjVzBMdew86/
9pPI9EXVmAHJNGwIxukfNGhQ7OCMzElW3cCiscklqh7u6lmt+s4psaK++SKMpQJeisxOpNxitllf
JHfmorfQE7N6vIxGvUXcgwSLjPXN1DNH3XEoxiPsF+pd5vQ+YClrXGcXxdZ8upsnOLvLaxB0BjCV
hzimO5YRHDkl+/zKlhNyG6HVTolso4B6g9+BRUEgOOeFN3aYSottBik27UvLD6luoAkn1FVdgUGT
IhpjXD2eC8mfAnIZEqM/QePL08VBYuVFcAD6FRG4In3J4hnodKXVIkwpyQEATcejmGA/DQ7Ohliv
Tk+mo/7LTv+LSbfiB9VwTVWW224FZGUf4U/aZlmerXmffnmw0l5JcI26EW/QcAQ3I9GQ92wfAN/Y
Q9tgSDgeAKMHScKhvm56CMTyi4Vmntm24FPjIDrFMPhXbgjVLVRIUDryIBz/H/HHgKjfMx2tRy9e
YWUq54n67hlzPApfSIOzSKLB60vavArm4sRWXrHckUR0CJDTdWpfySt8Z6MOfpGx0whmhsNevmM7
P1ifpLFCbuY7NVCRGWttzPZR+lXR+fcZS6PETL+sMZel3X9N08Q9U1GzgZWpIitkhZwvrPenGif8
kd9waPCwDSCj0A1Ci4vq2YqS3AM2K/Z5GLCJYunNmCDstLZ/L/h6Iv/v5BYKDhwJ9bD+45q02lQN
6nnR+jErpirxHIQpYJhCJrdFhU6U3Kdv6+Xq8hUqyGNeXe7amlEpx08wg4RrjnsXL8F6A4pReKU5
iGSR9sY2X13c1IOGC9oBGUBWfftoZx1K3PQvMy8Mc4Hg3fpF/sWgqBkDphiOdS+J7/DKZk2qUg5O
mhXxt45vVbgiIFjWpsHsqoMwgChcnB+pNmfztMIjyOiiBGbmcKIw+ak0gjmiCOXqeFgTQXQtPPm3
qFljKdYDlOxJQL/orNc3RjBBC3weriHZLG+Ss1jhYpLrA8cHhLsjxpY+IB5Jp23mZJfdc+Y927Td
eTGc+cI8951CSYG5NUiWEwsMP6n6B/lBTLXZO3HfWB7e1XCkg/ftkt2U0KbP4zC3eiLxZ+jB/Fuv
/H11RhAZ/64sUZZ8RUcp4x6VKX0nLi8emis8/lwaNwKJkmzehbMpIuU9RLDiDoDEt8brnGoBapF8
Wz1uUmLCm4Ajp+lh17L/ZnJAXTJklhay3fbw0VMZpYF09hjvMPe1qxUszUmwXCtXLWI0u+A5zD0G
cWEjpKgyuv4K+bEzF3mlolE6lQhfx5pUCthJi/XXIMJFO23ywQOabXgATstkvQn4xQCkDarlVfYd
B188INKAtjE2R2GMIvLuX4/l83tlYhpKpid7uyzUG+2XHfD3MYlYvCWMYA+sJIu1ESeAUo+Amc13
RG3NAtS+fNTCpecrx2rlQaI3D8otqA9jxop2GRIvnD6P19QfP6fkRWVg2FoTVQMqcIfLS0GD8iMu
3q9LINp1fZ1AgkhqdoiQ1iLUT7rBPOe1CfYUEgqHGgfdBsrXFHXQbEz1vmx6hzn2Nua5s6eiHPOz
OOdAwN2jgzx6ajkg4BlQS7A+nKKGthvsImHeHccWDpUKLptKWec7lCClCn/0L3RgfZX+XuZaUQtM
KtzsCmwScUYsYoLNj1i2UD5soQQx4842YKJiO0armi0HZovp3xLh89pFIBtntWNMe0QoqhOdGAFB
qHz1sgHaFm4lLJN78Wzdwhm2XukdEtCn1Flr3QR7KmQ8V+hQrfijhj8el46sn+zsAvxSOkJb6Stv
ARqYe0fla3ub+TL4olLhF6+mYdoU59UXlGaGyqYzo+W0j6QOC05AqRCFDZjbamkOfgOe2tVkxlRc
jtOt0AEAUoHQOpC098dR/35RU3e9MB3JMBCjN319AM+QoaenT1h65r0OIqFgsvz0vUdJqN5mlqQ+
ztysA13RFgCNVp1ETdRVm0I2FYIYWm1KDGA7EHDgaRQ+qNQiB3VU+H9PgkI4R6FLwGO2JFevSvKP
VoDM3Wp4phidl3v1OjalQ48HjbBRAkdcVFvzpIjolYQXBW9j1UXegutiTEpTUF5GyzU5HIchVHk/
Vus8Sv8vN91Oc7XC0FUiafs15OvoRaGPzYXjSVjZArbwq+pLsL2u8LXRgJtkVOvO616bI0RpSKVo
bB8zVCKwkFVoZiC6Wo4+DFy1ESBrRdBoly1Hncg17pAhpVqP6KT5M2jDx7+jrR2h1pJ2CFY0CMiY
06GagzCLVEyPtfn+sHIwy8Oo6VgvWhfv+EQHTNXU9GObMI0jKlM0k6gAEKxpXnGB8n0ecYObNBv6
9rzlaDKaLvBfPoUgF8SU7rLM60tl3nPObZMM3G574AUB02HhrKkaAditz8IJy4w1Hev0dznmeESc
mAG88UExpCL7jy7USyLpThp8AGVOUBeMfr9ITAw7auuufhlXShglTOBWoGjTouH1P0EoCHEW/AcT
lIspSmc23Tc/cwPsrQlOZgS7CGPiKUBuMfsWyTGZZe65LwWeV0ti5tBuzJT/LgxgQotlBcOFbWSW
wCreW7dmsj81+kv0pBG9dSg3Xd2CgDNW8w8j3G/wUi4rQLj780jhZs/5eCGrHHWaLFX3TrvM9TnQ
USe6rgyNIpYPS1k/NzKA7Funga5w3fjq2MhPBNIwrtO7l1ijfdJBfmaDATX5pCHtQGb4lqjMnqKE
4rYQ0Woi8OHkpum0vo++XiiY6dLnxXUe3USvJ1ccBPbf9KZnEJa5Enf4RkM+KObI6Ep4G5UsmXL6
QOIiuMZ1nh3uHWd4qXVZ4gCNsBCxXKXtclREil3jOi5p0GuF8xf7W+tCfjUCo/OuPYJhIb25aov9
mzfNReDNO/frARr9jOiQ/oAwWv8fKT+ToTDJdgnfeBC3k3YTFrtvYb924qG0gM9Dirpn0yaAoKMg
+93kN3Qj+iKzW62bi07liE0XpkiSlyy4sI33p7oejhKykUvEwpj7Z2xmdSjOqofDRmW6xCTIL3dp
ZGf/g4HGgJIp3dmUfcfLFcNFtzriUiDIZoflYbxFz6RHeXv+/0FOR4QHb7SVeb8kidWK3u9j4Cft
6AzzLBTetsyj7QnwJRLImVbnyCCty3puWfW9BWODcZaYOoXDF9hGoBhGmSWsvk6Kik7nwKNA/pNg
HoreGhOiJSiyRN4XD04xTaNeaxpvdWXX0Gi5tpIbDs7pkG5J6309e3w06FZ+Elf0sjCs50KjlC4M
id9w9CMPoqA/AkEUDxnEQsA8Y8mGbNx1vGx0n6djyPC1adDfbAaECWmIQhUop5qVhuqd6cIBMqbk
xYrXP3IrxkUtpZQc+nvkKcNQX1DSHbeSGBN0tswhX9gQ5WC+plnWtmyD97Axz1EfEUx5dXxKqxke
L8MEKFNs+a0k+JHpt3MxVsIB6qTcHVXu72DQRjNACN7y6Nspt/lXQ4+BhQHUW2nT9UP/OZIsc7px
e80JeuqJe2ImVytsL91l9SwpM08j3936x6LbyFkUEWDB4bqFuF2Q0+kcIiALS6gecnghdhoNidf8
sxqyq2p7X+YVSVihpAC7PA06XWKOI5Y8XURvjvtijBBbeAmMGKr2ynKK61h85+/FBGRkG7yqjwiV
lV+YT6b3BI5bivbwgQdcxMZPB7CETthhdHFbwkSlU/CiWoVdhaQPkQvC5s7Svux1OXamxv1lKvE2
Hrk9Curm8W8o4GPg9DuEwlo5MZNgqrDGABGaX7OOKWDUqru2M1eE1JGQZ78pQGh+WTng2qPQppV/
aHghAjJ3Sk/q6FTxHUTf1uu81dGNBP+0O1SMZLhHk89+Man4x7kcLvcu9c+vUe0uom2sJCcPsgaR
UFMDWNXAWCg8Qep4N3VePjazeAddb9kdK6ftydd7aOP8YyvVLXmYgjKKCvCFLIBrKIKv6zBmnLod
6a2KBwpI3f/sdth/YLm/Rt3zcTf112tghlo2l8Q3q1UR9o0qzyD3H2gx9dGbd0wDRioVtcIDQWnH
I1CBWEXy/dV0gjRIUVmM+aVT2/nGeX35EYCr+CxDj1gJK648jOmpfNDB9UOqVYpU850rpk2uYdX0
Ulm9uIuutXEChGJqc8lguaU/Jyzdl1tW4vfjp0/zadxfeuDaG6Nc9zmK5K1Z1EzOiizhyDRePLFf
zyfqKGZPzz2+mJofdccEgBc8jAOjwgwjNam8pT02VZb63Yix8LFRJn9AIj6OG7L8uxdiI4LPXmvY
4MGZtH2ulAJlB0ao86rg/d95+EUsRTfjVKC57hsu9awtllKZzslTr4GY24i3C+lOaf0dTgcGrKaT
909GUnWTCItzZQHP6EKMudTutSnqN1Q7HzqkaK0HQVrk3OhLyCMp0kioCXwSKWpphLrLMFOGlUy2
EjArsgk6Oud6BW/K8KxUWbJo+B4rtM/lis8sdpgAZiMCAYBDgtDTbOWrCjV5aWsLD6T3yo7pF8eo
GuyxXgd+N1CyXo6eWyMs4VT5ccEl4NHG4bxD8XTfd3uApwY+DtO66Lg94p4YfrILg+L2EIYx8nsI
IaLMJ4Evp+simreZWTASFf0j5PpdCDK1hovKadHtG4vE0WOz19EmxzuwyKnQKLUpZKphfUH6t4Bv
BGxcXNfE0mfbNY5jLcOlgY2s4IWyyluHPdJRGzcZZOBS+HpnLqTWiyYvGDNxR8Lcw+kW1lt2CRge
VEpAFhKH+lEZluCZwtNHOjIHRjUoQc3Y1Nrax33JyTnYtWBSMoXV6pptusaXYNEd+iZV3anG4IEE
UQLd0NNb+1RfcpE/7L7C9qA6Oo54MGGYDvLBytJ4Gh5qXc2V9he5OxssK7O5ktIN3XE5+ekLtuNb
TmqcZyYyZgb38ojq6oBUrmSezlL12BrBRG5R+iE8mVGvUoF+lam2eLNUWDcrZb33NziV74juaAnS
GAO/aBIbfOYwQYRumdCK9aHWL7TDQE7qgPdXQNgVT6Ujb5C+Y9GVAlnr7+dEAKc62iJCC+IfZrcx
sziBKxDLmY3/tML1oSh8oE83Ef7oez6aW8etGAFqevNj/ARRO42wx5qYxxLqWzk/8PphbqrlD3pQ
sagm2mjwGU5HrJJAXeXT9kYgPwrphpP3JSUwvf3OZxhB4/j0gZrF4hNBhTNCo7bzLTxvtWuzANXm
sW6ES3yB7mUbXzQe9kydFDB49ogFyxhTSSCyGmCDpNKqHdBpYTLHFAPNuBQI546cwryZmMnnknhF
12dsF5u6QBE42n01YrvK2MfI2GPvgOMIfGXPqL5Y+wsbsN8Dy2sU6maET4JdAAWgBGUS9kjNRSNV
0dNSKq2NfZMYI63JE3GKFJdcdITNJfFTsCY/jqXQV6nQZQYAv0x8bQpvcNa7tKuK5akZ22CvsLjZ
z+AYwVS1f80NiLpgPopVsi1X7zlg9eEfmVqLXjioGKHjXWolEJyLRdbhbo0bmY3NnxcBOy62Zo7k
qBqNwBs8hvJwEyUxODDGtFTnsX7nfLoVXmA6eh4SxOBF/SsWnVakgecgq5M/c3cflW9HxQZx30dP
OSI3ERhdo9zJCfLRzuTEq7xcFLvpJzq+I+GHO1GS3MdQ+yoKXeePD4pbEK8tpA2O1u5KMTSfNUtA
M1+rhAbXJsLm6MRbIC59xhNTCvtFGGRa26gEt+ABvJ4muWQLu3qRQGABptw2Zk9rimL/D6j16lAa
6II7r/RkCQXLIGrIWYthZo/FC+ZzQiSteimRVJBI9NyxHVsmHqAS+ucT46FHlcnV9eK8O7mHh1Lt
LUeDaykklwdYK3BdZ+UhbMQtHdtVGLDP87f0ypuRbf78yGJw/yQz62xLC42wit9Ldu57ejIH2Omt
A+wbwMz4rGj46xjYPYSu8hafhI2iinw8/O11SETOOVxpezZ4pCYyT4b4Sn19GIYQSBWO8AuwEber
zEhi6xIIlqskmWfcYnXCX3fRvQkDwhYOOIfCHN3EcsGl2s+ACAFHRClM5Efz+bLNAx9MY/erHOhf
3cdRiAO4ieo4pgiWuv/N7ISoZ1leUdlIJYyrZpb/oBxxeUMuxyOdB7OA0+szeeVdzCowTcRaPITG
NDpnRYoA4xLYQ7NCASNXoHeKcQSEBPRC591TeOm9FCTyB3z3gcWvxFX+li2U4pDyXQDgg5TTPNiw
QzSRvtu2e8tVV/4ejg1SX5c+nv2zg5M5Kj1ld55r5NGCeGUbn4zFLjzFN1cHbbg57y4CS6zVykQ6
2YtWLd8Knc/mPO4udkBSLuTBC+W1Eyv23PfZ9BXsYX2eIx3Td2w6u6pa3cGtdZa5hJuiECgl/PML
/3SgC9HX8ZtN2PcfPXyUW5MLc+e293U6X07ec2uT8J61TdHdZ2krL8r58gdO/5KklaZXzMtA28Qy
UFCVley5ZBV9/A1pZus4ByB6Mp8bO29LDWjmGqTXkFixtO5vzACpTmDWe3S+Jh1aHkiS119Wg6Wj
mKAFfPJy624iqAsBSWuBshxntfFJcYIcHqvC9hjdiddn/VORuAUDtrYhg0N8w/yorwu8ffSO4E85
N4CjkaqMgLG8/gLlAj83o54U+bQdKrCwwxzGftvXxbUCV6J1Tssfkq1mUqBkUc1uOvLK8yaqxTkA
xP8sq3PS706KYYiQG1ELIuh0cq3ZyOnmip7K6lh6HgbCRNg06xPxhqeZcwdHaw3DS5e+ftaWiNA3
vRbDVFdwXPAq7pOJ+Fs/9HuZ1X9DVIYGwmIzH0fU9PvVx63bZ0nXcPyIcN144tghpnz0yTM6yJJz
CYYYkbrZZwzeharoQyaXxwQ8IFP7NDHleKMQWQWciPGRnLykSSFjoysKP1mQv6cjc9hRVzbjEwM7
QXw9wio0xUAU9GYrzxOvGG59rXEp3hVZeSr++Zqsag9+r7p+Ls/NeeGvrQ+lWyoV/IqaApWVUp3a
jWKBxv/3mtQ9u1QGpj84v/xzIb0xFukdB+tJs5r+VzG9nlwd8YqXxFgy6haIdcoDyyOlKlWYtlMC
JJxPHLzTFt6vpNy4vWALfTNeS04IrQcwYsY5csEmhX/2aQ/hqpLz9ic7NanMz2atYoWqMuoWEYx5
1ZBMzNS9cdSh/AW/CsIuRiBLZ8AbJ1c/OOpFGw5GSSUjlA/MiNveK3HaCj+3O9lYLyAA8y8UXDEX
TLwzg3l9Vk1skCyBaFicF51xM83qUp9xeEG22Td306wf10r20tay8tCrz1b1Ie9VFITnEmK8hfj/
wG+hsj3VgX2d85Gj2Ffa2VCGem+cCpvu3XFx8h1MykbZQO/Pit2JPtiTR8ViA+4/goaGTGMGWayC
UQgZ9QMk1Y0HeqJmjIOXPr6Ry1kAl1FX5mkpjUSUFcMxAW/YT7ZfeBHZ0XZIAHvlx541vXFDXxCx
MEkaEQ4X6TFSnrA2eTxdmcnwe+XxKJllkR/K1Zu7d5xVZkYob+RBahoarTzWOwas5QJJHtmHhYHO
3WsYzS1OuLxTg2TzP/UccwY7FJ8MgmhN5dclTg30EyE5Bi4Mc1hgDmfg6P3/4O05MnK0uWiP54m7
1wQaExDMPcxaW1bv44H76DuhgwQREShBo1T5SW4YqQIVR4ErqPO3dkJtsv+p9uUE1QaySeezOok+
fG/W/hbWBZ7nzhphzH2/7byOmI9s/0ITBhSy8oRh92XTWsrWO6T4DmQ9jlNSm8WVBRlxKQvZ9TDl
bkxNooLywWmGP1VRrYPjYiJ9tTNVVbltqRmQ4nKcl/uAkm2Is/SFzvXXQw1qTIFuE9rJMZczFnpF
UxZ1fF75hHdf4XrvziAujuG/TyuJej4NN2SaHqOxrYOzQbuwsFY1lLzRonik8i4cQ3Gj+oDS3bIl
w+0HhB6tUGAMYhGpzVyg5HpPuXHMZSxitaqPWcWbB58a7QrxAR/HZO8xLtioFIb+9dmHmB7yH8w3
a+DDSGsiwv0PinErIxqWkKytG5SqRbERm0ttUJwwqf6lzHYhMQ0QG6jrqjZVAK/TqpbbxDwJ7+DW
SJVewbc6oWCzLkpPl7CNgmpsXD5NZ7034ijgRFMYD5lo6FufoxSerTvyTAw/m6BJuvTZv/xWB2WO
96mMUjm0PrTpfq3NaVNI8Q2rY5fzorENLr1JvZHvWag/QrDvch49IyS38k9So6lLjPEXooq4llTd
rXSrDn/IIXgOsLc176I649cJJSxIVzzH1GySm/TRvxo3hug8bd4HYIQhQeOaOs0VqvKLgl7bNCha
INMfVY8J0/6pbhiPvBXMHylhyy7V7VVo+ONebnrc5CAT3MG/1UaeuFSvQe6MwCw4N+3f+JnKVzIc
4x1JjLt1NV8VwnJh96agrDWWbwxHfSSSnhyhv2ERuAVAEsOJ8rcu1BEWTLNkcOcLcTwuzTevOev1
nzn8n7+hv+Rg4BEm0vkM6EdkwUZtkqct8XYW9KY33LaF9rghA1JDb1HAKobeoHj4eVjWQbv+3/CY
x02glC2U7cp2dcZJ1WSwGNwZAYkjrU0dLKC7VjmUmuO8bcEQXnAt+7FFMHMaRrvOJTg1T2gYcBGL
/oNBc7dk+TkzboqqBrRqPt9GzRiJexPKucilyJsg5P+eoTzhCrmL9WkCg/MekTea3B5oVxVpkrd2
Xv6m834DlCpdvenEHyOEuO/qBXDvlx5yNWg4AVDXeIw6fuc31UzDS0w9/0vQ4WXXMI39VUD5oiqT
A0EPbCypTzAPcbSF7ETYvVOFTwiiNOAITf8NaFRyf+SDq7cLlaGlMUU8V6Tv3eq7HhJXqb3N9pMp
tQREeH2cazsscZq9XAdcv3OW6Yqu3JfF/JrgWqD53cjIh06l+PQlTskZ8UPPI7FjqABXcGbdFlt1
GvRnaVw52GkF19GIMsG+3SIuuJePjrXGHhZYJAb8t8nplMFVrAXk7SRogC35M166x3ZFOSkXAD3W
cE8fbneNm0JC5ssdnvPTDwqFYrgavhzHDqUmTvjrcjJsa2qbvPotxojJIlIA8nF6cM89qJ+PVd4Z
8Td+fJlOPqe85r759hBlxU/inla2sbx2MtoQ/CHBHMDLoXci5+UgplbW2a9j7zdkAIDcNZ45Td/j
cIDIaYU8nzCAve/X6sd1MwJcKciTDzr1nu5M1EyUdK/bXSq0VTzLAcDRAsrtpGrk3S3SyWMA5Zft
yGRGsaj21y31uQHomXWygEPGjrOKL+RjCWF/V1E3ZcrnuRbSB8Afgr20DQpWHp8yZpgUP9wYPtIT
8J+hMV9eQ90laQu/nLSKive90ubK55k3YIbgPXN9cIJixjWR1N3lsLer5Jgv41/31UdFN5zTzQEB
yq4n1VSvH9JAb/rMQdKpZm8jYrWxy3+qOhc5zl+fYTziW9nP2V/a9m9dSwQP42IcGW3h8DWxRupN
dwqvQc1i6QFqnw3NPgCW4VABleeeMDIkJ3LPTL0Qs6IxHoE9Q8Iz7PKfjk1kC3+LyFOU/jb5d7zy
/oIosOKkAvJCGGGY2jAteUOoVvUw+H6l2j/BJne5sxmXiEZZlh2LOtaaQQh4VGJwK0MUhW7CXM8f
Y3qH7EeJESmWcCLKNhc/B6Fs6wl2I4KGdy5FuvHkcYhZPk5ywZEG1HRNdoRw33ulyJYnUeS49UTO
X2pNWJjc7ONgp7ByeadSSBZKLOmJuPrlayJXzY4Z5zblvdQ6Zy2AMupaJ3O0HePjQU9R6vxIi9ZZ
o/PvzWI8RyJT+fi+QWmSJojCD/zIxSoD2hMr1PYwAaprxglcQulE/2DPp4+pFBtvgFOlwS8cW/e5
xYB7ChXd/kCxB0CjIBlkkZO3FePFrtcO4UCF1f/672O5McsMNVe0HaWq91/4eUl8pa7uU8awOgeq
C4gMPM9BZ/TRbxytJxun9MaEheeDuS4wA7pGs9o3GorbvBISYAuGw5JlDrFB29joaGFmT91Anfiz
8RLk4oL3MMJZyBcTjS0ABenRH9ZNgGHYStUhq+MlI7EjMvSS/5bPZUMq2MXfcC+BsZJYIVx5IN7v
mdSTndbIjaKdEjd//oTnU9Ox+jBluD4HWxoMLDIWiieT4Te/r4Um7m2+dUzVbIvZTaHnaKYaVROI
myIn746PiWo0UIQe5qJT6/V/sVRLP0nlWOE7lxuMjf4K+Zw8hOOTjzkm+0beNNLLJ+jDr5E07992
kLVjxJZgGjPWD3Vi3sNvDAfehW728sj649mfYvxd/Bnh+vwFHPMaPFnibBpJhewmEmEJ8f98Mf4y
datHE3aPMHdh6oc8yTJqQym1/NRAznOZ8+E0UyAwLb1bNuzsq9fATin/0K0iWFUG6Zmwb9llabQV
2iJeE4Rjl7FBMWHZiWEIBG5jeGTozkEK2Y15RK7IfRjeQq4sXb2SZC/wO411uPYMAxlQcGRqMbWr
cK5alJHoZX+g4WghGItk0KrUeoumtM2i8qqSroXj+u/nxTCfzLYxmxZ/cjimY1GPoSPWHYh8EwMb
UegZCQTo3oa0XpabYPV2FHBm67QmTPNZIdJYOs/kT/1gF3uGso8lEwNIaQmMErd2AIIlK96uDcxX
gX1eLSOPDdCYayqTDiQQdVk5rFqw6EnkFk7u7po7l4IlaK4cA0CrioZ0bH8uwWxlHfTT6PybilrF
pRAsOTESH9b2wHFq55KPIgSYKIigVtN4aeMkYpBfzYhaTRfDGBqLRS6CC49GixysQxDdXJX70TGn
jJErmncqrFGcMW4/IW53gmCXAcsGqQLwT33UAzO3iA90ueGjZQJCZJ4IjsmKhQ/cgt1R6i7AqtXC
XBDvxbzNKe3T5kg0qPWPx8vlZfl+mad3wVaOsRKr6aV3p3y+2BYLfALBVg4heDsJvvY2TFdYEip4
cJs6iyB/RTdvmI0N126WKiOTsxo5MjcmGMIiF6z9efU/rbcJ8Os1YYU17i2F1scw095iTFP2ZYN2
WMVwRA/c5laLSJVbYd9JQUCQWfzshfKsP74cUxi6N/JuRROYaDsJrkwvqdwgP+UFoJ0kLckDbGBK
AeALRHHLF4OgP59TInQ3ZjMe+cyLialnZTJCg3SrcyP+lME0JxN2cNvha5+G7VwW9ei/7oR0H9kU
h0Kjq/RsWqXlDtwoViT11MKklGH4THPvObRU0aZbRXAYxbnsIZBq+i7ayPcARzkDOSXNGG4WhE9l
Birmm6M0ANfnQai/VO90HsDG7H/aBOtdoKCGytqJ5OQEK+OJ50e3Nrt5oVeEHWfGvfCNzbmwy5eq
wFzejcIemZRlY/SFeTOfhgjdRUOIcRNrNDT1E2Ql8OW0ebsGooRaYR/NEFhH3IuNortzsekRirZf
SrpglA83pkLCgNt8Em6qMZc/RDhGOvcXWsk1Jv2QbGmEuoCJKxGGOJcTgEKe8n80rIdYXyb9a3+g
chFGxfsAkL9Eb/2AN7VV7ebwmgudwe+jIexR1LLBaHb1L7kX1aliaXtgCdILpEubMchn7qu6g/bE
i7dQSgUEyrpmaBqDvmCgXYDVcwSeRHee5zsIH8C971WAXJBI/wy2bp9RoTd0Vu5SL5rYukmygweL
yNfYWeaE5x8pJQw+1IMFgZTG7Wn0XctIxCokBuP6Qo4lEongEAOTiRJSbGx2lUr+QRG9/6H9Hja/
OYsaI8+lj4viC4MJxHMS3I+Zu4o6DaPv0sNDsnTC9tR2YCTUceQLdtFwMoXewTA2PJ504/aPcuOx
VHKhGeaiv5hhTB4lmTp6WEoqGN48rpCM6UnprTL9DANXHYvaG5oE5mnS90KeVio7+aed+wo3FkPM
dDch+Z1WsbZ7k7csWitZd3NjMwuPw+RoAQT0VNfmY/tpY4xX25ifOSOuTtWkkY39/GiB3LExeWGg
6s4OjuPUAwSZiGgoJpUn45tKsccEP8UpH6dt0Qp2bIvOb4APVo5EqlvihaHJrcKSv6e8jQljCOQH
+gxyKqXMH08Yi5PDLE3ihLhD8ZHokDQr0qoCgH4Iggyi6nNqUvfPSyXxRJpRfs6qrl4vy7y0O/tr
OB97brZba8vS45/hNNI173qjHA+8rCBc8nGIYBm+2rgL6MaLzBmDnGrSjnxrYB8TuZbMUjSSt/Ci
cw0wobPu3ixqwaibtpeyxmy6cQ+X7ypASoJF7WHDP14mMrxnobqkIV6TaCjC8v8nDpVl6nZQHTG1
Wo03LpXkYHo9vWuRXBfO3Hu333SdHylX9ZmRuioDP6rqtYIEUMOKCR3MAh8LG3D3H5a/KZ+IRPHz
n6UPxYTXraqOjdX3fUoRUtpR8aQ7Qjuh3VV5NgapfCeQe3C7H9HqfUIr2+a4T7E/TGCMRUpYqsu0
aCESHT7YVo+xDFGBsFOQ5O1DI7Vpc9jxE2pKf/x8ZEvbBdZwjTk3Pc1VoOGL3oi5JdzhB21m1czR
sgF+OM6cJKY18Qd39smgrytAPe93wfhCrxBbui5wSP1Rh5+CGax8oVElzcjeGrs7K98sAtgePyp/
z6TA+N8BF4ZlQYEtjx97vWSEKWsbmNpbqtpBBh/LxyZMk8Qh0Zmr0hfad9/otpTlp9Q6O9qhPBuV
k5XEW0LAuMurQEaKGyOLWEXE1Cp5T076TaHEfJOf8A8lFzh381SHczD4ddlIyfd9Hpfecv/v8FPy
f3Xgfq/XTlDNnbfJ9QG2WsjKq5yQf6vPUrb5G+/am5t5NJNWJNv7g87ElzhuJ9lhNq3g6O4w1Jua
UbO6TGhEI/xOWHs0SWI47ovmcHyCtFd8hk59AuMV3EtRF5hBGTInK4vthVepuiDnIPwG5ZiexnNJ
Hgr7Csk0IYGT1DF9KfIQN3IJ3TOZrO7sa6yPXGLNgWqe8t0oMGSRU3Yb1i7nYIL2v1WbFxdle2wR
W6aWhkQJx8Q3quIDXPTZPTRWH6xJvECOyFAdug5c8x6pd6iX1ZWA+oO4pR2zfgC+hzcM16IPVgvq
d+23yz6eTJw3vQ04osY2/zZU/FmDUTMMEEBog1K6gjN7a3lK5eXEbZP5LLVVVKVhGD9XDog6Ry3u
V0FFbX31e+aq0pfp79LiFvHQd+zo3LXQtOAQOqbR5GQ43lQRAEkW+xsu9Vd1nPAAcnZNT14sOBjF
VyXAkDbjY6eUymgATV9BavYcCZm+nBxUut6ZKzwoKI09aLejkltXS+OclgMehh1wzz/DLp1jDHfu
KepI29tNgyo88mRacLao7k0n3GJe4okTSnT+Voc96fmi2/30cR3L6RwgbxYYW3cwqusdhqZp5+pW
bP/uR2yjJS7rgNHY/hmGhPrDyT6rGVj9f9x/AwM1n9uxOafDarTd/6cFPFpsTcm57XSSqgayT1+H
hJm8ET/LRvQI7+DERJvt4z4hscvXLRqGuqQ7BgX5WXmA/q7ai7a7mm2LK+hC2H0R0BmDnTEmkcXp
5EVjaff+1aV532t/ZRMqVAcRBPE4barJ2gGDJ66Go5OYIbCWumIg//TsTvrKCEUM5XkIF8goO1xj
hnmbYkdR00o5ic+OO8SGYbmwR95kJUv3vEacbgxGIX8tOyVUl/RFECYnb3I9PVGa5/POMJNcOrUk
mCONWIUQag5fmhErvb1DXzQJv/J7z2Pq4Hy3kaE77bX/Gpc1XXv1qKPrNseQcqTjPIaD2puzaiic
t5/+apM+A3gDCVyab9lBJW+xh2Yyczx/6mB1jgQg0QqLoZNd44F1MwgsqhAM1iMSYK1VEd7OhcKi
Y5f4NQoiBm/XDAA34ckzI3gCeYvUCBzjfDcl/TdbpaR6O0iO3MO/1DHeNVhcr0qWX9e3ufhCMpS1
fufS4/o9qD3K+0L1WzsLNWkyjqX3JFPCSN2KOhEHqHGvvheb9I/v/QfXHGbYMjYJW52TfpodZ19B
jpsFbU8MmHOGGysF8yFNrWhNgECx4KEuQbk7Oz5tv1yAQ43rz10hlRB/wNEoQJy/EKv4GAAk7VMq
OK6yyFXTM8TtgPJpOLW/2eAITSmCfhlHB5q8Uf+KRnOc+btI4wgLpEe+CODR3hQ58XsLg55XmwUx
lxjNaj5ozH1gZKCHhISRE7SqR5Fo5bpYBpjxD62ZDg2IpXviBgP4lhh0VBQc0HVOX/kblSL+mkWq
HKyRdUkIYBvot1RM96vyyEYZipktmRJHpKwuVcP1TQ2hUjDRUq97m60oug3I4thIsGfz1Yl+mze2
njIaIo837cJl7pOhmEwWvPUFA0vq27Z23G+ugLhG5s7R1J+CNPYHKGaI90bevE81Cf7kmOWPo5Ek
0q4mPbg2rzUeKkEt04v35D5rGonf8ssSCB4dqbA7VQUXniBKT1txsOVyMs/DTO80zojO51IxSNuG
tHWzKeQ3Qtod5WI1XhnYx7aAtREgAtNDbDEzK2EW3ul5yESwDGnMYLmRQhq4nv2D5bAjwPpJLOrm
iayyGAgjwXVz7rohR14ojvPIOuxyxPn2OqMWHoYiyuSn4QIMKl7gpJjnTqmczlsk1mVu1ljmXM3W
MDxsVuwAPdPzF0ogNPd4Uu5+OqekVaYKYLteU+PiwIzCWtdiiye+I4ECfd9qi26uRgvKpuW72GYm
3SjLiqzJaUxD+oPs54hpQ46tTeFUFkgehs0OvRUYp7BbwnjyW1qoaVCojc9Tam39n/WQ1xrIvmhz
IC50Cj1Mtr8buQBjonTK8GnaUfoDZgJtDMPJUOHE7qrm0Y7muUzUeEe1Rw28mhUDcp7RpNqAySD7
C6SbMDaowSP9VYrPlKkPscJCMjsdWYMjCxe1tg4a4ITRKDfac0mFLwX4G26ok1+IrfPrd6BXQhUf
iQerBUdubc0MrbYnCoW2MNS1tjo/r44svleUcNc739hSlCCmrO6vBo9eSwzKX/umb6AN/XYnVvWL
81ECESrEk3TYzvm8pfQVx+Fiks9w76tRIB3KoEZHakVE87FenSH5aJXMW+8cTSANXryGcp7qj7Sk
5Z+mcVknNPqahQK0tbTbImlrod53ezfeD2UoTn9bsDYN+0lp9Ns/0bkL3UV0exAeKAMT9uZevErV
1iGVOfmweq/gSGXRsLyJ7ZGDASQvAZEXE1AgsgVII+efasRThqEa9+6moMGVOVZTcXWc10jYhpb9
sXYJ/xCjt5725kKNw4zruSSc676p4fOSxo5R0FYN54O5hAsMmYjFPPZIriz4PNwqcSdZhFoeiGyg
gRZ5Ik/8bLqSfoarezBpxkpqQlMVH2wdPUEJD2jwzJs6ZT3bAg0dw93OwkeJlUaFbpMf3qDaUhEu
7P0NGDljd5oH8smufLRStBiYD4gHVFwA6FHhxlMSG33E7TJOKmO9glDzDaXIkNnzPWPhLGbrk8or
vOvL21fvmB4MmHLB2+baUf8oahUR1mAxhvVMnOK/TcMh7E9XLo21/LS7BuWnA2GjjD8bzQt6qCkE
u/UC9LIqoO+lt9wJomkmawNjLwDsnusrVyR7fMyPPEsUEBNGF4patUWotnzHCEguyVB3dEbduVTY
UBpgmCgTeBST9F3fzscXSosp7H7b1sflxg9wbuj5wlAy/Y3BDs3TAGNWEsWSZL7LEPkz9PnMIub5
A+bgRrzgVAEZ0f2bjUZ4ClPc/asAMEk+bHjdwMCLqytTmAYUhA+O3JijnaWZZaNteMYSPWX+7EMw
7nAiN+JwX0yGTManp5rAfeALVfrk0R8wAvXaSFtG8i1sYJPi0N6/b0UXfncC1sh046BqHhtdAQ18
eka6YCt3BRqu2R5myhlLbFb6+A+VnaE7ovAC7Znz8GMS7ZoflI/2TtDdEdQglpJBrbazNFtGk3A7
Dr0DGXj1QbB+YbUkpYicqZfmjGP9T+8GtMx3w2yyu0nXcnLWciar0dSiH6xiwPJ0Z2zEV05lxrLk
4z8jJRSAFLEJguh+LVK+xDR2zq/EM/jzWknxsI2diK3I2Yem0bxH3TYPqXT5ezAMw0SHtc6KaS3I
Gn7WThPpytp2Jfr+XI5dEbP928kyzD7X35y8YNk7E2gxq1hcH8NG1mKrSDRRue2haysdPmi/RfA9
q9yDOZLHrMwuKtPOqm+MOn+drc3yzfIPt6spuaBEUR1ZfvTMhWhYYlvPRR530Do2ZNRkOhMZtF/x
mp9Ody4vzmmR5z/1/0kH4wPUVoNbzeyPxFrb61xVAD/ELYLWg1U59eSzeMDMIQeOAutwNYopP878
Ym4JqpRiSs8T7Xj5n9tZ9JWOVQeHFLlb2LH7kS4zV47FJGKusu+BfgTogrNWzlODNVI9raiulcgM
J8m/AFpnIdgf4gRCIS+iSsEUEvEuYrtzg0QuiCwwkGV/62VUmfxVdLGp8yhQaTOKYZzgxoiY/8Ej
BhuOZntT5g10BXJGeM4oRDHReVlnbNX4rKlX/z87NoV/FpLeWgkeeXxt98uSG2JUt4d8ll2WWL0+
/mbnObZ16S2VY5od1P5KmmrZfsosza49nOvikAC/bghqsBWPJc7+b8u0DNbVdWpCNnN3wwb52Co6
tllOh9DL05xgx4KfcXh/QBj9vxJ81Ee6Y4smNibynvpQczhg1c/44dqHxDyL7oiw9hQDW2thmnlQ
1k0ikLuBQ1K2QC/XobnZf2eiahsVE75cfcQLyToXzp10SxflHGAEpe+Zpz/mM7+H+zMm6wqNQumw
ZoZWl0owC2PNjtI03K/jGxGfnG6B2q1DC2e97RJJ1mAUBbzAirQrNSjcDRkFr1MEQFQqZiidMGgI
nkBBiHTksR+SCJ8JuMwPDNron2qZzCh6Lr9AyC3+bzIVOMnY8g3/13VZnjdjEWR4It5p59dX/EB8
wg51Wk/x9jaCqQRh2Ia/PiCTQ2He77uxf5lGL/z9j0VZaTKGfPABuaSO9g9buPQ60wyoNJF3Ou3g
iWBUsbDJFkRxSh0gcWC5Tc1f8t6WsbncGju6i1YnLkF0Hhi8uOKvC74KvmEolGd72CzLiPPaX9+f
Z7Zgw/U9aeNvqh1UBXf7eJG0U+k2NP/5FllBrTs4EomHjigeL7WvbSbErBGkvaH3ZSvHQ0ABKCFx
yqUHcRBeJdoTlcfn7jLog2UTLUGsu6eK1uSPPv2ORt6ut2+kix3NepLM+4aqqVl5CLr+umpdjDzZ
QKxPh6LVBR/9rOnBRUTjrQvpnTHe1eY8SYCqFIOvCBrse9QB6oQ5EijwiI3L91dEMBG0begqa17t
ijHtLYBkm7BUCY3dbDDUI5ee1EyQtvuHUmEFEJoMPyKamd68oytDVAW9l8mYMBOUEhTFJ+hbF/g8
h7+zlvG552ts6MuObxkvxeDWplLzrgGkqWE49stg06kmutRJ7WSsCpGyPU3pVca0/WSALtoZU0o2
jT1jgx74ST5pKvZE9DBpTgrOVIVW8wDLjno8TxOwldyYQ1XEpACL6sDxiNmAVUiQVKlcevfew4B/
i3qTa370nDK/MYNcbnS0c4X7C8fwp0KV0hr54tXmLpTGB9cFAZbm8Q5W/kOvGT9y6cdV6KO1mqjG
R7yUP85yP51TYov5kx5JhILRiQObphatiwvw2FzlfMaTvgc9g1sS6DRd9SEUOjg1HIY5wKTCAcZN
ZHumo0yIrkRw7Vnn5lISwiAo19yAp8Il/43U6cs4Az+fPWHZ8KhSRenDti+kGG9LcT9uu66LhHht
sIpfkGrQraZJpubKG+WZHUFMW0GbeHKgBkDPl2jzeeHwdgXcb9D7yBeGkSeEqYthDuOIqPLO8Y5y
NAFszufud25PX3yvKLu++Hcce2t5+yceSBNJiKV6tjLbSGv+AhmS9USkHgpHTqdBbNyNeWJqQi8J
4ffOA6F8hnFIHGeBujIMYrv5s2i4CqiA53puhN5bcsYVCYQrgRqQlVW5+zidx7L+BJIgX3rZfEFk
qigkzPutg8WmhFL3IZcIIGITEn538qjqMxYDLXU5VZq6ZwLxUJURkB6keJWTIfGRtXTJ8y9f/Ymw
0ZTOqmho3eNSMXOTO9RtMuFUNKcFGtGmRKBh2GSGzWW2CL+1qy/YMGLKo5gT2W8d4TGtNOQkEaYI
midVDFLnCZjIYZZQY9da8+h5TD0A72XVvSyDwXAcYQKI+akAJ66rKps/LtHR/eMeqt3Bnp1Aov2u
gx2iHqmyuZ16CgWSkesG55Y9H2YWwmtBrUXntf6dYtU62MTZBMsw2LpJRGWIOoKgSpFzTSTqgVi/
uV6nbEuzSzj45iKLzAhhDW8Y/dLkVQ4Hd/+KezgUntcl4n4HjjlpClytumcjGjNFhzvIuOalCebW
2adp+oQPL9tu9J/u4Nh8JfFSFetUmnnNp2r6+G4RCPBCRpzBmgs/iPeruK0r6bXUD6UhaYxRIvX/
d2yMCsCinoukfqT7fNCaPegYcsDT2XK/iijOmkOeOR5iqQhV1tYemgsk8p175VKk+fuKP2t7Uwdm
SkBMWUzXJrY+/jLOS+VjeLpPX2wPn1H4g7LbJxqwsAyAen3yaXvzziGYiv+mjHTZokgaX0ZQGRoG
kaG9qr/a8am0vSUpa3KCtVLy50pYKBmE5llGO+mOw7P0MIsUMk3jR6/TXmHA2/4kh60OuzVPnaUE
8Wc87rA24pOoA9+YvlVNn/5So2klAeQr23fV4eSMDgnitoM2GBc6ZxHuWPRmCrVuE0B/2QSvBqD7
wv/8MC+JJ6Qu16MjmxztIShlY3Dg5q9E0dF6AXE/5Qrkoemx3X3nMZDCD6o6PV+mfYGqzsg4wIkZ
Ffse2hwBDwDmjrDSUUl3T133rRESKfu4hYWew0FXbnSy6OGJ28AM+uy8NxWvI975jEgQMoVmCX3Y
/x34FysIc0b0WglFMFNebCzx0T29MEE8q8uu38uAB9rGTCH9kqR8bv0n2Hk145Of00HmLdgA03Vu
0oRSGovJzPfQun5D/xq6mxjQu+FLk4ZhSpQTuOjXbLPV0/a8NqPeawwqME25tnG7kOXXygCwZkGp
2uJOSAoy80G5+W05WPqzQxLS7Hz7b/szclat1uJFxx4QjcnizMloKIwUuHjyg+tSlJP+2GDFycab
ipiJruEvR3H3mk0StBijeYX+EHISyL003BgJi7n0+IP32IIRb+9fbnDbE4WCI3lhPr7lpkECW039
NwQNjYbmPA9mJVADD/RAFWrYqIYEyz9Ld9eLRlonNDQVR0XYPujVSyiERk8+tTKOGcRbP/PJ4RO9
kn0pukg4UuybsD7zOLHAVj/xj2R4K8cozgSTPx/6kc+d0FRX9+XUkOgZkm5EdnjyB699EbMskrDk
DPIso9FeQ/BbjfSnQtJWuN1QKv2zO5gXavkhD6JcrdwZGEXkCpN5bRPXuG6lvL+369/riP7Jo8cZ
pfs+u8TkrMvR0U02zGz7zpPioAgBULy2r51oOoZqyZvS5kQCITRs8AOApkP5Q1mRVetJNbN1JedC
riXjE13LRt7mcsePVyVqa06tjlP6YFbOxvV3fCQlWS7CjTtoJWkLb6/kMOZ8Ed3kI7Tmcjr04Cs8
E3pw6Y/6lNF++n3N+7Qrdgzc79PO7k/tsGH85KoOQJbAtXEg05M+ygbkSW9ChQPtsgTrPmgwW8AM
g4HT4ky4LxEx7CIGwEuZYIPR038Y2VIVxfSoiyc0YHtzd4GJl8O3xVSeTFCymE+HhUVp5rDGUr/e
Tu/KdeTVUC1YaSv2hguCv6LgNzEyhqRn0OGGrhKCxdpTpcZLLZc6vV/wuGACuMseAy9V2fpOGDwk
5RAfvdCmK17VHh6goTcz0qL635LIYJ+VhhLGBAUHIZyrRV2oV8ViFg9KejbaMqMtLkRTkUgVemaR
uNayCXnIeRQYrnsQi3fvW2z6WqcaYBH32IPis9ErgqqIOyYDuyJyDK/MogVM2ZjeUGJwX3ysDimM
EPRPVASAs1TncJOfoqfoTAM5x0DUIUrTlGJPK4jcT06jjiMJXfwU8rrpQaU98O6ps1PLJE9g6SfB
OEJsrF9SybHTmFFMLUJrkChLp0JaMXArkku3MgsLhXCDENCtpk46eeaQ7hsVx/Gob2a6/0rGPZ+3
ueGtvxI+oETn3ZJUEQpcG3yeszdQRiYBfuxbQ5AkPXoKXsS0fKMBGD3ZVrsqH0y+bm1pK+9Xn8up
lmsFQrzvXOizP8y4AKKX1vrHMUsmzkkk/IrD9KNJBRpACiz7lCFIO0R+3YjFyS0C2axP/OzPvGot
5DX4UDtor61iDrM7N1v6UZ3FXhjnd1Rk1zK+jbdW320hc6BHxjRCbwObESfrSWi2zXCtD6RwZzWk
1UUH7thdGvumxt0dsNsmgdN3hS7LVBrZBt+6F6NcFcRXP4YWRGXrxht+ySfA3Mi69SIXVMBzWyjS
yvUb1UPfCssG0g3YXQ31sPn2aVUkVXUalhdHXu0S/fOunkkLF/9qX3xamxydwotGcxm1Zjzep6qy
FmEmJ6LQkbH/aBZEmZf5lDPbBMnPcOmq5i+43AUIPQifQyG7pE2FfsCZ5MrvaQZh4T+6sygjo0Z/
5jQuxzMQw2IHivFTVRXUPJ8QMWeBZu3CsMNF/gL0ehkDYjlXL3DpMUMgANggnVyyBtv4wAybjvA9
RedxxPYZAowNLzzb0klVXGG2usK8TLLU5Z3nPVPVzJ/lcBDbSvnHK+t1pNKaOujU93C9eo0j/klN
K5VEBrS5SK+DFOWxSxdsrvMC/IwpRLTf8dA7Hdgy6fTtrO9lX7CDwZ7PVTSJaI8u1F/eAZmzY6Oe
fgXDecvxudsYyJJbliGCyH4L8cfzzm0ECyebqKSyeHpU0RskiNcpjPL4TdHKtSzpg3AQyuFdH0Cg
KqmDF35CbkZW4oYEwc9pPStLja+bBJy5SQ9/kAuWP5+gBLC3Vqf0Dwkr0pm52ceR0avUozEKRr6/
nyh3SdoiQSgCiufYlk2GOGnWYmQn0E4vAbT71KD6d/i+uH7mHK6c5WbsZXLWMIJ0aiIcc+KjvAv0
yZtUQQvBPAG67wrP5YqXR1uPsRwPr7MQWl08UPrhLSPD7x7TxzsOaKyaLOsJbdaZ24haqWHctQp6
s1AcX3MQc/ZLdzRVkSN6MwZCwmldkcpOhwjx6Clm3hhgeENUANF1WjKGsEOgqhINZUYmGz2a2DsD
m80lxeTqDk7l6YhGh0tn5o6DP1NrPYcLU55q3vFcbeVvjEAp80bteLrYUGRp7/povEDqwGcS1//X
wn3Zi2N5AgQdexVcOAMZy1sxWkf2cy/wBV0llyvxRUKxOY5pQddlX+c3rhUb+j3CctwZaNvawcc0
YXVTbzLvxvYNFJgsipegutQsekEPp2wr9Z6NtOaML0qYc27cQ5JHo813x0U9/ipsGoaWXerzS7mD
83CkLFVwtKt4RN32Ag/7Q060TRIFVeeK0cPnY2YyYwqk7gSOzhytGndEsw7LSQaGVnD6knhnBn2u
kauibrKUC+vZFHqpk5Kl+0rfEGj98kZxYA2x1FQrd88vWP1cq+Qv1naFdIESc8Mf1qJydxmrLpop
5dm6DMCX8sKQ97vaHqv3eLqjV6sUo7aDpQMPwnfcfRmti4q9+UHt+6ArVeUkiFB9724Z8BJY846y
hqUiaiF/sec6ZsgStTJkfhPAfDS9mxTU3dXTh0zVrz3y5b+xN2LqZEwQd3eFNL7reiL2hjM8tcED
nDXRqeqkxK9KT8FK71fFTZEST4p8c/JikCCdiaMknNEsfOWlhHwNLNNiDFtrI+gofgv762UBOH2i
lgzDqlmJwCuOQMxswGCszaPuE2ArqSJCxGUDbUbuAscVk/fZOrCTFC4ViKWqNobl4S5jpN/2a38P
kaQBtaUMVqFZCtHuoMa4AZqTGWsm9vo1U8drGwpo8Xn7NLDyNkZP8cyBRbd5P/fNMSPCdTdKzRBJ
RoKEi0Npm3vUGOkyHIRgteVPP5uM/x0HlRvNXrqgcTgVtskkdQOKTYaDt6+Xq+H5Nf7sD8CIb5eJ
80FR3IzMCzQKuGAcjcP4MszZiEsp+/4AOcHQB3X5YoXGmYkgAQBT6ZO+ZIV8xKIVvtf/74UZmr6J
OTVvbf5OtzHjMWcFRH7q9Rp/MEjrS583RGkQ6eHdk9udf9D82PzzAMhoPhCcpMDPaqOoJZ3rld1q
ObO3ZPIRoQ5KoRc/d5F359SgonFmfLokwC8A8CekbwS6hwUhHxFTxLpFmUvS0xF2nYwMiXepMOoc
1WbjQRP8N+4cCrD8t3b9uMPotzeqpagM8OSTdszxq9A3EAsQLsycqg42OFYMMjKlzAHkhSmpEy/5
ka228JlG0f8l6/0ZkNLG9Q//ZeL0+aIMH0GRz31HkcJrjFNEVvyj09vtWg50rmeRzaBHDO5LXP8B
eE404Wgzkmq3+BzhRSqM6EmAydbvrNP2JoZtPtOXAOxAyg0E2TzzcsGlUdIMLA7n6v5ICzRjyDMQ
fiFhByH8RBeBfj5qzar5gg8/uxx/B9uhdxfiWjHHVK9ltqUU2jylLWi6CrtD6CNBF9HkkBGO0oBD
+v+4G9WDsDlgPFV6M6tC+CenJDqRrjYUUSVVTKqvr1MAA9Uias++I0LtB0u1IUYK87cQ0kO1RPYp
5kItb2NkmQlUm/YWGwbt69W4ozyIFgBxG37RfEr3Yc4AXg/YCtREvK6vPboIj0mRTB/VQSA5klWN
OeumVvd+MbxknT64kd/2d6rq5Ik+YErghMrU9K9prVh7AfVnDtKBxRMvbSE5bEbmVdNv5E9Ry8Mb
gf4jJhjqnaZd2IthSZRX6CVclNlcSWEFX6T0bh0+a+tw9bLssdPl0yTxH/OV7VDqSYG65B/5xuPh
YP6zT5wmEjePannlAWsV40GIsxCH+3wGt/2iOREmldoM3Ij8BPxP/+gjOVsAXS5XShjIng7GCvBc
5LrLkDwYvB7/kjaOMq4A/hv3vQIH5mjE6W6sNwI3VM4gwpW+kv7UJSI/AoeqKig+zT9xm0THAmdB
3l+0ef64TcZatkKCTh+usHDPlShtIcIiWKhQ/MZdyu2C1VbXFk2jdeyrXrquTFKdhkcF35ZG2U0c
vdvmrvn20jsgjDtKid0yzGUEe2UkY3H530Ql//z0lWOB+cHffKng4euMHZ9TxGf21Nlh7vSi612p
5s6yVM83CpYkhCquM/DOUUtTaxssGh+XyLO+gupWS//qSCbbSqUCAM8lX/hcUzmXkAQMxMiPqHOS
JHBz6vCJK9LNgtoYQ/cF4C7/kyeWH3O76TRQCI4Sjeqp4wGwWo2n9IvFEW/nPCP/CHuQcrxt4QoL
ZUpunXGPTbRxd7isaaHknSijYgbgqun87K23BcY+2ubfm6D6aOoHD/aww1ppvBnmkhf2hfA82nIs
5VdDARES0LWC2d5nHX9jS5f8lZl0sBxkAlTMlTLgv9DFhgDogDsRld291FzuAI3Z3uw7cYnJgJ8g
9ciL4HwcCtHIcIl4fZ5C6k/onQOZHmGRV5nbT68zPEGLZjA2QHHH60gsnEHXruwEPawlt5QcIDBR
tQnwZj4fj0WBpPdYCyjV80m9toIevpSPmwgX8K8/haY///KL9Ap8Dd/WSWzrHdrz3OF+L70ruX5a
NY9KnydGQnfts52M8S3XOFsq2fmWAN/ZGhIj6XM9/AhzJdGs+x3nlpntTlf2iQhWF9kZKortgImo
7zlS4PE6M/GIR1QVNhQ3qck0yL6OG4/0HyAuEKBZtaleUjPDMtvu9MqDRmUuppSnXVkYWy9bWXBy
C7JA/rA5GCVx2SuXAfblNRB+OH3sPvhOavei/Tpq+shrPFeG6cNK1fUZwPghbGJaX/ebg0Ve4DUG
FNlXqPI547r/6/WwtBCq2HBibKeOgRnZAhP25KfeAswL1P9m4TLnxqRPwuTdxsJz2Lu2yPjsBnCg
VoU1ja871h15foBWojF8CxOaffy6jTrzsQ8A1QvuIWBhoB9Ml8R9zhV75/ZZHOt0ZRAKTaTuC0gh
UtBYGXWgwNYqHB76lMaoH4lbeEfEMn/mhkElcV4WnlRrfcK8f+HgtWKbaMAp7xiN4h1HE5QkC6SX
4zINy7BK37gWuD1v8KyP9gthEaXDtO5jpsxWBZmvJJ0AE75BNpP6Z+ae2VOBEQy9DxaoCi54b7OF
hr0Za/hehSV+xQQVUMGKDkMgdd6sarOYAHLA7tkK6SYj0DZIe8pFif5drwonIhm8+t7qIYSKuZiZ
lIJ6972vTPqkjNJlwjUUJ3mS8BbV2bT0rs+ILr14o4dJFcBbBHvR7KOpbXLAoLF9rIRMTkB/qMfq
keixEf8zYpAUW6HH43zqY613YKUXMkrnXYHdrrQ0B+My4XCeSMqbwZRei1AWRkb3KyJi2Mdbmf4h
AupO+8Fbbk9wBkvQqbwKpxkPCU47noihtJTbHdgABqZ+XZ5Cs9fPliVlmnAF4F4w+4HwwtGfpviv
JEkmTNKxtdSDvadkH/iyadVGhbNHFoigy0POaX8v1G6ViefLhZ4KLY5L9ZN05Y3XHSrbrAV+pxk8
olPpCZKAudX2xT0VDhosk0f08SJlhHelyoyHFvD87sF2zsIcFas7NA6+SEtXU7DBZ0MkH3xeOvR1
4axzni9tI/9AobWgqdnalvuUIvE+rvcJR83TlaiB1+5fnIK/KkOViInwiGZx+jbHkC3g9gNgVKvn
cADKpO0HvIuRBVyzN9LLD2gFWyT40K9igG1cSdev9Go5uL9mzlICu1IjdgqGBVJBV2v7QGT3HIwW
gYyX6G8SXdQLOyvIxJN0Jp1pd628BpYsyi16Fr3CNxcSafpL3dqaUqLm9VGyfhWP3s7SdGb1xX7/
s92SQj6lM6wFcOKho7DWCbM1DwIrTAS6vPGbuPSfz+k5F9/q3dtHD9agtdd+PadbxvgFC6g7wmP6
TRmdDxRpa0B6FZ1fDiDov/eJEBgBidpalyVK6pTtPPboH5V2JuVD/w69SWa+815OYvt9YGV2Bb8C
xWFbnIc/DjAIVUJ7te57bUApO3BBAWn3+l/tiLDmJbTjMdgWsmeGUV4cNOcBp5DUqagdQZrpE3vc
kvTdfTQ4ieBBOK+RoWBfLtV6/bAN5YnVG6R3OFYhn20NgxXnZqgZZIC5Ic5OZlgSMgsvcT0/eN6X
y6gvEqKJCq2RHjN0QeK2cY9duBQ2sLIC/CnIIY3TVKjUQ3VDrW7H6zdl0/p+m60xj0X/CuRHff4d
Za0vUOiXKlvHXlvLdRHsu74jN78No5RiVvOtcj62Z8NF+A4qAhIfpn6RdLjxFEP6EvFcfcObSbGC
pfyI6aTXIYI7QKBYS7asMlE3IU0vQjWJ3abuAFVf/6elkfaELdzkUNpKt3ePGAee3ftcOSlDED6J
AtizcejORYWHYpy+u7ze/nCRJe+dXSinBmtBAfy4A7MsFbzFv5q1L42Go3gGWwqQSd76i5rJPqB7
dpdNxzY5/cTTGx3pfk+QY8q0LLC4lyQWMDfOf6WCc0ZiJkkMymn0RxDyQon//tGzWfNMyq6iRXcA
nkjqQoWbw3ODa/qID+g/HDjFIkVlg2wEXJ7zBJbx6PBUnaU1GmNHELJnPbWs0f9KA5Tzajpd7T+T
RdjbmOZ74hBtfY3C1LSQesDVBEAVrnY2SLmnib3pMUJfhgkALjaN5nmCtiZPebwwy56bbzvy++o5
ryfotsbkKoOt9i+h5pxyZ9bzdxGTn5siSDoRh18k7MSaIGzYPSC+pzBHTm2sociuO4k8gnV5WDla
6bUVfThmUGhZ+n0KdPN+Lcv6G0OReRn4u+oEYFbnsW4c0RZdvcqUooMPcNCoAbQJlBFck29yrhEl
wSSC3uAqHZVZeFDbdTrJ/onztX1ckWyQ5pUd3TaadD8xukOo7+f+0/3d1ORYmM55LUhCx9vZ/zd8
94XZ0NW4BKpOBY3AA2pq8lYj0lVmNE1bJoGkJxVBfKdVp93K3iq9HpDexm6ZYKSWh8VXgjCiWv4l
X2JLN92sB3aplGOGdATcpze7Q5EWEv8WkV9pvQXwjraGH06J0GM7783LymW5pVLN2qDAVxt6x112
fJuF1MvF7vDpT+Hvo9zlgpc9Zp3GKUsRnaLdmB3kRi+Plm5y+rpxalh95h2fKkrSBvBWhqooPqBb
q0EIiMS8241dzva8Jv2a+h6DJyBpB8SeGoTyWFvCWoLXblPC3ZD0ZXjQm2FwxEn2a8T7e5jWMG2G
jLGpDo40Ww9LHGJJSVcVzKdUrEYm9DR/Y9Yj2nJwwLxj2Dz3d6bhJ1Qmhy98YHJquZrITHwTU6aj
ah4ZBDwoXTSStnXWDW1S2IQ4nW3POHXtK2QjOKAY6b1YwFJ5fb1FrvRFw3Oia1cipocUi4Zrh2xj
j4uyoUNetA+A7ygO6lhkKaaVnvngKtx+B457ejIZxUm4aZ74uCjpucTtwRJvnNo2+7s3V6PQqzmP
FeGNrDSVBoGcW8xC9vKRDWDDLWRNNy/ynAikak/qxuvi7dXKwSaOllA+SmZgVfbUQot57EORCuNo
/p+ez2peNjzyw9oK3fR0Cx/CqE2Wyggu64/4D5IdN7OeWasINXboYV2I6TFVr3D5YzzdYwL+Rqeo
WRk7kEmZfWqmr7goks/ONtnKy34jAn6zU0+g4Up0+4Cb8vDPaDxF203HN05Cf64zG1IhNJu857cD
mpvBJqmfPoG9exdvDTPCTGWKYkT7E48UeHR2trX3GUhxQU7jUhBDzJKBTJ5lcGB3rvTLgRfTK/Mn
I5AhuwUwdil1PkqZiqUqtiXjNOulLlxUN0MgDDHqdr5A2rdsLfnkBwzuTUxwf5HemlNVucGsuFNW
Ur5sbUeyiXHyfGC69Xft4D7cvkf8nm3tqwtkHRnm938FxfPyGd68jBH47UF2m69Zg3ptMa50dImK
7L/6dFXlJf50n+c/oR7DKZEiMaS905qA4alUQdiRu3rGnFjdz3LeJZExjbPqhkJyj5E4WAqjn1vR
YJXFv1KVlv7yJOBFY2z5SFhmmrfPQrs6tbEkHVGYpv0Jl3C0MymQiEq+Bzx9A4gdCZx7kCaVF24Z
2qir0eeCLDQU7Z9lYjrKb6ZxGKRxiNAcHUae2sghPJdhbQizeDIUavnkxzjE3qikiUROc/unRoLm
gk1fjlYVYuqVxIg27MmNjGjbqegeyZlK/1J7ouBPpbAD5QLqGkkaOor+0SLrQD/hiTgpEIYqOYjy
nghCA15FqybIRredTFZnFIpCYhDj6czObC6AxlsxSi+2SD5Jj85PvDPSb22qXMfKHB2s3USmqzt3
eelLSzUyIdp8oCLGGHB0qDDiOL38OZOOBmYdv4/a5wutWDbQO1z2KaY2Hld+squ9eKQ+6f5Nlck/
i9Yh9icxSyPcod2OY6G99OfLNNSnZ2PtitScJnlxw6PMR8FIn6jLxPNyHn8XGmUEza/4wJzHAB7a
EXxWD60LMRf4MGEcQ8PVAGomk5goHp+xmkUJJH7qsCRyvcE+Iiq5c6hICQzADyIRxh/Swa6ja4Da
jrBRDpgQ+KXESlEaOwD2QpXD0i/uTQqHWWl4FlErCM95jR2n4TDdV1TNt98gK3DqMkbNbKEYnGJb
TaUzFq+hD6tXVGwHNnXK2IUA8fj7TKcppqjMkBoudpWi6YDSeT6kP0bBiGiuGXSwCdRUQey0uoNU
Q5LeUaiRc0VdXRmZ7pwnT+uMT7lZkEg0gLmlDu8TOwSPU2Zr3QIJothvA63ngMeicVnIhJ2VqS5z
gEHYroY29PltdzZ6T1AROsRk9mwiDjoyekgt7oLfT6XNMp8JK9/1R/uTMD7xe/Y9V0KvwSWpVwA1
843CwiMrXVcD2F3RDDSe+JXQVUvtWZq1N8DAII1NIE9FU9qGdCegVPLZNQze9BN/vpYWCVbg4xKu
PqR4kcf/0dmbl8oHJ7ffpiAaejaJSGWNBfnM42bPxaa0EB1wuSaQ+OvV66r/sYyTrnln4k02KJeu
MV2eGc0ttOlPqRnvnSMOF5STW+0PVpVxSkCfJFk5BVMiz4Hsbgjq4Ikc/bcVIuSzprVasOH8Hvbc
TXMDeobKvWSdVtNMAaLuoRrHxEEq+SmNLEw5VyXvEOq4CURZ8MwKpTFKWeTME2BS+HOtsa6ZDGUV
tMNr81Y4zVckw9LUoRNQSk700En/MXQCc7G9ifDst4StUNnDGKnOz6r/eTy+TjzwSevpog6tHNWF
VoyLTuRTCBgDayyiDDyZQCsbSU22bxrLjtrpEhv51WX8KnIPN15V9Z2eIGkdJv0o9tpdjxBT9j4M
sk4vrfgihPStP8/mDD9wDOZU3g8C7vfhd+QKoFdri43016BohhHfC6nj4hgzS/BjqNqXD/5tTHv6
nssMYYDrUOBxSn4hb+3Y/tFUcLzVNLes8VObUQj3yNFOWlCr5Qo7tvr22H+qKlA2KM8f/FXr0qKh
XeRs6RDn1KOIMwpAI2P7WgelfPapFpaZi18pb+TI25Bmd6vyoKdvNlnfBnfULPUY43+9XL0BYnLL
L9I6SsKsM7ItiX06CGdSEE8IACpp4wmM6nv+SKlcAY2kYjSS89+pmvinc83Tg0PqLqTscL9WrPKh
5jxod7cw+MK/ZySxtaAgh5UBjr0l0lzl3/uSgNF1Oxmcya8YFmy1abidt+AX05XO452qw9oa6Nf/
cpDmY36KTS3peXsMUko0oKFv4HhOcQdV+T3BZBFP9dJklEM04VSlJjw0ZKi0GJCHzDMn689dPE4c
9WKBEJB6thJRXBtl8HoNMdfajIy/y7hoVRXl9Iw3PfFlyJp7GsGXgMt4xuGvqBl0YQ+pehmAIRYr
xyqSp8Hk2v7katq7NMvxGXzSuiuMpyhnnJwpQVf1/sxpnvlxLUU+iyiqVKeEz3EhFJ8dgO/GXJlo
oLNJX++6P97QsiT78BZyt9uQr2X+OPfXLoGOZ9PPPypLS76DA0A/i3YsWkzxL44rtpotr76mpTxo
fy0jd6IuCWF+ZEJFBcugFDcY5tswAqUPD4/Z6z+c9ScVkeXyAK8FMyk8G2cocqT6VmDn7lDNoH4t
8cnlNU1XiIHSq/L/3T2Gs/PCxODnLVI/nMvXt4AID8YSjt24kUqEniLGKE1pG3PjUBkhxc97fVTB
pkR/3VKJ1s2bKMZ6z01zDvtEyplPfr1LjHvy1MMA269FVR44XkVxWmfEGoEqqQQphj5nk3h5589/
TrZjzTDtc7PQBLQHxWEuNOCWuIJLK1zgoMfaAxodZTZd/X30PJlpLWPLyzeArIqlwFI89MOCe3eD
hoqRfa1BYnM0FP2dajzhM+LVrp0RfBW2yR0CqbE/2wEPsxiRDhBJH7Zi8Qyqhkr91LunYF3ZunW0
krqgJNOZ/5Xvci3ELYYsXSQYKxThS0npFpCYdFTNdkeziMkw52scv/0LSmaaMGGZeHUSt++wOX1T
YyYEF/5KiIInX7Usi7pjXGbc1zj7imGfllRPEcEM25R//cxDaXylTQ/OUG91FsaET17+fvgpesdE
0JPg1wk4jOkEdJOXb5PLd0xBxtob5rl7gfNXY5iMfeJKpd62SW1Otgs/qXmUjzvESzf30WrOVc8f
YJV1uMLpyhRFN44I9FgUnhAyLTbC6jvDRVs+noQzm8lzkNM1ug1K70Kn5cIVg4fMFfchWwNQsTEh
VFI2lNWtX84Vhe1qD+AMkKkvELfbpuIa1sAdQ4OY06yup1HTN1XUU/hij/6LxGgvh228pcY2A1xX
rpkj9QcY4JM6qIBb++36ghlVh8efoA9IjVaszHq9TwW0Vvzi064YCdoMtWDGFbF850EUKayRb7iF
TEFoqZ3TUzh4/ylYXu2GTPuxl6NmDslcMJpIxgahLV5tmLW2nLur+oHKVQzlxI6EWaIowsXO5tLd
P9PZpBeaeFBF3IYc9tuz/Iw7tHt11S3lW6kz4NkXcDJaydAI8L2A3v5v6KWDsc1SGc2HVTjkLgpL
mruoziqbKiRdRmupesKX8O5xzismaU21P2bUYnl9qv6FvQUYzERm5KYkA9kb9UsqbeOfiEN7fFst
nUX3259lqxGOMFTjL6Pc8b1X/luEXPRCZx1Qzr+DkEfq38sADwtgUQxrVpA5MoTz8Iz+TGfUiKLt
9KeSJlKSHxHHETZRxqwoQiru2qEIUDc9b3Z5fiTIk/9xkAv08CfcjcoxtOQM+xXAMHIqiDMcseLN
3ZtW4YA7es+nN4ewBUPWwXJ2BQlgDg6fRbt6Ic5I6RuD9Cs0+fv2uCibJYH0GnqBg9LByMUilgYw
ms20hkUYKHQr1dPvDtd3rQH+OccMgEGQaPbgkvNjxtCXa2uQM9Y1bd8FqBHHoH4sDJWkghrjc+At
93CnFi/2A7K2KuzHS1cxpNIWfY4G1mbtIWPWGi4AVC/E3mif5NyZ7hsMvJqIni4ptY/bd67e4uTv
NpeqGAX5HYGoAqS/RGftMFy71dSpe2OOaVlM71PIlFrwU0kRBzReaRnFIfvNwSotKiyRC4DXrdxF
knzoVxr6hPt2z+dkXnRL0IqT3tFXgaVmgueV27okCnLLATLMgdwV826AAyj8bFYZZ8cJwm71dxga
jJhjuhBrRmnBMrCYh3lHrxzK8Vx02YEdLlzDgalYylpLbciFT4xS4fRt25CLzlF+GIhZyPkbeyRg
HN9lWracH2nokaO5rSQjBkMEuhAdmLnzmDyCCTfTFmM8e8+dxf36LteMZZAaxwEc1PakrmjqNTX+
7KMdqQ1/t86s/Kk0ZnFSPEcN/9PTOn8Y+Ldy47IBZ2zk5eYganwK2PmnbvXGUciEJatOxp9xrLO1
9G16K4oUYCfr1S/d96NKkQL1wxDQ7ft+3Hj5S7h2hxCrk7wlKtCUY7aYFt/83zuj3V8HjANH5+eB
Died1TY41NSKp6J7u3jAUt8JYC8Ud115VV77yKnDcVw6qVIxygNMbp9zAY02dO6W5/en29HmQ9Pk
GoYYJeUhqgOwGw9/L8YfGPlBsP/wsDr1xF5AegOLDQDwh+q62mMvVk4NsXN5zNfYNGs0B4XSw/Xx
bZat9eG9z4KmdCBSVF3TijfZJImlsg7Gy9vFiUuGXsiNYA253AnZjajH8inCvN35bMvBbLO1NbLj
hZW4UPDqSp2TTmQJhlZT2cDm8y9I1RV11dQ/o9vtxHTCvLzfwsEMJm2nol1/2wupIczkDi+npxA/
NOK8DzNHzBb6nOtoEKyZHdWPeRJrCyiWwZc6jzx3uGECCOeASvzLrXbgsQwuMci5EMoVYrCQ0K1n
CLRDj/FCoomyHUvvwbGfWfn10iOA6IQReTQE6HAnb6nPfVDFNWfYg6ooGjACEJo60mz21vSuHY0+
p+x6GUalWni8UQu5MG4+cciEWzp9Zk7r8mQOKbXeBbv23diKn9eOs7nUEnjKVsPPn8lo5fhU4Z83
GN9oLL3+pVxG/rKTJyKU1agq+ScZUtdQTqJsyJEIEsDhlY+cG44S5MKkcBFIifLpEQpOL1LDfRIS
fy8SRzv7W1JeSJMlgasTbZNYXarUSu/Xq+y35C2Wu8m8pnCODQCEr6jZ9kGqGmGpYQhCwsA8EpxK
my1UtjUj9SgKRsEctVWGXPGg4Zrmnoc0yVvoJSw8R9XQ928s5vOwYZDvJpv0rxyMTLfy+lbyV04L
Jz3aZ78f32S3Rt8A17QgrGKYDIXHK0Orr95m78XBAkqcGC/PxEfq117QInagjhR8EhaJer3g5z5j
Wpx9tV0EPr7qiAT/48+ATCp4HvK74jMUaWAGB6j35V7/giI2nKcDZpNfXrqH2ymgYKND0MGI040Y
uzjCkle9Ln3FFOJgJNjFWYYkdWP4VS14eA26tR2a6t7Y23U04ESRW5ZI89OLjo6N4UKrQK3Iodmt
Ix1o7HWhQy0Tn9k6/gSvXQ4d0ejzbLbXlPCTXhlG9nrIHoOoVpzm4ki6BeWEnndnGbpJdptfBek/
aov0X5Y3ZnZNgbbaOJho3yZvWiB7kBFJ3yGTZ9DHrJTpKuZ5KG3fX+8ntCNO+crl8W8YCdy+SYEX
uOlZUPLO5Xvf4tfR8nXK2gOQq2YEY8lp73xDTjtDqnFFbBiOOjetYwFPDNgDCGIHu4b/t8bXwFjP
xkTziDUZ+O60mKM/8/oy+KtkR5PhgfZAZ0YDf/N4SRMuM3NJ0hbiFyhe/6+O3gal7WcwIQW4NgcU
7gZtH9TTKwB171q/o6srpa0jvm4aBs6c5dH1dmCkLloN3AEKEVhHg61yPI++pB9HzLCKorZPnjXr
f9F1aWDQOAtdS5VhY2s9oZVMapBPq0kOlMJvwZ25ZTVhmjHlpOtzOirbTWUAR9VKNvfbjxMB3E1/
XGKO48Mt1xUMjDU4euhWjGyzb6HsyxEMLKJ6ssqf7GueEpXvmhlM+NUBfq8siegNYa9LYUm6y2rW
XcRrh8dPGoOdaB9b0KVZabsrbQIZdytzkd8UxH1KdLS5hkpyABwkfSiMyGPUWyNVNEd7rnS9py7q
/Om+BI50KRmgUGQijcZ+6YvVvhqcyOp8KPOg8DZby8l1El21G9V6MsO+hO/Cmer9MC90U9qAm+QX
ADs8PMnIONyQ4cT7sIe+RSCEhCHRxJGF3xO4401ZT32pj9ENfdUr2OLh723LQQPMpbVnkw11vTge
eQ8uR1Ruy1ViRNfgAEb3NvtrIp0oPxKMPF4tlkDvmPn23Rd/pjG3s0fDI9RkGPApjnRb5aqoKoVE
RY403dr2xoGCouTmqxKwY/Iiiexccxg2lqYG3Pv0A02PAzqj56xhhUzyLvgz2zItlCgUK5iCPxVn
LSWl5VOZO+CelaryXUPr3hlw0SAVATXYvE7rOHHFkFh1p/uaMB6R2/rB3NUpFS/75Ch8Y3YGEQZw
SvCtBF3xw2B6EmYY+NMJQknJ5aFfMnZogErpkGNQp+ZtqgblAsrb+AAdkjBXTgtxh400WZb9iCdk
Kfn0q06MBQ3KFcIl9KoNV5vfFwED0w57q+fk72KyfwYW8TTri+R2I0mXrv2maOePjFvLPQu0gl7O
RMi6SRyOmFqIMPmd8raq51Kb0c0g9ez5XxKGLaVEvHSp/JrIFDl2JBAjdfhJGYtb4OgV8iQhW/x5
rBOrLYMmORbMAhv9W/w1OzGwsPtpLIofbJMbHF4ImNE5xtShFiF3rebCOXq2cqz8VCnCCi/RRy4Y
c0Gp6JZllGvOJgSHQaXKWXr3btGs7+V0CTxw3SXVh0KUqVsM2BRIzYRLdI1UUvCqV8aOmQFrip+B
WByXX+sm99ctTXCh0url+RthEVo8vGcd75DSzcoGAsAR/j7kU5fT0QZ1DwOrc4wU5JsExYcC4g+1
8s526TUoHazFTv+MHC3/XEvF4GYU6Z0QBFerxkiSAmUid4+hv6EnuZ1L+N6Rv7o2PyBn1IMyW8hL
8PBMrOnPsK+NZlOr5XB1T7N8DyfLPN1WRCz3CYiJ+eyDSwvuzvGdAUKzOj3sqj7prZACb7voL8da
8TfhwokW9AELEsH8mL9OEKvkp7p9Z+vs85k6E7LNmB9r3KNKLZrIC5zGQISeVvfTc1+1wa6yYr7k
fRPN/EWbfHTVjlrq74VBQJm6evWN4GMGvnpd43e9SFgFf522opLH7YICkw9DHHZtYEP1s9yds/rv
yXfoXeE+iptqINSbh+4wIpQg1FQZHZ+7OinhnELtdAwemInLAZi0x3ONikjzNaS3mNOZf8kxSMWd
CP0fEsZskC6SdRoAiK3ZfmDQukWZ1K6Nfj3Z1JPtokorlrNx+Or3jVGOlBoj/g49KwAAnVz/06eo
uIZ3gKUj6tysgb2TxMitpQ5jW728TF9TxuR5HU/eLxxW7E+ZUR1N6b7jpm6X4HQrpvtpdNWa5jQN
ise2+N/q3tNlmyuC//GZoZ9DfalN8xHHP38tkk/lnynWi5AjDVgjXctS17E03Bh/zKhhlWV5m4TS
Q+DD+0cjvzlhAvwmzJrMydIl/lvMiuB/F+OfqqlnPGmSF+OAfssOEaTVm+u7ECziVRy9KEL8MFLl
NA+hR4U+6y1DkKzobk2SgwZIKAg+SMTbvel7nSvR1VklOZnGxD8bvjQd6dZ6TyHUTi/RHlzc6m0y
VjtAK9jlcCPjbwa6NBwZkL8TcNLc0nrDznG3Mj5JoeqqNC4kXqzVIYmlU1Lj8bBBwv1O42JgU074
x+W/Ac1caS8BWuh807jP7iayo36Z3rfBkY89cCnUy8WOuJvoQATLCdEUNoGMGKTAgXtLAWOv6cNE
w0hAF8+UFJq+jntnCfbH9cgWWUPwV+7Uz9oerh2Ent5VjidGeDXntkqmcCkJfvCdLeJ8vHMdICsH
DEIq9b6ddwFKq/eVk87+YGStNpyUzWwCGqrwGlUAwS1QW/q1GarjFmnsazeA8qoq5tm3muO3DvHo
EbpQL5OYDrDSUIuT4yP2RnkPiEZAA0kRM9iP0AazCADyumR2+J1sIcNeofKbU8AddlVcq9yh91vz
bJj5fdCIcZ9FhjRUyDuuQHFaWSk/lgIkpI+Sh05aqPVjN4Jrih/NRkhkZCGEkfEjG1RcH4XBTwbI
vzrgKjzFhKl9zWGDa/Lg2C1gHuaONusQphYcfIhuZhVXuJIr+A5cm90aNoV1ubviBP1GXQ8wpK5u
ZOwhZ3WcRhZFGlkV8CIz14TKF/2iDiFcUk4mtFXWwGl4pwPfB8MrELy3zN8ih8vkqFkfazJZiZpz
/5PcLP4bbMHtD3ffliyI2KRaT5xvShVyx71GCHNISWoCIWOofGM/wYBJUeplVevq76bqZMmGhSmc
bOiJp7N7YjSp5keDHZreLnluTbvcwhqi3zu8wyMy60D3hk83NvpoxhS2GExyaz9xKtjPHpqZBi7R
siQwTgJOn6n+pVFmZHoDuAVEuUveAigXmmUMMc/zVrjtbBzy4FCkQmagecZ8fMS5PGy10sBYLSst
YEeSRqmkELgOofM7g0jHxjiZioDtqp42aEJ1Q+olbSVbCjuGi/SnW3Pl/q/0fvwTrUjMisDwuUdI
j8/WnJExzPaBV65GE0Nd1WVV3DY6491/PsZ3CdiszAHMpdsZAfZWvHJ3WqE1Xk22dh+6vcraEbIh
9E4ANf38+YE4JkWfEFR9pi4DmejgrvUDUsjy4ryikELWuoiYz1uz+Ytr8c9BOQzkLqSVNuz8Srm0
ebjyTpU/b7DdTkqAjIHJkiaNYC3hUVOco80z2Ptydl4eBYHvUASRUCVc3lda7lAS8g1Wz965AHsT
uO339iYmPpT4vTFhUMUHyMC8/1BO1h1tJhWhv9vX3Lu6zculeebiCVMSmsRAZaf1/mPyvzd/32Gu
UUv1Na2QidQXgXxN7nIZ1usTlw4/gVxqFXn4laPY5+tjleisRRF1ElE0b+EUbtcXI/ZZ2KOzjNRx
Vodjrq8I4jcESb1dqUtyrYw15/Kcm3pA1CUhASkAl8v97/wxaLazxMIO6NQSUNTsaLjlb36K/hb+
a+A5Sw0ZxQwW7iWBOHlfQA+lZag245mYsOtcuxFB3NKO9qWtLQNsbh4Tfr5yIyjVziCqZ0Bly2o/
xn5PsgE9ktrrXtFLp97V+z01T1dIPDfL+P6F5PtsOlR8XuQmTUvvli7C25hVM24ao9na/8LTdCUk
sjOM2h1GxYNHEQfTyNMNjBX1ZnfQKq2r95ZonSgV0tNmNGMGRHo2qU/iQ5GkAXcDe3Ut05MG05nX
mCvnwvA9TdUu9kQtz+ukXgL/P+tDANmU43+6SbpsGiBZZhJ4pA8cwvpIsPqiD/welQbkDyKjoCfR
n0gvszMs9w8Hve3YhhE9cyS760Ewz0yKmNP6P8DEKYpgkN03QOG5v0dA0vigDEkOYnHIh1p+LGnK
RnA5WwiNKsVhvvk8pTznlGv9tdjP3CkJOHD0jjap0W7bBDc5h3pMGC/+4gBisaD0kBxLtGEHg7ZO
h+RcbK03AGLL/ajqaBOkOl4lhyXsRY62QrlW3DT5XV2YK+V1FKWiyaDM3vFdTmfljpc7rlIFPmi5
2NB7CpFwOKmhjUWt4S87tMdwOKODwr5Mop0PFbPcMzq2wk2MY1kVgbrII2EhIXYndNd3Ek9sefDl
C9QbSpKFt5EK2qJUOguCKN21jZz3hKJ8hGtr0EKxjUeYjDOpcsKFoycmHOhdWBE4pWkXK4HxdaR2
7nqA/rKiJ7qe5VvE1b1mJXDRETpPgWN+Px3f/4ILrQWidxwXqQHc3912IDR/ZtiPcbq4Zo4SAaYg
5XX4aGcF1kiE54HiB2XD3iCYG2FSegVWg6p635anyZepzRiIIFNY/qmkseK93lgwAfLT+VQX4uEQ
xFkW/QHsnybO3tkxY1knuO2szyN9/L00Mastp5N/YvJCIUDibuiAGkL5rQkZMONJRQtDxwFkE1Ta
VU8z+yT0Lw31iGpoQ7A0mpGtNR4B12vkedTXwGmXhh9p6S96pRs6cF7UXP/v1z6iFbeRMNjzbxvh
83FX/nDM9dvmHbVAlv1rX6xXM2tEY9gUCp5C8fMtx40i/F8SpFTGDa4OZLZh67b582N/Nw5qzW3v
HWC6g7DA33jvSggTL315mRfRn1YLMYQ8+0QfGCubzk3jlswYvQBbSU/37r2I/IIUOPuEIGejl7+p
rR2hyiUiVdJVjXsQnLtAJSJZk+JsDFTC3/6GU4JTJ/Iib6yTRliBN3Hy47/0LFk3gHXzXpJdILDc
DCATgOA5ALuBz5dtDGN4uHj0CHaorFk1BZ6D6svYt1Jntvsz3iD/L6jp95MnwIzwuVVNubRgrutk
y9tZOxGLzKrUsUhVG/fRAr64C2Zz0Bn4J5DRAvRAldIwK/a+Q0ZWnAFAxovY9qzpVbfQqUIk/28n
ShRVLOu3RTfHDdTjOgaBKdmZ292ST5dctp0lRps41nVIwN4lkt11UjnooCvRQfHEN3GYCC4utie6
/xjyOzr4+JMKBpMgQkj+QIK97mZ+gELYVWYc9sXU8PhBMsZebl1eohxPLjUH1jUNeuJ5otXn/UUE
I22Kz5UwecxOuICbi4+cWNQoacv05+GIGRtZkVSMCEanZKnxdXP8iB416kU8wqvaNAHdDC1UtCqk
FHH4O2e12lewirBNVE+6NfWBoRD7/Jinq7S0kIbtEUZV2yY4PY57HaSnnOvA4TcJtgXKzncAttcy
eUIX/ZtSabI+mgJ945so7InvMxfKFu+OuA82pmbUPIAEPmQvLzAt7FfZvtt5G4WM+3+rHUxTJ3Kc
l7S9y+vQ4/eYwWxXQ5SehlQpvq+SIhWKtvcF+s1EU80AfkCbThfJdtWs9vsRKcsaQIqqR03Abr1/
LEi31w2DE/08tU5GyY7YrXx59sFkMhhAVuHjHLEryTPoKjYXh9ikCpwHmkU+GE3BqeMVlxzfJ5uy
j6mUmM+puNN0R9BAiYOl3ixTaES+LzTZiQs3DDFItm0/bYWFQwUEHylf0RKCcQZ92FkiauK6ocxa
rkHw2qbdvauRCd1hJ8VAFcnlUq0UKZ8vYkd7zfETCQUZ0+5p26i4KazUh8fNQ23vphy8u2oJuZJv
5h4HTxzyKGOT9F5TffzlAGEc5vKlLB/bAH/Yrb1XPvA5fwFOkVJ28b6j19TIeMTZGba3oS0vVxl2
TEJbHVXae1zCGot77uJLqyNRhfFqeSP1ToTFxulAbNSH+ONM6ntGWYVKHrXHGSiDSSd/QK53Dp63
j+/oxytDCYtqz5m7zKLTLQk44kGFlXqC8Oqehmzi+/ZWWMVRlUqloeUzBhmpvbMPQRjcGUu8f/FF
yaGgQjG07uUBNkD2ZqzMcwiGqoFSNpwgpzmBddhsHKzf+LzHVwpr9Ar+M6qJevj+gC56c2FhsUS5
KiKFtdcII0nfRx4jZ/wCOoCatpymXN1KvdzVb/nj13cip/htoQbwQUr8wv3FeW5Bdihe1C+2+Ncb
/pE4fA7OBo/ogLmgD1oLcuP4eIxuaNj7rqRf85cJO2GXsGRxWqIjAVxuK9BgQLYR5cSfXsc1D/lR
Bk5UTrTy8uMW1ibNcT/UHIjAADUMLJhzU8UnKPDQDvJokNpyKJCoeFOeLuEejMQEfH/OAaduGy+W
5Mn8TuhiVq4YR1NznYwv3lW6672yCPLlWTkYzWWjxvGlnv0tWr3eyP4ETpIlRavGsJNEsQXZFg8u
CSw1U6BbSFbkuyrmO7LJECwOPbVlyGfsafz4hgS9W722TV0aUltTGE52+cGzDfy5Ocd+yCkrLsYT
E+D3vJb0nQWEs+7K8nqISjYbvQzqbwYmD9GQ1Qiwr71s1/gGuQ7nsSafIBEe38rD5aj2S596WMZe
RdLjvAf37ID/vIytFKzUd4zB5QPws06c6CQxI0PMY700DKr8tnCz2yfTQb9b52Qx98Z+vgAET0tG
XSiFwocwcv1trLNmbfG/GpRwXlwu8fnq7LO8QRyITxxnai0dFjhW+VCzJUxRSpWVYXawvzCcLSAM
Cj58NvLlQ/jDXvsHqgNTKvT3TPlhDLFlKkR1m/tWeLOBClIj2B3TuC1UeIKIbotPHvjYLEi/U/3J
xjcmj9Ke2g452CyGqIv6ffyoR2iFroH0c/YFq4bVpu6n78Usvd5WnuYUInCcmYeZyn1QnVc/Gt4y
YNo+yvHxAzuYTWH6mE3wZaB/uenKeItvbSkjaXBSs3uzDFex0AKMwSI78uIvqHBulpfG4bM3si1H
4XBd3iDvm+oY5eRQqXd3PUn5AbgaXAN1mNet8P3OR/zO8zkRBpXOudTP1x1uZNF1Koa6xtmWtmUx
XyagBlxvdZ9bhIC5i1oGjB2hPVLyMEalS9sitqLQvE5Mhdi17wiuwKjpzIoqn5iH5QNHXzuSA20Z
eE2INCUjGr4FQc5WbUgPd66+DkFS7f2tlVNqNTPzKk0MPcnjWl9DyjZFMNScDZdmuI7JwvnFvb8y
Wz95F0780rxEt216b3pOqbfU+lD/nb4qEtEQd45e24s+GKB6UZMUXAj6JXyyeKpyaIgpUuhBEy9R
JBipTW74iFHUYO/1IFq3caVzOBGG8NDVDQaUTwHHBgDyiPa64u7iyo+CJkz0YK2eyIz6hcraPm/k
eeLiToQo6Uc4Gg0kzEF1h6Um6J/4U+MWL4nADeIJVWddf0ErqTzGt5A53Llxx9iB3BJeC0ci2ukL
nxnOVL04t3b8l3iGzqVAgv4CUzeE/c9bt6jiriRYDd58nquY5U+0W3QujoC6YCYlnw7vjwwvr2Ci
Cue587ai2cvcPkcwYcIkJwgshSHFoG2KxWxzTcissjnG8GJO2G2UJScjBD2hBNZDuTjQbD6hBKt6
fENmAKLzzprNK0X19bW/XSlI1LFPgfJhDr5/9olibdei9/jNHUL5/lGl9YYGDXw98oVU2e5HAaA2
izMkn5RlTRPRu0v/8x8p7a4XYBcLd78v6t+GK776ZHJMKJvs4CRAEkl9oArcfGd71MPKJqZRLRRB
CnNCqZPuS7+K6/oDvUzcOGqfMavqdRwAsOskfUbOxOPwa9w2xRHX8ru7cNo3ARa4ePHiBt2qYrov
l1m/loBSu+OOQlAg4qJpu+0bRDFiyERzbLI2k18jPHOhOXggFblOjFz6GvSR/0Km1gZCTUwiGed3
CjunTsbyC2vMmoz6x8BLu76MqUyxDz3WPCMWT0td62sDIbl6LQQ0pOYbRPBE4jaf3TuTnrx3ycqC
ILATc3oHqG8IkfxZ484hHVqy92uWgO9u6oUihjjoICh+K/Vuvwxdgu+xTQBjXeBp/RRP1/Mq7pBg
BZsTA0JAdNTtUNfcbH3zKRLNFSet2LPKzWnfHP5feWp+SwTNlxjDOwVOGMQh1v8p9gvIsCc6sPWl
+XnAPrq8M6Rp/Sm28aqGT6SXbxXSnTLHZv3wP9AciQbz/zHV6CSiRlMwOeEoCKygFNAIX8xwB0h5
GIB5xnmNS7iOGa96lgaLjJkTzzmoV383g/YqzcaWB1tWCSQ6rzYpIs+kX4h9RE7kn+iE/GQOGe2g
lrpH/8WhuZoMHZM6hw+DLWpKW25LuXKm70fm0RHx0W+Y77gF1l2BSxPD2NzspqfIYcZS8T2wf7Il
gr+mfHaKozCZNgQ1GI6Qy2MYZbwdHd/4G4Hu2Y4Cv5OD9VxNv/FYFu6N72GuB7iiJpS24LXGIgrI
qYN4QtyrvPBlBdE7Vm/fVVC5WgYfqsAypdw+DMAhL6LipSQzPWxI8MUEw2w/WMFOpMWSFCiuoU/E
DA8k9lk5QPq5IEKSzURtKdZddIdSweB2B8AtZ98h3D49sD6Vc2yP20H8cjCLSjG93NC9x/UzkXYn
yAmS+lrirgM4xjUCusL7Y/yZ7kHA8GcgWXk2UbokobDFYcVe5Vpta19Caabq03ok29xLUZx90bm8
aX7Yr2HLq1oTuB0O+EFNL8iM5ePQHO9MpGEn1GXaqTYwS/mrGk2DFqT+loJangRhM1BWpS1QFUhg
XrX2xzZO8IckBoe5n2iRftcLsm0EP3D/g5oBJ9y4yBKJmTuoOA7ogvDHUxPQ7RhmaCD5NZFowZLd
rjFRN7RC+XtAyBPSCrzlvjQMnzc6tXgfU8me48rWziYdxaEYh7DYvq5ETQctI+QGvqlziqzLmBSF
VVy0CL6/Bxz3Rz79ICQA0XhBY8MgcRIcCtUUAc1CAJ5RTrXmlIF6xmT3D6I4Zc7bfgD/nHSwKTI2
9spkfr9yhF0Y1qFgduqIlFP9GSLvgtKeC54a42FWTcZLx3eWvcmkMBFMhkDycp/Omjv1amLlFy+1
/tjAEDqtiXbZcnXgcC8k7g+hb3fq3AcrILdnO3UJPolUjJbATc9/Q9ylh31kWHnwNb8C+VBeV114
+9EwM/K0W43Eis6/316n0jQGohZVTO/O1FEPb+vSLVsrTs+3pnBct01YllCu6oP3QE8bFEf6gld/
U4R7/I0yCmXhVfr3kcR2LMImyohxqJx+qo4kSPIn25wvIq4zN/NK1X8/p/8TU90cVHn2NnyALPbc
nNvdhiUJ7KX3hlZnD9mHQvAGtF1hDp341mGpupX7T4y2tn30z6WFBPddqNZgNCPnSMgMjy563cLM
W+G7s2Q08PUs2XtzBq9poXJ2uctxm69leQqZsqu6vT05bzal4z+fSD/IcI3vnJGuB/rT5zg5Aeyu
znJ1qdhrTXaDt9YXqG8s9XC2CiG0PZ1vr7sr8iPFTy1kyQ9XKfJg8IQU8RTz7pGiAG5TmEehHuMQ
VRjz/S4+fZ1CR2yP+L5lnR61QrPWCHQz7E4qR6ceJP34xQg8X96tmvvfeklv9S/YbXHbz9vk6R3k
iAxLwdp1KGFr/gdwkPgFXZZZkZBQz1o5j6JfpdaSOWa3DmG5CwT0mZcl/O97BkxpGpe8nDnDOZ2n
OX2pqN9AXDqnm3gPRxFvUFtPPwAkzmIJyRcuxy66aC4dto/3PEaF4VvqL+se4N9zKTlqOlUU/Nhs
QG2YZAvoFgbznV7YLKWtaC33cGcg+FJdojr2ZkpJVVU/hP4heutz93UP935NYXvxcOBdU1vDiXN0
wdNi6m+oCWJxYCfmAB0FyMOQWL+Oe+3fMZ+uPf09pDY0/x4W/YM6wI5TUdFcR+6zQ8qnZBkH83Xp
kHCOH0NtRwEecJ+kFcCJdX0dE47b8TPgOLw1QlmjJhGgfdiHwmjt8DlW1AhTFd6leFWja0TSKcRQ
5Xwr2TmP57OmSjxPaoMX0oJhRGCXFvRmQwnmECF/Qe+ayz517WYUqPm5WhqiUFEM8iO7VsDI1cb/
0fTPFvKd6XQxKog8scDHy9uQx60kLWhWxDfy6eSEvszwLSm4PNSpzwZo57sQu+JTytksSmvK4p/X
8/Y5Es4blnMlKJ2S5Cjry8ZyEDezyw4PacbSiixg273lHg66rSE92vOI/lDiya2CW6eLJU9ZKbgf
tSDIBnxsWhe6KyDiAIMoA6abJiGq8YuTexJxVjR+eDSlM6ND19WlzYwjnroOfghzFLo8cNMBB/75
YX2XbD4H5uSGX4W4wDGWFelpSkYJm6F7oTQvSu+slrqmoKSjvXJgDT+7OzNc+XU/0w+lGrZ1RsK+
Zj+jCiJoD+SvpPfQboPON+t4oJezHdwxl8POAF11qAyDmFMOD98bB16Vp1mQM4pSVYEbVC7wZiqu
n8EJf39SZgMXrI8p/LXxfKlGru9QpyrR9WvBNlj20RRogKRbzjDo4pnmsN8TFXtwxOiWx6trxIj7
QQuXKEFU3uSPGKKZh4fTjtSjxTxpVX9JRLBENTYOVSvfzbo3OGMg4qeVQuXQ9MO9yc3JRKORA+m4
+BAia0l75vJ3iDoHvKYvz/xrs9JElD1V7sZ37NESEYaQEcG8xZSN/zHNi1u32gJemlsq9niFH7iN
umde2Dx+vht/wIoc93xsmv4KS9XZu6vwSbciqBAzQ9dL3H+K/J4ksxvARZa1t3djfvrklnMPONaN
pLQUwWqiAc3O2HL3qLIW1FC9qlRj5EKEksc8aMMdNp47LPc496a3Dsm8VRsZ4USSCDcME7Oxvthi
P+mY2TFZgpulWQekbDpFrn0oqraF5oUCHFWiEAWQgvKMwCfVjXRqbM31nq4sPWeZ/H+8GohwLHix
rZ+6JBzOmKNd1YZMHdSEDx3ezbXylOKpqikbQJjeQnTJ+X5zyPu4i+5bf3ZrjOnnTDEDklDCOcW5
B/P5rS70/Nbb52HkQVbKzVdhyHI3BezLE9inlku2rYJt1wcT/eKEmEwbtd33NRCy5pxFJpYNdAWG
9J8zSQgofxyoktockHsMwB+swrvfE24aqoAtB4Zxx+68qL7Avy3qnbjj1pBxtzKFySm9UdayX9BX
/14gzjoXHbaNs7lAiSY6qTmWf7sSdJ0W09fZgpE8VGi7NH2WkR9V2weSBVZl+HVB85OgoNOC5YrK
O9dodnmW1BbM4DPOLIzi8s2Tjcgl8B5zXDmxIGGiX5ke2CcsjY0ZJTGBXjbqrAgEHe8bDDhOo7dk
qQGWDk19NFZ5ovpiUk2be0KAs/NE2Yn5ghwrmbSCTvu8hVAYx8swuX6ydIodidpoW9nVKqSxdiXq
lDF6i7/85RsSxenAxCD3A8hnwKyfWXocsVgOICM2bXGRY0IyvdvUrrgXE7JMwEPqxwcqTXoMbeUu
A9FiXXWPDDi1jLElSBcgNy84BVhgdgkvrxXGqG37eyoXMKeLeDbrQV5BjgLcBDqJw1ct0owuy6mr
FXz6frlU8hI8buIaD6DSWtO2948i6AAChdgCLtSARZ8fdFjBFlAx3AMqq0gwnOe5Q+0iNuqKsw3v
DBiqJ3C/bWcD8OjQUB7DqNLFk103kI+KRyqnwltkvbE34nDDxcDl7Akl5chXHIdRB/jC7Ue1DF/d
6ov9CT+REZ9H0/Vn2eymNbwG5Q1BYtjtbsAthTUOhtEm9vrzxMr02LcUXINZLz67h+AzD+lIqTpV
l04pmqnZQyXa6ovn1yDinwaeBJGpMcBFn2Co/LfF3BgeEzQUf9SV+mkvRWo4nKlF7deNI1foq1q2
YKVHyi3ck6mDBqtaI1jg5rjkIcxHlYwCessV5qONcDtImdgxA8LP5D/kNe78O6gLV7gUXC3ibIGH
DOv9lnRWbrRRa6X9HTOC3LRQwww/KF9bWj3MrevMxWyLeRzVe4PLr08sXK4h0XXIc4l0qR3DilCl
M31hZQw4si6FlK7tg08oPnLlIsHLe+prRr7mAyJvHFTwBWAKFGwt2VCxwWVEY1aMpISa2jT8lAxd
avtkJg2sDl4vwk1bE4so9QYAYmfXkHQbMr82DPLCGo+77roWSOiGtLKRgSzdjVKwnLeOkK7yjdhQ
1o3TCANlXYZJO8/8BKA6+O/dNUHRlod7Xn0E+CUP6pX9ptkSEo266htLoAnH760AvNooRwXra9M9
cmBg1fI/5vJYFlD+kC9UaZb7Glgfi/V4pvpTUswpfF+A5s6naZNpozv61Hl96d+ONH1DaNGo/ZNB
7qRTzg4H00iac+ZbqcJVpepDp8oqzhfDLfu86uiFkKl539Ul39r+2UAl7PkSV3Oe9u3brZNT8J8j
j54V/HlMWlYbxrvLXF3FtB/S+xe/dzzLvI/Tj9B28e1o6MWbaoYi/MdPpYGd6WSknIpZcH+TABZs
aU6rij38m1iu6xmOLZ+CRCKpT/ugevc731G1AYlvqeHhaV0ZydGdnlYC1cmW2IF7sRscTdrj9WpE
LTICtKWcjLgjLzx6d1Sce2nKdLgIbDJCYhAzxPACgXHDtQ1hSNfr2r0GxRKwJi/ZFi6RqFcnVWtf
gjH6tRIwM7gU6YT6I7zIwZxUQD/Q8rYOuY7WWZRZy0Ekn8zZ8vSQipfxcGEGAJLeAyJrjzK8J5OX
vEArAAHngcBUSEIAvK2G/CUrr1vzDEonMArIKf41B3/z52wrzX5m6ScBWcC4rVBsoaKOs1pTVBQZ
s9EZm7+xD+0MJ2Z5KIZpvCv5FJ8iYltSuE3hFmmV3t0VUZfKCzcFAuTxkI6tIqPHI3zPwn349TZb
Kpi0nB82QJzlc2mdFO/V+oIJV3Y5ohPuOc9eq0qRV2JxUMLQocGiIkEQ3kb61ZxvPtPeeIaK8Zbd
zzrO4eVXri04WOMn+281M4Xlj+18W3PVJ0W3ux6rA1rpneinPAZTptc0iYyTfk2Bd5V7eMRXrksR
djEx7eKZc2Xtd7Gr/GeIcI0MPWS/ZnQtcAX0kIyMfebMiuC2YbZBHJoab2C8NlITsppWeIrqaISA
mEv1KDF5XN7JVVPKiXzLX9h7R36WdqE2VXnt0f4oxZIczkN35Fbe33fDVRChUl++p0VncMb10RN1
p0CBYvuIuPxn01NLIG2INUg+zUDZsd4RUgsg60hw097xqJ/6ioAGs0m43fs1oBa/JF0ttuz222H0
0CNs9kPEPWYQRQcAwLjFo3N6SmZtkrQsyW//1pS7lKyzHhCm6yjMitjV4vPMmhEoDX3OsjUbrOv2
MUvDDM2Zoo5aozZknNH2XCQRHmbCa5xbrcaJgdJpUy1YgudHIwQzhFuqYRsmEtbOwoEYAhkC7xIJ
HRFYGTKOVyevYZUEKGis0wr1IVgJymvwFwrKpbbhkzo9qQuSAq04ToeXvwTirMXPAw+92QvE8102
tdlF1aXBuD9qqy+JqKi2Iuurs/fSW8yXs/m0uYdT5m2qlxXZCx5aann7fEUOvd6ui3F8jhnppdhK
CMN7xxCcT1irilOnkf8cTB5rgvL+utYkPOvYvRc851ByvK/XLAWJfb1f3miXrVZW+9uta39+8v5r
5+nUo20Uz2kWfx3qXCTkaMcqvxHKh3XxOCkLqHtgPd2nhGqVnZFIswj4qRnb4Udb0A9ekrK1ad5w
xj0ra1JbBTgYhmGYwy2SIRd19scKW24xHD8zDuqJIR5UVRDiPInINdM2/SMyGrANEI7ECmx4OAGT
80rriESZGJMkgzeNl1/KuwnwsKUl4bf4QZI9YVhf4+Si54SUm4k4cWPRMDvNxTdnMXfQ8lDO80V+
y6+he6r9FE7zehuVxx+581kmRMa77kDlFO9DCw+0yaDueq5Y601S7MoaIw4WKh4GxrxNUUfGyW8J
HUlm/KANXWncFPz6fNgUrIIM0EeLrsiM5vZeGF9IcK+xbkTK+JYNc6vMrlQ7qwnb1YR5cMDIOG0A
KX0Tnplkig72boagTya2IirZ2guJpsa/qeoQmseUna1no68S35px5fUfViUxIQIImfRo6UPsWJXH
Gvru6zO5p7diM0WYXhH03MJpQkXjRLdu5Lw11rL+GK9iOZlbNTfSQ2fpIc/njoDyBcstR84X4Sno
VN4AMk7KTQiK9liUOnudU2wQ3jOGK+B3iohxhAl+mwIad3nNnsHAoM8ZuMp7j9kLmuAc9zEViqDY
n+q5ARpttJvvQBQ+pAIlZf8pTEsdGDqkny37/j+8mToGfu9HsbL6clLMN7DRPaEGMNIzM6dZtB5g
r9zURFHb6TsavKcqLmOAGyf5Q5zu2qlzGz0KnsVQ4Ox+Qr1wIKaX0e6rPfcyjDyYqlJbtgD2mg6t
R24bs1p50WE7jLaceZ7U9RVLK9bwBi4x5tkqNRms/tLBnbmgose7fGm4qinZMQQYtWn2vbVl18fu
FVs34x9HV46/M8BFZe1hJC1Axeha4PHvaQR+y5LL5LgCSbN08bSSJLRxI8JPPl7L4JAxGEYD0jK8
cPdd13eMc6PNinoFSq1R143pFqjkV0PHYPW0qOY8EXS0a0e0epJXh40H05xo0gNYJW4ZvnMkzNpN
nLC99EBCQNIjH3Uc/9OyIn89S5iQs4qpa9CuOxYkwRsWeeBCPyDcZJ9LVHdOGgRjfPZXs45qN6V5
SJ3poKoFPXYcR1kjvQnoebUTskJnmctqndnkWw01s5f+SWfR9pAZsTKlE6X3+oPjSXks6PUlTZpY
B6T2FSMsLzhu5ETNaO8vW4C1QemP7Ov8f72DO5BDCzGPA0RdsKSD87fGqDlavLZqx4eaw3aUoE9U
Cxn+46trkeMStRVa3gw+9a7CzXglUAle3XJYUXntNasQQtXIj9qKcg1yZt1FiCdy9x826tPNJZpI
r1732W1fWcKsexCfJVu0jaltMPmMu8/rTjkw+eXU0mAK3qdcaCA+tztHfyn3F7bsaSZeSdvd0G9u
hWvjXZrBBNLy7qFOb19OLiHXxSIx0NllX4/QNqeZmetG7DkeUXdqK3TeOsyVpf4Sb/CKIMVUwMjz
t/u2O/ul/XllSREUM/ByCzHwFeyBJClyuNi0sFIosIKsz+gwZjwNUyc3i/AQ8TcN580+TPCXeWL0
Xa9DlROQ+5iiGmWTlTx6qrO3s0IFV9gzqwKNW6mdFAgSGIlLD8JQg0EHmHa6lbDrsReoVqa3QpyH
oAwGlDNKCTce2cpGb1G0A7y/EroDShn7bAmg4kHyExdEX0iVD/XTfXiFvtiCde47kb3Gjz5TCyqC
HlFKh6R8zfI0ERDP4WriVpNHLJm+cXAC/fuBOlX9nnFrfGhva7iBcV79v3bvz/QgD44IPdp8EjYi
qgqRodaV0bVTKgfcf8io0WI4JIvFdGNeE9bh8UQhb0lCos/5j+47XjGpdHIbiKdBBoHHyGyuL3nd
APnAz640DmmVW9wOqF+1TlsEoRijADTVMzVeHyyB5ETZgNSZik2tEetc9LkBoTdC6Cm9w4yPMyZ2
8meBRT6RwTaEv7vXMZF7iIrNOKG5batnqjUk99VnhVxdlSEbAwa4JCxxkHO0WsEtP8X+mmNTMRgI
PtPsI9J4Cdn3n/Lr68o0APgQ5aPYq9XTVX0Rc3K8sRyaEZHwxs4Aqv04EVxdPhMiY5si9MKfvdSA
LavIBdWGpCGnCIU3rq+DX3ss+cSyL+1OPOzvpyzCEXUSCko3gpl1vPyv6dbu7ymqSPPMg8FGkgSp
4l8elUwLnyrXbO8eb0qCdcrjG/RQxKFktBl6XhEsqwGYVL5qu7d4mQY8oaGmWKWhKE3TWxJnvWSf
r0VX//l1f0urqe/u78OTJjD8XeQZcXjGwY/sAwjHBUiZVd0oIXyx4sX6oJKuLozk7d6Oj5VhJzMB
6NqcKOaCGKa+2WIATgQEM55xHKp96F76k1s4I4uV27Ai5oTrVlAZ2dYe6XLpbNQIvmvCisEMSASm
COs3YejPf/B6+H7mFariLuJcJrhHQPvVp/xDFyLuSeAuDEhxr+8vwHTP6dFy6OuWxka9V87ponJf
r8LfZhwZzbws2rOIoE92++hkBvwU/A6+PVLzDExuaipGc5xU7TH5O4q+k7F8i76bG3u+P94vJwN7
d3dRTIBEiKm1cF1KVbcobzsoKa6gXFSxSUp763ThBlYc+1Pl7L8pRxBhqJs3/cUuScBFTWLeSbOc
cZFf8fmdj0HoGT4pgU+w9NlODJnkUcEdJ+4g9F4MM3USLO7B5OqTW+qnYyr+Q4pGa9rUfgCw9mls
x4ZQOaUtt/HIvJt6b/hhfKiYXEyboQ13MnNLisTM4Lln7x7fe1/NtHrsGiW7KiQdLal+g1Y6lk0n
lAvFht9rRdW13IL+tlV2hqL9JayZAajxSVVxoRpUw1V8ZNB/Bzu0N9DU83qlFYEHGz9CHWGyNdG4
iUUkT9op/cZ2zqesfo5VDEtrGAReE/dthE3nBBOcAkp1BUcKfrRuz+CicJUlkeL4BmBqFL7bRhxZ
CD1Wa/MN5ro1sDpXy7IIhens33D69GjjJzNa5c3uxTcQXXsKnSk+Du0xs2jNbKG6Qww3sOxFqQnW
hMLY+EJwQA/178qQttkcAm1g26Bu4HvBEwGpIAa5Cl2H7x0AqnsKhuh0M9KGAc0J5/dvqVKcO5AG
DAiVh1EKMRzP4+SY6wlZ2qbAV5Nb1wTUKW0jIBNjl2jwRUb5JT2tc4lVwuoFHWDPezd0o0v6wUpy
qSkhaPJpPKq8xBswhZPtlA1DdN8VeP0ddGWeFEEWP56hTaxLHF5zZ/PasW9tz/5JSYYRzrjD/Qxu
0zmygK9mQi4oymnmDynr3rM4IGNkGl6GXsJUErJqBJ39I7V/blO/POrK0qDm3gQ0rbDQ2GrYeKJG
pZwnYMKwxGsIk+un4FekHXNEtRndWMAenQgh0eleSQXtM9uQ/PDIQNjcRdoqYlOtWFRvhgYPOKru
Rn0pXm3qLvzI8HhkC3Q+EjFmQo1GdnJC+zKDhfX6hc8D5Ez3B3aFyBFN/B0PnpV0b90Gtslox+90
r9BDDryh1y68VTWFkfhcEG+yiyYLPDykZXNwC8OU54SNSJd8nfuma/4F3TXPu+l8biWI8ZYM/ese
6oHpQNUekfoTeWQJ0MSiEM9vBcLFwm2BZH7QIbVxWkUMKcrM/CIk1vRbdnie1/SJtOIcVsjlytiI
eZu8ZxRcHurAJdYIE7typNigNgQZKgdekF0Pc9ARAc8C3J+xzGsc50bco89XMVy2rwa3JgwmR9LF
a5B0oR44XYMvYgQ8LY3Bmv0poTEoLqj7ZrD/Q7vjXc5gtiNQERXTrmRjx5hlyGyrU2eFeaxlARJh
iha4yEdCzPUTJAAm5OKFFb9DzrqcQlU6Pclw35AssX3Q3oOiozPLA8MaKcRibUnub8GV2uCjHp2z
QD6iG5fnnIc5l42xnXJznUKzTTvq9GTOOZ9Gzg3MXC8ChL2Npx8LoB0FolQ+1xR5LLVHv1wdM3hv
YBBHA2xIZI3LWIvx50YBbQdvFnYKC5qRkvNzol4WWvunlwOSBsRocJf9Kz1OvykZ+6QN6fNpATHO
3+LNQIXgYn4KrmxakQL5w8RHXU2yaz3DnpaK1flC/DyRFfw+NJ0XIvV08MGMZsOrrum9IlvGdwG6
Wyuul0z7kS44H3aDmi2YtRG2y/95iaVM0oJ8wKqZISXyc3Y+6G9vYyeNylvAxzYAvq6a9mMc6PC9
BQspo56QvmtRlT991UG8IDQ1b6BuCAyTg0ib9MDjUqxHnSquXfm6Loluf8CY4OaYTGhidVO7caO3
kHN+stXKDaa0YLSGUsE16mT7btqDtPk3AaA+v98iF46iJvXZf2OplsM2Asne/i08/RfjhdLPQpDg
WlTo7rDFWxFUl3VQ/rCeynkYpv8NSDS7vFJu3jXdue3XG/wbSwZCobOE9irht2czZPPCSMjqcgn5
8mZqJu9siA4vw7i5qqgnaXkvf6GovMoYN5RwknJG7p2CiLffEcxBqGl373TcwyfmkbUXKCLGepnr
yDZvwIibjSRvoo1Gww2pb0blQCToO5s3yFOYoD5uf0c7Rcn6GWkH290qZ7OLfZBB96dSIVqm31Mz
NUVU2J+PJlFyeHS39p4OwMHjvw4WpV2W2VZn6EHYi/U3nGh7sSbChibFMjE/7aK8+VIjVto5ifQx
USePfxnZzY4IZ0HRNQMDYaCNCPyqO1WFn4otCBxPdOPRMLOc88kN+q1r1jjCKPPWpsYLk+dOH/Ry
Brz/UnUDaAIt1CVI9E6WzDe1ChlTerHlwzCzJFQ2l/chSqNoD+xOmvDG1Y2v1o+6U3N5dvgS52GV
9u/tcodMNm3RAJxBFvdOlCi7i/lKhC2prGfm1IsyhkCy/QmzccymFDYi59+qk02OBcevUF8sYn0U
V2Ry8LxphzGn6oYaBETB7HX9TrTjA2uzaHNhW7/gblCQSQiKSDoKT24n4en9Fbn1HTGEPLmIlEoG
9+NgogATM8duGqVOCFlDqIVX5ryp7HgxRhO46bKT4ntibdXDqxvbpYiOkeTovahRBEA1jf2ENz0Q
d0L1nuVAidFjsuyBMhQ7Su/Z25gvysbHodGR1IOrqz1ujhE4M4RJ5esoERKTNMqREY6XW3KYL/ZS
0XPeid9Ep8GWUDmqhp7wSi8i4gfwEvlS/tmzchbqOUw7r5XBrimJIEy7m4snwoHSc2ViUNGdwtGD
Z3biE26V8BgINyx6eV0nVRyfQENltcZYWhF5rzzNIoyP1h0il170Xg5RPFGxfGDGsVB+U1nM0mSA
QjhCnf7/8ZhFMX7xcORpgCMAcr95OwxAwLgm1q9WS5w1LUbD8c/KFZXF3bpb65Ry2cqjtbe6DAp6
pHn9dyGrMJ3sBApFZg2H5cuX48vC5FK/1YsmSmsO2SX9LPmkylVKvWFgrm1ZsBLqtVkGgeReKspk
g/Bi2qb0g7IqoJQo8n95zz+j/lQuy13PJtYOiqPX83KsH0PJhW+QVIFdu6Vo8+oZLizM8uEgAGrK
PM+t6RV3tfl1SvUC/939OzXVPgII7NHXtXKd/Xu7xIydWphiv4T7eZCMHdGVKVn/X+1tasikqNl/
KzPBmnLnekkEvu+PnVP7JqTUEEOxfi0+RhEs4JclnNmt5LQ3b3wrMtkEW4v1Kft+9doSzSACB3A8
D02qkqJR2+9LVGn2NC+lPbANhTDP+aHBhMUkGvgAXvS94wMYXqME1hHfRd1N796qMjvKL1RaRxo0
e7nRVJdnM7hX1jXtnvoXrnXGBv7poEY1exneYvfJHpqifG0SWYzlKIepnaKEatQXQUvxdnwp0KUf
ympAFnr/1VuwQI74z71l+TwtqXcWRM6QuE5RSJcPayqEWKzcTofxz7odwdRr2VTJAyYxDkB3ii0R
EY3MleZgGlMkoOKFaEwwHh0yLLUG/lzXHg6FJl9mxycuP2hvDzNxVv2vw56Hcge5+JSSCoYRxcVh
3kFouDnP+JruLPbMrFE/HbBSmtNOvdu74H4YbJL2ZyDySnA5ARIm2miPIxU+aGZWLxazsEBrvk7q
myjvrzszHnecSUhXIYDan3axaMT+61NzaYgjjMafGR8O/2EVAjE35KJqirBaMwpO+R8cEWJq58lV
StyiZiUKPFtpRAEwBBVx7temahJfv6Djc2BuuPfHI2gEO1mzrCTbNBoNo1pO4Qjt5N7jKjyj3SbB
b8336DBqTDKpcNUloj50xFnAZHJwmFVTGuKjwdG2UbmVR6B9xJ/Vm/mHA1A0wbzMA0hO4B6EpQae
+aL4tExsR+m1uN5wXHtp5AToB7Xh+MuYXN8+teezHrEjYZU7f0KUm0tBUIY13TOCqQQgMd64H3/I
WK5rS5mpWRhQYckMfdHpuwZiSsmG5A9TNYBfoHqPJ58VL2hAm4UW8tFxg2WyroGMoTLXfQn5rwZk
hKrtv8uPKoRSlSDBid6zrb7qx91kJ/576dN2Zf0w92gB8V8jH/j2rmLTyHMHK8BuGv5p7Rib3dHG
GMjjfhdDdoueVUhoDgHufQPiGq8YVlsBAL80UM4oUl5zdjJlmYSt378BMdQdKU3X/9M4XAbT3Fbu
NLOgB9wWf1RuLliSeNZsE6HRjwUq44yPV0R/lGep7ASEInK42ZQNj8aDFExQhGhoMRUqhUf1M60e
XPsJX4X47QBO5G5HWd7HNuNKQ4+ORt/PeDo9C0j/IOIuLCCKoKSvYQdMf3pB1N+Tivw+FsGU85bV
23yCig02WTgo7BFkQpM42lwwTwqaq1x+SOCkiO6DqU0X9z8VvLF5uj/M9oLklrQkky9O8Arh1iXW
7U8srk4xm2PMVdQF7SKdYFfe1ws2WhqnSEUD2BSskPUxoxTSEoEv8ZyHX+jOny7dbf0LuIwufFgM
fDXh9eZPLp0jRf8uvMOYy5Q6Xtq797kT0UfBb41kmRsQvEfJ2JgI5iRI/IiP+o2A5b4DUgL+Ubxi
ckcbRAABctjw7Ny9BOQi3Be1Y46fadKeVKj1oXQfdJLdbvEfoWEpfzeRwv/0TFNum5KF4ziFQbjb
bw6UwNT/wRM0vuI6lcmGLu3/EEz3m4gOF4NAd4nzr+ba7GOgqGgARFAPFNTQp5ZT6tDfI7eeSMqD
bA4kqNqz6nY7Vn9AapjBjkzas3AYWT6Y/WmOLLUiQoAhk97AW4vSxb6ri2G+EqrNcGlz7iP7aVmg
kPlUKgThgizscDTLPQVyhjaSC701W7zqBBKPAgqDlelORaYkjw5BYO5D7GoebFgc2Bz3L2sIvSRd
vSSwvsvevuO+p6oCjalWd0FaPVnMiKOw/rtuLcwl5IybSLMaveKrSe2CnfLoUNpXp9zqMUKDCOmp
JmxujvjVZPfDbpUE2k/L2AXkN22R0OwHD2vwYonAvJDQXKI6f1TClCEaVh30ZAyG9lTVLV/1rXaG
dw2SFf0Cv/rwIVHL02CYRnXrs9IUFe4KohzNcmr3ISkdHY0JheWiTFkJgsmTeZ/9JjNMXb4+7A8l
wqwDMefSCyXe8648vvDnsaNAMeSzBwqIxpDwDI3SghH2yGAHuxOHeg3PFXIx4sFVG1uYRYO4HtEV
wpn8um4KfjH4HQmyd48ybQrS1AzahVOSNzud75wRf4xrzUvWTgPPL27h8rwckIiO9OX2MjURRnkJ
rNU58xbjzjZBEoBnRe5uDsFAhpwnA4TvceeOkd6W6vHE7sr872RZ8aupLcT2syszKTnK7fJJAhed
C1z8Fql6VOFV1CDS3zVZpGxZb08SHJqRU64NJbKLUV6RwQDhcFurdkj9SnPqKI4DRU2NFIu/LEdH
SvZtVYGYsc8JN7ZOzzC5DBvyq7ukzzNYGexDOZB9oJypCaW/XGyrhODr+Bep1ov9Ig/Kb1U3Sv14
DP8rZmsd0pAzYjxMzGriZqD3RCYNsAIPWw3WboF6/3Sk+hMGBqAbiIltOv0qZE6FCyQ1o8wHa0g8
9ODbGZNOsxAI6y191LMyBuKly/az51RK6yykLSIOnDX13iYvE5US7HaLvbC1iLUb64zvfP5bh6tL
DaUcJNrIUi42oVbJe/MVeguTXakQp8/Dw3Aq3f7Z/t5D/0XAqcuMRPEKEcVapKC164WptdecJJ1z
8Y63fcLK85f29fl9qmr02Qne6Ku9hLzeN2YVJJzYtQQlbADD5RsIeTDjL6M0FQctZcDGIj5+XBmX
0O+PlbayI4V83HZlNhfUi0bDtFthoadndTDxhzvCEPA8U6t3SV+LxL3ZsCGorW2T92swZHIavtUB
vwEXIomzv27OSnasHrpnr++aWwJOnk7SSUtndeoAtDenkLUdWT0/3n4RpJFaQ8uq+4KFELlZGlA8
QtlY0JZY0E1AeOJyNOjqCPdMU4NE9qMmqMcb3B54je2zD84wWny+aHA1/oCA9P6GYnh72rEPWkKI
AGbJmuIRQbV+IFNEaVvL0vDVTFyLnLbtiASj5JYaJUU9sikarBZ5dGvecdJoTg0SZl6F93aMiICC
wyCTb3K5kNRiahRsrWrnluwYiietPZmivEZchAbmJqrURc0dc0m4Zh/A1ko8mrXRngG1VibcUxoT
FmPi3uqslUaqX+i0WXZDBq/P9gfZKlhAZe5HFSIuCiAqZTwKxTmxZ89J0wNWOlzZDQbs6uL95c9Z
oALXdvswQ2BFF3mZPidfD983GGx9wW7cvGxuE7y766uGmP5Z95vRe3xGSmv6IpBAJIVWAdUiotDQ
WR5GjS3Mp1e4mvs49Piln3ZqQlZa9T0xH3GwSywIJyDFmDz6bhKCBAFPtwJkx9jBMj6jVBV75Luo
8P/+Ty2xEtpbI9naOHR2fPrJ+RL/BgXLAzzRsZwFYQUNXEhFgizD/jDp6TEzsGWW9rvgPoAkWPBS
PkJEU3bjTMqSs4nRxrij+OQOPm+e4jUqBrrg6z1GApZOxsZj2wKsB+cQntgRZ392Gy7VLccp+1zQ
Jzgn5ZSX7Yc6VEHXt7aaqwynoqGv4W5iJ0EYmbMAtlRmWhoGPO6iNzXWRj8xm/zcSAgkJkMCiS0l
br9O+usuowf40f3G1HxLVCeICqT4ParXldmNtuAqkpG8O9IePzXLAl9pauas3cJ+wbP0ja/wGlji
2r6XhL83+AuTOAa5GciIB60zhCOQL/839mOY7dBSOUDor71xEjWDM/G91btGxdll3f49a1jHP9uR
jmWY9DKUoAQiPfTPDxR+AsvB6Fu2za1HArfYVQKJbereidae3r3fb8om2BuyrK8ohrKcs6iPMKed
BJ8bNww+QWNWQGSSdszWDxOTK5W5nPQagLwEJr1UzzpSfHZOAvkBZS19TCjdwcZ/LKFLbYch1XzQ
2DgWLrEybPpkxRDzgG7TekCMSUv5vmIhwyKG1C6aRJgniJC1UR9CU7NvKELSjNwu+EbDWFg3irR/
ElB4uVKIqrxjyym+X/aYNCnyK0TCXbLLJU8GJdNKhLF2lOM9Uh5p+IoIU7P9hWWwJEHoucJ5IBh2
hmjIsgxpGcCAT++IBHGft52adypp76USN+f6LMU2gqBt4ewGESTQ8cueq0eZCkUAu/As5oufo146
aSPleKiORsmUWkhKt/DiaIHgr9SiJfGSwyONQEJQMqkjMfEgGi/9O1d8HltMtMV41rmg11iaCSwn
EkENkayLmcfFL5Pg51Uodh6N6Ro3B/8mrBGm/dAr8G3RghG2MonLo2bsQQuVKdTivhbJkcX6FfUl
5L0Y6Qmtshi1UyzILG9RlS9qnw7z2JNeVJ2oYo+111LLMRVGjEioBONKZw65MPimXX4pU11FN7oH
4AODAVlz3a8idPjUCltQJ+PK7VSIbxYusd7Zddhr9hJ1dugbK0U2k+E9Qh9Z8G6fth2INAqalc2H
jAFS8j6qk7L3Is8FQs0f1cVkxSryhu97gdWU1eMI63lxwE5UK2mzQMz4G5tOSSsAFoywgxn9J4+E
0PDl6evFoDTqvSlXAP3yO3XWoEON8zfsKLzay36Ym+fgnw52I7U0jF7RTR7+5vyJeS7SG2HnjOIJ
ic7go59fxj9pTEW5tE76ZKYJqjGz/sNZkjAJhNttVIYwZ+Bd2ZkDkn2DjJ15MyCdhf79/vspNuGH
iN12P8Taa57eQ+5olEGu+jLy/srOQ1xjPSjidGiLb5fvD278PvcGDVWvSxXtq1RmQYHhXhtsELny
AtYimBLV7fLUVPuIeMjIsy9E2sZCNgrg3QFc0Ib+RbTXx+Q/7Ab8wPM8z5kdkSnu4IHib8T9u3+8
mwoXK/U2LB4TiI8g1oqgpMCiZ9rRAF33T8rHtRg9Ng+DHvcQrov8yPQiDhfOAUi1OLyMzmjy2NIE
44oxFgEhxvq+uxnMKatDjH4IEvJjDPLbnTlMY7h/NbNYTZfJwKe3jQk4+/W1rf1LaZ3jQyR0ljGp
vH5oFu7ybK2JyysKJlhgt23zK4rBflO4al6WPOvFCodgWblaKXi9djh2fP1q+Q/ulGd63gLM9RZH
q944zlNCFqv6mcuHv+bjtT6wb7QciuEt2+hK3inMwo0rv8e/0Ld7WPOtm9cMWNC01MjptY2Wi83B
AovXYng0JWwV07lzz1RZGoda8oFova72rYL6cQczmjeUEcT4AqWTK6dqhHrFwdihoo/5blvMOrqZ
PEjNaPQU09QxFtWznQYqWr5SSe6w7yGFwMK7u4uS109Y1FQcvTizQYl9Q31K9E/D6JHrp1uzmKgy
416SZ52DjJGPPf1+Qrhq7TuKuPXq9cdmYRyb8HpgIjmJnxRU0FHOsJX/XdIC7dnKJyAeY52AYqQO
C6p+8QjyK5j+FH/JuPI0UiarzkJgKSwycOHh9DUDZaahtF0F49a/Hsbr+oGKSzUidbunbzQrERMy
5iixjZ5x6Nr6jiDWZLMETTgb8TaHC60+26XdUKtZEw6fpmqUlkA8k3Ei27k5GZ17morN+tdsYel9
TcKg3fcQqot5cDe+VDrEKIaCrwV/5lE5yfFv1jrAsM508b0N+dKt2Zei5Q4tjWETFhQ8fMZP/hkv
gHUsNsbos5NpNOriToIRmyy9o/cQAEttT0E+f4V1BpGmkISbZHKqZlPGNAstrUtKuqjXGX0dGx5k
D+uJ5nAYng49Tw07CUkQW44FvjYWGqsZP3ZjcFIC7Yin6SFrI2CYbDvT1aEZC+qdDJceRhXVdhBj
4W07YpemWcyHDPuU6ZdMQxyR+8FMIGPZyG93S2fB7bRd0/Tksu5+V2OT0qC2BYMCwt5duvTkuew9
zxPJc5rfZ0GvpnAqk8P2IxdkYEPfpAX4yRYHJYkUKQyIeOYspgwIGDoU77TmQRfB6GWVht5iHmSG
fNH7j1XybOVB0GoJx0sigCXv7Exe3EPxZnpHWF7X6wnS0YDwK9RhaQeIGsBwLi59CM0342CJnMhr
P8/pZTaEUu/XMuL+ZlNrDtfW+i+b4xThOw5cIo+HNlsmxX6st5isflW11divoEyqVc3pjRyLrgfJ
djV+5VdYU4gP1afinxetekqbc/cHyDQ7sUYwiqf+8i/+MsCl9vP/ynu8Y9aTn10dLZydRKcnqZ/T
b4p+rGRVJzlp3NQk5QpHnEu0htkUTq2Gz6LSshh45L+wohvPZahdBBRvOwcAQkh6q4XARgtA/Pm+
HWByEjEEy7gfsKVIJ1vruNcpiA+NdwxbrwIuzEk4FSrM3fz7Gi8KgQ29nl3EjWmfMNYYQX2fu9fL
duifzXZ3sK7jq98Q/YdPywfkGMs46hYrbpqUage2a2f2yxqoVG1GqYUcX7pk6gUAa6hnFNlgqETW
mYEEgOWeSuimSSkcAogwQNWnuiP8GPPdZeAmwi7jRlcRMiAjxzg/XFQwy01ejnKa+libJEnLUX/v
IhgcE0a/nyViUreyBusYR6Xx4xxmnaFOM+zZDMBYgqJSMuMtlNf32IbL5B3lwwYLLmQeInBseMXe
301fzoidCBMQA0aSmFKuYow8Y9SE0KiTaZ1GYExZKtjkjYeyxiSr2RUjXk56vv4eIomltyCv61wZ
u1spXueO0ZlVVB7MAeIZfisiZZs8cZm3819snpaYQYaXgbr96yp+7dPFVUvBtAlQYnNsZbLH2YdU
V6x2g8lu1SOtHnIkiy/rbyXR9m5zabg+e7Ju2esvXAuq6NdTXzqvqIe3+uqkN9lljc7R350K8LeQ
lap1m1XAf7aEgCyPrpcTDbJBBDMCe7sfXYR331Js4Sz/UmRPU6oRsD/Z6czSZr/RmE6jMWwYNQmI
x/BPkoM59VdkveR9EeanPRV11KKpK4WZyAQEmWxS8uE7Xm8dHdiDlidgkYQtcwb1nfHownvev452
LP8afqiwRjIvhfz9Hc8/FuFPfPSgMH72nocBNMq++crat17gaYIhWhCC/rBiRXBAiP57wCPhdVSR
pJuzzteNBm5bF5zLPxpCcukECPGMbPybtuK/I2u51Eafg955koSDZPkjesHtwsnIUyprZAQ7VLU0
jciGCSf7n0kMXxEIDXEGczVzhc9j9tBVW9K/Lj3cPb3z3OzJhvL/NwwM+eY1OBLYmniOEYhKsXa9
PxycjC28P+1CwAPkWHPv4h0240fUTYAFGrg5FYliv0q8qS5oMWXGqUD7rDeDZoyN8tpJrEsOEhuB
lYYWDKOkgQJMjoxZcewZKAAd+V6rL46jGvTJYMIiiMZFboHZSPiG11J8LuALSBcjhAUWA8WkVmco
uURd/mt7Ut2RZ74nhQKTfFOqCgrmpMLQsjWsDlIMoUVpd/uHwmf/x9Mm+F8CtgBLzdl+g+kcV+yA
RJvU9HcJ91jtAjeCvXh4+B92Jgjj280GQJqY9SpstXV8YhG4AsMpzHxGBHv16b3UzK/E3KjEQMcY
7/ksjg+kPdQsj8OVjXyX2WIQzBg4m0+2KwHDe6zeZP3b+Z3zABVDR1YYT1PMgJCTph50tPdB/Ywm
5QM2mGTrtJk0ZAPwYvrPyrKpQ9AUmufKMKUhw43mWLnfSXroU2MXWJ5D+PrnWI1M+cgtsE6U0bpg
8MzwCaPJxjnYn76sEWgjUb+4SC7Kes9T+JMbgxGLpH2zsSYFQsiS6euQS2j7dNO9Cr5A/d83g5UM
VQDn0rweHnCrGm4SdTK8idFh9jtXODast3P/d/XD1U+LRSoDLviZNpgaXXNIJldAIrfq4SZmeMmh
RKHLLhqErzEcDaKDo8I6lfgMzYNiStnEqBuJSG0x/ZfIvfetk93iK93DDpTuaf7Z/6CflQa1ep7T
d+txFKJYSuo47J3RQoNDpbAc6ElEPZv9Z9Pejupd4PbLSzX9GYA3X11+mhrwk1GHzNQtcQib5z4J
mDsRRncsYcMI34Qw9b8p5UphSHjvq0OcUnuGR/Y80eRYZiggwT5SJyc67Vj4JrF0iaySBRZlTT51
pB5Ok8BaVzP5SVQJ1/RwPguXnyfasnpdKYLCOt/oCEPe0e6T3r+Q64PnC5bJ+zCARD9V+6jiDw7H
06SW8igvjjMbPdoXPzmMS2SKvMmU3+XqGbMq5o9QuRffM3ePklMSLrubcHURBMZfiOykb5WPvsD0
Nmeqgm2YAcGtUfT6/+Q1w2sV+qNi9vA8RUZ8Xfy/hRPgyL3inkT5Q7pQhNAhnRa7e5J9SS75YMWI
wt0d5Ck4K3hBuQqMgnjR7l9+Aiqe0ELyzDWnrMYaSa6GZ7bCymtfZ6ey7Cx5a93Sa1gam0bZwhbQ
D+KiZ+sd3fMM9BZOKPnUMYvGCWo9KRhmNmkAdKC0B3XCLiePC87MARI9CcWBhfM2gNEHN08XQBo5
gPMmXXcD6JTb99maN5FPdUHCwfLywXWwAzPvhKH0fjtajVkZiSFLpHKjqMMDhbi3QtWCafn9Pvaj
XGpptghM2Uq6uCvSS4Cd7IkAaykF7BF3UFJXtCLwkDrQnpkVTPalqE+qEGb896i8T+AqfztsvMuu
WSZB6BfGyUAsGe3N2AUa7eBSIfH5rPEJf9d8Ac4YcvudjxyVvIPfzs1bImDy3PvNoHPIDsGG91Sr
VdQmdF32c2owQMbTESMSdHfjGZRGJu8Bylhb6zQ+QfInu0yJ+qTzw3U5rXyISu9/WQpNrHT+DOdL
c0B7a98dw4X7MCqXbX+n/5uVnPeSrlKEtqaXFkssHqgypEPDEV/Thn/lr7peymbRTk22GKIcESj5
96dy3kb5GXU3Wvk1YCS8gbhq6Aazh6oqCVwuYqObIYx+3LJ58xWSK/zli57wFl/UYbvseRFMnvA0
yDgoWkwvbnF2rFj5c5SAuQplVatgaddi8u/EpDMLZ4rmBa7jlhewSDBJCL8gPbVLfIpIyUDcDZgi
VPdNRZdVFComuMxENOTzm6c0IWP4Yigh/ehhNs7uBpTHEkb8YJuvx8Bmz+AJvfvYCfg7tULcDxi1
zbDL5eeSQM6mAq049B2hKDAE2syQo6/UXdcDP3r5QZ92DaLKElKXNgAaiN4x22hPARw1gGQ1oCnu
+LQlnquJwxZPnvMnhsg03DpawLkz/pDg4m/AbcVEzBE3UgPBy3GZN2VbWNv2sUVoisExkHb8oiNv
Zn4c87ON3Jyg9pVMDT01SbyYWoUhw0DcqHiCrf+dUoT7oPTbryt8MYtCGRlNa4OOTy6wXpnKQMuL
e4Z3JUbTKk158evW6w0xw55X/V1+Gn/be9gInUVXebJwHoLBVymEvH9D46vmE42ShRB28A4gONBi
GJJO5ogCJ0b3UM1M3p51FE+OmUHm1iEeYzphPYXDcOXXEuuPeDACTblto9s+Q4hAOQKnfVlO5SL+
e1NIZg1VbjNCWXvnfqlJdf+DMb3eHpTQyd7XdtE52ZgZ+ve2dR2rgGN+XCgKY3HUZ2FHB/uSZobE
y861Q1WFjqoKB/WCWmtpjy0Y9SRs5J3HXcjLxsYviX1oY4afubJfLBbPJk9T3h2JoTkDH/stEs3y
rMT8DjlbUH/v2OGQmk3RIHsKOt8+7huPDq70jUfGgmC5Bo3aet3vXe4owq1Owu4uYMmuZnvcXwBM
b9P10Ftu3Xu4TQ6FA071tTyPZR0dZW30S0IFH5zb2gsGgGkkddr2Sr690H+P3RqDYfHGz62gq3oh
qSKLbw6jz+2DcIB3grgBYUEpUMx2LFCSS0IM1qTntA4K+U7hUmxd0z4E53xKKA3fBfg5VBKwQM1T
pYv1H/LnWhiDuP8H1CefZe3Q5znolL6sfcuFgwNbHTkw+WflJDQGv09eCn1vS7jDOvJKH02Q543f
K6IUdoKynzmzgo5AG0anjhiOm3FAiXeuEfT7jWqb6UeJkn6yq+l2F/uPTBvEuXXmV8tMsI/9FtxV
R0HEhOd0ZsT1kDtnVGrow/mhcy2lxK/ljINmzohosdMVACj66r4krVWZfmZuOTwBTIR5HwHaQzQe
Filsze0aa7vB4RzsjUFkc7Uns4yXmLOfTXPMBZ6f90/KIK1QHj4D1NgAt+7ecze4HsnaAr23CXFB
GixPkHeMejwOOEAbd+nfFkK3mqrpSrLSEcTR7BzFE+suo5qwTWZxPnlidwDY80KXwCbr7l1HsT+2
ApBsiZe0yXopyCbLhg2F2dph33Uv0cdrsQgCoVKjmF6r2ozIiJKXf6agtDkznZwyTiROLZICpwDl
VHiJSBAkDQNid7pTzyODRs49tLtW9ldO0IfggYE4Spyk0kP/IC9L+dn5LRn845TWwkBxCTqi7ONF
yQfuY7hVhFkoqgj6s0o9Y8EKQ9fvuj5AQVbS+Lti5P3YbD5Jxbr+3N+9oaXg84mdO2tPBp9oPPGT
K3w98b7LXJk2wpPqYmVjLAOM4k+eb6CiJjmglB6ehcU38fWmz/kl7wow7QCACE/i6U+3uDWToKcw
8opdWA7Su/jn8X8pLqFDMuURIZAjzJOa9NrW+lMkZkMetnIVC7b+2VSU0YGalhz0UpFhai2Nv1r5
i4HL2JJ9+9fwBV5lZ5Bsf39e8H+/b8hS4ej2jQoUEIn7yWr5QJtjJuZW/p5SqxJjb1fVFhjq2mLY
tsLxjlnA8+MvMyUMQzNb28Zy1TiAid2c6RusKqiPyqXGwAKDGRf2G4YOMZcUp8jsuW43J/BUFhAo
H+dXYtMkRuqKez2iZO8ktVdgLO+yXzD6jU7PHATCqI+BSdwDn22kILfW8c5dVrTmO5r1vdkI6Ym/
h0y/BJ/hfBPU4P892+3d9h5cBw7n24Et/JVjn7LzlOrQiVgr6wC2RPuneftPSzsPcjPdf4Bd2Cpd
IF1SJx7o18N5Cleltlgoa7VXZmo6vMLpQC0J3QFa6lPjP77C5qHi+6GxelLgR8RPl6pzFU47kca/
Y+StDbtiZWlDQ1Ax5redbeN/GY4J6qX5/9bx229XLE0ZF4b0Ai/UxOdLdJrUOjDsMMRcSH3Wr2Sw
rGk727KpwDfx2orz7mJikV/5Grcd/Vl2TOsrabld736YUcBy1kGItDCcV3cP5fxC09lb+TEYoqsA
QNg5KNbpPmQK/aTzciT72ewp1TPDqODAzrImMGM22trKvcAYndyjcGvIwPN5AWdyd5z/zHfH3T5q
W1RTBsuHhULpA9HxcF0B4kMkTZ+NZhEkFa8ZMdrNzvEdXzonXuBSo5Ffn16unw3bMW8hx8OXb/bp
SW/k+anaFfHniBc9s/KfpXzJ2gV7+f9to3gsseBsD8QJv+DWURnyKX4pNT6BOmFZclxXSSbo6BiR
mLkK2Lgcmlz8kMe0c2Y43eQh8s8Y76wBRU2MW6ods+EY1d+lTkb0PCZbWS0qUL4Pry2FaCt2txx/
wU1xpog0CQRf87D6Zm/Onh76aFth8rHh1k5NTevgrAtcUJjWYNyASonZkQExcTeB6s2DOoMYHcco
4kZcSrxpOi2f6G+m+M663PTkR00W+2B0zfxwfdZueaK/LtmJJWUUg7+TYiGyBymkJyioFDV+eISO
6Z271mt+eZFxUYIBxGVBDlHE2sFMxYY7PSN5KEkH+eb5ZgEQIflytmvkWGnIr1HtmIF3vFoap++f
Hr6CQG6foIFamJD0ZXdaD/R2bnDpHN0FwBvsmbVR0FA4Rz34IYPFu9SWtYmdJNow7D/LrBx8pPT5
py2XyaU3YNRnkFT4M6zQlpRHfQFNcB5dJ+pXOgFlim9oFHFYQ+mlskRAN0l1fsIDmrsCypczToSP
F4+RBV1v92hlkKxbz2i+XlGVprSNibqEt3nIdVeXktSHOnzzgz7GLa0ufRc9z8Vs1WKwnq7CaHZK
trXkNVcjWKQww11o3xuv4l2J/ZdASlT0AY3P/AR2ZHt8XztGdL5j54L/HFVt6HQjP7jONjpJZDRW
hQe5GTmpP20O0WwbJEE6AxR0A3K8qs+yMiIvtIzrxvAb7KpvGDZGtd9fxLiz8/Onkbz1nTZw/9H6
PNieBc8DPjL20Txw+EgU0XU6+HieYnwWeVp1+S+KmTVoLorg7XFsBNPELdL2cJfa0pXdsTq4l2M2
Ml/XwkkVSZ6dpsjGVHs5CBks/dxqFZ0kd2UisSWhkAKyNN5S22XRekdfYRvEX2V8550hAaqn+nTC
blJdU7mv1CnsSG7r8WTwcTwGg0PDTkbcI74pDirOcoVBoVyDjk/Im1Ik/zOMxDHXKC6rqFfPLF4x
OPANYqNblPbWaJmCO2wWG9cwOG0ySyiepDR/B+nLTIlMQJ3ysI4PlBNrahMCxsup2JaMcvzuHhe/
TB3AJBCuNMDhc7EeE95vYzoeSVtg80+DwDacQJOnPrLyFxsNEnVkUZ4N0GAQCshe15aq2zCgIWe1
/299RfneK/yTx1BlowyTaSsM1n7z6BGPsX+dbATN3hP1NxMGLh4NU/ayW4g8RJo2+nhTbImP/nCK
VBh1RxPmrE3g/gbgA/dz75H9Gkatknlf4PzOAPOf1REmpgTCZKx2D3D0pO4PvvvexeofHtV1uyop
vrb0cYIftRaHvZXLuqkOief8Siwjihg/0ycT+6nyA4EzXvO0NENpR8TC0r8rnslFn29tnIP/uHUt
wns10+YzXoAFpASDSclYS5jPhXNBJa8UsIourQaynyukz0tNRqzVlpqGtlesq1gcsjcp730zSjyh
Jcbp7CLTjbIFvW8KUL49U/KsbYp5Dizics4Nb32Xw9VCrNL9WvvZJ2py8+N1N2xvF3UeVfH+9hGE
iznXFeWYAvHxW5G769PxW3olmT6Dh71O1lr+ReaLSuHZIs71QpGqa7fwU0Y/UdQKVxGJ+1YfROOr
CoFWUiNmZe8l0mf+dhjydqezbaDGtu9iOnZsIHBKPzWGgpl3QoA6TBoBYsr/5xwodHXKyAMkK9Ab
cBRnBBv1ZE7SPc7H7RhMDY45AmhZX5/Xv/oSP7w2rBHFdQiiKRRfesy0yTJ0H2SAZL0SO7St0Z0l
fm5nAHN9M9FFERCv++Tt3+pHbZYm5IKS3NiQM+aw+D2DmGVGOisqtJW9UVeg7rb1pj8SSv8srQGI
iK0xuXKQsvQW9H0K44roylOgWMUTI5GlsF/qEMDSVS4+RCk/0toIHvwxIbn7ki5XxPj5torMIQsS
oMuxpihRD9yXK9pL81bNX+H0S14iLS/rQEsbPSj+SbjzDcJ+eyC+Uajy7P5uz0AAhly6SX2VfEsA
nUUly8o/9oRsBR2gWpLscHyUwsudmjAAf/DDY1oetkjhcm3XUWgMtYC1HkRWyVc3xhp2ucdtkANF
EmZetqjAXqjHj12W8cyVhvUcjLLsRYBpP3ESztgMDO3ZsZ551T5tvTuBQoPL5pnV2HVGnYb+8yLV
ETrPBwb/iqO4Fpt/dv5vc9PnppQgei6ic93+NvVxT6/egvQtoO35b5JhuS2bd9wA5zQeTlGPuz9O
JIDW3J9r4tAvxhUSKEESIOiFMKEZ6T0n1DkyvOjJX5iO0RdVa8+4xIsQ3LqfZKbd8WVXOP2FDGck
c0ZG3Qnr3VKZ2kpZ6J3XGR5Z7pS5G/rhWIA9CsxZwdtWJZK1cOEjRPm2V5VlHJIn35Bba57+8dr9
0KI0HDmNpqxRfpRGbXZ0I3K3PRsLfWfernWiHSk+aKgZ3Um72oXybAKAqBAldBK93ZjmLmNtDkhe
4mcc2MPt4lgLGn4qqqghnTz+Av8w6cu0C4bEcXWHh1tgMau55G3I61988RwnVL3VyaXRHJBeykop
eUsF4GANg9ckYvQOPAtOknET+8q5AVlBiFron6FawMwjkITn7fDPUJbU2AMdss45c8DCQE8WQHMn
xHQAVTFhwcFn2ay+Toq2i1zLcKZODQVo7qQwRKFJCJ9wPp6vxR2qIXdu8LuQZaKEcmxOU0W4smXx
nKHkydzRRaEV6qe8EI9n8B2tN5piydzx46Yo6QNlB2k1z/KlvRk1i6JV7DYSIJCLHrXrmUhDAnFC
LGYebq3qJNGpSSecVKyOxbRk8RY4yi+j8HUQqTV6QyCoFJeULS8zIxbTGFLauxMmyoHkC3q5XK4G
+cxbZxs+LAkybNiGDTra346nQHlYirc2k79yqU9ngpYN+R/SZqDur1Fxl4qT1SBrHEObQuaHOTsU
psFYVQXoFf2Y04mswD57R+V2twyjPu0NBpbVk2CqxHjj9YQSiY50P2t5RGH5Tdn5WEGpgoofLmoO
3YooY1faEt5t13ZeFmEP9i/32niSng4n5nsAvdD09t8FcJ7GbgcAk4Mf2pbPpkFKeCbb0nXUQ8iQ
f+GLp1hpuNXy8ZlkcBIYi8Jsy9a5Oa54hQpxTZ6rOq+p+k6b9P1uk/c1iqTQNDDiKKkOmp39eelh
BJ1eeuXhnJ0cBWEISfR6NH7BWQpE80GSZLINORun4TBBDII5moo07/fapLtNcd+Pvf/JqjZk2xrK
jWjcLUaUCpf4PlTHCT+JfRCnqVGUtdOIDXmtC8ze9aDptiLQ/D7PLaTFawoJdIiJIhnv1oQiOF47
xHQj3HJYarWYw7/6D346Fy1IY1rnlzo90EluscDSNiRjEtXvZsvcWDzGLiCKxeTzGd1IVBG3dyg6
1KH0oW0cbmyRqCa4vxecW+UD7i9oCNEBCK30cnltB+2eIGewGuhTxNe0YoR6AuHgRbd05i8Tl6WH
18a+sW9X6Zxb+6eif5oer/n4KWRc90qMOS2GPPRPfZkH/Z5NdKJ7+ooJNhoBUeZ2D+zfk1YedVJz
w+4J9tmSSXYFSe9mrD/SaZn8oh6IxV8KpEBsXivWeeLE4EycmK/nHie9+AVEl+GQFqzySp0p2fB3
HVPr8qlR358xMh25K0zda6dDWB3Jy5yejQdWqt9FuSsa2+SemRGKapAmMXC1aBXcZxK83UyDXbtK
5kkrJT17sC6OjS2Y8F3EGrwUNrDZ2I3m2TI1UCKSJwL7ZqIzqSn7woDpXYp29UyLDuCFVCuSHo6j
0YXcw9Tm3zL2fQnlG23TNRmMBLJVVobL5/Q1qR+/nAz/ZhEQFjrJg+rMuAx82Z1Tu5sPRBbuXbzw
+mgVmsFD53cgO6zv+1EbalfL4/aNO+C+MMzaywV7n1bbNx6MX49YABZW3BfcUzRoZ1Q4fmb4GSro
thitEEfthoCcyTxBhXvsFcdZmtbyCnTVNXz6w8mQFki8kB/Zb3V1QCPJPQ+PH6zqhor+i3Hslnrp
WDcd10PHhJnPifPp6/1kzYuNIdHKkM9a488VHEI+IVJiaz580IVL5bgQbwMs72liejEooAWDcvfM
fU+VeOEZVNqMZoxH/wMgEJ7lgcoC1uXdpCHZyqXfieFPJGPosZ+ZG/74H11RI9AO2gbn81Hht6Cm
TBPqkSoFn3UOtPaJfeDc9no0ozjnhamU5L9H8NJ8cKT1XKU9sHAPXiPjOuvH8DzVpDfvSe/yndZI
q7UUUfKl54sRIxoLzhjoeBDs8SpbgsTaQkqVjWaQxfTsFANyyObb86VXKnyY/UVN/LbsPVwyFHCc
GtjJMQzEXbd+Qx7GBGGLQEAqnIb9Rdh4feioIyBsN47sLHvC9BW7bYGJkPQFw2O9G9tytpRNhuHy
sZAKTn+9Sqfh1o91yyfrJn8Z38qtH/K4oWz3YnfsrnLEjNkfJwHWBg0ZXbObznoExNkJkMRxUaWj
pMEFMO769kdvGa4WDyzLaPIOJD104p/b64QF9ymKtTMxlXrXFYiloiUvRB+108ZaiBDvpHEvrEc3
wJ+aoL7wy/+YB85LSNSXn8iTW67pJejsWNAmBoWDHhvfFdkgoPHIfpXKr4J/fKO7r2GwjsyGZt57
3nY2IulJsvPogiFeK9mYjGVx8zHA08XmHb1uBbUmY8/Vkf1zrGjOzZf0/yKUeMFBadj9nsa0jiwU
5uVA/90eNnRjBkzFOVtMG9oGDIKL5i/agWMBElIoGVHH+IR6izQGLh/tYKsUkEtU7Po395c4umtA
o+og3NbPlqQ4anyf5V8y2Ltz0KxT0Ij187YMPOaZGMH1QBvbdapPfqyyPbfyj0DPVISAlQAtYA2g
V6M7a6SijNvQm1+IFBc8wPd61CcJ/L2atggPvO169iD0YhWa8+aM0ky7Td+TcU27gorneK/biLIm
uuJQCu1Jatgw0zi0A9SYtsJ0kXPSYxk55MkRFdkMuYzTm6ourr2Bcq/1EOupZcsbLAkcLVBtL0tT
JcUBQ2MgmDaQPyh21yqvX4fcqB+3xBj7V8nGjc290LOtA+zRLynzyLFGYlN/lvCBWaPE0QswAKVd
w3pVwxKHJLYvnyWKWnouadv+Pu/Qt3LhzGLhGFN6cac9rAZWswtJEjKHidoal7RJkP5Xjog2ibgJ
06FZfI7xVuxBx9F4UvWh1ALYLoLFRZFzk3SFP+UzwAf7jN3Z39QQn3PZu7Wv7trw1QKLqgyrFhDC
G5f/SOS9NTlY5yXGE9dPi4qY68YloOLNXIiwe6DWlQCMPae5AF90hvIFbOownQDMb7mOOgxru0xB
3yoAafuMBHj2+VDA7aotxAudSYTlsrCcyuPXh7SjeE5fAYdZ1jXhvRCbQCHNAk7KWkuV2yJRsDYw
MbZ71FZzafqFOguwleOD+1hCZDEHJnQYRvSu9FQVZDIowG8NDkr/9tEAzngGgz+LYh4/SLnixNdA
OYF4/KiFsHGABMZQBb3ssDHr/T0beVcbIkVRS9GqsmzwGPUyYs4PjH+u/6zFI5Ow9Oebdu5AIzBM
+RFKfpmqwRom2J62m/+nOF+epCYG+0dP2lGMmywvw0LQXZIi2kt/bj7C/GvyyItBurBw/HDvhvHa
FQ9XCjYCrhjK7ZEAMYFWcQCJRUHfiCdsBlnUnH9PWUrAlBwUisTC//y+TM7EGc9Jv2cnypiP2AGA
7DwPSolOPcZKgMIc3Hv2npUPQ+M0cft7+uzWj6qLG/Ma0w6I9sYwYkPkZiKKSmXtxqf7yMXMt//f
HTs3ta3K2Xe7bOCE8/K1ItgZLCxduUfMNFvXWBVm83cGS5VJuugRyewm8FZrV2gcoTnNdujZ1bFS
AqvQgAtuEH6X1IA9PwhEXx0CfEr5E5zxGE77j+W9JmdL89xXqakTRVova8/5dcwxqehZeeTaPQS0
F44oyN4MhtWFQxxKd38hOsei8341LCfOjrNeUPRES76jN/MAQ3xTrSV1ZJsczSwiNINZQxYl/raf
sJJCBaP99w/HD0zwKnEu/z/Gkx83h2xuBZJ2YkD8UfgcOtnujb9sT3jlMpo7UPmo2hy9PH6vzsgW
2yJljKYRXt3yGJLQpY2Zwzih4OsXF/wjcgBGg8vO99TsNS9n/2aXeZgkh0hfeSV7c7EdoMxsZ18d
Z6eEoKSTZcGG1SkW9pdSDW3G36CcQ1M9dxVrY+wvZ6Wce3zvFG3txWol0WVl6YQ+yfFo4pKIkpHy
X0TbjTV2nSfVQmkvqxvJw2Qh9dQWEciuyMRW29mdTiiCmkMsKE2/V/qFJ2e8CYdkaraHWhHEd9Vb
ajxzhfBnORP6fX6ucbQmsm5QtwRAHX5qrjqh/yCHK8huZwAnWF3Rtw69K0Yq4Xmh+TA7cKgi7eAW
ZuCvUFGSMj+jAK+Xf56+z4qHKGc/DmuYmgwjloL3B/y44iXhkg8S8xCV8UUgq+ZOXfaD8hBpzc10
Z2qztlSSLybjpZvBFyIgA0QShKTFapmYivQPLQy0A1TgyeiyFgt3EBf8z5VU8gw9N1XgBsqri+Oo
HR5E+dbQNepfw4wcayj8vPPdzMKqqFJtgGrzC5Ef/hjDNg4vGvhtXBrjfz81tK6GvKfPmPDTz8DI
dFMUiO/SvK9pA9F9MBsEOZNfgQOGh/X6+BtAMSX156B5nE62bvFpQJDPJKIT5Gmmh+etYfBXPscZ
D3uD0EBNmajQOlQaEZSPmgX45rDb8EntUTXV7ab6cn70WOB6/zqC+gB8g0RnxYroTvzxwhTudCfY
I5o8hXGnlnCLkpHpSihL4pbY3Bq5bfRYNWMERwGlugk5drQv7icII1Tfe2bH0BVx84E7vXpjYnOe
EqYTx3u3inj7TKyclCRr8wfIlzjxKIogmjfj1CzSB79aTtDM85At81epxFcdmOUUJtdy/MvP7PH2
4+pzbGWRdKurTeX9qLz+lojjUn4GlCxoEVMVoVvJJ7wYKGdK4vkgtP3LR85HFFrs3pRKIuNgVR7X
hH62v0OvRtHqqnHJA8EyjCARf20jVQzLklDO7imDg9W3xtHl7jiOTJsGHpWT1wAH0ln5CMJihW+N
MgXpJPLAOPGPyNXlU2brT6zdrLv80xMpltCfhZlzsrOSwN1A0d+yFINa45PlMoSortAKNhRU/1+i
0Wx+VYl9VORonktoixBfjXjpQoTrsLOmjR8BJwbrJ2lczRJvXyjw9KtVV0PNZvsOq/mNtcgvtKR/
1uRFgPf9E56X3Is6T4HBxxwtwDX1ROSTrxjctEHXyi65ZhAgTsW+DnUb2oxa8g7eRcw5zk59VqQn
44scE1ZQNwlvaBxiGabsXDJtWYRRe+EOiBeGw1o+chehk25ysVS2jkhTe/g9HxROfqKRFpCZZqoW
59SzDdWQp+/ycjpc3s0mosW1ttLf0DdDRL7QKHD5qPwHnl3Rsc6j78npjNRWQshtWcNyZB/5c/m4
1KU9O1RfZmHhiibZfscKPpikj8U7GFuO6lcUB1TSlef41J02OZx0NPGQ5ulvoA3QB4K+t+7KHhYO
+Clp7AV4rDCueJcyfpNPBXJeiVtIWDUqc+jKCov8Xr8ZITa6lG2Qie2Y+vhCelicRB70VJRPfebK
uHdm6tT8hQ8Gdh8UR39wBCC2T9gPT8I7iyaALws2mSGHCH65XxFg1qjJUKbNLgyias59ZnomCWU6
PbDIu2gp8VeUBDXrQ5Sl/NOU558e37R1Hzn1HrgiqQZr0cTZeBmbsT6KERaGyZ94T/qJEbo99yUW
nSvUQ2RrVMqAjD3mOKLqDjQ+nm6LvAG+zMwFkiY2wGpl6CCkyIPWu29Gta6LPsh46+ZidhXCWhXz
v2M7Sl+/28lSHXASGacPEkQx9Vs5Abp6TZo7/qzoCLW3fM1qJT5qwC4LETT2rAo416rqoBsf9V6F
vc4BBAN1SyUupoHX2QSHeib/z4p/IJfR5cEBUtA3JE0Rt1A2vixIxiZaYsiaf989IOFsbtP719rb
Jwv15qqpVhWoRBJUipWXAqo6+SVl8AxNTd8kE3czaX2BX9fjaJ5yqx4rTKxhClL+nndxSsEghZeZ
sstHMkkOW/1GibuEs5xWvoKHPwjufVSlZqb1FJQc00MaIKyGVuzMyUheXBSNlq/osm8MyzAajMV0
cTo7YP0RfedaHMKf4dQoum8J5DXNsj1BLBKAKju7B/2zWinZ74BS9wfv4ZCalNMdDivUp1Hbn65z
VyHULfV1v0srYovBfQnkmaBOvxu3GrZtLhdSsZwn0kCUhWC/qH6uN8qPIf6iRUqwCsbkWq/mKUGl
9hAS44mAoe0heRtJsN+DYX5Ry25RQCnO24A+m1g/0mE1lWQEHntb1zhCLEImC7hzk2Vd9u75aHP4
BfulJ9uDSZcIbi3lOQ/RHdYIln+WVv7sKPhh/jaghO+dUrqr2tKoHmWKo0Xb5ncIQnMMy5g3XYMO
67bCZFMbvHu6QJDRHwC8aKmFOiqIO8cvPLng/SM5UjPjAkqFXfqqa7v7LQRWulJlvnm2ZZoZN5yb
/DRMPad0lvhYGu3YnSLGwxVtf9v+qR1HW88n/IBZHFogNp8OTJDS0EOsPVWO1H6fVGzrSWlSgfqd
7VYBcOGIUNalQO8pX+oSmChidN63GTMP93lCfytuye/71UJ50E8YgaHz7tBWrX7n5QRntU5HBdJ6
zsnbnAF+yqJl7OX/c0G/qO68SOcOWCCIKWxZVRw5BLIYOa7yGQFD6kMSp1F1cGyrGO3aolDNo5aw
7TkPDsNb7TbiBhvK8rEkyPHSHw5K9myTQdIjq6TB/yDi1Iv8u1WZRCSK0JapGOxlgBhuaK/UkTBF
hrNIancACJ5VW37Ua4Q5hgE+u3MOjRsuCDaVl3+FvQSdWJv9CFrz6f99DA4EDWzHmpvyNy06/9Hx
3tNyAt/6wEfADIFiBFy8v2I6f7iBXxE2AwI5RjYkQdxxu47ATV9MIadG6JxF29QelW5tJkPWkMJH
YCMjDlKQUJDd4siZwBXYTFaRVmlRyumoSoVlISjj9SyOu+vWz38cNa9T0LSuIasKNIQbMrbxxN2X
2+K6k2E6UMLPiBXFVxmksm7ZoWkLuFo0W2rAf/e+SlDnBopeRPtKQA1CV9esiPVtp6oB5AxC4Ogw
23XvqNox7M87J0wKGm4ci2wJTIy+X8mfZdz3hbYmMN1VlZj+67K+DPqJMnvhqtROwrOleOMC5Nbo
Bvj9Kba7asCVEDJg2QOR0cDzqulabwiUOWbl4gA9hOo9DD4irKUV2X6xr9KD8/WdWYnH1m1u9pxO
vo2+9Y6IebGNh/epiEYWKDtFINiSVTrFZN8fndxDjDFquavsQvx6tHNr1mAKMfvQU/phdgvXiY/0
RRRSoZE9p9ro5LAa79ugPNOAdCfUcm87PUvs/S8ZO1RdwQrMp4BjBHV1RATyUvfB13Z+1hA8aka3
RGC2hx9ItA1ozm63BLzDivxavwNz67DijvP9X/tl9+YXkUs1krherJB094x6b/f51VfxJ1gBAT2u
8oJ42ujga3eiKKPC9KttjMZmBdv21Df7dOuuQ+666bN2mNWiyuSxp0/KxFLetYlCTeCp0s30/NPR
4XC13aqpmsUSkZciSvfT/fN0P17/typO7neTrDVSuRTYsqibf5C9WQ1/nYl3IAC2LdNy6L4nLLng
kul63O0WUmgHvPKJM1Hd4DLxdAVZmOky2F50GVtKUAkbrdDvpmt9BhfluHrSZ5RMS4tM05XN1BoD
CE3P4AU2yoAA9VvkO2nAqVjRbBkoSYY2bx0wbB1pFLBnsrQ7o9IlCxR6c3g5ulEz4FXdnckvJdjA
ytZYo6XZbaDTCcNC3R+sMRxo1zVubOOo17ZeAeeBgO1cPlEJlqX9Rjw6AFd77kwS7wXE7oAxNjze
IFcLkRVf/YzZzA0JHyQjIEZtmPqDBhozwQv1jYjF99xz3P3l0XkitBTVWrpsAOPVRI37sYeFYo7A
Ea/Byj6PtbEPvNmGW7y5iSRBXuwt1KSRnKFph6L5Ok9DBs4pi2gevPItBJtdg2gqvhM9e7TwzgrX
i1XrMSs5Pv9rfttMQfBfh/SF3RhYd8rOz+zBZMh/HcakCo85Jhno8Pof+XEWf2nWMJr/j4HQU2x0
0DjMQxb1KKlAbh7Iqguxk45iptNkAOt5RX0C5qfrKXBUiYVKPfwXOKWO15BM76kN6rmqbb8RKY2u
fDXwgptxAZL+VbQPD2hmchysuvPkNcDIVB9dHZTZqDtHeq0JMDaoHXsjUUm5spTMv31VHEDcalBg
BUp/r2lw2IR9aFrSf+xbpMtPMTnujUsWmEPBTS3IeOPR1PsGJ3F6EiGLlvRXHvorfLxqhEB8tszf
t873l3Z5F4SFZiMixCY9/cogUpQPp26nHMix6SoKcQED90P18ZhbUUaJAN/r4YhXY8FJyUv85E0j
ajwsCGESYOT6hQpQhejwkTjb7LoPejqmvW7ENDw9PrRUtHFKIXaUcunHiMG/E3Y2SubDm8fsc0xP
AgGprfXiBRkc0vLc0Gp5GdBj0pxSTdFcvYovuXIdwlxbZ9YqfQlK/rf5yhnoSZEiqVeoSM9ZJJ3h
MRhPJ52E53zoaFQNEmJmCjwzvlT0D3ZPTMXReghbhnhKdJ5u3UPLXnA/vwbugKF8FVJbKIL0tnLr
6y6fOJFNBHlVumfcf25EWze8w2kexQgHZOIi1s9OThNZnFvCBs1bZRfI8sORGZe3mM7VasRUo5YS
ylRIOovHt27aDqdRgVs5mhSydApy7SksZkTxeXY6vtFXy6rpJEYfjUNzGsdUyC6emVKPoOsFDQUK
Nxt99HLhMIS8wEDd/OBm/kEdUK1AUpxZypqN6Q82EkJM1JLrBGBaWh06tPTnHAZykokqDa4/RIP6
TMM9C4aMI2Pri+WqQTRZaCXuIxr+q+FscEde+2O+zqYiuL/2FO4TAhQKeRTRFT3xsNUr1TJfMiQd
yKUxEHQ59MKzGuDHIPRKoG9/Ka/p0kcsLeqWclHzL0bQFzZJVvESiOnzDCYDXSbFaSuTTVZbM/HF
4UkhbdCgPbJ3AMgTlLl/or2beSWYJXZRJClQvt4nBgQzVPZb+cq8o4vrRYw2oiu7bguhDXi/HhWY
NUk8jPQ66vocn6IRfXRoI7aMZDeR1s6El/9YKwhAjIs0/D+D0v1kY9V28DSCJ6PThFHBPBFm2E90
SGm+RH5kZ/qyQAwG8tJIxjlngYFj57u1labjGuJrKy+wg6r4sVgGXo023z7J88CzizaiRV1O8+/v
jSHOGZnL9GGSsd+KXAIbMqXFTGFBw/0iWEPAFNsVCmTEcEF/McwamSg8/TpQBJSHGXCFURaOPr4U
oc6xMHWK36L2g0kFQYe/ssz4zNkfBShElpMJp9pxfFwl2I4azPSuTAOpeg8pAhqLHOL6qAfjrPic
iFDpW8oBSSTETyfoQyn91juOYlsNidgZdKNyzc/hvmPHplYQQXH8JuFk/gZaU2Vs62qklEJX0Bxc
wn69xMEL/qk4ZorqvH71Q6W+Ou9waTvF6KuWEtrsodO12C2KsBaUFT8t6LnYyCj0I1Og7dd2mnES
aiUfdiiKMMFSFj8MVMjq5B7LjIJPHMgrLhOcrGG96ciIegnuAz4IhoKxhN0lzabmzZ6b/QYZGwZR
cRqajBDlebfmaYxhBxpvQk2lXuTNTMWtpgM9B38unNMSDxzSwWXXesQf77TasqPfvsEPk6IpcHtj
ZbvcvjL221LRaf5ooMbG3lZaG0KBgWBprKgs19Hqny836+9NbTOlDjp4NWhk3csD0nd62LBFP3Lt
qBorjU/X9uQX0LakIjoBGTzHMgk6fge67uqr9Gnf3dz8yLppB4CSTtV4T7j1py+uo9lUQattqUE4
9B3JQRls75XdHIK7JSLgUJp33KSvaAq0/kqjejki2TNOSZx2p+revuEB+qiFXOyVkjbTZSXzGqe8
j4ljyvgW8QXQ0VvTaQsiDeB2H4NilffPRze2KTp/ImF8ZCpjTEyC+ogVWeTR4pjvCSQl0gtCYBiJ
ZHfrVqIe2FWhisREG9NCf/dvxbZ/erTC3ctIhXvPPCVm4m1/n6Ky0TO1MP6haj3QsOIn01kIA67n
huMCEQITlFZBoEC0Uj/kX8mAavg+D3m0p5wFLdNdhMMf7WCqYC+VAQ5AUcSDh6d21tXF+gvwAdQB
OYqKvm7ZjTw/sWD8fnpOVg0kQ8Reql67IivwIRQ0GBfHPtjD5rFtxXD8GWkV8dXCH/oZe92WJz9W
foKXP2hFFoPqxGu2Eh9/ZdOcp0RpNv4mEx7JX1LbMcV7LJCp9E+QaneeSlrJFsLp9xL0wh9QzSsm
BJmgByl0CnEVwjezu5tAmUrJqSaipxi+V0r0ENMXRuLyhr9xSvm3stfEA3LwzzkzAQHIAOjGu4Ms
CcSDrjVC6tcWwSdB/2T+fJOeg7nh2vyTGr5OLIlHqHiZepzLUbKQ9UBthPA+Q0HaFfMZ/0IrSnYS
UiZkoTJ/kbeWETJSHMAgTC+H4C2tKl9WYzQY3v8XZ33pUAZVNPNUHmXqOFzBEnI2+CbYRwhUldQR
uk3HPJwUZdK/uaRy2ulwvGeEK9+CQbjKJ80xkrpPDXevVEGnx13haSFjEY343H5i6v4nkhQHB4IQ
XaqzduPNYbhKLkdslm3cZWLe83+3i4KOMmeklm8c8bmzksctUFUYKTNYXhnqxwFgZKxOh6ZApt9X
fRs60jTl4h9zrAPFcnmPPpxJvwE+OU5QSWstQwdPI5zu8XMrt6fsna0KFVFIAhcHGs2ok4XnZu5o
UQZ+wRAd1Szwqcuj3s+jOeKxgIRS33CMd4Qa1pQFZC5E/MpyBB9cDBWi9bWADRIBu1Xq6PSWABOh
d00QsaKcnucJ+YGZVLC8eiT7szjUT+1lgRZGJTk2tAP890F3Mavjb+i0r9I8UP2iucrjokVzIsPd
9RbvnIpv1huWms2HmcvXBFGPMyMBJxuiJznZpYR7UdV0IpSF+4BU3w7zOs0CFMiXt92IdvsbTTT7
ouVdSysIN2oYR6jQCkktBzX1Z4tysZmCzWytB+B9V7nPMLP5LL3VElOdKK21vLjd4PHK4h8zhky0
2FZDccuGetcnd/LcKkYcLW+ikq31go/1a6HKwXZep69tsdTiLv3SWnYin18cIIMHtIitZtMV85gl
Y8v0zR4g9B4a1/Wjhkm4RnkmiXDORnUzdiVuiDgMAQ969ofg/SmwFvTdee8Qpn3seFmdEfilOXmM
BQ9dXTpQUQ0JgeT2WafkkRIC6df0EUC32BM89yTUIB5oOlZtvx2jbNg4x9V2ELqa3GxBcpAh0viw
HT9Sr6SZhWeC300idKBfua/LBFvUt1GxzWs8kmM9jesx7JzS3gR9e2GqFtu0TnuHRYM0Exf+pjCc
kJKujXQE1VrHF1/xFmg0wkkWCdisOCYR1KWn2tuOgnqdyTiEgml+DsiZ37vICdFXA43BxNdDYklU
sKHZR/KQXA0FIyabRMR2uJFkSX2RM+W+BjpVtvoLHqkdDSY46GgupBb6BmibiyD3Bo9nlh1eluqX
JjuPxET3zkWn3sYkljqRPEDnkEBEPOlBzo0YXxPEr91sJvjO891T5VzM3ATU6MtvYndLk7ATacCt
K3l2MehuWaKiENfdJGz7xpV7+23/gYvzuUqzGSXQdj1e/cgHaOFa7Gm7oGxwHTD7GKGmORvljqO5
Pb/Y5c6KOlDzfnkT/r1J5kEEhcvGkQcCw+gxWijjIoMItUvKjZd63MrVxUYgTsXOdEkVALhPJtam
o5IOYzGS5ej6rXQV7exmN3EGU75wjhvKHf5DFEnJ41WrTzXuWh2Qr3xyp+CRwDgpc1m2kLcTfi9M
GJjwDGEUia6TJabZiC/WgFNozbMvLkMb/G6Ztuzn05rsJ4xhqY8aqSkROCdTIso1ZXkR5qhvEbaR
MXI4kkCefd7KSNG8FABmJ7OII67VV2JWshe3hRe26p/uUuynxBMDV0mjalkIqSQ1/eGhRsVKnfZD
+smdD8ridSlYpaiP8al+jPEm0aEidEsSekpVHPHJyqAGDjq3I/s0pxotB1EhuWLNkmg9nCL8urRq
QTQXlZG9xPIY03ILmKHrEPBubcm7WRDqKB3h60vdGrl51f9GBnat8IsRnVOcxCrQ6u8/tUgwn48V
gpH57CMX3NGEsT/ZWjDDZaYVK3Xh4XiDMgw7kyl8buCGyqLwGFpMOjMm4qwBsyoppgYbG3dgigc2
AmVcUQP9sWmHMo3iQmbk7lvQaRoD1o5YQgpr0kyYN24On2yWOGpcMyhh5VOd07dv0hv81fm4nWMy
iZpQvgbB6d9L7zGVLNiFSFsqSbNZReW8EwcsKklzdAeZa1MEII1rW9WtYmHLKwg9c9qu5wGK+378
ktwDPIIpkRvKHutY7kS4Pou8bJpI6PoPHLrjERzW2N1dpCUrbsFAoWcOkdVgOPKeBmXKr7qxsl9J
qmbxj7oA2Ns5CepgGheyjP5z69jomOeYHG0f1h1VT65D+Jm3h5DYdml4QSs8rYSmfFPJCR91xF+U
h1inHPDnk3wiG8EQSWEJVuo+T/cCmaWSs8GulYbtIM6WOMvqqLHw0zTWsJF5nBfqYNs6BocehKzW
nstrJMrcWfBv7B06kKXRvyRuxwCR2BJpZ9uq6toW+sBha0dA42sNhCfb4Ib4SX8aNjuq7NARY90J
MGSftd7NaTeZ1eQzZdP/jqAj7DBIT34XDSO68FNSGSZKKImdn4zBMEHXQ15eiyEsTKq/UoPgfogn
xsrJG4wbOvNJUkSUOQ9bX+EDdOTfyX/O8j7k7zNchfxLX3vCPuzzicQXJenP5BkEm+Pt48JVB1yZ
fZgPRasWjIXk2oySy83SQIYMZxhSMjH5NThsp/THX+so0su7Pa6gXBiCCxImbH0qsjpLhpDuyYH0
n8fYiZypldZjjgbLq9H190ov8VtrZTI5gbDi1glNcp2VMWwN2PJwXPUQpMf5swRTLb5k/KJ342mM
DyZnrNwLUMtzKt5zzLNHOOTQKYhvP23ge7q/tl2P8ZxCF9N6Zwtq1XKMFIC+ktH/ZYoFH6j6X5tC
EqAyVo/FfUT9153d9ssXvg6HIAmq+/3Et1+wcxIMSAxx2zaO3yht2ulo78OS3Hpwe6wbmNvgh3dk
aM6HDBI994Tst8+gQapqSWfbPxPicn3JwIGhUiQM9LZaiJOxcyIEdVoamk4IpozJqZKZ69PLoLFy
BVnjzTAaRiWVnEKoFp8+FgqZvSrjrxl54vaa+tkH/2sUMltNnE804YvlDLpElaYQs12JIgeuGdJh
rlvHBRgt3AjPyF0doPfFqUVuHkFcFkxHTGoBwrE62JKiCx6r4PO1ltVFmUHngVZLurAcztdEFNFW
FreYResWEpAvYyFsDdWvlQA7+uuPmn9ByUj3vr/XiEQdBo6/a02FjYpQN2H+PL1tcCVV/DhG0VdH
205DmFLS4rPDaX/GO+s2XDY3EjcKbqJ0y6P4WKS7uscu26odgUd+0sq4Y3Muz6SBPcXDksGWWap3
qqs5FzGtzdQ9/AwFHJAEryj0Wj5vusTR4IsAHV0P5QFWlyHDK9eYadvlqi5I5afOg8/LtM1TVkri
LG3tZbGK1Ygbe28W6ZJhRvsvgj6Xt0Ktx5INPr3UXQrZsYGLUGO4XwBt5YAfhBjYBUHFN88Qm0wC
gGW6JCrtOdN7xy/xudADipE0opeBGlGCUkp3FChtdOaxzoh6wcpiZFyyQKOkSr4Os7PIGeLZ/S3N
WcIeBUwCjuGhjEXmH05l6E0nJYN5MRzNuj8UeFDW8iGlfQs2YLlB0RAJ781OdyfOqRw5f8HdqoAA
/Wi4hKBJpB/F3+FhVMsrTVeLVs/wUWtvWG7teu2MC79XtwR63BK2doDGY690Z9KJIq2RZti8GCsV
9z7fhDxeVj3Cm6TlcuU65OUemMyR1CuAv/SXBXDeJ7LFH3hWlgZXgHz9w1rSGOYq5gHU/QWjNCez
6sT/LTNWZyHwVpW+ouVORtUB+wkoBqiM4FSlV2w4gG1beUpMw34ryaDPvz0qKJjW/BTUBU2jiMgS
PlBXVHQnj+jGG4dEkneSaMeZ15X5tCbwhVnYfRml9D6/b8BEL5IZwUKPIt1/PvRpEHZF6zZAjg7d
5XMfgC+FLtf9+a2gx9hgHiid7f/GcouN1qPHdCpy+IPmQYu8py6zzPT9fR7kZ+Ie8ZWzb2hT5YTx
M/6NocnXXXaeJXRANTsXAbbh8rb79kJ4TzUFuFvohq76ojhTGu07UZoRIvHJM/c7+50VcwiL4U7q
ATvLUzL2gSwsseuuceIKUXJv1rDIULJd5ZBkZTl7Ff4vPGB9vGR+2CZrMdrxiy361NPGJued3cr6
EQnKGRr8tZoqULfBaqlBSpdSh0HrFijWWJk729ZyKh/tgC+IAZsickfO5KKY38Qpqxukf8sc++EE
QfuO5Onl1Y/x5nyBwGZWgfJuT0ZXKXmkl5SDD0iML66i0c01cQTejUxA+ZuMjzfWmgILQ2xAsb2F
oywpg8XMS9r8dl69CjHdgCvElSINPFlE9aTLbNHBKF5VTVToeAedoxhqZy7NjDIf7EyjhUnsphmB
FI8TE0vM6vuxEYsy0Wb1BJ7mffcEfYLHhD7LGVfWH29WZLhJD25dT+Ll9VfW4wsP+RcqDEg0Ye6E
JOWyyLvJnoMgXj2EdvZydoketHYnT5Mtba8Al1suop4YR6Ivk08hutNFITZNmQ0h/xVtXg9CPd+D
mKgh3vPBFC8pwXNaqCbhIU87JmMVkm9hB3+zlovMB3OdkFIPygD/Z5J/OG9UpIsM9aZM7OIj60ad
4lYwnhbkaHAFptscN1QjRrJCFYP4hrmU6Ywy1/0VWiJLR4NjUvuI4uinAxuGwdU2m0BxQrDihfax
dGzrkmvqL9wXhG2YV5Nd25CBPHs7JUOi3ycGn5UtTnKtOzlxvkekNN8gwwCDSOaDnnpTcUEueLQK
Zol8rFL/0duP4VTWwtIq1v/rnxkhjvI1uN87Xgk3BqSUOtmZD2iNmf+W+XMDKJKHsf+QKTvAKs7u
Hg198Pnht6IgtWCebMaFvaY2L9MDRaJbTBu3hKvQzsDwkZ30Ybjy2FULurXrkDkAGpk0uS+WgQC8
jsJKneGcr2BwVwhuYg91GQD+NFzuVz7ddXp6JJfZr6vaMU1SPnNjme84REBNrkwnzT+F15HpREPs
k+kt13NA9rE+vPxOLH11UM7Fi+exXhZ+m/9twRP0DafV04SeYHI9X+aRIkU/uY0RWUtjvveSO1kK
bo+QVYx6L/OMHZFwzmuFd7Dpr84jc+lnBDBJuIJg4Fr8t81w6NyV3YzV+6Bxsw4ZKa9DG7cHt3pF
Hcw4L5jwhcvOaqRiNUPKYaIR9bJOV6JdIiBLJfWDH2f8jTs2JOvYG6oCxvcNMXvdTTA6sxgPlSL6
ly/1tvEOxlcDfYfZXm0FqZhPePdCsDH119oUK8dkMAVMLeUY1RTN28bctaM6/CILIhxK4h/MG3pL
p5eW0YesuQQldYzyDuMtE08blYFMkAt1YUP+kDD71UhOGPu2xNzZuv4m8Q1v5PFAq7gOE+W6lzpN
hfrNTmAQ9lH/G0cvZeIYT76telvkOWajEeO38kwsuNhelCYohh4bWF6aiEb8o9KKXC5olIKs/C9R
eIzPiDcmLUNvxARYJCcsWynCKjc2f4E+LQL+hXI6xk1zGTaY+fef64CEAtJAoNRxSngYEi5YWlOO
vRKe5hNfLmvheT98rkW+aSbb1fxantPu9fzFg79QtWnUK/vHS3Npt74P38pecsaRG1iwa1RB1knb
L/OFyLp4MSvsep7P4P26tuVc3X9UFfKi/e8biGndoZXgfXkJFPcHnKYut1OjGmgc770qgHN7X3aB
djXC7CdLOrMv4DjYjHEK/ntG9q5h8KW5yJuvRUo2c7pRc3tf8bgM6tW84UzfoH2h1isElM612bzJ
mONfTVfPhQ/couO8dYnrotnphOnEqdwWfZ6FtCT6GLPzyJgkwmBy+W+xEaXiL3ARRYCwGb9rocsj
ZrgFXophfsvFD7usJ/ODiD0OBfnQF2MQCra3SICjMAYOsm7vz0m5K7ROiHFxBj2BvA4RMvruk+yf
YxhBU4rLX3JRrx9DXmYT84TrnobMs1P2ihFIAMiN0Sj8qCk9+8kD0sedIyLJ+AmSshcjWCphmPw6
V8kE7DL9KesUpdS1uFlt8hokfRpWDUz77FYoUQQRYE24c3nMyGstvWwL5/nu06opZo1RWsbk+T6z
62Ug0Fc3LvnIcBjdaLPnHQpOE4Zn+4FTQ8J4eWfSEo2Sq69V9LWh7P+bEbnZPAIs6ebW6+k+IbBj
K/2lP1Q6JTmhny8NExvh7xaYjr9EXsT0Q8s0NSB1VRKh4FkM6DmHHSILxczGaUxdxlH6HRDQPl1W
HhvPpU/DmZrmZh0+edVaLnCmKQNCmfaOlCc34GUHJtMZivkOAOY/ep6sRqS2VLKMJkc6WjwSnfJa
HLzPfRR4E3btGTj6zHISGVCHrt2Pw9pJYE0e4hr/tI/io8jwYQ12uV/QZpu4R06TOqit+9slGgKt
QrzNe99Ra0wrmqbYZH8+8xKVQdDyFPqOWOqX7h7kBUTNjy72wGdlAKX/09Kye2PCFLiVMRJGZgwK
UWZ5jrpxlUP5b26Wty2xYnGLC/1/3VoFJV26sOrTWC+55kYO0qb9ANTNyWJad6HBEQ1ca94jtspG
i9rQrhqRDvEgG4PlWe2t3ZZZcAXMe8Fv1QCEb+hpiGH0DFU4hUWYvz5WmTZvaP2lPWIO4UHZU+3i
xVUCru3HEJIKtJChTILqzoG1AY5+wvfT7iLNGmAfCbSnFDZNbymB5ULG1srWANgp0VEHD8lmMS1l
DU10+s+Igo4umZiqU4zAGgCx7T6wy4GWm4y8vwSAGO053SIyCuvLD/D4CYZ5gXR/hLIUupOt4z1O
eXiWZE++yvvCx7bK8Aqt2jV840piD/NP+JsAUO15pWS9mqhmp5dg8qGwVU94c4WlVkzqiJXhbNmt
qZkeubXsQywcqrVRLilw4uzev+eRDEyNASF+Fk1Dsf8b29uZV0f9DFnFCN6O1zR7UJeg5tlApCWJ
Pt++HBrSNj/Z7E8UNJ10J2zWw0XTawmM9cZs/yNPYGp5llJj5jTmr2tGSn91K5sjPqEMozVQP0/p
kUc6XAHapFJ69a6IVGU+FJuaZ2YxXXlMKP20L1JWIQaSk/CwmmmKSr7xRdvZ0GYgQi5LDWMw8+iT
zQv43A5kqufpAfjLINCdrdyyLudoOhwQMT+sf7okbuLbl8TCF2Po1064max8bsJYW/dYZhxWYNYH
/FBxXOKTCjimePJCHI9LMJdxbyxH+B0dBagqcl2Wzsr1LWn+fEOE5ZXwHn61XkKs3tfmK5mP6gOM
ESuqF8ExKSZzz5/dzZHNtzo/fqyk4VqrTJ+QSLFXLIVbqI/W1DSqoUxotDfb0U1SxP2aLOt9CCw+
LsZAyj4wc2x7fTvduRWoslAvwPT06YC3h/y46kEwUbP5dO3AlgN7khXq3Pg+hyQkxjDGATxp7F73
CkA4hvrrx2M8qFVCpVMKLIwl+7fLLiV/z0++lIliKrkmSwOqQ9OIZPFEm6D6POoYearZOUeVGe2f
o3jAHuv5VjnjjfCdP4FXugFCaHtDuXSpQT1t6RrY7uBhpi466WYiMvZCIlZSpp1BIOt/QmYmU7dD
WfsKWDBiR8VfdkvllvLI+dhzvewA8OSszpYdVu/cMsuKUOUOw5UYmyCwDoM+YGmNIA3XX+r8LsyG
s8NUPGLpTdUaOhUEmsAC+UTvkLiZ7GzA9BE+cBkA9xSPg1NqVTO2/3ZzStkyihxyzswNE9aNFOws
hx/XIJAxyzD+ZY8jM4y5ZVT80GKYUoRfxfi6HeK1E4NIZ7JWoTt6W/7LTIKi70+CRTPLL8u4Jd3G
8HJHbl2cx8RGVlSN1MEuYOU9WRe9Fylkf2K9FhReBZTwTb3+GWkf42QMpCCkq4W5uzO9yLpuujZg
5RQ+d23CIPDsXs4eHUh29KLn4AX2bNWijimOhDKWOPOCUBAWrVoZJlol7lV4/niI8rnOOzAn+WPI
bM8qaREWuU2BIW2dhveTWQh4AJZ5m/SxUUGC31EKxUuwhVHC5exY/cnL60lnTZjDJarFum3FV+kN
wSFzZVlKSyLiQUsw/b0JO9WZJJ5LWBAl+DvWGbFBcUVMh1VJgqXwaEkKM0Hu3HXb9twTV9yYP8Mw
l+bH9MHuegl9J94+kA5MGpon6KqgpElJGvaz0FTKd3aIqBMwR/MBvlhrFM+ZD8gPSoXspVKlqmLC
pGBWB5bA83zt1xAcu+sOwpMlhoS5Hi6XCav1yOMqdw9hSv4lrCiG7Aoz6GAju8CREsp6FhqS7Xxu
T84KB/RpMpC+VqsYozL/ZhL0pPiIqH0ff720wdR7NN6j4jR1Pom6hUuocqwJo0hs5Sn9WDKXIPxs
1VZrIgIZFn5haEdxGVoPX4JkezWDhkuZYV3VsxzABUok86ecZo5sSt9kijakGjNx25riE/0/mgY9
gQZwlk6UqF1p0iexcmlPzJ8VR365xUGOxpTfRtCP1KI1gAKpjp87aNAedDgl6gcoJ2PzP1V/DnHB
q/vnXt9ZH9d6P6sdreCMAP4GQ5sBR99BP2x3QvrVaHzD7lXsLtrb/U+oo1JB0aj9d86GxIbbgPcB
bArfUBib1TZyyaMhi2r3+xzXri/A+oZfZ2LB4PXrNV3VShaseYbJ1uCEQ32kerNxlVyGq5iYwcR2
Kle/2Hp8e+6eLXNzDghDRUD3fSNPmYf3uAwU6JlB3ZH/TXps9QPRduYiR3um2VHXPUGZ9KeoA2Am
X15xj26MQddUjIcMRAXjRqQ/rM2rPaKx7wQkxmwhopIrwChCkVVag0qQg79UBMKCLCb9mTPk6rWC
Axl9WCEKqpPmBayd216PyUuvZbzPh5qs3wtsP/TJpqKSoWWAnd/gagtgLVkBXm7sQonHv8sV7G59
+eFwHDf+ZimV4UFlHLKG2JmuMMovlelCpmoXZj5O6IWi2cLhu6wW0PhVyUK9cWntascTwWXnAsUY
oysza14fhs3Ee+DjAAqsXnBla9ZR0zfKF4aunUyAcRcgkltgAuSsO1tirQjx+qiQyuwOaRuPteFN
+UXDpUbreNfTvi+4uMc+n02fu8249IPgirsaqszAskZcGKMiWkfxILzpj5uRUsdA5viu09akNc/i
Bj6U1O6P17IcEiLIVoQGg9CPoIGXh0ePEmkWMM992Sw44OSo/v41qrxity9dL7N2gpHzU53P4oA9
7NgiPRt9XZMefAuK4fxfdKZsFFrOK640t4q4enTVh1VgpSmJ5j8G8rqNeALd1TUyQ9Dw7gWZ7CrR
lMDjMWgdtLYyrRs577qPSbBrWI3m+7Zjvy7NgZ/S3oA5bQss7MLs79FB3XARXw2/cko4agZTIUba
U6KSvfStxu41bIo9UManmNgN4jo4XauoktjDpGwr0u3OsvusIGHEyHF5tbynrjn4LdR6nMyuhN7i
w0fKTwuxNMmbziqZKLJdVB0o5ISIhf/EZDPTT/mRck8RTtOPN0qoYR3qIpuQuxyXQpANz2Ntp9gt
cYBuQv4MUqb20nlMMQe4/JIDctHLBalX4WX1nBVXT8ofsAxe+V0z1/olZZRMxQB7w21DyuJs0CGd
BN/gr5N/fEQGQeWErf7WFuelIl5F+YhJb4Ni0TWD0PCdFxWO/EvBj9MRT6aLVazUQjPbSDFlTkPI
ViCaeRyvF9N2BJ/7Ng7Z8dB+Yvt8TTBoRIhgMGb+qxs/o1MN0FqrC9KMghnD1LsX+Ae+P7aZzKu2
ZgOOVPMSFMTehrOZxZUaC6oI3QHF8Fek9JrKMoEMxOVQpbarr1ba92eooyqhpTuthbGdX7xP4fnC
03IZk0EDYNltVKgpr8oec+qBbFBzvZzwsuroktBBsJ16k69mraNwQPm0daEErncH6VjPHm1sWsGB
JdrCYhzX7luaRWh+E502jVQUyhvznJJ3qXtxquW+jrs904Xt3jZNMD5n3xEaXM55XvYqw1LHfCBy
l83a1Sdf/uumtoQKt7aiXTfJWXVLXQWG70kD/iuCsSuHfEF0RDT4dM74JR2qCtewbbKhoCJB3S5+
Z2QvmFOdtqMrjTpvMtfcMtRZnaKQqlE3mgW6clklTSQlxFMpp5eDtU9/KHFZoRmBKd+UTgWfuQbc
Sve5Zmg5cOS9TbEeIz1+0hj0WvGCqpdML3Nn+WbGqjIkdtqeMdvDqf0EEy5d5IKwPD/IOeSFg56E
28SxpMSifH0JcCs6ZcRkBCEms3IJ2fOhTnLGpE5pbnWO5Lz+hLdHpBewG3a1Hr089jW/ba6amWVc
F9ZgqqlZfLBBvAEpVJWbVsOcOFAzqknFquD6GWUjGWYjWGAvSfWDLYAr1jSw7GTxL7ETXxEBR38A
dhompP2yMHKTvNJWacL/VO1OG0Z6hZIj06guZODEVkHq13BqGYbhGRP1X9Uc6C9I2Adm6an/z4/B
sTRVFIBPJ3PIOCG2GqlhOEgh/5UshkzkxJgB4Bd2mSjAtmK1Kt8QC62CE9GRTqMNTkAjkGbIQORC
tagZSNfl3jd7pKX1+aoFKz7QZQFRwM2YY7DAT3pOahy/PKsNBcj2qDsaqbr5i58TkPxF5btf4D1U
9yxfvjVGswHVYfKrDMobKwViRH+ZCBTAy0f3rpmwtwQTa/5QvMGH0NWPRp3ImScgXSZykNG50CXg
DlUQs1q4wM2F8fSkAPHeZ3YHz5IRByzOdZSfYrumg9EvKlKVFoOZyqOhLjKkkghJOzVmeuWcp/pu
0KgYH6vMKl2CE/i5xGS1E51thuCunv46LCPcdOibELf0wrHz4rSKL8A/4PpHiP4mxEzgZNZLnPf0
wvHyqB2X0DoGBP0C8d9W/IUy11q8+fzQpbcLp0XllRrKwAK+4lZLAXl2tCbJgoHrfm3odsYcNbpb
tO0asuWCPigDzdquNbyfL+nM1g3HhbdIbWP0fnCma9ftQWqTQpSYZc9Ah0mfbXOdA0i+0hm8R5k6
uMG919JvsbtoiwYWHKzRxzptiRw+5IRc25SqPOMIZEOFiV4bzjV5yHQnlkDK1JXzs9UhFrfdO7SH
6FLgV5eyZBSU8CdXFVb1GYkeSNPLjQqm6TMgdQk0DvPKEldcX6P3wSv6ruiVerkbJMqmIa2bOnQD
LpeWPJDIZ4rfv6fUa705tjtUqcNekVYe3tPpbboCbfGO0mmSq9MCO66nQaKUszFS1tblohRCXnhK
5jJW9c/4mlraLrXqEALQk5IPAPUxrpIqe1IrLNixRa4+suqlL41ntbjP+e81JnE+zJHyMlBXFY/D
shIolZ8rb5w6Zg2mFuL5rrdF3jHQlRxFBWWYkHQV1IK7xmJXU+DxVXgUdi7/xbHwYM+GQxF//rfJ
ev8hZCOfGiLbecu7kHT9jYdaTidv9Hgh+z+HXF+XQj/GK5sSYpVDYQT/Rc+4tTcEmDA6Ovcbxj++
veubFB78FX74ZN3kepSWEEmIBGaXbX8JoLk4A1C9OpexHMMdqbARvBt7ikySMk7zuuEVvzHQONu+
oXCqwpX4LqjUDsRAEsPMGcZVSbu7W55Lyx1hGLDWWbUinNOgpwYog4gVQhsTsKICOrLotxhsubxB
9wqmuKkj1rfEd8mxDYy5kXXRE0VKBbufC/vQLUxwtqQzvMvba8RNdjXFJhjJfKKUYpyJHecIC7z8
p1tUKjUH/SXvXP07Fq47RPrqAHi9gAguAvzdwnNZ1Sz0kF8dGYaz36Fo5S4rfYmm7WvjT47G9cTS
5ZDCz8G991lq2wLllSze4QEylRTV+utbYq/ktSV5PSGWnx66zMvlhXlTZt8NTtEZHTYTZUt1czsZ
2B8O9SWNzMIdImHAfo2rAriId6dcAB6GyEA9dDwSwIZknnw+IL5/+dJmRmHNBPNt0tvcG6R271ys
hXfLNY9n6UGv8V5kN5CqbsLryMStFrDQENUAkmH09eDhGVtQVrH9ax2Ose0UuHFBlKPuEz9/BC6O
sZ+OCGL/jMomFqzLd7pNVM09gPQLRSnGByJQoWLU/DY9FQGLOihY1AJnaZP2cQtAc72Tzxm4RgK4
HP72HArfmgnxRcckLduNO8oFguE4Z1yFtQIcQ32xhNuWKe9nT4TlSVDBrp1IPLe62cHeLG2njInu
Ra3DcTH15icUbdMyA/0DTucnEsQGmn3uXPXO687sAz9yRxD+JMo+MakpgI0vIJh8LNk9L284T9Jy
3OLg7lvEhSG7f1JweDd7A4jNpjPEgRC/s7dOe5YADVRTwmLvwdlUoD/29eYL68PuG+Z++RHLCHTp
wM7SHgx3dufmfxKYDXDCNEUu/YJ91sSmqyDsmOJEtFHtZKu96nMRtMVaUzAFd99HRQrK8GYEbVK1
2p/V9OCl8j4/HCphjExhbBwoEIYeKIbkwPue2sNUBJzc1eM5gyQyyP03nVJYgZLi7yE5TitpZqVQ
2OrxVYEjZWkR7T07VyXbGwzJwfJf24fzHpj1EVgoHxo2Mg0ctaL4Skxr7DCDV8hjhHROJRfPPMC4
3UKKfmAhIhmM/9Ad5sTI2qznVv0/KsSEV3kRAhAj3j3WNNabqBj3DAiMXUr83cFNJJLXf89jpAnP
Kr4nO3LAdwD7N/dxerLrGAHqFKCkmsw1M1A+Awlw/GrRtaF2rdQNymFFiSmnYDztqA+BWWcHonKT
nuMBQRkrJ7d8+65BTC1Yos3Ih76/vHVHCKqaNhYmOgpFzjPxc70rrCecegRnO2+DBhFu9F1vGQwv
fOHdd0WxYOoDxHa/hif0F5RPSUnsel3ANikjBZZkV0cjWW2VStULEMSQXXuhfA+aBAxHMrC7lE5Y
I5sFM49i3YkyoIIpojksbxel3KO4nwZgl3P7XVhUtazTiRNLL9fBoiUpNK8GxW/xS2r6OC9wLhTm
8+0UoVXMRs7DLSkFfd7rzf5VdAUOf3SE1QjokFFJI3de9OXpTyk8JDzAg6/LxGV8vesqy11AWU7p
3Tdjoh4c8kVuUsAXoaqYVvLAeEuniMN6pnNxLrDI4CgHIzJj6yYLh1R+QDC6wtU8q2j7QTgy4MJ9
jpQdxpspJJ21/QAAhuxRh9v6gfvfxI/e7IARQxe3r3yLnmEEpZwUD2TvgbfSW3FODaHt8XHI+Ry+
L8udFcy0MbcZg/9+vMMZbzTGL8FMbIkhgs+8j6D06ZsfsE4cHzRRCYR45FhmEL5MtfoNFP+m7jQQ
0Ii4btvC1Z+YyxNKYzHvBhWJww+PoeEizMWUwMgGZ0bVZvDemiGQO1yQvn8znWTn50Qw3AwyYQwd
0o+dl74OMB9ekNcB9idTXom/Lp4PNdVrefw+p387cuuTgtOKyTSjuoEpffNahsHbn0u6qbSqIsyW
o6BnvjIAAaAAdKqe8AETo39WCaVMWmhoYmFHBkcaH81suA9K2H7pLtw0cUtcU5xnruMBC0be1XPs
crUhdzST9osDrJtxdagtHvZqiA4JHt9PNh3V4kwKkqqUL5QSodFXyCb3lQ6M613XwetxkksnqVV0
NocpGdLrxUITQkFvSDsYMQosRfVe09+Xr/cBQ8LhiPHfu9yn5rzV7Tc0fAswYmeXcgSbSgzz6QAF
OrWtiNP8bANyKbjuOJi+lcHalBsFLzaeX8YmCXLAM0lj2T8Kg5MO2cTPxqBqWU5iRqHA90rVS5zC
AIlNElS6UB5TzUWBnI11+nwR570OosQyGKLPFxnCd/qeAy8PnRZps7h87EZcUrV6ZbmotdndjcOu
+fU5kk20FiRqOZ2KV4mc1oyvrkK59z+loUrvFxJ8NIkiTABZ2Bw1rjqiaa3WFoqkJ4Jt4mSb9gE4
uUHKdVh32xsHm9hUetm2QQW6z4in9b0TnuCMWMYhtcuhWCZInrkCcUMPIg5ajo+UA/FB0XVBKh1A
uZQIljJR2W/vwVIqX/avWJygn/6NjUade1IaZeHOlsCwWoAWFQpVAGx3cU1cGpIB0KDYJq0+3JBE
prCwU1wQBsk6RVtKtz0eMJUpqJvZJohX+sQ3vPWm3NvkXDN9UvVBSrI5jzkmKs7M6Ewh0ulGTTml
OdcebvTOuOkTJtRHcSghNwirbDneZz5LvjiYFBf+VnpwgWwkUWVj0MR1dX7ze5UjDppSJ+bonr5Y
JX/ecHW2HPMYLkqVnjAxVM2a6Ip1FPQ3FewP2yGxcJnZgyK2/RNy0Kce/1GlZdCGlh/dw9QX7s9O
Waq8BbXpNQk6zZErIE4XfEgkBewkqLUg/Z9PqYCL1mlYMCs/Oa/xq7fsEgaGukfwJUUJYEFWQB01
gWBC51nyUCir/u2DMKVtj9jL0I71F4wpEt8kyqQpIJtdnfRJ0mQebp8Tv0ibqz0a+V+IAt/N4fmv
7I8Vjp/ITdtQz+jKg9M2dO0v+/BQzGeqoURr9JpwbVdDHZ6CKZ79b8zkNiMkAUIPvtG9vuDGLqHT
aYdGeg9qYbig4Hj1cZu7CD7q2tBHOwo70/YJAuJra7Ppmk2a1mU6W44DOn6Z/fh5TFujG4n6x2vl
nmemBfvnihn0OSNsWH0aoMzUv48g16pfadKfih7uNOuz5nB9KOSmLy1dKPY6dJjfvtfzpVlEu829
8hKSW0ck/O+8fA/K59rjZifc8RQtbIfWGBzuz0+a60/v0gbTwVu2+66jceI5WbSqkI+h0YeO1kDR
4LsvA0jZhLRYiZOgHNxR5w/lgufloCJhPoU3KCwKCaor4iwTUrjKzh/cEMicifpYElR8b9Sb1SUw
OSoGA6FrGWm0xci3RVuBC0T6qgvXHCNv/58Kdg2NjtIWBKv5MbcTGM/h1zYz+4r90LMDs8X7WnwU
9uC2NOwGX233ONO4q+3zoo7N6VN9zVTiJ2mBgv7G/o/AlXI1zNTIeCWud1e3TnefczrtdRMvQMAt
rMnYE7qjFQyeiiWe4VM1zLEe6YuKAt3sCOCkcuAZH0gTIM1Idbn9Jyf66Ff98NzaSZal+W8F/uxt
3uLozF9Y58OQ9cvlXzQnljj4X/qDxjbtlP0lv09D7IHI9/S1BaIdIJvi31VB6XWMobzHPwNkY3cJ
AMnCWwK28y02pWM4jCVznqYmI0oI6SsU8a+ON8+XGXDp8LJ1Ub2ruk8KC+XYgXe579mBuwmtyoOu
I9t1NVODRpzSxnVOogeVwWk3UmRsx2QyUddT7FNWTCwET09+xvqL5a1miVqVQqNi2ZnwSWgkBg4D
ibDb0m042OKQGHKv2ZLeMwMVWfXpbAkmzoKYtRYP3e0uQY1Sn9CHJtxndhHlk3L9Gbz/wjVXMbQl
/Rf1qqVZ8lrE3gAo8//tvG+ZaMS/12LLAzNtZQBOOZPk11tRPzTFAR5DYhO8p55KXkLpic8S+Wa2
dgjq90wtFLYK/s+rIVzupVpl/IjQD2kqCsF+4Rxh82PR9/OdfMuSUPhx5t3Tce4ZkSm3tX6eUk2i
7o3JkdDdxVIYQZnSgnU5peV423SWGQ5KFasUJ7TcOMCT0GYhm7w+eHEPSQc+LkyHEv8lT/gQ+4VB
Hk+ToriXT/k4+H5iZ0YPnY/m+rJi7vKv8sB3z5h+aNq1MnEJJWQFnYTAykqfqZgnxC8jNQEqs7rO
rLooh58Vamswb3qD/7wwzdK1j53xp+KJ6r1s31kI/5ZCAAy1Oaw/zQPA0XUVKw/vvQsxKcWFG7vz
YSHkj4i9i89SkfsqkPxuwYpkvdJVZdPYqvdtQ/iTw8puVFmqu4lOyrAtdhXlKBG7sCr5mh/PI2hs
GxQiIMnehx3xWoO3387aD1mlxsMyiL7QJMYovK7qZjhhRFdSZFRlX+MAlAetRKrmBqxK6dvff+DZ
VBUIK0mllxQcIvl/OWz07B4rVCALVepDzp7SZSIAajV9sPS1EfzpVeFLVgi7jDfDZOha1YEZwyYQ
WXVxeKaHwLuHBQ9sFKjBTnpe1IsNx+YVpGmikb9ZLZFcf+66r/rSublc2tqvBaaktqgIDxZxEugL
YukxDRiWtWU3HQ093e0g8K/Qs7Z862Mm32hfHGyjXoQiL0AeVrUAiDKI9Ne7XFAwKYZCh9NghWOK
53SvRyQMwwd+nUH1ao3RgHI4eST0rBOcAYpuaz3ot+lGorIbxT/N7R5MpWdxW45w2ei9nMHfpO5l
VJShF+WNLuLzS40RIPjYCNozmpoeTm9/cJxGpnKNgZTyyJ0llLdqUYr0hCoBewIz8J18L8LfRerD
kra9lMe6eNVKYQFRCw6FbtBn2rX+9PnsKtWkMvv7bQST38SrMmMcIkz8jL1MA3W9dh+MgfxtLVN/
FWOi5SBSxz4ipwhWU4CI+MQ102GddtMbuDYOCnq7BinUesG+pvSyL5atLSVevqCFj80eZudElKro
S/OkWVuAgrwjAcZn3gHAapGC191ja9F9eCDBnl+AyOi344mFJzuw65a4flzxZ9vzz1s226mGGDYa
qDFvDyNFK1QsnJyR9TYibi3UPL6+fnUd6iplSIJblehSJjf6llNIUiBIsON8r4qVocthotNoa3lo
b+n14qMDaHVwHU7pGNbRK2OWwnNXxorNaYpd3Ts2WhHMe6nMaNOvEyQLJxHUOr25/xWhn3byZA6d
f+65maJNvwuq+VI1pVHR/IszxTqGQRWi1gCwTNo2xFFloqdMAn2yUoX/fsHG0a8rooqaV8cNzRce
nBf6IAvCLP4EGUEaG7vvhBTo0OiFMmV5sqAM37awy8AQgJ2iMPUm2vNdVnZIlkuS6z1+UI/xOHJI
V8+eISJ7h1/ttg0GVkM98tPdKKJkSR7Wru37sTM8e2Wvp08tK8PMA8RArd2ytwMnSkB+5oMJxgKu
AUSH17hFo4zpo1zJ17axI9lf2lPBhRHPuiiQINxxJE1WflLD7BEEwDqL6lvQUHn/hWsJ0XV9qdEP
yk3/6NEeviSS7OKokxJKpXkHzRrzlB11Vff4+nMQLo+0zdnkxx42JuUMXVf+mO6ntJdONNzgSGZU
UDlgLc3Vt5Lk2JL69Khtm+hYsYzVeoZESwe6epV9hkx/RlhP0Xc/Q+/1v8a/6I4B5H3rIGhedcso
SLypKB0ZubD+wUxGy0NRNmmqJJkQAs0jCjemQOT9BEO3JbvkmnZ7r+uKEptH1qNAcJBsfNSfMgC+
ANaZFX+4OuMSPx3+28LcsjzHk9QnQQ+nrG440QA1KjaJY8IB9ip8nvnaV5rQtCN7sOShiRw/dfOF
jEyu+nVnJHLDfAi/9Rp7EvZspzot3FLn3n/QKpSTLD8emB3pg6/fILSi88Ju+WTwhoGzYiZNYrBE
2TUcQDqcNymIlci3nz71nfVboS3DxIz2G4cLPeVKuE8baRep3OhB8vVIMgeon5QZsV3Z/gHrN6Qg
K0vc6crLx3561PkIDg+s3ewZGx+qzmKikzL3g80MDar7oee+dxFILfugsLOZHapppK1TbA5zc+2j
gyOHXIf60sLVfu4mV69Q5f0yr6awXSCaQ8v9xuiO8A4TN8s41Runi9SavqoSD7GvUe/hTRY9aljz
Wjr+Zim11EtKRES7jc6f8P7HXtXLbPCdLyihYGjQA9CTXJgeTYpbAb+2QTKIwgYPPieQpqGf+xdL
0vGIxZbIGu+NryWuELZbs43ROLRHCFUPuf3cZFwlKr+9RJ/a3HxnB+C9cD7E8Xn9qNtoT0t/NQBS
AY0HV1646ZVbcBVJ6UNbRk1/wy9tlM1yyOfnTa+qg57DQtkwBBramfjBpbH7Q8eAS2IHhrkEUJnP
yZuBrYpzBxnIz8KmXDfLoXiKjz4uCZOx5qecm0EtHDhIlFN/OD5u96y6lZUYo669JW/OuMmFyEsq
o0oDmj3tiNLWYKLwikg/SSpRz0eo9sPS78Ipb22uix2jIeCjXyS3xSfeXwHhALdIyj6AISWboWtR
7fwYXscZLhkIueSqIxe5ws1TmfKZiYc0cgpPV40cOVU8Iq9NqfxIPas/AVZT+fDCdup5fU64oBs+
m4UMSWHjlfIaAHWrvZlPG90EjaVOouH+xz94qKqTgEqB+vv62r4aFdULtm4ZgQIRRKWi4X4qSf8g
cJb7nVLfJGn3FMsjCsZhgl8AC7yOPi2NXun1kac4XNtjnp3a8RbKN8Hv/MvN9/B2zGDSFo22cJ/G
gHuhc4OsSTsjMAuJzUx19B3ubQo2/UCBC9s1YAqXkNNvMM8I1KVPH3/EY3gQEhPk0MLqa62YvrTU
BgbUPjpA9iocY3QaRA5GuJ4ZKCZ8FS/JYsYJjjes2E2IjPlEabBgXDQvKdALkdu7bu6JwRxRDeDP
O5VL0ALEeiUNuqT8G7ZcVEZ/qt2g3uMaWI+mWZUE59BDWEY6F9DJsaYzAkihsctOuWkr3CTrnedI
pwIdKHivGWXizeQo8kweWczGtTsfNvgn4ZeoDgl6jmXsmo3b3lHegcvr4vKGF1cSAEPvbXhLqNld
zWkqbNA3gXBOXcXNHin5EESOu9WwHUDFTPhDLE2Ze12Ir5QLY+1yNOTeAKXt2xbgFPilgHgPb1V7
16Q/S4n6f+A/rLQDnu8xurGH68MmjB9gbGvU9H8WowzgvLa/+5GfYFTcC9q8ax9iDipfdso7TDbs
QGdMYA3yOWU/x1ndJJdX45ZzByD274E/ZOKUeuGPGd+BAkA/DPBovKxdq8DdxaQr9fiio3Fb+qcw
6kb+SbwY05RLhwYWxWpEFeczAURmXQHFfu+HB3dg3Onj+kLZLwEWQQI9aNv7iMdOxxA553uHdENX
npGzK4489265/6E7/vzdY4P5vyr6C5E2uPaQ0XLiWXgC0+Ur4Pk9z7m6cVx0xsMOL8tMVO9uEMli
OapyeZlBtEgM+wv7Mx4SoE5WCa7cSz569OwTTogO8kydXJLi6U1HBBFWRx1oYj2xHCs3sOE/dy5U
vFh3oLAP41ksHQmq1artj982GT06LpeNCtlBnaWtC/neJmlS5fhWc+qJ2wkp2yVHm3bm9Bz63ldW
+mz7LlQ3A9WBF9hG9QStfZihBaLnopXXPkXxnTlMgzdegAnGidzUIyraURN2EWYnS9JttkCKMLsE
N1jr+MdNojg3QlrxeUBkFnW8C6jazUY8HR6b2HbfwUR9x3536kJs7aKJtM28e3tjjT7VcLD9jzkC
r40LYzP6+pOGJNp2neUilgfbIOsrwutSJ9cmzLPun5hGf53Z4fRF3bPhoqupMVNKExtZyDHDmEZZ
LuoiXLERmysA8Jml7kuTQadVsR92zcvGzazeqj6ejPViVcCKFGGgM464QdOEoH7HheZn2b7hpbEa
BvOOGMVyb+W1JAX/M+e6z29ThvRZEJwf5F/94hvBr5CBJE0cBkJo+4R8zYkutBHCkwKG01lVwNIE
tIE6ROLqZxbDA6qnsI+FOXlDgSyOrXer5597ifA6oQm0P7Teo1Kk7XkkM7bTLFIqAxn+KQgCyl4W
1SINCIsu0dFpBuDxe6aelBPjZFb/F2ksdp6gFwYB5eRs/Pfur/kDcQ50zBOJ8PUGO5GPkZ6745pf
biKjLa6qm5NWAFb2l1GdqeuLnX/hBt2Jj+zNOxXKHrCH2U5E+COD++pwcm0jFP8lgntZeGMk2ZGc
ghR+H0po91qZx1U0P5PYOWYH0yW14RX9Uawhasakh/Jr75YxAxcYRReeRQIdgNqsMD9YHYGGcQkk
rdUjSpaEildhEBW+LUXMjGJbCBeJ3vx1pqCsJG5vJ90+WchSAqmzvltlpvaR8PEQqJjmuL7c9qYX
FN7eElu0/E5tVkuRzVvWM3jWyOUHotVQHMtURY/7PGJo8eqGKXyt8wqEzWtgH+7SG6vQE2axLyjG
UNXhozH4lwqbDWEtJOE5BeCbw4cYRQ0dxnPDjCGkGl3I2Xn+tvrfyHzopAt6yAC48O9DKqEKd35G
7v1A3Kmi4sKN+WHFIpFYfMbVFB1/SeHlPWAGctntsZCRSpA8bng611sOtRnhE4Lg6ACWVVTRPLrf
SpyvoGrwEtKuD3FviUFBwyyzh/3fp80MEhUbcyoEOpBO8hc6SkCmWKRxE0GpMWkXkC6JJpXY/Hft
43jAPs6Hb8fj2qUA0QsRno02QOGkL1E/CPljcTj/RZXKJ0LF4xaO4Lq3xJjGIpJNjHerceggY/8X
3C4SEKyFovXmqNO2acXrFCaoTnCHBBW7vf1VskRcyyAAcc9XxkUMRvkZ/mzV+yFY1eIJE8AVAu08
N6KldkLKYjB6q4NXzKHeWS65ayEt6GglbDs5l9lKuD+9pvjqbqeLHQTzOTBvF7jw69ByD5ehinC7
oh6OFN/0iBUJonn2zZGhcCDMQzNbKCm+dW11jrwpaQv3rR0Rz2CsgZ7596AF7SMdExTjCFWFu1e+
BjUtGPj4I0C5N1rRH9d/NCsJJ/AK3fEiVdsSFleXDZBKNjmkP4/n9klJL+XKbYdjeduD0MG5J6BH
tOPdNU9MtWGdjY3uX6r4sGpfxnZ4lVAHQjWMgXJaRpGdgYYxLlz6lfQopMZdzMUmDXu4Fby8+WOB
SQ8G6do6YhsI6h7ilrHWmYLnW1hLWU+UZY95v81HS3q8pNSm93V35tv+aRcHS3zb57GjbOw/5pjH
am1dIpSBLc9rP4n5dtUMCcpLPv1pQbPqE5yvCHCy/QyBBUiCq/g3VqZPOC0KGcbsUXcJBxm2lf22
NByx3RkueMg09r9frdfk1+x6xd0faYHHM8ty0037Z5BiVFLjHIVQ3PvCuUKO4oTrnhzRGSdb+OBK
OfkHQfQrn/0Nh9eFEUOVGBSgQ7j8vqkhpjowSxLpKKsHzZAfY3Mqj+t7eymKR2Hv05kPr9Z/1sIp
ytiwr+VCEgLB+yVaLHykXogf8V9dzrI2O89+33hzOwGn6vDR+aN4IRFhlaSVM6eQbdmocuTTBbJp
Iqib3lKqETCMWWmVylmJnAlEhTVGW22+J/nZM43ecINlZ+xcMrFwD7JH3EXYEhQC2Nn/umI5OAQW
f66HpZvrKyTpCrx20+AxjhGQe9Rnd9ZZMOGBFbsFIXrjsEKaKtRmyif2iJOEzO4xy+ISwrd6NRXi
dIFzH9S7+SLoAbKahqpPVLmF+kmJG/4MRlAvDep4d+12ukdbqt2dGMgQv+Jd+V3H3AfEqgaVdswc
fZ/t/u175E+WVg1divxMntqJFBekQl+Bz8IA6i79+93nTXN+MnS1wbKcSCKk9O6igIMQOTwFSf3L
83bSAxW/CA9XgyMdmWIH25zWWS9kAk/0V/+KMuVTxP+7gmqa1u6Un7acyfQBde87ZfO9CMyqRXMd
jHBkqnYlHmAFaBXYdly8aGwAg8sbjmctSCQDcwwsWfEVwyH8AQmghF1rexrlOa6WoyygWgmNTENs
UwkzowNAzdmAzRqEKgTmbQLlPh+4f/2L8IDcMZHU8TrH9bJ7M0YgwarW4LZahNHz+tkXAHphSYxQ
lLtnHQgbTh6zLrjVPJ5DYl6UREtF+FzZWo+Pi7j/Ked6VRHj200GjV8Vy96LJLvXPPuedrCRMJ0P
cB1dt2Ou2Rdx33UBgkX0PSIOkEspUlK/FwUgsYqTJ22NG4xSPlJCee0zdkp3R9WiXjUXtCMSX0Td
EOm7N4FwaQi3d8EnKP3gd6dxJEApbP3kwG+UiSH8lBDgIxu4R4ua9TTs4YPRr0Pe596vQ6gP6fF/
KOwEyem2dbPLy0a7La54oZg3F6vyLFtCTVSPZeBNW3vyJ3fUwYMm/zzm1TUjeXtsrK93H3W3WQSB
8DHcmhPJdOuOC0wxt0HqMuOFJS3X3pL/FBtEeiGuAKbKoZnuqygPNGMaMtKQDz8O8yrhtByFM4lU
kTN8mvald34j/ZxbdOq8hpAV9er4k5CKQceuToG6PhqkEOmVHQe/3N2YH2GdJx3MJUbRCb/VAGxo
LPh7XczDb0haW8KkIlGymHodV1PZlEGUSrqZm3wYMKQjqkOdyXdhCumc7R3EHh4E6zHA+kXEAqit
R7nCysqK/UfvReedHLAti7LgjiJm5N43WIkMWlyALMKRRkjlnw5k8Sxp+vkDKhrJTB/JgEukYaWR
4vWv+5V9Id5amhyEot9sHQIEYpKCDbgOEd/o0Dd/Qc4yMWUmBr6aUup1SqEWqq1jGgkHYXRh46Hs
prvFUtsmWp3VkI2qYxt37xb3nM+bvL95mSenq6n4m3WQ1SV4MrtUfikVpIbO5TkPB/h1owey49tg
Aeb68FL/2AnOTUTn5IViJ2Uy3sd9mFx1QDQ0R1yPR6WZqvVlHkiej8gcc44dDUAzQty8l97gjG1m
+uT9vZ4r5KZytEPxkd/hkIgasP50KHOHz9lgZFvlo+mdQm4Q3Ib2Ljx48Z2I6Jqn+XxcNYJBg9Bo
R9k8M48BES164gl+zcBJ1K5pMvrixeP0IuHBDyh5LmsWngOR0sKFNG9lmNkT7buJErMBQfBeyZcJ
PKmt1J52iMnsQSjXTxcPm4ui9+ivgin7X1lnjLa2vMEu4JFLfnsqmCbqKxlFg2WEyZtWOGoUZeue
PoN5yuu241VBMoeq/wfMOhfW72M/JEU8122xEGdOfRwtTPMYSz0A10fEDkL1fmBvKtXfbIXJPOvv
kKISISQ7TIqgRKK0rEU5ARIp36KsF2pVqEODf+1S/xsjNaLxC5EMHjeGFr1slafyROPeh9YqU3Nj
Eij417ac6FaniQexBmlm+q7TmPiP2rRomSCrPNmNfy6NAnW69JY9ypRj4J9bq5CwUQ3+/e8/pac7
urKXsK6HtxR1Jt9XYM+F6AM/4369+Kv2cxiqPeAExQN2ptf08QQuAUFJMXVDwdgFSJ69+dgutTCS
cOXE7AtzBb9BQD9xKLay5oamDVoP2vrrETgVggKIn+JdnYCE2b68vJGv7jmP4YNwoSMypyFiDKd2
K7AWZ2SEXjksRXAHX7YbuYM56Wxyl53eKbfwrLXY5swgzOOiMuC5yvRtx0sBsScjBuQa6wsZSg/O
Cske6dLzEVjIe4aPqpGD+y8rOS7AsBAfDaqfPMRf6twr/wL97TmwY7U9wIbHFI88zPf/DJuL7ITE
O828UzkRWZjKrlcotkcYOYxkKRAlixN/S8NIOx0xepPMKlaVwtBQKaL4eeSNCZewBvAok7W9GgJ8
wU6ey0UdUMBcr3sb9QwU+zwT+SknY+4oxJpHF31Kh0QlTCm5xRNY7wPNx1imrOtk/yo1e5Y4YcZA
1dvHV6dDKBPk6ceaxUYPnO1aNqYhDEGf1MHhQCdwJEL+EKLgRRoWQ1Jb5kPPgYPScIbOUwmtZ3qP
BqG9q9xnJ+HGq5L5LT7ymWuhaOXrPpB8QAg/XuKGci2qKf8bJTgcPBgfC/kfAAWWvGu4pj57jEeP
ZrUBhZfxwVy6m0/BPx1MIultNRPW9lJaUcPYkgVCsqBBJtFehDgvYcXX9Mo3O27cVUNr/NlsLSTv
fwUVZpflK3/dnj3nerznyf4h90XLVz7rrHgHvlIHj9Ihr46bwSs4KPoxDN7W/3+n0grJFGtNE8XQ
VPuMz2jbxbPvOA+TWCFAX3d1b+3Rgm4SiFDsXnHGJaBPcTdskYddqO7iq6+YlWAN2JfMyMWzeU+O
AfAnty5F9mXVqTgSmfp4HlQJgPtKKstrH9IbMAF79VEID8p01mOVVzFKrHt7rB+GRhue9VHDPj9s
xZihNWuuF6Fs1W0hsHUbSvdPgYRib8kyhxwOuzWaWNBzXbAQAdFVKxd3MeSZfTdN54c1QBwegbkd
oEEfeagann0RU5bCQDcY7m7g4T3ja0OY/3lSKEKRElVgL8WrkKsaAkf/U5RjbAYb0eFvxCWmEmb3
7AeweEi+kEI/C2zkpZvoH9xbaRUJX971R1m+Sg3iQkxEVavcytrOmhqEKzuwhILHwOT8c3iHWy/x
RjTUNCPz0XULX+1W31L7yxcAu9XINmxUxxnyYQLofcBKEsXx7joA3vz/mdC0yeQH0g23IpVxd5/S
ok1JjEn0Z/PNFomtsCTG5evSAhli8TmavHgFGbe5M9solLhGqqh23po+ScwAwP4oXn2EOtJ/mxOu
+73WgRvsPn4rw5gz8vyNwJpheDH75Aux7/qpTLcwQMaOx9EJaVuNhYvtugsoLey1/yqQSjJBRXNg
ycf+jxTQxt8YoLkJHc3QNtX6wmlxdy5ejouQzXfKS9wcYFhhrAgUFuYlNrWqXQRcdcvc6iQFN/Ba
FQc/Ig/UpE6Vy+/0rzabFe0etE91+f4/dBMFJ8IxKP99AkaZIAA96zQ1TLK2nKyZvfJeED+KQhm9
OQG5951LBqtp+QyxZenHmKOo5XeWdWUtzXQF8flDwQAtp7dCKH38DBdlQPdyL5v6pfQhue8MKm4x
4Br1N7wmEpYe67B7jAWce2MxulJjkxEffqojjewHr1j2q5potukRn0PAmjHgzTzMPMBITbYfseay
HT3+whfOSjGTtGU7GahGM09YBGMk7M0RuR9lfGl3FvLLtt9CrjnZrVu5vb6RTUPZnkomxLi1cqw5
NG6IrSl0IorfGAMyct67wDU9oxvAidi2a096eP6Q0WZOHg4071bWICifr1HOQfKb7IV5Z+nAfO9p
c8305NlNh4KjCr/LGqiK5j79ZqGtglznbqPuCRWLY0JJHLiA8hG2cs2TpxyWOaDsoyQL6/BkHw4i
gBX1EOvRuhgezZAz5Ixd7fBPLUi2TpiYDQQI35vQSkJoo32MLm7jV/vwhhw4Q4EYzxTTO7oHaMpF
DcGx97Fol4Y14yKdPo6bZVsNHjt8v50ieapb7vuX1Ig3WmaeDvyTDN3UvmAd6jBpwR3onPGHfkTQ
2jBqWnkepNTWVnQrg0+6fkBWz8P2FcdNAAEabO0c0agIwRnkgGEjmXCUz0ywfkdTGuBn8JvtcGbA
ExU9YcUitI4OLOE5S4eRoU/HS8xDjeeYvistqjx/mZ2c6ZeluJQzaWojK8XD7Am90R9C6RsPb/p/
Sq9IivZ4ge3+GpAHjq5FUK52pe1Zeki09WNqvokJjHY98HwUHhaIushKj+VguSZcZFimz28hJ2R9
xDMcSdOE/j1arBENpaUxLZJZoEOX9k9i2yDsl9zJRNv24tM4+sU2vxaSAkuGMg1FQuhb+9FfXkOG
cIwypqr/nglMSHTiq3YF5kCubAvTHznANPhpIx6oOx1VYQ0TkAoBLOQlXvT83OmAC9wwC5W8hoRf
YpRVWTsljjEZYXONA77VSS90jRfJ907lku4ZgzwNRMsyZThZXSXbTnS7LaHvJmxCNYBIbnQyO2N1
OfCYPTz2b+VbofKTfKiV4l267zNtuZbYRd5OtKb/BG4jldltY19Q9JH76WWycbZNM7fLbjPKyPm4
68i3TH5fRhDZGvutJ33ZXcyfrBlfPGXJa6/j6J2k2bmnQHYs/KSQkqepLo7Zp/hJnMriUJgIKpgy
uul+AuNsRq2QlYJsf/65Dtpr2AF2gmGIV1mrNcIBj2kYhbz+YrZyI1njzm6O6tLh+vPvFWFGhff4
DELagkZ14P4D+C0Ze4KjpOa79OrIC4Vm85KAphQnvm7EYFIRVupFvaHYVGXww4UHcRmsEXaPxsux
s6++8J82yVNUpApkCTGSM0z/qMQABaeJjqKfK5+w/qIQnfTJv3eclyqevtiBVQMZY8S+R1TFBkqa
qa1LxERVAX3uNPrGBH9TPhYA/H9iVY6y7bhqADeDmvyPbydHrCO1/7gf3mag7G51y0abC50B6/QQ
j0fWZn0ZsoxJmPLVyrN0aKqwaq5aehPXxa95oPY3Rb90MrEHFSHmu86SQNMyw61d+x3PBE0Gg0QX
RRymy6+bYf1Drh9zyRRkxCiKEmshmfXdm0IqE9ArX89IcNU5N7hxitzgyGSH78Bh+0Gw2eq8luZ+
SjWxe26E0tJGpMbSWqF05cdJUhISoUwXQoDiqltUJJ2iR/dkBb3iYV7NZVB0AkskYsLA4+mGCBnq
BMq+Py1Dz5jJuSrdaDKysjZHsNwEgJSsFOqlYDL1FrdXjYjLBNfNWpC2XNpyZcOosu5WlSkfYLJ5
brgosnVnvLDx/YaV/98pQWSh+ky28NH5hAqhGOtp4+fvKegFmNXi+zEuulnMZjwrMxaBbeZabS7d
7PlooLSyDHckzJfOaaOKj3IbmXYCSRYxLkWbyXjQFDva1TEVJ//miqnxzy9Uwxg5G7r71M8KLxzb
QN1mTN99eJHFMWNzalZzx3QF3RngfrxARJB6TmO2C3lZUJNzCzSNPgeDsbxbd2MatWxV26GPxP7u
oWbfnG2YaEYu8G4QeAO7E9HQEr3ruuQG7k/gXu+nfHeLW9zn1S0+VlL9BZ6/suLC8NVjoAorxbca
FLvdvG/eq0gMQfTdSbApF+3//eoZyyEI+p/KVZEqqoVhIgIPgHljXx3inbPsFhbEqLGRnXztkF6C
hFUKX2a4C+n0Qy7JtXSmFz0LsiblPuaVTa0qrfXQ5e6XiyOfrpbjioglrORleEXRZevLLGp9XvAC
IJWpNbsoP652ju5ldDWf4NXiIrf4SHua4qlABW7uC3Z6OEmcFB1JzttXwcIzXH13ZrJNYsFwlhOn
zaUSQCY7orjHND297HjD4J6CyaHyuKmgLu7EJIXD9fS3THk/TewRIo9g9b0WI2/m03bEIHNEZZVo
+4wItvRijr7Y7Cm8405CqaAupWy3JJKbumDfJgTDQ+4str6Q07XU/KxxgNr9nL07G1cLRAQQlK1N
Jn/YI/RyDPEoJZfsxF+FlA56+t6NhpPZHPxK34/8AS4HQMMD/HdgqWm7/b4ABQ26sw0wbvR7e4Ka
6gk/x03zDOV3SDgq3pfwhZSeJBxvIQCpdnLsjbvD8V6vryM2w2QOmyTXZRkNFTmhEufoi/lDNgZs
+oWKLR6ZhiFRnCx1zKSwECzCPGaLv1ccGBtoARFD6+j96ScyRu/beP2qbAJZigrELN0wRxDPE5Rr
YdTe80XCy2bMHRDLu42s5OUW9F1IgDFO9JVrh/mWB/xLN+/8uHcLIgMXV0pcHK1RtllCtDxLiVck
gyBacXLzHlCBXxP9EM/499DMC6gk++fkD8gRCaFPzTu6jNsIkHWKMeZmqKnzYZtQkeLo4MyIX75h
LH1kDEm0HLD0X1qY/cqzMzvlTg+FELH3dy1a3uWAvK+Tr88R7PBAYUKc/yOh7AjJmUfUKHvHDT+J
/bN/4JXdKRuKyFv7ul5TOVM8qJYohlv27lWToLpsMSHlUXD1d+yZ9jxsjQX6QWAzfhKqfsvVM4xu
TzBlpTfce1P0AUdvjRmEwlYthWdlP0ujAGtS4xxBPqSeyfeHWXokZ142J4ugXI8oP/98Wjm41mcE
4JLlnTMa7sOY8qhfqTWWUNBxrub2RvTeU1TzYXKUFENwPqa4hYEi9hpawNX0Agmxoibe0Egmdljx
h6UIvn1HFQK5ViJyqBBgkG1OLJYWSPRnGZD1Eer95rGyHLKwaFHnsN3nIWFjSUSGlpFit4g6MvVa
4VTFFjkJkiVBzkNUAH/V0Va7mIhDbgiVx2UKL+3Z0BFH2Koz+kxnCSyELSY6NQImuda37uPCFzLc
3VeIbipp+8Ed763ZzWXVOa2jGgj+of71BkfAvJ4qAHCffc5VV2MXm6BwrUgxjIJZDl/RNIbRQCqr
MYuqNlcn5G6PkAMzxbDUbcZvTpuOkSLUlFs3AsZIiCHUGuH34ND5W2Vtx2QIskOX2kZMR/5DAOsn
e73dPmTEZdU/BYvL+B71vPpyyWqcKzoooNKwzjwOwKpFUIwiPuJ6f6UZFRbmyNF4AqEF5qwT4SuG
0UNM1S69JH7g0/U6Cv0nsD3olo5tIm/us0rr3FqniemWaltl9uYIt9y7YIRx2JwNDqs1Tc9EBFF9
UrHkxR0cY5MN3DcPzw5fji8ZyGKk5g/pxFg0rQQpVVzysxfg8Dssvlq1vyaaAELrPdj6E4GBE1Kj
bNZuKVLzg2huaPSJCt7D5iwFiwbZEqIH5UKtK2jhfrqEmN1kzaEfOD+meec8Ej0cygLneN2DpTe7
rrwMojnh1EkJhLpLPxrb7irWDKL10Z/zrLVxHmiuZj55Uo71baoGcH82a/4xk/u7s6A+FJJN3MzX
1yAXVbqR2RR9TirJAPHCdPLI1gJ0zoLKFl81+RXnNOCZxLcCfsPc/+f0pU2uORrp/Uhida2/1oEn
wqfX2zXcQO5iUg0hiOucUtdGbhnzaqQP+ZLmUCl/iK7/bDgKTmnmUth62qp0llyfaGfaCQhWtq7/
qfuj3lLCSwJeG1gx8dGGvo3IuqohbSvPHojN0SSGMfAAQDzYlnHrzTh0Eepde3+fDtLACWYI4kmL
HwWywtV7jNOEcMgodVvqxVPpn4LEZ3iFQBxEduKCrdv4NxJlFn1D5WqxK5NbMks3hR36bxvYk9Gj
ZgRILlPyJzYadubtJb0c/sTcNJVaJFkGWvPCmKG5NUbJgD6kFbgLoOKnzw/s4crjPBdSa5m4eC8d
Z7mEVe+Rbx4S6v5bTcS3mrIx3sVNsE+EX+8P2bFAyviRdw6wuVokS5ZwzEJ2NauPW2L1O6mRIUIt
t4zqR69n/ZxyuYOHOTl+TnCosQq7fEhx38/YY0P1cwXTOu9kM3DumuNDtgySmEHZxQaceWw93OBI
XrH/Q5BUnc71avFLu3hInLsc1bX/V5SHrZ1p0JDueX9A+GTuOzay/7HEzvV7kCybYbcbpDMFf3Lm
xp1y3FW5j8XJ1mR0qTG3YBWbX7Z9ew7rfPaQa4wcKFTkmeH/OSIprgIV8Y451H+frB2YI7RC2G3T
YTGoL9ZmDXiSjVaZIidjGrbxKlKCpmHAZB5Mt2SusFYu3AWCOi8kYvZOt4LSx611eTmvY8pXZ6cl
SoLQ3BylAHVdI+BZWvMjyH1WnWXXRWxb15p61w/HA//AFlyrdgTWhnDjNvm35QX5OPWszk9WIYQK
MsBE9ik/ZW0jEFZXu3ox952l6WwCmPc9qi0P6RAqPJzJU+q9qpkCiHjomTXVw4Bp/i2v/IHXkHTs
5YK8SoRRX+/jyszr2E/qCiI+AGfV9ToAo5hPi/X1PYpBko3EuxDgIUOCmEWzjYdnTShuNkH60xk2
QbMlTQImc3VgP5ua7BtSMMRrQ4YUFXyjk/Kekyp3YKiSXY483bWVwH+a7OclGN8jS5J/vZ77aJKx
RX7w7cNhK7PVn73o0/7m97TGur527Mkhw4/cGo4bQmsDwSCj5iyslzancRSIdgoYlKtlMffmpYFn
gd87qNQFamoQwmLH/jt6SYMwSnKpcqa2ErxxmC1CoemDRIp4ps4JlqH2HCxEeIxtRMa9aXEsdRWW
7QWpCjsVtw6mYAxCOO1vi1tm2owIKkUqOFwoaZttKdICiveoQ8/77MTy6BEK3gey0xA2Q0CwOXSQ
H9M+Q3ojLV24dqJ+Fzt9U5gPIUtACRTOmfG0gb6Z/Q2Fy4bGgPURm4eBIxZk48bYZqTBZaC95jVS
s+QuIBayI2C5ppp+tLifSL0tzkbs76NiejAAax+vxyk//2PMqE5bAMcIBkDP6iMI3OvTe4w1DaLR
BGsmjTZQdd/wpDbpgmR/ckUD46M7Dtlp9NsU6VjxmRvimLQuiZx7utvPrSX6vaE4T2Am7HsYDJI3
Bzc/g5TWB0JRnTpNkQ09v56qdHqeUqN1F6Sv9EAvrdLKKlDUetuyyvlw1ZHJG1+XiMg7sd7XN+SV
hzK7p3xRfIGVl07MycjxmMpt0Gl3PDdpck5QI41GAyDAM6nIXl6/ydCbNxpQi+FcR9BO8Yagsgrw
400G6AzcAlEMvs3djx45T9iPFo1dGZ87qnbH9Is02ZXzdwuavCoQBtqRc1uXTZu8W2mNz77BGrGW
hfJD8lyUJH7smtAr+XoVBlOwaP2QSjoPkp+rp6SvXllV/EWbDzAzTxNKnVlyrqkkXiObbvgrQ0Qx
drHid7FMwipdcMgDX9ZHe07aPgf7C+RYjVCLbI3b0NtSjjLr5bgEGGKuEJpgkU5lIrY2I21nIDcl
IQ3YPy50VwPZTS+L/LaeTj+8cyWlTCHmZciIYo2r4b/g1iaqIbFu6MHGnWSpnLVWqDSVToUbRZS3
qbEBHd5KrRoWGRtK4irAAnV2OnunuohPyA54IwkLViEUldSu5nL/Xn3xCghiQ3cc82sIfa7TuX/S
JHQQvPT7+2YtyvrhtYQVJeVyEjpblBBd51qeVWZ3oMiomdHGaG/AnzCUP4tUyGubXQ/51ZpYf6yV
H7OIYjWXl62JBW+785/yRjPNQ9Pufj3ZJe4HZmujy85N1WDe4ffOGHEYEtcCJbtJSc3COMJG02Hh
KFirhVtGJBgMz5Hl+/xMBxVWZkQKK6/ugONzQKAVpPIq45VWoH/r9RNLsPxyy/W20R5nAtkVwU8W
DVJJMerncy6W4eEdBL6uVjl2b96XXhaI76nqib1keVj/tVXYeirBLfZgEeWrpzkN1JoXZtDh0PYh
6e/wRrN4R7UIHNYqasddQWCj1tTa99gsWyYsLE6N0uqsa5pHCBzCmQ3e1oqm8/kB760qhotGt/Li
S6eSeDg0kSoBwbVPi8ZzvhuvTSbitpqoCe7h0UcUHo9ZKZrl25rsimmpdRCpcK7wRftiFhBG2B6P
uKRSU53h0f5hjb8j8W+A8Q03vWO5f4Zax+qNNUd1afdZB1XEbWrSetP/BRNMu8pUZ9yonCGHRYnu
2d36A0ixYpXhprdgwl1TalC0HlnzUBrenxhUT1HMiw89Ffdx2TPepub1VwMeTbMEdaVRmOPDQg9v
VGxSkb+NAc+CqsYWsoiwmNEAX1v/GCtIZFJR36Y7QFyb+BO5dTStlupu69swvRtcrVu9EuIp+p+0
xoMpXlTO9kKC8s1ZGGpd8shxyN2vknyYn3KBxGa/rTbK/E4mOrS5QSRQqEFWNAkER5Iq4GRpG/BW
l5b7A9++TfRO4Vr2eGEzeOgLlFhmJ7pE1BRL+Y8+jRYhVnsawFeGeB4cbLdGbnMwGuI18iSNIBHj
MWUArkBV7uacxxroiiSVxIBKVGV21/o37lylT+kGfVf93JsFVhkw7gJLTLWTCbk4OPkNTXergJ6H
5gtlgOYO7w1r5oRFxjBnzpUQQtjoxwtFBj+TJWTWU4KeYieGJ20/nkEcxN3RlEgFv4SceuTs04A3
h4atmzwnrC0LfwZ8w9n5bqhVIyX4z0wKJYYNPpUK97mJUU1RQ+wupZNcO09y1D5TMWk2q8po9sB9
9ARyGIxvJDhGAyMAnHfuOprnTfxBLUpnCSEnfpP7zLO/Wp/yeqEaUvmZUVqNdLPVCQKoUQW1t4OQ
tnidaFraDTCTDXOvAW6wkOcvpuGFKjDBOsAl6pMIS6vQCJ315ee9zFyjfMAriDAhfdsSHrq3eoIY
/cpEcTUPwVf1raL1mWZJ1aGQC8zZNxx/ITUPjmYzPYo6P530o1iICEp+F+BXLl0lsVMWA9L2mCav
iaznjzfv0pLv87PvRcKrrVDz2yU7cDLFhxgen4M67Hymj5vt10LuFXavVgthIlq9/vTPeXBUN/ic
1J/RqZdgOr5QZM+VIDSqICFJwKsHqJl7Mza7bnS1Q+sazzznYi9k73QiGiVaK77OljPqg64Q3pHA
r+g9pvd+L+6gaT21CvtNnfqWE0WrYBcgDyz/u74TaSA1VGCzQ4tIuXZBo0SDC1kTZ600nr8+imfY
ZKBPMvkIaiPqeXDnqBFSo7UrKWosm5pJAzgpuBYxuCsml79nkR9SU522HsqQlLNvaGQ9uXEWy9Zq
KLBbsqOOpfalQvgFRWCe8thIOf9e/Wnqr//HdHv+UmBrmFKBiJHblWRUHiU5VSCSnzrmzsKhZANa
EAnrJh5l2HfpcO7MvLYPXfrEPPWDKaq7bbFRL2f0acLU1olh0niuVpkMcJrKdDOLhbc3UaeIESGn
se832dQG2NSHHgZ7GHJ9iVuCRvO40tVoePwy0m1c5wCxNO8pNLstSd7Qp0Lm+LXP1dZ9/Um4T5sK
VY4xmHQ1PEgS7h56nBMJMU8N7v7DFhNg9KzwUdV8xJNnDptTdlVaMEPqPumtz6bICaNjc7GF9puj
y08NuCSQ00V9dAH399xkxV9sCs/NiVGBc+cwud80OZFn0KSYcTw5O32eoH94vubqZxddzazBcC8B
P+CAg20zAT0n5SePDmXPSYHTj9dA/p3pBV9j55U4uV8AGYm1f1xzkNs6OF2bCKjzvO+VkG6lkS9x
uNu9gnW2WQiWfMOm67dwGFnJ3ioukGEJbwFEga5eSbrzlLXARzuYk/lUT+364mYI433dvjZqzjju
4hdIxNJ7TXdmAzwUK7vLjZusKP9AD4IxI5HzVEK+AgDKXy8Hy3t0l8YZPbGCxeq4sYLyaOZ495hm
8i18r0nP+ZbrLWsk+f+nJo+LvPxgQmVxjsnTimZ1cBF+gAvKkj06T0bMudvL9Q7OwMSfb9i5wEPX
KILQhq1/yRZhJ/E7Q95rkpNisWgsrOBlkv8Wt42YGlrXnbm4xEwLwO1+eDP3cXvt0KIL95C1emSk
UPMyQx7bZ30kftyd1X7v82t7v1THUaRMCyc7FD/p5utqv1dYHxTjBowkZnzNvY0URVH0qpGae0re
KsK08l8mRWGJyzDFOFSyx1B2vYxRbAKZAp/ChldrFXfjHZWy/MyMKZHQpXLSjn9iBGVqLfoVlHKF
WCoN5EEUz6n7q/AfrlNZ40vNL9gJIsY+XASPWnVoZ8ST2h3K1jA6qTsm5yVNKIhIhSfMEZlI5rWg
qfd6xSSMCk7me+10kshPaDEv9xa/LrbuUnhqUczSaDpsvI2r9W2tsroM3vI0nya12d22rPS9x04y
h+KvlwapPihteO9HND3q0UtlqjRWfyiyss4r7NMaD/diIIdYk7NlHP2WjA3/tYvkSvYtxnrJ4JO0
wph0vCIC18Jk2/Vl0zcfnYhuxE7nMj/eVSKQ0SBWGX8CG1y0QcM4Fl1d0NEKjVED1/WYqD7x1EoK
tkGdPoab9M1SeYcZjKSgh8c0jCUQ2QaCiBFTnJ1qMl+U3V24c0jnn+JXmMHpbq+6tOl+SCHSCJez
EBKZkZOBlHBnO/vub4/WQBwFIUXObMqo0u8lAOUnR03erPBgeHoV65yzR2lxhD8Ihv4KIkDJjNUb
iodQXcGBIKzOuRjtX6D9zRMHU0BK67sQ9MPbL+jx94h4W346TSDOzLOUpkIaZnDtIgvfRkT0SlGf
ZCamppVeRUXRubgd20vFkI5I5wPTKIZqY3fwgMxlHDyHeaOr7Z2e7aVctbb0epZmWwSlvblHoIb+
VwHLf2VqYlHa3JeUq9sPRyhcW5W49y0O0ePdQnxmVeFJX0FTQtMQgnsnK5YOjy/oawpmS43L3M1H
AXsVMhff79MQyGgWR8mzqecrPfFI+BuYnauL7/E2kc5q+qfim5q9vz2aDdW23vUNDh5ZeKVpwxt8
wbmLZFkLr8Y3Pa4YFNCM+VXNr0gwApwQu8wf8EqO3MQSNAMA8PL8GuC9SJB/jN+MtTY7WKuXF671
Z4/8jQ193qKCoAQNxAOOEP41Fo1ixU0T97AgVXrylRCq3ZjvDPBUhnqZiaUqaOqvAbSVzDWJtscS
3SezjNUBNsGJTVtDowSbKfBK3CXGu8fuIvqo2JZYWg1TijjWabRrOKYvDXwfcf0r6/V+DvTHCWG3
dYpI2D9ZvwEvMyxkucEYXal1/pkO+FImDgRasRTyb8Ar9D76jeSVOiW1Hi5zxiFe2/te/07yoxh2
xky+HvdCdVZbLo6lz5dSSTBtO4G7QroTElKduXSAKGVI0VkL0K8mXV744jKSWjuj0Uid+1L21VOG
j2SxxJhoQAEp+T/2KlYJxNLXVOb3c5l3C+z+abjcnm4IbihRqvNAJfDWTfgHGa9zvFUanD/MpcCR
sFohN0qGZEzCEtzcZWVpCOwkANlevUuI6MSH+zYImJnmY3WHiIa3u3WRO0/AvOgL6BkpVkIN4u3f
jG9E0fYzFA+xYHnYpGSsGz8Y6wIDrtpA9DMGP4F2horplyoGGXC3HGdFLsksGqYr1rhMs8y6HdjW
74qNaxtcTbo5hfAcK6DN6r7yHj/j7ezIikkSe5NN0TZwJGuV/Ipf4bXvpeoY0L7WB5aEZ/7F5PeU
dpekAHPEyv5gHuVQkFnB6KwKRFsyMRENb3n0As+m89E1JS3dXtpWUnHupx/m681v4aZRzbOHFA9W
QpbevLMsAai8DlVRk30fd6zeB8S/YUjv8lb83Voud6Yzxo790eskSal9Oh2PGTY3bI46z2UIz8xC
80QWiQxaefX1RALpb4eH6OmgklsJv0q9aIVOMd3BEB5hsG3f4FYUZtdT80meOdEwMKmKvaXHsw+X
bhRSjf8T8eZLRDKj0VCVG77HlnKggNws49OrGlyx7XATpc4PGegKld27f8q9/eDJHhcRfflgDway
0TRzvrIlcghbZdygsQ8mLmMWxjoFRWirs8nMjft20r38bLLv5SvrsNTfbO4Q6+LncSj6/jVrOzb+
H80eXtXNy9/Ghe7+fCL++7oEdRjsdQmSiYH4KLjEce9YdKPCF3xYTdpWzyYTpbq+b8nB12aTUk4y
Ms9XWfCOk5+UuD9ZSP8p84LLknRLWWLayJcFXg4hbnRE8B779WOBSRBTDnmFf7T55dVIEKQ+s2QB
RJD2QGB5kWATFmAHK8ETCeeUrSZDwc8I5/DDc8iUls68+1pu2vM7mxx7oVT1eEdn5qFXPC3czV+K
kCwGBBVOdG84//JYzqUD6TiyBfMBkow/ktVoKgAerhT3cPm2Kl0XDUSqz2qV11MnlcB9gg5xUg/V
KbtEXklzI6rbDDiNMcpzSnQeouAuB93vREvXWnSfN610scCjjFjyjpR2FVTAGjlnmLqk2SAZrxnt
wgZUnwtCjpvDecI4a3b3j0fdNR1YnTmn2W64QSihHW2hbOLIeodF7av22jLyy9ZlUVrrwZzMzLgx
hKG0Y8KE27Hsu6W9q8eI1+F3sOViFw91UXZk0NRMA+jq75XnPEK87aREIga6PNKGP+4CltkEAbiL
SHDbkLoUkcDdGpTlXxIkUhKfQMf4AJKHQb6FRbn/6cEBQ25Ao6rd6WpsvYnXw0NKfmXDm/VLqM4U
6Sq8Lja6/uLIVcshNaFfwDQTTzjD46nMx1Xbjl0REKgTkOyG6BExFNWGJgx+TUpv+BDf/IIcV1AT
ivNkw5xFL0IwA/04ns6rDFIXN4dNO8PGuQBGcJ8ANGxcpbg2LkruPHmQ6HGAn6wR3fNneqXyyoTp
+vmRg/S5tAf5bMAurmqVLaQH2fJOPvkP5kxLnDLJVKw8UbyAasAlgNI5XO1SbkCpyul4ThUG8bUW
KfGPuxi5JYZN1hpuypXIMwFHRQIEqjS57wACl8NYZ2iAV5f06C1Uv60pZQUtc0PQwwl/zsyEzPpe
xlphw1F6eHOnSTiAS7LgWK7Amb9vxbrer0DVvtm0U+xcLg9tZuew7MFAiZF6hbTfi9vfF2PtbGfA
acULDzYz4GJ5GvJ80qUP6RiyT0U83ktw2K+fIWhdFwA1aRVAwXkpk6ISmdRe8N0sIxdpyodmRtQi
NlEq5qUTmQktpp4Fi6BRQw29EykpHn9X8h51D+6aQQXU+SSSoX7D/os4LWgQ8av6b0efkVdCSNlA
nyHhu0fdGK+lbVF6xUszHq+YUgyE6cKYQeEjkVBqvnlP0ZLrfwDZUFdeNDgf2mwMXzq/Ycc+5B8u
Yp3nrbG2FGR6ZZqRLSHjahZ6X/4C8jTybAUUWY0Y1CATxPxru5092/caduDXGyJzYKGz9jkvfjSj
IclHD/0cWHVuZcKwUV8n6uGpgVZHy3AqRW4mguUaOsxFLM4y+Wn19/zzZXAO4xxdDcC7W5iBrOHg
6Di+CPhLXyCbcHEJBRh5kzJkoDYjrYdqDBRLzMt1kkqN5BaofPEQE/+q6Ru+RPAZtHi5itxsK6LR
lztQwSoaYch4qLhrDbdUUXuXdwkhJceAJSxIkiOWrvyamPiZWjYzqLuB21pndBnGaqH4KFTpzwPZ
bx3Ly0NtSWlGaBQkQJnpNv5frHP3mAypYoO7eH3eqwYNetYdxlC1k+mPs66iBBB0VmPfxINf3n3N
WZicFRLda/WBSJw9EefMXIUE5PVFl8nSjjtIlxt0xZklyrQtSgxuzeNCGpWpUqlxyHH8DxjVbFma
rLdRrq0DKSnVdDCTRn8Kt+uvl3Y4bDsCKQ6XYyPk72VBsPiL+bDmlHoH1lf/ecfOxQqXnhMKAywP
tKVRTd/jour22Uoi5SWfnnuWbqNCZ23XDgZIAETUEvQ40sNGms4N09OVaLjt3GTbCRJ5D40m9iZ6
yfgcOaW4tcdCbLwEw/wvQzOChUk9LBzT8D7f/r9nLKEtKGTd1O/ATKjhFI9KY4Ts07OeV0W9Z3q+
a7NMW61r47BQhBnpEkuEkPLoKsetTN2Dly1yzb3BrvLYwaSZf2XVFJQaIvtJgpdle7XGPbZ403WM
k2GNwE3Sgs3qmSo4VwZSL2n0ASr54ImqnbZNVsdEG7zm1Rwqi+AUUOvBdlN5OOuonc44a8hHCTcp
o/zU4tcGvuQYr6/QWGZ6VAOHpHR6QEwlQrMmyE+b/+tf2KPDQABSMTx5sPeV3k0bthISgLUvPc6x
7dX4+qPEoojtqPJqp6AUqHKccd1p8mNBTk+yfL7vP7kUR7wQxPAWjdnV/ZaDDChVOj10YUx5OHY5
dcbp1IvQf1M2DNnt9rd8lpPjyzkBqixWm0D5yW7dbQhr6Qje+kst2KTjlD5gvjukatWRrR6xQr1y
7yf0dTsraNdEIl6kQpFx4qmmGzTxcyGb/aIHkrVh4DEBnvXiZ7+Mqq3aL9XUTT2ppd0VQadbGHoX
pBloQF9Y3K+GuV2vJYFs5IkmnAkKnGhIABKOTj4NZzevZVsTqqSweN0wNe33PMZRzXYyEbR9dyME
n+r6V3W9KN4AAfQmqG6llbynjLWGBwgT4iGrKUif6+dKVVtE0PVgaAzlryGmEgiud2LdZwrY1pn4
6Nzqi2jwRZnWCqpI+NLGBGI+Qh1D/ysCn9hWpPJhntqBbR1nwK48ORI4moVUbEqNx9mkrCKci+Z0
wkHzcbEEezM+dMP+k7CsoMpE24M5K0iQiZWUoWCZhpWaVhghKR4W9o5l5X0ExGiUbUWRh5G6enLd
KBcDGv2VMJi9caIMYR21JegebPk7z2iq94mZFN7deOCDWyIlMRfeFii9PXdLIIQTezMiD1vExISY
IXeRwIGrEDC4LkewXDpHbKnlcI0esPOD7xNHTlwRAHJsxIAqLbn2n4V81GE4njFM4gdJ1xdds4eb
0zT31DtKCk1foHH0/d0IFKE/7ui03LrCJ6Jm4xWjg9LhzibWl8az3JF4Gaq33Zn4/cXz1IqXU1PJ
2DvObd0JMO1UXXve8cpCTKXxzn4qhpcDr8PMJZ0qzHbPk1hvjdgAtt1B/0tKC1cb4kWtE8T5Lv1Q
QrbYoZ1RODm7VbsFlhodZPzD/TdS0LfAqabNFDadJpj6z5Z3ZZToJd7AXmrVsrJ7lF6AKd4f42RZ
mC5Aa/EubR2/9tlvBtUzzHZo4ZexTfVk0+WKytfRgj2PKUu4R1KcYJBnsJJeUyYG63ppwRFVIZsV
RuuCShVFVJgzqTZqLnRv0i7F2Idn+1IXcnVJZVNFfQI5DM1q++qO6iZwMDpoywO0pbZTEgFu3W8N
vlL9pE7WItPqacfSFv5fD815c0KE8SQQeJ5uEk5vGVauPAa4HBIEh2DFRvvpX+blS/GC/heIJ/1W
m6IxLgtoN/w3xgzKflSov19Z2pr2mB+92th+EMN5HC71twjgkF+jt+FJxpuqQTKyVAGld65LcE/y
y4U8ptnz1s8tmm5Cx38z/CRdoeh+QqJXKHZr/6yFSYyRzak3liXZLJmCVOePv6wZoEyxefer5d1v
V3faUf8mx8aMYGfTgshfOGzsYhA6bsi+D8OL6SBxt2miTvitS2/MnNdW3t8C8usdvW2/35ASpz5i
tzHYdyCABaLQ81Q1DAHIDbdUafnaaTgJVqJ+o2wDltTjo3uvlgvUBYEhLEnTXs1zS88cyo4MBLGL
rMlbsctx2Eq7kO9mWiVYJCgGcPc+HI/1nGlRPp3Gr5w9dqQsMSzPU1MFKCRakRigvqdT085ntEXp
rMuT5qtUXsX7PQtg0XCMm61SWAeGstK2uD7LGqX/PD2JXt4F1NqVWzlFx0k4haAw9dkqufhcLxzD
Tn9uYM9Ir697Q1VD6ddUc1VzxnIalzTlauVPJiFTWp88m3jRJU619k0caw6ucVYfV6ThwpM7k80V
1to/oSUcP+coixjwkaTssW13DPSPpbzJ8P+qfBA1zOMyZR1mBPOr56jca10ZkPcLoD0K8il3ibaF
4jb0L7ob1YRchVqB0WMUGzXCokDJjt3EI2X8ZLsPzdFXKXIWKpWCI1E44UlSJJp56ki43lydxBWs
73MCjZf2Jmm2bSvwdAjLzPdoBa5bwOOcW0fqz9kNC/xo2a9A7qu0JDWZqW9xyCM03UkVjJ50kRYk
nqTVxZo7zX06PFYFil+wE4yl+20CV4GTRlwuPFkIx43c70bTMllXyaeqFJ5kx7agsgpt1KaPQm0R
urTTmvRjmEvtc7JWK979ms3sLmaRDDgsKCMJnc0cZpBrOttNn7mB3zrs+BCrVFUZ8WDDZmN78k7c
VwMmTrmKVyhDyYtVx0mopxEyoe+lFH9KZZ7tRYcVCAECCLMtZRoXID+L0B3azQm8vE3cr1twuTHv
7wHsstLLFL+VcAe11yo+huAJ7uCCMJob5kZBJiqZJHXxZ5fToAUK9/sJngIAStiYiA8OB5tPu9Rk
Dqumr2DDuB2//FeFXxvQBGo0IpjqGxvjVQRQw9Y1kUnwk5GfKZEzF/TWjk80/+vYladlDBSu5GI/
zFOSg0JAPiOxe188oLG3CuURpXgGpX0m6bBsFuwZbLlFTwDBA7WGzQbxvdKB8dosqZiMFpTz0Hho
Fwgg+zqnUaATGl2ccAindPTKSUpFYqR4EWI1VgTqdbGgxjJck/7OKnrcH3frJkkppiF7b3YuGkiQ
oe2ssZJSaImWGrhlAX+/5bTDuRB6QRVAQ/yTvipq88imveLLBtVE6qdtCtEpq4buSx4OeZlS2VG2
ltVAc27ZHD1bM1sitHXeNable9bRzcZTZpshfBLEa6klXj1SfcTerZa6wG+3eO/sMyGwQukH0wD+
3Nnm3hhKzsi1PmyYwBjZwPLETkps04lgF40wUr1YZGeRFO+MmORHd3wS9nSedz+5GvW7hwWVDkdf
RinB8ZnsxTOsZo5yiWtBixp1tZ+KTeq6H61H3YMwp3Ssl//EQDUWKz5nfAB01gFLeksRhtz2kKwW
Y+g+MZCt0Gpl44XKfldqU7f9UG0A/IX5sSHjRINS+4JLTyeyBeicKRynsOd5+pssEsA4VOC/Srkl
c0IjAQKDNtJ3d65z9mlUJkB4gR4bouhw7e/SRDL/CANTRJjmc1xKFB2czg3ex1qHV774MY2WA63M
k62tw6YRt3O/o7WEl2ODRQncBLxrEI6b8iKyPtdM2ftHugFg8tJbmFGSnp6MuKuMjs/dr82q/gkt
Xd/SVu+MmfuO1HzAtlphZl9T3rae8JcHn1+6b6HfyyfZSpVaLww2zZEOwqgL3knejty0g9QBVP7G
AxQi8qtZGJuCW7R1V+N0Kleb01xxfDDolg1/e3MTarW6VhR33A+BO+zElDIrSTXZLai4hGhM6W1I
1xGTFBLBGH+N7Z8f8uGqLa23jgmpcXYpxdpW/Gm03rmD2CS8Iv7GAfC25Lw7XsFhdmJ5TJnPOfp9
wjxbySxGQWN7x5WckOCno/opyZOq//AzI2IVaT5ZlzsO+CeN+ESWrfjY4bn5ma7YYk9QVBWDyXYt
vQr3peKutQ5R5IbOGnUW3gzq7cKprrUVvXHZwfjjsNLsm1o44HatqJNBsKmeADHDKPuHfrsPqDs9
hVHtA5VzKByDC54y180UlrhAkGkAEnam45+Hxt4dB8j71fcvHSq/0b5qA3hQmQ74tN+/0HgMFYsT
Cqk9o50Kygvpx4yACcgbbxlDKZ/zA6xCjFMeVtD1A7+ol+oFbfoheomXM+TZG/hZNO6NDnwrUZUw
jNY4Exh+aEr+GbXUojvD7EYSlehk9NyuKcRXBUa3FnKYf473N4gUuG1O6EWB15U3/BtAKt/DbH0w
uqOsC96EEIDz2Oi8uo/7MKx7eBsJwvrj1X8HdnhLk3KHrsBivcsLZ6lMMwIqKNV4qhxbRmFB+mVp
I8JXnRv5gaAvJgTWYDsz/3daTV2LpQpERR/9KHYMEz+kr6ATBFEHY0i4nLeVnQMRHP85HS3U64vb
O3TwihLd4swHkaFn6kcJ/op3dmFne/Gh79N2VmPQe9dqmodYlBOaYjrHBgmVSB326d7dIRBiqOkQ
ov17W5ZHWDlWu4z1Ph8yr1/CW8SlyQcSo1VNrg68xHmNohep70Ww7W3x6yclyWjVl3F+i9g6Xwt5
bFnVd3SNpOIEfoi6MR00rSgWAEJdx9xZOIRwop6G7cC4LUpT7qrqFFhmwVRQUcJAlRVHMMBoQ7Eg
CqDddlPAmhpvi2oa4Cpzp5/OWjr71ICg1tTFMBKNOkNGBvC70JPPsB71v8esNGCzXjVLGcwhyv+X
9vtOL1eccWx4KBBVzrUuYgCmpV3C3mni6J+26WTCCaUZifaBZi/oeKQYs+/OR0B8Pg9sbZrN+ivE
94dcMiBHtaM3/i14xxcyp4SSyGd9yOcgLiN4oic0VkdVJCkIjLlXiinKV4mRAnILtX0tNdGmzR9n
zQZGBrjZzvQi9omoe9sHhwVOHbv38KrdIu5NYkqsd6EkwMEb+ASc5ARhxd/DOvP3x1uNKe9f5NOb
5WQW18YYosszYAblhEZXXULQ/OCugu71A1hWcfSOslL9r0/zd1XjDyRZmqlW5tgkZ0zAvCUraIT/
iWl6ADRNl8dn9BT9pDOIfgZ+8gG5jJhyjfOQhiZ7ai73xtFikpZfJUPjQqrCuxAjL16fUmGAbaX6
qSYkEAgkfukseWgOL5K3FXmQtadE/kpgNBsQKYtwxk3mZMjnYba8KIDytP1cKdqe88+1xXrnnF4E
z5x8D+nYa3SaHOJw/54M40fpC8LTykqQcKBei/vfJmrCp6pnKaoGEU2kl6V2qkwiFSFmwss6InD9
u7d8HdPZH2iVt4Y3MyuQwUFbUuwbwRBFgq75BVcGkbdaiNe1xBK4dioC071z2iukceDeKBN5N7Co
qOjWFZ8w/8txWu7YPhgke8MejotrAg9MEV+tbB0wi7OgKykZ0Rgsx7+/yDlVTeVMi5xvnQe/m65w
bOUrr2u2ODc1H6H7lcpWInOEK73BEmA49ZWd6d2eYnchrqeAB0YZn3jPOvul5rxCL17q7kWKDwhz
H7NYL1uRdIq3HLXxchjQxtE6o0c61c2/INi00GYLCL/3+j61OrmGhskfFCUOvDUoNutuz7j91SoF
CvFpeyiI3/mEMr3Q79ElZJsF6SO0HQ4yjeP9LSGxa8kYoxd2kynawgidKYS2Q18sJEDb2Tv4Lh7R
bmWhv7T4X4fg8SJTL8AIu8esAN/rWalghtbsqsgWgs+lpGjtr7k+LWO3zNmvb3j+BYIl8q+f2R5x
6W3iL4JIENYOPXF40f4MbPmydGXoPXot82xRen4W2iaPksYFC8ixaYkA1P/4IGGfpZ249eNdg2ez
126y+gwxNAuIV3kfcZ48Nwl7XxXFCCtJzTb8lbGSVrTxcOIpgbdl7udbUxCVfoc8CqfL6ch2OLC3
w+BqHjLAfpfgkn+/DdyllUcfw5x4vNn7kAQAW1VGVSCWimW+mt3+rJ6I4DEAQ/HiWdr5a9itUyAY
eOnMO2T2AaVnYHDzp/5m7quZyP0vtzQ0IT308HfLN6EdII9QFYsP37ogc9cLAIKXypv7tFQxiZJH
PNXPxpOlMuRmvz50J6KhmZ0lcd3hs59Uc4H8tuh3GdvQUrgX/U11q5WPmIxWYXCm9eweCoJDqQGw
b1soR1IlQWlPwxHdBH/FRum+RENOzt7/zamBnixQj6/8OrcPVy53ofv3QrMsTsXOLOpwzmiIYuSA
b22a/1E/g3iqrDnT0y5rQauGsQ3CEBhmYF2yLRrmfUb0b0pdNaP09mLtEhd699IewDaXisvBzoUZ
/XnZPMG/7RQ7kbmQnNsdu+19e4/0+KqEHqgKv+va9744CICh7XUGODAM28NwL4G9YrR73qjMpxeH
BkljxNEnW7k1VpFwc99fSbPV46KZXnqgreLrHi9MPWBc2FOw/CLy8Ht0DHdTMNSeiacG+cTc8ZFo
B59hQRcrsvpMFlrsspJDetn+vfr3dta4XffnKkZhPHmFTyZSNY6BpXaS3gyZDaEEcH59eKMiu13Q
IH51m+5jbXRFVBvK0i6a4/iq4ix5j6j61COsXNQxlWa34jw1HjPkhR2oA8pfurkrx+5ZP44ImXOc
XbkD35izrFMzgFBY9EJnrZKpmoU6iQXos+N9F+/DVGs3SKZkr+XMf6tgHN+Ty2/tonteQ7fzUOK3
bZtAqspZRTkLEZoA/hsv6VgwVEB74hO1hk1VF3M4PXgZb94c5hMuXnlPJ8HHy8iWQaDt/Kilx/JY
Hxpp8mWhgt9kDQEQHB0cn+M6v7IsyfY5POU6Yg0J+DO8jRFdYGyZrQHvHzJp49R9QODPX4em5eL/
TOaaQ4rA3iZY18/Qbp/ELnE3ygRUeTEcjZFeP8z9TB7iehrrw4Fn7SbkChij0bWyN0jDw5bRZvqW
Q8w/fio7c55xd3cbW421qCCX8thLF26IPPV1gUDF0Eth9v/YqLa3/ZlVn+hK6+BoV75T4jU0McdP
qWd83FXK6OA91OeS+JGh3HcsIzjvWUvhf/ZhNBeCd3LZRvaibMlA/oreUxgJb9bDOGNFAh/6GcC5
lYS2PgVrkZAI78BZBB79wcVpPynBAI7PUrnFQO443maOK6n3ptPPrqYy0KLFsSOZeru9nBobkop8
xrWa63Iau0i60Fs+b16V+bHWUDksOhBP/hOkx9Y0ZgTATC1IjYnH7sZTBipyNz0G19CUnuSehTFX
gGpm03UhpMrZPtjIAt2kWztmm3TxAL9+SVL7oqK3I7Rur1MksgWpKF4uIaW/6zh3ei6Z7Xd9p7jr
gBBy1zIEn68xxeRrUgw5gvCEoPCExZB8trpkQqJ8Q89Cxnqsixzt2CAK4JkRnUgtz8mI5zdrpRui
j5t9jT8n3b2cFN0egbN+CtRh+x6+2jO2iMhiDcw9vA8LNhBF8wF33ZmAWxKNMrGI8gd+GMb1Ef8m
nFBuvKeZX/T47TuzRm6X9USRUO5bB1OZ/3XNgK6MFd1yGHIvG0Q1gKxA7rkFTrn+/YZcG/9ort4E
OVc074qBIEB39xRJ+xu1IuhDBKVm8JzD0TgFRz/Q9UZzjFL3+SFDK2PM17SvsT957vUtxTfneQOA
hQK60hiQpCu5WpmGBE07liyVOOfwiG2FgeKWlWxlf0U7Iwwpt3SlpbfaV4L7fnQ77MiyawBEi9ji
ZU0swPfsmUfTMkKDTc8cv63LL2YM4g5tiK2rJZcWNOuzZGXXgvOGcK7pbzaQQhbnYjbRgAejNUQf
yq07HAABCQkwxRV+C4IsRN9RoTyBpUGzMyGu0KGxQ4Fl067VS6/DGCihReUzEev9wqEAY3udNbIZ
bPWD1TTW1JSzBiqlW6eEl3XvP9j22L+brWMKzlcTIBvkZeYd8uLppUe+XCvMuMUgG3anBahHAvu6
P0G6rL9hzgsx2QProZyJp4E9XOnll+7ammsl/V8YGDIpYEDRzEaf5PFFVall1cooxdtZHqHJ0+eU
tBTjD72qewmUyGxzcxp3FL7/BykpDfy4/HC98VK5G98iCksIE/fC1nxQtGb4LXH2iVFi4jQZOTwv
d1dMSv0PV2VPYmTO9JbMRk517l2BifKgsmWPiITrcrFwgShoUhY0YMFGy3Yrkxlgrje3Xmwo0GOQ
S7+cPwOIdYw3d4+h1LQSfAycThrijR83viwl6k4NUL9HPkAerauovnXhyKYOma79UvuIaKCl68x1
wCTCrMls+1mCYWaz/GFHLpwjiH6P1w0OHPYNsKoRVWsR7QC1Is4pJWqKssHPxUT7hg8JDrsFRj8I
E6CrRZtNTNanLq72x29AdAjxx+jNULq4FJ3ni/H6mk8b4cEH/c4NoMm+HCkhbltAcbzRcWUihHjU
fjr/eIZ49vEWf+triCMbwn/dUDA2YAzJ3tKzcgQ+mT6aEqw4mq5H3oowSt5piKw0rG2s257Eu9xs
CRuHZxzJmhbAGX+icyAJ5xgR9FxG15R4bOtzAW+StN3w9GBNO/GS1Jqu8Lkh6avZdKZk0/Q2Dls6
cSoUHNAr6znKmuuWGlNo5pV0uRGcL/pumoBTR2B4jNj3osnPd8mPqQ8JBYLdse1YWyvTra1m0JuO
gjIv57v3OFcQH57aZEHi0aQeEFrK4kcsWnTPlx/CsPKDLVGDMLGrhHOapNzfF03qOTQRpVuuOpKm
MM6RzQF6FKt6SXhZ6fAWnyf/BxHSwHFPVCtm2pcATWVe8i5ptP3cjmeLc0c/29KnhaNMg9Vge6+q
yd+46m0yYs1280NUKRr94b1A5Xwv6wOEmF0gMndfUSw4XjSHcPFTmCdm2UYs+N8C4NqCa6HjAEiN
3202SCNrBgro6fieBJqyj0K07LnoDlakuFKE+Y30Cl75OrvWfXLLZfevHTtKgmN50q6UqPY+Xy6v
Bn7kBfDm1Cd5CUcXb1++GUAXMvVmVUvFvS5VwmD6UQlcEs6+qSVPgRk2T2/FSXHuE3kqYQ7lGZ/h
y59YhxFrfPF0zAlL760Sm2e+yHLMz+r+lyx9BbsnrkJZt9RkCfOCvu/VrBB4LIu9y+JfHR0LY5qf
MNcerjlnsVwrUv3j+xacN2B4YRWqaZdMOGJ8os7Fqi36bx4Np1syG09csYIT8i/0zifEFSAiZL5r
NV5xBKP9kYH2tLyXZ/SvSQnbt9Vv9+3/LCfjKNPA2ObOj0sV0b4AlnOV8J77rAG9ZUauYUx3W6J0
L/2LpAyAcM65yU9HoZ1vBWbrEgvR5pvmMofNmju4+OXuywMOqqIT4hlQ8GTysIXZeg4cZqpiFW1a
ZtMxHnkOokLB9UUY0aZxJdYqhBvYC7NbR3CaXQALl1AHbZuYIgkB5qYGyck9qqJgCYK26GgEWBNg
RVYRoOnm0irrEbpnTQW/8HT0D1zaYwyCkJXKIfUvWnQtEcTgc5QQtfTpWy1f49E6X7L+OVCaKVgX
aZBC+HzZ/nbfBKE1gAbGZAgMmAm0uR5sCcXCVlYS2OYbqS7fHdO7Cr4iEtwET5fU2RRO/dN9r2SU
et73ce1qbSqGk5aUhdmKWlEc7lwnMlzkJHkav+T0KJQTe1iASsDFYkF1ZbjSVlfooYEOVil9cH2g
d3XjZUaujyjoWlLE055hjReRQrIUB3c46+bTQfuyzAsIE5II+QMlHPNYMg0WaLSbBu4HnVPsSGVN
Jm08sdufc0tHNNEBIVybgRAsxBzqXT9DRj182IIFw+nR/K/As9G513rmjxBzU1htqAUFMs6qHxJE
IehIjUFFoY/mouxos+gtBa4kTxFftxc1+wdhhTwlQXNVk55KxY97HlX36iZIiKSMlXKy2IX/U6t/
PhPLFhwuerYw83vKfMGljx432cGdbxrBLahYFeNeqsFydmQ478oVsegKxUy2KWyPlj0dj3b09VAe
DyLJLeZQIOzBV/Nhiwez2Jcy1/mXUfmkJSXz3b49Nu0t5m0AVayyiA0NkhzkDg8OucXjzPmBuMl7
qIPnxaRXiFnltpuQIUSpEPkMKcYQD5936eVUciAB7J9+QSzHCFMtMpnjR0pChj2p0zzAA3sfwFPg
yLcfwq+5kx4Jl0deSL9OTosl0W/MPG7hNKannAgZPgM6kKvtsQZ8pZmEth2qmTfjcMMTgAuZXP3T
A7oOU7NpwBWDqLXn/fWaT88X6WBnSZifPNaExUqLRDIXzESriLrrZRm4f9dP1bWWHSnrdm9UgSmM
KZVPhCxjiIUDTbKNb3ZGiDUy+2+q3IQ11wZ0898XBkd2BuWfT/tr6zBDWs19PXUjw2bj5egpf64Q
ePzjqQpgX95APjnOd8fEd8j1Ja8+GFt6vKQlIZPkqul0f45OJYkJdbt+ENf8BKjPfwRzkqRPqX5T
UQEDQ/lUFraZzz4g65LEMW1T4mU9sVFeEm0/E2VCMf3Hb6TUOkb+pdXMFUMgjmTUlyixF+LypVlB
sdfaPL9iLVjesf+DC3QWv0XEGEiF8hFLlqbVgiUv4udaovDZ/u6U1JvTn/MZrat1EunLBTf3oLLB
7ZaJF+LxXkd6flbg93kcShuPLBtXIaW5hI29kxNWydhMSiVaH/Phzfoe8oOomhIO1/NS2rzW6Hra
9kOOYRqiV5ItqQ4WWXRU71r+8uJPMDrNZZXgetTX4SraKR29bt3MoZD9ukBUUtAvQYauhlXxLUxk
GBH54D5OcfdNLUnRVBruP/l7yCG5N6W7yZo4peoXB+SpEy4CXVeBDcR86gw6ZWeo67+cWlX+cs6p
znqcoRX4USVvJfH1sVReRPoF+3TXmOPMMHxU7ckXY4Q+AJhrz+HpBYugbqn8G3kjRVZDrvqf2E7M
jjXJ7KOTbfwOQyHzd+uL02RxjYrLHe0HssYlRnbWb2O2guUBbsWsBKrfRBcAOARR/mxjrX6gvTPu
4u8bQNewnD1sBD4ArCEc6aGXCawzdLjAl84Bd98IkkaP3od1xmv8f+NwU8ins8jSWzffs2JQ+uB7
cbW0CuG6ioLoGqNsxznRsKL4BW3Xw05DrTmhGpFr/IQVx2IErx+Zt3oOvhdBIW46daKWWt+vHwvC
b81T+T592tF8l7/yR5caOGW3SGkH+JSHJ6voogZn2PGXAQkRw+/gNCC3ephuYqbRQpHioJAj5VPO
oggEsW4wvds0ghOms+kolpsVIZLpHvER/7OG0UioH3pT758lmw4DrZjs9PUYehXHpRGnXD6TceJ0
Y/JBbS5/d9uPo2rRHMPWBks+IrN7ALA5AXl2q27K6B8PlRxBrOZNvoRd0OAiYdddzl/DoLgIdbat
yL2nppWecPtWT34QK5+5zNEUrWmTWllnILtRzHhc8VSDTtK8hTWL1cxx73gxSD0EuF6r3dLsbz59
xv9T5jT8JXjkSwWpjIk4lUdoYZ+zkLfPvi7xuE9NMRvD261ygLU4FQhZDAmbGMvla8nSgNbzXGfz
mep9ENDNjUgzRlGARJpV69Row5RtcPs7KqIGH2xVQSVw1jzVHO0CiZwMX30roY5A1nPDR4AVNRUj
C8Mx44ziY92uZ/dUjrDMImVUIOETHdGgNk8bAX6Jbb6rLZl0nL7Cum3MmRXE4UWO15JHQC0Ykv+Y
WDiw1WrlvYNBF105ETsSdtJLwFIFpb/F4L48JzRKwx2EtE3UMXbmWZPWqsptmGVToNEMh6xiPrES
sREY5tl7LIimrX3ZmuIpLDuOq9ezSMEEtovHrbXO78UHQb1y7d0QN6ufawO7YvtaKZC4DkvLUQE9
u9E7lybtvaCZPv1QMlsNapW3lydnIDEHajCE9Lu12QRL6o9YaX5FIFFbB7ila5uQ5Rg+EICdvKCS
EN1CfN3YwV5rPB8QwWVGePzWL/qm4G1c+V/LVAu5XLrBbqoBaQGsITTvWIl/HyTGcvpdJjPV1Wc4
ROSo9KcIBC8k5lfoYJxDVvpejOMcSeishAcMpkhVUZGDYRIXdkBqFG5LxazzX1hjsPoDKxlNVCz3
hbf+F+yA5wnoZa5KxTcsIsyjkEk/XRNa/gwSj0jtOELUKHj/X6oBl6VdZwxFSHRH7oK/kpKrRgkk
+KqUEOLr7x0rUmMP7tSMzMkFQ1Ju+lsRlvp1gFLwjE/1qX92ciNB8JG6dO3QSLu3BoeURps68yjz
rrRgGywwo3JzXXrMY70cQltJm5VTIf9m6BPcOYkBPV6DdFPMJLA3CUm8roBGfm2DHgVzP5KoSJI6
7VfJizypJU4HXkK82p1Y9vVWcYVM+62f4yfDvQV6sCGTAANLL9HNPhadKYou9u8R+Fnaj4EtXqpT
L9euYKW8/gMdURfqHSZg3F/NnHFn/syLsbXpvWz1LsnxkgDwin6Rx3dJgnmxFd6lkDZL6jbQbzOU
fKuDfpMg5F6XTaqSXtyrmJboWc+zQ68WxdGJ6Bp40gRzCJoB4jDXME6o6TpyL2l3eDgpO8nnlpp5
h6SwhtDFM3sSwZZLtCkNQ5MHkqmrdX9bwnl8nEgHKnTP0rD4lMRc88kBEo7g3gwyLvoSoqmJ9TUl
MX70LufeHgwoXbsjJqcSBAONi/QrG1WRdng167j8fTyZPl14yzzTjchj29BsciatakMbHEx0ZpKn
WoB690X9teI2sH8PjjQxyx6nMNQ7ICzcvC+PFKoLIA9A8spei3TL3t15wIwMS35RAIzkABbm4KOZ
v5J7GzxgCqIw+7MyL+8vBtTxTzyPdvnVUOsGK4VCxcGtCWiFpPnxxEaj88h9RlziHMZSOaEjhpep
lLvKMHLuNhrwrr6+bauCJh4903OnRoQSCWpjB1fyhgeP0rF1kPYlO/FO2qR1Nyd0/BDKF94/TC0q
4NqxbA+5yVgsU5a7Lkg8/rV0nFH72+1rcjmMqnkX7MDlIH/URzR5wUMGVckuY8Dp93AQ+FmShAb3
VD/feXCZjc08PCp7AXs0tllCRVvZaWuOjzy5JJUq+Ece13L+9Cam4iwcXSSr7uuixSVhXSBVL6o2
9tJ/sPKX0T0ETA7Wo0QnMIt0auvDoQnzKBq0jK+3402BRJ39snQLbVU7HLthk3Lb45Qh0f/+3jkg
gTQLfev/e8HwUSNiVN9zvcZTvOEfblvOBpurABpBN7InIMHBJJ0xZt7ITqjybVqZ+zb498OdVU+F
hLSyV/yVP0TaVMbGpP3K0E2BFT014NibKhq/Ul1etJ/3evv9tj7PaKT6ERf1z2S53XhA/zkDoLdo
CZBL1gnzZ87NOY3IoJrqZ06FdVe9tSDkZczSTt87SAwGkMoqrYTDKHt8GjR25FBCldD6omgv1WBd
8PVkzsrP2d0Wx7p8FGsCZbyUD+zjibOo9iqW/N6koC3nHnMLQtAdSb8eDfcm3GtX+w+5sH5dowyN
LpyIdTrD1kP2o2BLLNv/ZtpLRtncqLdKzeVkO5CwLrqxGpOUabh4hpB96FrxExfh34pKG8gJ8GWg
a+qenTYhH1EK6dpptFYAwsRLGd0SbS68hDxO7mXJjCIa+EsAaEbYdNZmWrvFi2hyUFsKqF6ehYjn
N4eGWTD7SLjLqAtrKVNKsQzF93w8vr9ckGJjOEx8rDCGaHgkCtGnYBTgK31yiGf1roeDMML+QLSo
4JQEvUw2LcKsoPHSSzzFfc9gnyM5NIrj+YPqHG//GALxctmvtzGdd2XiY60uB/RH8UcTJIQrECED
1aFs/jP/rzfkyL/7vxaBhx/S9AYxcqL9Zoh1J8AsNgBMQ/Mdb/u+kwXEqWt9pFnZE3kBly6pxa3y
xevJOovEhC2Ncmmqfd9OePiXXYvGOYerW1GDH8q5TJ+yc7SFm2RTMx0ZRhVWaIDPaubkUPbpnUIn
H0AdxczjAPF0bODSOLCrA4xumjcsKL6xEyOKAW5ev6A3KogjIk0iG/quHh3oOuUESx5AqzS9LJBL
p6uG0+LXxsLMAwk2apu0JHAa2h7JqX5fMSoOwD9glz78v0usHBdMPLM5b6e3kCBLyzEuKk9Jigj1
CL2/us1Kd4KHMsNQRJQVm2IYlcXfkRPy6ZX6w7DjlJYtXL4086Pbc7B0bSsNNHn2HPAd+SfKl7FV
/gD9Z/wpM1BniUMsBPUAT3dco9KE0O5/5rT9xfL9N9KlRtwVoepvnSYwmcErttTsbkaUW75pwjH5
EnLIqlqG0DgMmWmoOltAWmW1IRT91/sXTZYiLW0USTGNgWC3GLwQzyzgu0CFA0RRKnD1GWwK3zRn
ksSjj96apP2/mIdaCtMpJLl98BN39pKrRX+H1uIbthlK8fPgVq+npOq5X66YMvQhTOrUm/9jzd4i
qymL9vjLzKG8hQTaxF1tg+o8qeQ6QdZG9pSrvxHEkE4yK7QqPUGPLKnZCdguG4eJleJXezeVZYdQ
hFLxT9bq9m0BLv8lTrKoZOYGrhedsplpShUTFlYPCw/TyptX5aXxWBjYEAUU1geW/YVuEE224dTu
RHpK4cDmPE4KA9au2nl6RKa6+BqEqLZ3X7/T4mdPEbvYgP3b7Hp9bGY8kGKSJwK/yQVEhUDiBpkh
vANOMoVFu3GNOz+BM9hUUFAkt8ZjWggbH1GM+S5rLvtAYaGTW+8Of0BjTEL2G2+D/BXsA6H8Jwf7
dSsdQ3WFHrt+R1JWEJHb06uhJXkHhZ2xM+Fj8JxhEFtVqy/4QIn+RwGc6tOUhmGsIVb4LelYmd44
1DBitwfqlBCn5yw+pB59VzrE0S64eAdUzA1GH/6FV5JfAOlyz8JF74pZrlH+qC7FqAFM3bRYks8m
tuQ7Tsv/wJGDHUuYuMdjOOnC309rHKPFlPvMxyXTloePmLQhI2phHNUEKrytbzu5+bJaXtzhquZA
0X2HI5Pm2suEUW7k78pnogv8KIvy7yamzOS4olQQpzMwV3C4ntNCP+aPoUuS6lNAbTKxSGrrnGmE
GMgTlvOxO9H+uf6oyy90eAJt49t0b8gslsf2h3gDAM3wY4xKO0h5Auz5Y2MEFJYpyr42owFHczr3
3kRa6YHCmYhatUsqUmxXh72g8rsxePuUJxmPr2hPLPbfPO/eb7GEjAtFaeiXp0sRBNQMWPXkmT1U
8o14+ioMrgMSiRHTzURBJrx+RNILh0DZysaKl+IdvSwfqAsZdqAAl5r6eINbUGk5LSbGKi5SXNrO
UlLpZEhX9G1GHPrfou+UN2utl4GYQsaMTwZcjgRnpXH/TQEdH+c67puKi2GFsHKq4IguIf/8iznu
fXVD/G+iCl7Hvl/FFYtI4H52zV4mNyOfzk3JDuWateNlgfbkoopSL3V3JL1Wj6J574D/jElOo0Yh
b0ksRnE92vx5+x68iWMtB1yEJsr5NNVloqLHJS7rb32oHFBE+hHJpbEKn84hcBdUnbBAF0FteKOV
Hss9WJyAoyAiX1b8xCnyvBKzhqxfPjksscJEGoIvgR4rSnLIkrdCVLHthcQl0I/BJ6+Q/5CGGSuQ
CA8Gz0fTwTfweMRtV+8cKEF/JdRriaFR0GJyqcXvRqzrxYKQHxjHHpu2XJKidkKLiRGcFmbrH5s0
43KcGCYTWrtYhb36O0tjvVd3ROQsXcBx+WNA8PDj2yhkm56S8CtPDE9EAOCtYdE+S7j23nazhEyI
sO5zgELniEUlMVdUbPumokLdDRKie+jF1Pl2tm5l/iKE1v7Ut0X9xryduZkwpTR1wR6fiz5GUnwk
d+SekI+zflojTLBqzcN6f0Tk972t35KdJneWZpxdx2cMiZPm+17fuw0GQT4g6ZcmSiACwDV5WB/E
1QsN37lrLOCZ2C9ovb3rvTPEGG+/rWH395hOY+O//1S4kVeNDTauzb1oBUoKmuX0TJKkCrAgaqvJ
y+V3dStwyvywnD2/Zkao8OWkGNRqZQQPegEY4HDpuC0iOOsIzZC8Ou6TCeWYqmTgQVf1bfq//Ktm
dIScUKywlOi5M1MOj08s/SaVFUrj8V2fOtAEMeYteKTdqkjw8u4xbfs1Xl4M0zK6+p4hRyoZBu9i
ht5M5l4b7ru0uf56DyU/WZduWW9J2pwasyxk8T/9nGfvS9XaENceJXMeuf1hfY5DOrsKtTY61cYd
k9YERt0IU6kZQSfdFaMqPnVNfzqKouLao5WkW9cmzGYK0WEPocsnZ3DL+vPEH8jQoBzGs/ppqitW
wzuyn6DupomEMC7HxitWfdHl5CK1/ojK+rGPsPKPE1/UVuMsdtGTbYOGNXjhP2QaarliP3sqI8Ps
7Oj5sSN84HN2aqTZHlExX0G/oAACajeEPi2AZaKHGUdh6Rxy0PBbYKyb+YOIni9kDnRuXQznQzm/
Zivygi94HkcOAyUqq1p75C8qHrMOU30aG8i0FLS1Wx3U9rUzsVGKGTGkh4msPoT4m2APCM6QE9k9
xBoxQ1/7QvpPc5jJyOA7pzTIMfHavN7aTP48B1SOWNtT5tUf/V/YtHldJ0A26axrwWYdvYa25QDd
jd/+WcG+Wf9VDyPPe39tKn2Vy+er9q/lfxucEPmgL8TinACGQr4qj+Je2cTBbgBlqx22So9Rc0yw
1eRkCUxouz0FrzcIEX5vvGXqAnALrO6wDWHtbm95RAz8cHUlFfDZE9qzv3HC9jOVAy3489mcloqf
yn3GizqsIyNNpxgDp4+xzRp9BhE0NwYBw43E/dq3KV+N+U6SOxD86AVMCrjFDIYJBUjDPHBewsBA
LRvgGtVBl6w0NQ7/412aqFHgNe4Nq/uO7t0+EtAFEKW8LL166/fo+ajm1EGc2b+GcgLiJgjzVYCw
N/jNbTonAdKj3eVZ+Yq0MrKoNq6wVbAEI/jFrqM9MNiFnhjtV9070p9AdZifWDRxTUzzwHMGEa0K
yuXLHK7WS5/fe5WH8GMmZuo+Y+/9Yuo2GrblutOhyDuVs43oa0TsJT+VnjAMDHaZ3c8dAf1WPlx6
Zq+dyV1iF/g2BwhKnqK2eYxVntRHYg2/8s/bX/p7em4ySd6n+D8qMH/ygTs6U7F5hYJ7H20dtyJT
0prjuJrsHFifePpJLLP0ttZQnG8Dz4D7X5d4F+DDLEumRLaWOyUJyblbdRZOmUQN6E/Xn4aIJXK3
T38kzBhSuZBvTYjDdmSNUcQ+OtT8IUGUQ/9+eviqKSIq7n4RFEVVasYKquDKUk4FjMCeZ0GUMtf/
sPvY4dP5MA+kdLNc0/0I81ZAiWb/+PY6L3/Afw4Ioqfnax4inZoGL0/x24Fk+KOwm3vDB2cAS29Z
DFrv7pNDw3L7tX1ODQNLfjFwIlnlkCp3S4wvKQ4Z4Q9Gq46iK+Lhd/0t1aAHZrVQaLVm/6SlVBej
yGVoYhsbzLps0HdBFeloPln1ihFdrTWEjrYdgJMHalgmGrAoHG8GBMM0YQsnAWD8SuRvFGfH6ISb
PHAiiqYLKeBAkVSIexsidCVVGNcoG3VYq7FohV7uU5ANsRJFqZHHMIcElG+s4vi+zDWpaOmsHoeE
hTTHuNIxqA+Ii7t19uyUvC8O/rCenNamiGlq2CiMsEIP5thfIpEjTDO8Qjv/KDof05Ur7DUcunnW
wzVTGrbEUH47kWvW+2yr2gC0HwUrzK/DUdxBqov0LKLA4iejdteXs+fWHNQH9Hp7vqgu29tDplZt
qnol0GH83LH+Jm1X5EVQQbYNLvgFMuymRG9uLoY5Gli5RasYIcVoQGy1PbrPL6Tg1W7OtZjUlKXs
gCaV/3XxqIGDYzR6mBknWy81ET7drRnSDSsXTV1gKuuOqkfcy+O/bwMDZ6JFU+VTh1/WK7Z6gm39
fdZBr/so2aBV+6q3MGSbyZAzrCG3FaDcMevsQ8qHTttMMt5Jmw0wbEOiON0WK5ubORGkmqul03MB
pCZq+a0MrVKHarfozZ/6oXKIe14yBzNm9nCg71+bOkqSz3TX0Xm82yRy5tFMtpbLluPL0ZPDJvEA
dCm2NfS63UViG5zgf64D6lHUIHUwi8BgSFVvDoBxko98nhkCR+OHmv6TCjzfjvTaqfZ28OW+7Myl
3yipfira6ntHJsafUY7ZRPQcGaus6iR+yl+SKq4pD1/ZU9PaDfe132Zk8PeHY3wo/AcbguEnuwoD
I41WA49fjfHn7+iU55FNdTI41e7+LUd2Y9ec7ea0rf2uJY4hbx5TcrhKZCzY0dWQB02zra9Xx9f/
UnhV/6VoJyBwG3q0On0psgTh1NhuzOuGqjLpS9J9jSiRvH0paF5pxmnWwjpo82FGuZBKlN9L2R7P
TYG2JaERZHdMVXQ8d7T0RcJI3KkFHOQlIBsMe54ykYoDHZMnmvkoD/BMNoz/oUyVd1Aaljb7/dCI
cfZe/NNGz/icU5YWpaBlg3T+zpDjQpZ1G3YYO64EzrIScz+4BOVdbYoAJaIlELJ0qoWrUMVCq7T7
4TfY8deRyTfkGOq42UvoQM3wpKxu0PtxUddismu409/i0tgURMFM0y+EX3eyvXgIkGLjeeqGIHY6
9qqaIXpfRWy3rIc1DV6LKJlNdIWdODpa5UDht63togiF0eHRc3d+Uly8UPOPzxESzwFIkfNKFcbt
530vwz0ziJg8gI+0MaWwe3j3k/qhPn6eSPzU0l4DIGV4R/DP3NvJ0S9jvxghAWIuQPHoinEXX/OH
cnkhS/m/IBUarGfoSBW+70rl/MxoGI4kEi0KgizKIXKUWyyMHOFv994dNDrXIGW54XlPMh5j8NOe
zAiMEIUVAqu7NDJ+vsbf5agwO8XJ7gVK73pz652o1G42yfHqw0o47i6tSTNb/Vc4ko4LtdCRLXoJ
Q/hsOOhi/6GVPD//EB5iU0B4n/J0Nj8ajI3sParn2BOHFPgLGon7C/FE4qCJ3n9Db8kLes6+ihJZ
/9Ov1D2LwCu1/M9J1J+QmK5/0lHwDOlZUxAIyVlcAZGeKqjHRhMZa+BwOJxii/OQCnhSKZkXmi4I
OHNQk+v6SCoOM0JHYk/Y66d9d7t9b/0e3xjRm0nBnrdsREdxHlkM01EvuT4Yv0YxyQoWsNBNO3ac
ED1s1u7j8nvyldj/0QpfymUH0q7T7t3BhPZxbiA0vApDCP6n7HrOwG8YPdY+ephnUVIvck3y5roE
f/B35KIIeKij3sXmdrNLyd/Z5h3BFP47RLQ5O/iccl7PYLeLPf4gUl8T4R5WIfKDq6FiA/5vBcde
lCupFnQi8nQspkSv7eH2ATeDMENRRMtUVzv/pZxSxN/DCgOD9qAoODn3LqROIq37Y9c7OjHvhewr
X8sUtCPEnl3W0xUOUWVn0EhWpLvElsOkwLvvNk+9o8pCruzLASTwdx/FJRLBoFEvJWwAL2sMvcVq
/oT3SWvoi5U/XHoKdHJ4Myzb3mL2EK0XvxtvT4JmVAvth2BsWNLdXu/qHBx9MwvjYH4IooF5UwzJ
cD+ojOnp5d9Qen4L6Pqhbnu64dufLE2scpzl7AzLdIh7pjdh1q75OViE0p94c1ekUIxxRRwTBuu4
OMfTA77+k0KUV+Yth4xWOGEwIwewRadfT64ZFMSFrIAiKI+bozYeZY1Dt+J4P3Wb7I3RRaeZE3/Q
BSpi9klXGjPyOetv3v1Olug/mvtVkKn8unqqTJBSsnkzX6VS5YSmrKOU8HVDBiDc4X3JYCP5HDBw
tesbeUrnj741rHofulMsDpk0fgSGrLTgGV5z9C1u69MihN7Drg27h6Z26M7CFNmyN4UD0CKcJe4d
Gy/kIpiGoFQkLxI4HJvKbZk3sRboA5SAqlq3E6Ll3HTJC2asTqApbCwaVEpuBppMmhnwmhLnfPFO
KFrKPuY+x+MTUvQLo9/uL6f5LXNP25EpGaN+lLI7Vob2iDDI8YYs90a0+HNcTiEQFJ/UDt3FwirB
2n+U8s9voD3uqvHtO14XjVzdMPyBZTGHL65EKb4hHtEIIOUehxUA2/knN8f8xIgeS4ncvoX1aimQ
YSrIpovSE4hTkhC43VNmvJdbWqsbTNKdHqJGdLTHkBo+dCPiapdzdvcAZseUuUT0Po9CNVBmEh8V
9nk5tRlrtnWDOpAw6ejLvIGkhlUsJ5c2YDDAQR6Mbu7C7Pu4mp46OtMUwTs/NeaKgdF6oyIHFbMf
RbYi4oUTBF7UTwTJCuyU4gTSDv60N7vOg4SDlJWG1PUQvT9Vdw1QA0CUm3SSvSV5+NYnvkJKOSXN
/nFVjiWfdCnge4u5UEpcZIUdKqlx7l1Gp78jI6g7rFXW9WefuuT89w7eOci6yLCwRa/yzfv/FL7g
18sChVYFsD/0Xu5wDC2NBQLzhFhqfyJ3geOeX1I178N1gFXp0/tlQ7ZoLC+dCgmo9ixHokNQopr8
8F7xm8M7JdKwS+lFnO0crBVM4DA3k3SMflceCtQm3S8GjwLqmnPkZXMHI2HNkPZr8EXbC7AyKUOx
DYb6ZsZt736q843akDcAx/hres1PNHODQ1jrxJyZ8r4FakRf9N8UJgagG3YkADaul7CCqaijgd4t
29lrRChVUEF8oXlp/rpLEBHVCo3UJ+kP+rmJx4S9zZZQysIvEZxw/k5aWRsArmN4JkQrYr0Ik4em
g0Oip0tfLGCYMoa911CkgobccFpj7mspzIU7xBf6LPfaqiDW60tsR+4xV19mkbStZ4sT5wgKcQHP
VUtLXQYXr8uKlkxpdE2ylX1i3x8LP1DI1kFoS4nDAw4DCQ3LvI3AaxodstKz8R99EcGmtH9sfKi+
6Xky8XA7l7etTC/Mf+BuXRQFwRES9mquyk1GuSlKTYS3gr58o0IhVmBafXLO6VapTShjHmv5lQz/
z3iL60SSHQMOJIb9kUJUutvtdNbGzjAg66TOvHqxzZeMwVINQq2332NOrp78Slk0Jw1V7xbU4Z1J
gToesXXkV3hE7OE+QMacQAg7ZZIekwr0aInqvhxUP7SzJxykgVB/0O1jDPHOyCYWS8xVSFUFJ/B0
M8EhsOxTaE/dwHoBC5oEDXw8pVCVlDMMbuS6mhnkXLqUSivXo8Adrdz+J6II2gTuMPFOl1lb5xWo
yMRQDQ9bFqr8G9BreZsmcfE4R/BYmmzfJuzSTiY0x24vkTVGJw3Bhz28ji6pnfTwHeodtjmXB8lc
6tgx74Kcbp1UHha5XXXSORQx6NKz3rnmla8NMpuQlSqzNvVJXocfannoGz2PQdVNiOdJ3usBpKFO
bkKNMJ6nMHrSau285a8ODw+H6G0kXksyWB7lnh34fLKazB95ig8CA6htnD9R5iJfuTfJ7bCJ/6Yv
DZmxwGlDUW/9MMABY3IjRCqxjdXsU5bfAjZwgLj+IvmcyJ7kE/VFVTJt5jzftDtNnKS7ZkP4rLMp
ADO1GHY4len43x7dEX8txA9BDXyp9ASbDz/A03I7U4ctDSJmDd3mo8rwJi+4xcob1KJgUL00lcWy
qo6zw2S4Rooez1ZFLmdaVSpsGj9pkOKTZloc4jaKrdX8lKRlgHL80oQRVJU0hifkrTYYJZATnKsT
KiDF5xjdUA68QpGTZ1oPYv5kX2TiM/4dj7rSmZ53PSuIMpdJA4epndDGEbCxcdzBRBufR7NZOH26
vEuccVlOqS0x1w4lrudZ+oHtTT6zGQXxWOkmB6pLKJeQCi/nhlutOwA6qaB25DwpQHWFVh81oQio
jVEbaGvaCiJ8KvaoHtFYT0OwFgKgtxigqJR0nJmMkinG0fkCGxvN36nw/vN6MGf0TOnyjrpavgV+
xkmi6CQD66x03DU668nGXOdN7MvvGgGmn/539qgoK+Yz2rIi/iIjhPD+qhPRBOTJZYhHKEm6RNwy
19+NwDeb2KIb2H/yp1PpCuSaucNUVGJ30LCd/baF3Sm7GTICz6MGK1LdfNjSwQFVGU7HJ0MLnOJR
PaRx4QDEJEEqjTfzLh1aiEBImu5Rsys85G4UA2hUPDyO4HNyYxzlcWBwUSWnGBHDExhZ5hSUIU8H
D8Rgvll993YYJxIWgpNvY4UR29GCWCj3EFu4OEBlKjXY3AIDe36iKtIeBdzrdlI+4l2BKSQlxrVU
MvBcfBabpAe8MoxJjh0AK19MCLx8sz6Slp7PGmWzWJaGpxHME3wYjePdBMkTTvekVIoWFQKlUCDk
PuA7sFDs1LRUFOwaF6hxaKEoqloJ2Gys8g6Q8gK9djss9Isx4ozYpOArfxK30uXTKd95fJIRqzp0
puBKhQvW1V0k9gzldp49ag/U+0FPnWzxZOeIEafk4txeM5uMxZeiJVZNWHybqm0JibTeymGoHuca
RZ7WAHGv6zet8mX3JR7Bu86r2q5jHe5k0TbD7mO53m5iECJmRaoqr8wpHrG3ua4OUq26X+Y+U8RH
4L/zPAvlnA/qNncHnZFXjsldXrPzCphKZ61Fb5bz1oHU0srETImy7ldas2wiQrtoipa+Ct10Yfzc
prUcheLC3ghLl9jmEXtMPGMwznyF8qdO1o62ryc1ZnDQ4ds7sbQJdtqfbXLUw1CV98FR74jK8kti
9bO6Q6Fy5P8WouNoUPLPiZK1myPZubelSesXrB9o1xgOHH2xFH99YgpvuSgAB5vzGeyVtayF8a/Z
jow0riVRW7cY9PJLSFJ3nPkEaF6fqRluljJFHatPw83jZ1kHhRUu+G8BDDMCPhJXhGIEpsEJ+UOf
zLre5yFFU1CsE9TL2X+FylYOj2UkY0QnORAW64V5RKuFsbBzq1mYPBSjUg/yC+oxrLz0sJST8Bwz
A/50QDCiZrOJtgOYwQw+xGD98Njn/3gYZYVJ4sacuk0VPDLi++0LhPX8FLpcfvtly5Vz1809I+Tf
6spgSX6RZnnzmG7M9S1JrAl+XeLRx2C7xKN0jIiXXpoaW9lRQsCK+3T3Y7IGQhHLvl11TrBUSxwa
F+yX07SFE9t9oeTW0LPsLD2GXQKNxpSZx4BssKX5jVVZKBDMk5CnnGK0ODBNmyEHe7E36+e1Orhf
vLvOTucpYKH1nOVeW0b8rGSyxPiF5huX2Of+O/ZFzQYtUpQHIj1IX4iVx1VCd9EFoMbSynyIcXYW
/bPPgZScbi8ByXAJCQWWldwt9Ni0ZzjZr3qvjrzGD9aB69sKP4FWW11mYeGIBzoXrpQCFr4jEpp4
uYZGi/KM8rHl5GySOMCTZuxg3Ga2v5pOnFMxcRzckvmnIwoX40sQy/yk6AWpVglrkjDVw84b59xS
8XXW3wAOQzZpui21wBiMaSvJeVak57if3XT5sQAfn4nRzrXf79BwkryGxTs33+3IS55YeSIJczA9
3a1yOMeqNPHuohiowMNxM2/qpp8cZP6FURaovgNLMVu1Pd0PP9gehJruNsQLIiWmDtrUESZvJL92
Qykk8jV8NmqVZ2ex+t17bLeYomlySgorhhzv+Iffp5KEkzvqyBlZh2uI9zY+jgIoUX9wdHOYeIqf
37/tr34/uxMzcAW05sqic5Nj08wGfmAaMgGHy3jBTv1mZdcIdOOw9y193i1Vfc4lW4OidBSmCF+U
1yf/xrSJaselZj1qZEfm/8XDIIDtoWZl12DEl9wyU2BrOeWd2r8H921/v4kHU5wCX/TwZhhfe0rs
nWZ+KAXwa/b9OvaXzNH24ZTAJdlEK8sQ16HyU0gOhfi3rsUKdfxS1ceVgjUlrxGFHvw4YMpKx6PY
b9BU9PUrOVfRL2e3awlv1DOcYEWr45/LQBeh5j0/QR20bOBcu+lOiD0EymlleJkjzOr/EjCW35gu
zMbTxGGi47yq5a+KTmLJkKxcCMIdjX/Ei0csWpw3x0Nxa/vlSOu2SGW9rEd3c4Ha6xX4cMIQHwE1
2jRILK3snB09N2m+BHj5bQlVecR5NEocL0HL6ejaF+ptQDwkJsGl0JGmMO6QlXqjXNZFNU8P5xhA
lTlTjb5MB8YBasG8bdDBShbADiSE1el9y+B6l4OUR4yjJyiceYC4yQo/hcIGBwTkixxL8MN7mtb9
RoVkdLIQYu9W6GmZG3hYQDMe9vF2tFpTmVkZbZu1Pez7mZpOOAi6AN+5wC997AvvjRHvpwXAg8eQ
HH8Zzh074rZrSy6pOtdyG1IS1VWcv6XS8mxBJs9D5ul1BrBrbDx9e+7WhDqJg4LjpyS9J5YKdP+t
IHBtdgh2kXEquQ1COqYSAytT/RP963VcY+ztyr12Bl2HSOsP737BwaOOc5NYkf1BfwzCCKIgqT/B
+3xj7oIEUhtfa1JpoY3P5zZmGZfsJZ/i3H5n83IxqzmYdwcgOk2y88g0jtbrmbA8RrlIssl//zrP
xdAtU/pwKheiaZKATHK6N1N0/SIQOd86C71SwhQHG4v9tTcwUiR4SyI4aBzccJaAEmzvOxjWjm1a
/Zo/d8eLFTYf9qhs7GXUZn4od2IrOSoiFivmwy38m7fBZAIXnxsJwM52AIo7o6Gz3IR2JJL155lW
YGEM48FoJsvJYBMwS08vBTjk5P9+xP8xFpBp05osC/jt8flTH/oFOGTVwtB2LMnqHgwOq9qOwkeS
hLHccbm3k3eDnIQE4SWSgCfRLy4APNVols8sbdpW2TsMmmhcMSQ/69/oWhaKm0QsNxIljhYt62yI
62own8LRVhPtZAFQ05kac+FaX6zeRDPXreEPKsX/6qpHNU6Q/hXMpvMQ9zmKgq8lVDMays1GlJqX
XECf/06uHlMmwG60iWYbZuYwd/9lAsTTebnKDu+djBqzDFiZMRDPElwspPTA8tiapgxwR4oks0BS
iwbak5s4pzAocnHS0+pWYxieI0ftH+LkAMUgaV8AMoRXJc+rZmczJr0F39wcYQHVsoAAE3RUDACc
pyAo12cSdZrk8we8dbHVXlp5QCrUOEQJnLQrUZJd4aHhIAa/yavl2biaBgtwKmDGt8D61ms3x/RZ
xOjzYhe0GVZsv96ylvbkTYFjxEImOWSJ3g9MelgQgI0kditPzTQ4nc6scR5xE3RSG9ovrgLxqlYw
Se9wU5A6LFnhpOGqsa5XVxm/nzW1gRlFJcS44+uRwmiq5fNftOmjUkXSZ15J8czldghPf/tXhj33
uez83dXstetJmOpm/IJMbPGfr7UayltSSM9hsxv0jlAqsHiMXD/XLJHLcMEDPgDKycrioc6nk6eO
l4tCZE2EmDL82CAg5CvsfMBiJ9mOOQhfdjaZTC/9x9H+psDFtXzsYugLF2a6+CKVnWXh//146sgt
HDOoPQkt6ue70wuScp1Lh+Tz0KlN3xr9ZoKbtO5m18DMma2kjEguVuMTZuXmMuBlD5vRTRZdsyWo
HPdrFDnc5yzuJUShCEIgRUOtglAmPudOdzSjl3iOEYLxoK5PehDjkmU2HNqOal4iJe9ve2rsrPl4
uSDhxTgigffOIVGdlDRrAjr45Xn2JRw7mdAM2QOfuJiFzkzTE1aM3Mf6iAOGhBRzMH3VjkS/DlCR
myomQoM+BNv6WYADcNLKT2N151Ll6Y/9xBMmiozbGp1CQzPV5/zwUx9yQRxVUSGyaj93ZQsb3pD1
FXlSHLz1Sk0klE20o+I5U+93diOoYgBG4mPt/9RP7xPDxoqaeW3+D3J68R0Ycs3XmpzfRUdg8apO
oLXt0EK9c0+TZBBtk7g3aKvDrSIr1yLhOeyFJC14Qaq9yfmQh07JkTJMFlo9SSxlxE46RvJo8vLM
pLWzWaFrkCuRDSBRx2KuEYKqkDRHGNhZ/cFVRG2syqdZ7OtvZ1beX7uAVocIqAiCiDibdC/8chOC
m7GDD5cCcGblMMREPkrJ0RLB6gq5cgEW2jKlqQJ3iqv+X1zeVqDGGBugVdj5sHQ0QV4kJ6egtR5C
fSdbwEuIzM67ijtYs4OK5J33EPqLCowrDmA/30baTGfOGQOGxC5pErUBtTQXjclWUjYKkf3MHB1o
oDczm62+BwfZyg5JDpXK4Udnk4xXNmCFfjX4mIyk1/yhLumG7ZjOxwoNPhwZnnJpEy6e9a64icw/
2NCzpfrizj4jaR7IHQM0I6fMeUFnvMGSLFkEaY+K3DjVn3IF98sDuBoIANNu/Yr8KuHL7VWksGPf
/lPbFrFCGT50589rGBqU1YCxBP3OazkCVygVZAlOgAi50XggtkDxyjGaY+2csGeP+c791kU9C3sE
M+j2K2SO5b8kqxPHU3tktIPJ6z82rli0CiodgUc7MsYUAptQ3iCpd06tjM7F6NjhprbdJMA1PJw5
/i/Cppq35Ku62eeEICAjB0nCE0aV5JzOqxQK8086J4bd/q8RkrXZxj39iTV4nETEeg6WtOmBqdTe
LhYApvKSMQmJts44JaPOtyek8kPmVcpj5VsgNUxJdHoSIK45LE8iXavvuSlVaqRd2joYtEM+7s7g
NlPiXnPt+T5ppKHDFvqVVuqicGRysEaenepAyssHuDHTv/MOM1H367knDDLC8kuNx7fjOS/NleHG
Q1buJ7G7KCMc7m7CnAtnolYZOw+YYcSEaNOPtoe3WapBmxnDncKGxeraZy3muljkiUnxmAHrTOji
eE688gwtwZGtmGbeSf8Gag4ytro/m+Q1zmJ7dceAN2iVHqaIJZxoVgGxHK2gfFwqqcvhnMoa3d0b
7k0OepNZ8fH9C/HhzzKtk1LUirdvqrAul+WnSlWTVrlfIdUEFuck3fmy+1ZtAlTj2MEtqTZEkkcG
//KiIc8Vr6jO6SwBJlLJQosnTlzr5w+jnENjHkCDg0YE4Tggf7ayB8E4NstZeLYeaaG/7RXV31Ct
8SBD4U/jb82fEN7TqkqhCWu1w4CayRlbbg3qQdGWgZM1Gw4QmAk//zo+JoYtOUhE+8bAt8BoFg2b
gBui/cRO0IXENLgwqUcQ1AEJ9jIAtWWTSkYOSQ3+g7Gr9Fs91UKWWR5WfpFdRz9aiUDeWu8Vpr2P
D9dgqTD6q74uhxAURTLVYOwkgUy3o0Ccw2tLDY40vPR74Yb9Lr4aMfDYwQLDMD3ypEuDFcQ0qZxx
1ZV5VrKdH/LTe9STMBk/2b4xNbMGt22BGt+1NxrKHlSeQ3xv+vA78HSEUVkvexuO0y+vtlGBBbB6
rp6PafuvsSgwHw8dG6qeu78XACNyZ6dqln0F6WghhlgTbmd7NRAVqKrhcPNO07Unm54Z7Nid6wtb
yrkv6i5eDTchPPKAqJnKYjXCz7VRVNxZfHdpynsN3lWhnopVqzTXaHAM6KGtWuPlvzH5i4aY0hvV
aUFxYxxnxZTfDmzuuBj2eHGWyd5ooyPwv2OT3pHuA8iJ9TsCYz/Nugq192ZMlmtR6hrMrJcrv/ZI
7W6FNNio77jRSITuuGV7I7jvgPS7rfeA03QCEJ4NISoFvvh2UADI0nNUtENCqvr0DPq5NfE5kPM+
u7TGvKv9YmPQW9aD6sZ3GbWiqGyZpojPI02aGpKFabd1XoxzeO1hrIMaKxAN9pd3JE7jTti6/BxE
cXXLCgEiIhN521szq+69tg9ePsVYXWVeodLmWSZ6oilTE+LVKFaxn4+2wQgGxLBbOCcRoPYe3EG1
y6o2W3TZt8yiG7SE/C3l+hT/hMhEZnAbiVjbdr6M4ljOrLvjv3e7CExtSyjKQOcMdzdWuYRkg3xB
9NEZ5/yC0SUd+wJhYMtN1BrehQpm06lbIxpg4q7NYuyVEUyKaTEGJECZF22u3U4TKcL3Dna7a4SK
vMMjIK053lfU39tz+MonwZ9COSSH0W6r8F+5eqwco97f3koJF4CsaY+CxUh3qkuz2kZTO3UClB5j
PmgudHUzC1AzUZaso9oNckI5ShV3KZxzyo87b06MWI/t5maEWFfNhcgmtPXvfigDmyvFR4auzX8q
APlFuhs3WJQfzU77dG0PIaGl6MQzq6JpDvfmg9nHzoVo2lSjaEGqt0dSZ0ypmF/S8+ciSPQaPbvS
pa9v7Vw46zmAbOAfhP/J42QAacD4xmAfJyImT3UhJfcgnOt9ZC8JgRMKE77AX/myWa9ySzFuisXa
FrsH/7Usc8qqEJOU+PNPBuQGcVNzEVEifJM30BRISLV9q1WiQWYLq4X9IyIZB4sKROL2NBxVtluo
3DLBGM9lcBJw+y8kdCt52L2BhFH7yuNuuFMgBjceGz+qOaEWAZIMD9z1BxjSlp+3ALLem2fceYwN
znpFg35DjPCIYj+Pvwnpwth1fDV6dLDJEnGKmDAIXdVrguvf87rKe8lKHjJKGU68Dc5fhBcAdpla
v2hzBzadb2Wylt9CvI6n3U7qSmBv4h8Fx+y2cuUHulIohMFbt5iQpJ/rOqkdAwi7SbVdax8ioHs4
6FPGv/YorC+pP+4tsJwjG2M7F/6AqWS2Jw3vbRd0WeQnPtkSbeKo2X/PvEpH8/WyyjCnFmxa1VZP
j8/2Jpy9TMsyoteTjqyP9Mf1bkR0d/Z1pOEJ1HyO+d9iW1Hn9kv58OnoJeitONcAJCpXMH3dhGFB
5RnriBIpSEB3R8LfCV5APT20CZXLnM86jwccabdYl0P2XHqSAmBPZUmYPokyAWSkAcWXxN2Af6L/
Jsb5CV2ixcKK3BrIAdgxN23YpLnDldTfr7OwOB3szF2gyCtOqU0meK6UpNAy/ZmADcJ30fchUIav
vSvckMHmwRUejC/rQOOAsP5Eh/yOYGdWNRptOXiubp3XEBHpy7j2oEgDned/wl3zuyakwvGumQHJ
t5PgvC60yTeGP1RokzUVba4OSEoOmoIqTZdkO4Lq3H6I0DpDzM4CamiMYmHCNytKngr01pnOHdLd
10fQvvSsZGlw+y+u7EagQJUnjrDB1WFZARQM9rzhr6H+uautqTVmEM/TvuNiobIjSOUgUN/9KlL5
SxMGnVqggwiT/SGB48BW3786qRVZpAA5Yjh5yanSu6MlWCbIOLc3YLrmiuFsFRJaZH7yPh3MMAEl
NWZXOC/qEcadx/DOrgHxMtctHBPutxfyAvNv76i8890PG2+djJdtdc9gZULQbEQDhNoaFSfRXVyx
AN9Y3zqH/hX00ukrqg9e3ud8evXWKTslxDUnD8LiPnQlmRZ89+rHUES8VuwNqaS89OJbYuy++U3V
5r/Cz8HO8YDq/ixdzt5RhAk96+91Dk89W2fM+aovmh9nRiT04UEYqQA1Lk54jAtp4yyzFZWsCVaJ
H2p37lBC9H5/zY0f7qFUEKQnydanzcEtoXRz2+cj0NB7FtwlDaGSonBhktvo0MQGHq5jZrpJ5dPs
I+hIFRXXNPS4FabdJmsM9UdTc5YKuWimxS3Nkr96NgftGM/2SPX9IxvntVYc+NiTlfi1ORAqaNS1
mO26nr9yBZwKJlmavGNcCScgwYD0MkjwssGuDzovEwaVoa3Tkw6ZEsF9nlaj33R8A7v12o4hj0nh
4puvq1s95Vy3kJcGD7NK+p0vIMnM+t7o6J4mOGq7XRoqOc8I4wAsoamqElO/mKq2s127BM7fKB4R
J7i0jX3f4HoJ2falNAg0l25Gxe4Q+6OJpE+mtWhW0lUbpoCoMoI/rOnWd0F2QOlRWv1JjVR1YuTc
jWOFgpHw/UeRgGU/67tnY/d5ZMlZSQN/fu6G8U2vY55HdXrBwl0CpIQ5BufFTfWf2BAuyfvoM199
feG0l5XvWyP7SY2wbIe957OI6i61QCcaFH+kAJiTTxAulk43BCEYmPPkIybi9kHgGg96Diyjwo/U
BjUEOBAmmAcCE6q9DkYHmvM/IVLDu07NXxofMBt+D3cN0VSn/E/Tusqk2h+RYYTrxuTaHx5vXkjx
dw0Jq1YS1xjxkmy06cUsh4Fj/741LRdSYktz2hA5kgbGKrzN9aeKNdt6sw5OnoMpJi7ItjnCzwqm
diVKMVerwpzGFD3nLmfIiYWuknfPeRCw3d0gQQ16pBpDbd2KxGb5GcfcsjInH5WHrdMl0lV7SXR+
3XyWf7cmwpsHNEhkzdO2XECK8OIUNXMS9YQK06aO7AEE8563QcZI1fPe6cjj7PtPJ1WKiNe0ItdX
uo4algRrFK7LvQqIiWelGT/8DeJ/fpOGLOZnRLrxIeqEKKEPBA4raXaa8qhWlIYbiDSZGkJnDndB
FpFu9Oqfzm4dv5y2Ykn+4IaZ2UVBbZ3f1fgOQSxqYU7AQy/WBk+O34kvpjhtEs36EitaiFiA3wHG
d9p271kZ1+dkrUwG+5D9yx346iPcfg3mqjvesBwh0nXX0niVevffZY2e/zQbNwXpTixJQtopWp0V
SW9+F0+hFsmJNOWFhrP2VMOKi1cqiyv0AXm+rYmzV818+0hXVbOnleTffb+1YCxC4cpdPH78+SdF
A5DcI0wri75IXxlhtayiwNMoXHzK3HBAdVllUu04Y5B01dvC+gK9lq3g8tnA+QdD/MOcedWoPkzm
/n1HcAgYYXkJCFV0hKHbt0romFbKzSpLWB9nbNCeV60bRbJ9/Q55f1zzL7Vf75I37bItMMe6gmqd
3AsQQbk0AhrcCCkPyN0gB0pJoDg1t8PiwXvOBb1P/WJpf93U+bwLwfb4atItyA7aq+UpGtYBGR05
En0HXX3rXF+qVyfG15OkWpmkXtMda9LqkyvBlLmzzp+VWHwg2kTXP5zCle8ADcure7T/VETFcfbh
S/bd8U3wXhQj1xzYX5MmUtADUWUxEaZxt1qHDdpDuDlQmYv4umzzIoB2OpkSrCrhDx9GlnsDypbI
gsJ0wutoDeHOXiT2AkR7PA4OZvHHCvhJm3Q9GyMeSpOhuJ1DY4SNgYwuYWimXyTxyPF1UURHTI9X
Z6z9H6Vl3pdLkPcluuH1Qv+nWkMHWKSvI/v3f1vK2Z/dj/0gwpcrgukZ+Duft+g3+totgTqVO00E
D6oJzLejGndosJmw7KqxpeuTeX4D5sVvLy7eBGLOwtCacoDghxpqTWG2Lx1vY1iTeg7hrZ39nIXk
Yr1D6tm+FiDATQ7GwLcuZvv9XEjgeC7Rl02QNfeWZ/Xj673bgGyJ289viMmSL6tnY3tdf8WhV1zs
JOVWPJyFZ1pg7DzlF9cU87OLohjbijNOubLjDX1D0SovFNKgZ5WKsDF9XcNV8imA6baiGI2lTra/
dHuB5WWpTeanqzqADe3p4HAkgnrQAcM3wgnyHemwAR9NFFGjjv4L8YzyH3EgiMiUm7F0CUwwFThg
cXygVkXKZEgRSrzeGn4R9/sXRn0Pq/ccsc5fwu6GpAODVM4fagtUr7s73UCsaekhWll6K2MUMdGh
eJayt7lR9spZCTDFGhKGb9fOU2RZpGyMi2yx0PXixQpxggV9laCZGBPekqjUOk7GYoreG1F2Euna
OVS6SudE3DBs1yocufWWtdj5vjJ5MIUBxkdurVcdOW3ZSMGD1yQ/HwtLy811cd/0UlkRTEtu6XlB
YB5/MnB0t1XRCwXjHBd2EnSC/elRzb/JJtFR/dhw6LKW+cG3bbJIkOnHVwI4/RdIIzzRF41R3UnB
1GLTiuVkklQxIAPLWAZdHV1uvjQWbxB90ZQWwEwFP6Nl77BMSYqeDWdUX0zCCorahwOgVvo7dMsp
9OtmgtLoQz9JLz7xQlVuM6gEsa9vFg+9Qhu/eVVwSH/KL0RaqYOBelS2bhZUhdcszV8fN8OM6lIQ
6QxMjhm1ulpDJrNd0Ny6dXyBPnJl/6ob6qc+syK3eekq/kH5xwJwMWu24ljqAZUJYIx5Xz49yQor
1OFqsNIk6Z9ATvZilDyvz4Mh/0B9LZ38pGpkqIsCaB0moN7FtxxDgw20w0jAh6edFYO5LFcKs3Ei
d/8+Yq5zET04t4nWrCX1AuxlUSXxdV+qi45YemFkfJZMyX18WLV809kq1vYyE/mr+yloswqMbf49
qjHaJg16Nf85edC8nSy8PPkim1Dc7wfvWZm5xkbEz4k4qiYW1sC2lEj6I0IboDXwEgP9ziNoq8hM
/CUTP8YvDQ+Yfey99Hc2BtQV164r0uPn9rupcb8zE5TIYVceZ32EELDs1BuIDNhUfmbqQsa9JF0Z
CQJNk9u+YuG0xUQiWvYswiu4/lZ8arGP6jOD5jnI+f5Je16KMz2Ap0F7oH8h0qKkri4c35SW+M+v
26KM22i0nKA7ioDTGsty2tIlvH3yKflOok9vaBVgVFo4Tr2hKnQdPpXqAkcHDwLNCLRP+ixYFdZp
3eAFjeurbIJGbPWIVK/DXlQ3VgYmw1F46iWNNMsZ9Nxs39iu6gu09cgbbRkI/IKk18FKg3aXcLrm
2OA6ENXUjZ4xsjteikr5E4b3VIZbL+DyqnxSxkVWkNTb2QVuh/HeGXiezXu1694bRbFlo+VpFUCU
nx/d1pS9V6YGjgfFl0QldxUigZ7xhcetKZjX9huTkjLBOdQA+c024U+04SZdG3ldAfJVm555OzSQ
ie1wcitm58nIfl0GzsTbee2Palmqs6SY/okkJL35gExlqt07rYK/ACqecTkHUe+LHhMAJvoAx2am
bGu2roV+wifHhDWu+0AoD9mjWOgUBPwitf3jRf7EQZLmJ1swdgsmnfGWBClamkgPzzKl7h+3Xs/t
hPCYCb0P1hlztLHkfYcHulO3gcpDcDkUY6NRr2CoxWrn0Nzmi2HRdbnp7uh3VQELr9QN//1R3KME
91uhUyclvEOuKL0bk+whmx/jKZKOsfYrgBv+vDO2fRjTNq4gEIqyghNGMzpQS+T+jhfTakvRnFql
A+Wxb46IPmo2am7SzXOTubEG3Ql2v+fZdvGENLSCkaSQJKDhhN/u0g+Sa/xnH6Sy8UDPW+VMysRq
xIF9Gw8ZdQYL+6ZymguMtvKudyZVUiUSzRBgMrm+uwuGdNdjLU+Pm0KbW+ctPRODM2jDKgg5cyAN
bNIvJ7azjotCf+SpE5KKvQB3xfwxJVP9iON9K1homRDxcvJhbq5J6rBfpA6J53M7LBSyVS9yVv8E
ADQzVhGy89qnTxGh1rwGmMBBV7mhrd9cL0wxnZqiD0ye1RuP6O0gZ8UM/Hzf2ffPMCG90FvkRxcT
BunPzuAf18az8nA77hDIDYejyCvHYkaiyACdxD/25l4spisq6/fvEL9svteNsE7FCqthqDnY0YDh
2eJmQBqCGA5YNcILJBu5y+xRqVuK0/5HwbwJXT0YyjH9ZIC+I/Th6eneq36RiPJ+uMTJ+uf2xlEX
Ia4R2CAL5oW+BaRVjW+AjwN6Z0MeE8G5+s+3fxH8GoPvCHkerpeBYCz1w+IJGZIhyY2WVJ6S4ONw
TH8CszSxic8d+o4Zj5aRl5ELsJedOH6ykdAsCvNdjV5z8G++tZxaxJqcns6ia0REULAxarEb45W1
xljhLpYHlhLzhKMGbRbNpqguF2++NQ9DQGD/okWRJ5EpszaK435tNIyy8Y5o10s3jMfSnSv47HQp
uVEcTvbsROhx8Cp4aBOcpyYnmL+cZPOrKuQ8nvSqoUTkJFvRtzhIVdfVppd7ukQxiW+L9bI2RkAf
7Hf5z0fxKr5LqAZrX69OzztMSLhTXp7ZjnUM49dUaRt3tCfIGdEynj+2Sk3cw8CC9TodGKuMsCFG
7705X9ld7T8j5fx0SiO37bARWoI6HqA4dTFnTVk6kfLDJmnflOylSO46FSSYUJ5c7QV0JWFyoBOg
OoakQBYyC39Wh/FK2TxkpdEhfMa8WDt4NDpMjr7bT9xRLn3iXKfBKpDzxABLy5hU0SVqh9mcy6jM
bYpRMkT2l+zTZOjflSte3Pg2XfG7u+f/7Eh6/YJ3Bm6r+VCKgD5iLXDx5WIIvCnZdDMJYKEvLNnP
3dsp3aMHjlgy1zk9QfLyu//EWeDFjPNb2ubaH+zJSDFPSfyHcXPGfCmy5/gS4vXzudQk0JiH9j3q
I8rL6a36k5d/1AzzFO9nflx/vMlCqMeHxCxANGQL2ftSOZ03mMLZ9J7sq8mwYH5bnc3hcP0QIVud
EnkFf3CyrUN31r/VVohHVJBqXc2vviZAwwUtZlV57NLfMRJdpfhXPTaz+W5T8hLwSY4TIq4qSxD0
IBpC3jn0N4DkJhoUmjLH2GW7IrvF/UiQdGibQ4EFlye0zTw5nsiCVuDJjznW6QbBuYeBvMopCVYm
Hc7FfKtiDOZVSm5hV8+cd9+RnInFNN9ulg51cgaerD44IPcrDEAxUmzr9JEsjVYahSu/fYNznWlG
xbLL4u0T7GxLRjNkzlQ0WLlNwuvxbVeoNXljqeKfQwPPOD2lXzLdXIbUalgtz6/PzlWpMvo12gL8
k3sX+pFnVWiIagHbJ5f7ZRa4bjcnHVZCZ9TvMuvHqJnC5O9jJkpW5BOpDTv4ifMEgKBtY+MuLjkL
ZqzLg6NwOVgdSm9y0v3t7RXzhXRC2LOLTmFw32j493eFj8Sgr4FI8a3yyilGy+aYBmFSoPxP7H79
aEqAJeycmZcxisSAL+OTAHTi3FkRdAtdDqdVWfGMAE35mnTZE9Pcs5QF62YYHp1KxBCcjCnsIw1Z
muCAAwPD22WEOUZ2/ZB+QNdk0Dd/ZMgcYLemLFgYr1t8D9M6TDAKA1DJwdRF2Nl0tGKEvCLI8Nhu
B2tJKw30FWKnUAWQ2L/y8PsMsnz/MFLG6d/ghKjcbOnjT0igvthxkmcVSqfj/UWekodVDq0rIDOY
ra1PZFvZSH5fyck5bWhNK3z2l64SA0w5yQcNH2xD9zfTurA11t2AZS/ax7aV1qE5raIdLl+A3E64
KY07evBO24x06ksbyXjIgSLdbZHisBfCZ/b7iK0tkT8kypsc22cu3hKqLyM0eGRjhNue/pIrzcg3
55yCzoAiqq+OQV3Dx+C36YOWYNZLvmpe/FmvLPOq9ADUmrbRDUwj0kxThWSZlXrtzWTzH0WnKkru
SutlVqObp+bTyzbAsR0D3BMomwgNuCGEIWBO3SjThrtMNJqk+T92XIt9yZVKkIBxiGdeBaUANNjM
pGziHBdYA6IifNPr6XPLhVG11OdGWklhH3rVFzre6YkqmLGKKiAGsw0MrtM2C+v+Hy1U8pK4WLb7
0tbsFz96tp5eIxlOs9/XWmYN8hI8skmyZbXu63lY//M09wmASp6xHQIEfRi5FiB3TDptwylGyxMN
ZmlH0qxexTCLmE57JV9H6c6ObUMdkD7/S+HOKmRZgzH4lkg5wpxw0BqyPZGanOMEwYnS8xYBtCn0
lMeU4DEzmlxORksYmRH3x0CqhPgaeA1bsgksrWG6bgZIi2ktgxKADUDvFzmSEttnxmPU1AZ1Gdd/
tbVnOmdF1qtIdFcXsJbCaKiJY3ZGy6piDfnv2pe8yxTSQ2BwGoDDJqmWHbrKji1Ai3dTjr6ShQHs
FSOLCWTMMX5zkg+mPpeU1bnJKMeDWPYCeo/ANjVxHeKoiNMazxqQ3vkL5ajc0XeePzODJjFo4cVI
yeH/Y4sreD4M1dWC3Bys5tx6iChwLK5lhPN21/5wZsgQSqEZdo8hYqJHycZDIvJxOwkoBSsGgKIo
VEM5zrn0Dd66E1zWUtkxOFBgNsnv+VBBmWXj7LygeGUsN0XIwKLiRQGrVQa1SZpi6eYQ5ZfU1IFw
OrHL5uIcDWIpLbM8YQgyyig3Svv9QMcgiMQf2POmUgKdquIr9DumZf868KTKV1AxZkwn2PgMvpeq
wQ6un+5FEI77bUjc60X51vXO4KcKAJZk3t/Tz1AOW4pXMoBx6ih43/1eolNn2lePjkV59zlp7WeR
SWy66pASJYxONgNSHZASdmhxSde7rc6bLd41aoBjPMRPT3gujYD8hszFjDiuiUkJxw+lH31IuN2T
dNO9ODdYDBlmFSgnzBGpNgJ5NweAs077yG9gsd7cIPM+tvhLrlxXJ/fYxg8KVVhxMEAu9x8xQAZG
JhESoublNui05yQkTX6pJULlfPvjDRZeMnqpWSayqbZl5KkDt6DwEB29lOvMc51RsFKXDANXjkWg
mM2Qn0s2vb3zwMq/xFbh0WqmCkwYZSMzXslxLq+nPChV35LFtI4dAfkmIQo0hcV0nLtOBKqV1j8m
coJcLZSV4y0d6DcgA1oBJCGQyrWHEm2C8/uv4aK0tjrU4NlBHbqz5lIay36i5zY+92aktV3kMguc
5pHeXCEYr4dDhX6+HBaRhRxoF7p8jeXcXHSDqlLhOLDbN9GbplhUzk5eJX+3M0iyXJc80vtXfriR
uRR3EF3VAQSMz3K2TL3O4pAvEaCGsP7iEVt0du4e8CZsTgios7PVoTmR2/N1Sg3WYhGhfF3ByrRH
J6j/35kc+x7Bz8gjLI4/9DWsTHdDhLzZ2YTAi0kBIZ2QllohSJ/Wq2uUztq/9fNFn8jW8OBtoILT
ogV+PdlRtJxrxR3xSxRYYRAJCzDJSo/vo54GPeJGGVMDC0JU7Seyk4dA6NmMA0DjiSukBtVhFWUD
4SNiJp3kJ3FhYA00Yz2bRV8N0bPUUZ3hb2AUCw3YwsWKnlmhe2N9jCto2HODGi8ca0JiWjhuCeQ4
imzilRfRyOkZ4qlFAeq63EaD4C5xG/Kts5uJk43575rb9cMiCYijRN5xTr8A6BUgS+Yh/bIwejzH
k1WXWPobw8fKjYTHqc+bb/6aRfsDyC1VRUQm4YpfQBkZ1JyzEY92Fb+F6s8IHcus3MykXlNG9+/e
h4+Rm4O5tYIvcvjB0bHmsgxLtDjOQIb0kRIsPVoX9ZkNnEKgQoPoIHSnUtiLEq+Td3FUM7AisBfu
Yeq1ZrNB735S6QjOqvOvsP4/iHHbob2df8T+3Zp/lAut1B7pupY77Y89AkLqbvvme7C6Xp8qRuf2
6+m6WbiR8+t9R+iVLsNhpgEeIa5SpAqc4xB3OhZIyoVSF4XPM5w3lVt6tjh8D7MxHRZrveOCQcai
/eNe4euaGDyQOdTO8yr4oxQ9JVxk8K1/AlwVb3D9WbdK8xsAECCrfZj0ayXKmxqCx5OYlZIeEIpp
THGZZ7UJB/4Tc6lttEjtnSbqqQFZNH3rlzpCMvyGR/4p8jMpDXEgItt0DjhQghnjJzKr9nMCcXWN
eG3H4+YTgFJdv3lYe7fx/MXP99NWHrGvSo49OGcBdhJwilWaDAfPEjgLZTC4bNney4Q9ZMt+Xdp9
66RE+9qbuFSBRCM0dDOcPKEYQYKRV3XHxf0edVkRkCa9enQ57hyS5UIqHic1p/L6Luz76yeBi3LB
FQwBQknMhLkEye42N8Je+vyrBvWPSGpd3Z3ecs6N6yQD/jq1ohYBHaJ9SeCymafblmhsXyPo3qXB
XrnQ0bA25jYn11FJ7bOLw3e6qBApShKCEpE1zQDa4Xx02EmP8x3lDHIx5QOwOZiHpSGz/qrkSDJN
ONqNanG5Nk/8PoONi2SDhUqTnuHKfUfdvkQAOK0amigUY2O8DUb2SYrhSLrOtei31xChoXVi/C4O
QLj+CdFovI9CI+9EeDct82Sjm4KxHWdWfrIvSGVAEzrnMbRdrMV91mUtHS12w98idVS8BU/1f0EK
lECjMgBkrscxxBGsyRyPyNRNWAvj6tgSFu2OSlAnEV3D9+Cr9e2w0t9S1gBhexb6pCF697mMAkzU
1humKsKjSFB2vc91n9YaRRBNq3dIF+9E6+Ooh/CtXoe5xu82cUnfjj1KGfaTQgEDSR9cc51YNTG1
D0+AHH1mQJatQutMiL7cg1/DFq1OVigXDcjBCROP0PelkrqoeFNGrHeRoaohaE+8tkSaO/fQVYx9
2cMs2hGe/Ob4I0Ii1Ge2MTK/qBNRA18Yh6KAEQmnMHbhffI20IWUIA2NagYhxXqKA6thZm8lHz2N
gRgdM8dLNTk36WmPyNpdm0DrjwwhxDpLNPobzqvlY4ink8hz69tElTUjzPcv3nA4wW4YgriHvAmL
0YeZrQsQ2zNsHWcj9SsF+E7sR/8O2kXK6f1dcOnQXEr/pnJHyN114dgyInwi+LBQrX0l8qklvNWv
d0ZV8/EcR/e5BvkCne+J+487EVQdkHEdAkfMsOi+tX7uhDYvN8bFfeyOOp5PespnDtU5vMW9IInA
in0aVDn1DaE5MgVFPytUCDxQl/ekcbt4v6fzW9gYgOi0bWWvpITHmetDN1CWrR87E+USRfqK0A7o
LMal1QD6HA5iB567E3nUS4BKZ/W3FbHS2ivjg4q3wYxS0BltLCFu3Ped55ntmWB5Ke1Q8pOBaoSX
vkp0ow3/4mVQDmAX5TdOnonw2jgjmUSbNQD70WsgfkaOQCMNJh+7mcXZtJ9wO4iwj902b70/QKlj
vDLoTrGM3O0mAqv2fnallRss0vzyVdBhUX48+Hgc5EM8/fujtCj5kRSU7tSel8Q/K/w5ACJZc9pr
tD/Glyr8YCsMIoPX10rJvv78+h+wpzF3qpkCKtv8UZRLWPMiAdchgv0YW0F67Sk31/YpIN5+lz8Q
kzvkgCqZ1myDhz72C9V7dFd6TnwXP7zEw1KfORU/qcYLB3LkSmFabABT3FIxCPJ1YW5v0X0yhBNa
3grqFOtml0LnD2VQc252fBduEvutl5bYTTNI6VI8M8G7lfn4+GjbNyPyHjxcf3JkRckOjyTExdr9
3D5nV1yfSH+CbEVZnvpfCuyGH7yw7SmAoLnN35JWwPsMavwY12KaKCC6xi6f6Jzxehk1mZ2vnErA
3zRO2h25fIl+ELV6+11iwELskEASSM3OpbHbdv6sn4/Tv1syLtNPH0Xk450TG/57HLDUCUVs1ZcJ
/0//05UH9MTIn993UsmLCp/R09Cwl405Jqrg2zzbnGfXnPNc73jGIhYWVEN9A7h4IsQ3xnC79+7o
cvhbGU8RWYRggL1FmnRqh3Rg107tY8tTCCwxuuMIBk8o6dDXeKMTtlgIWIKL5r0lcw3U5JF43pKh
h9vi4B8uUIVitZWVVd8NE1Wjup9ZukPVd4zmapuFZZLvSHj7VPmdTHVbFBL0xnPY+in2MU1E/iyK
0NguDkUTBDvJmIBJacqZ0X7HDESWYI6zWs19BOMqSfIZYCzQpXf6J3qx4CnA94c1A7qXSB8WPVmb
UzFxObVuY+emTrrr7nQRbe2ZH/AG9UabUduUJ2WklG4O9NmAufwu90KMN+3qI/9EcMBXBt59I8qW
9v+f7yPWq0rqui3PTNPFYeQPArT52ypjYXO+rFZu5RTZrXW54+of/b6C307+wxdlm+5njhQiisLy
H9AVrURcyZIVLXo8b8746HhoyJovF+lBlZHRxyuuTJsH3uf3u1rcqBBJagyEQiivk2wVVThGyV6s
TjUUysbNEegtjqImtvFUpicuPeQ8xf4/YNO69uSToWzmU1ZS7kR1VLTMw2Ye8IF7OJ6HVAd17XUn
2BtyUTGRA0C1t11io8WY0lSzzxnHG3yAeez2M3WPw21o9lUzFmaKCMFNPi5aEsQZfTIdrTVFE+lm
0BUxwwAMzOO2zr9v78tu0hRDVpcYQJdVa+gkXg8BeUBAHPxDtB/rsi7R9qr4vXx4Ym4c5FqhoZjl
mck/ImYzX4KZ8GsN1cGe9BYqIlqh6iIN6MVzE2vzA8geCwGmY1euQ44TlFpPcLt/4KsYxgdwk4L1
IQCmaSmhS68dY4mruiItcv9z6qZArt/JMUkXTl45ko3tnlSaydK3tHJdKgQ2SL7fvTbNA6Dast/A
m4fxBjsmwK766mSzKNp68UHNype9v5OU7yi9tHg32IxqQXzx/rE/3zq7Kcs/Xzke0lsJ/QqFNb5X
QE4cLcq7b1leqhAGZ0Lt1hMEt7wno3/6489M3mbwCTWYlXUcwB5kfKf4h573qUliA/9nj2jrNx2V
FjMM61bBKHgcc48vVTIMo7Olvzh6kuSH1wMHU5Jzgd5qgnST/Iz22GDcvg2tAvgRdIaCcUNp0oyr
sMDp1Mp96i3fargIuNkvA9QhbvBFJ6vkf6E+YpaGfSJBuAWl7McMTEbRG2PdgW8+oq3vP6onvrnG
b9+8xRf5stydC7jVRURoigGW0tHYEf6vYTjC8VeD5wEFYDyq0nlOPzljymTPP4l/WoMHdBodc2cS
7IN+aF1JKF/WOLkhYWfa3ENk94dpI7XCQ1nj59kzf0KE83K+9NP4a5kYDPxGNr5LBDmxRdyNqJgR
ZUkyyLmzf4Fv2TlW2YT9+W5TnjKguN7OuMGwDW9w1rWzmlFfSTkrj0aM45S+/KsjOkidrPZ4hKZk
MZl6LgodGsN4rbm/9ME0x214GcCN7qhA4JULD1BcefN0poUC87ra0xGzyZuAh3bKBv81UNlIC472
F4pjFamDJHt+szBNYJFWNvHf3uiXlKnE4wfxvhmYzxqQc0Ekur5dyyJBD0myfaEH9V1DxrVcG+1M
aIhStlMHOQpKb5VpygsC4ThF+ZcQqRWbBNOjD7EXnixZ8gqyLMB5cypHnSMEDO000MjkI2kg2vio
kEOoTP7W71Ud3c/2XvLGaKc4mnCo1PENHXQUZN4778ERcHX1PC165qLYLfFuC0XOCDHXBdDWY7A6
wuhf3CUInF0xMK5A+EdX6VtJauTUdU9DZWdtgS8reoMJ06jWfZ1HzVOx671S/lduLVuKoN54YUom
IJ5ksiaPY88DN0eMVj61c3Vv2a8qrYMECyJRLTdpeVfwZHncVYeA26TPBFRm1pn9uuFweAN3Si7W
IhYrQblw40nmuxaYeH2xph2+re5X/21Dn9s/fmlpsKKX9lIr1u3gaEjNiibNOqF/qzOv3/5A6csI
4B9ZX1IY3EY4VpqD4XyuuHTEqk4EZDwsXd3kc8sE5oDAAOcgt5xrb01roEhcW+yoO8TgFYTFGSdY
uBb/6ZrxP5UX6BUfkxPT5dGYNKZO8E3Tcvoaaq24rlvivESav49Zp3C9KEPaCgSvD3/8+BKizTWS
pyTD8lV8DMR5zvYeI53mzrC3ItykquR1uk2s0l3zbi+ljwhra01KZ+oMg0WnLeJJyHXD+MwJgopw
u4i9hcJpchbhS+Fkvvr2G0aL4CYgX6KBa5LYZQu2bmSdrhmbH75OvFJOGllw5blIRcic4GI3lVj1
7LJPUPeuTphS15ihS4VC6wSlL56N6kB5M5cZcdvqytU8SyvKd7h8qYszfk1ME7nrdSvsW5xF7+lG
V9KoYaMhehL+kJ0JR/Iygl2V9+tnXWh02gsTXhMtFn4UyGIjgQd5IhQQACLzIoqXW0OOB6cH7mBv
6ouhtPsvdxqWP5VgBtbLszwXzZuBi+zmeKdStGXMMxFwA9jyG9I6GJ6RsB/wn/fgxtLb0c9sIDhW
unmQ+ne/+MuMqvojkEGnkn3koDjGKLH8h6wGjz0gRdKzKhG5fctnnMNVCHkU2km2ga6OFiB/fPAh
iFRUlSr/GIOw+26bwfyEfpqTXjUggt8Ly6TyT1xNM/i1AlwB3WcAc7D9Wl9UEOlSFTSAQqqq7SDm
5pFpyKCjj8JxsQBxAlTt4YaZH8XFPfs3d7KNRgUO/JPyb6NJwreBGmqCfUgvv4si5GwX3oibz6bm
OCezEICe2izOO6c9vCYU9jgmFzMR++NcJHPJCAcwP2uOMlZFh2yGhoI0SR+LX8t/027OppasBwWy
1gs/ocEeiiwkJvukWocMrO3qDwwUwRHottxc7VTBHpHny0ymXwe1+78r7F/1BO+xMCLR+XwpJNAx
7umZ11ZSb0/AF8mAHBuDSXG2oUupmoNnO/H3JLdGBZWqWka2wMzzmYcKk1D0FKyVHv7xd0LsAGzf
kBXuGtqDtRX4ktaEqrIyx8oDFE5m+tgxKr0KckmfZQ5+qjaOypYwHSH8TpB2kLTyxD+fUOfLVM/H
8UWg44cT8f7fvT3W7k2exDOTuniF01q0W46Ta5KF4QnrrwCfhkgZ3gYRnBMl9z8HE14vQ9Ap/MII
OmuN/yXC2XR0eSBCTwreiojB7LQ+SBQVUGxIDnbFOCf+BMdzBfUJq2WjFxyaCRQbTjEeETwWoZtO
gwe/Jgkbc2PbKjWCRXiM6NsuzhpaP3VQhQpA+whA2lQDDcb/WqZD6Uph+S9a6Ieqleng+v2Jyvsf
i9XN/SjhIgyER1kYv+bPz41+RZwKXcb9P8nNpavJxaDdXxz7ZQllZNUnDCkzI54e6Zn9WSkAS8SU
ZMkxsoMoxXLitPBA5TVqdDB7gazzDGoEVIBVjUGk9xuyDpt5ftQTODeK0HliFuq4VWX60ZvVpDiy
e0Iol+MNoVhaXsmto7Moqs3oHPEoDA/2/sy5hdvjKzXsCjE/7x/5xePMmOh409glvp/HSTTVA3I8
AYJdLetwdM8YtQDlzizAAmSuSyNov/tRY3JDPKK7gMoLqZSzY3sV1YP1U9dff7ruUPmMgT+EhOt/
Wjt1OPW2//LtVbCM6R4R5Kd54OcP61TqcQFAKYtSIjaj1ytU0QaZVvS9TaRM75efhzaTTQub7903
YKoU+aYHkMhjWuhiKVVWo000PLmViknikaqGIwaIeKiqBTsrtFdoOqg7WGviQYmXT18UGGg+D3i6
TQNXf9jLrnZa7UKpRNY1+7pveVKl5jk38p8XBd4DG3cYrvyj0LPPhloGfGS10yUFI13gkTvoNehx
Z81iwlfS9AC9YjowVCjeQL2in9fxJx6zs+zcToFhsRrZIt87SVEJqTS9cuaPcL+3uzNPkh9W1r06
Y5XQAhmJWJOEI7JRXNUS6d1Cv4p0hTVRDQNz2KZwozHckcyqopJtfRhLWe25n9n1cET0/NfOQ7wS
yH5ejtzxHCs4ozSqa54qzesBS3QVnEenxsA789hejx2naG/gGstm+FXZYmsQX3PeoK0/GWQFsaZ6
hhZqGALnzTmqqr/lIgEap19npy2KZlM2n8yreSfrhe3opLTdfzRhA9nk0L/V5Nxmm1LwTr7uRUZb
D9HEvbsGYvYub91c80QwUFRQMDnFhmQKIsIbnzN6VaNFxL+y+aMNWROD2KQcK/Br7DYfEnMHySuf
TUuBwAr2c5iVSeqmhzY5GfYflaS1SnqTIIST7j5c13XEMX00I4mrYN8YU0OuVfLr/n5xc5G1EkEA
hH/hHA4HrTSOXAAGbmUcNWPi0rdJaOEuU0nCio3g8th3YAazwoM4b+wTPvyc8qoHmj1iIl5lOEJf
P0Nfgu6lwlum37FdUr03HIAchbprB3s0SP+Ivgx7cWfOMrqLxiztppAx5vis92ZI73sNUYuZ8UTL
e115hO7TV1qwwy7NbvgxkKQzPPlQCnv5VE2u84NejT45OzGHL8j365sg3CaAb4hp0XtVmyHn5M6N
QkZO51+9XNb3hajFEAASZVtFfEs1fJqmllxMHiZbYZ0sInNVYRFyMiVugFD+xRy/3UqVaqjD3reA
5K2WnU2aehM1JPiMWHLXUjuO/FsLBDS+mAQbA0667UYI3rJ/Y7m5sBYtKI4fbAdN6jd8vJFQUVWr
agDCx/4wPs9/ZtpuP55HT9EwL4PdyBNfdGXJNirFo1xLUV6vpMjFbXOWNsrStqUPy3PTJzQExQia
jHYCxG4UR0PsHSu2om+H5uvarDiag5KrG5Jh/bHr2CcWsiy8Rnr/PuB55xLW8k13aA4zzbpglUsG
y2Tdqljh4SKQNvB+99LJQGc4B8FYfDXh35cYtNcUUAUAk9zzm3QqqTuaqgMv+Ha3L9gvzivyx4yI
+SyaOx6k9Lrla4TmFZ8Jf552tD/3cuhoffb/o2yLWwNsFVfjWX8Isel0eTeVi31x+dGCkEvWF5Xa
oy53W2628ZU4Qn3C7Ncb1swwOl/EEaY0U4pDQYpfzN52cquIGel9RIad/GWZUZuPJtZCkKyyEJuG
q8cHrvq6S4gq7Y1iSDCCdRseUuOD5TndT7GeqiC5lp3hKZpGfU0wfSzDrovYWmU+E+02oGbjKlDf
X39fwexEuuzlhvIv2zIjCGjrqbKcvyguPFVj5ZQOL6VjnjBD9hlDgHjEU49cJvV6l3K82mSoRcjA
Z2VPrY4T8E26qrgrNhrM5cvtzO8TgT3pCs5l5u7zLtbZhPm7rnC14XK8M913Kl8MtsMgdBsZwPGw
MdGS2csEa15Lsy7ETAoWySD3+I2QZKZfiF2Liwj1dWlR0jGhPv6Y6AwJvzAAJbcR++4NdjeSoIVp
8ayoyEuqf+y2sOznpsYwigdFfv5WmkVqlDMNJY9XBhupN1xtqvmczYjvTmOPGWek5wt+xsH2Elve
yUdORLuulj2QUf+bCkEHxY4xp/s9hoAWDvAIHQ9sLR78FXjsk/QNTlnGp9RhqkdNDFU12oePGJ3/
iJTWMylsaaK0kyY/ez8j8PMCuwldG1/zR3FpjBdZnLKSZDIMUBzPcmfHhwNV3D8HDBKhdyeS37xK
L49xx8ma3HnBAmRoDL2y8hrpzIdVBltMWT9NRenYB3TbeqpwgTE/kCq+hWO3YRC6jXK9d9dsG6Jo
Rqbc9Hg03pXNbf/o3pQPSevRUevUvA9ECeGspn/TcJ0xm3OI1DYvdq7a6JVzAiRQi4vdLpsg7mH9
9Ep9Q97nQh9GYRxIJnCzD8X7Tr2IssI29GtBZl5JVc6VYhowRPtBZos8DHLzjNj+O2I0aiHle+3q
amT3n1OMMxftt/Rr2D5z4TlAOlxkogNAVE3gDqU0QRH2hLVlUb+xcym7Et1DHr92iv+BWVHghwEC
kCaYCsIE0JT+SSl8UKHbaSRCCRvTt1eDmFumttVU1MDLEYBl9X1rqMyH5cZIvNei3isa46YIk29V
pXNML9mwhkRu1qcYJb9JCKLdepPhbbfdQI5h60SpG+vTJ8J220G5EqXf/rZ1EmQ1k74cui/Idtlr
zgGNB3SeDIEEps+2cY1lqqDtgiMUB81FG/3YTh/0EqNso+eMa7ftufNRGJoEQIsYnIpiEEoojz/Z
HVCwkDEzF9PnYFLUhGFiIrrUlPOMudJ0amsEeJrC5j3OLlgVMxmfFSPlLefXfqq0YRdLnSiIb7k+
o+af7OrwPK2g9sokUjn4ia1yCCXjzXylqP10LAEZwNWVZBoJxclS9LcYkoE9yz2PEKgLAAd6kiXf
j/EcxhwVb8usB1d7ylYlqtKFORAgpZioQ275uZWmCc7U15TjBfXRc6QSk8p3AaSSKZr9x1Kvs2pN
CDpxkKigIkyTnODXqF2hohjv0JsDRtbTyHhgNpVH8OWu7W/UPfOcW54FSE0MlJxJZSc/0qOSa9ZW
Oq47OaGoCOicbhNf4ctQdzvVbNdAqHnwXyKqBaS1N9dJ9EJnpvUS/+pm2G2ap6lo7f8HgaFn7dB+
fV9ejk9tPqc3o32zIF9KHOgUSubiCea2b22K5eP2CyHaamOoiN8UzGAm0Y8+ldeJgEpgla7DriL1
PWJ14c1tKShuPNgFvvBkWn031LOX7lZSsl7tXhtcS1rzhkjN6pbrYRuLVtVX8hONZhROCt1Z3szt
kHhx0wDMizqIE8zTO1KGuUHpL7ZOQ8L5x8Pxve0XGLjMaKvJZnTiFV93AogQz2fFy3pN4+hkgz9y
Y4Gp+hfaQT7b5WmxGP+wCpl/XY2og9hHMP0W7MpdwPpRks11nC+g9JQh1A0+b94AO7rrIPWZ20bv
izMJhfkIL3om59baAXcNUpHyVG33DWw+2I+drgQ1FueAsLCOov4AekgKnhXOQitVqIKiV1jOds4N
r3vAAFw8UIrvFteduQo1LCiFucQnhHwvETVUBw/82g7aKAShib4U3BzSEiEC0aQvhY1eYh8LUvbD
b9JnHr8Gu/59xGetn1vFm2/gPBUy8fe5LqQz8dvhlbsnrnuNOWZCwbyiyXfV0PpnsjFoMRhDl7Bz
QMMQcU39HvATcAvA3YVeVMxw09Ax7R/7gMGlw4p6PfT/ivfUSfSjnyfKRopYPa2hO7FFncZL6+xA
rh+LVPD920DiLw0SwsT98NTwVLXioH0+G4v3tbli0d5bBMarYsz5m+tmdaN2eNXEVq89i+nB7+XF
LSo+jIgkhVFzoliaVa8w+NftZDwFNI/Bc+luGnQacPGRiN4znFHiLjeAGeuhmCcanJtPC4d2plxI
fw5Ckkgvxp1IyKZXP0Y6epwCnzM1hI+ZulNxmwezmv4LyhYcszJlF6Q+BAZWOyB+fa/HwIuMQr+k
3YGS8KApVN7KjdxBUtNoWz9A2sqyIjMuK3ZKQkggCzgYHDWIahlvumcBZB86KMD5HJLZjgB7xmzE
P3cYGHP7zFA/nv1q1aw8vftk+7X8Zk0X4cZXKN88qz5zhOeohjygW27Y+Qp0t5NmQQ9KC4x9ClLj
uxZEQaALdzZManPuXovHXrjvDlVHb9XJb+1S8MDmjWt7uwBT7OtPtT4LcnJbOJjrqCqZj1bptYpw
GkeTcTZPRh5Hca3NXMfMnHFfFiBzEZCgDnLgYnVjrlYlfbUcKJhozsbhqdD6vLTDAjT01O7TiUTa
+aH2lcecNnb3D7PBwuCsMWD5dqZdc/YEAD//0i59GnjnKLahu+7zSca2Owzsrmboyc1sUhUtXRiR
Ya+m6H41Wrz79HOQC+nH7npeEBHvjIpZBiSA85u+3sVcTPgmYiSUIzC7nrErvVQlgGeri0KREOXo
shsEMsJ9etwZ48sk8gNil7L6w5aMGvkQ8JbsEusKz6uD3C8sMtwe9WMcqtGd8FL5bEFnVZdQmHFf
Xp3jWi1K3ngxAPD/E/C18bn8sTsT9Dq+mF86qNmKGtJEMclVWwcEO22rhakJijK46SdemLB3z+88
a+OWBfYhUoeHbdLyh9zwpzV9CIRUoWXuddiZU2L4IJGNsT3Na5PoJcseK0KJ4L7+FwXoPQY3/NC9
R6vo/++L1AoIx653g5EJeRju1AV6dWbcdbQkddSZ5h0WZRpCLyB0c0TwDi3I7y2SMeMPTDEV5nSq
LG/ieFyJbmbKs6Ik/ZxwS9sW9vR0hrKrs4nGsK8SQx3U895JS/kphTdZtmx5nyzB8allcfmAaYkc
s89WPZMsMD2DqWGFyQoscZkCJNXVlmiXhBClV/rpDh0xBCRBTVEJwF8NSp9w3AF4M/NpdyVKJuRt
OnJE3Wz50IXGpOIpTcdpXZ6sDoyTQHNJQMYoDRqe8+xkTae0R/CoEtPm1j6d/RzThwOO8AoEzevY
m4ys6Ur0U2qTjJvaG2xo+h5wnQkHXBpkVCpgsrQ01u+3vqD5NR7WpRU8oxM5lRyNaBDYTJnmr+2i
7IDn5nkmddgDAuT06K7/Bb0+41UMy+i62R0w6ImlmqwS7GPaM7PhkPCf7QU3eIth9ogKcuoBdn54
PzmL6wUuKbFgmU20D5sWhCoeHLmigjQl27uQBEnFyW0vGRbee7XOtLawSijgbCCCU6WelTKrIqDq
rHOwZCHvwMpujPEydOdbyJCL40C1px5Xp1Dp3LUwqvSfViIuCXfSQ9dNTKX/BjmcOfHhlaqGLqK0
cwBerGh24uWTwvPWM/k+sNwiJ8wVx3+oqIjwQN/WFe9MpTHkKXP5mdr9eMtciBINPLDa+Y4uKnfj
mS8ct0kHp/d5INbh/oUFCN77XRybx9meSro9wulDSTvsdAywODEzd4VslJrU2shrzYxDAXwJia29
BVeepbILwQCPLHCONyGH8rvVoqx0L/JRvKu9S8IocCL+1c5PxHNUWrWDtX6UNbUc6o2KBoPdtLza
XvLDbl57H8KUdAzfTerR5vLqWvb/if8y2gnUOUewTp5lTSehqxaAYp1Sui4y8BErntTJffNWkiNr
16ys2dY7OX1QlNPNaeh/n56Jxv69EahIdkufpgEm+3n8SgisEu9lmFMe2d22CgHjvyllMCs+JoQK
6rn/SB1exJCAcAH+mzHe5CNNd2nfjqA1D7iBFy2BYgCrSAOP5bwQAZwhp/nfCg6KyrsGpVg0EPtA
R29CnzeseNBG/EINDVeeO9HCCrrvmIcIIxVjEO6lnTib0L6dIL8qFawHJX/cuCWcH2TfQtGP/cJ1
bEvXQRBHJygKCLxjHSnVVgA3bmQPUKLcgDKOCocIdKt/J9TFiZqv1yMSUYiC9tm+NzshUxP3J5lY
eFVwVom5btgHwZbUvozRj38bs2WoG8rJ+L3XsB87AM3LYxdOZg64XEpcoDdkjT9zS5kM68ppZXaW
osyft9VimDAqVxcN2HwnOBvGXs51RgXHln6gWu9Deqdlxi06Iyr7HVrQfNfg02UbdHoxs62StHCn
75ViusQ3Kw2B9HjUYo1Gkglz6BhMA5gpijF5JMxxuAMbVAKFzPjKh3QTMfKDpP5edjnNhQW1Yv8V
pRHKN0pjK8rCZoRQPlxlnsD2VK4ciqskq9PCIL2xYgyuH6/dVyBz/qkttbEKd/UQ5nHGJwrYFiYt
+Q7PxEfkFXNMazVPq3yU1ovY19DUglUqxPT5dALMWbvPb4H4FV8UrHTZj/B3IaTk2OqlSNgzAMj6
PAX2FQdC9897h18TxsyzCUrka+ctvmWNmNJ1ODu2kDpuLwqvejjSkE3kLiUviuttU62LugG9dI8S
Bu8Y1lTWIflQy/7v4g8WfjzNzLmiD7QqZI7961AYobYFAv29gsSWzKLcTUY+Aby3ATuFaTDlwFW4
/RW+zHbURNpabhSYcIftJ/YX4yoPad5aizuSkfjX7/YHOSufYOGyykJsYOtGwuQ1O9lMs83quXrh
AL1y0srcQKKU9PXeO2/O5ztFsgMdEqI3oXwAT6zqWWnYO0jI06yM5yRfInL4W0nlfhZRzM3e+0n9
Oj0VtrAoQBSOxHRVs8C7ye2Ls1dGDUMcv8UKCAgjyuXWSHyi5MN5q/1x9xfzNBGUuIFwIrrFsl3u
LOpnx65WtE8M4iSgCj4JADCLaLstyx/BsFH5cFmECnZAFjDyyf2GDlIF/x7c2Y0ErHihRTgRttLc
uMqahMGW0XYMtvPRRejSrGkqFqbbm1E+SWZ5k+cFfM4xxhEq8V1A9yFk1fWk6ZKgz7vbT3ERYTac
4SgFUuyF9Y4GVOhH6PhZQurKgn9x/992ghZxpPynRDdSVlpiMkf4M6gc49PT7TU8KlYUfwQI30Ru
FpOoxjzdmpOPjvEU+WmH219dEdoTo3E1MTPRn5f6/Kd//B/xgg0rQD/WA1sDNpMZ5DcEZ2K2w0fr
40d0YxrE61gir8Hqk+NHnehgpwjl41fLmcTJOxnOd4O0LmrsEGrOBhUsCC1FH9EDWTvlIVPGMEIg
rPCUiXOCM3Lj3Yrs0pJNZx/iiVZ2dI9KAiRc+AyaCsFv78CTYVejmbE9Ssj7VvaNGMWq4HC3jN6P
qq+WMY+03fH7rt7hYH7LuLI1LALzViYE6hCkPvB/fKdaivrAI5MMvRVR7y51PGtfE5VJBP8vmC3j
wmkUK/X5TiuYkZ8wCtfR9OINm8/jbg2qdFAZs0ltLlulC4ojbnbYhBXrpmRsBW9rfIwx8e9mvqUe
d5aMTMZpm3IplAjX8pP1Qoa+J0rIB8qsRVWYf7jGVuGjojAcjvQWBv4nr7qUsc1X0l1b4ExvpCcI
ugL9X0kPQqCax+r3/gYekawpvwTNZpNZd8ZdfMKI8h0zdLhu9aXcq4sP0l0As9n2nwcaWLC/sZhO
mV3lzKLxBxaHyq6Tz+s+w/5fzE2j39KNZ5z+yyfz1XvgXmVI2Rm8cHPrA7opMJX4/RtVMDpZcMTS
DKgtoDD55bkUajUNum+L/m5uZuRSqnK4MzZYSuwvqTYLx5AJyR/LLanm3PyFjVa3m4sP/d8/LFNg
/pJUs26AmYz/iWbvEt/La0bACT3ewHTHbNuo8/C6FidBg8XijjC7Tj0QtrxMaplOs7d1M1A4oHZN
gr79DLinGDC69tFWznZO/h9DG9k+IGPNfmofwCmoVC+EWDjNUtZ5jwlBwufzhhqbz+xEEo0kCOw5
EPEOYXe4ZSRVuuDuHyCF3J4m1YQehcAtxmUzu2UJBZjKurS1iCc4iIn9+h7xLGbK/8gwqfQtNNA6
C/hB2qypfa6WgSbf2h0ENKIClEE1RjJCWFfBzdGy4EjvD2uDMaxtVDXjERGknSW6JljBRVPlE2rC
x2GfBGbJaaGysBen8u/7eshO6XRyAIntrKrNZSV9eaURWYxZKXPlG0UGQltYIcRxP9t3egIeNyvQ
gIKzeNnbNWWcp+HzkXWCRG/8bK76qvBZzXNz4pS3SZAPGMPFzlQTu4GHM0PNrXJR+KlZPQaG+GX1
n8MZd9yaSqltOIxZnt3MIfD6M/E1DkFK8GAhtQL4fqsohnk1fngZlXMUbyOcw3yDjffN82mQIGhx
MvFBe8aJICGP/hi5Esy76ekOpvvBF8bnjPHYDur81KuOFP5bwKjdKbTu9w4/xr8UTRl72CApuk+o
yIu/TyFl82opXkPK8C0eaRTPQQE9piuhl1raHgJ3k5rK0YiKdHTXFofvG+BAO1XvgRT2G7ypR8sC
WZTeWthL6CMQUwqrID/a9rGv4N438zNQkpHUlQ71Dl51UGqCOMCTrx3jT2RGn2LdmG0cX4Qv5+F1
nj8V3KVX6ewOQTNChjinBEzkpiw+knTSxh5HKfAlmLsxXrEz16U8vV/PTmxLrHldAU1ngsiS8arB
qJp+xkJkAA6kkm0yWCA64765V/UbVlHKs2sYPAbONhi/0/Yjs7stOxZtcV3TSWqS/VbwA2xQxexO
FGND9qB7rQwY95KtApSd8sSN0Dp7ED3Kmsp1QOUiEiEfq5r6I9TEucM8rh394G1kjeQ5d49zoVIb
K4+FrWp6R6aHLR1i82dcb5vRRzLiBTMye8YFvVe53GuyZE8TPb6GfEu6ivm5YfTTPPhcP75PnnqZ
Z6JzWRKR1unDohJ3NPRdP3NxUinbbHIZF3SqVOjP6faUc1YAxAIPh3KuL8h4gdOAZqahHOAipu4s
opp1BdBmX28wxSdIHa/dIevCk9a10EB4eGUQ4VQd1zWk8Wo2SPtqisccN0FuE6o3PZQO2wsKwM2n
GBd6ZRsvB95Y7pgQ8Cdqj0SKOHpRWcp1yjCHK2wVxTOur80nXzp8L9QXI6bLe4K39j1ibpZ3L3qi
dqoCLxi6g1IzgtNWlRDS9H7H59urjLuMjAUsk5ezJcIYyzbUPktoy6HHhLR6/w8bqKZmE+SqO6Z4
QClTB3xmIk5/vD23ppPTh0EJLCPGLAlJW5v5TfHOPn0Ox1KU25UhnuK8gVV0fwjuomIVrX72I2YV
7D2QZVkHqk0X5PIrCaqAUt5/0gq9ALCNTVuYIMRoOLAZ9nPoe/tWIDA8lB43PLGIBh0gpvDuTvVt
bPyymIytexgYJ6M//GPC6eooTXY3UXzWheg44MsPBBWfP11efS1EnfI9xIvJaLKD7f/lHmWi/h9A
l2q3gFn0VlD5dnbzjPZp5uu21aJfCFsT7VUg395diFtrE3gu38BoqWxTRZ4purbwjtGQPjtqTbVv
UQgYVMppKY/lZ2s2QPHXQcrx0yFpl21GFA2AA9KAGbLcjqXb6fBUDSA+r1/r5Af05Lq74Z9OVA9I
/SGO8Eu7VqMnQU2LqXM3FNZJcH6Y5GqfAELrX4wtu08fzCvoBi4+KofDCwBw4xlS86GF621k/fp8
Jhx0Bj768DK2pEsQp9TJu7HZyXqC5Kp7YnUgIy/XQk2xTYqkDsyK/cq3IzfQGb19XFpTyl1KxPFR
5+2nKUGrX2HCG9/p8tEHOoDSvxxKyjCqJmDxLX4gM9bHwRq3X/AJZerr8A11HUV+MwArLWb/XcX4
O73sDT2+tWzrAxgf0DgaSsxr4KIKyy2vcDi7Y5vxm/eXXESyayh611SK1g9RlsbCQd2lGbkWCy0B
5b2plpUO3EJW2TdH7NvGibvD4jMfVvkQ2xjLU0Q0ti2IwLE3lIrr4vD7EVYfvYNbQDU04LRFcgJk
YetU4I8qRdhoy1VajaeICej6q0chvcLkkMup2mmBPZOVwdWQKVbI+cPUVrSTD7/w/lrvB5JTx1+S
JHchVnIQfzDxsL2u1FCPqh+sd5RwDjpXOLuJAqQi8D+nKtSAEqJhlHv7wFOmnXEN0D3mgd7tlcMY
Tj8B7cI4H0fTPOC4zJB6bQS43fSOKQqenFPIaDMMHSrTix4YLdDkTcfdIHt3Y5vU5/s42WP6fqCZ
N6UOyGF2+7mT8EQyJnihgj7739MbUm3N+1zSpPzAVLqS4Vq/8nqXRjM6NH0YHDfyJEMMhC5gCwgn
Pl/cuHpmWQJnKvN7lG1WdzUCQQbMUHKAMH2lpifNnDxeYDNu79EZXus2Mqjlw+glLY2Njh6rxcK1
F7ki1ui6oN/TPa+85PbnCTo7m4PtZ9+uX0RnLOWe91flIVAQcMILNF0qVDvfsCNWxks2gNTsq5Cq
BRRBfUK2a9lW3eftwCUUBwzH+YwqNMePAj7Fa9cG322sKqnlJmiXNbaup9kvusl6JhicH69BZPKM
gcUzezpu2jGVyeCjDJLelPB4JZokcRLRkjqExjzIgPEf5oSUPSPiq+lsyvivCm6dA9XLm2L5XsGx
slcRE9XpkgJX9+n6gN0tl/wkZCpbOq4ljiPtKnmf2gLWfCNiAo8P/YNW/FG+rfXAk62noA0vRCWL
2CLiQkKq5hksmANN6OzZF9LXNA1l5AWdkqht2bncBF8HKIBdejNQHcXn98oqTKPcwmkBEqUdvU+w
OjTlMTB5qvbE+2wW3WrVT58aFubU47sO3oHnbnbeTNMMGUr42CE9xutV/fOLPPQkBL2xvZu4UgxL
uyRznpjgEGNO/mY/3cmH/LzesphqfISNT0wj8/BUXbHG8IFi1xYr6DSgQugrzWeeXyuSglUCErip
lksn540WjOYPNfYFgYsxQbd7KuNwPRVCrbb/2MLYyP+0dVCI5YN9D7HJN24XqdQXrMa3ztHe2c44
409+StzkFNaXW4Clv6xjw5vJuy+4LFydeuSI/kMRKZQVKMHG+N7j1Eqluqsl4tVLtRmLkUbmvV5I
DUctZqZM8AxkRsiZ56RQy7Gp1cA2Ah1vVBbGJ/6eCDU+E6Ugyr7kTqxFCYvNHs+1AZL2+be8c7F/
N8SgZs8V59+i0BwrqiVSOCbo3gYHP5wTfBhvLe+A5DDRdts8RzuwjhV+Um1vssekV5qMmQpj5J6a
/Nrrn0Dl7ugm8hOPiWXZpv+ryD//q8iJBO4spd+OgLfbaMg+AvKf84KqEiK7PqRboUrAbT1mqLwh
NGrlYzG0BfufwUtFKeKOnu97QFt1uFfDxXfZ+jf33160EFPLeP9uKGUyfzApgMuFGPH6Tz0JPSbG
1glblLEHKwMJGBCsQzxsmoIYmGIKgDbJSZ0ftEuFRfuGtmkHFkk1K9IZVQypRVqSC/ZDxSD+ASyB
bN8/h3ghrlNnkEvNCUVnX9pTj2i6BqJzMCSbf7K0NhJURnBfwgjo2ZXP1auNa2d1ElTPdjOFm6b0
rKlly0xOszVorTfq1lP5i036RRBVRv+h41VrX2Cas49vksscuRU8m8qRAMjr1ObPaoSTzdG0HZWz
Qq1kMFdvIbgGtwfe+kah2RTAlFW8xF3l8RztZZ2w2RxeOo59Viam5hsLeGCKMNUElsw33gWSAiOy
ekogrrsZNhqtyTO93B7HW3DwucrXckgt5j0axtEd5qcxkZWyb66Y6+5UqvmsfLYaDHH06vXGPEtc
Fdzl85N6/kVwUoiuL4OLJ6iTqOgYIFyuGKTtyaEmpxVypVaj7S6quIvjymjrF73f5LOqkGlQUQGe
IQqa8zPCrzwgQ/W/aoE9ibHLWPJlE/i1QXe93CX7ZmYkLvNCO24gfaThARvfnXCgQeUvVqQbrTyI
5hckQuwWYGFLs9R/NpM2FLUb+iqkvg6jOjY3BB2vF06ezEm7ewzrqWKbWkkr5gduZBRN463IDu7L
AzJ27nyXoUxXVM5lBDMVu2evq9jJV6vX84d7L9uxM1ZvN+4FVVaMxQeCElWffIF8XuD1+uQPDLSn
otKznnEdKLcNDEwWHtzXSV4DsmwBKnXuOxPBm9tpND1vMBEfDiMchByWwheK7hMJEPS+BRm4+EPI
0BGsAI4wxUZlu7UgQdjBoJIMY/lB2A4SxCC9pkddYOqTRG4+sFJWLXkET4o7UCpS9hE49LALNT4V
w8tpqMKe6Ll1VSH3B2TJX4coX0N1eMro3ZGhx5jg+nK+6ficuPHN2wPkpSdO0N0WSH9scxDgpb9i
Pp1ngSv9zn36eZ8Q4OuMO49/Ai7l8sWlxbBAea/3BWVRD/eyz5yUenwvEgLh8BG85sfw75cZEouH
9OBt+KppjH3nWhq/iFJXx1SB5j5+7fL7idWkSSQvravIYakfU5FmAwLfKfbtei37RrVCR798RtXc
Dk9YBOWE6X+mgWiIOxB9kJwrx+zAiJ/l8RW72yKIySGKDMnbLjK82bfPEGYN2nUZ3svOVfv7zOxW
qCy7DSCpY8hy2Z7vqadn5cLwAjZnesy301XYiIP20feskxpOnRlo1pxt0Ko0Rca4GnkIs7m6erRY
amgGoRm6dTj9+F77lv1i2z1zcY+nLCjznl4l2GZXBEc7EvMQwwIH87AeHxKDlw53iZKTkT+5tncz
Wa9lzqgHfLDKMC7ywS9gFwlmi5/ym/B1BQ5i8VRblowTutQHo76sYISUIU/wsgM8bk/ziKlYKyUl
Q9LI8+qometeWoJd2IY7rjcSDR5RsFfDJtov/j5eFKmH6z6ZIDuVwge3vi6hUAuCFr8orvA2cGlD
mKiPt0q5Hrafb2eBy5rqrUbvZITYxmmP5JNF6gxWO7bc1+tjyZ10PymhjJIwiNUEg/uzJvX9PSvi
TW1RgxaJmCWdfKYT8tTzA+iyKMOiQx1bGpnvHRzOWUzTaRYVWIASDmqWPMoO9vdghgk/wEfq1c47
JoAcKmXujhCkb7WMFPFxmKIL5iCKZ3Jm0T3+Y5mCg0K4+FHpRpVT21HyBl7KNd8eZrzQcVdr6rTH
r4aFsKCmvtHyreW1Hle6s5nAI1mh7zLgS4hfevUG0BiBObhDJzhlcI7Y412En0hlB2zeTyBXh7fV
xEXfhjQv8N6en/NWh9fL1IEq+LE130r604J6Dh8/KjEt+zu3W0TLVwptV4xqAvxeQXeGRvU++l1r
TOHAl+iLhzfyD3QALUfvIQdoGElSAvQUXhOikgN01xoImUXpCtv4ATUFZD7bhCABZnMrFOhqJsiZ
b6ZSk3xQmSrrji4JX0fW6GzaCYnZp7LHuTTBeMy3KH/8iAbB+AvSYlMu12KhW6UCKNYdsGyNScHE
qy23sJPLDsEFhcDOxBDx15mSRIRF6/Tfx2vQpuX/mBG73xZa5OpmD64qDGtjW7ecOz3k1huUKTnS
zDB4PC9ZTgz6wQo3qsvkEn5fRNDFjGgo3WOoZggPd0aKBH2A1jelZ1y1rcoakLiNRqwnJ6h8oha4
Cu925YL7EtKEO7xWyv/Cgw8gaANcbnZBanFQeeSH6oVr6mbmFgqhELfnnELUpyIBkv1eSfRfmKxA
FygBtCSnG4S8v4bunzEzF9k8J6tSvybaWC2nmRbW4xGzc+MJ0tkhBr42FIPLELkVkXzNh1TVybD0
hM259OUNumS6XnvzeSdS9I+dxe2iu0w9bazALD+PCtysWEcph95bN66p/dG9axkrc9htfYfj+Ed8
TKnOIg2ChAZAUHXDlYuwWGc0zhhgg1o3lRG1rAEV3veKjg3N/dso6obgI+OBKbuMISykR42aBH2Q
guYPFaLazSSwcAd48xiE4dF+bcWNIxAdjU5ZECvBeUvD8p7kedqyQgedi9Pi1qqwwEBZ2RD81yji
6uhiFldPjXcXT5PdHADbZHGeLdTtjrOZQyB4X2P6rppyy83D8ILYglNbwxAZGn9lZ4FjrjYwM16J
HJdSmErP5mtebhPSH8PvuZRj+LoAhQpZFueiXjMIy8aHn6wgfxIiy36DjpGwMAQitZLqDS7bCE3l
ekj7bCG2oykfrkQx3koWfcBqgYLLjJBEeInDsv6M3y0CpIDROplvdKaqecnfHGrwrMof56AxVyEp
H72+gSTxjloawlVePUntJ2e1M+LsgZ+a120UxuLb97kGUXcn2h5d83fgmhdNbm6Ythx7HCmiEkJk
IuZM1GX3nSfA0wtL+8bHV1enmrFtYvaNoL+exDGOb4uu++AQGBB4iiAFSrhRv+Z+z0PyIRA7TQhc
ZRwWG7dinzH0XFfwzSVxaWVoGJqndEJ6zhpMM+SrYpjVURf1q1klEw8s02XDcEQEonKrPVVJDkq9
KNvf+8vtA+GEJ++1nXjIGwgaF9rPEaP+jpgesZrT+4zI1eCH3ZKAhvE/U/FSCqR37Nmi/DAS8dwF
49JpUkcByZgly/GdUuKdioDKiSuiI0HKPY536BTAuOY5HQL8rZuK5A+A2X/tprrGxSU/7mjnH3Vk
4D+Smkihqd7USCj/TWpCCabR1j7tWbTZZ7DxhipT86Rs2ccAaqEjGtM+u4Laj70S+yPUGj4rDI9W
JoAkENfUUKNm6YRhgYSFePqMHQpM8b6UTcqhupJ7cW326r9LTXm9Kw+qe7SJtVjmqg9g+9u077b1
NvYtPV5p6zyZAY0Y/XGBVeaudSRq3Tf+v81tpujooxa190jzeQIg3y0onAgrEmNlTBwuiwR5lggp
L5zQFAPrZEcw+El+eZwAE7F3TykGOZNffELu70Ry4dYxxOr7M//KMMVDc67LiMGpb5qiSLYl1H5N
xyZspN7mj5/D+V/WqmqtffFe/Ynk1BhFO1tblEdcPG5/Jaq0z3MP+i2/obtpIbCgKJ5nbeZopLHe
xH1V/mLHTGSQlVMDdvuGciQD20aLZDmsCjkk9rZK5vEo3SZKcTuqGpxdadIz2tLI6Zqzz2e72T/4
8FcBHp1yOjEMnMJz2d92wwqLzwqIs4C4Zt8/MMgn4V1mVCVAWBiXhe/ZEedKw3rO9v5h1MkObp4j
hDFDOhcRDydZjYsq3gaJPg+HhDa/E69XZB69++PiuMfl1tv8KzYsk3+XXWDUH/ejc660sN1xWZxV
qnSWGzCmxq0atiZ40DSkpm9NJ+ODaOtD/7/mB8YYBpImjA0GR69O4Qrgw8zb5eLqBWk3e3hEEMAB
lcj3Nz4GrrpHk76oPPQjBoNLicdYg1RVcpQ8OYne6oRVyC69fNUQH3lAMsskGvm6m2aJzKKkui18
O2tc94w8OizaUKnRQdkbReEx9Fa5bE7hUbM7191B/bIrShOqEDyS5njvTCjuNRbc3yHC1U26AXDd
ccSrLzykJNeqdS446Zf0GbKfflQrT5F1I0ynaSo6cYvQT8fWjLoPX2SxTmpk8FIWAD1mJCsXShJC
Z5Kej2k6kbswzJ8QeJ3x2/IMS2+eDQLoqYxPr9IDtkfEy588fSsAlEe2aR8j3mDYjB19+pOFr2Hh
+aSmGelOKnRQzpYMefWsif8kIr42UUxFvjJ6r/v1xBuFWn3PaV+nTiDaNzCKRc7Esq0Etpn8ccwW
pJOHHxhy6FEx8gQfJlNZO5FRKebsREmPoeI8ikhjgyPeflsEA7vowAk6/fB/juzJ48I9sjSGpgLG
JdeFpTqivcBx9XIN7lc6UwCB53bnGwfeD9uf2poQf10ZoUzDlhhqyD0oBUX7xjZQjM3efvssktmQ
kXSEKn8Pxin+mz8FqtpVI18JDCZ4slltyUaupEcIeraslzLc0FHfbh/8/GHBj770KC1ZO2JIEjvp
Hp84ShqA86UKJBYTHrUBHvpA2XUoyPUDnLRsmBklVy0woH9Mwpp+WbHHBLSDXYH54H1oVIjqSki7
oyFCUN5vBPeMLBMO189tw9V+bztVIcaLSutZUlFsg1yXH+w4xI+yasmiymslYD+/C3a7TmNHemDw
vG4kNYvCvha0xuEgY01mY0UdpQTcxmBbWG+mzqAG1FNEHijUEIrMp8R2hRfCkUfUr9VqdJBo+RG8
DMaXT4GdD9FEAuRftMSQ8o+x5GRsbkMO0GtI6O7pK4A+svHldikzHvFd3K6hGEwAWkJGMZIltGxP
eFQfqAkEBaHKjlvdBqSpuMzM66DK2z+1ktjXNoRxCYJ5KtwXdQTg3ZxwP8AXZoOch5byPfXXhUnV
pHPOKHif0z8j1+5R2z4u1d7Xk5BCc07H0V6Eg9wO2OenMeC27lnenYzfKhJ2MNjAdiyyyXRDvLRK
YtFlrlFcgO6J72pZOGz4lddNzsrC/igknxK6OJo/VYOV4RztD7qA3lYBrGoiYR9WTvFUgfn0sHAF
e/cpl6g3basFuDEtCwcya9beonH1ygmm+8lM9ZUI5+iT3NSaM86zgANAsjgU4xIXDVKIUztTseiY
bWkCxX05HOsIiMnKsq3NjaMzdnwockMdLgq2t4Fkl82RLkFMtHhs1gOXoVLRCLZUzn+6EerLW5Jr
LJ/yj7TENf9VQG3AcdZve+FISpsq9R4QqPun3J52ZhSFzTDZAL8nrntgLmILlMy2MvLLijo9fTTE
gkKfjhH8IUxUhJzQNGTg4pMAA2IxmT81XY5ZnMVJwurbYwvIoQZGj2gT/p9daDcR8MigO3/cZ4F5
jnbDy25n8g0w5UAq9AvWgzWF+ActGeboCCA+dfB4OY63d5rJN8jt+FQpiB9X42+T57Ja5MA4M3si
uTkVvK8FyFIg1bOGO8/NY7DxXBv/ECQDF8Dcbo4CskNWftx15QV9nri9bMBbYWazKZtN4BPXqbbb
BmH3AGpzKAJUV4zNpXeGiQZ8Pu5s9e+AN1PDuNeRAD8VuzrAo/2YhS+4KbBPpQv76DVw15JIWxSM
1foKboIVI8Zi3u4cWIw2J0a0dSHGRo7cLE5ciGAxYcjSXWlswxaz785ruq4eC9zm/I2D8LrCPkR7
hzFYjFECzt6twMvXB/Oc8kyMH8HBFvmPBn26f3X1AzENVDbkIjAXk3MGe49vosBjbkPvGxg1b/qv
Zv3jFIp/kRDzspwimfEKX7O5ONTJy+u+x37QBUgYv4Pt7ArfSw7STeIEuR3DZJ7rGoJYkdpIKEr8
3xhsFzdoaiUFEYwhoBge0kMnMLmdd7HR6hIZqyz1e7GIqVUrvklffNNEh1uiv7BD29WuT7BdDvVu
RBq6U6IkHLqJspIAwp+l8sJvYOuqcGKv9dryZoOuU3imRricaL1jVms8ITW0S7zskoBGq6TQSMUw
hMu4TXEAxR/2EMkeRkJQeCRDu8kl7mR8V0aJzgIOODFe7Wi395aPROdoGOvhMctKB+JqyivHppyK
Qjk2HtQ3Z5LuN4ErObL7JidptgiO7nDyjaN78BSbmptZmQn0Oy+djzCuNSm0yEkJd+hR1yLlwXuZ
ZLqa27Hfa42JQsoKLTJJNzKEDtSEXw/GJi1jvTSDf6tdG/HgS2KV/pft/q2SXnFN8bNa9CsDnFNY
c1n2YZfbAlgUt5fYX/gGL4d/iDdeMmHOdNE2tFUAD4lXlEFyW/BJzntoXMG4fObfkSVLAZQgpu4R
t7mQ8dxFxQJ4pDNqYG5aSy83ZPb2BXWY+LixbL2V/O/CTGuQ5+EIaBds7XP9vbAG06IJ9Er8eKyd
tkX16Gf7GBrhr5XTmqA1+6Y4G3uzjsmxE3NuUVZFQJFJ7noMTn6+Hz5lj34ALI1ehA8KJagd49Qz
7Jm5Ufilg9gvXfJxabXGfRNfgr4y/KQc9kgUIjP/rdDgByT3hFI8OssBAJkzUuOmS27Qvm7Fj2kC
3KuWgNe+0MGA6roJgCoP2vFQtIks8dz/+buxn+AGDzY+zbIUWfj+YYsQJ/YWgoTxcMLW+LtCxhiK
/v0Qq0a/WLwau7qDDuEML3W3Ssci1OJRHSlb233yoBGaNNjTqNFbEnAPlgRSJgnkarzh12GMKUi5
ieYb4XMx760tchY9qFJZjqAnnYuiEwGWUvSM/NHPYvXpaq9PecrJbEnFxZ69vFh5qG5v0kQ8xEVj
V37OlDmREl2TD2HbFr9Si8Pzc6EzVucFtKGstpmCwdZfbPdj41ZH4/jLIIKImojRS6V/MA1nX+h8
ZpApkWmfRyLbLRlMsyjSxk5lhDmx9y8tFyI7AAvPZ6FKANBHvfp5WuIoJ9dtG3b8rtwt/VqStOPm
4+IVUaBKuhtyMRXlhnkY9hdjkMX/6YJuDKest0Xl8IG4hZrI7eY/QnQZ5tctKzowWZXudeKbYE2Q
YoHvKZr5f+lMPb3nQHxHiaq8vSCk1ZQ4LqI4u0vPWrbo6KgL7QTSlbalBXYsED681EkVj9aJs2ST
Z/7XF70+rb7r2bC/sB6hjjRbtV6KcHJ4z2+cMG/fFxYo9Zo+em2g0jC7zpQlRN0PnIDoLgoCbt+w
DGJkPN40bWiE6PsDHwEckhjdTNhWdedk4bYbVCit33HqoYO64Rzf/jmIDMscM5/HyeR0p1L8XFEl
R352ADw98UeQQ+6XNOgeZr7T5KZE14HzqKgXiU4Ee9O2P9bH6JTBNV0f1CAT76Fou4VTC3GDFgT+
MU094WWZ3QnYTGR6ulODqIl9Oy/CfCyEm6vqXSqqOsU/28bYokkoBXQIsOd55yF/01/7wPH/BOzJ
z6SoXKQRqHngIJ8yj4ezjKNmIRpvN9HHHcYO0keOd8477Xw/eKZn0CdYTEe9VuVnu26zkmjK3mlg
fbYi7xBWsAgASsxMtAtGgtNoEu2lSRAmbqCo9ixsQirz/Ed0WebGuXWC+j5zDnF/tzOq2/WgS9cA
9svPzJk/GTqqPSMOHhALUm1JpfpVDxFehSUWl2+Sl32WDYYRaWcacCtrfgiA6pDVF/XyQi3j2G+l
ZWjEFc4v7FUU1Gn8L45iipWe/pdw5ViFvtJMfU5YdHN2kFicB7d9isdNGcY7uiqnmLbKRweerygV
Z9zqfRt1CKZCiUFZSIpJwuno9yYp+VQr2iHu2AfEMKKMzFKhanE8KvPGXUK+K+Zl3EOub3oFGNPd
HEPg38o6/2YAWyx3ZIkh21d6l6ivYXf95XmOy9DDKYA9bbVHMUUtf//38Qo8Vl8KlKhZhgFuDDd5
ilsvI5LUIYAGL/Fbu43s0cIj7JhBpIm9tZoFedWHF4SgZfWRygE+mYvhZgmM+16n1J20LT6BacEt
DTRXXPxTWtxcjorbAIwysmk09/aZiuvFM+zLj5nfksOtW3fhiaGC5UTVs6EFMsu3MWwpg7y3LcHm
vPcwybFUAbHD+3YEKx9l4kdEMKhvPcfDfG91TYuw3JqhLhhx5ouNqLWUa2uLeDjmi1RXhmYoYDR+
QRN6uCiVEjvQxmxvVxPbh99rcjxZvf3yca4Tr7NPhXcMc3+l4VdGoGTKG+87S79wWzPL4b6axDwo
iEiDt6E4p5R8Qb9tY8eIqZvYlcD3QvnJqdD6UqK4CJ5UV6gRpWe0176mOXfyEdyYZmaZV6C2pcb0
v/VW0ciIefP12r1UBKS7lfWx2oznEwRHvOZTYGI5zRH/jHobPN946PrYNN2L4vBmJJQvbM9XXBqk
bXvxCBcqSugTDD4HtNJvkHXBLdv/35EwEgc21af02MiVVlI2e0rKRakqYT7Aa9ONRKdqV8Jj85zJ
0noENHs+HkLtMzzVl7UPBqFDppXfZTXuSB2PDYGi0Y0x0ZhFAh1bB0jBLjuAfRXRLMIEB9UywfMH
LfFzKVWBIC8DC2krDAybeI9wkeFkefGENdRCMUHyBmqxfiARe69ENB9L6NnKtPMrdPh2683DWx0w
EXMj8KO4D2jWGbMB4omMo0Kn1ic1jALJ1j9efBrQpCj+SciU42SAVJF/c14XFMDEeD+QKnvp0gar
hi6+b1utey9kiTgBCmD4WaDnDccA0QPz1JkGwLI0cITMozL8lqOeigivUHN6WxITy9WDtSZc/Q5U
W2MBm747X2+8eWtg+SNjkfApR3hQEd6yhb2K7TSCBVAk3eLq+7yCnwsSkBLGspqhRRPEx8SlAYVo
vCaHiy0eTlaBd390Uu+nVsQOK0LiJdBCbjE1Z82ABS3goJwsjRix3XiZ3rd5Ua8SQynJC+Pz+6bk
2b55RgESGwdfcLQhtf0/T/Sbp2/s+edRu4gNSNfaoliSw0mlAwSwx6100CWHjYDiXXQFEmokBSs3
CmU3tOnsRykQ77YXnF5djF9apgQH75hlrVuZkQ7WUFyFui6KIikqaoyIORmwQeL/A4arBsth5UGD
UQjpJkT13M+8Gef8lreUsq5OsG0K468Y210cd3+nkkxUHRovcNh9LlbAn4uDal9uOLzNynfzUCwT
EsAv6cYQTM3jX56EvAHQfu+/qtUHM36KQOLmoyCFEye9CTO6gdXrsU2GoSjjpVuyqEaGYMRo1G24
kaap6mgcvj0bwiPXeT4dMoy8IDsddXhSx6EVsushx/lTXslgHxeaRNeg/BKZHH6qFJlQOjnli5QT
jfS+qx3PKhC4PVCUz9w+0TJgfmxUeV7kexno8rRHdO0BCgQDh2tqP7lnAugNiDl+eyNtdOAiXig/
ni1s1L0eHDbGp8W8piZkz2miWJfraFtcUUg/ixLpuNnAy02weTuN7pWlEeHD1PNQ+O7ReQw7khes
0XbwqndFLbk+Cob2wGE27/il3YLC257N+OuJz3j995Q8qisZwqU0uN+w3cWtZ4CGQj9DQH1gHkYB
WyreSNOnNVO40wzWb86inyi/fIqhj+aYAbk/VRMVus3sOToggkyjv1YXxxFpXXUR4yJ3zFP2rNjY
5iyxKSxNoSPbN1uBFfh+u43+66jdm7RI//IR3aDIxEagGeWdxEnZtpIf0ZHSbzH0MLwztmUw2LDj
x8rXcamPMBj8RgVAryOGv+UnkG7vDpMVU/Wu8CQBILoqf7aKe5PfCd+nzo/XygEsgdcbqhMsfxNl
ebigGWyoQVL8uNN8851YjRJen5VwgATnRIfEedJ1a1oRbAd96fAu1Ycj2jU46KJtJIUkdm1cgDKD
/4jaxnK7dmRYi5DQLIysh8tuJoBQKHyQDId64WZpOX8xkm06kby1VAC3rJUy7nYo8sKAIrh1LYcz
tgp6uqvUlprQWUYUzoM3iKW4jCgf8rjvr455e+Ua2RXmtkbI0bsyz5TldS6JT7dHyrQmEeEXt+A/
abKIpKC2bKpXNQkb5MuztN9To3E5xVBSrBHcjMTM2b4g7rmpG0YCVljI2HGK5EZU+rTsRomn5Hfx
6Er9aqwDE80j4qxjg/57WaZCH837HdTb1qLEd04KrfSG2Uavp9t6T8ERdXG57ypmcnJdFjfkfCWS
WQOZyJMKt/jwGgPg45ex4athmEvqWXeCVUlCBgt/Hh3tG4Exq4SrIAUruqTGVhM6aC2t5Z96wj1z
KqSMVA+5kbUNFun716x+XM+HHoE2zhe7s8pzv8HoweQOSNHOv+U1w3DmNCH9zNMXUlyUhU7Y7t1j
QJtQCbJHdlzcD6ycoJGQGtuZ78Sk0uuwcpk0YMFUxQNDJyEEhe195XLx2wi4NUVB4gSyc3hIuwpP
/XQHMqQkt6QGugiiQf3xilUE9PHkC7dbXhNudO+QxmzNekmPtc4wAYwv8dRrdcmrv4c8ORAJYXWW
n/FDXnDWlX+WqIzeBvFyoLtTsxaeY8jsTBUmZ6mW4IC64w00CZhutx2m+mx30zBYeMxs6SKJI+T4
5DnQVsbY1SZ2mU/hwsq+cN/UQTwfNVkZ7RMumUTLGNiTf5z+qgZwTnefbGjqQMrxP+UD7uUj+2cE
f8rcx1hefkL4UGYLOoRT4CCVc0MLpXbM4Gn/hH4uHNdZOXi6VYmQm1Br58Hoz67H1we21pkaaLhC
1c5cS6B95FjSFJzKGd1ygufvVngyweE6P1+DfF2MTPw9HZIRtcVLEejGd4LDKcQoOpi/qjm9WcYo
a1xkrrnOPiq6g9Po2y23LlXDYU2Xx97wCbBaC+srUt7+oGoJyeRicBa49ooqeTgGSHJOLaK4nlwF
I8KsZJqHB3TFByb1RTE2vN145mwHfjqPUTbj6h9olwpRhhhaSzhEmxbY/Uyxe6UrxKcoE4TVpSi+
mqUoc3prunKOWOcYgQx1/85drJTviuqC+VYmZxh9g+jiUIx8/6IFTSoQAByHJnoZ7F+mi/JYIj8j
a8XW45suuRuZ7WRnQTqPkGFBGYVrDhpFkDzQSqIK6XPyqyvZnn8+E/hmlQiHEcVS82srUG3cYSfP
iqc+Irv02Ep3OUFdq+Xgk5x2CWJJahKhu25K7Mmle35IjGJT7xi5VQnluvTQk24TuCWynvtHKmj9
zLcZMTN4sudHDtrkFXEttebQKKzBPwP10N07jnbhkzd15zyKS7eOcrmESuXyegezSVdq8Uhpe22I
yUXmL9W8YwnTvmzuockPRnxNzrsedLl/ErC2rqjsgWq+1hPXAM1StkHZhd+IpsqlPj/M6MNxYCLW
PFoUUP7YzMZcFu2I/+E9CeoRQOsPXsa58HUIaKstXJWbM0BkGiVVG8ZAloI9eqqA+t9nN89eWTRx
46rer3O72HLxUdNJM2b92PS586vh3Yh4eR1u/DpqGG0g93uXPaJEcck6cjnK3UX2d80PymqhGmwt
cbuHhFm75RTRHzQoKtpeB0qoFhA7UgeVxE6kJW2JdStHOaQOP4kBmyBGS0NNc9ApkVTtBKGtAXLH
LlVBFnEOqgz4gxd9PULabwkh7TMbBkqgh/o0d6OA02udh4FEt02lisT+S4AP/kJ4maIvtXC1C+ZK
zEbM+zi/6HkaER7/1VE3f1/U9mTY4qsYi/haE4Zeoy2vSihAkdkTHvTNh7Vz5A86MEvW9rpbJHee
oY3fbAX+Dr98m0135u5y7W4QOCch7jDL6Krr5rsYXLBE+xBlMsT5v/HKxyMclSDpWgqpbKq+lqNc
GYBiLeeKruMPwmOAlrTgxiTvck4d2xr5JYch9bqvSf0vBFoUldF/6Cz9Wf1R9UplxIOmQMtAX1Py
ByrOUUGs5MVAQHP+lpG4SiWWIx8hUT8v3LzGbMeAhOVAMwImXbskAj3rFk/TskX66JJ/tg3lf5Q9
F06xQE32/6DN0Y/LOeveSIp6Xy0DPfaCB6X2kf9Tj+kJBcFwjCjmN3r2ub0ZWRFkzXe/RXVtT7MD
M39bNworVz5kE9ABS8hfyvciuYWnnaREtjO4oAZ+Ud+QhqGPu1Yu1meSt44wm1Z5l7QOMGZjs4yU
x3J4N/e1bL50Tq95nsAmhWepVYuhNDDALSSk1rcG35Eu9IKXVWKVfGJcTvUAqEAVBp04a5vsCh3V
Dd+3Lrd3yqLnKT8eNr8rHQ4A7NQrW7zLPK7hKBFBkMvH6eoxyC34JCdU4aGnkWhBbctGdy52EDgS
RdzW++G5NsWsboidaVnasV/tk4Uane/wKs5V/Ow2PD+DdUPOm4k8OuOh8E0nCft/VTGt5s9TgDkH
0oTRWaFvFdS7nhTwOzHq2+8WDeGjRCVPDSnIRqJeWhnce+2tnaZPkVrtE0Qq5kYber8dLqyFWIB9
BMSlX3R+1UOQXmnJyCZXg0jXSylPdejDaNQ5zoNnugyCcZf6Ut7xIL3ItfQ2/9xVtQYbSPzz6Hpq
LSLxkeqvuLL4FqA38iQ6p5GePIYQGEp/7Pe67OF+jJrPHZQk+m236H9nkHqjrH+c6UVoYtS7gxhz
TxNHo6HvKo1xqkkmAsyM1g5liX8qQ0oRA4lTaFhRwS4baG95LZtanRc7UJdGZz6svzfBhg+WuVAJ
6XUCt5s3pnSXy0ZqkaF2WP11Dz+FGuN2O62mruXwt8Vb6rYHzDcoGGop+7/NBmzZ2qBEJ6O++q0a
ThtQHrdRKUhIARR0n3J/dJ/QP0AKNHhpSxd2yDrr0+LrNraXV0I6hYiVP3F43xqPyPv2GbNVb7nJ
AgGLo7n3QTh2TSXGy1mwGWywctCK9U6mlxK6zki85Yd5Q9L0JpdX6JYkpTXOOk2eC4M+GxSIZvgI
7S/afHfHszRuYGakVVfN44Ujy37ssXYGDpemEaB440Kvfd5PpMZx299DGhMn33fdG5GKE3Jhlez8
AZZQ06uneno+2FPNx1zkf+KO//UWRc+3U3cKxKwy+RBaplAce7IBDDxG5iK+Mlm7sR34vizXEgN4
qz8oXtdLH3jIWCRm8HBw/G4wU/wNvDAsXpL88Y51CjiDhD3oyLk5dS9zZGMoirMMvGg32xFqrCQ4
jnp/qxk1Fu3z296UcN2JAxrqlN/TfbI0PzlF44+jPSVbnLR64sV8BxZYlwJRDYYZXLU1ar/xH1uU
BYEsKE9rsUhOAyQUEgHKd6v4PiwPvh0iIqZGJatn6cf+1pnwwXVK1q0j3n65hW0YcY5yoIMyvXnt
QHufAkS6ShYeIWS/m9TWgVFK/gfkWF3C9jVm2wlFNKEEmQLgc2zMnd+FbXFEB3tMWm8c78jMdC4A
oTkzZMNCmAKbS8wdj2CTExlVAkYc0MWi1MizLgh7N1Z1LvZHOfnNeiGhKtOTDvISje9b65Il53hw
3Y5WHLXOOBZAP8S8vsbxTLW/CmGvF063NqxQoF+QcnmO059llY3K5Ez7iiXA51Pnv7cKFs9tfLM6
HGIRrhR3qJqeAAESCvRuXqEzUBpQJknh3BjuV8ee0iojXSQHiJwhKM5y+pDkdlRy67kp99qBS5yF
+6E71jXgjvBz89SKiOmpwuJamtS/4v9Can+ByhvgnNDQ0vrtd7lFIrgDgW/KVWhVVzO4262Ys55C
hLbGrsP7frSnWMsDwMwDL9iFfwrXsEv4YJyyTFS8dcd87R/q4c70N2g9tGOsV4wY6baHYcE31iQH
bLWjrKybzZvyJPYySTAuK4cY5tjbsyYVDNZP2K10rH6q2qrZ4Fi/uCia/kt04cRXLENcPUAIlf3f
FvO5eeFEVrFxUUNsewN9mLV1+27bLyIrTem+aN6P6GPsjZpaahnd9mnf3Lku/H65Yf72fZAleKYN
F0DenBHoiCbIq2ymCJZapLn2ymtR1YWSzsusvpFia94u+MEl1/O0MvPiS6rHsvi9BMUorP22iU9T
OOYJF9/J/w4W1fRcJJKuC3q4uVW2R4aG2D/6ZlD2hHwvm0Zg3xq67Xz3GV5DR9j9Ahkx7fvrDeFp
S0UXwNQAJYmZw1ROA0va8MKlBb4vtHvHSZMZkpkyXEDcDY6q5W6h9Kt7M0moNC0OZTwI1vfSqfQl
PDO4taORrb8c24rTkPKglSLqI61NcWPbdjmJ2FOaj7dtNjTJK3EytBaX04cqrgoNOs0YErlUmt0G
hWZhDVieYVWLemoAYem50XxEGzbdxn7JnVsprH7KNGW8EQkr88GIrdMzIsgpQ1FXuwPQlHdrzwQt
YS1/IamVbdlj3pudQXS/vSmqj2x5ss+/ICrxMaxzsivyD6q5ZnA1wkvDeHJucvmokhhxm7oFtzT9
ImuiHNUDwAL1K8z5bkZukD1VaIA4J7LrhRF6KZ9ex8AfI9LVvwrPGom9JaqYHFUZ0imzQksjKwzy
fDMUO4KfBHi5VQCJCC9WUPzCgDMT9/VgGpPfXCFep8dqTQEV2pepvGKNsqyPj+6X7RDeLZINk3G0
9Ri47AiDpUPM9y71CYop8Wy9OXhW5yy+xP29VMK5NbEaNwxoNfPCBt7+ImHfZMfpviqy5LjxMsmv
V5dpQDKdfb8lAjPxjAMrM6Cytor1zFrxjR8QW0ZTS0GEL6VLUkgIIGcvsQo7qEVu+BtfxV/+cLjF
tjZZqu0zBLkMDJIpZng6N45CWW5EGroCaUbZlC23YSkaEJgi7h1vL1oRx3OVPXww/g7rv2YNhb34
zGfrByzZ5a7GDmtrcWeVtNWxM60a281v/peTD5GO84NfHZTiNOdLlqstIs8ndd4mqZ/6x3qgRW+I
Ttb9+bofl8U1KcjKW2Xzo+QyDoVClht0ZeK+FpNCVXtaUp7NyIXpQpKvpj30281yf7CMiy5KedqI
Dwryu+G1ZdUd+ZiphX+hhzElM6GbxGZRO6V1HOEg4Z/LSX0xU4KiVROTTrRu6AV6GOZugS8+Qghv
6FYBVV2ywiYPPHLW7HWCDNJglhsCElYg+kSQjf+ogMKJK9ILZqem42ZPLROXhG5/K8izldeLh9zB
s72Fd00lRZ54FaPJOOBOiUbw0UxVlbUWSHKwjYUNu/ZD+8JYpQ3VI9YH8B5V5vp6XnCGLdF4EMvU
8Izj/qVFv8GXEGz8FvPFDkuGWM4oPsr77mTenO0/Rz4IUCSQHRTIKU7r9cGG62JdQRoHkMOcg+JH
JyXilNSVtRRKXrOfhQZgUp/ph3rYa23vD0NevloZN3SYqA8+1RtHLRzJVVjUNjYBjUtohOg+FsQy
ZbqCTrQ4S37K/trLC/dwgvH1c39K1HZsfqt3cbJxMlBoi/pammDoBRoUeFkayP4lGZkNddmm2xEq
p52Dxdm2ouvE1lytpc1nhuTem9HOsbH5OGRV0/NGFaJtgbRP7u3ji5e6SfJDaAW+gW/8d32eX3Uo
SbTDXQl9iDi75uv3gjN8xRw4kp+LcCE7E5jp+mWZ7UbJfSOmTARIHv9ohySUL6gff2tvGVO9hlga
Xo7NFobnPs/xY8KK2WrKTf/SqWAKOhuoTr4ccz+pKuEfoJXm+mFIrqqu8qHyyylHliqRq070qxYN
5Mgm8CF/l3wJ3GmSLs6WxOjNYO/AMevTl8Fv/+BOX/t50aMIPJSI+LFADDg5rqN7Ls4TmX+8h3Lr
XCaRnE0TN1UA/pecwleyBAw+Cdeo0Qdv/3udtmycii5deryS9Usloi0f9UpJes+YgLvXzEI5JQv5
91JZpXNmr49nqvCfiH0fVaw5ituXe1uRBShibpiLswe690NWjYAQS+DyiQqGfKCebcL7QPCISUjQ
KcDeiLgMoXfeGYve7C/H3DwfjUqM4mYF8gNFGY1OFQMmXaqHsJUI3fdLrOdx3KEBAjfyF4h+TGZg
+CV6eevNVzX4Tiq3gNqaOT8AVo+ppRHeWfhxsk7FFVEFpeWVrQEmMXW77fyTSkdXw+XgziJcMtQA
6oDOLZZBE7AYYRyhPiun1Q906L649Dbv7UwaJl00lroAmou2Kp5LTg5WDi2udFfu6F1irVT5qcns
+zF+o9iDHvjhPITvz2nORhgYS/dQIRcw0X3PLIbzOCDOoyhv/5uk2+/APml9aNULw+/QgXKelXcW
qh12AmervJ56Pat3QPwymBamAadoyzEG+Ta6emOTenmoxYoYEcDdpUBwHmVEoWmWCCJCQzxOqFUI
BSXZPRwOUeEMTGutU4DxV0uogI9pDew3LDzvFLxeiTU5nuRh7pPcEuID2hl43FOjqzLh6LK6i3Ru
65gsD4GYTBU03I30FheWnMNVfhFmmf+7gzJxayO5uzwtvTenwzRyT383J8yOCvkzCn9cJtqtDq9v
+jDtwWEl5SmTyvX6WD0quxce1MpPTGhwGlIbKulo/VPfZhbIBngtZq5QvG5OEiGk4Alw3xpW1fwH
wDdOaB+4T4Ny+A05bVDxHAk4Yx6MS5p8BC6boJQ12ETOV/Wks0qFkYIrTU1vMxse9XIsnshC6CwB
uC8+a5w+kviV0YY/i2w0uu2HgqrDVb5Y3zTu2vwPlyoaL5LZKfPk+4hRAz3KbE9b22KispN51YOx
K9AWBxEO9zIbJOe259ecs4Xr9CwjyJaiQEjqR9fYbhLXXYJUV/fdG1zQ6RVRYYzgDvr7WulEYgR8
kveVC+0WTtppTxcZDbBYGYULmf3+sTewRc4qV/Oy4hLsaV7/ngX5Fq5kz0DVinXzQS12MhIIKNer
MGlryP/Bg6O5+8KZIK5ia7jMRpEd4hVtNo6C7SaFe1IlGD/99Q4jRaL0Ywb07PL+4bQTMlpLw3PR
nAOlVV5EY7Dwzlyu5ih8b5lbDVBt7Jiaad/gXN6sUq4KL3G81dnUhhdgoEATAveMrQWlpx2ivJd3
KoyFgigxAYbUWJYGtIqqv2dtZiWXiLuNijmfWN+E8pNdkULYP/yk01f8qy6plXN1EPLPufbJS0E2
KuUVergdXA16CGjZx6iIDxKT63zV9It+haeD7JDzMqVgKaL1SycSXOvEkYlkRBTw4ailtPEm8lrI
//Q0mwJHvNgcQUz+hI0L7v9NsvmKG+Gb2ukEcRIYZLrBmlsHn4QuVS5PZiq/TJOhDOPX9Y0ojgeG
f2coNvngFgr4TmA05Vgx4lPCg58jJQiqBUA07eJxXquyjXyrMPEmkB22SzZkLw8R6DDcxxmZc1Jl
KQxQcPfBrTwt1jQzEikw1NKrmqyLz3CJ9F+/TD/UnExfH4g8QMiJVxL7Y/jjxIvZmSX1hCf7rTay
X//Ft1CEM4Vg4SJhfU58725/+pCHyJJfnDRB87uXtt/BNT+1M/nbWk+aeCTlKyhfanhQ/jcGZUiK
iGcb0gAcMI34CeSstR5bgnWBC3io2u7MxIod8T7IT9GxB/bBsIEgB4FHp+msvSVtscXPuOl7R6bz
h5OVs8JNsdQryH2QiXK19FHnxMx3Cw49KnQ26lTN1IAGxeFWi+SK53XwCWn+c4s+evvephDUnuF1
6lL0AqzvL7dk8bTQQK5uHWdbTTB9a8mjrVsjuLB2kQiMh0QuQVwu8i+NuFn3v4H3I22ZG03EqTUk
kSO0vzxw8OWpDtrlfFRh7fODLfWOXEALMY7D5alkEbVyEYCioBystZ7+cRqACy4PUtI7ZZLd6PdJ
hy7sMccelfBCf1rFhbo6oKF5x68bjLaYpXZoiz/NnfJnDHh4HBfak9SinlMcfNDxejgcx/FIBRIE
G5vER9qYHW8CFRh862rgfPc9Y9miT7gXuIPBt2qlOE+pzRBmAavEDz1na4w7pi5fEZn+tqzeLimb
fNHIJ6rP8nwHfcGBd8uID/qB66iN7ws9RnhaLPci1VCqTqT4UYrMcP/3SHVk+aaQVK1U/CY5DiS+
rXkIIvh86BDnF1sCP2ksF7c+kDPlBTFEg3Z7v1X8bVYurE3Sbm467On6hCWNAx9rDM31awKe+JtF
7gFyH1M1nRJ+uUa7Av27CDoqb+wFeFvjD7yO3oekuCvja9Q7VtRUW9Jj/R15D4nD9pexKhl7Wdz1
YEsvPHLU18OOky/NIxz7lVLt3GqbWUItI+BDe/ujlJbWOWqzeJSVRFLIu78McD8HmpXHsaMQABlD
SnI7CtF+CA99xLDyQDMVUf8pam9cmn79lYV29WysHM1kfPh5E3XYwc3FjHcHmvRIWqYvW3lp6iW0
LkqFWPzxUZ12ZpgByKCjlTYgH0UttR6rUnVgY6EVkxgi0kh7IFGjYijyuxduqVampJEIIfg2IAhc
llUoiACPFIgBEtsRrIyGanLbLtF3iKQ0s3p/dcMGKOT5k6tucGdebwAvYyUXV9r0jSZO3Md0P2lg
qIXIaN9cqU23nfIORkj0P0dVT2Nm6lwi2n96O8HRiC2QJUbmfqQFdi+h/jMTROfr0VNSBNz1z515
k/5s6a+/mlU6uLAT2+jEOBMI1YIXtqfqXXPzPwpjfcRf2hzbcwRQFauFZ3++kpVfgDsLZXfVRD94
V5a50mH+6sWI5dLJ/THa31ojjCYROT1SKbR7WS0hWrWo5khvJwSyVJ4+i5tMcUWNLS8ZjXyN9PpH
vQ2hrw6rTxKL3Z2Pw70bJCDz0h8llULcBeUSqEd7m/A0YDvzjt9tTL+aaumSm/9nkpg0hpcRtOq7
foXTagf/6uSRhyW97fvsxYPqpeIfLEWToLfMyJDV431fCojSzVbW3eLuPUFfpBoB+76LJYmu70mn
W1vJSbldFy/4jrFQARnNZ8HUQCAeDdz22WWhhl0xxZdHoV4TqDV0Q3XhI1vWD6svRuu98Hkv59sO
vrbW6/X2AcD0RUw95S0rSleMo8iHnHzlAUoDHH8/VsZes+BkIMLTvcduVnB8XS7NIs43kCxTK+iu
8ro5SIFSal0J6r/+xMhIO2EYO6yAGGbSVnDA5tkd9EmB/xWo1NH7r3y3NpUiUO/VSfwzdX7k/PpM
y7z5prfvf+K8lFunPoFFxJjWjpnJc11380dBEHNyUcVvEUFzE5z4bQqBqM3tBmf8ifzcsCejj6dx
gid/A7X0tyGviUCgFxOSW2107c3MVgdzG09dJNPLew3FcX4rnPCB0t6+gNhOHO8bRNoCE6XdoN8O
G2VmOTvbfFnlAhPsKsZI1VrYni/REvNXKfsqRDt+rO40g1MlrREAK53ojdGb/dy6JnZZy7GNppMm
JYU711xBF9dqmy/xxW0r3dkdp/tSRKXFoP8oOmFrGVs+vYZ/6L90Uz5DROMLKXzyLb/mRlCl0m4/
BbFmuQRDyABmOOkqS6c14igMixGyJPN6RSclHV5X5klVmVIa/gXpQSLofjEMgt+rCE9jFgNAetWN
mP4ooFccDLWhO7cCNQec2+/c2rGdk5BhII7ndxhoYHIkqlc2n/7tNEM4V+E8etcMEIubnznSLM3M
hTYgjwdvRCD48WGlXl6k3UTKyOaicFkCW4/cIdFibxmALpBD4x34cujiPws4KDUvhN5HjQvoo5Mk
uXaJb89To2pmqCxAbtesntvxjRPnm4QF1Higpo3YuVydEUvczqJ0XN/GiGmJKy+csRqlrkTbr521
gEWXE+7cZmQfD1t/dPcCFTzonkCkHfpfsoZzVlwCONmuLV5RnVGZJP1ATM9AsFqpBbs8Hcr+gLPW
l/FR9kpfeJXeJV2Ff3LFzBLmc3LdpdHoeLSCP3AhsEJ1PU9YYWTx8XUOMtE5ifzNlkqhRW1jVN+I
OO1hUoVJMoyH3krfmxa6fGZZ1JKzjWAMNnRF4mRfzbBTq221sFgzEwI7mCMDCpFBzsnYuvoLIiyi
IlRyxwE89kMcP/ndvjhJdVp31biTKbsJV03Y5wE1b9UfIPPZE5RGQX00qORf0nJ1jZuKSDk6J5WA
4dRY5Gl6MQgdYWmEtwOPqgB/bcbRopZqY1ynN0cXRcu247ihILMSIolJwcb8fxEBXdkzkPDpBxu2
aQ1LhPJp7pOfA5Omqwea8HIyaSjQBhFo3k7gmgXKY8/sz+QnMc0QNXaYcVI+sdHDxdJ4jFcviKAg
C44YePlf1AAT+Wmj50SM9+Bf6iWdFafrAec5Xp+nwa5iuC6Uhs1Hb0ASgRerRZKXdp0IFEP5PqnN
WkaHKTObZETu8ZTS4mH7AHAWTB7vMyqdBSREwOtS6bnGXesBpeutnst8mW8u6zm0uQl9itLToazA
fWIGYJR7oGvp/ztrSUBERpi4XxyWUdMEPGe0s9ea6wfL57+VZLf2pqSPhAIQqjjrkNLaoEBrrFw4
PakHDgZpgMpuI1oMpI/+7AIZfGTa42X813yjL2ig3ptbHItk5LUeDfM0+3fQf/Uhr5gOBJ9KfBuK
M7FoN+ESKrqHAAGNKQ2A5glvNtoeS6c3c09Usc7EKMGLcYS4X2x7/gTYPxRMztA9pRU+x88P76Ht
35VXwh3lVgmDRxfCa2kPp7Ur9UT49fiKfY4mun7tLmD0LqN4NIcjKUfDyZ7LBZfIzwt+uwQrSIle
qhAjsRLtxFtxyarKotzvfv/ma5amGNEnhGDVXZCdwIRfigAu5kvu9luk+r4/sT3mJUVifDFgUH7z
PoVaFN4I272XT+DceP8IoH48WQAgG2/4nttFE8BexWymVPJ4GDODRBKK6hG7XUpouQEqR5Bd69nw
MeTHz5J+Z0K/0K4mY+iOlOOI2QCbbbMeO9xv56VzGZ0JZ26FS89lQuZFbR6kU5RPVd9aGZA+idqT
xxkpsACjIcOMOnbpBJjO1U4k2Cfn34uflXFR/C3yKf4fxJ0UFvuPkEyBFi6eJqkay9RVlmNNxoUA
QJJvqxXGi9kAZ0yctPQTmmA5LA/Mqfz061m9qC4RQbGXDpoZaK77dRSOVTXTiCA3mAQt3aqbTCI6
Kd9ix32dBQOzfA5vGtAlqkB4eyRNnhGpmh8OB5ChKQl2qvPbymmu4Cf2aT3q7wvSg8qGrnfMrzk9
IhWNKRTJ0vePSHFyb/QySC5eLz6UL0ldaqvE4APaQU5cwAf0+HMDGDILyGd+kBAigzSAyiWDvOQ9
JfrjkhNTxEzG63fr2z5NM3mTSglZzxjhK6jEdT7XZC5h/dmppGfh/lM1u5cmswQf39g5CWfox4wN
Fx2KTrOCWPn46CHmEvGc7f39E+7FU9dfZUeg0Ksm+7E40thgV4A6JzewGV6+aJu3oOSRutWhQJdp
+tuFPhClW5qxF5XwPUnlp55MTTtb7LfGir7Ac8+erF8G4pSpsOfSVgdSr+jHYVKT90O87Lnbww4P
OoRAa/8d2Vi97gkvlWj9bB0L1+luIs8z7GeTy0virj5RRX7ZR/FHiBdsoTZVt+HpPm9Qwo0dosfM
Ao+LTic3/NfUXKbdOk1SfRGk6JCGLi8Ux+wF+Ua3r0znprxKZnLqgNCw9JlzQVqm8UMz84CNNy5X
FpAq/5qUXZwTyegVGypAVckTdUFeIHYuJ4JClWHjQmD1Ghq3InPzHkPTKdNcSHwA2N3pvmhCLb+Q
/3TzdmuH1cfPsJptG0J+yfopIqtWQmPk6kT4FoyKXqZvHS/LWAaLElgVS1TbZNBe5/v4FbEEBtGW
n/0RkTJk6+lWMM+SM2W813zT2SvKXVCboSBeKM2J+mT1WiCGTkUF++l/4L/H7gkFoyFGseeln0aS
dtI5pxyb0yd7+OxO8814+ep0hFT14zxwJh/fRgGI/5oPJKDkRF5+kmzLhtoJjSDX6zx+HKeqlmfF
+t0JAiNw/HfqDbnVhXhGx8yzXR5zonHIu4w40mSVfJNfn07wiQigoxG254NEsOpudwjCjc3+ovPf
ZiaVvj1OB+WHESd7BBl1lieX5W2u83QOJwzvMVIuIVAV1F8XVWcgdusmKtAsa1bByOenSJFmw0bd
Npa3zp19ijMSPEEdPMg2gQP6PtN3phX7Pq2A+ZuLrEbXj4Qg4/4s3L8eQGgcj/nuQ0gmaywTDKoO
nT7W84WcG2WFXjMPjsMBht5sU8CXIt2CHBei46hnIClRzcgaUYZX2lzbjMefc79Iz7BKB51Um87h
G0VFqgta8QGp6DOKTu+u2kTwufHp5JWQRZPcMsbYr+vpm3I2SGOcXF6Mkwoo2KtJ/jwiQMwIIWIy
93qiwLAzngwx25zvsXZVB+JJKeHR0oXOdNMabKduEII0EtuCBgzb22hFMRPXtpzj6iM/aJKFCx0P
EWHNo2u7wSxoKA+VVrtfk1ErogTeBI1IAhmXmdewhnzaq/2gwRhSPPE8S1SFg06GJ+S2hc0i4t0n
1DdsiCzMbpN8baauZiwWIPzQfZUIcaTxWBWgBUBP9zmhKELO8P8etUfhYYTpqsTbp9rVz2nOAqdH
VKWhjjFBgI4NURrXhdfZXNUt3Absj6Jx93hgiPU906WF6FfzNN0iHr2kLdGKUDfxb3HJWyEhLqsg
CNC+rk9s+N6YCo/NckKs2hPOPBthjYAJBjYykGgGPMnyBBU1RNjtsm0aniV65eFfWm3DPgsotwBi
v6vwUFxKuhhXP7ELSDEQDUbyJkMVQZn+TxH+/t06bdLjsQWG6c6+hLQ3rnXmNShsyA9F0x6ArPBU
kbR8hXNto362zfce0EQbnCZUP9eYp1gSczb75pW3/NMEU2GyE1hPsOjtreg6QPwxBsIq0TaBUObM
2DEspe8nITpldB41/Ya2Q2LJllmgIyfg7lWo6oQ8E0dfBkZb5oFzq7M0BYGlxPtGJ41wLSIuetAn
hFLpwmIXLGNY2yv6o4wSCixk98Q8qDhRlPCI2WTZGBCzSBu8FFGQ2ec77dLxm4NC/7Pm8sSABpQ+
Ro8AFroHVktFqSbXmPgHogC9S0ys5hynsWZ6BAblR3SJVWoS4thxKl2xpT/wGSUCxDfD4PoLcEC2
BgVFuASxlUdS9r7B5AL2zpI4vu0wRZ+6jAGhmWhS4i9pCwd6N+COSZZ1oRj66luTWkpkK2/bkYaT
EpsbGzZmxOQA+7DYTf6/pylbBnbPCyMEkNyKUStKSRtMxwB6GsTTIuVGA5PgMk8Osx+9kVOr6rF8
kuX290qyVi9X24Ln3Z/OpXrglrhAA+pn1qMfhsOot5ZhJrYW/aulVZCPIejlWht42JDhN3C2j/Yz
joYJU98R4O18UNkR2g47EIz7BNLYogSJjVRMU1PqyjhK0kvMmxoDhSbO26vcw6zj21LHF/czVxvU
v6xbnQvJvq6bIOEgQP9vG50BpupsNFtrOIid0CrvqCZ8ZmO9bBvHI0iZde7U+6MBW0zpu5t0mgK+
xV4czxzzUYDbyp3RzT0G1170S/NKcFYCe9bTk3OFerw6XAsDPXGb/be6BN2IiYZ+m9HygL5tCFef
uNgyOlJMwFsXkduh/kpZBglDj1WjufiMTLBveUnH/OSDrXPdeph78QePF7noddMw0E9He/E8YefS
ax2Vm39AN3E2/KaW/Ybq8andqKS6sDLBDfnio+EoCV9Pxu8tW8K2+fdBClJbi5KGx6N82LWiw89y
jlnX6XKwyiNump31RqfKakj+wbJe6IIeYIXbgmt7XTdebXD7Qa/fkqRUtwuvUzNu08JDuCVJy6J7
qbfq7Grp1PckEBOp9IgBosgOo2sojGf1JnE8Gd22stQcmxibNk14OmYJ30yyeKoz5BUcCQ7gWWmV
b5m2DfiiYbsBcqhwjSC9eJcRkF0t6bKNvIGrj79xzBY/o/MUMlMswEbOSVAuGpLF8FmZ/A0ysqRW
LoQZyW0X6ay93sfrUmVF6+L/BuNFJ1iUx24JtvNYXGtRAfKm0C45tRKGzxeJzrlCTsnJg99bJKl6
/r59MHp/5n7ja4Ig6UvNbPWvSXF8vzEt3Xe5ai85PK5pf0VjCKZRN+ihVnrDXbci50QV67ZR19e+
JVw+7/7s8Pp+phRgG1QfIjc8+63syU3ZI3RlsBSiv1RoSwBERKC7qZH5DaUicC5N9K5bznakSo3K
BbA3TpSAlBEqetzZIhnzFAC5DxikDDYbwV+WCpAypQaRbGcIu4DGh8GFJg6wN51QEIQL3xD7tTp2
CdyXyCYH/m4ccly/Eh2ENEKvyuBE0en3Ua/p96p5ueDHzosoJEj3zt1gUicscXxIqgQzdUrui0s3
qmXhi+vsfOkmXIy+ZcwWAbk4UITzgOXN8erPrWvKCyUa63Jcaw+fuYAwjEybFkKeg5hWDKIvpN+t
qVhGpHRiHIt0YnPQZbG4cpLfzwhqaGIQsoiqkANvftdqlFWJzOIOkOSRO38Wf1vVDsnfqg0uEeFH
+E4YGM94+P9KbLs3NTpTGHGFMy5nt0eKDcrpBPU2FEqXiQ8UN/Q18kElF6pFD8j+2BkpyoyCgK5N
oqP24XzZGXScZV/tLxyiKDrlA8UN3jedSgH/Jyz8jERqtlBTgZ/MeWKVZet0oszEFPGvjKD5g2NI
VwIWfIU19f15HO7/5y+DRumjWWrwmiQoc12UMWZI6nkJe/RBONt4JZr7Cr5kF+ZyiPXYmpH+Azga
iBOyQu1vffQ/KYy8JWgKHEV0WjnuW+OL8QxGkWkhFPAbbdf4uIbKPdY2/82lc58EVg/tUKbIPS+G
5fbWbNNJu9Rz2RiEECp7qnzxGctWVTdXdt5wggmmBifioiB/ryvVqVChVtl4e224ow+DGEGoK9Em
VmsWFiDiYq44zP2FC3bbBJx1i6kq2kFHJDXWDzD42L8CIeg9HDakIYvtO8MtgDPc3wmjAo3WlrPN
mxI47gN09uzPQB+yh3TfO1xBbwz3K55KRzP8/s6peZbGA+yUkmiBzRYYj1K+Ndbaair5gAIiQ+10
VFeLzjxKYpp58IdTXUEU2MUD+u9qGrMk4RQxsqL2JVNGBEXZdaJqC5ZcxmLTkgXslSzx++xZ85Fn
6h1JVCTnxMN/bHaMMXsihj1Eni8KV4uRIcPZmjE5v5VCT2jINecyIkEQnqD+1z8JsknveXHUV7vu
3ci9n9m5nvcQjVHpeQiXq/YuYtP/8OMQ8RsjH5nKk5E9XiSoCgk5nTEpiRWYxMxY/Klziu7OB0qm
D+ApdOt5PzlKl9j8CCSiUlTKxbVVgGDIaFJWcXtaxp02TPNX1RCRXfx7M1znktqh1BhmqpLVMA8Y
QmuJ74FpGklyoNPXSrQuLS4R1EkQRXegMPjVIBQfbWMpFpp/QUGHfcBaFtPKxezQtsgkiw3fNmTP
rrosowsvvoTKFVocQUkjqCXMioT7yNK2qWBWvP0K8YYEaDNTC6aoLMC29nXzUICMiGycEl08VLXK
bsYKO3Eb2WLunBl0AN+wKI9XmGA8p4F92J8MLKn5+UFD5fghnQfzqSSAN6KzN4dF31/B7z4ag6AL
CYmRSzgXH3F2F3bgI94eBeTiSCorvaztG0Nj7kNMPePJCDtq8jCmkNYHafuV46RYWYqIUwOx8bqt
tj+cDbGP4chAWMqg5gRi1cBteAV0hkRggaFJxR/c07zTCTfT7GAMW3ByFj7RH+ISVGNT3SkKz2v+
J70rjTUFhQdOZ3ZB68N76eLiKZ05vfT990zt+KgfcHzymzMzYCjxc0rj7fHgt1yu1xJe0fBAirO0
3VsiT7Ow6Xgl9bxijBJjXRoLiGt6l7Gl5YEA/jXv+qN6NxuLwUWDDh4e1Y3OEsmCcRT7AnhXHqTL
kTO2LbRjeSnFv5dir6ItrxhMr6dn0bBJr64Bz9rOynHBcVyoXh2KZ8dS1W3NVTfRtlqno1cj5pxu
gR5FjudB7LLDe3i+yl0Y7f722OeWNSknaAuDg71zzbtHZLG0Ky+XPgwIjv/1kEdEUIFH8i4V7/qy
zk010VL1hZdPVJCtzwOje3IDC/5lHvP5FiaVaHHqqoeAYFG5wblg/vbu7Cmk6ZR1ULVf4ItzEuvi
YzpYkPwb4CqaWy0Djc/QrteBaJNtLua5zU7TL9bDWrtuaM5WH9CCTNvrsKU9/dFjQCySO7jxRmds
hZM1ajCNfCY4z/5Rs1aMpjWtY+oMmtSaQPkGr7E3496dHU2VF+Xl4rwHMZYylQ0bWWDO3OMfAniK
s3T4lWN3ZqU5n27ChUIClVBfLmhUMxw81iJbZE4J0uXrrrIYqpnLWdIqkSS9eWOn7SgwezJVTVlR
UeU3b990pygYop1mJObaGe3iYjsND6pcJhoeM9cTtC9Skv5dajEKclzFh6LX3b8Cl1EvUcd6x/S7
XWXhHLUIA7YD/XpTv+rSKPqQ8zYPLldmxiS/s4rMH40odOBAgajwdI2ZbmJ35/M2sHqwTYU3hTWK
cvwFu8N/jyL9ectqqVsVjyjygR/c3Lbx6rXQhGysls71l2YgMMeXY8+IZxZHtmYTQ3OeBQ+eE2/h
hHXE2oTx5LsqVdKi6WpfFIvk4xHwdRKyAqcwECDXSKgx4Q1E3XI1jFZGe5nyFDrJy8CAYFxRRAuL
IIUfWIO0vTpZDbNYqFdhLgO6IFNqcBTAOCmS7TNEpb/DNh078zqR//jG/tarVILYitcQri7pe8RS
/VQ/0sXvyp7x75rfhNX69bT9JJ4Gpwl3x7O/FdD6PRj7/QirxteiY+/Q5VNME7RXJG3aPv3pdWcA
U2lrE3kLtboeaaxGDPf6U5tziOfvwLmNaICUpr1tm/6aJmpB4mMF8Oopa8h1I/FsWNIdjN0x+j9/
25MUmCgNk4tvw9IyTl+MDB+oHMp+o8uKp8YvHUJ5J5keEoVPetvFxcZgciNTgriGWKcdewPkJWJ5
uQQM5IWgot6hNytWg/6H7hiPbam4LrLf/UObe615bVLqe2UJVugc2BgDFIoYVv54ly9HwVCYgIl/
1hGXcM2XAPTEZuPunDbl8WbEoiV6BbksSFRzo7BcY8RQDCqHo8b6RwBSOqIITeVEWmhMlgbanfXR
XdXamIkv0h34FjCdgNy7RnQU+/KdeJOFT9f+aG67Soop9gNEJ6tvuPqJ0wYrV9IZyNxTk1MR3SQT
jAVzwiN9pwS7tcQbGNOsq6K7/8mpSJCZFGYFsLv4RQAfh3jlfqOY7b2OnWeocWO6EN+33k8x5ohY
xv7xBRiSN8Y97/EHQWOWac6Ym1j08dO7B3RbFuKzGhKVPYGBpm3kYInP9TBjmAxo9mTWf9Es4Ep1
EnncjjnvXgwY9J65ugM69NiJgTT8+XvC+ifb0YK2zn4Q3FVDEukAOuwtzH1SFjwuLsgdjcaC6O9X
rhgDtc6T8H2a1WjBfdV7yhCCoOiJBKzZy1cuwbLuDEQguquUFv7eQ6sFRlYJsVGJoknv9f/qZI/7
4l0U45J5b6KOtpS48TNVpVfBulvlMueXLxR9FdPjYNJPcf+MdjpjjS70V7c4S8hlft+hm8rt1t5K
iaDmVFXTLxr7S6fbRt1DAxe+Ymempl29GXULzHZ6HMzVKKIqYDHt/01PoLi2yqNKnZSiPd2oQM10
zE35m6szxPqWpbfGyAYRhJMcc0NK5M7tNsrnWmtzblofqTDUgnVuSyTXAhRR5I/UuwxaDnrYErxe
EFYlzYySqzQk4rm0ZIT1Ys8hM8xCVlwbu5dFqKBqgWQSnh/rfN0hgB/EgxSkgWv/uaIDx5oGpFVi
cblYG04MwYL6tBaMm5ySWeaTgtu11bzSyjAs5wKgwg4UHB6nPqbcoqVUJfSaJFKdbD+crRQXc7iQ
7KJisLzHnFts2IWYE1jOH0nBMoaRrgdLBJYeWRyBTvec7xA7EBOs5R57cbW062SbHQd7nY9ikYSP
jqFhaXRQmxZ2hFcAw95a8hEVSj6xc37xQgwMlAOhem6QVnHr0HN8ATBtfjPGLpOXWsOPjSW7+COT
DmAgvQMZm/1Tfc/2bJc7WopOzx3b7VBOfilBf0yGm9/sRvstWfHtP9kvYVjeo5S4QDykIa8AUzKc
JOzp5dk/LTj1C7h0dVaRDLQE7Lz93hZEDaUFCp3hMtYSuRBG1C8mJIobSCuXGzYTm1sHui3sHsW8
r72h93/9RoYQpx3/SQtnOArJmUJZlPfWYk/hIGa8/eOfIgVFZO+70wALSoAWe1vYwfrAn15+VrG/
Pp86T1XWrkxENQDluWM3juOepbi5AfcDesjMScYr2n84makY5z7J145oA5+89o+SmMYImpt3/rXM
KvPWfzkRHoNKHowVeel92XHwy1/ogmFYCkXy5OZsQd2YQPa37Av3waM1+Mbxpn0c6p6NAlvwus8O
235+U7GzoyXjgEKZ0GoB8eEHS7gSo6+1YhO8QJt1hT5TK0fLR3z4Kek3/FAGNXn8d+P9LwaqwqZo
a2L+u9g1HpGCfsLdNTnNevbymywsHhCFxhNnEJDl6fD1/yxx/bPaNE8xOVmcCLCiOPw/iFqmGYVD
jWXIOlgO5TAhFYCmxN++F7CEnMcpfVe4Pt2Xr6sKmjddSj9OMViIazr04pTiOtMN0LEiXb6YuZDY
rQHVIhRgMEFBpVIyRxZqXSn+EVeT+C9b+B5WT0TL5S2bbMm0uhHK+CgU1oNquBUpyVj3NVUpHwsp
YIf17LnWoxocBO3SZK4fR/Ez+clinOtTr5c4XBZxrQvhE6kFnxshDrh5pmDDRyegS4WQY1yd3nww
u7K6qcqeLwcji4lM8O7giUUAp0IWPT2DBxtDbE/lR2wH+Khz0OWIUPtRc+6yI/UlqowPm2TXYTTU
aB8189Ec9SplSOfrxSmtbooQA9BbvzQktFPDIdvb+Y+0RZEcPVCIVHdrQarigoPPOs0lrPduWFf4
f+kZAp1qp5Chq3BjC77/WcXujFRUMr9dxCBAXvsGwLtWTTZSUSD2GbtyNXBzM4QDmB9gWYfCvxhY
n07jCXhn5YRQYjdxZB1y6By6Df6U35WNoL7ljk+7d10A9DCm+BJ/9XGbwg3wqrtJ25oXje02Rbn4
M1eWZeU/i9DLLEmBILGKKQoUDlJNCJb1QwTIsBZZmw2ArTXbxNhHT7fDibm6MlUrEbgIaYgrcC6B
yP0jUzDS6+VGxtItMZ+vIJAex2AQ8Y7C0Tab7AwtBMR8xNX1xOGsq2QLpj6WbSNucpATr/0shiXK
oIui62/HH3RdIBJSU/cKjNcCHNNgZvBTKpkgJrXVbFjkLV0FdP+TKeaqQEhG+WhtPEKCPMWBU/Vw
lPQWxy8hZhGUzrC2KAxxG/NKYjDEmPXM7jhMTXNqmu/WD0ZdfqcyzSHhHj315hounWScGWbqIhPR
bQ+uT+gxZJdmqpAjAP9x7KCJxGWccZg0aS7SLLbPXjNvxP+rsbrTlUSMLWHqviWwTuX6mUJWF4un
pS7RWWDtCP/W2yBOan0vfcKy1N4ic6Ovo+QC7QYQFjFXSF3H5skwCIoMSO+cP1eAKEiI1yXc1wGi
I5yRvYLDeDdFiXn216GNRqsN7+QT+w+z2nyNiO+hY5cq7PAqaINmIOEHZXvrhL4o05p7N5mYFZPR
cBx6yAhnTepTiMxaHGA6dRrOpMPIHFm2kKqoQsTvwdUICSDShihMxJ9L49OzQmk+DbJqXACyYUlE
X5wgGmThRFpPycq9ptjFY6qlZ+Li8fnTS3LzUntLboF7vL9myLwBDzRIrBwkByi2sE6rS+Ja+/2C
pE4mjyckMf7GGaWx04opuKZ4bOXOsJqUjKD/ocg74pDwsj3mLIQU1fL56T9Ym4Do5XnEcJbC0UFC
kFlf162u69qBRksCBo6j74diYkuUHAfXWlltejPmiKBUVfuh8j6Sei5EgfkmiGVHyNGj9pYnycNR
MVGU/kr7EsJ7eCv3dTUOX6qjPjMH3SUvC3/vfRGDpj+6yzXLPJBrpKpCD43PcZYwjb0MVCqgHTuZ
/SsGP6FYK+qsdlxhOBeRjZ4wo7WmsSUI3RJTOWwf8bJ9gFwuOvvvNdg1nlySX7Xo4RyPMMYb3MVr
ueSa2+SefD2aBEd12bmLYbs9FQ0F3jwI8JxDoqMIA/Df4aVSYbwvzlCKTvpLooV0qJGc6Hg/bNMS
G9V9GmTBP2K+UtNH71rkPV3LcIvbiXt2x8amg13brLEfR3Ta2cGPyuEazyMyfCvBrKklkETkS99J
81lShEUJkvrwrHkuk7pS/GnzeoseZ77/1SpgSfe2TLvTSGMX0aP+2xKfYp5++Rn8zpwX/0RuJ/xh
A97wtFcHl3A365Rv54oxkAxgNePSY5USbUuQ9iEy+XiJajhzudbw5x0jCOzOV8EamdsYL8Cd5ikQ
t9TT25gcD6u9pHtNB134aoLEryogAJw77dCqDHw/9cgBLh3ZxYekgKvLdRt4wuBBAn9ti0jxVdlQ
1z3c2VZ0ZzswDg181DhqKb70PriBX/AXDQPPb920ZVAsOqKa7QEsuFyQrx70I5vFTqTXP2kizt7c
cjKh/YcVtJLtVYa1Q4KwV9wJzCrb0CcYTAcABVZGDsyLM3HHJKIrb8xG4ts04eYl5i5bOPk2tIXW
HgfL+f762JZhsvSRb0D+WR5DdUqsACjQG0q4yF2n1LD3ABg1KO1m9wVJJZU/5stu969gI8On/XW0
qNLyD34qqQyAh4ZNEMsF0Op/AeXW1wBlJj2dvg6uVc5GERJmeIcPCoZlSZ+e4Ko61Bt6gkwCi2St
XEIUnLi5DoHPD4/OPzRMnPtw48B11vlRMx26cU4NJ97Fs9s4KprLNH3gCW9cfrpsCkI0vOG6BJec
4y6HCPeRybhlTX/5CovLR9eb9tiIcl81YDVEVCxmarC7iAViuJ9eibMtsCqxW/IhGTakP1jZUAzP
CPuRubYjSAAf2hfOlADh1H+L98FAAy56Fi11YJ5QvVUaeQ3j3Erb19Cn021+LyNGWHwCOgHvXeoT
CU0VFVSzEPHITdVEBBEgtBAJJKmoKK4U6qXolUcWuXibzlDDGkhTMZzUCCAol3W1WqzotupTHGF4
0Nz71NcbRIb5K/jvciPDwLXIpd0pxeomBaAtlATAXIK2QhbV8a/nNEZJFM1Fr92EsoHWU0xF2BFy
yPaH7GBj4Qj04+B4pGBoGoMaD4/hVCpS6mCzbgLrWb5BuuHVF/wGtAJuBQ61C3kA9wDT/17nIc7J
dUxOUenWOWWmvig+twM/FLszypyn2cAalt/ksx0zwYzZi+EfRz9VczH3Ke7Kom6h5MUhWgt8ud0Z
VycCoG5muILjk7+D6Tud1wv+iM3MWSqx7lqFEQcNjjfdOJ21rcuuJQtGM26cz3vhh2y+b1dalat1
dE6vsx05Y/3raFPk1cf0lLXLF2LXOXdXC+8Je4pIUiB7gEhuf6wUkcqx0prhQ/0Sjcm/1yZwkU7r
BETy9nyOf07dhO3e0FujZf6aJ0+sJKrAMl3KScprsqvUhnRayZsytZ3BOqMd2v1dCI5aaycbQZB+
LgJo7fKa/Fp7wOEVu1sGK+ZLkZEE43lP4+WeUAglRQIV8uJVC/KiZxb8ARf85/czhjQiHw9q4Ce0
10fgG6rOxadRqd3Syx0td8quEwEN+PcpFgjrO/vd5zCHUcgrdw/P0Jte0Z+lVdQFpn8zT5Rr7YFK
CYVdLGuz9zvF/cpwdzQGr15y73202TlA6R1xm8VbwOS+gVUehsPNB8U+K8usnYlUsnPL+qRUpOKc
hHf087pFiP0RTKxiQaYxcYGo51Do1Hp+EfEozh13I+JYLSUtjFYtf/6zxFO4GBgt0mp5SQVOhcE0
f/6AO+Qus1J+FSy0WmY9lzvz6K2/4vPSaLZ6hV6DVQCrQQL1Bu/zftfc3zDwOXwaEaHWi+gMrzqz
DpzP+y7O3cs+Hun1P0c8manFLPZTP4LKq8lO4tRVX5axnDt8fldghdOukrjqhGUWG17isEjEsbdL
ozZPVP6PDqkZm7QZOXCG0XgMAjCEDyGJgp9ZxeoXDXq0PUH8VASILKwmc+9rliZLe30/yvioeWFy
YRyU6+1/hUhWN4clG5C/EBznQXmuwT1svVgtQ5t6Vp95rN9Xc44J6SsHfCopxW74OrWNzvnfWNgt
NNlOX2e2eENi+v5ORdtiQWJD5t1AgwE5blO9e/yNvtDPDbZdxWQxmLWZXILC35IOE4/xK0ehKfio
QO0pRsbm4YRZBGbY8oRqmulCuo8sIwHs0BLXEKi5zHoYQjCS9efAnugci80TzpNSW1IRaEBVukCl
riJdz1XMoKqP7AjeP5VeJIO/46ZGWBOSNQGvCPIAZKckQdQaqFEKKmrume4Wn4fbfqVUU4ThiA65
iHm0xcdFYyfOIahitAAEkEKXTUcxpir+V/CsFxiSrF8b0nPksetoH5cWXs9GvpLEbnmQK5fnlUeK
CWUw+24tTZItV9gcxdLG2X751veAnr/R7znbFIbRKmniNcpL7+CXILTKDH257hraDbmTnAl5p6u5
5GHLkI4pPNwiK0FBUEMbkWXNnH4pD0L9pPMzI3gB5je0xTGDBHK4uRZI6ZyoTcji5x9vrXr7Qilo
Mn7Xh74T4Lb7q4O0TKO+bBR7P/K7joA8e7cppKQyy7mLxqNJkFsKBU8beqwqFrVysmcdOtXX4naK
ei4WyTAzjzdcyv3LMEOu3Q3ICgf99hwQc3sLKTDwOsv52YLlRAQ0nVCcnq0YjUL/LDRrs75bN7Ds
NGr3jffedFm6d7TPO74sIMxamz6Cm9OpT125oGsqKZXMpxSw0+tWQ9EQ1dkJCzDeYc2p3tzUr6eh
FG0PD+10RI1q6hKDbmIS1iyEGXDzPbCwvUWToJrLsA8ZdR8HiHfQRaDznxolFoWJ8k+VIvSpg25K
mQksPPC2sbMJx/ozgU/mv4oRv0AzLbpev2ZDd1sNy15Oez187m7i/+V2uVjEqGvvTA1kLdg3lCEk
Ui07vP1M5imxZ0eqgAuStTT+emhQzai94xqY/P6KqojALl0jRKRAQHG49WZkdtfzu6UQNQ+F7HqG
3zAQgqJ6g656epfOmedHsNfBkufEztYTnutGXDLAtXaUy+fve0S9U65ooPR+LWvXbtY2NO1e6Frg
4S/gElXFSyJjeLmXKyIaT3nvcXkX34VHeMBrvqyueFOBFM3fWLpq63vcp3Gto/unqvV4St+iI6Gv
kW5JMgaSRqVLVi/MYsljGxr5XNTXrmGOyN/iPrxGWysML81Gj8nznUUfY16DwWwz3aOO8a92Pyyw
qG1JnJ5OKDvpGHl2cMOIhu9aOBgISztiAMrcy+c42CpCMu4tUX/Xmmy7YlVDqFDNIYpk/M+Z8aYw
ZU8oHEl/3bENu0ePQxH7tHJe6Dh8f1dlK6phob2yA6+9BiPNVpVdh4p0W6TU896ZsfghK44nccu0
iv4xF2zHd7qOTIHX3ZWfw+3zSbdzE1mH7cClAbIVfMRK2YCovuQVa56C7z8SU23I2hWCfFrgCIPL
chLyjAXCZeTiO0/OCLpx4mju47vYqUx5inNUA2cNY1BHJVF5eEn5cl1qMmzpusYzYNvecdIBKBPa
P556ZlPHqf1duJEZuZqtdXDLDRFjpFuqynRErv+0YfflcJByqyVJFDLU8dSJVgdKtBDPnxdkF6n7
KCj1A9yWEbqFQgsfmdD/d0ECFVZnjMh25NvZLgGNbe0V2+8DTf2O2w7NVk9B6HUB1oVl49Xzp2qt
i2xsgGUbKjweFtm8F+nb5qOgsP5IXuH3cWIxMc8e8VyUe3Jn6doXjYGVEUkBDy9kUmsnOCK2iA+C
emM8yd4eZbZKRA0MCQL8gIocxOAv9+tNBZCBNRLfM8/XQ8RclyiSZuiHnfwttdC6aYhEMbHeTw/l
bKMNahe/9fCXPswNun/nat0vonUmYBNK98CGJ+N0/pbRoPb16SNbmyqfLMJB3Y3cXlN3FF20ZX+K
tfawl9IJQ2RoLUVFehK71IVyAoU7w6xNpCuPhUkUKbhK9xj+7Ok0MLTy+2NR5DtNoiFs9pYRQVN2
XFv8pgdqLegjPKYzmtXpHuMjxjYSdJ1GNoaSknhfjvXWewnbvYPAxR0BueWala9m+Z8nhcAUpOO3
JRu5qJ6jiMHt0wTJHNg0FqroYXR8oF8qnE+KACbDX0sSYcCtBSTsjwXrpsrWAdgTs6SnzUJ2X8QO
XUdmSQZf9z98XNcwkcntNfHLF2Tfl9/3CXa49yF0YuJ581rPe8P7CK1pPDRyAP7M7pzKungiA+FE
27B7A2Ae3sH5r4yxKA1dCjpKp9iySurcYhabdpXHpU95yIZam2wXeXz3ZsjE/a0hgs/R1yuFMtoA
oG3ilYjpw3sQQolkan4t9kpQRPrQOxGoHBmzxVzbNLS409zNT4TlVLrcr/rAWaDH8E30gdHLNQu6
qsF20tUPfk4ng/rxKHQ7O6C9DdJjnzoG8UUw+zoZbsuHwh+JIcicQgkm6ZlSjD1XnsoNDQ7gju9T
3W+da2puso+QhxLl2XddxlvpsAWOiWdWrzHeZMv9eSKN4oRW2ynWlR3aNBJK4vxj/rLYEVKYpVwA
t3qd27ODmSkWxDsxyrSpfO8KLqdzWu3cOw+5OhZ6Xs3EHimkFL5QQOIoQgPr0OieGzj0/N0G/OE6
AEQAcUT5XsxyheOBd98gCDphH1GtCnydU1nsgxUhwuHw5ypU6NTKC9xvF5oPvQ9zQzWz1gOy3xlu
RBsYx0QMotIoEokvMAj0BibdZJ6hqtToDC7/F8YIuTegf1ZJxJSDWzzFGRh93k8Jgs1NyuaoL0OO
DJTiWDbStSqmCBAdsKyNgNOphQpQWkkBIei1Cs8CawmuwMXC2OOFWn4HMRt4kkpYUtFemloASjt9
JtdR+r4nlvJVeLg97Z91gIEtBFxTPknaqokRG6C4Mt0G0YQyDqdHYrB0XS6bASxtfnNjF6/hlkKL
6vgpzeqqRQNw+XjFrfdD9IPosFw0o4d/TpZl9c5S7+/KSXiQSeBfMydrJrKOY2moALt9D3JHk9we
9loIzyhMyNVgmLudtc0w43Aiu3GHeZrj4ZV3Krn0VARng+RnLGJRActXcqhx9IUF8vpCFzHPzvR/
SGv+HxMhlBroCpe+yKCLw1oHApjAg4yHwm/Nyh8iO0BBtZ07KbGnx7JqhK0SzE+4IY/kyC9cY/Cf
TV5rrr51D9XmjuNal3eHz3PdqjXO55RcUE/tjBrnmXuRM45xjzzXRjuxuiQqqkFNLPxquT8IVoI4
TJpJX5EIv1EVwLly6CsVf3Z7f9G8sR+uH+ngPkv0qMpPHdpsog2meKHAJxYItjt1hq0dd33jYV3f
8OA9OxUvsNB/I6cnccFZlJ3nWEVMYyAi4LPR9bj4OWDCwBEMGg896+t3Q3V0VX/oooW8ECIUdLY/
PgvkKoxTUi3iO7UEXM4JjnZpVtYtmQkgVwkC9CQ239RQ6yGwq8tliSsBwxqiiXUA5iXTWiCOAXee
/5KWB/ZY96W0nj8Y2WejQJEJmQogIqaCwjUdSXmLIxl6aq1CBEUxVm2z7bQ+fCx7cgXKIzBnpuet
IB1OuKrdLDcmD3jZphZv7W2F6swJEcDJAjGEoZ7dS7tHGtpQPuUh1HecrXwLjRu6VTJeFcgMfQde
UpaIr/AlZr1g5iKJ9QnYxx5MS/D/HBn2MRn88RAkA0lX2xH0qlI+XYBmCQykBy6rYLTW9T7kik2z
ok64Kn8ecl0DoHSIYnleF4LnLO+oyXxhTbH3LTOZRT/AYYJZmFDY543mCqXMx6vAVJN3qyC3d+7I
R75yeIshP4zbgtTw3VyeDMLy7XYGvM2mGfqni+RXV4Xfenxq7j/B0+37NQgimMiN/UYVIbAY3PVI
CR2unWWiP+BcZPjNeOthD/OtcY2v5xhi45BWA6CuhsKmTN/tfjJgoqU/aBe5GRXnEgjulbycEFpp
Z4TaPqHWRiWiRhG6u9w3U308pYrMQovYJAjWL3oH6MFs6ztMkN5BGF1IXif6qS+uO8jwmhn5D68s
NT3LO0Nx3Yltg7MPDqe1AdtgeYk/FIsaaXVM95gMKDUzr8dVzSbDnoJjIOJBkKg0Xa93gTGENcRt
Lp37owH+V7qM/+BxLWfR12GlDtkvGzrt7oke1YRXjBtMZqNsLSGB71FV9mzqKFKcmppMPrQEx6wi
Ihcp53MGK9GWoWMnuT1IdDwbR9ARYyzSaT6GTicffXyAmB0t2ADwadqPmhDDKt9ynDO6Y9svW1kS
3jByVn2cocXZ1qjhTjx8Y6j3AE4lhtB7BPRUK/sUsBpLSQYGxIxiFeW5IsNghSpbvv/msN6MwQNo
Jvpu07lIhapc3OQ+dllrm5yBqfYDpTmxlijJcyOKmWM+IGXxhpHiqVglt/q5Fv9R8CIvij2a5Io6
TiP7jNF3XQp4u20Ln7bx+RdqnGfHTAbOXI7Y2l14btDpzPCQCQ79oo21XD5quj6Rf8dfifgO+47a
SR86GyKmtTifNwKSxFXOKaBVUNm8W9E9yCZnDQGuA9hWdFVq2D6BKQlBN9XR/weQPYPWnjvVGYor
yF4VPy/Y1kH9kxdzJLPpiSUNGpbXXTUVVWDEiUGKZVT5bROoK0wbdhSAVsQImwDsG4u/5NPlXC1v
OUV0IoMfUjNpP9g1z24JmZUkqEeEgZW+usgAsUqg7hK2L4TA7M7H8uP2p8mSFhve2P39uumXaugt
D90aSMVnOY0Knx2PkvsDif03qaAYe9BGPqIQ7mvxi6wv4xa+RT8c50saqLTQ1F3XTcsuFFjMIP5D
xw3SVFZFtiry29IN9cclzdSEPrBLhZlw5+eBEpi3e7MOqAMWyHyJUEIN4w84W4kc241tSStOGkUu
M9LE8ADw7Dp+DB34nJ7OUCOZ6gQrwH8DcQR2oP6toHPRaYKDdEgSYIcY2HyGLalKtWLFkn06D634
k4BhqDlIsLS0PGyt2Ya6bUTWBWSIixEgpTqrR7qzj/5/3eCPXWzcdWehpvZfGer6acm7RgUzJW/Z
fnmmdWkWpU8lEbMOoV81FBTlvo+eeE89Gue3TewBYR2DqaCNQWt5G7rLP2OQtuaX4VLAeuZcybH0
rM+R1yQ7ALZ6tau8awiFRS6LdHFiXdd6przc6VgTvOApvNysRPp1nJ/jJ4kKBiAx0Nbjo9DsfSTy
/+Pia905yc5qJV/xnfcxO8NjelRKWM92amADRouzgHQgaF2+KB7NyxcP+LNG1/GpWcJhoLr2q57o
MccOnpLUO4tRXFfIbf7u4kWCPNe03OgwpAAtxyyK3pJUycqC8wJQK9PtZvV/NWwRtrn8AIFZ+wG1
e2u7akqru38N5ho1G9vyD/oD5JTgV2w98pIJuzmOkpl1U/5F5MDhwnj0g+MqHiMIRcJQUmS6knzp
9jqy0xnte40DZoWF3WT7kUpzCZQHjOv8WfUNf+V8glO2mn+UkUdzIkJfiIxNffGzMYOaQFCL3nS7
cuPp3gT3BUO95iV712AooZPcchW/OynApts2ySVq85/CcVv8Dl9HMH6aLHoNZLUolUNHIXFUY0xG
i3QN4CJfsP8qgmpXM1WhCB87CjBY5wVNyUJa73SezsW66rvYIKjVYymOmioJA6aox0wYk8PFiq/r
98E5mH3VSr0oz6oifUDliYQaM9bGvT2ALwX9bQ2AVbYc/V+da1gpEwV5XSfP0vVGRPgX/SMGnh6a
rce9Q6sGUAeg26Uwv1HoROc9qeEEvdKzKaK0n3M8otks9JGVcCnyvBj3T7JGrhGXgtaKP904y3F5
3DK08q3cooSc9LY90UnOnwSecssLuq+htqAND7d2vGtXH6AfaF/+GnAOQL31ougFaEFGzqqG0HpH
zOrb/k3qxmZjaolodG1UohBepkv+lQ9YpKm1U1DdmdUUB6o0WFqdEWawHYr8WgvOLaHOpiFA59Hy
xitlqRven0bQrvHPkDVZrff1/DHsGWCiivocTcAOZYLE1VlZf29e4adlzu851h3nQUucBYKtXU4G
9cfmgHs7cXGqDC3vRvpVACIi1oU3IyZjSJ9Wrkdtd/SP1Y1l6kUEbEtrWIYkmksp0MTgz8HcNNi8
h4i+Dn/XVyynHUds/n2nIVxP6w6xV5v76sRw9AvfL9ZEQ6AtOpnRKmQwmzk8JlqQbz8tAMB2geUP
eEhwkjcPNh0hisTxO+WPf9KOPmoVT6i+MTw/QKmV5AkCixq7rP20jHR2VsG0DBvGV9Tej48GvvCx
+ArDK0aE7ObkBs3jdMJAAWaki/M9xxvKiRB04kkHZWS3OQq8yzgOgx5x5hsaik/VEukUOaJOzCTD
67H3biDL8NNZXDUiV1taKlpF9nx+f6L6TMgDq7N9zX1biyfLNCAAfrrvhCtGGPW131RdN0v1ri+E
0RpuMwX7OpZcH1F/x9XvPP4YGZ/6bIl81aLYvnxkUrWUldGP0HAnh0aUOU98ku7yDQ3lzKhzKJ1v
1z/X5UfXcvJV3V+rMeOcevOqgn2UumtVbvECe1izO+9xOKi8si6odOTzzGDWhFicAnoP47dWfhuI
q9XXMpGSpYJ9epILgpSTFk9adsYxIPmPsJQT0Q4gS6z8KJUod7aNPuDAucmq4uIT5Oc5rGwU+oHX
SIJqgM7FVzshJL0r/r0QWhnvMt5srA4/Xxlm+oU0ORrvQJ6daiccP7Cs3qmlBs8uppauou2enRKX
4DFqddQ0yjHO9dIEbtV06KytILTh+zNMEKTXTT8OdJlgBMmflz5SPhbFLS297+jh19BNr0bSGV9/
N6x42apZSejDpyCx/6UDIw8/9oegPUQR1oOF2iSewi4a5KI+attqrQ9tadiuJI3YjPbBQec8N9aO
9C3zUypGGei2nc+qXevuWjPQpvPpmnOV0LXPEKv6fOjJYRZn7jDr0RO4V6PvHQVx9WFtg1kPgt/f
LaX2VB4705QRsU/0wEqXBILj1KLWtub8DLra9rXNO/q0Lh1n+P4rDVTdpH9m5CnA+sXqhdoEBdsk
6a9rhs0zjZul6qdEiricSoefmfy97gl9wfbPi5KL7exjccf57HFCgi91U7OEWQvzVZ9LslIBH69O
1NRjFsBHzJ2GmJDC5474U8VmO8su1MapG31noRoTN3Ie6Re+7cu0D19OYijFowXpWnHAE/hNtvtf
GvrEjF6T9zvGEn0i9LBE/K3/WFWd6HG+F4H80qU1z7sP1uVONlbdNuWVtoi10hMZ2mMraWxLAVrc
rdI3x3nlLOpqTmkNsPIgnM4t4I2r9ajBN8CiswbJvmYnZgpHoxXnrZ8ck+p34gDnthZ6pzk3mlQJ
9QKh0DDMBoxmb0QUxMravb9glWrOE9B7ZYlMr5VQZlIax+bu5xzSbszjIKciXemlsUMYXSBbYmzf
U9mNl6lv+TWRLQ5A/fVdWW4XrPm0/iIIfl2OK79lrD1lb2rkDJew2eZg5ik3w9nphYbMqMpGIqZK
qbe+Z4zbZwvpU9T5T61HfH1SNfS6YY7w2qn7kb6tQREDHKULSb08fWUHOkbKWWDNL1koqL8vuh11
YhFm2dGTpeKsEHsu/Pmp282aoEZdDmKC3GyPH1RdTb+jlIqjok3j/B3qwVuC4cGsTAZ6SEa/Wzag
CFJn1GI1yW2M6XaPAnJ0p525dqAZ2inVW/XkbtM/PK1MTXUNEDJTEQy948r+lq9YpSJIkIcg6CXh
Bg/O1DaYnA2mljeYMweUKJGRkSC7z7KIBZNGoE6F3wzzcnRC5qtYrcg21LJ5oF1EosSp4RRglVgd
EvK/MyZAJpJzULmJKLb8Jpd30Cr3qtnLBTUIts9jK91QOj+9XqMTVc6LERaZjPTfAnPiCUDidjqh
vrf1LMbqA5T4kpjtInyBSQS/e67Sg0yE7aiQrYA0ZqmMQQdtwxqFkakvNN4DNaI+sFNWOrrgvqSI
ORGZAfTc0VAjZYNc3K2V9nuHDhzC4yNZ+lWCPnwIpZG6/kyFYNd8u1NxmqqcFQ3UuO+7BI2T3DOa
OJxbUOoluQpS2kxtz00Q0kWPaSaj1JNjmLKkXNuibxN57+rE0n44VC1HHXoKjeX9lgPi37q3mmnx
5y475hQltYetQ/MP5602zdSnbxmEhOT9eY88RfqujQx6TdbwhuCK30TeKDTu92HQwi5Fft9h5WO4
wVPhen7uOen52YAQNu5Is9US+auaLUxrqhNa5UPPaL+eTuh/S/tLjHNz1+stJg3nktUP3GEaTRoE
1oEy+JUhEOYfG7Z25+FTK67JFmx8/Hz04KZnaoNhPO9LhBTUgI3zrE0zHYpYg1WOK2jI3+ljMzxV
kaiXFyjabwDEorj+7j59tbyStjBUU+krC414EoE4TGx+KLs5oF1hKd6q/eFSDM3ohNS21hqkflWL
jMur8ignJPR+xI0X11v1gCIY9RPlqPcAUw7B5BA55UMen7M0YCH4Kkn3mqUkJov04arK8fQTszI/
0CghFUWhUtdylFNEmA4a+8StWGlPqoo6x/PNJiPuB28cwI2lzleP9ZXe0tJ7U3wa+vPDLb/wQjpt
tVqbVMoF2XBzYUDQVEwlKjOmEmrO2H8hPjAJQY4VnQHHlOgm9YRAxfVv2z+Y3tUWY1ClDjAYrnzI
pZKJxBnJ8xn87XV3/xJ9SaktTqSVt/sV1b58Invzwkj5eg6J/NmimC6OS846HqlP6/Wsp06HugvE
meIi7eCUsxOYN60TP9qX48mEtCdtSq3lu7BbcG7Ht/2nM23G3XVHiWNRhhvwq2AH4Yz+HEtlc6oH
XxhozqdGLn2arOFBf6k5KS7YGP4H5jyzjADLHiI9aKtx2hvDGd/onAPQLzjNIo1Z6EF7xtSB/a7Q
bq9U2GJaTLvLl/YhOR5wHQwRdcV+D/Uu96MaclZUQWCVezG8+5xhCihGD+TMxMfdMXAX6ODIYLUE
811LrkJYqnpEconKGX7HcHL8s0ewwpmRLAy7vFg8NPnKbDHIBh70m5Y87cGM3tWtcEsxKt3XMVtb
/e4R6C5/YRs2+RTDtnjZx6P2anzaSTwGEK4ye3w7FLnnWYP5KQipkNmwbXmD3BrFtXEtLpMNJIBn
b9KcMSVufLjCxhIi+O9ut+W4u25350x3zV14wXSuIrLCR+m6lD/Z+gHPXKUcwpCo+QULTMcaOafs
wXeGoUTYrHOjlp0cRLlehzXf0lkZQw85gifSP04zDcItjUzCyOUc7yCy1raPmT19mz+TW/Ct4ke7
jQ4Gseg1C0Cci9WoglYwxWh6O6i93N8qq+IgbcNlo45LHnMqmLkDs3HXtSAfzlAp620BFcUfpXSn
cPR/fonveVAI8kaUMthNp3mVQuKNp/oBje2vCN2hvGvTb7r3aMdugR9TdYSs+Gn4ab3iV/qyQ4Py
xOG2ITHhAed4O/5bmAMnId6etqx2C/bhzEnakGcHPOXck+8QoiFr/I1AvZxdvJmq0Pq0IrjEdX3b
LfXoIaIwTpHnlHQI8syYq1nM7uDpdE3i98i3YXXdziFSlAZXIyG3yUrJ2JbshfnBU+gM3BOI4JNc
L3uBpxjvz84nmhF2UKs4HU9YiOVIXGaAwZgvHW/wFyT0fR9QOavGpCCXHb2/WoSCtjGtqK3genDR
zCgCFcmoXILFGUQg1UxUXyaeCp24Rl1nOAv6W5h9yqpJwswTqF4JE/VDsWX6aCuFPM81qoS2o+XC
kOZyOctmyuyq/qu3YEc/AB8ZKcgTAUj4IrDWz5K2gE/OP2bWHpK27Kcxydyg0ugsmqq/s/z33rwy
tcPisTQNo8i2zlpx0BEbYMiVKrTwp//NtXo5yem9oeyzssg37OQA1utUXdLLHodeCK0EEe3H6X+B
nRbeVVWhPm8feuEtVCvUrrsW3VGiRPUpVImIS9J60v5cYtlT8XsorA8sSQ/C4HSbi7C67HI5DFUH
ZNmlfTL6IoJBHlJ0mupB9ePZgN02vE0HFKvB18IDAS0yqd17dkUSNMsEYeQZOkGPRjJCCg5NZ6n8
+cdjSBk1V33eoHxbNM4R4t6fJhwh1kfFmrT6lBX7q+bBK489CuHgHbPqduLpt5GLxtewX59xQPt8
J0dEYd9CInoIoWsL45phKZOoU20mUEnksT1kc3c1Z0J1cY01KVNkv2yZQl5t/fFzctUUSMUZjFt7
SPqS3aCNPhr1UE+jE2eZ1K25uJ3U3RELC4UtYavn7cMVWIWlrgTCEQo6yF/QcxbI9w3F6e35xwV3
4PeoJEty1dGLQo9IM28q7Ce9uFrEKybZ409WFs8TwuRsYJwKgd9IiRNLHhyKI5DuV3WcE8fTkDsA
6glWVokJ3zTJAwwbRMiY/cnHMPj+0qXUsD7+ckGRkkol5klUFA6Ae8vPGN4eCAXArdkBKc044xMS
iuJNebisMa7hPnxLXngliSJMyKZpG9lCA1Anp9T/ikQ3IylBaORYufWovYxHJ9ydTbAMG4ynxoj0
i0BePmOcMQk38eVsm20EEeVLalUoQ27di21WWJKWt6b0liyhr5Q7HDpXAMUH/MPF77APM3Udaqdv
+XXt3V3c+51K1dsWWpqM59xZ+DyVFNCzPxDZrCL1VLmoi+K0AJPsFuHGaw8rHSnGDt4iXiHZrf/7
8Vs8bu+vx/V9Faaj9sq3TK7pNoBDQVEtqkHvJrFBM4XTjocQoGfgXAwOIIs5DL1cdJP+A5Obqyj9
T4RSkg1UTfBuCPLKPanAZXnKJNJHOXH87ulrVdKbqtlJly28BIz3tpMTxk4nXHFNbHo7kkLZUAWl
JWQyFLOFHrNYAYx7jN3xmqxl2l0RZ7flauFpv1gKKPyDjchKoS76HxU/byI5CxkPOXiwC52a/8pG
+MsGKnqEXBTrH+STK+NPq7qR4+zxoBS+wWJqIYtcY8pcG68m872DhoJoSZV4M33GySC7JtObQlYb
nzamaN+FFLkuimS5kxr4VXWyzHQEV0VLIAGPlYu3YCyjLMkvH+Yt+DImC+xG8xNfUDRYRw0HXKRr
mJCCR31El7DQpMVWRocTWgmkJPK/FTdyjw0iTtUqruFgs8hd+8c0ItjWfXwyadRiH2g/rkB8ozs4
OrRwovkdcX/uGH8LL7jntzl3pYiTiEz2m5lDOtbQ5vt8vczxK3pI95HLiXRNVHOHcADAZIII5tds
A50GJ1EPScsdKh5qLjhknsmeOynhTBovvV7MbBArfAa3nTWcHTWThX2f1wk4ftu82OU4ileIRall
+YgMEE5bRag4yS6iNbsJVzkMGduKBHUCXGwuabKNYbPHXi6HZ8y8RUr170+oWygGTxueYvRZzLQy
jzA27DfhK5lPRMwnkcRgTtzUiHrMdDLomOamzNPittzXfB8vY6ikJI1w5+PZmrqS7HGPhT4KT897
Z9OfqdKoME6XTVad0raX8NGCPHoSp95PoXiCkU+jbecHAEVaKSACvHvL70G4vgaP42VPdu/VO2t/
ErtW9fHjdGWqQLbTDuSopTtzGK55AMZaeYo1OYlX4XqcNaQRIS43nTDG/DEJDqN9zigSIPLaWmpG
mqnyAcOHsw0EIZoDMZi7BIMz3X5jnL/96VyRorLa8SUVUvEOLcnsqQmrF47yiOvYMv1tgfyvp6e7
jFvbz0+C95/3Dwx8Jfb+3iBzycEoIKPYY6kOfA/6FUVbWNzMql+KoUiAcvZxbdbglcNDmzf+GGnw
vjdSbN6BfqxOSwGRSc80LUsvjKHvMdXp744URKJCvsR5iiQVDCz5w3PRcYs2g+0qtbx+CaEw7wbT
snWsyoyYbKmdOtLykTBWpIJrZmGPvqZBWk7khdhl+7fJUedVvlqJbk1JjEyEsKF42xOSWDUJhIdH
cwutruC3QlBnR1C3MaQUx/g8z7U5Zh9nflJvithV2cO14A8xAB3AMhvRo/XUFx3Zt5IAIvBEoc86
SuM1NULzyCgli9hCajybjHPdIcW8siQtozWm1KInTu9UKayha1WSNOZSfmP45J1khprEUlsPZz+x
yq+QFeSq+gHwKn6lN138CBzwIL6RH4Fnx4J87k6i5L4Kj6wJiXD6JihRY6r2z92l8CK9Md0M2VvL
/Gu+ByHkvZaramdepPiJGyoysWNcQAIng05x2yzgad3akgLwMLO+LBLlrcpK71WA1H1yGpB5fV55
rYVURzWJcGNGJSHmCN2c2FgCTIIG70GXk7zplhitlvJPDMdJBhnC7EG0Go3iXDJcoFwNHf19V29O
3sQsxAQb0hkqcAYFAfrejYOdA/LFls9C0Ng4QI9ywMTSUgLmGQ8Dfkxl1h8npX3xgV6vpADygwaM
mJ8KSJW1J9c0kCDXxku0haMXYE0t8+0jZ73yV+WGF1vyUhR1/flx0rksxF8IIWgduQ66Cc41m2L5
N49abEA7iny4Ug9FVa/EmD38JjNp5Xv8+amerx/Y9lJTGGeAqB+gfPQZvThQS6vOK2s+FL+OhdkU
lJgU5RcL0X+x35g+p3v3tXpduc7vMGpX7os4fpYfyUAAZ+GBG9ELr2ak7erIu3flSZAl64q4Wrr/
acx78r0a/qCCT8pw54qx7MbfFpuKAgw7jOMKnquy6VXsviQ4VrllEFwj1PEw48hYt736MumdH2t6
xMSdJFSMptMrs915BJTJAMQM9b819Y0ghIAA2J8E6MhqE/UqLWaNI1AHLoGFdKSwc9KUYctcTrB6
/k6H1TM64lSkgDUmPabjzfKHjRSDTRmgAn+Rse0XUmnPDgbrczjZA2Ku+4ReF4HnkOzoeKpSNp85
coVz2neNoFefRLRZfIKMZiFE+uiGvAAKr8zdQSGcU7yQQA0Uinm/jaRnBVebSUVNCN3pGxvfeNBf
TXEewMGzLcIecSDBrkP0NTk3xgrFgkFURgz4oBrOsfINUZB7/VhnfkV5MhYGhs8tor24plWM256a
Zk6QhyE13WWjed4Rf+huGr8siwpA4O1pfC8C1DdhMD/cehz2OLoVtMru0CpDg96eyccYq0+SE8yY
1xmSeWoBr9ToloUS1C+KwU5iqggeefYJZPdwqy5u9+EB8yVrv1HEXv3PFI4w9zO/gSJWune8Ft3E
5T2/+3tcx09bGC+hq89RWJcXVd+pOmEBul0lDQrZ1Y1kIkMCw/HjGmc5M9Yq4/jSd82XOSlit7dM
Rv0oOyDTzq6N/b0nBRe0Nx+Jn/9bvY/n4q2Nu9BDjZK6tkALo/9fb8sYCIN8nzReCjZGURTyHOxa
J51hACipUVkQg1Kray7ipqS+wiOxmoztj1FFEB3PlCMqUJrySK7mSMD3q4d3EML1pi/KpNFL5tin
uNi8F5J+KXRhREdFZe+NsXUlJjb7lr2Jm6Anq0u6WtA1TJJwPYEtl1fDsUSzABMRKPEd2LmK+oHu
E25Q/7VolxsZFIJeAPF3J+IA6mVAshHgBiTY8tFcVmY+LbiUy4ddTr5QIKI+symFoh0HWEmIJMbW
fNwcR1QCCP/gaPxZ6h6RmprqNzliO+v6QGw/49wOWA2AFHJwkFk9ZM1aHBSh8hDN5qm8sL0Zzg05
ZAIC4GG5yDJ0Gw42/bv2RuaFqjjk2+bZfuClfcf4a37U9wzRiW5TfI/yhozwZtcuxWe5vk16r8Er
uGmk/mzIbH5wS9gJ8HV5KFNQFLb1NuyvWXKaLiRW6YlkYqrrJC7imr2uxzePUlbxFXxQylpmh78q
WaysgPrz1Nb1EYtaDHCdjXo2GukaYJP2WtqtyvQkAmIPb4JF5GhLwjLxB1c3ls8HTeHE22sP3ECD
qwgN4GTEPAuIv0/xDFIJtbnp8alTAS4xrLFsUznLVXDsIrfBBxkmJpVauMSUVfKg6Hvky+S7Mp/C
ISN2iFnP/I6kcBZgWBrChNEO57kPI8vRQAuq+LCDjvObMWC0ko2Of2bCqgO/8Ojm2RU6YH2mdJpq
3S7GfRkZvibwAIsYNou28PLyIPj1RM7+AWZ/4Zr4qRzzYky0T/+brgp98CYp60PA5pg2SdXtNa4e
JrwdyK5hX7GSACm2zYv/sEvK3wcmBbLOFNJSllZbDblBFIMAOgXpvxHZ0B7p9Tuv8XYpzeVNmU6Z
ksZH87zNuNDLBcT+RniQ1VeVmzLQrKrGzF1tVJqcijL/UpV5e56hpjEV6JMwBwde14yAYKp/eGR6
Z02dxLuHRDnDmE5wC6sTPJmpWRRfukkn/scTATFc+7akp3qFWikI7Lu3joGFFc1SNmUstlw3zgQl
UzDoWEi63DOxYXGIklJJfdBypu+ikd6OYfbFzIe+niIskiTFxA4cR2Jbz/9KvR4KrVEx+GY8E9ja
F+vjb96yNiEc/9HbZD9j8JQrKf9Xg9D12FFjaI8PMja8OELo2RHl/vzMd4eS1iZAN7uhI0WPvqqT
Q3XeS4L+4fqiiHUv+GQZE3P6xEvAInd+2Jh5rD4UOvMb/4YPhGAsF9dQR1yoc8Y99u1DFPHurJj+
RsuyCQJlex4R/AoSYibZEVCrHNZxSCU9YGcn+Cyz3chHd/BCmmCnNggsRsBRixoUgayf1GJYO2n8
2+tSv813nGN5oV9+rOOy1aCfFHaO3Xyybe4uOOViSq4dRq4RqMV5kQER3c9Ejhfg4CfSpUUkPEeZ
Fy241IjzPhXub6gOfxkU3NazdXXpdb+//uB8nQkjU7oOmcYfIkWSFjnrtVrRFYtyORN2VzPLIvm3
hk8gCsYi0ag0s7EEkOjDL9gl17+4A+rIczGdmiZu/vrQsBvmxGKnBakFVa18PQv8F99mACDTtEos
XnCso8KAjME7sG2qySIV+z7dEfO2Z3MrDcbAklSiMirrZzjTmeb9E6fcWkJJt9RLib5wx2NJgHfO
fFInXtyEdtXPJ52GG0ozIrfeR6/r8s5O9bjDZm6o425lTsDKicBfSpSPs1pqBY9kxPGX0CVjNAx8
XXlYmSjLIiKGFmdFvmZAv9FRvmV6N/1rTyXcp+9fRPD8XKGVmkRnGbzBLsvZUZlGRt7ivd3ugTOD
ejbjFPELDBnIYIGhu5MvlLvYA1/Nnu2v1ZGByoLya/w4tkdNeNry7j3Baf2weqHiKineVodfbrOb
I2J9+yMVv1Xq6M04og2E4nnTSzI+Weg5eNaUQB2Uy9A7dEd085+0oO5vb3ClWsEWz5rivT6DMaTl
TLb5iVZfVEyJUdUyD2lvdaqqaLozs8/HdIpPvCnfhYnMWV/VQoJuaxTBe+jn2QLvCiqW6EUX1gF5
UO5XWnR6VHWjnJtyJ9OXwuJWd0/SdmWdFj1PTBvAs91SiAbjWPPMFbQhEXRp6CD018QwTY7emEaQ
WuiP2jDU6TSw/PZQfRpaTiZYoUFJVjTR/ee7NWfxeL5ajOLY6mjWpo8jTlHYpdS1QGrVpo71Av9z
fJtC13NRWJPQaeZ8+QF4/k5+fHIEM4GWNWjJ5yVjDUShB7ye1Z05LHd8ZX8C7OdZSsmF6arVAw1C
UY4MRKM/DmFYktUhmldFjSGctipHvwStO2w3E+5MIGvFO0vU8M0q2+x8eKDRXU55krwNqiPOBoN0
wZXxnUrDBvgW60oWOaYWnTMmZv4B4YkZPAm3ktQocL3i3Toq5XNV3BAJzaISqeJcM//D0976Ochw
ITX/nfPISQ5IxZT/iIWJd+q5YpoKAT8nHri0pyXrB2IeizIZdVTf5UePpH/mDCDKx9C9IVNSn9iI
Kz9BEyKkXHXYHC/FD8Xvt0t3OM6yxhfCOCZ5IIfIvAKKqFrnlbOmYMU9/35RCME35S6DcOLCg/ki
ufvYh7JY797gVIPa8z0wU2ZwH613cVh1n2zEtVqevVdvk82KqdtReao9k/m4XF8ush+1Ghy6Y3WL
UHoxeyU01s+XJ3mF4Y1m/JcUMOrE/BPIL0fSNT42D1vGdSUmDeT8E8EVE9tpX5IsEEmepOWGGkSn
/pPCejTgigKijtvOFAZ5g6VWuTUrzlOPDYzjCtUnXL6RG1hbM35ILjrITfv3wmiisS9DtyZGEOPX
vFddOfLPodhj9Wk+DQPNr/RWf1C7Bkd9ofr0xAoahAmYnbxVxJlC/dCz0RakYUSNRLTqOowXmNVo
022uWBb9fMg+VUKJ4W3nsQOZyq2YOd5nZC8iCHb1wuCIdEwKQwyNKmyv/n8hRZUOhhmKElXBk3h6
Zs/u9IvwyMvAF9YyGJ26yyGnl2/dcZpV9yEO6jPje+QjWFIGZv8hX9F6/eigGVOL1FXKqVFrcH/l
aLusVfz3dwUAEUEtFcKburF1wyYXdFupognxcYcpGQLY35D6/EEG+T3rRjXeG6xoxTsDwPFjqkRp
9z8If9dZjtUTYtSWg3Zs8gObmrlb+Fn/3+Lo4hS5l1vMsqTOXnqhmKI9EPjNROsXajeD2bvKif92
Vel22tiKFZTyoe9WZbru0kY/jBofQYIyrr56ilk540PQJdhr713+ob+vp3HirahjXwVV/Rhgalmg
aNysi84F5xbsMbyZ2z50aOViZPajAiZQNo/X5kv8VHnCrY9nEck4Jq4lia5iaLe3sZAUoNmURPOU
BWKchBQHudLEARhRMtqSPmo6jix99tGkoQwm1Lfv3hyCvPxtdZde9C/82Aec9E2WI7Jd8QlEqyKl
3M9a2DqGJDKqj1M7U0ZhjjTwNpO2Kq50aIwoZvPre9j4eKkpixnuF2Wt1CZ/IddBcvohkP0rJp/v
U6EGDiERlerSzUxfhLTrDqXedfr8nz8rQd5Xyohz81ZvROIwQkvLV5cmjCqZrBBuorPfQhd4zfc5
R2HMu/y/lgl0SiOv3SpeNhzkxEXZxLbqvCEKDl8PnufmcXNItQZFXMVgCFnNW3mhW+Xr2PnX+D0Q
SxrL6THK5lFrDQOBU34WmN7oIg4taHx6wT2CC8sPdMqSG5ta+dxTbsWVbWAHoy6CRLuDOMXO2h3r
XDZjID1CIDruMnouAnFObFDM5iuhNjHoN+sOJ3KCDUl1Gi1sQSrrCvPLH5rDDXFqYZqKvN86OkHZ
pxG+9gLSVGQF2+QDzeUk597+KIKwMegHS6s/2xMiZBsZBHLTMA0boR/ZsPmon7AhpEl6PEkEBKSQ
YzlSOL8G3tU4d8vaWD8qIRyImV8IbyHNSsp/nFXT3xmd6b58pUD7MzootbxdLuRXlnxLgKE1A/51
X8gOyR+qWZMKFOhBn3MIpVpApQZjW6MBsrTqfWzRi90J5wEAvPEfMWbMLEAedKBbsRKXlfO55/kO
ESlP9pLc6bPoOGfqoN/bIKXrSJeQKZ4YqUqm/EAwBoh7zQWUFKb531UeVJmktmnegdhXb2cPRxLK
a9RnvGbKt+K8PW4roLu+bAkish6heSYqMf1EEozQ1bf8iQAFr5pbDjboNjTWLD7LvZtMTc/m05GE
EOV4gkJu9NDs7R98ZLo0cS5lc5ZVfZx+ZaPtVxmWSv8CIpDFK+cOWMdBTkHlUeGtGakq5uytjSWO
uJjBlVGSLFCqvmuI4BKWKyyTzGXU2fFk8TkVQCJHFSb36KD7TQo58d9wNeiKKblZLtLMvmikpvbn
GTAghvueQ/EYIIiW8BKbYhanIhQW05G31yFejBq+gt/4l8zVIhJfhWXuHOQ4CeMOErf4pniNCno7
Qfc51FKQJYAMvDei8EPNkpL3WUE/QxNr91jwdGhYCm1VNFavvwhfvOZPWsj6Xbb4KgIdy2FW+S8c
tf/Brf1WD1Nrju8c8czaRmaoQzwK8Jsf7+xbkyVF4g3icmhcEkIb6DiBuk/wI/gscUP+rLn34Hkn
ApMbQGNbKs+S+HY49lgA8xBe8TSbRdvvrPQmb78Ev9OqNbpGxLW797jIihfWHNYvblXKXXEE2IVa
ngtwElhWNMp8vfp0xj5Y63I0HN293849h9h6ZWw/O1oIMQTdKUl07Bb0y8UDaw9vC4i4WUQcTtEh
DN9JC++XCXeJz5Uub0ksRMxk44lX6Skt/6uC+EMS83WFngRwdTLaIA9JjqD/gYDFpuJzWqU5FDZ8
8NpNTckezZYdoKj1o0j5uja7lIl6o8Q5Rj8HeS/D7zeEDaIuasYxtHeI7cvkz4UJBpAwWzp9FNs9
/SXJZGkO0UQy8sQK1R2pob85crL8pLaQi67gVp0RdPM5n+w2Lj9RbNIHEDvXcPITgANlkZvd3N2u
Zh4Q7WPGQS1DsRHwyg5XhG/EQIWZw9K6alPTwJ9xZ3CZt1qnsh0CmEXhWws/aA0wg01kwGW1UPkM
zLREct0NXFvM3yZ6XjQBfPdg2seGX3rqaOyHSaPSYcf1Zdy9xBR1GZ+a0fBMS1Yyk4vgirzv4gs7
+OvYiK/1XDeX7EQj9quiPZGQpq09Y4nXtjG3nG+Tij/g9M/kinNG8ceo/pnJaS3/+ObxgO6UzXGI
jo9zYOaDYnEEq1AMydo9HI7xwPwxNe5sFqQhPu6hRSLj51uURlLC2tU2bAfnyHoeB/LYRfFRApbL
xhDh6HpYq1+Xxuzu8AzmJWNlj22BLQAZS9NF2pz+HcP21wOFTs/gy7wvl/kwbBwkPK0p7tSGtmAi
mpT+Gn0LHxbyQh6Ke9i0rM2735umCe5EiqPT8tUszqV5WHCR+4VysamHfvhPx+jB2o3csZwLKZU7
q3UNxZ8UZJ93ByOaKMkSkpdzyp3aVSMWvj931kvEGlRjhOgVYRSgptC6x1uqfe8MWxcV1pcgwQzZ
XMAsuyExpQBinh6pl5tZctuUQYstig6yyixXQXqYfoXnxxaKoQXKJlm0e8TnydOJv/SjeYWbNmxO
K6BY1jpJGFJaBgZrpJr4ADIbY/asxuvOpRyJmnV4gvy1YdwF11Ji/BPaCwsp5D9Nr4uxyS9/m97r
7gei3Kp3Mpl4Eol19Pe7NJWsX9mJY1ndrRSAThxc8lq/5W/383utLMIPGd2wpExouUszz7bihSdw
MWnR0jNagsrSWEQEBU6agoxYZgdo4tQVChpyA048B7J7ItlT968V81AZytujh3BOCexcohKXjqSu
4IFF4Ir6Y2CPBYwHcyQcQjcYZ//g9rldacOp9DlLSWWkatCj+D9FeYTjt36PSTFw52G2w3dpgpO7
4h7+INIW4voGQ+pdQWhRUMz6BD0iBf4XYIGaKGiBQ1E1dZ1Wd3/ETw2ART7TNT3BB52ETwaFzYvD
BBEjNXWBhj5rIjrtu0Bo8gQMFgzBUqqFml7qPUtkwbFzns4yw2aErCIW/lAOFJD/fVY/5nE/BLl/
WmjQLRqnRuoOBiBo0HBEXzNLuVjf4FSDzMTMC6kO/sh24qW+z9YYVKcaMYNe6b7BHaNlzDTqXQkv
UmtTqoxKVfx+Ccqb1lt653+INW/OlYgi2TeB2OQbdHIJd1lfppwpWEcDpR5IgRodT3M604bKygjq
5Fd/eLxjGrdhJPHYrVLRI/ljKHv49lQ5FbjWVsVPWoVlJGbzjz61TwLKpWOsUnoGEeYsdyuH0+qk
xpRyPIOxOFopCH3jTbVTO29GCa4Ubc1Wf4zfl0+WoKxn67k68qglbyvS7ZuBFivA6Bx/6ZjQuTeD
JkgGEWlx4Uec4RVievEMKC37/hlnBWTzSQClAZBHaOrbPuVlnXeDDXxg+o0gL+34/Dlj3DS7Hgmv
1a2R8W7AvhpuZSOJB2B9RV3bF1M6bSLJz7Cw/vgF/uSqozswKBSBfcXtvIaDdv21j/auXcWXU8Sy
ihYRnBNEfsq0VCQkSJiIRnlwSl6PAJxmxwzk7c11/0zwr/T7AcgWaeYvZUQY7OtqZbYn3ddfjCS+
cdSzZ+Oy/n4VZNL5WjNvvoNGSJOEHiaHP6XdjTZJAAx3a3OElnJRnUZgX59Fr9TJzjVPQlgFpx/n
Qz0yIBALE7sZR8O7REcx8wGXPoa092FobEXot+prSWTU3GoEcVS0KVbfxpl0H9ycqKlLI/uVqDJK
qKmlcGdPtzcf1qknI8QoJEkGuqDzcGSPhwoYmzMXy3QpLD9Xdv9X86nz+PzmB4RGqs4/9TXTgNBd
3Sahqp8C662p4VpW6gninq6Cz8skO4i1RmvB+gE7rmc2VawjULrHsR0c8UIiqG+ZhoMPIfCOLAwL
E6ciWbAJozVUYq+NuGrkoe4PNgCcT2+IyjU6CxBmyxvdahPh5XvUtOHThsqaDll4M9603tJh+slq
vsPwMo1RlUZP+EaKQMFhg5j4ZaESr+6K2E0wrc0IXgBcyGlKfG9/FSmKf8KP6QsRKd+MoILgrL2T
73e3by63+fnUTtrq14Por3f5Ijh2DxC3N/b/Ke3h9GLnc5rkkHThw+pB8j0sqisH7JL/L0lbFmlq
luYW/5j22+Y79GyrvePSmCKTSlOZLNJW6NlA4/sDxRQ8mb6AMTn8vlWCI9Ojy8Lm08rAOZlCXX0L
Pqyp5YzR2yx3HN8ER/VPWJ51HPwTNK2FV6lhzeVZcbgniCmB2c5r5BhMGNs15s2JI2QrNsRmv42S
/PSJLv8raclvwBi/gD28gtekj2OD8XVZHLhUsw6Td4v5s1ZX4M3zhUSXhdNu2EXIHyuFR5mdiPp+
It3HjG/QbuNJ6mzaDVWElDZVhbTcssW+C7fPgNO8YXsyLoDcuAuDJ0YY0kfjJRMsR0CCyKIV2CeR
PrCRic405LZeQ8fpGxTOWc6yF5slBk0r0PhD1+f2aLkgLouNZJ9WYBTZVB2dl40QMo7dqnERGRgw
wUQd6vuEQLBdWnFKZovi4bhBS3XH2cq4G3bfse47VAqDtE9MegxmzqfzxgpgWRZWuxC7PhggJiqm
K1ibSVbRiL+ZKrbyyJj2RDuPZxtEPI3h7UXNOJfsqohIx8PDkrtn96MNBzuFQuqyQN49VmXrP/X0
2FQIepkfL7G1HtVRtAmKQV8Cr/14CwWNScpDyie0ROCDFw1FYjzIYC/93c7TVyyFlXWhZiXd/rhn
Wa8MjRlhmyTRbs6sutvW0tYZXfKhDiCtns7yJD19w8yE6lsOMMIZZoC8TZBxdPIHl1k9FXyWbMFD
qrKEe3dctyabOH0dBRKkDHmOjCkyfwFWk7PtrPwlmQxqcYYzIkGMTe9tjIDiGWE15AGEFGM0IbKi
9VPWiRrEZrmUzc+0Zk3WxbW/f9MUTahGQUFFwrZ0NmSTGMny55lHILIuzKt+crgZIjSdm8cyISfK
5ljAhHHPsSFxFdFBJqmQ+xht+VrgVeDYOjJwabqxJBSQNkznjYNwleuRzfR9rFFaCrvbaybrg4yv
bEjjRyZ97k+nBYPL5lMMLMi89JNLiRi3htRZ9nxP8xsRp10goauwfG2LJHxwF3YkxXDa2ChujWix
KeS3r/XU03EEE+tWNRxEhNia2ogFl48QCE+l2j79cVTu1YlW+E7X99urC4tr+thIRHaNBJ8tiJ+E
7u29MJO2A3Nr3WbMqdsQaAjNziyiXbknujjKZz2d8YjT1wMsLpAf5lumsRuARWsdtR/PdV0ukUah
HE7UC2AXPdrEdYQugGTRb3SV3GcDyz/m3ga/3mfN34BDC4bSzhWpmTj3/yW58Gog1fB6R7N2ivN2
91O+LFVaEU1jF3djUADME/kZZyjeAdu8PkKqeolIThllMyDOkXfPcfB5kWtcbEdnDW2R6fUuAHDX
IjtIox4t46HVuschYPUUKoAcvO/YVdExX6GFRwY4dAZKQXuxvWSqVN6gGNIhL7aFDRzpeyVbRJcU
15NDGEpxXqYPP06Mquvpgt7iYNXZtXaQQPMHElB480VVkIt6+Ae2IxhZckPJawItRkDYD/JoCBGm
Jm7l1syWcwWaVvQCw1kf7ByfUWXeb3d79d3datELcSANlwLuZEWWYuyYZGuV7wV1Sk7SkS/8fHow
I4nhr6FbU9+zy2c60xZAC5YH+PuPA7hN9axbN5RasL6FFTdDLuArsiENsdeuLbC3shyxZh7Iu5nw
Jl5ecjCTtVUdqUMz93EQOoVQ+Q06c10Yp+3sFOlOYAcyNbW2HqiR/YIRnYeSRODwY0Mbc2avqQx/
pZcokSe9FhkojB4m3f8mYQQYcyddT9pjvWvtSp9X1v0kV3Z7tEMu4lvANdCT9oDRvy6n7TekXEQv
+QhzfMxc7JR+OneURz0GdLxNWFbOJq3Y+2ohuxhYOLQS5yaKvE4gi8f3RetV9U5/oSOf0kXb5X0k
oZa7DeeMWiXusBGiTaRlMdXhnhjO5/j2hDCkkHTAANIKSvTN03LZhxaS1pdp9k7lLS9o5X0Umr4a
Y1v800LF9hHuYTPf3yvsLG24CxQReJgUJCiPufEXnd6PnyWvNxXR4Bb7OpPYBvc1u+chPHkRTELJ
DgpYglIa0/JAc/l9b4FJVqPVK+6mjcEliWYO8OFxjgPOV1FNVGhXKGfc+4LHK59h9FTAMqa14hBe
1Z2Y+NBNc2qE9/0cBlihGJG5zs8YyB2nRWAc2mXtdiCwDPdQ79/Q0XeCdEBwk1BesuEx8tMRzF6O
plSjH7POu9cli3cCTffZ5xJ6gDvTKSiP6Qu2paY+ZrlPsgKjQR5GUbThx2QGjIanKB4cAAvSEZtD
fvYxkKZcyE7vLMlLWWrrse2W/naOBnUNJzA53V6JfFn3V6Z90ckioBXzvd4htvxTb+8dug/IhLPi
b5LNOxxW4d6ozRxHBSu1P6Zp3Jr/YSQkjFX+9+L3rq05A3f72E7rNsW0FM484RV2qNQuQRRmA0Og
29JgeAPqxUNFJlB7NChhYlCLpiNoonmvMpsdwuCB2CzCAy58HxfbIfgvD/DE+6y5VivykUSY34Mm
+F6RT74DFTRJUjhEJJoYCF3sHTvf1g69Fpk1++G4cAtCaC+mQ1N6UJZwiTCfcKs3TwC1Dl1AwQyW
pGtuBs3ZifbJUGuNPD8vDKml92RHdTXs28GVKnTant7BhDl5RToxfc/Tor+xRHBA5KQA31oYnd/i
1KmbKnR5lro0oQHe4dT5DBa60nMPsueH8tD3cAQqHa9M2rCbg2khZit3LZa4hK9uE8oq5hxSOvcF
4a3E7E6ADagR9u8Mfjx2MRAVzQce8y5lIl7/B6XsB9CMpk7vkRgPCcRu6vSgwtKahax5cstotLkV
ggxtKmuRernNOJYj6OGtuZ+90yDAxdjeN4rec/LSS2MZw2kGvjlb05PBd2jeHn65+1vRWw715AYE
yGK4Y99KslKvMLv8ZZ9jTvfNleZe/L/L7/91dHNaiLUI7/PAiEUTrx9XXgTfIs1xaj4f5rq4ZKkl
D/kqoSmFsXFANJKnyPdLHZiJ+LOTfwTVkdAL5hgBuFSGiVtaW3hnGsSR/1xG5hHqGeXfppn8t7cX
TOoVzfD6Zj+GDnzTjUs7HISoDx5z8tyrx2DLfU2GnhgSzTxu9gdw2epF7p+xBQavj161tw3zl6kT
i0upAMl+8WvxemM3V+NTIDcPcttDg0TxCzyNN3307Cl6UFCswKbAs+K/hVu2voWsR7ESyKplMizG
LTEd1xB+sLHVYLkC413/j0LjVDdfLqcbhMv5OGdTrdoOBzLy7UeUDbKjRaGeehpngdNnEaWS3FDm
K+S1r8Y4KfUX6Sx6yIKtlnvr2712k1Q2EtS78xIZdtCFigVwyg4ivJ06W2uJY/0cJBrLtTbd2sp0
g0bD6ed4IA58q4gtjnhiFUiSIbjYCinRkgxqyR7KLdq8fnVUKPxyHOOHFpSbDrJWgjLk6PBtzLs+
c+P0dGgyDcaJLJRZJfKeEmHoLZTL3Bje/0rEqy+iVCrID9uVYnQ8JAcFAtNDSq9A2P3KWktcpH1t
qSJM583876VlIrATszRi5D0UdgXQGGkIM5r804i9DZRH5LobZ3VKOkbT19y3hc4jfmlr32nfl3wP
/kPt8/K1TkNpqFwwH7bawr13XqhGrFsb0dnEeW05uyv6fiSAPPn1hQgm913YRAnzf/0UR1St62ll
TYE25eV4c61UqQoUYH+ODYYT2y+fDSsuPH/DNr8k3OjVoGfQINOS0bZyWtXVOy4xICRgxdhOTIJZ
FG/RE5/md89K1Of+gb++lxNd45yG3+75z1mVNmy5pBqP/jui+tYilIjv4/zaE1Yiwpmtj3FCacej
kpLpBEXg2sWwt5q02l9KDpl+3kba60oodm9EVc8BVJafBonry1hlG18DQuoYsQwW7PP1ffFkQuKD
6bidTPnI91h3D58D3iW1mILhN88u+yHseT4U2Cfg/1/YvJL7ifWLeguP7G+BZiNgiocO+f5aBJam
ek1RNeuKptfJ4D4ab3knZScadhet0gZZFT+3GH5DLxLTVZCUGKMZSTkal6CybUthU9LdMPgqiBzu
Fat1ot9+P7LO2m9/6t6z/dwG6bcSHOWnGJalHz2x2f4SxhQIUyL0b1Be03mn+DOymDTdJ3GPZeNl
0qmBUjHtrfgRrGYOuQx1VPTKrhGVatpLis2H3jvMq+4hIyBtM2yGUoqxtsNoOAtcbsreK59wDr3x
3FRqYdoCU3uhJL5F6m9s/DUsFXSUrYDfmwgrtX34aUWJZ6pbROZtAmpoj6a7jhlRS29QHrLCbojT
uXuw/0JIjnXKU/b/byy1drLE0QdfTdXSCUNMrmsOXDfFU/q4ssrqDcEWuHa/0vshym8SQ5GoDbM1
p5U3fHA7yVZRE2OCB0R0rUxVgBdn8XrZiBpIanT1Av/LRItFaDpcFBXeOVqvt8z0ZOlCQSZzVasD
+WstHQtZ0FLU4aRTgHbDZzEHZ/ctBxrTZs39RSo/PTvwXW3uSMrbqhPRIBILvSOU+ut4m5ciTD9Y
1tvy66pFeMqhjBcVGaWWk6zVJkv5wBNh0NY9iwITeRLXXSU4V432oUyQdELxfqFdUHxlKjO/oleI
EmdnTaDBsQgsKOa/cvfOBX+Ij0dNLzhRMiFHmzofDVbbqUSZSnIX/EE4qBYrITZYSkz7t3F5+au+
gfxYA5ldxy3H4zQak3TKDum8vLDdoELjnZ8IYuA22S7+sEkdELwusOrPq50swQLr/rNs/kswZiZi
aA3gnJifcKO7WcgFa7KcoMjb6KCMTOLJpzLrA9S75UcuFdbpOEhlDxPxIpkGFU5bWBgLn8HL8LdZ
pYByogOo605u+/kYm+RL+XKLe7LgfOW33XZOXP6DEoE7WmQBFMyM6w0IRb4tUgX2S9exHbikcKxS
EhgxJvyQl8JbXnoR+WrQaSvlS8rZQg0pNQm3J9zWfnsAn2B/QfAHzRJGQDB06oDMvte/Ga8k3WkK
ee3twpwmgUfaCrpZAG6a7BG8kKynl43Ymu+oSnqH840KAVakFNHvlfVxY5rb3W9frNTVL1/yuJzL
dDiMVEe9NCj3ZOSe73Gk7Yv+20lL9och8GjdeTqqaSfiGxMMi9cuW3qI7bKruxfmRjz/EdgtuXpF
nt6xPcgfQH4PY1fprg0NUHdclyw8Qmt+oqX9BpQj0iH86sKOlLQ0+RkSk3YGR6Z9zpIJd9W1rOCm
oY8ENAoda2FT1m4rH+BUJZHKW98MvH8VQD41rxg+boG6uKJv03RSeltLWGiIL/AaGohen6M7XZsO
sUwhgr4qay+qstVNjFlWVXpqFpaKMo33oneYpW9d4C1y42hnAqsIbUSCkhQZ8Qcl5HM782b227jL
iLBNcei59nS+Rzp4WQHX0tKwSLs4z91CMszlRsUsL0N6TdSDclQuRLjKhYB2w8xz9gt0zhZ3rcde
A12g2+K8+i1rx5xXEaBkag2ubm2lNHSfSOYEsT96bQRaxwnWB9WHqUDuQcZQ4aMxU7rqeuLMErWi
0b1DVCa3Qr83cxa9utFT8VhVzCPiEm05C9zDMb3PQdW1zbFIL2jhKK+2sDEy4GTxMQ5k24MsSZEK
VnwRmp/nRcPgJ+tyY/MjyJjqVVc40s4eeUzqFWdSINX9AHW2hG5rDHZes1kpBrUpg9X93VolL1s3
YtREGBqFGA/+HVHQuVKUWnvNEH3Q3UikxrfBhkB8aLhAhR4IHqjkVq1U25LMHDRWVQhXKFTUyFND
QeqVvDYWm1diclHwbzQ8kYFbL6D+1uHlERaFlP/pBK1e9PYHarB0qVQc8yRzT41dHPLPjXGM9jdW
JvCtbAwWOXpEd+N8qOTHhbE2DF2RbovjeJXp+ZSyY9hyiQFsVwE9umU8SDf3lH3T4o6sdtn32K3J
++/hN10HbLkTGnVGgSYiGht2Hkpt8maQHfdwoP5zgiHCDpPO4IvNEWZDu+kqPEVVAK9/e+7HWcMz
kXn3y5cu/GUthFpnfMZY/HP7981T4MCx9qYTonpm590Fl6291li2S48k2KcFsq+F0KR9jiNuUX7q
09Fhsz0Q7CbkXf01gsJpqOCpUbojf32gkkV9k+JY2dS9FHWGXl48TAaf1gPkHEGCzY7DGVMZzt8X
o82ju89wqhQvRD/BouuBQAJJrPDr0xHdOaVa1I9tkZTlnQZ7GGXepaMrjvv8WnU3IxKSkbE9BGzD
GMUJWsKUMotgy+UGKOK0GpR4t8iu5xq36qPepaAZeBjpoFSMkSROTQ5OX4Yqkyd+mTPtkeMJPTgo
kGJeanSytUww8miEtUH5R3PVYUfQ1/DhK7zyM1K9kdgyUxz43pCTJ2VbZb7fKvPHNwzjcq+t2VZr
R4ME+n7cxPcMJ3isPBy/WWCKxiRKKqbnqhfXE08CescDz4t7rEyhmrr6Osch8DMHCc/7FVirdvZq
3IHaNQCEeqfwZAF1rPXnOm6wfxoucmOjw1na/Au76yLX8f89rk31lHeGDXYVVfjnLzSXLGqbB8Jo
B6QIdVbg7yb9VOCyPlR5jXgmMoMjuDz9OU3gyW5YgEhsDRDJBNXey0u8DhBIxVkKeD3iDcSxH+Sa
N3sXsIzQaAnzl1Gn1iv7XBS0xpPaJt4Q92d/N6vaJMBLQBkspsmAne8M8bjTRCof275nS4xjj7ea
VChX3fMMMsiH70cuAYi7oVdDn4iadVzIZ7xva4Co83FaOsdanL8IApxrp/S4kF3Z6xv899O5GQOl
BAxrnYpQxSRE1PXbJXq9nS0WD/+eH7jDVpNY6L4y2hlHvSWyAFeoh+hKbsgS5LSlqYerVwglTSka
2nTM1Jy1XOqRWHMgNm9iFCX2p9YxryzLSweb7q4U7Jb0nbTPGPSEyli2o2XaCMglMpArT9X5JDbq
5B2zE9YR351DSb6rct0W2wBRQJG+OnpmqiK39jOOLgcDiJ14WwImy+SsQmobckrr9EtVyB/xYU7q
DlflzywX4RugVygch+ll/EuR9uFq2uZC77AhK7+/46dWjahYgW0kx3A4ybwPp/CLMiKli356R0Zp
oH856ZyklVMdL375aOjnb8DIlusu5NhxYQNlx9h7tEJ84Jw/AZ79pjaEierHBx9/8EhXdq4dzO7j
Q5RdPISTBcisY02XP0MuChUy5vZ+/Uiq79HDrXxGDyLr/GjCJDy7aBHj7Z98JyjaD2DkCqOc3kIE
AY+qqeb1gz0zexH9yKJ14j8OePuIG7kOj+F3TZlUCfUhHhWE18JwSrYvjRxt/FhGcNhkkvf4tEFu
6tvLTaEy6+fgTE8RnTp8wIj+8VdDUldHRacvyOwzeFln/S70zdgiJ3NVQrSBOEglwLw6Plq1TsgV
SE1EK1ayq3kz56V5sYwMagNrv6KimMNcJ4TGg4jJ0wcR4t64qkDtWaCAh14c4hpdRF3JDIM2arzj
3NNxPdYrKP8LwYnI0kpXyoppom1cYbtfOTraDeFlzt0z13YLKSMtDae+t6VJOGBed1ZtIcgzgR5h
GptSLWWQhjLqOjqwTEEze4DVyGh+6mXNPEPaggIS5ZJexEpZFK/7Hzxia5CYo66jbzfOSMq5yB/9
thNeRxAhqXDDtTJaihOEMPswiEqKneywiA9K32zhNKAKlK0e8AVPz6VuN9WvYnhw7IJ3zHtZS3Bo
gnJzJTWXCi4wMqyXZgVrj27YrcJE5dFcE4k6uoQzI30s93LHVZ0aRHwKZykT4uM07iFpnRrY5CHo
HzYvfcJlyqI4gC33wq5je1VFxr06A6NJHdEXJJoSqmWqGev3VMVi8uQCYFTK4W7ygvzE7iAnUAPQ
rCmeLUVvZEPgK7wjkILoyLPSaMYAo7A/t/PgLRNyPZ813Lf2lWEpfoPXcbX/m9ZoQZhMT5UxfVVZ
qBwuOlPBKTSP9gAHPM1tLTzsnLKYHj7MmHP4o9BU70WACruAaSBxrBvOsleWmwzj1+mc0hLBqZK2
g8FETk9PrpZ9kaj7tAygAkHFNH3bC4sgXuP7LCsrFJLFGQACPOp71oPMM9RtQvzVYiIVFygC81N2
A9luFNVhCo4mYtkX0p7SAkZ7GQm14daCpxB7+3fr74y+kPgYs6pLxL8ADpr2fQ8lONI6wEsd2VPl
4pC4DWB9eVDuP/I6cMCC4/IZEj3HJeY3WnEo2XDn7ozjd3LA9JnjbRRfddqxEHlZY3MytMJdGyFJ
CQs4RndvtQ+AlzpC+5VnuOGuH1DSr/DWhEkxQAE16GypXcl9Kp0uLKXsRIoSt4wwxVwDKQn9qgy0
T4t9YJaQF9JoRv/vUnowJo1WuEUWYdHF4Nj6EBRi5ee+cVQajS1abRe/Ak6jdafkea1UqovDP7SN
tGv6tAtQ79bSj8Fuu63WGpl2/vFsC3ELF9GiPUQ/d2/ckCrYwsTECNplzzQAYjWV18F2DJnPTDQc
VRP9XBewR3ClShP6szTY4qgfhUNQ9mgWZ31psNNM0+eWJzhnYWdMRFRjpKoihxFfMWIMsAY+NAb3
wTPduS0ognMscq3MCNeq+BQBhufooi58jZuJzp48vS2UA1ehQlT8hsvZbye9+pZviDgHGD7ruPCx
ByubwLBag/KdWmELRDQgRW4/oUcuXLtS65J5G14zu5r0W0xXDx+pePYMGKl+Ow4B3DQJd4YG6h/S
VEwopZZDGlHiOn/ThvBmhFH/72gA5Uoc2+1bVY37dO9qIM6mXge0vBWsoEgtpTvwK7mLSb0M8DVs
9DEiE+ZLqYm84nQmSJmRN9bqwW0FkzW1h2VyhWLGt4W8PeS9wT5sAMDc9gv99dtUlMbBTe7bTngp
d2PPlwD7u2uKv7wsQA9mZdNTAogXrBX+YHo/S4m4ZyQLM85b2u4AqJYo2E+FrzWVsB843INlitL7
9mkzZBIxseGnkIYUPrE0MGSGEi5qMJ/XO91UtbQmqiKog4ok5FQGrMvX49AmKrYx7zS05u3NB77Q
ciayZZeEF2SRgpqZt2qNcTGus6rQ+M4TnUWY1ljme7CMtlxvRfcqAJR6m/7cjR9kiJ8kZyl/XkYn
gMp7NNx6un0W+b7bRG3/xDUH4jMbXN2WZZggRYe6mrDLFYwDr8RSEfzx9nIgxaAHTYzaMdH2QY/e
4pVHNbAZ5uZPKVKF2jIGJKox7vsKnsg5WqaU+VLuvyb3St7/uNDEA21zeyhwfI0TbkKOMqKAM3Z5
272sj1pnshqto0LuvcIwkoxen8sb5bAFr+1alEpaINXXfQLm00AJ7Hxs8yDAAnlYgmZ8fLScJ+MX
nngVlQXqbveXEKzCMaEUxqORKYVXRr+4OXn/uf/vQDelgRu04Mc/I0WFnnbZc5f9kFiFmM9SgaOH
tdfLRUq/H4cmNVZ221fS+GqKbyNOp3jXKDe4Tk9RbwoPJC7nTd9BhCnJ7CMV6wSsU2iBhKeWgzuB
YRceEBqmHdXW+uObL4moUvor38/iyOfSTZwPJ10PDPDKHBfs/sqTVdPcjh99Z2D7HFNxEn+k8zen
0ksUQFiM2U0SI4i1hzfhK9WJKzQicFrOj6P+ieUD7I/SGAkKMTrz1tihwbIS3jwsIS+YCX7AbkS6
ZYFXP9Y3viSZZsx3gSFrFwkwB99kzZfH5pQaC2DipJLPO/l+RL38lNisxazTVMBlfQ6cKXCWD8G9
/Y83GS5cHokV0b8WaNOy9EGKpc7zooc7qAOvVdlc/2g3pJLvlDh6KZpGlTjd69t4Hs0EWwr+cfGP
4uScEvkD5wY9OnLXvq2R4osenU4oL0w3x10loHiqgr1zqh4Pisn8BBWgk36HT4eDlV5YES5YtpIg
ldMb6hvVmAHlXBXpSerhq3APEdsWosUp9+mqX2/5De/BreVcbqvqUq+TPkJ9kwWEtjCNuIUff8vj
6FD3icjypeae2Qza3eyFMvI8GBQlYMvltdUVpoIUqPULpljpY+HG1MZIhKLjYt0heLEQUuSTrUL7
uvdLa6hBHuwFoqEnM3AZ+YClH+OyoXaxIU00bek7J6KO1bNrqTC8waEeUEmrvM6rGb7BYMHsTzSF
qVKl/bGz+RdLNTrH2y+b4Khbg+K4wVCHOHUGzYQGuT/BuSaXpXdQ2MYZ9ehkKPYeEoDgi9CABZ0U
IpMUB7q+aNmo4l2zASkVoikWVYU3YXkJ3S7hNXhTNHPO6qgPQH8btEB4iKIpwTpcJekR44CXVT6p
BVpLRY6QGLawIQ31bGck2tAwWGoGpACVCxGm9tbWJrkzyGDzsHTf1ppBR+ni5dTS18pMJfvaa2cP
+PxIQ4b6GWkcfGOCYOfV+3kvpDjqj7n2Tsu9ZLLWOWVsDHMnBGLrRpZXbr8GRW0gMNY3LnA8m4+g
IJUNV9nxJIUPxD9BTVdmM95eacXBNPG6MtHYkqybrEoo0iSJoA0xcezsSVrD4fXQX+JfekYgDivk
LCKL7sgqqEuXKdacRsH6okjTK8rcslBqRNDvSOGh3xRd+9bqTisgdCjZWH9QmoUr3rvHwHjsz4/V
x2EhGSKTIFxwZ9pciaT5JLZVOlCoahhoGx50MvTnKeQ4cOaoNEH6v5yd+LR0kqDxWl3QdV4Qd31R
zNQvGYpSMIQHsO4gAT04pvuz4DCOYkpd/+9cJCaJCaG0Pvgc+932qm0vySleQsnqZJvtHn7bobP9
T0LMuEhK207iCg2xvkP+nphPZqD2ToPpI2SxC1ePxQ5go18xtfLpbukwKo54dk8y+w4oKxlmCvNG
8Rtj/1ZHe9s/XZy4/ae6a+gHp/q0SXJwv+Zu1nPTzTIXQQ9xMcO/rrGKU7tsTK2aGanXf6nuaNaX
+Y23+6Yq8Txj80nEA9hqvZ9fDE7i3SFZZmmqGsiyLANeSimfLnXGDEzzTIV9iS5t0lHspnRi/FME
DB6x0nJvEB3PpyCXBGyziLZcnukfqOHblrnuEVkcMMI88/tFa4kY0tBPFN8b2Whlgg5FANsuhQDj
nG5QKPJpnXqwmn8GIHwHJMwmmYuTm0JAAZ/ZM9cTVEGFdR/isufhXCcCTNqvXdiTBIGSRa6+z3uD
jJv0NdOrRKv+SmWlfjq1B4ejMLUIzJBW+ky1xxCV86Q9264GK22mt64WqwIBCsDplZeneE9/qlXL
AU6NoWlO88LdOmJRgefj8ER9UDeLeUdaRitdqoZUB39rG2gm4bS+K/VFoZU3OL9zDks97vAdS5Rh
VupAAXc+cl+jtHw8lGnVuA4epDY5jMEiIx+tvaiNb839E5SWZ+poPWgcd++ovgRGB90oJBzeKzN+
oMjHaMoDrSKzMBCUcuXz0EyLA/yfQeoAC2mLHAuIhaxeZTVDZb9BTug90rgrEux3TWe1l93vAdmT
SO6SDCSk8ldGT5c/CQ6+gykbAuS8uG24zoeEtLuljqF78aIuvXyG/69BaoBVYtplRZlFf68L+Vi9
Tw+wLcV0iKEughgpnesplVZkU6GS0kxh+llarn1N7nJMp9DGzGGE1Jn0bku2Zr2LuSrrjlQ8voNp
iFRKdshYuuvuDoAotJJIjvK/vXq6vDFqCeUxCMWwXg3fp7s4v4EbJ6+LXiC0NhqJzXcOgzxdo2SG
OBF+nNVvvfH6LzGKVRBTo1IUo7hgL80mUqphhEyCHuBI0FQcDTzHH+nBRNg2wFxNBPsZfKNyrS4T
UYsf64fJjnV+2RtydOSC2I7Q6Ofqda5ISc+P6+hhsNtWl3xYSYAWYzRaKQLTS+8wPqUKbHsusno4
p3QYlFfA8rlZ9EYkyQ0EiA77FvDoLdUUAZmot02wHGTc38ACgJCK6cfksUOg0uepw1bBy4qZOU9T
7m1wt4nvY9OlLO6Lo7Ahvxk+JtcPaPZ/628mOxbb39jshKeDAsJOUzhoSDb/mIqQRBmLYpYMwDuB
lsU3N+ST+RceuRYzGdG6Nz/tU0v705JjMHzqkIctvpZE6llhpL0eeAgFHWA5iyNejNTg3qrpjNC+
aPHhj4fXKxRkOYOtot5BMDxrMgu0jvA1G9IYzs6sxgbHaKlt2FF/XiPAoh8JLom3R7GkRaZN8GNI
PqmvMWLnJzZoce05cx/bOshVcescLOW4EyLhFnD6t64IUWYfpe2xUPNiTJMzGhWw91xwzp+awRxm
fnOf61/0VcH15PHDIliwmhvv0hM7/dKBuruTd/p6TIwxNSGGeH858/fo+7wikoSU52lfMMbhrMOW
GeeUKBAB5jCXg0kSXg4lz38h/RQ6c4Vtur4pE06oPB+mK560z1z/s+YRblnqiZ3YFRhnPmKI50vA
fhK5MEla6cJ7GhQMweQ4iM2DtmCkC34/Dt2bh2ZefqWUt0zlo3Bjf4LMzAaWO9h3c3WPgotYksV4
dZtiTTl5LkjErYGXb7769ijkBCO8BvpKiuabBB8gHOqwcTiwXUbLGit6UIsMa89bsBrF/2eIyr4C
/B2GsLWQUSk3b13KLMuS9rdydGj6sz4UGq86jteKUuR7WZf76NIV/OmoBWl3DCLeeTW5fmNEqZAZ
EG7RgxPo5/q5qOJGrMlaNpiQFdjseCdZgFBY0UxvO6BsiDc7oh4cuAaVY9yfKHRgP14YlhTtspVy
oOtG9DZPp4iEwus1ri7UWo6qjfejPL4GLbhxjmliLtbQh7U4gGUKHZo/652q+7Oa+J5gmU3xAn5/
ztpCGG1HOBuwBxGB7RSnqlHZg9g6na9D7wobKpaU2ckPfaFFGzBe1Hh6ogtg9KhdhdRNcND5NoVm
5+Q4/lq+ShDrYFhDvyDvaFIZChJ7TLbpnyRLOZ7K9A1u52qzRLSR17UNSWwS2MeZvniU8rUlX2Dm
oiSSVNWGCjtL/95cgs8RNh5N74kG6r+yxAArFSkuaLQDrFajj4AcSwxyz0TcSjEI67R+RalWTJ4a
lqOOxi17rhRoXsZOV+g1VZ7+s+W8gla1l7rsqTvGHOzxR57rLj55mZmX0b7pHxBSgpZDDO4C2t+0
sBmzktDRIYryS8Z4TEuDbYBKHneyA9RJBtyI0JplkqWpj/uKfYbdCXarjJCRP8T7PYipZHH+NsbF
NK0zzxdZzmvd0+LDk988IGeoHTuTzdFJJRndSdb+oWzfRq1WoSuD3lDLY8AAtui65LJ3XW1sfbIn
vAjXIJmWQWCuvlxixKpgb20YufZJDgAd2EfDQ77gVz6HF9pu5qOdKZaTWv8BGDS7PwYYc/QzU7Se
dpKLqt4hk2zfb0eXNdKG2MfS98pmVuiky3dgmryRMMr552IvLoM8DiA61W02LARaePqZORB47QPc
Nu1s+HmwRQlGnU/2FNSdvdfS4xZnMBbL91X1CjD0yFenPOdkyRqO/vAye1K0TgJMG7fMjvHBc784
ZUm1/BCLr38LwfQ0LQhp2ao1Kob2X/75dedQtXfsWODI5YWHF4msozI/9CYOLn6OcgmOGvWhl3JA
07nrsCplKH5TuZy/+k2snxz+MNcussw7uq1eJ8UrtWNlbKqXpKFv2GRX5ylGZJ+HigvIWx8t8Ci1
LF3NvKcHZky+MwaHh5iDfG4zxwKWNDgP2mfd/Ou1q3O2eZysdNqWRnjRd/Mba3AJXF87R04JvU+F
LBmUCg/zM/3CiJ3DEjkO0p3XUHmsikvRBTHoRyGGoLmeSJZRK9xVYF89Okqu1IktEWkbXdtlR1xi
29BOb6ZA8VtYvUuayHL9Qjt5NJmeWETEaTG0e2Uw0hWTbTjiIAmqF4zBAWZBKghY9Xxl/13QTzaN
8tyWZynTSrWL9lJSWGlqE8j7Se2UmDtJXYHzEOpvWU/0tkkTTOmIHzUxRI7T7cHugD7RrA/8MtTR
YMLGHZMs66U0qXwKJJ/hpXKIBJgpNkWeAPXEAg04xiRGnOE0UFFZum8c6tWrP5rZ98lpSbJmITcM
FFHlG6uhMEKe9auQAGS3NUwwfdEG79PsOsi+AQon6Z/l0Hi6lX9SygnwMmy9RxT53N8QjDn1891p
QK5BbZeRoUV9KeVGcOYSPd9PRa5jjxkv+TFAUpMK5DEpQ3Ed0LD0ToXcmo+n5xMTt9O/rmT3mNpe
5UM8WFFMvP4u6sDN1wb4hGHB1TPjQPwp2jgU7XvG6erVw8GY9K8Y78y7IXv7s4KNay52MEclVyWg
+w3ie7zzWtjruwM3AN6v2p9G9OwsMo1wJ3C8nN9eTg5AX26lgVyo5yGObKQzaeO+bB8o7h9HuEQ6
13IYrDKT/w182Qnp2sQeUNgO8Gl81Ex8pz3Kkp4mf4RS6D/5/J3mXkJq1K6mAhJLpfDpd5e83bc2
kZnLjRKz0RbD0zNNwihGMUMuTMSPh5pEEExAZqP0Nwag1oJ9fIjlLVbf0hC5dcVref9Ln3chPvwn
Umx/SPb89TsblcWbOQrCw6ai4MRN0fxXCsZY2mpon13CkggEulo+dccdUdCt5b2++28Zn3YnEo/0
8FmhZovxm3k1b6lpeObXDAFhk2SvGpp2BSJ0TY9I8ZXoWubxc2IBlupLSKRYs4nHmNeMBAq0gNID
SYgIG2/kwTbA+duOoLZCQkPeIZBDT9tJNHRfOWjxJKMSNkX0t4HbTac22bk/kGrPDAH8kAwOj2RL
6i3tihfdBzG2Rawkx267gObbUKyT4Og5kMIfcKdseZ/QQocfCi9XbR1L2oqWX0X5xluwzP/PPx5R
AZ6UfI1QQ4MHYtvvlyyGah8qOckzChpw/JQ8a+C7H/WsMjpvjVq+gatHgQqxgFSD2wnSzZP06s81
z90mf0gbcsqyyh0rX9+WuePUwe4FJ0zfbPUidumFb3LffBgPk8ebzfMB7KQyMR2LdI4CTNhn3SXT
aKPYzMEIhNwvsyf3fV410rERMT4DS5SVBK8ObRa7UCZ5j+Z7xcfw32JEjeqYyrZHgSTtlONWmRRu
UjNYvc1n2Vs2ngsPJGI30cV7JZ+654cw1Mj+xVEmqI3wTF+hghV03y7gopowsN3LmQx60i9BeLk9
kVjGyIWZpuwvm8IDAAhJf9xg+twQ3Ga0ZysZ8hlj04Pxha/yanAE1XzfqQx3cJEwecZ4u2aXvWR6
P/pb0NdkW/qP6NjY9sAzgOHayPpJ93BWxKqVNWaOjwFXF58wCuQmGf4X3wbYsLXvuVNiqJEz5J8q
wBE+Z10fhaSciM1cq35fGgthtBavYJqUUzXQpVzZlHqEPXVjtlsYT7VW+4Xrb97lVbN3ILIlZoDw
2HogozdZAntf6hPSyhGseL4v5FC2tsv8bj68UDntCohY1Pns5DMv/ynUzczOggEI3JysO2+8+qTe
LaB3MRFJMy7eQKlPPbS2fojbxD51Uk/NhDn7wEQgXGl+vZaNzDwrLsUZjxmOm9dHzfjOLIIXDjSN
mBeMjW0xwCXJp9U67/VSDXOCMC0fOT8nNF+UYQP7PAFuSbKKmwvisSr82fu46VFvMz434Uw9NAS6
8ao8VEztsJMAxEQJIwaBq/QYc06GhmLLVO1AsxssR/NsKKRsqMm2bCWkDqM6UqXY/YgXJNjly9mg
JnEkKtmHbmWML3zi1E9rQ1chvOgdEVLALx/BsIv3Z1fJMcLj9i2GA4VPaQE5kgWUZz4KQTybjX3b
6Gcg8fumbe3sV7fjiWiel4bR8In5PuLIhVrtw0yorYpilfvPhqPGmbn3rAbLdeEcfetPO1wA1AFU
OuO1DiSTIM0LjmVXRCazo5i5t76CLy7YkafONEU7jWEsBk1buyAloNlGzOCg1wNAJQC/medaYkE9
WhjxX+lb+Q7IQONdLe4KVIxV3p3m+hj/aMZimaPLfqjZYT1l7N5CTzGRyNtfUus0AhAfQJ8ykuoV
wTXkUhB3XXHK8pxB286xXr3qRKMVORjvWtoxw3xSSdu4dAIbMKUtN+U2hwbuHWjWqF5DjbMHf98P
qd66E2z2op1b0KmJa5oS86GTlreHA7EnbHRBY/IHBChErbkP7wZzaxAKvhPJUVbpwCfSYx4jyTfK
AtVKkt+AZo6o3H5StFPzI/OzoIz+KTmPDfh/wHgR0QgzxyVpuVeip0RxKQTuIwSGL4QkPt7g+A9T
ypemwuPQCu20fwQ4s5I5QzkhWFp/1gAbx+9XMiYbX4ExvgQdj+RNL3VouyZQKUPw3dauMg7KMFFK
c5ooqJRnIOMX5a0lnaVo/i1aNXZ8fF4FAwP5dav7pknhVB6zGrBsAkRMUMKaYh5lrBKRPQ/rlLTY
eXUva5Rpsyn7ZkExwVGuZO4jjvPPqjrhZ/VjEPWGDOHqCqFgt07rP+Wf/ki5waIm9Rr2PGxkp69f
4sryjFA/pUvBY7ngRKQvo4cEA/mOt/vAZMH2OJ9RI4elRzfB9bhSqWBcXE85nWgnICUZvBcTuhI/
OTqFV1BvHSzlFLIRgSdvci2VnENuRuQEs0eI1kOpikRpEhV3AxriD0PGMNlkM494BErPmMewdyFb
4i3/UeK3h1WzZQMqAfGcUzYuMUo5X02eVGWG43rjaxSaOQx7KA5xdz3NyXBpLr4D+dKKn/HEadm5
Hxhe7Npk29BT0LXylBFK30Os+6vF/HTlheUIRyP9+/Ld1eR3sDR+gByXi+UH/vZiU4xq/DTskQyp
CP7FAdMo6BfMg+Dqc90xt3F8TomF3TETatdd4ct8+fAMsNEm02M1ZoztrSjdduzT+LZrF4N+lRoJ
ez2R1zBtaRKjxOV1q08z0JDuwbaodUwSvfbATp48e8EvC7hth0VznAHhM3+ZpFyG+WqTb1Ad3a3s
U/2wECHEsih6HW7/RZJyW76qf0LCwdXMlMVD8QPRT+l1fL7tnw3JBueDdokgidbRjlC54iQWxlaS
rcTHzY3U3sCbTu8kRuVkCUFPDpiizanRjGWf3YmzPBlBJb904daFgwRXjlZrTD9PCMKupjeuRcxN
4K0Fww6rXeNvgzhv1ikbt9BJ4w/fe6gHEwpdGPSBfH+EGaNi7kqNCHHFivNiQ1+tHiSXRz77bl7f
iRft0mAi7HEw2rzCepil8v8moRumZIkqsghtkBXmmUwaBIiCAYWw9DQA6B/x34L0cXJSfFBD8sqR
FMXzUkJ6Axxb/zoykh1lqicHTCCoHhOIXMYqAvOsV0Yr21NUeoyQKppQIPS0eVFn/Vy0V5/3Jk+B
+fne0C6FMqSYQQ+LvtYz3xUEMH8n0tgtAXA1IUS3WHZWWtRs/9ZROyRWGlCoqhhh836SFM7Cq49i
u/tv0MUQUxDyHuT4Q/2HQ96DivyDfn98Htt/G2EL8IRFphnA/dVu6LwoFET4vWySlcGxysBbgiHl
oKjuntKX1CzcjNpoT6HcSBZGMzLBVXd/0YhpRDsERqEDqOSn6S/2qnmNSXKMK0LKLMI5OysHvcOW
BY0NXXbZ2eDtErIzNZcaa1hvqholw+87pyr2ePyLVenAyiWd8Ik2wrNfh2pvFyvQIcoELivL8Nv/
ELC+e5OkyPhGmRM8NSt1OA/T9vYLBe0fTOaU5WvyhagV/EdOkwEn4DhaM1kzn3kfmTuOzvVa+ukm
XToGpoikDeBLX8Kg5NLH54W64zWL9sP8pFRtrkunlo/vXO0R3Lhk/RahAlS1aYS7nh+zFO+deKyK
rkjUKRpSb5BMnhSFZ4q0gozSSur7/H3I9nPh1zB26qOBEFTQj5W6gcCCCsgt7vFbtmDUyuFPLxBe
saJH66DWDW6DdVX1tStAGycw7ftPFNhgTCrgeQtT7v5OnjoC83PMI/N8EWWAqDAvaNJ2M5pW1qeg
ewJWiui899mHRt4N/EzkQT9kxUwciKsBf+QYHp3SE5UyGY0kJP84FhE/oWjKms+UweqHCKDQvrFl
6IOXg86cQlC48sPFLYpXudNZBxw49Sy1SyY4JtLwKf6d/Q+Hm8m+mkZRbmi0nUR4i2v2oeyvP7kd
UYRPF5fMfQZVG+GqsntM+XlKzX/JwV0CnjkFi0R+4yqevxHSRw/SRGMUTmeS8dGTha9hI0yq6oIV
tGfVHi/eKwd/2KvQ13IdWM7vOcyHejYDeenLc6C56n/hgxto0WvOM6ffq+Kv236vMr6fLSBD5SRA
fsWXmguIM0bbu0p2Gkuw9zggKmIM74iowhmI9o2wJKkxDc9EAfiB1HNCDREPRUyGu+WoiRazbDtB
E9+IeAktLySfeKi2rZM61Qw4ecgLtKuHBQhBD6DLlqGT+oanqeU0Jv3gTB247vEwF1Sai6CP3rp9
EWdaiat9atO64bDbL3YrvpaG4sQi/Wu+356OuuUNpAuDFe5VAY5dW+3LGkK8ILMrij/vxAvljxHH
Q6KifKtw9L4o7JzY3+Qz6KdvVeOyuoeeWI6PeF/MQAJzbp/l70Pkjhxp99EbylBAIuOrWSsoqS65
Dkyy/TjQMQqFzPSAMG0Cvz1+hfSLuIiSK7a/zwoZv2ndoDV+9pkpGIbrBKX+fc0fineG7WU5+Yp4
jZVuuy5+N9tzpDsaBdhTSXSOLFTA38SB4SVyHM3n1uztvi0AMF9QxqrMYW7x5ZKWAtI31RR4OcSO
9IcHrCqi0dwsnyvNoHce3j4Im8evIUQXXYm6hlQh8DTW/28Fl/J1Kc9fs8YBys1gkdDRHdy9ROdV
jNhknIY58R1KawZhE6/F1GxlHSmLDkoJKMl6EQUKocIl+3GTb6bXndvVbtKD14mslel/PqkBQd9/
iB7xb+gozihjBsC3vlWYj95zpSvVp8ACB/YDtPVeqeapSbjx7q1o0GjCKCpfVIVVQ9xDuBkHKW2g
utlXAbKE9Yp0hTSYVHhtqZ8d0H0gN5B8JYvPMom9AEk6rpiZ6r7CumXS2PLoFT5kRdfAK9nP/7OM
lCKycB5/vgQ/rzURkA0i33K01wb91y5YmS9qbPX3e8mA6tPXBe/PrcnB8zcKUfJzKY3D9UwP5C9j
hRKtX/a5IWiyPhtoswB+o6lbLvGBxTULlBC2k5Yej5qdLhhwjtjqhMJvhIh9is5VXsgPtD5ZIvjk
jktSFFSpTwM/m3aT0kvVMhobam8bSjpeBt1D+c3PrtDD43mzy0Ps9unb0EUywHgkuvvUdR+p7Et0
KgiBHmQufAg/QKTvFhDqmmlQVjjTE9vN3xqICFROnOXhojQkPic27hUV1WjuG02n0xBKbm+mqdjw
8qf9qT7Knw9HgfZD3TVp2fX8fu4CGzsIFsZW/9GqzK7wETgShTUvebpndglZHOZEPzbiUYURbhJQ
pIFbHnYOPESdUlkOWbA4zKFThdYf1u709bwS7S0VmIrjC1X32/iScp3i9NJpwfVFhpuqKouMYo5I
lnlrcJMcC/zCyzD9o6j16kYvJui+QFQ3ya8vJ+2A1T3PmlIQBxRxEYM51fi8TfHL3YkNLczrq1gb
vWVUv8VZqRxxn+LNHy5ixehefyiiV5ROAWdT/lPjp+FyvPNmK7pmE7sC5mxuQUXWXJrphZp9stVH
8hdo7BTxWYwVRzlVr5b9n5mfJrdhz10KPqJtB6PlFpefsmWOQJEiOzmsOg/4I4NaJ6cZZa4v/UBO
3yYiMvRrO8RMIwU/6PnO9xk2Hw1vtI0x98MhsHKekcyY9qU5ff1unfwwhCWhic/KO8dKOY9chcgm
T9kUyDpGxe5sV/iuC8EuZWT3j8yDOUchzrB33NjNYqUW/g3IMXIJigdQCNcTX5XBkEDQ3h9dl1hB
hx76LQWTy3+qy2tSsthUTgzaruhoVVw/tL1FvoeWuewUHw2Zjl9JTJu6yADSjiu7d3bPTchF5NmS
wdtvKJZhzPGDCmQUvBN8Hl4ei6K/WcVs5o+1WdbqGItCyDi1dk0369qxWx3tHSpy1bZ6fc6IzFDw
NyGlHboif7KZXCA7AIIJuZ//DRRoQD4pOOmZ9Jub79NzH/Ctz2HP4d2H1/ZPu67gX87rEoeicOQJ
74xiKQLd9GdUtj3iu+qFmcrEsjNKexNvStBpXTs9yBzhojOHMEVAeY5UvlApZBoIkqMvunGL415V
XMNsFZyC17FOIdcAs/gapiImxI6bfDQUPNJtyRfCHUYGideKO7tDVEwaX94o6UGcNyigvp9kh3wK
MCiyzD/vtV5zeCOUH4u4H2cH2zZA2yh8HlNxjWb3k/3H7FhXyFA+1ItxXR3j5xKAmdnKSj05uYNN
NHOYpikAkRMCT6LJRWoLC5IszZCcUpnQXOCGv5kAGaR6X7rS8K+ByKd++zzmljCtar04IZY+8Sf0
D34pIPicoC19aFuryOzABrKwDUqVIynHTIyF2K9QqZzHd/RkWlnAghtJ87UoaEWg0GnrssU5A9Ae
HpI7BRqw6miDXBNWu1V//RUznS9+/shV3rZMy4Ef6rruA9Kp4PCy66lfEmrky2a5CKelarFBqtkp
0MqYIY1JV7rfrSjKEDja17OQQdqzN7L7i12NSDnTddGysXxG8lfKzQaScAwzbdFRP4honh9KBK5O
RXdjfrlC4dK9hA/G+hxYlkQCKKhIQ4kYv73LiYMDqecovUTJoOGCCEROHqlpvIVmMgOKWafF4DBB
EzJjKLv2GXwizWZnBDEZODGeKbmdJ4T4ZpqfLJFINHnlc/+gzcI05BYxGduTCbYoJ1bPOXXFMBoE
FMnryuXzOBOzOxjQr764NxfJuS7y32MNGirURApSxWcZ56o3kIVGUaHFNZE8/F7xRRjQ/r6o421K
xJUbFhJXmz5m0GTZcElkMqd093ZOXhhxb36lSzcoi+ohFg06j2Hs2YAkGm48E5qprph+oer31sI6
4SsEB53K6NpGDBl5o77ligeatg1hgRG8QVeTBeXaKVimre4cRY11oSFO4BmnEGy1SwRP2jv3rU04
avsF02HucsFdSo3Lg1stMNaq+55tFaNU0aJcsMf0Ln1BsvQTwa0TaGX+5KXiUAaCTTBn2lYQ+V8Q
pQSEtp43LBNUS2Z+MjWvD5KB9j71uv53rqBxcCC55XQ8My0BgIcilr8xSF8gQbf4Ie4XSyVEkvIk
IwwOdOLHdPXvu0mCJWPqlt3qWd5VeTzcNw2C1X7OM3mQ3x+8uEibdCT2mG51wSiNoew/Xy1LF36O
Y4iy9EiUJ9PG2AxwQiYOxHtEQqcS2EV9HCa+/tIkBg6BZ6hmqgCEETnh8vNZqsotTOpXGTbSO87a
ImRV07MbwV9nASipHaotKN2J87TG6O8CHSLCRp85pVno0CGWohjdDL4AEbUruJNx0NqOKZRGxhLN
35AD/Yb0XJ54em2P8K8tL+/JWgfR/U8IuwdZPscrMiRNcxQ+Fr7v5NmVUpcLtAZJHUFz6sHY8a5F
NDK9oh4OlMG+g5wfzSi1E7g9DYasj/iH+UGUiHVenZE2U1KbzAH77kYUIH0b77VGWeIhQiEMSNGn
KNL3Vla9w+zPFdcvCI0PE2svxO4ISOUbKDuADWdDwGRx66xp2pf7uYV94PzdKNXH1fJUs6EcB9cx
UTVue83nvGni39oitqzNz6LF9WaGEqP8OIezeH0E7WP1KjalrW8SqvDOoqd9aGRxaymER0bFBnrf
ezgkfKxlifl+16p+4c9vMoV5My0h+0TSbFiCJdjA8b6jzt6cOv+HV8a0PN59QYhLm10/f+KOgAB8
uDotD1vaD6As11CtT5IlyT4WwrUM931leSf/2ulQxrs4UjeMYTkodERct0rjujUHmYnrOnPTTjVL
DnRzjahXownKX9SBmoC4jJJWSm0Fb6saXiY09TLu65jO00HXRKYwCF3arRdGt24vPSOezirxKDM3
4yzejl3RYeS/s6LYUQsMuHuLBNpmuaXn3T5w/XWXjhmojXRz6lQryCrrVPC0dt9HT5QeKfY8o0ax
BzAKF/oUskChV0vsDU6r4si/wOjLD7cXUx1MEj/XPr1zAQPihQdloaaTdSs6BRp9hURu0oQG81fi
vdS2Ha3ZaICeHDaK2F/HniBD7gg6sdPDyk7igGbu/foeMecoxMzWUfxgEKAo2U7ajZiFn3bW9pic
S4H1JTJMXebwmrChQOobMjUpcGLYpVDtkzRxvWiGmDVRdaJfc4cLKSIaP8NjSjIgrIP2FxaEITmq
aIPTfk41/1BoKnP1i8yUHjJb+Umu1nQkSAPTUtHhc5GuDu5V7oK/fKjVNjc7Ip3MARBKC3pnXgnL
t1g6+iJTNpwwFfTOC7+jixlm3pjItDPuDbnOgPTMhfa4ucMRNlu0QHtLJtywV4w90y9TxteGfY9P
zSGySxaDEmP8XhcQU2yUHcykQipwa6sZqFXXByVtAxfwuh1qUVayRcEr8DEw+ju6D264AH3p+Bp3
Eo+urp8Nfku98gnvnSkWwlhLt2MGMoDDCFFm3MpwLNRN00DncfBN0qRsv8SCBCIpkGhugzmwIPDj
bmW3XC/h7Z5hpTA8e38FJ1FzKHAPtxXh7onI7JarmfsazL8Y5xbJ/q4FRX8tFLEHRmAmZ5N81LwV
EHc8kjiJ2OjXrO43VJYjrd3O/69fM+WIgb+zQc15AGtWv030dDuPWAfE0U76eypi4orm7YlNg+D5
YYO09Ed+pmVAqUIKLD0xhIol+O8GPivzEPmf2SZvMR17tuOUduzcUqH6G2YEkOca2iQufejw9Zic
ZESe8RDEVBFwWyj/Ys64R9cG/eqQ9uUFblSWsRpT4a584FntgCLojxME5Z5XFrZ2c9zFcmjr+nIP
fScAHaKY5E2gg+zrBLltQ5Sicspmw2nfOY/VyRM0yUNhwpjiBgWVCBuKSi1Zth+rLiViP+yHX/bT
FjvcpV1kaVKMMJAZUae1uDekXrSUzYzG2ftNEQExJk7dzqnuJHwv/k+/wGMGlLkfMfzAt85SuIvE
TqRoBsem581OfjkS84G25tjiMwHe8exXD6N6QlAhAVmcbfchlAjEGQfvfX1TwK5MCBpRuOtNVyxJ
XDNiYpcJeosngwNIJLEzm+Tk2P+dzsnCh5tQ2PvWdoj4dwbj5mPkPdHZ/feXFO7HvrPproW2wTIK
nNhIzI+dQKcWTh7oj8XE2hWalOVoerdLl99TUlDnJZYW1dueLzdhW7ziDnLeD5KSrEibjtlfl+cd
NzUCXhipa6mNK8UdbDAc0/8YASHmilxzooQ7c0SGVB2f+ilP634243DWHcHhV4eErkYORnWv8wUP
TWUMsTBPHTN9mGfllqJzE93F/cczNncpN3G5BGGUhAU6i0j1ff1LUno/+09DqLr5nl8eyBZB83GC
+Ljy2AXUYIC97nXWSOG6aJrCB8+dZYz2RTVcEtxpNLDRk+6zNyfuU2NiMxs6roKpi6gK/Y1cAFgL
2WhmCv95w3L3q1CkOohl5godJpoozVtJkduUb9R+lf9BEKd8saEiV98LAwz7jXHHU7FdFZLIUJ9m
ue0jKdbp4fG/ICKPPoqb0Shah1DpHDpVUYLkVfVgqpwOUKEp8gl8eBGOVrFE+gn/9s58zu630g3K
QbdYOJHl9mXAzVii8DxiJ18AtSjAMHuVcpLlqL3XoKBrN1EdUy6F/JRjjl+KL01G2+k8Ai8T7rQ3
OQhQ+HTddk9HtfIN4XbPn/TmBbePqoGc5jzY7dhNh14IGLUrHYj7bDzHzbp+Fp5qUr16qF4KNP3J
Cb6WwDcZZTMkEPzJO1YZQeIqzSAZ8G/fK8MtwRxbHPthJ+tKHGC1Uh+xiZnT1Ebq2oFhbN+OL44g
VkQEAxo1Dfd/5+0ZR79xqUYixUQG4XUXFI8PHRXh36e8VoRaoAYUhyJBYg2eknPQ1f1yGTnMwPeC
jcRwfm/GZ/x1onafhFtkpR+6Soapxt6/wRkA/hDfkv20q+koAgBmF94S7RV5k2zzz/8Yox2ynmKx
BWNRtDLwxz9lJTyCSqM3RbHKRTBbdOsmNmVtefRdQGPIQpfT7GENbtKDZdZZl6O5pCYE+g60QB2M
z30U4XkJL09Pd+ZkVE1LMoDJQCNVBfAsu9dDBtvRHHcd+OJ19Tj5Aqqzvspnb5QNnYXGU+8n5JTE
FC1qk75YGMbcjdQSsJA9xBUqPXowuclEhnioiyN1KYBNnGRKaediRayle8l8x9J5O1F1ed55JipX
wlfQkP2vS5xUtsvM8bKW8xRNRJMrAPkSI+Zkh2QoYE6NDKLpanGnowm6aCjrreS5WzcSSNBXAwfd
DaOfmq8yjfAe2BNoUXDXAL+oJgbHfdTL4uU2+yQe2xEGs4028zAPzRRHladRkv14IzHXVUeLZrGA
3Kkla1YXkDySlhlIom/0BRTBUOs2Swfl5CUMVtsR+Q/pIyDUJ25X/Txd+nHrJu1u6wiYg4vLjHYb
ZOiQL/ZrIwM+WWs/LJdfatei4+LxGtXB+6rNu1cFHxK7TesrOPMQnaVJP0Zi4DlDrdGYr1jthM9T
J77mE/bL9ICAa6JLaYHwL2EoRDj9BK1+5GWI9/tyu1PTc/hBWJoLbLa1vCoecjXhwhM+TmSDh7BE
VV/SRkqJFeIfzrHvSRLOoIxRADeO4+OCtZ21XlR8f0AzPJi5vjQRCapDZOcwLfW347lFbDrcFf4h
u/PWBihxPF95UuZSLbHOL6yz1z1+nGgsQsnBYc7bAk2mJMj0pXAUIk633tJxPeRKu5JKkRDCAwtb
k4+fqwPX4R+slcCpP8V2ja11z4kMrqbMiH4Rt6uxEhfO5nq+o6uFSSkF9MEIrk6eF0EzUldGQHTV
5fD3pOqAZDdO2KpvfxlfnwswUMiRoE+Du7AEhepdKJz6rhJPf27lB1BRlylPx4CDok3+Wztn95hH
I/naetnUo4g5gk6rHNlmdnfM/bcdRBVMR3VH1s1BOl8VLPTUKYPZbKRJwb1/21O3d+HeaADtE6lt
Yl+MiI+OjgMdGXz/Aga4rVFgnm0e+F8bb2bkkwkyObSwwGzkKGclzG0D5S2wLaqCLd3dH5B1M2zt
T8MjZY1VIernB5awhuaOATWMUu+oCMcz7s0iP3m1E1eh07AkK32qsmJk18Ofhq9rZUytz9lK8PD/
k228qcWNCghjzBwH8R3K/WjvpydvYf2lAiTDAAmhxbzxK33BFb7IGg42WWLApwrEArNq/XtsgpGm
pcCaw2JoWhG1Z4xqhRo22gnxoYzA7uGIg6k8f4kJFyDooHuqo5WnRai6Mv34mM7gmFX86VAIMJZx
iixRPWD7wblX2olFr6JZ9zwFdGpXaMx7hilEsiq7TSzINWwDk+U6i6yW5ubNFs/6iAQ1CrQ6hxt1
u6QOgwJfpjYXLRHWJga0TeyFN6Wt51ox68Qij1HCM7/hbSCGfhVcsbXwUF+M1sbyIU99rzq6zRIv
ikjKwSpgfXBDSWdc1m930DXbKxV3t5P2HAgNriB6HvOdHTLrAgVMFSLgnhPlNTKkdhsLC/Eih4F+
PM2Ordq3Np+lnLxN9WA4QnrWSrFuO3mDeTigNuD44yD+/wCu5dKyRtqriRsQV9PmxpdeL582a6UR
mXokDr0zKTwA8CU5G04WMV+665OoyACSFGDb3jQJhDtzGh0lu0fwInAyg4f8Sgx+697mRkNCAyCM
hlCSisfJmGeyG3MNLzX+GXJvoqb8xBwLjcs4Lzp/fVNyfytHaoajR280KTd/lxY6WK1yVArCMoXL
OVmykQitKjndbl1oe0FcQgJ+WQy18lYGWBRCAuCCqCghQHy37AInk+RzXXJUg5cHU0Zi6joibGav
/8+OvnB4Vw8HJLUZyKergSlvxaXwJif+LKkrAXt7w12bwV8VbQvU23d7IsvD87P5TdB8QX0A19cA
jTBXCv+Vc3cMy+oK8dYmleFxUNyzaY+0wF3wnEK71maekyANREeYhTWImZzx//QfwxKQ4uo1T5YJ
W/dobipgq/6eJ+YhOBCDOkHBibG1X6ToogSicvOBkDxm25+kLfV3Sa5jNmWAdfXVDGN1Z7wWZ6jk
/y+OlG67TVyvm5DngLOzOjGSpPxydf5wNWo1a12Ow7hfOUbzvkDhI5FHThJB39xmSYU14FNnDKwR
7Tk49JvCEm5OBaW8BJa8RG9ur2tZOA9LW3iV1O4XqU7tm4a8yuKU8ZqHcWYiIiUqlksbUBu6QfEc
tOv6F/f6kimGGFr0bggAiKOtQxg2ngecJwRjV0c7DFYUd8VtPQTffC1V9mQ8vsCuBzz1tT25roU1
53kTdCigX3dyy+8/YmSIm1EsXduXM47jYH5nuiQ2Y59tlpqYkNqAmKWiV+c2utP+4RcUWzWVGyA/
UcUOEhjQw6MWymI5R7YmcmOweTGGM4gUz5uwEzXfZ5QvXp9Bxhw2qmlUAEhaX3rCUi/oGwyOtv8g
Yad10s7F56jdO9q/zKFMXqYrCLzCiAPGaMzJuOGuG42WX8q9kZomGgGBP9qd1nP84h6FJ53cEVhf
0Q/YzZ2NI0mJsGEPPHaJgghiuMWmCRbDybqRCQxGORMIMSAgsBV3TGpYkw2rK2roJlcKVeMIIzaz
SPuy3CmwYtM+di3MO05vSSxjzQFad9bk2YSRli1wYgxLvgJxKtx4AWH9N6zPfKfKRCLakA7jaeER
W9R6tnXfc/KM5wI4NMRRk4k8LvTWnkTzOAZ/+uWYsWDzgLqdD41wa6We59KOLy/G8oT9OPu8PD7B
gyUuNcpCJNGlFlPJeMU8Shkn0YpqrFqRjeOKJOM84IMVpZIaxZWDCXWHI6IqlW9Wru67LWIAhXbY
TG+UkhPRzJlaD9uhyMbLe0BXPyJVDMlu4iGPV1ORSVHqV0ObuCPw+cJyJVED3v9IHgXX11/HWHN6
TbKNQ5R8MW38GVZO+9OR1XjW+nRBJkE0igM9Llw8ybq5dzDt/DTyRGnTvPCTjtbiY0PeM3rAJycI
pGaARrPrr+Vo6U8Pp7EHluX70Lh6RlsO4kCAYra+bVOUNc2erfPdj/sGGuhCyvU7EmaKT+riPLEU
MK0YpZ48IT727F/tvWeSPaqJBTUdxb7g8iNPSV0Cp73XYNZ7IlS+TwxqrPoM3NzMyEBhbJPx4r3X
piGzxn1EVqikq2n4xIM9yxjdHpIEIjQmm4OqINQ2j08iztbY2KwTGldnGuVmz3e5f+y4qz/jPyFD
26TVLlZCFJrJnNeodX1z+Hmit7XZIDefe4V7TzC2GEmoz92S99xwv2I4jM0aF4MCXIFtQlRMmTcm
28MVJuOmRTFOKrCy//ickMWh9dSZBzvPRBzT73F2sL3BuY8aMkGpsoyvLl0Xj/8uGBpuAIHwyeWj
Tw9celaiPSjedrA7TWbpB+Cgh5l/S6dxVpuDSBe4qIsZJBJ3qt0wZwn8c6sgVZL18CdeSwtuK1Wl
mtoQ1cN0kGIXD3JwaQ1WMkbraOXD5ygbQRbPNH+oOyaJ+y5uve1DQmsJhFVHtdOcQG1vKZ+N6MzG
pDhQ25syMNww8R2fdvLoPcWqFEjWRO07LxGZvyByphVLOPlzI5mrKxv9b/jeJW27f69A5sbk1iZz
7xCjQQgKur7Ny6DWpM+VWUtFs5T1YE5mY43eyEYfAkashygPoGXMcxQ/uFH4ugv5PWTFgAc9+KYV
GRMzvnqc6A6Z5Ao27aff0aHlEecAtj5M4uy/+CvuVOq6Zxnj2377pAwfBP4mJIqO/M6pSbCnAJdi
rB+/CYGUfFzXgDtdQjGTuIP5cHeX92xPeChJSDSrkscUqnrM+becMvoaqF0Opca9DJA0FPt22Sa8
r5hn1qEtnfNrveUja1i6OB70DQRyYwM+vOaz1sycKR2MeTCMTJlsBv9DNo/eWmGB2EKwr0CG0Fzm
nRvPxVpRrSy7CEjLRx/gEqEuHsusdqwvjHWiozVkiCEXPMzOtoZr7fslESPtoFRObDFPA+CgprGJ
Lu8SEOAwHVqwAv8CmaXqBaga2FoDPL0UjoZb8gbxBoe8OoV05yMtD6t5aGnlEyMc89B7u2BfzhrN
/3fUPzRSt7j58I51NPSm3L5Au4EsD/N0y6TqFFjfUEKV4amkV3SoXtWD0IjCwAxgMqrsOH0o8dYu
P/5sT+UoNzQulN8RhPlBAE+A+Xf2M6sPVGp1DoJD+tz/ipI1pmJP6vKRh5yc7Q8QyeNYZWI8C/Qa
2kkj7KO9DfjGrig5DzxFvLDd6S0p7vg5p392X6sR8Felagwl97h6AFlsjqXqw+CLP7hZP41t+J1W
NivoH8aoWqFHRRwmsgU9w2OTuLr/h93F/fOGZVMDKvWU7fCKDSXQHewuuYZZKbSuy2iX7e21s0Xz
9FboxFvScOQNcNiUoCxQ3NiFIIRq0/4YJw/BmaeTO686EwrvO6TdUNlLugyV2VIj/9jHoWr9Hq6j
n5kqhXyS5NJ02lO8LCepjI28zjy9CAqdod8+WFcU4c7L2wWQmsiQ1vgN3qnDqOrggw5Bv+PKCr5k
e2bcjQqNFHM7/2CJnkE9yP3yt+vmM8DQWa79ZiyG8VCYoeHd+ymXoDFpc8vw9ivKEpcZtd4flzp8
FTs38TXYaHPb2zCW3DAq8ts205vAd+25RT7LsxU+ERV9SYOFlZw8Y2Q6aZ4xPDnE35Oo1XKhfq4L
qInQsMP1CqT344AH3cFO2tbMnpQKiPNmR5B5Z/8X2yM2ABxIOXsX3ILr5jNwp77queE8RKvvhZV+
+oUmSdDZ0jvne8fgSYroATmF1xpgsQpeG91UoDCmvcbVy99sQSqqO7KELoUY7lYQ2FyKX3IYAj5l
vk4W8WECxzul+deePV8jcDv6QqcxE+zo4ilUn37MUSuL0DXJ8QJloLtOaY++j7nuK8aIH0czAGRh
gEtHPAFlR8FMLKjVso1T5zuUuPsIWJMrZWDGfFzdstMRdveVeeP6OdAxr8SG/zFXEeifsL+oyGWP
rHfZgVkb3UyBG/5AIxcYi6AskohuZ89XJ9oxgxWDlIBWryScCGrEcz2lQuITTu9g786LI/fWh3C7
8ZJ9j/E5eU0vYB+fbOyfSTg3lnP4zz6G5YItHnififgQFn6vIwnvHL20kzYI9AR+dpdvMJQncPtG
v6h3MwpKMu6vsF3vZohAeyaHeHXH+nuC3FZm3CMpKTTy9GtThF3vntnzqynIb3Dmtz62ay2HaH7d
gMVVYsI8gQ8eklN0f2E96W4m9MWQI5tPQrSfJiSv9UN0zT9FlWDBkKsv+8bNSQTooAtpZZsNZtRk
iH/ZWGx/3MlJGWjUf3TazIzz+K9DuVFffs1t4izhX4TdPFw3UxQErV89CUZVtabW+60D4X3QS6sp
hAvORxD6/9O5UgcB9RGuRP0i39iUF9YfWjQ1PHKIXj4rOZubhMeb0qPV5PTjUdVO1B4/WJhcBjZ1
B58nWRW65agNSZ6U3PEnX1aOQPS/Lm9mEzO6LHLLi9K9DY0M7rcbYsw6bKaj/+plnPASud0mloNS
ofqoipZtPaIBwYmj0hODm3ZxqpbEUJ0d3+QJJ9Ul640v6XVf4ZqeN9bsh38ag19pAaJ6jSIW+k9M
g7vIUUv7C9uTfrNRAiqVkDBJoX7aCHrU56gZy+bxw8LZr6ZHeHk4IbyXBmH72myn7BZNYeM60SNt
+zJneAedUjak6pLpm4LqA954KzkzfT5fPBUYxGrT1gL/kA0IqBJQ3A+zNU50ciV7m0dR3DM/fKIR
rdvXOEKEWCs3vOKGZPT0aksfBkdOTeHzwXSSSwqjTISVcstS5tOoJNXEDrmFIDGoEtsqXdNh5fqh
MkL2mwtFTbe4Ivlr5DVSeFSrsMXdxHYT74mEey/5SQfsEUK8k64lml7bCHXUg3Z1ln2RWlIen6LB
SXF71BUK7VTCiebxEhGHIFBZgyx0O/uj1N0OIy2naOu8wdB5BEOlvnGV13PfntOZQG2X1exKQcYz
ZwhHbKGqjJxWxcg7BtvY864DatXlMReJRkYz8kYhBZLh8TxpXBzrP+qsjHPpqHj+H32nAxSJb3Ko
9oTyo2img4GKd2K7M6XPqZPiLCwTyUOq/rwP5UujitI+JWwV6QHg2Hr3tZsmpPev1LvNhOmn9Q2j
MMtAp2XdvEFV7k10IOyuOFFlMQKO8HAuYSFz/leu/e+Dp3k0cs1sVBOGLyOOk82Cc4cLMc6YBrpe
NhbvKeS1ymy4KRZt0YHrjKg7fZ0N3cE728l3Sj07jhYAWlbqKyNEol73cO9YDmyFf+e1L6NDxREf
XwtSRREDDvotX+RtGZ2q95gDRV99AA48/5GROz9ieZr/AVLtVcpu6Bou0CcueLsj7I2O2+ICrSZX
JEOnD1kQLqTHdy2wFCAtB1R3zkkuhTioYnQeNktFOF7d2EMtX3q4kF2gjbhBLL6MI7oS+37UkXI0
Bw6ZGx+D7Hq9k8vcGy2URku2kUiySeagGz5UIpnj1O2nQHxdZCDC/cBl+1bh1ehtu+PzZgtUA40e
YK0jtvDi95fDZW1INPwDz6QEDUUbfEqCJaGFnxl+HQE6WLH2Es7XZoW8l/a6YK6F8gNq+TIvY+p6
CNTHkhcqoop0ZS8kodEm3MXrRHkPtKXaNfEiqXsTEISnYHBtC6M4X1Fs3gWsdpPI5cFzdaxxEnAa
1A0vIbdctXJ38jC8JSNL3Xf4RgMpSkX9HzaMF5k4GJBz3Mt0j4+sjMci80szlHZHQhdFFxnqQAaW
Ppis2nHz6Xz4v+l4UfMrhJ0Hou9gw05ElTbu7XmK/fyBuhLtuzrgMHDClI1px4o51p5CQx/aF1PC
HhWcEErTyJ9/pLWnLvA2MdSQITsLT1NUvd+4aiiFag1IcwUKVEBT0UUh1KVijfKpcfXiLzT0bzGu
W8vfq7zxwdAGho/eWxOtC+itNeUYxpV3a4McwOUowg8yrL9//yTAIUaGKgbOEftUZ80ngI9A26aO
wsW9OhxMUW2dQcjXmQPV10ABYHU5wcpW6j+AXQxvDNXW8mYjjd3H+fPkYnwL9zp7w9rwP1Y1wnLk
OECq+s5sVLNo3p0Hnc+kBigtXANGLiA/WaNmzvXgyWvmhuLnvldekO2S37Wepf2ZzJm2qrxz+Q/t
UzOUiVhZ3TBcl7GdDoDmk81TP/s5ScyLKOScv1nugZPcg8W2rbcpJCR2PRA89n7qRUXNR/iFNQTc
QcGFMyzu0TKidJ43OH2clw98JXBzh2pfj5IKxbxynmINO/Rh2LVNGNt3lNY2gK6WDxmxHF0dz2wF
E++iIt1J6dsRwSVjTEXZd04POgatxopTyLlK8Xu8U17XGv23yHkrXk5d3Ck4rjA2I2XhhFofz6Mb
50ABMnwrqvumU7qrHLNvXvoh5fc5CqINE+E1Ol+NsoQXylFI/tmIxCtR4rlmBvrZKDQbNxXp2u6l
hXoRQN/4vRA8CcFutGHAXKWrDV2iojm3iMjvFAPs3JzH3WhMuqNEwV8YfE2MFPb1deveIt5Mfld1
JYTRQcxYXbOabsk8MjVP6zTpuUz44zbWSrt8TD5RVNbgL3+6FU1YfjxNpkJ3Wbai0qhK53ZVtNPp
OL2oOC24OTA/Mj0nK//bmxKVmFXOAB4GDYIBMWxg2JbLO4ZFET086PMUrZUkzkv2eFuipkzLYGBy
pO4Qqc7/mkkXX/S5DzURWD7F2GFCxVbfDXdBunSWzdYR59yQaiwuu/I63yNwmr3ebM8EJv+T9LrB
g9HcRdzCB/adpxZOBDGp7Fb2Uo6aRh1XB85uKskGWx71pEicz7FP2kvn8848ll86+22Acwlxl7Db
KUxUvMzNIYmnFPnND0F1r2SSMw8eHXkGLiyLgFTT2zXUfpOODeZekuHHIWlsunSQN8/sxHghrguc
dDyTcYr+Jbk/Z3AUewvv7MBhMVo4eyV7khqs3VZkAFiGxdhEv5oMM2E92GQN+sRxN6wEUhbM44vG
w6QTwRP86BNbb0JDD5KjF4ZJiKP2xcjFN9KaCDt1Lpd+m5Ik87ZRg8jOQxzFz6aJ852PXUXjXUYt
9/c2dWNXKBO27x/uhull0Hu/NLBT0ciGfffhGrFBQE11zwE3bhQN4u6/2VlIykOO+Jmwj5HfYI81
GCVrTunDHRSEsPqYo8fMojYQ1tbAy3MoVRqCL2KT/tNr5PkNmK73oMEOsD9mb5tqdidqxapcHa01
zKdtdjIzMXfNBB0x7VmsJ5KkobHUeRCBkqt3qSwLK4hIPBla8G6Gtvv8hvqoDA9x0JYgMZPmZLqp
8qKQ9oLF6/e32TZgcoToGBsga8yQP9j7kCJ3G73Qg7mZFQag4Eq4k5tzDfdVnBljOKoxkLUv6ijC
U3y1B06hAVHp7O4gkPGjb04T3imDXuT8d+Zy/t98moD+fkmmEYk5cupqP5L6u9SvbHmbfuQ1DQCt
6qh7hdNeO9qRZH4JqIbpdZdHh4wl/PXExTHlMxDyz8Cln42KyGYZoTMZrnqDpDAPxlxnDYN7QcJ5
bjA+Y7JvaWDZs3cwDjJYUhoNwZoxMwxUyzhwnLJ9UMaOvSyJz3hwRExAPOLD2Rsn0vJOpBe0wQ16
qQZ9nPO3YkNq0cc4NFhOfb7PFnX7vg4k6ptNlVFuebywh5YU3BIrL5nvQKjG0YykRRJbd48DLxs3
RERZe5FoFYq2L2uSOGzkVUCemAi3uI7PrQOLNk4TdO4/ORRhqpO+Q9uU1Wi47MHtFN+t2xmVr1DO
AyTA7sfPG3GAI0pcJnolQ4i2feNvkGPgOJU62zgofNywAPWPJjG7+S0JrhiSD/hhYE9/7Ob15O3O
byv3bCRizn5jXAYUbIsNA4t/XHjCPnKLSkca+vqnin4S3Z1q4oBrKgfmiyNXs/AXBKjqPswg55Wc
qOYIXURN9aI33YIiVNjZNiiyTXAZwYh+Yv4pG8OamMyky8MfFWWdzV4iGNZk0pyDWPHW+BWWh9RA
5LIZdAwK70Xm0aXmAhCckouPbzKH3aO0Y4vaiFuQkGAuVjWMVzyTPlmYf5NdJeENZ2oBESoZD4BT
vTtihG5YVz0Kqrb1tpQ2L6cfklZsMAfBeN8rl5viN3lrjmsQqs+242vLEJwJhWolgCOwABHqLQlJ
Cvk9m4/s0Kx//A5bzkjZ4/6fUzvlLuD0sHM2QSB216cFTKXJWV2sJeWrzfyRcUhYVTLwz9rkFOxs
IBIx1jkCHy2JjEIANeKfCNiMujgD1TJwVZDFLOEuZUrnwxNuBRALOltK8yx3QycO/H5Ql+DmcEZd
8BQJI/yk0ALUdqvpjlyVOUZGIo17Y4XDNsZErp6ul4RPJnQiYOnw4gUWpF/y8ERl6E5AvhsTjMyT
JUuBrNJjDQC4vi1OaORnDcmsJw8FdloLSWpqh/8M3HPNm/k/G8fcLG9edUzLy2OJTx4dc4WO7GxM
rLEttYU1JnTD1cbUQV8p0acFra7CX++ceZaS6xH8pjgn3NEvOsZg7CTBavDN/P65T6ubcdqnz9Af
Ow48XePX/Obw4Ayxu65Wi8m+PTTZMu0wZJTYS3/c8ewsOZq4hF4U2ygWDelqBsaI2/Wlb0ExKNr8
huiKKiPMgDWeTmUA/eHLYhJDL6SfOQD+NyRcxcoOL7zOfClhL95DuqYdIsqIvUgPZGKxeSz7aF86
20YMJisZ7+QQzQY+A3S/RBF1A3NmTRpV4nFm0zicG5VhiCRq3JQrRoWPyaZePUorJmReRcP8t1KX
Nqv24Jm1t5eS1isoX5HxyuKRW+wq54v2Y713ZNZU+hermi0p/+kcgVTmaFcrHP9vUshVloZG7yiK
hxW9slaGyYoHHXPKpPHDIxdjwyPfHSv+jCc5Lbf3Xn7fg8FFzzqwgYIOsARtpIVOZ85szVh54/tA
7+kVyQwCZHChQvI3qxeZIuYOo4qeaM6vmjS4NtepFNUuDFpUUtCLB+BNox6YhLdX5/M95J1pNlA0
AGJhT+1L1ytFcqrj42jUy8UnkPGWoCwvjBkm2eEyHC9PVsPewAd89FdJ9Qt+n467723yxFpAc/KF
YIeNE4FTSFyz7jew+CedIDUrhJdb4AQ36Q2+aTqdkfS+pL6Vkg4+zc+5/nuvagzh7S/rKYYf5T8t
b9AkLXjSON0xSwZxPyVqAISb8D+JR7VqKSxxaKfpgwT9SBiTrYmIr1BI5CXBndE4CsNhisIEAmE9
TJ9iCq7CZKczCfRCvMhSkIJZcCh29mbIsNjMgXctWK8nh9cR4onbbzQWvE4HijoctZ83rRTBTlJZ
j+Nz7KOtYXjSNvoRR/pKPquz5ZyUufbjxSZlWZCRly65lXBUaeb04a0cvzp1OrT/zb7cMFTCZXL1
fX5Trel6n9ZeiYY8hqD0pUucb0W2sD1HJ6oUDgD1yeawRnfk5mmss7WN7MMvIvq/qblXFEkAflcY
9Sm1M0HEGYQtCbffOiLCvT176uTYxVCe0b+Jyr7xWlsnGF1oOCorgvrrPRaQIbkysz0GAv6qek4l
IVzvHgZmL1sHSXSO6O3Y0/oVH+y5FCDScGVLswM7rcrAtLnw8g0TF7rUhEc7pl2VXARC95JKNcQE
4NPJlp3JsDXlJpFbGNpDeMNZEpyD8K+GAiMX33M9nNcp/6b5NL8b31AXE5jnJzOq6k5KQlvBV8Ir
jPvrWRzmO94V4uGItN9Sb6VyBYKUryNMjH1XGspetPJiy6AwOLHvF8R4ilr8cczEhEITUxqGc3Pe
7xNaya56iJ2JQUVtOmk8qhwAevruvRcXSDvSQ8wKreRDuxu2zb2Df9Vb4lFgL8w+NKX1XIlqSlvf
dA3TRqK+s/weGUrHxB1J3kOxlQApNz65chuUXJwnfjCyN4xugGvsnk2nclf5juNl3/+cjzPM4qmd
VgpoFBtorE4oZJ4hfYg7OdObgMRlZtOSdwLE//jx2ebqyD2FTUTRfCrLa5MEpi4IXtZfQkFeoihe
YcxVh2nsxLAC7l7cP7M/OSu0gHYRKYSxjanuj8WgtAuGyPJYLUrg6TNyWJux1nduffSMFEr27nzW
M4lGp08XPJW/d8lg0uKLs7DfTBvy1dm9RRhYqEYs4/EDuCPDWfZ/gIWRZgLpLH1J5OvQB7DXWjEs
P6oKgOLEjbS+plbBEcyPH9GODsVOXbwWF/azzyw34fCcQzyvVKG98IUkGwHk/EGb42PdlgtM+YQ6
edDqgb8OOgsVKOiGZlug0UGLKIzvIXdZ4cu6aHb+T3Rk8Iv0MIlTcyST6l8UuW964ekgvBk9fruA
7ZlAVvQOD8B1sPTYamLQ9Zxm3k+V1yYWBFlN7k/F6EfZq0Vjl5+Uxsfghdct525/nGKTQvcCLI0y
oTRGZyRsqVJnMmhj4egKeYiCn8UQpiW5gbQ92BoeMNQGOPgfnc4Lz0rFox3nM3cIgG526Uu/moAE
SLxgxoeSOw9mlp6GZrsZlWmIha3G7ESctBXp2gmHNlWEJj6u8mKtxZH+s4fqqtEhSqeVtOq6nvKS
9Fwdk4Szz1MQ5iIhs+gTK1n2we7/J0lNhEt0tcaDxoFD95gqCNisc0nvg8zbsNkVYWZgxz4h2eZN
L6h8/XTHfdSg3KfeXN4EC7N+bWSvQVF7hU2iV7qQD6iXDYIIkEyfpcCVHCc8av612ibPtsufRiL+
KEb+7tzdgV6QAaKz1et+xsyx4srRGvTxeDwkokNLFZpMfJLiuam2lFQ1E7kpivmm4qimdTxumwug
6/QfDAsmRNKVurBDlOcVGZcJx2adLzfkCHIf/KcX0HR9O75KocaIArBx8J25s5BB3FP+RqZ6F80F
JVjJeV+O44pothvBaM/86JgGHqBeJL3E/C4lOm6DMB2xYQREvj4lzRK2inWTfjudDM6cwxFNccI0
oPGt9s0TlN910zo/BN7qKAMjeL/5F7rZNl7NrGCA+5o3+an6wYW1ZulBiqlNUkTuBk5Pvz41SxqW
zLMhjEhaXuccGxQHJVWq10cWkdaWuebkpunbiG9Z/cBY89tLgmQeSRFfzhvnAs42bxwlyb25SA26
1dj/MHjVcex6c1BAfZJAuY8hI94GszY/P47vohgTxZ0kDYgWzo9PaN6gVuP4Ywt3KMm9xIi5r44V
petY8SXzBmmBI4en8JzAK/GwfuJBcTCRp2xZM59IMYkNEyK4IquzfnPQmsYCPO8tMxXGmj9Digfa
ZgoxTsgxM7sbeMSwlvYKvwSMxcO8SA/m2WrtHFSQyohZESywMusBhmSbsPa2SV8TZXLGSuc51Njh
QyAF0Ki5vCh3yduFV6+To/H7UJLMqaxOvG9/GtR1JAj7AwuXYBF5Q/FRNiUO0C7kYw+JjE7JlsUC
brQjyYW97jaWP7Nte69LCeABsSR0Qw+eRaqm1c6bmXs1OqYctH430tBuI35D5SpOS8FJTyAtzD+/
0E3yhtZk2DjI8NYS3hRcjitLBtdcba8E3oi681L7wzASXA8s4yPU3rKALRDf9MiZNoNo9eK5HCp4
pBQcbTO2rdbeuTJjlKV/cu+tUVppfa7WbH///H0+qS6k3TmHE7DqP1W5U0jomvwBgaz1Bz043WOS
Cq8kibDBkA45RemwfEn2MqbyZ/usX11eyiTdPG1xKDxO/G/dz8Zwxr8cEqhXXgEKSUgLK5pZ4BDC
ohtANfh35xhh9losh6PwsjaAubkDF/3fzUlOzfAFTNss5pHLOChNXHeJ86WtmyRte6uOQRXsDA6w
sx/sLaSjOm6St9Yfu3vtoVyxGlKbAimONC+1roBovxZr15vRL3dAn5ff+hCQoFEI0hOUUf+Hd8UF
yWW/6pGmg5JN/fxMR7SS/gKQD/WNfhvYArqrw1td0WKzTVGWb6ZgdjdJuKXq/+/NlsGLcdcGDgq3
PwKGLBAHEhZvlyn9RHW4IldfdEz4h9WLm47l4InEpGxcp6m6wZQXTQX14uxawNQ41nTiyrcX6KUC
4FxfXOZyK6RrDf8Mflt1I1PjUWwhh6U1AWNEJS2XFTsCAWabFpb6oDEmbZBAE2EjbUjugqluMmy0
df1BFnIkkZx8w313eOvaUM2fega6zKi04GDTBMlDJ9VuYW5P8xPE/ysSwOaV9xy/E7Gc6Fq7SFAO
PGmQV8fn90FfhQ1wDv5AaKkdoLYMgowS9FaffkmAOZnee4ne+d/xEkVfcPEvupb7NxwDfJmf/QUl
JIvMpIkm3oIkFH0OHr9KcWL1xHopt/sMBG7aqIi1MNivlDFWJd6Te2gO17fD2AMLlqc1cBPGpLvM
2cmBzJ7G8Y7AS8Ho+XkLVVtEZfUsGBpYJFiLIMGfnnGhKfQ4A8gomIByeBHwYEZxLovs4qAr6zan
Di+7pctsJDqtZyZkByROcE9VvWl0xzl1587tPOUOHP9mImjh792QzsBFKsBhZCTdnJy0x38mL7pw
3GDMu3g2Q2K7l4oide1WtNwiGGaerN/O6tuJeZH8FciXPWjNJXgFqZ1unrugGrqk1SaXz0KngIbP
I2ZmoHoqjqUL9TBYgLIgQg0m6LSZa0hcbdcuyx5qfAr7fBX5dMnvY6cnGhFmHSiSZKAght1X3FOv
0KbjMztlh7iFf0c1JwkisMpo7LGl92W71wsqWo/9779f/rL0C22XlQA3ZdNBJLgDDCmMA23nQPpW
gJbDH3h0oA8NZY9SXHTnBHMamGRrMwgNcrrtS7MpwhqXlSUzJ0PqWKRVKuP4e07xk34uLhf/6rY5
8gfCfm6IsMH+uUtg+FfUCn5MO+Zf/gbmdYI97v8ZuQqpoX3AVSw8GvbKqE7sadEjHx7BsiJXNo0m
Alpl29J5DCuscFeonO5ExwmO/YxDxXhD91We2SVj1Fni4PiKNYxpiOkHq997mJ1Xg7eEUY3G6gSA
jn3705scgRSEfwiKMVeOMdq4BdSb8MYPOiqQcyWDjI8i06Ay83D/lSOfL68qIEtlC2s0MAZvt1K3
rNQc0s0mfFZirZmCt+YkrJ9T7T43BCjxewQB7IMX60GJyQGmUu5JP8byT4C5WnKjvPPrPysadTY9
1awhHe557K8AkwJX9gcM7iLbaiYw19mqKHP2hJTb8MEJPDQZOb3Jvo5UzYh28CO4Ago7obIAHBay
nrZogmod3qay7ygis04vsuoCteTRPdXa7V5CLTPGBkz2nb4opSuCvgtt1nY98ICGWfaOhqV57jVb
/3xO7ik+r9znOE1tQPEy9R2FS44CKeQx0gse062RJ3cVSpnMpU5II/CBWAqO5G4i4Klu6YrLpuSS
XkfkGqq6tgUHJNApB9h8MrDnEmN6VLeO8xY3a3MXMSnqtNVl6esaDEgHGFGOgjQRysImVLaLYhIi
c2JgxsEIReK+Es83QGDufHrHsJecIzKU5p5uAXOj0+Qjp3hv+tnNAoXVJ0M6cBrgTRZl7ztP5JnG
vqY4NIDRIMxTfomTVmrLRrzOyT2MGK6ZVOrIdCFso45wRDT3QYg2Prm0Ek4R5yr/TVD3zdX4Ulxf
l5DeofKMLtxhNUZIjnUWhkWCwhWEpFK1MPjmGsUiyzT6feL7EPuzUwZOgdDQDIafEyi2bSPfdgcK
Qb1P+UVALNxvR39dUGXIT4QHI8PE0ze3FzFEfgs2qqbw5LwbpeYh2vW7uvFI9XBYcfpkZCvVX5P8
G2GLpBAPXN4Dv8N9y4/EAnXeRq0juDnYvNzZ8euhXEXUhb2DRNbZauE44+9AoNvoZTTHfrSVX4XC
ZHvkPkbkQrTZ70Xn24NiiYffnhWJCfyUOPnKDgu809Ifr+7nWYg0MjOAe1HqehluFk4+AsMw+1P7
ZO2AkkmxWOnLkfGPhH4pN28YpeMf9f8+W7FTt2UvPc/JxcSH8VAuIfbWy8vExj1TFAJzDVKq7XDE
To9ZcHp+5xFx3bweW1ahtBfwF+gUztuXoripKzpR33OIHgh7oBs3oA3Y8LKdTuNLzKjjTsw8C6Z0
lE3Qy5LVYqTPwPDTyZWiB6+mZeVG15CujqFlQQMNYhzPC1KVQnlejkIJ06u+fZdSs2+GLeEqGR+l
UYX8JFzXPth2thSG+SfYblJvMVR9u4XOfzygs3PZHzKkJCxnTDhO3oSnViNMfsC8QGInqqyJZBdu
p7OGahmXB/9n2U7eeQzQjktOH4eQ5VkfPanRRB+4LCQASZ82CdzTpoBD/YnzyNS8yH3MnIbA1NLU
LLG59W+qT9YZFfi6d2D5Ed6eoh/HEg5PM5PcB63EnZzg7jOIpmGoTCtw9v6c+u1sTElyoCFwzuSz
KJktPT62KzDk/J5Dgey/GpTWLdwGVUk4I1SmoYujVcm4QQTvxdDhiD2715p+viMl45FUkG335W/H
zfUxkq250KD1A511HSxKA1kawd+nPPMBYN0FSp0qvE5bN2vU5gVLpt5hzPSxPORx1t3GaDb1Gq0o
3ZLWMpxbHaOo5TrJJj5jwcC7zQRhYWDg4a/lV1VczQydeUY6tp7mBxXh0AKAMm2VOpCxoq/7TD4b
yo661oeiNj7/j28JZ+BC/0SsrG64QPjadnxrbtYyD9H8vOLTJYNM9rpNTnNdN2DIILI5r5MBJy9s
TVSAnQe+m/BLBtrBiNDqinEa2be783OCCp9DVAKImXgaL+ddj98Nq2ViD22Xxd08Qyh9cNdML6Zo
A8B7JvJLAnmk/3SHIzEqbQxbMi6h4F0nPCOlAblv1GFxPbf/EKYmNFIcwi93ud8s6JOuxOfCBSyt
W+w2K+Ro5maaLH06CgPkgxQ7FY1RaJYo1Y39NCn1Zl2XPmUWjd9yFPLQWLsc+q5cxCtaMhVaQYa3
ET/b0eT20g/F3ocHUyKxFZlxpoys8maXToaTJWfOBz2YugK6tm+SF7B9RTkEJctp3ezFUnYI6Ic7
MiM6fXjim9rMHedQzA4FHrml59pcRZg21c01+EJFjiF0sjM8M6q48frsnLg3RFw6fwWZ2QXJ0mlP
B/bJ1LpKyEP3CSl352O5a6Hkpg/MfsTpBM9kJ4Tm/4WjpFLto3vpRqXC8o6H+LyKVGrFwUDnvwg4
tpf6RHuD7zl5Pnt8ig7D/6qMzCIkNp3KXUmydibpZa+o3PEaucJtprgN0x0C1Nlpw48CdV2Gnay+
Ebh9FjcfzsXnDwL6zVElnfD51i0c7836P1rzSo6iN5NumelgLKpGh1g1arFBrFZNuTKuH+zP9BOJ
sMVDzbSAtxU8Ss/Oazoi+Ilkpi2p3VteZJ18XcY+Z5m4I0OjVD6ZGoN8/WLg11T2vwr2+uNypBBs
BLv5ha9cGtf5s3Mc/Nag59j1KNUZTbvsxIGjFuQ5g2e7d2Qw5rARBcf01IwD4Vi005bSW3lwDWKT
3fKYPMI0WFcrLKHnxcfi0VrnL3c+yVRJRXbZHBXBozdEP8KyHnqSYQjHxMb63ovowS17nTAoMY8G
PN3HpT6+bEFCkSTrVXdvRvbD0tbnjxxtAbGxL2y81oWs6U0ZsBAwc+oe4C4Kl+0uaSktyCK3GTuL
AUbmooy7fUPCA2LVcGMCzYAxrjgFNZqzzsj1oWSRc6u3YRMmr3Nmb89J3Kr4ZyTAo4lxGxctdhCa
kQFTnzQaAggkK/4mTYTQNQfs6SQWRrJiqQtwtDqT4m8lPwBWdAR7D7fZlIO62NOqDvvj1FzvLe3n
Oz2C6vNnbb1LF/zOsT+P+CYFtvkXC6CP87CDlq2BCz0RPkSVsXYLvBt0gL+QPyE3VtMgoKwzdFgL
u6bcL0rGi9xibGqk3DUvLi1RrDHZABikfHsPotAHh3JJTG72klVb1g+8gTy2oYwco0zD9OXEJNTO
Ai43Fy86h91BMIdD3nyFJe8SIIiyZ/w75scN0si+mc4JxCpXW1QUGGaaIqnVR18IXKacYYl+BZ0d
5vsBu6Db5XRVbybsc/HAvo/yBMmcjWPMOYkjGSolv23TYr+ILiyvuULwDflFf/1/Z43TAK0OdlAI
CUhIOC95etcs5ntJjgj1eWzkTFC4H7RO2eKn7tgottYWFf29N7ehq4eGkvxgUKWGHu16KbLvmIAV
huuxV1cKE/pY+ebE9Rm5Nmq3VOWdIngf2ldk6QHwKtu09B7xtXGTSkKspvvRiS+fcxS/NF06ymAG
3v14eXkUSfJRB8p9lImJvrnC/BceFO+3q8wKn4aAmodceqCGSBS1iIIx8wbtzkBeG7YyoL7Y7FMm
Le1jO5IVMh/vkoz/rAsowdILNoHjckqhiiuhf6ua8Dcv7Gbvd7z0gYWMhiVMUVmeoDS8tSl/dJNa
mZJ7OJVJP1U0dVEcqTyVUypwI5dohLrl2yOLz6JI5E2kc68gvTqX23PJDoYKGVkegn44DgrSuCd0
NAi0HaV1CSE0izu+cVqGzbREtCEwdPS9DoM83ThLpgC9X97WmA0QeJS1YeLS+HgfE72w2gHrep1b
h9sfZcnHh+2mXLIm2sk4CLYc+HWAOnDpJYj51YfxA1AWM1lc0kTPuZVwHORun+K8UVGUGYugePA9
CkLk3vuHUfPug12aT7/8GZ1m7uzbcBtFtomDJLp11EHv0leFdOFE7qwNQ+BvJD5tzsSL3XE38E40
apdHcGMa1PKQwaRawI29eGljwZqJmlbTt1i9sGdZ/dFZUFDbjtVnNbZKm3L8ntmwA7sOQzJAe1c2
wg6wpPvYogSSbUOqZvZi9IbHfEJGFrIerw5FU/t5ZX9S232n7EFpPMbfQwZBmurXChIKzsBtQGHK
CKmkYiwuAPE60Ey6RK8dK7BTHU05LsoWzLfeqodhRvDeDCOB/6NQv1hu5Q9vI3wc+StARsbRRf9h
T3GBQ1jEnrQPbxSxKTN7rzExHB1bB/Px7VMf7FklxiCctpuazCTNZienpJD2/sws06Qd50vstulN
rub+cAFZyeJG1Ovr/pDqDH6cWjDCLcs/IWn1Gd01VoKAWR99kJJ6KEa34+M3eboiKQvVwIaBeEbo
6XdrfKbF3lxaymFBFiCWHG72fzMOvC0fZ7RtVAhlUdOvy1ixf7ozHGAQb0QOB0hFj11S1skf5/tW
rYoMHYsD0F1iiEnS5j4JJ0r+3E3h0XxnTBVtHfRSAz31v7BahFRP58xTLtkQy3Cq/LNKKYqNNaY5
dNqmMXq5O08cYQLs0+fYM2Iy6Ky5Yho4m7qzXrEsbh+2NFS6zxtn3Ix8pnS0bUjlmM7NT0tlBFke
hZSkIuoA7Gp7r7mbibsx4m94OnWZpQIMPHpjVteNluwqw9bciGZejtiF5co+M2T06g81fop4vXJZ
WM3tcXIv5JR+G8GwcQz7x4rmeqovMH1Bnm1rUSAk3KogMgt3swODfYNwwl9ZdPDsAhN5PxjaAHGq
iIXcIYmEqp81w4PJYgGllFOJN739K7hfasNf+mvNlbJDVTKqe13qC5mcocYZOkKA5ggduZzPhjHM
Tey/IdxHV8VMg+niCZepOurQ09n+KNchWSXzxm3xm9p27S4EM0YQ5UVAu0JakbItVqEfXCxbW6K4
VPDHgEjzUoFHUIVEzEfwd3+qgQr3S0tVtDuRp18VwORH2lDi5D3sXPfp0hodz9NYqdrj5XzA2Lqe
nmqhqpeiUGhpVq1e06+En6+Kk6CR9NdRGEJZMS2aog5mat3z5yO5zqQjKzsOLrk+1kzV6zDTGzGG
zkeXOPq7zpfh9CIipH8HA0guKZji3bDlPwYfdR6KOkUWysutf4zpMjjb4IFvwX/w8uVuFYieyODq
kgUX08flPHKUXmjVQcxG3P5+++yk27qt6+Mpf6SpW4TK0RKHNaGpJDqT2nUWzrT7Oh7OAZtyc6fz
y+oGec0JOIqcOz36kUjuBg8jYOiX6C2f5KS00VL7FcKVYuqxdomvyBNHX1XkdGwK5XSmabYP9DEF
sShnSfF0TBFBEcegBW3hadcWDQ7hk4v3Jof2OVkvlKWVCJ0rJIm/EbJU3bxL3xR15htzFd88LTFE
U8j513dEwzAYSVLvHV6e2wJdgiDR3R+KeYZSVknnpDwGnmPXteIIqKDHS6F6EV4R+i7fzDD9Rm89
FzVFcCUI1XBWhdHQ7xT45y4BskezEgQVvWp+XYzBVlH+pulMcev4JLkIN1G+rbYFugEU57QwWp3p
9Qjn/EQyAnaCSydZpcCz59wEbAUYIE8n08z7bFg7KZm32Vv1Dn6wfcPMtrvksMDwUXmP7pApkj6k
T5FnqJh3K6G8RCqytRz0pYsRUMwFDfDXGhZ9TSDTBsfvwTWwGXKbZgOsknoo72seRHy/zOH5lwWT
eI6GIPzg/f8sAvkqAODLa3WEYqsHgyg6zNWCqXUD0a+k4OOBXh7ILHMrsZVmluGTBBkcifW445gJ
E7Q0OJajE2pkgLrPQcbEZVys28FT1Anc1Nu5jfTvn5OympFwKED/dDtxb+Uwa11d4QGn5MpNm2sY
aM1wtP4W54bOjJXT+Z8XVmaW5mY+EDOrt/6LTWXFhZqhpLUpg6C2e1DxvsBVr8ll8A/HVK1QeXzc
xRqkqV2eyMeLTm7SkQki9K0h4D48aMdAtdBiRhtCUGgNgD/lA/8viiqyf94bEA9E0FrntvBlvJd0
H/TnwRvX2kGvVRPNi8aCpmJtDaw/708OZ1FAaq0W1fxm0H3zJFNg6r+N4mHZ3izW10+qAoHem5rv
G9a5wqw1wBkOmOtouvsehFjIYhNsNRg5V8Gr3oFhXsu+fYEDaxFg8HcKjtKXMoZYL+u60lNI9O+K
rR/8buff95jJL2HiiCDdnLBtCk5Uw3ha/LDaUL0sfSj7Zlr1JZOAHxkj0aaQpiUXrD1jNaC0UKYG
q1G5LFd6dg4lwNl4TBJF+SttGh8Q35cQ8HHhLdM/cWn0ER1YucbAn8qG0ju2VBg0ZoOC6Ph7QvQ+
Ux1l70oMi+ZB5ybEqIAOptZ0lW8ID4QV+xDb8HtcSJj12dlytJCt0pDs+IvE+wOu+J8isNriU6bp
Cp9yS/phHVNs5Vl0kvh+YROQjV9yLJ2t5Cd+E+XzJVgSqbOJ4wPqG9vtdAEbJzVSDnbOp9QzaDet
6Bpl4ro3iQRkbFDNGZUgp6xNrNmj9zcwASHWBNqQ/0s+KQiXf8LtyitZUwlpu877+16A17dIEZYH
uxP46b522e5NxW06M0H4s8xv58gfXBKjGKOgXhRPy0wJdsjK1p7PgO7ed9b6ElgbqdBuNIxEQfDy
qeSP2wDnI3SUq+bVjs/QppgNvtK27Qs2f3LobJHpwLqsZzTbKMk3dCkv9f6eKnfghLUkB/IsZfsK
DxUUeHdGyGKU9qybyUDAPKWXYzyxgRvXYSW4QcfY5sYCLsUMu4Y+DviHFtgu9XA7qzPC3m8MvkqQ
DodRj+jW7qp1dXtqmRcBDeqvQur/ozXG/lrq5GTurseFdA6EZCjZoQZhIMp7MHQn6wfbAW/FuFT3
Y80EQn8g2gy4sA0jMF3bcq0qTXd2kLDxnVQ0FyM8dPV+G5X9UTkDM3oA4K6v6+i8FhEBBTeMQ+FV
7/tEVRqHZ7puQyznBgeKnARGRdrbQWyk/CBYBK649A2oQ0k8p5ols1ll3FMv/DOEWH5f7F2yrRwe
vXZahqkl+wIPL0HYOeGF0ZbmkFT886hc8q4EW32HIUmdYd32T6AzbYMURNBcRg5+RUcs99w+t9OF
XwVDpuPxkXBueuOqyr4b44nV77cT3OCBcJgaBdZ7tYCScZ8EcX2DFXUHGZqVm5UM56B4b2w7iwfJ
f573Xq93VnGWcPtc8pLNQP9q2i3VujZ5KxHvmz7p0T/4La85hiDVoQQJa+u/7yfx1tPyDVHW4WsQ
VQRyGB8JDexyQpvcSu8xW12UNdK2J0X64OUPd+UC/XlI10dKajYTEdiROTLXWAMswy81i8NoOga4
JqdU+fxNcV83EVoH1Z7TKp7Vx++N/IpjLnK3V6CW2a/S63ETMQ9oOSrcGAy3qDWDYXoCCD8y22Xl
PRnAAVeDPntXFB7stRMJ02jW2o+MMy0Q8ZQ5wlNQm3M/yPEfpXEghto+hROhL6geFQkdxEUHh+5m
GJButL5wuiDjq4kFBQOrm9MnkBxKeEU+CfeeMt6+1/AHr2tncAazXDlx8oU0ZDiE3e46B1yiVLNp
27QmQZCfWxAsMyKyiBWetasvQiZfUzyXktGqseYusfROBmr6PfiH5O9MhlUekpfr04hb/YJSHjGn
f+rUPi2LbUHXPSJbdv9qSS48kzp17m/cpKtYk39dB1a8k1kioWaMqwQ+l0n4I1MUpISQL9Vrfnrt
VuCUpipC65Jh7qWU5ppmCOYgJzY++oU+1Ol7yFKmEhJG8cnyEKyMQMlbjCRBelFq7ldfYMmUHZuX
HTT2EKQVWLcTnZVjXvBNDzin6dOHDBb0luD9JB0oru5JJE9C57efeBYwoHBs7KoqmXGC/jsfi0+L
zfB2hrSZRNtCnc8VS7R0of5g/1WONrgqPU3xMVo/0F+Ag2MtjoQDc1+dqOS29KwzNLQTMh+wVATG
uSFV408teayO2aXJqDN1mTuVqwOpaD7zu/4yW0krZz862RKRQ/Z0zZ4YgKnmIia6mKppPu4TQ+H/
YpL+U8BT6IA0UnicLzF4bOxGOFT7JklNunDBt3Xe6W2zeBGEButuDoKS5RdqBpDCovkiTbaAHNvD
+DoM3rnddIswEAuDOJV4TksJDmhbiykXDU3ZVlEXaQ53ZJpd4EynGjO9Nv83i4cu3QQfilVr47+a
qz7HmSLx2tkpMVglLr+HhMCIK/vR3KU1nuUozZRnhcA5qcjNlzTMBknlPGS0L0egoyZRXZd4WWzi
OF5tX22iLWFLYKBKrVcxia70iCbPr4JTpufj334kuMKggRv/fj6tVNVh0cjgyrwYFu5Jlu6oiUPP
WGPMe7N6qcdbRBwjt4z9LnSn9mFXHlmfbMGVSmSVr1+RVGBRWW5CIYSloRsZTxTmdkF7XwyeCEps
DgdCXPEgfVndZKPaG6KAzCTPzjUwZKXrjJpEdOZdoeR4A+EeImPwwOVtZ8IeGW9qYQz+GuHE7lyk
t1WwWIHtDbZ/mONVnksBp8OOpwlCd98euNJCJjxHiboxMXnTRPY9Lpgvfr3Usi3nVa9TxIto1mzx
q8DSx7in7P5bK4dDP4norLVmqF9/mwrIYePGWyg92z3MOf9pcTF1SVl1uV/KcpORmckeDqGVzA3M
7RbAFRa6OGFwpCJpNqTdnnbifRA5eQl263Bz82Na6ljJ783P7Uf9uasJrhSSVwDYG6N2+rjaDDG+
l8oS0t80jCLEkIeci8LJv7hWgqD3cR6TRT46OjmOOwarI97AtzwEgSdABhjzSVgRzqo86At/Yqmn
j+tMG4DvEWFsRNl/15YZ8WwVypbn+DpBMxxxPlCxy8FDAfjfv996HNqLRUdg+uyWCHuL9QPqr4/O
jJQY1mylJmWDcvpGQX1+3CnkYj6YTqXqgV0BdLNsWADVEjRxVEq/VmfBqvLo8OoLdNhuWIJX2mLb
tbpNkoXQNVb4Fv+Q6+cd3iVpoGm4lo4RdzMIKrp26Jm5jXQB4lQoDjR0PXaJCtwpn/F/wJ19rqxK
Jf4Dh668ZrrIwWehHtj5WxJ0tiWCxDBm7YpZaWQlm8f0VNLI6sCri/SRirKtvgkGNITQF9BXT5sJ
upvSP0Aouf1o0Bw8/qEEhM/Ca9Ndk1aLCWp69Scpsi3dIAwbGLEtKWT+Qq67x1aes5e3xxtDbFZ9
o4oaQ330RgmmranBjKbscDolwjeB6Rbw7ygmyJRrtiVXRM3PxHF2Acn81I35XzpKUEfe9gk3ZZW5
XE9nMlsqAwhN3BvOlmEFg1sqI9A+ggqT9pUrOwROnedBAVYL43Sa+OeTWbw62a59hZ7o5T2F/AP1
zjDECT18QbYMZE/1gtTpsz0Nfgy6/fnVwbbFukz124/WljZoJVvxz9a4kEh3nnNbazYlGJzCb3H6
wE0zX3RArgDEKqdPseKuiMMkYJcFL/sHYhL8eib4ck1hh2s7ip1Mj1y0/evWQMWlEgGtl24zY5Tz
52wpG0Wc57IQ0nyI346Mk6tgd8wVuaQYxbfC1zg400NOZXI/7EsVC6J01LVY04m1XbW6p/cVz/93
OHiI2H1MfwL7PuHb/H+wZmaXgbdPeYgEXZsBuYRyAxa14X8BWcMC2aJb5fFAFu28hWgcb3bt8dU6
iRsg7ytfh2qCUvxrbK9OC6AK4aYZNEkchvvDjl6NMN3D9lryyPm/q5Lg8oYMjJBky7Oj9ppiz3xU
SB7TmXE5KsVVQbhB/jGplQhyW5EemnmVWVnMWk3e3NE800m9JLyGLi+iH0U4knp9RUg1OfzJnsws
F1yri+G3RIMMe01sByMGu05xpeoPv4S5FyjfyuHkwMd90giD7hZcA0bi7YM7featR2mbYa/99zXK
vGs4kHnfgPstLBFp+C3J8vSls7zPC9H3oDZ7FBLiYuTM1mpLX0Kzu/ryIibMjJ+i7vQFojd3+ho2
jVwnRZMUdOnhZkbkOCzjp7veGeI5O1ae3tSjKo17G82JwVcdtjjFf3oTyVzov7Tl1u5VMpGT/lSg
NUFqxCBUDVBQYgouzzC9HJ6gBojk0u67eGqDfkTHZbKtTEW5WPWRp+kT8uZggToorUMIrWK+y4JS
VfDQxnH8hb+eF9APkon3AugF33gV45lxeyZkZFCl0SuHJgv2DSQwf1sVDoQq7/Y568Ih4/nD5N1c
mZdmexbF5K1JUuXthI4lAjDrL6bEWAJaowfnG910CNdBgbyMiIn9uSYb8pgyeEbFvVTeH0RhUT8u
ih5MJzuE39wPTWJRsifbV5P/YiQtj0oDQ0UaODODks6Gzqj3uvcNQur7u3Tj7EZ47mIXy5qkIo6e
c7B6KlkvNOVSUGOaQtYM0XH4rkGgNyJQTjHO5LrtXOVYkOi48swI0HOy5IT1wCHPjePL5Wvr4AmK
gfzDx3fJqC52DrVYSt0tVjqojS29gHYIdgplAXNR9MmvVvlHB+tLtT2uF5J2RbqU7w8EYLTLew2b
vKAKW/hQtnmSnNoZVqacRa4a5jlbnOMDChFdZ3agCD6jRVIQxOg5ITM7izPQkd9s/K8Qcxg50hBa
wZP72XqkwS6R+HjSd7gmmuXQo4QMnSO/mEKACoBOZhz52MCJsd3aTCwKbY3zPeFAHKLlONhbosN4
0ksLAvgmOYIM94Kc4skFhKktzOP3McT4IEjbxuDkGgpIhG6OqUzFE10ki4T89+Y30qn6LPdlDXp9
v3UcYiGlev+auZvccw3xjaPxLdrIYcD6y1dx1h2zv9oUTiJLvBDZse015wmWo6lMgU5mMUgVLhvs
Fa+quBPfSHFrrc+5t0UYVKMYa4T8SQF8NuJYSwhJhZNa/HiKTGW70eDN5DOwFVjU43wq4UCFlmHq
zwOdPXASRnUFRR44Qszuq8UTNDjQM8gbaOKUwVhOfnhWKo+vq+gp9iQRj8/tdavnbgvmuTUSnH5n
lUkkPFWY775DB2ypFh7zZ/DJo7TqtGKOXVrm91oWYNvtYc1sps7xiqf8xuMtSQkTqMX2m9emA9SQ
kHG0qz8OVcoxtxqsYed+eS+i+80sRYeyem7welqRKHPyeDKc3LrxKAEXIAQ2irIGAOrR+JQBC9oX
sdvs5LJBgOJDkV2IoL/Vd4eDLQUHsMztwGo4L0rEzvlUpCaPYpcfi5wNcwe9HXC3/wYGDVXo5Zd1
eeXOUU+hlQQryUAVl1XKF6qOOnmnNJW81htDGAnWeBX3uCZbVa1/rPu/hfjq6gakcO6X0IPF8Ppj
M8KtAmVvzuZ4lHwgHei55BPMwWhXDHpHUkzfGYX+PI+mMwZbap0wSBT7S2+bsCQOzXRyJCiSNTbU
JMhPiM+9l/2BXox1LDfxutioAVMQ6MIgcQWe6d9M+cInTJybhYpQWfvcEXPyVW6KkkffnbH3c/dl
45opOcQzCtUysTD1yBFGJydBq2VMFua+yyrZcZFJX6rbzc4QMLKu51K84yx9sVXVHMYKaD57Y/Bv
Jb0PKNXOEI/T9nP4vLHyAHDGUARNe54zh9UIEZFBhFSoMwjcvF20knsyW7EMvKp9KsSTJAPVBPeP
wKvVX6BZ2wxUYap4iJBiRU3R4qKdFVDCNcX0HA+cFuVYlpd+6CwbUESJ9QlfzU5h/CC+9v1QV6bl
jFyHXEoAF46mL25oHp6PaxLl/xJFNoOlFav/G7V8DppZ+OPetshpZDMVYpUL0URDu5aU4nKcyjEz
aqz5bMBZI472e/Q7ysCXoMmhl7UYDF5CwinKeOlINU8etQhSClSae5aIfWesIQqAbUWhxKlz1jBS
hFlqdx0LDRvO5V2x0YFcvcW6uCn5caBsv8HHFcNs6971YnW24+huJ3TUblGKjBTkUuANbJcjYGFw
pEPelUFb4e7J/t8ISzAgU9l6ZJDYNdiWk3hb9gKuOMfcEoKaUOnak9yr2SxQrs9b6qXupTZQF/HS
5dNqXjBEegQYH7jLHYZ/EbmlNy3Cgc34i3f9sldLAN9/4Y1G8bHZRwW0VY4M/aIMLNqa2r4PkmLN
kFsVSvUIiCycs0KShrEYF+ZJHKoKayukjfPDUjIwh9872YvtYI9XjPAqIuS3D4LnNbVmT1+dFZv4
lbRUGQoOcMJbGXNQYwpBh9zZkAUMzNI8lg1A03q9Lb4G3uPiqyezzJQHEdDojlmDRJ8s4TiR8RMm
u8kC1zDBOz9NlYY4+GBmlHo74TOh8B/d5NaUzRRyLwsrv4Tsu2SEtnjv25GOKa8FuuIcauc6c/Gf
GPcNTsgse5iQ3FvnD9RJAFfD+CZaoQ1/WK0sfUGdUmAtejrSEZO1QEROi5Jt+tsWfXERCd/AYg9S
Oja95fwjQuvSbV91NOamaawRxfJ2qjNlaJdplAJDY+mLVV9sOCE5GYmCgYq+Ije/5N79CpH0KbqI
PcOONVrBCMeKnjp+zxdLTaRP7Jzwj3wdgrA1iFw0AcNi3yiTv3V5ezywiliHKKaQorUT5PBRuKh2
KI4q3E0pxkuvRWugF+BX9YAnkuTTgafgd2mSkp3tYiHkO9S56AgD+3rWF9grhQwnFGTu9+xpW+zi
Z2dd0n3i4tpBH0bqiXiGIVuCDjy2Q9ETEn2P1HCLC2vwJ2HgBqTAl+IJSSpgek7gRrldFP/NbyeX
2ppEipEGxQNHSQTKFy9TybZaHoJzQggYLcCLi69XYaXNwWcb3GdDh6RVleP0lJOwV8uEJUL/IWh/
grzRmHDaLm3P/SckHs/aB/wHIRhribB+o00oZj9QgRDHKto5OKJGCzJCBdcO68oOAV+YlNq1h7kZ
qjX5tLpFK6jgMung/AShDsd/cCaIaVrIZCZN17B1TmYzS20/Mpg3IPfujsxXe8r9XAONXsH3u+Hi
aZrkYvF4jCRZ7OgPZYEKnWahVMJOeNw7USsgkq5rNhpAbkMWk57Ai8SxbL1V2tLbiNyTquNFQ2eF
69Pd3qAgyuArZpdkirwQiXVhWQhzkB4Tvp1Y03f3PJsb0I1DHerzJZYLMfDE2oGxRdHpILJ8Tr8h
4mOKW55xG25H62J//RbO7IYAMPUn+UJgbtvZOiaMPGZ8NC6caDc6d54fnr/jL/Cs4hH0bhR2EVjE
sxYVSNffokyMAXXvH8RvKZXM59EWWrUhhDSr21DivM3yPp1hcU5dUWRqQ4QedOLIqyxp540EsWq1
jpgqPOk2uVxeSrKq8DG6xfDtnIsqu4sZzFTjQ4yeM+y2dd33js3KUSUX2hDIwZrZaUjJcDXfbRiY
PaDoA03Cgjy/cxQffDsV3naBm3eGT1AOSbI7wx1y/QGlB46cncgKFngv7k++daN9BYI0r1cp09al
6b8SkdUJXBBCk9Inm4bESkQBPxoWeBPlCL2qxBB6hsmzlujMj4V3faGl6u148YaJGusQeGjblaaE
64hrEuQPiaf/jqHtkakf+y9oeetwedIE4DRpSUev+6FIzC+wXhcsIzd+4zDwuPbtvVIfpJlcFlhz
3VE0gu5KSJiPl+sdnA+5oVw4VvRL9glC2y+8Tc3dS2DpH85migYJ+eYruKXgclt/VZdlw8mG+oFF
uPSn3M+y3pOB1CIr/W/sXv65OZMuyuJoTYgCXSVwoWjSNEXGD16H+NwVs+IBe3ipBxu+qBhwABv9
pffp1Cw+T+86Va+b7fJejCPJT/dO0sLH/2pg9L8LHPZA7w1Ms8rf0NgYrHzkVFJiWc1pcBCMEiF3
yLJTCeiYP4qHFzNPyVCkC1sRwar8x2Nr803ep55Ogygfb+AuOaDlflfUhIjLf7Q7LLjhjY3wibsR
jFsgy1Ye7/jqvcpMXbH7xp2owohUYuRls0IJG0tyFc5NtnLi3pVxu9cn+K28G6v0gi3ci2vHpbiA
AB3bhati+rABHbCaXkWOlJJMKfgbVGQ5I07SjcJqmkaCUQJ/x6vas2nZ6QszmJowk7vKJVUyFTkn
3SrVoxilaxEDMimoQ+n4B3VgX6lnB4nH/tupmVFlQhQpzpcb8XzPROIGFMImk3pK2M3NNBoRSRKw
of1X73WroRC9EG5VflliO4iOQbmGjT+XK06M/fmbPFudu0vQT6UmLThcEklH2e+OVankBxjYzzG/
k2DvCPkdoJA1FCKAQyunEDLmUDhituc8QZ9EbJ0jOiMG8JqWvLp3cYJFC9R4SeEi8PLqfcso6yeG
4bONs3vBrVvua76Gao+PmksVAOiLnCymg9vkuce8yC1Pfj1j/OuA8YCwFbZ3JqdoRNJA13Ag8Eqq
PGB+rvsvIhZKDbjjbS5SMtdw1OiHiOkQXNnIVH/XQoW9rVUs0Amsp6HNiAwYkhDMuT37yGr6e7Gl
KT3iql1rktRela8DT4nx9TnHl14D5jAXHuGyzifv9lcVAPKkyLxGi+XBgoJGcgmb/oDiTdqqqUqT
3K/ZfB1sbDaPgqWhkcBk4QTEAa7d+tJwulU5Qf8vML1pmWosuB/i0iaE8f1P9XtARPAviGnwdjaG
20fry3m9TbaJjpxnJKeMcYECXrwe6W4f9k6RNOnzNUlWg1FK5qt9cO4uEp7mWY1WbU+tig3/U+Kg
ErgVKcmelISXRwSNaZBE0/QcQraMaazgQ/7h8ewkbG9HurYSmTCtwwTWd287Uaf5vmFoEraJ3E5q
kPND6rd8rvP6+bYcqQdxKoGxLxetg3WblVjNh61GLJyyd4ZeuSnKVW0sPWseIryg1VAlGtM7SPNO
tqBhwEu/0vl8BZTeHe4+4tMn8XiL4nKoP0nFVTBbarc7Bf3hbX+NzfD6dZAtjkuww1kw4O9ABkrq
aF2m1oF5oOhHCPXXaviWxw/V0o3m+mnEH36GIHv3TvarpDT7TiltP4XxiQsvz3zL0/+4YfF7eZql
zd1BCRQQ8BKhW9jTumD5ZQXvXfjxWcdZaTGL+bJHZoeRI335TTJXxcQIb/y8OrZAfvXxJjk0O7Gu
0U/FzBFum7mMdvutSrRzpHVc3Ixfw+Dg4xgbYVZe3Qcx5SigYL+f6iyni5fbWFxDfVPZDMmes0T4
P8KNX6CkZCJfHKoLDVPRp/8d520qkkpqBwZ6X/PP89m7PdNSo0ZK6JvVEKjPRcZAsLKa3VcBGl9A
ZR11e8zgP+3+WWXMAGVx8KcDbcvENY2twh0PGQn/PC+fS7x1OFzEaff9cSrFS4iF6KZglL72peu5
uMDBMnmMuxERAFJCyy6/+C3ZnhYaIhB8+8Yea3M9FNFqzMGNBCYbwSTeVYovaVotsKqkof8jAqK3
UxLJSZo9bOFvDx2SaILcxQSCWyyoB6BJLfDxPVahGZKHhQqOT/kv0a5l7JgyaNrtktTfjnFx343N
jHZ3hbzSiw3b7sc7g54KWTHlyH09E433+v+mRYYSIB4Od5GUbQEW9JZOeUJeRu5gpWowciuY34pN
DzaxAO/z0cabdzevvCIesCwZLI8kUZxCZrtu1e3EuGGEVnWX4amxYetADpnHikoA6AFuCEJXyaqW
joF0dDsdac55pk4zX0MTD9BB/ULeMeR2oNX2bo+PcweJhHLUkNtLxinzk9ZjA25Sg266hX8Pwypd
QtHjinYwQpAEs6n7G6r02ZhDh48ku9tdns+IScSf9d5EMZosY8pGIBkv8zj3s34pzsz3nAzsqqH4
4a5356h5Rn/SB8k7oktFxbxT7Npv2tETh1gxQ7WPvDdU3+Wy5Nl8vQQCmu1dWPrLDyPSdN5Sof86
vPI/T+d+KNAWNIvli4Fyxln53bTiMSk77PairBhvIENToy4jn7hfJIeTkmUh39zPpuf//2udDjQ2
Y3Z97290MS6lBWbY0VXpBWEzCAzLAFD6cDzgcSOwwZur1vMgwEXUmzgc01c/AC0Xrytj+aJ9nWL/
Vg3HEfN3CXvOSPlVCToHmRI6wL98XTdK7H9MSNzzEBAzWTdkgQbWuRCt6JrztZXQJ2FqPjO6oRr/
tNxhRQ2vuuIq0UHgEXRU/Lb2FQNze/22pOrX+bSXG+xIfhPdWHI9Xmsg1G2/zDCn5tILZ73t3OB8
kBRXx/90AcVmwODexOpLobWiBMFth7z4iJHJEH2avis4+Kb7xc46+Bir13X893wtqcPNC7APFUDO
tUxweUBTicPbTi0rz6CgPiYfinsdsFK3SSkTtRcmFWpmlQjKkSuiWuGCP5PDvYrvF46uNKobGZ1b
g9WUhGn9hvwoH7ny9sf8DSNRpi9BcaBdlPJS2evKfhHf90kj0G3puP6k1qEbI84lyKzitOyWdSVT
ieCKXitxB7jywYXTsRtCQIULDuSOwSBo4EijMraoh9Ak7Rg+ZuO51fIsoazDNljO6RSQex3GL8RU
oYGxiizYmNKXFP7gzRAtl39gMMqcZiNws0gPFc63gh8ZVKgpRYfnTn4YbS8OP8ffzqXKtX97A+Sy
ywypWwRNjCO7F2uiaNsGevE8bE73YCie6150mtC1dcan0EJd2vrXHFtqKFndG45zNc+kxxKwI3Lq
rvha+gH2YXKzqcOszqaYy5HGbwfpFmeW/VjVp34Zd+OUu+PoFlCPeW+ZWije7Gd1JufCyLMANbX2
NtP2jmwN/nA8DWZDs/xYvWP9C7LnPOSo3sufxKhf0VAH4i+LyGmIgkOOGBUpmERACS3BVm6icaEW
8n3DmswegY4qhhojSvGpif0gMbH7iOlbNXwSsT2QoX7m4pam7UwZsJHqmgAZxRSfy90duFCf3HQD
PBPUMv+krLEMcK0LcVlHqPBsBZP2IpfRJG0i5OPsmwXbtEPRviyHYpXRcHpkbtN9eJvEEAa74IVS
i2q9aWJie7RdMUZOAhyeYPhLPuzrJrWssjBXbJYtrOjX7N6WMDPqLpVcC0Cpz6k428Ciu9/rc0tC
88TJGcRe96yGHCp7vqMP/Hkj/WOnwWNaptMAInUBv459+DS9xD5xX6+Vw4BGMnBdLvrb+j+atMIK
eBTloaI9Z2hbgVCOUFgRnz3bhmYo/fvCu9P7bWPPjMb/d7mbKYHeLl1B4eVyXvHBqRLgogce60iQ
kJynCfTWc4gF2MRCjFfuiS6nY6XcadPdOI4GzQo60JYFqjIxmHZDpe8OI33iJMhAueWWGfgWS2f3
3BDdrZnBWXkf7h21avuuvih9zQc2sk96L9HZnMrPcKcw5sPEDta/MPzDCNdgN2xdY7VhmWtNnMkQ
Lo+SV1ugNNYmvAMYPiuBP+DrdFo4rGpsU05gYIwFNzoLaFG0aMBIqbogYd5HY7gNu4zCU7yw+Z5/
uKFhmiTzHkRsmw73ZfoCfX33Inv9gKraeLfqvfV6oMjvxDL0T0VQbLYQWSdlkxBPtOfo0NS8EnF5
vsyRmBKLOp0z/o2WPpJJiDW/2kYvq1JIpDweQxJMOLb4mvicwhGRTs7MVb6KEcyuYi9wwNKrqzxZ
7mf/YF8EcGtlwMQpziULofNbK487Eb79E8GZ/cnwsMxHs6Xv7S2nI3v0BYNMwOvTjA8LPUWPFMg0
jp6I1vdB0OGTpX23WWBsBPqQHur/GbxU1BuAqFgKIrwfF16BCtbRfBgqvEE8QXAOH3rtPKF5NT4q
L5w/B/DKSMwlwZVmvCVVaRf5jewFDVZAr/5o8oLbJoZUvmRFHMs/T4fWEO93YTnsgC53LWQOWq38
IjthKF7c53aXyK6tWosREmOFCYXrfFwtkqnH4zVpRQKeKPpj0PL8ssbk5IeAcw73OcRiHiR0pl69
wyroP6qxs1Un5+/CWRTQLedXx/zdlPx/LNe5M6k7g2Ksck+E/+Eamoa3g9H4yfOGfXDuVhJALA6k
8FJ7vEDtK/WNfx5rjFONxJAzNHXoFfGegKpGg/N9VzzGd5Nyg5OR+8cMDtT4JwHewthDiP0Zl3zc
0JUcbvm0/fcQ5ARcA8FpZnDTsbggKuYGHrr2P1G7kljbwruLtb4Cv5HcfJBCwywaZtY3OhVpAp45
1E+PauJfUCMhS9kE4PNRA99iA5OKMPTHvcLH5DukITpHnzKSBITQIyIp1n4zEAX6DTBQ57sUo1LH
+s9hGxHsuXb2N3PqXIWVi2+AuOqg2Qdmyn3tnvZTQrfajSWMRulGmHkHjLma809Hl39Qsf9k3PL1
Cxv6AdltEB3YOyJR1S2qx/KF5C2+q5Xh48jNJ4ASRIiggwBIdCqe7dqL1HaDoyHMTyPhH7EtiS4+
5vX5Wlk8CwK73ZYzVvfGi/zZezBkks3VbsRudyzDOIxTMgJoQNt0tGbOzcwDmsqw8m6qLcnDLaUD
a8ZZTSDNLhbA95iyyn0JjlYTVJ9qQislZr0IgAlh1oxVAjIVydJdRc+MiU4Dw8lWNnub91ky16pD
vRBt49Df1VDxwaQ4WNKPcAOtJl8ssJ28iiIyCgrylpVVVQYkD9CazO+fcIppyPwCXud6Fj2D1Zxo
KpUOJxCBr7S7Vb2P9iQ5139J6BJP6GaB8KhFG9Q93LoYo8T8wOYiZeAI4BkVIlDEzaSuBvlJxGBp
/HvuPtOhx/WMETV9VO8BfYzd9JiLBdl57GnyaYQ4KH/KV1/cf3piLLoGLYifI9rnlmKVzHI9bKo0
qI7EegL/9evfTGwjUggJoxtmxTTcx14JJyqVfr1CVJaEq3EMnsIwdn2pwpcV8A9MYlr8Ijut2uSI
ZD0kmLCzsx/v7Kte3+dW4pH0FE02B+WiWYJ+DKnLf3W4LgXYqpjTgVTfzcUkwXUO09NpNlOCmOwi
wA45rnihCvFHt0NKlxsc4A/EKXNh+PttG3VzKBffd1nb09aWDnueN0s+o8P2trIs4L5kU619acDv
u5h/GFfKc4ve5Who4VV9yeDXoT8+8hfiVX7R9CV7mvL3QmmhoviP0KFgQ/vp8b3exxHTRI91DzEo
WWULag5TWoe+6ZbhiwMD3y4Oywu2QEh/xXZiwe5Un/jBF/wnz8B2w3O2V6y1kyMjJs2nZEdHQ5yf
XqryyT1sbLtjouQ5h/2YPnQcNABnjRPR/wDNBcPakIzcRUsR/rj4yewUxjjfJZvhkBDNqz/UcFsC
9jW0OJCWL3Fs8wlRpV2/6sTMdiHitaBxK84gEqRrlUjt4Rb23GF7HG40WRbfL36CZy8ca3rEy/GB
8uu3E6eeRWR6loubYp30tuV+CjR0vJ9zyhIJbSaEj2+tH9h1k2MRGOMh3o8yk41t5VzZ9TLrFKwr
GIPCa0IMRRZlsfI94aVJAk2wz3bOsjyxv4Kis8pNEgRR4KAhv55YbQzNT0t3Ip9vVLBMQSndA81n
8dLO5uif0mhCtEfHqVLxPr76uVSb6DTAb0P/ZJElWCC9Q1e765jW8QF4SPidCC179FRGEeLqFt/2
A6RIIkdXDQ4MpsjkdpjjsswhblcnpztVlEDRf/U8KBMQyMrTC4c1l34fwEbpXbixxvjroWwP0g8A
xxALSHEcNIvKTmwOtbEdgb91PRt79Blx156yLEFDXMZ1bvigX4i023e+IPwJfzvtm+It1TYDbuRh
iY6KH4HfSV8G1PbK4yxFjEgl+Sfb7zdHALAB5HbgvkZkpkgXrK4xsJHibH/rg6222GTuS3Kyxrjm
px5yDOmmq9DhJJgxpzPOEi2GNGa411M/jNhBIyDl0HBRtIrxfSj0oWpxe1xXbTyfr0fGkcfjaDLE
DCI+wFVHcZUUC7ZeKsqrXFcVt0RqqR7x7QsAPABc1rVKAS9LhdSect6SmE6J+81HmZ8sZDZTyf+z
oGDXLG9ViSFjwvYdVzUkjzYfwA6MI2Se/SkBIsGxxO0Ln7yqdXs6uehdMX/At6HtAjdbmi8NKVFU
PX1ZBc/J9bPa+ZqsWYrL3Kt50T0ceFRMcDQKIBwl6dqkT4sTYmTxMQc71sKMaitASFbe+fbxNej/
M1xKm2/h93k+XmSQ7bwArq/7QX+5MSpcKewI4O2OJc5st4EJTLmS6tt9OEujborO2+P77wWNbodB
FO7c9/hNItXZil11n7d9c/DirldQTDylcDeuqLnrm8Mnc6o0mNWaCJfUdUhThEp0MpHHCXuu4p9j
qBiHVNsquOUE93BogIfp97jpSmqppdQCA28vfys3PYgdQ3Tt6r9OI+o0PejJTL3uWzSj8GORoklb
fEG1kvr1eZkZsGec8Az6fg33jZww5oEP2MpkAbLjQAwXP/+W3FnbLnlgEaJUCEYZowAhggDTIm8R
Q+ct3fMpKmrHgwPuouEjDP+XgRxio3pHSdnr/849pQdwiszwSzru8r+gZ4Rayanlvgh0MrwVZg5j
FUzN6m5kzmZwXosFxXkfhhJSWUjKdq2KOOEfgHGsQqz9VR4li1da4ShheY//d+S3Gr8jzm44OWAq
aFlVCkutt8BMroiYQS9HHD/o0ayJaRjDoIt0JHp4Duz2DbVabE/H0ZzoQawYiEzUyyYgukiKsZ1r
MkC4YDlAJVKW3oXmaJQ2bj8arOv1txTBs6eUBc9miOcY+j4D8Ayjvl1qS53lyxL+rNLQr/UPOOS5
e1DU85afrreDsiuOcnLOuK7e1YNS7H9e6lvJFzPF4DRfyMy/NuEyKqQ2Ua3k2aNf+gflu/90wMPC
7wDNZ/KTjg8SbCTjkdD3M7GKpL4DgLis7tPdSSsQQCRv3I8e31bQQBixKJRzNI2K7A/WlPRJm2fm
NOUysh+aboTv3K1gmuCiOKOrRShxglLdDztZsorZO005zrz8CiyS0ZcJP8i74pwhU95/luyxsK/a
pRPIooxfOENJhmRBKmKuF6avG3doxbfwJrrUtH5flZEdTdeMixigRB46ec2nnnMa4WwlaFFZq/am
wO8S7TnQNnbTciA+7GOf7GmsbM4etMICvIszPu5BnDHHwiZ/2JGwVqEon/Pww9hvawn+WpSIl6E0
YNyeQd3D5Hl9uZVrDvfdgfME3EYq6iQwQQ+8b5JAXD4iUAdlkSzw0OPLA3uq6P+jupsLQV/Fw0ru
h34VMTDDp+M4ljWGKfxQkt3tuKrAJrBNHAgZPEiTo4slXn9tsd3bNgQzI6opx+//6SbDMmXkqYMp
ZEJ7NXYTy222s4M8caJeabrQJqWwvW7sMwXaTtQLg0ItnRI4QxEl3S4WL9JC5SgKyaLxS7HLDtv5
m+BpONmJgl8cifMmfL6TSp3N0TyRVT+GzC/b9Z1MpAZMl84PvKsqyJ9UaEwAnSr/ubTk01Rh4hy1
wyezDUASYB3u041j+n5j8VHEQaFk6zshyAioH+eHOfmHQLi7mrrQoJ8W1mgIekUexwX7gwfWshLY
3WjT9icnpdybWnXSHGDR0hCxWzsoHwxCS+lMo96cwNKzhjg+kNFPw9vDcbY32pzZMJhMdbdFzZcV
hhxhw56scr8qO7TWcVe6MISFPbpptdo4vFet25nGhjJRX1ptth6IAsnr7AiGUD5rqed+aKleW733
BkHu/y9SlpIWqRam/Gc4HnnXc4MgbkdZhwI+DoBgdCayI6aBsi570oxrdRiS4bkGiTC1IKaBQnlZ
VmQNDN7M1j7CUpJFBxNHQdbqwMuMh7j+LY4Z29fL4lf2uytf9x9N5lHTPZT8FooHCtpcdxG0qNn5
rLenIDWRgvCKni2l/mcXItGJ0hYIsgsyuUoYLhzTMYtHOkIPCq6PF57fvcDBbWarAcCx0ZMTXTIf
0HG3rCWz7NcVsuhgjJtcacQUTNidqU2ganWmqKyXMAgHCgMz2MhiqHprnkD0oPG7jGDCOCvjbldE
9mjEQQ9VEIQ3/Ogcdmg6bmcPX8SMMFKrk1irVHzI3Oy7crhMaQss9+LftIJAvy7gUpyDdh6mHg1w
b0UNTu3MEKE8pLSWJBgAL3mJmLNXNyHUAe+QD4p7iKUtno3JPic8KJFQ4AaKJtXo+TqiTgyLef74
kfJbGfupLV2tdgqqTjcrhwhG8O863GgsehQBy1hqdrigQud24AtN4OFE0F17/RC/ByEN2YicXyQF
zfOdTtR2Hd2HOlRkjSTuXUZzXmrOoHVLNVmbbSqxsOO61LyL/xcRY/I212znVf8EAw9ZbvG1w/n1
mNvNL2M3q0x7Ag47tvipk3T5yFlCiZ+KcPoI9rv2nn+0uIPmOxCCNmhSUwD5Wgf86OdyhgVmGJGA
iioNb3Rv+NtSAI7XveJPh4L+SxPxfPyiIzSUrdnz2eYxvnYeCwfqtLEsz3SPz0NmJmTulRpgcVy4
G32UzmdlSRxtbgZ7zvUiTCnk1ame5TCANBiDod3Xigo71e+xCY1ftNrIQdXly+uWvl7NNkneFnjD
g12sq9XnK8g+ak82c2+gktsVcJ72n1CgcbZsGsRO6z9vX35JWYEXtppcfR+fivjZAlrYxZMJY8OJ
uodgj2vnWaZVp1Yjo+vDI1eEdFxNDmouKmsUFJTWBazvZxqDG0sip71P3AhehktjRlVFIphCPwJU
Bt+Jqr9z4edsDlw4YSaa+tbIh67G443LAtmKRR0vTaIBl85+aQFgQBkGUf7jLwnlU3nzhLhB6Cff
zWMtMeOARsfF6KghBWa40B9lJANn6K4yclV6b0CRJ2iskmUPYyvXOjOem/64vrTlp6OgCBc6Q3L6
zlwGlKN7yFWO3m6GJPJHGTPlJIhmNuWXoIT7JoylkcqvCTYpPF6njAdczsbUga/4cYIHO5H6yyrJ
+Uf5BB8BPiXSehsOlzPr+sNuTcfIL3Qwf+agl4ATupLkZo1wj9s+MgIBkExp17BoeqUIQL3bQTp/
JMge4umMBDGU/9QQ17cQxgtT9ubkwkwHYKXHSe3A1sLDqwWHKLwm8TVDLudA6nDFJBRIk3BBLLxf
0P13NqQwlLFGTolBMcz2RESxY3txqVSOvElNT7m7RvrKJe9Pf//TO/W1kAMQjJw8ikPMMaTfSufD
9TXOuOjEUnSOrXetE1oe5RL63r0nBXbdEIYUlu+xKJPNn50RNdBoLPAyZICiiOF2d069aJmaLnI8
Xj1BKhp7/qoUCkVUYx7vpyvrhpniWdDGfKrvm6fcIKH5b7i0AegDRdkYhjOwlrn5CyAvu7sCNnBH
mlXBBhbErB9eg59Ne3LtDhG7lwyHAfBJ+rBaFcte37cW29DaJZaBGDZLybLONKfxYTqsPlBWHKLj
nN28XP+pYyZh8fy27m+iabSTCwpXpy9U0jC0etuPaV6KYN38+mNvqs6VsOAOya7KjartQVmfV7II
2oAPu6lD6wBP4lwtAMn5MxMUiWInfTsoE/oheDJTyxRRWhGIWv15+l5CUv/Fld6YaZs1p+l2WdF4
ZNrXX8BehM1fEALPkIVAKasQFK65rWPtaDIVdDEcpoz6qQLm+UVyu/D7dwKFogMV+tYIff7853Eh
nLl4CTNx3Mm6fANRLI2l+jUMfD1eg//zvz6CLB4+8xAVFXjT01VH8odsSOtGo1c/bnq+F0OfGzir
82Br+41I07MTzjifAQReY5MhPqPAwbYCG4UCM24UQAQkFwT2ohnNWamqtDensQui8djUFUrradH4
oREaMZCgNicHpY9aEiAej5Oy7Ws+rT3BpxWCM4EqA2wYIQdEY71bPGm8NnpKCDTK0EqjYgWUORMB
7vCrUhzxzVMPVBSbcxS67R/tYhWQ1hAZHKNHdax92nR8i9yp2lP5RJozXLJfHO16uPRyXDNA39Ob
T5UBBrXNUGA6VJ4u56bF0ynu5XWxaGvl/satdQKqJ9pkuwAOSTp1K77cn4Fa3kHLVAZUkWdskrhU
jQyYlfSHkizlfk+2vbvRMjBk2vM/gYSVOFjtq0jd/z0YMu7iDHAHw1gBL798KPhy35fs3xcsFhoP
WpwO9BPxUJMqRAPfpN3LBsNZQSETBioZzcn6zU4u1iuO6JSJcGd/wBEO88FIl6HoAnucJCAgFJvD
g3ff/eTPIdQbpr/IOO5AiJnLSZwWeZNSed3WbTBJOe6S5l21V9jWKNaZN/4wRdViEVdjmUDz2OUb
qwc3kxfhxRPCSLxpUzm59YYVP+bZ8S6rR8hokhqq9ZsKW2OaHvlYC4BfGhJZW+h5WYPT+RR0/tig
2KxRElekQ3ZnH801To+Z0xVn9AUbOFsVVKq+byCsyo/t2YygWfxOIBaHCH3IaDbxuyfsSlDxk/EH
nVEEeWVDYaU1u7ZP0LWGOnjqujkFUV+Rl7nWKtgk2mJDCbsk0Ow8bGq61Y//wURpYBsEjzNucNTZ
KbGoqXN1Q88pwvJRex+AXL2lkzl9dnqxt36Ji9nY5HuJSEiJP5rRcx7SFgTdLiMm+qV37bYHYoxr
HG5BSTYjQQsC5yiekLGQKE7aR0axuqZgUJ7tVRFepZppRlIUec8jHiWXe4q1GJ+0vZBekbD6RQvn
YFw+LMbOJwfqEJtbbB8xDK60siG1rpZpWUyUQOTzSzzeCkaDyjo/dsNm5XEbRxFjCi/GOEq+XKLN
Ioj0jN1E8O+8P57pcknFETTvb/h/FfPxZojKc5mcoYQrjuu6DQriC+Erffi+8vn5AqrmSLnZFV8c
pb/jXnbZlF9dVmhKNlTfmXGZKfnW4oqCHIdngqGbuVy4AnjRTkX/ixQ8BjckvxfzWdUcOpBc/qjN
ow+sOtIujyX9EvUnohwTwgEOtUj04sqy0Ynkx0KPMffeQF9BFXZMlDHpCmMPagDP3f7gvK3lafwB
0uiUCJ1q7ImidkM3lZfbfHiRaCyblhwr0lTvbaaq1hpc+G50Dycsmyrw4hIt6pHcO8qTCPkiD+oM
+ZXs9yxLe7HJDk62oDw9kKcasI74VmzSbrP/EUQQOMmhlD19C/VnPKuIkpAhTsdg4b2j4951Ebbh
cudI5+1fybVsXrE/9YSOtQONm2lilc42KhguBxvUDivgfz+ERfpbCq9h0ldwTCdGcnxoY2qFoEMZ
ap2xR/OPuxNa2u0dZb7jwol1JQthA4eOsIyeKDz2yh/ZhI3ckB1f0Hf6IoJUDuHnftfILG2aaIUi
KXSsSFqvQhJaRohuDLELWewx42gq2ETodssrivBDWyOmcaeEbXrZHqzYzERtZDQ0zeXV8+xotscx
ZPQ58xSHtHWcR0uVHBcmz+rU5FsFsJVxvt0N5ifYvBdYhqBt3y2oTruHd+8D+0PL0c7QfGSekxho
IQTNRHW9zherUU/SSBr2wArHlQ4oxZGdsG1hikG8u8fX+EbLPy8b5eIkrX/1Tqz6vL+9AHxWDQTI
GPMGG7S86XBBbOpC7U1zIDkYCqt2ug1yJ9gJNTJCikJ4NZPuZq4fmK0mIvKo3/X6O3t19XNLuXHF
259ENOS3WI6gzXbLZc6UQ67ZfHMgKT0ulxups+NIfp2WvCbrok6eQ7SIr2jIZ4nRAsjZvduVgibI
B3hgcujCe3+yc1XFNJUi8WKbqeE6JH9AeS2n3cP7rs2VwjbmPNQOlCRgBmpvUO6a/vgHVWu+vXPY
aCZ/FY0uzdZH+uiesZGwdVKSZW3V4iOg3WQcGR1bWDdR3FQmi6jxJmJ5mIhT70jABpL1Nw9R021q
mwUCsDKcLcRweYdU+VeglTk5hOsfmKg8JYim2dOcKkFQ60IXXenJr/+oCGccuWIHvwdZ+2fCTpNB
i5Cr/e/jjs8Oq2/NzRI1FZTzg/c7uFvm5RLYYG5aJWyX/j4fOOPnrknBNYQ5pc29lYKdc85ocJS/
PZRWOXeDl5kpDDs/2nBAL2m83LOSk1XCgR4v3zh67ZGMph30ZxGSchWTaw3+7yc03KUPSGCH/Aqi
GaUv5Kmm/chjKg/gogNVktiPF/I4wZHsrqFXeBr31IrvZ/DN0pVWn9kICxvd7Pq2Q73JQ6qpFu6O
kf8TWdt84JHK0N1CC6AhfkHAO994IViueAFKLjEVPLEONcd+VsIQ1F1m8LZRKgWztVI6QHPjdTPo
nVx+qUqzLKj31Qmv5mIJdUHUvXEZW1cznYT3VIW0ShW97T4Dar/xcrqbb83MrS0CdSKQyCNMjEFm
sN3LM8lph1j9CNcgmCmawa+FQZ0CExS1Yd4WvpVu2VmD6/fsYLBR2+5aEQeHKs8ZIZ20AZm2kWrR
xDY801cc3llZg1n6Baj/la5ss55i2BiryawT9lzYGwK826iyR3HNV0RbnhSWynCQvtpYTnvyhmjk
/c755Tj8yKJEtjoknAhwD19faneEfX5LLSXyo8ElzOcg2JfIwlb5sBE6mt9+PZRqMADRQsNDvpj7
bQHNmDKjAFCDOX/hfQ/JqxjJXrhsP1dT5cfZbjSMxzH5m4SJNkcQqHUnXxMIZhh57/DuC/NedFEf
CeTSPt8JFzccclCy1R6tE/bTedidOQq3OlqsyLe1+aa30JEpn4SJKUnzRVmjN+Cq22tiB9HkkI9X
DnXmE7Eq6lXfupbneO4ClX+fZYiy17Jg9M8mwJNHVrBVC0fJ2bGrBLpouD2UffCF1T/P37aMHY+J
uL7F2Cw9DcHM0RoT4w3LEZCvrOIZp0ER7T9EQgogIfjIXj5lmSon9cXiXjsK9qVmkEv3UVtvLEKP
BibQltAw+HKvLDfRPfvTgWDJXX3Dp02EQiPBjXiai2VKkfrfa7glXfKoy5ZV//nyfur/b7tKqXl+
Jkk+7cZLlqoKVl6weNvOFYSrSVXOvYQtTCKk6BzfS1+xrEGyyr5mCauFLc/PYKkRQIngVEVZppQ2
+An679sR2ti7s3fy3fd9AROzKpWM+5nFp6gMJgy9RUY+wCpI7GyHOwkNlo5ULcZYLvAbqpZbAPFo
MNGxO0yLT6cOgOi98FXtJsG6vT/jVYqSaHTUEr6snbO5u2h1qv6OESEwUn80U0hp4SDIRHqOgUp1
phADTdnDmNY7ExUZl+Cels9vICuQfuUNZq+150KhM+VbN+7hKSDa8giJjf2ptup1RATOB3L/uSYK
Do8GjGK0s16X9ATgHzf9V9ihU7A2qvJaqdbbPM+OJC8AcTgCyYClDihIBfgvPL97BQIq3O6dHxI3
fyHoH70E+J4Yfq9dF6cZp4fiRhG1wMa5yBTXDAeZu6W4DuCHKf4u1YFiSP78sAvwKQYtp+kfP/Hb
+9vjNqCu072assxNNyAmZnytcf+bU5Pm3yjMproSspO0Ax7yC/11pCZZ5U/lEj+C+TrZTpidOnSf
6Rzf1x0iRNybM9y6hfRObOPedACVfxgAb1UTNd+tNjoExjo8CDUTrefnjJ/e4UD/xMyZCLP66dez
MVESQsxzttnAmf+fVP8Gv4O7S5Je+RwScvjUIe7gtZ+OLwPTmmWDtaU8MHWvXHNR2ruSZgPgNgbp
UFr9h0uxcChn1/gIR41iGN/iwzXOEdzlwBjFT1GolBGRKr/4K9bVlnjqJpkTfRd1ahtYxMJkv7o7
+bkw/YTOrQVLACJpTd0ejpv06VdqbQQwMedCrdo+Ix9m7o9P3ln+kwANrVBPrCOC1N7Sm+g8Fihp
9Kw3+MHdQKEQQlWvUKy44UyJJDvexUmvp9FeHrplcJahJEFWBknuQf+Ojpflbr1k0P8c1qEF2STs
rNYiX8sXkoglCdDr4gIUnR54EW0pkBdxeKebVCKLtbNtFcPke+Vk3VR3hm1k/WiaWGj3CGicmcpC
XcOXn95sS2RsAXdON/seYOtCBrPjDVLsXQbVkeFXJRN2YXZKqJMwGTwqG/wO+hG6x6+QGPlaVUAZ
2rcO6vkiIqO7wlfJ++eigpbNDJBZZ8qfAgMAcr+WBzOuQh9WbhZEwo6Ribmd6WmIDeoeRMqLcN/S
HxL7svhyjf/Cw7lMeNNbEfyaxOGbkfPKvpTeeV8V7sElpRvMb/ImRN13OEiJRN2nx1oAKUxBDYhQ
5DZCEIO3gx9pFnqGVdu8taNS+Y2nPKQWbCjDHakgUSu7NEyLcJN2G7RDycaOA4+Roi5NtpbOlELx
79tmPnNIkpgQUxgvnMXzPOzg0PsOcdkbNFMgqQT4+EWLeVZqdvtayi1ATy8bg6rDPfOvCBVFY3ul
1DjmNUExzGLlA/1MThBnCaFEk2kA2c/naDhL9zzfRVGARTH8pd85bHMi1CefroGlyC/PtcwN0otz
uuMhz+7T5OhYi+s4eKgJPg18pIpGILw7XlMvQQ3sUUZlPzfPfIex21EQmt454xUIzVnF1991Hlbl
XV4X4HZTQH3YjP2fONSHO+JBBJWFEK8syZEu2rctQqTn+Z0xn77TgulrlVPoY3NVMLz0zZwda93n
/EtTCpxeUp9rnNilIFrpVgfRgZruH3Frkq2Kr0SDPlxOhURgQeHbe1FGHE5SQpuzbX68cjRECZDc
D7PU9vDr0WqBC3P5NMcWxv+Ji7qghV8x9NaN9ADYI+qaFH3NVzg68s1A8kiBvYCUInFlv7J/kl3j
qJoQ69wyCi4O946ZnyQ1dEh7psX4cJcWsK2mX6Ze01RSUOouOVC2IPl+CaLvcxkAAACuMq1N1n8H
U3GYIqc4bKqp1AVpIK8RV4A8kx+bYas0jvtcEUFu918YlLXRs+UH3u6gzbcUAv3+ukqOnfeYjtVk
8axGOqRyBsj2BUmsUjbsr9aR9D/Ha50aodzpedGByBlsh17tfnc4axnlePv649+S+b8slgjDOKAc
VZ/nzWBDe/k+KCPwYOQjMPACbEPlV5n0/EOnFBC+LU6zaUuWFHOeL26oqW0H2BjO0dHxLRxGEdgN
nBcWO/JqmtNz3M2Jtk/S+g8vUCDxkjVw5UgIzO6JlbsODAeE2JXVYi6o2m1Qfq0Jovz4iUuGotg5
rsgAIBt3zuZXnY3xEIc2ktbC45ZKkBcoEfTzI2zSJ8cS2hEts8SpjcTQKwjPyHWQs509UFp9QERM
dfvXWOxu15e6KwQ9E1SgBB0ON6WHALaUmm7OLWRMHwlm+QxY0vIsJkpAt7wiXjhMZAHIPyDSnQ4I
g/Fd2EL3TUpbxU1OKY04eyme05vbnFhd44Rv8q6o/eIgFV1n6WeApjHORDcSDgRcJovXZH1BWKAa
enltUIV/0JlWnrLl1jC5lnYaR6wKcvBvOie9lU77+dPEITOKPUETETtowG66OBdKKslrvtgPtFAZ
+bsScLfW291QLD0WXKZl8U5ByN6kSqKxBfeqWJLGcn005krGYgf4/ecTNl/wjCATpYZYV4kya6C4
IQjZaP1BvoV0in8ieKK7PA5NMVjQR0y/72tAN6JFutQPLnwgJRXZvriwQVC9fvscfNUvhWAw+Z9t
MVEq/9WHPXyDpZ6IQu5BsXwA9O/zm+vi6Kn0twQIectRd2s7uDlNj2QsUC5gzu7tHRDWuVT2t3dA
KhFwNPipTNT22rKiA4TghfP/fbJDeFeWqyRZrstGvsxvxGvHnuqBUcvvdalL2ZTN/qTnghgqwSbA
cD6PvU5D1emJt96wqFfoVkGLH7s+HOrcMbIOibv9UecrMWiDa7vILhg+2BQkq2N957iJpQhlMnCh
A4Fka/og+0oslZto/rx2zz4O1yxszdkmzvLO5xug/z5AaMbmaNHAeNnRBEWrXdRnqIgkxOD4m9Dw
cI1jKxchurmP8rBU4Qmjf2rmOOKiP4DkyAes2xCqtr/L0yXm5Sq7qQz1GRmze+a7SY1RndQTlq44
yn1DD5zfHAB78IhvPZWkfc4Jd8ffjQB6Pi+yFwvhp2k+eLp6DHFP8NKiYD1Rx+Km0KhKAdwxjk78
3tz7EVp7q1G5IN4i9PXH/BvrxhyZWy8GK69X/fmSOqIvZTUHl1xCVLsG7jqygijzsAPYQyCZpNZS
ZYmwH+Xry/E5/jwVKMbSkih228KOUr4bRZuGkvlGTE1E+WUHAm3MF4j7S8w8H1BJlQbr0AVyOrNH
6S/6uCmBU/kpyCXsVsJpUYzHjlQB7bhT5k0T1rFh5qLFFM31XxiUEioQVIwJ9CCURpCe8mp3QDxn
X8vDr6hWbxShEn01FWBUnWZLzIYuHlmxGvu7qU59tM5+SWQmQo81GpK1hyIBOmq2s+quppnmkYoB
U4iCJ1h3jTBRiJq0N3KuhVCohMTCbawNBcvLQj3dz56uhKcxEJ6deen+Z4W0n1Eqe1jxpPNPkpzo
3YR209bzGxtsDjLwm7WtciAqIcUfnNV9A78+bmTv2lIaTbTdYoDSzF/mgWpwnl0w9RVujzhTbFw4
qZN7NlKqCq3jjLFuk6iCvho89KhyhMPzQCP1fY7OBgxhAP1nglVcftWIKFuvz/W1SQeCFjM58H82
4NTrZKimBwcH/u2RGvw1NGCic/eGH+Ph7lmZOG63pRqUl9E/gl47VVSPQmEo5X6J2cqKsKbXQd6d
+hqFFnvfStXL3XoWbZESs+Myg7TOAXLP+Xph4OnAx0WDUmSHKWrIUQvx3qdaIfFqi1IlN1Z1xsOe
3mcnb7+SlCH0NDsmnii9KGev+0wX4d0kiKwIRs1jon+QhsojZp2UqrHNRaskE6eTeePqOePXEWxF
T/6rAp9C4XCYVsRy940lc5nwp/xaE3RufQlM05E3Y4w4VKT032etUkGB7n75ZlrKpdsy4QsgF0IL
nO0UfI4kK5GzbOvwIpZSFLQlZ9OBBUl4Kd4phtKs0AelCOS8FNs9cGvwch/EHl6CGA7NALo5Nfyo
5JmCT+Li5vODJIQeWv11FayGJIZKYt6ijPnrVvKmQnmilCuTeys0a1paUD+dROF01KgJjGpav4XE
dAycv7VYK4hdlFU1YjGkRmLOdziZm+cO7Kg1mWKaXAYblueeHY1jbqbtrTsiXt5JYXb1K8PNZa76
fRuDpS0Mvbiy7DzWXtwJ0fhqWwXg41NHDwcwUcvHMzaNtGesLGwYt6QNXngIKvZSNBkFUOxsa2oU
UPPKRXa7phOCKHUmrDta9R8ysV6QDIoVSt46BXpi+SdWoRy3XuW+UltgJTh9FKEROjGQrGCzldRr
wJN1p5ikzZhCp7tfaH11z1RaCgJXEqSUemR/ZU4B1vlR8CHxphdL8VLDdodZyHZa0ibGQZa6X9yS
nWv2C0i7qwPP5VEnQnLr4YaH82MhH6FhJmrOOxQwQBiDLirUpiIhtyQNuMtS94PVf0FksJMfj+5/
82tu1rI6fhlb66c8UPvRzgXGnbBh7/89rxy8fYdBn1zO9VLENVatnNuCgQM5Wq9CB/78q1gerukg
t3YOJ2IJIWm5TBfQ+xNl1hkYEeQrADINhu9xP7V77SQ+FIKhMOzabVtH6CL0Yoi3z1/Z7ZNdLXaI
zIz1ZGS9yWyWRw5Izgaq1dGL43fDufOsy0WxE8FaF4qo8hYZEackWEksxzrxq5Gic7jeDMTOkOtx
qIDjEG+86VzXo4kG2P1ZxDFWysBVtszMJ8iI4yIOHjtFnjsPaie8g9zvzUmTgD+13Kl+EnDkgWCX
/s7wImDnSqr9911LiLAA80VxkydiG8oHjJ4g7FKGYpnZBnw6S6zEAu7x0Mv90zt+jbWfouwLms1Z
5uiet9OHGB7zU2HvGxSRcoD6EgIljc+LpO0Fv1/W/iaPS2tr0RPGe79uKcFFqC76kOAai26KugGt
zio82YzPO9DLqncwfdwkKWRB+zx3fY4VkcbNuaNyKSZt19xjzjKPuxgOuyckbUKs+0F09DoESuAF
RAH2mhMoYdszOxQ/9VjoaNn4lEroPcsZpT8d8QaZw8iNa2sKQ7dUupUN8QYx0Scu75eEbX5P6mmS
QRFSvWYnpgPswlhc5BChdkz6r5E6N3/xBq5jyaAQKI0n2r3up2XwRk51Yw8l2mOO3X8G83MzjBPC
WtjT2OTxnugHWiY7rIxji0ncWaj67y3aSvqeHNoVBzufaBlPoMm3hk6MpWP7hvt4e7Res5QiLRtr
EF1ValD8f+USHRhXIa4BWJ7ir4s/P926oNEn2k+s/1czbG/bn3qw+X4ljG69lsuozDdhO5Ruwe0o
hiWVLzx1TjiUHUtAbBQJHJsO436DZD0DXHCMqGajq6H63kNFis2JYhUFE+b4LjO35+5nOrAh8Q71
fCVA/EHFCLIkInVC7nXCNqQrMdij6ouwyFIBkLysryfZCEaBuCI8D2pcINXQZZcxfrZgQx3Gku9N
fUJKRiOVNQ21k9BAc8QXCiOdJRMUDVvLzxxaVAvtD+ZHJ7qiJ7kxSEo5l8u+wc29mwWXbx8nsXSV
c338PchYFVtBxaRoE5tOU3bl4xzZx6TLd7nDzt5FHhl8KHgU/ojda6XCwPYRaO2pS4rLYw5xJVHn
iuh2YPDGznby7gR7BcT0QpSmbudktLBNEqESu8OF6UoJHrBamVVpoJVeTw603phpH8TwD98TKwDD
7zdj18UV8YXnIR6wUONPWgFhHkPhWPsucELU4XBbJcO8W1ZIQ9Ou454ySFax3aEMpTA+j0YMvgT0
45CebiE5As8L/AxSfFWYDh0SLUhw18JhmTlY7RiTgxROjhBj5jziva793JCLi7CQbMR3BpRASH62
knRDsk2R5rWX012t5oyV0vahfnbEvitwopoB6VoZeCPLgwv71iTiNxTV3ScWeq/Gbbft9Ih6Ganw
XhOku6y/+jOXJXHdwK2tH8m+CJ9FoVppeY5MfhEIEXsSnHY+m8RL0iWTyFp3U7g69kmG+sIzSKsj
uBinyctl6M2ZvOjHvU5xFYJjCY4oO9aSKl6YAKgNkJ/9JnzoqL62694b0gjGlthkn53Ewu27C1wI
w+92FRWIe2Q6vbWV8dHqaEXYdct3uFQAI0S6+0EVVV48e8vwVnHOiLtnUQ/0+cHPBI7vbT68Pfp6
/7AbCVAgB3FFXoB5Ndib0c+xRLIZBMPIJ8slpi3/ET+HgWWaUrlz7BDK/ZDNgf4DuEuAEhuQomcr
3wtk1kaksX5d6YEHbjYhuJtACPYTfDcgOhI0/5kM8NxoV/U1LEDAt8FZjva2h5nqmVBbmAeza9Yw
TLHygYRrUStWwcZjfArdmy8tVtL/o3EoVoQhvVmnwW9XoOjs4dIp4aKLuNH9GqhBt9Hb4ghN6a3L
fdImT8cmnTtEruNWNHmePbNFoqWSM/8mN2w/c+U4/OkfbL8SH7aRbM/6FXpWC+o0hA5JUCKKmDoT
aY8iMGvxqaqMNHsaEdQyIxpzglEGDgVZsuork4JVKQVoFl4sa8Ro21/gDoc5mWHEMH+m8aqncOcI
J8a4IPMdknaIKDbQZlg3XlYZyiGHa6q++IFMoC2t8avPxgYCEC9g9ncFT8QnmBdznhqEaOjTZSwW
IlOPVa9tElKF9JZpnDunn1GZTaqPHf1GcfJRUDUvQOTiEY0ptUh0lJH1zakcBPBeZVjMe4ffr6qw
NaEBdT+5jVYhnRVRvq5j37/HPrjOdSflvbziACYMDcOTklM8/MZ5Hh2TBKgBsh7mFcwTvwcL+drx
YfvJe5YMq19pKw6Owq1uCVk1KsiHU1Ee/B7aaFmMKVHNYljXRo7u4RJlGRXM6jkTQVqPlxiCiGWL
HxqeoxZ6kkCtu/plIVeFl3xin7uA4UeB7AykbIQMrY8u+dl1dGqxZ8OgXNkwUcDGRao2HFqi/wmI
GTI2Zq4tYxcfDKdUtBmGUE+CNPbLBT7WU1YQT739pifCsRhIk0TeYhFZuw5zun3Z/1BbQ9O/PjgM
CGlQccPbtYVTk559JeQZfyWtVsaafwr8Rcm+H6DayYeShx3GVO+IWTq6+rmqd/xBb3pwyLjDZkiU
7PvVqMJEaQyj7zNJLEPOfNEanzudLyFKIMA5Ake+odOxrGfk4aQ7iGEJTjLhImKHLvKeTAp1qnXe
8Ul8m5/rybv+UTdFy4ELxrXUrSeEb/EpNPt8cYKDNPoSQ0Ch8wKedLuKYs2X+0C2W5y7Ff30ACi3
+JrUaHSEaEXz9kHyfTuI5+UVb2MR/oXN6MBdfP+flVTPsrLC7sx8FILlo8fteSiFz0iAixEf3Icx
Ys3Oy8mxukOXCReZaFIc5TIF3qTQy/zHCB4uv8r4546PUdo4DtTRNHDC9QxQHxZnGsjVVjzHptLO
2bEtDlFySHvayX3cbbWj2V1lehlWow9wZsU4Xf7qZRLNjCjRtjh6CsWQ/YbZWu5kRIxxQOXeNbPp
rMwquQ0HWOwUHeFcAifk1PLqjvmZ6KeMnhEFv1uv3uCUK8PIpEYA9ATq2iJoa78FsEYaLYRhbH/6
JWutYvjgQidauGG2ig9m4TbRwdwV1819gi/py1lZr3jsaA9ddQZCfTp0LsfHiGKcxy74LLNaLN9H
H+10gv97WZ5XpHK9/j/Ij4kcVI1xtqhfrUaWQvETHUNy/f5FabhFYG4ofuhKikuyxEaTZLBsQ5w3
rYm5cMOj6vBmrZRnLMbKcJLGfdU6EEBHgXU27X2FQkbBd1TbDrqBACFpYd0MdNKwuEyBzCTdIjCa
Tik81so/nyGGbqJyINIvvnUuqV15NgDbN79jt04EVuZB3/UshxTR+PS1wBjTjhzs0n6btfWjn/A+
bIZkgr2wRY4xw/gtnnCzm6PuqnoDEVFkaamyOAVzIXXpMM12OckeFA0p6yHrctuA+KPL3/TGBYIF
BgtlQkso0jwCFt/98yNTlSFT5rIHRlwqC83AmvtQ8wWOP2M6N4N6zBA5ACA97q4do++qd30iHFXo
3Wugh5pQvhpobJfJf9ph/wfU8rDjcLBDRWUyHwZb4R5QCrR6vIWZnZ6XfuCKNrZPSSsWrNqf/Tgz
vbTcsCk+NCzAM/D4JiQmVuapxaqKwercUasne/FCf3AHk43I93JnK/u28FHfTsgQCgPjKYnHuL7C
tftPJavQDA2Yqj0Hrxvm21S9T0oDZTYdDtjx+9hnlOnvl59o5VVKJcTIu3Mq/r6gvy3AUrnSSGCw
PADQntmP/A0IO1qJPkyz/5CFLDfXDrILsJvKhxiYD6lVkxD8uuR95D0sAmFHKNWiRMQVaklZanJW
krP69YVN6TDGmXrwr4f9jHdg7mWPqlFu7SH1YJH32Wf/kLFJKrX8tsTefHieyWePBhtjMrfDymie
oiUcBuyRF6Og7F1m8BfjeFiK5NtXc17LOdnYvc2oUjAHfqogMwgvDk8ymGDDTH8OPDLei0j47lav
DntNMk+ilRP3sTMYng2CHOMLliryKbESLrE+bkrBrdd4Hp428xXTLVUPQOst09jEEnbFWiVU7NiN
jwuHJR94owPRtmVPQ66eilogdedV9qUKIsmXzqvOIv2XCgJ4/VCJm9w1UyxjKsXgLZb2ZtgJCXqR
XuVAipq9CGde34fz2IJceuw3+77zPmR5hQBZNgsZXlnOJRmUjQsQRJczjJZ3jqBtUdX50fRHkl8q
LcS2lbx1LXHC+3zSkdSkekEzeIi8ZiRRg2lSyFntW+91izEINuSSEwasKSTCi9r0BRzuAOi0RuGb
WuORY96ntQaYju6cAJTNKQkSYWjiDPmp0XFZq7T3fJqda8lDS12LSgotTtA+o5Ui/0CkZIh2yx8g
Y6z3GXB2sOawSSOj36Kk3fNke1K+mpUaqLY7KFRsAvCmrUg67jANg0eijqPw1lCT/sU8qJdbj5HB
rr/VoLMgRzGccGlQFuVtadHKSKC0PuY8/NLMPNc4Hn1/wB5Yp/AgHU2uOZTH+ykvJ3+sImo0DneI
7uT6PZmDjT7LkLPaf3Wifh7fBKz5pplkzSji795MAMbma9TFVOTuEJBkPcBG7hJFwCX57BD26oNe
bvyjLxAZAhTJmp0B4WB3mwhs2CZUX5Qcmsh0Fid/hTajwrCRwth0YYJPpBfLsjSSNiQGrMMdMMTw
a75HAf73SeiCb+gMHYLPECxA8fP9fvK46H1XDjs71136BoujGV34CAx0ara+XqidFI8CcFXRwBea
1zjiiau1nrUyuGMcKy8HXHo186VMmVHh46y3lTL+VCes1v05MqSQcmwWYkXM9uSUvrT4Ky5lqpt/
Nl+4hEYIRoC//Adb2z6qOV/JZEWnzzENhl6zfV9p9cQMcuHRiMXk4GOBQD41DzP3gwyrwIiuvWmt
UAUhMVdHNQ/vrKZ1ETZRP8gItXLVg8AokKpccfct8wczFeR3LxTaa9hEg7wswyYo+WlViGkJnJn2
tYmW2xsOMzQg8V0oG5mUNw6najNCcZkeOy0QP5MgqWddM6eE8cH9bL1nLOqYiP2MY/fDQe7WV7PE
ShVoME5UrZiZWuMOoj6vZzbkEVhYhgtD2CiRTMc81CSITaWHfTrrbC9wXFG3nRG2pbjeTRWr1Dk6
FabDa0GwHmzsVnkbhHoSXDVyTS5fZOH7UfssK7j5HEuaeUA/7CnrwvplUV4jt7mdcr0wqx4zzuaT
HIlLlQyNTNm4Bf0QdNh7WXuqz6mHlSWNtDst9J+/sUbnW4iXvF9iWmn8SXsoEOoXoIept3Ex7mXf
cRTcinnyBsEQjmUpAgoWYIK7jXxkFrW8HL3kF+38EKOWnAC5MHmnzZykk300F+UsBwbU5FYq6ece
H4XhY++kBJehsYQldNtiDkdSmqZT56NZG2bOEWIff6gsoB8k5aL6kjSjFY17SVkkgRpwVmy5Z9QN
wA8Idf63DxgHuisn/2o8ecCEMnWdlYTelpEtrOG7zK29UCbrVvU3b66p2Vcg296gb1KFE6BFwXWm
Q6DHZtobmLvykLBLuGxqZDMeD12FdzKCcy5iDmHaKFdQ2G4nv9B4xg5tDXvZXq4Pszfn1j/IhKpr
khJ+LqeDp5CgANDAKuMaZ92ny8D72p8GE24UQ7G8wtNOVIsQatdxDs5J7D1yjDlXtIEHBXE4WgGw
lV/gmo/kxfYZFi1Hjx8C4dzzCm1cPIyBR7ejnl9aU6OpU4WJmwIm8oKinvdDJG4+XqN6OjxaYsx2
TIAMx4s7pOOnCXJo7Lbdgfl7FSjp+AKeHUQ86EQKPNhCqZ6CzpXNGppqiqG6BI6mLBnM2hblDksc
BdEMrL3lxzUOZukIqzFiwchMxwz5LA0Hlhd4B48GlCeeDgs88MRKavA5+IdeOBkmFqpDkKce8/MO
rxAXkVwMxZ8WwKBg6wCeHmxwT1cHtw3QKqr5/Q7O6iiGfLJbKJclEKfI7v3gL2E4IuVuPKVnZCqL
sMvD9Qe9F4Vll+iw6fqOkLccf/xCPe/43UrKkT2NHITF/ooyG1n9mnWl+XJZEqoeljfqceHseFF7
d5UvNmmWv3xhWc67EegUMqQzhu5p0WrwIP0S9emnO8fe3NVSfxz/lQpzZH39WpmNRM2KExgOTI9V
PmawlBZc/dBq+EUrbhcmWwiJl53zQkm0ufy570VG8eC6ilatKL7A1URb9PRCFkpLLh8U1WqNKmDe
BDxSKTQAyWDLC6P3jJjYmFn9Tg1BPOuHtLt/J4TOu4pyPpsXwObugfU9+8FJBFTuIf9q15cVZt4v
uquD+cWAfD0ioaQHTNqtgd29ZkqAfkKnRaRibxvBCJYJtrW1+78eFvCiyavrZ8PVQ6YT1ilsrIZZ
8JhHGJVzFfhdkFVehg9vgnmxOqHihe4jNXU+RTWZNpKVsou/0yh6ZX3+DjsYIQzrLQQ/LVsuk9hI
GKaZhGIvxxsNnPdqUhZwMQxwZxByGn9YHnw5u6bGGca9OWRwpsf/Q+QhxC4XKwOov53pcvH/gZ54
rRVh59aOwD5GCnIwIC1trRl/F18uHybrb2jztYtws7lCezLqe05Iwts4G/K4LV0tZOcaFBdpd/6P
P9mGOmJr3AZQCE4Dx4gaKDZoG6mgVhyhEUDNg6cW465JQRoJoqmCDnnyUXHVFiq65jjXf4H0Mc39
rs5/rgBtjaoVBUvrQvgDggXM9QQW6fH58MCaGWOaL5DYuZmhN8jGeW/SXgiiEyLX6sMnGJaX7rhP
1IV23k8tuN6XioXF2iJIxw3KdTLoJFT2C+oz7u42Hs65jaer/TsCD9viMhtap6XQCgs5OWtxTM41
ozFyswkLCETzYcNAeiXaAbZ/kPGHrmdS8deSNE1jEE6yIN+4OB+RHVf/XN/8F8lGJfW586v+dqEx
3FNXtTcd04xMPPhGQ6uyQk6lpSpClh8XC8dCIxey1kQr1Xt94GxnmQAqEeGNamoxglA7/1c7n0lQ
KRDOxKPSTfKO/vaqsxw+gQoaDoh3vKSxKX08riDXkyptJIItlOOVjVXWXezn74if5PMnywVXD6yE
Gk54zm/mDKBFRvqCw+r2rKWlsgBJpcceUh3PuKoU8uMxGm/YV1raJtCvk7Th094Uik06hlynPzXg
evg4QI8Xn4MMYnKmvtafMdHuEsKj0c0qvVX0WlDjw/s0P/OOV0T8mwmd1pqR1AfL3RzNog3KC7qK
olsvrkQWqLhyNPPiiWyDPH6CP0VUbMPBbl2zJmosi2Db2VpIlz6velqYgmkncfC+NzpATt7NIbvC
IPi6Oj7WU3HUs7Or1Enad9tEhUlZH2a1Xjin2O1XzUjs0SuYSk915BN7wCZ0t9dq7O5t4THpAbwR
Fit4icEJwPOSFQj8ZXk01nIhOj2oA0nVe2ZkDaJPbBMggdlbXuiAVC3bZJ0L09x3sQsuFMcLIMEu
ediC0TkW+x8BjaraQAeOvE8j47++9NMN2rApEbvFhrok/aMN8/aBnyuuTT3fabbnOqw/UEGUrcS/
llni4AgD346I4dyri/SP2H1kYua92H+XtpPA01P52Zkqq5ZnpottSknygQLwa4attgBWpnfFXVQF
0T72/kHM2iceyqzQ8ZRy6bTQZoGUKeb5NDJ1lSK0nE9/9p4xEcqKeHePWCcrQKtAWD1GLEhN1PzL
LRJxwfm43Wor8r856SzwCnE2P3rop8bWGDndv7bA3EzzPyGfmLoEdBlZ9eyNc4yxi9+atnX2egqL
wndWB8StXz86R5ngpBytWEBZPnyNuHjgzR91Or5g9lcsrYnHO+8veB8MeygLEVlCjE0x1BUFExBY
Z0I0YU9lLaBCO9ksOO4z+cpg6zr/SKNA+vszVcF1qDz3gwIQsgpWVImkp1WvvyddoQq0hRaRdoB+
96K9QemCeeBY4+wJ+9vEg6YqnsXMoQ5kL7arTZ/kAJr6pJnLVeEfx3LeYQpwISiip5TAYlaBZb95
W6/RuN6a/U7r3MLITLuvwmjd7iwZRtaLjTCAsjZMziSaq+a3pHmM9jVi6BU0mpFmIyNRhyT/vQX6
hInT4phM7VHpn/kfv/+7NxjzDupv5/D+5ubrUPL/Y/d++cV3t0hz+xOU7e7RYn9aY3v7QtX+aD65
Ss3d3Cf9DPcxN6W5MZDqpaPvUXRus3EL6E+rsu0X/1WLw1SdTHqS6KSR1GGkXUpCrIybJ8qy1v6Z
i7nVWCo/dNmdlT8IRmMYKlwyPpkFv6IkYew43REb8ONuEiIRPigxHgJFZipbyKgkKed/XUyvRqzP
bhSsZW4du+VizizZEJ8nvXL1byuReFTCK6CtLH+vW7wZ3pdj5RUjGcZS2ho6n1OYt4JAum6LLH+4
TQZKwGzbtvCb0HMnl1+0fO9kEJanDeR/0bCCj+lgp8/eI1S6SpvYpbAJMdE6RMxt03e0R2yhIn0y
IzwzEu41FhgI2IpyVehqX9mlAQdsb37d/zEA/I12sspGrRw4IBuZyHdtjT2UUUuE5cxbU7ZO1Qrb
s3tsks2WESEUxsUhU1VPx10C72SBt5vMRx+uwxVPMGJMGkW1vTJeNe8k8hTrW/SV+oV7bVT2OeNL
aKdM4LCmRwFJnAL+csmsimy1zI+YC+eYKr72nFUNklFr11JN0ovDC3JdUcPEnP+HeiF3oI9l020y
iiRtfzaafdAP1ggPMpWEblbXqbTIWLbAF+HXxgPov/BtOBSnXMK+Zrmy/OeGiIAf7aioUumSkrOd
lfeOrsH7lZNQUnv6HdaLB5xMsa3bcDZdQG3vzstzAmwQ3u7fWvwMHP5+anSAnMkUtwu3jHTDGzk6
G0rPcr0gX29RDs8rLAVlixJwv0WU+WNJxz7NCb1nFY/lxeVyXwb09kVudYwHYjmHTwgm7y9NFyFy
YYq3AcmYy20WcSwdtNljN5mZEZBjG8+vjKJsUX7QKyuP51haY2QwjRJhfE3WSlms6Nu6wURbj2I0
iS65Lbo335TdGbkqt4UmlEw3euPjB2RKsEpwgW8Zhz1DhlK+2tjXDSt21AteY0l9zPHuG6/kOqcH
ku2dseGGj8QMInlPsTknVNTXKccC1TYfcTK6selC9QjI0s4jISNIm8PPc2RSEd8Sti4NkahQumG2
Z8IFu6St++nznKE8oWfhlQHPMhom+O87BQcnORC01wQ4Ivjz8RbidL+yqLZIAOSETSPl/ceNh1vp
iVAovfsBIeYj9MJ/0NShPER6LXJilLLXgttf9K0yj7i9YBH5t0EtDX8iU0Qp3pTyDcI7LrUeL1tk
U7Q/RapHmesRzAMAsp8176FSeTPhKEdCRLCcE5KpSefgHHdPaJcjxK7Rxp5ULh8irjGuRcbb+Cej
ILRj5wjinE6/XLonzIlDFOJMzoDcIcRvzi8rf9+VU1DehQOEUCTIT11uVYEAtNJLh1E+LmkFWXXk
UkeDyZZ7LC/R6YybEq0u0i3Beo6UwMS7LhkncF9/5/6518yg+MQ8oPnFLrVzGeNk8tcJMqqYfNSS
dT6kxtXYuy5tHcyUNC8ka5U66HxLww5yN3LmnqU8ph+jG+J+CS1AXZaPJaYuRlBLPlZdsXTVzVPW
qU+9H1sxrwk4YPMSKQnFSu/Sol4r/RZ7q/rSSXMvQbFmQjQwZ+QoQ6MX9tgTdKEyvaSIeSPqpyWJ
V0T+2ZTbWwDOwQ/nphsHTA+ahvff0oclMILQabJSyVd/yeQ/oh8WWNxmSmvYwoPDwANeBK9aSoRM
5ohe/rbBnkb+5HSXL/gwqYG9QWk04Zq4XdU1VEGnXU0wfgqXjGXEj2l23OjOPba+DW/2Sh4Ac0Zi
N+3o0dOWoe8ipcpssMfsXbqGS9WVNfeirPjYWGyfL/jIrTqcyhZK9gibI0AK8bSCjgVco6lL5CLR
SGkcmfJXyUh+1XEXuBDIDbkD0QR+ae2fucwNAvfxgtHrTFKW45hLWc0FytJVXu8C569Xpw04QSR5
vOo11qlhmBO8Xiq/rNHMCZKzjMD0fRJmAhy+eB+maH2TZW3b5j9jzhsK9Jd/NgomqA697EF+BTZG
TW5FoOBbFRwLPKMVMAUhlFQnlT1MM0HaGFCPcvOwAjQ4JOdYj5Y+S4DtK7KtiyGFrSA1IAuRqs7E
q76l8yu+hJ7SgXxJrjtku7Hku78WB0HayTZn/AlKSTGf28/PobOPs3IbsyOqcylMb/lyfMccU4wz
kaAV8RIRL+C6o+JX5djw+ipdWXvVl4q0bvT4qY1nF+Y89Ho7JJpGaryEN0k/nUY/G3aQT4XG425Y
TIeDdc+XZKiPvK8aZQhxZX8k8YK6+mskUekaFC6e9GFYdUvqhACJJi0GqEgb7HwCpHn8HPArAFrS
rdxM8BGudXd5J42FjfickvwCjfndL3mgqm8iyfgQsySREm43fPrKxGn6H5tk4NvEV0EoW+Vz43ba
ybk5gTOqIp+gqF/ZM+o3abFPWAlMZhsx+h46BEl4MvB9EQ4NGrNlqzZ5DpHZ6r90qTXh8FOADoDg
F2J/Ef9caR6J84WPM9jTyxs7B7gff7kUzG0t4T7KA+XxngL3hkbbsZASx3bSlHpH1hE44BmXLn+E
A2ZhkjEIlfbTJj9RLSgy+KKCghkG2hMh/joEysxT6+cWFs6anikAOaeOaQd5Ipf/bHutrbgz9TQk
1QuF1rK0WgdL7LAA/xDKbHkty0Er95ddv44TCFXfcqIDW+siOuoGt1+ufvFP/80bo2Svy0ByPMPo
66dayfPRhpl45Ohyc6iyjK8XMPRwSY2TwTm6ACz2y9eQiwucxxDojD+BTr9GoV5gt2B6HUV8ttLl
e2gIqFqMcJXsGMKRBTe2K6IiqTWDBqjhYQsNn1Tq6y6qpmB/AYIoFAWxlYnQzPrzxymlXHbK8IvN
n9zHnnfl9jR45kmrV54GmYaa7Kh6/J1ZqAuHtXY+/fVxA9a7aHIWhSpC5Q5nkp59s+cpNyYbIJ/5
9B7G5gsX/01p9Dw82gGqUiOveHl53+7+TUCKyh35MaT+nC7Y+ubcmF4Eck0kneKYR6LkzGm2qkCk
3/kslqZt5+EfdIuPm5h3nNJocz+0aXricWK17Dg06WeucU68iHXlG2Zb9qJav3tLGewOJdrh9WbP
JAgRrYVHngafAng4Py6kwnZjjUYp55VzF7EQ/2sddeJZHj9FJANzBDjGtFDC4F/FwuJnjxQQF/kt
7nvBsqCM4yNCzkccnvQGbL3welysX1/CreQtWARvQnyPAHcrjpYeDviJrpOYGiQ+ZFk8QtwfxOB5
IyJM10sg8Fp8SigL1ummRs2YYd66hRHovIada+6r9zyV+FxaZVzCHWB7Vn/eAFheSb+Yq6sthpWo
dkFGAflBLZqwZiFbo5FQShy/NjHy7DSkgLWIdnZukbM4Yi+1SDTsEOfeKQRxWquqIt/gvW6/ZYwk
LIcpEzhHqX0ZgDOWMcIMs/iNliMLfEXp2FXhgXh1Ge/YA+K8YjVear/eKDErAAUyyGflzC4XuUGo
NWuGXb9YLV5x9BinhRjuxqk016jtI04W5vgHHkIoDWJKc+fnLM5iGVfyJVSmywP+F3RQTbq6K7NT
lozRre0uuF/AR9HZ9QNx0fj7dA8r1y/u4nBUdNCsskxUKZ4KO/8iwc4g59xGnDqWuQJnNblUwoPL
4R1GLOOXIesGVHxykBpfzjw/OE33IW0tUvoysHuYgNi2FuONXBgTpyCMD4X5DKdrolcGD2cy1BJn
ykiSzPxOeUExnFIPLhpCS/QhpuTupAXPcp8L80clpy/+5vnt8iGMeehMdReUPZoSP3ezok44rRCC
b/MxIwmykKTRTyQQED0iww3evPIXeiRd2RwzhMOWGNylgHPFCAhODhVrtyoI1OC6x9k+2v6LexeM
7OzMUyXwA67FFgfR4qwjiJvZ9nZ2d84fgDcUlF32gzvdoSsLNt021NZy6rh+t4b98ofAnIDjSwu6
4XpfHxQ/c2j4iPtC9Dzz5mRVtBfBeUWnFeMLm81MYBsYeJwDEkG0qDtZpb9fiPHp3fGzXJgAZfX8
cX7iRQye12jN1WkqlK4x/jFKXxwIe7uJG/J0geI54C08WnBIkAwKa9ZEP82Bub+El3vNBVlcbaWJ
kfW331n1KZpkqwLm/b8iymkaNfF9skN1s2JkMuk82LJfxNl1er2Oiyo4W83Puc4Z87xISzPNg+nZ
t2bIw3EmYg2OvGIWvxG3FD/W43PwEM8LqsfCKhKGcZ0bwkOfGoL64ukkLwoWnAL0yrDL/kz5zv4V
YicYqiVFS8kPncBVuTjEHENaPNdtVJB4eCJjO0OCOs7azlthnSHV6ZVzj9/dE2mU3sDv/T0EcFPi
41KeAq261MPYU3xvfGALvFBqH/O+MmBZXN03JYB5G3K9nK1OAkCn7gXLwjlBW/vEcvpwSFQLI5WI
VlyumpOa5l1p5bJQyIfqwYvpSmQY0VYweKecqy3XqBJFtU5rE0aa4s2WxBv0XvohT20xqoHEYmjM
ef5yDOhv4VIpLwzbZclAGDXREolqLtBJ6QegZopQjKuAZItq7EOpjB1hz06P8l7VKJci7y7loirR
mFW96ynZvhgbTvEcwYYRyf3j5shislLAiffTIPw++AYjKiIYChBv0zVNEoBuGITJwMSucXCKdlL0
csMjSj3PSJhKZgTBKyH3fl1x3R6g5qFE8HMp3iuIujvWx20FdsIsCdxJLSszn7Tpuanz2PP6VGMv
3DK8aqHqNh3J8qhAygBmk9LRc/cDnjSLBK0fUzdnZSW1bg0RT9Rq1gwtLb0UmkCxiX3NL73qSLZE
zzSLSAvmLm2IwzAE2hRAqJuIxWzs351DEhVUtf0XE//40+6xq8Pm4kjEztiPT1+ubQMIrk+QXJgJ
zPv1D4BABg1fHBI9YvOTZDigoXi01hBFvKZCYPijpYQr9no99pcVYBV9dRDt1vIoGdKYX9lAIAmF
55H5dk23HdD89o0ND3OKgxFbaq/6rYhTr58J3/latbPjfsd1uf1wJXxAKeja8N635WSnQ12CNsCI
c1T14beG7S8PQNIc+aarTJ1CrHM6X7SEcSXIqiu1DczZ6ix9xfM+qVASmBIDdCLMcrqxUDttkSWh
juNCaEa738D5YQqJbBBKm2QnBdzQMPuy+tG00GvDes39jJRivCENDgobWKxUzUDFXIU9tR1Du148
8qEOs8z2Po88sCJpHDCgDqColkMaTQ/dTNi6VqCQKG380y6H0mti2yAbRH/rEOg37NM9J7vDQM3+
M3HmosHfG3o1E009RPtxOEiijeIpStRn7+4vfnSktXZt0If/8YDYwFE/JnoXwLzWjV3yuzG4b4hK
Vr+kee0vBf4PVnl1FOFtg5u9EATpFHo6ozkyP1b5Gib9+8r0zuOVJbFNJr+fa8J8tl88Cs4GOb/s
eMmsbLB8f7MneTXKQBP5EGYRiQQc7jmKdYNoe8twpYYwddM3IRkP6zCARyv+qGRehqlyWZx4sr5G
BURkhrU0tDJfTy75W/K8OQ6mZECX5ddAsNvWSjXLQIh0PSmczCmiJKuZTnWJ0bqrbJN5P9kHHSBi
bjqB/ioCVTErzQU2BqsnWxY66NK3ubFelZbQcikCNJ5Yfokq1G0yl3jvPuqlx+9zimAqlDeFbI2R
icgA7Eyxk8JdEyfCIMuq3UsLHUXiFlgp2Oz+Nzvzsbv4lEbFD7M/GaumjKZJ0mCr/FtdRb8mX1V5
Y3Co/OQDDa3RBB40ojSXNATFajfDesERKk5ucTuRgqVTvIOZzwJQ+JTrqfyBBIBhpLTRlVUyTy1P
qtKmO45fCSPVpe19Q+HTtdzkJZIW1T39L9Hrl4CkaACyA/b0dwL0Spq3CAOtda3EF6BzIDjA0ebi
Oh5hoYs2ycY33frgyAjCes/YopHwBFR9I3s56FVvDkhBD13OfzTIuPBLHI3Qan8ZkOVGVnEB315y
htKGmDj19hRum7hcmSvUH1w2utibg/eTnu6wVXXXoTdHMIASIxh/zaIgIwY0ZUMO6ulmGF+vatr0
r3oQkSlvWn1KHJ5oJwTahhz6qdMF+9vM6seXmFYVsuZdGjrnDFCPSVsgnNvlIWi+cCJt8yDe2674
5JutYWuPGCGpw3yJtWOBv3l5hCZmFZQpbVr7KuHdXqEFmh1aRfuHD/U8tURkIrJ7Pl5jmsqD1vAB
SQVlqRa5gLi3ocu3zM8qJbKnyvcOweKbM7guJkDWx9UgpK6lo3jRT0MpoCY/lr/MPIfHsPiyXIHk
73tP9izjrub0oivJWKgDQxZbgViBIidklTt9fjkWgX9DGbHQJVp6D3+NfTRVq59KZhD71fPCJcaQ
0osqfpyJ9HsP7zAwqsfCy1owkUFmWmPRniW0etKn0jTmMP/QA9oEWFT3wWxOZYP+w+6Bxqov54xn
EspgSbvzvlHvohepAshOhg5DPT4kL82UrAuxMApWJX4jntHwscLYTfmjkqc0gSCvIuEiTvtC7FJM
rKDOlSfsg+2qzdyk6Mx9Gimr7euZeiSCzHEl5ieiS1lqSsGc3rfOkvGjbkKZPtN9ixDG0HHp93wT
IJY/zz9fBsI2/VhXvZ55sz+GH9ntVB2pJWFW8aGGma/erpwcSID7kwJJstIGidUzEJn0oJ8035AO
IIJ6rFHrhoqFsYrMegdkFJS4SgzM3TkPjSs5SMGwGZjpLChjy9MEGp5X/+TZLKd93v4KOGmoLUfd
AetIWBxVPSg2WUSLBpro8Qcqb8viyh5rA0q0tUK+iHfV0+P21kG2LnShcg0XZM6eoPWC6ijJIa0L
FG0oLYGdIgtXb06rquyqh0jLPZuW+QKKLw7UYRjxgO+/LSjomz5AjC56rfpwIhMgs+Ra/cbUyH62
o67voc56NKIXt7xzzjz1CIuw6tY3KRBDXCMQvp3P/3Z+1+Q/FqXh3aKtIAS5w0OUs3pu7OCwI6xb
zwf1UgGmAraVQba8Xx7B0+DDx4G8BXj6PALCDKeNHRfcca2u2FOL365yJzWtAdtYV71ssT0nlx9g
09vFHmZJMuM9tM6wt/V/wR8PQqUAfC4LtsfInN6TQw9654C+skcU3PohsLOigQ/xWqvbBZ9nnuFh
6PnLImLY9X3NBkCxRddDnYdYfFrC2pCpRyTekWTG5GIVZg5SAszOnV1zpSs8HXc2JG50CSTLve/E
d/REty4R+vWO3MlAbVm7r+CB7k91FSrChBc3p5suWKkV1kGEf1vSMmJa7TqmEPifWBdRtE9gVN8V
Xy63YUwyEwE558LOBs7kJ36RWr+i6Apz+LOR3Eycr8mVx/dlTKgGKCDm30gRHG3n60o7fkMahy5R
F9SE+aRt48HF0gWC+1PECRKx/3WYND9efws3WHCTBuKAfGHQo/TgrDOMruZa1G7/jU2v6HuRyAI4
XXlM7PY0iwWOqdaiNgoPMvBEQoIF99rSviAu+scYn3tC1uLXjG50Xd/WJx1ejyMD155kYBRGgt/4
gRz4Y3VNBBk2KqeuOltD9yGFaJSVyk7mXTtxGcTPZYbb8Yahd7Qdk+VhiILEROYyDWNeG1tho6ia
UPrUaIYTanz1SpwaDpSKhWa8hpiRIrtm1CHEAZHXNOLIpb4ziM71rN2QSpKpiQSCcehnAc35nTDi
nYzgtbJGZkNWCUAE4iSxenVfFWeTt5XbL+W/p0xBwoQkw/sYa4bNgUyZJwtEibXPrK+OcDhExGRp
jml/50tl7YgU1mhtFWJGlQN9+CGaw6C7HDErZNnr1DYqZfl4Bjxc6fmfA41wKLorWVNo6PS8Dfvy
zhmhG6EWiPiQI6JVZ40qYSRbwz8xDNpz4udTB0JWf74j+FZGfiyCls8oD1IVm8oQRa173+xWkhba
TMDXJJp/8cgSES+3ZIgOPYzhrpQqQjm3GSfgBUamAq5fvRM9bqMSE8Urpqzphv0GM2uhUQL/XNQ6
VqeAYrt5UTS13BAyR/r/eHoA1xA3SXRZtWRXtGxVZTJ5Qa0RbdaqTICZrdLlVocp2hhfatNOipnd
A6q89gLjJWsecTmZanQgHpXmtf3w9PJNlTzp9QpEyYxHqaoAJHBx7inO3ZetZPeKwrI7kylhr9+A
K6Sckm0j86we+sCIhTM/FOnjpUicU9rKthVtKzTQ7Iz8bs21wXIKRlFLbNzWLWsujchvGsJwuPkv
QbEEqkXKEkhG49IlJ7SssYPCifPEL/UL1YrnNhAroO2koO58J7xA/PSpy03OrmwOWE7S2tUaRhSv
fUiy7qnYE/H6yeGsreKsvZEZA9q3MOUxM4uXScjC7ftay/oLdF00gUFAyYav3KyqIrJHKrf4LBAC
f5nhiK1poawyRpxF9PGxvBsUZGbiW2CGBAOfyDuu2iRyhuogBwVz/FWCSwNLJ9wPsgU75IBor5Lu
3AJNcNQxvoKSGX3lQ28bkOZzv5zeELYPIvoORj6pxVLJq/KjnxCUN59gorqNJw3J8gpxxKEdbtKN
EIV/VYEbcsyauFqSjWQeFm/UOS9m5ODEgikNRhwbwm8N45emk8WxnKHVqdqk71ZM0LcCaYefnSMK
zFUQmoT78GOIPJW4bvIoQCmVg0bDROtWcncPjEeHnNVe8YeGZBxTelYdsg8i3uBK2FUF8Ys88fq+
nX+pVI0mm8+BnaLMG1uGSyU3/cnrSz8jkW+OrAh/iKdmxun42cPx44Vs+KrTEXTFQmXW0JOeXYc7
6ZO3xy/7q13lmA8K0UrQ93n8NRfgOv0ioZiyu4zw2WGd5aaXLkPldqeIzVRPkAlw9rKS/b73hTd6
r7OUZQvzvPPjSqcD/kRPaU6CH4R5NVkdPfhClXIwhpfsvi/e3sNJ0qUFeOm0RCRhndvXfCRhW1PV
28D/4rXtkdHKx8iKAC7Z/8KlD4621CcfUELxhgP1FOzuyjS1QjspahqrVzPrxVK78pCerhP71U21
myOTPZ7Sk/DmBy23oLSiK2a6Ks8qqg+CGvd2f9mQySP0suq3tqLd5GqL38oUOoN6CS8OAkkpVgAW
lFTB0tnn35TNvRKe6rcWhl0tiZSBTQ1M9YnGzrL9E3ZY936C5pKeM4wTVGTrva2g/VKSukJj084z
RvWQPfHNTam4TU8KuE09ENNwbbvhD8z1z+q9+K8PeCDQat+0o49FXZX2DGFXftG9KVqGtBRUgHjB
xg5ZhgZALHSFS5H5vdthZvCOjWuuU0M67NvZy6AwGVDa6BcWZmbIY8+MdKP1KrG3tiaPuz21DK23
VHmS5zs5WECE9M4BVnImq0jSzs6eMQhpOD3t7PzA0wGn3n7OYL/sW1UPg8EGPEA8LwSs9zM8eTow
G2yLxxmdynE2uqertl1I+VzDZ6CAa89pdztl6EOdlkKuobAp0bXL1eLL2rX8IANKn+x8Rl3PBcoT
oMOfI62KYcM/JYWoosR5KuxGV8rmq/Ed/eR0KNvwoX9kdhfjquv+cRxk4r8boGqQj+HvurEWADkT
f+p70JXmK2SvgiZB/Je7FYWj0VmiORnevGrrlThofxECQpFTHFwoCagnUlngZpad6pkNd7lKL3io
5/+baZknAo7NdRt6g8yRkXb1/qS9RvnitNGw5xSRSvAZyG8h3tsSU5ZCkZSXDc/KMeEjIqo+SWRM
EYXnS3iE1sjm7oEZx74Lf4bGOCF/KtQkTcN3Da6S+LLLXziM7c8RLiKfz2Aw6TiRhmAwOCPwIGJJ
xQkgplt2rb8QUA4meGhWov+TrJuk5WMYeT4QD2LooDYKMjY+wx787Hdag4sOnsfqYmX/vRBdi/dl
zmjntRW0/sojv8b9D89O/3fkVcwIcHaFhq7Ez7UTLAY5odNxVVkBByHqq2OcUupMytLGMmBgCpg4
RAVALBLx+d9M8shlVouiSe2bZ3lN186otAOV6iWExHIk6lLmivuXowpOSD/eQBgziK4FKN25BOqb
vWquAIdl1rA1Ami6zEd3K8xGLK491JBKbSJGBwIo3Nn7gLAU/Ah6h8NlbMow1Eadcpwl44w/8cjy
moY4TGgvk+StunpM9pCLyhyRnL86X+51W1zog3vALTJ9PBP/WeyaYHbjgYYS60VCv6CGFOSXF6ti
Trq+uaHs9veBSXu5JZC+gSqs8PAD36NF2kq7f4yP65eXh7LzbiC3p5pNYnZnPABhuBNGJ7zEFf72
Yhf1Fho95DSM9QL29Gn67JljTlUopjfYdvcPa9YBbHMfQN8q84Vw/n75NkFuKtnf9Lm5pwD0RaXh
nkARL+V78L50Qn9rb/XFL8g1A8Mjp6KZyZmKghAEmExFFLc+9hkKHvKL7XUEmXimR7Fxp444Q+Qn
dO0zs6EpO7RPDZlEeqX0WgzozTznLP+YyDppnjx63mapW2ym5pDWJYAdxAgz80u+UiyQtR5c2zA0
GGIce8EODfYkhnhEJ0mnGI1AC+JbkUmbC5IIxU5H578+pZJlXvVGk1quY+rGktPPXqcgCPuoTYte
Mu/Wk5iBlVcJ8z9VP9bsi4xAzgY/PtUzachyq7CrO3aNj4YifV0Ls6lez49WfXkf/tRcYOBSM3f+
4hzvEhPH3Wj+jHdu8b4DRQd07uxpSV7b1MzQUApTapA0hJszt9I67DKwXtJ7lF7bkj2gL2Ngw+vq
j7Qp98TUMY8G4UkYgyHlw+FvyefNPrqDbW+EzJds+gD51rE2pCFxyAAJpnFgRPiR6EFvbqCkgUNY
Zsmz+fPetM0o5r8wa7migT05l5M+VnvV9EdaCct16xCKwBX6qdhpmKtBlboGoHHdZlavixfLT5e2
ceFmf5OhHmdWYiZF6FiPEUwFCYxT8liNy4KplAEjRH0bWufDIuu2CjhjQD9vkSiSm+JQl/goU4gx
8QzjZhBnpAI6jrM7YV0BOJO4HpgGkScE2+JXEX/J7PNhFvzgcYAcAqg88aGReymRsgJ8X9E/Ci0E
hMh0E35BUXL5SwVmaKWBZRAiYJKWbe0KdCQzTIbbLExY8QThRt7Px+yaumdFghY4w2hkETcpyH+a
chw/lPrh1QIQOMNVfNv2Qy0iV/6YDHKQqbuuk9tKdpD11bWcaU08UrKOpuho7wtVYF5TF0SnflHy
WQIEoG0NfGejtYdPV+naJe6eBXEA4QChtN4rLTH2fDhmBEqAstH71EfLBWmDZQ+4tkf4d9AHp3MW
JO7zY3sHhAlOwzMqEHl9qNMEp5Lq5UzKBFDWqo3NbCmDZhQj784gZX7rlI1shjenFdrDZV3QwHYI
zQJt6wrg2fDiYFqakuBYzw8z4jKLUDWCbbf7FHYNF+mVrioJqgVvLx6ucVdLMV3vfqpPn7jvhElF
SFXeicrldo/lbN8tfmGQoF8x6MbU2HgdTyNaxTgHb+z6AQbwMKjQT42Ji0g7TtUgXMVxKXdqijqJ
H27pTn6rhK0FcGbGuXWem0KS5Gf6Ylw6iaGXDUOLUeXoQn1kzccCRWCu1zCASUbikjP7oz/8BM7a
InFV/+4QAko7iUHkVA6v9bzrldIoFzq5ikMpZm/HKDPKfG6u7mOSY92ao2DfSSIN2qrOIQ+dQFhD
mllP9GFfksudMK/EhFzbMxpX1QNqoy3mD09uESmmUvQbHPSeOh4o4P0X/wODTigwCKj3bYIaG0Ov
hyzLJd0cofKZieCVDG8Sap96akK0PUSSd8W4mj5CC4p2TvVgFfZ9TbcSAef2GpqtZrhEFjbgQB9L
kPRibIN0quD7iZOGBNe2EjeOTsDPmcNBUM3KlRlr9JF0+Lwa8t4YqwO/MFnUJAtA+tTZKSovMOYR
eVAdGpu9QTgw9Mz2MvtQn/d1cOGkAOBiy+ZwNDDtvGZcSg92g2D6NJ0A7iwh+yvmxC6+HTAgDHi6
ICOGeFWQi034m2knrLwe3ruJ3mNOBtVR9M8QbvefosvIvy6yl8F4oZiUEpMGHnKA40tWazLRio5X
Gbq7mkxXr80QTk14ZSmTzqZOR/ISqqPfQRAkD7d+xZ/ApXkQfckpx3y/SNf3nfrThnoR96eY19Yh
2yFs2t9W6qiCnIlu8yOq60u+76Qc1yLWYPc1w2xaWNn3McHcW5Uf1WzJqDKg06OousEWkxXXd7f1
p6k6ch6CrDPKsiWzo2i0i+8FULc2FiCBR2VciGBs4TH3g6q/ICeFppetMu5Yaz2VCnQ7uYOB7src
DgOIpXAp6dxM5WO/PcgfroZxkAc9a2KXzLZPO1uZtBTdhv3QZEqJoryEvXmr5ZZStz60Bs7ilkkh
Gh3bMXYaS6LQ/EyjSENzduP0YnvA4356L3rgg0L3XNbizas3wszzIHFmZFboZamvweZmgvnon+5C
YkvsR1WE4QHg8iWwZ6cwR5Z5/l2+cC+VoeEnl5ceuTGq0x4mGWnC0cjUkboJ/4ug9S94EzMq8MxP
lHYK3jfCoVuM7MT/XnGK3POJxY7lpdg9agAU89OPZUXhtpzFIljbjDkLvNSmcrpKSgqob/no2Lia
1rFF9mtThnZhBykPVphnZknotYsuvmI85J6SeAhQpiL3JGAsV6qU+3jej5fGD2+R3FQ9GbKvvpkl
FOxHYTvztarnDlJgZ+1b+nO5q9UpuqqkuUspayDcUR8qSNJzw7zrOcuMB8Qv9sYsBWfnfCQqN0fk
+8Ld9sRZB9X1xtqRmzzPJ9hmCkPmMIgnchGMM5CZP0Q/GFkvfdm531BQQO+jk5toJGOoaxS4lRkp
7J7qfc6xQdBWZuK2q11PFQO7oeajfdXuiNeFQsH+jTUtEj3zG5DjwD28YB1oUmejjTXzD6Y5P91l
OTgtwQ3Cv/TFX38vVIvmvXS8sH0NSK8r5oXDjMwfoftjRtVUpCOb+20jiG/MXdkecJ29eSaEgQSS
u+40KJa2V5dmXNRW60WFrvsGP3vzchGnvCh/WUYtZAQnt0IY72PsaCl/XjigmXwleWr53G5RGIw9
arQFJ5A99k+XCbXatf2biIc74QVzarvJ4NMuQgaqwdNUXJn9z2Z1KLE2ir4PlljNlgYqHZSNchjo
m578WuJheW031QYWoRoprFi6QYiXx4aD0J7wquyoouK4vxOZMpPg7DTI7ijKbby3NjIxTZYCyGwJ
dsEruiV3C8IkedFPmXW+9qF+Vf2eMahyaoPUBMJUwAikv0cFAeGvHKNOW9NZno0phtrgo0/r61mD
1ilo5TsNi8wjcneHSPeMv9T4ITHGQr2EtSytSfPZxtWL/deUvZDofaZ6z7d9fTIIk5MVTBcGRwGZ
DnmjHPjJ8DyfKskpLoUAgED9722wRaXDnPAabLqCYYbpp4YNK6gtyB7v/NHftoktWiGDrqU607Kv
20gyLcJ9HUGn5CAn64JsIZfq6sVYyLNUPGXSYnkiYw+nncO6IZ5goqSLbcMapp2XwyAw+27D7uMY
K/Znx7yiJtJU25x4Tj5oBVuxVfpdVazcNeqH/puFDDxa38g0zZQWC+zFBRzSRgzRUkSXYBzJIJ6q
rgF1Zk15lsAX4Fqzjekz8p1MK+r7uQPGdQjCt0C41J0mio2ThBwdUTmHBZZrPi1v/mrWS7sZhoNv
mytWj2Lu8JlAE6WP1DCB+F/ifZGWvILQC+bBPqlgN+jybnX90rBH+0pcMwAiEAyKx4oLtWFLK0Hs
Byooe1+CymUIjIsx9zrqeuDUDAmubeG0VLjXeEzuXKxcGRWLV2u2Fy1OhaOeoT1tNfIUMh+BraI0
OemmSnoHXc90nyK1LnCzBOAjxL5wfJNlSG+PQ+Nur5srfJkhwLKwrMxH8mhYxXVHrtjlZwu/XdR8
Y8d5Dyw+ljGu1Z4OTQdg1G09NBBUSaSgCrP5Lbt3YGhdseB44d7FPL+LralxffTbkMlDGsktrwkG
o6RzTJ0fWdiDGpJmeGydaVuE2yIiWuMNgsFoLW8pa+NF015nPKG8QGMvAN4fYO8desdEqif16MmI
EaZodZGIDp6fBC6rnWY9jaXWe8Syj8KwlUi6zqw20KiRKDzyGu/gqkVrIoHlr2x2RRYtrtiPjMDO
oM4H1vgv6NroMVR6U8zWZFC/jPZBWGYabwQfDhRP48MKKthHx8Yl1sLllIUjVf+i9jktQXBh1yGw
CWq1L/+ub5FNuvCfdaVUwppRDnIua6pgMLHNk6v+f5+qeRU/gpcmtwEW7FGwWHvxiSsgZX4cFhwd
9jmI5TpOm0UhKmnmr7UFVA+Z3Lsrdq9SIqit/dpVAgt/Zp19151HXoNt08zWOkZRJRvtLYxHk/VU
gY3+9g5TYyR2jOBCG8U78FSsOZbk9F/JgRD1pVkV+2p995FAZd/Bvdola+PRUVlibgikimx8EB3Y
fq3MTabDtzGcsJU9Ax4W6/s/UG3J9mZqghjLC/UCue38ma2xpyf+fdyUjexrps4T5gz8LtpOh+yr
awsGAA2te3+U85UvzmJPrYBjH9Pr+lYSlhuoNfvf7gcYoym4CqieYMQIhl3Hhgrf4Jepju4OC2Lw
YuLdtJyudZVHiCzF9ce9+mHHf1OC3FH6ybsmz20maJQZYD/5Kv6EyXLIadgoz2kcC8VvMbVCj23h
s00DKKtLmYMuli4fiBEBHqp3wq9DZr9Tqg00A/8fDTOOtDYKr5gENDIBBn6VSFWhp81Tl7BJF2ot
hWO0ch2LWd1w/DCdYwtQ1lq4E1mnsL3JOsvCzTbFDXPj+7IfH0ILoN/no8C2m48AEb6ozD2OuYyo
W61H1K5gts50SFfpCOiqYME11Z498QMXjtHZm4YE+mMkQ30K08BKPhrzcMGlSo0Ytheg377lN04P
5YuudZisZl9RndjE6Y+ttAHznAxN6luRvyRH85YNBrRzcRaqN5Cz0XOrwu+xPlluQzUaFjkzFJdF
b269nhfDEowVFp7cSXKvpKL1gQqIYjnNJ9IjnyuhgU4M0DvEzRiH/j+XzM76nmj+HFOSVrDArT6D
+CXGtknKeGJEmqidQzlJXCj+jyu7+WTdUyPkPbQJbjcEtTT26VjA+FVXaQ9l+bnE9M4/FO7LRPmb
VSq/orcosIvjKsXMfub1DOObdJf8tdwrr0A4cgKJajAPbutWuDxrql9JdzJZbRxLE5BH1xEZFYfD
idGLU6Jvzz8h87MJQPf6fdP3he5rbiW7P5awtxWgMMgWG4zoVf0dcAXzSz14hX2+EMY8iArGekLk
uzucRAOhmy3Fkjq8elW4gPYYyA+pIfmwyfW8cJ89dARbGH8F6CQutBnpUlUxMZ8Vs81izzmgRbz8
6s89u10E+LeM6KT1grEAOskYAeWfvvHj0ozir9WFHEyY9V0s1FKE4Se0fNRN+Hvb8vWAifYoV+x5
KHDIUI4EYVPL292cv9J7+O7tC9IfFhAJrJlSQ4jjNFAnUgWK47D2JViaq766MFz4rQKbVYpw2uWW
zJaAMYdivmxTa5j8zznvXkTnAYTLoTmdIerfzQjxDvUZdeOkXf+D3mt65jZPcwzzbJccsq6xpHyM
o+nfibAxMEAYzWm2aN5MkfT4uvmmlbXJTfirBxFx31rVGlNUl75/FYJoH0eP6QVNYU1OVQfvYOAJ
529qDKuN9C/9sDtrUPmQPW9GARQotDUaN0xGpNq1WCB3xDy0Wq5Kc1XbA0AD0p8cZFt/McQ2AZ8P
iSd391hxvWyq1rKQwPUxF9arKZO6kp7+GIXdVFsHvaxK3ZAZi3B1jK1Bt5w+9qnBz1lcEzvnfpYI
NsqlHiYIBrkbbki31l4zbQiCcrnNi2REWoypC1R750ljVddwQsKtwrVJVQ1QkRB/pIH1pVtX3+5M
OIMfF+ez+NBnDCQST0rgp7W3sIQ8nFf4v2yqwswpzQ02MfdLcL3TPfNAUTqEeO7ixntKjCYjweJ9
7t5wRC/2O6ggkVBHRhe3WcIiKxQ/j1A0NKrJxkRvvr2ggC/T+j7twK3nyKyuNBVxkZDAKVZB8iLJ
EumOmaxguWVpswYAUMbt1DukmJJV3lGwpYzYMhXfw04zGXEi1m6E50PaAt07+6dIWrIlNj7uR5Rh
CIGiyMrYwv0QhklIy1i04pZERn7NHhGnzJDEl+bGsMy6i+B5AJPFXPJWf8C/7hrPocvJu8+FIj5E
WF/+o8k/Umd/8249sofdaUJ+7E4LJMrf9PLRrmge2CITzCP5UdZ6vJeCiuG1HgVfUKSL3jrJXAie
YtJTJO4/tjebM6imE9daWTt5HCkxrqwlCp6W4rm68iZKF/5Wa0uxH4D0A4AdCf9pSNgztYNsLsfC
hL5TLpNIKoPmhObfw0ZwqfVs5Y6ZrvDPVgpOB0UZeCPt24b1KFtnHp0lCFcFUtAAkrDGZj2jh06f
JHR72b1PuRtdOm0gMasKMHVpRlmR18LEVhWrJb8fnn6ydM08a9tgT9GjxFpwOtt/dESZjnfWCgoe
XG4iPnGm3wmsj7NV05RrHEwR8UYdksT+qPHkJnDplGtACrbDbkVdU/0pzFjlF+uFYc8Ow89WUgCg
9k0al6oE6f9mzXEWfUJ6AD4JPmG5qqumaUisONqWW9cSZLJxyWJmPoJyqXYgI6/RCj6KogbOQZC2
I3PADeAlRXeOjWucxe2BFtJSPxFbsvNpEhCzk70iX8IjudyFNAmykAJgEIZh3dwu9ZVmjCYseopl
f2fNK5LWycIYPWFAktP3k55InVYBBmudn8f50WTj1ct0aycA8DvrOODbS3mgpE8rb3FjBBJHfWKQ
H+2Nisg+TXN4vcbCN6UCkF60PoEvSWUPBW7RTOjF7Eei9W8bxl+BhiuxAyShV8P9of569hrJYe/g
OwLXmyba7XJQ1SnVFVlqHMyPIp0CYuY/pjOn24eZP3Gs7LWjps2mWJbk6hLSzYL6nFhdgM60nA87
S1VspR34zo8G2iO7jELy1Wh7rNR59CEdyd8zk4CcofMI3jAHfY1VJRqB1IdflMawKU16hPrkpTwz
PyJ9JUY85wj3HrC+Vn4cY5CcJPCllIvqvpjOSblaKesa1rQtbnEC0Tku6o9DQ7GcbBqtP+MWk0tw
O0n5zvmcgbAYW9cQlc0gyZpl1KNeSB7YFCn2oYroNMSHSIfc5BcsY041V7DK+vYx/W5fJsq8lhyy
P0J+5poKCEoctRWe+PaLqoCJPtTV1dKME5I8PRLHn5+TL97qSsEHtE9+6OI2GfkFcNUEpcU4z79B
/U86t6Q4/6MoVUMqhFqHRZfI2a6bHY2MvzisTiuxIIjbPHhu/bXfa4fNj/rXZbpYEabgIvQfNnBk
M9aKOjQEM7Vks+BekxbYIHP37g5TyC8hNTKQihnzRgYNlBYwIMNcGS00k1QFuk0fEakAnLOrSPp5
RAdb6XuaOp6icbbW8QRi3KPIuO/8Z1Z0AkqFnyGgbQoK6HhO8u3bSZp+HVYHdWUxEuUbuO1+5CaE
RcILOBubPLi5rB1AoMTPuV9nbPxI8VaXWCgDasmDMmiP/8tgzlNKgneWoIPQ82XmRB1XniW9sdKX
zameZY/1CP4J0ZgRGsqISMk+ZE7+dBZWmqcGtSJVxi43n841VPpL3KR6s4PhXmG6bk9ihQ0zsD7Q
tG1hT2EfnQHcGLMwlIzPhF+jlZfuTJROXlSPTNNcog3L1dMFjh3+/KzT1UlEXnoFOhKUMl9fTx6I
rNMUUpfgunSB2IJUSFOxgJpWromNc3GafsERcSZAU++AeHLZJFm+8SGIskBI3Y5yDFtqtGkyh72b
yyyiPR8ar3IGX8AVtQQiQbqi24/pok6yUJ9B4k/RWAaSNhtqlZvPkHmg1U+SViuacCWlcd8nVZSa
DMD7s26wszDi/Uj2RHHiuUt+QPwjbnNHdmBU/OB2ExnwBAGjseeC/ZAKH75P6d0b8WOQPZriE4HC
yIuE/S5DH4t38eDtx7sg05AcXsJuRo8UCGl6qWRWDK2d63Eg2aFEfuUjiVD6E9+1oRj2t0jiowdD
Kd0LnrV43cFjJEXXEORn8Smedj+r5SfpKRLNwqDnCxyjz5Q2NejWNuhZPViV74yzdUQmair6CkSh
D50oT2irzOmao6kaMUZiUvvsSLq4jEFeHaW71CQMCgkOynMpRLjyP3YN4t0h6PlHh/Ru76e6iD8Y
DhNinlztz+igRL0tDvemri3TYc8u77fNxEJmYS18roUn7c1NQdbwpRA9FZ96XRsjWInlrX0Q62Y5
Y8qiniZUKyTI1ZOGSr3r5ikOp98TUgzcy7Sf861YD8vys+pAauVbcm3GjPnHd/TFgSa1hT1aSELP
s73FqXSfosYjfmcjTb3MNYSrRW9Av1/kQ1n5E3gBMP8lewei8UQRv720VIDrooUGcr1BiW85P/Rg
GjThSBmfDal9hsiQeVN9+wh+G0Y75uLkMteUQcUnJKI+/X4Wn5PexHqGosvKHbQ0nWLMqRLXv5vR
rfPuBPA3/sYqXpSRGx99wNR+aYwCyQwqgIthDYFhmOHZDszSB5XT5kaHi6ipNZAQxZXNgWvTH0p8
gayywXqrQ2IrspnnajGGS7inQ8KP67i3RxhWr4fNf0zhu971SOGvW0k1JmcxCeB+AGTvYol0Qcpf
E8/HwJrf0g1XDIDXuKonVhO99g2pwihfFJNSsfCL6jzY94UxMnsmekHK9dkrIVb6qzSUf971paUw
i/Sat3s4iEVhap64b7JZlHTSmTnDrkgqHtTS3PtfMR50ph/BsuBfhJwr2kZwZWh//frpfw3tlWkI
mEGbtDN7gSCx6EjoPo5fexNDxGVwMlHNQ1lQpT1qmNptNPlD5G1VPXvFCeRqlfwmXkd5ebQRhqRH
RBx5RQ+C4LiZRrp4M3WO7ApDZfh2Jy4CJ+lSOODYqG5KO3KhBxVIkx3dw90uZbW38c54llPJvkmh
L97Wj1JB/ytmARxCuurLuqiaP1pNeO2krxaOa2LLzQJWtmXPzch3uhxmA25mEqoQN0T0du21L4UN
HHCdKGi2v5awTG88PW3uFQkavKKKfBlLVbHYgrWVS7nA1OdEjScehROiRrIrSISz+WwcC032Yz1N
05nqcoIFEqJN4Z9VRBoQxnERbMbXtxG0d/iIn24MGXDWJsXXvHotlqIv0iYIrY3VoE6hepVA5ka3
CIhw6yBCwZsfanzEGUPWx+1bUwOg3yvK6ExHAiaqXlV0uopyVd6RSKK8KJTAp8uFyHu6+7rJdGz4
rrnjLP4uPwwQLb9LdwQTCgX0GkulRQDJLEHM7T/qbFvqbQLCX7Di3IthiyDQYoYYBjdMy922PSgb
Q4a9HvDIkISsWIGhHP1CrKxr9q61WCB9fTXKedc8c5blRVgGlbE1pWIc0yUteNujtD1JCUr1cHCQ
Bgf5wQdZeNPDzmrENSL7T0sWEPeGZ2eRfYREZhsDg8JmnCCMzgHpLkzLL/ubc8H66zqz887sq4R/
HBtHztYZccATrHCoCpJbdDAzd21TaW9hxtsJOhH7AUm935fKG39IcnxUi0NUsW6XjFCGiAHsv0XT
Ouda46j2zKspdNO5OGdno+ki8eTab97Nz8aq97Yoa89KBaTAGtab4fjx6WULDi+QIDlkpA5fgZ2b
/8bXw+ispEcqnAORUPO3SChvS4JtftbhfFQBKdqMQso3UH+rwdyJtXGJ7vPbhwF+IIJgFdKx53En
UeMcQqYG4uYW2UyxR4BTuQkxFlxeoN7Ld7oG+AcPFBmk0ppllavaaS4DSgq8CzEPDJhS40JlX0fn
IQFFqzSeBZ7Od10wcPPanzmbIIUgDIr1CjWAl970vpRt1XIJTwzGcf0O4hQdQscYhxAkbQKOhniY
H82AOP2ZGKd+2XoA1MdluxNB/IttOQEo5TzPsdo7jsuvOarPBCjETJVJxY1Mta78s4nmhv0Sc0ZK
nw+Q53PEj/pCgw3smYBfaF6SbCtlwTOQ+lYz+2idZ5PPattVcvGgaXls7vXOnRXKNgR3Os0TuFHf
EH1+OEitahhEWV/pHmqiqSHRgWbdvFKfAHc/u7atQHx2OsiJyP5fpj5/7U5HT84UV7NhXbWE9otV
fn4v74Bk5YxiTWGlHaLLwM/vpQrerl8qlO3bHoNHFeYzXozpgG6Y/ZQ7c7KhwK7GCW/4AI51X8gf
NgcsENo1/V1yS/KNPLUcPcyLMiaIfqqUkQN8qSrxBqDp5zEzuDWk2e4uQInyrkG/KBIigsP0x5fR
8Rc3rfl365KKDuxaQeX67YJsSRHV3kOyOzftBEJIQ3IpwX5RwOTwjqSy3pJueXDYCk1B7s2UkvN5
y7irAXdnHtBVSg4umur5n4Dk/hy0SScjAqnWeJQNpA6UgYJypCcUhw4M2fEhD7xRjR52BuSoOTzR
HdBDwiYvmgBZ8u0D/btcyee4DA+DYmS9CzJZvRWsECXdO3n+zR9DVBoVx+gEDfW6rsPj+2geXTKc
hz8sfvXlPB10vBT13V1XoI9oRJj9aY29tFAjioFUJJHHGwUWKGdo6rnorB5mXgpE5lvR/B11eoGA
muc/uYpGHUjwiXwN5zekJctgLn7Tco9I6KFZSevxHXI5D0bB3SA4QXZ8cDlgabJ1FcHKGOmt2YcG
g49aD2TygIc8FBvZMx60OTNadBT0zj+GtUGWHbjjtGusCvFrRCsBBaNx674AaJE2/msmaVjqoGgz
CxBosQJJfdaUKbQhfCp0HyajJj53JSHG2IpoHThgn8xHT0WgsuXzZo2xgwfKPXAuX7ZMz8zK2Pwr
x516IvM3OI/HFv6CnOC4w+o2vGO0N+/hNV5LYG6n9X1qUaij/nUe5+Xp6F9j/SzmNGqMcz/KjOzg
fLxnEGtY2c6TV2cUc3pRhwqMPwTiToEHuvHGXaowyBOYua54HuWiAUzht8dvqLXqA+he5VhiJ8C7
+6QD8hM6Vmsff1h93ON0Fq4LbH0TAGzNneyUYXVTDcjKqik4oj8BLTa0VFIUITL6/S/XbDNvpsza
RA5Zz4Q4pY52pxHp/jbXMki/PTzI4aYNsZyZ9gORbusG1DkZ5cZIz8GCU4TZaH1/IUY9KJQqrQQj
ge1QlVQUmn2I1sUAlsubx32fJwb8L9vQCsNThifOhRpz7UWFHgOa9qEFxjr93KejrM+M34SZZfqf
HONSTTeXDfgpu4WwXMGdp4dEE1RLS5ALZbfFo3Z8FRUjlkQQV+FBo945uRxa3hfOyevPot4l0OQu
RzfWXIQ+fYyAv7xxKGE7YqdLrOTnEHVk9wcsmnrGXQLmGjs60x7zvcDEO1wCVJb4tvfWw/Le5A24
k7Rzaap2aV5eXz4lJo99+5vW5BRG+wmetIfNWEYJfemb8KDlSKUp5Ulv/6P0dmCFR9uJHYR65poK
vBhlEDcNR96Q+8dhGgZKPcSrbdbYcuEYBafIsZ5Nr7XJlCUhP9HR5ahi00KxcvEASHe5Lz2Qyb++
1OkkIPCPdb0MupZsJ+0pmHYtfZhU6BRAm3qfFrkQ4eKB2fzq/U3or/kVRmYCNMMDnwBV9Kvn3TtF
mCBZJu0OF8SAblwNBIQaypBsE3eBYGCPMd+khRWuL7b99eRWdo2JzkOcKc85xM6x23exTjLN6ZBN
OKoWnssZ5O1UMREg74zLzszY99hMPy5/Xc3iNOtGOMH1ugVn2j/qpL+evH6kBWztYtSga72uBdao
nhzoA4ufsXiyy9lfgszrS54qadltiREtBMdHhP8tDjutAcBaHtr8jjjVm5GsESreoky/dWscaLNh
5CCWrL8TCtAsJc570/QS+GOTYsgifgCyer597QH9FPZSs5AtAp2l4vAneCt27h2HLnDjFWe95wFl
UMYjWOl8+LZmgwAZId11XXk2l/gJSc9DQon0y9eQeqXiKJFA/mBALJC2FlYF3VdTGIn3ALyzbgGy
UykrCOz6cdaC/EM6aKUyT/84Zy/WnzhXgU3nkDMAc6qQMf0iuM432HQBcrkQwXmzgbhtu5FAl31i
8IupF0z8s7qzhaCllYwAWv2UNRsnCygGPppwMi3r35nX+A7PDxeZSX5QZH0JeRdaupr1JBDzJjgO
QQfuKuM3Dyzo6C88RF9pD4VCinjbgsnTeA8YdbA1RYNHwBUnQ1UI708XFk9kWG/Jv/gR3nFO6lL9
xEBNIsApHLy3b8IuCHTsOrlfJXEGonlNFv9BOTv4/Bb8Sh0e1d09fqZsvr6gkDELsOZxJWQkrqbD
qfPV7yRw3L75ABMU0rGpVPhUxI2tJ2uZ70dMhbCLhfeirXMJgBt+xtcX8JN6aId98jRTqehcBlhq
VJQMxqCSa7k76XGp/wjUZbt7UTT4EbWRPxv4aE54gcjgzeXJYv3bejhbG1eUf6s19UayfppY3dRC
1mh5C/79WM4wOmyPm++tZI1dl5qBxNgrZKQ8CXtxXPcnkh34v9TDtFSFcY3Hqp+DD50UxipgL6dg
Yi75IswnNDabGdS7jXW4wPzvfERKt0e44yjAkDy0Wt+16Rtnpz6U4VJQFsmaRZeVFuC2LYUYwCmh
eCbxa+64FDDgansvk1MJMQhN67Au+ZLX+OehBz3+e+o613KqcbUZAUiVA+L7NKHursBFPV0LCAHM
oGdlfOlZbLit1OSHZxmaW+QGtrIDDrdAisc47n8hti5Vz5leacA9DOnG9AkBceKqa/HsbiD4t8yF
Saa7+gzwJ/P/umO1Ilp9ciw9MWFe0Bo81yjt9U1BEYIpYpu6N/WLPW5FJ/UU/cpRhouQi57DCYUW
BoBTUHFEqeC4t41E/wl6gaJRt0hgG6c1eUqFY3J7hArKFXOw9pCc4uD45Bmyjm0meDXYTgLbe2xV
B8ehAqDhwuvtm3it7ZvW5Eg6xYogCZBvDaxR3ICUMttT8Wjbyur65ljmFHdxCq1IZHOVVggi8LJD
G2J7oUNNaJXJMH/+PE3+2DucSBJ9gJuKKAKemT2SwpLddbZDR5FqzhAUTyXGl54BDJ0+sAnTpGzl
Cs3cXAlMoBYn1N8C+XJcNksEaYdhEz+UoGk3d8VkJbfVtcpFjecsC+3xuUtKmxCI7HuAg1gYf2HJ
AuonqYSuFUgl3GH+1GBQLiRNmHkbM6x+yMtllIImrSWNB65HI+6iH4gRwROuiV2WGgobVKPFVMvu
ZUHIBHi4l4IHIYgPCKlZMcQBEWWFNlybil34op2Ztb62bA1pLbvtKOKjosa3f0Ym7f1AFTMrRnKh
iWC33NI1GWPQ7JeoWeyzKu0cMEhd7FXOcxSFBDIcLZbfMq+ys/R/6JNOnQUuW71C2bhT1j4KF0DQ
XDog0psMTvkH4u7iFgfQz6jz45kabaRA6B5FqgpksLXpuFz+k4E6v1/JKyu9B6boDQAmzRBbIqw8
HXHy8V1H7OEqpv9XPN4T0R5ntHcvTeygyk23fBbK0S/9ZADF5I94AHOInChJOOperkXtpcgO3zbu
5EZ94/c5Na+psKsJBuVJvLyX/mtW/cb4gFb+wF/UNF9E8R+/w7WCv4g75uTvw4Lmo+qwG7yxTVai
0bcy5g4LTAEhplNEsYeCWICHlmxsUyI2YEkBB/uorrVpzKc23rhRF6uRostspl0cJQe+rO0an8GN
wRA8mZrhEDyA4QG+0na1vIIfvPaHj4/NX8TJ7JJthI1pbXoceumPQvqQWdqFZd1qSUNsQIghlMLU
sBLevdJQJKDfqFScjSJ3RB8le7TYUFBmZ63ESrfkhGDfiIg7AmaixApDXAvz65WDo3AW2410JINB
9M8QZGXh6SItNhEF2ldXpgODgXUD/LD/3b8evfOBofclIaHKeMLygLfDHfyDjOZvibsHgdaWTVzh
pUeuYyKSibfAXSqXDndA0xVCNGj/kMHuN/TRa68TkPMNOGsz2I/aE5mluKX+6FI9Qy+Kfnuayk1c
KnDyN8WnE0VLgfMNO/3vKae/hd7C85K50TOwNtCY0Y7RujbPtRiD0hMyNLbGehDMuP9vAhjFr5I5
Pqe+STRwHsoKVttivxSMhyNUU7DF7Oh3SQ/asdEy9kDi2+CxIEl45wf8+7fYG1iMpObBDVgR/V1z
Brl2y9SQn/BFO5Fsz1P9S/moYHcZfgsVkejvlyczdCvahHEWOVGzmSdiOMvgG8NKw87cBNGzbMiz
+MkCVGvNjCbl7JaEK1EC8RA79Exu/lLNeRDP1Ib+Qjd3qDYXjKWKu2rVK0bRnN4Rhmpt7C84iL3h
LHswPPCbXwncawmqUU48yH+Jk3n8yfZWTJN5KDC65N92qEf2WkBNVX+gvqUVjqhbKJQ3NMUfbXk6
UI4ySjm9Q0iLL+81N8aZ22ctFt5zgBmxEPSL+GaEwrwh7WpJxdgxaizTJQfaB0x30bqKmeYELW93
eM9iT40crVlQisS+wRhkaTUs5HvuNF5ExHjIQmOZmqtzICBhkw5OrQU68Z8BWp1ui+MT4b9UDCg+
f44z4sG+nICmBWSXjGvasyPdbzT6OYvBkWISiH1EzMXBNlh4yi+/BzcgaKwH6pEyHERoYRiI/SdB
CA6hC3Uao2zZ79ILofEjSilCRWxshEAm+a98JsU8tmsTvgEOcfkESj9GUZQyw0yz2TndBx9uulOk
cju6IdBMflnJ53n4HKN8oYeasUOT6EidsAlpnZOhkkD98kK9pg2vHCSKcQ+P4IKsrtBIFOjJuqm7
94DZf/lrazV+RZye0p/nlZl3HsiJtoWwHpGTlacyHEGO1aDzb+70TttfZ7TQr6um5kqpg38XQee+
ZdcNSUkB8Lq2VGHoVTHCCq/U37dMJfu0MOMJCB5LeuZLutTzagpLbt1t2BCp35VPGQgKTSZSKtag
zDN9mppfecKwLs4WEF1LKGT92yAJeBbjq5jb4IUVw3BW2zsW2cjd1m6dCcFF9rbZJLmFfTtbdPt7
qqvZi4fxJ39EGo1+NrYLAXopFYJhL32Js1XlEM8BOa2rkDpqg97JvPWKZEUlYztaEUvEyMNd9NcC
Tb9DeSMIEpoxhL3sl1a3z6krMNGAZpjQyqXYmWyu8CDashQqcDPMHAhKsDJ1ASujY65yIc7Otdf9
osmBJzQY766XCxnoRJXploY8x/nULq9ZREE5zrbotgDL+02yu13qNiTn7FyFcpca0V8ycXmy9zuz
dFNyxLB1h4EVGsurz6DNjZSJ4yCgOJuIOzAAmUz7mFMWVAKvYk+S4bOMApgfSfVpm01psEvVx6Ai
ZqmEauFsY5C+4eM6MReKiSmHe89wztoCTSwb54FYzqPiZYgw4MfDm6b+GEwwunqvt6xZ2SYQKMoI
+pSwGTcMr0rCDqe1YmLs2cSRjRUUid/70QnLVPgcVJ5Kxhcl5hNTSialqK/JeJVSE1U24hkZgpaw
mSEIoj0hb5T58x+fYCWBW5K3IBEEgMCobKfCTaK+wRVsyJJv+Rnqik9vB3vOpz5BSTMo18+PFNhq
2sydnMpdcI9qEYiSLfImft1wH51QqAWDOnOIr6ZkPDj7oKX0a5ogaXkJA2aR1d5UBseAGWhfedLA
DfCR1JNJk+0g5QNLtx/NjOoO5ju2Agk+BCieiWn6AojDAo/JjJytDz51a7f085B72QUuriievMzO
gPtVZr1VcnQraU+CQfVOxAYg56h691K6pSgA656/RYQJ+AB1hutEyA6VAsvTHEAeGwM19DNCMvGH
H+CokprepOjOXFPZYkvlGkLskPJMyZ3bnOuGCHXymhrpAyTpSNbtJH4gv7g3eU5pMUzNrwJJ9eOo
nEzqsTAdZ7zBd6orAgzfaI1zoss4p379SWEpUw5iDDeu1PJuBJsZ42OxYZSglCN5LR8Yga0Xn4jo
JjdChb/6MXUFU2DydzCSBz5gjJcyQcGQfkaXWty0erKRVXxcSMTLciZfTJtk3LdgyP95XWd5zIIf
VZKkgVQz9ARaQP+7ZUwWsoKsHF37D3cRGGNkpqpzW205jAt5ffEnrVX/2zGwEk3Ep7+HDHrJYx17
F6VL+1DOjQSiKMF6ULc3UeZj3L9Z+juEQRhbNchgyJMiLSTXDaU4euW6Jk7iE0uex4pLSY+y/MH7
ke4bXMIpl49JJN0GjS0Th2Ak4/+w+Nbl6CLvwYF4qs82dUOf0vKnLoSz6TW0PNS9qsoLoVSTLS8L
tibf2026eCipfwjnFVwoHC59X281m7nxT9CJDYjrP89N/R2CgRACyYInbgHDxzRxE/uGxt46K+RI
XITpe15GpkPCqI1LJ1mbHR/zO/GBxS2qKVXW2AyV2Q2biKIZ8feguX2NUmw8tdy/a3RIzckjSebD
gnnZa3uO/aNV5uVBrTbTLInhWhcyZPM48zuPsmG58Gn+DvPtx2hpofrhr9uAzymVMpiWsMfn0k0t
GLHXe2E8XtDQrWJrFYjicZyA9KYgcAMeIF+uw9UkcPGrdHBqeb9obXWR+AgoXU6Q1t3gGLzrYemn
kU9wfgaTM4ICQNHgJcyDV2o8I4sUsWvR4HgWhGJ69IFK+U7g3xGHh87WBSPYHCVMQuIeaI0uDkSy
T+coVbMafwVJmHomUWYCxwp42OkBlZ+sX9GLXJDWsZh1AT3pOboHqDvyRaO0aPi+62XCw4Ox8AaU
XqPCQpk1HxpeUa4aK72oUBc6QZqsBrZTlJSJJn6q2lsWIikpnbG3Oj9He1BD+35nnKAiX41/0TPl
7t1mHSVUq5qX3yEK7Gwd6oOjKsuvPN8r6TXE4+ocMJm1HMUeD5cxqpoQJCU+PHJ7iZsZEowbg1Ej
8tCkYJHQtEQtY8cA6z1eU61nczSQWMk8xQEt7UXaRWa3RexiE8v2kZgmnRAaR7tj0cxLbepVCT6F
By3m/SHKP7IOnyJKMvGS6wnmfN8lXR4UxJKrXUE5oyAB+wf1t88tgljUlkduK7vJDRH+Qk9mhpf6
hiGz2O2vAcwWtuFKuaW/c5VTryvlo3coPAxNLS77nOgfqCpPbidEsnk6qpAkNyuHhN/d1GE2QRm9
lJ0GLsciCaWYiSC9i+j4saFeTS98/LcBzGV2byzs/wseAo5nojLsXt3fM31t67k4j4C9CtCT+pL/
/Bl5BxFzal6Y3oYk2RJimHatbpCW3AhYRQ++hrhOztiS3KxSRZK6j6wNtxNAWwP8ho2Nj4KfERLp
yb0Ea4hLbbZt6EMfnB41bSTh8/UhSzCgEB/4akpnqsF3HQVTYGOHV4eFQE8rppVNyboQP+W5UnZG
16EUNyoR8ciJAWc9rSzFjq3FPdpmYpOUTwyCm8gQ3Zt0vxJVdDyi0NMu3Nhb+aOZU8Px3aQK/tJ1
Pyj5DL9rBJgjmsH5n8MgeKzYh93KjzP+28N91F4CgcEbgaC2qxPZHmh+BYSDv/w7ori3Hu594JjY
0e3teFLW79QBE72Fd/eA2DblYO33El9oXBlqsZb9r/aj2YzjfVoKsWP7t6lW9J/qpUdzTFsDbVpm
/rrN4vd8vf06ivyYjGajlaz6dFKaydFsrBh3P4Vz5C+kfwzZn8uZYzJya7zXu7eFGz1CVOjdIouc
6JxlSm3cjI+UoSgb8bG997CqZBBrLczuNAPcaxvUIXhSlmqKtojPimubIcdAbXYMy+tD7hP7nD0+
TqqoZ3hs8TMMIP240mtUdcNNo4e8aRHQsILRkov5WH84M7losoxw/ywCoRXrwsovWAJwKSlNA8Cz
BL19dbGgloNthaLb6uxmhtsOCTOOZP8UX2syG67O9uQnJ8fyc41a+/e/rCB/ZByDBsTsVBDFo2La
XO/hEzPYsKdhYlsD1DnmwI7zpVNzsSG4Du+OfmiW6n9/NqZdwIglOoGBTNRJvrt3yxF+vzJNaqT+
zOYgWaqnP1cnlyAaf3al3oKuPKiZv/kZeV3bssFcBwfkvCQXOJGWnBpy5XuYZgvb457tSeO3V/vr
3qbljxkJi/xnei9X2DKY/vhjU6Iz/p2yPgXUdbQYxZEdBryF9Sh7Oohcal4g4WLVGdHSWRdNZUtq
Q28K5jz+OTOP5JrLnSjd7FmuMsortN7Af6ulpvrRWEMvgh2XdNbW9Sp/mVpQrDsnQkL3WCG8y6AC
meqP9BgB+vLYJt3oeDRpaPFt6ce7i25xX4v9vdKXo7FzL9hoa2I1jQpiH4STzoEKRJ7kAafI5Y4p
A65osgvjHGC+EPPkTt6Gn5x2JXZhUJbOZSFOlFDhI/qeeSpgDuS6eoeLX+BZyDVkitcmFXWv9xgB
VRWx+YqFNuuKLJ7MglJzHvYG+g+XuDJq7mo/Kq+TDq+4ENrwXrq6MHD+amHgr2oM77ER7YCwiqsy
gl8cRcVFH+O40GaBcD8wS7aQeczG0/YLPDgAiCl5tXGx9P6Vvzi3Feo2QdF9tXsooTyXNr/U+EBg
CrW31Wirwd09454R9a/fWN+1Np1qWzE0117h1xZAMZXx+wQNzK8fM9ottci45FUi4vkuckmDTk6J
+TMARSM9HOdKCFSTIttGxNENAKKJqX4eRbBzLUirQA/QfgjgJSe/IiXfllkUTpEAsafQgka2oYBw
YOuoyl57pN88mi8vdioNnKHJ8QkUzNUaJn2hJZGNyRWrpiepS/ovmYFYpcLVZRIbXAh+qKTpTvUF
YbczR5q8dyPhNZrx9P4Kkqc2PG924/vi+mpAky/zzhS0VukMMjoxLm0yFLx6rq3GosYpbVQ13cdO
Fp5QvRF4jcUYBn+7tIvHKPoP85CrH5MJGYpMXfAFmpY0Vx3AqA1JdmkaRoGeXeX5KHhqATPJarRv
hnHWQqr73jOLnjxkLm7Ct5oNaFUUh9epAyIeGfFxAW9S1vniYt5cTU+mH4dFUe7LwLfyIGD9mEsU
XfX2Blch5KR7H7tFSWFkXW6kL3U37OnN+2CU83ZuFuplh6degWJhOoiOUX5rOkCV/Pq5VzajNlg+
qZW7j7x37rQBrd4s8pm17To9O5iwatL+gyqc81PAj+NNUC8TnmLodiZzU7WxP6dwdoNTV4ZnTLZJ
NkUhFZa99UeMwJb68DQgcIdYDBRjmGVe9sIXATtZIeMSDiyZ24fD8HW8BUU0WS+TU/oLmi0272j0
xf10aQHSIXrktixBncZVGUZyeG0IvMl0FALzwhNKaHNB8+wlwbd0iGcpSLFE7DQZHvfldyXMbCN2
q261/KnXsre/NETU1/bwkU9jhUpuPYz+lnnF7FdGnL05EHjFE9QvrRks2MeODIio2wY4n3tfdor+
/pmgue7wacSClBH+lPugP9ZCGD/QzPLqQWSa8qBkjqgLr+86O6P02dG60HhEdpunZecLmUdkU5YH
in+7SFori4HJ0HNxebBxy4S9UeiOqgxFZh7PPimIOJvXPSU5OK1nY0jPV0YRcBcrIAoVgCpPaoZy
2/llEzYOM1bd3phKjJujA2VEqByELQQQaXpreWzG3T7csmSmU5I9cHLzdH2XOttvKsdnCKTAAcQJ
W3k20ocCm634Bh2mVFyr75V64ZAXJ3LPMPGsbajIh6/3qTCiZafVoU4NcFb1XKCQrDaTBg49WHzc
8sKBe+cGV56mA0qZUE5wOhM5NXMXEUp/gzDQvcDnv2z4OzpohbKm5sOywlRtiSxsNbSxb5OfE+6z
9Fhz4sItzVWo9ou9dBAfs9pphkFrot/eni5AlqR7jYl6zY05zD3Nbg945L+RSx86JJwG+1uTp0ER
Jd7/WKayu4DODnrHU5rqZ4i3xmCF3PTjN93c/pDWLNpv3yK/71dTnz4jdeljDZtxrKiMIXR5cb6z
pN8n/5k+FfdwMkAYhJfVAjOWULIZjYXz1omT9AmOYhUW2qTjj9FKAOS3aU3w9KYIG70bso4v05/t
BiLqgc311t6NQtbUVa9nFq1ZPLjtd1Qu5QqmwhHTDxfEbgb7WVR2lCybdcIudFxQzGCAeLqn0SKG
iNHe7C10qa4f6P+H9oOxx2vrxHuQMt/3yVTG00VeV6E1LCAsKnYk0i2Jjrspl/LZdK+CLtruIsGA
N8nTy7AuYu8G/IkzcRGflf/j+K5WtlZa2zU/R5g9pC0v/+pc0TSDupuddhD97afVMY86/HIMKIeD
akpwHBAvxexKvTkQTOKv4b+lWGNeB5EYz54Tbx32vQ3MU1VntEiNVxJDlG+DCJrm5tKjVRY+Mzvc
jCkyTE9/2SR12XYTS6nsUoN8P0Wk/WROwwppV+ttJrHofyQiCitfSZQx00h0A6l3N+QLiJ2lZTI1
Xwsm86BuDhjtjz5Xi2qDEY60z5mP64RJxOLhyFaaMvR/DnInAFOue9E3nBCSnSBbrRmvJQpvUN39
QpJK2LhFd9dig5SsGVt1Zc+CSMyjCGsdnPWOay7UJIIMMmAJx0hoW3m25KJkd9qOUgbLxlE/O3Fz
BUJxLBBqCCs6/uO4BY5yg2ZoXzWbP19wDXcmkRq9AC33I2XPdg8uqy9f4FPmNMaaN52NFf+XdYJQ
sDhRDg1kBMZ29sQzddvRtH/A9eIaiNV2BSXCqTT9r3YgiVa712uV5plBkag2R6XnFXxz/lBLLs04
6wqwVjEsfLflGuYGbdMIKTAHkMkLLyvm+GA6eLzdvqmUNltQYQBXtPee7zGitcF7cuoJaYKs3S4e
P0E/xuS1E9Ei55DsRNfKyH79AaFQIRGkBg8qAVRencwol/qtFqaIIlxdKZK2fCviNP8vvamD9iD/
oIRsX3POpAY4rsQwTF+VHBTVTkrreqoCUPZL+OYZ7lK+tGCeTVghMNSyz0Hv6eKWorf7co5sK+5h
WHHtfkPXE8vM5uOu9PekbYKMtN0MhlMnNRb/dczSpgsJ2gr3F2bPT7OmjGM9CZx8Wynen02Jnagj
trBhxoN1ZZHE/hl/51zE+zNznSn+W4Sac9miJS338IHVqfSqDYrumyV7eCjbx0iXpTIAuC6LNp43
ndLRbFZfhylsJ/MybW1ZqUudUCgoDnM6bMDL5w1bd1+3SqLExe9c2k8HyIVK1aC6nNYqyItl/OW2
yCtwY2aYihnueJQVrvvlSnAwVLpD7ZUcHLm3q2Apmf4Bz6YpMBXjRNb6YVWZ5M3Eozghg70AO9er
9ZoEj8soWGKCAge8HVoOl/6gyU+QTvYtssNaascfLQ4s584XxIiOiGlUoOsTRXSQa6cqJzv3Ttfz
Pwv5SWfEO5V0Ge4Pgudao7awJ71AlTS1F/oWSTgYFpQ4FJJSU8JnItQzlOUjZiBL1oKb+6Prswav
S8mZCiVGbXoN5WhEvunG+8ZCPlqNsexQ9KMmBAasGefiLeny8rPLNhSVsh65BwIFYt8Wp5puVBms
3oI1Ihih4G1a66SXykMYpjt7/dp/Y9wkiyu+VuX8GlodQnN73fNxlH2+6KaLv3U24+HfXcijAnyB
QGdC+P7/94Ypdxmd4HarIhdyV9RoUtO/ia1hdf0IoZRSPUvxcmVnRxYxXOhiyIxdzOBxBnGfTF58
rEFjZI7p0Y7un2r4jSZjWlE9cBeRbva+b9FOHhsIcTqGFZQbIDx1Y9j3N/jEIh7qZk0O18CfNR96
SkcumBgch/daPxk1E/NAMJUlEBEdHIXhjLL5EoK+I98XN5mCZbpRlHL3YAEo5W1tayPyHfJeTgDO
ORPSmPWJp/qdWDqpA2zC9Ulb1M5PLA+Zoa5zId1Zf1xxwpk7SZH4rnHDejfzc1NAIG57uyP3M6wm
TH80+sToYt/QzzlywpgeEfK+b9EuyEwPn5ZQmPyn5CeFxu1v0plPxfs69GN0oI9QagZVw9PRNaGA
FOBsmVgOdGah+IN7ekM3mIEFfKuuC1EfKwTYmw8gnMzpAjQuwZGqMittgWL4S4/2iu0oZgeu50ex
d1mbcxiBCRFT7FUmlhqCp+QFYoeIiXvXKkqDf54LzoUWAIRq1wHngmpNnzHibtk2rnpXJiJjOuK3
IdkOt4HR1iMMvs41FT3I/G9poLOH4b30p7TFGaLKBsG6RDToG8AfFYuw/7nUfUGzfcG5g0ymgsay
n1eNK90wlzY4FYcxOVhfy/zUMJ1j2tDTNuAOGWgwyzSAkTCDE4MnVOgMNBxPd/CygBx+RRhUjyb3
3aklACUxLQL/7iTKIrdQyh2+IOTMFYEWMf09Rd35LtH0EcbgjB4GgyBRpLXJGMhdZEZY8Ul57aPn
q7tjUrJTb3f8kFcZY+vypPoAwaK1af+s6X1RErVjtgakL24wSPY1AZDiJyjjAZ+wHbHhJnNX+blV
MqoxO0o8Fsw5TFT8hqBSzzyAQg7j7ZnN0ck+mNyi3cy2u9oc9IDAoQA0Mxcw7SiMhsPYDt8RHcBU
W2V4dQPMc+KKXIh0T5/sLAnoWun0r5tyI45hA5Sv/TMPKwvGblklwkx5u9PX7O1Joop19TucV1MR
qI5QLg5mNSWLubpgvIyLhUJy1j1LRu5byfyD30uQ2n1HXrBnEy2TwImP8ulkFk3Yq+sRBdUMvLfr
TDVn/JW+3GgSg/2A1EDEeSAAh85SP2VSEU/3qAmLhRF2AXQVQ1M8YW9m6lZvcyDke1yoOh+v9WFs
wv2A0TTW+pb0FITUeDALw/FmTTLZKExq2/OVkrVBYBcC6LHeVLmrm/KShf5+Yk/bfUShzzJkE+PP
iU+Qsy0cvkP18UGfmGtTJF+JxPodvO5sYuWzeKO96zdKQfirGvtKusi5/mykeGwGcidZ/DZRroS9
BiGwJ0exkVBY0hm0Uuuu9T/x7O2ngTrpyMlj3erPCY3GDCf2bG2iHrNrQrazXLB6FC9SkZb7Wq0i
Zd//nvrV3fzMgXMCmwCOYNaOzr+azTBv2ppGfNZ8+6TTqvs22A4sMst+Aog/Se3f/EyRjxM6SbD5
dY3Tl5aUuQh/Ck73DhFhdyyWmiFlvjNoToxLFS7YTfpJeve+rcdIjA34F4ppylC6n/cGzA6W/5+w
ZrzjHAqehVXxTZwgjc7HidIkUeZKT2kvdptFWoNwBFmKn3uRhvRrQrlp3iPmmd+t6a8jpthtCXcK
dAhaCWedYKm+DoWfsL9/qwzbhJqug6rF+4UMfvpJaptJlJjiQ5PIA2leOnYPbpZTyCjKHCciapTM
eVq0sEgudbW8BfBa/SnLevInSq1HsQUlzkGdMM+n48Bw8qIXvMCaxfQDP+PhjuMAUh25Njw18ocw
8h9ctd3vL2/ao9J2J3bGQC8rrttnWOweagpCi+i563G7pEHFDFqLZY/XeV36g5f3n18LzNEVXmKJ
/iPisTJLCt8g+jhP5c8DEilJ+sxH0VkKlg9sxZJkajoJPSRkUxrQr4Jt/0/KK937YWPcbQNto8OC
NMYJvw7CzxHHpH8Tqr1x6evAnW0G6K4EPlC98aK/q17ApZybAeYBjVUhz/PqPDsVDCmiyeYrHisV
kzit/zJN0Ww9e49kzQV9KLNWFEFNMALxsH4IuzkPgiA1jTAIwbnbd2o8jZPK4AC+k1aRJOT1Gzc9
wsXGjHVNKKlgtVq+TEmxnwvWTzyV7EKu8bab7yrOOYbqZoB4ZwxFrkiG7zhMCA3ivmyAzyM1TO2c
REpUD8QII7JV136neD+E1Ag4a+2J2+1gAFA7KW/NoKX39b2s40q6/z1jl7T7xifT+oHwrZGF+oT2
+MWIUULe+uy7ZFJRyKB9Ms361G634rvX/z/lpZOtzCfoRcymaQDgzh8X62r8rvZ3WloUSHinBxHQ
7pvCxleJwFfHGu/sQE3g5USH7c8fJSppgwll2WuEC/8NXYSrBosXi59XF9xa0o48Ey2d8cjyfhlS
oNb3v/rKAZQDA+IooRUBt3dcaTDML1K+cnqsrXxxORlsh1iwM3FAIA0WPzHYILLMZFoJ523/6Dt2
ishC9k5XvhN3hvdLQGi+By8o8L1awCrnPr4DGmiyr0GD8SBILfLIiF5at7TpaLR2ZBI7iPRb5QKU
+Kdx9cKsxCAjlXIuZ8C74LYb+L10Rmsja9g9Ep/8yhE7RzmrvP4tmT+73rI73ffxPCaGw6wX0Llq
AhOyiJDu3BhhQHFr0Z1pvIm6W02Vgtb0NmEf4ryvgwX8MtTkC+NgIEbWNjMpw8SILL+NZmNvuuSV
DnRPY2a5CUrqsqzeeFqYqbrQdO4VT35Ngsn+5rVwwpfYBwZf9kLQUZA7kMCWocbaPK4ygj9SI+/7
MdbnKpR5SSGS3AhLyL+WZyHQG9+Hq3/+qKVyWJ9mDmBOkBnzuVqO2GCHw1/6+ThI/sBBTihg2cOH
7ybs/nyq91fzl2nDlw/G6tUdltBtwzT5JSs5SPmMefurVrwyRVWemRXHIhxYLpbVj6EV4BM2deol
VdVQF1e0cp/f9d5SsOa81C8Jd6W8FCAleERqnmmrrnSCgF8lev/xd7GiwvAoujneo4vsAWtJFhO4
pNLpowLEy01NGzJ5QeKL+F01DaoIpy+k7tQTsTt7Jdfzv1oRkIuA1CH4LbNizawhR3w/+MWzg10F
acSbFWgUH6kv9WfVxykSSozy2lrUOYsY4zfNJ5qCt9PIcTnkd5G3qFx7Ao3veQVZBST35Dnv7jCf
ppbdxr/urdwtWHvFWLRXMpAtGcjvbDbBg/+dDlvdiCpBPUrvmKpMQGXXYsVbp9rLD6oA12IEodUc
qfbPCTcw8Kz+IjqVWxxysc84G3c2nmPpIRdv3kbYSiu5jm7/a/ymxGNxDzTjEKLAUBLtmTdCB8Ub
Hd0b91bJHjXF7RPPmlrgdbfJFRgU4NrNKHcfJ1IyZxl3nIjmFiaKSvcybUza0D+BeXGLkF46sKcS
FOWlpPIt48NiJ9CN/E40d9jO+MmNdYbz41o6rFCPYewTuew6RLHpbaevZM7ZayplZfsmlAe++u0C
8+21zpRqqf42PF5lihnoYuEH74xuEkAK0h2nq3EHeDExZF2sdYdKdzWEwbHO+CUM1YTm11ut5/GQ
/VBYXCsJhd66y+Ky5fNI0LHWvG8eApAWeP2lR6Gd6U7XAjluMQGKfP3uAlbogOl1BEKY5qH3bp1x
Cl7axhhfsdTAJgS86YVKsnMGuyDa5F37g8I6g3epDmH+Hfs3KdbMiQN2HLzA7plYXZwwtfZynibP
DvEz/kHJKWlhyPs+MOjTWJO32tPUH0av+U16smDla7Gpayj7pgoz6baDhaU4hhmWARH7DYXLnETr
PHfSCBETCca2rarNQ8fMJx07Id4CknZVpsM/ncvlYGzoXVmmXdabhWLvRohpn6FPoGBDXT9uB276
1npyyEJNgBXvCvDSSqqEnPKYd7ezSERf3oAZmz0yyMXkFQWKXv/oG66aTw69m1+46YwyrGEYfbLg
9IyHkpzmnLgU2LAxWvodnUS9E+MFx21Jfoc2Aq30pBWYIIbZr1PWERYfnLLFL7hZ8vdsCHnc4YeB
dPkmihGrsWqRbw08FKDE+JqA8AQP15pNPrz5ydldsoi7OV8VTOXoKVP2mOCS8zn1Oac2l9MkiHNo
OPaxvqV/X1+rX3PqIKFGef/V84mon7YfD96Gf5X0HLylSPh9RIAM3vV4YYqCEse1P7iTg6nTsFV0
PyumVKMIJsoiUjnBWCrNzofyCCcS0BgkwZZfXoMbP1qoWG6rYFZ2ssRZnsLx1PH/VFNt4LQoNTOp
b4kqjSFGbSPumGIxNfY7buRPqjktEy4/h/I5NQt6fezwGsGtsiCUoMl2Uth0+2e3uV6I1kM0DlhH
le4jwQcf+GjtUohoBq/4lMKne5rjsBbU/9mrHJofeRxXlYKKs6wFcw5uEYXeP5P5WfMECqsMeVWX
Oe4oZ8+7vTwVsN3zna18pEjbP0teDRtiKO7NksmvMi3UNlylzp3nYri2S33kUR7VIsEVT5EFK816
IiIQp/pNFGS2D5BqQY3n+O4B/1P1KNkphrD/e1tYg46puYwTwUINBoqtmVK6V7uZjcZHnTngaAFM
FwtvcD3S+RdsqQKVjY04IGeuWTyzIabB1qvZFC1sk57oHR4YZRahtKolPoXODthLA2D9YhMuV8lG
pF4Flr9jJ0XVLDdQa2YF3vn4PWIp4mhEULJlzipT/fDBgFaNQ0C3yjdvsxpy3PRPi3qS9dPQdCAQ
XY+Yz+geFa9F58CCHepd6g/rA3UKjWKb3n/bDyTNRxV7YHZCJ8GY6nqWJgRlZ+Ijw95dHB39dnoo
7we+d/aXPpND/mT3SQ61iCeeu7l1NuW6z1dwwnZXaYIhvNEgScJr1PyqQS8PkcJwgKgwus9FWRxO
t7d9ODhSL2ZCD2ujTMRw/rAnOus0jDuSQcOk7y4TTKCZmg0WKyheYmoCxJSE0wlzMvy466SJNkLT
AwYIiQyu6verWP7wazy0wtbSfDeoHuSr5THNOMziQg8GXhbU4KiU8RIpeDmHhe5GjYxxqoSNP3rn
7iq4oAg1obgPsyS7LlmL0fioFbLUyz8TdOQyVWSlGWVlvW3yejTmSd+S+atHJYnM2NPGC4nvJcgA
Z6kfoV4KGVQGgq+9f5QayKfsdsAf3u1vAWC8v8NvGKaaiQxG1WybuNdiyFUTCjqHo1MNaiLS+Q0Q
zUQS6RY3Ta5aNRvMSP9HG8TvhnSKy29p9kcLkQsTcvMq7saQRNcCzPASWCOSsLC6dqCAkTqabW3w
erwaul0viWAjT/BXlPPhw28XIAA5w5Gaw8Ib7BFXkQF3AI4dH2NYnbyTSg8Mfnoqwf1/Bo4SSvUJ
y9e2m4CcZ1C1FL8lsBgn3gbN8LrY7tcnK4PdD/L2hrPqlFtCt5vXcNSobVc7AFXsfiIQYp0TXcWW
lSkIylc+uC948Kw4Q9U+TSWuyVXdsx52ZD2AmAYk850xl9OzH0Hmq8hmEMrP/K23Lzyw4TqAOFFM
XEx6toIPt/phlteysAiz/oaOnOL/HIoVrVfGIokJsej2meg/T7C1nG0QTOxh3D59cO149n5kxttX
xjH/JtAhzQ2ZRJtpKV5EXkFlazsKcHYSYZZgHpqhbySUuFBIALxTsemfEb0kKx1v+UDOLpaaj5zv
8S+FU2yDyNdSBjCben8ROZ3XdJ6oeWdsU1qV57JDl65c+buBuhj9ZrS2uTGNNQij+Wojhm2Rogf1
TrAn2Sjmpj2dr3QIS8h8NYxbaGXkAYmjtJIuL89Fa5BppPw8e9R5sWD/20E6EAaKAK4YczXAf+Ns
XcS4IcGLtY0zmTVRUA2AoNf7imeyjGAfOLP710okvU4dm/VuAQwCvGWwtFbgubGvxt6BggSY4Kyq
HOtFwqivca8COlTI4L1KPqWiw7GlObgcT3/5GYWAf0FtgcTPsJIznyVJrVyIZTUUa3QIDaIVOEiI
OK7E+az7v+aXyTxeEPK1DI2JIV+Bzlt3OMR8S9jTdgA1EDdZ2Jldt0RUGeEASLCJ+mCuukoCFja7
iZ0YUp7xOrH83xi0oQtHTIH8fGQIxBFewAdKebDtx14RfHHcwlu0KeBdCkBd9IiKBVMuqACGK58G
JYkD30TDxMzJbqYhYpRTCXyXDebs5K7qLO01o81JHYhMMHT8rHOKTFVcg8U+shveBZfadqVQhbaE
XwqSx5oj8TUQs6Z0+GQIdeLzudM/a9mKI6ST30MxzITH+JXt47h9F5sI1yASSkwAZtCJ+BjVMh0O
wne5pAwhanDch0WdnAU1kSJCz6CnNYNT3YFd3mc1AGk8Its1OsV8Gs7eA4DYimfuYH+FskfL24u2
qN8tC8jSSIcd8l1x10DFlHyYcNzs0pffWNl5Yowovx5ozkY+UoVhSeoGT/6TY2tTf5PYqqaDS1lj
4spzeegIMNlPyfhlb5/7qfu+CDOc4EZHF0pp1xaMghEei7gHPFfqq4Nunb/D17IGtgdDrD4cMa1M
F5DuXbtQG5j1ylritKVHUVcBRAajH1+C1LWL8NBAflWrniuYoDTTTh0JyWSpRsgRLFGQS/vmkRZR
S52XAkx9uv3Z8gjfJ94auh8OXzSjQceCOUDRmQcQD2ABf16QO30QJ6YaeQmEjXUm1E3he7sXT/x+
il/y+at8mv73hImCCajSQAu0Z0M6U0hJnfnhg76bbQ7RJB0Uy+IPF5Hbp9yMuVp9NwWZQF3AI9rZ
qtHcTBAbLQhD4DGa6k9HLj6OueiSaCveaV69K6pTp7hE/zMC0PkHXKY9pTFFaCLY/E3scVh/LW9K
pBcQrPi6TPll0+x3QyTUr7zGu3d0gyA0W3TEARaB28/ozvvsZrlmzRyyo5FJC8TqKnbwpaVvxZOM
sCMXa2JtlotSc8Jmhbb0CuJRXN7f9/Xbz2v2QCGU2mF3NecYeLliJ/nC8rmIBJpUh9j+Ioj6YcWS
FWhP+UBv4acISl2ZKs5VUQBxmJcl1Dy7b3VW6JZSOBznNY/6W80kZhVp/YUxeNYjGjVVT/vKGFXf
9HEcJOXFFRJskpgRh9gTrGGLhZiY60WWPQ5Z9PMy3ClqRDk/vy7DZh/8td2mgFu9VzggGHI/Npg/
EHlryQSFZ09rDTk7ylcMTBvTQRjJb2VXHOvKkxGzz6hXaLTXzHE/maSp6sf2Pc2UoHt5VI+tl2zs
zX4xfS1cAtoRE6YtktHK6XsZT2hcXmEhdP+ppo3QRK+/8gWMINDtJNUSaPwlejqlrC6Pde0h7yJG
orBeXgq/Qb/x4VeBrfK5D4xJ+Mbv+wuvUZ2Mo9rUu1UGhRgjHo//CQq5vGtMZwcV4Th3c74PFKhD
EbsMCXK5YRE5u8Jnz2ZvRii9Z1t9nhdSC2+22nEH1XdmAvE+mQEDF4JrSes3NKyg2xqCxPdgl0Z5
4WUX+0xmczuWMzUMObfa97DHPlWw/LlQa8Mz51i/eTdM+9hgBxQ7Z9hdvYQZzHkMOn3lXZyIDKEl
ZmQlmmRspTmwQbDzmL8s8Ahbn0h1i/KSUOV7/5tpfl8qT47YnecjjBtYzNm5HR2LTTttMlW2GbMS
GZ+FHxzQmX0SByOdiKfY650l7uHpzaRPUOnMjmWdKh3+deOgQsODuDe5mfZTCUJtG96YdPYwowK2
0iP7zvwWHLYuOqSz0pExnzcl4944vXNrl1o+9PiF7wswUVMec6sHE+Zkvj44HYJZfW9pWGySceKm
RffIPnFxGIoVHAlvyYsIAhrC8YaVL4giSiKzAkN1C3QKMfPIi/8lMGFKmtvICsYWvzZpQlNSc+3Q
e6FRKPKoePQmA/5ic83sj+kmX/bvHbzFX0cuGrnDRv8rkbzPaE7jJ3vAXhmUxmTbS6zmUZG2GUST
JEgxzLbOBSKTtjZ6NqcbQg32HQfZf7yd1GQ67ddlzlf1RM21fC/vJRGDdC7pp7kwJRnYaGU5Ny8J
5CdNQLNo0gHScwip7OStiI4VEEGwMPd/Mui90SXTd4Ajt/uRh7YhtDKPH6TMbUWuG3QWsvindFR1
pxacHFAWk06jkG5bD99dkz0zJUCe7cb/bIaAS6zNccXV+mMXoRBTwrArMYjK4WX5af3oSv6Wv5ab
+hB1xzw0vwzdwG1skAdd0isWaICZC3dI8HJwPJd5LLMjk95F2liCsVNOBPm8caKQON6qEJdhsXP5
BK45QmBpiO4QJb1ES2rqAeiebuLVkEchAHW6tMgOh/lyBWQtNU0J7R54unaQSXkU/+FhbDzaC4VO
4Fj4AsUcnZ9ijdr6ODeNjLYz40OIla910jcDYzYuyz1YPKj1N2wF++jf0Ti9tWiAKusc1+R43Cjd
if5xJErDiW9NkbGu/PFHXar+7xGnHiO7qLmJK7uSY/4sTsoAVI9ZFTooibeLEDac1YoKfcwbd7RD
2WWrm5GbL7dtntXr8DbhL0+FilHW+KxQiSBqcyYJQLxc43SrIVLlcv5XXt3JO2DO7tPFgfDDBjq2
FHpZdmYwcc1LgqZFTJPf4IDHDbRywfUCLkJzr/5bULy/76gJHH7yiou/GkAtIbeCZkK/YdV67lUo
j5E8fbMeawLspSZARHyK2jm9Xn2Hlo27x116TNJOHi6iTOV3Rrw4mnMzaCN8MMGION6jJbOvdW6K
g61ofkpr0r/lNoq+HRQ+sbV07OuRafpTotxzQtyvHIEi/Axeago6/DXPNs20oCBKTF5XOrZlmT1M
HAyxy9QayEG2NOHJDcxs489sFf3AA7nLqj2jZTYzOw+vyI9elqO7cUgnvXpCWA2MsWHRTm5ggVz1
vnwyLtoqBCj76qNjI4+6ZPkOi5pP20o6XiKzkfaL43FFeMK//iBWA65IIE52uGW6FMRHVxO90Jo6
zNVYBuGGEF57fCv4x0Q/U1qhMLzAnif88vX4tFHo+7427W1QqYeGfylOiOaUcyGmb9ZxINqhNUTw
KskT1o5Q9AVSmxc8KTFkbOVix4xzolRYLJoNMXVYdcHq0OzBBdGOJS2pYDhjmbJQVMj+QxGsJpvk
KxEt/TVMz3eGdVSp8KpAyUBvWzM1Qz0a2egdU+FEzNd7BlWS6tKSzFkIqrk0NqZLo3QcAoxhVjhF
MkE842L4mc+/QHMD4cA0tl2lCYwIzvaPDbGJhAnP7+in6s1VoYIV+/RsSZmuinJmvLuy7oVE6zAn
P+sUSqIuAfQMGKQtoxXEcvKkk7SxEtH05HdIY0bhGSHEEoNLLf1fQ6AjS/BFH+e5blRALXfXeZu0
VL2eIUU18PMmfhJ35S1fnzxj+wH9ykgA8uXD4BkCExHeVSfpU/SypYAkyifhEMtOMY4YtbKCyi8w
BWaXvziLkWwX0fwlaQ8ndK5xcTJ/PFN/ni9V4yWKWCpssuR65ah4nTkcOHR//iTfbEYcogcOjCxU
wxtpEUNruU9pcqTJqCyLRVEXIZ3jumMcOYdy3VN+PqFOoPaBtjrApMFDye4WqXPWU9qC/Q0IIEPB
OYOhD6eLq8HsvnJ7uWEi+ykTBYqp5t7DULnY170HB9Lx4iN+fUbwJfLc34FYrbAhrZiw6+v1j94Z
v9j+MAHJoiHuJ7U/aTAYQ2o4kZ/zWKqj97u0zPMGHVOjQaE2ocOol6ygUZcG/m4wEW26FdFkpwLy
zbKuR+fTQpOzB9cp3lo0Yrv1KymOwRUGTwuLUp6ptXYz0ACxKhN6VaMdpL/Ndy0pyH7oU1bxGftq
qlddvoXwFglQtB+Wxjb7BDzxDRoFi/ELbtCv3jqMIRncXYGT98qehmjoTQ6XhOjCFBenlspXN+Px
iX24ahbTivndEcqGAComizzf+QbtHx2eS2mQmjBJ0ncuXE6TQ4K3a8bnvNyo1V4bDzckMxqjbmFJ
abaBamKVmf3iVHQ99T8zuVGmV3bxSr+Nf7mMG+o/fyayztd5c+XrIqY7u4vMOcY5HNUZXExvAFf/
i/p+4PtfUMx+imvUjIzSQXpNDJCNXE2kXQtBuJC/xnFAPkUBvjsGAY6Weq1E0F2dss0SVTdH9afq
1/aPlmqhZaj5XCzDAAiAeGvMJ8whD41zwsvLxvtztoR/JAgMpeFlgpcaO407TcOxnURka2H+2IJ+
I5CqjakzevQKEDiyP1V7URy7wFdrHrUkQ8h51BnKJxgb+6+HpdyPNE/82Hw+OqUjIQnTXydst9ba
k1WCR1LjD+m43PpAB23Hm8A6mr90gQpC6zQ3Q2cATlyiyTAyjTUX83FKJUK3sqAB3TiBT2J3u6ld
Lc7dY3SK/f3uQaZ3ZhjB/zCEFVD378VgYso/S2dVZuBseQXy2ZNdZOPjKHF0z3mS/qP4I2iLOA53
5fF1e3nhl8di/Dyv0oFzvbT4tPZexQMfrDuFohvP+I4rOMOs0CoCl/rm4Coz63r0qLWZPOHTy7wU
SQ/P7cOvZfK6cpHUh0J5HoTtnG+T9iQFjTvPBHgXy5ImeBQgcoxWTLa4vSUROWVAlaYoRa8mi2Rx
BDWRsAioBdZNqOqABY7lP1vhTZ3lD6HH9pOvZf2auOsFed2mHWLgaZ7vbTUYCwtmsrDwLRqu7Ew5
3GORoE4fDRi4LiSG4jbQrRiaO9heAc9Y7wWCSDHV/cPhP4A/yf0sMn5q3nxCOJ35uaxWueR5Af9P
qWXdmvECJMCu4ARDv/dN0fvIH9l9VzYFmxa+QVN4s4yK7wxm71Y6dJdO1jOjfvDVmSpJvv6fi4t6
bRKpB+H2+7/uRNPHUi0OwGqIGakpGfH64UX7D9RDGeo3QOJFfJ3kV4iFr2Ey257z4CRS6mli9HOm
VMohRA6qFV5f6TpKX3ogVS7VTSwhKIIrpv2Vz2wXg/nSL60fclpPTQEd9pKf5cmhipECGg5omjD2
grIMdXGrVLDSYvwJJWfsuJdI3RJDos+4+gezuh0VSGOo+AYRqCBya9TYESx8ZQeSg8U92MvG/VZR
SfrBOab+KcfxOCqTeqcCiGcjlbu0L/Umx2FWWhlMOMVv9LsiCTfMzSv7wubNEjp39TtwjqO+CP/+
ZMf0hORKzwJSbiDOo/GVB8SqWzn+DMpXwjNTPIfvdjAdqHx3jaQsb4fzz+wwwCquyXYVfbg9NbZE
mZAwxfxb7s72XpqBJH+xijEOG06HmYU8IKFvUQzduvhkw1RMVY6C10nrH0L4XSIhuQ638kS/4LUl
Nd4ysrCGxdwNr/nnQl5ZgnKkuiBelam9P0BxqaXDWQ/e1T9XiMHInb315D+z9qHlDlfEpP7PgSF/
kUaX8bA4DnkK86XzD/V+G9GKr5MKCiOQDbA9cF9JCerXcVdpv0ybgBlL5cmH28omMiZ0CsVfx7xr
u/kRmR0+N1cml6TkNcQFsFJ4f3WluJvhpvzOIFv/XVFq1RwQ5POfk0poX+LYkxwuVzBM4zde4yBg
n+88AdlgXEvh1im2EQabhBqdg3Y3wamwu+k8rScK/gR9h1j/6YtDtOXoHZmlNxgeg+H46RsXT4AE
ozANwYeMvo7zPvzhpEDcdw1A3H7eb3siB1wbxSQX4y+K3PuCeKb8VRCSII68wG+y9MXkWsenUdZ9
4M98SwIYnPpVQQzV+Bx5vNzJPKkmXxt7tH8/C7kK0RStHVxOSuUNYRmp3ZcCN24qJsDIoVfuzwal
RrHQg9K48y5UOhO2ARO3j6ElRjqVjpyqvrJvVt64fwX9nNXh/MDihaPDhnMBy3l1eVgT2BLrAZyj
zeGXdlYk92c46Wn4xGYyeaXdZUNPPf1kaGl74fea78JV6ZPCSvf1W0wF1WoHSqeG/l//AJ+w5xdS
FAB+xQYtE2PFmSp51TQudMArwffJkJILQWaLy+tl/ZSI4ZuVA8dJxrsCL6/psunJV94ry3BE4Onc
8vtVB7VGZlSZIdI/xqR9HBrkmSKy+/RX4oL4sqWM9+Xhoopf77c167tD3YrW79pr7xe01EBslGeN
bOYoVqa9Zgunwn4TDizIbWdbm0eOZ3kzqSeeu1Vi4yayj2pM3Kw5G8PxO6U7PHzyOCM46NjN4whY
GjRSFRLAr9qbsaqZluNLVgXmkpkSXxXqN47a2uy9AS2VEOnXyWsbrcc5cJF9+7lbId2sDkSiuGDr
AGos2Z4xn6y9avYMetg6Pce/7nBvWobz99dbqhC/cPfJff9l10eEdKksQwb+OXWa8x3XN7nUfuQY
C/CBUDpnPhN8Ata3eGKHtDpcbpwAtwhyQunCR6rgNMQJV2sOE78Ie+4NiW3Nu1pArtq+K4eQMYgy
KqPGf16lec+SfUIfTRDEmx/my63ZXjE6n1GC6buzaEKckKRVUyJbd+P7nQLJEpQi2LVl9Vl+dj3M
nrNKrS6t+BKPMlcTZYw2JqJs4bs3tir2LKFMzw9K45LvDiO+J4Wm5ReBzZti1Ch3Cg7R2sZi3mv1
MgB0oRifE8+pXsy8gIgX7VVRSgGYrKF7pEGmtt0lldCTyyIqLWL2Qt633OO3G2RVRXVZzb+C0z9r
pfYWzJIUbqEHrMIsV3kkd1zLkzvB4WLNbBXBBI5dCKmnTmHA/4/LPfVrKTYQ8RB+qWsqm3cn7Gzf
1p3HOlJsxV+/3cs4Xg2z1fgCEpYnEa2JpxUpnddRFLRId8M8C3zGh25SDkKb9tOQ3yOm5Fg99FA1
UeBkQsDpUq+LwadxK5LiMMnYRtEcFvVeM1yWeeI28aUzIN5KOdYn+4Qu0b9wZSBDiuGhnLUR9Nwb
epB6lXSwIXWI/cC1Yqt8JlvYyyJ1XcP3+lMTwl11qVeXRO7qsX7VdvHjylJX3lkv9xPFV6p1HgcZ
gBIbhp1mnwJg/+bY9fRrhlxPg4skkmEdQmw6m+RkC6RuM9ClYt+QyzJsYDY3fdQZ+Fsx1Jb8tqxr
tXfpoZey0p3bX2gtiGCeRvVG0twePekKI74ADRGQ2Hbiw7se4CUjjlHT6YWTdWC5Sghs4GGtaYQN
XX0qDsC6iFnOZSBP9hLEZ9d63FwKmkUhaiGRqNZbJdjsqwJfaEi9ZUI2Cj9dLuEO/JuQXS5Z9OUl
/CF80eejzef0WfhDwaRuvHpcSX8Pe9lhYImm2tr4lDafGYT9nQY3xfZtCUD2w14LFiWJJx9NSrPF
l+zL1+KBSR7VXAdPvTFq+IYdAUVvbTS7wUNaJ4pgc7fMWt+5rIC+ySAE6biwEiM13gbemUFVqg5b
VjVFM29iuZWEwcd8UXOB93G97bWJ6VcHgc85wihagHwnUxbXucuh8vWLLvMGkxNXdFGj6P1HxDFJ
fJ/JOEhhNrUt4dwBCz4o9Hr2VB0U2pjxuRXh+O+VPMIObpnu/HeItdcONm3aKn8eupnp3NkidErP
wRr1VXGHtrJ2r+GAGcUr5AQPbDbNpazX1+oiM4H6j5UGzd6FOqwZSueF3FCe+erCqgb0WMgy8wSq
4FklwdzUCdi09Djl0EqbqLQjTg3nM0oHwhJD9TsSTytazfpqBOwECfwHHQOybBQ9CL9CZ2s9ITU1
tIB08RDM6YSs5ikUr0IsM5o4gvkmkP0ZIUeKkmrEQLk6DaJ8Fjrb+B7afheHvZtad72D9ulCQArj
KTO5vycvCQuLs5I6hR1K8QPRYwsrKMJ20U5B4RRlHdBzynxD+RhYwOLMcuyQ2QrMr3nA6mPcWZyp
CJ4TEvPoSMA/hwRgjURgpNbKYM+itFqWf8JvA01Z1wm9yzAvZ8vLXzjtGBDlju23DmZQlHoDbbiW
lz9v77AXqiyiApKcBJO/9lJyFBwO14HPDcXJYe/Jzko4zpq4h46z9GNmXo3mRJnemZB/3QkmHB97
eFseQW+i0ieiCEnHEqcMkKe3kBmFfSIr4VfCjjEgZLraldoEYgBi4xT7ZjbDsQG+mBv9XbhmUoo7
6kbQ4QNNAnuko723szcDmtxAbECQC5BcVFt7CVrWwCC9clrEFw8NDrdJHrGAtFnkBnbCbTiDDcgp
mPl17lh2aLoGBkfYEDyr98ivXYZssFajiKnmxTBJRze2M2rDn2csGuixKo1QjnsAv8dNiVkZPfN+
Sy0xDSZxAvys4Gf3e4C414hRVH4V+rzSLSeSJKRx0+gJoYF5jDe59CeyjoQFIQFcJp/xitlKezHB
IRFBRcKf67Hn20Fi0cM6jiIy1f7xJBnwmH3o6RcLwfI/LFz9D9EX1tN/uFGBD1i0JvyZSP4DB14y
RMbPuN0Gj4xEADnRE7iZDt9evAvKL0/fXebJ9X0sy19NLI5jC3kP5kt0OgnZGF6XUGsPRqkIrUKT
b8IdRTca6KAtLoyBaz72cJrhRNt/ZL0JEq8m5Rsz4xriAz1agdmBYPJn0If5AMMGIrlV/CeW0hqP
wfR7v6cU8D2u468qDTKPvkaZ20+l/U5alHuRX+/DUydRDrE8gNQa8aRlah68BfB3zqi7Xdj7/yK0
soAKxECbqy9/a1cq0lUgSYM5mwxtbnRxPg8BhmA6En5CQVogcyy1sZe9iUtaYi2FFlbq1rhYz5Tc
6wQVY00tohKazzXu82nenIem7HMMJRTJJwuIE35PcRptlfQ0s3cEVYLeP3mmhSuJyTw0jyG55dOE
9A+pakpbkNBjFc0LxbjgH5CAhXVbmQAyLUKGlEh6FyocNmF0wkJBmJsTKDpqRmi6npM4rt31BPa/
sCI5gF96EXGWt8Z2unURmNvjAKFCqkWRnBm4sIu7C26U3GbjX4x/0+qZrtV2qKonVhkA2TkxaM4U
2lgwHPPWkMBFFsG4W+lIOEiIujXtQfuzTZaeBJERCEmk0NXNi/x2XGlXmL0tEreUQPKxPncUCz/t
ii9Ox/vIABFuIt5so5U4CjamKHde7AYa5uyTsQNTC6ByXLEEhTHRQ+1KMYX5Cd7sr18TghoRcdk8
aYFDMk9JpcZCylbuNniNBjmuAs9mzyQRLo/7vYkJDzcdei36Vy19ihO4jZpBneBJjd7+dgDRlvq4
Y/iJ82NGBkr/4ZYfRdIlEtkrmQwECnfbvZBhZGGPXPBzN3WwijD1n6zJpMDoNT7C7QlvaEAY2cv6
vU98nSDUeHi6z71J9Y7ApTiL+ZGHP0L4Sr2XUQMJ1Xeum1AVIE0tQ3u18zNgDMyPlc428NOd0RMQ
zoCuVYEbO3Rn7QwEcasxpQHUC6Ly07NyOj8TqMGLeEMaXw9sIyvYyBGj54Fhs52LEaX6xK+pjMNO
TS/977wj+W8+ru2ltxy50nUzOf1Hq62nxrlYaC9sKccMPePpC9swzzLlD0PzZ0JAn+v+epTU8GNo
+N+RXtW75Qy53hK/FJ417o1kFZnQrW7N829eu2eHoDD+obiyFMl681cvrO4wTV8aNzQw9ma3YNhA
DVTD9BKu6sWKChPqnqsnjef4O4mAf+9T2rW0bCcNQCxQVntnY7uauC+c0IV6WmCBhkAYAb2dKAIC
8rg/xj9qnX7Z47jgop1xFGNwABmr9iP9MWVS1AX+jtOFJMPyJZdAG0kRCsF/xXIS/bXSy9l1RAw6
nfS6DWm1h4xMjbIGpvu5J3O748qppC574VBD2hZr4S4AJb9rojnZJfMot6CvUlsbJxEZJO0tIcDu
wzPoSBMauzv3r84UNknNzqD4M6QzpvLpxVWavel4wxTConujK0XzajWArElGDc2q6KXbhcu2zJDS
tjuN/P9E7hYMlekUvZZrCE5sn9a12Rh5SpkvyA6/htbRWPvktnqILVGhfJkx9bmhiew+07+bpWoZ
/bGRJgjw8ql+pK0mRRI8kXFpLBo6nvQgkDbZoixSC9Ci6g7MZl6tLVpEw7nYZ8D8yUDMJmObzDy2
DkxBBFpLGCWBIT90IYCASxXbBV1L5w0JsTN1E+qTEwVxWwK/trsuOpkL0nqY/BkR3R64v3OgTnmJ
NuhqsTTrmY6B5HKjga6VtNqBIKqf8A5y7ct11/dVp/zNd2j4pcJ2S0PGPdkAbsIV8rtnBKl/MzPd
AN1KUW1nrmlrBp1mDHXUyzoHRVFziCvuKqnpSPBZ98Dvy8JyPzAt646PTx4Y/tdGfBknmanw1vVm
SaXRmeMu8B8iUFzPUNk5BNAOZabgoaotwvRuVV369MlFlFORdsIEWn78HsqJDDsQH2RuhEKnefky
z2mrOgzHJBAIRYS5kAKXM1OYSJb/hhYuJ6WAIAknrDXmT0B9XNnvsiIVaTjmp8qaCgYdQ6zmyCRz
l23GicicEjACvmfeLf4R+1OQbE39uaf6OQmOfTjNTk/2O82EjVZ6S1B9fhc9F/L9lWNbCoR+qcJW
XWcZJXEiGdG8wY73tSlIzqRg3QQUhdKxN/yC3FGvrijZefVLlDlhcEUGN3dSIuQglRa1PKsfEnON
WjGhw2YxzqIZyux8z0x0HT5sr1O8WdPpAGrcXXoAfyrCbrgh95pMaaaUDXKsQNYnpy2ZhjAq6eCB
v1CbIYkws5giA/Tyr68i445QySVX9c03RAJo1nh0GuBsOyoYwaxKXIHYcAaLvAkkOGlFjsqQkGMe
jT5a52UI7H9NC5IQI7RJbZ/h9lKrUAwC9GaIIiNGCd/yZNUh33RIsdlr9la2ApufgV64ygCS0Ika
M+ujpHKkxALGr5v4BivuoPza7E32VYirF8t7I9KXSdj2Q9oi3MsFZgb9uXFte4tZ5ZnSBHVyO/Ti
UGQsPriTU3DaoJxdOck/rmyxcXFrs/Dky7d0MTIWqyVFGynZOeT7ULyO7GuxOxJX0UzHp9dOEfpd
5o7ZnTjwCHDM8GV6QHbUD/8y03JutXppHXUo/JaDoW9142gOCE6fqg7rlw28KqPtDVONlh91ZNo9
LXKfSonbGY1B94ivYcfrV5WRlLRg1gaIBPdhomqOpzX6f/Gxnsx5qpueLvIyD26U1GaVcc9JIuxp
gMvFvd5vUetaeaODWDBajTwQXdRLRUm8Kjv7KPeDvOLetLpCn2bTXZdxTMUKw+2gDnsKwvmwZFPh
Ng185UFwFAuV2oby5RVduujcDJT3HflqfR1opqKseB7Zte0LgC6yxoyhzJaJRcbrRT5fWPq1LnFB
9tbAjCuW4IPciDc64h1P4fWL6DHMKGO8ThD5VOBoAy5VVhCg9n1ga24Ltp3YNG9hs8F33qNGO8jf
LRbZbcthUEe3QnhvqSyJ/4o+P0KuApupihi4wCeel4zHLllYATtYdlqo5M4AEhBNHHvzYIb5OjsN
X1E/JAzVuwFXzOdJtV8W6MJSnZJNlnC/kkJ3kzL66djQOJw3eYUCGqnAR6Mtdpfqzncj8jiRoqWf
hbo6p74EV4e4NKOxLyGb13lM6BXwWDWTcdI8R5bqlSAUMl6IVP7bSkrVhYtIRJxoHWTi0CmWmA0P
TEQvH17EAoPBn/ErJqRgT1DxmnpsadVB3I6IyWeFoJdGlRX6D6u2nmCrf0rcygeS+N1Z9HsvHrxF
8G322+ETh/7UDOr5Im1m7Pmnmu7sN2lhzFWc3GlVPN+iGTHmRiXUY5R3JnkDfi9W/ssnaMCE3LEo
7+KlpT5oy46iU3Mh/0hO3GA0YeY1507GUrHdGln64DVnxshPfE5fBupThzubtBC6K/LzYV0F0hfF
1p0JShqQYwWESK5xE40wOmbUiufLrha8XR08TdeCCCAuBYrMTZdu6HfvgeL+GI7UHipprfWd3WxU
ltIRT8N8v6cxX3k76jfzjby+9+gILVsRor4tz2/q8CnOIFsGI2L6HiHMt2oC5nE5IamTuBBOzrEe
5Pbd7zUd7Fq0VAsEuWJ5rE+ocHvUMTwBj+OjmzzJM2dHwhOyRCYydMMJ9tcSbYz0mJBQDp/lpzSj
xZwGOLUhsU5Adx8VeIzcFKUPqhRlTJh84WcbZFervYMJ2ufd6cGxhdQnKiT8XVT1AT3dp9YRDy2J
v37ysvOlvBYwNzCBcqtcFIgC7LfYLG/KrN3EjgUvZCYVUaRYojmzuub7cZRi2Du3PFTI2mAYJ+WR
VwCe86yMubCYD6kAaFD3+0MW8hFMct1L1qfayMYBU+BvpcNpNDId5jpg2fFSOuRIEF8KqOxqo8eV
Gee0CseMZLXQAYzhU+yIWVyI4uGVt0he+jERqZGb1bjJLhHyw+qZUh2eJyeHtg7wwZ/D7ZqIzu5T
A2h8RFCDb0/kVU9SrVA81EImaK2E3d4t+4rTy+BFCkYeJ68o203T9bGasIFDV4YXdh8ZLFD7Cl8s
g29nlH1CEYXpRbG6VMprb9G0nRROJM1ClI2Z5c0/2gbuTdgVbN0YdV8Cm7jTiIhRRwwUZsPxhZZt
uEkDmTo3504xvbHuAfIUOsrmqdqghYG0gr/S6EZEwcecqsOAfbN9KpGv5Y9GqLmtqmsODsdaxj3R
8D88Y8HuaKKTDstnN4VcjUomiGYuWId6xTbfQHy5AOsX2hDIHrN1YWgNN2nyCV6vF9DD9FfvwvmJ
D/+6kkjilKK87o9aLtBa2Q4vfm7A5oLpfijc9G24cpNozy8GKPx7bmw7GJgIfHmjpGSiohPIe031
AQ99LAvHi9LtzCM8p8sRHNMzcIEnKoDqn7sgE+K+p2ETq/WPwCo+7laKMKnql5VntIiLQZ/j1GZb
a+6y5hMlot8+qtGRyTd37sUzO3z7WfpBY9XS3O4I2i05q04zegqOhgA3mWv7iCBYOBowzl60SqtW
A+YSl2fWnI/pKequJl4UhnedIr3cmv/n1qAXp7oMOcayjYAOHc994KiZkYzhdZ9PTSrbqyhXPMCo
2aSi9jebEOidbk9Bf47hoAzdFjziABpJuzgU6nhVR/mgsi9luGNwpuxt//He+BOND585Erhx7SyU
Vrf5JjOf89quV2+9npaJcE3tFmwjX2AqIjBvxcyPQDQotRi72UaMerfyxgYalGe0pi5ZUNGkT+Gg
w+sji5GKOQl3bXhB1j98E2bba6BfJeEp53+rGbjS7dmP/yNWrn6ph61ZGSBQdBQ+HctrgdDaFJAp
JbhHu3Dlr7guD2PvAtvfwBGImY/4xDhyyn7sy7uHtZ+bFYa02YhnoLEI7F3Km2+lJ7AEbJ2EJpaB
6YamU9IJK93SmCmBSbgEx8kuLn/2jLh0AeQAybaKmGwF2x44yIib1aabZ5B6Qxi4uWWyrPxjZq1h
9QtWHgEv8hHrateSJY0yqY9/TBKLNJjbfeyMilY7nlBno74XrAIX0SGltU3EaX5Y+CJ0mVLn4bhI
7DKSDXxKDXwi8oTVY1yqJNBIUFt6ID5Mk3D9HoeVhbV0QlO6EgJrqOCuGiUJgnd4xWykFVQTf3+x
z5EJEMYIKOtbhvPrJbatzSpCMLWGLmAkshmoh8w+Ba9cO93AGK0MRDHoFtp9p+yh9yi3Kg9KgGEM
BnwzVWNWP2Wx0tE7+UznvhNuH8ChXn6LDLbdVTH9NHA7fkpy+DyB40aOnRqvxuGmfN1SxF81fLox
/ZejHEQ3ZxIR9jBUQz442Ek1OJmHn02sxJl899/vn6S8LGzS74DrcbXwxIKxixcr2FnoCxs88x0q
D8Ph069iuUI0t9Neo23Dq4Kqb5cPDvjWoakt8rD6ILSl8ENSDQ9GjqZbnQtwGAQuzpclQgzmHmJM
HCSPWxa7SEmGIMCEmiytFtRlzcsBWmVuBobeOjm1EYcLjRxdShlSJekx/SKxkB7rrDW9oh6eX9X5
x9qKl0YzeeSK4o041OZfUX9Q4xOuhq5+7tPYO7uzYnNaxdtMnVv3ogecalGGsKvIjNnsCD+TzcyG
30snC8bm87d6qoPhRh/ccsl0rIPkJFr0ixPcwP75bhMgTdxrsexVP9US3y9APlTpSCBPjlt+fcfV
fMLD80zGGd/smmIyNvg5OWgmgSq+DiRd2mD+Ojbw5u3livxyoQvc5BR+PUVq57fc5fwtcEFfV1FW
nMvS2lWn0thpJwb+QeIPFYVFtftcGQcfqirPPbpT0H6v6Hz9YUjL0H8LW0+AWm6m4z+s70DYpASa
fSlnNXh2G1s1rrOCE+20aTl6kFhEHFCJ3sHo2ach0ZCvAzR5K3Wp33U4MTbIznFinYshRf5XDj81
KjbTPAGT9IP2+DKY+ePHBhBPrfVFw0UqqzofYmw5hsfDDJmc+4Mj2RohvpMOtatjvPTLLYSgxaXB
y12+7hi2MpbAa7hMZstKsqh9FDMuMT1MFwbm8X9qCte/410n3jTXGETrkG7wM8jOnDc9wQgJqrMp
JVC8UP3ekbRhDftW9L4xfwbycZTzWPrCwKTr1udBnQRgBtZMhJy9BkOH1CV+yYzB/mLuwmZylkdh
nGZKRFyrYJX+liP5KG/FT87yTSQae7wjoNm2bXxKhSlrfNQ+Ovo6GezOuFA80ubQ0NOJ9DJNAHtH
qNAqlMBFSTGoN5elPMxvCo1atRDgjrjJGIHEoaeizf5opXPHJFqHicnQf98w+QnnFPVilGglvqQs
48PfmY4QZlp+Rq1YZSsj22YGfZywmOE/ETyk+a4Wm0Kte4pQ1vIqgJN9dO4OqlBRKbqUkQkrdDqk
FCVehKSZobDL67HGVWX7mtrQzL9qkqZrKq+x82Qb+w6qZrR9HR1EuAZ18SoY25vFoC1iv6/7xbaL
69956LbsOwgtCFJ3Z2WSW66QZEpwr6Z5V59SH3YPSuyZ5yrZEhspqZ8acIwIDZZ/HH9tvUYUgutl
8vOfVqp3RxGK4sMMdOX/vgsDyWzRbsvaxyNWr3da6o/0slY4JHDqWPgFNXJGg5KymXA9+x/ZYM1K
+qULogviUR0y1air4aV2W3RjLQ5/6sBPW8XsBfHRQF0YKSKRRIUDwXC/YC0g/PaTTxFKnWqb+Wmp
GxmZJmBzk5BSEvm5RNHjXuKaijhJQdyKVAW3Nzrg8fjKjdkDXePNtJhqU53bt0htTQ7zXxnkEL+r
fg9wxJ9vLqoc3mNrkvigmoFml/DsG4kKTMF1fV62tIqm/NCNk4DEw0+DIDlWbcpsFKkxj6BQnH7s
dJnVQNeFLn/2hmY1YNOlBn4QssLLJTFJoDhwXfWBOif5NicX82LzljELQP0J8QYiuh1cWe/tZON7
r8eGBuh+8uQvWBTYYQaEHTxM1yBMWDUYL+i3XP4qHB6KAmO9BywIf9RGvS3vxwEK4ilePKeSCAfc
W3pfqUlt55ilgZwFvM+dFuRMp3dwtwDKluQtdzrgaE9uT0d2KaZQaosenVPI7y0hinWvCAQ9MpMs
a7hUsRH6PTxarfwtlHfIp8hIra4lEjgk5/ybrm60ooTyZAFq1s+duIENDmnzgIkb9a9KY9KLKD7t
FMHv3KQ8cC0IjxNKkowVb87w0gZZTBBLF3O1JvUbM+I1Lm/N/4i81hbq5sT2Z7vtN2iMuaGjPVKZ
Nf5NOK/rzge+UMdLxSUSJqY2aDTKNQTnpx7fuOXg1yFKfh1MKhygHLPq5BcRGzXpaUCyufweeVkp
OjB4KtfMQdHu6mx1tZ/416GF9Nwp2KYOUoP4GaluQAL2VZLDZYV8ASwva8gqolE0UoQy79HUWI0w
yqPo/VQOVdmeoqOZ3TIPCQMV3KnellueDMwBXedj0aGE7obcihSqRfodDF9WoD5Z02JvFhMluxRg
xJppP2DncAmIMu0J0QjzTt9GrZYP4J1OBF/2tDXNck35uHhHus5mOxcxKKfEWe8vdh8++8NdVSRU
Lbp5fQ5ORjQAktFZzbevei6y3e0892+jcwbYF1i+Pit7SGTPhQc4NI1bpP1LWMC2oIezdSmXsxkD
0/LPetHEVXrZOcLPSfFMg1WITl93YS19ThC5I3FN8cJ0N276mMjFPbr5Fsj7FLo8U27BklTK/QnS
JY8LPekYfwkQMO1sGgaNqjKRewVzy6nm/xGg6lw9UTJUfc40BgU9wJoFyGlCc3zTOokTfn6mQdIU
KN6i8CQreBaZGC4nRQN7wq7zVro2zaQysvUWNtrZUHtJqg1uyLRoDif80Vsf933kgNgW42ARjw8g
Q3mcMy26V6Dd0IDPpJSCIVfRJvYzAbwVu0ruZKnb7t/OtXW98YRdQE6aD+GgioJEbJ24aQjH9bRv
MU2MmQt/Fetj7hySeVpC3APNmaVwBt1Nm2SPEz3m9tvSWL7xaN4gj5vIYQ19tHP7PK8sbCMZg3Zv
DcM3Pfppc7fs1lxp6d/YR3a8lYfCd1P0igh7gCUvg0hFTou5lzrDgTYzizxarezwvl2lgupLqLsO
ZniPdsBeIsY1nvVCCRQk+aZGL6EUunoUJp/mAoQ+Cc0jf9frZVXMaST7B6Hwr0iaaqT1pczBdxBg
y8SwBWaB66LPRgGR1tL1Z5F0R+jIcSDZ3FbjxMNgweOZTz9iGgK/pIxlB94WNtqJDbv6xUpHYFg/
td2/I3kuEk6qb8DzNpcz646YoXhSr11zZ2FjrWjPa2PNdrgnFWUHPqjKgzlEyha5+ux5Qg8K3cbi
9ImKHT0d4TXCcPUGJMoA5TrHvEVW4qpBzfNglMNoNZRc78KnrF4bZMI5Wl80kNRJAv0Zmiov1CP3
moAYkia9zb7AhcAZ1AUTF5FCX9RfuZcBdbJngUXT71IuJzTpXT9KfHFnoWHr/YK8kaLp3w3s4O9+
xi+NKmT7ofB8Dnltz6xdpihAHtbw5HkyF7YMgz09/zDPrE32CUdFmgMS4PGAxW1SOib0l0beH61n
l1oXksthYjPoodfCsp8WOKnjk4NjXggShXOv/CsgfOE9Pi7Pl/DZJGlJtBtM11hIM3bd641U7Inp
bVO0lkn8HOyX2ByWsP41wu9Jre8lCbjec0/yKU7WxUBd8eYlMAIQDeifkXACzeCceiuDs122Smle
OVSno6c8EsySm+g4YSsBne+p9LJxyKx6AjjX77FMGMz8HSpE7PL6oV2P7a/0v7su/KFv7mxHlkkq
tq1i8gK/F6iB5TBdfx7HO81BoINgmH06FPOACq0kdnWVAHH6b+3RIz7cH8oOnu+iHJSK0d20ma/R
He3+UMxYF+NJd8aPyLxXz+hBy4vXDyup6hI+PxitviPhqXGexlScTGeI0pUhfZU1jhPfQT1C6mDu
+M+EvgXQGZcmV/OntimiZNPUj4NBXAUMV7VZfxAdZMp8t/xWxy7XYsenfqINgExcc4anCAOJkzGm
DbDuw7VFIM7bk7Go1WuUKWj430ulWr9WnN/fDRFi1AJIL2HTQDYSKrpgVw92gF0AUk7Xph8PaQGG
ASusrGgAJvj0ax0kXYffoO+rgZlYYi/2U24/Ta+6fV6jwqVPmzjVTi1KnVqqrhKHJ9uXh6RRilm7
jAbN+BwpXVIjolish0aYYfl8jNZ71VVNt7QQfN/gDwEdIZpxeHjpKGQoKvUQupY2d6wVpXS4B4vX
i7D4uoPjD6qT+viwQUYqHghxM6cOzhLfauzIOIs/P62YP7ziaN3+HRksrREzPZ6pKfD5+ymN4C8n
boGA5KnPV0QJUutMV9FTHcnjZMnDcjsWWnkYm9IgpwC1KHcWxIcUMze4FqPNPLFSeTd4vqmEQELJ
cfY4sAbZCdvykG2sQMd5wrg7F/SinPp3CKiKSmhAkUm1MR0z8Ka/mQGd/Av+vanRcVi8XGRZBsiB
sdy+nO3W6aqU+7USESKYcLVIL2du0xzxZrVbDJ1fzLNQ10idJNvN9CcnGCmYzR572JQiknGLxr5n
3XoRb1vgArzw1fbQd1XyjsRBDE2QGcYBbgMBQbTpnsowvDqFD54rGFHuvbHJ30D6F5fJgobl2+Uq
Ymi5pKI6vXBTc/2T8LrPyNv28olEo/WRySn8bzy7pqTMpIomYuUsGQxCQZ1lSKPvOVZpUzQOUrG5
lkXAeV+ujDaRSxd2EswWWeiZLPNiIfmjl07HeJQHVYC7XjkV0N7UnH6RffDRTzdulIvCfrkPzPYq
8FC9Mi3QF6qGC8tNSF/rX/d1rdTrrDzUs8wKT8SRAouaeSTU0vwI6i7lEWmVcU7ilnilm0n+ehqs
SV+Aw/ZN7hPccy5W4aGO9bZ3aurshDoY1B0Ogtm5QCp/wrO1cjqhemDxrAq+TspeFz2Xp0ytBI2e
O1e3IuQ35NYpVNMTsuhipz2J+HWxJPdD/dQCTfIvgzzBjNPOQZMidQGIOYckXufogB85zBsYqniV
cHcIJaTZCw3s7JTYRlIOQ0UwDAZihPNn0uOfuqEJmiDh2fMelIWnYwvfZbwOgb5y+pVXtldLNTVb
ZHhtXlQfq1ycstQubkQy+Evta5PWuq1SCVBstBzQ5mlHxlSw1GfIp74c+ZDgHsNmHRmNmI25VTlu
ytgBgfponppFjeqzgVK04v6EQ80re9Iz0cnunVdaaa1IMFlfx4dUs7pb3wgCQR1qKIHLbSpo+lhu
HOgwih1yuQ4Ma0cjv2X2NtLPVETipcBn205d9TSTcaiWrzsg1DTvp1Zoho+SPtcQ9zffjTG/dAaU
lBB2BD+ecoTg2UrgqjEw0fp+c87kO7pXW+5yDUyvF9Qy9yo+X+Yoc9nNspHJ/XKM9Ht36Ogv3NSs
by952UEmwNrR9i5Hbv4jEsotjGB3OHN+ToDpyEYtQ1koiI6pGWXoBIxPY5OefrclQVsfQR8eGxqG
NXohwIqmUR1NwYeMm3YzPsvDIcRd0lNbWbxlT5kAAPfW5vIEeQS1wOTYaeKDPoh5ECfkwYFniKa6
865vLijQqZG3mzWAjRuVLI5wJ72NWYHt7fWG13da7wou6Ku+7v66YfFkw+FGYnW/ixJkCafkBl9W
59QvDsRJ/RDNBoacnbh7RjLEtEATzer3MKh5llLqdN//iwpMiTf6gTlNGldPx2LJO+uKWR6HpB/u
5ypoeJ4lNgT1MwkDdbc6kDjt/3ZDxwjWWjWFWsGnsM0In/XJmA7VzaHacjK+QHB2wK9QGRLVsdF4
ZGVCgg7LcSzOc1wddfrsqAhW7XQReReNjJnOY4//QMcJpKTsXuhImDpgjjuTeZMxZICs2gpwCD9i
KaxT8je+kyddJyJgduSsrtvXgUjb/7WRxZOsED8Y40dx959mItlmOc4aLoYq3ozbsqocLkVI+Jzp
gDrU2nleEo7xBVUm/V02+sEzov5jXJ1VtbWPdzyqi31T2kheBIeOVNObyBMF+qPV1jKLYMxSpbCw
CKS678xGFZ3Ylu8VlLhfBwUeCC11dJwadLC5X2GEAK9ULoLyOjtGGlVq9F0UgBn/y7XfoFEQXqK8
bl2Bz2giTv/eFNj753uo1UPK0KNAwxMuAMUWFIpghB4BYEqDXaFCUpPPwFRhp7i4GFKHvqPaXtCR
0BhA/CG0Q2qgtsUlN7pg4bQEWilLqBmrBMOhxH+XWUU01FC0b6sqyELP6qs7E/I7LHBRi9jpxSFd
pgnIWfwNcBHDr7nGtEpbBWW1/ZAMoc3z4gl05HmodA7AtzxpWZfNObMvlREPXNKQqntCGpBj7Leo
X2kS+8wjIZK9kg2b8axeod3zjbqviXUMk2e/NIpLSTSJ+O5cnR4Fi+UoL7I3VkfpvHrjxFq6ifu5
yFxPInQKsXoSzO5JXJRXVYhLZsy0PkVqnoh1hgLnUGwnykqDupYbd7BaxmPYSbYZwWqsB2b41ybV
LcaGWOGJGXuOe3u3kNh8lAEehu3WiHg37UQfVJetfd4vwTYDQMZ5avR1IcDHW8ord2FMgLVSWQIr
Sk20sg5l+MaFdB0LTGbC2PON4RPtKbXwXYzLdM6+xwsB4A+aa/mgCV1ksyHbGbTEDtuEqLz3Ur3h
eqJhUiYrtL/QzyK+MNgCzuajkfMA7YRuxDmmAOnRNREbssdmhPCLjFe8g77l6tRmyaaDlQAHsOQ3
wVFCmb7QQVe2MmgWKhHqhVkTkhisx5HkNWa9/6nLQt1VwAeYTUO3+W2ZWXkAup4CbeSuMUcGnxvJ
HWftVjNV5pGdGxyqdYVULOEYnXtLj6YUx1pY0Dk5DSFK4TzOshFQ3XicdCZB9x94ZwjeZFFFhkqJ
Bt0trgl/cxD9xY/GA1TCxylGqg46QGnsx1DuEy3nahqekEdfKaxrjX5EtAxc5HqkXfyHAdeom5zk
iMWlEBHy0bzVWHYFDZK03wPzXRvy/LLdNXtR4d/DBlO7ON0tvQST008GLJI9sqZDjX0d/zchSO0P
/wGiRvLj37EH3ii4NB7B6Cme606TAG+65KPgZ2EUgsqm0MEjMH65BdXq67Kbz1rQHpsT5eHvUm2y
mctNUlR7MxN6FUVdf6BJrUkYSQQ3BFkZoU8hZDKmKEFNtxr5YDKSH9Ilv4H0FeD9HjHKFKwdmY7F
TYdfnKig454+al8lYSbGijpBAj9TMm6JkZExIJukVOJYyr38InaZuO+3yEUtEPreWTRaHyeuKePI
KpSsKZJn/fGBUgU+JC0mUP6VjJIvmKcqbmf5b6iXbGGt6ZmQ/3hIfEimUaReDkblqfyvvW1z2KIT
ip82RtYCu6Ppccy1h3C/Q0bDn/Lx211xdjTWP12l/nWXceTVX4PTsQRsgoY6vW2kqWL/DMTyqzGh
Tnff+azcjmsSI/k2ESlM2B+Vfk1mSJMNRW6JOge8g2kGIHKbz/5xFZRHCyZOid8sxpXBPyjwOj+S
0GKOgWoqilFp+K10TIA/gR5y+Lu41WJF0RcHvHEM4Q7JuWnQK02gWbv25Ba2ZIiwYWiWbU63C9sh
Nj9pK91drUMwr0FF/tcgnZ/9/p5kFixh1Ochtlr2/9kPHsn6S03JyAF18XEl27ygA4QQmDO6y632
+hdokPKePbFy5rq3dSeYzoACH0RXzHqCfbDBCJfM+rPIbWACKAnx84o3Lentt1P2WnoL3pw30Nho
Q5DAyp4FmkyfMOjxuohxzoObGTwXt0bytEy7lD8bBm4MUk+arE7o8Qe046z46SIRg1nwriXqSaxM
3sCiDyOLMGoBYlwQ/o6ACSP1YFu4Ndj9E6kA+7rNQh2sdI8lCkv2zVcpIOs2IXo0kofPhKERdH9h
1JospA3jdC6vfy8IfC+VxK37hX5vMLuXYF7ECvyWtYyywgZI2NxkZcKz8AQ0LX5KRU4emJZlaEFo
N0+Hn9GZNRln0iVlTcLiMlTYCnm97YwnzUzZjLDk6+CY2RszhwgrMG3ZfMx4lCKMS/T7584vOz9P
i/xrX13k1RnQ5hx7V4gSiYgari+dc98opcWJlZMnP/t7h6QxbyFjbf7HL5CWvV9xXYx2UmUq/MpN
PHNmWiz91erN+XSjCe11ET7ACpesaSpDmbqntAmjbjVn6SPPGpue/E5NpNtMK3SDytNaf9WmqCnH
jC2WjUMd/0WMU4eiYKmQdGfvjU6G5H8YCIdgjVodf9Y8ZryvlpP2yPQebI6BmCov8SQTr+x2ER04
bNVG1KGB103DH9Ma8ydgVp6wNRr5cq1QKKjfRZnOG5lcQtaN5GohDL5C24T8y0/hqFf5jNJECIDP
3X8evGQolWdou3DLNmfle/BT0JFgFSUZLoxmwz9kl+2RXhBMH/5VXJwmJ+gMl40bMKTcmo9hKhdy
sNuE8smH8ZRc6bj9nn5aq3NJEaxwWOyT+HB5SA7TTkakgwsrlk5M/5LrfZRq0ZUU0JD4+bhqRPBs
B3buN/42LTktqiH4Z7TBjuBWlLYYQzWx9kRLVLFUuDiw+fB6lKbZ+YD2uExH3uPrFI3ZRc9jDipa
MGiMVZZVYCT+xd3OFMpxbXlWt9nyVS0bGIJ6ShjpVG0w9QcULz5ttoTimohtey+PbOq5frW/YkIA
sgSDd5NpKKOIu2gWTOwSRX8OfC2PXeqyg5ZUFSeiENIuZtYv7tSTXNxx4oogt3cyXefkTxSlO5x2
mHcoHTQihihwAVDFt6nWTI4ckJlgf66vfoHFrXdaw25/Yu80wUFTpvPNa0a6J84mEnbef9KM1mMM
ZI1cc+blMvhMvmkP7lkEgH8LCFchE5HCh+Gph10UcH6/Lrh56VGzCZS/8lMLktTZDwGTOKPMLuNw
zFoVuQeAc6kFUFYhkqnQs2kshXUUvQVCZl64gR/s2xUZIMy3eqUzJDY2z9lgi/uu8UMMw7Uz+TX+
IHciP7eF0trrIDhxZYpKGPN8DAFQSwfQHlnSaq167msAUdeddqeLtE0GTG96GQ2Rg/2iA7WnH4Xl
+W/zJ7+Gu6PhBQxAZ8tTO5XO+knMVncYtHZGbrIAuji/oQGh3+Hv0e1OuCuzL5aiKJMdZ/mANt3m
OGiVhSUPd0Msk9+KQD4gT3jrtWNxLoRVG/mcfoOmJZQ3DXSt3uEshjVJwcsNyvItGH8k88sQW8V1
fGrUJd81UortGMkNM6fcmLKoux/06NX6f6NZYsllmAtPZwuHgvEwCDlOeqwKzm0rckyDX9AlLVHw
/xTbda6Z+H0WDLGTkmCdlGqwSUovUvOBQJ0R/BCsn+zX8QMeafX1Qy7ZQ9DqmCrcZBQWAk/C0oDZ
XsYkPZQ/2GkexobkOEtsX5c/OgGvpL/f/7/ubVpAwJoj4CDSjKOl91bIsySM8P4hTP7CeqRSaRoW
9U7fgRJ/XXhgz0s7mvu7GM2mSIfLkvNslGKX4PG6np6UEh9OIBg07Gjqw5MtLBB5Jni91g2yVqKF
DhMqeMVZLCA69VxAx+h32DWrJwgv9QqOV2F1CQQWKfxcRD+9wgWYMVjct/uVd507c9eediHOeJIV
f9jgXHGqhj45Q5WptqnOR5FOGgdCaJNo+3zfsTR0A6iwc7Ybws0F/NYoBKpDWzLTPuzceAJNHOpg
QUE2IPMHUTBu1ITvVC4Gd6VDVJbBUHxg8QtPYZOEqyFW2xr7j6j31dMlJqnGadw8pdASTe+gkEuU
jaXReH+FcjqchLfTFyQV7RWPbNij2CS0lxU2VjOPsSWnzFhzsaOapEdaa2bdRWXZ2JR5ggTBcCIV
kkdTdkmfAu9VIm4xcZNHvvODRaHGDF1x7e8viPH3+yASGaGboQ7EsNQzxiwIdUq/wKaQ4Pg8NyfA
Nqcavjv3skZHpK3hXL8ZLV8S+wdsPjlzNEN+Cwie0J90U3/o62hA8+asJkP5Y7t+tOT5bPiNfmMK
sE2rAUZrONq3Mbj5NRq6tinFaT2sTz4ePB8ZqybTYXJ9a0zf/QvKMO2XoCfLTzIH3VbFo7IF1FpA
xUslVUxwiQywrlzNAKzyz1YFsOOtHA40OnK4QNdkg4/tjvxZFNG7B18i8FvgeT2u6OnVQfBgl+bL
CCCOFtK2SEAVAvPESsAn/Z32cBypKru19ZcUl5UfBDr6iaq+s6UfES+dbFMNqzfZz0ZEvbDl0Dv7
o66qy8FI0oyHPTrF348NPsng+xTon6Q/jUNDo/CstAyyypBMeOq/5iqv5ligBmtlGJ6uxQgl7rS4
u9By57dsmkmXfjxuMDzpZSgKCOYEMjcUje1iuqFbw1W93Tn38RiVdXi6MCeLP5QgYhoDUUz+XvQq
gzEpUsEZOn9HW3Pr69dxBM85Q3t2rgpPlQ2tYXQ/umeKUizqV7vNdc/72R/PC5qIbtiYxb4O/ntz
BMUUSKgKH3hwgjXsDd8f1qkyHUDm1md9ko4UPG13mFZpHXCCqAtAgqnRhAyjkiuFji1bq7ZShTqX
qVQcjHKfoSJUsqoDoU41tEJgIuDx0jgkd9zgTZ8C1snyaPSsp9f1dwu1nRJgxu260DC5r4jy3Pw3
e1qzprYLSHppLOzc9cXE1FcCtA3rbayVnmArMqOdzDX2pIne9YwCndwgfcq0BdnV0tplzny0jh4F
yRUB7INJ+4/J2Ue5HXsdE3GEl8rAWb6Zwn+Mxy0qjMVE/GcX9xC9X7Bmv7Lfg+hx0FrpExNgaV/j
O1Sv0Rk779/PcNawPtw7qOOZXKyz0f/umcZnX6O586QYIkTiDZWTGFRanj+4Wghwq8p6ddRrJ7oJ
gzKLBICmc7pw2EDAohw68XN6lveWneURFefRFOQZlja5wT6Ku/exo9Sk9TcccMlsRheHS6P+xKA+
r4E7mKwnrKQ8OQytqoG3YExv0ARUN6LZLuVAA+d56wP7fJPSW55TJh0Rgez8Lp2cCC5Bwue+BtBz
pDF4L7ycc/wMDOH7AVqifpgxuNe9hp6TbyTDZlXcKod9ghKdt8jhnQZQgf6Upomx5f3fWuGJWDvn
Dlv2AFHqjQazuZWi/uD85NLwbpAkXgUVE35vTGujKIQ24dOtg8ty5icF7mWZAZCSh9hwArlRUKZa
DIJ2CZDOJV/WJrab06xro1gEbdGiQttcmJtnib1jceXoqxKBt+quPcT0z89qQtiS74owOK+4+zA6
sbzluFMgRaSnZDj6GQZ8FEUp4lBxK399P6CKXHI4lBXO2BRjbYsDyVlo/odQnzmrvhEHQNZNc+FR
pfeg4IaADXdPn7Qbb++f9HWfa7qTfAnz3xBZ+jpOXGIrH0kn44F8CYJIeHXJFBFImKAyCz8IgqLG
jJMj1+1eE7UVernao9C4hRcdnDkuVmg9iRRrFdawGMLfIjF/NDU9OHc8I1CQBPqFfR976br7TX12
1IvXEPLyCZiHkW1hsEu1UZf65gmNzxZwSjW45RqsyQzWKKyyIoAtyx2he8r+ypVwBqkoHh2aYeMH
Zt/teJqGSF5cKV+1gwV5cjzUbAl+f9Kt10F56vuarYvP8/BLmGLnrscdN8AftvzrqFt3jMCaxWrh
TqPmFohygjwBbZQYhO4L7naUu8MJPSXubrI/KuSxyhSpc9sXAHXEc/m0pc7egrl+Q2clHUrVyKAb
c2vrxSf5944Wm5PLL8hm7LeILjbIE2daQHQT6gWTKX6KkZCF0QSYkoQxDRhYFbc3bROxLb4w5Ezx
81ohFZryT20+7FFC46k+CUILEmA0WLfWRc4UdVRh/9jgbgp59EUa2WDDm8ZtD3mXlKd3omvbOHaL
WYNwuVhc1kq4lnf+NVPaZmPRh1Kpp6s3CTzmJUnDkZ94JtvgOJH2OzWt454AXymdeA+UrGsr7YZE
9D6rsIFJPH6VQXtiUnA/HW/5WuRwm+YU9u3MA3Wstmzd77ickrL2tvRNwDqfwMUImQ9DDTf6zfuO
nPRaHH+gF6L0DG5pzmN89wNOCR+Oh9UKzR/1iUaKTwfIBxS3PSBdZs5YCDKTtWIFleMg0m1o7Gz0
8vHB5bX3PXQvq8lPXwx+ZsqHDGn6XOqVL/9o6OsK04UvWAmqMt1x8JS+0+IOMJ5OZL7EJ6d/JyJb
LRjNDd1XgxSOu1q2Fsil6yA3DFL6VKEe3LG8H6gMjOPH1KlMfc/U1XT7eMKu5y1ep8As34TKHWhr
62sUDm0ASog2s1ruuN8xpZZJRVQkUtx1Da1ce+uxxUGc0XW4WV3YGXB5DhsDxh+xMb+19IYfc+e6
9n8AgeEQUjsG1ETf6dOAknh1/CIIsJrtjIdPDv+psrLxsv8nQSBBuwmOOjqm6gLQMk66EMQ13FM8
jckQsac7v5LD8WgYvHiiX7OXsBR6ZPjDzQhUaDsbOcbBXnrnFpV2/pN+MwT9h2S6ryeqVylu5l06
u88y/HsmZe34DRA06Zu79wgYQPER9Ua9XVJAsR8Effam+pQJNT3OqeEYxmCFyGPNw0At1gw6R77w
cxJ085kM0h8dUKWt2wNFfVbRDJfJ3ekZRQpJkJ+IOtziXsKsCX8rJ7NURnfD5Ku9F8HFIAmhE5cm
JYcQoy1XgHVW2jl0SXcSjYskS1eOwguIEKohZnpkPf88bL4ULFktWsm2Ioqk7wNWyB3PNl4df5hz
fKLcbie+O0OgbiXDbBlbwBnUz5gZgrji537GZD56D7dbLZasFFSXLSXVBwG0jKtogw7RVWTVezwI
GcTFJFAVYTaDhvZO1bw5UPWTrAo4EDYgnUaqmD4lWD4XfWUlT+5O1cAIneHGk9IZE55Bc24RVRew
+WMmNAGHwl6f/I+l+WdZmK0Q3DDIslCOfL+ENfVBfkiqoNfkq+Xe/4Ge5ubYPNkxu0hz3wTuFAeU
OxaIZZe3GXnO/T+EKNXLYLM5PtmDgIZI6Vj3k92sQVhCQcbm/8R5/eozN0mN6Kf5hm2DNw9+/DmE
KgRc3+GcphUmj2jM7j32Vz4w+Eb4JXk4JH5ztCVD/6PbVwh8WdXkUueVvDQSspKlGo6ZIGkZYK+X
3ww1Gn3hlQkat130SHU+c/wYE3cbm4ZZhM2U5guzRQhkvAmQlsFUmVOWNyROg2ymObZhS639KiAx
M8Q4kKRAHnQjwzYRFtdxdK5Gmf1z40jJhalr4e6ouhWYE2aa2EjQJeYRSjwfPK8BPtoeFFrK+YaS
N5EiFZOq1GlpWKPj6cg3KwvwCG/MTAkXREXkRAX7Q0SOEbvuFLn/51zww6b5eXKzlVEZcIeCoKjC
b2Bg9RW14nijdwv9b6nJIYAQgz4HlMf0awenb1ENlfw9Gd+ZkaoxDIyj2JjPUG6vRgGzomGZYyEP
TjIE1RquKYzTMThTyDtWBQsOIsHulIgODVPxiZnAif7qLjRKav4d0rSepIiraRlYSyipfUVg1u8z
bR+i692UcTnAQMxKhHcxAjPayWKZf5+RQUHiVu4UZLo66t2dY+/UJf1nl+P5o7KrtbcG894aBzpx
cHRshseoIQc1ul5idNyHZbZ7YNa0Q6aBcu2Q0ACdPPVVx/inv6EePRrRY08grHVOt0AOUzAaJz1x
ecE22dIotismSDNS1YCo/v8FJ0b2CKyBFR+xjgPKDYnMnoFJNgpqWCoOSQDsFLq6mMiibMctnlC7
/jmJu5eNn1XKRg8gos0TJKu+2+by0BeCR2qyCBuAfxUhaKQWI12GdRMJKnoDTboNHHc8J5tS3jEp
kDScFsKcCxfuhYCnyucCQ5IbAGEkrty/I2CzThTs7tvpx1G3TUjKBDlHrcJebkFb++/CHXsN2Kyr
0HGx6OzJbdm9UyZQA8XailKKVlqTZiRzB3pHk9Qep7zo9c5WKe59PamVjJfT4amOhfdN1yI30Gxu
hxHE9RF+hsc/ZNmGcfhp04WvrYm64MZRgBW/VeDVJrFc57lppTeiRf+HqUeB+myEzQaivRZwo5Gj
+TEno8LZwLI7Y3T1WHpMnS4IH0P93CBQEnA5nPYtfeIWAXV1kWfhRwmMbeM8x1Ml0/uREWZ69+aF
gED8cLqT24gGhU4zIXhbUmNptExue5nVqUuUT97OQPZdN7HWvY4LQU1ZQO974JfRUZiMKJtqNPda
T1Z4Hu/sr0/oD5r5Zg2NLLfqY3PvfelA0PejcAekcyIulFWwhzoMRlE8H2gTWzv0Op618vcisOX7
JZvdBLEKKunGr6YW48a5NQ6HWbMo09TZxpaAx+xcojv402Eg+CU74MR2iTajKCl0/n6cRxhzQsxl
qpFGIlXCXv1wabU62vsEAjL1EDJV4AvZORym3zHT1qxomX4HPjpdoQe76v6732xsVp2GNgH/aUT7
QG6GAtNzowlSZfsjoY2/KxvANeGDUeh3t/WoO5qVSy+/pD3qaspM/m/667hgB91+9M6oh2XBu5+2
FZb9YsJQAnBTwQr2V26KUbuEBVUDPoDzRFE1NtSNpQ91vEm5iml26z1dBncG+BdAmEScVaS8q8he
wWV/QJ6sSqOuQHhUc2ca3z2oBaSs5WC4H2ePNUG9AwwdjwWKHMIgBGczDr6ykcRNCEABXTe9cO8U
kSGaUUQ/0wZJbCOPIXhzEQq6tmV0ehJ2OmfuZslDvL/KN3xKf4itpqM0SdOXf+n+mmw0dY+C5acv
u+hal4htjYYLy18IHlVRk7KhPtVQT50jhtrOb4IZ+DaKBxkr1n01mfVEx7gQ1GFzMLwQ931XJyke
uIGaMFGHMz0fkJlbYBD8i5I1qmwk+C+ck0vVf3e0z+B0BAFPvzeFPZX6Lye1Zboim6rdJuqYUYVE
JYM5w3AxgmZjX4OzCpbveI+xiXZNKhM20K35w6TF8I4ZgK/ufOuU7vTQHZHnHh53GtR0/0D4vfOq
qB+YSheADNjT1zq/eU3aB9HPXRlMEvJaMlwLf4gzs/D1PCJDXa6cKtY0TmQUzBfbLWyfJTR8sxqq
F6IZDPB+QqMbC4+cmKmcM5rhhMrBP2SYUjDCFXdDOzCYqgqM7itCPT9H7c5yEsEzTUBpe3XPTz3o
1yfJ/8eWCbCYTxAoc7HCu8SHMUQXEKc0qeC4fshgcw1a+K9ZAcpsppNwKM/xLpScLDnwU2lVHupr
U4CQW0po80XGZcr65hIww8P5hkBx9/RQEa7D4ZPI1fm0FeDGlXmQS5hlCIoE3OSbGfqBIEiML7cC
PiDEH3unmFeHT3f8yVczExijcqqoMsvAPOdknTog8StqZN+d14HwW2ziPoWtzie0JmGmAz8/usUc
QmbgERrRs5TB3iUW70gVn9A22WYLCJuRUJ8/GKZ/IeE0oVrIUs1k55LsoqW+3MtJFvl6gJgEZhDY
lsa0RZW/o2areXql8dEJBzHfHKMIylSZsBYe+KWJY/nCXWMfdoc5tgutyBWZjZNmgwJTxaVcg5m8
MzdyGsl/NRoMHQ2lnnSLvZ1Dglb5U+6l2enpsGwiE92wPEr16s+8+NzS+38c9eMN7uo13zIBe6DL
14yb5XN8r0AHinRuGeRfGhnHdyAh/qfn74yEsui9hS0te9rwbHuEk/ANKE2fJPHMPF5PKQxVMqQs
RdQApHyuC1e8DGwLD5adfI2QDq48K5JHfuAIyRbqqUZCFioPgsgPWY6X73fHzADF6albrCIXhibi
Yia6RbLln4iv4cD97Rfnd5SMbF30/nBZfOTfTicSsJugK9FP8Q660oJtnn4OeWPoUB1OJvP+KWYO
U0Ld2YcMn025dEEj7A2qNKoWFeO2D/lLVYx4nYWTS/UJg/HGfHOpLTnuVruNRJGjYelXj+DJedVJ
wVAmEYHHQUuLBVZsiR9KsZETBPEKaLIE9CllHcpQqwLwzWHEjhhbl9fwm79iJ9ZlN2+jQEqjHiIV
J59IMcT68ln9pZkztmcdQWN4BXirvd4SC2ibed/RMELNxBaVAA69l946Ylv8raNn4ZNl2QN6QkBY
qvuXQkNvmDqdzp8BbqpyBxS3oSd3RK/w3nhbNVP1nN5oTTLt4LfYSyEkqIbW0ApMVkE/6X1ZNjLY
nexyKVFOc0Xa5UVDMsw4a+ewiLOI8CxHcw1GqLvxglJHcPwA68B4M0+Jhu5udKu4jDTeTJRy0v/u
1rPNg7SAWf6Akni2FB9MndhepIjFyI29hs0uNjj3I+G/fpITizfY8auGgA+k76fOB/BvUyh2GAAM
inbaURAwDJMUC1ayn02j507fBh+AmVNdWFxdgC85GI0mqkU8/H8fc8X7zqQkFpKjVRDV2DBQ9pW5
SGfzuqsNfwJjPvhys0tO693pAoIQ+YiJfeAbywuUGtlVp62pNSNY4kRsvS8tlym8CeKsUDpHg8P/
MbsNF3VCXGcjAQcTvT17t8HsIQpdj1q3Bzf33C49f/Pu0pPG3Egh6dowbMlTU8IV3UAEpRIPuqam
S6D2Uum2ZXS+HFujSuorjFAGwQTtTphxrv+Doz924JjP1OnR5Jt/EECtmB2Q5QZTKv9ErRd8fgtk
YC+gOKg3ewqm4ND+WmZO9W/DzgxxMAYlvdLzIjU2ZJWeVzmXKdCcgyIYplBaDqtt6ZyBYWYHpk5t
QXnXjbwHJ2POpJJJl4Axt54axmjVsrLaktt0LTwf503wijroZ4Z4J4f5Is/n9UQWIHViGykwSGw5
WON72/34VQOyaR/YFCIz556Vm9Llu9NwjQxvKhxvVpxhjZv88BodVk10zMlSGdyHj7g54P5ftjGp
8AxN2NIV6m3NxRqcQL/eqyO6tkDUVUjWbBPXvO1TydvQTyDURkZBhikR+ZRMbXdB6vwSrc6MK1p4
xEWTKeEcxqhF/yBnzdWwc/DWmQ4qGwxhnjJZGqMfx+y+BmELC63CStbYIOOvSddcMsaubDqvWhCv
Tg264l3XyUaGfR6Gnp1tN6UJ6xRObzp8caTTiHzFOnKCh5vPd1DPE3u3G89nNEBaCQsvn67m3Khj
BzIB378iVKr8wFXvMfgfevLb3Wk4oytH++zSpS8FwgTj+sC5qGW+L/ULk9hnTbblQtcTjj1pn310
51vpappsit3vU61ndQORtU0v+g4YgPBKj3Y4BXUoFQ2bTP5WGcS0ILYeOrx5E55zP22tNUKFEWZm
P36izXZ2eJWnXLA60SQZ5wP2PrGR7ADuvcRI5zEgLy/Lo6clU8aObSLuk8C8ILWfvt2KNoAtln9H
S74WPG/Yvw+bLMgZXlM9L8SobvPUbf/2kE7XG13D4rj2aRQBvUirgDWTJV7htxY8jS1rJ7a2ix9t
VRyCww/QpYux+Ch4UxuDvNRkiMBeVwx+SXf/QxKWhUMUFtcyb+LX27GGwlFjAwJ/WGEEFEjQN+p6
bFn16J4gT3F2aY8EBRz2aWYcCUo/lxbOEzglLUKkHl+HAuJriXReieztY1O1NYwYUUT4ExpI8QmL
sx563gUonSa4o1RxYBV2t4bG93P32hUqIQbLoQGrwQxAq5k0FiqzT0xMUMR6xVLKnmQBYJ1meICj
gxS5CzxLDKFsKPx6ZdS+PBU0KM4RGvz/L10BrNgZgc3B9iH31mXMu3HBnxUYzfAGj8K2800n7SSd
hLcS8XFXpDc4ksqiIau2p5mH8SqwUBV1TbbFXoRR3hGU+Idd8aW40Amc/GQykVHrceJv5u04u/Nn
nWT0dvwhkqHPlUP5KFE8fsjydPaU7gmPnyMIK7L3qANEpHWtzbhDSDpRXlWYZ+UFcJ39p/LeptsM
p6+6V+v5Ko1eRGPEYWzY1OsdsYYL9WUWVheCXg7jD3xw8UnMldmXeyqkuOUHxjn35jxkj9uN5+nX
PffAHi+auxrU1z/FOvEvZGH0gLvPlZeWk1P04GCd0qIxpq9IaNnSPRfBY4FM3AKW7QJn0KmP7IXC
jT2qG+JW511YSGAxjHnC8FACeUo7uai438DzavKFrUy8LWt6EwLgJ+BWrX75hXAII5tVkoL7vjWk
75ZR8znklDYVgo9qOLPHiNe4aUaVwOuWKpYbpoZcD+VIMIVch00cA8PW1m88kxi9Hv4l1l/wGxOV
Q2WvAMsLqNv11QBGggWYJlalLLkUpzEUcpIv9OS6Yl2jVs/ywPgdBkHrb6Nqt34XcmFUc25kWjyh
h/gDCbB/VesGuSSbu4PTRtQcFbWNlEXcyvhYNO87QILo34yLf8dNU/1rV7trAvR+e9052vOgYe/F
CrFRRepSYh/DiYh1A6MebS8Nj0mO2uYqZixKrnFT1K0LHD66RhKhCqnzcO+/Etnywb9GP8ZpGMKf
wYrEP1at5eopApAc8rnvVQga/3iazL5N8EWffOKcta0ILTOeVqFY16IIQtfByc95yMAa7Es+eR/O
KiO4ymK6b3q73zuvAaoskAMo39kkqZbKg/pRPT7uM9fivON/qTuKjQFtv4HR+ql0tEwS4+B0MuRs
W9qYVYGwVT6mDZoeIGITKk3DnDQv6OFnHkS9gwUHArsS3pBlQm522RwzIqXMFGUNTEIWH41IwHuK
eoCaFmiDb8psHNY8rucCVvyimiLi3RBV1Pg4RH66oaEjfUZhLpvAuleyZbSLYNpf+7n9vDizK8cz
fEsfA0B9CZDA3e7yNgBzuYFIdjNOFWMz5Ng+RCpT+VEmCgNbrwvkBRVLgZOdPWnpOJ0LyQqZQFlN
d2XBVI5+rtb0FbauG9T3J8xNgEc4l2Xs0pwH+NjLlI6r7k8FkNa6LVaQklpjisggj5g+ywRMmDww
LypuDAiaAAH8cGjctUBlbSzVJKPwdxIbWEkQD3jucOCIfQjagAdTz47cCRXnMsfGPJmb4ROq8ICo
QdShyU69NuKC8PnsvbHVHxUOwvwFuQUNsOVuw0kwHp5/tUMpYaNsNHcrS8FS7in949tCGdPCDzDa
TauqhNtHXnxDAbXwG1IsaiE9jrhfC11ng5WMhVh4Gr7CMHxOwv2OD0KcQ8sOtQhvEB1QRf7MIxri
JbpvHiJF8LS1Mfg3OH6c+g5X9kHbzgVQUKUQgwBV39YJqnak5WKuhMFMACuXE53akuyKTY3w5kgs
5CiQuh18QeTK9yGZNYx2pTAgTF0NW0zInx4+ib/7860TKolfymDoDrIhoFBoBRKOZoTdsqw04FR9
q8c2zZBt34Ylirgg/GdGETmfEEOgBpKi7kU4P3jIZgR527abknlAyk91Y3LN8igoBo4QxPlQHeF5
8nLDMyiz64WJOTop5eYpgRisGd3KAlGyllFZoUeHoWrbQRC27t9Bi4i5adZSuKPs3O4UjjrEQwzP
+s9Tosf3drEifspgJYLc4wklosLuGjIMUbJF4D4z/PZBn6aaeJI2m39+++Oe/I/tRosxZCtYqR0F
vej66uFNP7dR+xySd1JanMPKJoCv1vOzzEfl2g+5jBYEDc4zrIOnFBkraEqrpWuBhQUa/NUI6l/1
d+rvBlL+Y/0NQ9fX3RA8ryrVEXHJo1kR4jeUW7qq38I8+OyIIXn4BZnk5ifJ61NeMZjSl3gqmgAm
NdFeZXdwbtz0av3Om2/0LFBf8LYIRiGpOavOrdw/aS2E0zlcr9oceo8wc4UkZvu255SwsuYz2vvK
lcv4CqmX0ZKJL/BaaRXf/ILAYd6Zg1c9jKo++QFMInjvnaRw42WzumTv1b5gM075QsNbrvYBqKiw
CAWA09tIWk3k+jSG4wnk4eFWCl/5Z4IBsJ+7a8rpFfzu398hIaUbZoJlqrWgHuAwabtk4RCRGX8p
v9tCW41b49V05f7S6eJQIJ67y9jKvSwar+xQqiVqQIc+SRoYar8g6P7xnAuFVsiPIxzEenjDuJAx
nHuXzsIvARLBUZktqCyI/uaIORePMlvoEYy2tIVYM8Hvc/crnlkzt/q2tz/lFToN1M6AW56pVK+X
O44B0lN507CdKVDxygJNBOjMuzg5IWlQyXL0ghfwjvthYZZyTS3qTOjq170hnvqqhWOUxNLitDlo
o425fppDHPaeHuYRve1OQqTWTveJsHZZ2pqfKi9lhpFxNYfdy6nMqCQTwof+bwrmUhZdVnh2te0g
6NrCwlqeYmIekll51l1JHtUmXAEDTjZDfsmuSXLLDgps7Hp0u3yOUPaE2k+24VG1HIBfR5Jt9yQz
ClCK4cIV3+JA7KmCp7BkbpmJtif2RIsYF73DGnB5lMvYd4twD63ZRkyF2RM9qslij1FUcSseo6cY
z7eXdSPf2NrnOPHfO9nwdbTdpBtc4n/+FYIlAV6ZskqEONyLWh7bLC4Rk33nU2S9Ji2SjZq+BYpx
oNnf4RzERXJd7pILvlrBPGTRxdqc/mLRakG9Sos3H+q+Uy7lANiRwpp+wmObFtTamQYARVkFi6nz
HldHnls2YNeX61JEMzt+9CLcMxe3geKClczV3n28bS09T/qzPdk9cpKIoWQadajc8KAxh8oxbFPL
93Y5cgE6MEDGNxCM1hH8ld4JaQSbpqqH02cjThDQBQy5KlfHBr51eu7ljqxVKsJL2Y3Ex+mzWpTO
QdbE2A+kSquFd7R7m/UdeWnv4zsSkXaBeUmk/Af/W9GwoM8RJBozT600Bmh4F1utcK7j5J/dR1xd
8lkfFVmxMEsrTQOn8HJgIg6tsNxUwNtpdW/MvCATj+EbuLBT0duw2o9g4l637Za5XIK30A0II7g8
3Pz/4HRWAP7Q22IJ7PLivNWe+cgG9J+emaAnO8ybyYGbwBOIzpLSaonR7Kvh8EhStG0M3jUM6OuR
oXlTAqsQT28//bQPxb4wWS62KPe+Vl28gHGbNevBZVy3LZrzLBr499z3sYQK1R+ynlymYSLsJvcZ
2eGndEpl73VJmoHE+Vn2u3MNY/WtQy13KT9OHk3p/N7sTr3CkkoDapakgw9cOSfsJuwV1OwQOVmU
2sFwLsoaHGO5kQdQD3oE/PPJOpRV/wKU0uHSZiJHx8ghoPMgoi/6XBFQKfSXm1vxUkGKtc1Q5d4U
HrdSuOyYxZ0BfuELw3v+tmSZqeeaotmVgjnHkHKYaY2jlnWYviGNy4T/jBcq/4w2hA20hyRdmhEK
3LTNhGGzurGtsClHbsSvHfAtTnrapU+XwfpBCkKzEZ2BvNUHwWQ5t64Fon3rFVBko5WcpCJDMWyT
MK/9CTzTpjuzw2iBb7CNFL7T4yWxd1Tkt91yWA8UegEOOA0+VCtS3VeiM7ZnpvPCoH3rAzheZOkC
BU+qlW1oY2RYlM3GuOSJsfeA6xLtv1EyweA7fMn25yPsj9y59eRkoolS754UveeKRifg9wkqqRXC
fxvtRXv8ysdAlUOpfnCjrvaeFcNfEXjtKKX8Y1HYB/q30sv6NoUSHRI9hqjzRvYJqiOoT59UD3XT
wA4VEtvM45Hsu1i8k9aYiOGOrD7yorB0hnw8PvIMOUtDsZneVWgHGoaumOh9icr9Z7C32CzVLzJ2
3dNMyvabh7tOe9n8wo2dpZHp2NzN/386Gs/j5J7raAKCtvORGfMsudKItvx91qiBp6NWtwkYtsHE
RJbW3Hix3/0WvimP09qKVII8wWyTROzBrkTLv0DggZJuWuYoT1WGQokJbhRlvJ2kzWjE25R+QDoz
1s1Nc/kKhPZq17/q13HDWao4fBO2P+/lyMgI5CVTfQjQY2RQ+GWPqddcIeOLdTNN+Hk+rHzHDRC3
DBMM2INblue+R7O10xQIF7E/hHh9BVFaQ+xZ0UNev6Ioqsl//QoJjgWWwK8dDq4qtSpCIZqXncZE
JsVBlDYkLbULoJFaklPXx9FaDYiFYK+d1Yyax1SKulmWBBsSto6qO92fSNwk3RsCgZYYU9Yp73zn
tFDD55elzYXWg1YdnrdLA4Xmbjlu2s284zJykTwG8r8BVD85ftS5/08B791Sdtg2mfcUbI5C1MQk
IYucrqWEOYVDBTSE5Snx7CLD0ux478Nzmec9+JWmVP99L8B6jMCaXT5zXdPSQYmpy2XpZ6FTwAKt
pqqqKwD+ZJI8RZdGgs/KEi2vW9BHktg1cCwZIFm7I4Agan9xi5F26XEOC/1G60/Aer7hsrXI1/R0
RSLUH48xTBxq1rTghfIvX6LfhWFrVXFdQrdA2YJcRBAD2mMWK3pYd4jfxYic54adgjoIhr/jpv1E
MwUX1C3CT3ULv/UwH53Z0wpr50EfeMNPRfipbmOZhB/40yRIy+wO2M9F+Gs+OXuPRzmu6a38mP2h
+VLO/v3IuGLKwD4P8bssQ/PKhaPKm2DPuiywPtbXMSCLNhbrM7Z0hz716FBeyCPtoEdeivUTK4pe
lFurD3JZCPTrv/NBN6W44ylTQo+2eMMaMXnN0pf5mYHJC94xaR99VVAAA6/b3jwI6eR4DtOw92k8
A1ZxlM0is0LgKgdyUf0VuE0ys9k623tmNHITMSPfI7T4U/DEpT4ta+3pk34JbpJbH517Kzi+jVrt
+fyZ7EgeIDVQTPEakaURLZ4r3XxY50BPo/Dt+mpHEvY5A/pCw4yIAkBB4uJmYKydUSO0pmN59C45
YQTpdl1L2F2RZkQrSS3uzRbxN01KwA4yRqh7rwT88nEYAd+V6sAFYdfNlR+/Lr5UdqfteKt7Y//p
x7ZRBbaYJLZoj/G/okAAGT6cJ1uSj6DLUg/ZigdLX6polhNl7NbRKcX5EfF9FrOZA1UMIaN7oJTE
ijrV6c8cm3xDL3H0T3MteWow5M8Q6ddsH7W3C6wZJDduKeDTxtUouN3MrnA5Unmqw5YdQwtwDsTo
JSwkFCSP4PtX93PyZTKz28GzB0zO2wdjIGpolm9hnN4/8ee17kK3SgPgzox72IX/mDTbx8kaBOop
MMlmG+osysxvTdr9fnmKsLFw80Vi55YE6pLicfDdP/9PAfPa4yqhegBcjtym6DgKAqdeiySVYd/d
kYuYX0PZG2mUdUQYhaPpJ0/IIRziBkeB1/Cz0X9jCWII8vo+C/jeGz1AZGiyjwkHgsvQdkPPrFSr
a0nbkm0iFT5xKqUGsNhylK4NqR/tl1vWtZ/cu/r3mdioTV2PipB9nqLpe4iZiyGDbHnBYvFnDY3M
Pw7tU3welTUimUO6c8INSueoI21RdUofnfuuWUzklE464c4Zpcr00zd+rE4Zm7mD5Rj8lMi83vQT
9wVUIATDRzleN0nB59dICRQHwPj/6ENZZe8gH7qqafZYDLHq4RnTxGvUi0Iv2/jtn+aoQGVP53oD
5QQCFbyKJmcuwdXor8JYsuxqBhPC+mh1I2AO1+8LkULMWigWH+Ize8gB4afI9LD2qfprsOMxFoKc
nmocfUrXqQt4IppqtF5FrP0jvqPXjLA9zxOBbvLBB0FCwpfjivonp3GwHMjorW5wSZQfA/pY6yZe
J8cqrK08BXFka+8vzT5XwWef1gFDyoeD1hQSI07Xur8Kdy/IWh9JE2DAU3LK2w51IK1LHFKIT3nS
Ipdzyrpdjm7iNWzgxcYfeRKb7KiKeYU6Ndg3iuW0zKCliLjlFcnbaDzhk9vdeM2hg6fpM8Cl9LjI
t+HgvwaY6qR7vsmOLf2CpGca/f7HVxEHeHTzNFoJ8/Xou6ILqcp1/L4rszw/t++Qn8bMM/EdTeXo
d4KrCQPwukJLlUDJYR7GJAaf69kibUkKWRRDTQXVwcFHNoV031fgXvb/T3l6ZORa86WFfRdOTsOS
FkjuY2+88aGswvruUHBiaC762znRDNeEilteCRfqHZe9Hj7rUm+A8fulj5DsQXQhuCw3S3KPHm7L
4yOc/IO3WIxzmxR65JzuQebAlvgm73Om/wHT0zKm9ihCFFD5w7DER4RP5qlUAikKV7Sksz0SVqrW
2S3qg1CRMZO8b+u1OYfv+NmR70WN1aIk7dOvsQHoFB4SWCQhuTa3G6IFs3JkIkIw+3zVt5XULrtE
XEuOMUIYx0vqBkqN803BnHXH+LwnAULEJXzaRL1v4hTvLqhDf16rwWuLRj/dJXzfJuaokGwIxjyd
OWNrI85Cy7M0VRUZ0EeGZnpHwiiA2+Uda+hzJ/1hCXUgPWVW+RoGzvYvakPqwFbz2M/oIzLWbWy7
YqrsAkwcVLs0Kt/Q+xeLgsfWKo/Yi917cW/xHMBy8hvKMXLPbwqFv47DY7tk+ywvwSXHHJHGzU2i
2sVqeVjb7iWjDVmYBfETs44X2Q2/quaf1akdW+a+3Wj+n7ybv3h3hfAhkebCZ92zP5x7eZb/YX7A
hwAob/290ZNuWQ9eQtmh9YM0RKAJqNqx9hKsC9qZUc54jWLnl8LgZFF0RgYMVtUq8CXPMHujtCgz
iEHXY45H86m/elDoSiSUPwNzE5n44RQSsilGlzYZU/TYmXM7vAKMkukkAT2ub4zyBUePEVyOCwd8
JOBdtpRj1ceXsER4YOsA+akVrFnAdlJC9/M29chW9xA+ivlSXlM6C4Pq/ShlZnvJzvP/VyCOZbov
kxLoo4fa8a3eRZeEmylcUJFtjMaRTbCegy6/aCp8f3WMTzZSFjdzKMy1IQyMYCjny3Vwd3TgrinI
NeRMwdM7WymhegbG5052n77bXIHfYqkmVPAeMpSD+fDkkDm/xnwC1IIZ30H9PORz2MM4bYTycFX7
DVDalftF61MZsOf1uMAYNYETTHs009Tmbyu011oI97cudZdzD+gNSxt2rQoF3LtYW9CpDZ5PLhYf
fyAnNi/NIPrT2rUmlgnMpRF0P1ctpjYBVe82k0SkXNnrx/l718nlJD3/WrLCV37S9AVZtS/z2TBT
xNEKD4LsEyMffYf2MVuVpAbj6MkohKCo9LRRp8TooBA06dFI8Ih3OmJZOSb7ljA4aQdH44yEXX0O
4R3f+gAyf+F2raI7lv/J7iPcQSMd6yn1sKa6scK9WoPZG4jPw+XB/1mSA7mofAy3Sa4auf2FLbrh
BcKBtbouyxrjWZSjFJ8qZzMzQO933v8nU46iuXhRHbjpZ+hwQDDW4QKmhb6fYWr//0xoFYevG0sV
vTc775hoRInmq5HyHeIyDA9uvsBNzML+khHMC+OOI/B0WLJuZ/9dAAMejBWHrrxb52SQkEr760t7
2pO3h7UK/SvQ8OdOtlyJM/zAgqzqvN5inu7bTgghjsPXttH9OxguwLE8UnazYf8yMN5YXJrzIhd2
eAIu23bcDOMVKnm5++8Qg2hd3bowlA+R5O4aKtwm6t5Hlxoq7gYBv1HeJ1zzdmivkMTa73Dpirru
uNJxpC9Rc4cYgTYFJlg+A1wyULyrmgchPjqhVfXcMiPB836RjfJHvbbgEeaUWwA7BsvLkBpO/nAR
PUSqZlxTvKh8qNxpcHSNS4RGM45O2pb1ckDqz30qWTZAconqEXzw83vz/ox8pC/FiPWuG4oYUGP8
UsCtxyeMCP3a61MODgCiOX1ng324Cw0a8095D8N23ot6aZGk4pHB97V4NN/Fu5O3yWXjzg5bTaxI
rNlwsUG7/FGwWxZ0TWa5/x0/VgequuXsMDlyJAF5bcJBZyAecvj1LvvxpsOZVuIsc4HWbWhTdtWr
Pkxk8L8plxTlhgRcB/8FFCxiVoYFFfhdOspNh7qyF6E50aCdRoRw0ge74oGi7Klwdlvjw1bBcFK4
FcFFQdSPgSmClkNn+FnvBAM5Xe/I2va4fOunUkoZ8/1zudkdS8VmU4rB8bq+cYgF2wuXiIBDjnHi
sTIZuWX+ddQdK6lt56UMGX1b1ryzd8FpG9o4+2WjPdQ9AMYWgnYlKkaApC1g2+ML0ohndLX+HDFl
zVfAH4SLIlzdO3czd5qRXYPBpEA63go6ecBzwuwDAKO06qjjK1oLmL9OJUSbYJ1VBiphPXPUW90P
GCfdBdaKCvhZUR/mX4sd4n71OhfdYpBgjNa8TMGM21fye1DSpNFzaHWcYJSSrTvn7d8r54vV+XNt
VxJIXwzeKL81jIFdzZ/PphsWhtezOjsOzdeEXqhPdnpIfTtZ2ybKtC487JOKm4lye+5OONcdL9hf
6J4uLpBPwErY6fKwvnUssKX9fGZhWTqpFQK07l7KIo3bOO0ep7ti78v5F4gAHZJs2m1Fe7zW31vg
UT7BKgV7YjLTnU8pwve63hEqDdzSVlel3lIB/V5Ofb+0Z5QG4RyWHP/PprdXFm580ghdYisXIQ9k
ccWmSDllMVJDU9uJHiqsmAwKPI49dcUUORc2vHoIQcuwuGpg0AUzo/ktBHnLPdYrRYxlKi0UbTb2
DWyLGmlcMudq5k2IkV+egKNqkqI1iguRVii6LvGa7lR938LfHa3SgsGIbqxZ2L3kjraomVQNrbhZ
oLf+++zkSxJkAl0WgeOLDCH3OarlYiopaFxczkjkYBxfhxySLrtaLkkFi61hcjsjbM4FL/pZyRTh
Ihu3QbNyI3qIUfL2r2lo9/vWkFK6AI0gvVakYgtpzDiXz33tLC0iEEOFLg2iaymrY9OCDQfJnle9
aBwgl68OtwxMvQ/sY5B4QWRgaIDpkdNtKrN3hpyPkTjsVIvJwj/yd3IB+IhkhPqZv1eX3RWa81KG
oNTZtGw+AS0CQJAlejf2Lmh/2jmL9JuzhAFlfHFsBGa8jtHvcVdKjIVKqL767V7XVisnM2B73KbA
vzIBW3a63LnN2nplwAbPtO7/YH+X6zrU97keeKhRFqA+aCY2Q7CqPxPY9E88PGa8pr5ACuEmO8Mj
u9iPwqAMTvkXRyAczB0urIqWEtC26dhUhaIkGT6Iyuo2teH+eS7AxL9u9u5vEPHp58gzQRvzepCY
jFfiwgEwyKqK08P07YHAMj3W42zDxV6190U7b5wtpLOc3qqAf059NWpYG8u3rMOminiYqDA5B6cn
r56S7izv6pFWPhZ+UE1I5y9ufBXSMFRrQriM20xJVfGBPfZo6869BnfEUt+zcdo+ZC29GxgVu/a6
R35E0uK94VE3/4NuzALBzqR2z8fQF31Rca7vesdxb1/fXrtZ95oX9DAG/ynS+P2Hr3dPXvBWyqrr
UTrQx4vb5TicJcFkjihN7SNME3NvldoLBTdiQ1FUZQDu2+lsYUbWEmgWmVYax8zvOp9Mbs0jZqa/
gPFnnKv1u/nzXgsixUzF1nwn5dmdrxZ7PUZLDxPqx5aCXUAt7s7NDrtH94QHDtYtaF4K6ZO3i+oJ
skd4jgyx3bbI1IusuFm8sAm9/DKXCfZNi7alUqsf8UO5KRXH5Xrn56Y9yNIgXcwpxY5gs94TzRcO
M64R3mozi12dhF25LT0YadFnKw3S+ZcGMPalmrkTSHD0mxS5h7K8UqOBhf6rRDV1hyLaspH14wz1
teS65kuX3Ik+fVZxwo7C03/Voa5Ggu85gVVpO5zbMUz/z8WnGzyjRhGDRE9MAsccMVDM9vluSZTp
P+BJ+SdY6ubY5Ugw4rpBbhUJ0RU1yf4dBOAL37rQlGesOml0LReo+w55DkjmbzYomtM9r/rCjSEU
HEw8evlXF6XY1RondKxHk+aaEOoKXuDyLGdSXCJF8tNiR3tCydglXlgno6E3rZ/8tm/HOCf9N98R
NVIhfBAsYJCTKtNOd2rciXrDTnIbw8meTGgiBiurkPXOp5pgDUUf7rpHcwJK6KgFBLS0x0k7OgWu
UIx9398xs2oFQe2VBFhoY9VW2epdiTtBIG++aznkEWxPR4ua2baBH/9x4FbjiqV5KOVsv9VmfozR
YPxkXuTzaPgLIKk13L7+9B2scwz2DSpYnf/gkb6W01hiBZ7JYwvuYnb5xJdO/kU6HoIG3Dz9wHV7
KS12Gw1aefiYGZpesVSgNetg98AHm153zRx7+5FgJTVEf3BfI7bzc81qPtxsF4+CfSJdx5AgdWhv
ef7aj6QNJmYvAjjE1vi0FBQma6NJiRv0yju4ihOmI5HpzcyHGYIwYYtUvtq+Pb8NoBgf0MyKurbh
u/K+tZhJcpWvX2qYUQPfXMCs3ggEC9CVPRsWpgUO/1EFF5EV1YNGa1TrBfrGtQA/R5AbpgJDGJYv
juMiNI/IazmwQwK5jCN2aNHougFPTjWwaHcry+RxI2AUemFzP+5WZREDXheXi43w83tnpnWUZP5u
o3oQUl/Ne3VvJ33oL62n1O3tGn4V8dtBnyw42DbPxqNMxCG88eRkBhklJPQgMerhJjeJ1bKJTheY
5i97pSpMYVsSMu5FPXOVcbteAn3B6fytmFFMff0lu8aU1z2x23iZ6ORsbYJU+DYlMdwFgvtAxVjn
8H9gkU1Q/+lmD10QyES4M1Pv2wmtTLZBenYgujf6EdHRcWFOETqNdMjXLFA432g2Z+L20OTj6k40
TtKfKGYsUUqgOTKzCv+TYCXRF10CXFo7gHeV4gAoB8zO5Mg6pmlossLEKWNHlaE2yecDT+HMBUC4
BFA+Y6YCU2Dn9pwyCmJv/upEgJqIenTuzgp3nbCBehDSPTjv6xLCYjGo4akTUwmCXTOFcS77iP3J
abBhTev/RgFMbKfIcNH6JMfOPjW35OBpfCmvaCpQyMQ9grKI4pKWsINA0A35L1J/g/GQ3pbrVzfy
3yRceNuvOxI8/Qv21r+u7nmGf5gv29oL1Vbs4K5HJeL8iCCqgiA0iUCBjYxsuBD5U81T6haa1Xbh
9YAgSObeFh27SddclBG/3wkJ20BUhgfF+iu4obYwZtjicUdbojXXAYgGQIcWt6dD5SzDp+kNDx3r
KZApN99JRyVNdNZR31v4cnMwNnyK2v/olHHoYPw8fI5zFtyLg5BxxKQqJTBSxD2oBkB1Uv/NMGi9
uzJuGc5JVEvbcigzU7tKnTOi7DZ1BL4Ae9OjR7L+tAn0/FbSndUrsB7P5RgilnpXYBSuS/yA5eu0
+GeloVnTIPoun2C1pQfFfODPT1131sbXrpWqrkU5MucVztVITL/5zcqw00rsRl0XqylccT7vK3VS
TVrbAMf17WBBJ80R080q9s5bzE1bDeFOhkDa0rVFcxnPSQfoD6Qr5Tic0ofEFf4ivRE33exjQvvS
HgGxVj4TLlNKGqRekUGhmYw8IGOdPUFQBNGGf+Yuc53W4f5wpOIxg/ezYJS4sA6FBvJcO8kBODaI
+9GJVKWUMZ4WxbjPrMASpQeUQSwE6wMHMuslZVVgcZ0UWqMHBlJFtkSOg8E218mf1ChUiF5lHPDK
zcFnrQtW1gQeMM7CI6WdAbXZEj29X0sDYiw/+hhOo/wpjlm4AE9lSMoG/1wHZIiumBsF7wlbQthQ
2S5uFwoMTywsZs1Xw6FVaoF1vnZtWsjOWw3ZKtusMSnDJf3DzTwsSfK0U45LRD7tIi5+Jmi+4x0l
+jiDNvOi7uCVBrWdvEmIeehDW9jMBnS2wPy+ON1OrRGjCzT2ftrid7nTun/exGMctgkDpebrSSf3
qcBO3/Nn1gXKhm0LjLjYL19gKvjnsQ9WiHa9VB/2tExJwuHWBrFYl3kT2pJ0G5/5vwXxiYILXOmJ
m0NbVTB5c/3UIGDMm46l2ONHDX8WFpPLB++PtHBlhz6YzmL9Jsg+o7oZg2h398Kw9IlIMNf+Urhx
hIjTldUNwXDwK5Ftkn7QHxjt7j0AbqF4EkRCFgACRIQqd0umMoo9y2hRZ9SIg0rrgQ/qUFJulnNV
GWTAWa+GGCw6Cym3TFedG4Q6giNkTq4GvvnvwQWnb4KlwxKATVPFftT0h1RuE92kmlAxSAFigMAw
kWb7vvWwbVoBVNzthcy+IKRpO20KNuSic6t+4dufpHUfd4KjpG0Cxb9Lcf9ELHsNrLsN/j9NAFtw
NrYMqebwVDv7GTWE5Vv8gD1wczfuOaRrDVU6qWp+qOt+uykeWMx19sIjXfnsXNWAMZXYXHUhM6Lp
+PqCUxn+a+9wrJwHMXPp8R8QFm41Koy4T2RzpNBtvipeKJu9uTQ5yzNn06vAxXOpZtav6e8GlxAI
iEycSdMM4OqxfU48o3vNYNEx7kMwBooku0XYjePnIpoPlcds6hIDvVPp5qDDPg7nozX+qFtLTeOp
wSdCzWQ2QystOEhuP9EOAp6+ryFdppSsmRIMSd2ygnw3vb52oUFjUNffAgt939lC4WoHvSb/+hPO
2KYDZQHZs8xCmn2VozOcsib63fEzZec13rK8d2ZUq8vDC/ERaZ+022+rt2WmPJhSpiMMj5L5swwn
MgYP0QhF0qELH0XCIFSDUCHmXhWOwU4XuUSUM6rnyZUCRCOkXmsPkRoHWxzPJ07hucWArmMnboEt
ZNlIsuyfNb6QuwrHq+jfCO1KmN6HMdvdvfW3mojuFBc2VJ8CbGvOvp7//YCyMlnEGz5azI64qfqx
UwRkIDLTBa4ncX9gdn5Qrsftsbd5dwP5ScaAMDjaAZmK5g8FRFonxX52rQrCWxKo0RNOaXjQJdFF
C9acDRtrrc3wSi8N3eW4UkLvEv++WyCEe2/wCosMUP4oOricyAsHxZLFhwtAkxZ7+kwAgvsoJHk3
XKq/3jwdIMweJlgXYiKXjPZeMYIVfOg+SmbS51evSLakhLjLmsLDUsXp9oU02CCYvPUCPLnNKOnz
4WWlRP6GDX9etvxT1N7PJv2YMMA5lc6n/rtiUJEhwcUeAARrJKgZgOAuLyvZwlUogHBIWQI1w5AT
FcM/cN7CVUtQ1VqG4j1giIqheEcLzVmD+Kji2najsmroDhckd0stLGZPy0va8fAGFpTQQrSGimOh
Wl3jgX1Y0lzkNnD0qRmLxKgjnPEdPMJImoFyfuNhZqyYE+fyKbIlrzYbY6TE+rz22jHgsHAcyPa0
q+i3Bv1QocRa/T/DSl/N+jNN8Eq+qJ0xGJBz/CurH6FMYjyJ8v62TeWJ9XpUBp3Y/MrDXKEbOj6k
oO4FUYF7xhMl1TAxS2rzVB7Wf9aL6H5qHQFUs19xXyreBGIB5v9Ba9nSv80VEcfjGYXruDQNTrQ+
wApcRnOmia55ovBxz23F8+D2xlwnLVtkNukrwvXATuQtPZEzP97J4SKnUdFJFwQpo6NlpBDFSuk8
lAkBOwD/Bvift1zlDNrwts+CWD5wV8lQxfQV+50I5aTi0TPCp2NMT/mS3NJkgHNazOtzDFjlSWz4
9uEmKHDl/3YEFT9J4wRwwnmHB2Xi014Qb5Z8Zy33V7jE6dd4waoMwb/s97Mebh0meOnA/w1pJ9y+
LegkojB201+t0ikWDPSSn8NXp7E9c4gn7DWRZnVGdDWtwLplb+BJqrkVQPPkmWUnbMl+22UEEIeu
kBYpC1aBS2cdpMp31niimTqCeuwtlCgZMYzK7/3xX0Gv00t0FHNs0bx2cvxZ6tg29UdUQzWElqtV
s+mH5ADlUQbcQUEbuuPrMsWdpBwFVaw4EnKqvWWvf/EE/M0iueTE9GJz4F49WgmA79+PvFcIO0Ti
qEm5cKM6mz9/v8x86l/kLiM8Lf/+G48ybQmtNo00LEMHQl4pfA4Zo0fdMyS9WrjZc0bbCSG0lkOg
OG9AOVPMVQye+CmGfdNGev66DjT6T46K9jiMO8wNP9jjswbCIjK3zRlvFuxwsg5bJROaObzgr/RZ
gKV5u4jJcfA6PTnbPq7YuduMcvXkRxGHwHeOMI2ssJ3sxgLRMfLCKTUjEGcfvW0xgEhOuTZFJJvz
b97SYlnX7X2jafWbHfW5lYeaoxdn36yznbQDcPKRWUlECax2i630RBpxpMe6Pod9ilTkd7YUqx+l
eEMN7z9NmNC9mtdiTFs5m6kvde+7ZauKQURSOiqPQIYpTxRWoOlkI+IfcukdddjYxrrFonbvwBrI
CY1G2Z23amGqB5khW7cHrJXFCAidd6Huw5fs3U7lHmLlrUz1QdgQr7elVAPTMO5mO8aoCGoc6anO
mpVJov44OqMjIrFNKWoe0tRruAoW1ZY5hiHHRzqytSLkj8iTQFE2MFaA1ktDwa8aUTreT7lILCU3
rGa1q7rbXPlmtcirnmWkxE9Ixbq6lqEdhE9E254XB/pFPoN0Wg1T9wyCQrQXwlLVfLbtJZvTktMn
IAfmq8EcYIA9BYBAufi4c0AsgLmEznlUZGO+4HxpFJbXoCr5FBUoz8kkWz1WeKlO2hL5v6SydFyR
fDuEdfmjS8+QmObCntSGQiW0nXadNmRfnXUUf1xga9bNzEW2S3fydDN+lzh+LySp6NRY242IBD5q
S3knXEf7eVBb9PFO47fx8i5LxeSctYpOTxSWSm7ylt+Trvr3kiIkQY2maTMM1obMxxXZJXfUBouS
Aj8YUs0ekLFs1TONmNXC3+ctZqKfOCrOUf/rCSC1GVI971K3sbSwWH4VFAdkJlJhQ5H5XPiZyTQa
hTspahKWeZe4RT224DJPgGUbzjuxEacthTjy+amJuRBi1j3O8iYZsoLEfiznzvQnKHS5SF6qmIZW
T/EVgmZEsg9WMkzJX3ihdLcpzpAYQ8/47NC7saeMkAhAiGoIgP2fDVWNtBTjJqeRqoL9kvKnCCXQ
Mi7CcNTKstkUbJ5JulCRilF6IXkndZEPfh4fltlkTHrTObQsDpyRR0D4HN08HQgFodG2x/SeIMLP
p1OcPy10jH722qb4SntQndndsANtKFajP+qwrWXTe90rJGrAIHPxBxus3Jm2ZylELqi2AXe5YXa7
NviMD//ssVehWMaNIJeatNzUTA4Bh1xuRWaT5EuxkXyln12WDtHCaouRgQrIr3ctTDncGApwfbsQ
VLHfqv5qjR+bT31P2xVwlMk/gd9qelJMzKnEmEts/gOj1gPupznyztC/SBrEzbMsPCb3ugRrXFpE
k7pobglXFawf5fAOlX6VjjV0xGPDp2Bzl5pEFJkeU83AsjEyboYzZeA+DlMUvoOcjm+QT0xZOB+o
2SRFZv2I7nDOXaaFllEvtdXAYb9r2Voje3EnUiBp3cW+dSTcaV0gzZvYZuncE4bR31lyz2cs+PQj
WH4FL4+6RJkQtJlXovhllBJwueooeao+278ts6Ykaf5vcI8vOrY0kItliLpSvmst8Lzxk66NGE9F
E9rGe48zX6pDxS9p1KggaLYKCSzieR3rOZr3mxgO+ZPtcAUOsn8u3q5j2v/L/OC5Mbtt1KN8G/3I
PWtGP2HMkcBUH/s6WQUegVjH25RkEMeMZ5U60oqKZtWUqS4V+4nJUwIg+gn1wuoPuxiJSPurFnpi
jecWa9/5RPyeJlCBA8n6VGuXRGu0ubMtkIW3uuqfz+A88/DDoIfd+P54yq5tKF/nikMGGDq9WLWv
Am/JnDCiASmEyCYMi0bHb/z2hP0PXc/2GPk2ue/wY7C7b6fvkREFla4NUWIoqiAizCflyadPfmMY
NcdY+k43ysCOQglTjR8LdNmTfnaga3zaohazbuk/8Gy82RKlCXti+bp8hDzWKQ+jV5Eo7zUO5NhN
d3msMz8Z2v+n5rd2yElcZgRlk3YaLtuUqQWucZqoo3C48tl+5It0bE5rSBHnBl0EalOfJKn6gMiz
KYe6IWByH400MYHzDYvMS6r2PP0HTLYcDjRrh9mEJlvuLrNDPDiK00I28Hc3o3agPmg7ol27XrX+
SOjHc/k9kuZPGrDes8mAW1wa72O6t5bPtdfkLgDWELj0of45vFMCaEbTf2H6UY93DoHQeBWaj4Oz
39Fx2m7i79jDZeLg+fAcKBsEu0xT703TKS6319QKxfZQYfctTUSkmY1iouEsVJQVPXUsNWcVDNMs
qGmcyuYsWMEGcXPTZask+mhl10MTzvEimecI2SaILRWdhHhUssv625iyjYPk1u9FqTK7/FJlNkVW
dQw9z1C6+RB6GyIjz7yiPr0fBeLeUOfxvz3aluEZ8l05SyTQW0isHV9znMDk2PdlbmSH04I498Ma
lZtEYNMEvBURJ8PI8xaolzEsgelR9IoVZCs5PB7Xa8pA1mklZ9l5kKtusDNtAUYlj/i9tWI9XyXa
vpLA3lhh6YiGLI0fMVaorBBHLV15RmfjOxzN9bSgQSfJnYH/AA8RbRYpB8AOdIaxT+GrtuhORuqt
JWLvRkKZHTjHz0u7HG3KeDx3yjGCt4hdpMqKOp16UkuWaeAnD5NjLRmhMoebihHgOeSyQZ5yhTEu
aktr2XNEehl6L/PW9OOLPDmLUIEqY5/MBHV13riRRngWf3k7ohhqc5Cuw92kQGoe/sWf6G7V7KHR
AF51j3JvgR3fs28Ei2gBfodPJtaQtEG0/+2wGmg9lg1XyDp+x76HpLSIqZ/WwudxtXbUyDKpwgDQ
/OptJF7d2Hh0yZn1Ha7qu/IIFLBZLg+cBbQDvl+uiYFA1lmrWR2vKtY83+lkfyUfMWq32jz+8qAT
asS/MkR7svMyPo0+GjQaTcePyZY1kdgQz4s3hRHVEyh/bA+mPKnOCVQDmu5MX8Nc2DLVCavh+gb5
vt7+90Gh9XORSje2iKdqJ+KDy70moWEyf8uk4I/NVnV4F3dd985HSNLvMlbk4dqggKcaLOgzPqDS
CKg6vx5n60C3v8LwW77t6xMnXJiHTmO69JEFbreNHf6er1k6LrsoQCr8KADrMa4aG3qszWBN/pb1
1qR4NBZVJuJ8R5JZpZIvpdqfaF7LdMw+EN0O6m8EkHb0dxVBLVQfv81uWf5fqHqXY9DsiOElThqY
A++p0IK3NDcWvnpiodxeXv8lDg6U60StymLN1vh6qFPjzddHPvB8zS+fhRT9IJ8Q7UQ1KznVUMVX
nYK4C54FV3HCO2RIuY5GNsqxLnNz32zIz8+MsEwHPEy6qmoEZ5bgBDIyoU+2y3TBot2oggSAhzjz
yFkXpjZIcD5w1KJVU/3TNJFgz+rDwEArb95lH9/WZS99JvLBK/SlBlmM6IRW8fAXfZASqZtZPr3p
byUEBqGHKgKYQ5U0eexsRFyRQkMe/5UQdLDOlW1XKy8oYo7R9YyW/u320fyBxkJArHd28R8tGvri
OCoiYtzPExsdS8c9dKKcTr2NSkvKGXHBLd1XNUfhBeDOxVhtnapmabX2b3QgoeODvDCo9hYAk66u
7tPNTKwHa+wCYr1mGc9tnkLjfy5wJ+1R0BIJNtSnw9wPPBUt5YI24lii2+pslyovdJ7IyTyMyrK+
SCrOk9wIoRXLTIvDROmHg2T+1h1oIpD0U3FSJt7sZcstxC3ZLcp0nBKvMsoxFANfDm3qiIlYlN+w
yvZj03aPb503FMCXgv1Rs16WZihllxZBeJVQsFj9ETk7/km0FF3foOjJox5o3AqAKrBKe3UBVffw
JntHAGFFKvxRcJpdZrarlYYDw6qXq5jpP17nS9os6ZotwIp6ASzAYUgv6cGMNSShMHgl4rsSre00
T4VRO9wZ+rfNBU16hixEjwEFOir9BhJch5/WJKKnAA4hSekkLdf4KJ2WjLwldI8uCw0VW9N4M2LR
JauqsFFtmCNzGyIn96COL4sk8H8aVlg7R+XYFZREfUeL8Sn2OqqASkRR3IRQcCYy9MWGasW+w9vH
jxEv8lFQPtVkh1nluVPQns8FN4U+/LU9DwF3GiJNW4QnKQqaRmBmEJGLFp1s9eQSSmg6rsx/XACj
Hm4tABc87+pDixf3spypWhtwH1FbHgoYpeKm9fdpYkyF8t8CyQdHkObjK2coOXs4+yNNtJdbFPzk
DiA/X4d1dDR838f7cbfzMWyw0uUpIqCKEdkUv9pMU3xnsuiwoVn5UFEmvi6dS3i0OFyPOLSVPe3K
6F5zrlobCnHsndQEdxSZgrr4FmsP6TP9ES4P6DCOwBIz4LO2/BNjWiZImwrcvKKu+AHr6BB9T8ru
l3RlOSZcpl3iG9jtds6FVl8alj+Obc+Quf0GSP8Ue1KNJGU6jqQgKQvA4cFtbupajAbaZiTdRUQ9
IwCUAvo5u8njyfOD2Shy/2gYXF7HGetP429CKzO49t+5Sra6BqCwfqyC8tYuj5gwHhS1NIchnArj
tnJjs8jbnZO1SPDoixiajy2fIJwStj9dKxZMB6N68OTCleMA2bn0hguFUCh+xJxfMgopfOsuEYSx
f4reJsmoKvyj3mdO2g/uYJKnp8LCT1jSChZjXF+WZEsdyWKoNyFSwNmNJ95g3+shqZMQtyOc6izo
sWRAWx0X4f0DrgR/1ygTmODIQDw6RlTG50qyVgTqa5rNKHoZ//B+TOjx6G0gtzExcJLZgA4zzeWG
XMZvqOTteVoR/YisnJ5Kw6/Kl5NQhnwD+1U6r+rnCHH014BuWQBub5I83p8/KWbc1Rd7VG+DPctg
w5oDsgEf3AJ56ntWMBjhrkOAoLGIdT/Cz6NwIY6oPZmA8E3G/pGWHncSENYaJCF0kvVwtGQVKJed
1e6FiYoR7TEVEbjwbfD61CTLlo3H94km6ADg/mkmsrj5/j14/sfgSc89+LtMurzv7j8xH+ydm8ss
2cg1bIMm6XfbRrsB3TXquxK+fWzPkLhFLxUgDS5H0Lu++cpefS6eh/kJaoH8Xcusa33Oa8ln5Hz0
naaNpXMCEiw13kGLhHDKvH15V8a+S5A3mMVQypJ2EoHm02mADgK39G6wpdR04I4Zh/YXgUYhLokx
05Xz+N6jLq5Lcr+WnPiW3qMwjfjMz5mkTzCCMe3LRqyHD6UfRSe1P2xzzkbpz1lRJgK4eBZ9VY5i
9HV2eKDvfL5rZOCrQB0TiHOBQa/ZxNZyS6vg+eyWEopeAsfunIjuWTCZ2Ww2ryLSDoehoy7cl8ur
4R7cZ/RNKKBGzMbkck+r9I+2pPDWYdecUPdtn22Hd5W3hG30DXHrrgiwAXKVadJ/pspXjE1xf6kD
XAE13c02kZb6aVmYMu8AJulv5MWGt0qoxOkOrqVyq/litA1dpuAH5gXoPB47JQDg007B6/7Tre7z
bksXR/8+nS/zWh4pZhU7hZvLiSQ7HyjNmWbRYH/gwBP2w5GvKATWn8T5GlY4QcYOTK8DEMRvK7hS
rj7OWphlHbH06OOKxvv5J2eTO5WQZUJ1JvFTHDvHqh5SMxF3CM5vy9DHGks2keeJON3REiO6Mh5L
94IJ/jOiznFUyH2l/Co/84aKn0Hbv1FOTjvEyCXYDMsFsvtr02RykyxEK8MjX8MMZi+5HMhmAyjv
kEdb6XA033C8+G+mYU80Vh8g3ENojDfpZ5soKj3KU8JCm5e6zYmgK3n4Fxpy42vTaNknNyUJMiRp
wHZlDrSC9oVf8CsSMGrp2LQ1zr8qcXgJowS0Vj1+WA0gGiIyVbqXrW/W0ZKfBdsFuHqVhc+f5dxt
L4OcCMBynifjp/lEWhCan17zDX21/Z9Ygpw+utqioDTt9cPIwgzmUnBcmeQONZnW7VhCoiovj0gQ
wbB02j9Ub8hmTRlGFyzqFyXf5b/aQ1hxVmlmPcCz3MopZ/FEAMuXopznoyKAsjuDEzE7V1uAttQ/
pW4Y0kjU4/AjOPD75J3pAh0+QfEox23eDGaGILr1+7b8pDFDdkW7gAgA27q5Ybpeb06uMYRk2hTp
D/byknjGewWnhfUsIeyiQWYMktHm4Z5YY4sx9JZPWxaYuYucqZEzs8HEePFvOcdHKyngJ6ZZYjIG
2cZEL8osndfi4GUmyXpWTbzrY6jwUw/SAEEV2seOWsVAZGoi3ZKOmSQHGjpzMcZ4v1BeRub0Kd2P
LkvCP851I31gEeApZfzJ4JhTmX2Nyz/Zwq+cT4ho05NgSSYSgRCjiajwWP11ZzNX6XFraFVghIEr
c5P3si9nFZCttbuU4oK6BGKzWSiK/bs1x1Q2Rsk9gKQqheLUx1OLSQMdXIJPNMyK+xSoWJmgVOMV
agCtPtKBIe6VXEGLDHdQX33kBvfKawDv0U4eFGuBrQiUucBFHqNsRUuV36EuphYqmHtNexWCGDv/
0aU0KKK7CKNPbloyrUQiM1SHaSA3eyvCAqPNY3e293r0HWHhxtF2cStROx86rNd2m7L+EF9yIJaw
2l1H1DTmi+IdtNqZGLy7d2ySPTxcpdPsEE7DFxN5DltEUwyAFuDOSl/Jas+QcGMwQ0AbuUUjtDvg
g4RHAULj9C0BWfqWitFau/6B8XeWA/6snr4vYYmSIyCdb0nkwWd6fryOEC52Av6EbwLWvNsc60kx
mIEibNuUalX8qtF6jpIMCKWFs0dg8Dfn+vhN38fRSwbR4M1H2fPtWuNB1XIglKvPRtApWmDiNpCj
VhJEsOFgRS/Whgw7NR8H/Uoy+2Mn1itBNjdvPo4dD7TA2LiWLx2XWRiVc0v5b0hiyxIN8NEa4iGM
7dUmU3A3tvfM763lsdMCf5yQjUQFNW2d84tW/ZD7FPoZhEkAR8aVDj6IB7YTQUXc5GCpIGo4d5jH
C8awM/S1JT2OkVuhusGApvR16J7NIeWEwWrRMPZM9ulN0k/ih0JZs6yZgbW1aP1Ap4hxxwFf0xmH
34Nadqv0FckfAX+NHDi4ASQrLQKMMXAjPfGHupD8w6fWWktcT7EpSwfyHCRJI0YSvqH2KNQtgQrC
KtNDmntObo0WZZbdHodHp2Ifgyg7MDvLz1SMZbDfZYPG3Cp+NxToDI1eqrnxx5Z4IXzwy6nf3fZb
PIBHGm/D3Wx/OIF23aBeI6JhqAUEBDyt9pKbys3ELRtKdzRBrjIUTi31oa/zmpuak3voMNkfvG5d
jXrMspGoUmeLA7H0Ekl5CP4Mkt3/+t2mxW2BWcXDHTUCUZkwe7dMr4wJrTwoYF+hRIcwj+q+XS3f
dJpuPxqM4TDN4bgOiF4XqqvyBuGFZDZIv20QkRYDjszNn+dNRO1GMshrhxSYfg7Y8V05Vs0HPqg1
IM/Mv1WTLkppnSngyyaoZgwLspcb2Ag2szspCL8UKi6uof36N4riBMNuJ4NjPbGh544Kl0Tl/30n
MvoyXzMcL54F9PymcXSITmYZZ4dTvbNCdFb5OqaPAEEdJfq8LdZM4m8OVtHXi87yeSk1osB4ehr8
xoZ7qFBHOG45ZuJ8ESFZTiIpXnNqhtO4Tc5H2Z+tPxs28AKGp7GBezjxzpPZhNmcxHYKxcgWPEE1
riy188GjxZuAZzv3ETyKJiUE7WPJnsRh0BdxK2kXq/vF53PQWdlajUXILd5uwx8yEC39l0/ZiTrz
GFeTaPaoUbmuDrKZQ8q8qUl3thecRdvgjH7FPpbbEwvoDgqtSzBRkXzKXrLeWYTZXFEC02XNwAtr
Mk+Tuc9u3uNDfYnzHMlxT1pqVFcnro2awdsjcrwfqvbAL/nZly98VeOiIYp3LFRXhf/rjsyT2qQi
ScsBs6YuZsEy3lnCO7umrsRVmkhTrV07z1A2ATUPCX5dqJBUrScKEE8vcKjUM7UwkFP4JyiH1Lcz
KaSkB20iww4GltUemxDgbrY8gPS2HR5ZMjoMfyT74nfrIC8QzCQ2f1Ow+A7MLQAR3KgRJzOz8/GK
01k5zoP/GrkR3lLIf6fLdJC2u9MXsP6dIfA2PWhbwPCyCeZJpxx9C8tF0CG6kLrii8VnsBOxa4TO
nOtUS90soU34gTB8ySOzB+hIE+h6LGthwLXfdLX0dh0l9HpjBbJ4qQETNuA2DBOHMzYxOOqb/YIy
1C8wmGQdJ/4AfDVob/Q3iRBPuFFC7nxvAP4ukqAZm7joUMSIrfswH/kpL5nj065Jz2aShPsZyC26
tLrMor6TIZFLpHrCwDaIbCrPDWET5473Jp95J+iLQfuTHL0uKMWyUyjhrKdJ57L2t+rPfJHp8zMg
wHwINdgQ3ncAW8DmPyqn/NBn26LrCa/7sdg1G9G3f+Wd4g9jvUN+Uxs1BB7A/YwiwE/YzGcy34Nd
o51K1aCYIbVsj0krsJ42tJCyIUaxhrGT/hsNpCUW6N4gFKypnFG3mBZSuFnMdtM7Aa//cuIivVTw
9UA7HaRkmj8mLTasDdQE6QOg3KoQ1/35syYvuGZ/rWzH69Jb5XKmHH8/CdjDbpkauka6qUvkYVjJ
CYcbYpH/Qcpkevxx1rPatJ2e9a0VH6uYo+JP9MzMYmfBMoB0WNH8zDcGKWbfCLppyWbeVG8dD80y
vdw1LdSfrDZNADLHfkS9JmHOP6FBRFGVXIg2lTJbyMqjE8C5cwlBezyDctERAH5mhgKjwNsdeDU2
8MVKbEBkZu29tN2LgpAL8iZETdXH1kBIWTrP0+oOyAfzDyO4vPVMaS1NMd7oKPN3SSJhpYyBh6M3
2FOzlQruqWT6xWQ+82SMV6kRU6nI28slGEF5HN0m6eTPo6MltfhLwGMocM5VKi653FxSSDb9P0E/
96qySxfAlWsZobr0FQjyYMhU3PQV78m7Y/yRcnl0GNKIr+UEUR7T98f0+R5oAyk1lcYgOyQC0PWW
mgnpAHiZZzodVOyv39RwSF7dcQOr1OHAbKA/fLPrGEys4z8Qg/xszeOFd9INiCuCPbwgQ1Qu7Y5o
L0AGctThreZnyLe7ApQKzTKD2gOtNI+Wh2VNJjSqX5kwCHAFaHbXRCuAQtKfYFUXEcOxGvsX8CGt
76kqR11HCCZaUUu/SEUzsBAOvA4AbNK4f9WDPojty52OAeExACevorXviUDzg87ppM5OFKovW7Pc
8T1D8t2s/3n0yNV69xPTUXLDftlXaOC6yAB8ysV4y6VaH8+CakZdJl+mXbAIAUkkJPcplFvKPDIC
rjXONxQHJDCsXc2zZaPIWFqVA24Hs9+O7ZajcyxonNfZyb00HM4E3cVOgaHydwjKvs9FyncSCCwh
pPZx2fYG6LKhSG7BWwMIdhgu249AIFm6pbuKtKGpKw0EL8E19v7M+1rOrprKRpqql/I87fOx5gsO
kfrJTzVbJjx59g5KSJZKCrxo9YbRHs7UmdP07gwZCwE6NwDyUHj4eiLVpM1ryqIpmiOezIZoPyJY
asNu3V2rdYYmeNrsLRZuEyHFGaueIIgGXMcGvYf4UYgf6DOiIGh6aNdH4rA3YRZMzGcExCjjD+In
EVjVc3QM5VB30gnH25xTt503yAcuT3gBgMeUIXZiVR/iCbI1ls5YnF6RB6f+rjGE+/LuZ/hqGu3s
GkTIaj1qnTXmTLwWSw2qCkkzDVbHzUHtGly1lrsZpxLyXSCUvGaRonpuMWToRmDLehOs1MkJ7Yzn
xGwhE28Ab3B9qKcQ6lbL96Lx8hjvrBmobn0t3B8c2UdWVb4U9dwAUN9YsgP9HF8xHsI1Ne4jNQZZ
FwYWQJGKzNBcRoNt7tlg29Fs/6Pay5egeR25MX2Uzjya00Q8ly+aT20AYBspoInYVjkJsNzkAcJW
zZslBBO4TsEhcYy1VkEw0MVTAtbSyZ8pzwPaBygZw0AVfFJj+rDa8aDqowKIlBxuNfQLGyqq7uLn
MLuxUuU8RPDQDDUgfcMAFknws3I+wkszDlSU1Q9jX+jy0EqEx76Oj/+bNSbRrYCkRcr9Xp+okb6k
EsVDSnc7CwpHh5UwvZsci7dukcov10sGNovz9SqrDo1wavyduW7HTCS1lIUf4Gqf9ZLKxei/uKw4
cC2gkvZxocbyQZqWpQSHJlXq+aDANTjIHJSX2JRdB1x9Sod7p6RVf/VZH6jy8itTSVADIf2kriGl
+6nBQcmZO/1dUpuJXuaaIteAPvyKCFVPwUwFBpqvxjBaPJNfVsmtNdl+hmroXh9jy/5osmwa6eKJ
PQHPVegzFm3yK6zB9fpoJkJEkcXjccZ9Njf9r2loqVpevPs9ED0Cm7uUxooI52ieQVbuVXhDaqs2
UKyaQFGBqu8uE1ivclxMUUc0aGArBhU6yvYcK9PcYYn3q1EqpWHqrUsHaaRTQI/6GY8RTK3lYEBx
dY31OTLFaZ9AukyYF3C5pne7CgW2iZma0Ge7dE6e9FF0BaUyo2M84H8M0czIdLNj+OkvJ+JpIrry
1EwKHIytDljrb294cdHVTPxWWKhn6eiHKUEkSKUJo/JUNxiSmYjyAD767yTLpnj3+tqrt1ZbDfTw
33DsK5mvl9o2SNWnIv27a9S9cBSS6uCb3531HjMlww62zfSRVTKpTAPaPvKZO74VaIHDrsW7asRJ
ES+YTc0hwK+IiikHt4Tok/ZY7770fMUjS9CrvLO2AMF5vOrzcQB73VluhXuovhaGXarpK6J53MU3
147C/n9ezTiRWwikH4MNsKotL2XZpIt///93FxN+Hrb9ZC/Poi9/l/ElO5KVjRIAKUUCpGYsO8Gk
ETIW+WxppwjB+iHUtv2tyHX9utoDwpDc/qQkV2XDiLR++jr1JbjQ1PvTM9AFIPTk5RdIKMZD/Sav
RmzoH8xndSeQD8Ovg8V8UPBP3STH8aSycn9m1BwSnyqjg/YDV7/T8dl5J4KXLZKgVBZyn3OI5fXp
igR5KEweVDQDFG7yCaTUzBxu+kGE+OFK1x04DpEcFAxPnn6zoFFsaGTifmLohCsCeiD26s6UHBPa
hG1hhtFHwnTL36LputwEGIzohKlgMthTEnMnS6SGXSayl/HgRnHTex6c0T97FVM0a7ZwlWLOGoxL
bnzTlYDbwIU4z3TSu2fYNfCd8FiOkFayTlR++frp1tXWYax5IzmTW6QTmC5DVw/odhNBY+kOGrme
WUfstqs2BEDaSLWugmXcyVf/jVsNDH8QuW4VFwFRQnFPwWhnhN+/C65TzNoZLPsyx+1k6a3XaKpo
7lDTcp0EPkgkyLH7h+wkJOw/JhivqVl+xIubk+PPaB53APhXN2tAV/5ork227oZueR+vVectLCk0
N3A8fhrw2/NWIKhNiuw1P+wK40/v/aGDlf5pdrNaNyGwklmB1FTcZNxwNEiHNi46GapjvF34nXSc
ZXI80eEn+FhglyKQ15R4KGVeX1D3N2SspYFfdeNWGMKFd+Zm/P2OFZAeBTqsXQ4xp0mpoNZ3ryzy
KUcvKCsicSmc6Knq14175FzqfkEVNpQoqI84PMsP2jhhWHeW4cBHL+nyqXwJ660JVdoBI4/z6fLU
mv8zEBaXjwFPAHAmPARmePjrzewtjffCX40ZGQywQKjN6F3JvRcR5bAtu5SRmA9ovg/+uzvKPR3Y
vVW65sn4eme6H2ZcPn+JSH/qZrQJQIvz7eyl7k0UvYxqsxh4iNP0tRW4bkVhKozvYauRvoTcKuvz
XXifg+HudirDQmwp3y5jBwNeBGQwRLCfdL6qGgLuph3gbKpq5yUBHEeAdBDokaoOqDd+MpqRQNZ7
gjlL8h8tj5qc43vQjiWlAF3O65F8QjdwgFaLwTZ+PUQMjUzOV6CsBOcTKkNay/VUJnif03OrLoU1
//Vw0L6jw8McfQnSbPxfMENArjVenISE804uC4ToKjtbfHRkZT8j7hpGvnBYGdd4Hj0bgGI1472v
1eZMal/Xxks3RxDH9YUf9Lc1uPqj0KycAYPdAMgmh7l8Xa84tcWMG6idjVdOYlFUhUl1p91t+sht
s//oQKvElSFCwz/qDxVRvEGhbPy/AQ1RblT1oKTj5dklaXbDQq8vMFweJj69if7YETFytthWNR4f
3ucrEO1B8g/NgGnhj9AlOMwr6ogMThSzgTDBipWLOJn/vglFW53fysLZT1cLzGyMKfPTKTh+BEmz
ooXSPr2X1PXiMm6KLOQatuxRTz9DVjO9IEOwRk6380us4/WY2DR4zVhmhaoB2Zs9oxcP89dMDWsf
gTXiPKKriSQRiGqWuGR5E894hVnYBe5y2SfAnWUMr62rjyvXbVzRAYRXLsmIASOGJAk0FhhT7x0G
s6Tl3Dlm0jEwh1PtwdKZVLuB78ZaI9J0zqdZn/ZgBDOY6EtN/MG6y2IICCCbgd8e8dvBVKCuTg9u
gu1FtQsWvvnS32iMf7+DSSXnFlKXdhp5bqt2qbBZdzk2b2CrQ1llZWBkNLkqUI00vphOcmU1CljK
7mFXLe3LcQuwS/1+ZocRLGK6lp3G9494v282ACHDYa6QR93fpVCx6YVhHJstbaon5ST4aIujhjXU
CV0tqjOFRJsd156h8IWB1owGyZgvMeIi3BJiDRjD5bA5jVYQadiXXwAYmWJphKOsPM6TMc0O5+y0
szyUDixzRzFiL4nQnkKfwbpGeNz9mF9KccfOz3/LQGxSw9NgCPaTjV6AbDWMdOsxXnYOA/H98ma1
GEApaQVwyAXbYCZOsvjwqvOIecu642dvYKkISTVDkjKF1lGx1Dt8khGHdenRyRe8+rCmnOKENwct
ikyyp6JxEISfSUU/lUMLbgo/ViFHEk29kxHBxjWMrqUViK7hA78yjGkuZj3NsAAsmCt8ABULWBg4
goPWgStijoLFxXs7oRaG6kj0YUcfRBLX4dRSisF3LqABiNbm9xqYbpICZY4jTjmsVd7NqOR2VtKQ
Cqj8hIjmtsepeLOg9KMvFlgJIuhwM+LRWP0xSj8rV0zxjzL2+L58VGeFO4euJuA5BsZbJzelAPOH
fD/dw1kVhjGm4FnvpswzfZMJbKC51AKheDM9d732hToPgBSyeMOfYYlcifmSkD6m4odF3t6SiwmB
bPUxIE4ae9dJuPwkevem1MVSN4j3H6x3E5IGnAt0bQqyWOlmXffvZmuaVfSRwzIefXW0P42GNFSr
h4NTTKPnJU6aLNPObknsGgSEiemxIBvzuUvj+70OCcm1QV4GNqVXHFH8P32kNNzJ3P+rCYsRHx75
yEtTu7XOWoy5clNfxFvyIwNhIjgBvvfcqaNrUddlk8is3EELo9RzdHdX6Fnm9uhy2c1Skx3Spvy9
9eXn7Ahh9o1RpuqUh7CgliWUhfh4g1yByopR8V0pjE56oSohff7sPQEWOhbzdjT9J4nyv1cG55qk
hPzpcXO5+YVdswCDvSt/jWYFVG/bbPwmm9aXhImWldNARi4p94tvbrvpHPiVsgqYhbom7Nx9nJ1E
yxI19an0KputsjBjXM5+LsM63F+jnC+kiDpXDH2LJsMsMeCM5esai/hsFz/RQI/RE9nDSjQ/L3xw
PB6+XiRuLQSU3+6fe5szWfUHmQ7cibkuC3YsPCqd/DVkS6smj7ADvpU/7mUQzwo+HGJcnyzJvZqb
GcpMlSjBXUTCyc+vL2eGGS0gqWpsCUWdLM73+W3YIYasdNP+KUo1VUNvgOSj342ruCJqt8VF99sF
n9DL09VW9lCOUt6f5JhEze3YGHdxnvfx95OYn1A1cFrq4mVWV3h0mz3bzi0Q1yR44ug+wYBvNkAk
kvthlWCBob2qOhekUoOb50CHvGcIkgpFEUeHA3OLSW5sEnUtsfLMVr4nAibVNJEHa7//+kq2ydNG
rRy0qPS98tm7QPxkTavWmcIM4z3B3RXPqqSRzpEW5/CcU9QDtFh3N2zyilGZQHtJJtFl9nVx9tFP
UMb5SI1WEuumC4+M1VxaAPi42HaynTNOXAaI4WJ2ATCv7n/3dus1bXtk51T8kSwk+C2W6ygmulZL
p2Cb4Inml39M8LJbXKuu+mysixqsJNVknAtbOOMXyuFTojdMg5UicoXvGyV97xMsFfp+lClbeDMz
r0HQvBtYL5O9fDbhpBzRsjLGrmFOuYVIUoCxMSx3UniW+z4aDs0i0Bmy4rSp2pSBWybzmwXAQQnM
qGyZQrLNQB3qrQ41oODs0b54fASNRwvksndxgxQHB82APywEghxCJgtQiUqyQhTreh71T4KLbIDH
CL8QLDuRz08U8zt57QZLFs8IIFFi8p454EsInydWAGi0S2IJDmIKRmZqqnOxr2dIKMnFjDz635FA
S2o6CAUUpBmvE8VU9eQOBkWDf1B6E1AFlP3aJOFSgZxrN7K0awaxXcMmnCMph23I/c3gdWdpjUbE
/1twLa3WxKuC32T/ZNMg3w/wp0zf/rMEGwpNdelo00w2dlqHP6Yhr30lGlH5SOtVpccm7j0zJQFd
6gag3/ys1wZS9FfeJw81dkq2fTJmqX7m47g8ZHns391WCdNQiu52bo6NIcdxyldYrUszDXhECSE6
jSyDfhBSb6NPXy/d1v/4EpNvZWIyMB902htCkCaLq/BZF2CrO7vFiurJzRq7xIongSPMLsOkH/R3
sA5npp0MS7GR0zt3ciZE7ru+3zC8AkagFnbxfFtpnhKDScGbHfOZE+0upiC8nYnDKm2SwdetvK7m
QXBzR+BuMv2k4/t2Ia4kaybX1MfAeZpUUM95fhUGv0wbOsWntmhFclCJ37h+qNJ8ZmXMUa2FCcZG
pSQt54w4162rkAtguC0MmmkY5LRSPB3VaskLOdio6/v941tPWByf6TBksOnWp8FjwGNri+Rh/Dl8
0XOaJkBYHIelnWt53ywA3ZVX3eUL+ze8xhQ9Gwn36mPyg3uzWq6SLwUJcsU5Rmy59GmmOBROziS4
9kcVXGJ7K0SzOI3N31TIul12q9uKnyKHnnVm+do9c3vnK3rn8AjPCq7Dacdc2VGkcIhJ18ZA610I
XKpyLo+9XCJbEHtHu+5akzrLpg6WwKLR3kezNZ0Oj0z7wl8wyfiYEE/J5Mqp42/Di+3oOL/7U0WT
8aQu6TaJKZsk7/Jtwgyn0teeApSsU1diZ2j53djb4DOzWW9oyt/nHbZYP8cc5f1T/loyryW/xJk6
cymTzXHuhh6dghzBZxTT51cYgDa9y7j1J9SxJf41pF0XKRkSg1XUh9eIOMCMYNVvST/U/x1oU80Y
RyQCBPc3IkP/akOUGO5SqFN+LM70wILwhitCKGrnCWSG4MDUqghSn/oajP5iUPcmK4PpEAB7FJ/R
b9+bz1vzhuFvdIcdOXSeaslRiX3st5YuT4TjvAbIwvkDDKRlwHKIDcQRC15du7RwGtXLATqr3/F4
IjYWbH4OzAUROMHZ56xlxJtxwILyA5836YznYSKuEHBz/fZ8QQdR2wjBeKSxgSyXd9FpyzOuoQrp
4sREHt9XKxf5ZMLqjjoFht2MEi5DXnvo2pEw052uDAudJu1ma7ScU68oht/ONanWmTy6kEeBBXq/
iWgdDFKTI9GZYnHuOT6+agOBGZEEI5WquM8/Tk/2U0787ZPRrywOKp6fBH12n45DvxvmphpSecLN
VhIZUVADXYXQGk2Iayn2ueD/lwerdjhS3bcIM24FTufG3m2iIyWlp25YbSX7K1zBfTfyqxsI+Y7i
9frSzKPRtCODjLfN+sPhIe8P4okTheXn46ci9uRLkwHmzmniILW4K59WBHCia3annwhtHwT1/Yro
1b5WD9UD1KjpdMCasmm+j1uGHjfLTSdZHgZPfGRHT890kd9QUtEDJroFkAaf+AkL9ye9Lh58nA0B
DyyAxekgTFa4MvCgh9yF4TH1pD8EnubZKy1sFAd5LKhPA38RJG8YAqw2X27oSCNuStq4clpK38gs
XG/NNhjbvqro4g6eOHZg1I6K+E+65Fu2eK0hMPXvoLagQ8Qv6xsDockdLju041JshBCMaoC5Gv+f
ccggH0jF9xTQoUfkEcIEpz9PaRn2HXQdLMBXvv3qSrxdAnITVh2bikj1P8oPaZLia5Vhjy7ALq5W
ChY/9evM05ItkTne7RWpETZp2F8kJfgvDYxQCbmibIAXAxtqhJKthQ4gsY2i8Inf1z+5I+uH/tJM
kKaF66fKHyQRw8W+OVzP54xZmN8XmM35HY853A1Z1rnXlawmKMngrJkS5bCOXCHBcQuotzUkV9jy
E0zzr5JNWtWgm/rLxCa4StwB9rw5pVnfAzcVDwJ/ZEDDR7YnC544x89KICjxWRedrdtGcavezZ+b
j6maheht///7JQxv4mpz0/nNDTlqvRDMKHazs5tS/O862iI8X/eP8bTDfWb1nIdHCm41J4gi+jg5
KJEisvKrKeugUFu70GCZXtrhVqBW7sHiKv55MsxXSq7UM7FFg3mqCl7pG8yeDj2p4C6ssF4RSEqd
9QPkznULr10NSA3J3JGRolwfmT8SiIM+zZs/n4i3HJNnE8ZTQzXT5Qkb3QdIAaUg2/ZFEzVN0XLe
Na7H02Z8TMGtKE0+ZxlXUvlCPnu15YFA5HIetgbk9j9NZvJl/I9+u7MIZtKuQgBpm6KYvwHW4tQv
TCdoaOcBgewDCcrtjEpYxj3GaiWsVYoVuvD9Jls49rXAEI18QP80ya6s00jBpY12ossR8Q8GVhrG
nQ1XgkrjGJbK0CyeNXMU7gvw6d+PPUkmLtitYQCpHNT28FqEeCu6L/zxQEv2rkQmS4qkIa9/W8ol
uigc3J1JXOOFqnFbj1DCt3ApFVUq+z99xgArO5M8FljWbvaiEbAZBUEpzC0Tps077QiVkp/RfZ9r
vygYeXd+GFY96fru8dQIxgegJLjT+BoRzYmbul8JS8KKJQIzI7gGvKATJG8KrTV6YIWWjds7zd26
mCU/ZRRZYnJmowPes2cbof1TiRdgNpCP7ZRge1Z0fjVgRPaAaNJ3+fY5WGl49+nejn/Az97YYrkq
f9bJQ8xILCvfJiGWvSH70Qi0HOcYiYDbIx9dfnzkGC5n0xB4bE931cdUDuBJKXhJiOld7dstleao
JnJjzdyIjhwKWWh7TjT8T+e0H5Pc3G/vWwDRxMctXcZLj6LgRkYo0yRqPM4HBM7aMdSV01DkYGtB
RQN9IUUYK9+mqR5vxfVre2b9WaOrR3LjOJ0cwcLjfaL55DLKomxp3QrvgTtIUF+n+EUII9wPrYBQ
YhE5G2SyBdwqFA9Z5fidzZfrHAlgd14MZ/8vxbKw86thznIdXDJId9X6ZeoyfOL3NL3l2gbXSKkQ
m2EQNtac5JEWcokKcO2K9IrH6j8f5bdm6Z2rSf3Hxz0Iqc1Dz4RrfxhMoG/ozwu4LZL24CVF5P+1
k/0hLfmsTUcbJHzvaBxn5G+gW1vjjvRAuhFILTxLB3uJFh8r4i2H/IzyB2AGIA96DzhYRUstoCvv
tuAQhKeH+yDqD5Me/3d0e8GmEglSWZa00fDnvsAo42PX63Pk6YpPWn30RjnY+pIFxWYkNueplOjV
P9FUnJvrGDhHf3+LM8xfSiuFOM6II+iqk6tmXiBufJ9hFXHUKO1oEzECI0N80uI1/+giG/5agTDO
jezCOXu4GAC+0implzU/+mac2CmqkMwAphIxWHBN3iTefI4K7Wb8zC5capTdHEcSP9TpUkvthccD
qpgcjNie0m+JqWkEsv5ClVa+r15KvM3j8pRa94t2NU5GPB2GRopuLpEgjWXUmXp/GLNTHP6e9IN1
Gku4FXmUn4DqTQe44Q2tHK4mh0bUTT1gdEdiehmPeQRgqEfuid3oOe5y3qNCRDMrl2JRJMLTUzhf
FTD9B8ODe7v/Ep63P0B2SufrIUWgHTh5TkCImqD5T7pnpa8n2QpwVEnNX+Uclh/RKSm9RI0eGU53
+Ep0kReEEvlM0+ovgYE1MlTHSkeJEYiLhq6rpiuF+4IFiG0dgIDSC7PfETjKxnoM0IgVByDtWvKr
5SczQim3hexSIX3DrSJJ3cvB96WxwFQ23t48VLyXwUNWbzv2qEx7bYG91HYVhKcfZyZafeNEo+zK
Fzj6nNLDbQTRk5OWR+Zkc+Fu0h5/0ehDi19vQIPj21nxAW1ky8sM+mfMqSqBw1JQ4v3khwsAjmZ9
XHqdmhqN1KD4NJkY2gUR13sPP8EC91k5Yj2hqZAuy8FRkKcExTI01XN2gXWf3HofPyQlGx9J52od
WKPnNUwOUYJvZpFEU4rWf3NvcSSkvN657VjCfG0zhJbvmx2rLkG/QLSZGgMFXFn3+K7Mt9iC0eI2
vn+zywTBBnspNvA8Rn1he3JhBbQcvJi5C1etQBerXky4B+je89AZdpAyip+chU2Gxlx/i4BSQzCa
0rqbBVmSBuHhohcJNK0XvJED9zAPInxgP1saugJEtauPer+F2xxW0RUFXXWFIy2WqZ34G3Tv+3TN
Y0csFW7Xj3tJ9WSPnmmsmo+2exxL9miPlwXOZPaZJjQAJoQzkriK0ZM/qP5Sgck59wQHO6fsgnHx
8rXkzT4lbFPCEHQ+oZgFWXLooRBBNwQVMifJotCyrKSaPclQ6fGh2bO9olueVIXvWhLcOwX3jMgI
PpBzw8Z+1VXj/8FkVW6M+HfR41Kz+jnjAsS9YMDD+h4NYCoNqO3Wyyj5AE2Jw5m8mUJcSjrksMOd
JpWgPXSww5cFhfd11Icx3omxNYq0wDNRRxBHMtiTyoA4ZMpNhyn9+Afe2Kcwplq7/7yIiwrSX2vY
9WEGYwVDx4t0unQ9o3i8bZCcfs1wP/0yPFgPdaWUpfkCZa9qlLb73RZFMTNIOv5yxPnUXsBFngm+
kTWm7OdNSxu4YxGGMs0WdHJuTe845m9odU7BSLdzyMu/XXQJSYUn7AUajW8+rIx+jo3lbiPn7LWP
Rpb0d92E7WA0TG6dYG3IcX4G/BeUug6e3R88SWOiPDcDwQy25/vXRFvu7zosArkSpRwpfYWBamxc
KM8AYu+vzK3eHtYGn8k0YYiD1QJCJb+a+QoYO4xQQy1TXl0mHiaf+lGf/xwiCkzizzMJX/EwFJuQ
msIhJtJS+J/2FQtxi2QMPK43eDb3r8UNt5qsr7qX1wb6j9cAq4AOerFh08L2oIHElOmABrAe9BjO
P7tb1lDa5aeGN6b37nvWTBFKKRMug8X2ZFe52Q4P55HOolxCONhGBbHvDDr437Q3ZQgQbrkrXenG
OfoP6Jf8XjxD9+Ju79yociWGEzH+DZ/7c26tFDOcnBoTg7pxlWtzFfBE/tu9wKK/96gsuWN3DXVJ
Py/cSKRGyO49teZizAughwsMzUN5pb6TO6oEllkdLKnlx4pcAPpvRndXiEs/aMkNe7+Ss4rw0PAz
ghoRcxk0AQxFB7wqkNPs4u7Ps4K47LL+/JvrtwZQbmY0BB45tzke+tHKXjoWayEWYgQ3IsS9HaaA
Y+sxAAuuu9F0Y1l/TTN+3IdLsjL0x+CagHwJQMgUKWzCuBf7y8vrcBOeiRLnR1rKHHuRtqHyRY7G
p7KIm9lGRI8spISn4vq4aq6GRC/zzmDamg5s4uZjDLUrad/8f+7uSm9xYUEU+AMxM5/5TpKaGYcK
RYfLE3UnX6165iTvdCcW/pMCTv1v5tppj7AsnwgrWRp1CpZfrnm7LUFQmFDO3+D2yuI27WmoDEfd
EW+tiqK6hcYIqniCYJoE0RHQ9rEebzOiMpkt1R0YtPrOZGcBuOWEWPYJlofQcQ/MD6vxHVPNGy3+
PTn4fAX2kCkEnvqvvuEeahNxXGvdF8jzbazhTbnqpQPMAO+8vHxHY38IKxYeOaGLZp9hbzoy8WoU
1fmDYtFromirMADKNbd6/T5D3PMIVskXnK71LtpHIEkf1Ea9ec6Ih85RB63HE8J3O5BiwUUT6YL9
m42tfcpfxpO34CASozhTuJCUaXu//ebc+zBOTihZxoymX5VsWYzmyxr7UhJ2mLTkKH3B7/C17oAJ
Czv2aLlnYpBzWWQyszyNG6UUMNU5UsroxwUFr7oKAblx3XLpboLcy/5lngBqwXjmiesP2/joZkSt
BdUDLZadCKFpGn039nuaiAuErDExz0Sl0oaKAsF+PUNUTIIZ1RGrrnjkECAVBZN4hGFijHxHTSe5
GXIAegUOfZr9LXhlUzPy2DcYgzrwjpnsYtBIJAl1sRepVJz1ECCHvmTusMgqgChJphe8mhyU31F6
QicwqDXU4KlgPVXyDjq52U8YOvRlTjeYI7wQmc5kGXmUThgTCN+wxIKcn1tiGWkLYXu3nlEawxTv
KBl2s9B0vTFPjr4DaaaZW3SYhPF7apcnk7+ix0OQDHvEuDNYIRIrZEWb1gqZt4CULqybRt0Yqpft
F5ML3UJkV4b3KOASu8/TQUadrRZXoB66x5qqvnQnsJuYFTDjklWe3Sc/cqx6rc5ixafLT4ye15V4
FoEw2FCWRv/RQc4on/grgRkEcFKiB5k2EfquNhUba0iFfNbom3TaPyniXbdSN6mpdE3IvG0lLdDJ
xpg+0TVn3kq/BoNkgqEr12tM24jeSvQilhMjdTNHwpM+9ck5lppqI89YhiyB2yNo//s0pGlwE+6c
qj/mwor5oiGaci1Hieyye6IJXvUgPp+jS6IAY5TaVjSiknbunamsJDytDVnYT7jasLjNvp+r/3jc
mcAoRsarUHDtgLcx89F1IAHlBBgE9Njisz8KBygll+VtZeiMtIQal8d/AGh0Xu9hbFef4qP1fEBf
fnFPVEg7Hyu44hmaN/CDv5BLMzrGdVqWvG2AR9DpDgEnLXML0NYUDlXOnGi0Gmsp7dXjVzQ6ShHd
Nlq43yQRnHAwv5zMFmSQdYxVpg0P5qa7+GDpw1ADCwthgedukE0P6rxUkY4TedDyBAX5r1gBqV+V
Bm//8iiaMdufLXt/JgneoBZNFbLnt5a7pupqriLKjkT/gYZUyGIkwfFaws+MGIUaIxzD8PijwyDx
fcmNuGgQh8DfuZqCLVBSC7B2yfhOxRn/gPjdzRzqpzlmQGPPgy/Indp+T/LAfnqBfVfnUXp/Twj4
+gA1TiOjwGc9ciQmhKSW8N1to2tWyQk84GSA93ZlCG5ZkAykIU+MaIJTfAmQcnwB2AiIE77QhEJr
hapx5JOY9dtJNx12Ba6p5NDnMq9AicmmyIkVtHYV1VdMm1vnnZDvW1NfsiO44I2s3afYyoAoYXFh
quKxNtmn43COaoaJoTko10a/94SLSe8M3PJfI4AOQgT5b9j5pkzODP/LGu9pii9VRli12bq67ZHD
GyxcBWCBv7+V/1366GR5XL5wpqtJlnMIg4ffeF+huKdPLAQ2niWRdnoYN62ReX/LGD1TILiPDKts
W+vRe7HulpqRgUuwgWoPKjAdgeX34L7BAHBTK8xK4ZoeyIm/IRFjOwGEadbUzAxusNeJCU2v/EqZ
EepgpDTl25sVyCr0QNzYIE+KftPcuniNzpXDwYSfMjmT3Kv4UIRx0gGHTnIZpoS8pJRlLlmiT801
LDIcLaYj47s1AEn0fjBPV7foO78vz98mhzXMEySu21hZQX670ph/f330vcMKqUZLgEQbY2HRjsxK
PsUE+wi7rJ3aDQOD6cO7yXK7A1OjviH3LiAkphuRhLY09kfYWlcmTwxEfkOufB6ItxEp8KljRsoq
Ijc+UcjNFYY2c9fOBNCPHYEf2mz8115cor/b1eksi/bODbNveicAJ9HnTan2hDPh6jGKmv4nZi1o
AX3QfEHKxkSO7js4+lZQ9rRAM8pjhaKdYMCEMqrr2q0Xxm0w6OF6WYm+QkohoQCFWFsQFl1XMNnD
CdiCtBjcULJDFSAMJDGmGVcmpO4NEuKBIw+ADm4IRNwXWNFyBufL2rlqC5rVCun5/Aqtu5A7ykNS
8TqlmrAfBuuMJJpvVLtMC2WyLUVY/00F/GtEvB7LzukNeYferxJYEES/N9gyoLI/dSTYYMcsSkng
BPtAdtvwTxJh1aELiHlS4xgy2/YQr+zzEZZ9LOhLGRFdZOY0tb+gFj13OzcoAhecCyrLl58741fJ
BRCyO2YzDvNxnyY1G7d9/hvHjOa4Ud+zL0D5heusLw5Vu/U3/A5FfG7MN5ndfOyrjLarJlAVsoLq
FUU0jqCHu3jfmGLDGyTOMk3HN5X7nCKdPxCZJUPutuzPdaXLRAm9hXhFqSATeVOaNhuQ3QoEvRqu
Qf45htWOzLPsoA9ZJ0q6h0oMbEuSnEbcb5tz/2Rb6Yc00RIIU9/6cAY9y0oRbw/+SZvA9dbz5cn7
w8skMaGieIrDHbvyTAhVQGhZKl4RaPuJMW6c4tEqIVVddIK2BNJFFAUAGVVdKLZIh70NnJq8nX/L
ob+IU63TWUsbo4y2HTtkVTSeOxu33Tp3a6AVHI8hvFKL761R+F70ZixSQfdLaYSj6uZRHGv1DjMA
bd4rYDS5McBK4YIYYibIjQoQg3zcMVcNd1iXX1bGdKVCh+l1dwiYDPWUpSsbZWyz7b7k+jBJG107
X20rZ92BC3nCY62YykUk9AQO+4S+aMY4mvpopP/Y5rDVqAwLVm3m+o3Sh3eDiTNPwe1LftgHy7aI
fLryZtd17B78CMNVk5NGa/WaiJHtEkdsOxOes5v5Jk1ZsmNWXPNZ5Fij9It9oE/LTWyDW4jzztWH
J4Gi83qhUayG1Y5227xJo+Dg26TjdBP1x0NC/qw34rlBPT2TyzzDHgxY5wfyq33CbJls7YmMoEho
swTMcVO3bdn8bH0pOPgmQFohoOlOrPdVXzp51CsNCw93gXMXq+F/hG8+9lGBansv3zs6QUhcde28
5mwnlc73Rlp97q5KlJx/16y7XaL5y27pa065bqga/EOj3G4t064AlPLD5IYj08jOMKw+YqfU2SaN
5ZI8FODc0ese2bsoL5eFF3dBfTykEnaump9X5iCmadfFb87BzYGIhUwem7PlHo0Snp/4S/H7un5R
22EztMXeRc/5OorOArzAm7y4a08SHfTZnqqqWDuEFBaKxDYGBFAu22Yr/9no+4WMSmiFuTFWP9QP
faDShlPOUYWQEzH2dLFSZLinw0cQ+/Z3FafWhpqZNsGmShHK2V/Z5Wzbbrmm8X9EJ7yVdHK9kYnw
Vm83RNDi/RHTw5LDvDoukZ4dj+2hrRCoKwIftUT1442WBS46R0WK77mZiIOPCNzXrbJej2YHQIsd
ELf4zPEJvAwVQtR5E4sL1CD5inDqyfP4MjCk3jlTqzHrctlxX5Iem+t4LmdNRrKWE6xY7U2F4tPP
sMEXJBpn6b6d6iEaTJ8dsI9FzpLRgUUyhgqVxAJN7k9E2xbr/qRRYFJhZEpyv7GNbBS3Pg2Xf1X5
l/48RKnz0XfkPYtT6CYppGnRXQlZeR7NIciZTnMaAWKe6NrfYGAqqdGwuzb166dJ/GtynvYyGpvP
BkabS2y/jKuOid5IxajkEJLlq/lME56XsBhy4nPoMXdEIWzXTAXPD7y2Yqi2bMiBGmmG5tsZJt9M
CrJxLLy+HF3mO/kjzzvXVF16iRvRWbBeDFyDUaumdxb5KNlTVVG7GIf5NLTYnoFk1+fclT3YEw+Z
EGMh7PwaPpQvpZ65+8/DHr4CV/2n0vESz3lXGDr1ydsXw9YJA17DKbHOSB62iTJPtgkGtuZ6Hw/d
VMfy6S+F2UGgAgUfO278t4V8LeKbwpxuOi6SRWPhavLyDAJfyanOtnwLg6+GkZk9mGSNxmQsGsOA
U6UKDRtUG2sQs3cJ2PV+lkSJgLifeavlcuJfRYIG4BSy7vbAWAP6rkn4dFUtCIe6Mj1sT5HKc3hx
OZjUx5e2KhfrnOTk0j4MAw+JV4mLfhqYXN6brIVPdv1SsXsVvPL9u5ZIGVw6MXwXn8U1Q4HWDTcc
VmZqxEgMzsCAxeMw+RyQSeDVeSxu54E+eZhUOqCE3znUbf72qrvv5PKWYqNW/wzZK16fYf5i12ge
XrQVMe5u9vHExlUepQ79m8IWRIoNcq2rprc0hh9lY+zNcI2fh8vM2OLObYy4T9I0id7A1qOgY+ML
aFKvm1Bl6gzTZIiq5IqD8kAJ3WAVHEGYJgnQXHgfWS9tKXonW9hZCj+jjMvZvl5jOlKZZADkORzI
oLgl8Rj3evjI+vJwa3WWyNHky3RnTVqMPldFGDJwtVocijlfM+qkz2JOdEDGXTnH/I3q9lFbxxxR
5gcM0Y1AP+nomlQ9VigCj5EsvtL8hx0Vb2arAzp6031Ot7EpGieSQmTQkfQTkxdLEQ8xIQY3J6Jz
dFwVbBKJgKd8eT5pDuJNEiACyD/hfZuW3Rg7+X5EcQ4/V9vQOILl2YwYWjCTd9sshSPN9t/AbspP
GoXGskdepS6lLhno3t75Tok7KyBUe+MYHDGZd2TAldsLz+tl9wgJwglmfn+UV3/2KSdyggn69jdR
L2LZPnG3eZgydArYeEl9B0os9OEVGugrwRZ4NV0GY3O8cvK0w7EyKyELru+jsuA4PxxUMO/K57XT
7gjW7dY8UJR59bliF3I4a9pxrVrxxw9V/ypeF/8v7HmSvZjG24ozwQkxNNfUxFL3hyklNVW9QnhB
CFdzILC7xNHXWjzuKQciKQhiCfBWQgcG91cdRblsjGqs1gtZR7tBWPrTUuCPdbXXk+Aczj9BjIXD
dnlA58K5x6jsdXfiBfS2CbupvZDGdsDUul5cU1uVPGRgj6Zvhi8OR4Ql5wgEpSAQ+jC1VAMhX+Vf
xT2p8qIH+vy1fAaYkt3F6nBgm2+6yaAdmgvMCv9FrafeGo6G9z7WtRVE/ErA05Vz13k8yLx+FU1p
zgClM2XYypx5feD2SCOnALEYJbrt3kQBJMXsmjf34uQuCvGbM75F/Bh9Qx4C010ioqc3IxjayCmc
DVK5Ic9i/zDK0ZNSLs5fPyjNC+4BpM9qHjJhgMCGyNSOh/y7J8NNVUOrmQkzrErVhB56TbqryPAr
RbJ24XKE92Uyt6m+KbSWewz8ttqliaq+dVeFhYkukRocZqJA/5sBBUAlJXjEvO3kHpRPp+gmkTYp
mzeWEGdoEZlr+3J9v3xR6VndOcmrg0SpySVd/tIjT/P3dw+IXzHrKc3x+Yv9dAM78ednu7KpPzNf
Z5vyTsaqPPYuzrSbJmwkWvPNJ9nPj6YkihNobbAnA45BlELidFQvIb74gMnDH6lmODJilVz5n3ii
ZLlkjXT1pJqyaISMiXY+kAdYiuDff9Oh4YNnuWx/6iKt/eMD+IsMN5nVVUmrhJHBv2B2xP1naUmG
jYOGucMP3Fz4X9/OPGLEOB7I8jRgHxfUawhzqD3emIGNstMAhpvel9cOSPz7cnDWFLVxsbCnzFbn
utqkzJbqg3LGdYWTe7NOUexpDGOZ4eguvJxq3P7JjLcxXyk3S8shTqrkT5ASdX/lg1QClrdHr0N9
WmDCJzgz4hNgnCrWZ/m1YISCNztrdc6rx9xUcojkFrjrN3bdH9KQviLZWmuLl4QPpyZGCgdp3Ck3
vcNjledGb0eUrI1eezX8q6Gm0EJfMJnlYPpWrGnWzt58CVv0bgavCuAVJqcNhUiBsSI/QtMF5yDI
LobaMo1gfBDFAsb3G9w3UMbuWxLANY0m1zgwutbnOlMjzD43W5KA/EqZR2pcB4jrD1ywCSdaGGXR
DhLf6IaePYh/mwkaI7Sv3a3jmEkaqtOOoHvKyanLRikWH+/jPxU9yIGPAALX8yNv2l66DTW1ppL7
QFiNgq1Ufep5sKdd7JO5NcmXfNWMbxjKxN+ZvN022SJGTw5Q7OLr5ahDBe7+cSD0tI7yoS1ySWi9
xzQKwqzsEerApIgGizIOQwr83d9lCdtRYQD3cOT11BvM7EBVPnySRfR2VE4yO78y6IFSPkWGJhQB
BpvGl1f3rPc99iGEWgpvBWmRCIkBfVgfEjDyE9RKby3mtjFsZH6EIR0O4R2b4mUYcDuPpHlOGu8d
WXGkR3iw7Sr7v1Pr3ZndKC4iZvi98JFYcbByV7NbTGO0kynWDX/B9J1MDTxp99peDzuUymzla8+j
q/Vwv+h3gamlIUQF11Vw5b+L6h7fmk8yWiioEAI12RRPGteMtHJekm3lJGd3VmgqyykXyRUcA2zN
8/NiZu62MUsGcUHt2uZ/XzLEgdPLO1CkSPMzfl63MdnrJqBXoA2k9zRMGdexZtrd3fl8dbJYDo1E
B06ZyMs8CdCAWGHkezwW21JQXteyLcO/yHPSD+JiKIiKcGzgfKDm2QVgpytR3sPKjJ1C9AnQVwuj
U7a08UFz8UCy8VlBufGerwu+V0FA5fD83G++enmyCQ3huMVSUvLRzdH/JHVV3QyyZLs+qu+dd+m1
HjyMB9K+8uxjyYB7IMAK9JMYGWsl9G4RB1wjHB7vijFLt/DusjFnSAfpLUinjlfIuBDScoghFNZa
GyW2OwfcXuOJ250Qw6Ogg83utIV+egPiN226IhImZtOfKgYkwjJUcPGDrQRU3MUy/BOjDjaFHGWU
wuMMsw4vdPB0SUppUXNHRXHdgse9KugoO9tp1QBqc0mr+r0AdFK42GI566dQyrZPb+8kjkaLc2F6
12xSSffF/7DFl9D0+BXNGVvjQKtjo2MQvXFxXlAjbLEbPylIO/7WniE0RweLkVDMY4+G69jQnBpq
k8JUumE62uv7buxfighOVmBDpq6yv+nOM0VcEha1ZRx0FJWnzw6zejh2oziakptyRv9xH9MG1z/D
6JJfO2o7SKjxc+NeXDIYwW2+hq7fULCeiRYXEvt5JcISI/uP1vNqaB1mcVGBKONNuSiaaXOfBgtE
7bOXhktE7BKSaY6UjvN+3t2QMgpV+TTAnkqEXbzArJ9adX/Q60ZsXK3xIKD419b/ExX5FGDqQJRU
cElKyREOyUy5Zvcql7zL8gEX3eWQPHj7bO49YTwVgWJmnoUUaXTR3vsXNGCDLCtXt4Agm16HhdEo
QL1KDP/czOVxYarfVJycvKz/4ouUv8hLO1iVYixev6w9JevBKZ22fI1vaAfEQYa9F6yvANQgw0fz
hz3bUDEccCAoBNAiYpoUeFSNYl1wLaIiZtLpEslvvVLRAVFF1WVXJhEYVYVNVjTNZBtwnpHji4fF
OVO08S7Wz2zwXmVVRRgYWsJ5JgDaXnAlrrmZmADqOIjafayBhfCbG9k88dL81vl1BroUwqDewlHD
FIaoba6vlDiZPVN1fs1VlA2XpPjoKiKEPQexlrg/klkxwrQdwOc6mvjAm36TcX3ca6x5g2VXvPCv
IV6JdzrBbQB7JTEDfzGrQEnN97PX07MZWkqtrDpkoQTHp1+6soxtnIwOvSA2WwH4AK3zGxl8Eaoq
hwPfV+EALgWDG/dr3269eoW0BVcUh1QMigrKTgkmOBqrb8oGRgapDvpa9h8dmLhRsYdxYX+2w/QS
ahCXA+vs5/+2HMarAOgTdXhvE85Rlqr/xjvFdrs3gt18gwagXFDV7tH1O2spChddaRS9AN2NsRoO
Lwrfml+3kvEbifMVkgKygmxt2gff2hvhvaXiVyXAIhsnbUmF2Gs2kDaotPIeGEMkKTYT41xWh/hJ
28mVEXwlfwZFfawMJOgDNmUNUptdaqI3vBFsxwp0xucftPZ6rDkoKoe/Psx2Y2l2rxApQKkte+W4
iZj9n2TOX08pFHZG//OFNqzdCkUBMbvJ4VgCxhgc1t5YR5tJVQ5rYEPKcgyfD13H50/b4Z/V9VZw
Gzk/SGxnP7MBs0fl2TtMgmf1KmXkigtKfMWgEir2rcOx3P5q+os6GYZW7DWYGwDHv4AjIoI9g4cD
HUZoYC64bjYwaUAF6UfaQIPRjEIJULCz9grBIoTUwqUz3KUq6tWLtgt4E2Wyvn0mQ0Y982kHx0/n
2heYuLC/wY8BS74ZUPrHPwDybvd7J+atBP8p2xud6uVtjJrnuqIxalahKemMAq/U0Qnr2F09+YMo
jNzvne6XnWSod/WJimqNcRgbAKhALJw5GF1jLowv/AVxtiLAVcD+F0KTqqKeqOk1+/dJQJDAXGUF
gYlQpuomV/Vjr0kueJeOFRQMDUSVug7W6z5XURe4OKnC9xw3U6g41r1U7k02TtTjGBdlEI+0/xHG
IME+CzwdNYnHsbvPZ09YcOmK33jct4mSnnyvDpVvoLG8khr7/28xXswJJx77tpPj6TeyedZJE9IL
XXJXYcggZvML+gZLs4aCkkH+NSA9w26tLHUIZDeTSwiPx0QZkDFTyfymypnA5T2yeSaXtzexTnJm
SfXEJTWSvdy0DU4Zn3VxVLoNLm1NUh7mdN9fFIh0qxTNNrj9L92TrAOwcR4saD8YqeFrnMrDDJOI
oTlQbkFdxp3ROAzxtqp3jNC9Lv50tWO6USrU1JI5S4rHpK/BvRxVqBazXJiih90f2gnP1vS0x7tC
4O/RKJLn5jk+NlOp01DVxZB0pRHEwnZgXpsGgKbgDHiUwBG4uLXvY1QYJ/K9uqrtNhi4GBuWgHmD
IDk9db1OQ4e0Ua+o/w28K1o9wi/nP5nf9hCcgBqGcNmGxOoRRUwuqyYogxH/an2onlTCQR1C143Q
A7tDpk/fPQUK85hBqxk1F9S7TsbMZ+noZXouqFm62Lnlp61GcgVBCDsXseOLN8BofuPOMk8+8EfS
mDgp9HJJf1zwyAkTDjQjuyX5lWTNEiCS6z0Iyh7ywa0kCbpVz3AvxG3wBCALmdkrRaKXyF01ISq9
MEnR4/OpMNxLoUoaISIda7LXedEMi13SVvD133BYOt0Bzd/PTJGdOvcbmkRMniaRdpdSHEh9lzua
e6ZwIEGSSbpkmGPkiO8yxyFj3Iq83qdGojyRH53QeTbkJrvgN3p8mfoBpFlUvNHUkbGIfBzMrhiF
YdMYFS1KTGCLDgEymo6CKRP/S9avkGSTOs0wvVGDqNJK3cQBxMT/SmtzZ4Z69P8eZxbs/VUAK/VI
lbvm+wnfuEmHA6PtdenepL0VARwsM/2acBi+AScIF89ApfofyszgE7yxeY+87iVDnhpAYVNHsDXv
Mf5vhmNc1ks9JyR6aOOej0ksPtg+lAhEDgd4Yq9p0jTzh0DsIaYH+71TIK9ueokGVmIGGJbQQbyL
hakhmv43OiL/uABJpA2tnffCcU8BGAFzPxmXXb0I9cKsegaX8rYB3CY26Fnc/7nhiCpFYbs/01aO
wkYy0TsadA2XiaporcZUt5wW5beGYEfJgM5a/MLULNCAcRrEJ6oeCXl9gEcahy8r3qz/Pz7I2d6Z
OEo4EVU5kpPGgYlh0s1jUCltwOq7c4S728MPoOgUaK39o3f0NgC2CaZHTbtIWxHqBxQCIzfUfega
5CmfoYoc79vMOizhd8sgmXrZ10M1ipRav2016b04TQ/Axdll5tjGn01+emiSefeW4p0tnO06Ms3N
mupj9XFEbbIZU/SqYW/VlOUIgts53Ek+YLaoyRzkw2XuCwARIM5F1glzpU9rI5M+GH9RRkP4QSE4
7AlT2MKZ7DBcG51a4+6tAw0GUEDXgFAw6A0OxY795PXvWJWF4NAiPFT4sDdegDA7ehNL7wMjJtuf
nB4FFl60clOePCS31VhB967Umx4jZ00qttKjEK0xRvxnAk2WXsee3wbTwVkwiecrWoIefQpeYgbq
+1xJ27nb/yWxIRwl0LE1hBvehJ1+V1FsgdEG6fnoK1ri1Q+MdA0fIUlv2mrLG/JmfNwUh+WAiWx1
v5ADgAKnmynVMuhWbYW0u4F+CfYFNRbLnvievWJ6s/ANqO3xWQ5XpLVcbZYgW1730zr6U0bL00Iw
bRCbf6sWXtHI/Ccs7SuTmin1+VFoPH9hxccAj4YExEUwI6XHMhFpb0Qp/UcbsxwSsgcqmRJEmpdc
clbzW0u2avdOyCqhU306UEFmqaZhp5AEVbJUZoTcqmy9WBmMyGaiWc5dyLULAcQrJwDBzgvbTiK+
SRNfu22vkjSPc5I4z5CJIxLhYgfyHo7wwZySMd7T4gSVNcLD9Qne1srRCAEqQUB4nj5xFCDIrV6v
zy+HuNG5H/y81ioIHhGgjCP4Oj/LzSWXsUnTx8G/UYtaXN61OAuBleG+kQoBbDU2TUZB+MVkTrSc
3tvSKbruw0t1QhSzUMOyQotRsTxOKQbqhhzMRQp2BlT8xg90nL6aDVuPNJtEjgir7S0Ei9Er+ctH
hUiqY4cQuhHUZ51lbD90kZiS47SXfW11NWC4wWp8N7zdQsXWO8ACl3+WAq72w+SG0BZ0fAiQhYCy
VkfwNKOYYxOCG48qfQvxS2LAf/t+LRMVNoQECngvyMkxI2iKYMJeCjDP2WDfvc9zIFkvKD36k5dg
Ke+HWbeQmZ+D9FFNDIQWzJlgdAQ5Wf+VBvWsQ9I1tJmrgOsUvygfz/tk7DJQpXYJ83rf1fpqiC83
zG0oDz965Kq6vUUdKMqRRXeBQsSdEiJiKujsdcUx9/6QjEiwt9ex0WeaSzUOUdt02Tx5OoWVeBCo
aICJXLP2ajHX4wxTtRWfn7QYuUI35pS7cVe0VHv5IXjh4iMuRKVBIuFAJd0KuagBmWJJQCAAidmq
z0hfR5jGe4fy+f2OM/67eRaDqm8nwCIPBPoFqW9rpl2KJnC8FrdE3qEk/ZPpProjnfj5Ar/dOeG3
0mcI+8AnPvaD4f7v6Q5mD8M0VZ8s03p58TKUi1xosfHmcFtz4Wc21ieTquFuBEWjvqiNfKPbl5fw
FAC2rWmogS9tkRf5i2/CKijXS5uor16E+Be3oVEo96MbpCHDhQKF67RapyWHvy2FV0wKKQHsLgt4
cVTeuohIGHe4k/BpxvOFM4US0Av481DHa9+e09ACwIF/NONaedKm0xqxu9LGBdcbAzYleN7K2JtF
wM0nJixdQ4axC+1gQu5zdKRuoWHXCpVhAlUaUpNxfMMLibtWNtm43iY1l+hChnxRc5GBAWd+1UZL
acfYVl/jnGbYiPGEtF4F30lxgyTb8WYH0e4z9Pe0nZ9P8L0ihZEP+NGYDEHliBfYGl3/1utvY0gd
rTQo3Sf0alQYsxCeSmhP0WLLUqFhvL1Vvl/+z+2eNnDptTbdEbdxNs46DqRk2tvnAWRUSB+iM8WQ
9250jaT7FTMTgEuz5c60GsFSdUng3YsadyszAtxH5lSuu0cbJXFbEJCHshbg3QnBt4vF7hHhA0bj
pUhCSjE7vtWdJDca0mYUfzNEhkNSTQHrCPsTL9xF0f0O+IM7abgHsNS2/ebJsgDPOeEZ2JjbnOCF
HWa/12qdOtz/Ov6jIEl0yKPv+Q8YROWxaVR9kI9jSHWL+kGyjvcZj5+9E29eXIzdigE++bZz/puu
IJvUS3Hh6lrxOpcH4rh14kD8I7XuNBlW4mIbyHNCi4pXNBCUJZVgV8tkvLV5pWjICkyDKKfaQ0Ur
w+1BqqEkXdocdJPZUVu6JyyLUzvpWrJ05M66Oa/fubyZJatgkT/7GF9sbleOXJkanylPCI/+44QJ
568+6VvTUtRU9Xhl2fi+rB2whFjVMbIZtdlZUbkXvD0nRN7uBJCuyRcSMFqMYX+Powq7KeV08dK9
ZxHW7jXFbvygCTNFoJ6gGv4l+ScDCuIorA36bGtFeIHYyVGqNYa0bQsRnQ3ACAhnWayCaLWO6ilg
CI7AaZBGBh/OJ+XEU06s1HjsdmYwwQ/8mreH2N9rb9hvOjV6Ny+8Y2T/F6VFjocqW7p1rlZ/9cD3
Z0aapzOf30fyS2VaBZFXJ9AlDuyswb/CxgXQftOX5KULkaxBcA63LQ9Rh+AXPaSD+kjR7PsWHYcy
JSYy4t7a86dQ80oS7weaz9pYOzsQho03olP0TIB9AnS9xRDQhxE4vguqMC3WfhFcYORjalmnrc0v
b+0oGhR8seI4eH5YxSndVjpThJ3ez1/GhiFXVdvLNrV8TwJRVvyIts7BbZBjW2C32D76qF4vc3F5
jaJycS3ftQee3q4I1qE6qdx4opsmaOhwAFIJehFdRv1ehQdxFWuob9c1hSNnaemwzvk1Dk0MIx+m
Xdc75z3TtZeCfT3xaUvwh7GIp90jf/VV3Wnwi8/sN0WPM5/IOAiydk/vBNBzJ929rkHPoWkmV4jw
oyRu7SlJCfiJVfWm6epHRC6xU/S2JdvLYmRLblCIJ38T3EuzwIXDo9Fpf8p64srLaQCV3kjJAmP2
5coh91m+gT58DJSVskJORpJXNIbBmtLHL77qBNrEB+tQhyWZMC2oM/+76w8ocgD0LNKjuJ6rtOfe
cUz5cvQmRvU+fDkyXo8x5/YHj7eDLNqsZ4ezLJ1+j7edcnPF4bvyQdpeZ7RYCwCVNVxMqR+p0fur
2DdM4Z6EXXnGHR/Myhs1Ypl1UDhDRWGtJL6a5uUiok0e84sgmmCnZvwJV/QhiIXv+UyCk7nc3umg
jaue1aCTJsB+t8SZQYBiKq13K3I5SvWp4aEMliYqqw09Eo4/ggp9nUGP1av1Nzg9wxbELYBjkEsz
grfAr6e3XLBCXNbblipSu/ZwMYDJ0SxIjVHsa6QKuZQWTEijFJerWPqpYCyU98SQfVn63bBNcUpQ
LqtpA6i8ZXzK6gvWPQjUjX5tx4F+t0i/4rwrtOUmVaqb9APGdty0X/b3pVy4M7+VCsNJzUXYDmtO
1ftyEjttFhVa+H/Xy5d9d0FKwjZfqlS4bugSp5IBvDxt60Zp1jx5aeO/VILzDvN3U3B1Wyx9zP9P
EXBKKnQAruB6ob44XdUDCXrm9hkLi/sG3GXIcA9cNIR4VWnrSBhimzrmHupwsyZ4HltaXeLiIAWj
Aeo2O5JgYxJn7FbI3SUwn8Azy/tXwBgjxy1kgE4mek9xNyHxIP6cLr+FC0/Q0TOtmCeWphpDVeW5
YBktofnaFToimSJR+jc7rA5J3xJz49CzEyvlVED6EoHy1y8Nx7vYCRwCYm6pWoPz1d9X7aCFDbur
RPBNKn7A5o5/nJNX8Oe1nRZwhSaqkzxFmVLdoSPX5BrHuly1sYuvB1JeDgXwYQ23jfCnFHzrf3tY
frX6RES26VkSkwvlG88qg6IqItQFvPWGXtYeaV9dwxkkjvEeq6bZeXblFkewiVsMWYWGe7lvtDwv
pPONJRVfOGUHQ05SgdeDNNlGN5HyA+9Es5zDSqvfwELF8ufQXGc7n4PQjBCztvNojQEmf3z/5LsI
RjqY0eEj03fxZcQKdp/lEQGRISNzp+KAODsMsq6jaJ73N+vHvHD8Wim+BUNBoQZbBa2dg/AU+41V
n3Kl8blbTX3rbXKBeoreB3QC86dCxUOZvj+uLqn4zYQJxUPQpuAdMJWJXSuK98LjfClaekECvkYf
3R5EnUssk/27GSNOLT/YA3JpPZ1+IF8/CrdyCyVQtwbDwPT8d4DcS6fCgU5LyVcpVxWjhLm0SyEk
aU/UMPMUtZFPutWWJ9zqOug9hwVhiZvibQgIqmV4qu9FRstJTG26hFgv1kUESjvRJQ2mMFpZCJ98
CN5TQWFKqjN/+dbBpmkBGxRwYC3wn5mCSKrfbcxwLGZ949I/9aqeatQ/9sIj1yJCBfxr/snAxmmY
i7rMICs20yn8O2ET/CyTaSHycNGyqF82G+iJVjr5jp29S7v4X40VR1pMkq6E7gbrZdq1VtITsBrk
TAjhRo8MhoMPLugez7jqimIMm32n0kdUNPIRu3DvJ90JuvrchqyXYQBuxFnuz1gaoqtZRZlco1JL
6C5Sa0tzHaVrWGeJm12Pi7cHZCf7rvDhmsZpkLPBfhoLzTQSr4fG9WoGvzSjO8lNxFDoIBWvoXFc
MnDYfDcnR3BZm0YtC6gOEV8kg846GcU1URkcXOLDj1j424wW63DYJmfFMcCAy/p0gkHd2Bm6Kwos
mSX2PqqxEjhMM2jgkUPusOfMZ4g3abXToP9Rl986crtWa00JWmuCqJHslBgEv2r3/5tbrE2kXebl
RFwb56hk+3/xfl2/wem8kgScXBXJwoGDxwYKai5B8YBBj7MM7kA5SOD33VxBDBM8HjKrmgfIzUFa
ga750xtsDPUZx1KIe9ZBS5QFjHVk2YQgBg5imIuE6gRD31oAUMWx96QC1hyak7E8cDidN5ZfmFYC
/+s3v8UApttkFExTO6+xy+GOReOuYmc8eJWa2zN1Oq+nllFQ6CKZrilPIgRxTTFXcLDQLc6Zd7fU
uHzsdbVLG3uEpoy1aHB9qDtZraJQSW6e4+p7ira7qfohnrzL85Sj6PdjLvuXVBTsqu2+7Vt7o04N
8JX+uYQa72QkeWz7ntAiFiwtzARTm9yl6Sw0dDZk9CYezvAl3mQoN04bYuW7dQD6WSOeOVneQr2I
s2e5aZTesU3VTs46+tu+WEw4aViDjs02KDseRL7SSw2qhfoiRsK3iYcCR0pPtKsBxMNFXd4NGZE1
HqP+inrwKbFTmHowh4W17vzXdK0qmEpGtrKwomggWvAHmheDHSTAk4uKnPTwBSZHAZt/oGe4TOAZ
8KS2bNHdRyNwv1acHaS/qhMZaJzxgtBjttelvl94U6rhGegZjWiDisiXDKtiXc6/IQorXTfF3xwr
o3yJK1EAzI4Sh9goVO3T9YSEPuubtMuZoCpXCd8ctctWJb2d6a38lhlQIr2DThIU4/8OEERjOBCw
bqgZhDD5Y2SpHB9N0ZXYPKskaVa7hcQOuEDNdUprHPABeyVUbRdu8owBXmsE8uwhj/k0huqUCMLM
krwfCIxfZreHaslGF1k+i1Geo5azAi/i8dvP0hWdwPiKOMNKGWCpxV4Y5b2SuBpA1xK7RIAKs++c
2uW2kxV3kHG7JxMf2e571q61N5KcoJ8FZ5u/1YA7GD/sJ8tNRwYGHpfobeHtP23MHfUPgR+sOddB
YRk3INpNjivn8VzgyM+JCXqerm3DDMy9/oq4wa5aKQvKlgMC/yh89QrRuU4PMBtbjxYMgmw5Y3yB
yDrL4+Hr2KPE8VM5CeSw6v/QiAQN0XgqHUztn0XwRu5FCId3ON2+1gMCSnq1h+Koasvb3GaQyTjc
0ZqywlS+hDJy57Z0+Jz5TdV9D2opjcJpdps74OA6CsnoYNOYLMo5JayGMFZWc/0qmVEzkMgs0NcF
0AfehLzJXvCpcbw5q25u1ZiX7IPvOApv1n1TM0DvrdEpEJIjs1Darv2MuMRPDUpElN4eWdyhlA5u
6e68fVocj+2miJszP7sQZsxQWmEA3ZHvU4ZOUPJUC4aFpZS1dDyVMAhB7skb41ARvIK6jRrpR02p
0OmYFS+MAOIY/t4b0e/iNAR3o7FTZxQwWBlALae/c6GwytSZGHGH5XhS3rZzCyUa0pO5nlRfxmGM
NB2n2piPMNT7dUXg46BCfAXTyc2rFTfAZuly85tg3FlQQesAGFHh1Xj+dstzwUcldlDaNtLj/A1Y
5E5X5OReTvdB7EqobwoSoxpH5hVl03+B70gb0sYqn3jWuekq6kchwjavhsZmFRsXlxxjZL+pP8Rm
lsMi1BIXQALm9NC54GukLclMq/aXRO9ie3jooZrsmMFFIWa3qzqLJE31Tz+5QYSQfZ2UtKd+Qwo2
6kuLDbtUR798u0D97Vw6qYwEbovHW0+0dRCkDOgbbPf0e389ey5oOctPmr+QGm99YF9J7lCuHwJb
sRHVkHiNg/I+P5USCqkMjjaTRY1qdVSPw7LmEK+TV/2RPH/Y2cxXOD3S2XSwdmnTe1rOlRP8UA12
Ab1vb6orhv13FQuSm/XqOE0rvR7ZEd7DfCK7wj6kdAR/FKcZofod+d+PsR0F2dzHNB/B1Mxvj89L
VEzmS+x12JK9YlV6ef3MKjtH78huPMuZoS5ra4IGfYcFQbwYaIol+bs1Vp2TYY8S5uazWMvd7+5v
JcTQMM380OL59S+pOlhxibPDPk1kHps7g30YlFRbu+Famwi4840WXd3WbitWKcdaXhUb/ZG0Fu8f
J5NCruBgMPueBKigecDtz/PiLFnleTQfGscGCdKLPXOZm9dqRvs5ongtqsrwtHRYX54T0uMnU00t
ZqhhCnGz0XegdJ2q4a45gQaBpWUEZD5QRjE9PmHHbXylqDwG2tEamXmtuT86ySncKCU8aeWLCDjS
egbmPETdu7UbsQTPfsiag9ERioI/df00WwXwj9i3hb6p5xgZjG+BadiJN+ypaYak3AXReQNkhTlK
ueTE5Apf+sw7V1Gpf95ibL1oWyYmSJhvMj+V2/96gJCNTdSYmSC5etyA7wRgFvMcx9t23wpQV6Fp
8yIhM/jPGhTxmk99k38BMHsRsMxhkr2LJD2s6nRNn2XLf5Hj1cWfFB4pTNOWePIG7qiVLmzSL/BM
e2aqw/AQ7d9pxH98otk1PM7/f88dUfOQLdIJ3tHfaJNlBWEhNCX4VNUdylx978Ito+JgxViX3Z11
Y5bu9EImPbNu4+xpxf4ZuzJJG+Cig8ALtFWGi08ndlS1lu9fKNLSl2Ddezs04zvQ+SRS1bp7MPoa
Z36CpqnzKWqPoVwQZTwtUfifyTxZ21cbvQk4uSBxaNnrV9h9Mt5k7BZ4BDXEgkNCkOnEUL/qzdvA
yUH6e1JXi2n3b3MRjJJ3je0u2n54q/FY1yaYXIZaL7RMvTvajlipyIoTlstXXETkGWrcQJASVw8N
Y9ZZjVMDsowgWdzZ9qrYUXhQ7vB6aZdBNJ8XK/ZmmnmsYGoAwcSKvVUEiigdgj6CYJOcsdSfhVbo
tT4V0my9YA3Is5w0iTn/oPF3bdYfLzMQ8fGFRFtSq1mWDGbr0IXh+bNlCMpisUYjmhVAYbucoN00
VD/mQ4o34IME1Mifx02KguY2Scikg29fDeO5CsbHlZcd8VI3+SrCZylBGp0f/tDOE4v8lwiZ0nd+
5vdqPppv67LGZJU79y9hoCGvD/kFW7C4BOri7xbPlG9HWur3rLEhwSBUqGpwFisVl0HYKm4u+SDp
4Lh8Cq7XQTY9q5Q5QVow5AzhYjIK26z5DH9JdsGfIGYsfBE+z1qSBS/7hVRxp/MKvvJrvuSF9yhj
5X+igqAEoBTPEguebF9R9E2WbZJP4W3izLi2ndFjS1PUfBsN8yBdVP3flA7xpum7JR3cx4HAmhjU
RM6paon6JXe3pCshcMNIPsafkkem5tFz5EYLUA32d6WbyqAM1LsGJ/DkQsDXtDd00S6eZ8aYpeLr
zqS1NgmwH/OIulDm/x4Z1s/EUg0UrU2mAe1km+6JBsygxRIWinzr4PqJJ0Pd3HzF3p0CH+tIuj+h
rdUzwFIEhfm7LiaAw2mi7V2qdG/XGqjHaqWMeYunhlxJg/l338ExvSR1fAjBVOSrHogXdQ68KpI0
o4dLSJh9nEV8yzHNBlSU7R97bw3kGHGHySN2XubmEhptqsD6bueXEb8Ff3f0kC9U0D0nsCfsfdDB
tvowcz4VQwc6WoFlbGNywYj7CuH/86Ni5LZiW2f9swciTxfigo/j3rm6Uttv2y5yM4l+I+GGWHPw
ALO/oz2aNUV3hLQNIIf/df6sGTLKVYjyICNeP+f4zZwktvUtyuEwSP6o5SAL3Jr6c2ypMldvLBPr
aQCFmBqAYANDf0TYUtEb4676wYpEAG1t9gDp7rC/sdEky4bdPmfynGOkKH7rMPHqWRGtEAVIktEP
+3TwQlrjC6L4yK1siFzbgn/vI2BbDSYzhtYPDaT0G89vgpcQAQ3fx1HqWQavsrDKCWVKnwKMmrjN
rAqQVgZTmstPIcVnvs7exvzQztyntGnmGijW4yHDl+aamMxoHqWCAPnBHNIAMZe7uy3a+mj9eko3
0jBiCBtfsz99Ft1WOlDOug94+/yD+jCYwIPNMIDDLannPinUbPCet2xCQoNSaorAOMiyBMaaPFHy
B4pgA4gb0fdqV4mmASp8wN3dqCdIX1tPe8q78QbE75wkIfJ5kzxCsT8bnM6djBaE/IYW3a22pfB/
XDEFvAQOdq7xs8VBg/cICxbad76NntnhxZlrFjygSXhNtCqzJ2PpxNZzW32snGUOL9joecObYwdd
fC8TgOp+tYGvBwyFXA1PmcHEPJNJHDKTIy5vDtoTpTiQnvPxxmKeCdcCTFDmha88j/cXZnUh9cPR
a/9uYKIvUvVj125EcAtYFVDLcWcI4Id211YARpNg6+Vs3aWRVNcgB3f45SpGW3Ug2rTfXMCDuykc
EZVYMFBzsmwVfqMJ+NIP66nKCCIJzP4CM1e/+brKDP40I4wL4b5opy/hJSKukdGXVrM67pyH+XcO
ZiY70NKPiBXMfvoFnR5i4bVZt2PcjbvMFJ5Ol/yEoUv4cQrVcrCjAHjwmKtQTEuZRcfrdVlNP4Sn
kWstKcwG4P4r6BJYQNigEjUVYEBA+FN1nFsdZ82UiI8RNE4hPhqSrRjmvLEYoln0p02y278OECUm
v9JVJKPf+iGMG6zoMd4lsKD4UY62l9KO1xsf/letUpcCqxG8DlNcxNpwLg+PtRQ+punx+ncA7QuA
2/T5C0zrWtX82s6YezPGYe7w2/K2M7z7T+ZcAs66mpHb06TgJ+E43g6GQo43BcHRfbU2PX07/Dhr
7ou2Yc8645IjhYULX8EGhdUg82X29nyOMtaOQJdZhmhQCdpsYZfUdg5qYAG2inVXkjpNzQ7tpRT/
MmbgoMUdgyoKNoxMCbO9XfIuM/0ZeHj603r6uuklKkT99JO5MGy8adBp3tymRdK4vIH1mkqIDayr
fzzvjWsu3KkbilFvtZrmFiF1oaru9GRDRe4hiceLIfOivHbSBXZH3LHjSnFgLc7Tk/DjSXl660jB
vIqDZ4fuO8vI/Unstq4dWJoMyIgIx7VIopfKT5kicJHhJ2cyUzqJQeyYm075GFRD/Dx+XxGJuiQJ
911IKL5xhImvDXEyqWKQegYs1bC6RgnJzz9wFfML7jYqbUruio1DdIu0Ph32sBzcCbcXOi8wk3pK
qLUHXuRpr4A4ao7rhMaupSsSudLbBRhyPHXSL0MwfUZ42QppmLK9WguqoTusJuGW6HVWRc28dBLw
xw9Ls1kOPFCM1BUUIXtPt1fwrUzBwk0qoOU4OHMZopuJRwRldlwYA/kAw2bEeQK1vWEUZjKyzlvY
RMciwuJ6EUlx4TybvrTp+75ioOMXe3LUtFSIz2S1/e3g8G9NknoqZntWxnPlQ854xXbeA7KuoxwM
LwKr8PSRYUoerMZsPZzEpSNaaog0loEidLVQ8ROdSnuXJNBIAVIaZHzmvvCS5R5toTzqrnaYvBEy
ZTq2vQBC4p9qblO/l6k+DWtEqGCBUG6QmJqoLUZhXS6pSCLEb3t4j0TeFu7fiJqEjokjcsn5xjmi
obeFi4NE0tbTiQMrw90aTMxvAHPKiUpgzrHVZbudze6Jsm0YIhIhUDV4WCa1ivhjvuMNW+26hNBA
ZSWxfaXMaxR6+cgXlIAhxRa3WKruND7zX/VKHDKpadu8CXrYBlbCGRiZ88/AHSD8/gdo+GkIp3qp
5IGURCsXrl1hbyRKJ3pZ7uwrBiSBmC0dKKrDUdayYfDXCxr89MSUuARaJqc4ZeeTILeLwh4WyGBg
EFpzglGAVc3TRLYpB/PGVhXP4Q/i8+ovJ0TtbJsv73XGX99++Uxe+pdm2pqv5s5z87diSJeGmC5o
kSlqKKdhx3swmCWwyMM5A+/5WElfvJWPlZljua8zwano3kak9D5D0QWvilIKWkw/8CeatWk2oeGl
mU/fXNnAVbo2js03xFaER5IqE2dQYVsinAUUT9IJqH/fK/sQgibTB7GycfgE1by/KK/9U1xc+Zbf
nJwb50XVQUCyU/hrV/WGwiFCYG03/Wa/z1BC5KspnlVev37VPPpy/boxVbZrQzUmGEVmqBoD7PkG
BpHrmIgtldEPqtpvKdz45pgi2QWx6BPTUdpCv4ndb9e+i2YQc+74y5Qep5REpdBsUvRW8d6iU/dH
d0KjvuoQTbf/wHc0vdIDHmmjeya8QCYKo1d+TRgqNnWjjM5i49ONUiH8O0S4sVsdYjobYLx0YJHQ
1unZQETPnqYtH+KFBcsTiUg8yUkuuw9UBKheRusJ8YJTdpgb0FAaAWjWwUJDecLRO5DxzXen+k6v
aQEdflPA17PCy/I/4wmuT7bhkJDYTODRo+HXcpZ1rtgJpoav84z2chSWaCZDAdFYZ7uzSpsE3wS/
gfAidcxBzGxn+tlpc5ia0+wCDkJDAJUjGdONeYshIyHn8ycgNaZVdJj9/CcvBojC2pIA6UmJrkPd
TT7KIqoMUvIDLqLdsJtrjUAh7bQuPoujbkArJzApKnq0reTvtQN4io4OkMxbCYRUtAn56d9HYbQ+
ZfHBUzEhjN5kvsYWKOH8cVRFrE37X18eVT20DTx+PkdUBSJp4hW1PpFQtCyXszwAcMOV6FRXIOmT
7ToJsRXvvs4QmF74mKfkKOZ98O4GWBaSMMGo5v2mIv1C2pOsnNd+sMt+LXlyjB4YfrM9nU7vaAkG
ojcuOG5aW1MQYisMJgPT1VldQ50RqrhFNYpMLSp5IQC61jkiS54FGFA23B2h2j2PavStWpx88RBo
zaCYdw3kJbsXHjLiER+94o8/9KeQL7DNrs/iB8w6QbP4idgijnuWQkkgVi1o+H+mtgu2/ZftzKyV
uV2Erkb1b72FU54v2q0WnHUb6kXLHTdwd6bVzu5XcYgyaJELolmPXAeQZnq1rpTNETsFC8HPl6rQ
RruYZ0JqPcofjE7tXFR8s+BrsQ1ZlztIy2NKRzntfUvRwrW+TFPtkOy+59TBqnWU3CTlvmunx6wx
JHNJ7K+YK7rtFyPdp4YBn3hBxOgUw8ClDljG9pNiUuwQ66vE7oS3sGdXpHT9txfGEEgLK5pyqGCK
THOHbK0lEMNeD5jEEwUy8tQK8dk/I6FdeNHB89i7TCbwt4VP/Be2A7GEnVQGEgo5q6Oh7nm6MFRQ
Ob1WjlKy/kE6i+QvtWV90ed7RKH/PRtFcRWe5xMpiWsCEMQ+Rd8rnWPbhB1ZARzTdtcc0xGcNbCW
TxhKmfo9gGcDiuPfZZyWj1cReAjm7Le2l+vwRJTd/JAeiSZ/57qZDbRpZbjhqK11aagz58FFl02i
RbdlmFOKFKi46SrOx9uBG4zztrNcFMYyoFyVz5fSyE5zVeVSb8tVA57A22j9HWMaspX+YOFoS8rh
2qXgdbYbjT5sMmO+zutMn7SklgCMZ+HOt+ubpRhjKIwevD5PIptiJr6C56/WH8VyVcQJpfwX2cbg
muNYZrFChPE3tcRJhu6yr0ET/2/syyblnWzjycFvUpYFqvgrO5qng1l0VgRGF4aDQZjvR7eTlPUg
5z8M3OeJZqwC1OVcpEP/7YTDaA9kuJvSbc9hUtsvTougktUyZfnX6CzmSj6t0NXCWvmuALCXBmAn
YakdVHs1L/3GQnqKv77Uvt+/JeN+BWzaCYgvXxcg1Y50DPlvbvyKNx/NUCTvdNwJDa0apn9nl0Og
P7TswclpzClupGrKkyixdEglcKxt0wLCcqUv0qbJ4tvPxteEpGxRj0u/vD1XiIZacMK3tkUMw123
Jd6++mZddnDOy0w1uISYXbJMMEOlp4x4ielqlMSWmHz/qwZWxuORtW5lliXEzyRkVwpihkSjIBU+
W7g8506M/t53sHzSfC/ybIaGna3E1LSbnIhvXJ2k+ilphfKdxnZd4oXV1VVEexn/VSvuyGwptLqE
acfk0rJRWY+iBOVRWtTbvUSolGXIWYMb+UD5EU8mQzc/U1qzEqijsZjB9iRyvpgtjFIcvkAzUpif
8LIXx5PoTJGOLukae0UA1WFaEwaB5Ydin3suzPH/XS6r8kEK5p1aQvOC340UYvKkD/VSNHubyeQY
BdVfIi4wmKx6B5BClksNfIUpRzVrituohfqi5ffVfI11EAx51p3f27fy2NR+lX3H9v4uvo6AlkdP
Vh03trENUPkf/u7ks0AXX+nICoyL5E5b3Bfe2tGcnGRvJKoqsVXgtyvSqFXPsAGKDdI2DuF1UiPd
ly9TwX3Xz3SmBw1FFGadAPqiSCZX2FD7GEMUxfL9E9lhidg3dRffPSf6giWX0nzKAaFgt2WkfJPT
wgDTMHY/U9INSCZgm6eCQCPvxEM5uO9a9g1PwUAqRh1/dD6/F28pZ5DdIiBOgNeXCe9t/blGL30e
O21GmnCv8MUcXRFRup5kM2t+oOOiXDwIVyeBe36LQtxnCQXVXPLqJzUwO7oFzuxwtLuuK89eWEhb
2w8k+7dl8MmFlLiaxTnw3B0tGO9Wta30hSi2RqyfIE6puz+ZkXo3Pxx2eP1Wehxu+6YynoI3GnJ2
tO/e4hqco2npPjqd6HvFNDVbwC9BvEGpYw72/nB6G93Ad4MuM1DoU5H5eCplA/N9BDP6u+rH2vJu
c3IqjJWIiweZUlhkVFHLsDZgx0zVFOoPLFQfVIuQMlrDJhhUQkp0e2tlOUI6x/rRMYCvHKX+FcNe
qq/tib/M9o6gLv11hXRbgDrVNft6qHQX6uVfa60xWRhpK7ixojXpFiKjgS9lmbCv7vlqw3e59mFp
EQ4wRBBN/wYWffvDWLF3tsoO7r0Df2suMZzRRgGCrRk26SY7kGNJhNfBBXP5bFQJHLIOQo44Gxxx
XE1uQ5bA14I0f20QYgJ0UUXDn5VHKewvIa5h9Gac8Zyas3Xf70yohPm3SdKhBScbXy5Ymbom684U
shrMwJm6hCyQk1rqoiIjlG7QK2JvbqMM9KLxJHFKydcrxG3qZRs3dQuZTBDa3XwhQJ5trNGPCfAD
s3jJwyM2VCjnkMwEyQurTjJJUpBQIWL6gF5OcG4TIKEQktPkczKATNXnjw9f2++FpNFeawtbNAOm
Nry+6wG1IDn18pRh8ZjkFouHCj8NgiYT5ldczNTfC0LZGaf+YUr35T3QxzMaOTWbTyixrbXG252X
htaduP/IQHPkM+MvHPF9D+azsgOnn+LpLZpPq27ntaUwIVBpy2KySjBNsEbPQ4ysERgdfxfBCWUU
NVN2EBJosxLBC6MCu2UuGgoYA5Tul/UuracSIXRg747v9r1yHuA2JGiHF75cL+4p6G2vX4konsTy
lS6Dsf4gE0Ig9TYygiUCZAv4Y/lrVz4JaWrpjq/+UrmZzF4Ek5v9Bb1lkdHrf+mOCjImuWVLTTT8
b71w09g/mV7UeyhSCvK6qMi9jeCP5T8K0H8tfbzuo7bTjwWCUP5R0+0sfGac5rAO6x7yLF7yY1CS
srm/TzI81FP+TxK11O+4Y/hVWp1rKs5EeEeXCeg3wky/19L4VmkuEDte16hmNh1o1R/mQ5QQsIYf
s4krPdmbg134MqyaUxpV3sqOFFFMFrDGvEPEcgg4xarMTPpMcya951JHOs+3wcgvQsQ11ezKVxWB
UXwSczzExlgQt8NF+HKSGGojIxome+TCQSFN68f/mMqGyydfxo6JS4r5RiSdF2xEsSPV4zQ8UnWU
O7Gmb36f4qwp4aExhVQe+9sVU4hCed4tE1DQBeBCKEVSY9jOHL2mV1lTrPh2l0rbc5/QenUj2O7X
M3e8TjiWlJuk77wV0WKqg93nouq9KEfabrlzGuX/Bh4on75cO06ka6EN7wLFrURUeD2D2XzzAzfW
iNF0zVa4hmLPORzxOLYkr3DynkRRCFjQFu5fuD79+4pGZwaIjk29FX/ojqyyvhoczQ9TTfCLjcLY
B4zePr33IoKRXzC1MzW04zk0RTfnNuVcKN8lbTITazctSczBPHAJjiThji0b8fGuNZYQ9Tnt+KMV
K9bFXC24B0VjcL1TSW/5wjBKGf1FQ/5xcU6dAKyJ1rlutw/3qHDzrp211wq0DY63gF06N/5EoqAI
y2McOmDnc5m6pZkCdcccTVeQuk8Rq905Fxfs3imX+aUBr1UONpm1MqlcsSZsG9kywKFktyTF8ekV
w+vFzA3nocQa/l6Dc81AB9br5fabhHfCUy7HkDTS8cQdAMQZZ9JJstnv66xrc5MVPb95s3oPdaJg
QRljd58OlNrz2bBJ5/ctsZUZlNY4jHgHNptvhY1dWQFtZ3XDCexOZLPix14FkIlen4S2m/jiKkv1
P2ofcCdb3LLc3OPzEBKxNesiUqRpQYPrV1Q5jyJ3SX5Uxh98zvZwKMutn8DWvxgr/XJP8T8fbH4W
EP8TU0n3NDffOOmUU1CvvKflFNzHMDPTtZ7gVfTyNEl8BR9ocOpFcTvy7hO/8+2CuESw3UTLU5ql
1yLB5APsBokieM7ln30ew4q34J9PSpZuAXEP9lxQJ79UowjYKTGtAewf7PD9QFaXl66yQrLERH6p
hXsFWtaqlhsDoSLO01amc5NBNdbTwilC6KELq6SpcjEKF6wDbAitZYoomNbHjL5uje5r0eUev4vW
fESwN+jLTkeVPw34MQ8ppjEclaSc/O0WU7VCjwQaN1+Yls4Lvfq9OobbwpJWuy0lN/YjGYDxhuBK
RXpYDmDJ5dbAC2Q9Icuz/0ReGxtfIQq/anc4+F4IgBbF0MW9fP4OmWI0utdVBPT+nFyaOatrxWvF
jV+OXRvv0inI6PGzMUgRHlo2lsodHNC26kUPduD6TObUpC2N47xvnhoANeFMsTjXbRlySqwp+Ta5
SgIzb88I5pwBVR2IaFUo4XkskZWuV2vZK3Zzq6OkXJuPVh4IzONrVUHeCulOrnZzzi2NgNhe9+Ek
V2KYeF5M/8nePEvj3qfyNoR35wRyFf5OW8tZpd6yMnHCIO/PKCGDR94ye95W1wPGf5ZGmLYeCLoP
jXW6HxDymo0G8oyaW6tcfr5UWbY54I1TgP9OezYVhecgDr+st5GWe0lwWd1B2pJaZlgFHhIDLrB0
55YGcB27zk0UGXQgckYpvIDibEzzGwlvX+qb1hL/KCs74RoANDLRmjzm7iy63hsrx267AOpVcwFw
gsoc4j7fLkkPnf4eRyCcMDgP75AvPbBH6jn4rHM51pskdp+kDi/UWZtZEurMGY8dqsQxSuhlLzro
ATTzqooF7sTsIn5BsDGK/vt+8U2cdOF9FfHHDxJsL/Pv9XS8h63+VsVAXDVr+0A1ddtC2RQSQvzE
QrP4nqd+f3R0qBj5q4HswmM9YBWQVoxKTMtdHTo0O36a04PYY8ipUkgl7wrG//5q82sF8Hyq3M87
XO+//4jpVKwaqvf26lVYkrmpuuVpFpyKnpUXfEODT2f4eQvgrZv/MEcDEKJ7+/U0Fva3p72W5PFL
MAnChuNu4DQBCQre7bB7rdr5OTvgfdIx5UvoA0NiHnNd4LLeSU3q11mF0nwW3GwjyV4SGBluEmWh
sdRB6e2vRwmdpFumCS+DELrWUBSm6F1w6Co+FBkF+ACQxJ7eqScPJqBvB9iTbazvJtzBBt6PivAR
a21wA0UWGBOWIBHdV7S8FjTIPK+71ATGrwvwS/oN7jEq1ruSOLKTn40vq4wccLgfJoQ3+JmmC4pF
FdZ0v9BC5bxVlPhPN32davnSbHcE/gvh2XkJWM/O/+AU07YTOAaBUVzwOQFLerHr+YagzYW9Pkij
6N0TEE636CTgAooQc1UmnjqSsRZNUmAM93fi+mjtpkHz11wOYJBlH4+7P0H4r3AgCHkhvz/on8Hx
KhaaXY5exFFxcQnq35cw6L7pF9t+Na5N01yX8duZhdIZ0NcrYq1O+gCXrXlvVfaxsvtLg/oV5qnS
L30lAF31O5Wcm5QSlwriSfuOEUZk8dLJbPH9hNpZHI8vMufo5tT5WCVY60NDDCGVorGQR6LRUWsV
eWaK7LVa1hQdHOhIhM0rKw4SstiMi34aJlODUJw2p5r5iCeKYgtyyL70755+4jq0tqBKC81t5ka8
wkw41BtzTPx+XJ3ixFfYugyaIGEHII2MSWH8q2lOPUBD2i8YGqeRDtn4m7kVvRHJaiMxWhWjwW5X
p4E/XTVdgWIQy9ZEDKeTt+TgwOtzMci+rf9tlkF/3S4etqq+umDSEMT0k2ly6s01/sqZLbdxiMgw
TuDYg4P6lldU+J4dH062sJWsWTOjzXBYatdHwe2BFaavVbrHLVm5JnsGZC8muf29wl3GVUgBw55x
mWCEtnTvU6eKwpOpM046EGYws/HBKdx7ArPKdBJ5BuCW6ZfwbWp9lLUUgOVJ0XiCKtbKIS5WROKw
EZBAJUSvcHx3P6pHXZSluxxVZ56Ss1W5IZy+/nxyGD4Dy4x22xTQMWpCLQ2tTJ8ni56+ezvgiPk4
U40NUYzQty13IvYVC+wRy0Wu4+PT3V2ANfwINPigL41ESSUeFVTWShI7VHvOAAfp6KghhEMIb0aG
hGKlHadvZNI9+phl+ME3sEtn9BZ9aGGp9SNjWvFAxnM8GR/cg6OWg4/n7wiH6/Orl0eU51XE5ziT
UQHsGYzAISNCURyRVX5R0xUeJ2NDxvqg7EDEAJFAf19q6sK3t0BwQ53TUBO543XTbYIkVfHUmDlX
3in/hu66QwSOt8KwtJ0HvEcwjk+iLcaXLlFt16WQJBLQNRO8U5ProfEc68sR7SgQY8jBFEmbaKUt
vy7kfefePffbI4u+OlcZnSxHxis1/3Ld3+d8D+piC7wZJP4Nu+WVosjr52G1mqSauAp6HQdi72nX
3mjSPFOyevA+hfDl0oPQ6pQFv0JzAadh8GvsDghT2+kEY4mY6ZzZ+oFT15NsPHI7tXJQh2KFmxr6
JYhgWC4ckweqMeldiyVWruz0hWgS48KiSL/0YrxP3fLf+f6o51t0QJ6In7+FXdvGloxWSu2+N8bb
BkEXMnRri+VtX28Uadu1VodisLmEWK/uDRG4eL3VKWvPzmmdpU9s+YxZG3gYkPaT6Cq0iJUkYG5i
SDETjEzG0YCBlE82H+GRkEn4L3PVN91PPiQ0XQmVuba6Jmy4FmX0YkI9ExW6s5w6xdK85UosepH8
QYGmDNQnbfKnZLYfAQUgmbxTKYV//FwwpaIe0+OKocGY5XGSDzzVPrPHHE0cjp1jdMDU2ilxcBFE
+rBCbpOtjKIAL23wZncxlLULjxaqPWO1Kv5sQ6b0gnRYdElIHlTOhnBt8Czipae4j7i1OS/RQ0O4
a/nmz5CYjz4WBO4sb5aopzHtsERJVN+8AqBdUGivI4LXT/sRHhMpWlki+z/Mnmgi2PsiN3TD8OCF
zEmfLV/+hfe2f+JkWBk9MQj1h0m5mpqj4F4OTBpNgtyGIJ5+FV3kPu4ZwG1YHN50DxAOU3WPiRh9
n2dtoma1USjxByzieQz1K/+OkeiR6EC1PyLQK23k3pvp5IQ8O1EBpafRY654Qx3g1j3qp54BHQbj
GamZa6+UCFz1S2y/Kbg3jg0PT/OBEbG6mCESimA7fOBvIYZFJAwANbv7wxwH3ff4Iluab0uyn3wE
oo4hUYfPueT5ZEdJ65ninb6+pJhC23TdLm45eaxJGnPkAUBYo8kXK5xmdnPLJQtLJwGLwngF7ksw
9R0VD7d5VvzpRozsdMgyvNGQbpidHDS9+Zo2tWJuysKjMFXR9wvNgXAcJK0omYaRhsvBnRd4aVXv
LkNOsvbt7OK4dX1Y0Vk8swpXyGaXQ0jCCK+1MiuvuRMz9dxlyNfHPHbj4RZ/q+8nM28F3QDmbQ+8
ni2NGXQvQIm0xk6IW/iKNoaIbvXlVhbbj3ya1yEXNFewwk11aK0C9J3uVpdHZe0bYsNGBEYtXBwz
2c4b3z6yP3o0OdWyRpYWoPgrI/oGzWgO50p8RcGeeZc+AOO8Wz73hGi4KafCw5MYlzNuid+pbENK
RDllbAsF5dN+q5tAzlLb+j2XySb9z8MC/Ac8IbGXMVMRr1juZp0fOviv9QJzT5JinHmgWjnfKwbR
qTvhCc/nMOzSTwIwwnzLrtTOoj/iN2og6wDIXeAqqwKJZXhaC9hCLpZYF+2IRmWOX7/HHsPUzJOw
DIjVqsMphIQdgs8mtdRaEzKzGF4+GmQHU8WRYpYkEQktnANcGbph0KXBxz3sMQzBl2jHQgHoRbM6
XX96O1/ao14J2Va/3gzY7cLbcI2FUdstzrF4GpmitC097ubesGtqWFFJL33EOUPv6Uek4CcCFMjT
ua0uXO/CSCScWX6i/NFg9rWCarNUuq0A2PZlklpSeTxdjYLG3X6K5NZS8RAgs7ZB4+I/hZZOAZDc
8HN/3GT32zKwB18iEXO46+rRIqDB5YLiBE8KZ+OZI34irpRFjEIzOtlr0LxKB1wVw+3E0mFnqwPH
tXHk7yUlXlAdKGgczVerT0T3MaSiGG/kw9RGZ+CeJfgdQq9m0yyiV06kup4x2E1rO834mVVVjoko
XKieKhGLeab2XjPG6IvoJEV0rWv2rNGJiiiB++oiqnanMISeLkC4KCLzdYfzHidfPGtHQorDmSxk
YKD7mDFWypSZEdSCgJI41g+XfTzE91g79GtO+jKOLmi+ezK0caGqKdR43ihKM7TqneT+VR8236Ht
zeXyrbneEcMJEz/bYYDOhm4numjrbGC4EdEtAgf3GHrQQ8ylA5xMKsOB43wuba2bihY4WfHpjV5v
n954IKGFQe7HwnJHDrLMvTjwxc52cGCEHOUy50JpCadr0QS56Mbpd50XJ+cuvCn1Hu7EME27P23n
7PTBPoj1y/fUa4qmozOQC21ol+/6OracDUAvd/DukG8Py+Wl0MZ2kwjUpl0FljF8czQ97zZgJedK
vEPrZ0jtVjAlsU8IoJR7IF09WgHpniELaYytXBv8n7I/5Ek1QPYPg/TpFxnv9s+22WIg/WUw/9tf
jqwNwr21g0F5L4Wm97CeGbSc/ZMjCd9UAR2oRBpjDeyRtd4HVekl434vuodrhqxHNGGOfAiA5FmJ
i8Bi2BDXAcKZn1+IlsxzFKIMrVI6hbj6sCJveWfyirwbnHCl8cMRbpDSoAD0IN9yQz2952UtoTnr
+cfwwbOg+Cg6J9xDUneUq4lmDGXITyLqtTr9gOmktQ7o3OTO57+P49knMs0hyZc8iEW2sW/UXw73
cpicO8J4sr0WPk9rjW6HdBcfTsNdaTKaLb8sHupdGGwJeC1QRzPjYrok+KSnYtbrWeqlAIWa4xXr
FBUE9e9e4S84t/q//OSTEzd9nFc8wLNA/zJJzQIy6zy+h6RDVyXZTKi77WKa3y72O7w1eXuDekZF
se3hTuWNHdn19K0VxOdwqxJdBGzdICE0YgwW0NQe04v3LOKzzc4BgrSCp4bGYmRO+78LCveL8w8W
M7GIQMqKzrSzhHzCl0ExCCIU9ysiG4wGQqpSWOTWIXsW/bbhjfJE8B24PqDDhUtALFWuaTWUmpET
kXX7WukMc/gX/PxQxUHSiPNi7vh9ANh/uD7ZCLqDTq3oD7eY1pXcyjltsGhmooQ1Xntu94Q9bcQE
FjudJGpRsVbz5MmI//596TgczwxanSokAuvFqbJS+zMweHZDhXL9EjP7PxepvIbkZ4nRuRma167n
tChtTOEN9lRag87RF/NpfOb2RFZbM3IL8vXBCCI+CdxXlrQbJqt0LCrNRA/lLwuxVINytNCUr0kC
+uqZfunr5W6CpWjdCNDRfiyvnyW2Tk6Uw5LieqeZEq7z0HOLWTHxzksf0s8CKxkOTWv76cBGZyb0
QYZnLeL18gjH9W+FjKmxS8KD3SDsSGcqk6wnGrusV2A+fYYkzo+0gGqark4E536NSgKSooebtNBL
eSVnA11jwYHPaIBLRYmPjjNbJm1bYKIAqp7DsVm/4OncaP1MoqJKYG2TSooJSpQ0oO1miUdTV2eN
DrHz983BMt4/AyN24e/ouHOtmaNTaO4u1TfrQNi+7HpgHHGN46Jr/mtsxeQi7FnGieWAywGkzZ+B
IlVtPVCOx3JElEPfhPTCeNvIztNyvwInM4i9BbrYWk9OCsL5f4bvgLZA2fRek8MKqKkArs4wjfx3
+Dgdmmb5NFSdKkaxEt4xSZyOjFyQKZXPmx281pDAAV/QxbauGi1PPkeDAW85TMKuBkFEHuKCDyIK
QaQsoljakNdRKRwhbnLklXfmu/TZqCl2WIjrvGYiVLgrJ9ANmtjras2kRjbS0N2t1bf5qoVyHEkI
UvhGaHyXpPECKXbRudGWa4k7Wrf/c7f6tEhogc2xLPMeFT1LeHW+VDKUhkoLEXCfphsVl+8K0pij
wlTBVipo8ChQFvUSSxa461YqHLEgXbnHj87iv9bNZwtfaMcxnOQaem7ZJ4RokGrBRKjKeG1onYS7
f3/pDxqlMhNC6UPDqILTEZPPRIZBKKMn3MpU1bPBui0Ycy8WvTuLxxBm7Gx+8Rw9FdC6UYGIPoff
Z+YozaWbT+rYmKbSq5FFQpyuDuGP8y753Yjb0rmbftk88/CuiZOsw1PP086/B6g0cGoOXDjf2gF4
U6ocys8/jdu4m9oIeLE31s7i96iJirXUEaNNRvgBiCMcXz3zWWMv19fF0fw31blX+ScfK0CEpmLZ
GZK8X55J3RETQKoJuBhGH+1uvY4CWxmyy+4U29g+m1xJVGJR8Vi0JHJRktuefBeZ5p8FPBAvpTe7
LP37MFdbxqyZKuHSEpyttssM9xXVnlAq/6qTFtDzheMoO1SsE8xD9CRiDQeHnuGFYhY+e7wyNluA
F8qWj7laIFYYDE4UG93cLhkxnMK3HD910g6hcBBIslLPIIrQ2YNDosaDOLOEAdbHnDayMX++VOW9
id3BYibZag9dcdxPtL4RN+FBq1/A2bVIdeQ6V56m8ONlc+1iXX+PkXw7/6qIvuSXS5t+9ksqtOuD
0LEIKWtMwP/2JDUx8Sr1zgTf+8ImhfUx+VVyxV7iagnkX+T3SLwyp1yzjHGLSLP6vXmVxqa9ztD6
BAbNSjX64g1+2pbaLwxA5KBHoILBtejVCN0hCdggPZv1StB8JwTr7ClAHtEJOYkuTb0s8mZdM82/
6M3iJuy8a2b7qUNGsBIsrYHz2a0xMau4Vy4MdbcdCvmGPS9Db9MgL0HtXc50UcHVMItam/XhMlDK
LFm3lDzNKg14fjueDfsxOSlD+BMqePz4kWofjw1vzcmtUbqwqej/EUaO1kA4eaGsXL4Wr6IkXQCI
qPbSeJq0qXuc459hPNgCmKOAbGouDc2is8DVsJnkujqobB88vpGryCKQ6ItF5lpMIXAFaQpukl3j
2ge4ttEpIz1K57NnFQwFcAtx8bk9PsStySrCxjwuJLnbIj322YDD/qE1nvBvS4dGwwFGmOW1F2ux
zN9djDwgPRukO9tJ7BjltxsYwLsNjbiRMbDeh3EsTUsFzEltg3jl6y54CEOnvKL7V/rVkUft9HXw
klu3jULULCp8op8MMz9UetOgxVhtDbj5i73NmSl6o4bl9M2viYBorHywv0ovKceB//d+QZyuwaAs
mB7C26yHzEmQm9XpXC3MOBhbYiPU8vhHJlrw9gQQdsoPvzeWv8VE1cdJcpj7hPd2gL6hOThbHU7z
O2ZIGS41d218U0kk3c6ucp6b0kfjYjbmXB89MC8y0Z4KkRFCUK9xNcpsIKQCHde8J5M+y9k37ksZ
xpf9BX0bc76cdvDweZmvdU0Q1RlM3WV1n5Lt0j9MBZUNiCHTltwRJ7+8gDKDr0g9JsE9zw4cMjn4
cphJjzdMWVj1AjTRdJTLwX7IqaQq0uP1JZ7B2EiOzAVJwDRbPlxI9Igi4heO7G70IAcxo+oQW6Rj
jWbb10p68H3OsXv1nfJVwcvlW2LIxrMz7SKhHAMTG8ktwpe9fpHZ10h7SBszN42P+s2d6G7uPNSH
PnTk4JNDORlvRGX/QbCdVUKAK7EZlqg16vFP8HEUH+Xwmo6zXVWfTENBjTdsG4MPu204e7uP32B7
r0FFgQINFuHQMTMUDClXvT7e7O/0st7dXUBmhKjUuNpHsUY6gxSy70VAkelWOOvz0RUDGcE0yxla
lFsbNBMGdzuopy5KTX+UNw/2/zKba14ignIsUwLBcMP3ynXJH/BETEzg9OUSuPXtrn2aHdyToRrS
e0MRXLvP2tuysgLcxIKa0FlMuWj8K0d8k04RPGeDBkzKy7y8WUNgyBK8CHiL/sJ3dld6QTJEl/VD
UBvfEMs7K0R0Amon2ARMigSMMZ3z4cyxlXYTiWyCH74M49H2FgFoTN1guT8e+YOW3RK7L9s9JH9P
CsBInGPZTnn8NtK3r+ojO/uXae6AAH8KMLTprpop9TvJg/1O0MwN5VfItK7RPmNk07MI4WvHT8Ul
0N7f7F0zlyaEDGom3F6kHo/ZixOOGOjWPXi4QZ8p4YJMf0F/sTcp/6U0YgVRU0qwUuHT6psS3IgA
8eilQRp0QyrB1jVh/8L10jjLRnRbhpPF4D8VMJU2HIosksm7LT/ZUqyp+t6kVUQr+h0THc7qBfm6
A4c2pCEGeZvEv3VzYje14VV96y4+L2xTIMlmwJtqfOlJX303i36z+dZFN3wByyR2P1rKHxwjX3Qr
wfXYwiandDyT/syUjfsjoNTVPDpXg7oVeBRKHM+3/Fr9YoRIf4m1not5D09ppxl2aenHu1hy4ek5
7Qu7vL39fH61+5HwrqYEMrVNMi2i6xhmaccV/CYuf0VC6aS0Ve7dnDIrzvyRTBE+04so9nEcRZ0L
K/2LCcdiVeuOGvsSOIy6agfpbX6ghVeUjPNwIWX/j/r4gtDgPfvBF/l4i+UbzRvbXhS7zAuTih90
YGMWcGe872NB/OzVjKh1Fsi/QM8bqqZTDYtkjmdwnhBtDORQPirb/HD5W4KCZvQBA1l2zNS99VRo
ccqF6Cij+g/wGBHFdnr109Nt78cvfVz+s2HiCeJJtIeppK/SKRb2/V4QOW+HJLwX2qZFxs8ekBhK
FUK7ihlC6swxLkiRiC4ng7DcKI7UqIMoSpFlhzXjatNiq5VB1R+c9YprxqwM0ZMEfUSyMHXMyDAq
UMZ9E5inAA6i0HZ6s+i9df7TPXwzQdoPR/0okyJr5r9oYChkQri4C3mXe64cmY9rdWsIQA0OC5/M
smWQpVxEzrN/Fw1SrXmXiEpu3rfGV4jOuZe+xFm8vcYdxW5GazGOSfly5Fq4QLXgOMgO1RWurQhD
igY7rlmVsE8S6p3J1SQUjbz14hQsrYl9Yc+cQOARMQLvM0R7mbhOu63hIqY/OR81nTIq2vEfB4EQ
DHDLqFRWqWhSx8d3gBRCbRE6jwsmQ9hNYwBCkLJU5eti7A3qzNbnN3rvFb8XtxiD6kWgWXydeCNJ
nkAK7pkSCOtiIqWsIJUNNO5gcXgDtL62dOYnjbFj7CbJDIkzpHgFODrYwty+0sQupKN54I13HXCT
qfCF5An6te1ZP/jaVLpMBmJLJz0QD73OlLkKIg6EteUFPOWjJ8TD3rVgmUKo4qZvOuty/EawNV2W
VtT9ESH+MvjdbHEbtOeYaM0I0ixzZerOSeos391c3Mdi2JTbFPs40mf03iO6oH+ie/8fpq7OUp4e
SmOKeZUB8iyZDBAf125phBA/wwOOuL122igETUK3ZZ8lyjLqiFsBW+dhmyNR3nTX2HGXm575aC0E
rrBspeg+IvFXMqlqFRDQYVldtMrwTKr3/AkMmgq5Y00w1jYwDfJG676iCcnZrHeVbId/aBRXGvcH
4CSCfH1gib43ULo5nuZ/vV04FzsqaEAsbt+Ey6jg9EflRESKnkG/aWY/7UEftXrZ6oU5Sykis1wa
7bgb55uONV9aMu/DsBwEqWM+BfuAqWx5V/y77mG1NEmrXyLNqe5wm+Yu8IbWyZFeYtAdcqfARCBV
hDvYUtjGad2CmT7nfQoGInPIPIvTslbfFF3l8e7ESpLL2DK33/88udgKO86h4Fn3HIZhhw+/Tfmh
/sWyjUYYgmU8uxJCAQTrmJO+uEgJ8xNzSj3+8A3z+nTuavuF1VfKcXdbxupx0k2qiaBeuGK3j3Vk
sYG9IUEhg7zIluWk0tAPdb5EUAlRwFNpISFCwycDQnLCteAxE/X0GBk2m+DzZfzMVWTvry8V5e29
EM4udv9jgLat4hA/l3wWY3WRtlPowmfQ4VG4XkJEUr/FOki/jVeZ52LIUCX3OwEioVPoekcLvSY2
/97JRw5zdm8VhBX6F/dS3wn68sgd9NeKYkzfx7EnK6KONRViOS7oz1MPsn7U5+duWfeoE1NE60QT
KumaW3blNvORhxiwl2mah8GqlxvtHzUzCWnAG4nxyM7GYRyLdXMeksbwHtl9APtn6kTmMsDANk22
xEWhC6arJeAzxmKOp6th46WANLRq3urySbvSTaZhyHD7Z3KRzKqy8305BxMTXBAD6RdBDDni7pXK
KPycy3UJytZ2uyw+mNI6ydNQFtSsA0DI7UkwEDfSPSXrY9SCqZl6Sia88fMcOhWx2wLcN71Yzqm1
+3KovOTW2DxYtagH1wHSf07wvMYP6lqDUxaFbt2XR6gKyGoKxtMb1iXNgfOF620tLEwpB8lu+m8A
d/zrVRCg3oKNr22Z8h5Hs8MH/nNqziAY6+eqtEAC0ar6Bt5Ai+pIgbunqaAZkCPySEqOfm5+Vpkm
synQ7bBIEgzEyrxL+iGIQ1bJJkMuG9bHEQBX9AGRFpODM3wf8CkuZ5OWq72burr20qhYIUIRWB2N
DK8kF2/ocb+fU/o5J4j71u8UgPqOWQAOpk52e7C/6MZG0stF8juVZeYgnK5sRmPlLQJ5NFpVA3K8
i903C4OpNJfv69ENYaLV5VaemFX6uA3/nar9meQp0b8AHgLIBVZ0Gg3nV6sN3rESaPIhXZ0dc5Dp
p1UioDvuUMTK/GOjcejr6Xb1oCaFssxChJV8gsV1EuXfFOK9p5oB97VW6jeoE3ldhpWULeiHfIfi
fH1zd4ffob0bP0qHiI6sdcbXyJga/ZYp9g28tkdvkePH/62PrDsHTocgyiZg6SAamK9Pz0ZigFrN
SBCMY9EU1jl7R+er8RFeo653NW9ojbXDmG9sMf54SOgDsOAjhmttDmvrafepMeAtH06mYNPFvORN
YlGArCGZJ0xk7JnqDrUEdMb7yiLMS58UtqKKAcDuiota6zz17gdChm+zU/jIpbi8xlkVsep427TX
zAwG5brNktfma64MBiFwuNSDiR8o0RATEFC7fij3emkQpv6PF7MQ3Z2zcp60bjhlRW7j09QQbNrS
i3XkGCJr/uF0UA+d4jBOfzIyskTFuRglgBDmYLtQJH+sxKNK2Ld0p2kC6FKeVoEyxghire2jXL88
Uks0Rn3IZDhgRIa2T1+19dlr/DKd6PRGVqTkujqtvrPvMbvxRcOe5ba/NVO8gOEI+S0hFZP7lHtT
VNampgQ10UcDqjaDBTbXbjDk74mgumUrzTJJ77kVAPXiuEXpYu9V3P7ExtLvj5lP1GmK0G4sUbiP
Ekf+ZdOXhntz98QfvKFPjD+Qn54lAC3oJSwGU+tc+NZ/oNwLd9PNVSzGWq6L8HL6rRkeAHkBJGxT
Q38VSTPPMxFmhAu6OocBDtInwyGy7Tm1uTkl6Ll0hg6avNYgk5kUQthoe3wQRiJo4cbU4w+ZNo10
rokA8QWJgcAGeRDhC7RNmlgPVLzs+1K+JZVGmgnDZjo0Q/vtUz1JCKjDmxWJzG72V2kDD34sZYtQ
n7Iv4uDM1s1Yes6jawfS/AbYNhbNNoJCv6MEf9D62kDHXeaaBRNAH/95Tmc2loBkc0TRwb0JyD/6
+CZNLteme6SjBHtlpvfJTAMxWVA+T/oL05ohjdCeoqi1nbomneeqH83QHp8VhPQSuJJgCS4cp5sd
cB2CqHbSirzEMO7Mii+GvcOLxcb71bLiX0aIdj0yoZc1tZBH+d4AMI8Oj7llmgwAIH4EKQnEKNun
aLpmZ/fnkZABBmzpXOz6MPU+J5GzkY0hFQ/u/UXtBU7eIyRY+P+2EDIrwniGs3qp2m9zBnIGetxF
LiQWEBajBIEdGovXg1Dp1W3oYaHBDXcNO0mV+ceFbcYfVuZpIfhbiUuA104NSk3bM77Cnx7G3F9r
bL8vnboWUjeYowCCqEZzP8JMkfpl/HoN2ktezf3awia8mKSscmTuX10Itvf9kch00qQyHRPx2DOd
yG36RCVUdrvmvHd85CCbGBt2o1rJpHri1///qjUqNqNGV8mA813HGq0/K+4TGZs29CySHhGF34Dz
xvRBos7Ek6+IWYlQTPKQcXZ9KFOJgnxSmztgacYR0b7IjoiJP1uW6V2YkEzkINSI9t8n6AsLhwqc
UAZld/olfK5ZkRfMf+mEBnh68lGsOWjGv3f6dZ/68K+aAZQshLeRaLzIRv+4HfNWaz2wv797PTBI
zLnY8F3VZiXn7lrLL7p70PZXIeVg/e2jvJId+AojmE7daiCSgllNIV0ZaiNk1CSDzk6VAb/XJhZp
0OCgWeOWgyIOBiuy0aTvwj4a2zHwNkJYfkFky+UeZ4O7ktzb29q3HHo3SVArLXHN4xolPzy32Xpi
aMP3Xrbeaa/KSDj9HLML/hmbNC1CbE4CKvOmIPVEK235Ys7/MRIR6R8C3ZzdZ3yGyhe7Yb/6Eg9z
Fs5ybskXs7r3qkFt6RYDpFveeifb6S57MF4MyvJtlASgZ9+3An/lcL4wa4m9n/rsyXmEsgM1bzB2
HG2RDfQQH4AsjncS81ILWlWSEP8eaadJES054/gDNY+7zjE+veUm8Od+HQ06Xzhqk6uRYuVZFE+v
iczOCheEDxYYvWI0mL/Su8Cwru6NeI/+vhiC0lIovnbLmNNji6SH9EvauMnH/K6Ulz5uccsY0eiv
/VNfRhhpuIxLjtgBWBY1JtC4Ub4JHH3HiMLzmhq5PvGZqfQSP+ZcJAcL6jYeB4YUGiadF405WgOK
+u6Xb+csE5tEka8AtPyQ4mBQ9UPUt4r3B5AQt+dPgJGZUBnFBYxm2G6uEgk571nrhYhm2Fu3FTdJ
ityl35IOgvI1D8ids2LFdZEWRIYK4dWhXV3GgNaFtGzN/d/KSXFPXzcAkLz+OqdZyWIwJSByyPUc
I9waMx88mdqKBU6Y9VXNEGzpBCEJvMJdl/qho8eYxfslZbQLPqj3N8qQsJc9zbBDhhRpQd03sI+m
9PZQ0XbQMH7I/Aww3uhP7jgEXwDLbybRS+GCzGHpMP1QhUaA4+tOVoHCLjLAbTW2tGVomc2QvpzB
jgX6cKMhD4GCbxsp88Fe/s56T9knncl52+5U0h00v8KQ7dHGFAAXlzkq4FCtx8jHdPnDXmzhB3Ux
thA4Io+CLIxwbxHZ98cxxJOpPFXkNkVbITc9yFyRKHM5T+XXaOSEJMDYZByQAUUv2V78rdVLFqCg
njbyF5ek390e9P4maTyVlaRtHes4giPemdvjMqhbxkRwt7Wlj4oYDQtUAZJy/x9wDHby0s/sTlS+
Pu9eikouFfxHTZoncus9FJl4MabN2jxAIU6i8Y/8TFrbJr7Av+1af+oHHq19kEmuy1BUyPEJ39YR
Xb/Ln1XWgF1hUaK1Ktz1hzr6UE7dP7fT6pGiR82moPKl4DEThw5krFWxGHBdpde4OuExe6fSars+
1xFi40LbIT/Cs0H2RZgg6ULFAZpXkJYpeTBxwjNHMs6SfMa2eOdaSvfkRlytazWZ4ZdoFwcYRBJo
sA7YD2HYKeEwzOclH83+Q2e12WpkoWFkNWKgOnOMcrGk4416lIytgT1dUXor6k/2ECEK5yP54Aoz
UspzV6lifbHVPGDwEZw3wIzTmhEOJpKLd7wJLJFytQQ1j1RSH/mPSuIsAsdhT1W4uUavzn+tjgdH
kAl7dcTmwsIZixMJgx/6WVbmcrf3L4PEgvADXHTxOoz1bTaYtjEyDfl6C7bmd2e8wjInzMj4yZus
tnkTvKutOlbBQQJ62AHFNQmjKNh6HZMSYCeOQKmVXZ0KodMFO/Wc8e6M7ZPs7uXgo7PSivlNP8Av
7uOIpfEJRhf6PdPvdNNfOcGvg9gU3odCjzjd/9HFc+S2cfcTw25V2qlhWXX8+wK0h91JUJMQ4GJk
8g3psTinPdiQ1LpxebrLT0Rk4ko4QPwzcu7dwWzEUZ8S6QOZtOojX4l9GJHe6vUqjrhgtfocjZA6
7xLBkvvl4T9xazTSASABWDvGa+U+CLiEcBqB+GqXpV7ZD62eP4SkFb+x4UFoUtzOO+9qcT/0wyFj
7aObcCgYuBIQVQhRbrP1Ewmijhz89PuzObfaw7DdxqG/TaulIGa9h6LA85eq6MuRQ575HuuHj7NO
lTu1yPD5qOZOL3/8ovfRG33EC7s55F7OkfjW7NRw9xxk8lSFG62hlFkUp1qR4/HbB1Tq6yGkNxmc
x4wIZZD+aROLZbxQatLe09EDvyKxA+77klez8kRwQfT+Y/m8paIlBBT3QiDOs50oqQ4unLTgX3n8
E7GLtPUGKqzbmT+IFVeUgpIqMeitPj4Yd7/TLt0pHLS+O3o1odbB1SYXtzK4EYSvVVx3FiQWm4GS
uOer7bcsS6XRxouUGVx45KWAAJUdLlC/P+IJouI/dQQ/B0+hjUXgyiDSl7FiMzYmJ+Em5DnjK/Tc
8mmtkB7WAbHvz+PuDsF0vD77WFkux8diUv1EtpfQvZK+X9w7ggfEjq6YBdYQxn02JkjqsJb6A4l5
k3W4tN/aZ3dI/LTOJHY7hsLGi5CQukKohf/2g9mLxdLDHcVUHT2C74BhC4L4jKQ6G7imOQfvzOUJ
NBWUh5QUcWmlyZpEniJQt3fk1BbuCUQcFh6x17JBjJty/J/iuD+zgcfMBZ3tMxy5gAwdPw3wYY1Z
SSNi3m03fyCGQvddAx3z24E7/dRccqIEdmuWAruYnoSiiRq70ukBaj9gbUgc3fho+oMOx3VF8nqD
9SxWtGSf5hSsUocNKGNHLASprUHNCssNFv2C40+e6qwZTKRSVtHYN4IbSsdkwlYGGBQzyji0vGxy
+I84MQWwNVmSdkPsExNIut/YKxEH/302OfVP4EUW3cHcNgvdIEHVz/QvPpcnFsIW+qjtX0gYOjK2
TAO/9w7ypcQBT63oohszlcM4XY/kqZP0GpH65ZD5V5FhkREHEdhdzD27pjLF6W2ArDiKF/qWp4Ji
HjVJEzalRCz/bJRojZlCfFzCg1+rNwSP/+1LvSpSpZrdVVk96dlAihtrjSkzxl83J6+mPNmzwB0b
j8CM426fiVzoXRxyv7r+xUYA/KbADgrpJ0k1tvGrJfHz9EBHFoW80NWC6hsWufcEb4tgHzLIb2Ev
FFHSGpVaa34gLHgoizejDDnhGVPyZkS0fh2outQpiaY7p2jfFkhlK3Avs3VSZa+a2hLhSi/l2Hjz
vVRrtmr/LS0nd/kl6X+ojFBvGqDbRzuoBTpDr8TNFuEQ3Z6l7m9DApJN/JISat8yAhW/7VfTk7K6
LDePDhUpCUNuy/7td+D/ikLUq0+k4CWWsYJwsgiwd+Zs3VhY1axRJ4T3B1VwS3CSr/QtrphJRtbR
6o3eZs66nWeVlZAIMpAtPqR6n7fhBfMx+F9JnNobifzHDmHEpzqsCXdyJvNlUosD3KXHUxihx1w6
PjgKJj5l6cxKDlKARxgD9VH1MyiEB219UKuCep93TcnilZfXHlJW2nSiWf/lATSwhvKSo0zc/aF5
eFZu8hUs8dStDsgQQOpPwuQGLZVBSJjSUcjrotQyU5TsRhcAUe+OMqX7NKIvRUD8Hzao9CDh2X62
nYpdz6J8XZr40otnwGp61lp71m0uQJYiLeCEGtimhgqvjKmYljImFSVzKKuN7oaZ3MBtCaaKA8+u
aYHXFoxbTyh0yBS9Z0Zz7iHCb0nHYRDwFC+E7DpswfKOZx3qiGuRxvKwAKytdRrMaih2GRdDbu84
pL2JxMK0XwC4pL+/xj4Cat9TJ3syz52dQGCsqlu9sdVfFiIBuCGkl24e7ZPjmk9K1Ccz6IFLPgDw
skt/7rw0TwFXkbpaTZZ2Nd9kj/g7+vd2OUdwA8+DxQeVMp+0u9ti6xImooi5jDgi5SMrF+jPVXhn
gB2fzM1KFH4PVERwB/UEK+4/BhGFJjKhXw5Io7zsvR2zvHkiLmSFa74t1gY3YvI9MLXooEZSMxv0
WaS/qRuBJPypq/LbBYa6DdxdNXKwjSeyMuWCVW/U6KyTJ2qlGvJFkZ6a/Yxs0TXesIIUyVcV8AcN
kgqBXFhzjBYqxTAkCD3JNAS8MaAObLmtCpf+GkJuvyGYeYxYySzn+UMiM5o0DdGxqLnJHbCuG3yO
BSL9+DsXMvJAIYQ5OKJruPh7uvcETvJValOgH0QIgeTtRJmn+KyVB64SCrAaCv+drAM8lpawciBe
zBDt6C+ANhaP38cGlmHb/CgO05Pd3SrI0E7J/QRKxdhiEqvHgcmKCnnV0OBYNfz0hlVnDYZK/WHK
IovTjbt9l9ho6Zc6qOH6unADZfB2pZzFSh9yB+X6/rNNbffh6gGKOsjDwf8jroQfQKpPVMYddL+M
aW/zPhDthmDQCs+gpoWotZf6zc+Te0b4Hv8ROoSzjyDzbty7Onn6MrqBwMlyzQIx0Yp5m+d89zYV
FAWdjwE/v1f3acBlUX6DavzCwVleDXHZ/R+ELaXTa1Xi4woX57gtAeiOnVvuWABvjh9ADQZrvw76
0bCVnTfXtgIMD/DD2MXIKXaG3gfiTDHovqjlb8RzIbcOYs92TYjk3nBLxyhG+GvPpSYAqr+91qMd
GdJzb59s2RmTTJlMEQlnTjAJdPmPDhUwO1mqiI9n2PZW8XNm/a5/xNbf6nbmMBE2qq0hUaQdq6X0
q7HMdQ/x6KhQ6DqkATZ5rTZMMhWdAab23HkACjcqcvn8682SHjHqq/zo9ueL340vBtjJ7mAzjZ/6
9BhERiB85eVvhO/1ZrKmgYBys/A57eONhOlDNk9ZeVS518jzhky5OzT3SM30V7+FBJKU9ezixI97
vXn1ATkAdXMKhJjjITz/wOXZwk8qqL4eEn7Mz67MBRkqqvMtcvx0y1g7sDwBvo0eklq6VaiESmTC
Kw2VR5jYoyj3WVO07oXzTqaabeJngdmyrS6SWVpwNWgIsjgxmEwE5jHCDkis3FjYEO0Dkhdbw0Td
zMi6jshls2Ad0CozQTQ3n/LF9Dwv36JPmIruZ/8Yk76KewUkvcyqT30nK04HnHb41qujyN/OIyq0
PINCV3M4gXP/aUJEelJRXBdHqjjHEG4NwdDIB4Dv3ERPAAN7t49wQX9uKFzgmr7B5JcVp7vERKFH
Plz3305YnXVagikLGrPEGof0CuWbo7G2Nks9Y/MJ1ow5eFF6SVgzbjEG5CjAcimo50ZjZh20Xmth
i1AZ7o0kBwIjxZ+fVeXDRvh6INgNsb2U2C1mLDt0yvmo47xoIv2pGo+9c75IFgjmijFHeGYM6TJ4
hrAuO6jbIa8uv8Dm0QoJ5SSd/ZW82iXjaVLZrH69GiNbmZVLUjYwmSFtNr/a8s880J8qb/raU4Pe
+88QL/MJd2NFJGauozV24yXEJNzyOPjdCueI6mdUoZx6Y0pQfCefSObZrAtMq2r5cJVeOXGGU+14
U+ZCjrOYGmd0CgttfcKCrc4bWSSVJjhQwHyf/2PJl+P18F/O6QWO+cYxYCqzFKHFuQ2iIeYhESCY
02LUNYgKZm0HqEM0+Kf/t/jj6r8AkqfB2DXLlvO97Yw19aDEBzkkqVH+sBG3OuvVU4ZplnpeTb4m
36f87nmpVvZjv28azFj7VomhkU7ZXbroE5l+dkaTq0H+NXeN4veOFzTLNlEwEWPHR7w35jCW8Ys6
GiAbK/bYGpdccIKeaypWIyQBVIHLP5S6/alfWSBw3K97QyOG/fnv50SYGWAZRGJx23/7eSg1KBFg
lzvkGwSJZ6+mmcRhPbJdN5zhhQSdPkG4kQCXlccn0krc5H3XqBy+w1rs+wpScaFGlIITwiIJSU+/
Q/YxlmqYRG45uaGky6VmXEOB9ULEmkyS1c34TCd3Tl+MlEU2hfjyoh1vQq7NZ4Am5nOMu43UpGqz
XtbeWMGUyOUaAre3c2kK6uM5koW5jOM09KHpdCBINZKHIhv/fve9dyjsuuOeSWr2Vl2zowgt1eze
2uea3lgs/NK9lipIKguLQVLPhgihrUBi7tMHuJmKeJsxB1TwZ43RtvMjvYVBudqOWDUBybP1rD2/
fP5uwpuSvaD/6G8E7aQLnhWoEXgAqF3sMy6DMZJjE8Ri9INlBEOvhk9Sbkb3nI0mg1vrshROYhTW
dAE76sEVTiRXStmvWINOy5QPfI0xpXl97TDetQRQUDGnBpoJwVvKKnynXGNl9KPssdv9Sdu/xbBi
HIaexUwjDynCnY/+jam2wvDfmZoikXfpwaCdnmveYD1/SGGhMjXYa8gfuKR/x08xpFeHOf+e7rpU
RS9ztje+/YKt5ZVwzJYbC/uYQBz/o/NVjnfQwhMrMUaRiBX/dfmRmqMXyzDyy/RhUeIuGKu2H9AK
2vk3Xg1Rz4hp5nT5JFLHeu1JbLG6RPU/+70vux3bd31qjlmoP7XuQnP43E0EJKyxzpqogl3Uctqn
1jCEtbXhAZGP1I3HxaMMM51ONz2M4BRjn7IdjskBoYADHkMqv77U0mqxyWzQHnFI+pj0T0OHlE8w
6PZr8x5Fof6JwrcU2bFfHzGZFsvH4mGDHgWocGrVEALqSko5iT/S+LHZL1TMOlM5EYcJ77i1WUcg
SqMIHEqxv+iZua3sK6URISFuaIQ6aobOMgRMx+cFPagM6Mpjy01jj2N/Ma8L3jDHNS1Nchg/oJGN
11T8mbQbViad4Dh64otYNRxdWjHOmJCYUbiebOkK+FPc9RdJjP/0UkOhLQEeyOC16ks4aarwF937
MwQIZnsFKYCaaEqGvQjTIwV/6JuMpSWT2USQBPa1ZPH0Se2w8h5D3AopI4K5Y1YCq3wHOhC3Tjw7
2vCjfxey7nv7PDylkNjGz0R//gjojoYZmqtdHO1CkpRh5WqoOUUwoX48xMvXvCCyozsDUrmCPU7K
HgW5GIn+g58riOXjnb3ynNt3ZPqm7qPK6TBueqPnvcB/N51fdV4mSuevr6/ocKRfqma9JBYWGrJD
Lc0tWncdY3Y52hMkhwWlEv8vhwNJFFXv4FERS7MeLFTn1ak1+DmH+OifnAaBWZdWWBjsPcpdCoBC
SPPq9H3Tvg7ySt//iu3dElJWViK4/JKA707mv1kIqI5DWAvubJ9UOosk9/jGgWO31GeNOgEOkfLz
XBpm9PnnjaNCHovFFHqsux59Rp9wc4WCNFidJJ3JOkYcI7+USnC4ELQIVsFSqy8kGcUd8eO4pjCL
uWLJID3a3n+pdTAmji0+whtAq81vMDv4QvMETihXfKrYS61gCGPHdew0E2m2qxRB2wSVokR1o4LG
ons6znowSAmoKJ6FgohPUPa199T47S6jExd7WDuvIv0itvjYZR2K7h8t7wGD1vOJSiq8GO9P+D3S
wZwnvG9tKHlvQLin5aH0PMPmZzV6wNtoYB//NodpT0i6Z32xnvet85GVZf83z2Kom7Ugjd1dcAM9
LUNCsRObmfHTZl+Is9AepkRqfID50saVZJwZwyvRChYTZXSTEVb0+v8ddXkolDtXLHS48mSXW4jg
02vjHnf5Z8nO8UI+SwrOYcE6PnE4l+voAga0NSilvQZEm4vhw/oXuM+O8+1LBLSwJF7Tlf97cb/K
olK8wkJHNFopUa6Jt6li8R4Pr2hHWtHi6Lbw9xmF3MSgEzhbXubV623UU1kbkBhrU23MD2XVWqxh
dGjW0mKoQS1mTGJcZ3FDPWpa/Wz9cVfdwOW1DN5JygqB4szmbb/4q39K6fxkRccmLHjHuigIoaAt
ww8P3HDrhHTB4Bgty/a8VdUuYubFM/pSl3j/Swlx/JFSjKhd2TlxkIMRnJmHastmh0AHbNFuAoX0
Bnf8xs/USAx1h/4Dkjw/agvHEmioKX4Sf9WQ8LUqZ7cU9mRZFt8WUciXFygcBXk5Syv+Xkorp7m+
6YiGZiJFyJpjG39Joy1gHDW58S0wBGYC6mzWefGXl0EUp1RCRfBtZO2Jf5mHHWZ7IqcdI1gp2w6e
lPiQgsTB7PQQBeuiF0ajn82xnZruH6tTmVPlxgx7E9u+7KXYl1wl6BUr9J1Zg22JuZdedjthBsEY
+xnUsEv8oDgkKnsh5VfAkLu/B1TCmrgP6RaotBW3y7+AqI8nZ/l5X7tRkmyTTW7hKX4vZCeC5qU6
BgHe1fXpB8lmbVcM+46AIAPkB8PVcQJe93XDqJazbjWqSdYZEdguW+bY4Jg3hG1VInXvWxHE+FN1
aRRJzTLavBTy556QyPj/YwoCOorQX56uUKHkPwQy69k32RJkTJnraXoobfUwKc3czuRBWNyqtwAY
NzEGqTFXMpVNGbGXXlxFCu2x99q1tIwF7DprYJ4LvNduhhJraM8dTtbAL25gM35nL445qko6E/Ij
34K87vGc0VVelFqkOmtJhcm4P2w2Wse1tbTe8aFlHMNWHoImI0X18wOeu39pOyCDJ83hp2DBu2IM
dx1b7Z6IcNSxueI2WQelB5hOgUSxPU+r/c53Blmc1x57TYHDTl6Hy7TwEoqpLJZPXPyithL2rGIa
rzI+I/YYdMwKHFQqq3D+Bau335gUJ/30RgSqkx/fztQ8J6UcWSZ/gCkh7WdzM0H2/vEMeumhLpIr
C2tqTjJ6KqsoosHZllBqNFwxQGutbNP7zbRd2VqY0TYuiVwcdttpIVMQBnuIm2gjBiZEWWo1WufC
2oqG9/RTf7sCqoqbqBdaG8069xaftQgvOwNtnxNXGvpKKJMMq68YgSewsJLi1hXLP+GgVN4PyJk0
naJ4/Plvyq/7wkwQVEgCMzIqU3UDBnBZEdvwTASNw3YUtdtXQ5aAzxPhruF+zhNd7nQ7sAHwkb8h
ffODwaUK9xN2sbe6UhW1B2C8Jw4kLP441l0WEiN0kUi1sQxZ0EH7SdZ29kVCIDJLOkhKyIX4H0qS
ZcdAnTo8RaJ5RjKmuKEfIrz4GU1ozM6GQozaeOFz9CqDdTC7xBxIuwyteOcMWFCNEa2VBZpZZ06P
ZPeCaBm2J55aXnZFXhPcpHC92sDF5kqFtJH7OcicoVAh111VQiuMsdTU28p1eqTTwUWbpabhZ3qa
1q1BwVyG2JedtksaE6iRgoAq+eu80jmE6YMgryGah82PSjpeDHYtngy6mJLx8uvHAAF1yIjuTHW2
ImkVQx3Ul+CmS0f2ii0N4489yfz1MOHsCXDCJikA7gPCtYejsFwj60bofJVyjbRv9p7RbOBYc/5i
eapPR8UhTVmX+AkhDQNKzZyZGQTUfBXTNyENK17iEKYpF7fW1Pxz5TWBHzH9OWuY2ryULc1KFWzU
PWROnkmlGD4DZzETqh3RhwyMkxuvQ5tefAh+i2y83iEAnSb2+tKFi3LorRx8uyL9+OKfwmxM8/zD
IkUlnbv123FD3fGiy4KjoYj7EN+nyR9Ka22D6e43cUOhPWw4GJ7RiIgd+EnkcWgU+UfFrjrUHyaI
dKM9wgmSAbd+g7UR4tPOCI3EvGmlqnafvnpnpXTJEJVwFKStv2GoPGxKZeXwMJuzt8dLNed1SgRk
54jasrk5C+8NRfYQ5qiORTWDwIN0U8gr9SYbYocvgMJdd3Qw+KjOsTkw2nS0Ld3w0Knr21lyEC2k
+M9w/b+FvqP58/ZtjlXDiAfcGVbQAjM8GhvmATB1hHuOvJaYu6KTmo/pamn9lvZP7t7BBlpDEqs4
BSZt5CCzTds0kzDkFUPbYjVolCY5oxT9Pd3joLyil8nj6nPLkfkTNOaJvAwKbH6SZjx0J7hp9tQ4
rawLvkIunsfPk/z3SL17vaLplY36rhhvnNnsWLIIGaGMbQUd44Rc1sdL7oaq0y4rOLtV8fXqGioA
KzS17JhLk3dhCLV5q1eGuPciCBjo68TxHl6TITJ+s77fv43EQflmN8DG8ak7psoi86hB8wBl2yf5
TuQFpZBswvZSWvhD8vzI6GvTdAtcGYmIZTdXZ+41wi7A0PzX7jWj+yDJi5kjJGxoVuJFTbemNhvg
thJtm7YKKGRzf6Zpcxr9fvv5KYyOZJn+cEcs8/em1yqyq7InRbnUfOb1yxA63wJvYxBOpBsS96h+
JYQwdcrWoBsOb0JwQxnaj6g4BHQ8aSejBWN1i1r71ktQXlNInpf/8f6+dahjmOn9UkUGoArzwsVb
09aLlbo/l8vsjmyRTXlSEPVxhg3uHon7JVu3Rb1F7KKDSRpymNPhl8rg8pNiWMJScYw1gSb+tgFL
CMqunAWm0qstENPQckAIxb0BYmUkdNrNXXjRZp32DnBFeYnvgrgayFZWX05QVi8xPrtTjFRhRrXU
CHwgisxTgSd0OL/s/oaBdXqAhYzROv+mnLIDZNnDfUvKj/eXbKzf+gVvyViJ5XXOip2V2tAnDRCZ
MKSfcrdofAErH8fJw2ppvChWjDMBxJbtdwUsGpfb8xaRrgrbiWC+dniOnO+jIQEZjg1DU8mIHjin
LPVHaFM6fr2QVSVb88u46fWFIdVVQgPiBM8VmAgeznJ/Jf8ykiTm67UVn5qL29dXaHBNrYPnKJ+x
hQE8NF64+jM73Sj8tvdRBTlje8rtTMxhdhOY586xt5Eka0wGuoO9nFbU7fFQ8NkwcE0pxYshvAKP
xqmZX9w6Sl9CCCTs/1c+vylWegRiqkTJIB8gb251c3BIRu/72QfZmI3w20vLOz7stvKnJutGmCY/
PieYBismKZbRnW8/ARapCSwduVnc7GovlswpTIpWRUrws3AAlpFDFE2Seudugz6rLxBKIFFfMTkL
VnOr9o6hvdp0sBDBSmINu1qkX+8f5PwUWdBz8/yqCgSvVyyIRxYWrMc5mCVY4AeFY1wNgVkhSSaY
T6ZRMfNy5U9s6Q5tax3UChT0m1gIhfw/r23ckk7QbGAFtObikm5rG49d5fPxvXJVTMvswhStctIr
nzVz8r8TlEvP25U/UWJbAUWQj0wlgE29Leg7dFsq6ncprwNErztD7O6gIrFbYk9rnDdamuwPiTNJ
UkzNLueMIjFk0KIRUyQ/mYN9n+gKrRi/sLG3vE+woIqBR1lidnOnyLFQQRK0dD1soEODEQpJvE0u
aAgvWoBdqcf6pBjP/q/RjLNf2ruHAODUtcLrccTmTwADtr8VFBdaZOsKuFWExzeTiDRk8CRfm4eG
IVgXYrf3h1wBwMjamBMx1fNrLVOLQZ0k3OVTCYxx+WX4HXWSZV1VSOcBJV1TGSmiBAu8Iac/SfJL
5m8XbGH9NuwklIJLwanX2HqryEWe+WebviQphn+fOb2l2wW9ju/2iLve0HwRKMolmOsBUyc9k5oR
A5NsW2igeJh6hnjhUiHVHPMjHzL7m/t/Y8pdPno69mZYacsXVDcarBtGaXiDV+ZcavRUFtvQx7KV
9kyePs2ebOHgUeBL/QZslLJUkb5Uf5xJjnIo6XT0MU3yE1v+UflHE6wInOp3VcKfq14c54+RicgT
tR59IvSy4/KB0U73M1B3ziZzzofMnmzNZw6cVrkKB6XECZ+MQSUy16pHc8k08fzAR91Vgrm4n30y
7m1sSQjBFXQjQGnAiejZddCobMW4sJn56vriOHywLSn4XA1rU3A/YqucPVftljCjRF4TcUSXQdbc
eKLit5CuK2KBnGM6Vntf9dhJadndTDeMbzslaRTtGeE6zRLaAXk1/7dkLOUYSwHtfoMYgeZcXEqb
WX51MdfeWElyywtOj5/asmrUcqydEaxcLLkT3JKLoeXlTvhCzCTnmoIZWgQ7ISagl/kmXXKTO+Cd
vDIgijDzTojUMTcu2LuvKzc6Sy+2xwgvsLAs5zWbiLlvtEwFe6suuYyxKE004XAVna8K6OCrljIo
ePg2YVVXrB86Mn49IiUnwWnIUFZisPBIThtgh0UoNbU0lx9aXjEWpkDL3a4WNF/h06ZyRay2X4sG
P/5lQNroyaq9bVE2afZaZbqbl6+fFQxsHq9jtRrCH7R86nObOBiJXIDH1QQ7vBqb70jVBJ0fq/pw
R3LE3cPtDDaO6RuTMxr3Df7TbbJjeKbX//lnMdMtCm9DQ5jEKJVR4ayFggAHLQv7uazUzJ5244xO
ZX5m9iHZwYci+4G0t2eNJbg0rwp7bDbjYMt9O+uamaow8Grfe2RMxsreosfwoytvyI7RkyHqmrw4
KUMg94S1G49UAFg2hKJGZOHpaWxSifKkNcBpQl7I2/zjUqDczVP87T0nsPMK6AJLuFll7mgqVRMP
49ryCrV3ux5mKnwC8ccCZ4Zq1nSg5EmR6HyBN4RiPNpnrb4XSRMIdeHlq0Endy68jgaJkg8hX4cI
Ke16D4qZNJIAnUpJ9m+mj+lhpZoNOIxTUTKyZMpaBhsAmWxqnOkzarORXBKfQPbxEccu3wIL1KLq
Wq8dZXM9gM5L5lwQDJucWSMDyOD4QvPV74oOTDShUzA89afEYZGC5s9Mbo2SIwfwwtSqkcipcaLI
KGE8xJHlDe/D31YgBBMOZDjayCyxhc4tom7+cUTFeC0w5+/AkccNZgLRYEZPDw8thtSv55d1qIXD
YyIdUlCEXVVbaKBcxPXVL+TZueQGsQoPoxtYZk33ognAMBWIKUrw6C4Ym2+8HXiukF0YAFUFKgeH
wY5sBVGl15KoFxy9VKrtKTAp/GQWp5C1xtw2fxTjv0Wm+xNlOgTp5ZOsjpfrWkicz/Dz2wtr8atk
Tr9iOaEvNVr6sbi5+azKmoyx/egeviEKjk/J/5LYEfmRzko0ZUDccvqazngyRd1ftS4tQoWbhhhc
a/kiSpTOgUw9otBEzf4twICQYydcyXI04ERu+L666j2qVvR51xie2SLR3LfCtVfscVLAlbDEjzIZ
COnurkV5Oa4f37IMOBdDy4hOWjDNePpMHmNdjRI6EB6VGUV+qYdcZd0RtJYCVm2kL8ZRMgP3kVkT
V9/+8Dk8zW/uyPk5lNVbEDJ9TeSG6wQR2+tT6knNIocBG6LcP1CGigNEJ1STn8Wdxl8UUkIeE0iv
9QP5bMiR2eXn02Wk4Lg9iKOEH2KDYxTJDi7iiLeaDFgIjg5eNP0oFJcFigp5hdzC2CXcHKsAyS/1
P3zy+rQCVeGM3BHbLo38Fxr4gPDJgaLBFXrNRWh1pUBVXTR7gVqWHKsAXFQdQ/68pRxz/qglGH/w
TLA9N2N3WcBTMS0P/gBZQuMOXtwO0sd3KpERQnRnX5cKClG1/BaeGplrqIXMt5Yhk/VyIctIOHu6
K/GKaEeQgnyfdLs64EIkckehAXz7qczHFgFR8I5IbsGCbzM4o3U4oy8meVSm59UCxZe1xOpwaMJB
oUU78Bey2ulGH1668eiapbYPp0lIQDzJjcLsa08R067fe7ieHYGyHMOFmU9Lftxk0dRLmcUB9Ipz
654jlHfbFV6ACyL/8lBopNjqntDSSi1BQKusjL1VAxhXOLQ43641ClTK3GLyRN3g66xeh4mWsed9
3iYxybo/WfQVRB978vfyb0qSRmmMmNWVKhkq5ZcgX+e9A8w8KlsSuh8/QGggtMAd2v+w0ohMjZf1
5qE2jCbJuO6Cfk5q4AaF3QIkc8sLjYPCWCfGEJb2fRQPyZRzpgZkLghkUngyW9ejbHRWffCu2z4m
9MN6owK9m/B7Js+nfI12KfWYC/Ov7zwBsD0NDmQxUb8FB3dLDJXIl5jiF4H9saRpXwPqiJOPdCts
Jws7OiKwBOCJXFUeo6g0GV2hnOXa2XpITPpTCSWGEEOyNOqO070UPS34eJDYc1H4ghaDDqFD8Zxr
OLgcZeVPCvKHw2z/IyX+bxi+FDWWYR7wzUtEv/zcsbMd6ajGHi/7SchKdukF9qqE9nPqHycw9SgE
Yt7LAHBn5q7GxR/YE2AUMLNzQUXfBBAGT2jaYFIDyTYttOoA3qprrf5kMd49RQ3sXyQCVgcHJOe4
askNnFIEs8IgJcJOazX2muxWlAJQ+4RpSe3mQrZKt/MXFpg1kVpWonunf7yhkxbn2fqrmuQMGkdt
PoSmd2q6GJ6a4Ta6ZjMia9vD3qsh2VCu2+T7YKFCC9KydPMOr7oFEbxLJZnCGIVeeR3k1APVwLIp
hWalaA7EygmF45HormnJmfAFKbEs1IdBkAWayfhTyuLr8S03/frWYpM/eUQnd6B9/+7ItWeJNVGr
nPc857qqRu/8jxG3oYMCos1d+psM47Vo1J8OsBnjv0AkLvRAh4CDJH0MbTbf1RW7ffwq/8ZcE420
xZVCLetV3nAlVSz1GVmMlzmKAA5vm9b/suGcFZh6tIWXPx+mCpVnBx9uh2gMsOySIEM/zE14pgZe
FuDbd2gtXZYwfn9k4FfZJB35oMrSI3wA5TPv9NjI6+HWmRcy/EoESzcb7Em530HtSXTTN2jjBUms
jXDybT5ZN2TazMKZlKiWeFQQwW02DN9pxmMTL1/NQil9IdiE9Np601//29Q/T5J4qvADfQOTvAta
pFGPoXWW4xYKs6HUwulUmwCtXnSJu547Q4OwwkZFnZ/2CZsBzCqhxW+VO3FL+Di5cuyy9fLa+EQR
rqGT+sZRO+6yl+z/uhsJj4blhv9iB0BOZoxaV+7aPtAmEh594Pl4/FwKmF9Ix2YIIXHqKwh2al+c
SaV8VBtoVzirqN+g8/nJZsyhiFFiJoM3F8lxxd29htCAtOgpc5sge9kQZm3HcaarF76gCM3E2KR0
cm5wA6GnZe4MHqrdWnMH5EPGBdAYFOtZPgr30l5xj+SOwml1wyxxll7PvZBMXCrDoDm0ydn/lFGm
rIR25U2WL2pqJgkFKl0taEgU8nQYS7RqEBQ2CZWP5+BxkpOUD0A/rPsxUT1biVdTgJzgL4kkvbIK
2ewMa2Mns/hYcEBgdQkgHQso0o+dQFc/TZUR/P+8ufJSBPK49xfBrIT6ZfHmzERD2AAQsXN4hVMf
I1xRMaYVR/JOdgw2ESCNGU4VNzqZ46UZXPJHsITwaGDBNA5dehbS77ZqINx9GumWRsH0Xc2C9OEa
zBmYsFfx2bd+eLLArHyMI9kutIDey0IPSt/tJwqlbd/NUg+Vr4yktqAYLYQ68vaxBK2k6vajCbuX
QB4DA38VVzqxAPV2S30fggzzNO0PlEP2B1pYa/S8AzTRyTKuyoUZhw4eP9Xzo58gaUzsT4SiTpW1
wnHv95CGUl0zoitc9seBE3FkqeyB2eF1w99uepLwDXNodhMAt9WEr40AkVZPl27gTL4Csy859Bgz
8a5FaDzRJ9fvEvxYCMzyBv8AEKD92uFOTLs4JWiTfSfftOqksRVnTP5w9OadknLn3enId06FF/oy
HEdqDQUqQsQS/tz3fdj/T6EBfyp6WdXmxIbpuNoB6cwD6ytk6C3ewQitf7yJGuS7SKHQDnITeMwi
VmtXNBFJyJAbSrA3WefTawSMrLoeHJRNVt/zPG0mIocmI75170jj43DYhhhJJ3d9apHJbIWrjgFM
GdtfkY1kyZIoJzVqsxx8v5X/+HRwFQfoFGJEMGuVcnwnAjzHVAvvb60bcAccvFhFtoVJ2Fwn5zhO
hVxsSb//Ha7nabAVxIvUk3QrwrtPaas/5a1FK6Vt0VaMHISb0aTac38vxbu/fdlRRz7MhoFnPyRr
tRMde+nxq0WLHodH4tixzQdcbpyREsyJogREDYj3ANqivrdgPkbuztOeGs3yCCN8BgwxUoTdD9wM
WC6V7Gi30/Jr52TC9XvWfekeQNyVpC6yeLiQo/0sqrUFosGFmAbH0SUuqwY4hJemacCZkQ0ED24h
zEi5r3K24BvovuAnZO2WSQZldpC9y1wYVmt/2EXMfl/zeutfg62QhYwDPDpv/vQmZ3cLiwvQQUIv
Y13zFzB7AQTWo4e2MgPuP7wYfdIKfIfI65AhUulYPoQCMQ/4e7O0Wk0iArgJ74766P3s89Y8FJ3q
gh6D0efbSBTz5NSlyDHflyBK1FGUr6psgkb2VujHfNBHiL4dCH495CGW0qjNiohv5TL/jKuCtt8w
u1fuiLKem6TDm2UYv0lvc6I4e8wu+FgKUDA2Xj0EbaXbh3voB4jMg8mQAnbUo+95kMC8bl+//eRm
s7lVYj6Vf0tNpJgPnDW9NXIRijqRNlm9ee5UXI9O2ZKL95pSJNF5b0QW3vtMvaAe7W4Wmpmtp5eu
9j+JoBz0ns2LcyYd9TapWxqFx3nmKZkDH9FERSNWxmhc7oknZIR3OHiHo+SwVE0GJbpOjMvdUbmd
IqLNSsr3MC01u0/AYxZjr6dqCVeLCN+ysNSvkGUO6xxl/6G3N8DhXpxm6ljS+JKn5ouj+4iBwbdu
kuXwpW4CUBCVbmzUyF5Qz7zk1MdQlq+s5Aj0pZfJs8AHWgLvvM0dcjhGeTAAkgIYRjc2Lhun1H/P
/ys5rVH+3x0pAseP8vvFXle69HKOx9X8MtwQiMMVDgfdoDgVgbVgz6cXg9esZ8zRhL/uX5CnEzMo
CsuMCNuCoG+PmwaQcOzl4OZc9sep0YwVa3tNGS05BT+a9Q1tMUx5VNT967WIBFRYsGkmnfMeAyps
GM0hVOR8dqADysyIhrg69FgC4PBrvhgvIj50oMZvLLmTK2vZqr7asWivVBa1I4MJh9Uv9VpPwQqJ
HexQZ89D9G2TnleIgR2cZXoqqvbjEIx4EhCUYcXWZk0eg999yBYVXldNpzK8yKgsJyv2oHyrAxgK
+mvbv+Nov6r9cY1fN8PWLOlva8FbTu9M1Oep9Y2sX9FPJGpPdhi1JTKcQfwJ6rlyPsNTbuFGyhoe
4FOGped/WFkI1bFGMxDoYWptUWgm7fv5oV2mUOphgGAtUi3prsm9hBc0Rk/ooHlJAU0yd9R2VCJt
8aI6AM/zkTcfbOO/qlj/akso9TGgdPvThDmtoh5oRnQ2NTS9Hz3hmQhr+daul+L5UK4r6Cgw+99K
1KngvV/uDQZ1i1QOFYA2mVJZTq6ieGDMGTv9BBL9ecXLDNUHqXe6FZRGSY+FgrfuJjcs3nfNzfzZ
Uk/S3jpHfkyeWnsCszBHwDqszYLRwfcp4E5NyTiKnda5PfHtfLMPAqnEaTk+lUhMDoYbp86VLGTk
Let1mFIWaWggJDsOA1KeZL3yJF0cghQ6TA7uFFIDs5miG8Os1MQsQORQkyQFn032IvVfh9+scxyt
hhPstDDjSzIsl8IWSvNwGYiGkMXTmsU5Rqe3zWyDeAZ7oYZJAOk59z5l854/xt1k9os/GJrv44xm
NrD2ajeVV5rD/GJexDx2Kx2OO3DoxQ1S/s51Pd+P0e9Bz9CC19Xaw6Mm+H+KEm0qhLSPDmjCfs9E
Zp8E2I29G+1/CAf3QK9vE60DJRyii2JbBtxaxcg0IHKclp2tDog4HhklmG75A+UDJAs2Zu/2stnj
OSdS5UZ/iypkJ8xXNO9m9DOdv8lbfAezJBBlPaw9py18f5DCaWpQvoQuP6qOSTZWUnsx4WH9JuXb
cSli3HU7fAEEZGTIJqq+hbORgdKsk3vmlUlB/OBV80BojHrG+JCNC2usAZzxw3drYqK1vToj0sQp
Z7IcLJpD1M1c4IjIOyQOJSzqkSriqkLhdzeuTRutQalp+0sehvSVBsB+bULPbQhBqvu8jn6ePEZ7
77xdf5wm65ShCMxb9P+XZVfCRVRAl4DHedcD2h46teOz1T2i1Y5AL08c4M/8jEoyGBPgae78quOG
au94c0WDmzSZ1+gXbtf1mwvqfX1ACAupCaDX/el0Nmvlo47TaB6xyrtyuCeJG9YH1p4U4OXybmLd
fnAZxzJ9VEoCkJ9kJb+071Q7n3Vfkp5Ckvw3nkb8yeVtRkZvFUleO0ZNib3Jj3ual8Ndp7lHpQY8
dXStXyqwa0z4qFfbQb7yuGbu0dMGT0vjONacyWUQIGKE3Ifn69MMpmlYtxvtFFq3JWEitkyOR48k
/xZavoEQR4YfEgmmWLA9FnBFVQfzHb+du94j5Z18zNnwxOcjvFr2El9cCG1TZNBbGpj3b7IODIMR
pLRm/gMHWRN5G9u3vmY4tRfCpkXX2D4SPUaND0spZ+AV+2Zc6EevpETIVqy57wxPdffw8k15UbRK
1TVhtHVF1Aq0lP0AoiEar41dprDtonzyCNWKBCYDivk6phOE8yIS5WJ/LrfWJdtniFaz53MmZ/GD
axzLR2RGQIqX1d/w/kvXMumNhKTAUkw6DnB+mLMkRNnU4K371AnKdb/6PVNhD/x5IJ22n62eAF6Q
YLXy8h2CiRL4QWf52wUlzEJuWE2cLXVyhj3KP1HGgU9/ZPnlq60B8wiSenbuxlPyN6CdjsD9OIE/
8QGd8hYaeN63PSMkrK2kkifJ7qZ1rjbyZeVeOt1o4MyJcdq/EyeVaTYRKTCpmyntKEweBlqxcawq
H33gKnno78HjDqmbWrIIgt1bGWgXKsyP7sHa5apQS/GhxEMb7R200ZcP634kDIR+XSgnujBRVJjM
3aE7Mv4vlikexlJMUGAjBwxAhD3Wv1VyYTDACR3Pa8PrALlU/oiID7cTkwpOF+LTobcuj9CovwJQ
a8S63i7HVRYcLMwEe73PgXTZh6PYNjtZAJaTlNkCwBgKm5xKgB0QhA9tyqF+FRC58OR7kouFuQ/X
ibmKXJDhnsN8kYegCnPltbExcXmc5pM0HVaEfXot/pfSYsoh5lne9cBNDS36VujhwwXe2lFuZJ6f
LZZGfon1JtjnjS0rQMXFy/MdK0B+c60tG1WGEswRC5cyOhnGR7qULgOAIJeyH4UVGmdN1UsJi5om
PJWDOCFW/nQijRXANkpKjhN+8VzEbDvKfCGHCrulPYZu7cdYBf0GbGtFp4JInhRSNaBKOcDluiYc
GSCKUPclJPbYLI53iz6wUOYgM5NlMPH1m9AwbgTeZ3hxlk61LWgDaX8EMhyJRiLa7xbFDFo/FLpe
7Xlji9vMZJdiOkDoe3A7Hu9oKuLxIe7tRSa95pnPGwhTde8OemOmmEdlLzK23Ga4qpofRL8tqsqI
084cfszWHhBEMYNwEN0oG7U1Lf6USGnxmFVoatLVbHbMNF0bbHrnjjrOu0svJsYdDJ18MN66/G7S
Hp51ZRzU4GfmoH4a+Tn2G95Zzii7nX4KwzxVeFRvzMQcGtpzKrfyKM9T9CzkA3EDX5ptkmV6su5N
nCSJjq/QnIz+ZfsD+IWCaZxsjd6njurkOM2AOYN0PuErgRLzMCnPjsOp8PVHo+ZEWOqPmUrWm1y0
NgGao97ySWHffAmL/EI9UFp7fLWcwcNZhYAvSyRqTT8LkkvCMnWNwFc12prFvsTa3ejW0T2dF3Tq
GQCVoP9GcGLJuNScVPa7tdAp4TOVvrtVtSBZH1IHJuCOF87qbtzxqe63vL1QPFaw/rVqYwPRMHPn
GulAIe7goHkCrPlRIBqZloBPFtrdiV3hG01Gkth33tJ3kzTI33b09dsLem7osSS7K2rj0nYFbioR
7Uz2uJDCnUOA2wbfrS0tIJGa7IyIQDw0nAWtFtSotrW7uxR9kNeW2ubfWirjNaRfqGcVCpWBdsiR
B1HydYbIwffaDX0ZTNIVSRKedlsMsmhxvqyNdgxQcfJAWvDxHfPhb6UVS4oFbG/42U8hodDdrXux
2CJDce0VQ+qFjDzdebR44jK9t7H1a1AYvOfG+xeVBO0bCU/uW/z9VlOT5xATT8wbrWISQI1SA6Vv
Z35wwD+3tlcb+gn/29r5Qr1qGn1++9SxvT3u9kZgP5pNJtgXDxKxaRBI5MB1Q/zQAXPUKD5nWlHl
RPrXDBc/TZMh91tzQ00Viv4mzGu8w0gMyP6NKI+f2m1YrAPuh6aM3SAPnK/z3NSTeSnhm0t341ji
fZwo/KzB4K3oqXpWTBk76n/GMwBQjvqGehmuY3Isfvn+Z1fk55GoMB3EdugT8r2RPcCgoBzTDqA+
Fy1rIojQmYWbT9od+kZyakUwpKD3aylvRFhKRvK79Fd1p/bG+24xpt0zWA7W0lXg2x3QF2z+dxCj
h78GHidXa9F0eQmBoFW9MVFL0yvbv9SZ3zb6LaBHt3P8GZneK/q4mmEtadeXRnCKKwq9mrDtNCc8
SFT+GB7iOKTxVz8nOiV1YcB9sl6o6xFYhmZSynyPQsP+nWGqydtwotVtvKk2Fv1CN3iB9nhx3W2c
NbosXF3+uB4mbmtWjvv/FZevt2TIqWqaAPcLLFStGUvlb7gNuQdoSdC59wppi5Qgp71O1ITzWcrz
UitWTVHBSAm4lkDIn8+AIc5t4Ftdjfdgbo7A2L8pTnDUcyfc/1+dlkQYXh+Zi5gbpZeRUNqyqBMK
i0BT1BlCQKrLknMGVFm45Of5Cr3eCMpcQtSv1FDZXllhBkd3cus6KkQdQ4UuCLuDuLc/AFLEU0fM
+GMDc/GxswTNhiYT2nTVP1AufIQBj3KrKxJasHMPgLQLJzuHQMrB3OQMR3hoYmVs9Zd9SwM6+eiA
WgFIEav8Y77So78Yr2QxMOPR+drtg4gJ6WP0TvgpcuwrnYmZSGe404Bp1fjloO1T4aqpW9gnmPKR
hVKnr6QxCuESsz2EPLUIknV7VmrzFkq6iFgNNEpB3UB2mtJ+cOVn7PZUMaxkgot7s5NLXgDKBFqH
zGCU9iDJHgz1ZQxkaM7zKMrd105NoCd4uk/R0OZLlfqZmRQp0fnqXJWOOqUBaxv6rQmM0UU/2dCu
/Vn4k2NTrnESt/H2CDWB/PmmGYwua0iJRsczTzWgK/lFKnQC/PKoURroq9NriZhkJJrqvxQuJ8nB
AAXWMcytoLiwzbVwySZAOyFOKutHiDv+AjEKKR9Wn6he9iW1XpiUVqpdzPjUBPLOst+ibGjspR/t
C0/8KFa5kQw7lVnaJmxJsvICd8a970vpMBKk3JoMG8qXRe5zN2u21RGIBfxUT/vhvCpmrhb7PpjW
V6Y7Pw08PivHK+/9mrnU+Ztud0gefIagRXQ/M3iIHHqh91P3sUrA097tWWVCz64xe/NgSqcC6ttT
/b/m0BcBymr65s8xmhj/ixtDtg+hcrfRZXbKP9uhSUQt8roDHwocPDz6b7ppM8zFW7lKwrXkqZOl
eptfv3lnbZm/qlBGVR4H/GndjjIXTklXaF5UDaQPQlmOZRuC3+W2qpo2KUHkP6UfSLpXyDxASiZq
P6YXCdpuXEGSd5bzhEOSnXgaMz/raiiUAkDPyfvh8OAN8FAwjd/4gEqSQLmfpQPizzcb5fW+EAfg
Bcp6TwZhbFCNDzgWQa9P1+kLXJjjgkZ+ZbQwx8Cmp3aKvHyQIxpAedosD96B67rPuuQoL5QGJqpn
6kv2l0QDDiVuWp34FaT0ycGAEvIUs0OyxV5xu/GQzxZZ0z0hd8xjtaWqMoDrhv8fo930JOBL3val
+D0gLr+PB5wE3suVI3PAR4t/h+8da2g7bRzOdGS9C8wIBAToVKsWgTJosemKKoaxAWZ6+mbXjnOT
0eFSXw9FNpYWC1wKlVTf+7PDahnb/dFJJIba/9QtcaJJOIQMAWKa24NkAeIUALoFdNu27DYu25pK
PmA9/uzZnDQwtPOTmw8CFcCQYnx7MzQ9xIQOugoT9HU6cLaBTdPvsSq7AFkvfKFXtCMh+GZkKNP5
DyiWmbmvWF6PFr8hnYJemg+5jt3SAGUQRj6mb+QYxh+uB1+IcFDjHScb39MX6bjjfIPLvcir1tic
/DNEHgplQAmKkZL+M4cugw7gSI9e2TktMuisiguNoaDyBjD+bJ52wzrVy/fRKchu8pfKaDvy0jWF
F4hw0dG9aL6lLLhlHk4zndtzi25Pje5oi9dbx/mmI9sP7iq4mFMYz37x7zsnIvRh2kpmHR3YxXMt
Ev/mjGV/yRRe9cs/6WSDfgtbcWNuoXSMNW79P58B+5DkBzy9aQB1N+HpGbM2Eepao+0ptxPktKkI
sWzm4TVZPfaMBLosUxQznHIflYva2sQKjRnb9Dw1gsujauw/AxMwqYvEKLUqu3yCCpBxaHh2TGjX
4j16l8vduG7+u3PHWeF8OwQb79hfCi0GUqFIefnQZplAI4TGe4U2U0teLua2ifYhdGgTFRkdrHvY
ukescPg4o+64gl4rPQubJlwTgvWkIck3Wp4vQMf6Wi5PMuQ9Wfz6ewForI+RkVPC35DSv9yDTINU
VfxuzX9Rh9w9UGP4CYsvNs1+60k3sRBjXt+1s9gus5l1Mfle3AW6cq4KS+pwVXWOSQbRSFYsTSXZ
0h87+Oxbli/75Y/8yShzlBgdrWIwn58JOo3OBqNpdHYgVydw/aW9P0WB9RBcD2G7zXZraoZVLSyr
0f3j8eBBZAkYxTpL1A9b/kT9bZp0w97tY0p9ls7jG/JjMfdMUc85ZEmItzUTtP0yABiXLf6f0QsC
6yk0Zk7U+nLxjd7z2W6a7g05cqPo4J2zCMXuDjqyxvK6OBakMVAhTgoACGhp4SjswJnoPah6X4Yr
WWACMiQQT5xndRHKVSNvs/E3hvRRgkUwDEl0Li2iXdyNlSpIIMwKfeE4C9E0RhMuFmM8q3yiNe1c
zJqAZb8NMgyyKtlC4W+c5RZmG7xAxEQu0NpnuOzL6FnprSj4XzcR5dgYS7JfRK1ZubU0MfFgyxta
ZIQYfa4XH7Ixuq5BSYlOhlNiaDIc5PLtA4ihwTVa/l0Ee16e0aYc3txUqWXu1Yc8pxOGR84fvX8d
SPB+9sIk/28oWbiq3OX1GDXE+WDQ1U2A6Kaak7WUWhAlnzD3tvgOJXzBnzyOx0HgojF3YInpv2+F
WVyOKZxgDRlehNiLiOrAo+JtZd0Okpt0VZrui5ktB2psPmDHQRK9lbdo3pENvGRPhd70KUiJwBFw
RpzN66VEZ62uj+tp2PNpC7c7LBY9iTz3zd97Cxmzg0Mh/aBcGj62DEyznlTosxpBIcZ7Zm3p/E9k
ouahy4A3cClfpsYMplVGnbUGiU32cLyCvnI8mspRUN2HbzDbY7YlDLrC/EqWsIKGaULpD4nS50KL
kw5ChdkEBg1Ml1yKpw7x3/dsXkX2VZ7PTqrmmrNXdct2wTI+j+lzJw/iPuRN3PZgEvbZe2w0l7Gk
2cULL6pTBIC0JH6K9f5VI1OfVDF4rEhs1/elHL2DbfeFGGxqmtPmMpCgWjVlB+HN8OFjiVfS2RlD
5VOb33CayNAlsAVKGHpAF2tkzmOgSh628MZLuZJM368FVCyO7zGVk+VBFsrlOkepLhp47UhBWMS/
zK+ZxwHDd/iTWO/XoqETv5bAYs4yno3VX7XIRTqCkultIaENHSFRfb7yAJi0oE6ZjmVOE6Fq+KHh
XdVJ5JlRUWU5ScpXIG9r+McF5pFfVMq8WP+6RdllK2xX4Vw6Cg4D/u8oRhYVYcyWyW+dzuGQgOzV
mD8uHo2Qf/MgAg3bvyGbFxo4ggTD41cF6aQvH8WM1QZl4jVAhPIfTWtK63yrdReWRGAJugVt7xGk
u4Ay/cIfgoruOELbXJ1PMxU24GthZnaUnPGakLZPvBJqhu6mraFqpKV1lYFBqcmzPuN+6fYEW2UD
Ngej1PlyYJk5HfEQatuaqK/RT4G9N3ie9JQHMA84auygI7tSP7AlStxeMIPWDMzON+XamHbGeyMt
4rHR+JD/bAN0ksSrP46X3OhxS14PBkI4HPJa9JFesIM4TeQ5CES38IVvyLOT9+1d3lCxc0IRfzj6
1eU4hgy4lVdIMG/pZ7HSAY6U0xF+b6WavOJYru3vuZ+ocB9LdTgGjWsF0/SqtHD7esUv79CUs7lC
s2kdxflcysF2LA32f6o0zEYUgX8lxy51Yr59tp4d/ah+W79TH0E4I1KLMobNCT52FiIyH8tTuqLW
4naAZjWEWp5qvatyocyol0FLBQ/jdW0y8u4KPqrJz6ONzJCBJfl7cZRTAet6HtEMmaQG/iLrIQ1Y
8XRr+iS86aBoAuhYLSMmdGyoPI4Qnz5D+IzZppx8xU1U3P/Znb9mIwn0OJf0eAvxO7hSde1Iu9H5
JIBU3DpyVyTVMglEKAeQIs0VP1LmFXEWGQ88bmeHyG1t7SNcp+gNqjXJk84EXWhWTjovlL5wTjUl
Q1FSXKxSWnw3YZUxLhhkdQEYQfoYj9Z2osXdRKaI74i/sUlJ75N8jGYvqo1Lpe+5RPLvSVWpKsmd
CbDywQzz/tP9GEU8tCNi3Ynfl3gl+c82lxU3LHuvxcK7TncRFYgouCHAl2eOZTrfgJg81cIth7YH
Xu2wWMy44cpCMnBoLZVx2+eFKTcPraSQV45KnCwO9YqpntJbCU2gAtkZLgnB2WxsyKEsx5gRiAxY
l1osxN4Yw/T/XDzJDtG0itWd88TYQmq51GOND3KDlhvL7waytqACYygiDAhMYXmSjwykXJdh+kD7
vJyXKgOqsL4+Nxj+zQfqui+SqZI3dAnsYSFGuHE2OsKTqReFNgYJ53UYdX6oCv/N/b5s34/uome+
m7YrFIa0nH3UC6QXdVDjbmHM+guqUjTJ8YSiKYpQR6eJt1NBy5xn89cxENVkd9OXdSaF8QBOMgbC
wkPwn3/MtMKK6hIlueoLi9UQ2az2JecQP5dsnNozR3wJDWXdXn57RAfnql/NabQn2t9r1nNH1Rh0
53fRVINEb1U01vPQBznk/27UnPGpheXok8Vrrmgs6Zrfk7LRJROb4waX5MQEU56/nlXXEgjrm/sh
AlJZhFRVe4LpwXi3B846a79OC9Ue16odCt61s1VEylDgI25VKpg9/dE9x+sRfdGYoVO5EtWfd8bp
athZi3tV6ct3IKxb9BJdWRr+CwlZ8dzIW9lIZxueg91jAWJK6ooVL2YEf0vCqBELrkZQtyvHR660
DOyxcJV4+AmAxkwdZJhJNbFCTKg3DhzgFzwOfKpDQ4KW7sXNAYAuP+FarWve3TYo1X3knIluUnkw
TL1JD+T18yScodTz/xvwao2yw/FP0doc+HUHuOKwh7Yi95TUoeNLHLBFlZHXuwWWsgJfJuyrRwgE
ccxWYDcnGCwyfCpoYHAd1Y2bdNheXVYn+mSgN+OuilU8McgJKEISzIKlpC97jKmfqZaq5gJ23VAl
EcBmJq61N9OHPeqlInSGXrgtDB6q5mI5BpYqHgOY4x2T74EoOrxMdvnxuaYjJBSBuYiKwkttvXqz
oRoNXukusLw3wWJncaFQLPeoUgTBffpB6g7VhL91WI2mJlAXitF0uoIdZe/HEAl4wgn4m+n6bQUN
cgfJgfnzoCL6cNFOKAhdporPSzrjEK0kTBLxHB/+RF1uiwAjT2TUIDBWNDl186iMZgsQMId232IZ
Ay1BL2eRefTehBZNPTMNlGZYzNZcvur8XMyimVxauq22VTw38q/fgnf3YFLiZ/hva/aOKmw1h194
kMINmJ4E75NA1HozRIZbnL/AjXbIdwu7pwDuXMPaLLhpRUnXAjzU0QcuV78k8j8S7nbUFmZbqsjx
9RQovtxgk+ROqzhW1gpXE5pJhWQ+F3ribv4Rda8GTiekF5Z0vSxZ2oOZ5jlyZYLVAezke5Gd4b5A
ViLFlPFz2jdjHP3mDRA4adntjS4vrFnG19soLUkf5h80z5D/m5bNYZM+elgi2IlV+t7SdjVwjuW9
MyEBK/ckCooLiJIKg9zUCHlKpJ3V2XxyeAes4eMpn4ZizGQX0/7uAg/BGpJj75hpEiqeUj2np68D
qpgfsVIukMn6/0ZmVG3fC4xz5WO+OJP/VTOkgLqDF8qsTUwbS6YqCiY+vpVIvlwMJA7SALA/xWk3
Io+APjLnOxIy0MHEv8TvEWzfto1p28br8TMd4doWC6RVjr0rOLHu+LNgwYkr5I7LPpna9YjkCqSz
07wjgE4Bpy0Sjz2l3YoxNFhIbZMWAAvB+koJW1+hEayb4jItt/SwnhWH4EeSTFqtyLRztus3xyzn
ogJZbEiS6MAic9CX3Vsafcg3LrM1wSoFopaepBK+Up3CAJrvIeVPjpnhtm4dd/rC7OkCS8d79Jy3
JXiuduUvF/0lVS7irqB0C87sUtolCO8/TZm1P55dvydkG90uA+GgTfNU7Ct3og7jOSTsHTL03FMK
VLzOyyYMOdeZwORRQrVBWgqzjBvphU8rgGSxlFoMDuftOuqOL7nwNMRN1/PS61KoRwEcm5/NUqKy
Wj2TROq79CS10V9GDNZqSVWsK60PXi9w0RmZPQITIkPrkZm+/gfwV9GHODnnEqQ7J7+XbcqmaD2+
CHFz92+7MDe7mJpQPES8Fiysfu9RvEoJGqlvDxJQhQe2dQ6fabIhqkqS8Xzs1nYkwj/Dtoz0/DTq
fWCNItDpKHPwssuS37JzYfaDpC0H5FghQSslZZB7JdtmiY3rwD6oF8+zMcppShsVT3blrF4XEbZp
5ZcGBHehadtO4Z2wPf8DIRu3ZiVg8Jhx+XqXFJ/37cP7YmM0j20UCwDhtKO0/xZFgTffsdhom0iq
maN3D5n2swCA2eJfoZgHtrmPJB08Wi7rIbTtHe1mBqc2YBMzB+qMRCSpV3jzonEamprtIo7l5zkW
0+I8ETikQ473QB0JlgV8G++BkUL/kOaNgypwPbMaL6AEHr32fCytoTXqi1m9IVKFYzvJ2+R5LD0x
291i5wJYRHe9DMvwUJkGdWcEVtuLP83xBFy1WCELcO8zdZMpAOQxsd4xFgvHS913JNnk9RE8UJ26
PFDt3Vb8AMf7YjwElAxMRKStx0ZZ3Pckim0Y1h0pGdZkivVpeQpxjV0Tg0qA7JMUV1DBVXbI91oT
fsd0Z43VcwB6oqpGEQYhuyLzuJfA4LY5vZHK1jdAfh0FDo8lp/ZfF2E+kfiUN09NQWibWIDSovKn
qQ7GmX7DtTNtVpsL7boyW+5Zz5ByhfCPJuCUmgfWjIPTrXnFE2I1XM4sFytbFx8fR42Dv11tvDQK
DfByH70yviQE0S02GdAA1vf8ICJpInt7jBC23VyYua1/8UE8DcH7y4i8zstBWYBvZ3LnyBaNtTkM
G0iroIYMRqXt+WurI8gwYsFypcrc8Pyg8EbIteLTR1VcrbQZaowB0KDe7HNe5jZbaQQIPefrWZ40
peMmObw5oUSj/WnUs1D/trrvmRn/tY6Mkldzt80XdKacvVec33e1VcqtUaqptdIylptGD2zEDotA
3Xgnmwa6EBZbnJjseOlCjzi8OWoGZ/IDjBqrjde1JgZ16hMyGshyu26RJk6GGnqwEXgn1yOExZDJ
GOE0kQ5HqUyiTOZ1gfS2dwjkOaoQ/aqbTJL3I/GajtDz2JmA0AEkiX9bFobqK+5cOxGqvMcZ+EbN
cYqUvrN8FmtRaGoUjTcXk6Hy4bE2KgMNmxKXt+zy/K3Nosxkjv9JhIrilAjuTx1HgJxRAUyt202g
AOI4ApnRr6WzpFBoU75iy5yT6ZqLENJ4ErPMmQyWAwHibHBbKekTKjNiarLsz/sZbhrwl5ryZT4e
MAFuMrN6S5AKBtn4F9Q0+WDhp5FHf6cuYjf13fXWxveqPj0axYWg2tuVR3oNmmxE55JXHpVpBcB1
o4M3WAWKgtzL5zSw++oI1UwwvWPCVjUoXdzBkbgeTCxTeVi/0trYlJVNVgC4hj2IHKqazIPzap5P
TpHTwn2ksFKyWy23jQxT2pQOg3eLe3Hi/Vls7ftfKoyaPh8R5ttKaY883ZF9p0uoHaZFNoB/0d+H
gSJf/oeV8WQrBxaKr9k5DPikkSbDrIlDHWccjVMkhBFGvFhhkKnZbUgmioHJNpCoHUpwHX1zv+Fd
57hjJkA0p0hzeAWH9zse63+dSK9u6HmuKF73rAEUz/Xg7GrA2MNbuRh5xjwf/fwDH/WsDPlprT+p
+PVcQRLyiV3iEF6gvR9DoHjpelB6b0ZQGQFBFEbwDSUDRrrw5r8JMhILHw91FjR171pho9gk0d7Q
li9aK+vRPBlpU907izeBU0Q/tpU4PbBiJnuOaZyxDdFzx++7S2YYnZkUChol9DrrDuMIZtcBFRjo
YGJeRR3E6mxopKxmXk57NL/kK+OzoNQJ7fgcKcrGLXSPd07LvaqFYamrlA5DgHpAcDvpAFy+e3X0
5p9zqhR1FbVbk8yLMyWc0HDI3Ii6I3NzgFFpakHaQwNhuu8vxwLvCCiwEFxRSJL8JKh0ZIxVqr+O
a9AL/dQC+cP9a5xaEOCQwUh358nn1+Cgjxti+Y5UycKGCKK5uvp4wBHkz1RvYb7PFcMMjbqQVNq9
E2yu4u5cdlptfa19uLVUfmUFR9fv8PiF0scDXj6Vh25+evSWP49oMF4eJSQZXojpaEJrcdmKLwoB
W7dQNwKbvicX3Sj8ClDYgJ5UZOj3bkG1jrejy2l2W+4cKBcvNguCFkF197TyTy2YDzuQIWVtaHoZ
WS3CXX1PW+Q7ncBEKZ13GZEMb3IFtlZKb+bTAOSaf2Qb5Oq+kYHqiLRElurGz+WvIkcZIEe6/pwf
rdSIuEs/DeKkp9FUSrROKqpW2k/ot+pSfJmeyl90wYWZ9kbw0GRgz2SDxwOy/Ixu99xJ7t+3C+aw
QLEsnHi8xhCWe9uRAIn5y+ooXkYppasehxYoHulfcaaY50s7g8dcvJfhyPbGDPGDjPjAtTgEJw8h
PzCnJqgGzfne9byR8eUnNepoW96lhMUJ18cUxaLnXhlyWVEy/UAbIdcPqyyTviBYUpapEchgZeqg
ADBC9mdodyCfUJRAJxO2MGag9fxdsxJbmIfup0hsODTW9UbG9wSSz5abfpl1wOByCKvZ1rxw0Di+
93nIZi+szPRXAIUbKyjDaMbaXtq6N7Fgz7ivhw0EAGrKcXwlsz9hfNws6jndpfRuDeeRL84td8ht
9UH3hRVkCH7ICZmmG2ui2OEYiHaaH9g03ppxJLv1eIgkJWQtL/5xVSAv+gix2WvMedSJGeFAaWpt
6WDe8oT3qtd0tbR43GJ877M4DIHwqxxcN9u237VNOysu4agV36OmMl1PJaY+gAQiDgsWJfZzmDNY
RiQMCK69t6QpwHV8nSQ20U9KWICyxsOliC1c6xfnAOh7ypn3/s+mGTHhkvYt0ZzUisOmP1wOqK7C
Z9LmLsb9dew1d9ZtuokHi+NYpwTcIsRfVw83XsqfKenlyscocNfSXqBrYKDQ8Hk35NR2TcfesCsO
rb6FieHV/bVgnGmGqAgGCyqD24zma0SzzmEdW0vtXNaqV+wEzduvrw6NrKJMZYmPhcdm9xEtzJQ2
+M8AIQbAe/5hkj4c3PJiOijzMnnEMQHjddzwwfaU/HzNyDmDPYKUqOZdsgy/XXobEDCU5lDSAnoh
o147fGwyLD0HTtXalPt8vCzy+z8oiU0cZag/XufQAniSCVWGXerbJKpv+GQ5xZRtJZwDh0n1XoQB
SZ+DNuamOodm6pVS46+t269hmueI4bgJXofdgS5t8ef/MfooeL97+5i1/i06QA6JnTJAUYd94fZD
gsXdyIxAisCJ2rpI2x0A+U5iuyAWeD1UEzfLkevOoz9+tQbKvj13KMbc3iTrwzfW2z2ngK//X0w9
kevT2YC5rwHABtzFB3kDDeh+dCy4hNg/J0gYTYM1vy6eMLaH3Yf5/QT3IamvvnYL7CY6fQBm7AK4
lgrxs5Pd0aN7ExcEaNVILZqjbSYDTCME9KF5en/Hsof5XILoxFqA76i9hqOIJZDs5JVoNt7/hwUd
boOJ0teDqVzEMn5hx+lWnKpiroLBzjcTL0vYLK4Cn3/dTYmR/8xKCj+6IMuJ0/ZXsRpz7vkuN8ZD
3nX7uEtuDU3Pho3MPpsJFwqNTlGHRrOIwDCaZFx2zoxjG68b7FtE12PAsnKAGFclknJVHnzGOn2D
Kr8byPugFoj17m+RcLxnIYq6zha9nnhib70rfwk9IQ78nFV4POwiCuE1/41hHwxTYt86BT+J82Uz
Fxak7NFFtuz5OjUteGj7OxrFmhb16h8JezOS/TnOIc3SPpB82u/IAbOsfAzu2mVZyvJTYwyv2JZn
oVh5zUiwJUzQ48D/W5NRw4nEkXQ4L9moiWcZYGleUdVX5C8bC7qPA6C5HnkzZCfTSEfTfvFW+Zxo
E3KQ3MODBn0vSGsLnCEZBY/lHvWmrkh2tQkvlvs8kdG9oFt2cJ1Aa2R1WIbQj6XJqNo1rnxOaDTt
CCIBgqGZVLYRFkxhlxjeYkGa5rG1+tIlo6e3GOqx6kBER4cCTwV7h1su8Nr5qAVguQIh0Y3mJ7Fi
SHwm5cZHDoPuiTd3rh65TKmrmwFZJXS3djWkAiAA/fzYIUqrPUbaccfuxSYSM5ezh6680dOeWCd3
OjUphFJNv0oeO3NSchqModFroFEzl0YjPAfsQRHWdEAGNyPXByI0N5jA4XvNd9tD9W5pBzAH4AEK
HcJpdb0loTWaUAXYV0AZYjiyb14u75eUxlmLGvd2oZJNdvthTZ1J1p1Imtw0fWsJIWAxb+HE+9wG
3cRKgF2gpUZ1U1HdYcFHhPoA/Ppqd35nwKKaGdjGvhQkiXaxTczt4aZ9hSqxw1Mk/ZgkMzbTwtrn
/JqVjkWk535BXfh7l9W/Ohc0Wm8CRCqKbaMTSPwH5f9JIjvD13gQBI31Bko/OSNa9BFtqynTofHb
/ozwxJUzI5GMEU9rkpP6Mp88l3UBJ8kt2W5Rlu6nIh0X44SZRqH1D7ezaGHTO+Qsv76jSWgFDPXb
V4ielGmR2C49LPCOlLbZLldWbBhkofoKMgAsSrviXI6ikyivyQiU7bDqCmyYotDkCSRFovu+RREJ
WnTLveNy8fHys+PYhvPCAK3luQizZEspUdQtAMJ846d2Ggs5Ze3YwpVPaNkQUJZDCy7plpBGvBY+
TNu6lFbvsZh88aTEN16hNFTJ0eVF0QkE+suaSmq8imQoLJMwiFJtxV2+gL/6NorFcDju5VieI1hA
HrTbZ24fKxiY4xlFAobyLsIvja3jbh7tFyVLjW60NnejsFmu9IEQMRl91jDbLHj5BGCXKGvByEHb
eVdOaBlqS+y1RDIhwqpYgem8ljmSrXzL4cxJhCm/eWt5o3mZxiZHoM9e6bzIhrJ8s5h50IjOjHNe
5I5dxNNHakYpFAil6rEZIvxxjC1EhmbdPMgzBM43Qee6ZWIF7J0JfgVy1Ip+6FA9270/DCU2Nycx
dr65wJl9Jd3TLkGsAd/hhL+uZDD8Sw3veTEKwpoPWRKfqAUgBrgT6HdScg1G/NXm0gIlWfB021W1
Ju0mqJpUn1cAXxuMIIiGQN2rcGbDP6UdTx7cKfqb0UUu8dpP6I7sJULVN007wSCSdcTol8QPDUW3
Wht91sSrHUrhFlnYAFNQHFX6bFBiAlG9ApLKYAhhj0N7Jcl/jZG+sy/FkokMrx06nutxNzKS4Uac
nMBaIZVW4yWSTesVvxEoSP44WyWy8HcLeaFfUhd47YR9gKLo5eAcMuqej2ZqeVhsUfosbDeKN1+/
UFsd22485iCJrjLqTCwXAmOD1xDKsXumlMyU4ihIGQYyTNPUu0IKW/wDziN3EcVIwGCoLh4v+7RI
mYHObtz8tvJa1Eh06OR7xtHaHRiLgR4Wa0RFjYVSGlF4tzzED5+y1s4rhgXq5Lq2OOqXBdLP+x8e
wETrDNpNuqL/w1z8aHegxBM2hBxuWqSY+iIOtTnkU8VItGUJ0x4H7yYrl2S6LnHzJHef1S1GPpZH
GAMpSr4YIny0R3ufmlF/ao5GVPpHYVq4elQQ9LL0DjP5SJ/z0fZqDXJRmeycb/IMEVolqJsWzwir
cbkxeIiSpQJOsKLWyS9bo/lFTMuiBEQ9rh52ZLrv69vIza5i+4yzrhDnEpRALqi2UqcFuHYz6YAY
XnKZw//qIELRZ7BSh2YPgk7pVPkjZb74LY+DSz++YmyV7Jl4h4YssP7R3J8Y+/1JLIi0UwWFsxzt
7e9BXFH8nKLB7N6L6e5S/LCO/49NDsJl2M/8WBxFk+iOm8QclknExNSESrBJQNzpMol1YM+G8RJO
ThiBuqTAZwACQdUgWGyePophuQs+YIIIiMr0kRAke951wGcSJeR4OceKnBRT2ibHciuDOCGSGAQb
eLIN6cNSxHRjSxlWyqnK6fnT0yqzihlHidpys99KCPm+TXQUeg7gqjfHJReQMvHaW9V0DsbQoea+
geVueAMy7FaxdgYO3zZalvELJVbXbdwAkFA34TZzgwzTpouWTRllESgcGp7C5frNgPhPZwPuoLhH
k3sqt763BzQIfh0q8oaByoGd4lTx/TdPRINKqbNmF3Vhh9Xxd1u+/oofUoVRJUkyXe8GqnJFb6zR
RA8iZo+731W1LNXl07IfgXNpnt+aZAFMkqYfPJSZ2TUzioukjSTazqVoSaOMRyayxgZt67vocG9O
k9GvINJuV8g+9nTIEqjZfLa+RMZR4BCqQlo0kuFXhD5Aghhh7ZSQP5QxqQc6fqbXXZi5cAVXao3q
sTg2XcwMGNvUxu54N2nwwr7qtnAMvjx+3f3rIqlYM+4KWlgbbAaPzi/Hz4hXDhmdsbTVaDBu5oOv
A6KVUlHjvvygf0KhQQXuO0lh6A1NlUjfzoAdqxHhQotPCL5uogCIlvUmdCb6clYUi24VL9VKIIna
CJgAjJmWXHr5Wy4P4358GRPg+1YlYzrBbV9q5VbDrYvjeQbx4QXZhvSHf9aEsaDgK/kpcIhmG6i1
HbK5AP79zX8hT2Z4yir4Kk4WxlbRH0yJ3nuSZd+cst22ST26PJBUf69B3Zud7gw1zCvk95vPi6c8
PxQvt5Zbv6UhLfhmoqTy2mS7p/yUTZ9wQteMUvW7+LmbauKnnTFnJtuLtlVM/UX0U7yLnjQSpge8
eMhw9XeX1kHE1pm8iBfprsEJtnW7bUlFQvmVL7y9RzeEfzzmadg1tGYIiVniMP3CCWGtD8VUKaNj
j5QZ8CwkxXAo/LonYAbN0qJhWBEy4LVWUJiwzYmVRpu0zoskI4pt3H7KMs4G4EW6GOG8cEqOqMu/
uq/oIgnDcb5sw8Hwz8nAEiG8SbPndRrJCktQt8ZdYVZOXlzV5W8D1uIp/pCV56lQZ3SvMAD7kUHr
e7PsNO+ngct08LPLk4GyD4v75cWgoRND61PomL18YfzjpZVvluj6lHnb2Zu4hhPymKbq8UvS0fTT
0/3/Xa9XJ1GWnPds6I+PzZzGSyeW9kB1dOUottTZQppSTxbW4WAqw7XoXvmjkcVPdP7nCeKLuLLb
QVq8xyhfccZ58HQvU0VKwbDbyphceEDJ+J3sMaeDpotShKvkGHYr9w8XeJ4H5xBcX5Us8PFPsexk
2XnNARWisM2KQsdAJUHkLxMClWdA9zXT0uDyRPbT998ZEqEM51Zx9zNZI03ZcRcViYxcJtrM5zm3
pPueAlCtxZRmcB29TAsxpLzwPJRZM+OnwFwb6/P9V717U/rrJdNnrEtWpncfJTyDKV+xa0yk/YHP
cC9mzwcsiR+hCfUr+sUJ+0POukfZ6Ij6a+2LNnINnV3nq4vB6IkRjl8hUVBjrgIRAGOmTj4KYbMS
litRy9L9edw7tzZ/sf/HixnsWcds2iyt9jEy+0PiXu8k9eT02r6gsho1Io/xvKex4XRD2PXc4J8W
m6JI9o4xE4rmS+V3FGvoygUo66xqktGVcDxtvTSAGoqZf2rpSfvWG6Egvsx3Sq/vWNfAedAlWnY6
fqEVpQXd7J9OUM+47VtL8n9uGfP2lh81aNmGd0Tv3OIqmo18h0LjaivaGVRnRhRZXD7fhvy8e/ge
uEQVIJW2KKMYoC0b84LE+ShY6nN7zuSYs0E+7/99rF5Tutw5nw9ZI8ZYZDmNOZmOtwGv03+2w9KU
g5SH4n/t19/0ZHB2T9GYv1xDjQcrOHeleDSxQpHeXgqtsIPpYerbU1AwgAW4vbK8XmAXVa55dFQX
3O+XHd4KsZgLL/9Gf0dR9UKXJ9P7auTkbSwgm85oFSzv5O/7wkXi1nMHliE21NMnfUzcExN0wKII
SXYv1HGT7m/hnD/IjX80ZNV8dJiED37M3xVVciq/tj5T9C2tSR4B0w8vZUigu4e1YmzJ01YZr01l
nVBXpZ7PPokffE3Af5M3eA03/OMw90giQHbjod4XwS5rNBWNMs5HNveXflG6uKD7uDWFgOjIAcgT
wc4IbpHn3BosYjv2fvSxot7YHrewvuIg82i7D9NiE8dpmlYlChMVDPaln+/VXi1EaSF9no6WSDAy
SkaE2FA+mDXpm5WATax+Fr3iRrpsiBe32DfVG9CtJ7K+Ce2hkDymS8uEzxwVG281AlVtRTLLQwpe
l0WmNqMMNP6aWN4N2YaQ0U3soz2e49wNe23qtTkDwta7g9G+CXHgJzTaPiqJl0z3WYCMlYCF0oHe
GlxQRtTkNHbPI6a5J24ga/R/YMYpkkCnemjt9+X8e4DABHXWEhwfemoX86Bc4+uZ2c5rIrI5uGIi
K46y6Jx2SCuuclFlOpOHfipLy6AEl6WIETIyhOPuNCTbekqeDDfYIQDOV7eL3e4PG4ePCAcpQIGm
tkXIGjW9BFc4icyPZpJxho9y2QuBhp8QhWn4s3wYpyvFftPDpScXvg9tg8LsCg3PeTfhrckCLKFu
CAvhB8heGYaLgmyzZ60c39RZr9bH8D0os1zdmTU8NNw4e3oL9wBTVaktU+qzgjPiv1z68cC5hPNK
g8C4OZk6Bl4SpTgU0SXezCBHvbU7RVk9qEEjxkgr+MW2CUq8sdx3WVORLAJ6AgEKfgoG7O3gNYUy
TP96qkkX0v14ii9ClzjI9rRdKnw41ulgfFMQvjRH1r6sVr6xwQihQRZ2YudZ6A7iqVak3ueQ0J1h
psnGXYia7ztf09cwUZxCNb3gk6mQ8AHLA79fCaJqYNJL3Ru/kvwHA5/TAlq6JQraTHk7sy2Ds0SG
pDNujrZxHksDNSNKqlXRtAviL8d/NzCIGhmwWbnQ+TbzelCjWn+xx8A2MJFJlKht7RVWF5eF6uQ+
eNwYGYWULp5RUyj5Vu0XDWIZfEE7Dk4gXwCJlSOeUiC7Dy8hcbVM61KxtEMG71P9tPQeq+TyEmMO
NnRjkS2K/4BGL02OWKhIMCXoguQLL44R1kQ795fC73RFFvYc/45ygdQSCAQxZjd4pQ3AXedX3bFK
qfe9NMOV8/UfJY+/Mc/HXY4Vvgoeyhg2O+zqEkhKf+AjL/961pgb+aRC03WRIAiqcRi/xaZQ5Sly
t6TEBmb9GUnw4kgjm6uqD9r78bwLhluBefzZLeMNbnnDTvG+09/+9GrGp2cGnx0tbhkGL2kWSIGq
9pGPqSFDR+H/wqS9wjCTf50yw/fMU3Bt5qSYxXJPOpc05/M7Xl4S3Y+ZLM2/Jg0+NbOrEAMrp8PG
wOUkku6yfHyS1u8YRjRLLmwUA1nlnlTfYcEK52z5TlASa62LPUc+IURdXspYzyrDoTl7FQj8zB91
q4wupliIIqCH0ZE+cXT6Y+xH+Ch0mCqHeTr3CGJ/x24juixG50ZlqcAL7m2jGBakd5R8FPBCf695
7LZtVVWPw1QLnl8AzR6LPIReEfpK3r5809xABVhkNjJsdL0gCSWxzMwdesOoOFmHifjyjce8Ka08
n8SbTWSNtxdksaVOzNOEQXd2G1SBKSHYfWr4M+3wl9momb7n8j4tC4XIZ8EtF+FvX+AFqTEiET0p
5yeMmWY9qdKPUXa7yXXYZIYnQwubXF/HJezXHL+opYWk1JXPO05QmSMXvrZ5OOGoRJRyD7Tf4SJc
+fWLzCc3AJqbBRdw35JRRgNbG9g/qHtEt+evig59Z3IeC7+wXX93kWenqUej/GVh8V7IW/mQiLlB
rJfpdJ6gq/v4BXbHWwTmTrTHXD+6vPtEO+S/BvUBTaV7/+eTtFwE6ISEQP7+/4oO7GzM4etVs6ub
rEf7WW9LZWTqmrCrIIZo7q2L0kM5n4uPL/4DwKGt6umkXVNnmQNVJw1nC/qrznHsxRQdD0J/WyVt
/AjW6w4MlE58Hax3t3o7wQn9HuFwQO3/pI/SLthynhQo/o1jHP55/7yfy4tkKRiN3EUj8nN0OtjG
ILP6GPlIzj+tCmhDAmzTKvrdJUkV9VSB9N36DKAy6lnngD8kYsj3WL5yIAnlO3jZQz91D2/g0itS
MYMwrdw16W6TLDB5vJVRupltdV9ka0gK8EfvhkLjrV4h2NdhvXPfoE+ygY/Zm2R3nEjOgoRY2ibi
AUtBKtxcR4/fdGWfm5DGhFa2xvt/auFvzbJLBHp2BXBdhUDVF2xIWZ3P8h7A0ZHCUaWXXrjLRGqx
5zMVhHk18eXQBXQ+H6RA8V2TtywQUXGwjUMAhN0TnyHx9ynSe3pAIZEIif9ga4y0r74T6bHA7trT
3utznFUKWuOwMuGsU6/zhQUgIsmGuoI/06J28uML4PJo156ABg5l7NqqJsoFRzhTgCWElJnvfxlg
Y4bYWr+Q/3pv63+NYyRU/E13wiTxNYzfDC1CA+yMjc1+7MjtOletDaUOvy4XLcM9NGpX3HyHwkQa
2CNXiaaGu/VHuNFpaDzijQWg90A8xoM8CEXZT2ydN/rzsYaYuxOkCdFVBniIPk/Ko8uShj8K4euA
nyzow5wkI11AP09uvTkndZ0QCt32Cnhy2z7UPDnZ2ZxWTOTeSWmd8ZwRfUlbLlNlLF+ymZwqu85N
Db9d4Cr3NwAxPXBjTPFm5x5p7lG07mqjt/zP3CRZ8ZMd35dLtjScQf7PokKD8eCIejZFqttASSdy
+8gQJatO39bKO8hGrO6lmkk1XauYPA2DbyL9ftHkmEi58ybqaanFjkJqXHujEaTwsVS0n6Scl61I
NGH4fFC7H6YhcFgmUQSD/AyuGr4Fe+rtOujWQ7/wt6fV2PJFacrJjfKlgRvcLA0Cm4XnygZGuN/0
FvrX7jE6Sj84Cdz/ouFFWLp5X+onXhs9Y8AC7/gNbEQISh2znE8c8GQKRMHbJu9x1ikEWQp3LH2X
sbj+W+AFlecyotHMmA/sKhVLuVFycCwqYucv+6+1FbLNFkHODcBLzuL8dMdybD4Ds5mrqzQtChKN
20y32VMJXaGafkRkSXZ3Q7B3oBueUR8PgCSmy1nEePNkUdF3X1clJvUzWi526Ag8OonXM8WGLLf1
sO5jbZqdi8qAh8zEzNYTu/mWzxctgpKg7qKcOBPp8Xvl6aXHrMWlZ6u2dsK31AtVjR/cSoWgP0zR
u7s2jlPZwTZFcF1o3eE/FDV0WUmez8B2to3yVIy8QwPu6Oapi0LhMmNagC4BM2WOtEgaXdaXf4yw
VbJK9jzOeOEr4MObPx9Lt14bYv0g7EmYaodvWhz7eV4Zj13ZZ9rodaZ7LYg9pI6Xap/LCNu55hTd
6qRF0cFNYDwn1Y/e+ws4DiczogrCzwHuCWOSUEhKCmkNsqcUf190URI8w4+YC0vM9Ug0X1IdjkKL
AM5HBCsmwVB+3F/cTb2siOT3b0WyoaH1/0UFGAtzmqA5UqtgvpMdnC78ZtgCh/ZN0cD3HbUxeWuZ
ji8kUSQ+mWf38wABvdhdTBd/Rt3tE8UKw2iHYxwlpRnyyq0gT7ObsAZsIt57oleOcTIxw6li/VDz
LMi7v5CpIeovzWHtPuurbPlYhuH9dj890RGIL7IePUHG+HgOSI/x8ZUgLUT1Cd4XEcWgEITlrLd2
ywZDBUUrsX6XyRaBeLMVIG7++QHOWjtqssBBCkK7Lz1AM6fMXUspU3qIMO0thu2fQLWqcMNa7sL6
ec4er6bHrqx+lhHALW9GZhUC1S6dGPQpvh7EFsBO3uE59UBr0wg+bWUTyKlNmON9Fg6SpimMfAju
AmXcXMdzy9idotk5VlHvIBHTjjObQCbvQJXnJq5E1F1wObPTY/gvsYrJZsh0iwfXLj9o8R6G9ynt
bW1cW7ZQK2eQ/Y+qwUu/gh4AN8NfQq4fHnzwLs5THv626+QbwEOM8UI5BL7d7LvNSbAwfSgArUT8
TK433Yf2CyrDysWlez4uoaZMtpPknNKFMqgDxbkQl7f7IL/4m5POBx7EhtyF1/uYHuOvsP7qEKZO
d7UN8efm4LEf2n5ceMkashIwy2EOpEl7m/oVo0NRYC+xdt4mAQMMJxGa7fCnKEXInKH3hmexVA5b
9T/bh08wXcNMpgQ2C8PJUKGfcEA48/flUpINxz8KFQxTclOzay1spth/1QIVHahn9FK8OU+7vD9I
VEXfM1MhkrUbU5IMXp+ExC0/E9SoAyuXWPvA/IIvGF295JX0j3NDAOsviJ8kSe54Zqy51g89WZBO
36mDm2GEPKRKW23QCp8s1hbdb9Vcbl5T/ciOIwNpZ5b0TggzeR0TMyKBafIyAaOFKhVwhGZYPGPc
Ly8W/wUagNCaEK90L7INHV2oyFYvQ5zVEsOgJZwYpzNqZtVlnIkasnb1ALgUD9HMktrAvXq1Saxb
fMU4TZampQXaOU/NbKAPuQuhclUJhwHc1W9f2UpkPJq7adJMxHJpvLYnzEpc/0JiMh3+a3ui/g0l
1xuOetYrdLass+Pd4HaTYESzPV5TyP+DtfajWr6ERiip09j2mH776CFTPZ7AUROxMYji/mgwnazT
MdwRmvN44U/bnJ5Ott5+6tDjknjNPuZ/i/cM5WdEuL0dXlFTenX3W4NetebIs626Um2ykMKoUFw2
yqQQpubdISNqrhLzXEICqO4FU3kuafIPzWkOZGDv9qmH0Un5gigOvYqvMJlPeQ2hlgaEM1b8ob+i
0a+R1QGkLY43Gg/Vna56HGb+EL2vWqH48wiylDZzZST0A1uYmEjJ39Kq8hxBndXTDWqHWS3h6LNj
w8AOKXSXJr+bh5QQrXbbqJes5YQ2tQTF+BN54VP5GJTf+71g02drYuJJbKb4z+745hZfVInB7DdA
/awJ9JOt8FvqQFXRmUotHXK30u7dZH3m/ERIL2xf8TrGfONv+h1+H8RO3sj9bsbubekqbVYp97Qt
tWf4DkjfsqMZEr+/MIhWnTmMK9BGfiqnJscAj6KO0fyPC8d/GFiRcuf+yUbFqMs9OpgjXIkpxzSz
pJbsLoMe/EG70LVp9K5WgSD9xoNrFWhzk87DdyQDiCaCvcDj0W7bfwT75+dXJrsGDm3F4IjyoCYm
SWykNKhPyqG+jaqthUT4FvgTpMsG587WW8yWVGjku90Xvj3XSwp9VSmZP9Yrar6gBvD1/FrT7ovz
rt5cRbeBqxw6iSqFYKdMFclFHHXNnQqX5uKbloPPLPr9KiuhHgdzFCBrfcsb5EMKHSGzSQQolm8x
1Rewes4WyvILxO88sR8zJ5o3sb2aACHSk23Ej8YRXLIJdM1SFdmQU3ASw5WQxq2qnQ3Jk2EFKgWw
68vcyanMz9w2APeZ4R/gPjpHBYSuEQ+rhh5p5nveZtEJix7DIsIWGtA95NtF6JLIx+nK4PsWFaX1
xi1huovgdnN3dxmKmwM8k0uf2UFJKjDKq3kKZt6jsdBbZDKsnO2EqE93c89eP80C+xr5ZK7g+imx
DprpAFpfCni1dCKjvmT+mYJRO7HbRol+GNEpmTbman1JWzaQdIewBMxcrljU7Foi3Os2wXdAH6+p
If5/ScJLTG8fyvIlN59OCzGX2DriVl2y4I4lwOKqClvT1G9Y9tJPXVgwnVHcAtPLn51opOxrNuv3
mxAPoLPqFbeuUSEb79UWNHD6L/jOYMijqQB9U8lAnNDWWnwi/0efLnwgoJOHWE6OZhBNZnODrgKQ
d889Gupweux7VrkUVu0gD9UzSzJc8H7fUyhw4O+vGJtRZqj6m3m4sLWrnIISrzm4zlQykZsKaoqS
O66Pjk6rN08dRyFF/Yc2cxvk58CEqL6yR0+SBGT6/6ZlA3RrdV6tH4Nll7kBr2R+myhnYzQbq/dk
XZB0rQ7hfFgbBKvMykcIAbnTtpeSCmp6oiPtofeHnz6FuWs6uBwOp2GzLyo6kzVN7NKAL/pBqLAC
9+CAaKUY4zZlM/AegiDYHaqNqQ6EgVzTcDozdqDHHcsloCRfmyT4GXgRDr4sEarxJuB8g+EYKxPl
aYtYA5E69B/zA4zYXdIhzyJsQh6m+y4JdNQW3TQaUVNcfpipltFzoiirtJhKCz7+Pd+lY3AOWA/Q
O56Y3Nzdb6lvEbEQa1ECpGUd+rsAqhQCnPC+rlJbUukDW3EY7JEIZh++kAnZbGe5VBUfQG6EhfKM
Fb7RuLrVrUPe/mhFjcBRrWfN+q90HLyc1PHPY6EpxG3MRROB5xmoAXzq3OgU265huns3D1O2ttPc
zAyC5jO2r+bbjRaREhF67V+p8hfbf3+uJBAj7cdlygxZ0kFQFAaoVbaGJEhrTdEg5lyb7TJcbjPo
Se/nav75cJPyOnqr76TjuKRlRGskrVh4DAL/IHT+BP/jsGuyK8Bs5Izyes5lyitCrr/qRIHLu4sx
mbEbgkB4VgpAY4JW3otQxlQSKESCXaTat250Spw5Nzzcq4xi3+hSWBgURIUi0La2mfsx4tv732Oh
bgaW1LkhIoryiGbdVzreSdJtVgCES3BMn9CVbTICEp61hF0Rb6njFnj+zrsvhrCmJNllk2nENyL8
HDUEBV3iFzWvEfD33xycCOLa0BRft6eWUYpUNYVYtpWlimc16RSC3kMHQwq+UU3KVgMqNgFx7MoA
Ze+0fQdCmjYdxKHk2SWYsTidE3Nl8kZccFF1Am6kOzgpdUQTAx1Ph4KhZQDcy/kK4n+banyM8gzI
sCpcoQF/VlgfWmO+qyrjslZbafswM88LVuJ5TDBMC02z21mN9UjDNdhciesaeTMQvQdjwiG42v3+
c+qUmRr9B1uTD4nUY1+P5xEET33M1XNIcXurKsmA9e+LJiUyb4Yy4glxGTchjorpostE/0ek05lT
XAKY81/NDCjWaQvoRhrtyT72Fka80peqMJgFcqMgolrmyuralGo0aEMs/kAh6J2+9JEqHTHaO5/r
FxZVkdvXL0EkJvEym2M0cdBSrzKDGfJbxJ1uHLkXczTEO9q9rCzZevBkgjV50qzsBvEox+lSixcc
RuoS/esp4FmA09lAjw7ZWhs1PvBRd6gpsVXcROsmqCMsUAYdARj4BLQoiI1axZvJsHtcY60GwhCB
X+QH1wfU2moUa/fPlwPoVOsH4+sBfE3laXdzYOypGOe5g+JmAYFH+wQR33oVz2bbdbtL5WIV7Ewg
H1aC6NK+yp0NYIzi5ERoh8oMr3MYRg/lohkhx11w7LVuoCuAP4oLNrj6vaIdwzNAAYFQCYftsX+d
Wubus8YGAqYukCvyE8f4uxd5sBFEhCgVpBjz/dlH35mytyMA+Hj4Df3gU2sI7YWKgfR7rOG0VImS
zCZrfp7mCMMy/22VxgfMWtkSd1FwkR/tuGiCKRtl4JerXCnL39971BlxHt1MVUyTPyUB4JyFtKPS
gkfj32WzbtKuBS32F1+r5RpQUNKNXgzeghenAHcTQaF+OHP7B94swRYK6kKUTB++KRaO/HPPy+Bg
4TESXW1JIY2w2LLDXmYM17KTTxdpCZR53ZHffybdgGBycOeVUhwvXP5VjLL4iB8Se3zAMZX+3GZD
ABwMxPUBn+KQhV/xtJsPNJdEhc4GGxGNiSGHMcn730FS9WJfhRG1d7sE810Vn5PFFRb33b2dijfS
sfpa0D9DCo1+l92JmvZnw9S4PlYii1VemyxpbHtMmLbuk4V0vvxK0GnqdzsRt/xRXlN6azlkShPC
AUX8m0JYD2uRGKMTTUFNaaccrgjSUum3Pvq3ZrnXQzGKhTK+zNrHLZhfeEVYI5GqyhOjsFwbvYHG
UfRnpEa0yRaJsFaXgE/cVPcf+BEs3pOCLX/KvS632WqKkCFpodftiluHTfcLOTL0umr42y0V7urJ
gpJHMUo6o7rUTpUOunDVemmiovZuJieX8RuFi/Sj8HDwpSc2m6IxhAtUKLrQkjD1KO7Rxh8Slulx
daBKX5AN6NeezGXpesqwqtPF7Bpvn0bt6u3T7KwDK793KugffIMs/OHG0zX9P7FiZWh735QMo7hh
PszfBkHBYIubH78nWHmpkp9Nk5wrHWF/yVINdHVGjJu+1kO6f2DkMzxlloz1VhKwsr/cpn+ApThI
1XMegW6X0oLxUvdSFntmhtKhWae9ubkDZF55MN+0SFwTfoK+65aB8bBmYFuOolmsjZJ2Fopga2Qr
qFVjv+6P0oeQ4icWWGMBiPZDjyqeBe6vmx7P/BqSBxTDms0EOF1b3dLY8uo3IFusT6pharDXJsp5
ovc6iRlgeWFm5lWAxVIpSjMSEYoEDdyQfAJtiGv/juAgvOky480qC8SsErtKltjOxUfmrPAncYiI
BlXCdcFps7/4TPHsJNcWy5Nw/MSVj4lFTrnqnlUiAR6grNQNx6N82lfRWsobY2qTSXJNnRE6BbwN
jH0TO5AixeK/c99iVEfbGtO8Li1c+SJRXBFTnaDygk36UbXX8nnryo+JvbV52ZPRSPF9RxWsOSz/
00/wUC9P/6DS5lVYwSL9VYk9RGPkJJ+R8jn2GX3ZCpOQtuHV+JVIUhzoFTzTCunnHf42X4zsoTZ5
Innniv9xJSmymKlAG+cYlpQJR19TSfZBmbUccr1y0+4musvOzBwI/4Jq7laRrYPHFJ0lctJVetzI
Km32ucymExwGvwl/jM+JIxqGviO0C+9fFQfoz6MGoiBWbTO3r2GUBTtaR2eLudHYzbsjZ+iB0aM8
8f8qEZ1h2OqUpqqyNHIZh8n4Vx7xDz4uOVoRZ4NFI/S9uHPE/X4EoPldmK86hisIPBywSPxivXzH
+v88E8Fvb4FgyiA32kz42CBGXB+U5+MTpAtwd1YIbDWLqkSEsgmGEP9JCLovdNc6KTr+SpkApPrj
t+usaWyL2CJHPtSlnXcLrP/068kHIyaLKqd1LhUcJf91bCJYTaUJ2pOsmFx1gHabHOX/PrDtsHtB
f7Bytg3UGha15q94ykIhzh0f0kXuoxg4nzvEtlPUGr3Ybdr5G/bbeav/yWpVTHsecozMVCKjdFCa
M01+94ic944UeUNxHRLfad1YlOhD2xdb1vq89atbXquprxFKGmMPRm+GKtuskmtl5KdPKKxyBbfP
Wat2kxTs+eMqJEVL+fK1XBWbtwTMgncctm0dW3xMGsR8XXhV3k+9XweVo55t0+/4F1svA7hDUYuQ
SlMMPj2KZyzhBXxWmXfdHTG8OERr32EfS7OL5j2WVrW3MhdV1N8+aBqBh+UxnBlXY+qNQwEUWlSv
Kddix3j6PeZwTuMsd0OX76LugaeFsd/IfYExz/xysffbLPHJCSRnLMIY34XIQ445hXkt4rLakrFI
awnDxTMVd+CAciDjzhttzBFIlZn68fbbdoI8zvj8TFoN1DAom3ln1RvQUa6+hCdm0Y+h7n0WsnOp
/FRM5ij9Qfk0H/+PIll6NSlncyMJPkUXiRK/s+ZMSwI1FAEWZ5IbR7LH9vOdmpRsgPEyIVwAJJds
Y5fEEq439bfOi3QZY0+uj6NdFKbSha9ap0fWLqVSwa8AnKyK9Fojiyw8t9RyiXKXqND2uRaq5s9e
qq1//BuCpZs8VfpmMS55FVgUPighC7qbq42BJwA5Mk1Vnszc5CzU9wUIFXGnST1uDJ+Bmp2bABQW
sH9XfKl1kFMZANhsFBfHfsntHEU8ckz1bj6frTE3TSnvExi031RTfcYNf45dwHcre79HFcCjpq2m
PPBFOULc/rfay+c3IjkJTB9orc+yfYx5/xyIR+oKMFruZ+pZ5DOxBbyeyzKLZhqyuvG+xLPLjdE0
xw9pS0vfKa3E76Gg4aJ5bX8bHU3eEzmGPS1ZegOq/G8TJito7IzGxVbRwNdXkuHTNSRgrTbAekm+
A/ipz/VKsrqTCmsMT7n9Q7HUsl8ey7XYk15KkLO30kPhiQk3aAhGM7IMtoxVGpQOlLaF3n02y8ws
sY10tfpHXZ3vY4P1uPrDzKl74kv6fgqeAVHQGS/oy6APOZ85Ijcg9IJY27cBeLNKJm2XTPY1kxCS
+VR++Fo1k70oBbkAMiOruxIyV5xh8D4mDjWwDqYJVdwctbvmRAYWkW7Z3SZnw3P6/F8k4tC/mMUx
Hz2hlusGtcFXSbA1tdlpXZNirwMa7Oz68ovzmx6DUmB4YUrRprQuWipquOXppkugee6w9QfyapTb
FYd3r1vx5nOwKgS8F2a2hDofw0sDYUotEYlKtQhwb3dpHRchM8DTS53FJ/EA276IP2AAqOwI3j92
WdLHXwDEbtib5jm2PJTOr0i4WKtFUDEgKoE0CUCQeXck6TENaYhFf9jKAq9AmF1SXpvHHRosyzYA
2Wh9LapX/ADEFZgy2zv5apaEfrvMoJvknR9xq9FTW3hZc1nV/hd/45JpglCGNrt+L5lkGQHbOKkC
w15kMGpfdcoNKekJE+IamKuGzDOFPCwNXS3tUnNuzGW43k7kfQlYTSXFY8bG9Dt40BwuU5CaBNJN
a6AADXBEYsHBD6tqQ+i4fn+cjR+bEpBfbCRNfFoIUx/CtpgUAZmxYoTekbynE7a5rwEDM04tNXTn
nrgP7oGbO6+R7kF5b5gafbStD1eii5bI8xojo9viNxtEXQnQwW/t8VCEwLai5nTvpB3XMSimKrgi
0Ml/iPWRdpsRmcxXYVCkPI+5c7d+Kj0njSz1F6JaHUiftqAjBEWVI+CBtqJ42A/iSNfzYc1TBfwe
0XJRRkhH560E50BKxQtWDiO+hSqJLe/veuXl1kLHOf3ZFkEjMNtiD2dFG1PN09WcoaYr5c/1+nJz
DzsXjIfJWt/nnII+AxEc8oqPF/37D7JhFEX19uQCoN4mEVm3rVoV1tPMScO1g9tG9FWRsVlFt1yt
hiEZdg9Jq6feHWQKn97VnnkTMMQMBqHug5xFTgiwCXxnnsIoVu65/e1acfQ6OhNvbLubicMft8Ru
8i6yZ5rtlOcX4SZHYmM3dooBumkNPeovMWtRNoB7BNK1yvrakRCVJB3BOVPjTcg+/iOuwkZpPUJY
/wVI9sIxkpPVvJ56dyDhJTQf3B6iQmJxPlh/fjhK2UCJy9icxhdSBifXgz6Db3tAiV12Z+KMPQuu
VTzDKB7GX9XDfyLiwwQe+jJk2iECDJGdH7ADz1EQju2IbXBlDgW8YO3FM6EERUlW3BT71VsbKs5E
B1HDZR7mXAtPb4ujIa8LcFv/fNzc7CCJxjq7Z3SqS1Oj71ZSZ/J6duZxHS0/a2IRaoF9dZiw2qas
2JtFwHUwOkt/j2SBbzlAMxPZWgtTLavNho4pQjmxMvUMcKTzkps87qiJmk649GwrSgqAdzkIBlpt
THaLX6roIDweLzYISkKb1I4lZlRyfZ5iSwJ2TIlQ36PnQoOZEpXgsu2z5LgE/zfMAxgEsgBEKTAh
czcGDff4o/3gHSls2KSv4HyZDTeMdJN2y654Kbtkcxf72J5cFmSyRt1mULoVdZAzLwrJbDu1M2TP
+hTiyutG1pyhH42p9RNbvuI7JkyRPvDl0mJhJpq80am4o4l9ismdJCFq9PmdFbPko98GRTcARfT4
KEE77njEesYbh4KkiPpiO9Uk6KQhpXcQ9bZ/Q4lxc6InKqzg5YRvDQt8XfGeatmDa7bOmTnOoJZi
KPTY3fIUoEO9TzE90lMIOsE370zHwV2PYoSHbdsmILE+rZJcWu8pZWZ2H0T3UDdrhoYg2prafdF8
VcWIbhrkV+2nFKqFnKwf8aj/rrIOpcppis/9haRyRTuTZRNeXMQaaSIUc3ONPEiH1cxmeoXWozWf
gfjay/qwnYZWqvO0IyuK5F/SQ0/c89qFWV/0ujkRkztDPzBXRx95lqjTp4oUyzT+C5oUaLgYNRE4
nR/6zlsSn7KcxxNQz6UbSos0b8Mx7GcZ+ijEr7TJNJuvsdx0rb1MCiwdfbZfkjUP+5jqSLQnkrBl
gkBgMyIEoLWdZ8sNextJF56DDtk/IJhlK8UTmSFvR8gt38suusyAnUYQo5xGPSB7jbSc7+8RHWbq
adYhpRXyJAeUGX3gpX0SmHF8A3QG95Zgy9VSbgA4gWxAzQV5/izVRxIKc36CNKlxybxJUbGo5Ydt
0JzL7aYs41GWZP58zDnWmS1jeYpWeMIef7Qf7E1mv2HOrzZxCQe/bJaal7DBMXottuuGnQcCPT3x
rG2QMkEx6s5roYotHpOKmVEdouFN4EDMWuan6QJZh7IZK5Ed3L8oLZvQTJMzMVABkHzoI7VwOF+N
z6zr6oNsfK5WsUNpnPqgZ1xqFFM43Nd8ybO4H7qvKA8L3+Ks4kZoovhEVh9VYTSTve1CcKgY9cii
B6isBvE+5JdkXrH2ZlCcaMrA8Etq487hjHBLcwtMNLoJIqNpcEgj5U0gnL0tGBGIV1zcWC36mq0v
YL1w2jpx5wOXyJj4UqW391MHpOVchjNKcwOdBQTOjctVgo5qALR+u9/T2krzehtf47xVd1LzA00h
e0lfWWs2qttV+VpGON9aeVLP7SMb+F2VDUAqhHATgZQyidfn0iv4GfkJt+oe71nLu0X27Pyfmt8r
Fv+BvC3T4sj6kUPjAJ/8uw7QS3vPfdcvHB83HXJLqj8j1Ll5gMdMdTYTos8upVRagwxL+lSFQ/0n
Iba6Dn9seVXGMnZCiQ2A9KZWA40fHaab2/gqmgjjysLODxAKRzoUlsFP8eKN4XtlUejUZNML/uY+
N+0zDC49Dz9Zu+fX4G7FVZnPTJjaywrs4F/Y90qvjTUMpWkfPfBvTlUubrd64KrSqh1GVjMis1Fk
IjsNXFZSA9IVBb/2cZ5QV0YnxDI1vwfG4lfIn3OwOMHFMCynO/YCqjxiDEhAajzU0wCdrfF1ONYa
mBFovyzYzRn6zOwfH10TzNgu6Zd2zyW7aFLzWyJAPb5kSyy4EQM9qCXJh9jZWSubm6qRaAy+/zAs
wm9saPKqrVSNRseIRe7P+Q39CfDCpMDnkwlyXHmGuO6rkT71d1MetUtEqvKjKj3eJMkG6ozGAy8L
3rF5J+Q8PhfY4wkNQoFaBAkrXKb3Oi9uESnRoegRPTUrcOrM9ChBTlohhXxi6pIFB+GwtQNkrVCU
i3KPUBAtvux3ITosj4ESmhnKFgHFwd+ARh60ERDjcocJDSJmhAHbfzvxwowST5Vj+iRVInlj0fwN
rzszuBrGmfblCMCPl22nJpQq4bOCoGFoAw9HSxAM7TDqDIpNwT0CZHLvU2aa5JiAjiDrRtUS28UP
0ChllrBgWCIEEPKW+aXI8qe+8NNzOh4WSrRha/JTbql5oUs/VWAwDvMspqYSZB/+p4DxDlTdyyPn
VMom3o6ZRHX95DTZD+C6TXYGNEPWVP0KtdjLzqRPcmSGzZvcMie6MrfaIPpHlmrrU+Qp1fcqsWgy
/GlAyPKGauASrHpcS8DYKiJYUE/vyC4h9M1jG+cDDSh7Hbcvr4ePKANpEb3C+cxakytFmBGC9A7j
VnWkCWI59q3quqcdoVaC1VIfoQuOY9RoQgIyZop3zovg+6xwniTnDeDpiuNaJkOp0uTgWZpSqjmA
EuzyHnJORdCyQkircibv2MAtnt71CcY0a3/ThSS890JmeL/+h4jesRzdP03PVYJErrg1aggU2lNu
xlgXNt04IuIqXeH/ogjlIz+5rjtWvLceolz0DurXfFB4HfYXJJiLRhUl3ZxYRn5a27I8Fjo1+ze3
ZvgVRDxk4iI2jPcGsz3+AC6Qt7VsffeTDnsGdIArGRgUBza3sZ7qnkxhnq+ZffeP//iTW/yXYRkF
fk1FSxhB6kRkqLtC+zoKlv8iqGmRoFHz7arlJx9sV/uSOWgFMdCS5Ovc/sIUloxwvYOOr3GWsc7K
0Y+ILRFpDTz0cwBj3zfS4BVhxs6oa11+K25tJ6z5g9gM9CxfQLnzgSPvuCzdhkqBpj+jkyqt7sXm
AaRTVg8qDyvol6F8iclpbQCDGTh3KxkxIAZD1m+APQZH28CYRXvtQBpyHx+CdgFP48MbdZZtTOFx
bPBIFYeeIEfC7jqgA86/5r9LyehUffHOFoLl27eRO1d6KExoKDco1+bCI2IvxVHjbgbATrMgktBm
wUj8w1qteoPd3JBu8RyM0LZ025k+MfKqHwvKuhZ0WpG/Y6prx8eWgs/v2MHskpMrSTyecGJSvMnA
m7B5tcsemfWa2YbIDe+mFkD+34uLsbkfiveRbAGLqLcPqufOFAxByt+j6MkfJZ/7vV8+WUGdkkGu
nrzyrwO3p7EZTZSs8XVSbkiyOxa3QiooERAvxBVAwXGZRUHvicQjKtzFVNg+3x6JM3Ix9mKtAW/2
y4ZBLwy9rLYDXuxKlyCJ84YysMWhJUB2n15/uwnG+ADqmMMbpRQEP4NGMjmL6gH932HhyPTdED+O
KkiZm0+gDCZZ+z4ZGak8P8T+cj86OPOdO5mk8TvDdNmebyjhxKapCG82/zzg8A1aeLQovlJee8Fj
0U1WFuHkYi2vi7d+dZI1vmsAhtg0ytXNeqPVVovefSaPcIXz1QjUuLpZ7f3+essMt1C2+1AM4y8Z
5Izwik865icRMLPt7A7/g08zmz3ncwLZTvqpJDyETHwpyjcEFz6mwBHS/XfflH1lmMksvSS6zyRl
S8nQHtYAhrptscWHWnGFOwjhCo45cjxkjfKqAOqTei7kPJQ7qG9ddk9BTS7nY1kMw9NbtVDIHbk+
FBU5iMTmFkpA6KA2YRt27Ngkp2lk7/I0hmDy2M5Nl09vhsRFxQyDhyiKWwodQq7fsyqgwyfUWjrg
D+vtoa9q7QMU7AQNB0N93CKI4nqRIsBwkyswUYfSrmm+vNrzmJRnbRSpg7xnFhsnMnTuCk0w3dFf
hdhzeLjXtrIRaJz9yNBhCehWqXJcvbxWXbumJ1okzOoOX7bK9k3RGIwL3JTwyrWG9TzReOIRdgny
ZNxGLHzVE1OP3SAaNLlEuR9Z0OA0rxeqTGDne7XWKc0Xem9jDlYz9dg3q45b+Yq8d3uCoDQCNG2E
lvvJhJPV3CevR6f0hLBF+JcqdtK/NqPgL7kBTxPZbLWigWCKjO3Ei4rwRdn7yyP+tb09pF2vDpvv
nIP8tGf3bSvDXxOpCqSvWlBs/f3138yFexN9y7i5oHC/bJvdC/NK1NYONBDNwd6jALwhWkWIqPu9
mhqERToO4hXZF2kbuIbU94/IW4IS8w66baY5vkh3Cr8svaVnQTxeT1PnZGi5gYnhGl/bh6VFY8l2
77Z23B4MEWSPEO04cRcGv2nLUJ0NKLRHdWSt/x3rSsggYaMWzlWN9b5006UWLSJG0QKDJg76YCYm
Cir0h401Igy3ZtStZHly3xg62I+RPG9zfFP9DmTEdLY0Ei/L+i0D0Lm8W+OgjgH02womuW6fa/uu
1uSZVAarOit0sI2sf90jDCdnOjwafdsgrIv6nce/MwE9r4qxAqN+aYtUWw5NiC2iInhUT7hdthjZ
5DR69kmbfe7hJkL8qxXb7YJ/5ro5EMVlXe9Ygea+6J2j28D6pS8aef8uGPtXwL6+Ep90Fe0rV2bB
Tv4EztFZgtKV3J7gmzJPgLZrjxNVoknpY0DLcrUHbfzxFykzq756Va+zlRzbXUufcS7T4Afpr45W
lDmINdn5nljTyElvxJPhdixjOZXu33lH9tPqnRVm51i8nUJoAQTz7shQloJXGQwPEdxJRU+GqJcP
9zplddPACynwkKviAkFNYyVjLaylaUCc5Oyemb9Pt6enGScaRswR1ZN7Cn5EjzKTzxvA/BVJCF+p
sKfkQkAAyXQH+rnQa7q8McanBC456zXigjccq/xVGX3cSDXgCusvyEQf5Yu0Dfvz3aBWrjE3qQG7
/T8hKLadW0I+ZMumjFHjg4tKLetYtBfRnNzIu+xpuvXuteCYzDWmzpMmlKAgp9Vc/9ENrnZcCV8a
svz0D5yOvAKKzV584l66hNf+SzEUyfNfxNzhA9gWNHnSJIWiCeE3TfwE3oJIqU+4+3pdqOeVQdZb
xybN7zIXpLXo6R31xhX1HSm2pgrsZfb/tVR435Qz2ugFpZs9R/stq7diQuXzE3ecq3VDPxuBOTs6
jJzntNYP0FBWJvaAg6EQfhINX3gCPa3R8CjTBkLijfSPN30S5Us4UyLD9+2nVYLYzNyXoWYH1BF5
wPMBtLxfHaV7HwFTPBH//r9bTnsrc8rsTwFbHRB+oJxP9yM3XSDLYychQuEsoqMEmDBHUtIRTXqy
8l039FojYh4bddR2If8pAZiNWZ7ekkRfLT1g1UJREoGvFcPxdyF1KvSWOMTMMI2mT9NZfbOq1Ygp
NvEyl0JLAAC/SdH+JqW73KgGDcV9g75Auvimbnv1WgYyA3d/CiTO0Q40YKJuD57E4WMgOdTDGKwF
VoAnUv0C1G2uQ1bjV2LEq/d1vUjVAOSxvEorn56M1fCxAJhZliVwYytrAAU8qRGX6P9xHr3z+X6m
kIcnJqAuv4RlECgl9tvBpzfEajbHWb3oOArFpV4G6DavTGrx8x+BxRGlOjhQAJ5jZQN4SQLJsLy3
XFfuBIQ3LMCVaEBvOn4uTRXZ1QHCNRrTTxaKukQd2IQQ5KLtUngUmWBKw6shDakpO9yZyZWDm/if
4DIJH4tERFbqX3w71L1Hic1NgB2FrfjJFEq+9QpX6Emo+jQwiQmpelrF+25xDK0ut2PcxcMjPGEe
cdb8Kv+MGx9oaytNk+KCZe6NST/3CpyNDjrVtWt4lho6PwU6uH08tBL4c6rLWLwj10vidY545EKy
ZjGq/xSfh56p5j6usa64/a0PYoimBkmMkC8ozxJ5GMvvHOGeH4CMW8st0sliELEI+bQBQB7vX0Df
WIkPbxKvjA/xxARv//FWMV5I1cHMMwLuuFwOlkeUUZzi65XqcVWRxq26J0Yt0iJDTKnqr5hALXZJ
ZLoVRwtO7l6Lg/kXyqElKSAHsVMfgtcFFrmJTmpvXl+wNySq1m/Ip/d1ycv00F5nfOooUbtUZ2KX
1bYX2U7d9//jnhRJttHoKUaSk7YFUP37e9e73rM2eM6b8cBHCijTsY+kavHDNgRcAmvQFrQzmYZV
PJK1gHgXzLK7z4G0gXYR30xCdmcOfQYJxdAcyZU6o4UcAbWKXubuBwr54vjcDv+6XReXbfEpv8cd
VXQkzybGt7Wy02Lck9LK3uv8ViW5k+DVNyxKbxRYntwyxzskVnREconG3G0+gKAUtqZFSdXq6AA8
S1J1JUvE0GIZai258w1jScKQyHP0+s5vdU2DVJs7J9Yao7WGtCAI9qJWcUJpAFAot9jtKjDp2CJx
eE25wNb5x2pCTI4ZZ0rJiB6AAihPEsHVZleP1Jx6asBpkop8wpG0lVK/fuertxAErO+NqqY6X+8a
0ylUW2oaRfDKCnYvyCPOfBqk0amFZbGa2LsDQJPQUsCxK1ip15YrrqzGXu1tre9ujHh85X8ou/LI
nSXCJbsiD86flxpUpGnVkkP9KVaVBNIjDbc7/4naX0FRlI0kLDibNM6DdG9hryFE9kZ9+hGgSi3B
XX//3Ejkyt+yStU2u4E8hsOHnM+L32gmUCB8TvmjgNAh8pCK6EEImb+41tqDwqyv8MZGZ3YWAi8w
M0CMV0GZqt4/h44uVQiaJlLBXsr+FlZg417v38Yh/6lgdYDrzX8+5d8P8GETRRthlOFd9OO0LEe3
DUu5qSYq9nxUlmBe0jo+0iOZJjkiTf2H0of006+atHGnFOrpLh1yIaDKs3ojLHgrrBUpHXZPRu+r
Yr20aXcGoS21ialvTu/wwJILJLKnFSAd3JeeaeFFAykJRSsfuCXbAMZssxe15oF7U3OqVIc6Zv0a
qpUzkA89VoFjlInoSVzQBOWB1Cp1iFW3E/2fifrwV0jsq3jEHXTwl79n2b14NE3HK4/3uAB1OV5l
VynTqoC4O3QgbfyvHjthFVbtc+4oX4FL5Wb/WnUvQzB4Ibj5G+Yv/0zU3XFiXJjoVOQqQcExJafd
jvg1Eo5vT5QLPsvSlq8nDDfguEiln/nlZMdqZ1tHYovcd+dDW2mCbk7FJSO1Icm8Fn1LFJ2CRtSR
+ty//doVJWjhyqRXH96XjG7Ykc3CIx4x2TImWV3w+ONOJhGjvyDlpWKBXX7yfPFXaAZ0qdXv4kRX
SmB9SnC3zLN0kqr744XYC8bRovwVnR6D+gh11WveGBs9aDukHcArum5mo791qGdXP7mxN/8/brZS
7CdN3So1j4aA8NniYp2FIc4ucfAMa+5bVcTXS0SBdG4BW+RB9RIjQL1Mz/RtKfc2B8LyZ7MfRKi6
vcZA0jao5EdJKDxBWyg5Aaz3xv6nwLsMoYfDqgR+OJsmrx6cUurdI5EGs35vb26dZFX1pKb0+DPh
nW9gL0B+o0aMZOgCie/bNGcdSJQURqg3W3hC/rXRyGVIwGTi9b/uLm1LQBcj6eyh4qt9XLdUerd6
fpWkHT1shhX1bP9k67ZhEqACKEk6Unn9YCcGa89PiltxBWzWYgh3YLniojWUCMqHmt3ltVVopMxo
uFhL+Qf6lA7f8hfOV1b0eQYGgRLN62rIDsuDMOtrColSk0pn+PuUk+L76pwmfkAI6Qy1x7Q6zaQK
KZ/0XT+Ju34DaN/WP8vCPdmyaZHGBnNjX/eHiLrF2/eSuI57XCF5rcsyvCIUpE7iU1AVV4BE2Jp/
05b3s81fNF5ilP9GzUhU+hoWYD4RnkrEeC1b36lUczGsNGNyqT1bJ88j2Kd9iM5L9SqPF2drb5wq
wpOijG2vgYxigZMmac1scYs5fl6GBmM6ynJE2yKFnQV5ZmbXvp9O1ZH5kO/iKPOi9VtEYRgRfSmD
UKjumZ7lHOpaIvBjocNQWmqpIje1asNDbgq4kFGVM6SZ6v7wxt9mILjF+k/4TxegQh4fLncf+hY3
nBjDa6o/XwJX23gCFM5Eu/i1UQSF0T5ET74/gAarHj+sjixXMKQIwBJLtD5Earw7O39YDfuICdBM
/dZmmnTcHxpDgcVQcaMw2RYHeSLalALlm2j7/WQVEX47vM3jzluBtXmchW2cDILfzMSGQhPbyRij
bwyqGkHL6Q+kIUpKreMw0LjSaN98n28Dk1iUN+8uwogmnYoPS3hF8a0P6aDBnw06aOrsJmWFfJtd
Mobu3CDj8yvOiE4AG+mcVVH16Ja0zRx76uRGD6gMFcK3e7K65gzTqcsLnrzjLA4xGVK0hJ3g9uPE
VNN/7PnIP7PY/CBJ2p0iZVUDaZFmPgEldWBbOB9+B6/NkeszLZ+A/IHoO1hk8UcvqmjycY8FvqwB
ctmVFsqXnA1tCGduTa0DoVJf2I+0PAkKIiVkrYZhudZNtJuOKB39xgTehSuLDdzcUXxM5TnnEZwS
nHZgzMu8Y1Ydfqg+KDzGa0eBgnnAlwqgUM9aux+qUnro9bexXKMCh9jT7Zt6c/F1NGovz6Eq8IWW
6bKv9MolXS+n/nqwEcc7cJ5aBd9NOO7yfEU4DovV7HsOxMwADanKfq4bQhOPaa4UMA3e84T82gmK
Sx+RKgb6h85bOEM4Px31/U49gnoawA2fOV+LHLxvl4fIkYBGFhfo6FVX5SnOL3kz7lITeDb3UM6o
WGdHYbYpFZ4HpHrkg+GMX+/BeI5wRCqmHda/5sB6fSQkcGiEHDgn81c7dX7UmgKuDyptCMRJLpoN
YZyMpcYKApQznC8bsStHFQMf/f3EkG1Djus20QEYR1Qfc/3L3UHwfzix0py9kCXkTF2jpyUSAfsL
YNL/zBm7HNshEOsEJ+nEPf+kcKkcda8rVf+Xgw5KVNBrwFFLmRZ2mC5f/ltsTgjBC9pgLjpHm/js
bmCjmCECk8WlXiioNuCCJhrN3nRZoAocp1noozk9TJYRiBuEza9gQ46wjl8nNN+VxeVhg78nXqcr
E+rAYeBaCwnZIqhWrWnH2vkOXKJlNIGjfFQlge6a0rmZoI2iIcBzybq8IyYpDbM7Yuu7TGyjLyN4
l3btXeScB6gyWCbImagKu9+Upl2UEF1y1SaEvVr1EC9M9M0Og+hlHeT9yPY6eT85KLl2/8UMWYrH
bTBbOMQMecAkc8mMcWzu6fnGB036rnIJaeTR5fsFfnBk4Tm54h+icw4XCC7xwCSAocLliTsu7WRq
5BeIWZruIaVuyjVFaw/UFJ7kVfInutALWjrVak3raiztgpbksClHOFTR0smEnnkFETxZvTHSY8mF
w2ObtTDBBBqVynO5U35ZST5psrJsDUXtkseYr+iKxWJWds3njV6d2iU0zaiFwePKaoFQmtz9DTgY
jaB+edRCcE+PhMVw/K7znkNFUdExVawkzOULnE1tV9HcYJr7qfL+2+8RCB3mLdpge76c0eIvn70+
vm7FhUvc9dHtchshRC2lWXCg45CaxG3OaGE0t3lraSPk7V7TgqEW0c2FSj4UHizfXODsMIYgSDWj
kMmzrUxpDbawTKqJUa6l7kKtpJAnLriMl4pWxlNqzrtVZrSINPN/ZP4QxnbrwU7+oF90q8RfV7oJ
YYLdxX2hS3saoH4z6fuy7ifIii8GR9CwekVjOAcuqee+q6Fbpmv/Ssi+3PrJpC6hZK5iPn8O/w67
UhLcbeuRbhR20+T5/9boMKZ+CK1WYeZdODqmsUbpF5SYCt4FKdewQ2kRpnp1GAtMsYYcMu7WYq1p
AKr+6uDrvxYm4AtQBVFuh7U6mhU54gSJ1s5jnZ8/zyU7/Ueqtb9+UyAHUjhJYTh/TdWP1Di8M2L3
UuNTFkK7Ri6UzD2ZMTi++FPhCXhc0OYkPAi/waoXH5TMtcPzLyJvNxVow9wqvoW9XKfo9jo60rco
Bm6FqUYAWuCVYAYVbfvIwWr5SnGGHz5QyoHYF3c5/ESfRAuf3VZOW4e3AYihRUFMOxeQcMNnD1sz
IifHe2n8dsvwojMKouHIK5h/gwLFRmfPRa/zwQT42G/eUU0DXP+oT7bzojTs11xNb21kvO5O2cG1
WwgegTfMx5ydTrl4Ch2WpkqMJ7Y9p1hhmeFG++SIwUR7xTs8tNUC0wUUFD1Ta38Qf5fgehNWx0fu
bcJW5Yqhb4r7TDXyIoRRLp57h4wsQX+rw0amN/NJEa3VND2XPutyNYUOrd6RaDDiOvSWQyhVagQI
UTk2s76K5yHYiGM6b88OJMIcxDN1ds6OSgguPiBsC5nLyLPL+j3tdlJWOqRG5K23375Ce2KC5Xdl
G5hi0C1MxKjwbd65BkjcSuq2za26OGnqlHylUPSO4fdj9nWRY5WkbVRkx9ePhtbEsG9buPHxf8Mr
vtLzxhTbjrIdi1AK2rXNxa+9BUNq0IwM6dZlkx0+PfsYT2ZkDQNq7uyRCjrpg3Yx6MnpgQHpUlBj
mQSJEkK0FnAEuMoPoXBTojZvRa24tHlmnjfRScmWRpy9fXTCr1qLNPkLQDX0hoXUSZAO5MdI7aQ/
IMcXq/ZINatlCOkzY4siIafsf9pmvcsKVDnF6V6GOxPuUcYHO/zkGoATsIt7keblMBx66CveGp25
P6sPYuVDt5Aje6HN+MbjgRggAQT8kZhGRK7+5ljJHBRznuugzOtUeu4hpdx/FLHAEhlxsz5mM6M1
tvClVeU0tCzRPACQzvnY4JQqtPM7uLZMQWx7RVSiKJZ8xuaX6f4GpzMXvsTPMWpTa8kL/A/lQWv5
YQ6+5jqGl1SFsJl5dy5N5omkTjzbuVBsGIqVsJdjzmxJaimPpwsO+swZVqMzkt5zG6bZiDtX+678
ZdoF3t3IaWDvUUNHEcI7BuLmMHwevmfdYu11yLuy6K8ZYcFwWPHVQSEgXg68vzwhJGyiyL0wSPvg
yUc3Hue/uY/b2NpFbVQ3YAvp/pnqLFEZsWu5FUP5T450oKB417tZNOMEGF6U9P61kFOTGTHPoGJK
stgUcfYl7Dh9zGbKR+5RkkcwBaF0OkqQNWVi65lOxhTdUB4H/4DLRh+spj+PPlGsq5+7OZGbVARn
yW/dX846CFy3OvTzfMegmdtqWSU43sF/hPK57VEhNUPJYGSS3TObMxqI84JtpxvFBZNRpOM/BF9G
UGgPy/+Dwrr4To6xhV3UnlKfptUPWSz1Kyb5ZAhiEZG2VJfP1vD6aD2Jq6Ol/5rm3Fnvig3F/un2
IXdURpAAyXo+wTRuWjcjzWv7n5s8ZWJWZJBQNjxmVDvsMxKlfpzhW0nvCw6XIslXT+a0jCc6xprm
BZN8yb3u2qPQxCA+Q2OdYq1LQlAQQIBP1kXA8u3wFOt+r8dd/4LJ74n/rKOaZvcEXJ98kg+hLdS2
7iWiGR+M049uIKIoHpT1N7byiZ18pVNEsac3RBZdG7HQVGumr/jlhH/COTfBatDs4SvZlJzEIxWz
CxvjKdY6+Y6P5kyCxRbVAXBIOGQs/2Y1hIEMpZJCn3/3iGHsM9mJBlhq82v2Wscasd6rQoiF7BHD
7g2/ZMZ17F1TVsD0RGxX28OnFVcMRva8H3wMri8YJ3Jm+X6Wl8CzdILshE/mAkIpJKnSNyl8Y2z9
FXJap1YSzjkbQEsmmvD341ToepdU6B+z8AdlFpn9MLuy9eyHPILNZCZeF+joBa+Mrj/HBnWVR/5o
Dgw4Gisim8QC9qEPNDF9g8OzUZKzj+r6id2nLzSlhsS8ZHGpzHslD5uCawoJZ1qp6TOsPUjlM2Tl
z7H3qyTx/wSl6KXHlWDnBAvOjy2uk9kdGyd9SswUYDAVZwNuthEkavJ7eEfzvRAwvK1dRH32EOkf
XK9wNKBhi6WSD03wRmXo4vZCPNGBbhToRFSWRedDjO/8oy7pQT4Gwtmdd9lDvfDMh5cyS3+nFYOo
mqxbDvTE+QPFW9gE5oQv0khR2Tos/GQgJh0tdqRemytRdBTFQSziqIFRb9p/xQRtmSWi2iTTWXiP
rl2aEU7Ejvk/+Pt4DLCJzaZ2pDLTGRTz9ppvmHL4PfefL5AblI5BhSdxShh5QKbkuZ2KxidPFxsB
S023hOymWDKbvAaB1jMn9JqLLJIRybSMMLMtOfqxYRxzAztYy1r/JhwSIniZcET0Zr2QAEgPteph
1oqYRJQ1jpTI2CS9Bb6+7nPX83/t0nQHf2DHFB6IEsOyBeYhjHbRDS7xDyTL6aJpW35AgEEBpp2r
u2JYP0UBON/g7WsanR1AS2Fhb2U3FDWNJpQAj+RbZuD66U1k8wqbWnfwMS8UvRmuLOInK8HYiqWR
1KJAY7+y+7EuKuxbkm3gPW3T/1UDu3RtDtBw7vSI2LqyYmzpJ/uEfjmYvmR14dWPFLhI8CQtcnYx
TCy/Fo70ICJMVXf1rdl+u0XQcdGMtuFEbvqsFuRsn5nvHgfFg5R2ZULF+db3Tg9nw75mNyzqgEQJ
DNrw17ERT3iOY8Wg5VwxfMpgB9atc4pmtxf+rBNlIDLC1uJvvvsjxmibJh8K19T7fERx/4tuWDFO
22yDtgS3YC+M2RA38msD7YHOBmVlBfHFPttgr2PzS4QqvDqEWxgrEOw1FkpA3Gy+Ix4sRU8s3ZjT
1K1xRWGJsj8on9ACCvjfriPavpW21p+BEjW8er3MKg6C3wCAMmk5OAJaYbIX919wIo/cSwtzMR1M
7OcrO6FJgUCYJ9xtyLFwr3ecKuPUYRZemgScDIpUSGJKy9UaIdrui3MaBr6TrEpNgZ2T7mCXDzYa
URHD9CIxvWRjsjN4p/aCRuy8A3xAIQfjqh8idYw9/o6xCUPTysZjmwxW7miTfL48eLwwgfxNox6w
PB0nvUVBBB17b9p0lePobMZA8SPiJh1QJ5t2pDktVKlXDK57glCWswgX94FJ31QEgIgI+vvGMAOX
0PPk4ybiptHKTJwudHpf/2DDwK/CRx1Y7YJnj2uYPJSP9VgHZqfIUvYPWSPnEWvpkGqjaU3rfeWl
ElkK1YUpLKyPmyYCZwqFBs8dl/+CghcL/GnLV6MDCaXvu1wEn/9ejaCg5/jaKESESRro6kkkAf+k
v6m6NeAuzQZ9xNSKedoVvTh69kNKxoSa8HaqEy0Qeem9G2S7AfhWUxHv6MdVqmfRhmjHv3j+k3bX
Qhypryh7yqnONJMNmjp+KgQzTr8zdqyyzSFi9T8XuZTPbGJM3/QZDSjyPvWRV2r+HTScaVWHbIoh
rvr6wY71OZHngI5nR15IpqXHCcLG/QZKeWYpMDKuou2EbGyCSkPhVBENrZi0YUa8JwQGTye0D+wB
Z5p18tV2cg94A17xH03slzZjAg0kOaanxVkk9wMLxAoq7GbE9RdFJKb8qA/gqolpgxe3jP0jhDOJ
SwTCIRRfN9L50geVV06Mo0bHF05qChCXetXJjQplToWTKX7opOm8xkxRLVpEwWkmNYg5z7tlnu0W
zsmgxdaQT1rAkPH/Eqvoa6uoU3o420NX19dYo79a5Le12N4fT3+sInm8E1sWPw81Ijrfar32bCMI
C8jAOTLH7ZbVk5kC9mAtgFActtJsAuohyexJrMjoAlKRPs8an34RLtP7A5qvpqABzwe1+yxnYhU8
Qhy0FMBj6xawEfk9/n8+PuJcyI5ye93pOUOuK0/3OY9Gg2B+4a8ujeuMxfCk2H0rI79tXSSb7vcp
iRukdzhgSw30xBJ9KdgbAtDugRZ2qsbsrlHW+hbjgK3/vdIRyGrj4UwwolVL/C8lbDqB5VuTKvzP
QejqDAt3Yl+a8lNqT9AcEskH9IYOtHiQmdVcnRY4jDQR0r4ecL50qfrxp6QTAIi+MTn2k+WSaEKY
dFCXRcpAnzsL4frpyJruWoNVavwDRyw8YgBQN84HjhIFZpH2p/nTx3vpTBbqPaqFtdCMpRpqthdP
MSZFol8kjK+k9Qd61UywJsPolXd8vokwj/UvQBKCwLEdPCqkvMCV2gw8sAsZeicLmtGPszGcOZR1
1Z+V+unZJU1cJpPvgGpczrssw9tRcQwbxPn6ar9hGvaVK2a4/ciVrlNT9r9GaWBHmJvjUyEJcFz8
3RClnDx7G3mRfbG3H00cZYIxobWMi4884kgCjFcFN81iXtLWbHRUpissfPKY88st7qCtilLgyqBl
itRi9/fPElTh+YZSEGi61NIsHPMf+bcFFWBkD4Z/XXIRJbE8oLgS+EUwe0dMO79qnjCnGpv2o9mc
8MseM6SvZyVpSfFZ44o8RZjT4rHvfLfrRR7tI2ezIncQBMgdcnNtQQCS5kJDT4nBec1K1i+0F68E
6KB2sxUCXkRXQ/PDICBp8hi+V1lhoMk58O+aWohaQXKOjtbXN5VTsoYDq2GOrrSnGBxwIh5yiC3u
CTHrJINdeLlbf9bXsKfkOVGSUDTSCx5nANbaUg/DG451tiBz9dcp9H7W98mP+A2iM++P5D6HT+iD
YK69ckypb2UDqGHnElrk9d1Na3bIu8evAwgmuR/E/MvFf8VmyGNtwIhJxQGDfM51qxcOvijR9AVp
KytibBmcVBIsjpz4j22s1Z6pssbOCXUjHjDtpp52aL4hbl0e5yXs9Cs/3lbSV+h34bu2VY3aDLE9
UZZgXpXkTW//ducxRiGeXEevlm1AgsRCjcbH6gkM0D+zj4Z5DA4Ian4dVRoAVbLpMI8ZTTX8ywFi
rd5Xlwic/yo0HGQli+Tp/ANgU+wMA5inCNklDkOdZP7F4FN0xHkViFKvZrlEJn8VgfqMT9YX738/
ia4eewDSNaQSCFLF52d3JXHspDMmMb9KXLEL/d59gBh7+K3AHiXiqQMGZx+63YPTuELeJe3MSv1E
vlVHMyrqs8cqeYaIgwLI985ocFTrgwPQCUtPpxoi8HtR9Uc6txyGglyTaMe2HHTaGQmN3l4vCpoa
dNrcnMSa2DyiE24Dl/iyWu9U0wpGhOBMJXWx+suA/gBW/coyHRgHfpmxnQ33eH6qnqGcbUdr5/jj
6i7I0R0obKr3sIYgyjX9MO5xFXUqG72EClfpe/vAF9tY+rOabXrCxLMn60A8B2c9IGvQq068pa7z
lqCbZUCkGhw6IbcIjn4ki+thamTaGHGeNHebSBqGTeAH+zubVcbehlzNiKd7d0PauzrCm5k0tz5r
FJwMtKDX8TAPVMguf32E7n7C57XtPCkcaxoPLtzcq4ruwR0bt7TEVaXxkjdLtyE/edmvp+kD+Vtd
QYyJ/2VBWaL09GBzvFSXl5WqPIjKxz3xjVCTbM1q2frHF0NEqDZduqShHUSc+rYYcd3PTOG4e6as
wWXdrhv12zy/nZKCh+/WJgyJp0dDGc8W9ZxPC4Ab6rNGFE4g2EKeAuM1eEnNh7jk2eo/cWcqEjpr
UKTsXeXo539Mj8n36dFQe6QI5eMw8J2veMnnGAq30Iqi05klfN9ppRAiWqhr29PWY575ZWPTfuLk
ImxV1Mga+WmCtHfHbsqISYqEaNWrDzOJXj3yfwxr6d4YikR7y02tJuCNUeI9YS3yd5jd/VV/g4B3
ZNBXmqS9Qs3dnBSKvCM8lKVsKIw/6sCf31vEXZmcBVcyeWlito5pbEfFTcqgIqCOzgVONtu9UkX1
Zlyz05VfEBn4qPW+d82jO8sVE3UIOZErX0jFWh/06RECuk1duFHcdyDV1vyZFPpwFJd65Qybu+Do
wy7lTteKuauUjIjatMxIQz8lhWi89RzeFZnM5WOq+HSPX/0NY6I+tiG6kxnghCe5FURdHstjmT2F
EOI5reTbR6HfR4skIM1IbgjomnOEdJ7LCxdIiHM7y4/QP3LEGyd48ZoijEtS5qfy8NFfzFE7fqdX
/9V7eN7TQmIy4elBrCSUL1IrKoPMCe0a/cQ+s5u4j4lGLeKZYmXU7kHmxdCYjpCLtpDkBeWpCaIO
yGQE2BweQwl1g7HlzPHGSflthisvFUuJaGDnynOrQEB+N6D3/uTxhRvDppyHKRuLnvKk9iIhspgn
EXb92/FWxMBtkJ/inuBtwiMq0LjRGMnOpTJmOOJ/4tl3KQSpNq7RlvTv8COmHMjSlH2b8XGqiPQX
AT0H2umdXWovh94+lrQidVnv33hiN9uuAF73pvXxqbJcgXOqgXALafxAw4/vKZv4YGKaKrT6Xhkx
EA8nkpFRgzT8d7WXeo/3fI3eoSPCBaVwIKhGn7fSRBXXItvkR78SrUX5jWz7BvSGEQOtRC3SsSOD
+6JQ2otJlg/g30U55ATR2q/Llv1EDxJ2pBLpV1J7OVa7mX/ovwvBffwwh1a+JfRxPhhRdl3JsnZr
KCAxmrlxXnppJ6YhvKqS129SXN/ac4VYcaFIyK1SYhEnlneMm6v2N0VDevFwFIze0XO7TSGoG6mN
tT2iy+Kbzpn22FAXdVHjJFPWybx8XCksyLYAjsTvoReM3rVL7qj2tD+ACDx2hPVWf7YiZ1n/iRhz
Hajym141ezxTcjTX1yhRKeJEB2eNJoo6nQMYtawnuhoRVMCY7oYAHuFf80k+NPA8LTt6uIH0VSmy
1uOO1vAfS2MywBRhWGRiR1gagY45bHxuUmAuJbR/HM0P7DPWFk9786CviBrQrlxTJ3GXSRcTRTs3
BDvy2T02wLuyUyou5a8Rs4nK616lPHa2skzQOrYRdSFeqKYraymy8HjXINgoAbl9fASuzJK83GO4
KfU2a/AW9MW4GDWtdIg/wULuBa3URPSZSAzq5e3HynNs9wMeENUSo/ISNS8uI+g3CDYLqhMkRexL
zE5uAYBceU7U4ySpYug2pd7BCcwgJ7faJv+8q8fJMdbGARXzmekUPz5J60SNU51+1No3oZnD6Jme
7cl+UeEWDrmwqYpzOnldak1yRBiz9q0BT9ajpDdp4eAvqNdCyBr2qN9Ng0zcNXzZ6nGFMt0WAB5n
LG2Bccj9TBbZTQE/+Q0o3TtOJsZMck15Di47Fd4StiI+VB0LIReAw3OXuOmCtEyuGpTp7YSGQ9uf
lj8PTq6uBx1nHG1rs4eoCAmeYUWDIhigCW+QfFvIhXaWie/D0dt8PhtxvdKBAMDrM7yTPbWOwIlG
H0sx28H4iR38W6jtcyD2tdZOXZDBJrryKIOrgjCcBgtoSTmKK5HM8DLxylnSLG94Hm14FcmLkLwF
yC6ePPFPBNn1yKKqLtKPgyE1zUHMBYxKBNMvk/HvfE9c0NHw/Q1fhlvbmS3GOkzrdz37SPT244D2
41G2YU2hCepWUv0Ygjue/lneWWwJRhzu94I5D6uXrJBldbi97zdrGfDBXEByAjJT82+K3smuzbhG
ZDaPizgEM8wPygf01tA2uLaVwiyTvMyw+nvwtJeGXXyI30HqcQBsTYY/jOiii/+7VG5WyKZPUmOj
R/oc2hbEh2pGonXu8C+yFna0+lmenpG7KqFm4VrVtGFyLJ35cbfAJsg/MaSFdYAUw5bsIE6zRwx+
jbb3FFdS6GJIF9Gq5HlI0TUtpy+uX0HrJnFeRXtVkJrCPEHr1Vt4txcgPg195dGCb36R5gp5hf2j
9SSqMzSYz+RKD2ablAzPr7mhpZsRXVYNs6bGg+i36W8K2SgpQpB+0AFPEtm2grglZCWho2nbaqzW
Bf3mJeJxWDgbTF4MJzl3omQuRC23psGOOCbgnPcPeW6NrcODrGdBj+Yz5T/pPGiklj2uLT4xl92g
NfyAgkFLJiVdlKS6DO8pi8dt0DE6X+ZEY462pdfTWtMpVh6sH7MdOzc3HixnYcCU/mokGA7OS0lx
elwUCQ0WSIxWHJyH3G+6d07K+9xywsmaS9vvBHCMJOK3lU+ixig4l9dT1KIom4ysrbTbZwO5rs5E
gUFvw5qdRrSgF0Lby3mcmkwDqzoHcAgSa8Z4Md9uudp8KZfUBK6aeOZ9jJj0UX6JNGwhxugHZhqU
+V/bY3RXvYSlBPZubGfYh+FarekC5fg77ZoUv+mp45nv6/QrhyNlO+WT72T0sNh7co7BShHvutDx
Wyash+D9zvRHaPd2/RqFUD86O7iG+fupvuxzPbP0vQRY4CDXf9MmyXI6+fN8kMcvnEJlfSK9K9T0
v/MnynCpmE4pIjORlr7u7QYMrrQ4X2TPKA0ivOVlHoS9qcq1//l0d+c/0fVfWBTRVfieGu0gvIqs
26YQQXbMJMcxlr9zBNxftynhEL7icKbalLLnqa3VELaq57BA72SGM6sfzmcd1FyPF9iXGlhkQooG
13Rulq8Clg8ewCTh7W8eD71diqzLLBeLJPs+qAe9XDYJLDDs3mOIqCH7KYB72Pch8P4Cd6C0qKJx
rl5OXg005G+DH17kLaYCX59nmsebxJm02j15LGDnuoPPi0Rg1UlozhFAh5PUIOwZ7+lm3infXJ4i
z0nlDRdE1yLPIRSuzB/nz8AoLHsHpmEoLKuG4tFGWHZvE4csgMxsFIAdH7bBRVItzb4GyG7pWpXi
LEtKW+mXLzDNiGl1raL1ZQDa50T1XPv3XQ+2v2KmnOIekAaIMbd/yneszTl8M2+jiDbAkYC8mJiy
0RXGYLL8oxOlXEr0AXWHPCZjyfa2z2LZ9l2spEdOrKCjqrupOaC7kPg5uLyEgGaqMUHOxDprdtSW
7Um2N8Wn/FuJInGz5pcAPBW4EGkSZl734qyIDQz/qdkoD6Knj+6aRvtB6ulR8ZgQtgfJ3Yp/SS6P
v9dvWsnQvQNnr0MNEbw5CcFXlLIAOCIUSdO+bhZYPXYHizgUmtcumto1R9elCDiMRVn3vC3sEfaC
jKsNmhSCIbU7XL2Acy7a55QZTRspGVzADcm+AzfyR3ZHuzEYJKLoj3HRr9KqLTaFKmLi1VltGn3R
RhQ1OxRGQ1lF7KHx64S2dtORAW9vQsNH9bBoQo6ny6ynwEoq4gti8eWnCrmG05nXH0ZYVaqkZMQO
0Sr6NHo06er/mBCCWu15iNqmTCpyzoKBc6+GR34nZlpUxdZbwolebUPUZmGXhQyoUdViPQZYchcL
8oOvVmE6xMHzwjsSDM59DCxOBd2Z/pNQ9IkCyvoqL4kt29iu0kaenhoP3NS6lRpm8cLmTnKPmC1/
PrzDBNkjJzUb0UqcTauLHwaFH/naOrTr+LjmTWBZ/ZVWQ9zN+x+8M18OKv1TbQgLVUwmdtwDczWV
MN8dWM88FyKXh2tvDxm/6ssMcJMrn5P6+r+LGSUfXxeJRQwvG7KKiasXIewKnkxnw9yXCr5bg6n8
wkfIb5KbFfzscq2UKQ3D8c+4Kgc2jweThwamx0dqVvv1lPJBzQBtl+XEGXkck4LyxTywI5Ahhiet
n4mYG7D4PNrbmOwZNkImUDkpi3gaEbf0P9p9Co+76eymvPxM5Y6hfMFKCvyLFOunLqTdZ7pb7rvc
1DQT/xoZzZAPErl3ikJUPX/qD+AygsTRb8SUN51uXxG8RDEFXiEoMQSjSFFDbA8LpmIrns9oB9sI
pARZbX8LXG1X0NIqHehFTEv1zx35htTmtIyqP2Frrz8HZyUHJZsYEk+0QB0MoFcUScjdiPVxvBFE
ajbN2p9gGKUJPeK/Je4NKDUy94Eof0/xmc6Cks6L3ZeRdNd9Ut80MbXlWRjmWrcpIAp0AlwJxrjT
TDFqQrEDbzY3FWtROHhHLRJJZtqWPo/QVOhQEZIMn/152pDISbgFcO574buRh+dk4IMXMxNVsKxt
mmUjX45L/aDG7LaEOl4jATzxH+o55cP+XOWpiSbHISdA8bNHG4cTBxzFLVaLlnfijaMIXA7VCxcK
nA8DUhGkjQVbI8pfnMbayR6gim9tFkXu8H+fq8oe7zlCUepntE1ZiBIgU8g96bkGFdDc4zKLfBtO
pLMZGxK5rmqmEeNuYDxv8FaHScoGSCqCvFJhk7i9/h6nF4ZMxqmSGEBoJUuMInw8AQEg+6nFIDBw
FwnXkWTFAxq0KqlibWAMmOZ58hPflyBF9KsPf/ZP3D1KHm4YRaNijiDK4Pna+VF+RHr1JN2qWv4N
d14+/cHOIjAPRTUQJ/CrK30x6QhzJ3cJtSRr3EPdiCr3WeVk5TN2SbUw/URYA0Z5Chw0yqU8Fqwg
XdTZOf054FWm4/AFYqjhjvPYRnRW7eMmEqcG02A5mP4nYZzpOrH1lI4+0rkXPQFERKI1BREhmU6O
U8+aI16jIRFHKBjoeQid72Frs/h+P+fuDzPvTBpejAVN8X4aEORcgQ6I1ZD20qFqMUZHHgPPRci6
D5eQQHehP8kKFsFHEsUH74e7dFlek/lIVMR1e4id5pF+21ccThPOjnMYT+jG/TawMuw/L/iQl3Y4
T0anDR+RITKls8CWgV30n4BVriuJ0CwUrr2TVMagdt5zTzQjQEQrr8LPvQM5QktGwR7tnk4rvbOj
sLyxYQUYVOaehhV+9ALm2mZWKE0bCtU4HihVTZg4esn2JIIyZI0uH8/bkDygSqjzHb+2oh1TeMje
L6wL6Q4POFj+ec0493xvscXSBcX9AKBcylJsJ4TpHJ1cYrCAG9RfiDyETQLVX3oQp8setotiD70J
/uUIpeAbfbJZgyBz1bEd7s/tlxCVHC/NIN/CuQSS63eaepwG6Unr/L3NVoJbJoyfWY6AFct3pdLM
VcLsZrtJK8PegOvbNfUSFBICSoijCnoOFlWK8BNg+FBfoBX91k5QmhqoNw7vnJr6Wja488e2gXkx
oJUN1VJlHke+F3vzNuQdHfQ5gdsejkdiYGK0Fmtm83MiKU1yQsVOiYaauM2Lrtg3RopTHZqez9F6
+0WAyic4Ufot/NUwvM//ZwlDf2Jcc2QXNEGenA9XFK7evRONf+DyaZrHIu50IPj3eDcO2PVwFfNR
D+sgMLQZJPX7uXY5F/4p0QC+3bujxQe8U8eSujaegCH4VPzRBnC6J/2CcYZXyfqB0/iwMFuF3ILr
IsmBER5jhcWwRkW9VVkdYEjMs5nMQ8E9WoZxzUx7BKBLvlbKPvIE4+xhmWkUJvx5AgpbczguZ4Mm
5auSka8eB93YweMlGtpUZsjpaw6EAbQl8lnhV8a/2uP/5jgLNcqcOmqtfNfWqAE6ew/P8sS2PRW3
ExkqCL7R/yBd2VKQF+HGisFqeebr0bK9SZKrj15ki916xayOOUHVJQmCvC+J07STY3V3xoNiBJ/D
HcFSFq1SNtDIla7MbcLqD1FrrAaU28C5aAxAWFScpy3NNFEol0g+7xVBT4tEbQdVfWp5k40R+0MI
dLJwJfJ1k7aOmJwywig+Yoda7ZpDBng31nR6hsxSNTsA6rFq7hdf8aaZl/erm3m0pNxQ4zxyHzgb
uqc3Pp6xG3xcZDQDOiuNH5BP3THC8otVAyyLnCaUnZumupV+ROCIZYUPr49YYoumjw70/ywQC+Pv
oF/gAFKTrYxMPj4nFEAGcXxKlP4GysT2DL7z8lff3pWLdNS+w7HpZiSFF+3nBW8ZeO8JHjv3sNoO
s5odt22QJO4zPNgrQoVBzOXHcXhKfkMLmFmxQ59dTberkw7wddBIfu20E0jg43zojpj0wRGrvagK
+WZQbXrIeTAuLy3Vk/AHWG+mYf5KpyhgBlB6Bk22YfjqjsXjfPe4HdHBFlWgZYg0TohqfKWfoa4M
X8NnNbdL2UZMjfQtHdr9jO7w+WPyVwK0wxVKoAUS3PbiPe4dwabmpTTqKyZW4lNpAnWB4rgSEjlQ
D4d1P3SXQW/E0c8sZO0519h3+Hs728MqNH/4MlkIjhWkRxRKet5Ki90vDVAMVhLkFLj167DoMTcT
uYZwgaeuQPGY2ofxKya+rSMuISFFBmFmpziPDjxvn6zkJD5QsqS1WIZlEezEUA9EKQqgGi5/MmEC
YUJncWZsTwNG1+0P2jLx00MT80hLWUjxOXO4HStghKWvgjOpHYha82jPDTUy83x1fulNk1hPB2EX
pdOmK5Vgt/mja27g2uqmBsbbyaizQ5O/H8noA4lGs3aIgPTJBIGIj6a7bsfPkp3ccITZjpv9+li7
B+MCC6P8ngsIHV3Z78OF3SI9QFuDYlgoq3rW4+W+AnzNOqglvJf77CVz5dWAh6UyRwPTZZJVhneA
4OocJzf/zDU4BqeV9/dgN6jxsU6fssqb5AZkOMM1aFkd0yt8IKBbBgdrxHIOYMn7VEPp1KrrBNX7
6ydf3xUaBKmd9gNt3afaPzFMWVpE511Gf38qZ9BPaJbbYrv4vyugQYAwGOHXAVjfFJw8pXac/blr
fWKcEBU8Vq0wlss6AwKazpY0c2srlxWvNa4sTluhi3agRSyxST2YT7HT6J9NJqLPa/GkgAWKi3h2
aMqo6/6x0ieJ0LaoB9YEDKE4W8BjZg90dPaQvO+ICDrKdI09tckRb6DsGOaoPCEAVxrbaqmC+1Qv
rc49vs8ZkdjtIuzvlHxWvK53R8fDBJYp/NqGHbBI93qBPSZm+t+FOOx7IRy53mtmjFysLm8z9iCa
Emi7WQQbAVlnZe5Z4/mvTcXFlGIs3sdarRYWU6xulCLMQ5ohN/oRdm9WqtEue4mgyz2G/ZoHtrFw
rBo699o6zwrthMiF62E7vdGjIFUOHhnBgqLCEhh78FpZMbxVUCKAeheRdEu/FBj/sFNJw1QbXN7Q
GGYPS3RVhOPM7eO3rOoqq+DR38uCMJog3jY66h9CNMOIwGLkGzR/F8hCN6/OlazmPxljO9IjkrBF
gCl5XVUPOxZzEl3tYwYWrUoQoA59grEIpEyUqmUUT+K2xo38X7eyT5lfip3tm1MHp32L9hDEcX4Y
JF08TKOgqlox1j9QsuJZzw74s7uEYuxSO2VgfTOORP1cpS6cqmpzQLif3cw60Cz/ry9Hg1aj/DqH
iHJK+YMsk+B60wwHrvhwVZopo3ayzCBYRjfXPLiUu18wm2tMdNb9AxUdlOjxS6y/aBuagCTvdUN1
qMDdtNDLHUJ+PEiRXHbbezjnaBc2MuGNzqPTQKeIX5lCYYtDzNfnMwbSQkPiA8alQjRn0ZQKuiyD
AI8TA1CNQV1ansDiFgq4BN+Wj9TDurO8Cdw8IEjq/Uf5f1caIR2LHB+nSpjLoqbfsbv6OdvGOToi
xemhtw1s0xj5hVNOGhmQTmT580Ya26F8b8iI3mHgd2cVjkxOd8kP1WYocSpmQKDOSc9M8Z1huOMu
cJyi/MUKduEJkDrL9sDHSFLiQeTtnYtw4liD5Ucfjct/bB8uNUZILwa0rnQQNDEenOJu2GSj27jn
EVvieV+PFrbR5wNl1f/iAoT4XBJs7DtPMvESdYMRunVTqUTVybGRl3rZnZFA67S1TTnJ+92KkGxV
Zqw++Jv7W80Md90GfJa0k7TN6GYJDzlaawgwRvHNoDxyd8gnhxyDdk+MAozvsjSTJJkXliQ4L1QL
ZxZKjmHp6WYXA1h+xrhIVnMKKzmkzF5Xem7vba4MVOWtoVRrrqwPjUiLkQyOWFQ5esrwF7sJdisn
iwUCkARNDUyX55+iOAQbcOJUmnrJQ1r/HM6SXYUyQehjbPcN51LH/1/bbg5Yvb6MF0aMv+pm06xs
mFXrjQgTPve1evcnXuCQ91lXIrnnPV1e6/GX9PvfZ3LM7NNXBl7OEVtF5lp98JEWwuAq2grwT+6M
O7KYd5cZOXLB83cJOVw8nfrHmhVUYRdwhVfy+4L7JuT3PEEPXhbyOyuClWXneJrPthqrbmRSWD83
9C5n344OvOGx5Oqa3N1HLYP6UlM5XJKyyxEgGdYgfW4yifZPrTaQIb9vowhLWsIfk7Z9XW8RMhs/
QYyMKP1pB68afr0PTHGRS8kwx1SrYTDhMlqTM9IW3xRWr+etViV73MEffMCQw9t5UDl2vrBb0uhA
eNFiE1AmSRNdsMoJk9Pg+sivJOCxo9ZGn9oLsO/dK/P76dmG19byVKs55Z6uWmU91CbNexVeM9vG
0DmCf1Q9LHybMwVVjBYIOqUPJxjIGnMDwfrZJ9VvmSCw9IkshBzFgW91kJLVnADM114W01ssQHsl
MJgKqc4w5I2pIj6NjWuQ/NMhFnB0WSfRKEL/iIGq3hnZq3QS2zzRl61kBg3KLgZLbgsh1eVKNbsj
FdkAwegbmEScKrqvzusC9Z6ZqYAK6otF+WQeKyiO8STq2wWCwDVWg/Nv9G/EuIGCyXGSM6QfmtI/
/LfgzsmC27NBEQtVQHDKu+IOa36+BOkMNcbCrXVdlWAQhL1HxbYrTbHA3tl9VuQ/nQ8z89090pFY
h0qe1w2u1MWGvza3c/3u0YvegDRjVbmMjPlJUagMy/rVjpqZOy4cPpTraWE9ghluzyQ7RJAB4raj
cmPct9UIbcaBMhy0hi9jc9I6V3gIWsh/7pfNWVBurcZUCvFUTF73VwB5TOBu/VeTgSYfCuQggxrX
BwvJQxnuqyxIwcHhQ/ZtlrWAARC2hJprA2V4/AYbnoUUZOfzSiycXh21W9NaBVZhv2yeyD9xKnBt
tpnmzEEsc9tnY5KJkMRkPk7H815jl2cWxgnzpcKatPjxmnTYHwLkfqrRphtdPUBO8oCT7glZMwWw
AaD3w7M+t0RJn2RzRVQNbbg7QWKUzIP81UD/Gsk1dxn0agvc31nvpeo3/oqCHAN32yv7NNVmNPnB
IwVGFdflosv2I8dOpk1ez3ySSY0j5aliy4miX1jYCZgKGxKk0K1CnR/dhcJfgQMRxXf9jqvuMrxq
qlNb0eL72jR1Yg98fTeJ8ZVq+CiFj6ypIhwdz0SgXBIsAzuqcEvP5/VYPQBDcmXby/3+KNpmzsOQ
0wNGQh0l1vCNKyTi7tlFCXap7SIE6wClEKqLd1bf5pycTnUFzqbfDRlc/SfxeI2tlyG1NQR3zMTn
auys/UW0xqa+6ZwkUkgfP/QhNqvi++BxxYZL6FnfcK5I0i1YtncLCWdLamoV5sNpOidaJ8Vmwo5k
+ecRP5OmkOY0nOQkrr09q5EINE8vT6ssrkMhSo39MmIkW9vW1Pxs+/91M+bTlJEw6hquu8+Ppjlx
gKOW6bae58p0oAsEqL8PyTV5hatpMZ3TmjhVefUcTfTaNsDKL3hlunWY1ldR3xU7w8iTNfHJY61Y
2FlI1k3wsNWmRtugXWnxf3jcJvyVMx215QWm/qqxTb60JlHXge4i4uaSLgAo61JG4qTQnrrgZ++3
vMdDg/P0M1vi7HkX7+LMC8qIqKBrjTQ8AXe/04zpyjYTF2dWkyUAMDq5OL3lFPSjc9XqFGMOaX7R
iN3ajZJhynlLE9aZ26dCgMfPlZcuV2RJT5mKYBBLNNUF2TLCVVjU7Te7CMN7g9UPT+JK257/JDh5
OkwkFgwbyRoMkJFvE/jj4zpSFkLnriEJxzsDo58o3L8ft5gXcku0t83ilVM5NKQQTmIvduwA+94b
PVpv6gPUvziSxkMTmme0J2huyYxPYAyEFOTM0JOKqX4G90JmUO4FhdZAislyqUcM/brPDbBlyhSa
hx2DATaDcABDOE81eUrJhS/6rcNbzpcN/KHn86mV2tUtNcptxDSkmBQIR/ItMc17R3EezBDrE3od
Iq0XXf7H8/e+tRAEozplmfTel9ILRUmQw5qVGzP1z1uLZgbUxnSx1f20uzFcc/JZF6t1K6DdlEGR
9N1XCw0YsndDG8Tcx+rHqB+tEZwnzYm+v48UqJJU03r2JyM8/Jb0dwOHZa3NwuqOTFB+YR4izZTB
kwH0FqMEnTAPIYhiA0OAF7abL4ur+sOZ1Lhqr01G5Oh1ZUCWVS/PsiMEi5UMuMgjLFt/4k4H/DWB
qYzQJtTsdugRlXpnlsTzORqfjwwj5dvaKfjFEDE8pjYA7+7uxVPrKm3dBdjJCTJLD/VnfmQ0rjEH
Y43QcZe5rBSBdN+dkJdNEhRmtS7kwAK6cmK0zmHSp2nspNb7zYok0QGInQ17s51yBEb3K8tLbVLw
AN4S673l4kB8sq8IxYWRBTS1KLsWIT7KHkh3A788ob40ieR1e0a8CyOlZQxuOr0Z0/9kH4+ZPokT
RYUzKhHZY5B+DRzAV0Dga4hYE30shdGjUWW0pAE2XnR7+Bb5NZeF+qVcWS1o5D2fYWWOQ+jwA8rG
Ahrjc9+ZUh3O/iijASQD9CTowwfzIn8wmNMmc1R6XhQzuqj08nQWTkWgYTzkRcVwMNZYULpJ9s0C
K5+9rnKI+Jl9QMM06avGwz/TBJ12twlST5Q9Qe5nBdGEhyBTPuoIN2SD8eKusClH1ODidsms1vdW
HaZjsiAZujr+DZDNJ2GTa0Gef1XrI6HSh/F/WQzS2jOPICT9gRx/IwUxeJFfgzLQNrk/aoPa8n8W
LIZqC4enj3X7O9NhhhNqK+leFosW5lEyY5OeTgMCQ2ZCrueMnUTXLWzYDjBN0OYvLKk/8FPtO9uD
7jK/KNm6Msu8cX4X0sNcX6l/e6+otxRhA+nGAapFmv48e8ommo3w5auBFcdCBYwWiu+96Ah+DHJi
3N1QivMFbYN3T2mwXHDT5CoMKWJfDLcWTXSKvoAlAWkGjmUBuA4FReraJNERCza5OASgdsJgMyZD
pinXfHwF0KUXFEQD4221nMTwBlNNc0qrzukhEi25T//VMFmk+l72EMjM2Tq6sxW1r2FrPArloHV2
9QFyie654G6vlZoGL7A3CyQno4OiN4Bhx0Cc+NEMss23zQYbKnG+4h/KCoNWET0aaY71jz0gsK+k
+a5crFt+lAz4KmC9rSTyu2g+D4ZGVGJTXC8VB7M9DX+5/zaBFD8UhrmaQPth4LSSM5x9xtY8dUUZ
YU5GvQHoG8rW1As1krPcDswqxqa9mBpihHFIEVBzpJojmlHdXyFlH/0IGUZ8/oW/XSMIiNHbxYWU
xNoK9vYCJTd9S2iRtftMnJg1x5toCOhTRWFtTgw3Y6DDV4d5QfeNSOpDMEf7ll+GcL/J/R4BG2FA
AOIOIhNTKPEiyFV05Ge4YYzJWICKhzKa+1zmwT/lQz/PIwboWfS+6muwYtJse1D6hcHuwDTGfDAT
SRygeElMXhYYS3QBL6eBAMwqFRhJuFg0NEneltr2EsQZge0e36dRmmIFkjqeoDqJWUvAeq3eamuY
GyxjCPrVY2gfAdYPSFaA1FVeABfHCDTrxb4Rek9Pi4PCqYVFPh/ZJ5saH9e4n7bE/+zbJqRo7udl
XTy2ATt+qnK6lCh6dnAKdwBmTPHwVM3er4CLIwPMAa77B5bmVK/IZN9kP4ctv8FYZxVBBLEub3+J
K9I3cRmWSsoJqPE7Ubw72Nb6BA3N/bUuBCdUB0V1bvpMLhNiKYMJhmXylrVo3bZs+8VIxYXepZ/U
Ah0BnUAZfCbdBBx6hReua9al4NdfIG2pYV4Y8IZyRrhIjA/QAvsgBLb+WBHwQZ1ok+QurSv9Lupj
TN/skbKsPfnFH+6iabPAQKD4HxVNmuemulJjWeNne+rVVHxHUfk/yjtUtVEuEhTy4VenXZBusLHY
PNgm8beZ8CqPiqOLm8BLPTeNm1PDSxyBwQngMU5WNGqnG6/lQ7uHtm5b84AvS0Ot55xDXnPj+kWH
wJOBZGIDQ4MhqvLcp4uBxc+SiJwhtDbjtnJT6kIj6Ypyr6dVM/fITnW6jYKwbgRxjPF3fPJ9Pcyz
owRcFk9N09hgA3ViGPAA+qigZk3pN3Ys78S2c5Y2Qn6/tLCm6JvxF52bvuWEkiQWXHbywS+N2y1z
uzo0WQSC5XzBOlEewLkGrlVDqjc8OyLrVl7D1QGGweI3JRnoamS56GeUCVA75TpTGqKg4HCgEWtY
WEeiJSSurcReOobHR7wcsMwDoUNkrwgcOKH3qj8FEy6YMWVgknOQVkY5FP4RkASru7yyE3q1bRcV
6pWC/lCGQ5oKo7JRtuKo3yos0TLu9svE/d57IcWgmpbweTaIXX3n7o/LVkPvZ1hq/S0FMIaKb61n
Efa1CSoi+iEP76kSGgKd62Ir0NZZ0QfkqTo2OQESHwjjjjrG/H6SplMf1aLB1U10pFuOHzI04ALv
774vMkgk4xO5C/SbjMhZok4WTzvAl9Cn61VBqzSD8TJHLls14TXIOkqqN+5cyGlegk8vA24bnFlo
tnDQ7u5nv9l4ODvabsWk0Nn+c4NyeeNI1OL5ZW5hR8WAgAKEIgmtHRNcPLvUxzUevZY/BjvwM0L9
Ad5M3mFYQBLFAaj0sPsP2iGI/oWpju7Bu0u54w/gnB8wqU6fy44dsJiyhGj+b4+4aWadiTtCE1QS
9xJRVlnUlq7ng212r4GOfmd/cnhguhqLDkhF10uegKjCzcqF/uJ6Ixr9maJfuYhQ/EIjgjq3OEZg
tcfeiJDwhC2RHNChlo2yDOcbIq0GoHm1Ln92S8vCbkuMCV+tNc/wCbT0XT4eyVVPtquG4SJOz61Z
5GYh6DrPEwh/ArxofPWSXY2k/97BCoMSfwtgbnXHv5Fbo5+6IThY78C3N94CcbthMU+s5NXC6G+t
sYtzWksGyHmCHqSNULJH6942OdQLGL65bPqNmRs+/BdllEdP/loGMZDcH6YXpQuZqbYzooDaU02S
yOP0+sAb/lKRC/ySGUK2kh23SFvGuOfpUoIfZD8rD8HukQQ5Zxh3lHqcjuO1Tx2csuWPg7QHGa1v
esORxh4ut6YQqHQrP8q95w3jN4vtlPrRVaVC+NKHajPGVf+H829+zPvocC2fIShShV76qFtu1xG7
T4HXepSjRjvu6OK3uID8FR/MtG6q4+Ba0eLYvqGMhEHdb18ZA64TzL77J6Yhi+JjZGA5734MwJ6t
H7vj+WNjv+AjVk3/JBt7izG4Lpwa1ERxRVKK4U2DjiLhvbSsS7UQKURBXMQy6BAjXRVJW88iKoHf
mZdGJkW74tJhrOqxmMMc7kFUHMh35496wLgTvXPqg0KLBTMI/SGpi4aoaHPcXmABjJ4gak05XvHA
8GmHERpdvfTq+6FOYzGX0tDuxmVCyq6ohFx8ggAgaTRIzMEsQt3GtTvNsFVlwrqGBJZhoUbd31QF
0Ss80PpDOPrn/7tPzFTnKGoUwriTozGZqWP65MHZx2zdFK5qmw7TsfWrao8elVUbhZZ7DjhZo5XW
Y/JASqmzxp+vO0uLTbj+eZz8ecTCFW6K+xoUnJSreDJqXrUl+7sRTnDOo6eVseH2AE2j+sEgXept
TCIxQjOXiHPbwoGDgjplLayv9CTJhVuDPsLrFysbV4oMSx1axWQdPpRCzRz/e82Mz62z3LjDFqe5
lwaQHyeLKiq15heucG5oUmg32KocF3LJ3idFBfJ3XVIUALfV8hXXpOV53xtJC7cW+XqgzLAhwFpB
RIJzb2mCFyp9fNbP2DmdiJgDjhWLPjocqQRevTZYZ99KoOKsp7CRIk01GoAUN7R5zS4bjaBCMaIh
6BvAuh6nsB7yT/kiGwD8AFaXhAaN++QMbrKadFs/vtVTBhR8yn/1P98/+N4rZ7UB4jcUR9eAD0+t
lx8xyg+er17E4nDlf0oT8M2CW1fAY1EkqMPjqdnPchYFs9F4v6FXgKOL5uaWYCv9p0SDpTqAQQnQ
Z7Wm31Ks4eHUTLGESgY3MEJiEpbQE0/ON8fWGOznKu3H4bQA5XL+uKpXss9sb1eRDt1oUYiDxXRd
hl95iTjWVZdMQkxh3HFn54JTCLqJWUqzoW3MzHMGE6Dnht+TV1YQNKbRpIqTpLjzkRHWdKRKlI2t
i4h/RUg+nHDRlBoLJkPcr0DoE5G9EUkFvhk2SpxZPm1gtTYnwcyO8ryn3nt7B9+ohwsAo6314J/s
uXC/piVBMiFcpcw1BHLHcpFLuklb1eQUypNQ2H9x2GAIqXHobEN7X+fSHQ4NWnjwMxrTCkeNvfkE
g+F/qbKlJXCA/1gTHn6I9VE/UALbir/NmB9FQuHDDY2rNBKW1AzejiuW8AnV7PhaDaGnT40THR0O
OHkcCENsblBums0EyECcb+J/Q6Z+5vjvhSRvPb4eREgxWM3wToLdKykTtNY6utPT/BFlv+daTnj3
GooPLZTN6+cmcPDzeTLqHbEn+YBtqwnkk4ZVWEjIH0AfluPJygQGjwrQ0DSqTW5rroBrGSGyicna
WRfrizQK+vMdYgMi+awpSyk2sViC8HdHJtBspLJeHaUkRLlx9FY+hZpznpIiOl7b17DyceE/AuMD
ehSJ3UzAVgee3chPIej4gPPGmWAfbdYh6PsCpIZxtTrY3Jt4FyQVPVWWX4bzjvcuTOVXjxrzF1Ir
NYgrQfjpjWlDP2juNYMJq8sXznmHPczcfO0FjUDdsZBnOREn/Ry7nwVOCIACMW1nZJSpua4qgIXv
rjEArZObXEJ8s0FeMu7DNYI+WPfOLYS2Uz4ZS3CvuBhtU0p+7Zvt8LhiH1xWvy8cgInZ+9oOoEZE
eIjs26Yf8ZpnevpxwhrTcAD/nGQC9DsDb200XKqcPjmZk0Skkn2cxSpUzTVHDK321rH7jUx3ITnu
uI/eNZrKBEDz7UUVsCY0dt14JIQ0lDPOtBZRMwzwfCVdhv2cx6dfJ33AN2cy/LPLhAXOwK01+Lvp
PUWtkzsN5MHyFEG763aBadjbqj72h/5RyMe9ti93qmYUYmDG2a0wnU9rNLwa0PXrXhz2DafT/e94
Jge2nMzhfPv4fM8AccHFQWscNMJcy26PczBHOM1+BsLHHkFcJkiQ57h9yz+aP0Lfx5GBfXRE3iRC
EyY6yDmBjElovv4EoMrT+kiNZn7+Bn6HPzS6CcPgZQYkVa0wR9zJETzdC1w5TzXvB23qKa7Pawkv
PYTJM1wvaU/MzOsm5+NcU4bDTHRIilDFdzL+cevF6G/PUJVrKSW5w1iP74VPhMHRskqyNESGvg0X
nVtH7JPl6iUkM5KsBPOevTmIuof1L8U6PHOfLyo8T8ftBq4GiAu9q1Lhj9HqbhllVmxwb0mcJSuP
8JOqCregwOim1b9DYvafaFHTBzKtz4Vx6KXYYgDnF/6DuvbGMkNqX087zlaw3Ci5VcYUijlEG0uZ
9Oq1ePZy4pbrvxa3eADupOfuoRF1aiHKLMDGzHW5Yl9ySZXEYyIpKSYhMu2tthuZa0sgfWgzEAli
akuHwyqN4oIx2X4vPBry2o5m9Ba66LoDXQNtAAUIceIMQq47qx0BNcl9dwkt77ZWumhqX6rVEz01
vuMLIaHuLcQlAGl21QejHOtq2zvRapxCkO66nFkxArjQwYjCq4/Upv2E7056r2N44ICBFMPsQtZM
GCJ93qbmHmqJFhBINXH3ZCp/jTx7VBK5MPwtj3N0+m96PQ0tmqru/9rqw7RZUJJ0BA0hY3REXPuY
wfc7jjhE+8aW6kYSSwTCGUm8fo7F6DU/IQTsfE7evMbI9w0m1c7mM68fklNH525XjhIg9Yxq2yGo
5PUy/UZLmos9LFFaXMH+HNKEIe9idnbMRhUKy6KKAUrCfHabfeU2yMW8uTY2ZWyYyWQbI4QyI2Sm
Z7L8S3cgq+oflfOaUuqDkbVii5ATH+SdHC4mqdUou/hZvqHxT5iHl9ObYE1f97ax4dZgHxvSGme/
apRYIpjTdS4iMkeeJ7wGl6fvq6tD2DPCyfSqfy7/iHv3qW7BwV9XyKutPnfyu03pHIDQpV4D1oVq
32WIdvr3esXtTfg3k1TvdY+BRDvLOlHDFMWgzovpET6kFHLwe2IRa/W0q9eE5x63KrC9U3mwxcQt
zXFOLY1Dmu0ZrbkY+ZsyCq7c2GjPbyMtvlZ8iTUkrnp+75D1RK+M1wUmx76JtVByA1RPDWU8665J
27HFBsGjWlFh4zQr/4GcyQUHOIS485ghZ07e5IRAdNdq0taT+oB8EHpUjY0KKkxfpOsSg2THay+s
FuNRrXqZbR1TfANXWLyWW+QTqMwm9QoDePdGzC/pEuD2ylGTRSK0/dJWFA5crcPkNaVARocLt6gg
oULTRug7B3T2m3k9Sutt323VQCkMNY7olekNOa0iyi5q4K98y04PKMMKmVbs6uuA3tJQk5Q0GtC0
2we/AKFrqqmcKeqpvezBVaArMJ86PL9s8B0d/h8BTDYm+f2dzNXujW/HoaDAhiPKD55WURQw9gMY
C0IR4w/W10dOIS3x6qepqfH1Qlv5S3aqmHYCAUxRFXYqHOZjyHvV04OleWXLav4pcZ570HZmYQ6o
q2eK06oe7sLFXZxP4v6csJNqKApoSEPkyUtbUv9i4tltHQURpooggY4aFQtcqGXgoBrOcfvW5wtD
6JwhwHnUTc5x4RgNou4xMsZh+0A1T033bVo4HT4nJ76ZgTrkEVEjbo37Kwp7GFSO5WYGAhOo0kU5
04NErSkem5k+phzH9tWUYDal0JJ+u+uXCDtsytmT8s8IO69irso9MDF/B1VGC9LhpzTlO1DgVO9a
p+VFp9Kd3ZCbp9U3pCZrg3tWajkANTnaSFawZUoBNtHk/TSr/RpUTnjXcSdOXsjIvJkOszGObPLS
1lt7TMnTdL3SGjRxtJy5pwnl4heRUr+/IRIEAqZMcMLRypHipeA7U2T2KrhktBkVC+jVFCb2Cs4V
7GXmPJukREQbmIM9JNpoTZLEt6FPsM16V8FEjqJuIC3eltfIz4CurBmBEZH6votR3mOQJ7wfKime
eTL4Gd04AtRb/HUAR6ZNG3Pca040rvMsHEh8XhBWIJFUck/Uelx57WC4tf6/P2xedo08WbZ66hmk
irWhQhS4w5wEg7iLW3idXO2k1hDZN/bhrJzbb6Gy5FFP0hnQfaOKDQX0xDH5qNzp5b+C0MiZgtLA
7poM9Znim7G2SPen96ku2oXbATlBLIe2SXrMYDRxkHxYdOjSArJd2KeBUp1qn3VbR5tDW/o5RvOG
bURhxJ5C02pk+gcJajZlaNkUTTTovFCwaj+1pfAzUOl+bXxmzM6FnH3JQlk4Lm8SfbCunBmLQjvt
Mpp3GzeXOjXm3TcC1tz/TeD4CRYweagXyA5RB2qLQMBBu/DUG6ocG8sj6XdGzGs55cVbDm64YEQ+
bOiLMVAcDfy4cDDDOl4Em896iypLVElnTbTV0No5BmUs5Ym/XYPDPiDqts2apTNO72BUW7xQkW+P
6T89ga5zexpswlhVol2l3sy7YAyMiEXdcUkJ3NUNFN5kffevz0qAfgWtxOW2alT+VULhURzbugTL
mVqAiyvVzcsGLlZvNXHMXb3cx89I/sP24PqoSdHR4Yzn5Po3AlQx4qw4dfwDE4/HqOxIV5/xxrw4
tnJ+1wMncFrQvesWPJmSSV22M542KPI5NvfyYEg0gcxD/sPVHMXpwLUtTPgQ0H6dPd2PXPEexJVP
SmjM0fe4pX0V41xVmDPQCweIjm7gFB9bt1Xqo3iLfeb5iAA/UZvyQfB+RlPr3j2Yj1DugzSiPiEu
yaLgs7sEp4VNdJ7AgLyuAkXTnN50RIxtP0C7tRw7N1dZXnQ2x1598c9QxHuFCEyOP1LJqJiKkFRn
tpFvNswRQYHe8uSkoIwhfKB3WbgL4EjiU1QArEOoFXHfTrk70Iu9HSyPY2B9Qv3b0yu8oTWabbis
3QPOvvfy0k7KgzdzZSvIKFg4r36GGTgCJ/nPOBOgjBmikW2tRFBYiP+3Niq8IqRArrZFEMU49GaM
2FvuKIDGBMycgIfBjoV8XOSXm6bKGf3rQMXuqnwjgDq3FONxXxF7fkhgxtFOQVRYSE03qLrvApGe
o/0SUuvJv0OvWFWt6e6SXYit0SNr/09vwGRo2l+KI+n1elylYz/acOxw+5I2Gl62NwYQHX8vbeOy
K31lTpp6rUnS342ck4qQ2A+1yckhtuk7qBnsnaKg/6B4t/bjxJsjyiGCyxzSeolsgflX+dHdXe0j
Q1uLG5MbHaZ+UiEAFEtiCuIBwx+xr3nrw17IjDxb1o+euA0/ojBi+6IwWcpFhvtpGew2oP5ckp57
qDyj3MdyLFZoCV9x/qJeOMjoyTrNfG3TlFuOC4UII/nnn8OY5YVXLXbe8dVldslNcJCJtDlG9ZDy
8icfggEWAVRbDj3wGei54yuiPrEYp/iEmQXcAz9VYY5OrKMF24Erv9PtGeZ9zZI4tI3urO7RRoYC
Jxgs6u7PMdVLmiwksjKQVmhbC3TqnmgPl90zwg0YmZCSGKGCXWwCJHrBkRb5aFLw7g8fltRgU7fU
fjPXnOj9LtyyAqP0FIAdx8AHRcM3djw3w3ViPu/wulYHvih6FYe67cjbQ14iR5DSKho/1QS1wDYi
pWu4oHzCaav3ikNyCv6GUbtAjYByMbC3NM0nG8xSacHZCPYJptGZVqVmLtOj/3eOyfYwfRJqi53H
oSVtVL2MPeUeR8R8NXjwBbtQ7RE+59qvgSz7LJcn8Krs7Np8aX7J0WwwfFJIexsjpvzMmr7F68x7
w80WGN/FQTJEYWyjTevHLZbuUdc4l1PBVtGZq6fVua4ToI5lFtFa4mptKcPK6Wn8jzZDZjGEhvHx
oiCgz+U+R7H3N3I5ZA9/PO85JJjauXctggVMyzwHlkVl22ePT2JnqpAoK/9yKM7y/+u13c3m3MvN
7XkH9Rw05AAAGU7efNMmk/Iz0N1BE7RM7oEwl0G5VxmnX80FLNA1uBqv/2DJUpmP4xZZspHIOc2l
DfKs2Qk1yDcCLwrcXe6bhg0oPeD7afEeHGqD5wKv+htSVPV+IyR+ipcjrgIaEwC8EwkVQXegW7E2
sV95I8Y3PD/obv2bjboiyxPw6fTgidYzWE0Fq1tIwxdowgzBqOTyyueBCk8z8fgnJTw+uAbiRwtS
GFjtyYFhDqqAPzpEbi6WNiZsw06w/rd+61A9j3md3+UUp6irCtmf82xBnpwNI2R/2j8tv8o1qE6B
vi30VeBYs0XaK8SVnzaa4/CP01xvUiixwqIbE3G+k3rDAeGvy1rFfTBbjoIfFRt+nTnd9trWX4cg
Ibv4bLhdMafwjkgJTLWtRzccY7NspjGo7OyeaKW2Net/4DAqBSe8U8mmuco0XKL4CrXuNFCylvTS
DKfuqQODxfaZhHMHWRksrgcbsxnhl8TQlCUjb37D0kdlGI6CMD8oN61UfYfRVKNdsYLi14zdCeOp
iVKW+N0qZpOKKOzbzuMukZFNgJ0POctC4puXdrgTN67d4/A9aVxxomZAsMsjn1TEIdRji67VaAGP
PaL12l+MB+XzL84AxpF5xNQq42w3hlrpZx2kjN5v6Kc8/zqNy1CcbifpOdW5TUHqA+G+os1mZunR
rK0lS1Okcat8AKqlV2zMDEQMRLmHjLUqzQAEFepmugK7mg/CEgKsBICWDTZBvYC3LN0EDYdYZmWh
zk/MYBnY0VHWR3x7Q7CWw7gKUQxFTirxsS08dPtr5LD7CMMy2P9Nzbvsv5N4YombLtR46BdHGqoj
5cRCN4EK08IS1sPxA6y2CjazoNgE04o5lcVwFMZWbPUlZbMbO6d3oBbfZFnDFBRtxrTbptro3VZF
cjG6w+Cis7v7MGauxYIKhxoYrJy0wNNgYf0EGwdzZU9slWn55Zeoo4FcKYRI4dS96kUNcFRXJKbo
HeKq8AC5Eb4YuPyqPwrgs0SC75iFx1LvtY41l9pdUYAXgezuvlM0Zrh00wENEnpsjlsmpLHeH+Tt
1PDUnZMJkHpuX/1dlFt1QR0oXCefqcZJan32ph9aFeyHNHYDGEEnzOe4AIO6P515PJoJatBmTd4K
gV8pxjJ+TLd/MsWMWZidXJbwNQ8CIPepGZDtMz+YdbfPQliTybolvipSudasHF8R8WYA9uKbGLUt
qvb0YuSY6DEs9mLiTZxWVu1qC83SRQVsDt5NvcU5wjjnlpqTpvIt+jAL/R9IvBG0KtKOFfzhqdr2
vNeoc19ISeYBbteaJFp5ZXK57HTs6ZI+punWOK0GQETHgtEI+IbtXS9KQ6p+QMGC9R9BSlEPLeIE
y3urpuz896j6crp+2oLPMNfsaAmf4s64ZFkduKu0OsHOJiyUgZh839NZXaBVN0YpZOfx3gQCIUs+
57S+ljtMrHSUKsf2XSJUHA0pKoSc1zu0E+uPcUsvk7UBaUqESX93qy9HUFv+METkjhaYw7FbQlY7
Z05IV4HJSjRur0DPvgRkOF+ToUb9Ziso9j2F7gncJI2SvZymJKmpyFz74LOhWDtldlWJHMoOHCpm
BbghbrF/9CtFktSeYXwlkD1qt4/M2fgLYCfUYh2yl54uukwmIuF5smaWYekdNHEbdxKzFDACnZ18
2q475BuUFZ9avBcJqR0Ftjp4jUHteFJdt2xi1rhGFX4HK4HpxmZ+mhdoqUrqnyf5mrD+b3ITi65Y
JsKaVuKKirl7FTMVSLru+FvYOopwM8juxSkGW0N9yEYqq2saiSaHkqfSlB2nOBEpPtBQ0axQuiys
ZiLxbVKhb+q+MnbojyxibetF0mbU29RRrFoNgRW/uu3rqA7mjJgXwIqxmaLK62jngWsDJbLTMzP5
6zO2G78Dppv0VvSU5MWn9lom78i3lPotgYSpuxpzTNQKGx4Trc3Z2JcLwYAu/KM5mRD0M0LlasbW
pyhRcIbkPts8g5cuL9RiAeJtvDN/sjp9XVwLxcdtMbtRyTprL8A0+xTIp1eiq5e8RPMh+CtF52uW
pRwDgPG51zZFvLPZLyRPj4ClcMW5xWSz2pvARqzqd/Vkf5wXrqyDGDBS1cSoYpQZCpOHho9h4Mnr
NMByzk+R/cfNyjqrMCKJdtC0co3iY4NKOSmXpA+ApkSsIppx6wo7MYV4Oy++PApwRiJGDbRwTMu5
vJzNmElhq4kqzgAfKuzMIWwm0hBdKuCZvZUVorTvXQ5ZK9PtCovAT/5i7g3Qq+cmZapE5V/2PX0T
8CovJT9vrgJEPrfsj2IuaJrFmjoQAUWLUbOv7o+nZjTCYyPWVbC2Jgz1wiDF4xa0BAXeISoijiiC
C7Cb6MEZfABzYyf3pWpYnQhRT2tl2XGj/I6xUXhlb4eu3TTB0jYE9OV6pM+Jy+mxMC2KEXx+k1bL
bY/D+77n/Yvw0+N5rgl29Z8YGiPZdVaS/SK/DouKYyuXejjdRfzHBFBr6Bb3t1HaCXKiqMZ0Kw4G
n+iYZA9eJi2IorGTGlhYprb9KpqZIAzt/osTolD7lvPGJcZ9lTXwk93pDKFfY0mk0tqaFPYniDND
c473EgDYbphAUmvZJoFwduPLkjiZZiT9ma6saZxWQz4FabY33rkI/UWbM1lbdFERCrpc+MI6gaHR
Y/mPQMyzsHSzLVt9s6le+MXTWD9bTjaauf0E+x8oOc3GGI4YUxE71nBN/9kJMRRau+KGuqsWGkXR
jhbiDcE9cNw8v0E+rHDrr3kHFa7VMSllKEKyybtwt8Jh/T0RC6csAigKJnKSI8R8cQE1/MRTqM5T
X7zEObztOYAcxnrgqbhMN+Cg5znG2ZhoZmW4jzM8FO1BKRd8Q6OUaBRXOUJev6QR8KHRKriaQkI1
OzatcFZMgJ+c5nQ8adpBVIUmscmCax+ba0dyK2sneXbqiQpSMc0JOxncAZ8GPRp3+ywb4XXJaKIH
ELF9FRKNheUV8VIVbbxsFRGoJ62dHq6zc2lfNkRt4dClibE4s66fowkDETyTLyFG3m0lRX/SYcBz
lXzvZekk4L+u4yJRudp1wXiRs24GBGEbKlP4kAEY5wGNaXevkWyB16MSLs4zaMMIRauNciOu+imC
Zz0bS5IjBeCGxSPYRdUMRVlMZB1P0JUeu0BVlIaeAzc7MdT/lBLT3OYaSDvD9qH+tQqQjaS7xc/6
UANNBQHM2ic7XO3+i45lTiQl6/RueWmqYnzRiFv4SmaiMJ/bcBsCO4wlzGW5k+BsnW/VQL6HqwM3
An4tVuJsTuh2GA6UH3MhVrnrXTRAVff80KcnlmvmBRDW2gl+TiUdNBoK/BhtB/9IFsNRUbvrDIIu
qiCgLNF8oHDVNUey5QEbx5/624IzTcR3YvyY9aUXVasPf9JTG4XeT82R+YVMXYbd87UUDjVZjdpC
7xsxT5dGdnGhAG6qnLpRBYKqx0AXpObfm//EeVrXt9WoMhlG4RB0vrroQ6bb3oUKxmJZ5RzscnhK
S2H9xskl/8qAxN01qK0q9afYGYaZUkwznX38zBU9QIacpmrw7dvG7WgHA8+h14WdIDf0hCxOztLF
GIjzIWVrgjBlnfV57roVd16IhGaV94EI7T9X5xldsOqNkWadYkedtQqMM4flM6F/PXGrWldL3di3
PAMzzEH4cSqag3Md57Krf6Ld3qm3FD7CrWqcrkJnlWn05xtnZE/OnPEob8mBZGbt0yiXcMIQxIob
uIV6Mc/uA+4QHpigAlk7bJ4a53pJZ1VyexC/3dB98WHizGoha5/kppfq6lg2SOfS3U45mNy0pl6g
6gxsLkw/i8j4DkmD1REmwKGNnJ44RDO7yBD2UODs7zq/j5GOZblUm0viLMvfQSL880phmaVLz4nN
teXHVgr8rlB9odTRJx5McO60Yt19//Omo4UTevWUPO/IpIPa/+IRn9iL61dy+PLmNUS+Ncm4T07c
CLXyUb950C0dD0pEAoSoifkSkzYyQkZZD4q1r0x84Z+2tA4YwYOB0KGqPInK7oAIdFIkaT7Wqbl4
VqhJ7TYdo9jDezxWNfu94RyQQdWBritGrrQv0UVpJmqkUsmBqxTQ23Fjz+7C7hNBSPxTPxXQoIhI
sJ2wDACWecOSch5iOj9UHDBooVqoDAk3vozXQwNMdnrtTXrxmPCzO+fj5Ggr25BfBMpzDvjYL3/1
+rympVYFGkP8Mdb69CmrjRSmecIrbEmC6C1m6WIw9nRtXQIVNVDZ7/pi6GVJHHl2eNMnw7XXH09r
W9cNzeYdaacCrbw1WGTG+NcdS/4CsoIBFjFJ0F11N8/OnrNkuMLos5U3GVdPghzULzuULKSN0jOX
e5HlSZTOXe6W+Sl4Y9Tey5+R5ZVy8OdLf/hHMee2KP2HelqycmjT3tUFOims7V2s2HfcvRqOcyw+
pkbFmj05cp/NYgwo1rEsIDl7xJ1hFo0KNsZOVxawMxgikqlKcxDBtVdsvdnJDBZaEUWaodlQ5Gsq
08SB/CJWBkcFRH0+/obcGinw4zijPPdg7Iz2tUwLNpbTcdggZJ1j2MQfcOEv6M9BsGZyYuB0ypaO
slHHvl65cVXiOZ+8+esCeVzYioEmzaegGx4mv9SEQ4dNhrLZMaR585J/HsofQiizLUXaFnusum6N
FWAkWQwfvS11FtZG0SwJtJDUHJDuhYI7JOcqRv7FgCnpuzj3rJWYPEEmgadduSzJ1R2pw2fOnXOV
FYC8wzDJoh+B0XLoL6HoGgdLoPMKeIq8N8pArpsBWQfLuQVLIupBbJoPKzgJ7HMnsSzihQbNbFCO
9dQlAmgu0y6s17W708nUdzvMqrZP2qm7lWd/Y8DagULSXm6ALgin6NCFi94BUhJXegITMrEFyL5P
uzTWk15Bd9SnDMUL11LXCndqYKcE2AwrLX4QKM+2oR/NQ+0sxSG2WuG8w5+0QpNjOG4h+feFae2B
6sJ15l2b/yjRqR5rv2tRocrMn0fPYwXKDc5LQx0glVSTowXipacaSYfUYdDxJQ6TZMnLSLtidpSs
XZ7fnz2f8Fa63hMLjKEVG1vI049dNy6K9+v1+Bp+0SXS7/a3vIwK7tMj8rY6/qxbEKn/jVxTuB1L
pT2hg+fcfVuCGPRs9d6oNkinvJdfTXWeuwVnRE+5OJlfjfbuWVA02ZI5ux+iPKdcDpsqhayQ/m/7
paG7E7TyfL61Lkz7FDbowWDe/fvJPXhG1Kk41t05Qww8Yx0/0ZlN8bNY1gm4j0wwKi1srgxMoWDR
F9qjh1+tA2nNJz7wwlyR2454EjK4JCcB0xNUCGtmAVdPwq4CvcQ14vP2wayWAXDhj0wsT50JnllM
okw4mv+NRpu0KpuNA+Y8dKFaZHCkNHI6FlVFBwxcxBiHr58F/s6l4VfF7ZG9Qf+bj/GVjyDLq3Cd
bosGOxWZUAxWJKCkoZ7azYORNa+gArvmvhsiPQu+YevJ1nNCbJrL+wdJBO694pCPPSLyAaORTWtx
tPOb/ks0QCwmiRmMldLQ6NRn5y04rZAu6gNd/qANNmSYjWd95ERnYubX5RZNC+DqPjm/KFHFT6t0
URFzMxEodWqRP+UJZSd0jxD1/oWXsVzEXwGkGqJs/5qd5LJree25qc0+z+YK014SsTHV73XHkqfY
c64JRJIrCv8U3oiuWedFxaAAhFgOknpewdN8IcHd2YxNfurGKRDXD/tCCTXFGBRYZSPAMsWAejFv
Sl4EqcaFhPS6ujgT4yVT4qrm2QGrSkx7k4CEwqxEoel58646l1QWmg1el9ffd81jkqtuA47sfHAq
XYpXbIMhnom+Z07pJlYPbeJlnVKB/6F6Cu1EkVZIBGRr6JI8gyC5Zu4aR1dfjxW04QLZDjn8Uv4E
EJLNkL5JQvwKgsGiz/t86OB9GcnbL5QsXLAXaorS4Yq93F/6T7gXi+pmm0Xr7AVvyCR/DhlyS4SX
vco5mNGTev8RBgo3eFA8X6CQGpEM6zaPXUcv3CsLzwrbPW81pCJJhXeQmY299EzEc0yXY7AmbmpP
T4PDy5mm+5f2CRnJlCplQcPbx8fUrCURpKEK7NAQXWpz4Dja95V5WNGWztnSxiMjNKirJWvA4wJI
CL/nZxrA5C4nxPlpZ6eL5pAKrZSYPDGrgSkmHaKH0hWOZqLciySrheFLT+61JZI4MsPGL7iAMC0w
binAPes7qSvfOq9ixMIi8xTI3H8Y/jhlJrfmSNDEc6mLmLt3ImYHA1zjF/egzNYoQCu+Vl1ljyMM
3wOH3y6lnUuZJoQnBfoBaVGOUmAsJnEefkbqwG5BuwOwwyMQ7h6BHKPN318Lf1dYQKDte4928Jl1
PBkDj4Gy55zQJP8A4jX71MeY5+HecYBa7M2GdWq/N/+b6fd5rAOEsAqPXNADjD+u0yztDMWZleYv
YUgS8/ZQnmSLBSdNxbZDFVw4Qs7BmXBUNSbtOiz6NvHTP9W7FTdAXlseUqutXfokrCP7FgTGVKHc
T7HmeFXdz3Y4buXBE7rQ88ZBcpQ++nbH6YzYVavLx+Yc3JDZcmUXHZAGT2eeySFspBKfbxYpfI/c
hGuTeH7xetrtwH5tV1GIBop8BzsReA88zUp8FXAiAdNLC15IPhnTc/RzR3CqoutkPKSR4jdZIdTu
oY5b0/jpe2lBxDZDdERmYPK5geNN6riB/f2x2k35PlaHcBxdxaGqMUrCuITwIit71C8bnozIiisf
vF3RygUIYg39AMQe7wJIP326vozm1qcyp4CReaK+8rmE0DYwnG1NTuHgz3GggCeAveWt3NwmXFyF
ByQLKemJjcWy/6vzoXoHHASID6AV98Tv2xyFWBRgs141O9h4NcvxvWptj4Ghcv/wf3caTjXpAbf1
rYMfr16yMuu+h5K3ldb9iZj2j+n2HuMOkNGjfdfxRKmAjf2p5az1O9yFseGOWnmN/E11jSB3r2Kg
Izd098KQEeWljyQeQY59NrroIGCOerlKqH4IAgK0/MaYIM6JgzCz9NcWuplugMuzkb0hVF48m04L
NycssdoK3JHn71P49T/yGeDgzQND0V/+boCyq3k014sEVrv3sDSgmcaBgNDFDB7C9kz2Ym6WzKsi
fUGgDaTKSTAEuT0gh74gSs9IzCXyNUBQcIbUtgVrMeHSpqbFwzPGQMPhcjobbowEOgIDTrU5kFOf
NLap1NwkgKPqzvhbg9Cp2euDavVLRMl565Gw9kvHVH/L/Z5AQUn8vEUyY6P8AgRsofBPdqwxTs1b
/jnJsDZaC6GXORInnT9WSxJ7Ckvxh3tlkcGdjUX3yihfjqu/BZmal24LE0JVoZqpZ6kGxAgD6RgR
dPva+NfY9wIFo8W9PYtOp+2MP5ctXfuDabMbT6i4ppU4UUMP+JyA0pkmiaeJuDzsE1F/iMZzHZ2M
7sXXe+KIQFBeoyLFKp3cNWbsDFVsHKOQokS+Kshtrowf6EDTnEshhsR/WYiBZt9DGsrcWwhMTAyO
sCxadQtkgLarmIIhMXcFbf1QUdVF3XmA+qnnvlQgLCXU3VugSh2SsYgoH3ZB2QXuqQI8RC/yJ6ru
Org8u67yp5wsjxXZ5dL6JAbTOSbbOfgA29EDl64vxx+UtPEw2cCejQcaYEiJnEmkekpzea4zVHm/
yeA50k5EAXJTX5nGG244XN5dWBv/fBSiY8U2dSkrQ6NiZA+qFRqOcxeMkfuoqGTt+ALD8SPNfBTz
c20AVby7thmgjeCx+N6pMjCKP7jW+vJC6kTkbt7R1FLELY+q6AAnkWY+29yvQ6jmHWXu4HcIu8JS
nff1UD9Tz1YVELBdHfnmK6FnDjQr9yIafi7G+Vxsw2C0wiKueOjUydu2xsBOaNCga63xyYOQcuUG
1VQcy5WH07oAyLvTggwUA2LXbMJV88C2kTb8dbLIztdH1kauVkWwT2o+3L1z30uigiQhVTxsLbXV
2L1lRJwjjseD3w1Qt9YjuMRt1S31CqAh/UZfcOJ8LnmUQUDPLAqtybLypPOvR/B8Anfj58A3npiA
q3XnKTe/qwmpxQRw8pxz257psBQw/ipkqiNSsxTHYxJucWBlJG7r6k9Pa29A0LRG/R6VEjG96w/j
yQkdulI33cnxUeQFSABS89A4y11x8NgRmzmiWw1+SqG9uSeTA8i+sCQOc4sJjOQwF7vH1q7FDkjM
kZr2KTeerlkKJsNrouFO62rIisI80/tQxyqdnfLd3hhfdPNuUtlb9c801C8uTu3+ovfQDYZLGRJU
HkmT2iKN2miUSiOW1a42hqBcLC2XvzEmFkN09oT/OIloTjOdaTU4QQII34NRdrmOe/jVwg2cadi9
CaQN5pIgqq6khCsKDpB/mE6OKkz9MN7mAMJLZpNmnPQnwM0QIys3se9I0mUAADxml9MCPyOPn3/I
dY3SXDnYQNybriCcmjOHc6SF2d5FImdMeMfakBOeyqmkor03R1u2CexM2tEH1NqmFBu6rL1SPJ5H
TsY4+pMG46YR6x+TtYrci/DbMfaSJPFpdNL7DHsmMMtI38/9x4BF1KRYLm+DEf9bzX3IC3Rf6Jq0
ozPDkgh9H+E7bs6Bvt/p+2JbLwkOK3cylzHwo8c5zf7iPlWMoyPssDVIbCGmtWJb3SCy7a3rWRHh
Oi9FbmLpxoR1sLI0UHMA1YOxAIvqq3Gkwbg9fJGtPYDIk0wU/M4GLPKU3Khy3NFVydq7jB3viHPG
8CKvrjdIkxgeTwR6KftjmZS9I9egVOyOWNV7uCkSqCG1WR4VE/MEAO4YmmOErMiXsrVPRHHK10dB
jrKHgI8OS57lNT5t4vpcskGle+xkuMB9QAtVrhU86ou/vyNq2c1gFEpqcCc53goM1xeyoIm0PUSA
YcVIndUOEELvFFp83JD2wJtE3xXCJbWOfgWvgdazcoRv4mjqbd4vYY8MWIV9h1dWsjCtAcgfTHNg
hR9w31NLDJFW4jLKr38zxStrJE15zqlqNhc3J9toVB9tiL0fJKtK/bhaRkC4zrdEofvusHaS4CJn
U0LyS7eOKBqX2PDUtBxrR0UCVsb8MEltRz2v8gqRaEqg+sypWfpguEYxkTCDoG1mQPnVEb/iINpk
Oukk1btV3rUIB1ZIkweFg8yxup5uiYbQMeQRIe9wQiOa+UMBZmTU1a6HOWtN7hHbNIZR4YmN1wkJ
lfSB5ySokPjGFPJ6BzOUt0fev9j+z3Q172AIiVXaGLm8Tf/MNk/1YwcuRKcBufjdil1/WK2q6r7J
Mdb1MslT7vxtYvlpt2Ahvk5r6dVac9L8DSRwlA641ndOv6o+iQQpN5wwCNDRlJt7A1IYP6GOa+ZX
dYAXQiI9HLsaT9a9ZwV/ob1mu/3srXAX/Zm9H+nRjMvQ+TXQtRaQWkywrR5qBBpFyiDChyvkQXSu
qxj/KXKBsDBTQp5JA5La57HVJtZdE0ijN+PYexqeV+UJ7zd2H+b37stbbV+i3nOucidQUz5OzH5j
DMlrA/VAInycTHl4zIpastSBadh5DmyXz/5/xnRKat7q80CH5/pX7IEsg78vH3/3pyRCRXamcB32
NhHiJCYX7kYhucU2hrltUaEbxtLu+ywYXNxhI0lxIpMbcexVsNi/c6CBKFBmr5LEdEEfQsbBuAEr
dEfiryPPtfLCMNBsupVyQ8caKQRbXyezeecgpQpIEtzWxXYBTaUozRvQUXH3xdbTF4pf4qERt+rf
IZFTtHE7nNciFLsGdFQf86SPrXTXN+OwSWus4yZieK9ojfXY+3JTQAgmZtEH2hLrInsnI/++oBMu
ohX+PH4B7d8/fwwXjKP+vYVO+06selZeDtbcQnioi9ywgMNEitZxpQFcitvdYWdMaeDOuqRJgSKz
fJvp+M9ytP5Z3g+2fK72sVmMI8buKs6fP91KhNbrsq9yOUR6rmkgEEuLkE0+8U96GsxCheQVa5nl
uKm1jJ3MX6J0z6ZFCRJMC3ae/3me+z7EeYndOvEfxg8u4Ad+Sf7Rkio5hV5+qGkPEQ/2QP+nkcdk
0qiX52lbJL/pnGSud18KbiuYukrj4skxvrVteuTYQcKic/li6mxjRZ/jdSv1//+kHraQ+MbCUC0I
MaUOr7pbzOghqDuxdN4TW4RZq3O3HSWjXxQtewb42VvQyqZ/QbKhlHdlJrDvPN4sjgpDkCoIOKZS
4Ciau9+Rl0z+ydAsODcpiNBYnq989x1EQjOBwUk0CYVTe+5y0KE5kRFOFUWzulQtkL2NEg+SUPsw
qEtTTfOyPtZQbPWcuV9sPy/UgFP+HJnUuLzZlpIfx26Xfg/01bqho/sJiyloFrJknwsVNm7ufJIr
h1+SUimAA2FempxVVRCcntyGp6MqUAPMVwNyQUWx9c/aP6JZzXk3p9vRixHaWaYkjNpDGCknsNI7
G8eJQIKvIBwvcHJcvmYX+TMPATsKWJXmfYqIsvFtS7lrVAlIVYwzgLpGkpjHBNvGuvi3lu/UwbcO
rivT5PBaM2IQKS7XNTKCr7wlOkR26/9pJ8mQJqvDZMdWasEjF44MsdCytfKjAdr02xcsDEPd5xQD
hZbwAIIVXl1DGs1tS/S9VWiWY1aXwynAdCRVtA82e5vFMeaWHtpPswk4gQ0NlNdFd8kHDKFHgSl6
udeoH9kZ0Brytb9isCdbhgYHIWxsQWQumZ6b1t5Q7nyneqqPZ5979UPsSgSRhuMz++H8lJ814xzb
zT3jRdUbNSFUr5Q5ZnkU7e13EzMLVQbFWLazPOVXQkTUriEqUIpRSfcTY4kq37jjmN0JooiC1KW7
ArJT0tmw9Cggx3zbgRprDn+47uRgZQP3FtC3zEcpydYRJ81zR8fT+uTsPkqcHeS3egX+3ajEdjSK
Gbkxa32fQIWszC1RtOWIdpBS4IPpdhINg1ul70/k+CVaJJwVZ/RVnmJ/EQIH2Ipc1mDCH3RPvbEa
VsDulomD0TwbTt2pmzH0mHjMDCrrqvjhk8YKVjDhBueaezeH0BnGYtOqvIB2sj1EXclv8z56aZHe
gqbCdOy2Nie1FFdSB93FFM6MuaVealiUI/Y867siWeSYs9x2+LxumiHoNGI0nOVM73LmRQnkSEFz
hApLgRP8RJkVtyZjXkT6RTpgyDtd02l+d4r5KQ53SrIpAivgREhJpCsOyQ0JQ7GZZoaDbuVqdtVU
k0861FT3wLEPukduLVUQczCND0YrtgAJht30pgZRMgF5oay9w0wpwIoEIETkSYYpeK0pVNt048gG
HeKDAAwpTGNi80V8KkqBkRR+reXLOfOqx/2L3dGldzoR8Ay3c0j0T6VzhvQzubMA6oeg/bsAIL44
635fb8r2WKp2y/MbY2QaI1Dcxm0cuit913Fc2vBQ3WCaatd7kSyO/CjgK05q4APjpef3a0rguUq/
MHctLbPfdrY2XTMh8rnEFYQrQ4/l5OaKjA87AfbIz8LQHArokyMKomERTaOc1NfGNEoBeoC79dDB
v3jx+KpDYpgk5gTMAWF4tMZllFcBYTqRRb3dl4pGCOb3GNhgnKanNRi7s8zqR6eNqdo9QPGiJQRX
wQ0ahCHqA9f6BDHhVNL7PTTmKF/rc/ozB5xIdpeoNKZi8kl/vV+oiMTHzftqy4JBmbG0XMIrzqy0
jYzQDVd8eD5UwcGew3yQ0T5TzU4PxSpDKJmjV+He2LALJGx2JgKfZ2XSyeT5SuNUQnML8H94ylmJ
jwkhNzOewWWbe8AymE4gKjwnErJCfA9RES3NzlQqV6nml/Hn6M5BlvjMIy7PzJApa+suNLNHJ2hF
9LuU4yUX5j2qoRfJWDsy+DGYNSYYDAPaZoqg1VI1cAPiwFUN0xFreNQjJY+iAwZHNfy7mBQAUFym
HJRSBxdrUNIyvZdF4m89c85co5UgrjAK7hZCkXefNn6/eNugm2iVd5oVBCmxfaj9GFBwQpkrhwJG
NZC1mjRMq9Y8+Q6/0urs0kyx0V6UTUd9Q5OPHVxvLVPnYjVk3VDILkAz9jlU0ZtrgG/luR5LArLy
iftrMuzCmpa/8clk7IPHLDsa0gDIEhu8PvHoZNAE/fHC8jory1B7YzgjMFxnI3GCvgpkc6lOl5gl
6ivJKRW48njwLfStjs/1sDqpG2y4hs3P5cEUhsJnFshbpgsfncSuFDnYyG/FVWXqZc9qw+mO8yYn
Bg2OJa1989Y4kCLn/VkA4m3tuLWs+Y43vuKP68cMOlOzYXjrdhb9lRl0SuqNPilmKWcmm9rcFiLh
oD29GjLJ0WskUFrgv4Yrn/c8hYFSloyksqyqYm6IMbNDlJIz60NsxNWoAFQAtSvxcMCkIpoFchxM
s2QPDsCKMdxudXXlU3PiNC9P/fomdvG8tv9i2GKCxJzH5YEPd2VLJ/f2W8c6QhFxGw++dgY1cQ17
0FPziI6qHqzfjLGDRmdLNCQJifLpXaoGvfqlTvhd4/lOGzJf7YiAiSoUvIpaiW04M3oIseF3T47J
LKKlx5lU3XUaSngbseLzcP4/YP1T3p2bkFk4Bykw1CaZnZKh5cMjTGM+w4hgGMhRH0CtCdPVEIWD
VUNQU+hWggxlg24ACH4LuJElFws8tryv0Sloy1cn7Q5CkFBR0XY7dykdjqOpCqBRIIfqJ5dCcdiv
8rLozSx9UaT+TvAGxxeYGqcSmGgMSt6Ql4TZzB/KroNKiMmlEosxNXvcVW93vZcEKjTm28LqqjfV
pdnQAY/G6Ub7kn7kromR5N86RBr7g+FlDhv7ZYtJupsms/+4/h64uGtWWBgmLP3GQj3+gWIs+myK
/QBYi994uyKtcDWjIqIL+cyVvWZwep08Nb+RU4au64HXBv0aez4gjszBa5HpKTk4LBmcyN/TcW3n
tLGeHxDwH18wmLZN5Y5NfltmSJxFisJQJYMDycUJYs8VKzxXHvizMa7WAZnV9I3GnG36SFfFEJ8I
PAHqKTLDiEJ/I5FQqvOZ9SJBzp5DxpcmQlXvm9nMOk9M4KXdzVljGs2aAJ3bIPsVGedf9Ulw9Iw/
LozH0IIr6sxn9Gv5iCIVevLoyOXVz6M+84SmHfDB+2x3bZ8DAS89Zg0zsfPbBty4MR4n2N0ohNt5
BF21TgmaHsbCaVAiszDacoxUuECEteUzOrmXBQ8Cs/X0Eac1jYGSPDeVVyr9QxFOYMrp4GOPCC3L
siNDaN3/W+dLPVFodRWVAvEWNgW1CGqb+30nU63+3szsbjQkGp1dGcg6lUajg0wVEzZBCKitQ2+l
7lWkWzgVvvDEMMhDfYoosVGn679czMdOB4dSK9FDWInvsIGwvzN6OR3iMsCO5uhp/s7ODIMxuitq
yBJjcnJhqGT5oGXQSisX5MoBHDCBgIPjEudL1Ex0tSC0ImwmKUgX6uLkJePNNcL3oBkY6alBV3TD
VRPxvYu83alwC9Fad2ey2JVPI2HYdUxiUm/8YDeObjLBGBuEsv9Flb/gkZYu2hBFZx0RODMLX/7d
We2CYyHv4sWxW98fD3u4PpsSmCeinYeRTUiQBjm1Kkj2g1KJjyVcCWEDo/Ub/EWb/4zyLbiExec0
TS4fKUy/CDkZfepAr83pqUt2b/EgUINNwq+XurJdhXCpxIeiAdKsaV+IGQDbOq+GSPX/VQ8rJTBm
9QxQBf8AcQGdiZGXyhosdbK5cy9hFtDIc985hfSGXNAoNZ91kxN4JoyvD6g5KBuJMmFFQ9XIkQqk
n608hvFXadHuf7puZGAEBd0zyinVdbOXIbelmnEa+gjVfxzy2Upb6m2GCkIkAwYq/ghdmO9avSN3
MSpP4Tu0traEG/3aUVAD8KUXlyUquE5kD13LyRC//OTHmhW0MqOMfWL31jXsDU1aN0QUd66z5Mms
pvMVYYO2yuVhtNC0uPSL1ztpEuorGOZQtH7XO1SITljkq/Eammfnwxaa3MPvP9XHM8jY6+iUXQzh
zCvyGIPNb3/mc28U70EPS6lpoOpnxkxohNd2crFkaEMfSR5IxO5/PsMZRToNgHeShJUSxbzI44fA
cOMsmYlU4SrBTTpX9bbVRJOh62ID+zhC3wUW2Z8D3zY9DbhA1ii5fz5uiS/pk5RDRhZuM8RB6MV7
fS5MDeF1ygk7lBVZZQv7vY9Y/eaQObS+N/hT2/ft4iSVQ2LH9ahNSw5AVDUqf093I9o6YgkOTuqs
K8LSRlL69jqDIZyHMT2+sunLsGS9LjOZSq+nHB7tGAG5Mt9j76lI3HDrDPYFA3ckod4MATTvllSj
trCdWaI7OvJZdc+I5abn4DATNnG8Y5PrTiOQTeqB2cEE8u/O0LL1l3kWxtV0KSo2ou4IK5bOFTLF
+caU8hKrvswjrqhSwzQDb0LBhm12RYbqdMDF+uqJwbFvbeGjw4AuREVBg2uVfBJRXIjebHtK6Znc
ypCSLej2222gyCYcZzunBWmGNc9Qcn+3b614ybXg+djo5xLu1+e46sIgKo5jTxzEZ8HcLlclElev
txQvjpeC+heQQGPLHjiyXMIo4+9Dj/ZzQatpGxws4Io1HgeGlbwNBo09C8kLVKZ9zGKior65iU8c
6Ql6ydZBj1TctVFhkU44ZU2w2DiegfULOf4fxe+LeXr7LO5mLjAT95F11s3KdXO2kAR14wNeoZu4
Tca6FAzDFFNbABEXNWhe1ARXZzWbSl46By3C3OwZqCEvow6nvyU55N91az/0s5alYwRsOvqLURGa
1F/B4KvXx2nVZG29Wvrwh+WLZOkpJE+2H289l+QWQuCcBYkyLUkxSPEjX1ap/fciX/bCoLjUf1zF
heHo3piQWNyopKhZaCwsLR8l+WjLCLEQOvehVmD6mks7lM280MklebnsdryN9+qjaWq41WtungWO
1pamI5qe7BZKddRt8KLDfSjt+b4FlN54N/YIixjMMBCZG6/Ii7Qvf/e4hvARqA2iDVatW5h9SKOS
p7f9/Mu+OIqO8nqlVeu62d217JTJTEs3iXINOxSEU6mhtFbD8+YshTrYNhiNUh2Pp0gv+52hVi18
qUcZdoPyJwdneCJK8C6PIvLlMmRfjXidY2ZCTfzoO14uDw44NQYOT7fODFMVSfcV7poFQ9bgsIDa
6aZDQvH6ebxjeZjeoC6GRLgiiz/OOLrkwrBqGQ5uGNdEnsKkXKuol/FxBrLTe6tIn+1o5bFX8uwL
ogEaZFs+V97SH4ASQpmRFMGQ+674CgT5eTwQWf6OByz3+9y0DzepWVHGCYLmOIbP2SG+4xfKPs5W
0bpnFU9DeChokYGSV2UuUpERtmwi3mNS/KB+k51P6/ZTaCDvp8OdGKwOXX6jZbhViUrJzo+axduS
uDNLUoC0TV/j1JMe9/iMX2ibkrloVUZ3Ia8Sz0WMrXqHsUg/ZML0VKrNOWiVAOOApvSlmgmXsLkE
VUMBHo6XEboYlYDvUwPLkBf+5w5kMtMW4wZ9LbaCmxghh46ZQkg4Vl81Psvop5h1Jin51LDhMMaZ
P7oJ3n03TN493HuXmsNMCCqj7cX0DqXhoYgpWT6taFF0r59jTqyr36kUiD1txsVi/bNMDjBx2R8/
R5gKHJUJ21amaeBqFpVxV8dUa23n4WXIYyBxYirh5j3rrU8PKHyBkO/RZmxxqNt81o+Hp127wQJm
gGu1fAa5Se52Da3SDDv/ndPoBnTcpActsasJ1RCWh+fPiQikKYNTerdcLvzeFYPFkzbX+idikRLY
Q0CFb3fTSXOh9LYnqxz+twGMEwfHtozcvWpKRYltKBveGBsJU3YMnQ7foYfZBOi+Nine5RHQml1j
qC9iek0chFfCxzUV9a1N0dnV+L7GvlfIdqzKPCpR0/gRdp7OkG9Xn35SBVy8SFUwhnOvDtkfbY9x
PG3lXpXdKXWmopntONKdX2JG6mNJqcf9EBFxJzuO4KRPMLIb4n1eUNLPvGje/737gIbNm6POQZ28
WZ1D8gVe+HQzbSGi1Jz8EFnpnoiJI/rATd2swOO03fM3zR8nRUey/DSWaaknMh4I8Dhuw6M1FtID
Di6K+81fsei+tfhsJvMzZwlYJ1tLnno/N0o6HYLfckJQnBNToS+PJAuOTlTLVeS+eVQEB4x2asda
2hbCJYIXzrs2wrMvwV4w7q4nxBGSSKVqIAj8tXZ9EVxIw0YFNqY0LfJqhzSoiXBwv+hleWXAPLIR
QQWWtJL3p9cHEN6pvAUW1KQlO/Q9P+81cd4G/uJc2N/vrzNgMGh7+LrmI1y/TtreHjqlp7ETSPgK
Kdx1khll1BDagiU88xwn1rTWJNdztwAtDj8cIcZY7Kr8U0VCGfGNAAbwGsO73gCYU0YpOcb9zk5b
T2+iNIoKMwdijOR5SWu7cSUbtiKtXz6vnzsAUyC4NudkCz10abZU4dz/cu3tjppB7Yh9cmzY4MY8
0xQ+pgDD8dhKVkMMrPYFf6+UHhcadZlXBAAHokW8syiziMrlwXLFArmiNvpR4G5Wu2otEQMRKSV4
e1DAneVJukolnX/BciiMkE5AuMyzkhprJNJCbwaboW9lBjdZwVTH1pJR8lnKLaxR0GNvhnXrxlzO
ehnFsbL1PpyZkrogrSkvWTL4A2hivNBZkLGAAj+fAZK27hMwSWUb0jJMv6rvPjUx64XHCHkKm/Td
vL/043pq7sWL1KVhVlliEqfo6kT3z30u9uwIzj9/pQuMPF8kHuB8XNhXRhwK5++viL3/neB/52Uw
RhAzrVUEcVgjnIiZ2RxPWpTZ94/0ggp89Ckm0i1BniaE4/nC/9PvIZ6sYLfo590Vzm67+CXVucaE
QHs3wLSGAd7GQ1q82CJPWuufkdZgTQSxCsctIgBxMlKAjukbCNKTxYD2m+Nn5GLjeTkRhjZVqSWl
smkJhHlwxVWhMK7UnKx1nX2IgKgzNGh1EqHRA8stzHJ2yV2I/VPaB8CE38hlSUog8MGgJ/aSktXD
6Cdp/gJ+caSOY3hkEOXd/S1p3WA9rtI1O91nI4m+TSBnilEj7Yqstgk5YnfYsZg8I4oHT5khPiOS
tX63HUGfvOdGG+DKlq3FWO/q5kkhTsh1AJ58UgNPH5Q0V8GpvC9kqP/NjjYaLxXa7y1peBnYMW4E
+JTsx1GrM7QonDOoNXaiAgEBJesC87MvvqZa5GwoJpShFQ2hQLbccI9zoZw6lEf5eYQfaEvFP1fU
3bb+x22ufTVutpL4gdxsiTHG8oQzEP3/S5AktfNKoSDYBBSRq1RZzyW+1F/Xdl3tH+7TIJyafFlo
vDV685WoynFu0WWefCUk+u4kW5+dTYtNRwxZWFbm4jiwgucVy/HYiXMnYF2zT/fRozkqTp4cdczN
v4Jiv2wKGTdRLvt294AiqTMvXFHN5fHibarC4SzjNNjG5ErRe47jEJD8+mgcUHnR5gB682c1kd3N
9yj9bKqhtN6maFGhV7tklKPWEAtadTnXsNpBPz0LEu1RI0EZB6vRI0zXggkiq3Pju9Mhp+1Bb4wK
FKq78u6t+KMq8DqmwKC9n0pUh94dC42qOF931gaEy3nAxsmm1XNiolhiV74RwycTKKOjI3qAhuMB
2UmnWc4y/EKGumeShtAHKtlUwPR9XUuDdKA99ckeD79rSFVJKu5aD27WTbfZ7uxMQhYuIab4OaTV
xx/qScLdE4SaoTFMUKtutB9bNe66hgfOCVdrvaVLjle1P8MtjLVBYJ41H6Q0FMa/JZtYW/2a7S1O
wx8uYkv69UwM8SG6N0QxQBxxuhdygd78MGCCitQek3HCiuXtq4dv1bxUBfS8Vci2Kj9cc/FTdx0D
23Yu+Ut5qTyK0QT8n8o96DVILordqgwTRulTnhTd+FOxMa/DC9uBn3wlYBS0xGZISanGLnWLKIFr
E6d4zqIlORKCCwTqs4sci7BSkLt9a10tsYm2ikkV5ORNjqxu8lgyKCaH2MJY5kyAo/IP6SJabYCC
YSNv8aNlFXMIN0wQa1i240L4iLlsNKqYg67ltoxjFUUIPbGGV8GBRLkEWA6XbaCx5sdRr4RlyAzC
RkOZHUq0FV1mfcYdls508W1LQPBNPP8oU+1ENZTPrdiLldDIYPBgrbngK0sVI8PDmNlUD3p7K93L
ASgu3R59E87PWHrMVT6VXoKnkKPiAcOS0pl2H0mLk07bsGXnlnS98+JlNpIdgudppKbr3IPH8zIC
w5DX7D3xLffKO4AV9im+7m7vH2+eIbhjxyS9/d5ogvUxXG6FejaU71TGvhGyYQ1XarxhHNR/W9yd
IMZlmqf0kUpPgB5L+G/RArbl4RBbfrbQy4iz/XTvmcYJOXrc8nP0gQGvq1dzP+3TigfvmWC0OM2/
Tw8dQYC85Sr+axVCsYE0s3dV5qM/6ovHL4NaFnElAN7FYAUYQFdncUBawAqtDUA9t7+5o8G+tg6j
NS8s/0UXTbSqC5bWskJDpNSQsXzJGFUeTnUJkRoNSGyMolN9r7SFbmJcDZXNODt+dKxCOkmxBPBm
bvXwkGnXQccf3zuV9XwTVoYTvmi916dBf4PgjIqfvCEyoUttFGiOysJRLOiFDnjKAXKfpwVNiuj9
d4Kx3Uo0xbdxc9XfumjbV513O89dEJSOiR4DRPu7d7PtHnhd/2eIzsWX7QxGRnklu+xA/urNL6Y2
qdWM77Jr7U8RWjcladFTQ0ScQ/Yuu4H72d29faN4F8c74rAWHiy6dLPQxg006ULj6XNYOSf/0Jis
JZa6Qdl8rKIxg3YudIwsv4jWihdYRMtzvEmda/cueesx+MYRMnLaBPj1mWQgwXuFa+YbyyN0XUr+
15/W7j7I6TbP4Iokhi7PJ8KX5GHl0hvtQHPBqZbrFDxy43CIc9XU8Ag6X0Y1Dc02utjodiG7lfN4
unuaQKLuWcE/ySCWECnGYZ/9FwfMKdfZs7Tuexnf9XLlNvengx6cpp7sN+HRgDN2E1A+CmCC0jdx
qT5+re4GE9DSF/e2TYS0Kg7OktVUFkG+1meFTarCTRivLSLLNBUAmBDhjnrgpom25B9r1592YhB+
GyE37ZxNxjtYWG3kcpiNFb8N+VLZZThFMr6fZqsC6AOtpBI1r3MZJJrF0xj//tbUc/dRl42rLotB
NXJC7krOHTqW03f8+/eEZf6n20n3KTw1BMVYrV7aqsLHUtN6Jhdwa8mstjpm62+bnGxkkyRGHeYe
TX7NQfy3MudvcJOK/LbUPX2HWvCueR7txpFQ/ZueocPsN+ZBiivDd9TI6WIQmTbGz6rpnRvsRxZX
lJZVeeUdZqEmRn/td7giSnqH4BFo6prEFA0hinAtmvTBJDYvfmSM5O0OlrP/FVFRQtAWPCNCRgAX
nZ52ldyWRXQ3SXKJBsENzQAwzrGoqlLWxfgbJBMcPeeLucrPYCcP6BrhrsfxfQyhv1ygn8TV+Rky
8yanKmlN0JwEsT4Lu5AmLR7TSeZ7TPIS6di3HZuNwzn8gRN8BOH9HjLvNsGDz6aAgBdUA7hZ+Lmt
YdkH/t3SY2k49MFpl7+jp9P2c7qVnJMFFEFDs1vax6IJ0ivIBHj3PX3+iTGbPACGOfXxP2+d4EP9
5aqzhQSSk/mABSMF9lci7JsEHRStEEH+imQBLjylPaS/0QN3yBBNbuOvFHjDlUtUdc+16yj/Efxk
WbyrVGzF2z1ouLIx6RkPMXiC0zCXQWrpYQb42TDcXFjZmjJUdl5JYdHx87MZn7tPK330sliGG4G2
rosXAMimrB2vCaWiPjKGuZbsYC7hTOpQ36lOsJxB2Ym8bThswbQhlqQju61xZsne5D6zxpqcKjVL
2m9SWVQqYggdiTStgny0Mtz/+GGoRPiizt6VDLRqWyK98ru0oPQBd9KoHvhr71iqexPlynS+bvq7
RfaLUL9Qq8Rt2sDAN70JBf5vbIdSW7wYPrqy3cercz6rpjBarOn4g+B5nqYYCxeinVbZI+e3oKxV
RaoAtdBlim4P3l0AP2A3nMIfmLvb/0WU1tO1IhTgV6g7BngRohhYTipnUgckz/D+iEEIosUNtgzH
ZzfYkXUEtgohs/lfQTbmZA2KQH0huTlPAyDNTh+/A3dtNnHW8elJjRrhUHdgtXD+yIXs61z0/Eqm
m8oLITgJfQ5drAGR9U/+xopuf+zmVhh536kkZDIigR5Z996PY46acUpfqS6nKEwRyQEOXWBRUqtr
s12BWZGkz1U26JvRkXm40HdO5q42r7uzOl0xD7YoD4bbbO6WeuliIFB0djxNpr2L8MzaM+eLwDlj
cffVYlK/S3WfKgFTbRyTxrWKGVrtDsP/zA3amj+nfjvT7wk0QSOEU35+/DpiCsaHhCTi449rWXlq
8ZB+x9KWxRCaeG1sHekrPt7o+el6tEzG+vGXl0oqtH2mzc6X96Vr/Un+mxJ+GRuP+uxBSFQcCsfF
VSUMd45AWwylQL7dz4sZd1UhVjn7qoRt5uZ7kTyZrSzVpnFTEEt+HHgh7q8zhXi1o+P+fhGq8yuV
1QmAwOwKJPTmmcTUDGz1ZNu8X/XGN+jFsLXRm1ztd95ofK3LUiT1hSiuS3bJjSDhU09TFbeMrcGZ
K3hgYcMz5yrbNOovX44LS7SeUpgdl2nqFyzgexP7A+2T8BQAyRgbgscxu60pDqQ9HX3asws5t3KI
eYbMRWOCr5/y4GKOTNOkUAWA91MNzput2bLrWFmvohXis/DhUAzHHRQkcBwg2tmqzwfi+6ahzByv
Alc9Yr2O9Jg/98Jg4HUNkkMZ8Gt2AI9yz1bQjLhxGXKCQBhR//YFN4PfB1OOnKIJahqLx0KbUTmy
4PwgBAJ5irwi0MOkg+sTpECgli/BrGZD8nC+q3DmO/LG39b2iYnGzQ4QekMHWYJgPc4qbwvA/Hm9
63GkCrHhxvj4zOv3gH8pndRl1UPsHPtj41BxBUam/TjhbbXUkwNVMTrzb8Zf9cHetvcywgruZ8ch
Ca3TWskzXU/t0GLDx7zaGRUbF2awkf6CbjmWhOl4orWprZa93SVkcvBoUpz8t8Vr647YoG58OUoK
LndupWtyFG6TaGW6xeli+VA2WsXQZ9euFGRh6iI9K55Avqbkz2oaTY7niHmJ/B8foIFYuXMxx6x+
gz4vWuHEd8iSweM8ZRJQugdkLbBUOpsiYjuszkxus/llplSupM8jt4bJpfww1trp3DTBavl8YWlM
JJrkdCWmJpEcwCuZywGd+rzn5YO6z4/EBSQCgqiRxdajFw48X3A9Bo96hYpP+kMrEZQvm7mRt3Ml
vg9bP1W9UWFATR7n9KOwLvRLNE116wOsChMEspnvBS7yQwkDRiXmWSpVEOX4FJguxCGIfXz/SPFn
AoTT+6ZBz0jouRLcRCvgJOw/3OP85Umdyzyid3ijxoL5QSPxEy/bFixMcN6fE9mre2clbmKMmKZY
lwFPyJlzO4F56EAQa2RZrxlTMOJidEoRlDXety3r9Bn7NAkDvKYtOfrVDz4OBsLIZhLE/tvVHpmi
Xu3sJB8rZYxWN8bFXzjL2WaGhXuJwvLwe7uA4N5rcVWr8mFziahEOoya2iK9LxTp5gcCGagq8dSn
Tkglo03/woCpTM4sHf+lRQ+ihZlCw5ZzH3ywxFBHRuyb3FltMmFAd6uWTa5LWxu1SGELLnVbgKIM
TmPx9n7lQuELkltr+abWQj0i6u3qZpFeLfzPPj+gJakJbBPcBTCr6Igp2KwmSBfkaRUaDmq4Y8WI
kxrZcOnqGldiaF4UVDHvPDAoHVM9eNdBdczXCDKPWFxwUr55c/bPiMFAOYQOhGluQIRtM9wNUTRI
JrO7T/5pq94pKPixK+f76raYnwsQHA6ePUmUA7ZaK73VwLQrrsNZQwIIWRVwI2+5XVcWhezW056X
nMTPrnVdY1SOribLIMfVH51ctEwjKXx5AwUPoNW8mKYTIGQAZPLBXjL4ISnRMIxR1y7NWdEdsAM8
tPMlLcCxdCS7OIBQZWseUSD3A9x/xASg7G9MguydxG2MPTYfMi+mMcszQA++GLRnHjrJ1GW1tz4t
FlkfVhk5KRLoOk+50PmBXj8Y9tFFNI1uEkyyI6HZRkqxZlAcFEglsmYUcyulcjJ4NN7d0st4O9bd
Ue0c/WiaT3PuvO26H2A1mgnE1SSFM4vtOVAA1/nJ2kWA46af59Z0zOSFxtQ7GSmPPrAHq8dSqgPz
79uR0iJTf3K2Nh1OLauXO3a0wX115Jp2Tn7rMAy6TVy0DGmCzeCvrrxO8ODAxANu33PyTc4ot3sx
5H1E0Y1OnVe2fMzfO4hWIU7uaiH9R2cbasvBTnTAhK2uXCM5oqcZHBxHEEkoJTrT1RXFyHTiOmfG
GwrXw5iyAnOIRt3oBv8/qcmo9Euk3oEmQo7POjYu2mqbKTvv3u54XCy3aO2hFCU0JTHHh4o32+rd
28F2VSeOosxEHp9s5JkiAPgjddup0MAV8AWKsbOy8c6MJSlRbbde/u3cH37ogv8TokwPQUveXryV
uMRxfzm1TACSkSqoOHTZCEMaA/Utg2W3AqICJuM1w8sm3xkwUSWbggDxzg4L6zHbmEcnqQlAJ9q3
Kk8FqglSIgRFiqdHRjeDgRyFZz4537zlqW+xrd3BAkp5g+qgNR+u+MMpB6Smh5xIp0n+SOBuL8/u
EJajDECfbaLXyOyXYHqKABBMJO6MPIzurHnHbNiFUqRxL2C5OB4bkQmxDTo4BMKOHdbsLDJ+TCTZ
chfLgc4K40O7NMhABFAB3Gd5BWXu/a/kMypaC4RpPaA85MjnnLPCoDRQPS49BFtJHJUDPvPF4m0j
JdcMYvNOFbEOjHFzDu0H6MQ/OhSeALaeZN79yDaGau8tKmSA+QZmmVNo3NLE2zFP/kKtkcDK9TLB
T5iBwzpJ6B9OKyvfSBqQPOGwZs1y4t1oscQS6dWdsIPTwUmwq6wXV7CL6/DExYZPa+yvWp3hmKOg
eyN/MwwfUl5rF9bGKffJiWArXfbweaf7HBmYeKhM9AixUf/xJoEL9gcgsiuAIh3MA1Jesf9wriqs
lATxt6cRtvRDCVr6k1ZWR0K3WfAiVIfa5N9pGeHB2WBwZjBeXiPR8uk/8KQjqKgCfEg3vIKfOSwK
3biFbuzf6XX9UKP3bNszX0Ppj6E+LNsvcU8EvY6ul/Vl3p9YHiIrVPvv4QLqq2sdrBBYDucvyrlu
TUW3QcsJLAPZofH6DIGNKLWNoq8QaS8dUt3GvIbe/hq6Xw88GFlWuGABz7PdbesZXS8sz+8UykSt
06HdM0fTdK8WgO7P5vpjH3LKRW1+eo1407KfFqGoDJhTJdR362pH/oHPkJy5gexQPmxnEmIHc00Z
CJvUb3smVXMGeR/HDnLelOSTeijwHRNBVZ+Cl/FVbgbgnfwYS2pWTTdgULM1iJsBm/Yq6KOdtszb
iVtnQ00e1lm+ExEQ3U/ah35JqdVSDAp3Y0UNP9nomzN/TrKQ5cLhUlT1JVnv3Ob7u6CV8IVYXLxV
8fsInSFHDiNG8qotazAqf6XhzUpjaYpZuUJgsVq8i02CcbCe66wmB5ht6HnWkgA5upkFsj1n9Rnp
zxsYIaovGVJkIizmA94n/j5vICI63fSaslyx/UxjNZC2IRuSd4LfzDu+iC0p9WoCaG26kF4FoJf3
MjygLPMKexQGWDdsdQorpfkmVUSVbhObc5YdMWd1CjjUJ1jWf0p0J3B36uocejJZeHaKt2F3hNlh
kvQPZ460S3nlhUxH7hojteaNMcnj6RuLxNzs+UBkY1zx5VRe0OWEfK4glChWp8juoIhdeGo//VCv
2kyF6jceZ6cF5tCj3kpL+rcBO1TNGJXlHpo6rwql/xL7w/HzjNHQgj198MCpRHs70KpSpOmlOwkZ
edQhcthjt7vj49WUgTS5SD9fUU3ACdlNr+758tmaGMHOBVn6jfy8DjwOAZdDel6jEy+GAHNnZ94P
CwUWHjxkPb/JJqjpqT5uoT6RoBqZyYN7Ym5z56WTiYFR1tG13QJSGXz6EWGM9zfN/++6wD7Wu9Ls
rrqxZG34Z4LbzLhkxAd57Z6+UXD9ED4q5z10FZQFm6truRWT5R6BycHy64eZ2IPU/LtbiFO0vlJu
9fFKyyCoFSnyqm2v6k6ATDbdGCnrO/gFHpxPMHagV02hXk7PF8RWDtuaKEGeDqv6o4MAFPa2WCCr
cmh2TRd6EbLwNKvpPGyfcPLMrxDhKHQvauT1BdWQ/zUdqtyYp9tUiv/Vyba1NZ/rhWOwzlwfej7v
jbhi7m25NNENL03VTkExZf48EfcMFkjkUhYXWGAFrejFavWAabJMboYquIkzElWQv5+3islsTCYf
1Y1J//Q7y2VeQEetCh1bv+NbcfOJIvr9KF10GkYI5TOH34sV10Q65GWG6jwOCijaE2wcwiAZfrLw
TmdFEEOGicI4zQ1EO5xaZBgzHLXS0A14Bon9RN8RWEYMDa8wrxu8CuGoOedRn7ryOrsdl9QDoNVy
JIIpjsOkg7ZZO04SQo/zXfssQN0LOqEhW+uWN+xVuyuLSrHwjUgNTNZndzc7H1Mdl2b/BlpFk1Jq
JRHQEibvH0WucLntSTyVylApkPvcLpmUHGfJOiugYVm08glbGQ0JI/iTnu3VPhpmoZR2eq/H+NEp
3+JFiW0g8eJ5m3+dXZX06wOT1gFhWGIVarJaPWkiHScCt6Ad5XHPe9B2m44kq43c/BVfxxLUkVod
JEad+WPYcRcFV+3arAsJi84XIMYdnKnv5jxvhRN0aGqriVucnLiBEbrbCXrlQT3Gxl9N95rBFJnN
EBk5kUZdiDwNKerTjgzb9z2jBiS+fYpanSVp85vIklOz5ja7eIMsBxp7vitRlwlyEy9I2TRR3VQq
Eiw9NPvazMZTzSj4AP5OqEk0U+L/cQgvBG8z4F41/IloVmyLTZN9VtNKi5XbimSVOjpqgYNTXqzW
34VX9ehjKkABlqEk+Bd/FFwI+iXiZfO/3qm7gHWh6ki1YMVCFyopuElOswYqUSvuC6JpH1j54knF
r17ZnLeeLyVBUjhPwLlBDJQRVHNvZIjVFQYhUkMPJjCVirL0O7wfJihGOcukzKU4Pyg2zpSJOssq
YtvvzHFlIYbDVkJxeBcWHoQwPe8H+BSfA+Fyln0zy9+68S/qYRPuulBMolSvQnFXCDt614d97h2G
/OqCBlKkZlRBQI2ud4s8OEGVlUPztN90VkdpnU5uUXZUWbNOcsNVlHyr2I9aYYAHxA8bzVSKxuGn
HJI6tXtV6n5pYAV5t/tPmaQofFrgPOYjiOSMoboIIArWpdpID+la5zVfb+jpMHiXyG9pn64Ym1yV
C0dcS3DPfmUZHqO5IwIQr8Bh73fn5ij3M/UgqrgDdXsUiogPtwO8+hCsFUGiqK3O8JR6laXz+lHd
EF8Wrx17OX8r/togcWht3A915M6/NSv4aSFc0iq+wHtV31Vd1aiJAxwpNFemzBQOc8tyUm2OcDSG
uV41Owdju4dcg2J44CHRHmfH1czrlfkLi0CxKvH1Z7iygNR0MCSEEjWFvmjvLTDSHBTpwsQuV+So
U7PiKPnksRrShlMRuEEE8TK6c2jVoQ101X2KuHbYATd3zNVsrQxdTdngGdmg/BwUMeM3Kl791A8s
FzknTIqXtv3dMsfu2bkZvd7kBA+R0ehucnStzOI72AQR5KKLbAUjErGfV+6T2607McLUliTFYq05
EkX8gCxcHhcF9qCN16ptH1g0KIaCHg6NFfuazNctW3N4IkERlo1OI/m8Qd8lQYuyoP+pxZKvE6NU
IDMqnnA4AAzFzqylTJ8/1g7YMqBF07uGtl6Mba/lkm486XMoJ4HT6Tm+0YJyyW47g2hQzz/mLPA2
wPGCLit922S+zmmQ2wlIWXGRh4f38ATER7bIB7igd6M/6mjqqPXV9LSSgoY+ZX2BQVOtzqqtmMCF
nHf+186vQlqpN0OBS3GfjbIs7oPyx/8KX76V8PKvCa6vGkRIaSCbmxqeOvDIwW+5lKnOR++Wwd5H
jk7HldxrkZB/brjxwYJE5fr/El6fVjbN++RZ5CGM3JqzjcjbTbCzXu//3p+KbLXZLd+u73c/n6ZA
ZCuCoOchwvbjFCXqiRL8mt0HxAjLavHxEbSvkg7ncX3FbcugrY6dRZbosMARkBrxeB1kNJell/mD
pUAh0SzLBblY2HuikoH63u3F0Zo9GCofGq8SMKtLRjjODTLDQGEImKLNYsYaemhjK8MWpLdgyw8j
f2ohMRNK5+A/X3q3Z8tH2ZxqvkAorwc/b4+zaB/VCCDLd5c7JsUT1n7Ubshc9BVP5njilo03lTaK
svLOz+DPV5wzZsLJ8XrgzAvRwnHmlfxWGMoeasfdMuyx6MHKa3NzvOKMuseKjQcmwJnGqBL7+2CN
cCH4ZeLzRJ7Ss0ehOYYnLrMAlrwwDi/oAZKlYtKZhvsc1Fpz8+kvoSiiOG3ohMwEWu4CMuU7RcPV
YF0tuKksyFmkYvameL+LqWyWDroV+I34al6B7kUipzipDjOYNfFFVs7ITyDZyCNVvEymsOSTZxdi
FDy7ZIIfpV2h0cFj7j/WrP/w9dImLSGFJB2Vz9TbhI8DYWzGObPxH8yDlC5neI3/Nemoc0henZzj
wHTgsZ+F1j0jIfhhFHcOtwPp4ENIkVVW9TkDbbKzFymJyHMxeKowlBAiNZwxedo3oSOHel9A1bZN
yPvafm8wDuLj5UaPkxahIAPAStegHstoi1OQM6ZZOT6pl7IRiFxFqofW4e6CcUQwhnexLiQLUd/T
MQh2eGJIsZ91r1EjFXePOZ/2LuLDnk0gmqN5XKDhyk04cPK7cUT4sLFedoPlyEJhlAis0uD0xkgS
WyRPIguGne35pobWEvt2KVX8GsksUkOCSoEIoepSDIgUcsJrRePE0SaLF8W9iet6mjbC3qSMBv5D
siAlqMoj5v4qqTtiYwA8Ze3IjvoIxFaFktqU/YZLU9PY+L6OLvYJnbbTvxGh+oDUd/IlLSDg1BUI
5sneYaCbc44MupRnW4MYROuvIqnf9Wa/FuQHNcY9vfrA4El+iaF97mMCs0WQhGQLG3EdPtS0uybl
3IikZMH4ZLPc+SjKqwQ8K9EJDLJ8bVzqmCENPgReaugcvK5V6XGiQm9g3uJ22fgmTQD2S/teekdN
k2KSH36Pu7mWW5Kgf4nt4pLNp3+W+qm0MNyZ/xr5sSmKvhS8dKcQVmvJ4WP2HMP3AkoM/bH0LhWc
dkKfmVljBbgDO2E7RtXNFb8XAbdFKHd0fsL6HQTxJD+a7cC/J9PkwJY0dCfyQoMN1kTlXJwFkx6N
MxwXnwNSwaF2CChI0NQ8Gr8Ci7ib3V4/dcExXs1N/d9gm2RSAxK+7vd6dnxtRX5pWBpbFd/TFOW4
oVwDpuk6saTxcPr2CXXfxdhsM93SfBLe+Bi/PeAoeaKHXfj7rG/UMtFiHb+8knYsmA5hckx9SEo3
o/mH+IYsRjDI4WORkoye4amPYdNeF5jJbWyIcQLcfcUoHo4RoOoQMMJIoUYlasAK+YFguVKAwqrB
ud/oXkOWj3RaLXCz1BS3NsV5SVLolLRz1sY1HgFYoP0ZXBsJTUP2hG1n2TUHwXtH4DlziHAv+Bdz
I4MqLx2jzfV951VX6YVVqw+/a167LiJ+zrjfQXpsH42VzI25/bq47ttlJNIUzCaFSd4+9noqoQqc
UlDsM6YfXRrxX5IDQQn9uoKaII5gBtADo0G2Aq10yLzU1tZM6/tY9PCgwCL6JX930XfCuAWLuFin
Vgp4KQXBen8uC90Dt959chJHYQhsrLLIUTh4tMfAUke9rncPIdCR04Ggjs8TdYzAbzxJkcUfxmF3
AqxqGC+LU65TmVrqaXxjAOMnDdWw/K7TYj2TEGrc/PpzOL/2B/fyJOoy7xUrhAQTQdbqYmBRwSxy
yu1StCkOUM3Y9nxYYyTqgXgaTO+U92vpWlqTBf4Ub28EPh4LzW4lOoNV1D3oJdoaGYsTklSvVnSj
xxGg0DRpYAHcdneE3CvcpgHidQBtqZBkxPb7lZL9Qrwsf0l88hImY383GfQwK+uo+8Z6VV3fLBoI
2hD0p5pJGmPynTE9ucyns3aou48fLe6YyZS9S2Xc0EmJGQSSruFAJfvUucdFwa918CkTXoEMHtGO
JBYtLyKfQCNjWqAQs5NUV/KomdYyevgBUXLomHw9mh7+TUAWz+1r/fE89wcEie0haar7yxI8p8lz
KJT7vh6b/XjAcI6zL7oye+i5eRnfmNPTN6HT7tVftKg1+Q9DuH2BKUQKqMn376VSqKC7e7cz0qio
IP/e9+We2bjsxVKE0UX5OnO8AJJlO8/208d2si1sE2oilTi9z8Ns9v/0BPISc5UszhZbM8D26srt
EWHEh21bh2JgwukXlXV5zCeKGI24jCLIYqNTrjMbSX9kriISuAg5FArjU/zqr7Qhu94nZcJ2xLtU
dDPOZ0psEmRP1m6x7xtR4M8ADeY6VeOgAMBTBCGop3V/RD4p9y2o879qaAoGQic+2vrtBJDr4+ir
MzfEVWu93+4zK3JBtHBUCK+skbSVNeCty8yZyIXcc4WwawBHZL4ZnMsmYP/NgoZAYTLybp8U/kVb
fINDmlgfLsEF7lNMPZbb+ePUfFQJPnJxLE+TQXYfC87UbzHO0Ha523MUmaAkV5Wv6Imq2WMFVNLm
G26hl6VYap6dWotBiP0M359tFTGJoXoskgmaOHt/iqFo9syzInyeSniJ6TFYVaR5vk20A5KukTQ/
NzN4ILPgTh1d/IBr0htvdyA9WK8CUM3dqwb7/C1s81GtG/fJ0molxZAOYIX6HwElRMOe3BoaqXKB
pxzSsvlr4HcODAtOyfE8QEM9cX3ZwMCfN+cFUBFEOTCEXBTq43S5NSdH9Q/ykN0MW8XUi236EJlL
jxivrj/o0WwqhevI4EUI5L/cQNjWZkXx3uEmW/Mp21XKJRi5/tdrYUqc/+CSZsfAcDww2qqfHm6O
SBv4ly7NI8DWtioJmxbQ9Fw9jzT8w/Wz17OkZPBU7SdFBOF8xM7t6xtpEpIcMfM93C5KMhV3ehCO
5XddLn1iq/UpQcKKpUFI9GCMWBxC2LPy7pZjUH02tYdErioVCsW+PSwZaeZzacTxrJAHAfBIRCeK
4BTc7Z9DeQFARvJ8RZNPAZaV6Oo3fofb1fsdMklSIOjTayvEg+4a1K9oJ/9bmITIprlHxbYANj1y
q8asuGyDNjhAwXqsQgLHDWh7iK8BlvchcRy8ePkxR5OCjdoXtqzQEVMPEjkNa5d3DuKcatdxZw0u
YwtYrUEyCcRuDqMI1NBNGO74G7KN1sOge5RWKQr8x+BZ5PcbXNu9zgH05GVU5/B2KtCz4p+Gf9r9
vxLQqHgsecT4/3gBvsH//e/bNGdFWKzTFdXrEWPHtO3bXEE6v5kIYmbP+fMis4nNP+lP64ZEzRKS
V3+cHIQKG9vZQRNO8UlMG3csGndPInw+GM6IB6mMUyxoR/G3oW+7uGMWD4Ex2e0BFNjSuYK0XkKC
+LiE5d9thcDpHqn9XKlMjIa5gnhv0tr7+l/WkqQASnLeSVzqamgMnSulxu4I4fqdLl1guFHB6VuE
IOESDqYK94PA3lXakwoIXFEP+hXWulNq3TSJqBO2KiqFuCb35mvvjCVE19zUr5IKBtfMBFkhcVpN
XoKb0fFquNMu+bvthDNimlQfoVqqPdVlgCWBH3rBeAWmkFLb2nr3ZLwnTJ6MZMjXiN5NABexapM3
S0W4G9Ap5qR/gNtkQHTd5beELRi+Lni0nZrh+j7Jk2brjVCGCyABctzB/Mu85ydPtgWEAnNV7vf0
YeKpod+43TjBecqQydIY8TZ0hTKvpwZPgIsC0LC6eef9TgdAGC8hpSYzuwTn/VfReXuZcgQs/c3S
wsdNAPFgKLRK5f/Vl/m8s4vvPhE6/SJTC+LBfaJImoVSlzNRCZU+nzHSLX8v7Wbdk9V1FNndG9JW
7ZkqtFJmI+kTiJpCWPr5Fcatdiuc0iaH6bCCDSYyzdhARJ3p/akX0rVnz1SR2R2sLJufCEA6eMKl
0bNRQDUr1I9BU7c4WJO40pilNbI+RbSiS3vjHNAQaNhObglxXAJnflDVpHU57XtmCsQugD+I1+al
346VpN4Mu828h5C7Nl+bADxazilDeRrwwG2zfpvD4Wn3bRRrDYHE7rIq5ZEhnvoLSs0kBnsPGVpa
4pvn7Z5kRgvLLUz2ntw/9rE7qzAqRLLZWZygwpvpspNVyG+Jv4qdYAxRIGQuRa3C2hUqnS6LiJF2
vHNtYXHLRvcNi9+Rl9vuQKxh0TA4c0mLaMA6CL+3ahaJkkxUY4kGS8CnTajrtBsGOp0EIELzcBdp
led9jwnqXmpIuynOYzdXDEn+o+n8PZR4UyeOMpDd2zlDY7qJLIE9yYCkDcOOMyJ5/y66qQ6RtVcf
yS+PIdNd/IANMEMnAgxowJOprO21s82W9cYOf5Fa/x7qJDt6YwNmlfYVFVAZ7zNYqthkDEmEU/8J
0HS4LAeF73hAZkXiC/K75Uh5lxBZtmjRextn36rYMvKDuO3ZLKXSa6/wHzTo4aoUuJ2bHLgab043
GU5qDcyv7oqGQyZQvOwhAT9tPf+0WvwOWqjwO2xv3MuE2dt+T+al08GCmJwfcVvz/LEy0tEi1OEA
uQ17ugYuHdPuI0QxKb/JiArmAOcLlgYyGvJI3TVMSlMLxDTUXL4TBtiXxG8aUyhhB7Akn++iK5fO
FbHq9AOm7GX6l6+2XG1TlBsYqqCgADqSMBO/XDSxKMSAzSHFtVh5Ss/NBGTVTSD164RiK5meAlq8
IZL7gb7r7BqVHmp6UFB44bh6EU6Tgsyj4mlAZCKamkEjH4L7jKqbfhTA8yEP/+hS1ka8gxM2aD1i
y7QtH+i/8mx2AIrKOF6Vc1ZCHv0Q+zbPVcSSt2J4AoQlH7QNmxuuP2k3ZPLAm09zE9CK9B3xXUEK
IcyHEcsfYRO+oI/wGA9VsTcv7phUrDzaz1ZwC8lv9O/dsZKOiHtvcj5hr3zUwQP2vD89ZQEAPxG5
P6qmIncafnIl2dBj4ysU/0rrJyzEHW7IVOMfdyg4FvEe5bbm/8dZ2fkZCS38YRaWPUXLbh68+DnQ
XGwzf9/bbxVwbsxBGlj4yhefIG7w3wUn/zLs91FH8iAGFAjFFHJUo1z1rb8VRGusaHYQEGVbJwsX
JSNVJoXDzuohjj5erZDj+IZfuIei5nB8t+LgfDvLKB2Jak4ZVkV1u9Oyp+JWxj9UO7DlCQIq+f8q
A53CQ/n2Tc+0z7vXb9o8LTRKmhtUdj/w3BOmB6ahvKBI68KMUe8TtQ5AjF0w/ZzZj7//z8TbK0ZZ
Nl3mQdYiIudRhqS4/0vdzXA7aEdQvWh2UTz42m/Drl2vJhZd5vsP6xfwBfHBh0LVtSdcnkp4fpIS
FcdbicPoXSToxV/nL4XyjQkEtZDqpa3/ThiV3A+41vBf43RjKDKdR6g5GeDDvw692IyV/eanjkjQ
hu+bSjaxo7ZtcNognmqmTBj2zuyZhTJx8JdAJQWpOZjxHefII7vDXT+dtfGdf/LX9OKEEY0CYOPB
oC7dkrF6CKwkB9VPwIFUDS3vW+3bDz9x8Ysu6AjoO3BSSemg+OluhuCU0XorPtsSgisRzRMFNBcq
khQgQEZvJKdfLMFjZEJOeWu9HViDo0PRZXD3+RbfcKJD9ikvPXW4iJatX36J7jF2u6kEOweTobWR
nIMWkkxz5CmyK8tEASUjTZ+nq526B7DonicelrPrsVZNZTomevHYblt8l2B+QKYHlx17guXJjt8N
5pYFvhRw3yIQGasO9E9jo7m26uC1GJTMMDF0FQiluDJUafL5QM4xfw3FM1sTJRLmOcLc1gj7hYDZ
JeAkPkIRD70PG6Y2Sr16/AU/lmFiX2rIS+mHZuLcKf3seHdBkwwbpOgrO689ISX+a7xDQMeNN175
SoHgzye2verRVEN6qAiuFUbn0YgZugGvbpRJjPiUI67771dI82wlxtLUBiq7IfDqdqlzRJRtSuLV
igmmwpN0d6braSjTbZQWNisbSWX11iLndboxbxYBsIX4lUJaEQ5vlamyoMYx6fuooT0H4Mqw/Za1
9lyh3DmVZYsBT1BwPVa6ZzN1f5vY99AwG59YVSwFqttH9qGU4EaLfhcA+2AFXbOUUADGjT2DviTt
Dq9/nulGac6/eCbPsvH5MUYK6ApdqTbk5W8QhWw+KUtYU5OOTD1vulH4YB+RUA30zIlHdp+UNdpX
QLx4OAp/w2ufBOowqyVtgBAKIk1+a4eqPNy9nwU2MT18bl+xc4zb5FiAPMIDo4J4XoPnsqnuU7kq
O0rzcyHZo5EXPzLOygp5AD+HBgCj6UqOZpZVuBRFK9+Z5cZvWi2ZeHilrf07zmMvwJp7BuZtt3wK
DGhZBPY9g3NDFzC1IlD/8/lG0p48ZKALPD1V1kmwefj8DJSvT4ILyt5/9U11/5W6uCxjv4G8Ba6T
bmtLpJLCmvlJF0JAGp5sQHgOko/N6RAHwRji+qGfbDdMHgcq9sF2t8Ub9JJOir+F67bJYZvccf6c
xui8oweY+To0zGt86cEWSR3f9U5t+FyjVN1wLT3CV6YRJHFyxLILGqozjRltGIQguX2IpI2J/nmm
kp4LSIaDY3p/QEfvFsYttiAU2tbQbJUNI41q7IQIr3qL7ISfeE6Vev7OJ8xiesDOyDgEj82/Rwos
bCSEhMhoXfd3UPOWntR/80WFFd8krE9zCK7WbWFEbIRCpolZ+8Fd+s3xHyneI9rrhGIbdJSzNVms
aqr377ab3hZ0fJEHX3LRkvFWOufhOw0bmp58BCPkZqbTWWRhA6rbxl4eSVnG2M8hMMEzDucLWinj
3Tpz/tDZEDYJLOESdFslG53KUFZVGoEz11oTYEX5lI0ZRstegtxC4hpfAcIAMCQyAJCseWm2Hpa/
srzrPYWwCvUtV9lzY04cXOFf3rPE33QbCqjXpP0AUkq6swcFelIJmTEt3osboREG56G9TTCL5jr/
I/VhZA5n4EayxKCQ7vX72rf6iUlyiSCJTOxqGpEvEamGv8m7ey/+DrU83cS+mS5W3cMdKeQv1XKa
8XT1DICuun2DKMTmigcynwTlYnWjDRFSh7hiqOVg7cmSoD4s1yMUY83FAYUGE1cpnp4K257NKBjd
YZ/EzAF4sywKAlz3r3INMRoxuxjptm2ocRDUnV2M6xD+v9S5Lz9QJA7t0e+lMf8yfER75m2ceKip
ThLdi2a3ugL0fzxhS3++1wx0lBva11iBeIzlAv1BX+0Q1CMjK3yKJ7FGs9pALEHI8c7b1kerfKtF
+yg/J6xjotmLWD0ApA/GcS77QC3Zk0FzxEE8QmAxRDqDHPeLBLoly/Wpoz73CTXKldfpHsUppMW2
+xSMX7vfVXnLfKpll2tJgImLv6+wJZTtJ6lWlnlRZVa8riOs9g4XRAv7CQRmm3OPVunbCmHYGoSi
MR6YSoHRzyD97C5OeTKxv05/g4rCjQKMv7o+++zig6OV1a8tEprPzkc+UTJ8XdAXTozTIFvXBejv
fLjuczc7M4NLMKBMxIbdxrJkF9ogLj+t8zyOGCj9XmIlLow6XN1LG48Er4S6zI+natLHl5lMBSAZ
7vEFQwTIwrf6IaQLs+eVCapF1ZJY1y9rLwDCr/MSgCJnPFwxnKu058GSsUlxUq8tFhe5lZh85DFK
1YEZk30WV9GSJX/WJ3vd9PgFTJ1qqFJBu9BQwzs3Imr6Rtb5V1dHnBY1jlUyQ8TvDlFIO+asMwcP
Z1jl9RTJkcFSgvuYjfDZlELvD4gV2SvEZr8JGo24udVAEf1jBgpBNq39DPihR9LymCZydbVVOJLA
G7x4nox/TVYDd+SWys41T3h8hA29joTwmTiRzeQUo2kJP8UtZrrg90ftG3NkBXyuzzkz/pGEnL91
lr0fY+bkWTBg7LOJltgb0PxY/O1Fy/QFKZuWj7yRYREe4dihPRwON7hnsMkafxHysZNfm5UTheEa
ME7typjCPyXamiEIRYM0G44+uquWOmqDg6NlDj34lmT9tz+kSnT1EYWiPJasURA8KMyjpSnmzdzn
FZGeggg/BYYvWkDC/iFv8d8T711vy6caQrIqmj/ESCFutRNgun/ZXIwN9Tol42oT+uthrBgpqHKR
ZpOXgR1R/lzIuzuWAoG4aYy7voYkc91t24SeFJDord0CsU0ScG2SY+n/on4DB1p+TwvwsIP+JOJS
XB+bYP0Ua3pYBlfkgXHgs5pdJuu7YO/qPa8obPd0X2flWSLSEfgnYvVZnfKJFhdVbPETJFlSnomo
PJMFzKdLALV3CTE8Mf9uWhGT2bbtpenJ/8f1PUN5/OQPAEOvjeHFXbVFynx38dyC+I1u59632Fh1
rwJ+2S1QemWi++PTz9hapLR6hriEdl89lYzEQu135qOdRUz95qQjY7z6OFB0/jI6W7rem0uNn8pq
8kUCn3bRptxv9G+SPCkxJXsLtEZ4xN8Sq+ApoVvT/XHrgsKOerT/AH3/Ig1sMVxn1/ye+MFWNLH4
xH9rJHH2AczpSv9StHmaPwa470izvtQSzcULQr5i/5x+gUFAjTkZSqUo3f3OjNK5i7RuWDoaXp4C
i/YQF+HZO+/CWOe8zFnkRmzOCg+kZwd02g9M+xLZ3AxUz7iBl9NN6l5MypO+ItlYr1KE/wvfZJJL
HMMFnMU9S1FJOJ6wdtD5FsabrwD3vhh2rLM8JaYECDUcLodlds+j5YIMUfh4zIsue5CKLBUq5hEA
AMuMPkNIilpPs2IlTgCz/58mMFV8TW4CP2qpInwzlZIolhHLW2cGnXqW2MxnwwfqT7Do7MZegSK3
KB5AVrK9ULXq4wHm38kUVv7cIE9LBH+D63/MYeM5jKTynB0R/3pAMmVIfE+hUqBL7AFKIUImEPbD
7KZEu7AIZXu0JbBJoptefeEqY3wCP/kXdi8an1rULo8K1F7jzO7fEVQYj2Xw5/xbGCV6368uezEf
frQ8fscdhiaXXiyajTp1nJqf+h1aHPdSF3jxkymEtqostVTI6jx/Gmdy92cRGmiz1JNYDuOLMPku
mkCib87mgjBSIkicZZGDeKdIKgpfS4tQKQ42fsVGV5zFVeSQpuB6J8yuPKqDp+Kj5w3uzop86NlQ
1bfdB5/SKAQs0ahsguLDyinrExgezsUAbvDTUPHQIvE/WaWjMMyJ828cRUFKslje2omgdJNd+Ou8
3/J7zJ8GYsiiKlTZi6r7Rw1oLk8gIlMUwKF1+aJKEBKh7/3ZDPF+D9el13U0TYLPCI/E6od3c4Vb
QvGuevLFD7VfzH8pKaODR1ywPU+WYgcCZ4OvrADKlF2KLdsFr+D3VKRxOYJIED9ZowJNjsS8BLsx
l2jrr15jVzWGXW+Ba56loRAn9vK48ZnoEAp90a752M0fASZ9UXWWOFaCduzfYjzwtpqFCuIK008B
ksIR6Kli+VliB1v9S09Nwje07cdMC3xJK86sjA7T14OEpsS78nStkje8JImh67etniT2Ogm2JVry
ZrSkPM4YSLzdAnTGGSOVrixbgPoIF7m+CaNb2KI9tHHiAxhXTABcDKNcis8dTUkWYAf0pu+OZgo0
o9cJ0H2OUzGcmyD91BCFTys1LpSS2Wq4wHyLA/wuy3NAhoVkOBeUoHACtU0N13O7jLSzAz3IObLN
YwNnEhNt+Jd38bJv0x4gFFAZaa1agh1dKVfsRVIZOwU1Qf+V2VPtJyf0N1n3OTDFzTCnCxwmnm1T
dn7GD5lQTC3jrse6OvTZW5TvF3N/6H4iIguas/VyhtIOihVQFgEUfdTm9FkPDZ6ANH7k/x4ro9+w
7RvdP+G614WyxqRB2ElrS+AqJenQFZfUMRYyF6RltiuFoeN8jSKcuGNhVUxj7MW15QcxXNoKypIv
u9nFrMAY6FQhcaC/PlEXjYk32jRWgQL6QwVyNFDhAxbRaNXGkfsCnLB3RimmxAqxIJv0O3WifCnz
bnqAz3YrU4jkw3duC0VB0SyV7x5SctLO4yT/Tu85gMM4SfE3pkmM/5H+DfbC8+M2U+mxCW+b52wQ
BRteqFTUdV5UIDJtT8G/3UAdQNU4fFePDSTrbi9ZQRHp46ZjP3a/Y1hqAxSGbW7xYdR86IQBSlwS
5WRqdMr8A/W2lHhMUZ/bFXxSh5yPXAwlQ02eOxb7Ny82EbYHIt3MUY65pzMqdRZott1eqZzwfXxO
eNxNAJfPVRytxwFMDtvuiDbxOHz0GXnbdyn1ESDcHih9rFoNH8dXLudvltmImb/FckLVuPv9nHn2
KiL33EtZINf/6jXDmFASIw1FduLoJN2baifrmYQ9avJs/V5pk6GaCTqGvgYZ7MXTmD2UafyDeM9z
bO2B7betkGS6L1k2OUY460OndnjekAEXRNdiAk/0drjwL89dCBtlTgoOBirHszAx41v8DjWp6TEK
6c+H2lXaadIdQJcr0HtYcUpqpECVfl7qFv3LHmXqkABG9ivwsQj3bZ/e7397LKO9JVmz/VyTA0Fp
6T2ByVoxmL6V5JsSwsenRayRDlrNU6voy4/MfXtrDdlvYSy/uFD17IwMA27yuCRtf5+qIKPNb4O/
teKsFUKrQmZFXccZ2JPcnh6lSbGzt+jMj0hMffe4w1JgZ+hyGEOG2KRuwDPEn4vZrxXMJMFSgUDW
oATZtqdGQCr1IwwumwNEXY4uoNQIo6aTNn+XxYjP0I0Pp3/22jg6HOYX03a0MOpEDpcdggfKZdH7
RyKPCfGvMjYTmJF32plDOMNYJzdfSlGQ8QItY7joZX4UAH8V+hwGgY1uOftGQ+0PR7HwODw+YD66
Q2TwBA74b5png4MlnPvzHkP7uJkXBxpan3ekASlzuFHLXaAMPPBxVctIuiD/+IsBn521ZjPfbsmq
QJjsbAviEF3+J5pa+vHi0MGbXHip5DbZxihnPb+3b+Ur0/S3Pq1hJ6VKlNQfbibPXV0atlEBbQ5u
AqNLR7C2b7nUJ+2KrIQ5rJGRk1+ssWdQWXei6WRkwT2+iEFB/ET+cSCYMCzxaJ4OPVzNbFd4StxZ
cP8ELXNE2ELMphuKDorDkA6WfO225STVfBbFVIF/ym6Q9eRls0oS4C4HMy0UnZE49wa4pQTBVVIK
VrM7t8Ge4xFaIohao6uIm0G2yiTWOndJNR8RpMp6WjXdfhf+tKTMBy5Cs+NPi/uHa/6hc84xSv7Q
BabgGYk3yLEy2g5mWFK19YGv4vS3sXjOtWQ+qdLLS9gvsKTJAQQQs+3aeQh0v9ABWM3ApCYgv3VK
WhyPpx/6QTssTLZc2wUUVAI+rrHl7K4Cw7LIlQ4SgWN2omSmbJeLRYYDWba9ER4sXdZwbz0c0YOP
KEqG+YKfLCDBgGRlSK6NqX6RsJy/kqc/zTztlaYWO0hdF73IOgVIJemp9wQV4mnuEYs5mmrQxGOm
yN5/f6QMyLK+j32CRvjk3dmbfYGNWglitmZrOgJBhrEnZrlh/hE1qX16nP63jV/ZqUMilgUldNTc
e63SanKjFdnhh3GsL77LOOLHmwtbQDubo+Trr5B1atVqUhyKOGKBCvgtfIFL49C0GPqajeLqsQfN
sNAD+Pyz+CAYvFtdmfEhJB40NN1WBBDr8bX03Dcs+tWQnPg9mcbWFIqmmEoy1AWrlCDXQHhr9Kb8
3EuiM+NnhhcXJv2Dr1ukj3juXe5BVY6yCqv14Id2uVf3iJwOy+44GevsKKg2HE8IJ8LiBpA6ulf4
KN8qRB/cEZXPJ24r40f76pkb6qAWrUw8deUdAMPQ4wlORdBWfUUAZ1ELfZvMm9ZDw6bnuxfbjDYT
19f5lofYAaOcmtNLtnYz+uoAqRlQxERdwY190NpjcwtIIJlsOcBv+LuEOY6XMWW4r2Cgxwcaw+/4
PsHC/+6aBGV8Vyf9jbNxH7P0l2CAnbLnDAkM1FJDqF3TIalsuDJlZ3mtCb+6LPDec5BKAXcQ9RXp
5jIeJDR8mSHa9QsydZqOYC2c/mKzB1cUTqDPeh/ib+icR+6DH6blveX2yJ8Czc8pa4d1W7G0adFg
odx5JprNinU/upTupJZgQb1A9fQDyMppTw/ss28B7xwwzcjSozgmFv1xChoDYUm8oAcUfPSJ9BC/
+iS8aBahGjonTQD/Kx7wU3CvFXQk6DVbIuCdeuJ2ex5MMQ5FwTongEMz9R36wW7ohD6SK92yi1ev
X5NyjNndgEmJOeTC4EpqpUGOgwHiuIFTIm9UvFWToS+7rCk0tBaW1h9ZvX+c+SbKAk6stHNE415S
eQxwhBhURVUTzsYetMYo9isS53CAz307NJcklwWA532WY/NAZsCnqKwQraLDKFx5Kwjr7IqVQX8C
DMszM6HgAtXaXSzPtHKJbzKmZ6b6tNTQCnEZbCr8MpsQM24DC7xalxPIoL8k20QzrqtnVbUFRuvW
evfHPsqm0qBSKMXL4hUoW6X9MUFq4gpzF2WqHLwnfu0ihgEHQ+p9Uon9PMRo0TYHGAudG1kXreZB
MshidKofCkPSQz96QZ+HiaG3nAictQJ33/cJ/YLWrKPSVOaBjYW/E4SIXbGFG86qqfcYruycfNYa
F1sopG9HnKMA+0M1aGEGAMQLtNAaa0W+/TIpMAeVMc5f8I8IyGTIu2+jZeaz+a7FE+AOX5FQ78jV
UJah/nLp9wTgm/xvajDdQaHja06PJ0cRXATXQg8jMpROCDRhfLjo5AI2rLTV1VaI+BaGmUzj+Y4E
p+UccpJWhfU7HQJT6vFrEty10lRtVQpYMOfgXdyqTJ76rsRAfXv75R4/+64w81XvsKOV3gzYIQ9V
G3qu5JZexbukvuosqKrw6PskDn7fTTZJ+hg+C4qaq3ra+Vhh+qetOkFwfKX6kaXM0YeVWBiZaT9q
ZyY7C5nW7BP0cDwhX03VsV4IMZEWNSKXcBXZkhHHRVCzMZeh8HQKXd5naZPJiSCRwGeTWde3rEI3
Y/B+o0B00Y/o4u3NzktEVbqrAZA5BrKkpOG/ZiWg5nwdVXPvTsuXDTtlPbIDXuSNWyeuyQ3loQvj
SyjxbxPcRQQJLV7bxiWeVL/btPmudVj/TyuNX2nQmu3J5J+8JyODLMNiO6sSijUujgrY1WnMfkqc
98EdfRO2FhYb54McNSAKJbtksO0olc5TKzYwrKz/lisj70hmKYdAm805k4Rx2L/sm+2FkirMZzbm
RGCoXc+f6kToHJ6gveAYahHqvGDYV1HbH5RNmksDyotY9oDU5Wh38l6nwnhUDnbLcstwoky9e+2K
QGE/lI74l124GYRzEp0skk6hjoju9DNJpkRtnPsB3D1Ezv9pvxpGm+7+DQQBMDv9nu89fkpGKU+5
r98uj0m57gHiMDaNvKKuitkCWA3wzETA15xZ+U9gMWED2URhEDTzAhAA+MQLHFfBkwf3qgnaiNsg
t8utDqA+g4yqo/Y4nYKzTsiPsIAT7WkRCBEDoeT6Tr7HX+KJA7pFveKldt9Xi8m9INr3AxR8qdvd
dr+SFU+5Re3ikZWzPjLsM/Ra9vKH2u0lrCX9QOQd37R4zg0xdlpU0vSMX9vVc1z7E0VcqcbUBU25
807lY54ZX1NQQOvL1HVDw73ccgLVxW3WvcQ0iPprw3RE+KkzR4Q+0Tqk/nrW2wYkrtXDZp0BQIpJ
cZsEDeYWr1HwY536HUmut9vT8dMIR5ENrf0Stto7SWA9UBf00aGCcRidjN7ssqkmqiujkNjBPRck
NfhT9LbhElYclPMCPIqFq8wa0EH6WkDz6FLJwdVdIWK3ROEMe9YeN49nTrAxLfXSOo+fqGniuSAl
uP31UOcSMRhTDma2ByeQOcUDHfDod/uzkTGDoML+G3DGTLd+wMacr2+sXXFhkBd/SuUTHkbhYkko
XgpQ64sFV3hXhMnY5PUq08u0A9A0EOaWRWaMAMUGCoICA+1gO4lUoKhqbmxpaalpojeoSz+7NCNW
2qXHMVgEBpwsyWh8l2pFu46hOkeSBb57sTb/faeiy9OSO6BcUZlkN7b2hw9WP7XvqWcwd05daDCb
TrI7xleKM9dcXYTQmi0oeNziGBzCSEmgavz7jBacDtUdCk5z1I3v6+pXYq/bC5vz6kmBXpYKlOqk
gK8E59qIp/8gLseQuil+/nbkbiu9nA1898Wkf3CCycvhuICxJEzMvvEUHsBZ5M3g+xdMu1pm9K9G
+F8LVX4VDZwJIVqzgux4U2Y6J0WFfyEsUZNLPdrE5a4WNePE0cpkJ+ZUf2VR30LPTZM0/v1AMUmX
qYHAfOztUz/lhDW09OEYZc/zA3F+ktEM6VNR4RDLUGDvUavUuecDEUIttfqXZdrVZOg9vENXvBze
RPHjM/UgAIDefoUvu2DpZSBov8eHx8irIhmnL99ofoe68QDz0vY1ruizlIM24KnypFJmwtI1s3Ii
N5WLKFrM4ryweocBKxzvzmObzBBjMIHIAylMJdkDr1E7C/THtGimaXyIZTbOtHnj40/MmjuFq+P8
RBuqGyE/KPjBx+phh2a8aEcy07jePUemi3AaWTbJV3AfMmKm+qcYrYfSug2uCnMmZ/Lt9vMUudjX
pOf7Bc3OygQj9YK/ArFe1kegoMFs/TDWNOBPb9UG57TR3tncbb1Pqam8tIogLWt1GwoQCVxiRTkb
0QD2soINQvdlX49UTh8pfnGh8bQghBdtcFCF7y2sWdeXkBit24cm2sMPFZYqe5ykxvdirFEF4qvv
BG8n/KHsWgKnU8tSxAwrgWT2ACJOnHaWC6N5P5Hqdrg6/OKFdiUJIdUeQjqul7rv9kqJQhk+FqZU
wjrEy+MSDZRe3MKOlEOuxrVRnBbM5QoN5ekbFp4dm41WlyfQ9bDkmg0EZhiu4+edcOuBJXt32FiA
vYHkFyuzMawj/7a2DqdonJKbm2bUEHV5TW64vJqsl6URyOF97cXSJ9qaC51vRCOoSQivuuAddZKf
gCcTjOg2DSgHsoYvxWTST6ODqKV7hk2DKPP7MNGXqI2a9u96FT5/n9og4sAWPY/OMr4PybEaAqdj
IU3e3lMGZ7Ok6bGAHWpS9MBI4Wgnm5utQ378msUnn3IPgqrIUwQsYEZyDOH+jAqBMqUFmgDp7nNo
mDjPCgPdq8G34b9G0VVPwzNx0Th+Z3CP7AY66L/8jfvwjRGXeOBQA0ruMgflIVYLpiQMFCT6cXVd
m2WpnyxaKAB95tOQ9I0UhrH3tOlAmiKwU1EVgNNbXLTDf0ABK9VHOAedwgRoXDueu4w9tZQ3fBPj
UMY7hF5W0HH0l1YWd7ahca5zlHMiLaDDm99N+VzsPO53LPgxWElrKbbxTUa4CrIFHiZkGtHYuzOD
L/sPLm11HQ6AA7Bi+a4jbPEe58DF63CoSbef/2DbjcQGss9oAkwzj4kKFJvvwjdd8+ZA56Ilpixu
0jGvTfFTJjSt1rbq5jruChwVaMhNQ4RAQ5VLJxSDgUp5Qs0YJB4DeBzLjgnfC0DCgBgtU+H+TeNp
FaEmCGO2IgLYhu1/c0bmiFCS3Hm3Z0sSmhC9YGsmT5X/0LQ2MMB7O0+5NR3qpcibBRVVBpE4HOYs
sqgt4jh7dgWG0snv40Abrf4m52naXThLwn4eBwTqdRIeTHtTiLszOSAgimsGV9Tk65gjN+Fa3KB/
zbkMrWL9rUNZHqtId/Yc63/CXpO75KEbuF7jXEthz3Ye4C7FjZWTqpesx4xByK4H3EbKWzFaM+1t
2+nTa5aK32hOC/UQr7QoCW3P/jYHkWhgh5rXVctcmIwQvachyLVl2CmVl3nz/DN8snsKBUnkaMQx
OAlXdbrUUvnJXGmtbbFkqf59LhKItxyuF9i8jrA9z6cMLmih/MiOodR5iR5vXHEoH6gtv15agasx
B7q+ic7B2/yNMEajN/trRoJ/3KOYF+QL1djWDxZv5NnyWmLURP3hgkiheSxIX5YHanD7onnZxJpO
mO6WNWbRWNcaWTTGrw0Ff1ALvxnIuA0QDf8Z+945jsNIdAxVBPoBGn7IWMdXEwHy1M4RuG4CFmjS
47B3AS1Vyvj2y5+VRYdoMKr3ALF7hQG/QLB1eMUdeLGsmoVzqSOgS8H51sDZueqQk+Sa/a+QOlys
wb4nDdpktAvlsZrw7bGGhP+VlCTKzf40St4iipWN3ybtWvTuMcCTAwGUvsBicRl6TcBLBUYN1f8/
Wu78Q2EotUGJQfrmrKUhPLj+QP0KSVoy8LsWCMc0RH9vLIqIEWRXt5pkSWaBdFzoOzKIsH8mSlOU
7mPBY8KVva1BaN/CgBaeJTIksV8r/RAN5cvd62sTr8zSzu3Tj0OIgbfQb0PbG6nFpSfJ0f0e4FXA
Un2ILjtaw1onNO6l6vo77piRx06WPCSAOYwkGj5frgqx9b0sfn+ZtGkBGiyGx0wPfe0QuRdNyrkt
vtGobObEgE+yhxJMwzsGtywg24iG7cAD1KuSp/+0C2vl90kgmAsSeJFELoPVqddOkz08cBGpskCt
olIrt5lcI1QWuEWCprKb/EXuf4jn1XOUqQpsFvTmtrHmQYvn0/bcI59rOmW49qkpKPO6us5x/IOh
F9RczjqO/3r+AWRxAJ3jDkq+a388JwhxEF5PAS3hDIbyGkNi9sngLVMNt9QNqmM4ERYH4hDUOQiX
/euByZrqXsxgIgwXa3Cl1dihq7QWLgSC91WwgsJFaNbxcp251p7GgMAQj6UronASgo8zXJMCF7AO
pM2kayfVGIEffT8qjgzRuDl7okt3eN5fc0SHfzKJUe+e5qWLEBUjHeAYOjmSpgqwyB7SCWE68veM
Gv2zQI4/p7HOgjylKauwgXB3o0p4xckrfRBAu0F20vltshjCXjfa737mhfKRsFXfLrtYGjg7igpj
lnXYZg1v0ENks1vkf5ojbL2w/MQy5Yn1cmIxcfoWC7ksws7+2EezS2xBNYWB0PTntVsMjxBsF94N
YkyQoRT3j/tAR5QXJiSb9+zPRPVV1pqwjU/VCjfSueFWB8RK79vCmGYOMcvLBUCbczlxpg16C4zn
t3jqsjsNAkZHF4faho64blx7FEk/AXmkyIVQVpax3KDki1MQZF6jz4svOQRqQksP3UQm8dYmWoQ8
W/jyL+DeqUutl0p51HSZzsWamhOXKlxPCXcvVIQuB8a5Xx1jCR6Is6lQBOmb2yBGs5jwhN6sPFUa
abOSfZ9bUPbPbwA9OySATIovqyrAw2qnnWUDyc9O8907N6mMJJE+Pd+bcRiMN3vfycDc9LMv6miO
rDVZEue0QKdWeymdUsWO3s0+S9A32lFCE9Qm80Z6sO7toWHeNaPt3kR4VzUduglthL69sX099Md6
LdkTXq0vmY9hLuN30XfoNy/LfaD/bRIqlSCF77yXfgSGiwNAkHJY8XLrElJ1f8usKqDdzk9OOC+s
juUNOUvGmFhr/tvORHNiwiR7i9dLVHVYExAGqEXXLUgtV7CLbLdQUGi2CGCeeuzt+nt8/I6FmH+x
xjeEzK7VXSivBr9rvPsjxJL7N0ziDxkNhrws8evpBOz+Jqr4BYuBgTaQ03UaHeMKvatYVvFFou4b
hARlkFS0/2aljZy6GPLdPRWBHM1ZTYs6iEW4K8iVLfcuD2vUU2+ybtS79ptAKEAb7Z2c/pV0mjPE
NyIkJKEIqIRNXGijTI4Q2x3trZ+mCfJiwOPzKGMdigbEoD+IYIumOhIY/nevFYV3BaMn8oCtCpqB
Bb4jRFCuDX3feJFyxjFxS+MfZX5pVat3hkliHSmFjBmWSEIxufRARgHDluY4cnGnLOypiTkaPrSD
tmjJ5AOHEWxIQUeer3I7nNVpu2oBsSTKsxwItGdbYV4w2wCLvrH1H78ZdMJ71LPzyFpxVkuFo5+e
xBWeyzmgwhkC05/58KTRduA3O6nuXXKQB4YiodLl/LeNXLrMhFS3v8+YBozMF7nkQGJhh2d6TRBc
qKU9DbTghR6E10ps49C/mtW12sOVfRYnZVEKmEpg+ItLLr+QaNhN508eAZoy3ig77WJnebZPjd23
u1c28uhZIZDyggxy3ZxlO+9uJCNixfP9kWrNkfZU4s/GlffDBbQ1868qZrFhfmH+C3thlHH1+P1p
8kAYuCNzKsKde7+UIyecIGSivNK/pstwkXV5pXV+b2E56Q9t2Gm4lZzQqmUhOLu/YptDe7VDNpop
dYkW7yA7gEBjEmAXn2yHILqONF1EwfIEWVxVoxcC5Vk0aIQwek1zku4ObSWv+wdziXfnny/7GRPQ
HH3LT1zIPxyyP/I12x/yTJbzB2+SGtM2rS621oieSVzYAV05zb2jcOyg8Dxk7lkWca45gW7CeHiC
rUYxYhvg4MmzHDON0alR4E8Lyyvg7kRvMGEtOh1Awjd7Letav2ygNCGPADxdZcRnZwROqaMd2917
udUakpL+EKSr9KpG/ut0dvalxZzNqiDadffIxkNHwzwok5X5Y3CzL02nwbxLQmE6hsxRYkcbwhay
9cfPW+X0lOrubcUSQd/77LT2Vhz3wkQwjvSGcLLmM+DoMt4yGhemYx3MQCm06r26cqjwIS++sp43
Qh4P/PSRDOM1Mq3web1opuEkNvs2USeRavB9GNS+O7IEqrQrCJ9Vt8L5rcarXJjBOLexh0OZBTx2
rOPA/olN3U+wlusJMM1HL1AYGovNJe+3Nc07B1OMCzM/2s0rXbUR7K0lVtwaIX9vg5F2mV99FhyH
26nVFkg1f/BdY/wJcRNflm9mEx3hMwFKQI7iG0d/VcPuHg0RjZni0mVxGGy8KTfGw9dmdGng3u9e
HHf81QENSIMIkU1zIIRILwnGQgGAH/UoYS5sXLoPBVo6rGIo1w2th+YBIT3XT3WU2ZiJvNd1H32R
3QfbVCcBTWUVeiSPXhxCDJkbNxymxFtz0oXdG9NFlfX5f0/q5WgFDJjIobjzT7urbdENUogn9U5X
IdIouSYulwSCw69VQ9e6l5gqCdWOLBFJthYWsIjVe5YGU/wXf3VgpuRk6i/kj9KxEd+a1/OKY17l
KD/xOLwGAKCKsC7Lc0XZCn8dsbLDG9y5RYdJkiAXTeQIrKK8gwXjDlSpaqvukzpxmlIdkwwg3/xE
fA3Jriy78fyScukZhoDusHLo/nVRoDkUnWxpkjdTD1Uh0b5UvrDULTeI/gaGhmNGBe40vsP173u9
4X2FkOymjTVOQ0sDzUHuszgeRPyMICyzlG/7ZLkWquRA+jv6ZvljU2bGn/E7KSiD7i500dghGWBD
AtLwUMDgucb4aOflvP310TLdMI5gpR0msnFcEfVugGweZsQlqFEpMVsZ028p5FUmLkulxkeIPVu1
5frfcHBk6k7g2LaUwfHX7H1CBVyZ+T6JiO12rNlWLoWKq8l7nsXOAE9fXvoZ3q5xGfRkVgFXfMRA
QV51dekeN0vZG3tYav80cd1XPMsQbC8yhIdR1aB0HrpTuVO3drsPNC9atjnz+JRAUBa2Ca6QNAZQ
qN+rExjbpjzQ+aVUZ7P6k354reOkE+8/zeHOzmyea3UEhFR9adDQI755c24JjtSvXf/YAeLh6Kzj
70qDxobghVXdI88zIkz/hgctCl5kidTUYGXmet2MBmxfTKWCS6cchXw/Nd4WV+4yORrXBkcgfTfj
zZkWbBzWJ52MPbtzASDQzc5HY7410vTqWFX3NnAteG8FtD5DB0SW3xSDcBVJs+Nv42gRNePhDbw3
MT+92erAvsraCuxNdT/wK2bREtNHYTbN6i0iulJCe6xEcKNIlZc6Y6Wr+neK4Z0+/tbTJgoKFcd/
4o1TYjJo9vXekQomHDq71jCEj1md+0mxJZon/QazA7ZCyG69hOXqOxZW2lHZVeUuFo1dORvPO8en
hsvvmyEjU8LQryELrrcMyD/dvlC1RydxvySiLyOs1BtN6dYRBJotU1g6hfbt6J6mnc39wU8MqPbj
QybWml0cj93Xqw1xiKst6KzpVT5yH6tbFtjWWckrfELVoQaskK64bfET0VeUJ8hRqAri+uFclHfk
+zZrb8d/oRkJX/DnE9nlP9QnB9z/6zwlcxyaRksc+c9/8lN1sVXrKQpodNgGeucGmz9BDDW8I8Pg
FswSowqN7bG9viQeG8NGuXTQJrAAbHEV5cBSQuERQtsFUGVJ0dxKOGy3fblYwcopLdmanhkZl69V
VIUoWiNnseo+WY1hfR5aafw/stwDi2tEn30RFNHahpF4SfeSvrBkMsdiZp+SG9m1L3MLRJzS41An
XDtFShKrYj+P4aISWZ9/M2/eJkfiE2ZQRjIloPFIxTlk0ubX0JUy2gTDLMQxYai+Sx0RwH86XDMX
9AuolQxi3sPlrqIMEcu4kU6VtB+J3t/NJGJmkTcVgsm4W4bjk1n0k2DF80aVGM4rtSI+EIb40GK6
4KlaSrnhENVnBbNqrvR9ygQAxZZKR/Xu4ipKX8t6hoPCHCq2qp7dslE2+oTIg4vZrrzHW3BPq6o8
lWc/ZkMQAGC1ww5uoEcKn+o3LO+rBJJxSpgUHpp5MmqTSSNAxWVgYkwC/39IRMFBPAqHorvdnZOE
+Bl8DBijwEWQoWHGsnxW9+bXozQpBMLIBhcr3dnlZlK0YjR8NCOtPJhu0LHtihHTalKdPrhYF3sR
Qwb1C4fAQTQhiAHx1c18TnVmkKavnv8bx6pzZxbcWKeKaICDX+ZcX8nzhV5pCre2eJFmf09cyibk
+yYeCijTTuVwu/IE3au67iHDO55pNSNjH8eca+Fegq5zt9HDO6xFSkmaIjEv5YOASI51wC5/mvLY
Wti1VKHCSY6ajlBorUN7tutURUy2GCmFcZnh5vp148v4Tb/mePDA7NBW3ZOOFTSTmrf3iM+Iirxy
KVtNLPvWX837fcAY1zkqhPCay647VufwpKlLcNVpOZ+i9alezx1Xuw5Tp5LwiJrRXKKEw+xn8KRG
dJw5BxYH7pRedm5tUHuRm0dSvLPKQ4yi/baiGQLiyEQItkcZNeFctdBTE28BCa3j3J+KHchRye7K
6gtNBFk6OUWER6qrM7PgDFM1TWsZAgGJ//T5TETpM7yFZnXSX5dLmLo+zO7DVhCN750jZLBTKuxb
sOplyZPu0jozd7q1T4NIrn5y+Onl2tbSLkptjc4rX02v2tssKDIalW/TzObtvEbPdBNxvOFVFYJe
d6fDWtmCaa0iz2QL3SH+tbFSlYYpdkjuV+Y9xaVflyZqVd/YiATa9Jmiusb0jrRM2cqaAsQVbCfs
jGWmwRH+v5q5HfWze431IeY133HcQMrP0GWRLiB90OW6LpvL4+k1Qd8U2zewkvepkgPP7cnHIHs3
hAwg9zKDN6Sg3gSGaJS2UGeYmDRxYJ4AcK2ejeMQyFz2Na/3pQe3AJJuhG93mqP2ahml2U0ArsTS
35wYP8wnUiVVIz/nbEelMe1xMXRRpTw3q2Xd/PJ3EGUWPFuTzqj8XfJGOfAqmgKWOulHdrQXlT0r
Y3e6cexy+FAkHQu67wnlfKgcZOZkwj87c4BwSlb+jgDI50IPBlhK0RbgaVDaXfvOEMhuLRgONN9V
TjKJIsEhTQBKqYL3hyDoUyRMhe40B9zSIDTH6R1kPVBqxwLDHa705PFTUviMk/uy0kzT5RFmhzDc
KeDNsbdCsup+ovkHfvHlurOj1Bwu/nWn/NofQfh6g+/vc0fF5Sh3lToNA1Od6ySCBAE1F3zKpN3N
cqPtly4hwsJDeLWvoqMbi2qWTCv26LwUXmccGfZp2hUQWxPXOde9FFPAsH7NF37nzhujjllzrfJx
d9LEJl4/Da009p/k6eLJJ+iW1Ncu2OjaawMSBhAdnznrYC3xVVBKXtlMzMLi5J1zLmO8mEBcpLh5
YZOKHtJbwfk7Ca3sHIiGTDeJcXLEAvvJ1zursjVY6AmwI37qMmUOQaG792A2xZQZptOKVIq1b2gd
b95mLvkwPLP/Ei5mkp3wvhJCb0MktG7JEtsv86JBvH9faXNOm+u0Z/ybgcU6GALqrkRNBRzCObX5
IL2Mg0CL8VPru61RFMZoHwG9B4/zzVyLkCpS6fB1MtJns7ScDQjuBffjMmzbIfkWATbKLh1sHZND
cozLj7SVG5RA8Ck+H9NXYwa6YSKcBt0Izg2XI4RAbR1PP28eJB2GDUaF0cJrURV2pevUvOtNZ1on
mXD4REhBPmYBHNa0PbhvsMidHChNseuUNe+Ix7EKKs+8M0Fp2hEHD3pEA+0zLgW/VPv6BJS0EYxk
lCiqKsrEj7wGcvgq0AuvacyQaBkoCkUwsynZ3k90kjvTaqxcgmpznvka3kFc/hV3mUAA6sVT+p+v
/HRJZiMJLQZJCK6Ga87MzuxKlTn1vnIBJGCX/n0XjdMA7v9YxRepPqWD6E5OPovD/zft1BIquB0H
8yQPOyiUY+G590MLeXRZE1eeIncXDIuehXPMtiCQIMB5VjKjtl3AzVxBRigIo/Skx3Eh7nlvil8S
6Jbishx4fdQHyjGCs/KqpNk5au1fFMyRyXZnLvl4Gw/vfFG7tApIjDV0hY05TJI1+g7zi83Wspqc
F3MUuggohY+EV5IH3vU6KnMHFqCHvUnbhsx5Ta6vXyjgo1mjkx48H6X1CsYgc0giCr+JR42wlNja
tvmWbsgZ+gvK7rSReckvxKB1jiqQc16olbziVQOc3r/6ZAE6qA6mK4buHGNFNq7hNwMRVmYYV/Ae
S0BDvkjeSO6ppce4JvzFJyPOMJybDqIYgi9iIBbnWwXirg0/n1QyzS5n06zc8YRG1M8NIa5ww8Si
nhIGj1Ju+lDr/0f3xV/hXT4YfGjMc/E42uOlIMyCijD74/UYoSj5aYuot15dhO8hKDxrYlNJKy6J
Tcfwnab4qu98rD25XEDvMA41oFeHGCB4m3lDlUkgP7zMvQpB7WMi+PFE/aPOPjGEnAV61OC2Xamp
mYYOnXf9WHE5UPmkkSJzZPjz4Z3315y6ILKzMg5uY5TFDm9O6afo/kWQcZOZ2w7RQKGcnH7OmIuZ
HObXDDVUQg9yXSXX6tqUhzQDXAuZqOE3T5K6zbEfEUAHXsYFct1G7DQM8QQrPcDJTSEI+rMZGA+C
RaAssWjO02Snt3UnlOhuI0BOQJYHUyxtnlJa2Ab5/2WOJ22GmWIhlMi+NaP2RI4ySsarPO8dMk1v
MuGJhTrVrVkkN/ZWPCs0CZbwaC7CVBVjlvrQheagJ8bUaBeevQfAOJ/VnNgKLsJSp8fW4eR1Rhi6
ozz6m6QIQNJFFo3GQJkqGS3wTQ3BikBVuCzJUdjzq1uQepql2ltzQaDK7wpXJ6+TwVbsn52NRZda
LWduEX7BZDGnULruUPpydLQpd1xnZN81TEe4wjKcKXZOE7CGSxNuR5IYf3PZURZLEAwOpQp1/M5e
J1H4mSslo7aYf6Sv1pNE187zY0NTIgRTKoiDQxWiJ7JBd4EECp4FUkn1BN1Yn2j13sCbp+Ad/R9G
eyizXGbthyoYn/DsyMJ0NJHtQ3qvRcmYd3tpruO7iKIUQLzQTMl5O6lHJzlF8PUv3X7mEctXqzAt
rMnMJsj7lw/zBMHjw15NSpYrdhAe9UL3+sD7sbiELK3NNKWTyU0Rxj2oY8ZujvrTE4fFUrMKkddb
jjeA08wfOIX/4fA+zk6I2RMVUM+Vp8PJFKIgDUPxAtCVw5QKyJhha05cNjAzRPcxTM+hrVKeP4Hl
pqA1OtHSRiFOJCu6xTldE6lq9LTYiK1vEZFFe58DGzktyW9ArxDLCIa6oUnETpSLluwZHomQpPns
5Kh4gqw9SiM02qMyuTdhdF5vpLEMESAQdWdOJTymy6bTpb8df1axsHQ9pSDSV17LHKWntGcpvYbL
A7//xaW080rIA3ZpP9hEzj5YSsMhG80FWg+0k+2D71vsQPHp8tThflkthIgyE0YbehPznXrKD1J5
w2/x3g9sEs++n4tX7fCp703KcCB3JouEB+YDbcvrAF2dbQZQsF8ON5cqmW3GxNefjWsqMMBynuK3
wchHB+MMOpbCaDPBoSwXs22X60+aOF1QhY5qkjkWs1WJD/VlBig8mEj1Abry7QUPQp52xjWFYADc
LzKe7PvTk7tuqO+/cV7DLhDz2XAx0VKS9P8ywW1fOc4srPE9bCy+gURZn60l1ze4HH3RkBSY+KEl
iJ9aBkade8ia3KWHOUnz90d/RP5Rw7aJcGH4QoGN+5vMuK5KGjK7hdn8jkikU89+k5FETb+4pN/v
kTp0KZvIeFJRxS1IvHCaJgzzar3ZOOsHl1TyIDvFY0F0vAK+WU5fqO1BDgkP+dmP9RnZ5Ahyjixq
ILg0pxZjw6zZpypZpzXgdWBC7cCcAPEMxgYr4Vs5srqv5uis63jsyAWk1i291YiGaLkjR7T1KzYq
xSDzFwgb5KkMcN0fV5Zr3vFabPA4t386OErGqGHZOWbi4qYspjCRLP2OnBvRYEKEGSbHmX1vuvsM
nqe3wWN95EW7EhY6u02Rom59OtTEPQob9KRgcbrE1Kh0twUjQNQGrtTpQ+Ho8jIOjyKfkYPg7Uzg
PL5MPq6YlMWOWLGrfpGswUIQXu2MGxEpK3RJAFgfcRFIfAF40wDD+1hZRMGdV4CJNSnGOQ40so7E
I9mUKG5MjtNm6OoCxQLD7EvweiOjkd3qaEUj0bKDW98Aky8QQPlMdyR3LtOwXR9L/stcdTz4/aHk
91mZwy2TdO7iyyjvdyBW7ha/jVDhC7mTkZzcLtd6V386m00V3F98iKZv/d11H4u0r/3UX3XewLSU
yGru/Guls519Gr4finT1q+YmLhPJK66KHQRAalJo6XlOTTJJgphiym0D/+9GorfQulwym9upWv5S
BuvbWkYPTvP5BUGel3cE49JzB4S3WM87gKQ5hVZXk1KLzfUsNcMrpfMqIxH0G7dlwyMFS4GmeC3H
X5LRSYhnb9NVvwjVFhZCc/LuSnUFMFIownAJ2BYZmpPvmieGyrk6Y80bKiv29xSHCaV9at/8dD37
amqXm/jLICzKAU5+W41mC3iVc8csrFg8PxVfT7xyGyd5jqyGADi+BlPzHwPo4sG0/3arS1tdmLb2
leTk8SshgaqVKXkVlaZ0LngEc4f/9Wj0KBFeFUoqhTh1p6VAJCq9N+DNLBhorJyuB5NIqnWhJg+5
SMz2O5hxz7S/RKOAntLLHxoJ82gXC/WYBHMrkk5T5ws3+tVjZ+gXC09prPL8okuKTh2ttIruVNYw
saHdCSeHI9Rnf9GuexPz6JycgL+77YZPou6tNH3DmD1T5On/NKvarwqPDP9jjA5gOhBJq22SiCgB
m1PrJPaNIWCZQ/IEu5QonWIxAGLEoGz0le3SDh4sHuLZVAidFGoncWE2zT+9+Isytzmo7IrRWtHp
0KPsBoNftErAqzGE5uNrdnefqBamHPoWSj0n9MJkOvoVdH/eycdjoft9Dpm0y7TwwAFkPR3PjB4O
Km3zInyQ8/uHrIxr6en8RK0gkifRoZ4wi0wDbdvim9Y4kTwLX067+L+KVBVakGjh0XVqevuzPu7s
lmkD06ssaV5aoXpQ6uOoo3hT2AzqcNVsaGgA3Iwncey3RL1ncM5dCuPcEmyJ/0JqBN6Zpzm1VRaN
3YyRmEjJ+c1kFabDQu8425I1Z8PYW+FPXUzgyVFxCmnvptZD4lMdVWs1hFaUMYYvAtFcE8qLZqHI
irt0kEP2KTKemcTO0PMEuDYkftl1F6KWMapcW8iWz49wkXK2b1TgTorffp5XQWTn+qjlKVqzC47b
0gPcmqRY2JSX0X9NOm3CD1veTqXQV4Bze4k2cBggBq+cT5IxyANznsD4Rz7i6wHwtcxhDHcnT4ER
k4yYtHeatImlViApnlPgUQS8f0QHL7ldQC5F0/jnf/2Scry5X24Z4ImS1QRmUiiQT/822x57LOWB
J3HUG3vJKiz63k6RTT1nUKMqVZwnrVgmZkqyOx1EY7FyumL1+ZX0pLjFoe0yERBOr+i8UPAu+/Z5
qLMW6ld0GKUxOXuySs+8bDgyqk/7gckG9SJoC+D5Vwru6dehUXLZ2lyK6WoHZi4QErpQYDv5jgew
VvQHQaWcV9d+tqqMnkAX+fXQzKgPDIT4tuqkPlDL2HqAnrZ2aDQJxan3kOnQMvWg3qDWbCCI3Y+n
0Mabeg+w4lYosC7USYU1k3opWNBdd0x8antSu/e30P0frC+SVXtWebru9gteGRAaV+IRcvfBxmOY
sMYgrYIQR9bwOc+1BOFqHVZir/WjUxFalY+XtQR7K6VGy8HPqCSN1G+esx5h2Ftn48b1NeFKvoNc
3vX9K1FwXEP4odkQmBs7nLBqzKZiXT9Ef/nqUc5pR6MlVQEk5Gt3OEBb1d7UjOCYPyGq2+6r2zpg
CqiEg7KISZFxnQ/ePvO8YYVmFAc+IXRV8oFD6uFCklzFCUCEYeuJk0og1avFU3O5CqJ8xtqG/Z5/
PRhjnkhJ9taHMBxEYK/aucmtN4Du4qzAXEs3Jb4p90/mP6wcbqpOakwAmt5WkvXFpU/qx+98gAJ+
0BayAdrR9OJmhR1aHPSyNdQrdlNVBXvmd5szKWOfsPW1+KD7YuNwrun7glTDn3j5x80YT4pzvvUs
gV4rmjsp4QzBXfy0JdlNYt5IGEdCeBPt85rVTghdhp/N51fVfaWbfOVyjha6lmjBiFX9Z1P8Mstg
4QQkH4tA6ExwT9ZDFh13tSYr2hqV6C/nOoWqQPT15I+RLvtjtsq6IHUDsGgGl9ctZhfB/LIu3ka/
EPzf5oobeQ7AP7h0L8d3Q3qlm8FvNOYv400/OUuP96EgHolea4Ym7rJDeta+Q5LJDiY68RT5DD9H
y+oA3JTl/DPAbIEV4tD92Ie/Wx3B/6PmVOHPC/kNHsxGb01UJvIwnzRZR66xHszLm1bzm2zVDV9i
UOds2+0dsbxO0D4v5Hnu3CYu9xyc4RaghKv8g/ff7gDxyW1bs7RAEYaLcGcn+YLm7yR6XbePgsr/
kAsLveBqROCATcPG73y31nxSa1TWZfoAX/NAHMj2DGSsF+vno0kiW7WizMlOzZznOEYfGKqJIi/0
RKIY4Whj4c9Idxows3Y4DJRM8B3k4tRCuNI/9UhmmbX6IKt1k9r6u7qMEDKW+QOO4BkNc4ziT9ir
L8kwj4jWXf320bnkW+VLw6aiUsC5ZYG0s1tfdemty0Hpng9qAh34DeeksMUpLCidGP/B0dTh5NEB
1iWVsbI5H7w1kicyNrTVgUq96XfTqWYVr9ltXvrAgL8dqCa/1OYeOGY3jzt3Y9fkPmlVftqrU46W
qeva+BQ1loAgBYMmrSeElSoD1Y3nQpkYZK3k5ST57wXu+DAzLo/p33Rq9pjStK45uotD6/LsDvWL
GfMuj4KdV9kCS4MJHZU8swbw7FF5e3tEA3BxIJpCp2veIjLqpGORRkUeNrKxBAduwyHsIDecl6Kp
03ajL5XOI1vYo0Sb4PTlWj/ORs3PaWPNqwN58Mk+6EbLKgextii/Ob7eOruunYq5XOxGU+gXLwHB
fnmEguofmH39GHU1pqKXUwglV1T5j6f9yyJwXebetWcBz/KDfLR4Y9TgIW/9pppwSqx4LMy8oUeh
O0ExPe/rnqx/RlsOvJWDwTmM6uWQwOpck/FA0UVzvt54aoSxs8dzG8umXRZUc01E1Y1WzUwuWiGw
Y0bdtYpaI6VzIcpFF3DqZZj6Rd/MrPK3ieTC9pPeJQt6eOAyJyOGLTAHlS+Vt83xyiRu8b/d44S8
DJJghNbY78sPiQ+3rJgQn6XiSVc0P/ms+0si7XvYXkminWY9cw7KLQFPp6PMPjSnRSaT3nfTx+Mt
vE8JyxVTUO80fXKX06vaILMGA1DR+SdfFKC0iex1AUkU5XG/pTOVkqS7QRJ0BcmPXiiFDIMwvuGI
ZRBJkabpA08FFM5BWabr74w5QNYs9rr2psFBUaQtODSjNUlsRHK+VJS0ErBtLJ3gv2zZpwBnWNxA
2280jR9J9JjZ5RuNT6Rhn+YBkxLlmC9rUFGmVadJCGmxmSCMoriwQxXTgNxV7I34+HKNWnhojGoN
Ez6equeWPViWkYAOV/31BrTSSSqHFD5271Gfleen0VNG6MJfk3QrUbNpqiDZhaDUiFuloTQNaKwf
DhWeiOq1dw7Zao+Dj8KGjBJ3yjCSr+/aazFZgSo4OWdOU07+sUIfvh8XAHlbAzfdh+zlvmoYs/wG
rwRur8LSa5zOANVOBf91bvYr9qqzcLCy9EQx1k5GZ2mKwnfk4nYq/xzYAim5deyLGdXrMJdiUASl
BHkmUjYSX/uOZCoqXxG1qUN4EXjcVrSxW82kn6yrHT//4UQpb1m48rEEaZueeihhaLw201oputzf
0efgx2bQmXB26gpHSYU1cICQAU4M9fBDTZW/SJbJGPLZii1w0sULTVvHK54U5jWNEyWA3grfbI6A
I/+ozVFm2y4vlTINLZ/sYYQWq5yx1umZ3S9JwQZM+lJCNKAXPnXtZEJ6KaaZpH0tSRyS1iUz89Kh
xjPNjIjaGFhmKS9+oK8203JkJ1hYOzl5CNzsBcrpCVDwI8QRi7BZa8KPcE2HwDvPom3CsbN0XGUp
MoMc+YsGWAGF09qfgXcJ1bXo/aiwC/91pGVbIp09NB/dZTdy4Nvn63dgTp3y9fUZQxCLmDK1qbAQ
boRwIrPrOQl6I2529f1RGgVDvKnmH1tqR++UHUmnJHUHylQ75JTA99SdvcWlyP6jUj/WnfHEd4tF
UZV3s6etYcLyqCK70xxw/dkoKmFoHDK+LK6Ynh4vqQpPcGE40b/KF5HYk4hc+hWFr1niG73Q8yU2
roCpYqRioLGZNE1XHVDDfMbTFm6jvTVJbE9byzNtos2hBtBXWxJwF1QFQAtm0XY7tsdWo2hs+4Zt
sC3Md9TP7A/Pe/coGEpmucdn2/5hh85sDW5Y0YxuN8hUC/SF9anIFWR/cj2fgeudNkyMIV5+Ivy0
nBP1emLliimrwCy3S7oqh7LcXPW0nxb97bV1ZolcZj4UwboocttG2jMKDGIHXL19QN54o7bnRaHH
F+Prq/uC66KTZBMpDUEbcNf25USkru/VHXgsa+HOv8j9qSpuKu6o7h5rZzREZB+4JiVlajan7pBC
Obrk+poa6K8lHNJ1iQv+YJ3esv4iBcaQ1ZJdf2f2/36MO/uY3+8ddgZLgvQSVR44yv5qbTtkBAQr
VUnoy04LhuGsCGGganf8ZZfvfNiDrA7IR4lHMO1ifrx/Ow/74SurQiCCNfGs8+VgKNUDeEm5GhMo
8hYGz5/jOIi21bwfDSpzowmoZR4Pn3mtE48QwkTwDvIsGWX1KkjyAtpQ9JVHzNhcHHO8HlEjJ3Eu
QX3YveCVLcoAgZy5SjNEkPCHwRZxWbdm1cpc/AgzXBYz7ULf6T6WWV8qK26eHi1sH8yeAhM8HQNf
3X2KztCKW5rORWxrOgI52qrn2XXw3qB8b4rNx6lP9rsVikLus8htwabZKLq+r8htR0FU3A5TEWZh
kThoEcG6mDPMbAfQbtbcZiyxOWyLnZ32/8rOL/JmeWncSnZX7Rzj9DSEMcx6HaTxyqilVUqIHjeC
kC3Dp8irpnyvn3+iFOBu8K0o0AXKi2j9toO341Gu4YNniT6vJuz1ur7vUCdIBEeRNLSWpCtZALSu
UwWZ72ba2znRVN9Sq+p370Ritn0A4oA30PK5iNxPkqCJ/VztnBVgaKCLbkYr/DBZtUDxfC62kbv2
Cfx9U5fYbpQtuqxVGZfuaV6aIlLWVq5eOORuuo1cDDPgkVE6kldHGkh9f5TuKTl8yPjQ9W+qIIBl
B726UdjAxkLjjDsAyWqZd4qIsNr+cofo8SguMy8ES0Xk+sMEkeyBDkAc//8aay3xdKLv2yJSk5Ti
x6p5ZaYx+cQFtRn43KtnThJGPzKt4UjD21nia5sJE93nc3GBPA216mAntbqZHJgKFfss3Up21nD6
4ugCUWna4+hJ1uDSYIOU9TfybemS2gXRrD3VkhszDOfkOP6xsQwORJwXFQ0/AHimZ0ExoPpea9GF
C5Z2q5M9yhGFhe0nb8eeUzIQNpwJPfiNudY+YkUfYt/oeREkoGvZvDpMIcIXkcsO1YNueTKvfNh1
3oyjXdXBj5n9Dm61ijEW0q1Ce+EaeBYc4n77oWCRbSDf5vB8YUSpt/b5irSI6hUieApS2pxJSrsz
Kwnq65K3s42m6EFF7VX0ETLtEL9lmsgnwOXOp51bpU8errVlfthMwhDYmJFqD2++IBO1sJyiG7Q6
KDanOrkJiDkIsqSVCeLxYTPEeFWWpHdpl3gYbDQNZv0p65nUmEuO7LRzGGhRzkFZMFwI/KTUqIXc
+k3lmTm92OvKTe0Oklj9x54V0I+/HZ6eik6a/ghh1QBsdKuJyFYAdHMob+D8Y1nRBcKcW8HBOn34
tYrqsx6mO7g+oI/4GzMQulKLV5RV7+rgluAFJRvRRy1srwy4q7NP9azvvilhhMMKljY3uwFD6DHz
VOq6FOq5ddwCathjomHXPzGR/q5woY5QSasHFTWzD70WeLMK14xNPjnlKjlgrt5U/nx0A7jZxMVS
gLUOMH8e56XGFrmBIUTC7Em8hLNosVxQjdnwXGqjpoHmzEMmfqQUXg6Iw+iFEtIA7uxshTIcXGcP
LksVbg/Gv1c6hIQee/jY+f8XY75dXihTC02N0QYTUf+ovZGA8WWvNguLf+4LYubHXWG521u179EZ
TYwgDRvaj0b9BC5YsEhT1WocBkaUAwkXU7hh6uB47psgruY7L/alo8X1KJqGsMjB+F9B5MTeglcV
f+ebJEcUreb2fJEKTYnsfG6vhZMsT5mbanJGXzuayz9qfT3DzObTl10snE0NlrECWkM765RxKGZk
aPrieAYJrIAJtaBUWb+dxOY8CvmPDdGWWewNtoMtqeb7TenvojRqqfMSzCBcLUTZKuUv3UUEr3Am
EZiJNYt+6HRD/DnZgtLsWti1Z4E7IK2EbNRBSAnq9O8FtgXiqAo0pqyNB11RSWjov+mQC2TpxNhu
smmPsHQ9n30ILenJyk9YwOl9S9+tfle7AGFPYKIMFqF9k04eF+PjSfTSOyV56Y5CCT8hpPoBnxsx
nQNUdeuaQauuF0SzbsroG9GqrsH4LpxoRCS7QPmoPARaMZAC9O2c6c3lPszgcew5BBvCfBG7K3DU
DJAknIFw7Z/SIG3Dqwh6BIr95OTaORAiN+d6QvmvK1AoetgLj7sKrkZQC5q1uLSh0EWbFZk2YKf6
v+4KJOA5NqKopj8kZ5TnE/Q4ckN8vLNORnVei3ysqPO2uwjS3wLkcbLPaaU9I8I1gf0+Z8PrERok
tGpMFFLV08Dwu/inHtSnXPfm7qmROohAxT6nLML2JIZQqjPrcvkg90dta/T+CziLN6WGpRUtuAd4
dIjkpiyzXPP5HUAtr3uPfyxveB4AxhPV7xhJVXJ81TyQ1GI5UJ9EWvgSBse/g/tOG9KaXPWT7zSO
PpOVYWb57TIyCCJhHIcHx6JQZDFZTYLlAmaa6VtNqG/rQAFMhyth/rcZSPKIJurqolTsuOq7uIO/
RTFEYr/593KnkZrS9uwL0sW3+wz8yJxpcver2wmZzeRvDp+WCT0lVgITgvw3XSEcm+cv5R3bzHmr
u119QkFHDH8H6kIM+vVfXyOl9nzvP9Ry8tmeecLmQswUVbIFu7N+OeLE8OdYLH2jtPdJUryyHhnh
icMpGXXMZVPu8KWmizCJ31VPG0xfW8q3faIofrtNvE4cQE3BZDusyXnsWXpXljgz4DIx0tLlKGNw
OW/0Y6pUCOkZyeSBMnM6kubgrYkjdsUScY9f4ZmMl2kN8PbNfGteSiIFtk8kP+7RtHpjanFs9lJd
1epYYHSEzdcCMKbEBmWcTmNdweiyyIbXHGJLfNbwbttgVNaXqVLdGc4GHKMst6GV4UqfDHJSTAI+
E34/4SBmHCXVtIvv/oXMLm9a4RgiT9VGfyDJ9BAqkw086IWWwv1oilg8D1agFZuAWnNi5dWthNGF
DQrh9XKtiy0NKsyKLojQjsrt0YJ55ye4MjyNdDZSUYFKqJg55HSD2bDoQackCIhqTuiGeXIX3vOl
Y8V6067MIz6iy1a+SCUGv3ZfNZllML81yxJ4x7Vlcd8WMKozgL61RXTqewoouG32MSOvgWNLgtVt
7f7WSp93ciPnViK7OyOYzMFbLmFrMRUjmZQYQLkcepSnru/lIbnA84mp297nLUq0NQpIN1NX5SM4
bfsoi/Q93kvWCbfO+J31Lugevyu+Qxqam60XowXYw0BWvnME1kvApm17q9g9qpMgecta98hcR3zp
sQQBew2uiqIVXhNWyU0BSnAuTexQc5f1cTD5LflA7WQWGEAGFJJNwYCYOnQVFbDWpHvp3+ljEjSY
7+h2rT0qYDedPLZYKXcE/IaoWxuWXzLcv+AoRDS0TcMejVKDx/ypFaAm58TAjsJ5z1J6iifQfqv6
qyjIBxDm9+G9RzJLkrLhYK9Ph0xfAhVcK6m5LAX0F4TzZiV7zoQJAA4aRrTAcLSunURc1UbCPV3H
CNvS73Rx5R0A5fG/zilndHxymT/XLIYowQJnWl0jl3elEWqPqp2RS6PsIf0noAn8hXyWyk4r0vgB
VUrkfMrMpNijKsEaeO0iechQTgM3Fts1m0ELCTcfWLw5zOWQkppuyqH41+t3lQxwJe/LIeaQxEhX
7IajIyv3D9jELrwJlnDuTiYTSFHUSW1Un7Yn0duf/HOvxxQxssS97UMPeYt1w5l0Z67PZxGY+QOx
j4nx70RGI3qtHxq1Nfic9Ojy32VhcwtBkbHl11QpDlIDGGEuN7ks5vRxxU++7/qor79cOYMzR/Ge
E+tDiaVR8dnUs1uo8eY8uynyMvGyiVzJ0iZMt3uVPDEBKzKI/LGCmg6Zzod48MYeF9ESJCQjaEpZ
3NCY7ZVrRhxznsrR25ACPNicIDIpotz1DQxEuUBPQzl2o0QDanqi6bfL0s0jBrzv/LPXDGUKn0BL
b5VBw0VxIxyDMS+fMapJKvZCi38Hsznc9KsnbmKX0nIpeuoFoqhV0+NRJVPCHytKdWg4Nn5x9tGL
73G7IdsO0XJGF6tZRLhZqEh9+rbSr5gWHZHOJEr6stTcrp8X/aQhtuY8tLwGjFMmXQFZlpk+bhB+
a68kZ5Q6yB2Rh7Pa6o+5sVVOGA7V1u/VzD0g6t9O8tYlWjKo0p+wwbeLpOJuj/3zLRiY4RFuXKwH
T3NqY1zctYkCjxa1vurUQW70We+bilbDm/loR1bNETHT40m27lJ1+QT3PSfTarOOwDKl14IzADp0
1Rfcs0MlgZffDzKcdxUxyr8yJaU66DkodnFrjBzLwONPdNMQaYithY2oUMTt2LsGVILql5b8728i
WPZtDVuv8UyyOUv5TUXBoYRU8PTSX/TLNJlJyDr3cExrJ2PxkKDEZ/C0UsKtW6roqSTsADllGN+M
L58gH9VKIG5frCL5GqURYfSmbSYSR3O0V+nDzOqYKuhhhFW92f3kMBCE1cbXotN6/Wr4R9dS/0hV
gyUTz4h94M4cegVxZykyqoGuWd7vNY/g7Yg8g/a1FfBmHsjUrAwarMnV1UbJoITzZ8QitVqzvFzV
bjD4XAOaQzNntIJFbf/c+YGxHtFaQEDm17jzY1BvU6g4xGIIh8pMmgLFwSFrxqD/KB6rJA5JIe8L
nAvi1EzAV2oUwVPAdU1dXrJQVCRsgJqwLMnsUvW03D1MwvlonSWLdVPvgR1l/3Sm2U5qlVOC9L3R
wt2eP4tfwdtT/9G1kupDTzAXLg5KDDbqeIpdQLIxwPb9EJL2piWk+3yPQLvk0E95E1CixDfkxabi
TcY4GrmQll4trZBLJYBibDhMlJG4XuITlevTODMRQ2LruKFEXgPe6yHqUNd1bKFpZmgg8qA6KffP
5h2ulXFX7+RT67Gs9yP+78GNKH9sRRmQdld6iu2oQd5PjC6HPAdwsEJ5zLArWIhBSJjGjGovyr3Q
Gvbk/uHJ+jQ8Fa1mHVqEmqInLLGbYYgRuzr1zM/6wbPyREpyk9Htxm28I3bQtnyZaygTF3bQ2aIA
egKJtxRP8aSYKVj1ylDhXVBEzOOdUzIcim/g9fl0FBEWOtMCLSavxNf5UQQnfekxVOhCDassIuc7
KshDNwSUuHNgqrVuDLSbK9KHiM0SdZqzOtgWaiHQxVRJt3M7So6fE7U+1DfkU/H5UscSb08vFtcW
M5l0gx7Ls41hQc7/gZ6zB7/i9QYbaNAjSIm2TgyfaajVr+MAIpMhro3u8mmptaqkzjJhuIHqGT6H
nc1RE6U/F32mFiKzZDIOFejWtC4xjKnVLJltvL9xofZKfe+H4Jqx+CXnY53wheSae8lb3l/gERv5
Z7a4b6HHHbcg5kNoPaSWaOElJYmw4JgB5j/9v2s6bNWZCpqmQ+6535Vf096V6Mnj4Llq8bsZOblW
KYbDIk+IG6qM0mw+817zO8E3bQoXpFtuPvieX/os41N+0bYyfuDoxFCpbv/fYo5gJaBlJXghH11k
w1h8I2a43yC78rF/U/qgW5GweuQFl9k14xpTvnb1gbaEMavhe37acJdhA9DCJri66zynbaqECtUl
3MD71BsHngKCXtVZvSI7/T5fCF48LHWF4YDfIrr6H5z1FDh4+idiFfKRX9Oz1sv8FON6whNAt61w
De2PMCJP4mKMN7rBS955lXgcYb/GVJ61cRwKQn/HqiRY8VJwIHSX1zY6pBL+WUvvDVjD3tYdRE7K
l/Ueh8KfLdvEuF4p1t7Fk9hCZROxCvT3kbLvEZiFEpwb8uTitVwQXUZrMOv49Q64tBhPnsrge0tg
twe9maTKbFhiuzJKBcnOBlNm0q3wMR+Iq6sT8yx1VDDZ+KkO2cSYONEs+PCMJF71Lxmi7BYC0YXn
+FBZMMJomnkgjulAfJYA9UwN04tufibMAUfGx2hF6Zh3K9CZuGlL+DsaAMogQv01mPlRqTB+3ETK
7Z2wGgCOPto56QWWdyIxufYwIzwwcCDTPvTnv8rK/Mlg7I5vcNdNwm5Hp6oFjy4MNmaoab8L6Cp0
L2qQMf4VspExr4zRavlNNaj9ksNBMjD/icVtHvnJdkvxPwHlVJayAg9b7u7kAseMj2rtBuMvJAFS
X37beuLfuI1J4Xs9I/mq8q2G3aCP3fPZT57rueE7giPptvbf7ib0lehsEYxb07i2elK+YSjhxGjm
KSuovrVcbGdquAoQ/WxM+zjkvvO4V5mhJINhR0nCO+kpOhul3oRTrq37+15rAD5ATjWBbwNHaw6C
TJzXukmmUQYnkuHmU78JkMzEwJfNCbUY7Oihk4OrK1aP4VDeyQmmVGzIopnTsnIQFbzG5KiymcYs
fbfIUjfW1eAyebDJDPUA2WVMj58UkElMVSKz1Nrl59OC5CUAbb7bgdiyL//Fwq9jf5JHIrII4NlL
oVTu0lXaNMpJH6mu+8FUsx0Jiwb+CzhdlgbqOu5t15/LhgT9MIV4Ld6MjAiXjy3YwOT/cM1HeT1J
hwVPM9brVns2TL4Tq6OwUMl4gXBNStZ7cD3juQkb57usQRRb64R7up1orLGpvhItpTZf2vUyx/gQ
hhHQD+t43UMIzxBHTR78UXFLWARqFQ3BhDZJdmBYcNk+WXybuh2wpdhgH42rBDBBg7kNRCMzmweI
143LydkvyFlWnw9W/queVGbLRcY/N5GXO1wJ3dck4mlaPFDMtkkiAkXTSfNOTXi5R4iRV9a5U6B0
+llF9DaPjOuCUUMSZHkwOK47A91xoOgq235+9DgQNFBDW7DhdU1vVi509Q2KIHMPS5nlK+mzHSAN
X0y+DaHxlkgeNsC+CBO88u8S9zKDB9CZaeJQaK5kCLEIoXftvYfAlfkm+DM9KMctYypVsA7rn/s+
Z40+6U8aBw37sB35e8YF2Fw1wegldKeDYS22wYZKZZJwSXToYJq3ZhohsrLaVVt+lj121RDp5dpz
OI3imlJVqNewSzzklbIc9BI37IEB6QT6HoKfpq2XeD5sxEUufC+Wbb214A5g4lvFOzdoJyPJazB4
fXgQIaxl7rudYF9zaXn6TnnQfScAotqQOrB1aexNmYZyv/uW7yyINrOUd3jhOjoViUoCcWJDIvD3
ddWM3aDEDzhz1ce6GnUnzGTk9TWUGeH10GNsAf9TWjNCM8LigcLHZqqhyYpvYIYsoYHKoTzgnHzv
rxnS8TTQzybeutApm4shoncuFJUzBT1AB4HTbBK6l3/XKfLqHKda8GlOG+nIUf+dEZC063PYaO3k
TlnOw2kVxwxTP2XsPJjDdPVP7DbTLn9M8pD8fxNoDzV/deveEQk/wYPkrpviNWSNR0yevqIrA5oo
BLTvi2OjOAYd1R1IxRRREuyGnID4hTnvAjggA2rX1+kw6rPcgZrCe6uZRRJDivX4IaHx7EJzdfY6
Ls6vncCCvtmQ0HDqbeDX80WFHcaaFQ+e/4I5vzS7oOJ1oYRBB0S3mj8Cekt0xg4ziOQLSPVQ//Ya
QlLrvivSGOo+AbzZgQqQ1lRVeDKidB9qScYAjfRjHP6bHMY1wYPWqP2a0aCdvBImCjWNDUEwzjCU
GMQKekEcLsDZg4gpqCjFfQXV5I0b5Y4F2NiWGj24qsycTw3vAHgqpBeicgzI64Njs+D6hWU28ivh
lUoicKenWZkpsmO2Av/dtGSH+8WWEefD3hWNSy2P62rTxuXQJ9QOnlGO7teak+uhCw9W6shAI2n4
2oj+0V7CfmceFBlxi3VpRJre1iZjhMvci89lBpyktYBI89lrJ2JUunhpGIjlL/kd+aqwYto9ziFy
dMZxb0L2fv2FciymLgsN5LNNnAbgknqgDCe+uJKFM3Z6PX/K0WyzdBVPzPcoMedlvJGiO4yiYrcO
xjhiM6MRrciDJ1h9Yutyc9rkQhksveWJ56bCpHowx4MLYE+FDm71BxcZqZBE7/scuHueCQBw278N
ip1MzUKTiKc4C4oqstgAarAtpPgcGGYLW0bRNuz0xV7hC3BXjldHqw5/L3oSGkmbp2HHt4GeAXab
rsAJ07T5rcuTo6VI50I4uMEkAKtn4coSpUtDXwlj2lk0wFAlaFJL1REmBVMmhSfilc/6345KI5Vn
ZvwyrHyB+8mle1RdRxwo9ozyuad/PfzhmM/b8p3MT+CNmO+9+XLPRoBXJN2YW3xiSI4sof3RB2iH
BrIFgKgmvuRE+tz0Tuybg/GKi87Q3eqdcGlJhnysd8/UCEQppa7NEVyVoLhSg7GLRyaCZlg6UWyo
1RdktDijb3nVrAIfyLp0zcm4t8eqoVktgumipssnw2A4j/1+T9uwVaiWZyYr2N4IfV6feeegNhJj
HCYm6Gpc+D+ybGKB60uCZTvUheunEQSHYyNAuDhC9xM+Xs3VqPI+NMvh/GyFW9HIRhdaWrmU3arZ
00klWhgYrO+ZsGoN1vfwofOV5qSauPK7Ay1zDY6Lu/zqwuFkNZUo+q94IlHfeTYHI/GMlg0F/rVx
avSVzp69K7vy3x6HomOJwh9a5grquBfLZwxRMr/wY2LsUcbPlQZXdW/eRlFK2y5eaHYwJTFa1GGN
m3VLjo4hQwaYV5hCFPreegIUbTswO1+aRoGCqooUTw7PG5/CfofCaKmsbP4c/kfD4XR+nYdyJROl
g/pP5qMsQ0n4HPeXObcTdXYi5yu7vTt/BHkmQRW4Dr/aAqg3Ar2eqCfxy3u4+lxx88YI8fTkncBD
8mldWEQYCNcTBJBSeFls/vja6H9pCFTQ43oZ6WyL91WHdRF6kZoJQDtZeIHBAE2zvGGxGmXVLQHN
bDtesnBxNF70AAVJnhXzhMj29/akbs315cveoue3zZoZGGYKsEITt1vKDWg+RhXM57Iqt3B98USQ
RbcT+L0b2ZTS/kwoeIt7j/xu+AjeHTwj4bhBGmWeSqvHsT5yXgenuhg9IAiayHEMgoLpDli/Gz69
HzaqoQz9c0NVvhPx/5+A/OvFyT7/fdM6Z7jou64tZurzlgh47Dp11jpldseaCJCJuE9Lme69xNJg
E4TIsmHieJLDhNKXIiAOcZbmkkuBqVgFogxdLLZdco5oSOKTdXG6vWDLKNMlWTRQ5ewtZ01Iu6KS
Hun/FZ39WTE8gY6p87rHCMaCwptk56hwxs32Az7FZjQCJvdMLrKcZ+P1T8GcDJNArGabTvjXcj1U
GNcJiWp5aaEHVZGOSB2NyLPGBKKnFNq/rQ88tAgIPLLN4LZhmhBYoC11bOmDJfR3WrkA1IPmdUre
vOZeH4PoJkoZGb7yzrSmjjTHXduf56yCXzGF70Sydrd/9fZXfm6Qf4pSwx9EC+r7PoZ6j7twjWPS
gtibTLxgXJqY8IFYhe95/ZlrW3fU6mI0FxH4RUMVjjbmBqmiubVfv1Ufcw2pJnYHw167aLZLNeTF
2v15NjX1fcfNpQZmD8+zaxpZ9Gw49i0DY754mO532489PUJbowMpzpCL6alQipnXu/wWuw9Wlvud
IpxNGeDmzAQfKglRVg+AsRIfPlswbj6bbILgEYmZvaCFE+I1PFWIRlYoB/3vxLny6nJXLag5L72m
Uq6f3UO3hfZPVKJeOJGDcKDATXcS5MBIpdvKSHlKJwAUqLH2UvHO/rsO84d288qSr2/R+RDcWPyb
9yi9QY5shkPVxiYx2lvM7iL6L5KC8MkdMHrul4FTOFnznqzz7pqcM7h1GeGCl23p2Hl/hbPzG/IL
ECgISA0A2VQveypqr22wIOiBB6zeDQwNtQRC4+Mv6bNhc28CwH4/k/Y6JUHnawc20H1Z+ShONX8N
UgcL489PQSFtEU8IDTiKf/31nJRNz6PYEoytsMwDs8JBkORw2MofShmBdI0K0A2rsFEmw+jKezgz
GC8GJp2Ij2/FYnJ0vRu1dL1g3ZSrekLmX/orMkpTUgZilz8BD8wZEfItu1yAqCmqNKN9+7bmV0cE
HIpcnhvK9IlSUPmh2mQwPipBsLPriDJkDFs91lWofhb2yEzkypsCoyV2qsmgdl7O8y5zyJ35ZNGW
Coyg8F6SYU7M17Izi1k/TUXwrON5f7T35bEN13wfKc7gtcSPfWRNFQM06edOsBtNPO+kQnzDCwhi
46E60FEc9lPtOeqiWz19YZvtKTy1D9oyNVOyL1HikcnM2Fm1E+bycJJxmtL4Zw9svcBzGhvbQuui
vht+vueT7gjL3puSIjEosNM8ondc2K3D0EjwqMegZVXSpjMK7CJI6sYA/S85e6khKeJULxaos+B1
EKWGf3FUnUR+3QhnEj9DW5ng9cenk3q1/A1Gvzr0VvtIHz3jcctxVfgMpTK5605dtstF57bjaOki
53gruA8HMmcgWsrP4zvUMp63OyYR2e601ZxNvsIAR/u7hajUJdobbHOclR87PpB4cmOgr42OGFs8
Epzh9NkA/3bHb3/XFVnD596gOMDZ42RixleyCSCxA510gKt0U0mLdr2lWtQ85AyjgYyr7pJ1tFQy
iUIE0es67jYuy5RAZMWZutJPery0kO5RbfDlU7we73BXrYYq1+MuuNjxCXzbOpD4M4U5KDrBqKPx
aF0rQl/8/WBB1sFup0nAAw6LLDqSg8Wp8yeNo2Al5ywKj1K63wvOt28p4OuP5nIxeQjO49Qd+x5E
fXkz6wP5tfB2GwoMK4x4ZLa6CplyGrHlkSBQBtKRGtAcyh4fe+B+RQZ59As3WXnxToBqqVqCS3St
EZ+2rmgVNp2ANHey79tiXqvzbnbtML1xXk1xHEo5sy1LQGiEDM8R2aThy9ujOuK6rvqhC/FNw+pu
PxDHtbM/eaWWIHyAy4j9MhTfBTRnpPz4hHfSqa/VY84gbi2GoanhnF0VJWVApBpfI3Dkih49iRSJ
89c6ZDIHkjFPGJTQ4dkQEgyqWdaEzUexpAMBpaEB5z+4j5pI0SbrOvpMJOSZmIBKPc47/NlIpG4w
u79OWe10zy7TpzXCVKbMLD0TemA22Sh4U2pWACYL9gvJILhvm4bSm7PhO/eaNS7ADNUywABwiTR7
C7pXnarn7I/uV8gxk9GdAZEUyskf48/9vEvzY+zwaJeGQ7dgcbLEp0/NXPo4td4YMQbvLjKPLjC5
z8e5Yry/gU2kU3mGElS0QAbRu3d5OjUw/RAWD1NkIrfPL7+dclWLthBR+P7jjTHt/k8lBTaExN5A
Oe8f2h045n9LH6sYra7/OQjXfqV8sWjXz97XPVLt+jGcTv/GQnqwgH9x4cdoV9MwR2HfbB/PLJlA
/ZNrnnnjcTWpZtte1auX4olNrFqKQLV6VPl7fOz5rU7ubYGch8a23jGn4phGcKSmrBWN/hclnvAm
HAa/SRaouBSJWv85GhwJMne+6p7GXEKprsPBZWL9mJPNZh/jokhR4cFPejCJrKNzjFrTBQucFKXm
il79OsEhU38DpOsOHhm9+xa+269GZjdJ/fz7eCNdWz9cb/0lG2+rtXfZiwpMZ3iIecvtVUipp9fb
RXhOpdbxV1roeD4gZjx41tF7sSgGPMFwp8G7m864q+0wHFqDdAV2kaVsJoBI4SuO6BHuUR4RFXw7
bqg1rIapjzEcp51nQ2SxqYO7eL2wiDCNWumjzMZI3018dSc+4+YXFFmWW30D12tgBvGN8QJWou+5
oF/2bEUcH9ltIhogS62ZSOwiF9XMp/w+s6oIycnL7ALB5Kc3rE9JQ2Dg2C+97cOeX3Ob4m/Osr+Z
DPJzR4RCwEDCS7b+LYHy6CMcQxV/KiQQkBCD7WC8myREAJ58NXncoUGsi1ilGDVhNFwlWgYexOcG
F4VmjX/H1xPMruaciEZmIwLSR4+/v/H3hoWRxkJ69/vTxWoi8GKvm4yxPhXHU60jorgNtpVb+yKF
HKcp1tT4uvvm/A7hrTCVgXJxYl+I8SSTFIvPZVZ0VK1xDs70Bg0prQMA9VVkkojzRRYTiHg2AAwq
0MmMdF6auv6+q4Pk5qlNiKKmskwf6ncFpibCoXgGC26SCsarvgyn67j1012EZpvlk7gwm2nl6IRN
yrTYJ3K3u4BGBgAtK0btDLhZLv6BU71QImXf38IZtS51aUqsIElnsukyQJ8c8gymvIPF84tBpKE3
kmLwRSmrd94qslds/SU1JW9M9rUzXzA74WvuBZccfdcN7FiqvqAQE85h9SofRYa/GUsxqEVf6UZO
IlYhWNJ0ygcVeKdSCqnaN7EjmabLFsirHNJ/+Vef2uHuEdLXTCqodS56SCBxJ7OTQiC1H/y1jz+y
gd/824JBypcomnKj4nyhjJx+sgLdyZx7tKA2DSJ7ZO6570yMzk9yQPfsP1KBIogjq6jay1gMBSFf
aiCvwdjAhdSQZRBE3BI8SfR2xik/FwXP0dW9lj3u16aogtvd0NEAePEwnXcUbGbGcihzvXwXKQj3
sGNqESgoeI6w2DuvEoasH3OcR/RRtIejMAQdIpWDDrwtH0bgRWMOpO0UQHw1iFt9Y2Q73asR3xjx
wxiNBJpMXkHhufrfcb1a9gI+TnxhpLTkOX/LdrENVloZ90quOTV5ZpjILmIJ1T8woc3uAVvRr18H
Z2ZL8YUjm2vLF2QGe4p09mAhdV9/+2eSajf3SJfsnHeAXFclWPFssj3BuG6ks6d2t0ZL2cGo0w2V
nR/zXxV/JU9RHq9NkNHnAFSCFL/rOfi8+WACZeZJS2D8kC1NEtAUuh37EA025KbeySUvH+mEKbhq
NeM2CaYgJEJ0taVFAVh/5cvs9TJlCfIyyMq211OAn5Ib2ZyrivC9KEZIW+7pTozK0jso0M0/Mmjn
DeenvIAXWPvdV+zq+CYl9cap+mtN5uQBPJsNkRc3wuJXr9MCxQHrsxWV4aZi/kMWR6E+ECC6yGkM
0qUSO6oELMuf9YEMx4Ui9FuyZByjUS13eJVL+4UmAz9zemBHm6+006uJa/3dMa4+vnKO/Qs5tEDM
J2v7b7Vea82xxLM4rgvV9CHndrD85Q0clk7QhDEOkYJYWIyfDxqJTLdiScTXAEE7nxx5c5p9w7s5
oyz7NwY8EjlufQo7bSFpbSJgKyzG1DElXAtQPYhSwlBKFvU2lEITvPvur2B0WRNZweaeSI3tl+ys
ACbCJRrF5Eja6P4gaxSWkmpV1TxwQyA24AiDJdvisGC6xBM/mfMgFIeY6Iqzhqm+yPI1oySI8am5
vi0nk2ZNsswMc5HEHcMV66xFFFfacIlNlSx7FO2cg2oyGhCSy2VX0+ZYrsJ4Y1oouVHnQfj3cYgD
0xSect/jFdbUQz47e1jTN+Ysdw5Wv9CVcbqw6I6Y7gFPdNGLAppQRXtebat8m74FAvP2aMrWRciu
oEeC8NHdc7TJHML64OF4DeyLgtmegclis6c4FIh3szKGXmzCixz/Bzz0E0biuZNKmTwSJYNnCzE5
Xvrk108SOFrJhPXeCwbJYbJIjl3JTMnw7AJPrzdwiA93m5PjWpZSkqyzGEtHYyvyxPJFLeFcu3ea
YIdk/J3bbN8Bnl+DwKHaTJjIUYQx+mlnOX6mlXR/IxjoFLBoRrQYM+E1DeJl7B5UI5t2s+aMTih2
crvZx8DGtcq0w7uR05oYI4+5F9FEhm4i0QlmgV3HIMqcddlWBozc/R/tEIj1NJ/7w6ryrshxGAAV
2M0t0xRqCutA75JgTJy70WHF8mTmYyjrBr8wVpnca/cgOGkF/9ZZhwoZNeDqT5qnbRMsXfYSYRxM
c0c/DtC3WZcUhSDYRIQaExpX6R1P4xWTr54KjH9pNPgJ41uWYGZ0g8/tjMTMxkG7MWQWg+TdxUQL
+rrMPdc5cIhAgjFEmm1ClmSCJ+iJi3oQ5HttEEPrhLFxe4/Hs2X4FhsySJnOyOyyup4tGpL9hyKF
zlqXlOwBGd7w1ODKTZhNR7DwzJM36HIp/4YHilbbIyuIICm2ohQ1xYRtDoFwHYGA4qsc9a8Neosz
Dol7VyFLdq+zcQWrL6nncMesJNS32PU0LwFxD11KsIGoVxsT6BnAHS4hYdKwF/oMpBeCbCMpIm6Z
aQMYuumFIk8HVwJ/4alRw55DPBKqwI65pF+4p3pVOZS0BCq9Lzwh07GpjYSxshiECirn+1l7fqHx
UhFgxWT/O1x65Pr4x0vDX1q5entZqHo3uFaFC+2ouw6VQc5CsiG0Q1+QEASvaf2x5bekeCOZpN/P
2+/0HB7263X3jxYqWZl+TAYA9S95xjQ+9xplBGojWcztoRcdDXJElZ+OHq1eA66nha4GLog0W4YH
JQgMQVMfjpwcND/txcE4zTgqOSGhZnoOiGtKjVvCSYZX28T6oI4CdI3Tdb/Gekym5PkOVKVCl7cL
YPiH+EQyrBlA8UgSSykwLFBpSZrJG8+oMRjIMxvly3rRORu99/DYkLy0yzdTIaszFsePGa41BVOy
N9k9ZYE0KDDvAb0/ToLJEJBddx8hGPDMWkojtmE7YQz/gstICns8BPF1Z6mL2rfPZtQ7sDfJ8rxw
fr1Dks1ZRj7taJfCaHOJRWUYy6sdb75ZCOkA2s/S12+lfvfxXQc5jbXXFLm/XMpbWeHEIbO2fYdE
4N/nj40oPdn+QxWNuq9nRimP/2/2tStan/TwiFM5RHwYWt5bosE2wJ26E9E4zfE+k7kEqVztYqPl
nnHF1+9Mqpf38McXbUPFGU5TLK0ZAFtKgNGw/miyxzcbQJfDRrr3uSyGgidPQHNSYaAbQZ+2azn8
ZW4YuOmcyXlz8Ci1aCXqzIFspSTwGLW+XDaQu801OYNfwLCHQlUmo5Mhf0A6GOBZzPpR1NdSP+9/
15bwhNz4UbXvNZYBzCf+G4tSgafiLU92k6/EmFvUy7HnCSP4EMl3JAxMv6FLLrzMnVep5Jv3f8qp
yp+UXk/00SbnMXwzo425RG1dt/kOHAz/iywxJKNUYfQR/9djyDadf5bjjTqIiqVQ7CiigXyV4JX6
WNO6cils843RIDIFueH8SynI7Q/VHwh8EHBy2jpD4YRZQQ9JnUAGkT27jWTLhjogZXeJdx41j4cl
oqA2Mvy/wdxbR+9XVPIew6ngthSE2O94jMaO0jiCV1+o0X+RBPsxusAOgThDvqsC12ci6OcAUlSz
AN8QUXdwW9k8wgtkyN18b/iMF9AMBr+qZjN/DNl314OkrB0xTNKhV21WZs7X7COEZBQBr3+Ame75
MAMmzQRpoQeKN7wxO48smTLHw7qyeIvCcz++22+2PsM4VyPa+X5X/rLky+K0uz/nU6+nT/nyyYlZ
BYnUpUKdtMm6DtFhP2Oh289jzGEpYywHqulmJkkTtp2y4O72KuL5thf1CXijvWi5atJbxv7xb78h
AkjsnkDLWi4FvFXDaJHEtXdyodyvqbEdg5N36kUTSv33Btg0zBq3K6bnksJXRl+7QpspU1OAuwUr
5iaF8agBdEPJnnE0Cqg2GZCZkDahnJNy4rqsfj4AmUho+QwDXwQO0RedtEx5L7sOAiMn7FBRi8Ns
2Q59+LgsdXsVxCVLKPaQPZxA2ydN9fAJk3Ts95dawnaSNTSFpRC72SorHryTbZ0+oTyIRPTd2Il7
a5alECu3zDqe+TQjKkTSvLbsNR1tIjhPG9erm7Gx+fuBdDPwswdzQmA/AAH9OSZkrEFu36NiZ1LG
aloowV9cWeJ9jlCGS8Scs3Lq/zbOcCGyzUfm+A38YL18W5ex9REsByjC2pyagHRnWr6zLjbcbbVQ
zePr6frAfFV67V842Th6AK3JJ39B9OtFRqO6zALOsZYOUjlDAwCobmpay1htvQDtv6JdT3XGB+u4
ekO+SAOqa7Q1gIXbVxjo4YrZSgVKrJcbPxjGeb+ZIbah+bomxPhUHTPkOaSQx+qMfnerDNOi/Q9M
ed0cTn2bbkxg+4vR8VtyAGn3gOm3b9cfyj9p3zqmnoIHeCLg6nilqUzMnKBf9Caw/nZ6vEMEORKu
2Rtd8leTRz9tatAfitQMx0LMkHzMzD+V6dZSaltqq1vyfNEnYpBi6fLFYJZdqXe94EBTloOw7YVO
dLXzslB35Z+dLfUBdJevWaYCfhTiGqn7bV1u0qt1iSZf1ghcCPiTHXUD7oIHmeGIWqLQ02qs7DcX
vMBd6Ba7DyF02sBqQ/sYULU3PnCRRg6BUSCYreQSCs/h0/dpKgj35Q8lXWQCawmmCKPubg5TQoCp
Vmo6Lx9E3Wn6RQvDzYmwBDziQNn9ftwmDHYMI+7yD8eERgu/NxueCgpKEJiUhmig6+lgCFfZ4q+a
Zw06mhNY7RBTkNwL21uVLnJ1pLTH3eCBZyUWUap4Z0eIgunapqXQC0pkeqwFcn5bH4ObpVTOqaih
zSjVZI17l6gIxqO3cSbopsaIbtHiGWUDsw/b8AeDmNoF2J46fs+NaCe/T7iAkq5vbvMBgTlXBQGF
MsMJlLNO3kk6vtuUBcNqxVdq21PLFDtIZ662rNKpbRo1vqXAszgBu/94oyWfillMS4x6BKR3Adi2
wJebCIW/+uVw+3zu/BwJ5E0sQvaE9yqv6yAIh/FRd8vCs2i6XhTd1ecssorW/SvBf9lUCnFuRZm9
qm38jqvqczSjmnIrKCv+zjK7G993asQtp5+ngsqFoJ1jf42VsXq7x4ENog09WN3NomWj/pEAqk0x
JXoVkqqrrkYD0uTQAgCZ00AzhStQ/OADYqMJuYbd9WsHJcWM3xDdAhR10cOLq6ouGclo/k0vGozC
KHqpVPsVcSHRboCRRj7qTUSj2yeuHDYZbkau4WwSB+REclcqhfcGYK8ciDI/JfPs2FG0u5LXbRjY
KpKdFRjWILd1NZIi4d/lnDpmpQ6Bx7PBrT6tO+NbYBnYsJESnafWEQ9xgzSR3Fbjx0Xl+FRRsRyc
VKysSqHV+ZeSl4X1V8RsVA6SvdEHsKdqtZn1vf23DUO6JzczLi9L4BjsQlZlK9cCy57MaYEZs6qq
1O8XwuI3QP9w7bDS/9g0VKKvhm4hWHfZf9Vb3y6LMYMu8gIZbYtmdM2nTC22fC+pdn89qhn9A3J9
HgQ5UDksz/zFukEXW2Ci8kf5/VgKuQQQrFhenda+hByWItVaxooESgKAvZJEsBQ1JCAhqnct8u97
1YZIo4AqIJy7uHaLvR3eV1JH+fxRaq7v8FOMhR7Mm48TGd1aHdnHYifmtndDXOX3ObgR4ieyzldJ
jxA05XWp76h5bsOwRdVj171p1BFZFTIi5uP7K7yPhy8HHa3zPW8LefU4ZADgSnfXNaWqp7/3L0C7
74VbbLnXGJQlK3SqBKlwNrRBm8LSCG2Gyqs9l1yw5xy8RGNFreW3y51qokp1JZN3XSyEqR4rRfCZ
TeaBy4OsdwqD6LXsomk+guMzOUVWOhTkJ+VmTxBJu8zctuCw07Fj/Hp1lNWfbdxPSlzyaWd3QMST
CmgMscKx8NbKLnMW9OdH5Zg+piMkWQRfJOpS7p2UrenVoPV+JLuQBqGa+HpgSHttP9WLElxGHZW0
O4dF5uYAgykOKLKxOieu/4vNq3HJmXaXGzmaD/FX35O7LbsfpupU99W7qJZeRq3YRiSewdL3gFpe
/DC+xMfabXKvHY1eYaHbk0x7S8RWuhlTJFkB2/CDIMNqdB3sZHJTu7fN8Mp6ULDujwP4PxrQ7Hf4
6akcdg+45vsdHn1wdcigH5lLkzCVtfbMjyz8gum8neCkeXKl05fZLVDm2yKfMcJD0zHZHpBuUva7
irWcpI4wQK7pKh9al7BBP0B0H+r7aZRSFKtnH1vW+LT2iTGsjevvZOu34hc0zbp95KwLagorovxs
tGofPG6/yPAT319Jwp891QEdUn5l6Xr83QAzcyKpfpvqW7DLDk7SmvY/2ObksI8cEd79quMFDVOm
f8DMPWg+/jJD3MPfRxPtwnLZ7P6eMCpetJk57s4SBhxKkHzOOZI94hIsEHW+hvcV0uLLeNVvSkmP
0j04prUmtjtlDr3kIffu2HVA865CHBS8jA1bcwSjFZwmd7YftiZsru94XY2Adf8zwH40N3ENqzm0
jOz6eldiHrZvkd0UU7FvBHiow5vUVaREL+ssGKoToM8/b8UEUqp/+nPWyQ/T5n9pytAyZEKSc1Ss
kIOpxDiRQcpnrFOjHujNH5a19mJ3M6FLznWf3s91XhRT26SlDAZwXheyQisNxt5tbJmyDhnvJ9zu
ACHyFmlqxL/JFxAnG5ba2Ii7lUfwKeyZiWeMQ12u2bcysNhaqXoR2YWlOA5ORcxU6PWhtuyo7FIu
cxTleS0PYaATuGPvorXI18rtNlsQPVuHA3Y+vzScMiHVGHs41aP2m7dnbIREizLVeeJtm/TRCnma
KlLxulZA2/bUwsKOt9fAbXRsDxo6UsQIjQBXNY21AVNAaQMW44ruokMpuaAXh+u02p2v9KznYJJJ
7czwyqtiDvioBbteiPy5BKOoC5U6fQjAp3xT6GGlGBBqa3SUjujOLuoCTART8Lbr6Xtj3exM9udd
HaRhYVwwhuu7t1hOWrCS/+kcIGG9i8eYbg1pn5BvtDUO28FDLKIu53JOSL5H9CCcftn8IdUF5yGV
1kvZKo3AdC0P1UY34WrTKRkvVXa9L4201nrVWUH3KAL2XYvQZF2v3NDUQD9c+Y3c6OfgWT1OEm00
juQ19Wn2CSvr99EZUEQOMlMDhTg4Pb2VWxMStfckBqhNgLLEWBa2Ipaw9VUAFoNBi77/o+bcsPTy
kBUV33Uqvt8kfpK5EWkLwYef6+GxMbv7/D0m/QZsfQ6xFsBMzcWPMEqBByGvIoj5/xiTZwDvMhN7
PE4v5ZIirpsHXtvBnmM/BddeWdeMCtwKBbiaKDxIkdHFInAqW46k+LG5g73SuJv53pUes3YaAFLw
KMHftPGFtDF3/u1XEubUfi5zJSFZaHi2mz3zuk+IXeNIEAR/VsEsFz1Nv36oN77ioHmM71DGdG0U
+WGJvHrRsVs57UlsPLyV0bwN73cPKkAI9yF4aTeRqbQO4gLWIEyF6SaLU1q/clOkjfmaUr1A+pDL
qZe7GItmMVNxmzzIl88e2v2bOO8ClIaePa+fnj820uBPrsCTrdLG16LtRmgTjdqGfbOIimXnApwv
qMV6mE9haIQ/MU63cdMan6eByXEKjGz0eZgRA1bDG4EULy61O2jAsBjAYTq7LZJNQSQ6YOT5e3uM
IwvY8IyM4cBB5n00ZOuYu07ryIrcCb00S/mcvhLmipaY6pWoTAfW8yxY5sn1FPto3FgqGHWmPjju
z1zxryqOZr3y1pJp0uak4yCruTMdGEwkUbypHXhzMLZR1xPZMF85yfwBc0Pu1qkdJbksd6wGXLe+
XKtrwSm6sh13ZN70+nNzvbvKGXYzoqbXo4hOkObQ8+Sx5uU8Wcw0ywwnsTSPlOXyarhgMr2K/WVY
RtTniViKkd+BZed2qm0wRRprO+hYL028G73KgirXRlbdKQ8u+wkoMZnlX8yoiNaT5Szy9qSkAnGZ
olBPxG5jEXC4gLQo1ARMmKi0cZDtsM/SEGcjBbxQNGaVj9nF2UcCK730uTBrfnM4LeL+lw2XrFG7
gJPDmqXgDG3T3dmdCxlFckn/fuG/S0KpyJqf/XxmvSGNxhqNs+B2lpWbVjfHq1xjEwdatWKEu2M6
NjTR2/K88gq3CwryIB0Cxpfqlk9ZxRuZtFFAl/oPBQhKVbQj6zc1md5DYflAv8dXkyOttoNa+9NN
zYaDAphInVWR5Lkdh8neh5Gmr+RuDLGUcWbocqqXCuv8MW9eviVx8g3Ge759p0vxAnxhc+xTEa2g
pV5pRx9PtU3/CMagFZi+jQU0hgsoQpF/2E8P+AmQRHRac7ccMtYI3VWU3TWMrwx2KWWgiZuqL/Il
B3UOi7qdK+U1Q6M6lozm2xFRTath8lmFyrbJrOWb6lrThTUO6VfwOXUGuna2jfDksL3pKJCuwunM
t0t8s82RILekN6XYqy3l1bDFH3cTMz5ZdIC/JCH6EuPwxZnWUaOzmXUqlE/qHEOi+EzkQGIUIymB
YA3HcQYcZYqQA5GhU5Y1vY6RgWsxUNt3/vksRQzVvbA0/uVS8MCgAyaOWc6+MoPaotMvAs4uJk3J
QGlftzKmjVEFycVoQJgbjkF3earBh5ov32vMtFieAbGyZTSge1rJqlNAwfE/vm+6aVdGE4UiPTdW
OCxV4m+ZDMkHuQ41P7KIBwa/BlKkumEwLjC3VN3bMXIdUi7l9NwJULTpAPNVBSM/jB0EJ+ISpR8b
3KM8z/JEDdvRqTGgGU3DtXl9Mx+iS5u6s3Gq2U9SMcmq+NFtmB4ImCzdqjQxM1zQpaCIOfe1PWlb
F8whjQWPaSuJ3YDuYFXAAwJxi4BvSwIrsp4PXtiapNYoU4I16l/AEZes7zllwt+0VdCjoCMze4kV
zDYYyG3xkywzZRxqW+90pbEsvzq/xEd9/ru22WfQpd2PZ/1Rwzbg0aizyMSN3lD41PSfMV7T7pBR
1LHVmoU3sagHthXSr31Z2yIJxLMhYK+AFAzDm+yOCQEu/7NmIFjcduHc2airt+9AwODFY6Jnf5Uz
rY9DyRqTHJR80Ljj4ESmgxsBTWxMkNu5Rnm3xamLPM5PqAI28gJTWWrTbC6xiFAdHJsK32MEfCV3
J7qacQZScBku3CDIbGjhr5ua3V6TjhhZcyHOnEzuYOWjYQ3yH6YP7VKMf1B/Vk590cac6EzLRzjX
5yWrrSC6WgxK+lxHsOBH14Sxsf6gz8EDDLKngLroklYyvtmdDKqDEWXkREWFdCQYjZgAWOgKKS+G
agDkQWbDXPi4Md7559V6bxkylrbIfySwRqunH/zK+LtZdMzgYJ2jQzRCGOpdpkwPZ4cC/5mlTTm7
JgBSrwVVjzfAhDn8sZ8pNvhkQyDwrYdAr8r/I8Y9Assag7BV7sS5LYyMjLAFwTozAnPspYT4fQyi
mBDfEQYJFuuwbkPNjl+g7AsuxsPg30RcXUie83s1KSv1T+gPNVF/AvL61BsYuOMF/2PEZdPxWl5w
rJYlk9iUSD4jAW/Pb/4m+oT1uDtLSL2fSgV83FhmT63KJtUEtMagoZtGYrmPPLQpL6C3SckH6oDq
vWKJG+/QcZFVmXz9OckWf/Kx0lAKxe3R86DfndIugrVcVUOWNDu8J+6yVEO19g46ndgnmgRKC8jz
cJJXwmFMxRt9ldB6Gs598j9K0Mbghsl1BmOzLpEeTaXWRhBN9u3NiHE5J+WGA/fjzuAKbtTip6Wz
alTisWWd97Gr7ribZCGyaqj0Qz4yAK/FblXqPPKq4jUZywaTnVFRwHt8UaqtNNwctYVUABYh1maJ
wmH2k+Q13fD0o264eDU6zWgLVY7QhDwW374rA3B0Wodq7pIqnbnovMJkHNP4KStXFIJ2nI2xRfZX
N5R0RqcHd2jWJZkdz3uc1Ix+Of1dnkCv/e7L3a2Q0Jt+Pq1gDe4RkjjWMfBJS4Y3fYJzlbnB5+c0
q1JnMXqtQO2KT7izzsv15Mp9a6S1645+T9hbEdsS2w9Mm8IkYvhO/WaAQlF8m5KIi0h1dA99gAmj
cm5kmhDjGrtl6H5jBTzcRIBM2/hPWL/v+hJfyDk55tiS3ghvKiGPG8IQi9xEq+ymZ7XxZ3hIIiBV
grN6UbDnozC6wHwjTdwts1kytjPBWcCsk6ZI3LQTYZTvqsbxeshgNReX46Gqcih79V3pNYCC9M1u
18cxYlDLicnO3PuY3n+hP6TrLRcdvX1XQE0My8DifVNXCcVI6+MZ6YkzAY415+N6yUd74BPUbrbW
w4/Z6tXqZYHmF9/rH77VlUIyPutuuKAgmm303HJfwZm31df97nHGyQGJag7VDLM+LjuEKdIcfAda
jsLwmqabsERLqejTZ8apSeVcdrw7ugaYcAdEFv1N5twkW9qldtNeAhTAbDLQ2u1fLUmAA3FB7wLo
pkSj2/Wfr9S9FevwWdIv93K0V2YXT/Vh7hndWXIKHDGlgT8iLKYT7mzkcBHeiBOIY+s0kZKmmjnJ
jziXFsLBTamri7k8tazKenx4ZvqOzfcVTn8sUJrN8UIWp7nbTj5yxAkf+7cwyRyQUXn2+sCPZexP
JdFqWZJqpR4jximBMOr+v8leMJMFYPqF9tR2l6NwBew3Tp+BO+ZEtp7Uk8Pq02nhokauz4fgRFtO
gIG2g97ggT3e5FZSC6i2kd12g+ZY2ifdb5zMIWB6AXt8liCj2O33Kargh/Za2RO3JbuYtGWIKxpd
l5HwrtwHhuRSdYOc6GCZ7BjaLeikr0KGuwR9ELkPEigEw4DoOvOH2cjjXR0sY7tBCMdvPktAnNaG
cIUEGv0I07izbfFeAE/3q5ADWBhJTv4ZPwNYMy0gK8ME66aZSddu7zlM+WdiAuQ7/0qRbkdsB490
6uML9dqG2l+RSiRuUR6hKkFRV+eki/knvWM3XWh1r85rDT1XRw3UVS5UAPCY7nHx1gvou2KVPBtC
YtOB2Tk8Cv8s4haHzu0OGbF0UdUw6+8HIJr8ITwFfOku+36GRWkxO4mG6P6FUdmrT0aLc2hyx1L/
KEZF8JJzybR9wrsawIhvYDFMP5sjIJ6V8ynb6s5S5yREf6Tb4U21rf1SJNVR3dUfzNQ/2zHLkQ3X
6zNKy9P1dLE3y+hDy4dd/ZCr52AUPNXSB9UwnngLvbAOVY5l7R/10x/L++Yf1QxCs6WXTxn+jcUF
0E8lGGXuQ3xCmhNetRuLlmsDg95iXA5ISt4J2uVvzF9iHTXXOK2Tabddm9uReAnf2i8bHqrKr7Lj
T95tOOiC686t+9N4HXFcLgTMKb38Y3eKwA46JmeqVkEcNIaBQ/GYdTRZmEHicegSjlFyT4wWZSyK
gU6Z3fzjjxsbjaPs4/9TV9hpPU13tmBOY46+9Zny8oW8/ysOiG9RKHAN7SmpP659YdP+df3ZNru1
T9tY61c5I5pg+BP4PTMp/S7p9KkVmwjZyjcRlLjmtT9VAJtqtd8tBLIADKFG6kP00oT1lid+3vVn
8QyfpZDcl2OOVkNJSMMxu4/TH3DQm9bRnpbwBlRgyuWOlWdt6wJ2bV51UdpSATc60XX9jM+43GHm
uG/U1g6eQfRcabOCdEA0e1jHqtS6l49+6j86C3rZSfCncT16k9qCmW41LM5ntJEzsZKiJTnHj4RI
bsmp/t4TXfYw+PWkBzRJKtDbF9ZKtybZkB7k5PW8LjWw1MeP0as9ZCkYeyyvnIaONPlUV4JAmui5
5Cm9ruiOD/mdrIaNZj7Y50K5gE/L5DbQheseMHethRoCQPhdoKw7gmjEGaUE+rHooqrnSss9Cv2G
ithVqBh6D41ILxSii//ZoTzEMz1TqAF0gL0CbdvmZCSLx3sDzCxUvmkFkzltHFI35NwAkgkk6N7X
gVppRbzG2iyeoUPwwhgK7/086UlRb218qVtileisNqDWrU9lbuE08GEbwDwaBMWIfy+3i7C9kom8
lX3KPoOpc3UzcUobQ/TcatW1EcT2Vv1Nc7Lt1iCdK+f6FymoXi1hCXGjb7l94/PI8eQNNeumJwcp
WcMVUxxR8L4UqtAaacYpu65oK9VS1yHdamCLZEk32TaFDO26nHPnsXfh49ircPURqU/HqI9ZqsLY
GpOkYabJNQ/W0BvVh+nVA4yFRmYagzKoFD+oDeGpc6kiP2J+p9QupfeIU2z033WlWrFj6Oph4cgR
SHgC++BgvwiTjcF7En5AqcGOcUymW57w3kl/UCb6FnsZkrjQqynkwer2FHt5MqEt4VAGDEbUTsHW
2IHkVq2jAiXv1OVKYcLyoW9aJYNI4ojIU3N9KOrCzJjZORUN/cjcCs9n+w3a3PqGJQZvMv16HkuX
GObYuWylXuTZaWsgXDB4Syu40Z3AHezhhadz2UWmxI9GAxPrjo3QU3nsg2KPA2dqm+QhVULW9UEa
lpogz2qr5dH2v+b1lOcdMtAGXs+DYtZ75Ws4sUuhn/wIK0q9DFNV0aWocfLu2F2b+F9xSVpTA1Dm
5lzT2ReQWl2kqkBaDL/g0uzdnB+8/3s8kE5lHKOjVYfOj2icGWhO1SLi+mHuMWY91bZjUz5xI1Kz
ml/m32a5VGCElUuh8NkstwGNLpKdfVMcti/nv80Btv3BjDwZSCDfNBhjAYWKua3pBm2LtE3mXD0C
PK2WNxbA0vRG9zfntNgBjawNrbSDedOCba4+CG6Ts9Aihs9GqFscp9mQq2UAbWthyyAwSP9oUYRJ
vkb8AniCoh1L24YwOURTN1A5udpJizp84pnKadOtWkbMu4QYFFZIF4WG7fzLY01JZRHneBwkadhI
5FMNNv5WRwnc0KbUSUrUHuzvzBjVfgrYREzql2HibKqoxgrdypCVNl6+M6RqwPgFCx/CFXSFlzfz
oH9+zilLPYsFbGXuA7pvH/UbZS0Cgp4tmpJDax1homduqEgcgmHqzxnd3QlMv7wQNdUzOmazw5n1
ZJiyyf/jvWT9PpR4BIQUAqBiBmteofGbBgBalxQd2mWMxqNvFTh0CAhn8+B87Q+Md/gQDabxilJk
W5S6H3+1O26sbHqaFAsJ1iB1+flYgTVPDYIdGbT29amkQVunEaR9X7UBESfeTVSspJ2IGzlSyCz5
1LEDXSkpIjEVfA4TsuCQkKin6FCEwTJC/o/B7hwIdK00aadEPihH5uzN3JQ5J5hULbjjrIlwzzYj
2L3seZBv7Fq6fe4rUC78+4PyhMlsp77LyIXWxCPHmNxFSRAb3UmuGdD8XYFWdgBmUFBKA8Gzmyb1
txfCu79B74AUMaOTcLcZBYWZO9r5i4IuiJpIWXkWtuXNijAJgVDouMmRCrrjPcDUetNK1s6ul6Iy
Ap/39KK7DyrI8FhyrDYreXlM3esf1JpIAVUen8O2qz6cua247UOIwHCHQ0l3zQysOnhBc47okSW7
T6EoGMY0mPNUi+bfMW4yZVByK54B+Sje7K0PYQgPeR9gckAoPonnfUQTVOUdSlPFZ7RglrkFtFkS
3k6iYas74b/8yb+/1tiMSMwgg7o4nh3z8OYFXbOu3UaXhkshab6heBMRCib4x6pVRZRdf0z9GTE0
c8IDGQA9UGoiANBkORiG+kvehiuuy/5ETEeb/w+ZChebbbRRlRWmEiZuYVKvFWWSrmnI8kTZ236l
4F7f2zrUTi3010dGBWVe0xHWehJawe6Wisxa6G/0TyohciBJhb1J1yUU7Tpvb8bbpyz9gFAzXuUA
belmH+bjw1ODv9yTN55iThmx0jiBTCx6bcxcEAP8hgJEd7dgz27XZsdy42/+fiM/GCRtdaH3NnSB
hS0H9HgdEXwca2itGo0FcfDBGFIoMAjvMPqxO8Luths8FYPF/Yd9rRPk4nlFcSIWk0ENeXrCdoqx
wqB7nggk18MdjAyiSCZHtXajkYgHLG8j05YhOLpjmQphpwlvbclXOr8FGOJMqiyKzCAGWQhSLwoP
2vFQhZ5goqJkAC25OX65wWFiwUTYQg41x6tpWoeqgMGniXAgsTcACJwRylnBDV0QpQircPtIxELJ
AZ03aGvGgneeQUmi/aP6JKIbVNgNTWcFyDSRVW9Ku+vOFEGX39dS/cmGQOlZONm7U0CxZpocmr+i
8x6lMkZVDX6YqcOexqsEAwvflDDUZFwQ97tGiG3jZz7EWOp5A5gQ3+HqW7wNPH2ESMOMULdluheO
A9wjuXnUM/DPVRHWb3aPj+vWexqAqLetKbSEfVoFzkjiYpo6pqEkxKd70r8v0TYzFgyon+eqrxfF
VIF04pdq9HqeV/e0aXH7pXQ/9EI56W9rekdI3RyZybdUK1fKV0i1BaWI9ofPlxdR04zCfiWexdvH
jSMRv7VfmLgWs0YSf/2gv00My52+TyTVBXO7+g+bJrQiyDIH7oFBcltexIg8OAvy6J0kH/5hCop0
zIJ1SizOGW0ocb4JWG7j8ZiOs+vuPNZfgMogeaqdLM8XPwxBDI0f9nV78q/deivm+T/2ROp29yLw
+x+L/b7tf3OMXOzGLDJO7491OQCeGLRNIij2DAy4/dVuCYbIhDyvcaO+KBdtoQqeEyjDY+sN2Tid
Q4Nd6GKMJQCoq3vDP3OJyQn8lMz+i37zUBKap7z7AlUmWwVDp/JUVUPJoG/bPRFGu82GnZP+NGYD
ykxTpzbBDpG766pPmdwAfYxW/i9PaalCH1YTJBb7G91CqAiTbizrluJWDrn1b87NUxkDZHjXhZAV
4pUOy3b6vX57RJipUrelArGUC6M83hgmLzn0hakDSb1XUZerGDydQ8lcaSRxc0RlhDxBs3AUb9oL
SKEBFT6jpv6/36ur9fdpSgowtizp+BiaUXbkuYmlFFPDQ5Tb0EppaFsCWX+sWY7eRqWI50C/Eb8V
Xway/BxgeqXj6I2xD98LNrX580Ydcl6a8/AUTv1FT0VinKJQYopq1FUgJYH36q7VHwnrGZfPIBCV
GTratwA6K+1ePqazEUUkzwNQP4IkikyK/kUq3T5ZtEMlgbKHKG3K5jgWdGfEAlMkzW78/nwT/cdL
t2qd3+IzRbneoMhIyL3oQPpWYV/znW+dpScyL0A431ZBwD28Y5YFSXHc4mfUvef5sXJTFE+0Gphn
rruPyUaDLQWY+w9JlUOOC9fgAacZoXa1dzcdqEN5Zx6Y5TX5mJF+Jf3hJpxB2BTVz/tKQ/O+6/wo
mNvNtavCikSluNiiIF/BMF+MjF62a1rOL7vIUaPVP+QGz6U7wErifZ+J8CmFXiCM+KwuhA85TlU0
RzaT+zKVZ6dWfTYx9BBue6jBZS2gScfWuHuIlZMzNv0bW6KAjqzTTpNc3uE9wEeusoUd2kBlrb69
UqiFyM3lKAp+wWRTA2xcEH5AzSmwf54CcT1pzkYMHTDbh0xnYL/79BSC4atwh13pi7TbvzxuqQFj
BFgRNrXsENnrwJkC5bjDPLfLVLtPrdB7FkwyL1+dFTToVvLhW7mTd23LhPbzGDjZ3UpLUUcQ4Srr
Jqpxiv5zIuc3TNBElTEXtPOtykzBdIrLQabk4TqMFHgxqVLfGs2RZ2hASi/XIUr06oAlQ0aI5jkt
rZBlNT/KXXGYo/4EUEfZHLiKX4iYFvhrwQgdIl7SUoHqS4kZVyJewcvqYxzmLUrjW03nyfECFbOf
oTK/5T+/s3nMYUx1lC4oYyk0qu+DaOE5tVbfW8IKx2ytcDDcw3Hl21j0eVZgYRwkaMansNMI4CfS
W9yL6hWSSItrD9GQ+Jf0Z6nkS7nRMKQwwpRGTRsx3jo/F0imTT1oCtpXzCKCyqoQszcaA/QE5i3F
gOGSX/B/ud1FZCBsjhwGeWXmYS5JjJ5HQ6U6oxyc4OiWOwNJco06xJAcE3yntSaFJHRwnzZd9H4L
3bVPXVda1MlaeZ5cp0tOfcEORXhODv5ktTnDHD3+P06+hSa17BhjkDNq7IK9o6IbvPO/9gKNFrkL
080bRXDKt8jg2AALtqCpdERGajKCPWPYL6/nijoTkEX2dmOlT2dhTSHL5dzQ9+CEqBwmOi8/uAWn
zUXYi86OWrRngmOY5LYaiEqUm1XZGUwUX3k8ivYwg8ZuXMk6L9MItdjSKQb89q9uZPa7YtWiHJki
Kqaw0pU+QkSWNNBwJ8TvTTdtiyknamTrTgUCJyKC7hAkuL1xuwraN54JUV2bSsffAfEgFywvBY6+
xrH2SQNp3jk3ZGUWLbbun71YDsHEUbvXQZ9dXBDrjU3fzpvNCr39ruD69QGyysml/nrwR48lm//W
voPaYkqQS5jZNg0mkeUFobFpGtUsMmeAfQzVNe1w2werQye4S9nFKb8GY6WaFwIZBCD1jGRftdqC
N0Msj7OWMDlY1DSzAsgWajluXZxxnIFf5SCD2SrYo9VmV4+lHmRjZ8Jht78mUMppu71/kqWGn31M
IIzJvoffLFNc1zDpKmCLQHY+985LhZQRWjQ3SZKAg9v+UOL48Uy8Lg5xAbz3ovMkDc7oS6AJMFdM
clgFJGy1QhjvsThD82ssM1pH68CgpH+KCROs+BkO/4UzrDgdseFo8IlXxgNZkuqnc9MEN/UvPe2B
zZyHI+tGWU8Ccp14bXYaYfz3HFP6XyBX8A0cP1NMCF0Hr8cYhgiPXuTjFzlLFSkXEtok0SU5HYnY
gO2pXZR9XAthyLKhasP0qaY0kYMSjzDPvijUWFJJ3hHYzEytSQIhRNfDbgJdCTBxJuBsPNH/ojRe
nyN+SE3V2kIJuMfhrKGbLsRCL4O1lKUNjODEHnnkgCjxAROAOS+stTzziTZuyMKo7nu7DbSFC5m7
zHjL65rot5JIDzK1hUcZiTz+SGpjqLCxaceJASf9g+f6O2i7QXS6utuq9ghNcp2jCbnuPbe1lLcr
5qFzA5d5qNEsS+QYWktBELpdel9Cvo7DBwtD8F3iickzct3XlowB05uFmrD9kyf1b6iTTmu5jl5Z
IutujTcCKR/lIEUKOh/wNi+OHj3q4eQbhM5mwdk47HL+vAjjgeN8zYzWLSP1lTBTXeI5c1Z1kw9x
Qp3Am2YIxiqwHT31PiSnTWev+fIz6sgBHQMdCSW+JunWkaalcBl5e9vmqdrQpNx6wyPl670eaVE2
RTN3RhSVu5+gAmFtwfAEc7cfeO8SngfkhBoJzyi2alzQbBEteKGCCtyqOK0xaTvJONESP1VRWYZx
G7E3psUI2oAbTTgDfgU8OLl0W1pnXMbkDWFyEAZb61Nn5aTjsHQmHyyyLw4cTSQjNS3x4mmcWSix
7MP/9+tP4hsIRYWSthl95ILeBDgvukMjsd11PA3EEDmVMqofGpon7jvzbxJGQkWqnPv2OqXrcB0p
uuozZyjzLa0USB2/GG3LfHO3wslW79qn2oW3MapJw8F4/eWrH2qdd11ELn9BwBMiYcwAk91M47hJ
f8yvd35wRWAv5+feJ1BXuP3SNbkNfQtOJvUj1e8q3wXgASz9fVCg07a2XrFtm0R/ThZJvEdNpdD4
BIP8MZGrNmd4izES8VTmvOn0uLT5+CavoyA8g7NBiTDugEZXa/lh4yDpxKoBnb8Bedurmk01WgxX
VizlQkTvgBCph7bDVREdLaLMcEwT09QOGlrCeEUmRP1MPwUla3J7pNyjdWVibhUkBUClJjcV/mMe
xcoNC9DOqaNG+7ExYhuv5qn16o8RfoSjLSC4tbieHf9wMDhE5JoWq7rFA3U6wCcrxWRJuGNg1qhE
6CFmKMsxQNOzI9Dt4sTsAbimS/FSwbIcKC8Y1vhb0xsxVFlM2skYkn4wW38td5j3le8ifTLKuIO+
ha3PcqeMvblXSEUSk8G9pExtXIUxP4YGToLc98AXFRwhb6bGgQKQwcfgw2i9cQIDKk0u+xe5X49F
6xcS71/hRkHvOiDHdB8z4QmSYcknJaa3MUXt3ywKGOujmH/OGTbfqC+MvbpqF6X0A3qNHT8RHg4H
YM7b9z4kXPJ+5TecfOEYGqKIYGfUzLsRghzXcRSObtQ2I7A/idYDW6WFMKOTToDbXEq5zIQBXKb7
erEEe/2VB3211NyhutZfskR4aiYcAt3mAHrh85MU2BfQrhJzF69rNXy3Ptn6XDJ8m0NZkbaBDQvS
D19ie+c3emOgcspWenq02dhwJLCMVWj3jFzLCdmarymI9ddjctvCq4BzqwMmSQr355/x6R6knqdF
fUMbRpes5p6sKHk1moTZXJLbs5x1bMhKpkd3hDyLagQuUdQAV3fqKpQvaK8gsChSSkqzZnwJAaJS
MOLeM9Cz55UCRPhIOf0rB/cuIz00mrUgWAKcPx3ik6SlMYU+dySW8fdcbq1yWXIPA6Q79YKczNy4
duxbseOxtzOrcQWwI4bHE6Sfeei0UBo0KhArpHIXnwwQml+DRZPW+8THrs/C5AmnjApmScMLuqBd
9AVu4/aaLA3aaT6TEu2wxCfueSpzx/k3T3Ppq8c2BVqUcCFtOBIjVKuCNAV4maclCFBjhNtH920B
NS3WdD4qf+wP9hphlx2v/j9fAnBNSYDUI5yG2hy/WMSoS2rvoRYIDEPFrpfRkktFBrNUp/zgYK7H
UNCFo008Cg4uT56i0yC1PpUlqR48XDQxI99I+LjRYg4f8dFPwdDGiyNn5Z9XiwRzpCt+OnTDwXmj
h0hXBHbPGJMLphunblrXE6FI5udr8l/iubxzk18VuoLAjvnz29GPZMEpAocdoDTBC7BMhmra62nz
5bLiRkJOspreZDYGrLQnSQZpncrx6Nh8lIevMX2bSfA6oDkeMRkbF2DIxaAq1TugjdlZfP3TgsZM
FfmqeYG+XN7KsU8/C+sC08izzC0rDGC4z5VFyNdBBvV4hUPUNQhjWlCwfeDhxa9mRnteXTpYOvtx
fXUzkb2iqSDOW1C9omNUuqDfD+ntNcFOIkNOBaSmBKnEaX0WjxAdYtT7ZJeHEEn8uKcqeoDFRkbO
PCNRkXBBQVj1tMYnq3EpcjJ2UPZd9tb6gP0AQ7By94cCFWbey2X2InHOeBCs/Z1NYr8nT6rP7NQM
PtglF/Un0VEi9JVcvFQp42tofFdKaG47A2gls7sDmmY4FCy2Pqm0kjW5dO9iKP9Sej7BwuqXB0bB
NQDRRRFgjwRxPxvbsBmAFbgqSFVY7u1SCrinDPURcDtdwM3blJiXVo87bMF2qfL3VoL7gd87DEVB
O487RpKUO7rgA5HaO2S8SMb6gzc/X7pbCP3FSIb2glXmA9NITZ2knoKRx18lQADF9CltR3MnEkOP
tOQVdmI9vlCsCdANwZekCLH3KUgrznv0s3mayI2MtiwAZsyXoJVUUWYcwfflVRY9Mza6Eg+iyc+I
7EcDYB3t1ADRarN4PhtL8q5yZrf15OUxPxth5Yy9eXuPO568n3RGL3yHMWr6IdifBWx8yEt/amFX
sgwQhrii9ZIgARqGlUPe11S5foKWHf1q/QCqzQrduf9q5lhSxfOsL+1Gu9O1gdZOiVmu8bPR6d6W
Fxj3hOGNCRPR89mAf8szSGqL97UfMtTKG/xR2GKbHfVf05F8wtNOMxCtFF7F8PdH3T0cuL9weMfU
hpz12qfHUUe2l+kdPputhJzI0K86FjR1zwyYDKRXOeVmi4PPTuP4BBpNkr+LHBAD3hC+FumPolgQ
t9nQ0t/yexEJmrsARJOA4VO3Pse9IpCh6FL4yAQhuJME+sbicsTzomNNkIDePNTl2dchwglzr6Er
1xPqUi2K0zBewzZyuUPIpY/BRwXgGLvHIActnA+MVuEhSTgFo3vEILjslnL/zUuhTg8be6VWiktZ
Nx2C16mzADIOpzBF33Vyynw96oz0sRRTZIaT1Il6fwIcClvapQ66tbFuQ6MsBEX++y8G9Rqt+n6r
LaT4wVRsGa1kEtFHMPd66fMSZFBjL+1U6Iq+Wm6kfueGCuvRBDGunxqBg2vUbMt+HzPpSVnqJZN+
7Yt9zgTVONJCsoigT7lZZ+QXtNDTGPBvhQW8ZQOgK8zabV2BTDVyCap0TRRVRhA71vbrk6WrDV19
QlTEcRhV+KwpD+xuGddJi06VdsV4Gvhwnbn73XiHPlSq29TYYzY6iGqC58QjHI0MStZkC+1PWKBN
SAVE/YXShDkKlhKVe0XR4ZPz60Z6Nwur2CCF6ij9gshQgqEfhF/r3t7mm6FMJhB4K2TtXeDQJ5EP
Nj+pCwa+X6ETxt2HSVEJdZAgzh2+RGJpXYpGcekjWlv1Btv/B+E7W/8vxR/sHwjGwIJLNyjjBLqg
uyQLB5ybAE8aVpgG4b9Br6UU2HfJYrHrz6vYAtN9T67OblI/gylP94T2oCuKS4IbO9lYIVPN4Hfh
9WNq7KvD05Ib0brt9YX40XJ7yKJJeLkiCkh7aAzrRiWytnMcDaty392GTXVhlqB9rPmUJNkmhqvg
/u2+MMEz3uq8smIUxUjhJ1hT5xlpadobqMrwoGmv8eYeou1CMDDwa8GOdut2ORUMh3Y1x3nMVCYi
lyelwnNCOPh44wKbKFZXrK8154huuvoUbiBFzc+KZksRUCI/m7v8HzF1bN1P8Np6eS19NUNa9Gmr
hjkija6kQXKxVGDodIX/x6g7WrHCyRt4gYXyHvlUMLWuulqTlJGsS8GAGuyXba0+lpPcQk0X1tjl
y3LMy+kS2it1zoqKVrcfHivkdx4722LH/z3AoIcKoC991IIL5m0xan/pBCwGLArDPn/Cl8vdM90S
cInAnpu0gx+/whvskavYlhovygiNw1gr+EhWqPiVVQVNzYiEr6bqcCofiJy1YY542Lu7dVbGpDeW
llzAInKnb5cFJuLWNzhBA9Dc366QM1Wm3+5io45y70XpzKyXInk3XD+Kzy1HPzr6fnzwMxULtqxg
Lmg5e3svlVj1t1Wxg8oJCV6Gd34awf/VltHHLd2wjm6QUKrxfOZ9lke8qzIhIlFjPpMB9q/ldhCC
4Ci+MoMKdOhCzTaINFaVKcOQF9yIq4zItUa9YgXrj1p81uX2UU+j+F2Lknghie+EhQefBrP3Q20m
cyaEdKG1VNcBZHCsDTc80z3gWe0BBmKMEfV5BxHliR8MqMaywhhVz0WGH9+H60+YXHy+uJduvCSw
KfGggwz1wNt5LcEktjQY63I35Au99IQxKRU72dUac+dBBgGelZDDwl8cSkthcxYwdMjMjUXt99Nn
2AhpJ8OhV96fq4mkQZ/UnbSbN6Sszt11KT2LoM7FJ0HbqBwi2o5rYa5+oDqGVO/Fpqun16OLb/V6
vgC6F0e+BMWWKyR+QB6FOXiDmCreqKMpZ9cVb/TEyTOlWRsclmo9LloI+MUOzJhMzgkRPi13miAD
kPfeFYw5UGBiS+50SQ/lquk9X2G4MwNw0QeRYJSfi9qFUrAUZ9wH50m0h/aY7utOwaH6YMhj5Fgi
qwnRCfoWxGGePb96Nlc81S4DO6In0PtQ8gH/2tpvqKKVkT3EmxcYX0mrkP//gTDJEORJhp/kde9h
iP3rm0AL4fxmcqWwmYJ1RpE7qXLDF9poqdp7uS9BYBmH3zkptDTcrdWhr6sdlkYk1W0c0A2c5F3C
baQdGKbiAv7slL961DbGF5Mo/ZtQ6s/atjQ0jiYmVijCT/cRrcksQYuEaH80NxnwG7cDsnj5GhGb
ITgY4HncfrfYg6dMKij6VLHmdrGu1qYlMrBxKfvxtEKYlTSqWbKaR5Tqk/C6UXmJk9AzgKAYhgn5
/xBz4Xv1X7kjpE4AJ/JqA+uURZbr1BiEtFEdXdqeSn4AONO/A8zsjKEzMJTGB6CAHdWeoWZuZixu
I8dWLENE2x/+Zqw+bpGo/vRpbZpe8JywHQs2K0Rajp3ce/s1noSMkRCugdCeWxBrG7GLkkJvuoYC
G7bptBNi1FDg5twdtm/8JI+zom3h1gAobgxMR7t8hUKteOlE7iU3iDc0tZTNnvXAdGvWREWCVz1y
Q0F7PZuhk+7eGfkd1A0NS5hHlRDSJbMN5XPV3ppc48hq6R0cSGfhXKZN/+sZTzlXWSaKfHvhkARx
9Ix8HHOIEly03/6saRDv3PqwVSTmMy9whhQtz4ch+/pLEnINGiPnu/SQ+yqMBn6PPO1niDTJQQom
JbO8UAc7Nj9aQH3gTa3dfoVRIoUsqLOHpJD64vMR/7hS65eMofhsDMl5QutsVOH3UH26yt1TQpQ8
0rXbWJS+IaYUkNh5CjOA4u2QN2LdRUqdUQ8Opzt9edREdBs7prLvxdvujlsz70cNXOmorHwhwggQ
9i4rFRUHcJL55Z6VXfWDB/LD2gCSttW7v1/1COj0emXobiZMHLtfFJZkYf9dOPF6pHPlBFqmQxbx
TXXomqsgkhVwO3vpCz028R37OWTOF781Ca/8OJbMtGwK3zJONlV8XwUoy1GO4NGWoZ2kn09bv+hs
mpwB2Id80/xwwVayTD5sF6qzriRflvKGrPc2zaHKktNMa+3gHlMjBX01yNBmjMWkGLS/kjqbDTmO
LVOeE9wXbicOMNZRquipTBbjGrkaj2sQFXCt0THahthr8yDe5DBQTU+Fs4zUFQ1XF2wYHn+ADlT0
vfj+e3JL0gwFynhp7SQassa4lvT5gkTIdMPrOmtFjgYv5S1tShO4TGFsz3Ou9bRB0eHagP/Ldz5U
BpXGzf672jM/45VEPFE6vG+LTP4Ed1w1uBHmJ6UEiEg+E6MzblguHEwq6gBIzE92NNDjS+sGITzA
GuSGhlhXohhUJ1CgOCF+O0Ihln1JlYDGiFWAGKNWHcoG5n+WwJ/v548owtQErmljCf8ZCvNraIjH
T+AAFaGbbrcIolwq/SwgplKoyChAHV20hoVultoYeibfeCV3oC1SGDt+pEfYNjNkJ+OvMPZixiVt
HeGTB/EAW4YJAfGYbwBRnzSk7QWy36xEUm6dwRvNENCS9q7saTXnOr52J3X0yYD3Azis75ZCy8tF
ClXLdpmYa/ArXIB+l4bGezpfc0ZzJN/JYoWmhcspom0Xggs22VHp7+aMW/Ij50xLvfaHCw91sGYd
0k2kx7cfgHv5LHW1YNdc+kq/ymI5VVPkhbjbExg+J89KeLYP8uKtVudv8kzy3OHwSrTKGa+ajAH/
rgu5NgpuvYnuojsStnZ2ffl0m05oIAqmDfrAHyIIZo76imX3gogZY/hr5gzpM4FaKlV3N3YMpLtx
fXxsBl/29s+vJ3vH+JVzxz4eEiNbcbJIh3AtkwRfWP8MvL8A8mxRqkSe1s9q3cDSaGpe0DWXz2WX
C3APp9eoLyKNazDtwFkqoNZMRa/2FGaA03mH3QuFEv1pVk474qIbxx5JMxGNQgIp2P1awLoawTEM
N3TV6ybn5ENSEEbcNLxUnR272i9DJygW9lTBX5QFgvDXoEXUok9d+4MbFhmwH0gp27PkkEHKHFiU
a8aOJ0+GuY6JVX4XRyPqh5lI78cGUFOsZLzTwQ2fqcfC2kxxYLawQW2eixjHrMQ2aTq7xL9OVRsV
iiGu0anNEUZGnYpERvcs+De97Zk3TvW8beTRNeBZ4ZwDfh1KHxfK5kyMPbLBPusG06AfdgoeZm2U
afKtu+D8ZfohMuZeyUqtZbwRKoDXR/U/18Sfz4tsIW7+ATDyKD+mST2tkRGX/tn+5JAma7w914GZ
iyd2JaPfJPe8POZfRNwKZTzRfhEZSo+ZcxEY2KgStnGNmV1+7YWiRHLJJwN2YL5VFDcyrIXiyzY/
pOco+q3RLXdyjVP4DIMm0NV3VHj95ZF5BeXnOmz0xjcMfaAwb9819u4aRJpajO6cKSjEnRBXQUSc
lFzbYqKrZSYUrbez9E/P0owHuKtLq9RiDZRTLqHFzpcYfpioJUeJgleYnWod9CLdftwCXZNmvW/f
vL0rll8zc0aSUEqdfTp8o5fMnpokbEC+dpVllfg54O3VOoLticoD74WJfMUcy+tKIQkwxpmkCSha
BjZoTcpMq0gN0VVcIUjdEC6eZmX/IHGt2kLxHxJniHEIPFqmcImStg13nXle1IC7jMsxjNVrUn86
hq92EEuJFfJ3P4bHAbSo41jcWpT97wr9RN3Hy6UhyrbwvIeBWug1occACSqjc9kVSfH4vfiUDmnp
IIMMPhUD5CYVpn09xBDA/jR7xP7A/wLtRIDjexN5B+lvdo8TglY38UOoxddVoVa7b2AdN2K+llsD
ppIs1iBe0LP20Kv2HKLpCaIokKaNnMRpqRRLmiw7iUg0ZOPF4d5ZlXw0EpDx+reIQg26+9VUJU0y
SAm56l1gEN0w9C9PGrqbYRwBYPzqEVp5EcrR/1lh+AT/c2ZPzr2Uv8bbUB8CiaJZ+cKmDiseBnLi
3cM0o9B8R98HEB4wvOxAz6gjzN2mRCs6skK17cbnqWmgrtKb/Yr6CFFsLMvOSk3ODkOHjKuayg8I
FF6YAzqRWhwXRKubv0FUlhQ/xdVOImhDFgmrCTys910MKnReAI2OXclSv1pmkgdI0T9jcq/fBsx5
/phbZT3r+980cFsWmvCOgZ8RJ8ySwYnYX27MRS0nkba+K7x2Tl2Po43PQc1YYkYDgpkTtv835q+o
mEiLWW+ZaxuneBKusHiC7mDPE5shxQVKxQm51k4vMI4KF0d9JCzy7CebcsCaXlEhsJAp9GUaXpdl
da9SVK/k4y82XPKErMTuIHFyvP0er+P1B0PkwE2F+KsLTRHUIykZ51MmafbETurGL4PsFdJcz28f
XYDwYpYeJF+BAYOFGsqIp8AWRTBUQGgImKSFp3Tnd9hNXhmvz63aze0vdbbPCKslO8EalcaKh10n
BlahK/ZyxD9KByqTX8tmNL29nQFz22VrQQE2kyHotaBPNVi8praDu3jVXWWP+JpmEXtqowsI+aEH
7LqZrbjx+5VNpFzoAe0Ol8uQVYEWL8gDL7/RXAxNefuLJPBSlnPelUvWsUETCw5J4Bymr4J3uqL0
LRX9ctJK8ZPkYdRqkkc2kVv7cbuXooODZh8cAjI6mKVvKnmIX4dvGWh9ioh+aPAkBRoW+LZ36zvy
h6lT8+FqlMnhR0s5BLaJtNzQfRn05RKs+Km9ZEaPopna84ggGCtMitc04V7Vuzdaee/w2dig335c
y/NMUw2e3zto7OjVTfv1XvrlikpW1H+xsM+4R5ej2VbT5tEx4Y/ruptYPjqw5ozEe1O9WD+wVGz5
XswvpZNFlZDt0aI4baOIVJH3WOyu57iQWMwPPacFBd3YXHN7VhFqI7Bw1kxNofifv/gHS04bMTGc
e/iHdjiHFCIVUMoInWaLOVzi2573TuIBuEMHsguWKPnLU2O9gkTfynxobwsULV43kVAw7xhJy+cv
0yBQ2bYxzeMIUpcfW7LfNfbc5/0RUkU1SngqmfLfLaSMXeu1njx6lHPpdsnSQaICiTsQ3Jeq/So/
KZ3WbMFnBe/+9aFmITNcq3JkyD1ybcdUQkdQx3kcay4IHHiTvO08Yoh6OBOHKH6q+MSCmf2Ngs0O
DlYyOoZWL092+fvro3oOK7+MHS8BykEoJ6pOMR0mcG8QA2eP4FCk6yKkpbB0WxSJ/JXWcNOT4R5j
I3YrAUkRg1GBjH5J2WVNnUHBOlSLvMjXIySPqYXRxH1pD64YRd1sVdS39DoaOcbBA3QjyXX+jt9J
lRs0MinlbOnTnzdISH332ZX3lloyqaQCVOVTSJppcNtzVEGMvOf4dy9aHhD4cYsMEPuVmB11SVWm
B5S3MylO4hQJUCm81Jo50YerOeoJwt21oFAgvPdP7dJfyIQtCTSfNbNRxHFGfXmYO1iQWI2zO5Mo
ojxCrgKYTD51i5G3tRQvihEUAjeVs8YhGqJqiKP7jaonJX5BbZlYFevoDqp28i02SxtB9O8vgZX5
OjSJFmNamxWiFlYUWkZRLZE9URnnqY3DkqzfA5iespbJJ/NhKVw+qLdUe6z/Avi/EKzo9/aK90jR
QB9UVEjeetrNQGBKuzwUyTE0lDmkLhYB3JRKgweTtqt+sjkiA724t6Wtmpn/DZFVv7QJEbHkN86T
W1pojNHD9ed9Yd4IsL9xokBlZpVgayceXv8F8PnGQteJ7kVeH0lznSaPpRiYXXVLNPTF8EfQ1J9I
FujxyVEmV1BTQxUqptPZ1xvHUKUGgarTDYXAehfWt1GZmO1RENRk6/NSRvAdzLj7eB+obCMQqlZr
uGSTslKUkQvnEV9T5bA6KvkKgxcM75DS1YjN9a5TUDiZ8LQYWEmK0+S+WRgNdOTsd894Bt3gA8hg
EdnaxdmuLB/4EXDl53QrjbBBqB6jaFYQx1hvVrDQ4paUSfzharmZPCpl0RYJv2WEouoMxjJN9S86
xH2kwSuRPSesDBNdFbhW1PValrlJOg3B0tpX5JH82XhLhlCbQYExFN1pW2sErrz68asw9gukg8+K
MPKaDAr1PvRr3I1+m/5hIRAQAy4cvLJuH8lraMyXlj+QILL2NIRDNPmyoXB+YaQWLY2f2wtcn2E1
hFL+VUaDpau2I6bOdmPyK8HQMTP/sN/4IU68d1mc1Q4kGg52Y0CUz51Gow2B7CNNz8pWKmAHX7H3
Y/Vc+K/nEm/GFMcqbdK+eU3KZS3EpUPO+h6ht42jFqF08wkTIHtG8RA25eaF1oMKyCzwGp542h16
4LZIpXCL8Xzw//R5YBh2MnDjOKPkuq/awZ998VEEHiUQXqqY52LXx2H+mBeHZACWNH5tXTy74nzY
DzPplO4pgGEG9MilejYNOsvDjgwJ1feSp3iRWxbXZO+QDDApc0pPT/JGsci8tVSh7xKEhDfl4ZIF
5XwJV+qhQsGISfzOy2DczwSwN/HZp8p461r46lZ9d0td+EZehVdWHQSK5+krCf6RhhhyGpHlqPyK
YeSSPqtEX2lp957kF7bmZ8RLWbplnwSXMTOVptHJ5pDfgAkJcYzbFEWR27RRxGm6lW9P05bneZFy
UPeuyWOkgpTWusaQPN8py4Oe60pzChugSu+iwEh/N2R3/j3Ff9Tjhjc+Ds+6pLltcqxvGJErqZDS
UOGyibxqG1CqazrosD/wrFuxY8dTyj4Ri7RFQRaqfrrGLgwL4oB0Bin17LstAzU5jQjXQ1BlnHgb
LnKgQqyVclCd6saQ2DQ0+od//WDfb11LZT1ukxmIapBoevbRZJo0NvSZcPuyAHua8M0hJns51PbS
Be/1iNYsqKm5osYBUWJ2ujSSvoOt2u8y3SkLfreDefjWUj/3QzLrvOOUcMeD824SDvPnId7q/mHc
UkIqnyhIwbEx7ONlfuJmGuOOgJM36WtPRlwvOwQJbp0tPAFbYXMRgAmasvEEJzX63g3tSbkLWgfv
pO+yXYMMAIp5upwJYofpJ2wDR0eOn8c17chy/jlA2nZpLXVHAkj8OX3WAd0EQXYkn78BQ/5SMcaH
TKAHfy69sPX89InrFk63HE6C6cVYKT+MkWcl2xCnHzZb2q0LN8cGWa8kN7Uqly57kP+qDfLULjFk
EdZzCJ3MggeDNdjCnnRwQ922zI57uhkTQwGeG1dpp2gb5EFrRl7U+b5M09+tPzwggs1MIzBorDHD
XH5ZXlB9YMPIz2iCpgwPqrlhihZXJvakj734jf93n6tCkrFrqi9UHKFxGhiwfnHg5ho+KFNpT+L6
MawdvG49SNVrVqaWpY7sGZ7H37OjaAFCA9TPrQ4HDQMjTJHZhNQoS8xqjFh8d7mUEmbGuE7gIL1e
j0zjRz8SnGDAaCcn2E9A1yxxbFCtrrrKoGtBpTOjb5dNP9npU0zVjAKEMCdvOwcHp+X4JSvx5A4l
Iyzc9j6oVfhLiUjhtlhAj3WbpUM/XV6cugI+qL2tSZCNyJRVtAR8b7lRBThdnEAdc/Rbq1WMR0My
sHN72t97agbkxEsPaWBUHvtzz7oCw+OyGgmq/EZL/BhmGscEiMSBgZm4zj3qBrvMCaubYhZ1sGVs
tc6Rsw3j7AUXz2PzOUqFJqNDzNib7h1cUt7111/wMYZ0qt3yplnKs03MXEquPpvG+kKMaPhTWMmF
71uMpdwtfV0CYx4ChKK/roWNSTuXk/MaPF+r0OsCxkvKAQJ64ezen5jfFtNihQGk5JLR6zHASpHl
FceOe+uhk0ldUkwXUKzokbLhJYY7A78s1uZSf50mX1HEAOnGnUe+I95wdcm4XQftUweq31UGWaNm
vHHImSHa+ubL8CBRijIKBmRtu1X0cRzgl9mfWW43FWDocjXZZ9JDH/3JUqL3UgdGu16LBjYfrVIe
dGRac1HhcHgOscdau7c+6hPLgzoA9JCJXdcxndS3bR4dA35wkIIv7227mzKsZC1R3iNh+SK0SZGG
Mk072CyHUp8IAucq4Y7CF/LEUyuOsCcE1Xz7hFvDwxTi/5ZA2C/vdUeTFYjdrfASNin5jSdRxQvX
EjGTdcgul8wqoevXcsP/hkUinhB7AiegaRKFt+ABr+Qq1QaULL3HUIe031ZaISQahrWi8ZrnEFSr
cuhKfhd/xIX3MxnFkByqm54ozqK9bqekDSlOpERUDT18Gw/87ulaCEe1Yjd13nw48snAjCmRZFuD
LPGW6hsdPdXWlP3wMYfjJmdr463AptndHjq0H+ENtli7q9AyE5vt7LnI5t0VXn2f0T92AntwulTR
bnGhd0Z0BaJ3D2th/2kBy2Lp1euxtKNoR2xCKJDZo0WQ01+brYa5FYCNcpE2K+qbCd5XxqkfGCJq
OKiEwl8BboWpW+RZ8japgsjmT3gOpLQW1ZrGhtU43mrj6HQHb8xDHFbqDpPJFlliwP06vO8xHAtd
FXfTuMQshzXAQxFcdKmH6joy29LvDKMUy5IkETl+0JrUsgUMNr2SgaGr6sH091Y8d4TdWpLVBu8K
nZJ5sBUx+MkNOSdY2c4RZ7R+uKwAYGhAIZBwrXnkoskoHXQ93Xhd0kUmR6armXTXXxyiN49P+jn0
pt8ui+x/xW+xw2QiiSTBpBIuhpSSh2UdYfqhbL7LIUrkpZ6czE8/6XKcJ7f91vqoDQ8Ecp2DdYlg
fuweZlEEcdP3tbdOOaO5t6TY0xhAI6tYd+u8pYO72jQKZy/fB4Aa3U0XCF1WtVMbfuys23uDqYl4
7KuUtub8xazKM5cKcJCDDB4X841TzHOVn87V0pjLGTYPMu9+3gOyHGHvevCXtrvg77OJI/L7Lgfz
xvyq+IrAsSK4JVYZSRVax7pfBckY4Eefd6WwBciGJjorcRsnTKtponn/ng5DfpVSe5Y9+X19ntbL
BHPxHuFRi5/o/VlsiDKstF0IcHVvMR8OgiCAKAO/VZZqhNbSDmW6SXuBLVNhGmLIRli6SThAY2np
l+utWzKlZhqKjWUk2miWwPZCaazZC8tAp5FFKAD+bQ3+dUxEDUtKNj76DrsxpRYWX3WvVNDDjUgY
u4nR4OuT3Fjtm8Q4u90WIySQ8k/yXh1p75smo1l1wA/cy0358d/bWB+92V/3JvDt8YpfCxntMM5t
5gBrmka22IRDurC//soBoo2Kkb8CWkTcd94Jk+V9oIP5EFeDY//o5D5Sc1K9eli/lD8twpGY1bx8
le56lZ9NEWPieC5hhB7dmfk6YUzOzWtcuitWBGP9lbM4uzUqey2qKDPObO0xhg1vMeicvHfCFDzP
KqMusHlRAE7bZGUeDTlohS+IBkvRzrm29R4VsCwNzjKDRlL4V+bE6l8maqQIEbglKUsOtfStJVj1
Be1kEDtMNbDfCyZGTXC3cbiNYXDbtdCMI9o37sAqWO4lQun/tS5V/uBj7zQ+IADdQffaJZIi8Mfs
PZgHRzFuWK9l+C4D9Yz2D5HPqHV+kJ4GfxW+xIsF09CFDTcb6Hl0KKs9509O8vHPtC8Dj5DbtSG3
gbIvx6v68gn7HE8sEiyiC5g6O9YfUnd92AMBuYbskW4RMSfrL4oUgYConmA2SjRipyYj9mTzg8lo
al/AyI3Zk0bKwzcyKlQfOiHT0YnA49oLbMY42FIxnS1MexFhMSYnbAMfsFQx6xZi8JoQOu10guQS
77qLdpVJJfGu2XFc14617uVOIKjCu/ZD4SvRqZO5PghZz6Ws3BVPMeExRGnUz7tihq1xPy4/oMR7
+sxvbkl+F3JbDTZVZYVyNLuE438Q6taxDQ2iRCL/9Ps3DrPUK7xK7SXIK/v81XixOwENOupg/9bT
+rolGlN2dfg/FArZiBuNKGEbBuuopzJxkqCmufCA4QkkSC5x63rr09Ioty0CQ2V6LC6rTdjN5nWa
LsjNukXVfEeAGRcemWNzTjTC/FatAgjl3BHRNpQULuRiw8rM1j1AHfNypRASuEx1iB4T9GD0bNKK
x3APKVpHWuSMhwDZR2JU/END9xDb/IofG55rHK9GpAuNrIH6Q7cJ8Phycsw+qGh4jeHwb59UQDiQ
J6tQUK3DvVp0/taJikGA4n83lq3dyJlJNLnTVvZX7paBRoRICqC+iXfHyZgTzzYiR+3TEbzQLEjn
5no/8eXgzBem8+tATizOWKV4ZG9TvW5pJVSDFE4pfe+85rwgaX2IIxiBMrOnwWRncRLYUZZK9DUV
5zCdkBtu4Y1i5kD8notumasZfsZhPHueyUJs5k40va3rNb1nBrKm52wC/WpIpE8QYYCvUixVnMka
PP36Ba+y1PZjzOqqDoNJjsuZeSS8K32K/84y5jCQlh6AGLfke8dKd4CGwGC7+cuzvSfRivb/EISZ
K/D1aAoIfH7MR9hxr/h8WIPt7mwUbWSx/rGY4k2ZiySwbwy8ijf3O/rK0RWmIdNHP3qIOUmzRqkD
hAR0xn7GKeqUxDup45AvUDhRaacM4QfzRHWkj5yL9EdrFPAXHZLTIvjN16vwMnWgfbs814a0ywr3
Ppyvs9bN1t6+dpXsqCn9UtVftAH6nOhyrG/5gQxIQvIdqQZUpdKNgXFMCgtBHxMZIgoc1fAw+Sj7
Hrgj3muXSZIOMXRTctvTPM+A0HPmQ6jNSedvKnbBNVGlm1mvJ1ucjZfKGylJ/DovjVJbv9/vzxLD
t4bKw4GMaigaI23+3Lg5rtYkZuc19C2mXG2/PlwZvtnrhsGkG6OD5e9VFXkxKE1Kf/rfiH78VKoh
J9/uqBhKEPXNKg3maS5Uf2a7bmMORUSYDDMhM42yT1apmzJRaOHSrJAZlHoKw+qBvFwG0VIsSQEl
16oBwMmx6cP87Zeu8cAlj8ZHXRqdyceWePtjoI2MfAVB3ndnr0dlL2EEdwlGqXZ3jbLlxVAoDx+U
Q9YURFEpNunmMFxa8K16uq+iyAjGUy+6bTXHBp/QLoUG9Nqj1Ks9pp01PTFqPd2gU1o8VBV4sEX+
/Wthf3t/un1Ml7Ob+rF4ZnrdxfPuZ7WRzOcKQ+GQMnWhzMJHZFIJjjoBW1gSCazEAu0uYlllJixg
jGwMEnABSk7QOrVLUGVgOwqjxWlYTR3LLeMf1GUw8GxRUzKkrXkehkXXczUdShkzg/W60Ib5MC1Z
8uS5RKd9KMBqCewGZrizAeLvBiUuTYTeFyb1/tQTASz3gLNrgAAY4EUiZVE96JPEjIzMJ+rS7jGu
OCImK/0Jj273l5JiG8FXosNjEvpCmdcKu00q5uo05Wot04Z8lHBxs47u4XGygZFK5al1eG+AgJVZ
vZRh2+RMz8dR7wQh/kOlRMrGZTJJhG7U79/lgrFpG32qKeNULer0Eih2hlcAma2yAVK/1840n2yJ
jSSIvI3vziTGo82xEXE7m89GSGLjqdjYvKGmcUyXDQyBkt8iahQNMw2d6pqLPSbhgoaxD15kou2S
71omIKHFRY6I4thlX60nOdGPcE5wh+IoWIr++R+K5i4qxipdj4EtHu8fpDKfCFKk4IVw4ue8HkGo
PwcWsjzgn/VdphAoOIlNwf6tVlmPs0uwgWuu9tj3m50qJpWYOTAABdJGW4vtJqCZ4rJSBGO2asJM
9LWFUBVYvewpcQslmTWYyFEt8WMQzSaj1h681frFD147lRngH9PBwgYlpJhYqYLm7zA42lXgM03p
UYik9KUWB0NYhvmQi0iTfCVbY42CNkkOxx4V2RtLiBdab56KEQfjicyhEn1PfIipEJRotJgvCfgp
wUMumm27hXTq1JjHdAlZ6DCS7G8ZQEmy5TC1TLsLehZ7snExbYTC2tecixu65e+3sOBDFXEJaNJg
kxVm8l3/uOb4iSCPh+sZtv+Rv0fwF7v8hMlLKM8aRhLNv4DkHszBxtL/8ht5HQUe4Q3Miy0AzMyE
qT/U+Jg0/ng+TphNvkYNRNX9Stw9Zx//nGlJ5CJyhdIdlXiMJxoHKy4zm6J17HaG463z6q5cOq3u
yWeAfw/enyNb9MgmEeAbq/uNQlgvmphv+0BKmuKvQG0TA5Ub08Oir5eksQF+sIbpcQv4yOGRmd+D
mc4Hlwz46nbPDon359u0UFvUXgtwF4N7/v5kl2/X4zkbiybiScfDf5HZE1/tFsAK9y3Pk5YDU4US
e2EzomRaZGrCCg600nRtgSNEyMealKVYxDZlUQXohkWpuGa699rB+B2DPF2ky7ryrBVHOaGDortF
uTJF9AP5WpktOjgROdqdGvg4UROepkIUBH3IZzFOMiMcCfMqurI8qZZDOTVlkAece9YkK1e/nL63
EQ0Loobrb+d01hGOW9tjsxM4gzwS2oizsxzWyAm0hpBPKbqgXa1K9dHXTbRc/WDF/TRW1oyO6gGk
DCQIsgg6vuROw9fK/erP0pwtYdlJcwwaOReEd+l6sBhfOdXWXMbROMsxFuMONSQGpGE0aOodsAhD
UXS11mIB4S7eZzUibYSKwXI2u+YbnPhjKfS8Vw2hHFyDMId9EEzSAqNVGeV7Tjkr5+y2SJWBte4h
4duftWOFe8AAKddb/xsrthwLPI9XCrYeEUX6hyoxS9NCkJCHlYtVxVh5B+2zfuA0avh7wp4zCqxS
FJ29QE9mz+VUT+bvKpomrGSptgTY9Ea/w0zuVg0GK7uYlLNrWrXLqpU7FKesryts506yDJ38FJ76
B+0H3+pAbM0k0/u/nhMBN9hAZqEC31p8nI2jO8vr1zi4T49GbYjYQuLKS2Dzio2KbNPBCfcBNdio
g/sXZeWO/nJDoXS6lle7Wm5KeB917wqNRKvQJBw5LPH5d96wYFQGyikzN1kNf23UBVJC85VYXGbi
A9SbVAs8m9ym3rA/XwKEamFPiy/dInWcnkZtR5b5bK6GjHyjE3+i3oA1IGsars315SOANxPxmdm5
nB++dky49hF6Sk1H9R7kt6+MDTfDZhMBXM41C1vPc81SYhnB2A2PMhNXizG8wA5AqbxMJ7CjKLzz
9r2iZjQ6tprXkjJG++zYl/kz9yTHEFOtCOP1V5iHYM6aDWKTHG2V5GONfOPbN6GiB+qqpT5bwSji
OsUOqGzJXVj1UWs+Fu0PqXKIuYQzBznXYzSWAIm1fgFky3isu5LkaFTVT0xS2J3baoc1QnU7MBRn
WwoZkyTZFgpZT+PIfvdU1AZlt1KYIcRm8kFlKAhfZAf8f2z7+9P+7RmDhiakCYt3oFrbw0oB3JJ6
Y+rL20R6YSW0KUIXTkwo/ejRNdCOevcst4C3e6YpvYZ79seFSkqnbtuz965pIN+vvStw/RQbJkcN
fT/NGNM82DF/SGh2s4qaK3o81evdyOhQdzhg7q1QEuoCuP7qAlLj9Ix8sk4BJh44HlNFyM3UQjE3
7IAcCjWnPXdMPf+6hSUNt4Ke3kasluqy8pBPAR0hOa4fCtateuMT5/YFzLmJxILNUyKnfXtsomua
DZvdwIzkJRAQAmpaByqvc3IYDXjtaIQUgCxqELfgKUVwATlzRODHFYLFk3mMdAyGLoVh9vEEIQKC
ilhGgCoK5HP/x7XRfS5HpT2CRY3nBdkE3pkxnj8q7ffB3CiPRD9jnbL7wmG0JbD8CAoCCRWt2NLU
42FfxbhfSVM0G5U9jq/mwRS/dylKWr532B+ErY9Co19jhKbtpsWoG2kZB2XjUsIDY8OFtM+UzsL/
GqXV4vir+uYdlAMR08dpl+BJFsxoEOZzMu7PPzFAPozvxUbFtAhWoIR/Jzz7d63G/wmCmW4Jv8UA
wl1/05Ojs7DEXJiTg2weN1wAnp9M5XQA9bWhaxYQt6A/5u333QYFVGBGFgqBFB/R59xVGH118+Zc
Bj+5bCYyCwzQOOCn/WVPzkPn6T9rASJTO8PYanXdZAMtgOk0CqhMTXFuHqNR6dnZGVzUXqx6ibx7
4shZ2MFWXwd5Rc3mI5lOr1H6rkSEQGlnS4iHFPCTMJculGGOKN+SNmnqgSwhaIQpG91vdziydwIX
9BhCmVtWa6oM8FP7OMiVTSiFZZBefYCMn6KBAv0DVW/bf2zR2eMbF7FPnJX+WdkbkVxLPGkPXsFT
2g4/AuXVx1RmRsVRSNH6p4plDLAT1unXyWWRsBeTCNlClXScHpk6O9N/5iJsFh8mTR4vh0jrFmg6
kPq+WmLRBdDMClU7Q0zHHcBionIBbPfF6PUsvrsGXr3YmzZd/abUVWxcAunZQUXT25kL0MRvJsuY
LZl+MXFdm0/NTJch5nFazbBvES3B+N+btxWXPP/o3qZnqnQ0j6WaFbd7T3xTVK2Dn5dByVUpOx0d
+Mmq8bEINWSo+xLfvK+BxSkRfO35aN16PbcGipxO32bKd/nNrlZkD0/F3jgdD2naWIlc9xIvgeP2
G6w0teeJjvtwUa99KejSe34Ahj8nQsjaELnnADhoPOWA/9YeRX+qWXTvefILgwm4ShgSurGrQ+Tf
7bYrDiovt2AzdDzoJD8ys1+tsV0XhA69udS7YEEpqGBemeaVeDZ2N46P0uWzjw+755WqGwgvKHxL
t7TC0ByLLduXcLEcDu/rbM3SlmKiHxLoKnUNJSRtUIo8Ept+KJy7E/6aMtBHoW0VH0Uk05rJ583q
3/UeqXrMKm1M5ltyVmYTHXFEboMTowwQxVsU21YAluAvri1yAd2/mCdk/IWWPn6xFvCqDz27Hm7V
rAN72CJfEEJBF6Uo1iOcXH77jLl3eaxg7cerwMPhiD4RIGTL+Rmc6nHqJ/wa2g8otdGxo+UTZpKy
kzZ0qTsirOryz6GtBe3PHdKlMGqKUq3PDPdpTTmKqWzDH0HlfC2lfyWszorOWT55gH3PUhQtiOLQ
hY4W+TTFnmxff8D69e9Ob23SK5yAXgNcd5iW8muqjBajo7TqosGgKucP4C/rBiEV6bJhpk0ilNsQ
y67Y/13XGl0U7YSL+xXD69lYtOadFSoub2YlIGu5la47CQkpk8pmXNUfdC/wyZdF3Ke69A3+4xNP
BM4zj/ZkwPNF3XPGpapMBHHozJXcIWcjTm3BWG+MjAqVIPvuRFDlbA83LvwYdMCOmjo1Szpn8CAN
DvvIYTY+bKFszyiJMdgN8PzsYhAE8dqBUCg8YC8z1q3LHAfzMzRKO4BrdX+4vbCM5JtzqbbGpoVu
tt7LHmiXSvJY3UzZ7WtB4EQLOvTYeEmlFzsy15eGWH84pSSZmmoGQF86TdddjjbUlknpe27BhxNV
mIC9xlX0PztflTmzuUmWr/FBvG9elTuYVKEufhQsVQ1f+hqH69HLeyg9H80JQatYjMIEWSnAVK70
xnW016Ih2q8wUH/oM9LhGG6XbmyH1x4BIuWUsJYgkrtIrDCjyWy2AfTVVWWpvnEWcSV8EEeICB06
ESLGSBcOdmaCAbfNDCVYv5jd5InVxwF/9oVVywX5I36OKHhLaKUT2yYouEPujuSTjbS4r+PoIItF
Lv43jrrq0iDgcKPsxAqFRDy/NvBQBt/G311mTg46VH71X3ykoQEAi0925s5N9d42eWXcYpw/sBcu
bX8lF+LjK2zt8UVvY+Y9eqrZnh+j3MxBVhUzhp1omgqglyjlx1rzYVXgi9WxGGPU0tItGESbJpzI
tRMNk/Ks851XPoNyowxDcSILWk/cvS6J+EVM81atGuHnxKjv0OVgMBujsZhJGA1b229yHYScXgsP
TRG7BDpowUPuvtK6VBbyYWqwD0RUNuNNZ3ZkVwdThp8PRotcuxDKHVNEdEafl6P1x5znMi7oMlrM
iNIPJZqJZep+q3qvWGKHiMn8e7pok2KwIbXrQiVYeFpNX4OX5wP9SUM8svWDk+1LQlY9wtSMGb0/
szeQ7Texr3TpT80w1lI76L3BNoRovSnwpedHSv1RhmJouAJjuRmjElD/qWAfwL3uG+OMdQdOmMV3
k+KBuAocSNF/MD+rbeh5R7T0DXDK0Ol2qbTE4MrD0cdKR6MCfYu/yAPOzDxVuzQ3/uHF88S49/PS
9FvG4OmUodqcvoEwjxZ0Jsd+sshfuDmiVM8bx0xfogzPyKOJWBTmMHRcdq1WKklKZFhs3/1l12eE
TPRhWL6JX+CMZKzYIeqV676zof/R+uvpAF/Hl9UPR1Ke/9F31NB96ojT/lxN1Z61fY3syzwhXdKL
yFtY1HH5O8N5f2h+YiM4odQzGwb+eX2/mP5EdtqTn9Ayfjtv6k//9WQJFX8F+5geXJjPdJujdaGd
a3fmUmHMvemEp7hbL148szSVUSNw5VIl6prACB+uGKkqYvXQblFH1WtzFctxhX8a+gPMj3UAnph6
Ld7Q9Y/RODmHrgPF81N/Ny1O9xoPyYvwUdf7dicJVibCpYspUn65/SrVVd85vh2ZBmVkhCHBH3Tg
/MKoyuBvOx1yOcj0DqP62ZwqQ41dNXXzQ49FxBYopny8pe7nsqkTWQhxQCLakoL7YJlTBQ+yRSDd
6iFUwVUZrJkoRO6Gk7ELA2fEuHUs+/cGi7POinfIDM7wacRTJN66yO1m+0c7hWFlFGucdnGaG3Iv
O3btsVrZneJ2eSGzXL/rAUgBdJ5rrww1FI6aInxvat8VQvQ7pONXe2gwi8tqieMwIGoV0wSgiApT
6UlmcPYvsjQ1OE0R+7ExAOcQP3aU5fvNzwgeXOZAMbomd9H3KLxeBgpJ7Rs5b910H5Xf334uRZiL
dwJbQYTb7LVlMzObLzzL66420wsGvfPNMvK4ml4ib3KChqPWm2J4f5Lh12NKlesP2yfWdZWwMn7Q
tYikSJs/BWgoJTF0Z3HyaB0sGelowFHigV6kg3NQ2SUeyFq4dMvS53CuYuIoydXzG6OiqIMhlK2F
C9O4TFUEuEYrsriDcVXHJd5pCg/RVq0Jh/qS14rqqAtLTCGyMi1STEAyrSUJZHcjghEaQTQpQOaP
plsz+J4WlPpgDgzIs/MRguor4ibz0Ed245mrd72k8vgXFTS629V2jrfUjPh7bl4OHxcpx90iUTRS
uRufd0fFFEa8UVZt04LtdoPYrYIIme32DIU+aj6iFRPfzCmBnVv8KSw3gOU6E+InBUEnWoyHHkiW
GuN8Ks5Mk3el2s/6Umd6nbY3GZ4YNRBIM6KhJ7RhQI70SmBOdIa8ozBh7GPRORP0cWuo75wdCAEB
kpOY+VdA7qOSYA6Ptkv/39GCCbrRJIIuoKxuDumR/ObPgTsSh5ptudBCv2WxUjWpIO5t/HOm5yVH
ea429165L1LjqmlGCjUVkGdi7ng+IPGTtAuqGPWOWIyEQ1h2GCiQ5R/w4ZhkzSyOnVwRDSTntGJV
iSqRAM8G44kdYPVtqTeX9k38M9lCDalwuXUKvwzZz3wPPJGn2wrPbXM3EsUtMxtdsJapXfVdJJJV
wV1sLUk3Aqxt5+2O83tfcw+yIeCnArvu+GPtp0+boNKCKNDUofnkAwAw3HjO5/jTcndJ6fr8PBaI
lgzmy6Rxkzjg6AUEguH8oHR/CVTD/K/uLllaF310Npmg9GJSMQzN7yr6XDWBuHutw8w6yA2soYGy
VuZLrIh7OgvT2MxxNQk6nBHB14DY7b0ZCcn+Lw8URDiUg6C+ltiriDmvZb/y6iINQvaP8vyYbiPT
ZBaphX72YKwZXZmDk28QKT9DvD+pZG5lqi1X/ZVDstSS0WHQgIC5MLIWa80TVi7vqP9veFL0agMR
WXQq4t3+oTQbzp3/7wZf5nBCNJBvmgtXxOFEYJqOx8c9FfKOZZf1ZELw2rmGLSYzHl7sgUnJx/f6
2J6iU/wTLOyT9bEJ9jfio4HYXQIbWwq6Jx3InqG5KPTUzivSqhUfhgxqaWQpZ/lJsMP5GsLpFa/a
+RCGBwDhYxqw6U6UoLYUp/7yGGgS6a1iY3JHOm8Q30kBrFakNAsfRInOViBernZPGT7zN55yEJQ1
/0fCza5ya5QMo9znHpfxVgu96Bot9krrknyLcApaJpZT3LSBNoJ9OH/beedHYCwZgE130M+tAZ/L
NAFoSpNolfAm2cbkBjPfCOuFSswgLX5mUeUZVPdx/hIY4BirQymRxnoNfaqsr/8zYoipBwPaHVf1
poiOxJWyDfFxaB+MfcwTlBUCN+ZllzV84ac5pTRbEcpz5bRKhSLaYHKuwXbDlgK7t6oXijrSpdtt
O4/LsT7bsqUzJykS+hJmqWlsy8WY+VIqedUosVBJNsC7PKY6D+6dk+dqeL+WEQkX0tgZEwZ8JItP
0o3PCcc4bOhUeMwscVkCIn1Gc5H6qQN5y4ZG222xnbuedd09JdA4fn2DjIQ5VMAGWgXnJJS531OS
IjjWSfrE+3PyytLZdHOKVuR3aCkz2vO6IrPsZWwoyTP3qOKwCerNzfn60Lxsi4vXjaYfARSf8uGN
JMf9BoKcMYen13vprEO9Ghu+kztobS2LCJcCd5hRhufWTljriFIC+KQjYoqG+InNq8ks2Ze136YL
6YNGjSrajPCotkdYZsVcDA2NVO4LnrAjLed7axehPW5wNSZP2GYSFzBlse39Y+9BgCs+LA6dUFHO
M7NA/jDMwrg3OyywHFnUkSAMDbNNfhRSFYNh4q1omIU7SGi9bPp+omV/0cOgHfhdoSK0ymVMvhhG
p1VuQ2Q0rvc2H7+ja9HJ8ItTOuM0PL5qIwZq6iMaX0ChJdb8xXZ9C1ObIreEcBEsQxuhtWsFpCyq
EiQqXwq6cf9KhJiAP8d9khh7YPrzZJrQe/M6wDiZSqJ3uH7lGMePciUtbn5ZNa6w8r21535oOs4P
xhzCPBskxvR0+ErI+i3YowACcZ7T0ssDmDwVN88QqA8mD0QpF8uXEkTo7KWWx+CO9fFoLy6KUCgA
DcvM4sLD1sOjrTM6JV98Rk5bC4MxIo8O0LDjMyWhVmQT0up2UVzKJiiMC7gLL+p12Sz3vCutVpIO
PaWRcE0Y2TvqTuY/LW3YsYrf/xrv+d3jpm7c7WYKE4HmfHpzI+76t4Mp0byIMBD9bgGOcVF7f4GR
n9nqJeA5RM7WVRDCZaKiK3+42JtXhBzRixbYDjK9Ae1uNnTy9rjco67X25+aFO6es6mZ/EEUJEXI
2x70uCZMLyZ9c9j1FwW6mfI+lZjusTSQgmYb8c0hTU9xS9boUJ8vc7N1RleZ6gJRchnH8ocpMbJr
++9phDy/VhMZjdxu6kyYCQg6RGhpxEB5B684cnBsTDZOsyGd4QZH5inCWGCvAvnNT0Ntl4bSqZZl
vqrYwQRC7yLjFRF2H6DY9l2uIQRPI91Ws6dm89Rd7vq0KcShbLVNj4COg6S1jun8cnh4mJYT3pW/
3sbEgAAJdMeQ3gUs2/EHXk3XIt7qX9BRYOph8Vx/Gvm1JzHeZteO1uQ2AoMjnPiHcsas3b2qU5bN
3VUwxRbu4iSNIYI/XCgwnPKQLt+5sd8oePOE3pQ/XeTIKnztvRDu7lEq+/dsfG/DL1xJ2oXYGa5C
AHMj1+PvmlyUvzp8BCTQOCnq2zBq9HDqssusv0ZWyT9OAElPxEMuuKJNY2BHdL//t04hx1zOAUBU
zQcht0wEJdmWR7jIlHe8rzC6MvYpQ7G8duz3tK+Pbb828Z5JRs0URYyveT4KHjkZz4P8XtGHLowl
wOAiDeD2aTzOxRoVtchITP19smXNuUs7v5sVAwf3pOAoDSLUK1pHs4WpapRC0kWVfka+JnNOimk2
OfRCJCigCStYLy1oCXlyUr0hmOdeVc0+VViLlVJnoi7IcBen6KdMq354KYHN/gE7ZFUA9W5DtYCe
ywfzch/2rYPFV8tagCptKhE+50rs9+HRaMegf/1RoR28+KgUFlxIiDjetPD7pJW4bRbsgI5Pupqz
5Za/0qmByrfoxRMn4e2EcHA65XX2uQ9aHV2/DnjPwNIcx7LLMzjYyD5KyAaQanu23vPOdMTi6FpA
QqQo/tck2lSlZjzdKQfUrUqITtf8t7ON94o96Sp0brmO+JgNfzFBXtmFV5E8xDgembYMOHCF/c4s
04U52tr1sZxR8R0FuQHxU/UdQWgqeSZ5yV4xkVUsmKeHrgu+zmLjLywX3Y3Mbe6pmKYxXLYiG4DQ
bINOLSk21VkSvwpHgau9Zzo2+HXBmB1QtQdsuAFLcEAvyEBlEI2uKQTY+u0jMgtyUwG2RE+fVkdv
ZiQnEsQhwD6Vyvw3j8emQh+Tft3vUlMq+yneT7ssVj5ELFf6zb5hjhTJRcOyc3tMi1dooGW6UsuM
otz6lEEtU4/LHtqCV621XAeK/Io9lkWhS29QVdoZRah+JHspjXT1PYjURnarcmAhTkUteVVbSjgH
iAl/R4lxaNW3zlwgiJMdH3AcJvyFhW+OR1wK2XiWd0Pc46zwu6YKdfw0HqwsZAXnR7s4LosvXo96
1d/5OzfV4gMlJTaSBabbnqLwaZp69VqMW+4FIZRX2ziAjtBgEZIA8ESYAGEGy6ktBwDSoh448vjx
DNQXUKN4MCYBL825XJBKP4kClV+RG5J1ceSNtSZWelaFlw2Hj9UZP02nbvCoWQIK/AaIiIhMN+lj
keSttFq9HIfLMRvNce4gOTHicyPdV/z7tHymYy+xPyR0yuZtWyvzgbyWIvzM2RA+It9u27/oGaPr
2vpoITKPeWq2gT4ocMr3TJygztcDVirySzr31ZBtxyBvySR6pLf2eoyklXN97ue5RjSPqpc88Saa
DCE+llkHB8YzAsp7yS2dQPL2hJ/eBfyXCH8LWsKQzpjhTJKOQUq6S0Yr+ycO73JdU6Gvoq09Mkzc
qGFbGN5+HGlIqjkT6ew9pTbFceK889/qheQ0JL1s61jPR7KdxAw5B82i6+6mXXw10/lCFAJNa2ns
xAE+5LWlqhdP5iacVh8LSqpVfRSGz3jEJCZp/qBFzaDcXdX1DBxuFES3vuQKNjYs9l8+W0RWgttN
eDmBew60pVz33f5SllhcabI9o7UlSuAWUGsYKqVvRVhJ0+CA+cRbiW4emCR2POo20Y5WUuUKDFfU
MixKECPUkbcqGtGWHHDBrAe+m3I5Bn6LspToWaMhXmt8eku6h3qFtPbFduR4CGPhqVbUDSp1eU4L
vBg2J+x86wgUgISw75UvWnslcP6fApeFrcIRL5jzGxH1G9/aMnKLyMqMBF3SwS77cz8W+56ceIsW
NcwmkkRhnWaBvuN9u8ujndQ8ICAXtAv9RdvAiTitt9tOUXcA+aPfUiw1Ajj69RQIn61qO13FsDbA
3lA1DQZ7wU5s8XoYvlq+XMP3EfmgHM2m5XORHg8A/DBVef4Pq5yrpIujSqgr8Khh9ORoIHWNIi7I
M/uqkHcx6V76HeDO5skxSKeB3mUlmcdvLhsfH8aff+upjafRM2QI4w+JX9rOitkRxcJjhjOJK46U
rn6xtqeyUmLxWx9jMzpJBPIun+ipAFnRpr/ZQU27gatfbREB1XehouCIl0LYl+sUCkyKLyzfz4C3
qxlqETyshOIkrtVXt/ZI2SrbKr0tHxij8N3c/vnZgOGEOcZ32vSpczD0TWOGdIJDFp9LEdTCa+Li
h3Lu5pPpDqC0mnN/0zXrxvK37mD5zHHB22GoI/L+ST7sHqFmWFKBnaF+SNH6D6UZPMBXSuxjjEDA
+UrN2CJkLgEsm92ZeFiGcfDiIDqHrpcavmX2CIUQmIVOrWcic29RSdCWLu+hFE407dFDUH+9Ac9g
uFAayfAJ1OKjDjWJG/QWL9PhYy/6Thd4CRtjy4C4LUV5jY0prxkuGUJP8eLDKRrbm/3QHtPmQgrM
SYwa3taOZy9KOuj2QGkqeFqf53THKTr5VY0oPTvRl6Qt1ljOj23wYrHvUdpkNCfgb+JOHO6ysYDc
l8Ws8lrMlxvQW6OOXTCg+HBsZk6Se5GiZVvjUtCcWN9PHS8rwF+gykookKikErTfu3sMZyyoPXDM
rFcXnYufjXhORcDHpfoB3RYB74xmAoPyL6JOtuIlgzGwCX4d5yMjdR5jtubNw7+hbVzok+LfEN7r
I0O+TbN2eoW4B4G/OWWhkAn+nZZw5TMnB+kfuoF5OewKrLPIPNGGrUn05iGKFGG5tCG6cLMZzOMj
4MS/wSae9RG6lUd6mibP6LagLpOA4hOH+Qos4B19Avp6puLLCL7ETP06XQF52yoM5oVHjb0UkXV5
3kPZAxdKbTFRUCIYDjtGVJHMpnX5ysnO8fWpxxyUQSVkI1pEhO/QN1TpmyvxI/bND+Mn6CYZQLi5
ipwE68DwOoxfeNfivDKEy9eNPvECSdtZHxeASAgbPbxYNJAkG8PsZ7WqeZUNRmCvduqQKeqGICUd
Aobk/BUlirTpGKoPu+V4NMLUgveu2m6iQlib3IKmzXQWRcbT2wuY7GfcjJKQWd7rpBKQg6OsTOWN
D6+GXeMAtPzSfMFPaSBteauNhdV/VY/8iZhn5UUuyiCsLRzPAK/xhQ8IGCSosuACLlU86vdbnJ8i
1KBc8L6OAAP85wDES+qCoXU8LgGvTpitcIqG5nGCNAmAg+Een/xwSQcIwYY97OLhuoE3ii6mG9VQ
Hjbo/o6l+73KVoOIv9YHVEX+cv/ooQbtJrH1D0ILiAn+uORP2QvIHPVRzZbGfXlhQg7+tMqURbvY
nETgek0/Bd1pCULNhB0lSUjXhQ3VOAPDkJ7t9lCv4jxcOKtz+HT+UwMMtyZki46VMeF4bNuMyqrr
bwXP+coukJVgoSM11oy0XvpoxWMi9TH+L2tF1uKJkNgfk8t7WSt/WvAy6f85wnztcc5Iur3PxLNL
X90BuzUEC7xuQqmgwg5WGSIgp/y+JRRTJz2po7qGM5K4U/FbdFZkn+eXYVB9G+S7ODZx7CcWv2a/
7uOQ/erTKlpL+KzPeCu0hLAQfmCc26JUplmk0N2jOyWl8UWmbE9ACjQXdiSAFm9oOSPg/xsZu8gR
H7GMEcLCsQBKPFAbh6itcQ5R5rm8gjzYwwFB9i4dO+5uXSaF+i4h1q7Hf57oL4FN630C5HVQVVBe
28i6HTU+0lzcrcGTISZFj8ktQyR3nLyxwQIZ/rzibfiOAqWKOpt6aqH3VPjfUtdzrSKyP0orBxFN
nEtsXdhU8XxFIBt6KE+jxMIMauW9IBl/t6Fx0ufaeqqUrE0lSyNY5MTtQ4WMRT2hH4MrdJKhSWa7
DnJVbItf7yR2PWpIiQQil63IkdfdmFWy8V9uIdz1a8q92bDYkQSHERyhMb+WDthEnDX13kPPqf3M
cyqSC37ZlyPBoYdlh/551FaT9V7x3SE1VDlV+gMg6WnmU88TO+31l5darDpU88S+SNYZMLpofRJX
r5LDVW5Zfb9aE8LvV8sS7s7ZIgrhHS2RG1l8B67Mhnj/kxSDS3H1zbXo+3/s8vvx9QY07+2UNA12
T4jZy5vhRvxz/DhIC7qh1qykuqhZTh/btR4Dxo3y40ahVoDgicWC/EPXE/VCEsDToimhaAVVjD+d
6V7BeEdji3e4osK1HzqrHut9X9AIrVKGR4GzNTC4tf63wWTtnk7G3Zxh6ayXY94Awnx9zt1E6c/i
9DGHtdb5ANv1KZTp2gFEnUOrIkl/AIp8xY3mvX08iHuol38wwUdCzzl6PQlIRf/Vu9IM/ITM6Tlz
pwSxtzwH6bUA9EL5cFEAWp3buoQPqAdUWoqD5L/2QACzjzMz3LvVJIN77GAYY92Su2f+1aCzOjd1
gbtYe2m5NDqc9ZDdmGHE/UUjv/pOJa1Ku/z2gxaatL59WmNkFXaY8GwtX+fuxvIZBHw/da5yvyyZ
sMfnRrjs5RJLGJJImXTArkZCNpzgDtaAtRa8FiRd6jhBDH8A9VMRU6WNgHKc+vEWRZpZM8vDQCN6
uIpZusZrp6ugR9rTY1gp5X3e4JVQEAvx5TAsePdwHHVMUBp90BxkCZmhEdG7zUeAfAVO0XPpWfCZ
jj1jO3rfuGtNwrsfHvNF0e67OdScKU6pQ3nFIxVx+0WHOU/sRHXLjt6SvIrIdjNRQOPVs6YgMo0y
p6kXOv8XCCrlrb1NcUbhF6zFKZK1rim3O6Ji25issPFsDWLTBT4f0I7sfeTGqlKIYhxbp8/wp91K
cy/cHNDULKcEDtLlEnf2SlajvF+oWxh53SBGZ1wp8EyWYUwi7ieeo+WLyiuU6JKxZAZ2qji2fOaT
FAvXNoVsyXdAC+o6jDtCWQ2lcYdximyp9mzBJk/DpzMsR/6HPwrhcBDbb6sJJEWJze5ybABqNPne
SizoG0rOudyc0RrKGWyfO4AfDM11SqDsdf3NvfGoaRkgT45qqCjIzVEdNsWfkQVHWTbny1ptRmPv
9YLd7qAlOcsYeHoQTrKmzTbwZlyDM35EbVucy7dfxu2r+0qccEl8yPDCRzhJAOJTYvs1cEm51H/v
rymXqO4XEJHArng61B/FiFiCJLmdhOnnTCeO2tq/XrnzyUTub/BcYOoCBN95GUTPdt1ntvKNcfWO
ZdPYb2zx9yPd5tcV5dWV/F8kdHt3VIa/XJWD4uIHwlyk79OoB6Ycku71kB+q/cIambrXnQpedZNi
CLdeDWYMPznLfxMx2YKxCH+fvTorvVCRQ2lIDAUI5kvHt4EmUPI3WQHS76Fv7D1Jykdw2XTOThVH
5HiUEhTJfX92sMlnt+sHIScafbD2yvJ6XLIOQBMBsMb5pAQ7gKg6k3SKCsX5ofQWZa9ogLQlIS7k
+RcCYvLPBcEVU6tgMi2usZGHpmpuxPRq1oK6H3v8KOw3dsKeFFvwdH3sTZ/OQAvua/xwwpr7vqaA
8V5E+SEFc+qlhYDS3ino1clx0TXdJEWndiFXxSvsQxU66+P7qoahxL/pommBC2boFSbxacf3KLCV
dml67W0yUMHwBwPF61+uzLmF2peafa7AWLTxqX2kqSesAxLVig8pEnNNZpN81EwkAFi+DFoLVsEK
3uQiCSesx4aUGhFHVmBNx67T/AQK62tYWUtoMFzv0ArHgIZigbSU0OQkTfQbTVCEeBdqAASuc+Zx
gLYG2winLVZD92BAJnm5/TSuGIAIuIv9i04MQ7v5dnhiWzdrzUMahTZF8bF/B+rDzWsyu+UhES/F
R1pDGUgqF3iaDis5qUCalmgpPhrtZ7Lzkcfj4hxvXxsvteL6SmbMjjwrDn2kc6R3VOzSDNU8umJq
O+nG7xTmoyyx7dD8mqYukmV6Rlyr4U1xbtx3sxydqAK26MnKWZV8VT2rCGZWbPI8el1iU8NN8NP6
H8YghsvHeJ8qPddAzsfg4m93LoUhWjyEkYAowmuHGhNZhA1P2t+d4y3DAWQJSAiXZGG9LVAU+zF4
tn70GgacrIpWXMonvRdDgBYp4InIY6PLQRPRaE1n+V+0OWvBOwFQuW2agJCRn06RYxpBy4Pj1CnQ
Y/ubszqS7DpNyH1gqR2uVbEKNIJ3QpqJ6YfyifXFR9vwqDCW0ksZIny08zGX42fLUT+qLW0lQRDD
TGgpnlgS8HW8+lo/GmrfDeP4t7v1476KwSUxuRotmsRNfUL3BI01yQ9oHoFxjjPFLf3F/9ol5HtE
Yl5e/K7RJtmVZMUwX+WokbSXWbwomeAzMJvNK4AkwYJhvzdIN/b1egDY5IuPBPj4hYJDSrUI60+p
yHb/yjD62STU7dTr8axz5d6FSpMNRXaQnAHtZlLqiSAFH6NwHI24YAlrxW47GvbZuR5OFIwJQjE+
NykHfqSRH81OhYZEZj8xiVvYnNTGU+d9qo/TZPbJlFLDvcaIImqjNMtQJO3HPNwl64/i+YWfsSh8
Nbwu7Ru8GdTUz8i5tTGgXKPNKdSZ17dIj7HQQTnEQKyP4XmmsLbWTu5K+cHzYhpRoWavWcItuehB
FSKPexM/OlHlvv/5+U2jM29gwfa7rZQZzHiZRXguy6VZZweW6aJ8/kT1HH//EegVjckjD+dRbbPk
V8FEoBSYfpwjWf7bNqTvQPXru9Y2PT9D6088p0gdQ+R4RsXWqsnepF5OhBsvUeveauZWL8qJBlrT
zCAW4jZOOhkJmSS0m8PjV47uNKWHqonTOKQ60klcZAS2bce8QSb71LmfF/aML4gK2v3T/KSG9np7
j6f9dOJBVNX4o9Q1GKsJAUlUm/7w/wIIRXp9hIL7mvzrBXUZwtoAEdS0g2TnqtbE8iuiz2aZus3F
0LZ2pFqYqvlUTNImq4KYzomoICYhMF5TXItPR9fRomEavwjv1ACQsdSB4AF3Q+FoHR1nujDo8cV/
34CouT+DThdDpICpZpho1LX2WCLCHJdB9xWDUXbPg5NdV58zLNc0Ye2CVwfXivi7GGrmZAAKQ78r
do7Gh3mf5w+vDHPBcz7pxRA4OmHL+Ls+G931W1n/DY3Ue12VLtzZWQH7/jWXwt7A+C+44urLewt5
+vNSeCjnYdbh161fgqHm4o2f4eBondc7oIw/i/U/by3OUpBFo6TRYWxCFmfo0FSPY0vhCWGVxxyI
YU8CU8Auqkh6vhsNV2zPuE2E2QTj5yDJdmdbwVmDue643icoGnrtvQiJA1iWChkpvMTvQ2bq0a6x
shTz+/8lU7uZUdVGZNrD0DFi1CkyBBrMSESa61Hi3WQC+LgO/VM4sqbBg/RYqQNNvWvL+jH2+/kL
Z36/pqgbh9kpxPtkJsDhrfUHUe5lOm/7HLbXGa0pkL52yI2V33oLexNnTqQet4LqMs+QcbSxK2+G
ygS+4ICex22hsEiC0j2/LVaKEx05rk9IIvet2AI5/aNw+R0yNCuJN5SaEkVXNoXIw7URy+lKnKTD
qrj7zRPaZMCJ4C743b4yR5xRj7VTH0oK8+qw/Wq/7zgPeZ9olTkNjDEfT+aXaPe956hH2Kk8t6yk
JO5o8vO0scAVnSWrTMWvPP5lNkhJHjkY9Pkj6PidIyjJmAQTXytQuBJQ08sjm9+TkqeH5cuFd9Oo
8UmYQcu7QziEl3FRVKRjHZHLGA0L2FFn8Mas65ou50deThb11lzKDv2kNSS64xtqJd1CNk8hFG3P
48FxiG0ozSWUF7S/Snk7yGaptoQFp1AxkXGkYWJ0r8eMzKcGcWb1QIY4CxbozgZlMImo+16OCnu+
nJSXiZgNAnvmYh9ssKCIn8gis+MuLyqosraO8bUcZHAtbAUKwrSyEBdkUjgUX+fYrbxsum4QwmF6
g1s8RxsgYopPMX9W98cZgfcNRlv6pyLxe+m4ddbcojk+9rafTpsWYETIZ9Jk3aYOnaRL9PvzStF4
sPzSc8H/+q1hYbFuGL3zx6OAjhgMZkWTnlI5/VD7FMh3Y12IubdE2JGQjxyzfyY583uCs+F2jsMP
qnMYyqB/ZmfSZ2ghRkzPZSdjcH8H9V/r1gpGmSZfITrSRFswgBPnzP7M1L3/Fx4PL+0CUEb4zAwc
eIj2nVhXeg5gC/2CVEmeIOyMF65A9rVnahr2Qwfc+ZZ7BsKf8jtD9WkLj3CRgQKRSbwzf/6TKfRP
5sunYSdAA/uNQW20c3rzP7J7Le85bSOjXARKTB91tEQGyKwQn2k7f56JRk/0UHT3XBd78GLB2ixf
Stq0iClX0ahtd6p24lU6Knsn5oe2sxMjWfB6G+NpWhwrQTKpBiZKDYw9ppWPOVYC34O4QQ5vhJPJ
0KIcRGqJO4hRm8bMVjWThYqAvjRdKpqYhLFJqYuMCRLfUXcBO2R991+EyOxWcKZINoRs0PK6SPhQ
a2mawEGGJIzJjTj6OniEWAJqSK3IwpfST0jIDpxQbHxiqw7uV4FQuyTjOUoNtTu0bC4cBtO8/zSZ
/uMbn8eNIOiwZmFXKnqbxRaJYslqALMy1IYb7bEjGGrg3mPzb+h2AKEKvHQU7dx4PiaGwjwh7Qt4
PI/leg+mLTBkK5bP5533NL9h20Im9sIEUPFqvUOHS5AmALQDR30J/gVSj3Sg4UAJaXzZgVdPARmp
XRyDMzwD8+LxCDhBdITXkwmdA7VIaKvwJiI+M62ROnL3qIjeGUFHUblPtW6pY7tltYlYTKQY/0SN
Eo+5dg9pC7PqCD1VzqR+hcO9QF871m+RPP1EQ4S3/zxxNLc86U65E7OzyFLa79EjA56BUwsUqz4C
RmR2xajPCvyyKtg3IIxeyl2v4aGkxwJIJhepTP2UjBzo6N4wRgEZsPEqqPPiqlg6wMXeUcUDzQi+
N6KLTHjp78B8eObQV5hUl07UjtK1t2ro7OpNY2bGXON85DJuKIROiVnnxotXM8F8qJIwpuk+FnJn
/1R51SegIqmOPuJHJghfAXV3FrpdOg+TWGiuisNySsDXfXerUzvg6Bn1AjIf25DrE9eO+p7htSRV
yUkOG4om7ulMJNNEGIJfYj3YUYS8LfcZ3rMeOyIfMCmaxT5IKyhiH5FWZ8oIxNJrtmRgJiI5L0BK
CrQkhxtXjDKlOrDDHlJKuH/sM3ZYO6qTWmrPYsq4c6Zo4nkggJJqdwyNcZONNgdD5DH26T8KpWRa
0hWz25Znwuy//PGbUxUisyBsa2pXsr9gZAMSVJK7rwXU17SYv8DLw6Edf8WEtuEKojMkobAxsv81
DB40TBANBzHEf48AiWVWNq1F6O0/HasAHOrwuKLbYXmXzWC6nZEO9yqqV8j23CXXWFY33nMHTvG9
kFvkq1nPvNUtdKUGzpc77k3Ss45j2KusPBHS1BuSZwVoLZX1x3BrV7s6f4xd0n0uwgIfXYUw1lw1
q5mOQMVpdXzv6VsLmkGpmTnmZfBjxUJNJda4a1cPg57NXjMwHziyKZk7lVJe+cip7YUMO8frxIKP
dmqyUzbwsDfkaS7yfHnmyuWwVi5gQdKCzYv5c+5WBkAF8SnPrtQepk4gN6eE3++lWFqq6jsRm3JQ
QwtC8ciNvEYWZ1FbU3CNfNDE59h7rg4/JyffdSYhynmzcmYLVu4cESFdyKifKTp7d48OCEm11U9l
5voHOQvAEhjT1Rhrk7tAQBocETPV6ckh/9IKvLSzQd81nDVxHJXyUXlZTArxnWiDv1f36aRDATCJ
B/WwxF5JTdrVT7AUoxxjp1QAiOmNBCQi4Qca1x2xG67fAJghTx1qx6RxahEnkRRExLHFj1Fs/rn2
/K2I6U0liRKil5aurV0MGi/4RmOCWUaT9kLi3fdpqDaFawTNElHJlspvNDTbgjjX9OVSCoq5WBo5
4aHCZlKqgKZQgYG94gJhU8+OPWlMCHCpWAWSK5X/fXcbfE8jlk7vpisjePQZrEfuJhrHurZ1oUMf
T1BrOYqAE4Twu8jBi1D8vM+7qTHErQzkpA905tKqYoPkvvDULxIoakuQVp7b87NyuKfvjlPgtbVy
pbn5FMvyMhttTa6qhUmAH/ITTS8Q4Y54MZtZKl76uAONNXxCZafg8wdvQCStsKa1wtWYuRhjcC9Z
uULZfsj7+Alz26wH+7srqCJFTpvo1gDINJ042/taALrDsTGBPlJfFmIpcL5XUkOAwTSv2wVjj8Sq
KcgoeGFYDHOc5/tKenG11AwhJSSmLltOLwdTftosIA6Eq9C/SIxnT22Nj4O5pEusl8lgxZwMeOMA
HjBXZtwhop1QGb2IQU2ihDGNZViCfLexa7Fzcty4PZQ+SrS78MUnqLtE4UTsJziFdWBYFpJoYxFX
SB9NoUO7LT45HNDVXqLnmeZlmk3uEjI59nI8MWLyOcJoKHDGjma9zAjZKh9Wv041NrZ5YDqzy0gD
se2oENM3YNOusTgqK0heK00pYLyXi4kfyJu01SW4/vLQWnf8zknIkmkNXYUFMHCn6tcwRnl5sPUD
I8aRybZ6JREQ/IfqUzOg/aYOdIOptr6lgYyBN7TW2ZYUkwbjaCriPxVFkGz8+bmFn6akk+bZ6QPF
tlZ90n18MS0BSuCtCFAAy+6apqtsTnFO4eF30U8N2brV1lQTIWEUXKIZMjj9vvTFfn1OUuSzTId9
F/BdMl3rl84pgDlROEI2gT5izNiO4Q6tOVZt488hHbMJYAYeTmKtXBcCN8n20wnSgisk/nULyO5C
mcsP2bt8oUQlsKt2oPaR3HgOsDnuYDAzmuIaV8Ndt+xT/CsQDH5TItRBWoWFkCRbn8Z6JdcuBCaB
TpODV9FXx1cLkgrOC0YrJfPutu5KdIaSC8re0ptg8CU8CDAm9Bq4JWz3GBsKFf/GKTVslH4V9p+e
/fRD2+M8ovpq5lpyVNj6TL2DYtmYKbsF28coH0PxD4f4/1nphaFM8t1Wu574ScTqHJbRNcvyfUZ9
QqiCsXFSb93Tckikt1o9csRVZq/PhzA3OC/NELJlBjOlnJesZNhi3oOfEuqqzJROmW8CG6p3MPsn
2EzcjuLl8DDhZ5bv0U8c21LFZEUio1jW/EBrqjkLSK7TSin726KvgnEx5PBdWKIiLZc+08FlOpCM
X6QF4bzl6y8qmGG99Hju3RyeMRxPGDi6LMuXXWaIjdqJzBFKZvU/DoSpWLWX7AW07NIQYI17E40P
/26/4SmqXi1o9iUXD4LJ4PJ0s/IpbuAkYLcx6/pB6uomqtwL1m3atx8vwayVr7CvjRdqgmkOcdsR
tlmyuHH4/rXT4+mjJ5Zk+v+hqjmrMbreOsJw3QsOr3MTEvmpUw4LPX4e6hOnq8DQNuxngUD8A1RU
nW8G1tgHjlC6OyzESSeV36nfPl8q/5Kk7bVWGiSCbbcv62UzCj8SoACvUw9Dtq206mxBSMowGkaa
hnE9DJeidoBonsxou42Fx/UsziAB4AY5os65PTR706Qeml1Y0w/8+3imn1qfHYPPDqna7wPmE6oR
N39cK5JN1XeB6F3Tba+9izl9shf8S+o/1tzSJqR64NbkcAgvLLhS+zkDFzproqRnGVz4ijjxQtcC
ihOMWp2vciADh22/nZhHYlMhbS2FmmnhrMQRgYLs025wPh3dQS3ooPklCh+/sm4rxV7F2oquhIcS
dXSLoOVEB1eK/IpRykenKJwiZik4OEpx4e8cVB6XA3zQB6MIQwpzCdokHKISJRSZcwmEYRZZ7KjH
xRlfa6lUdNhDraJdSoDBZwF6tTdQqW+9ngS/D0AP6DCsBfMvaxW55wh7nWJwYx3zUq6Mdt65gK/E
WcD1Jr4sFj7vdwHrROFRMp6WOp+9fvkj87bt6Baxg5H2uLUOwgGZinptiWipWY8XTG8vp5QFVR7F
JTuxbgH7QJVQXueaqir+4CT6CPmSPuKeUc11H1DdBd8V4ZC0ILlvBzLxIoTB3r0xUBLQOD49PIyo
cDyd+qYcXetH9y8DwLofzNP8esVsIewY9K5XaEHWzJmOl1uzfel9oaSUhANd0MGiXvAaiXkI0KMN
n+c10US3kJ6bRiEH+q66ttqS7JJEJavL2UX2oAzpz3cZB6Le207ZrMdSxFB64AF84k8oB/YhhB57
FIwoX/sc4WbzvkezL4jqTa+a8e0nOSsj5QmULyQkuqxo29cmrHodZoxr0BFiCQyhDVi0ppzwFCtf
5LtZSIBBPSDAcfman1qYoIFK87ziMBIK8mufliAY1bZv57aQO3xnUBurzNc9M4u7rviAMViTlB7s
TdaaSfDATfaWXEIH5KObhtz9BhmMfbwTRT3hhmvd0VpXtGUie1wffIEoR6isw178t3ZEiHxun6OL
GUUJ2fpPaNNKHQTd0cvZbOfP8LsCy/J4iVAjrDTUsc7MLWUhhvGPnugdHCfsO9V4sji0cPQRHUhg
58e0Fd+QaaXh0LzJgQ3sT0XX0IMV3n3djSiEslVIrVfEBv7063FAd+zt5SypxjHHz3eAeiH/ADEp
Bx4TePCEaHrdQGA34SAUOwPwV+3N5XN+g6myVM9MlIGQOhEBubPoMs5HnHbPQMiPTPlr4ehlU++O
Y1cfSQnLjVX4C0kaW0MWIwEJohQ34LQcnxDxxDoFhyVYdwlimwgAdhXyYtb9mIfLkA8O4bARbQCp
UB8pM6s/2TGrF3G1bCtsgT93LumbATXcnq+NGdahYNt3FYzA60GpgpQqjF1RL0lXqp3fn20z8wto
GrC1qV14VM1Seoz+Cs6BSwZkxhm/UoEbn4GbsNUG+LoGdVP7PLIUUKmtjv5fmqKoQYgRXyZS8XWz
5aODO2EhlV5DiwWeDAmO9a6I7J351NQFhoeFKPHbv8OuRd9NUWWtuufw4Dy7P4xedVndGwmGK8b7
JVOs1fhLshlVPP2ObwzBKY48tm88CyX0T9fxANpCPzm+ja9w4wC+/4IwwH745M63gmIjL1hf0Wvm
E0GNzqplQINAmgh7w2wgfMC1Km26e2zw91yso4YkurUYS+6DL9BHw1LiXG7rJJVEW3kl6TnGdt1y
pr7EVVb1v95HKVTpDZwUMlwQtptd4nUoq6msX/fxY10tl+0UplkZiFdQsrr2uMpa7hP4GPBYCRum
GDEXxaCGGNqHo+t3S+rqWSeFuhksMVRHShImgriE/ajnYvrLPVDB3HEfMNw7RAa0iLmzRujdFhMt
4rMYwd5DTB8MI/wjE0rgOu1BNZRGkdjxKFvieiC12hBhrrD+xIqgAipU/RvBRpVSumKjuZBCwyEg
mKcSQ3E10g8FNawLOQZixVDq6jzdVATJURHT+jPWoxUpNDXAOajY55H1lNYpsT/fuMKbIlqsugpS
t+exKEI+NairEJGpwUH+1oPIw+hggm12F//LzzvnFkm+qyQTpqnOaLeG9WjHKGP4bqiYUj4R7kjk
Tz0d9N1eK+HfxpQLX74bBIhsjerynkgN9L4Twj7xBfMEkAwWGgKRspXIm8HiMxVuKTwhqlNMBcYs
cHPZfpqjMjq7zMOPuva00wfnalrbw1XH07kKxNzxBaKkg/DwZ4LQiPS9gpgcJrPIJBeKcnp5Lxfk
bbruvRxeq+eXbODjdZwj/SJ3EJ46GwrTfFymtPAZZek0CvA6ZWfMV3C2MMre7UunwPFWfY/+Il+E
A37NOZ8aa7kKVBq/qsvqE8mgAv/dmP5wQYbiDMKBo4YI2a+BlCv9MJzNgEdoDYeMy8w3mq071FRz
V7RsxSJDhOwPuwincPaGQGNwqBgrodB5vYz+ltGepms8m9MZEAwtpi+Bs036bx1HTCwkveCtYOCy
IQfmzIxaz1EoZxLHpGm54DzDTbzFuIPmmLztL2TkVLd+V9SzAxREp0MqCMzfbauabaGm7Ej+Pdtc
VHnW7L5lXJ626hsK/Vf+ri3sLaP2rZuZcqC0+j1sHEJ7eEmBNPAgE9+lP3QT4BUb5eQoYDaOGKRL
TZYaKml7dw4++HQ3AE/S19T0hq9X9Hr+bE3u1DjEgDOXBNUb/KeM6MGughPuzKxQznD/cZlfOEjV
xiBUUtu4EPPVIHeR/wSnIX8PO/UdbUhXEOYtTNuSTvFL53UphfF6+MInyI0jS/tzQHWwKAobHBvC
VFJtQPCiOgug7boGehmyT/kWRGKMbCP7Y4aaqUitPqAFdVzDEvvgGDQbKVLTNiwBrDBXV7OB5/YF
XcvTYaMWHH1It/fo4rKxymmW5FD04HwNdRgr53uD0FR4VUq+cvx+2tXLvGEHesCBDSGPnKAql+m5
QWpxPdhddpJoy//KI6/CqU31b/39uZfPFrfB4mBP0hxilb/5ZDwPCrFPVxcEJuO1ZN4CTWq5Cg92
DviAtgrvjTUdhfoJ34WUPTnx3Njha63uC7XULuiIU18lLVqGD6Z4JxoCeQAHqm5ZRdcTr6jsnTp/
arX9RQn9BlCVQ9tZl40W/ec/kTcUJm1d+5cP05RXStRF0zpL9BeXq6Q/RVwDlJGsYbQ114jW8vQ8
g5MqyYD8BR2wRWvyae+weibI2PFlh7TN7Og2BgUFPouTpmQ2FPH1VmfLbmhrudjNCsdj/DPYUju4
rsA6Q39YBI25ZcN2OJOSEebNN1htROjy4hpaGfp5+bsdYUqlrslquL8cRLmLdgaLCyh+boHIZ56q
AaGwrTzwbyH5i4/C8c0DOfif6NKKx9wG5ikcUhN+leO4quTzc9TMwGLg/IZVcBu/cYNVDWLikQZY
tYqSKXXaJnW0sBtOoCZuMoE7uayfdBQAn9OTfOVj2dGIYdrEaodU1xRYzkLhC57WoLCfQPCK5HcB
onDU4N/jJuMBdwR8hENBZanPLNVZnrI7un9K4PaRlLqU28XMZtTaTNox2qOySHfV6IlTvd4FdVS5
+wLRB/euj2ztXbDfNqOc52A9YPW+4E9QLnS8i/82B1muiQoQqldkshxFbBBxoYk6QMCzeFS8sybu
xJjW3pk6sj8VFcTfLvN8Mx/KLR9G4EqZlQ34vPXIQzmStSgQ4Gmx7Idsx7+xcxad0whjgGKpOs84
eHlY3D+2TExqQr6qbWRhTnsAXuXG2Zrt3QYzhEPzdeh4rMgu86zjTy5Ox2gMU9LXZAISJswTJSol
jtF/sEA+WF9stJUMs8nR5bk2SmlbJCqgJ+cDuY8uMX438B2+8NAAYcvAwYBHGTI28cj/tTqzHXfM
9GLpmKT37+QbsM5PfZm6XsTteY54F/ZntVl3rP23QXFIiOI1KE4XyD93y29NBCV4+uKI4nXgtkIg
PcKywpeCnoJgub0NzH/AHmpY4XmAv38Dk36UOnueHLvYDJ17/ZwIjhn5vybNeS3CaORFVTsd7K7i
E/SYf4D2+GasAMqeWuoRDF14uBu2KDlxMO90naOCkms40Gv8hu0hbLkIwSXR0nbKcUPh+zksv0JN
GEgjDemWLEjUZp9gDjmN761zI9ocXIeT16/6l78RNRzMj9SgvuFK9fmLmLnibUBD70eiPF3M0Mzn
vPf6ouVr0QqABc+8M7spBGNNBgrvLQ0INgxqcWOUA2v0rpSIwL4WRo7Q3sBBB4IwgMfvDcYe1I/+
AP37UOOcJKXAoS24pz1w4j4OpPOiQkTOrqMdA9OpyM+NEDZTfhXaL0mH4Oj0LMLuv26Xg3keKMYB
CrEEqcNTGthhmMTitQKoUUsug9Q8kVfgtoG06r82qzv7TdL5JCicZdPSmCUONquFV77RC6jLEop5
s4OJHQNc1/dzK/UNQKhEadmeUIOplz9q99Ot4SfiYPR6paCgcykSWwk6Fw71W4yOPC6yWlXKztyz
EHgduHHeQAtGcukSzpHa8vO54JY0QOiOIZnPAyxWaQyDE9P4j32KrEKp4ZPLWSj+n0GicLjffVso
YoUTutb/5EWuAqJKSET2aNyn8rt9PnXSQXMgqwAm4e3zV6uKrMZUyicQA9zh+2b1jP2g+KSuCT5C
WMIlHyXAYRGCZrCa28e/L+fV8f32kDRXsrC9zoAdf3uw/IrNUld3S/hsIeehgxrE/dAAr1dToS7t
ohownZngtiCA+DLDjUIOZq1Acg/BEVxLcWh9ATyWpchrDv5mZJ18axmHDscLTWF2IG2cmXOqoSoV
j/MhLE6B4x6AMSndpsw9KvA/WusfHly3Rr5Tag57iw1UVkp0ocFghUpWoSLYPWIOuInw02eN1cW8
lCNK83t23VgGvyg9irek3BWl3vz+U5/cALg0Qc0wF/2heLtL8CLjbbVZ+focy+yvVOP6rrROGcl8
q4HYk57RgQIRMlEyFbpRg10DnO5N6tvvaKyT3VxSF9a0QRhlDUOphKKD3INTKeoDyDkWqyg3ryEy
U0jaQZ5L6tlJw5GEDrCdxDEzuwnfILjNscY7m1iyrf1OCetUYYa2qbCsCy6bPiDaaECtBO+RMmLN
FkWPdesh2L1ZIWEYsRBQQpKSKTtcEW31x1G5TCEtmTfRcf8ld01uJRrCZWve34/11fDwEPfN6haM
6e56yCzmx+9KEuW87QMaZTAfkbkO0BkMKBInEZEAO1KsbnvbfTbsDFB8DZQ0FIaQxZEfwc9P0sh5
W9rqK8d6bM/rOSH+HgxjkI1Yct1vQto9665qeEzbhTuPOxL1fBlBKU304p1yb/R3L0F5nsY8guQ0
LjXhL9f+PxI0cGdSKk2Jn/1PjogED1pTr9iropKNXySV3g7yqYS/2F2i0jgYHsqkFnyA4pIVaN+5
DtnpeLjATT1+MGNAnqPk69rPf/NbtSEBjbRSHhRMKb1dFJNR5RKgLAb8xF0YDt5jybEs7/cGK1uQ
xGL0Hy2spCEMggyfqIxuv0WaDXxwIPgmOsW2zYGcbn4kmeGcWY8MHyOodySNp9HVuLsU4lXscOhK
SJreBAhl81b6Oh0/lzDe6cL3goyOA3A6ZV9uwrYMLqF8wc4rSok9du4i//8XDHtSHivSeAZ5Xw7c
xko/Vj+Qys5PtBEU521BtmrkaZavZzsQbamvdR+szzMlMVoHECPLHRevZ5iaS5k1VtL5BEkWdj4u
tbTDYcadt0RPxyaKrgpqPA3Ku4fdP3wCfgLzBGEyaCAwgb1v4vw05udBJVQfGOs3YnM2L9aXIu4R
CBM9uOj2kalmjzZmyS6MxO4H3ctw3GY2P1uiGjSwHa62NCpeUidX5XAOwRbEMAT2GDSGmygNzogE
tRDE/s0su3EGPrr/Emxc+3Frt6/J4If/kDg1PTSm9+XfMsVhG7DTmanaVQk6Lt/KzAkW4515xy+N
HQg1NUup2MliACT1yw0Hf5xey2RZPWNBypEPnhq/i7dwOMi6eIf6ifXKTur8Sca+Ml0a7rMGPC4t
8Lfdl0OvxaSiPxUUVX5SmqzNowNQwWv+rNQT9IGelezZxUPsH4iOeUp4nQCZ7yzyYzvjLxNRk1Rz
KP92egggbIxBFYrM4jnhtxmH1RbNFnbG5GQWb1rOWx6xUxez0kWpNlgMOztu3ZexEh+Tna1mJYk1
3gc061yE39f9cOLzzdWtVakWhy33xFlEL87GxIuRh/BtCe5E5X8HkY2J6KRtORg3EcZiRFjiHXpQ
jE4/Op6mGeGY77vyIu/rT2pBkLChb3LwG/7wasKAKcRQnwZAZuIzEENM2YOH6ha8SJ983ELR6WTV
7RVyt7UgDWPnxb5t1PCwUXiXFk/NMpepsCpmY7sn6jgkNH+bSJSm+WEjeQYB818y0rj1pHNSs3ZL
C3o3vxIAPLlqr4fynx4lLi2nCH1JXlbYhLE40MUzQjjaN67rlPE8+EF0vxEKDzvXIQYdecKuLMkU
xoKFwKo3zZOs/y+WFppmsIUU3hCzhP6W9aEvjCTMs0xWkNGdunMiK6P2l/Yo9r1WsRdWxSwX5xVe
UmVrnZfZSPsnNzNMvtOLceuzl35bd7W4QrzexC0bidZ+fgBPDmCT4YRrpWBQvbVg7XXKXlhfZpbZ
IkipCtT6WacylOL6fsK1Aps0RBmehXMF5UTFi294M0N+ZqpRJfQWkwOWfsq42iYYIOUU3sxHt4+P
wDr7Drqj9Loc/Tel4gGWhr3x59Sp8DGKW7d9YH/hsWjkvh+bGO6Qd0BbZ46XjNNzln6Wh/y7b1Zt
3EeEksrXQFhSf0+yuC5yDohkcORbhqXRS4itHp54ggs9nSUJD/7BIr3fXGAgkcAq2Oe4kw1lUA4Y
aR/4fLXM6sBTT7oxAVDCehd7wYgh9GVHdQfjwyKW23b2etfnpnBqNAxl/PlnJd6hHt3YwZ3/yl2f
AQwEcouuvSVcOToV5JrmDTJTRfYzYQ6MtyAUFlxNGD0QWDH2jNbHRH3kD7tdeQJUTaMHD7Dc2M+W
6H9/2+N290l6+FZEcfG2xaulGDvIyM/NDMZN5hl3NVBK2ELihgRRCm+akADQlCZ7qJcXiL0+LpcN
EiUztLk18Al9Kgcj5AH+VfVGMvHqlNyvTF+gmDIlKreW+8mAkEQP5H/pzPXDLqQAtZ/zNbhP1sck
7pDoFMRahQ669MUc05phabkIrDua7mMUg2Jw7xqbZYoV7up4B4OqlyPcEXCTiq/JRUcBlZ8wko3i
j9R/hxjA0W4qEfZx45xcWtYl+ILrOeo+SklgOM6AkZbWEX4zRBHVFWqtsRkVT+iPDjKXbL1L+AKW
J8mVSibhifsqJyBICQBoCLq1i8shyuYVPGqKbeUZk5WqsBlSFqq1MnZN+ChhxR1gIz8DhyrU02/a
ZpeA8Dxr3UqUOQM5OmrQNBtQ5H+lP2trwx0dQLSMz3QfzDOl5fdSom+glLXE4WcygYeHfXZHeAnC
GQvSklV0i3y+2kWR4vO4nRegJ5vZascrXa2BX2/T0EgU+AN1JrNDuEvtpSgx8v/c6sOdpbswZqXp
m02Mbo7YC1w3GYn8oMcNXoxjjrknII2yhaxcWv2MMm8nPEUR23rMjPpeZnwM704nQ7+5/GGGokf3
uXY6x9bWIkY/VIS9xCXAG/HY7vha3ErnjW1D6G5yEAM+BUjuAZZSJrIrFbGjStG8YEf0WpYTWX11
v/Htz0dIBqe4ZbSHySIzW6zBsG1jxo/gRLk/wqFXP9MnYAvPQheWECfbErK73miSpfg/+SNqt63N
Ff9rrjua0HsNfGW+UkHmMEr2Zv19ilJOULHsesPLxPBpugrnyK+R0lsZKIeu2sEuDJ3F4x466+/C
k8u/7D9VSsczC2KCItc/XcqxQF5qch1kU99H/UuNMhhTN3ZXH+9GaAEZB8FZ3JHrSkluDwbcyinL
RigAP2F1bvQHJvIV/uSkGyqukctOWRqNPWn5LvJ4l48OmriY+0AaNMaLtqV5zaVo1tJ/rS+ApH2x
Zw5/udK2BoKteTQbjHpTl5V9l84EUl1mqRj20AcurrUoqFELV5W4rZ/24tTF3DgHQjyQhc3G/7ej
k+m9f+PNJtsWaRPeOsbBLdeVyW1ZKReYfW58K0+pXTfLR68gMF05+BR67evhU+hnBS3ElADRkqiQ
AVaPUIihDNXkzh2slO7LZktHaOX4gVDEr2JQM3eK+l9dUtNfpDdSG9rvLppMi4won2zeBVUZE01q
CP7KMe0f3CmDyaJX/Fh6E29FF8JJGARXUNqVHDoPTJWdI6XZomiWcKQPftwzSvLMfTs6jX3cxYkP
GxFD400EmAYOz9BDjqFr9E+hExmI31Myprc8OsCVroVYY8DXA0XecC+QUDsTtzHJW59aAYTwJ+VQ
5F/8W0OEqwj3lOYW7aMzchlHEzK+hu1kJvXIbYybAnwnTKlFHc1ogxrUs1lzo1m5+pqgKFaWFB5x
+Iv6TWO+ZtrWhtqT4tLyOy4B4CjVrOtakzh7pGkXhx2sYXciasmdqK8BR+zRBqq86WddEAxQJ4/v
homP+vFpvvmFiBAQ/JWLBj9OHYpbR75Oc9BxhjV/LK3nt6Xd+Iwm+VyR//BJRpxozRzLVkk8ptHB
Wo4O9wgSuSG/OHXufu/9rFaXW9wOPV0pFBJDMXF+MY+7JxQWGQ5Feb42G8GpR9dWOF+4FpBOJE5M
rtmHb6xkzzwDOyrs6goWE2KKobCcqEAAY+WgA01/fUYRnNVu/Nc+kzUs39+880ZvCPjUoJh6yDA0
HMGrDTpH4NOUJR8SqwnKU7KtVaFP3vGZfZhZ3rnXqYNed7rWnBZUPmLxgdVLN+b/T07nWe62IYWN
wgo3Sjg1ZVJQmPsf8BXRARpbaNs/69E/e/TgXWxffsd5GsFNv4DlSsMhh+lnW76L82DtPyIbptVJ
xlJvLgVHOCVzZ/zH2dyS0Fg5hYEHzdKn5//ERD4gPta/uM1TyBJEhMb6YDJMZLXEHOju2u7CskTB
I/tNIk08qT1Uv+tHqS4JhjUKHrJAEwqClwIaVkTBYXyRAkPfPq18pDC1wmGdV43Y4FVvIt/mBhWZ
Y0jRtF0DSDW4purUIL/hQZmFFWs3pTT9vKKkc+8rOCrxADpqpsTh/xR3DuRnWQFWE3A94GG6FKJL
1yIIf/VaFxFoDI02xDZYx7g7DsQkVLMv86oTMQrM3VBn89h0WVs8T0NPla1KKJaDC9MW8rffA/Fd
fJ7NY993dmygth0KMwNRtq6pmEHZUh23l2SxOVdFPFl8YmXEVxg9bfxfKRZE8b9/dx/eKT8PZd/S
7SHpKMvHQ/MRtZlhA3vVwSDYVpwdHaCTfzuBJLn2MMVISwBQK1E3q259DTeQIEpPxF59ZOAelht9
cUtCi5qcMlruFSjsWNCWDu1hk/L6mRj5VXLheuU/oKkfynrbOFNM/HKPaV3CkFVzecyn+wLGH6FB
fY6QIyxue9hDCbqMI+5+O2ZZcVt4NbXekgCFLhCN3gmeSO8Tokr8Y+p6lb6es3x77Et9lS1Nmv2i
q89o0TPNZslYdxjaURz8d1EGEVj1R1bd+6v7LNCIrSUUTvUoxuZwksz+lCTKM6n07bTvcx/jTDAB
Ll6iph5vruecbrVXVqiGXRZMtk+EuV4YNUpa5i9GLd762ZKXWIQ4iOsFhz3zJ6JkX89v0o775ybH
Z2jpR7EODCzXEqLwf7+XKKUdBnjwmyfOZ/f0eEN3YMLdYEmzW6NjNRn4jYpj4L+6IGGXci/55vj6
w4qm+ZaiLqR37MMxCJDftkDhN9i9vrnohGfiMT5/okSeTbWRNoxF0U6UJ02z9rfO3ErDkYDEGw7s
XSpuSb7Mdgcsh9XQ0oB2waxC6A6MrNLqRHYGl7D87lTes9/NKg/JbrJkTO2zkp2Lv8fhDbxHnEdd
VP3pz9+2LHk9xi4S5+/hf/1u9lh8IKa0WJZZYM7f+NIy3dEeQA3WMwjaHF66v25/TTs5Y7euHqRP
/Msyy37iy/vMcoKo/yxfrq8ka5ToWIHuKvrtGevDLzKOdRDbg8APm89TSkgsidBsMPWQGYgREz97
Nn5KGzh1sv7Sj+5+p92CEay54htUHj74StRUtDu86VSTHYpGVx61OXJQr8BHsUXVSorr07KgonR9
y+jLuvkzeWg0bOlGCe93/dn0/SlZLujMmfHZ6ArcPrEGs0+KopsHbZxiaZTYt1OWukCo0cbupZdo
0KgsDqoIUgPXF1hFKdda2M6rQRQJD23rCkafhmfHny+/VlsCpLJL7yUzEaMzgVkfFCvbizalDD62
+IeSdPcdrsa/8FGya4EcBqOjl5wTxMlMvWiIYNLkRHPm+0RayTDID9tMw3bpQoFE0yjUGcexEOr5
LCbMRF6/6KTDrlCKPp9f4LZciLZZDjhbRPFBXzDlGgrnsHt9aKLLFozzQlwoLTvVUgJcfXwNS02R
njqWjHPp2QwrcbCtcQ/8MGHvnIo6iMN7/VqTnPCo6aLLNeTFVsCYxIr7IVT6X/wx+jljzFykgyB5
/1+eJYdzjGs1ms0VCw2J5kfmMFfGkF0IeD2x86PrBYvZwmLYn2jXqHYvDCTqIkWwrPWLQj5HpsCh
TJEC794t/cBqTI9g9VTtxIJrBl4owYywEzK9c1jYDnewMRQDnfg5LK7cAxH0UJUUGEoZgDh7lVK1
BdX1BUM4+TQJIKrZa0b7SKOaNt/3OB/KFL4feTxtmiAgXcxNzie+L5CLyqGHKsCYF7kq0Td0Ewzw
5ecQktWTdKv6M2KuMP8qcviUi7NxP+baHK09UNU8iQ5A3WVmg+Th+pZaUPSI3fZL/NrIduFPd/cC
x6X6+gDTulDzGuh9Sbhle/PlCqFQxTYzP4LwgLm5WxJPz7Wm/0uxGB3b/Z4oYhTdwcVsKHinh8yC
YXGJZ5EpHZXJpeB9axYkMQWC4yBFtCDcTFaJUuwFxjMhs18gNzaHnVzbGfhB2n8IAIH48oNM7QeX
WBcMVYnARERJvAx+P0lsjwUmcCmfevrllvsRK+SFv3pApAng/XJRMp2nF9tlKIYU83eXsf741Qjy
CFV90x33YosRnhikHRjmjAKwEJI0XmjIlP6gOSglp3psXb75A87M9YOGfSCoMr7aQjLbwXZrnc+5
q4qJSUrfZQ6+uwIni8LOhoIZhoLu7+eXEbyGTiZm6MI3YN935+5wvTeGZNhUnplWDC6nvSqtzXht
sXURHUkWAAbVqeir2vpeqXZ3V5Z+d0xJ1TC2OoS/M1wZef74Kgzww6Rg5a/KBue17UVO+4bDVnGL
K9R7pqI3W9k8ojJe4JNQ0dmm8zjlOUF6Wuc6g6OftkBcyFdjzKTnYcsCr6LiJNa0dF4NU1ss6hUM
edXeuVnMgXS+Jvcn6SaSanXkWaaUtYHPsqk0oMAccccGwhxTo3/jjrJRWb/LcbPTPIL+ztzrn2xQ
+93/9guTf3UJce7Br9GAf6FC8sgJr1zwBB/fHsGzXOzAm0OWknEcyZXDo8zrUqtJDHsvF+ky5Qk6
7Z7KbCrH5sIgmjcgu7A5vGFUD6rFuKtRvwyDMhqNMPMfhvmIFUsi6GheVgbWup20oOkhLMG2bPY1
TawfdZaQRKyUT2/j/pO2U+HoTidn8N2yuRiqh4w8uD/Ho1S+UcbUZ1sO/s7QeiAy+TD5y3TKFrpL
bGAx4qc3t6bcwnf7irTtfj4m+8yah0eKi2E6iwgAEoShTqj2xSJSNnrYQDvlrE4wMs2Bp+geYhSF
sHfB5egewXHPemueJsY/lix0XkoMO0uF/ozHN4Gj+a4dul+7gWsKzEjoPDHXdE9hDThOZn0d/TDL
lugrv3EJWZkr27HPN8NfKh5ViOgizRdgSiOZa7O8WHvHO5B8t+AQ6wicoLLr/ZpXbXZL8LJ3IZ1X
qg4mbm/7yNsU7fp0Y5517nvCmGdCyrN/DJLFzwxOtdV0cciAtUL2UzXL1WH21Yqly8ZyFAme2IKL
yJ+LfzrGvpdFsrKVV6qLb+r4tPpsd7jUxE3JjdVo23ljymB/XgND5vHSs3xKRjzJHXWAyOjgtM0g
NRj5YhMnlgUGexCFsDU7SDet/7QWb7LkeBjsDZ+LKCphebainfV906AqRx8nPAaBJpVkhdLlU629
oiLdkZA2PyPSRDMgM6dBNzwC6dXKOFnLjBJKhVnq+zCFxGThNyBEgbfQzwrq7DOUOPPAA52T4Mws
JzOBvWLvIiqHIOCqABEY7QiTB4+X71x/8agZWVc9vZIVUz7DMwm6A++K2C3caqBUhpfQMzfuHOIi
UEaLXeihrH8VNo0vnQPozTnk8UTYm3REQrMAw3GRNk4qvDq3sqXiyB5n6Hgj3VzTH3C/9T3AhUr6
mgvDvVs6gLnGMdqa8JKWP4yB66wuJL7NlKPWfvz5K9KxtjLJhaHzZljS23nGOL+xGEsTlBphTUld
yXKZmL9AdTwGmVV5amsNvVccrL92CipxswJcNwL6hDiqgRwTdF3cOEgGDyXcHpnbxtVv3vyQ3+TD
NDD0EBFlKsJa0XmMpAHyRflBnuJetYd1nE6hCHrapxANqV7z1etrwel9eqTXpo2C9JdbrCRinsDG
W48EaO/1UQ9PNDI83DorBIXp+Qiyq/kg7I4UbggfCqeQidDFvwLZ0mC2rVq7tgMU7mCCghkBtYc4
IfJb/3z8asRTZusHONoUjWVlIQO8DOesbsdG4M88nCBDUrPEvoqtLTMi9RipuCdJnqefUkNvzZbU
nmfFB93fwbF24fiFMFRGj/PWAjrmq7yiU7dxHBEa5fPgQgUgEv6rJ3WfTJDf1ApUMuDkSLLPsfAF
KFBnQTzzsjOminkpcvJcQxw2pHxGOaNqARCr226IvOsU15v0pE8Kzq9ApKK1TfcXNGLNYPMU5o0v
vKSttmHPBSBPl7biMpmODwXCDJqNy1KhmmBI3qsW0wT3qiZQ8Zib4+hb1QO5szIgsxa/iGjfY9iL
Lb42OC2KcwS86Ya9DCmSRtZJgZXqD+s5VIoE6mZp6Iu/8jgaJlhaor6/8nVdr7x8nNnmBqPpAEYD
SFaBhZhTX3QOAcqFRLylin+myoqRMjna1cdaoG23LYLi8nRP8bmIJM/bjegdOB3dDRd3xDA4GTRl
degA+C3miQy9yIxUCLfZhIoymXQSy4SUkI8oRqPrHcC8qrHG0DeyWS56mnKZ8LjeJHlx4lWZPOvt
V8+FiSUTbVYy1gK6hwK4Ys5GB6nLAtqQjnBt8v7+7fUTJPRhb0sWHIa23sUEcbv6Ff+tXI5BpavO
0kgR5MDkmj5ri+AMRbJgKOtjEUioqk4LdcRMaTvFxJ3tG1wzg5Y9Q1cp6llSC3FJSRE3k2AmuOCG
NRdgv9FbbNC4lvDELU1+mwwBC/VLT0DfhsrHOuD+Sl8qc6FkozZOBQv5kVCJ7o0URjVNYdU9GB8X
aLLMOt9QR+H77N5Mi81G8/kKC2oTy5717l4fsEFVBDz8QfUyvYlF1PugNL9L7nK6TJr3KRNMz85C
6nhqFzTIvFvXQqz97xmsMEdhu0nnE1Qd5vX707eDWDbP40LNpwTFpiNPjGYGXP6mUnpyVI+Dx08U
v9yF7VwlWJzQcrUJqVqDdK/qCJUJqnTxIL4yPD4zm+0TWJUE7rd6oQnWxz9Y3oHXqzYGVafVo6+k
393vR0BIorwJxE+PU/SFW5/2kvLWT7bxooD9IYFCy8T9YQKCTtJY/KUkjL30I82K4BFGjw+XIZC6
/mCQPb3eLLCvzeIEwVD+nUkgaGVaqPJo/VxKICQdx/QHhhaHb0z0dvJAVhvqMRfbOeP7HXU3+ocg
7IOT+CGqctDDv+Qml8s7O6k0Q55HqkX8yfbYdkG7pmtruJ7Ab0LCv290jVUqCmhB++PPxFmVmD5A
e0TYRtzurs7EEM770e+okhDlbRRGyn/YEsegMCDWJ3DTXgjv8G4JVMAzVfIDnbYZ8mPsP0BKYcx1
cjKSzpdRNy5HtstMclsphLrNfJNFfT0nWxRtjLOyphSf7+L1jTCVMlAQocHp4tR6s5GZpvIIJPHG
4pFjYhdHW7S9t8bZa/7uiMWMHPN6U0ZAbMvBNRHzdsZnSgeHrmwm8NYt2DYXSEY4Wf9TF2aq1Yo0
hADpY4x28HMYsDzBcrQONMiuF1oLBbv9BsUESLCqdXFLmZmLJ9pOtSThbu9PLFRQVNkY1uqKFQeO
4Gj7ddVH2t4SVylh3t5zu56mMLoWD1CEqC3cBZfEIePM9ExVfkp8pnHMHDSGM+Ezy/XUUUQHCJMI
vm5yYRDijdk03vr7/mqvBnG17NaoMEf3McGb+r4KdUbR6rLSiD/O/6hNh35g4JqSrtfEpYudkqQB
+Zpt4nSCaC6Tek/+IBtv+yDIBiAMtm92EMGEskhgvgUCzJZH/t7X+HHn3sAfS4d6r+U0nskT/uk8
ucsToIbCBzV5t1YoVq8G4189APy5nukBxE6CZvfVks3G5jLNuHgujfwx7rLEykYlRmE4zjKBr2NI
8EiDW6nR+Soy1J7Nd95QfmktIKixKaZGY6bNOy+iGv4PGOwgXYFALBDiVfxs0+NEJpLXutq6Gn0k
6SouO/HnYuShBADxWvotUSX5klioy7mvaMsEsoi+gdcEqSTh/2JhRxfe9vgTdRP3hNB7Qdu9CZJi
dM8zTnIXzdKBrknRb0NBK5kLHuIi4dHAh2on36QiMWe4sbektYuqKhqlNOZyQrkyWzOiGSDsgKzc
gWdsVUxAUCXwYmy44kQ1P3qSuOcOc/ZD2IXRXQRMb3EHZEK8VFPKbSLZi5GlEnoqg0NXkyhPmSqB
4XukoU6T5p462fMZKZ15gL4ch0IVjPY0byN2iIemwnj9i40Oz0ECRTLYAFjMAWdH3gBeVA0TABKL
kcYTD9UmaW6euPNdW+l2zc6IPBhNW1jVPesTyoYOG8qDOi55RrLhR31fb5Qofy3FStI9jaAN07hd
nN7f95deomSnpXmKUvemOi2mdGuLjcii8ba2b3XdB4a0SrwT5PaAET3K8+kBP7H1BIjJwQjMAsED
eihfoLOcs8F56wTTQyFRyMEUgmstY9+WSpy0n8xAdOke1bMhbbs/UiS9yjo2GJH4O33fNH/jiIcJ
nHsWrArlZLVZOu8fc/BT2T0/2gyGprylt07C6nVXuqOwgTPKYFM+vRSI6WgyD6Aa11ADpu00yNb+
+No29/Nlm59NGQMJURkXcMZm7Ipsb8a4EiwP7XgE97hBRwWDJuXgNzyUSas+iDVs21NWlW09F/TJ
7YYSPQ5wLpa5yoNJeLsE0eSCT+zk0uT/Sr/M7xFwux2riiOmCNefJKTJeYE+IY2kmTg/4w4BoRkM
4o7ePkmrJ/oRbsyKjGhwDcFkqskoarJBrOA/MdyIxsv07wc7cxhS58lO0wFSppHCoh1cUmtTC7K/
o8YWqDnsfBUShOyXtVRQKqGdWbTILe2aretBYaGAM01cnRX2huZ4Pi7C67uFteMUzSVeObJP3Mdz
GRmnC1rXhRyqT/uXNIGkPOHYx76N1z1LkzcQtVMsCLJr6gaGLfTUG6wr/FyIfQmdVGVFln0R3Krw
SOvFMmvcEvbssiUS69mMDwnJy5YhLc+DlYtX3gkoFnQ9xeqHRGg9EZS+rK1YaDplSm+nBXh4Yrsr
k0si5mtdgK+VTTog0SbDbre6b3DhdAiG6HyNp6vDqY9xGmtu+sHy0cDZ7m2+kVUwZ3KGVNqyrlKk
5q0ZCJeYO1A7a2qcXfz+FL3C5sucLfoyQ4X1XyGnAfIlPegdysGRROZL6L2W3Sbbt4pudQNNtn87
qB7MyZ6o0uVBcSOLViBp/ebItEC0g4NdTlTq3WyFe5Lmt3qJrkg5EeR8T6+knP/LHiaZEB3v9F3E
VUZ9uOupCr0a41KsYXFrn0konZ1cLvPvw61xT0dYeX0MAwQjDeOxPU2itnzZYR5Hw9Vthc+RkrJO
wBRZmM6/dzBLyIwRdyMnh8lf2gZxJ7+LXB2bLmQ7c1fmHN4if7ULSDLOAT6GOzR+PzoVIP86veji
1lw+TOC95Y4qU7X+yOlMUq/w7yyuQ6bF9ikBRCq09X4Tehw3HDNDPy98OGowgGnKke44o07JYtri
tc/TLkPaniqgS7iR9k4QvZxdbRDR4/Y/HIK5+G5KjIM2eDCVBufd5eGyWnWCHYVk2kly//0p6w4z
2BO3E7Yecy840z+UsGYeDch30MGXUTDOtSfRBgE4BsOOCuqH8GDOaZZWqCM+jygHucgRLIl07oGM
1swPlWtmBhiie9i6CfScCEJDr88ZTsViDnnkcRTeRR2uIcanrPou5CN5yStZ4GAAhaYqXu/A25aT
e1GlW5aIj7F0VvvPYZto/4IUpntkEfrcHjbwFbULG0fnmQFVAqCba1dD0ifPKMdECk8IQjSKl6yq
B2y9O3t16aMriCfmAN5Ctas8Z6pieUGoKXJ+qI1s1RDynD6CQD3XnmQOwsDueQu8Lhxtaa1dKTbv
8ERDVHWXPfcns7b6zZJiQrs2zsPoTUT2z2L8wxSqLg4J/7o+Z5JoYRXfAZ+Hz132R1z065LlJOST
Y2BaVfHIGDv+fWi/YUsxPn1e8ABYq2Fse6AWzBK2Bc3seseLUlgiAPwMU3ZAcv7fiEiK44yCcPt9
/ZpLmER4AMVdP9h9UaXVql6WN25ObgAvmFP4pEYqLFxm7Vez+YZ91r1o6WRGF5pzr3kFHvKxBjWt
0cpUelF9eWZNwbqPxrgddRH8uHu4m1Oz8Bz99pPGbyLFcZObneo10Ig4HlcA+M9QxzIgzgYmDU4l
Ydfbv1Lfgx3C3yHZWdKqMI8RGi72It3P4eP3VkvtUAUEKH9Y4YUhVmR3KwN0eSiN+0/h5B8BPaCR
S9NoRfOINrlOyNriVImZ5Ot0nyz6PDi1gRAtCErya0FnoQeKj9NsKKOh0IeOwdFX/9SlVZjEnYNP
KLP2l/V4a/gV9fdbo5OQjydEaXCUjEz0DfHYn3wzaWDEH+my0gkWESvKt7HYAD4hw093kb8nygwE
3IDYuIu6bwHn2nXgYYXEZdBHpDTA9rvrIzixZoewmL+opbmJCSjulgwZnRtezwjjtYJDmNmHO4iK
YvqJH9t5v21XedgCqlEzQdzVZ/iLO6KKu2PY4GN8tRlkKDZkiTlsvOg4Q5mrKH7ZAtRL73RVfVO9
f40qYYRUt4g3bv0o4960QOvsaPlC+wXsKgbSlkCu2SBIlQZ4kBlNQJvNETGYyuQGhbtYikQGnIVU
uXL0eSr840M+GKOENpp9dpj42NVWf5bruXYuThbto89crFeK1/UVjeM7De9L/073k5e/MDPEnvzI
2cgJcFAhVUVmfMC8Geal5abKrKnbitIjm2XPOEI0zu391n0caKmka2ekQxemJTAwQ0pWF37K1e+o
cHXAMBHfE9omTB3GTFO4TUFKGhOAex4xXN8UvQgTPKz0Zd5fVczoXiR4fjpeUKN/yT96M7WPGoGJ
/QgjychhlRXZkLy90peQT5FbMioHVzxSykYVOw9J2Jv3QXgU1XL7pfckNAvVtqK37149KbXjzjjW
LNRih/Q37sJ3v9HvUCXC79gPkRw3MaVoPc5OEJH1IpD9584gOdhUcPlqbx7JECmbCwZICJiQf+fo
Q/F0lI1BNawErEo5/28UMu4v/h9Tt1HkAmI4DFy/SLmzuq30WgqMiUpUG6Qt/up3Dczngz9mXWZU
Fw9OLMB6+mj8bnchWa3DjJaQGD77TbLsos1KGINV47ZMWK6rsC3dFJYynrgYrLRhtGXzXntedNfa
FyXu0AIT3Tz1/9uPYxykNDszg1nKjAk7FrHTS1lKBmG5iYzbHchssyRhUz+YWY/3q7HGHskLzICC
1b9sQHRQROOGFWaHCQNHkthAXIfxfXJ2JHFitPAmQqHWhAhZp3hMnw1K5v7+wHE7OAUHGb+PyNLk
rZ+JGcFGBdR1+CE6zf+aRhAN0Gpgkqfa7AhNyBG/oVnUJ9SVU0uk0aRtzPMZF925YX+gZDKsXVhu
KplSIb23C01+ueSkgYMuhl76Ur736n9sNEqraeABq6azrtsJfOV2TJ/DbMOxQy89Ptg9M/H8Rwqy
nSrcsPx6KAido1dQfdVstEOe3UMdZaj2bDzWZyPpkym8mPeUJutvcVCUFRsPZ4euubOAgIcBkTuz
idWeLAeo3wfrc+d89QiOfXiOBXwtgrSSwgSMnvdNQXFnTFuNpbUFePj5b6Q9OeeUt1Oh5oOh8xDE
I3IYabQ4IVIZy1+dKTlwvpJ4gmlo0WJqgXLYlbmlhpt6QxN2zRAxuJGSqLmu0FSKg8jfZK8gm5n3
qRpiPBpFMGNeAC0jm2vUthcRIBz65YtV+U+fbbb/3FYVp2nAxWrZBbxuGzR8MwFPjhhiTbcAwcDR
vVzIa8MOLrvF8mQbbl+921zz2hITKrG1jOMOLFLHXHNu1E8cH5xi6PeJK4yUDIMrT2zW9aX3U3QS
M/dp+SqlQuS0o2gFJ2l1yGj2FP83j0J8tYq/piUjUqay5HGvJGEgGKFMpcYUkrqjHpkgU6u2iVnh
qoa8QgzbyAYtLk0Zrcw4KiXHTtdu8ZYwoPUS/oGTZRp7BiG3yTdbyk5wVqtjaEaza93z1AEPsZoc
PNmIV3N6tgIhBm5qDakeDW/Dj0c666AcpR4JpnmuXRaYj5hfWjvAG+Twci6n74RVkW20YSkx85As
wCfXxmi7w/xhautSD9QR/bAtFNEg5GLvW58gUtx2spHzhlRJ/5Y3xAPVxftD7OA+BWm/O+ueWP6W
aNp4CdQdh2HPqkRCodAQqCUORcWWhebnyrulNuAGvm80yvhyMXghUy60xKsscu7/dIro2I3Ds5Me
esct7KyKBpyoOsugFqBMFd3DBfvIJEPIsG//FyI22omKPotUhP3JOEDrbQs0wBaW09Yivm5tWv0c
aQPAoOwYGig2jev2prVzuwxAP+X12qV44jpKpbZsBvW16ynqlZlYm+rEgqZyn0LHwsXzTUXVKRsC
GvZKAjXgAM8NgidkrAxVkgBtRBhvQ1NMCxQVU7s8+QKitmSpnehTOAM8lDdq1VSrlqgfU+GAwzoH
45lLNWhCgrSNTUcXTGU6rYvQq5yjYrFofa4H4dzXypujOylWtt6Vy1x8A5iikvx0yNVfwC3B+FQe
aFMQRSL8zw2p6pJkJYQc2cKoERfyMwhC0+D777P/+qlH+mhzENfdeLcbnjH7rPZKk+cWH/c5cp1c
oiVelZnNbk7NbxeUB6rC8acs5AfbhFfS+CiNnrqXaMUjVL91tGhRVdAYDV6kPJfekvbxZlTOUPqG
7sdu7XaQk3DnHUjX1YkP1KRvPGO8dGizgdSbo1ak5Pw5t+V0mtTGe+g0apwGfeKgzbsHaHjV6qLB
6gY6bQEO78jqD4vg3GGlRpQKKKP2mGGx72I2OT1ceAHu4A3hN0TDyPRwseAu+7PikmFfn25BHKeo
xlDrPcAlJXBHlhHmuH2bA9FurVdHkBIzLJGsJC3kCiASRvSQWl28kBFBkWiRb7tt4r0IdFhTnyz7
TgOegbdZgDhWLthIOWjTx6kZo2p27keGbIUXIOwLoda5V4e4tu70h2clM59foD2isHbnDcl3JF2X
a67Nhb69xBmAfr0/99FIko8hRikYg+K1I/G9HmnU06ER6knP8Mo1CPvgfTzM1Gg1gdxM04qn655s
auvbo04iKzD2PYv2cvwYmz33vWAFku/8o7wg4lzfe5/Vbht4gl3QpTfVMq5aVntUO6UhJFaSMp22
OBhCHLWUUbgQWxYTkA8S/tWeqTuB8ND+j5S7u136gxLYtXegNLsAkoTVQRaxAVrA+bHNmAnjAo/b
POOGHWrj2iCtQVsiWL0uhiNE26SuUwcQ+KxqPCBRjWW1dYCKhSAmUDbN/pDKnK9nPNbkl4ycAK+B
7W/RgNS7qin5KL8k89b3I79FUud9/Fa4RmsC7RJIHFZhNARYPnw58R4kL8CmQlV93TJBUN3fy82f
//33DB2KCPb5/eGhFueY8eszHFtdUZEsb5Ti+piV9mct4IbwpWajk9WwdE8quXA/4mKcaz4PZpYo
7gbw6oeVCR6jNfR125HKpizxn9MKRUb80Lavw2yoSPiPQL4g5bkd9OrqowvAmhvfTnb0T+PVk34E
bmmf//Nb7p+CCgG4fswRyPlEspBRPiBg90u4GvMFXt2cgpXSW0XKwzWEERbxCL8dL2VxqZjT8vnA
K65MbQXsBwjvWSCLJ5T5N+APcQi6y5EqORP+59BQsVNmS7+Sm7s2XOQ97AzUXVIq1I8y5ocAFALV
+AK8jZM/Ny5yw1Rop5QxCuIedgESKHsvr3hIG66hAV+9S+Bn20M5ceE9kMm2skU+4v/AaSaGwaUW
cG1SdJpbYM6UpLCbSBjfgo6BhyrG1mApeAxfhhSnd502i6pSw5qzp+5lvVK6xXPJG6wuBumr8inE
l9lNjt64Ic5ZQ7NigU23TLS6XYppUemXazqM0AaL4w2BIRBFq/x5qo3zFcAGBMzLoab5vea/E0Fs
axGsGb1oauCYOlQeZ8OUdhQ2qLKaHHzWJKYhx7+ugh1Tg59VqBcJYgBpiuN/LdqndfVZPLRSztTp
i6ZwsMUAjgVQiKmp7XBirkvUYt1gAvjg80Abb+b/+dgE+UWFgDB1h4a/WVYdd0sVV0WsHyHgAla2
my99mss/b9mf9zM/hyWwUUTVvqeTWbHqxhye9URsAkQjBJKVV8LR/n18eYoXQWrZhCrGhKHyxq8O
e5cNRjCPCwf7i8YwViohkKqdVJcvjEsLNs5nny5F38A4TjMjTAI5Gyul2g0kJ4DzFtgEksrR0ko8
WWfknPVxJavZpiwhxNFza1vFo7MuaZ189cY9TC1AriYwNtn0bIbsPs8LRVagSjSePkkfIuuSXUEj
qoZt1h+O4YBjHRgLNJFfbcIomWXSOMnVobs5oX7iufQeVimo+KMoiSwPHi9klzQKBmcWt4mdkSmp
3lsUCaEz144XiEMLNiuD1OcSk3TlD81Pq7rN9683x5eTC91Bn7DvQ0m4XkTKJMzksxdzkS1joWDI
OtMoz7AkEWhw+lcysO7ye/71s5blmNlYnBBno5fClNU6JkN1bZvJ0WCB6TFujO4OOiO+tE7SPR5o
njGcgZASc+ZzOJZQfm+ckAUyazvyuStPcPJoDDkDC4FXdxgZ+4qiIcguFaPj0KfXPH9evCG2xDsW
lLMGfn/n7M1W6GYwI/PT4KVraz/KfLcWjk/04gs1f4eEGKQCbQXzLuxz3kmb8tZMOM1M8lOWaeca
DTb1K+C4OAtuYjOrYe/P8YzyW8dDtyi+QVklW6xkS3l0C1KV49qm5q0phmrRyyAztd0N6iYfnWyo
SsdlDY4dHOzivSTrE0aq2KrKHFbKH7jSsviFqSOWXfDlLHwPOHTGMczSWgifh59KtuTcSUO3sWvR
SAGVeXyz56z3/q5pxX0ZsJa65/7AYdLHeWpVtcMmAXB3El8JpijSlUGfhKe05cnDiDwzuMrLjARy
CLkSqT3RGMZKdmxbdi61l5lnUEPI1Dq6zS2JFQ/++kO6MtTmWv1+O5lETL/QgnYerxcx8+2KDno1
jF1Lx40vz8h7VJbN7fL/3M0IWl24onUxFS0hvVtLhU/J+wj2YI8c8Ba8Ib1OVno8nAamqz1Zg20A
ym8wk362ynOSfowcBIOji8TxNfUZp4TZsYy2N3t1oWUbM3oZYEvc0pTL+HwXkBkyPWPquip5R75j
QU4Tr2/I7MZqeGpt2b2dxNChNigkDE/Yb8zfSRLpYvP7TW6xMEgnF2ZDfbx5hW/eokkaegOV+AtH
dg4EajQ5Yx5loVFLG7I67Drwsu+YC9B+5Ndxa5V6vvV8GX4h5TFWDjPfAhmoY/MtXnqQGMOw4wwx
RW2ivU+so3nYKZ7YnWPEai+ow3CfD5HG8CH8RCQzxNfV7f/eukpvYIt7nSIOryytNM+doCYAufQQ
ud3f/GQtOqJnUZviPR/ZAYGTB6MEJFEKS47UdpJsvyvvXVKyGLJQXTWcc9QmsABX++T+4Myoayhm
loBqjHkYKWwYjxxkuFqwJVONAZsyz9eZUyuuCWp6steY0NkptSDVfD0mhDctb2IQ7blnAMyZznwD
crjjqvjuMVHL2xbV64sikzYUe4Kji3q4LtRS5TrmWkzc9eTwwFzdn5PSNdJYlkKPNn3/uF+ieDDF
KQMeJLsGzAieWL398AhUtSwA8Dc2NW1A1thqcfpQMeEd6nYyArLdE3D08ktMaRMB2joFNc19UcKo
amcwuOTOWK7sibLK8feRkPboOYoH92k9Ksu1UQujVEWq78/87Vhd9GT2AiJygmEM14CL/ImRAMJ0
r7VhzLkFGMwxpiwmBQcAHLGw0nts9CiX6wHIUBrCVwRPyBiBT0KDl/yi5Xs6su933Lc/vyBBYXin
v/QROxbUeUPCHaE25U3iHc1XqAG3T5aVGqDEDN7OBokMvqzCfrw+S96PJVlqeTDfGknMJxOdodFy
J8lzrP3rFriqylk0qDNDixF5LT3pYmca/ahbXMTmTvmD3V8t5hDY8tERYWnVR3sMglhotcdjOFNf
nVJYyQkWGJ/ahnMO2OSjAitkF1OBmpogsjB1Ed4EWxyLPZFACv7s8yPUmKrA/1Utzx73qD5JO5JQ
axD2IRzvBDg8tUOzK64ec//0A9V1TnULv3NOQF1g0oDdyiWHW2SlU1KuyKyU635gqBglk6YfsIgU
pv0sDchJhVT/kU3JZVruTZeW0vwALgyQQU7PdXFxKa+bhzOw/nX4YVsBwAJci3caMr4oBKxjCkHE
UKM1In6upALiZY8azdiRgEDTstYIC82j5sIQxxWkMiF0Ida2OBRlom7zJ7Rl9IMfgqMVQz9fNUpJ
GWyZZLPNiDZaGTTTBfYFh/nMu73v+5SXa31prenPLXbxDI7sPZxpZcKKrPLW3Dfz+qX9eV64kZq6
d9dxOhfXiKaHW9K4C6VQw1DzLN3rawpUHdN7PaYawakgtaLJldub7stEZ8E6SpkwR6aQeMjC3ilR
knaHjkhHVDDV/y7u/MDZ6T3S23bYTNfK1Dbcs+jlObZk+ALIMP13nwIm5dtqodoFY5dZTPWkxSTH
Z6mPxWL71I5aao21KXPuBiNT8xb+VQBusLrOMusRzOgbUI47flX1F/QrHuglJpwAEA886uyp4/0W
NxQ7N6JmbqEflBI5OYaQEa4z2FKh8YNbhS5MgaXD4M9VJno4cf0feZ9rQtRJBmFh0F6ByG3JBgCx
g9EtOyHNmnpZYVW1BRp2y4vogmiK3k3gWhIRkeqkkAea12aBtDBHoX2iQRnPZUjdvv5w8sldNRbr
+AYfbhyF9icXsLbumo+UIh/omLrxFIZPLHFim8udkAwph/BdmTYDJIHbdUwXkApf3VbDEVGYoABu
YU6GwsOfCQxAK791BTrU7ktOv+95hBGN4EAq++7o17j4wvWuD9aK7ooF8CFkrIP95fYNx0O609nw
HkhFgcNWjKNY+oEFjZEkbw+ugZ+X07R5pg3cZqCD8DDFRXmtwadE3UgM/LylRlsI4Xuir1Ad1qFv
inxJN8mSFHGpwUW8a4j66zwFuXtRrbiXE4JjGQF0h3ksu1+4th6XAv5SR99TzbHDuhbAtRJubPvc
iRzsu2V9Bmo93+GFn/MhPM2gDoS9BPZQwUTGypDam+Mtfu0S8mKdNUgEo/WPQ2zUDd20ZZh0gtoz
E4vnNveyliLrN5Tl4cLCPp+M+dEo8NOKR4iqR/SwcsiJMwU4WWZl8zaQkpq1N1/YNfcz3j5JEWq7
K5ct9ozuTPSRzHfEDVZmdx8G02Wp4llyMO9bXIlaOBQ3cViJHA2Eo5pUm8le5+ASHvyrfZJFj2kK
h6zDs/geQe+XLKdVxOI4v5FU8qOr/3CgnD/srm7LPgwziHNPoQKTcdJ1DZW0MfrEuXs8uw5i8p/W
rrUBhzj3o3Fb1BDY3oCVnrBskBWIDpcHqGih8wsTOK2PnKgGQ7KUpYdumLCq7Zc9ntDFAnLTgUwt
WDWSSLxscvETrg2CxlAUs1TA22KSNi9mr8K3Z4XYwlvtFt0TSEjqrJIHNvjOb3asTvPw/3y5w9Sf
XdAVwFbTf3NKHYTCg3h4XKcZAUIFIujvRSrZlAoOg3jzH7lbbZDa2r/iTV0aCJCtpjgMOTDBPsCp
P2qFMM8c0I833ogzBGU9+U/ZLPCa+UPqRdDwnYPdfKTyXHtTA/4fLvwjp3sms8oVc6DgtYl168KH
QcGVTqLK18AR2KpUwbMDVby53HYDu8jRmjqcUg+Aoq8MtEALIREKqWCp0hJ46Nt0vzUuIQGus/ut
xg0E5iRv0PGEsoJUV/w3tfRS5WBYpEZ6uruiDktiPYcb+kymTQNKLrQYJHcsqwKn9XstFtUGGS/U
RR9/3tPMnZZgNR4VUeVKwlerlzdkkS7O6Me4g1uCz9MGscGFRWE59zhQ0bedHSFdQnftw/Dbqer0
p5URllCsKuNh4/ae1lbtljYA4vj88Gy0SWcBVQx6N7q3OBACEK+kHc9TF1Ny7IZFj+4OxxpdKV1V
7tw3aUq67qyj2VrDmaZiWIo4d5OOIFR/a7+rbPnHJcARYpF5uw5UOt7VK0h/oPtvUastrikn8+vB
/NexigS1dQgmf+WS31wlnRzIQhrFeBji6eoocSTqcaByhOWe5JjfnrCPdQJD4iCedNW2Bsrh+PXQ
hGFDAZFIeWe2RfrgoDRkB2zl9nSP6+dqN2Sgf+lOtr0/Chd4iad272sU7fv+OBIC5D2DmE7/HEpM
i9aAqxxEiO97LPiIcvN7NXCGdNKTAYmcgWrRbaHo0LMvAMj8GYYTinupDwaQEquKTgUoF7zQuMJL
WkCqo2wPta97MTQQ5z4x9mzlD2Hp/83SuVa17Io8FtqJznZIhNaz6QsjGDaqQ866tmO4FvKFQGpr
4ykYaWDYQ6yZkbN8An6ZuSLRjh+7ctK1jenmT7koUHTFHwYgHnEPyUxUAe/3cya7ROkJMEQCcut4
S3KuAd6NXapU/RE6YPLpInMPjDXkf8tf3RVv9qUMVLMddQbEwvIUJZAvjA3V10Z5hE8jXV+IRTjF
Z5ufQSqHXDBM/qmG2E3FYa23NVTRA2a8whMi8LVVqk/85pPNbiB9uD8He9sHqyLBixqZmLHx6K/p
thCV0uSWuPAYAeK7TIZi68GjGWG2JCP2P+Xf/G3KeLhMH1q/BhZFB5J71iUItMRa5Z5MN+Is1b61
5Uvcb9ZWnewlJ7V/duAKlhzlxVhf1Eh3L0IKrR2UqIEnGEZt6sQNYfeDHQTuBi4CpHdxji6OrFsE
FrQlS77i0E5dPIskwXv1TQ0YudmMjuozeMR6DdyD9zXrmuOLIwuOfi7sJEmafT22gbp/rtCaetoM
2XUjvY3UB9FqYmOlfhrtYahf9yvJXG9Tkzqbq4LcmhlPODBELOFak7T1v3B2VvsQ5+e/5FblDcQh
okgX/yQPeGe5WiTZS9fI+gvI/OuWxq5TQOW7VEZargI2uJuVtpmBYdwbS9fo+ACnwpLSoEPt0BSz
shI3x2E7ulT6kcw+1756n8IOqKpvpFuTtU6Wcp+ByjDL9jqLJGNFvBWRBf1Znefo6B7gZBzN9uM2
m9iZA2nEgmMibJLMSSLU1H1VtdTZFTyKo4lyBPzbhWNQ1H/whz/K/OPub2r/FTVu+YDG5vCKxjKW
QUpCUhkC2dCM3Y0g3falnIcXgpKT8ERi8YStuwkybgGH5gT6oPzmwGSN75NeHzxq6C25crT7OPgo
3D/HczUlBlIpF086Hd/lxRHtNFX4X7sIPKivpdCQDCqQw/fXPK7j4bK99RKKl6dYCjkzuUNWu91q
k3m4orA0OmbkL0GrZrUaQP3xuOinrjCZ7ML/WGd0dq9Km5bRxfqx5o3whHovfakgaIBnLiqiSCKm
BC+4/uGWycjkKOpRRloirCrfut/ENfhb2QNohFi7sq8Vo0TLxpD9Y+dEP7MrJh7+i6nfphmAeW0U
EoPBnhyfb0d+luzwnKAZiMY92UtVE5lTPzcSZjUwxHAiEHKqnTXMCI2TN5MmtLlCYO7kW5dUY4/L
wrdD4z/thhhRotRrj8vUNC0d/DIyYjrt+lgMaeBFzaqWVSfM1DIS5G1PJ7UL3wpa6G6VKxkpVSXk
ZhIHNInGqIQL5BSVISWND7UNieG+Se3uPn7CSj1oRpwFmb5IzOGB29LI0UV9TvBZRGBxrLlh24ge
ATCbrAA67ZP/Qmb/tB1VqTtSoO41RK6AMCcryVWApSvGdEksUYR6isdbaaD1wYhNbtK1odRlcJnq
fB1v9hVd6lzkUgoHa8oJl86z+Jy06hqNsWvUQczW5aH+1lxnPWjDENzOfiauPC8+qPx4pCI2fW5N
WvXKWmLqeUHGBIon940g2T95CtYEFX+IpKE1UoEDE1+ZFQR3TCujiRb/Pd+3zOK7yLESDvN3oSWV
tDHbc1JtGdrranscspPkTPYQMEA3IkNAnziYPs3iij/+N2HXVEejkwVHNTXLbxzswn6niHyDkQUn
g2Lnvzq+wsw3wpJXuaHsTlA69xwm4AjLPdniEs1HZkG1lTIJaJlWl+csskuaL9CXpgSPedgDyahS
ClNHQTt5F0ugjzAM/R7G5h+3M0tw1E3up4SVYa55O8WJC/fRl+qbB0hHSJx58SvOUw/6lZzYLuIz
IPB+mjfbc3bOaXq3ujZVJYGiKMEyE/T58mcm8SdwNyJxfbUSLNGirANtPybe+JOq28LqmQ2sz9jJ
BaSj8b6dwMeHgYX9EgdBJio0mxieaBiRkwhwAl5mF88GW+Y1CdnAPhtBRowmxBaym8eotZuugncR
Fn1hKpG6IAYq9tJ6RfatsoD+QT1/rmd6YQkiKCVh93O5HsxaXNVKWMohRMN3GjW8zzmKPPxkmzLH
Dm/hgc18I7vBbIK4WbKljTJcYI+yC1T0oSzSM/9cZNVU5I/J7QC1Xe84M12QJI/kLo8fsvagu4C6
deFo0vO8NNHjHM3h+bAa+9k3Vhd0PsKui49oiKbtg9WL4HBpiD5zSbsNUAZZaEB053VsFNpz8qv8
HA2wxSanYMfzrPJyeNjuT+XelosK5PK0FYanWNiRzNdCfw23jd+CJfPBiBx0V4ABVjibt7xmoQHI
xAybJ4gZZ2nc0yMT00DjavQWnwyxKb5XOHYPufK7lBrWcR7xJLEO5mN2kUIGUoTSfUMcP2JGyDIy
9KoecFUlr1KAn4E7Pd5SYSWEC5kDP0LXxmpSeFqwObg7ZdKnfLMEw32SdUwjcUb9XWprW7TB+lOb
y9e1KIX/uZMXBXoHoHDTpHhWNEcjC6icgHv1yPcqI+NxK7kQINAdJ26z/vElxvoI63VYdUtQ4GN7
+m3sZNDvJi0hPJv5Q30HyIRMW33RT2f4kQLmmvyiTLt0SDdTuExGEfnaKhMof1YyBrrytLLNZzf9
NJ5QPcUlZrnKqywL9wMEKIZK/TcgXPKpi1uHTjsNbRHoqKHsX9P0Vlc+WciChNiAFKY97sAm4oFn
nD0BMy0TimSfkM5gPQXzMfNHY4HFFAYE1Z2RhgUvOb5CDgMuHIQfp4loumTl+08QhBSk7Hv+O5lG
r41XYs2PKakofImp5MtwpI0O7c42Baoa7+sUvBu9YCS+cuHEPUxDt+pIkKgMtv7BzC647pk8VVKS
dFIcbBrkv/56qpK0nkUMFwaX5IHM0BeajHy4wOna/Ns+SIKP7YhlY3jq3VZWzDNC1/7qt9SlUStQ
PGvts/JQDAdpVi1f8ZffC31tvwBJQlikQ1qiKl7Zq63si0T8h5f1KplanLriyx9tu+kKvJaPAiQd
lnuxB1ARsp+D/rTx5dIuJdZQJNqA/+Z9Dd5gtkzGeHGPJjcgo8i4xkuQ+VZ6yFJ4uoA7CmCXJMvV
RCNVs72WXHZKYb6wf8XvJksnZB4ijWTpt/EdXdyNwKQ3rhsX8NY6ivOyoChSEnuW5ftpVqC3luYJ
L8QvxJItU4XfP3eXKpb0h3eBLavwmNRytbF2FxnhVfwkCvP2Qadf6YQrxJiCWgP0XMa13sRaZLC8
Flu3O5RQLG8VO6VidNTvFXlXARC0KbEOHRKAT3qRv8PRJVRMttlPBtFAtfQzcNuzTXPVzBa3c4w2
VyvmICFcyQ8cxHqDvIcpfmLPHvC/wwjVEWSuj2fkMbU3TdKh8B+AVJOY3R/azQ8Fd0f3hqpxWM2V
YEUVOnC/ge47Kuleu29Ot21nkyfBViny3z505JVoznvCdR1tYlJNxgIq2+nyb/oSSGZwQyn209q0
QKaS/2a2h6nCDeI+E4uINjbP3SWOW3kI1qhz1bK55vajHwCuyQe2UYpn1zdYWFiF6Kgd6datpjyx
sJvs5DRKpmJr71w9T9Qyce2+3cpJxwehIhHmk8Id0WIpnmuMqMEDXkr9jdWEp4aCm4INSzsjJxwU
luB+ak7ccxvbtol/b1GIOcftUDzXwRWU8WAcbkqoo7LBHbddZeKTHV4Ne9Tlgs/gQLqGbSiP/seG
v1B67FAP2zS2InyIiWOtVJ/M1eH7u7qzWofAIaKRFaOqPNUT0XMeVLvK/RKiOwDDrgbi3Gq27DCC
WVuQDJp/2ra1KeCssAvQar9SLgFvLO4oV4j7Fuxlb7TaHPXwx0U8kAblrcXaU4Dua6XtZiqaS96M
fRTUT7BcDLbzpy1YvQQQDzULO/XzgXLMbrTJIy0h2Z17dNXcXYaC8l6QN8gLrBhJT8GipV+bUpY9
rqhTD8MliifStn0yYPtUTUAL4IsZ2lSWOMnhLJL5cLvNJp/nMwkjSkLgil8gBV4x6/BX5mZJv/Tp
OfE2eB6D9c8uhAk9a1vJG6n/fz5kBT6u9XuM6VCDn2kZZYboBliuCgt0ETgsfFlPG7T7jpNyI+V9
79NEylkSy+p5tKB7NiB71kZYYCkq/y8VD2kvPcA8glprHusUzks71GxIIGcPAXI2Agabuju6A6jv
Svi6O+UmBUDst4ucPJFvGistySIYLZuvqh7zLrE98k5t1ZojAmxkjbh9r+cWdJHLsRclqgAxw/iJ
Piv9F1Ct6PSG6mHfRIS5+SHbU+a1i7nAJ/MREHgWkpM0Tiqp0k2Mea/++fATHeLMe893y36zq076
Bu8Ousoo9h9Aze9uNiwDvfXGLDiai2fxU2V6+ZXa0DZQe7s9ywjmf1ygsZfXUACACmj9Tcctfes4
tY8MGy/aMkvGVC5EJdFXtcJs1klybwl7HzIXijoIGMkWJAhHBjMfdx9EDIaQkq1bAas0lSWmeUWk
KvvRP/FVtfUHwIkTERqg9Zqgyry1x4QJ3Lgc7Okt41Cv9CGJFfgUuLmqRw5JVEV1l10WMT/+2vzn
BBdjigRHwWLnaLBIcukU7iyhA7LjSS0HAMmTzeK3MD5ocsCnvkMU8AT5Y+CejK4EDBmCgRHic/6A
spfi/YjjOHEGVG5PeGGZNXmSRvxZqR5ImEm6hr697z0igyUMZrpRDyUCr40QHvUt3R99JCQptzno
eKEKuZjRx5Ai2oszr1D1+1dfbnRY6bciTuA2RA6MEMxinzZU27Y4Xf2LerJcfg0PTu0GDhwWIHhW
nlM5BSF3A1oYNf0rO2+4rXxfz42fsL6HbzdLtrqJWF0SlUeOCOVMTCEV6W1sgjmMMMeSF+ehjrSR
91w9y+//dP34cCz/TnyWNcJTsq7Dp+R3GAlQPslAijbpARqRHrG2cKAiP4/0gYw2U2zBn9ithUT6
5ua/m7fL5KZpIL60Juckizg+0wwvNaSquHoE4hdssa2DvY1imxl/jORNJ6coUTEEV/OnqLFHAcdB
bx8mP6p05dkp8T2Dn2y3d2P+wpbM9T05mAK9UPq2ab0YTgnKnBFoQJRYu2wE576FBG0TVkHnwDj6
fbJeZx4TLcPkoq1SpsvTE3TFjYNIWqizAGmT1XCgTx1DR2pg6DdanOObYmbjbkVEEJzlywYAK+XA
daQJo43bGiNzV9M7XVvgfAmL9BQnFf5d8QAHbBg0s8LBcJ5qh33FMuiiHXI3lgM1LQFBmyRQxGS3
b75FfJp9g8Tgdl40DjnrDP8kGOVP7Q/3/RYzS9vpr8wHq2eVQxqiNDRkN7gDUZWrWAhx1jQnu98r
UDGjYLD7fd10h7Sh9MWN37raufi5ljRpJRJEx80Ko4+DGsKy0j+eHj9QCuDDhHG6CojuPOsJOCiU
ny54RonRIlMxrv+pAb8wCqtCxy0Ke8bKfGT7CR6DU3y2F5clRWj5tK4NBTmv1moMCGN90btTTfTM
MfcFg/0CBYanzzXYGEDHHmcwq5I40Oqe+RnOF6TXK6ZY9uEONu0w3QWTdT+nijm0qbLXiUQQm3be
DoMn+VgDqKA+OrogUHI6CIXT3TCmtEwWfPYChkQeuC25+X2sbiyDW5RhtddrUxkCB+6FxeKF45zU
/0zZ9Yeg3TEPIVP0ohdL7Qz5NHsc7fmVF9uoFngAoQN9q+E++82SurP5ztcJwFAL5e1a8NJj4naD
Ix48q4k4EvRmnR2Ns6L4wjpTcMYI3N9sV5NWU50voX3c/I2A2omuqAOkxUsfdT2gXPvh84fpEuNa
+3VJl7ycxVQoj50Mbz1MgofjMtiRhIZyQLgLyG8nV/Vk4u5pMp62UtWKIkHYFSFEm+fWiDi30+uP
7EogR4BA+H5JLhw/dWMQ2hxbaVzpJjdmbQE3sgjKApDVLMo1EWbfWPkX+q/roTxUzUbh/CmPt0A5
OwcbTngQN7/S9p+cBgj9NnHBjK2Np5jfVKjy9XyBvSPuvgIsiHRQSivzN287GRRv9oB3WQIGyrGP
aEk3sV9EV39P1zb0RzOKFdRvu8KImCYmbVsrWVzieuE/97MKgf2jHnb99yq0rYObaAxB2w91ykg8
qNoNXZee74tgyeX3kIkAeWeDge48XSXXnUAgeuqoirDhZFML5FXrpaUdX69xGFRZFsT0Aq26h4nT
vucQXQ/3JF5TXkILANB1chGkldAsRgwN4XLndONSBL2MA97RESarxbZwNwTLYrRqAPNpFXaQZuKq
6m/L+7NZaeoiKZluxPDF88s5OXT4mQ97YeCO9ATSl2fnLonFKWplBCrbEGGmehQpQLJBfFtuTDpK
uXXF/gtD0EdsL7+3ZZ7iiivcmDmpbfAniw4z/4sxXxWd+FhtkRWQSuVokq5y4g51ySZHVOQTLPlx
qc5trOPjEUEqjHhjgm3+BCcmaegov9Cd6oSsPbSQkEbFFfmRL0msqSkF4uehGUFWNvWKeF8LuC10
KCihUcNy8JWcv92tCQIApKIuo2yS++yey8qCMCe0tSJD9vU5e5QnICIP7NG+WlLOcn8n60/Fw8Iu
ZiQ3zMvQjL97679iy1tuUxSjYgKFu/YAAoJVt9J7BMXUgl82MpDK1zPZxGC34JFNeCwApq5X6Mz6
J5lN9yxaXdj2k/Z8vSW54wU4aK/8V0IBWCANUrTfs7RKOvHs5q0OK2i8DZIL/6yhZp3cdT3xRuUV
M83gn+MLK9aVQ/3inQbK2CpCK9sD9202iyFFe0nHXzexknH8yd2XFh0/lWzF3jcIsW7kJpLovvkT
OgIHUCAaR6OSYipnzLUl3duZ3Ip0VKN+7neMI3gD/XoS3E0FEbLI1ucMjRnQoaAbvklR8YaudxbU
x7HKJ75S1T4DkCCMAzWlznwwlKsbew/zM3nZ6pPkzKDTSnM+NsVDBvJa7d3IMwSRLoZP5/3kippA
mmDEL+9KZWna9mdepR05CmzjjllOEpXBgBr94U4k3dXuc7DPJxWPNv703tKYHh5R+0utgIKIJPwk
wnYZnRChnODQ+4SICg8RKDT50sNLa7/H63XZxtCpOtoy6hZpQ95hHnYDgAf46TwLhU6yg4VV/xHp
L/NnZeoBfHb0+jzFeeVBf4gkvk06hQAJbLmDeGyTlAjc7czT6nN2UgpLeiKSQ1iUNx5PVNr4hy91
h+IZAj3StJAHaGe0BquYz6YSGBQpw7ZJbW2tLcW6RmO6cDbUEtFx1nnesexcDoWHzVgpVCrSYBVl
x76ZPS3NCRps5xRqvO6nPiOQnhqj6gFeS8NCzi+dMprcR8nlTpLW3TBBnZE0VUa0MDDygVgqR2vv
kZ1cMgJO5ZdQzhF2jgCZfxX98vYLS5h5oxYIIe4TgIxGnuvtv8Qd4qZ0qkLkN7PFw0TuFwrLD/rS
DHwALpIBhjFHEQPLP1uoHxt3/T12FQcPsinqGHx4Sdgpf0RUveD7w75gDUJURC+Qrd8Gefp4dtzq
ga135pcTR1dMPJt27G6Kv4cfjYIP1Jwt2eaY4UnVPnmNZA6JtbBJRJh7UtDyvFegzxKmeb3Bcoap
sY5HOMXm7nysFjo9lnufDectDv+CngMv3t4CTjg9x2z021td9HOYGgtPgEHLv6qkgqYpjCCE5Adg
B2S5kEVqjgtqtAfmzOsKPHl7/f2SmlMk8KSWNpI7LTT1psujlVkx9FPKAKmu9UkDpSOiO2HRVf82
E1WtWfDwEI0Y7gNlOtjpawD6wUlSRSLsKWDWQMRk/SSiqfqEOw3q0YcGQyjmSkYJS/Qfi7IJ13+v
Mqqk+QzjMDOxsAVXbvmM4ShXIlYuoOuweK9jzzTIV0zK9SAvbxs+VKWnXfVZYvfvPJ6ub//iLowJ
FGkHp3G2uCaHR2vw58yATJgURwkWc1PF9IABP/uTB798mbQnsx4TsbZOnXELU7PakY1CuPNJG2mk
68M8eRGMYp7FcpDSQ2N9dCovBkEProNCJRPxl5rq163EUirtHmE/2aipS0zkonNgZg335K5urv+I
7raVjVtktHBwHfPRhs+fxcYA8XFhO5MdhsCuT7FRDUFuDXvDEop7BJmx/kMVqous8K7Iit3dDied
1jIlbZogF1U8Nq0GsXkE2ISma7BGeHqukmvaGt0ObggUNSQSKjLWQ5/45wvbXWYzuKapLTaxLNyO
ZXT6TFHxS7tCIZv8rf/KchZg3sImuWun5I/6pmkFX2DjS8hGn09N8uDDxRru9/qmGdokuU5pf3Oo
VXt0s2tb2ApbdXNPC9lOaIIQ0j2+36vkuO+7ezgJ5oblavQ8QrBE9pedsYlRf0M3hi6bBeVrt7x3
2pJTMeNbfCPZw35Xr0XWHbViAoO7MAG6FeRF5LX4Wn49ANmVoZx60TQQH0aND9aFTcjDv4TwtODM
g/+HSqk3058Bn0l7WaWq0vcnuZfb46v7VVoWAdOGVteFizhNuQL8/JDpO9oONtUb4u0aRXNnV/Zs
NfZRlRwSLxgo82VQbhrcIgg9vq92Jtp+Zfpva1CXc2z4MZbBcjyV042TBdRL9iiP/O6hCvf1E/cz
FkSlmgzWnKzH5opcYi/xnxgVc4+c9bZrEKSBrHbHxNKFHJ9QPwK1Wl9Pi6iQj/aIUmnQi/SrGjGJ
kNAJoGLyVfR3usptviLu9ckN0KAUVP6EjKV2E6AFnV8G+M0ELho9ApQEe0+mDfW4zQetiO0zdYWV
QsXzIo5rLcoCiFWvgzXyF8BO4IK6zbbo0VyJTonEzOkr5JFVorVpsoehCKWm00XXZaS6DmcEsEdu
4jQrM+Hd2RCsuwyxeiY9O10ztoBbnGjsu5K6rIItYMO3MJhevs5TDggiqXm/87oTug07Mg7UW66V
AOpwxva2tjnxCu77BIjQ1LTd3yECURM6OwpXZxj0lpO4JRouPu48pFQ0Lj0qcdRUDVR47sSGC79H
ryayWoZsKTdqh2Lvsna0UoQ5IWV9HL8D1Rsqm7d06NlXVhob3WfxtQu6pWn89PFk1DywwJkW9365
E2iqE5QY57wzYWWEsmYl9x4X5+5vNFDYae0QzrxRLnfd3Wv5tZixP1Ls16ckBqidTYQzZuNznCO3
eOKlTcFGJnm6iP24CPpz/tzavosGQ0xfnqem7/HWTgMutl5i+wQ5jtOvqs1JkOfPJapDjL/aAsAk
wsBIAFpc+NwaOiIZPpGtZSCAff+pzNwphQ/3lDU772Jg36papLUGKxUYJ60s3y6Tf0p1EVY7/6IA
LYjjBIWJw8DJKrKWtTm0LTGMO0gDcvTD+3o3TLmOWdp8iDXU342E9R6lfhsRm+UZYBWstSlN/GBg
EO9WBD+mVB0YICd49YJyTaex25V82xSYuLLCsUSeU1+kcMRnpsRVFqEfmOQZwnvfhyP2NvdixJkH
8DwZJ3l0S63sT4k8nq+Mol9EB1Y7LQTRzwzNBbc3aMRt8EhjsqmyvKLAg/OaCWO/RQfeTSSe6cpO
mGAWdyYrBtmhkqYZvGHJYMWUMF8z4vB7f+obvp/pj4eNx7KyvztB45wWsHClYkEfdEKHfKtsaA9J
1C9YnWBH0655RDvlvXmS5BlC/exi6Q7f68NAthfNQG+Mh1lRzpzqbVRBI9DS4rgoorvFrvtkI4UB
RoHF8UGxoKMLYfYVSCLZb70rhd6njmH5xaYQpdjbhAqhQoqk9BaQ+vxZBohrH1cQAbbDFPOeBtfx
Fku/YywSTXWv6LRjXm5ZE+AD+3rucHRI+AEM/BtUVy/mlwfFhbvR9PP9xG63l/paCs7P3RPmmP7d
xFvRd2RYGV4rkgM2UabOqT16zQutK4MDJzNWSC5fbTfCcBvj/5BFrQd7HCYbZjjDN/+Xyt5jI17D
YHMSB7pTkqghEL7uxPpB15Qx4q2KEWHh3bb5q58Pji1HLFPhGrcwaSflpmAalVk5QUvGVoFFqiMB
LTV5HUcIMFbnNwnobj0+LmfFVvziBmrNs0clWsOcbFCw/oIbc+PM4nbhExlzNunWY6ZUg4+6noTO
QaJrbYtjBSt7/XOFnupsvvqjxBAjpoA3Y/1lU1Q7FUB7Sk+6ntrN+fBO7mPcOqqjK+kPXnzsst8h
eFAWHKcG9pq2wvqKzIuMVY57dbCEhaiYB3w3e/MZGiyev0S7sBLutYN2ce0nsIkVeDPinpGrMzec
YrUOjA92GTwbKZpvw/ZJ8nVdypK2CZGeGbyLaCCgyN/ZL2JuxrGmVwEyU00YhRVv2r3io4A5KDid
U7alX5/pSGttz77MHKue3oVLBbxD5nYLqkp001Fhc4UiALNiaeci6XkymfxVJXHMdITniJKpbTQI
HDJuQKni0Ob80mkOhEhBhp1khcY3mrsPpk5BtmBbq2tMQycP0kHnALVBx/xQ7qiwz6UVM9ApVn9M
9bgBh4Fh99Un7TvXhE0NjYU2FJnBSSDrtslBp2oYRvbxyNRnTW67avE9vx0FmXCy0XRcSaS8Bnsp
Tus3pZhSnmL3gXq5l9MJV7hjPSKwm8oGv8wk/2PdpkNVW7dXw/ehl4MzD8tdJ/FUw5AiyqmcPEG5
6l1bMrjBFBX2kr0ILXBKBQAFHcTtZv4f4fe+aYadNzkQUIzrdJAhnHNqgv0t2dr+eTZd1sRUVIXh
2HkFOqO+IOOqVbK/p30dG7WVXquq+JbCrI9o5UAshKTkFGmUEfdQ5ytp0cUjCTIF7xSOlCFYz99W
5sIX5VtPIzDzfeHfloO57JjiJttIGS9V1v/Dk+VbyM5Zs9BeOOL5Q2xG2lXBgIwi0k6bZ9zbNCxR
osQY4pXHRfjM5GBGRREbL5hT7PHj7viYP1o7M02tyav1Kx+g3LlHmnXUpuDI92slgmMuRt7yHw5W
TJSSiQlyLCxjdLUqF3p2QMqxtMhZlYkMtzBgfvPdc9UvkWJ29gGffAkJU9KGyaV9dSF4Is3ftIiC
aSYVkQCXsWmBfoqw8KBJDLg++tPQ5mxvWrSQOtnv/i9CwnAKun5ZzJdYnym4frLAb7/aiDoXE+aE
V121Tv7li/VFwKwqyy+VXqCrdYBUaeQjyVrgiSFuK/Mnz5rnOo0iTsAMhbzJt91arDgsPnNrGxos
rrvKzurDMXX3wJ4ghOHgEeW0yEdtTG3p//y3yZfWTgdYG8kKfKvPBeyA1n3Ck0gNmsL7hrfWjVq3
Y9vZmD+AKL+nzIhcs86fP6O6c/snE2J7EPTmaKXSeY90lTp+xo8Ze0feFNeeQw99WvIO8CZ8ZVk9
54CNFieA6QbCtJfLRn7pzpMgmvcY2q6K0hC+XEGEVw2iTCV9kUPsDwNsIq2YfHlg2A6h48k9RCzV
O8XBPnlvXze4h9uv8qNvLWkpCARFwL9Nq9Yn0nBS1PMVI6HtCvqWDZJpY8kyEwluulq1QDOSTzBk
dg0HytMbr8E3u9jsAu7/BoY7OSqsB+Caj/HtRh+m6aQFm9yVPFz4/+Bj4jdaXdaOyfoogpqa+9y9
yfvbFIgIJAM+rSlqB0kzcFXFqarBA3RTvz5mDm637ZP6VOjef7w5OGu2G+LxQvRwv40i5fusZjlw
/Lu22oFGvm+dIqNxFxGzGmHP29uYxutL8v7nfW8+wi4xCJWjuoxoqo0AIPs98GhlFaULeCOVxX6p
PqOd7cWmorzNm9CzWGHeD4B6D/s577bDsaugBf1e62kLCJxZote1tXv5vsEnR7/FneBY1driFv6u
QUOpt2oekJ1W6R0SS94w2tQdp7UHKF2uUWK2Qcet4CEMSN8Fc3Z0YhAC7M3GkKZHV7D79NOmF5Xw
dZ24+Rlrc3MERZ34mZwdCuVU7hZuS+NrKr4a5g5OQ2Dw9l6NB26T+zaLr0KwmtKzI39bPvLVDZIi
Vme1UAo4bwdb5X5Ued0M7VHj3KP6DNpfZ8GZXGXA/R5iDM9n3bIE49HZUoZ6b9CiwsmfKNe8XexV
Ix8sEJkLEA19CBsHJ7eBIeokI1f/iY4Zrkzr8tX5yAaqUBRRUwsLno+yO1tr5ZOrHXImL/e26zxc
SEi9q9G1n6cUAD9kIPrBx0b8jQsXIyVG1L0dc7DtbA5akTUNSgvK/WaacMygfMz1+NMCG6J6PoAu
jc4dqyW3wx2t8Qbe9pMosUishuSRwgS0pPy9qi+NcuJ6e8Lr0nEVrJBfICK4QHuiy9TlWOHGSz/R
rYBz3ai6X1r6xk09ER2lukSPS6d1tPKAC6l8kX81sna7AHbOx1Ksk8iobcv42rbbvNVYgSjhUCkb
fvRFMQxpYTUUt0M8Khlq12M++z2IXpzhEWqp/vLlhaSS+fHKuCNK4b4iZhc1sZxvf00ZLwCQ/7rN
Z3FAPIgbCIKTBfCeYT+mT/iU5HCy8t7Bq5nrr3yPf1vFt/2SF/t/UWS9YvFGPOJTFYjHrxvBNYlk
NSrm03GPPjCFjpJeGyZ8YioLH2Dr3/ln61Jd0rptLLXHmlbiNwi8zP34d5ayOLiRandlcw54cBFO
27VfCdthRB1HBH5qJv6iUHmQumqOg9HCC7RA8he8muPtGQVzHZw8CZPt4bTkIpfWx+muyhbpk36j
+gPKLb4A2LYKCbO3unISml4c4WTchUE+61J9wpF+foDDeHYVkngOFtnLUbpsZR4QVOSK/lmokUc8
L/RAosQfLBjc0QmOPerCbXGWAKanyeUDTjitPA/9pvNkPC5HIXXBxsGFz2ukWMUAaAg7pvjc61nJ
JcAj+GLnzyKyhwKMuxPOBCIldiT34yZZ3bnqsUcV3s3LPZpOuWlfArmCSYnTEHCuul1PvE3RhN5s
mT3ZkkCOGR2MOxe9K2+q1oo3jGi4hpRqE6b95AFSabFDnAWhQho7jJNfmnTKyKWkNs8Qw+m1I93m
SSH+ew9GDWNijoonWLA6czPUz2m3kBPxSDP0FOAwVCWgUs+eeB2gQgN4BPd2zZnJ+BKLZwv3Q1i0
i9rpkVDpgD2esNgvaJnr4hrKfScfVMxblKdHfKFYWuHK90J6yZqut9AQ7PVKpUEvg5tiOQbVsjRy
+akTjcmA0feVzeKR9vPOo7QqUsvUK4qPKIbRtYQ372epQF71fy4WGpAxcclYP8xwxbHZprxwBpFQ
WoN5BSBPzBSrL/kjZ3MSdrqxQPDsSLLe/SjYmHMJemNi5hWZ9npTGsBqJrcO+vufeqmsIagwPBI1
iLo8r0aLfDh8L9zmiAgMxE6U6vBLN+ZID/tKIvji28+tCAKmRIxdrrNenoLt1PDsdz90EglMHyNd
gYda22fxD7A13Vzku+b9T3BmV6EiWzgk4lZRvbSIMBoVM2uaY2lX4lcqXrntGvsTeXDg2FZCa0yC
WvIXSkugBFd25KjCbwzO2e5cgGoOPZihXFXjqt8/vuikwgV9mbmr8RswBGUBhI0+FAtgm6pIwk2S
vtV59aU3AMOe7FfITpfrt+ZZk2+qS8XN4nBfdogU3MLCEgVCjxGAoBhV+/FhyRAVv3/zikxMFFTZ
H1UpOjRzNMamPsv7D99uVQLudIvU8ZI2f+Uun4SQo4oy2TzKoecebFAurZKvlTyG6QHCBFelisAh
PnHxhHn1qdr6p3XHCe0PLbvlCFtZbYcirgmeUBWWMJYpo24XpEWqv/lveDd0NzVjkiA4YkSffPDC
ngMJHiOh/9nUvqPgL2weVQlpl3kRD9+82j5NN9fCocLTuM1u+uKdV/3lCcTQGHpXVnXMQ4fE9nW3
FgPsUm+uetc9pUns4XCy108LE/IxJRdi1gLJJ8IsJ/iqNWjA6YTlKPyDjrdcrGa+hmAlTLHTh59a
7tP/IYOSycw8YQ9JBuxIrVhBeR4L7ib7Zg9e5QYfcsxUUjCotkGx+8hLvPUg6YJA/T3Fe90/YH7d
jnW1Mj7dCVWroFwI7fCub4Z+xmTBaMl2eS+DWhnjMfUeSM7j7Xi3zpzI7mWKFi9MH/lWbmjD2U6J
1MgiqhF/XE72najU2WWmqqTZjt7KiUimWE2ydacXH51T2tgrvrODDRmeablgEFlMbhMycu+qFtLc
I8tR3G0wsjl/DyTZdkjKTqmvFXtaNDi4Yf716FoGJU+CuQSEmKi2mTT7H4ELR5oHD/v+l6M074ei
SVbbFTDoni5TBdD8BrJH5ATfibVzAsiVjVu6PXjREZivEkbeMorWlQeEE8UXk60cDMWs7Sb34iEz
GZS8d9BS0CsvZOVnT18kHS75rq4bskf6yynqJ2NKclquwOAFcZuIJFu1JarIqmZbIxqq2aA+Y1gN
oeIdseIHFr1HieCOcj6c/Au04829bcB11DMnOS6e+RxFIdLKAAzvekhT9qyCg1rZXm2YCfoR4sgo
1K+JouK3q116eQkhqAn2ANULs2J1S1gMpVuy/KW+dfqLIUN6lFhQmMn/4EsVe78EPp48yXQsD0N+
txmKQN5SfFD0XqXLopHmQ9gLgmlkeoLmv3y2uO4L+QSbmmg7qPlktiIcUl5d4CZMa2e+NYwZyFQr
2lSLbcTRs3ViE4F1DwLzXI2Hr+LKtq1fR6o5ecoFW7jq5uJE6PYAj12FxD1lYCzOCBSkBMVtRKem
jJaQpT0SrpV2CgyHjA98UMeB73EQKMEjINHODLlEzniWXXV+gjydyjhMk0MZiV1UW6Pfx4HCSiiB
1wMo2tv0PrZz9KyyqzYydKVSgtDYdK6XclAfVCzD9T/l3JpwHONTup0z/XS8Gs7vnYkhECilZEAQ
3cjBKY66Dz/IEy3NLs3U6HnilUOF2CDK42KiHKIEs5VikVbtSTiNl5qTrPRK+WC+PVeeKz3iT0aG
hcM4JIvlXR2pCvKXRP6Yv0+cb7jRvzdpsu4rv4yMdPUCkJlM6x4JkTynnrhpSqt6YG99xopLuQnl
/XB4IJiFPP5/gaZfzLdS0Rxa27sOca7zLOqCB7JC6ayJXBifJiRkTNigRXrDnrwFf+2VxpTnMUQS
stPlJ5oJepxBjtiiB8bPDyplxm8PlqF6nro6p0J3CPmsuNlhi4u72jgNrvsMzJynEVaLIpazSLQV
lvRXuoJKhk4O69P0G3V4/Ilbs2NjRPkUE3eBpmtRNGlf1sMAsLJbXy2anUbCmIfIcKkWYKkKSyXE
CTJNPE4sUg8etzWvEtk0zbX4VcDlDc9atiKRZA5R5vUZYOeyz5EqRK2jjYPvRg0zBJ+fv6J36lKY
pGxtGfI1IyR6XDA9r9Y1YpcV/Key0nfqSaQqZvQwfypItigIH5I+l1QNfqIH6bxPE1sbGex6uncu
R6UEOVWAVFjCi9mUATb0TcBohc6IwigGViAjKHD7RBJNTgFNVep0idBJh2SKh3Q6CapEk6qvlwFs
HALxKALgyGQnI/XUWyX5WPcJ6cI+ifq8XK1DTeDUVEEHIawpm9fj5HfVsmeP/md1HnUlLV7+XKSz
fXnJEQZT2E9VgT9hpOwhlGdqzp7fpBAmEKCrOCYjwHPmj/gCgslvaXxMXsvxLiwHHQsfgmA76cYz
AGY5XxVpO7vKBXnsyXbd3zUARvJ/g0BzHDmxeYppo+I5abnukBSJL17ld4GDXPKt6IGwYNzY6Rxb
GWc5obD/r9mdRdRflxHedwkKLS1y+pG5MMQ0y+F3WoAlODPvrt8Lb8EfLOXSZXR28OCZ5SAN8Iof
ZlYfHo/9ZdlBddTRGAUjsYoUqlhJi+VI7f+C6ZzPshN0QYmUtKVBEmwAzjOWwXVlG6urZ9R1r+/E
savpqjNgRgU9LQjlt0P+tIbncNrvuvjfc56eJjYxrkCxyPwQwJGIyDfaqpcRWhhmq6mdPFTOA88q
d4LmVsvqAGAHfPRpygwZha2C/nNgAwJrpQVuRwiAXOaR9AknoSNRP8QgdZwal7qTqqrLzndh8t7U
ystXiFENuR9WSbZ62hkxjM5/e70nQXmoWXfeJ3b4R1MkHkUXBYlB91pGCo/TIKcqDapvhgLz4YUd
vUQF0up73H8xGs8yn4gY072jwmniWlmFdmgiW55647lMe1Hk0Ans6OLqdI2PYCMo9BGl9fgPVcqr
0i9UpzTiz1NIjbdg8vaIajZn8KmNaNHZ9yS0LIytQu8rfwZPeS8HrgG+104cDD+kzoGrgl25as/W
tXl+6Tu3iDE1zEBOm3F9DhvYVu85MQFcm4ynhSG9Nf/a4n7M5yBj83ds8PoNH0nn+9gcYlRD/xeK
zDNO2xWT0X6eB4kwJ/oClC7LECSlFejZBv0Ta/7kXH4nqq6w8ncAxL3ADdSvCl52/w1XRPo/8Ee3
hYPsglV6NN222QUPYJX4q0iQnfpztL7HxqEvSVx2HTCgkxvBrRqGtPItUojlzyE5peFJNRrJChSg
uyDIQmHx3YJl/EXkjyjJKH4s8IOVI6wjQ4HEZEBrC4U0VT/ukM3w1hYWssS8+AoEvHmtSuw1lDq5
hp0coDlUmXIENIblZE9B7O6IPoEW82rh+V/KjlIYq1OxK6ogkBZAfGIp+rt8uXcJUPX/NJdAsxVR
B6GezC0DcAPcjlRDbv6lfIGU8qeTsZ5CkrMgE+ml1ov/iFS4vX6QET6U9jY6gXvveXWmXspkiLhD
+LmxipAfyZQmz/oKRqxwXn4TnxSf84F2sSb8kiqUswPtEdTlSEOmc3vyDjUpfH708vwRAPRjOt9l
oGjgz4IxEzxoXXHfNYGiqdY2/WHSZgjiANHe4xfDHy7tdkwftehU1oeQSo4RC9+tnw3Rs4e24Ob6
KcWcoAqTJDtAJuBq/Ufr+/nExe6LxmBzwlYnZHEPfn5mzth3///+WokJh89Q9kiKtV0z1HEPRVQv
rCLp9FLVgcU87EHlByHkNpSJXLOjrTJYpFoM7XEgqc++NuM8eZ6eGrajN35SEZZ9xs3jECh9hbOp
f2uLp5/2NLlG/YFAduGSbtmOZaP7dCWcOV26jj6/Vt04bF6js+8RiAlhGePTABbau4tlXOrW5WHg
hX5TjxuCZrJdVOZ1DE691GZoNmPhBBGbJDCyl4/N1PhQemaCu/izD+m8N3KA8Y5/YH+2Sec6Gys9
uw9ZFZooPSufxMRxJHutTbOMcw2wLazIlf37qjVdBGV1pVdkdbb40+GVUWpQnt/gnslz8ELUuwpC
YLuBLZylJQ9FcPf3g3uoMOFGN0ARcaMspIywQT5c0XjEXvO2wbw4+nUO+eQZriBseFP0RVj9FX1a
SsLuefKMiBc9yv3flCCr72YaUBKd/Q0EEanpzNEHjXsuHbeuAYQTbPU2hnOTxjA2kZVXyAGn3+/V
dDDGsGjhRiRd3YgyCi3zV+EFh5suTGEAtgkSE3qAG+XmIUyW26CblOF8Munu5QQKKrnRsVgPjrqV
leoJraCn2CfTrSldh3nbPMlsAcFJa5ElHnDvRK7kL06d8jh18dq8B0wrhjFlga/Kg3v6i56t1xi3
k5saIjWlWTPSO1vdvTEQmMAq+wsNVDk7vF4YcjW9U57TpTGo+RNdVzeoVbAD44pbjvst5elThWxx
EVaM4/3DiDQBOqZTR4op37HMm0WupDYwsOVSk5yQqMr/PQnZnc3zmFVg2igoqVOlks2V/FFmAWuf
VwUTO/FNUTczKKI00CmkPM7bid3jqNptgyITvYxOl9Ch9F+mLYYr3XGYU2b22yrIcrMz/FYCstMp
wkYt/zCpj6isDPjyr7LiV5zKoe7iC/kz+rRqxMXDe3tA/E99up8busJQTQA4emoEzqIWs++ZR6Ct
mhdfnZSZSjhsrInZrQQmQHFyfGLw6lhU+YzznNkSPBPB+Ud4medt1nJYrKF0BpSko4RMs33YwaFu
zDG6TaY8lnea9gmNihaow8elSB78hzLr8AaTRdjWsZumyQhaZ/MNYiN4RDivfq9T4Uz4+12jKY7K
ncTpbXzoZU3sE19T9joStu4t7SUDVG0HCIe6b0xdenHLyinw19B4tofGL+NCr2l0EgjTLyWh59o1
FD9DBtvcAZXxa5OVnzSXfR1BL7NMsSLzOf7AE+Ludgnu3iPtVPUJeODKgg1IUqxebSJcqYwvkcRz
cWItwemRy3O2yl9H7CF7YmxsaW0J7jjPMpDAn0MqPlNIP60tYZ3pAx+uYm1myF5i4qRCCBu2Veqd
scxZHVwqo9VHxksibbYdRcmL3BGx/3RNnDlHFVkSL7PxdV8RSw1Z3QlDXhZBtOCvGhxag+a2mB2B
etof+r3CcWEcJA99SMt2gEg9tyZAWE/dh8Rv4FTBypilljqgkGHCV1y7dIEeMfMEHgvZ7NZVemwY
uiACKhmbu/HMaPsBvpr8e90MZyLckaENqfJ/pWpgjY/yR8IsNjeFLllIn7ZqbN50wOGSMhmf9j8u
xArxGhgctgVGTgzUfUiosi47BCsfGwjVXEaNzEBmr4/MC/hm/hJluJ6VFTsgHkSJ2dXQB1hMLNrc
EM3FNvpcKoy6BQZAqWw/3WifBjCbEYtbgKFaoa5xsjRKbrTJRiZ+QU+scObQLhf1A9R9ONY1uFTr
NpZ8S8LrlFpCkghO2xAClqQrTyvTIpWfFcw4FpJwnjInBlUEM9r0DFFyM9ZwgzExPAdWkPvzPU1M
hi3eU5+AxzpZ6rplP45KIiJXDY4OsOkXpoZSDk2h7Zv63bA72a42/D1z7IR9ff/tWKunSecSbbBc
IKn6g+zkEKu3ASFmTl0/GYiiDO22VVqGjJa18sJofx+kyNXZj/NjeFIYi5IzpGR7hYCcsz032KIV
P71CiteTEESe4w2Vi6jyY8RTH4Ukd7IRJIpB6vGEeDT3l2qm6sStDHVJwfzthKoUNLy6R5L0Ldxv
ZdPkP/7lN0J/t/SbE8NXAL9yy3j2aUKCX6b6uWA4uOtVMY1gNihXuW4PHX2maLckTj6A5Pbfkf7p
c59YaNtKGedAN8sActZWQzupRQebs0LK+R2nPtM7EwwzzduTbx84ybcb6Fy0ZOLjjxBHafZGRHCg
PX2fVN8+xGtLc/cyH+sQPym7uFHXgov5SIMIT4KyZpYz3MFkympZ0kytNoi87us5JjUR+eVWmN2P
OY0VUywKHuMQ4gXyh1sfetNLC8suIdqIbzhVl/tc9+vP/BDnhu7jvUudhoSw5Wyl8qLV1l2PQbBj
rcje8W/60Zr6VxqHjYoJbXKBLVdOkMeBMvLHobJIkjT2SqocHnlu+pmllN9HqU/PQhA+m6mGoDEx
JwdD9xRmkuIQgcT29qUhgyrhmDrEIk+uj0JFMFlN3kBZNVP1rHxFL4039k7cyXFDbappljcoeMXQ
7vNNyvPJY27LyjJ0BXLQ5vd8ziGffSMyVzSpOVe3CahFxo0TGXSL8lj8rLxtkrrdB9WS1lmfcqWR
58KwQ18oo3keUbrrJS1lTwX8rOF+41Hn8USCsrGNwfGQdnXCEaKGVXKHMowzkBjgb+qfKqOmkSsG
N+KHjyNJMDIkVxSddXdGDhAbFf0N2Ui00SWcefhKwgg3edlp3IjCjLYyh2PzIIaaIK9jmsZPxWo7
Y2zLZyLeif/0vAwtE3NXaBm8JL2JrCP1VQrjLS/2im/UjxnZ1SL8BpxfqB/JzkpxjkpTFQ+7wgLR
9xznCdYziTBBwcHpeyQvpODl4gcptlzg5s88GRIEW6l6bhkg77uniGnYwOmjgLqDzqiyBSx1BC1c
pTDZiodGxJ/Umj0dn90w2cRj3kKEslj50uHyrnWCF2aMnHEMFFNTNfFstnccad0p9zXEXgdKoLC4
1ZuLkY7BF4xJXuHCu/t/LdK3x5FQ6WUZRMDANT433tagZkVHskZFrB+J+BRh1fMu0ZVIFvt/lCiy
OIQj/88HPNabM5mPT91EFE7A1AIufsszZvcMF862wfRsNc9ZcPUNNnuLnGYtbQM1YcDxA+0m8Ebu
nDwxHE9R0zxhXO+PznqpJkNkDWUUw6EThjarolE1A39n7yKhREtvlI5KdsqrtMGYFPLWpoqBX37+
itU7ogFC84eEe1k4n4A+85yGt6XI+S9WgCwY6nDfVdMcuYKrZBzwhX6RYrJmhGKeVIw5zD07rQSe
qzpty0sPCYBwQAuH79IiuMz09qHLjRtmPHJA4ky0PhFKIaIVQNQaHpoTndW/bQ4XyHSCywO3FpJM
SVXpePNiBl8aGg+04ruJIB68hj+r6TPkKi0M1tG1tljZdNgBvZQOukOt8P1UCukM49GzmRJ3Ndmr
lfWuQvdE2S8N5YQYgrljqvLQ7nMZ7SI99t01bsMZtmhQgo9HUcXBi+n8w8MiqcYR6V5lzHL4VPW0
KQz5KYI5ykPsd6Wv/0QJocZ9/Y6UAwZpW15aFe4zNW0lYcgIqltWGGamE4ZTwhDXZPZhuSN5E2Kl
0d/LOBUHIvagrkgsCTMZKTVlbPAmYVw/8MERwxhRPFfFwsjeaOBMZXv95yjjzKcDhze0PCkYooFE
fsSCBWVGxVSbIY5DVRWefyYyya53tKlbRKr+s1DFOcAVe82IyLzoL7ydCZdoEyXxHUVNHPdDbpgG
zWs8sJYLg82JVjG4Nmk7P9OH6hkwpIAl3TRuhbnZns5o0jlGWlhHTk7PMo1tKXe+CK6uOHfIRSWs
+uLhKYYxxydSYWWH3MX/3WHqJ7IsPNdnM+LrL/4FM9vASzvTtMem9GcIMnqYXZc29jOix1gxpD1m
u6FhEaWKwRbDEZ9lp1fgB4ILig2PRBdNEaWQBuiotOIZsNazvCmVSb5I7z2TXY9IhWIwnwN/xklc
b2TRi0Cqcs7ZSfteY85YhtIvAEBleUcWSMedQpJL4UqOBtxy0NVc7sCjTLMiNhU6dAZag2c2nVIP
tgK0MpWQBio8n2sP6aNUqx7amA+PTRE+vT/oFhMSrR6eyuqLuzvyfFNLGpn8tfCEJouEjnu8VWs8
UnEWLHL0bNPGDEc7IWhVGxbnOAaswPRxE5wT/4pJIg+JDCJhwmnkkXAx795+lTg2Z35wz4BZbyo0
g7ueAo1l2s73miLafGx9hxubQ28XtxipTK+StRgBQi0o0guQ3uor2+6beTW7OCYrRvKQ/iy6YS69
NeLGbPCX5B7I96y5AjCMR8TFy9CCzUBecgz7q9lwTYvDd8AzjkGb0fWeHqn1VVnmJi6tzfox83kv
e49dr3Giq6e4ucoiTy1X9XEyUnVr32JiuMkbxelKVzoeooquCXJEF/ayYvLaQ9L1zcrMSHU6JD9B
D1HwPqHZTiOR8PxEsqy0d0Km75XBFOgupLtzkS4GdJAzTY7nUvLcTiY3NxBePRXlNM1MGR8/SSbs
ktqEOnsCeNSeetkasMNcqUEbcTVxH6xzTqGU16dI45YjwDxgzmzRGHjy9m/fzUgX9QVY3XNi+ui9
8LdWn0uz+kL8tusZFvknTx7Q+Ygsgyk8UoBM7tQMUWNG1n48smuZqjzWh+oLnTtA71jkHb/Cu1/r
yRvLJTsXzjureUD+Drz50rlgDXPlpKDU5UFnTgArklE0qJ/7HS4dtF8dP70k9jhEtAtiPIC6s6Wi
hx7wCGwzjRPh6yrC7enB9g+oN/rHCWxsoBL9TnDmVORylFGamij8+/R2b/Qv/+HPXWqBoMEWCsiX
kWkb1QwI/FVJazx6hP18MViujEA2qr52/KKsrxGcVQqlvkmA3oaL2r3jrUt3gfuDlLYPovsjhK1h
kBt5qIimnVxoSLVXA9b+b77y2YgHtZLUSnEKlWBlRnMWedx8tYobfGXCaoxijkReHUIV7V12XvDn
fIzctHNSn4TdFbhKNzPOQN1QCpaKoOInGMBYyXK0CIAoAVBZzKFuuntJUaRxNTVdNGjgH7UvS4ik
nPwlvCdeZFqqm7zso8J64PGMTqb3vPRkxZB++f2herxlNQLflUtz8arWy8Dt3LE+VZdEr7WjRjZ/
pOA8DrJb2wrKAnbsUU9H8dlMKsbumcvA38gGnp+216nFMAlYZInOSNHL6vspOf+PJLhQDhBtof1G
YSfVP1XX69ktwXKlcZ0kldy1hH0GBq3NpYBjVMuhLpx632BIXbjnXN/Yh/vICQXKH/QqjaQesxBR
gPt0wn8dPwwJyeO3dZyoTu4A48iEtLODVq/YcHuMeWiAJLFUedegm8aSMODVEPlKBO1pVP0wicCT
GcyDChRalAcFQkJpNXbspo/y9xeVLAoMGzhmJKRPRhqrTvNfIac7pbo3gSdCq9LtR0nywCxqoFbd
eN1QzitbNbdPNwvTaqdsF+rtKOq1JqhOJkoJu5Ex+Y+rS8i0A6oNlONcSDIu72uEfg9lSF+OrbZ0
m8vziyG0dsGtkKfmaBEYmCqtXYXlu2lC02rAYawrflvXPSw7BF5zU0cwEPB1S2YX/T7JlOqhu2h+
4rw5UDq0+Y5gtlskrUKQcNyahxYu3ETvgA5PxEx5YSi1RdJyDJirzfuk17R+PowLSyYXNkv5z4F3
qLnuD+x8ZXMfhEXN8KORcabDZP+3Q6N6OU4viTfjKyLz5/Fe4Ixg9/jkAzA9xZXii5bdYCBqH7N/
LekCfZfNb/XUcsgaNYxsEFuAty8sVIwOuA2F+gc3uc5DsHsl4DTvirP5u0/IgQa1/BM/TYIBQsY5
swBWwg/Gn1nFbP6AbOovqEUA467J2Tg4yuUABDbofWxHEn2fZ8z5r3OS/OaXfoW3DmTVfxAkiUEk
pjQPo7nDgdkOb9XbS0sqJqENrY/Bqlv5oy784Byp0H3Q20TAPUtLPpmvpHNxETWwVLBVRat95zZZ
uSkpvsfV7Ouiw86LFSTz9RLxckAiwraNK6YRwp8TsK9rdUVyYTuJT08ZyUrsVnRUjbkA4kDPxDGC
VgvIQH9oW0YgZ7+KBMTcXvpRJ6B1UnlnwkP2czxRuJnrOCXbqgfeke4LlFo+8HfP1qRyUtCD/3Wv
bS86zgUwu/8iwrJapIX3KRI7Zg6zV2VEMl5YsUuccJdPNnsqJY/PGrvmul9lv9rdSMZzuXacYc04
V1eaeYzxQLGEolgifKp+zGNmDYdQTy7ugMPj/q0plnLoq40gyW5cIURF4/AkCJ6NQJddUii1Mm4a
B9Sifm69iCYbs7RGqhchSHAQomrw18reHDQbk0f6syp5Ypz38DtLAdep1MNOGgeL4+H4gssVItBv
yW3njYitys9TkC49HqHxst0mAH1BDgXOmLTKBalx6spd8PekXVI2/upf1GkjU2+SV5kpa2zZ8hRi
98MsKD9FrDvNR//ixptLmWtmUJ3xEuoID8RCE59f7L48dj8+/qmNSzwGndMVetGUpjjlmq5FiP+w
PaIBNkhnDZQOXjKpzL1uBki7fBykdXD1lNe/3ZAQT4Sv+CXI/PuQHPp6UeHRu0Byh0uK/qmQ1JNl
UshKDJkwNhhZrHQesYQl5fOa67eRcoUBbqoMakk39f/d31ncrgmgHQIGYQdRgF31wEzRqjJYZmS/
e0xV4t6C3JlGCzzYw5LBYrGS90Ac1bUy8RrqjjBp/Zm2OwniPMB9VoIGywEpIfOnffBNTXQxmJb+
bmLbWeee+lJIUd8dx4ggW5Q01vLGPJ453Wd5YlkeYI06yzvhyAso9V7Z7tG3RgErh6di2An4/kFT
HCMB6bP9a7wFj+H24K+P96aHhDOCRJRt4hIUIGr5X72owIs2m6PmcsBvFQSTmvGbTOsfa5ScG9o7
wAElKqIqy4iblpd+iUVUJNY636qGvyXkeowrgPPWI0Os6Xm6o9zM+IJ8PipNiKPMrNwTF2TRH6Nk
rOfJiiD2sZaijhKYxP5KllUu59JbMqe3O88SOzVn3gBQPLrAcik4PaxMXVO1EclcJMI0ZSyAT79e
yweLSPevvBIguhqxr+XvEhDkNJVfglNxSc75P30cF9b8CV/YraTSdzXaPtJ6VSO+hJbW57/JJZ8t
gGc4C50Bbb8ZBCv2w4kAGAkUmYXxRDdBlhscvwyvslbSzmQJWz/tcRN9keBisKwcLWjWcC+1bZyK
OAd7mE6NBK3Vg4585q+9qbnV3qp1XEyguzNamym36XNra5sNl+XYSv9Nl87UTCwpsFtHEn+Ou3GI
8e8/sgcGrdtVLhjkpC8TCYBnCSE145uwBx4AF2L2xnlTMgSIEZv3TJrDS6Mi9cmYBLtUNhS7c0Mm
6wxuBLFhEWTbK10v9iAjfvz5pZhLiBrEKqTTykl03C2FDZghGZLLEnltZx2HA45Z3/o3C8Waw4VM
JC0ZevgsGT435pfBviiGIFCi8nGpABV0oGZZNA+QtBt36TYh7Knktpm2GCT0HkkswChYJ91my2ME
ga8XQcZAcXa/IfhIhdc8VgsR6GogOgwF3Di+/twZKhXqzaHMAajJb1kiWOsx91D5gGpL6Y1XM/Cc
x79OOwGUxWFghfOmJdQP6QsCB638r9gbiLUGO/QzwS6JBNDv4mYIVhpepAmHl2CQ8DeU2Oi+bYmj
SCZwl38SAtJZ/ZRG7Qs7+Tkx+Rg0mtO4Sc2w7EkvBx3aGnr2vM7mIIx5I47j+FrQhgXD2AWFesdy
UEUDvnbA1XUsDbV9SkzK9kShrH4cd4O15mRG5lrOGXP4TU/dTJNkk7Na6bXmPg0Ej9XmihS1merG
eHrq58ofyGRWIEjEkZZYvz5yzThdXVV8GURMgWYDjVkFUb68VIONwlB+jucua8sxT476IHpZkPYJ
5x9tXXZ82KIFv/iIvdmIZzsCbRzvAleYRT9vuU69TAUKLUioh/3STRnzWS0jDrAiQwmeafoFyFcF
hIb4+xRVC9cVXuqhZQ2wzDwwsbMsjacfsQbmFsN2/BcD5wEyawkTmiFJqINVhxB3IMENR+zwntBy
cfOQnZHvvkzrtJH4dRXjyGf+G9dNXnUeWl1R06fIJyJo1WVd/GFQRg6Qo5V64OfxcUztOn/NkuS+
xrYvmz/dWlj3edLPQJEwf4UXxERHO78mFavgMrmwv2tucrOd8WX4R46Fu9Phc4AcAoSYHnbJJzJD
CDYBKE75/+xVWnd56f8PCc6mTwYTG4P/opnt05oNP61F8OW2SdQGVyPLzSI0FXc9YzIyzoUSkUHh
6iOAM/iB+6rufbdWsXA7Od0Gw6/aNE5+TmOo8Zq+VCL9YTuVAOxg1iwgPVn/atG8n+5Nboavigzl
GubdSleEqJlKbRH1vlSqKn0bIk/MphUu0c9+NXIr+JONsTwJm+MVmOLyg1JJDXpcPFvs1f/VCsF/
6hf+WNqmQkSFUAjMUVrKtqkEgVYFMKnuri4zMFy8Rv2VOCtcMmATt7I0Qjh6EM0LPCujEh/3zvGa
MQy7rOerZ5ehPlB3uPQIR8NarfFksCzGcbHlHPoQDi3n8cTKhDjuEryKRF+NLapV7pvx46CQbNH1
z9+WeKJeU89FjW2DBA72fOBIE3bvugM6XBD+LXKuVaAPnFXrWh7KvAIuKOfv78b9LeQS8c+/c6ay
ssBpIHwB6bnQQWljGLP1zC91M8gp0KPFIznF461Xu3m+wM99y7ucsigpS7mCekme/0M1knsjuUZX
K0gi3+CRY//U7Imvm+ND6Utazli27DSCrqEEzyYjR3IWfsysWKIePjWYZzgTSSzWWyEKDKprNsUI
MFqHch0wr+XbFn7lSYY/xTaq0YqTlN3j1Dd9PIR3YU9iSzXTNW2ZUuCP0E+f6S93YyoyNgsOIKvI
u4FDWTiXD/g8rDUeAVVa0gGJNJ94r64mE5D07/AwbE2zzLq4iO1EQs20b6FXth8DJiTE/AEb7uzv
5qaXpx/WpPX9UNdXkcrTy6btubTMV4scZp1FPOXcoIffS9R8vN4o17JzFJJF8Rf2p3TWTiaGvYyB
wWh4i+8oZyOl71lj/dRBWuDYTETo8IjYMnVGQ5uORl4woF+tTEI9bpK7pKYwNHZmrGgQYXOhzrQJ
bhkEM/u2eFaAYA7mYgKa3Ba32ssNUarI6Azc+57sjJpBNBpAGGOo7pRhbe/b1cUPPLsGiKnNNrNz
9e1UlmSxi3hX0mxfFkVf7fDmPo+hODQpaWqG6Nx6CYRh+OQL2+payABCFXuFtiza8py66VZuZ6hE
hH6yrbKa9iF9QudRqFu9JDcBuev5TIEgOKs6k8yHhX8jr6qfIEMEcqCGEzv/LgkaO8QNAeLCWHie
0MRJ7rzMo/X4GMAoeRqWraQA7IugYgtAZgOL/mf+tnT1E7E6FL2+vQ3aRrchjrKc5dd7bYK0jJd+
3l+OlfG7dZdO3oa4Yg6/1MwUnYWXN5HNNz6AETP8MCjQMq4cZHiHxGrvmz7VrZC4dNzMayBGdsdN
WyLj81EofvY76Kyl2zm9ay2h62qN5sXJtY9BdZ2jWC3cbknvXM/yHBJ51mes9xm1VulsGZfNXd0X
GEbv22FvacbMZPd41A72TiBHt96+g8LQu4/3/zf3iBAOsYjEBJclPC6v84ObT5S/M71rZIEUE+2g
xkwpzov9htbPHFETGBIO8tFAILqG783kb8NqTuYh2hggvIRgb3kJW7eHosCu63t85KmP2xmZ3yJZ
SL6+EUXCjQvO/DzqIhCT3wPjlxoepsoNlgFfDN8Rv+Au7qjwir6XAFwgJXXbuaRwtec1ghS0Jckj
7RoaXqjMzBXIsu7YmSVDLRHnBmM/auqBBjz+TL5jQi8qSOgaWaL4kV2U/mBR9pSKwwHAxQ+zYOiQ
mRb6Z9I3gk1J8ou0r3z+Qr8BkkJ7D3WTRmtnSz1ZQYRlIuWmBAiniYT5cpnbK3nim9TLT6tskRfY
ewz9YI2xiRWwKQntlQmisLyJ4VRGaz4DfKRQVJ2Wpdeqdc2nyhxhYisUGBiB2UpSh3zxcGqJEWh2
wJ1uldAFK2C8L2CNTYNNsIpX9XxTWuCeW79OP2jDOJ+QGyzWzVPM0OA08IvcSNoXo15ub71wVF5X
Mg8YCPPLiGO44H3XsuKt1xPnYorQ2UinUizPr17WGN4q1UsAZfdtFo7QRzeMbtEurZy1uUfcOysw
B4JdR+KsSiBhv3lMI4LDy/wQahf0EBXU10PXgT7S8SBDrHmkz0xNMDOppVi3h7wR7VpMtyM/1tph
cdIwMu5bdEldglGzJHTTO0XZwMoCtvfQHCuB8KIv/MdqYphMlTuBNh1GkkQfDNG6QhlUhnMwVgRE
7LFeKKLJzOn9JUYgNqkFARiD+AR5M6Xet9ptrHsKMmzWLDm1nWy1K7JcW/vXpuNDngrfepTQBoys
gz/UXEqePKrF2cwT63pAB5SZ8A+/6Tp9acbkgCbetwiH+SehnpCbkW/8IjXbh4+gzcghOWWHgdpK
hiLkqHS0Ni/+vysO1cTFV9CRztNVswGCcCgPU4IsxJhYHfe/7XVomzBOSfthW9nRLQC8S0548uJP
OK2jNbxm8LKQ3CGnpe9mjOhcRWRayS3Eri1Y8Ykr5tqJwH+PmpEEvgy+71Kj8XHY4NHR9hy7pRht
bFxCXgFlP1h4llEK8Ujktoe9F0KfMlazLFfKayh8cfhRjvdgo1AUPE47o3JV5ogJgAxTLpBLOkI6
bT5a7IvIxq88d6JiyVM/khuGw1xZKGPj2rJF78TP5MQWGeKE6pnS9r/IaFq0D9P/MrBY0R2QuFdc
GLOkSoyedjT2AkPuB+u7QfrAGlB+zV3eUHfPcXjec9nktHtdaSec/mxULzsnAQiuGOPB93aYqpMY
CXApZUkDQRuA2qMWgVd60PUSc5P3H2ID/N+eNeFR9iTLGDqlkcMv2YxzZ/2vIEFEnxAI8QPOkr4m
F/GylV88xOzBv5687vOo+KG9L3ADpLgbC1WOJJ49wUEewg54LAgkU6XmfhQC5STrr0hbUrENPP/W
wTBofRcwFaf0Z3jZV59PEdOuJDOrb5ZxPiV0ZVhZlKRvIy7oi+pdtovK9PKAWz9KU5x72FQ32bpW
8/DzL2n/+spyBfVv0/cSc1MXyUrEbI+5JKBEpeitLJzqToZjmUqNFWOy7BbvfvJ0X0XmkjT4cFPS
5zBqeeEMlgiwWG0YkVzkt+8Zw7JICm1RKbhSSEvJaM+c0zNMj9ASJQzN6Gw1d1q5S+/ct+01dXoU
JwDjuvHPgybPKnzemNSOYjEMWOTAB49GVaEEirTiZbyZwfj5gIKVmwrN5Rmvaz3OxtgoelOebFbt
E9a0fldvF6EpeFu0wCpt4IohpReMFmJaCefpeg9n0U+ZHHIXe+2aW+alFWi1207EYX/e+hNzEIOX
eQSLvXkUoJdZFMViGFPod/SHd1GbzTmIbUROCloYNrkQTP8R/IszHgeoeAa7ypqnVRHRYSV719CB
sVG2ZqyO3gxFxMCnhKSvLYgnFQ6ypzwPVgkxI8Fn4nOloIARbY/njIbGQbW5iJSRP4h1oDJD2Gqv
rOTAd7qNWIXHxrIxFcLxdNQ5QLomH0Pc/sm0ILqzMYOvycUdCEU5rcZJbqtWzPa/lJ7OdElv57Dq
z4aSYKISj1BwAkHmdgf9+qRLLL9PN3KNUjFcb+zjEpF5W5Ca5bIj7rIkwTlBY/+4DB2uaHLNbMTn
OfStCDJEW5CEh2ao+iIMY37Y6Xm4zJAa9l9tTrInKnBnhYuGE4egZhCWcnSB+CN5DnlF/JjwSJB4
ken6p0PUJQw1A201PwFCiNIEekhaYko+J+8SVC/J7LCLRLPFRNmLI2xV55UC3GulbAq4XahMCIT2
2axq8kAtnRaBoAcdBLTUI7jp/gTjxM1DGrs6+e7fyEiLh0i4lIx3wJwvnIWu4L+csdGZPgHYJmCa
XFwKg0D8Jpw5OpZ0Je25LeastYeWuGy21xLtNZbL0gh8DRV9lXsVWv73+dhlX6y4hktbtg/at+Bu
sqXmIoYgVSNQcT1ip0jJNhoImZ8iCFOVivwfnfB4/QdOPcZ2dycc+nXZfpmEoJlfp2IC5vpCpQxH
oziN349czgNwkmO7XgANGZcu/fKvIQrsxoLYhprrr0J7Xjb1y+wbxSLeiTTmSDw1nAN+WhkGiDpz
F3nR09fXGu9iHpTYnUf7SUSk+Uv7pa6JxqxY2LHZuQdNhWXNZjNY00LvpgnJqll87YHALOEoB18O
245c20Fg1jcGU5Jk6dG4gRWWWzdonbSy07VUrxGv6MQL7gH5b95uxBeKE2G83YTkrt9cZOFG9qm3
ZKillDdLEVC9zwF+1JHq7zAXF/vQ133+3/qr0rF+X7ml/PAQdq3hY3UofI++/+MG5bsi+rcXTYEo
t/gMtCxbODh4+FkqB/zXGcPpobb37//bGEpN5YLLt0oFmvtXcwahyzoBevkN8++BYwKfCLVTFKe0
waCmT+k4/Cj6Pk0zs7K5Nbo8Ba0BSURt5j34SOrR2Gn45nIBXRC+MBOCyOXdvsGo44Y4NccZf5oO
oWuddK//8X9TDVJNEmWchcvBjIni0VVqdXRpUxXdbbFnzb1eEsijcPUh0Scw1h/RsmUor7SQ+NjU
PqtXi8ekYWERMB7kmKvv+5HurroIokVP7T+iVx+NRTF9dLtZnaDIlcg50CORwFQNTHMct40jxnRI
m2HMNMdbQhVJzijuFJE/fI+TlJHW+w5AuLxGCa7KNrKQRAM8HeSqeZ7xFCWJPACnSkUpS8AoSh5F
gSuZEihqDjrkzwLm+/eC2S4U8bEuQRQPdtIr+1WS0IMuLlqrFFuCL+YvfvdwE44IL2RVvyzRxDND
nAZMsYXvqD3YhZwHH6KTBKKYuw5i0FoHiyDuDg9TTnM28aLhYsCcXOuUos0Kqa4gTd2tHVfCfbT2
8mxMOwPw4XPmkgU51+U82de1Fd47etcvpUFCMuFTcpg0fUcRpkxEj88y3R6lMLPrJmo0DuI9KqRu
4TSqgtxoYzl2aJwXf3rTXiPTbMzIAUBmyIiW2Ls2ZhElp5gbeOauze+jULdYK+b/lkyiYfyF1yp4
QcYAuGvn1MZK+AJ+tAv4rDNG2m4liCnLhDW+rkuVinbBzGplFFHTvGqozdH5TNofz4Zw66rfWeF8
OXrDSyBaj8fYzrqcI18tiwFCb0g5KFryckUtvRbJ/72Sl5uPe/OUL1AyPS6MgemLz7rHVO+TrDG+
ETl6wJy5haV/u5VZ35M2TCu+HLQgheGGY2mA2eOPMYLQ6XzQcUgPU7thGVvRQeJ9eEC1/LKZeVjs
KnfPiLLdS2U9aCFDt0t9Ma9Ewv5X8VPS/9kRMzGg8EYLFBtWeyNDBGB674QhywrhHZCvsONSJWMP
FUgjjMyB9P+YmK1tkd+MiKZq7/EKqwR5is5osgvnDBxLC+9ufX2vLATf1SsU2Ql1bdx2e0zFCBVg
d07a7QdjAZgdEKXph4sG+d38wVn43HSACrysPEm06rOjikpNjGUQW+zlJfO1QXF5/gbEXmojJEOk
62226WikY4+FAAsdGd/vUz/wvrAdsQaOglZ0B0zshM1USve1Q4WihvVfeXCIuTdCEbfRdRFsnueZ
7VS5fE6p4sVK0RJMEOo9qXzCdw7ysxBtH2lDW3/KyOxuZ+Vz/ZY4vIs/VFVdfTXgynBlPHM2bcJs
4QOSQ6nIioIwAVN+S5w4sm+iL8fPK/MX4ZMBdS/9O+iOG/qHDDlKtYx2+01nfvVV+HFHbGrruGuT
F1WBPynsTOvi2MbUrk4NxbC1RXfdFV5pzWjr5a/Ej7S+7f2ft496vG9os/y7KFZJByjwf2uu0lnu
QVSXy+mXVXY86eK0zeBdzAEg1eF4QwCH0Yn/AYWaCiVVDfeXdkLeim31ho8sxRcQWRgMg1QcIZMw
gNF4rPuBxuv5zYbd6rRKo+h/dRmU8yYsuv9UnUYSzrMSoVM5BnQcJlEXSwK/DGRc+veAlavY3LoB
IqkWKr6xxsIqN5tNL/oOaNjp2usSMtxm6ty43896M4xCQpatVYwItCn2iWmTa3D8hT2YM1TlA/4Q
rfGGqHLJhSppkmo/QaX5LeATzDSgzDtq7CgNhHv+zakDd55ZQVybK/heTVihSQyh9kw3+IlxtdEs
7mhcEViwEf51/o8mGloyjBP+tkSZU026s+jhVZlc3HqJY5aX3/LkK6/zoGP6yNY/GzJ0klgUWYfk
KpD8k5D8MKnTzSMNjrEElOrLCmHGf7rk5IhxA7dy5bTHNZXDFidMfCl4Uiky6dKnvXg6woY/T1hX
HuIRRQCiP/lA56rfjQk8QoPq5QA1yvdUKaUL2X7DOjwPCn81zhA0Jl5WULY9Jq6+FeZei+QNJEJ+
xYqXD78EKm4OOrjX9UF53BM3tR+7sQDj044dUrUmhUWT1yDpxa8bDWJdH3IQtKfOA5awVeBh/7zA
6AdBWjyISzFidLJ2dXQpl9x8MGdw/RmFFiOJ2CPKQlzu34ITttELyJonwRtaodCD/zF4PpvxZDXp
/ZO7Lj3NWivSjjUZL8uSeOq4tIdK6EtVUuqVMmaqAN9gVK6L0ScUErCTO/ZXw5VpqQTMTosLnDiU
BNkdcUXMCfBQ2G3dWhyTFtkRMt8zkxinm9Nf4Wwcbp1v25CtrdVs4wkEETZjvQEiPZQ3mZ5hZ7WB
C+KgfN7X1ammQKtqbpZaZtUkpj2b8cPFtdNO7wSsOZZTZKwLSkcddxRicMS5CGOq44J6BkmQXX6B
mhliMSUSVyYcOcdguncLcI7LbTkfXEkV2AoKKGJwl6f82vY5gTJjGuqB8uKo+EiQfIbpoC8GtEc1
/r7ej0qQNnl6iXxllV6K6S+lBKGk2NlB6UPMBoBnxpYHW3hMAj1aJG//yJR/wXUsbMj5//B3QrTE
2XqBZtwwE0aeTp8whF+zVkDA80lebH2Gcw3mVseDVBaFLo1mscbKPWjufTj+2qZQtfhNqgJzlW7r
hwuE9c4rRhtfwE8Ao+3HKrUcK2s95EhKRn3YZdonbN/QrezaeqhpqXakQIN7lx3uOsX5Is8aff3G
X4IqQjohlK9tlJQ/uDuYVYM3wMYLIfAtc5BDhG4YGiXh2jr5hVO6VBZUxWHRSKm3Z2UYhgHL5zEk
ERNfXFPgSejoFVZABTABHirUkjwuSfFcRiMgE+pH4V/8Auvs2Po44WTi0xTcDKqQXSQFTqEPGmLT
2nN8n8ys4CSoGpdEQflPy3wCIaypRjEKiBn/wS3rfKSwQSYhjouoK1lYXQLoj21XnAOcst3fI1OQ
kcSjNFK8Wwj2MePsJX0UXVXet1rHT2gmjV9h4U+9TASVjV14wZT3KXNKRSM3the2LJO8AGfLSf+G
RFxf+IyAlZOMjZtp2UqD+Ad8L0aBxs+UvtxgOOXPhX+K/EubqUBi+0wVe8DZ/DKe3vEEmFCuzJ+K
f4X3MxIz7UznkCXl3BFIr+fVlFfXHuBIvfiA38PzG9QzrdZS4a+RlgO9q+U816H63+uMlNI98CkL
8hsEJ9TU/NtfGBMeKPnasjwWHtBJyRbabCCvWj+r1cbVdGRtsaV+aJWexxZwJRsZ/mY+Ctts7qU5
S53hDaMmOlaYu6ZAUtYR2dE+IYztSwo1ur3QAI9joZhgc0zjdOMAWHBXrU7K+S5wR1n6G7HO7/jj
GcGF5BuhKJFrBolfXrN0ROrBRAJS1W38SgimcdJgJ5jQrIizKSL6waoIEmTf/gJz6QnMG504D8/J
VReyx6GRW2mRM16QKcCICUnyLB2jGffrSh0htwS1WdAbBffEPAwtW3RgPOUl5wrXCLcyN1uQqTWC
h33SitStLIhKq/p5+axcD+QUTqS549+uJcgf35Ir/WsoFPVsdjVPGyEmytEv/4FTtn1zh0CU7SKO
jPXT6o6NEZMt7E8/itMSJgkPrg6HBCci7dcfX81+L4U0RtgPwBVKSPdxMCs/dbZacFjrfnDU4USX
yNLVFhBS4/IbVknKN2L3Lt1GoP9EW0QP0O5xoT160AnwSGJCFs03gAUlB71EqEBWDJ1dWAkt5zex
oP+NeZVCLAmp7ImK5Na4z4y4DSfR8XPIzntFA28uPqwd7ZBzEtdxJY3ph2sHJMI9DFaVvF+JoAA9
df5+wj4wRcgknBZLC0OZbiiXdgRjFEkCxCVgBdanpGrjjFiPnT0t/ZQVU/2PbXU5jqekzvxN9B49
kOzNiKYlD6XwkimZ529my9rRh/CkDxOt3RiVao7lAETc4itDsiiQelTERWaQXzgCqtl9zxgCwSlb
IbfHL/Y8DZtPL78Aw9qYbU6GwQop9SqAmrXGU49W99EDl6SL1+Rne5E1LkL0GL7vFjp0gKYoIezk
2Mer6VugKbDxvPtFdQJTUKfLOMYDCLnms7q311bI814vR6132dGq3MWaMEiB/D34HcjGwzgUEpOw
MY/dTzQ26DBWBQKqyta3VjSLvV5mb/n3bSUEz6JzTyoepj5BJVGMxVfJsHqv7mR/O9/Yzc1HMcvc
gbcuotAr1eq2baUwgh0kYPfgXt2na+khGCxvsL/ODFbDAUAvyvc6JOUUkbPJq2uU9fQw1sWrCccC
gsk3UqZWBKV73/+7CN5Ip+umILtW35J+8+0BVrF8QnTn1lJBLQG50fiC0wqPJ4vuhr5TfbAKed4O
JX+e9z39PB5vnqWUFFQmUfBDnG/1n1lKus4FFcERfQTrpZs09J1KUD44HTcMXJz7kBCuy3URzXbu
i4fE1Eh3ART+0Lw25eGCmnbEQG4ZKTIl0YfuBlzkX5k5ISSnMdRLC93HLSXbtsdrpUBDjMMAxju8
6JrCTArcffPJe1ruHiLb3nJT1DfLTp+tBLF7F2Ijf7dtdgtkLSMJ8z0wu3qbWiXEx200F1HSmlZJ
iP0IIpqhS3Q9FxVBqQPIuRyP+cbf9V55TqZVA9Gqog6V7n5jdu9vnzRZLg8w1E3PqBXgtIhYm1D/
ysWWQAv/JcQYb++3sZY15g2Q0amf3dN6xBtWgqSDRUBp3t1PYb2XSxfgCDDx836LIANvF/DnpLBr
IXpn3q/Po/SdjX0mAvRPHDTPs1yNeL6O+yryyjkCTUPqk1YBS+0ncCaQhkSQ2YUEpvurLSybPQd0
mChc8dBTAVP//clMGfpRAeCzqYKMn1+JS5wOPjgtlZoZ+aTU+oz6P/RjXOsQjQGjF6/0ooYP9kdo
sgQq/kcFBtW5MXM1pEOqiNx5+QK9DoLSu/FZXc/MOXEgtTVs/F8OelUP1HSUBmWPoh5U2+Y10hAZ
EiTrhw0N3kbFfTGSP4Dk9Gxy0XnS6aO//k8nYY82n4ylra88IWwS5TuiocbAzGa6lvt+tYq4Goip
4Egcg2c+CCsGDNbqpvy9MfQwBT5pg7VOZpoDn8N99CZsQBP5OussuCFCqvZzxaDmYtwPIVtdsKtA
kfzoY/kIT1y7qQN+TaZFqXovxINbef0dH92wW0tMxK1B0YyQRDRUZKXanj6n8t16C4ExZeQ6V8fH
s/jSScBrt/rHC6WI110OGvIWWEdBYiHBMOTVKMlEwG0DX/tiijTE/jZarAGBDvEg5hdpjrhLdva+
oam4CKTA8g6t0Dy5hFWYfSO4uQs/ARUzCQ95BjXNZKh/StXnHY7QZpfKbqwY6elG7zIBmzpXlP/Y
07vjlIst8sb2vvQtGM94OLQYNUCK0WHtEfbdFbc7Sj7cIYYReHcVWyVsEDluNaCOQo9dEQgGsAww
eZ21123wEw4SxtWklW9jTwKLzhxIgCUyPF9Ntx2xDZX2koOle5OOKvs12nP3GbTedLTm29V1P8jq
PA2s5HYlxVXh+DzFaBWOz0/eSRA+gsOAtKo1ye44D6xOOsxL/GTnko1/y1sTXYZ3kxhcNoI/s/X3
pcXKm0vvKcG7Rl98UeUqVnqv/TsXih2SA3G1kj0tTqq9ocLTML0TkzHYGSBgRY+l3zBVR0hl7G3S
w1Hlp5el9KPM51MVsQDJ1xmovo8EgVr4LvNbCTvk5SJn8M4odN5ULoBajaKim3NBIlJQ11LrWKzt
6OpDESdoMDXWWjvudDr5kQHGnfV3cyxDJwJ21NPs6SqaJELcaUOsnyLzutpqEJas8WvCBJhYHCFv
28UuyQohgmoBqzlWCrNg04kGIxNusI05KNc9d3Zsu2+YftXXCtqV9GxDhanFJ0JYss0PNnX2wOYZ
XmPSkahk/5IpdwRqOTP9oYDAy64wS6vl45WcAlbQe8jOedfg26P2H0sNsz5spKxaI2R9Cj6OIQUG
+dHFCtqR+r+9xwrbJCO4MCrwabhzJOyVATkr7BKXZGeE6wljSiEZCfM3eGXJz8ZECCwN8fS4joyl
S7oIsYW1KDdK4pz60AwXBNE7oSAmHjGVsnD15UR4K4bC2GITp+OejMkHxT8IRtW+2D5WKrCvnRC6
+qM8ODlHnmUFXNW8/kGDU7s80k1Sep9OCaa+5c8tqnc4iIa1a2s3QhgbdrTl7rWeO3RaWb9vktvC
Bg1twYIhw04t7afO+rart5KNoXa8Djvl9HscahrE8Y3K4ctgc2XDXGjdJYG5pZeYod83FN0U97YJ
JRRg27aXOUfQshNbxrKItUGdI+jpPUqjbzvvighrqg699l815mTwVxDJv7uOKo/EcOrUApWSs+g7
L6IZmjxFXHqQrkzC1G+MQrDdaJ+Bdsa1phyhTGo8kUVTCZ0cAq+IbuwesHKzphxmKvlnRcjx+ROi
eLQRBhsgc+SG+ECHQb1xGhEnDIxq1BQFEzlfHZBsgSTM50oSbfXcO+PK4W1MKHao1C7QxPMXMkx9
mWRBWa3d86JfXJtoiJgxtcOuo6cLH/Wko3VQEg5qCy9tdRJ2Gi+gBy1UD/u4FNsEjmuQyUsF+Wd1
LkzU/zDbBRI5gUbkV5QZdTsQvkh39bZNXBAuBDiDeC+Zl3ycNSQFNKniDW2aZZYyXchOaKIyTqjh
QdpnFhS9JpKHxToJBQWJ3lZ675aYfkyaMUmnAoNYSKrAqXNlvdlgux0wKvG+MhW+lNtl8Do2GcN1
F+Z54w9s/wZpUuLNzF/2KJbADa0DV4HmYOxVu2zVwwR62BbRaRx7/3wTJfZnoyfwP8ro7k+u++1s
7yCJkEkLw1YCJE+MGa1+0f9zzem2/PXlZLfjrsBZUebSq6NgGejHPklcUt/uPfozZmzSSySsmJsq
p9/yuC1SvQJN48b0adeTZfW0lB5uPKFtORQc8ljE4GmqmJhlDXR3WB4hSnQf/ceXcj9R2NpaoUrr
v+NDvT+o3Dhl9NL93a7Jg5J1XDWokRF20ILjtUNStKJNGtSqSLciejuZHHixENCg/L/E6eFgSysL
O/oTzvxrO3nvGI43AaGDOjBU6QAWbAprJ9VnWicYGB+JogTnNZn7G7goGG/TG0Hv8SZ2b/Es9c3Y
g7dLCmHjhicO19S5bMGizmjCUechQCmTNCcnAJfFa7T/S42c9QTrRGw/nlWfrFs/9tMolc91+l1W
iJzqa4KS1GKajkGnydqLyiSd+DfatfrQN6AloIkF6nCK1uAg/7C5FV6+MwC+gsqJ/wQYmVcbsxzx
btRZfDBcexLe7bg08+YxnKStjY/rHpE8Zrx2yvsUEgBag63Nbpd3jLq/GBpHdUpQ0w3R1JRaP67Y
Dw+Quwn37I6zH/C+70HS2kiK1RoCv0SobN1jFBbKjxAW42jt3NrXZAKzMqWQ3PEjR7Bhu3ti9bNS
mnF8FtQIqtrbRsS6+eUQYWBziwxOZR6DXeZTa5FpHtPMSpQY+CBTdr+2DZuSPKIgoEzOvQa0iDBQ
CuuiBOfLSBbWsc+Cx4nfayHTnn76KvTQTQyYMHyEp3DoOzyebeZqXiXF6mbGzLsu4eVsqIgtyCFL
zXvV8cEgX+NMPPjwqbn/qPdKLbhgxHpZu4ffJwiZIOGLoEFLrS2m+x1K3NYe02D+0khFXxKpKUXd
3uBfXCif12dIxmAz/dRvw8yktqJznlRW0B0yMCNUZOO0wtBkfEk/XCZsjBu3XzEKjkrkWXGBsNnM
lZTT0CbCFBdKv/9jHgusk/Uma97RvsBpSSn1RJKOatHX7VsMyvipiPW5xZLi00sunihB4nUpAKeu
fzcNtWSt7mfFM7sZg/srnex4NVbEhviqQKvmgzpBLJ87DpCAsgnBv5o4wr3WjNlAMFGLB3Bg5NgX
Q2fFi9Ew3BBrqgtG2xiSx2pd/QHdHj4QcfK8SQdOXeUsHsjGGYFYwJ5uzNh2q5U6KzfhhEGQoiZZ
P1rjwKEryvKTr8OdUvxykjKUKggw3XIzNzxKvxXfukges1yAXj5zPMrYJg4Vwkxf/GaB8KIZcWra
w9xvJpEbrJjivIooi1JVDjqwXPzfbDMm9PDGSzuWfDu17/kxEM0L3AWtXtfDVCNAtA+XKIyx9WDu
1IqR3bupa1X9vCGfxOe0cSRAjA3Va24qx7NCZNvZ8KvLlnIm+zqSuyXb0bZkXdTTJUBbJDHmW8Tn
405mNy0TDkmK8aVuIGi1lCyBlatdVA4gRZRKTa2VoDYz4BqEl73WcwQYpfBozaZTbBpqFwDDUcE2
nVv3YgJMDYXgSOL0jfZnQ1taHV6H75e93FtUj4nlSW7bGx+07LuO9e22b4uDswZMRqopdn9LfD8j
0d/Wutv5MtwOKdl7dHUCNnMQHrUFmqi3NrroPao9QVcDDfrCwDAWXDuXgDvkHuS8MqD3MRuLtkR+
/TG20M9vZUlqZsa8+q7v5tWFT1W3bM2XCXSne2bzIlQT/DxtADiVGxPAgfamwbz6NfEUJIJ0Bvv6
yFYVm41dj54UJ75tB3G2ADVxzInNZFhDui5Vr1TEUV2uBszIcHKtSzIgkevZdcId9beHMcId0O4N
mKpiLCGUJIEjdPOyKvBLdhg1s77gRFlFnAZkO+Zhdb++P61snmAsb//GF4E7xb1M89o9w90vede3
gf2yYk8a0wmUTzFHHU5VnBZyAns0LdDMkN6CjyPm0K0YGRW+iYIXe2u29CGGnGnNTK39dGqNZBm1
aHEvyoRGfOUlFImM0C3R5Oq+Gr8Omrur1Bpmxi6BKaxShRghJDqbllgM8AspRY+Ad6OPkTlaGPJI
k+fByhN+awzrgUlPGdvDSRrUF98rafvTgIyNqii5QlMmjtMy6N4SDe21ir/7gfL3UwaSNle5rfkd
qsPD/TX0kMZwwrSLw1WZwxmBSDyu9COvqlnlrqw9BzOOrW31+2/gzgDbMvB8+GmTHM1qt1scx9da
ARfFOHIe/qM4BZNnDXhXipdC+xVL1eCILA/t8nmwY79mL5xoo7GsbBFmkwqtY6uMZOo1Svn8Lvl2
p8fQv2qk6/v5PZwZT3PROdW/TkuWrTFRCcpiOrpegHzBBiHEGD9kKzEme1+//FphB55siV+6A/Gc
n2mpAG36B89CSr6J9UsuYlC4oMjbGQ/kZw8Oe32zyGt+gU4gK+iWRc4SZ608oE5cj2ciroS5EudQ
2EXKWNc/JlRfmXy9Wsf58Un2l9XIXt9aEZ3PoJonCJpdxG4XAD77X5hv67NYc/+Ylh6DSAAfOfCz
x8BVw3rU6e62bmjeYqhAaM14jWlhQq8EuBGGDcqPs9v2z8F8/CCdb3JBLzbydcE67Z/qtvLpsBxV
6vv3+zfffy9gnn+VI4EfpAxYsds1mxyuqNYPkFXOhbPjIA89r4g6oJoHHj60iS1HnSHTOBoYYzrG
TAF1Uom+dIW5vBDX6Pp4AEYR7Qm5O0jrFIIr0YoYmoYTcm4m0bdMgOOQ0WhIT/tqI7ANnKKwRNvA
OxM+qaaRI6SDqrXyhbxpHpMjygXZfKrKRBSOoPYECpVEitvSS6MvpOwbczElsIp1bNpVylReyUXj
vx4LhU6U8SESqHoOAD66e7FU8a/aabA1eJVpXnwRZOxYVCH2odFCtma7qULFMoBWNziGB6CI2AuM
+/cb5shqayr3bcGf6rK1Gkl6s5Zf52rdaCLsr8r6xKK7QLaGIwNmrZLlT8rQXRQrnSkBFPVhMGMz
UNa8ksxPzfmwnS5qJfc2+dBUYjaZsra7GFtHKv+4c7QkiLSTXyJHa2zZiZADwzgGP+3o/U6V2Q/v
E9QUDYnVMOI5XxuFCKzfRXMg4+8nraSJpcZnuV0Ak6BWL9oiVRMqlrb6y2ULfthE6EKygCP2zB1j
XtbhZsxZTNq+2yk1w6uWFNA1FN8MG+CP2Uqp4m5QZ+WDYhFXW17ZUXhHuN4jenTN10q8V+aiyhhn
Z0PAKflk9zMUY1Y2H9eJvqtcFGomeWCrR3tHHNMv7L/cwX5/Gbu/BhzPh2d99J9K+rEFvb4VmwFg
YUP0X7IzCOmPEmRgHBqsShzJ3mw6fMagQfmuH84u1mbmq9iJRONcNQStN+DuHkaV3CzN9rphV12s
o47p7GznnpS/GlbQw53jrW9ye/33A788kjTU75GeKlOEQV+1ikhUn1iy3i2jWB2pS9tpHhJ/uK3Z
g0NBsdwFCxHvXoOwoyzQ/8eMBYj+OiDN/cdfZSt92BaBmwJdlZGeSt0/TCG/7rp5jLX3/9fC2vBs
Vj9wyZf1PQGOtms+HsWQpcMGE+nBqHq0ab61kKUVxWPxWUo4983GaN5OAh6zwIuPOSZV5BxcEtMh
ezgEn750fcOsekObeKayP5KJhECxvEPbrG25mQrCFQ/6YGDV4Rwbb1pjvURFEyS1gWpbKJ8m27Q4
Fv5UnxPnO3Rjel4abBG+aPET5XKSnbRi60IhLh2MZ1A17WT22iBQKmiTVE9X/OW/N5b0EbnyrALr
U/zvK0U1yudDi+rfgLvh8JcuQJeNB49Ho2A2sOxGXmgibDO7SKMSfSBrpkTOB6AiNz53XfZucZ8Y
1KdmMb4kMQtAb7HAwLyrPlMUzTRy+he2YCYLtuhD/xgqNRe6yC7R2V9bnL+k6QXBjvyOVN7/MVpy
cizfL0SFBGyJoTbG8mWk4LCbfVI92uoITLC7WL5Q92WduMwA4SvfqtWTPpXECgIsQJYVqij4FteX
Aqs958maXR39hyDI0i5OLujxtDFMy99EfnZNdnRqtEj0LZ8vzxHnCufOXaIpTy3axY74oMH7jifJ
wQF0VCAFZCXtdeDJ4soywgNti3mvszJUIP/KCn2XuP9y7U9CStSshBymixV70LpgICLWsAlLKJrS
Xc+oFebh2c6tUFLhe2LQBdzZWCV/25vJp9o9L9ZaCMzkHowMiIGVNJlOQGBt77ayeueTzjQoX/KY
5eAFHiE7lN+4mVXvlxGlYE6RM6KYpRuG3REVud4wmyVx2csG4z80IGHvB+jz8bAuekiOD3ah4ctl
SbJIvyppo3ogoD/Rlm0Y1KmOWh2w2b6f3EDTtlef0wwfXowYN86AdMhb1F9AmOu3BcbhlxlWfZro
2sk0o6IcR0eACV71ppcRZKHsG9D7bbmuwrI9lvp7iXGVXQP14x96eQ4K5/BNz/QfKawa07JpgR2S
bdlutCG7xhdwwFKjpGzD4ibhwhHFFCjRKFmQtd2tX8T9m9E0b89PXSrxSCm2nYVQFl7a5cISPXh3
qGVYxvoksxvxiT6HHd/Uv6YqAscdR/31r/VVpvBogLzjzfLuY0L5w8wYe1+Q0czAFw1EyN4v6LyD
mFRLpC6eV+fgeGUctIuE0YnSfF3aImBre6jrnFhwKl2VgVuP1uPTxP/W2fUOwn5oa3maY7RLQ1+P
Cs0MaxaQVNDtbWZCRJx4atus+WBokoD9sHQV0+zVpx/ZHWUU0e9T295p6a1MezXSlGR3BWMlXAG+
2LCgrQGStt2CLGZLADObBX4wEah3r9t91ZESL6RQccextsE1YugLBCbzofpjHimbeYxFAXIKV4p6
zLBgvHQFYjnlZCJHVzJc+CtTe7RXGmEDFaA8FLQQ5zt2YvwsxyR0/V9qirAwrc3W6BTSVRik2++g
FKQTtl9QzH874yknAx05VzCVBgTuYXfV0y35qmNx5rXMxNXLR7GKGtLxVL7smAf500Bam8gnCr16
PWhBAusGdIrZnnQh0eDgNE3PP474rZzU1WSx+Arh2+uQiuRrYYzwRbyiD8QdginKRkutUd1Tnx4h
e1C26fUXu1Bvn9UOYrP+WxFB4PQhIt3EoNAt+Kz6obVPa4WPrDf8XIqGy1qEhIzYeL4MvTjSBa2s
5gDTLgzoVkHCgbyPbUIlIDLPLN9y5SxbAaTelMjtlJUcTunSFw/ZzbmFS/T1wboBkC7rR/q5gPYv
q1vwXmW7/E5qfRkc/yBuXvzJRz64Bw9eeRSI8BQGZs8lNxw1+joyoaps9wk/M7gVVxaOCCsf2qrP
vyK9eFhiNzOFDKfYzEcWh2mdrxnavgxESaPGujlgp4eImQWBsjhx88EyTxeN/O3eedfJ7utv6hds
z00kj2K8K88Lw1FpfAzzlF0CnLx1Hm3oI+plommMj41dWfL0UoL6wx0BQi6mKwprcATDgmulAiLR
6ruN3FuSFQivJUpgCMGnJESIRp7p4Jz+xHUrAgaajC1Tf4n9dTn1BaKPn7AX/zZqByy3Vv5T0crq
H0ZU3WVWA0qlQoMdGB5q4N0MD8TlfZ75gqs6qHTET/xTRjAqfjugn517fa+0F/G2y+IIox4cpK0h
wA3CAzjo5/CpUotNuHKIC/6nETmKVbApQVlRa9IhDdoBdk8mB3HCJ2p28mwV17Q3vV9vol/1KslT
ur4Nua5hrLyraeaLYmhXKmUpA9zHjtkqTk9L/DSuvZS/b6gp9rmchHz5gOyepKaguY6mIDz7uFFB
feRL/pvixqcKMZ79J+XYYjTAFia6MIxAQ8ReDStWdJhGVxyXhhFE023sqn7Prinew/twyKCmpQOX
0et6qCeUSOvru6OIOu+W1ugPRUd/6cSktMihcThBDVo9VTMwPa+glIO1WueYFqHfwWJbbI5Yiype
Ym7pT0/PNyMlGnQr16rLq6VDJwCPIlzDnS2J5btDQK0nksk5dJpUp/kErZoERNXrjPn8yjSxJ/jM
kieE29gIG/3fNMCeX57qL5Lm7/fzYXJWKnd7SXgv+lni3+Mz+ttT5vhpLXMSc/SG7Wr3YAGAX+kO
Rv65hrbwjAbWkLNUNh/x8Ax7hgzWPT+yki6x6FemZ86XqXl/P6aSVr0kQpfF8AOlbBQIBY5tRLX0
cVM3EdljkmD7LHfytJ94Z9TRCjBBM+nHOKiRz/pq1yU2V08kdaSltmj/V5N1NokvRnb1h9Drno0j
qWq6bhb235C3zlSwKwSgLD+c9KKVYOKkLJ43BZqNyNCGQBbTn+QO44kqhwSx5gH59wjDEYWmWIj7
sr7B03/Q1XDEt1eRRYoikbjx/Ha8Fr0l+x8/zmL0ewCA+c9mP0xJxtgBRcyG8vxt6Ly+sv7lHy3p
yDxm519Lt5JSb+8ADdXjYRj8UvdkcMzzJomFd9P4jyJ6l9+vro2TYI+b8exn18pOaG6PZHUfC06/
mR66aZdWwNmdLEaKUhoDxZPWbsRUnu3FlgNPJILmJydAtHKar6o7QrCyrAgpdg4ajs/MMc9Rn/ja
Eqmg5nS0YImvKPspLEkrENAgXAPnMJODWzFh3ZBm/uTQJF0KLCkJ2N2e1hfr/qRopCCCSXG6Vmsy
7jSwn9Obf2VMDblH+r2deQOSH3t3z2rML/8UuQGiBV3FPdyUwxaa+L4CYL5Af4gPU7CvOIFYxBT/
0ia1IbCPt0tfYhiweNTtDq1nga57/RHHom7AdKFRcw5f2dzoQHMSiXgjHBWqkKYNPDJ8OxCbEKZp
MdQvr9s2KTIVF4MJ9ReK4bqyEFyYCzpA21+OZU2ZROKJxB9M+Pz4e0WGwqfh1IwFJpr9M38iHFHL
q6Pc1ewWp7Ab+L6g/P8c2oqK4bGrG6kSpymnK+uy4ozC78rZmkTzyFIhXz5ebMTTZvrJ1SRo1aVt
R8AeczQ38gkApYcVXcSOFUHyhJ5F6GK+cIBd5DWOpSypF4iEVK91RD+tl6oIwAJVyiIbvwiFMYVS
72EEFLWLW7XPWqK5fvUFHAsGuWse7b2M2TsoNQtUT9XiG1epb2G9iuLshBlOesZYh6O2i8SE4s8H
gaVX5NmqdnPnV51Wr+PSCixSgSP/xQaA3VbuAi2ZiKwmy6WREm5q0J5qtEIeDt5R/tIA3WuBAJzj
t9HqUaJTZ3Et2u6ZF5K8Rym6JNDLxZ4nKLoL6VSU9SyFN7U/wdkKJ+2QGcmy/nRL2Q9qXLtOJuK+
NIKSVgxPrggM7Dso6g42A8huaDckCHMM4SGYGaCarwU1ARGPcjQcPGl+Bye8h3eE3qyodNUShBVi
P1y65qzBcZEheTsXbHZJWBimUuTcUZaWNW/OC4c82QSqDhdbvR4B+8DIUAG/UIT8+gzfsRAohJR3
HiPRSHEOBV+PMImJsrQ9GT/DKs2Px4GQthgOV3iGBIhYa/mBAdJ7IVHHuAnHaoTcGzGM0si9StkC
i65qBVj+6cQkIMRQTpUDCUQYFKfT3bfNHXcJ6ZrcS90Zdk6o7gkeE5BtmHnnrPYRgPOSH/JIFjqr
mwHpyZwSNbtrB3GtgLk2TuSS3wLU1ARZh2/2l0uwVnbPNZn8HN23qMM+jscYn2quTOW8UbGQG9Xk
of5tjGoIUx8VRnzdu0Wb0VHRa37Z/8+J7aes3MRfX6MosRoPaobCgF+P8oMWGD5ULS7dVbQPCSYo
/UpEIeWMNvs87hNRYq4mDlztdDIHBwQ5CDTY6vPFogZVXmWXR+1QlG/3Jx/8hWEXVdpL115DZhkV
MH2YXgvhhsIJIsytjQHq8FYHwbuj1TXQRXdOeSOAlkCqhL8elBNaOUHRDbA+nBYVsLaFRA9k/sH3
bpv+KEKAx5XYl2qvHAQ/NP3U0D3LBbkg9dhOjhpRqAw1qyhKfRFXR0ez/cSef+ICFTcnpdxXBfw4
1PvEueZZhHz/+Nf7reoh6p+kk2g87TUVXpwjz9MiyrW403EvG648wrw6k55+dJ+//Xx9fbA97F+5
elCJeAZmQ3AZADe8bLeKGA6X3je8yN0io5cYep+lkUhCr4MNd4BhAzPAGxjIOAF9erx9nbfot9yZ
lBWUUS66XwpIqOwGxjNnwJLw8MSfCZjcJHbaeamIyQKVHWvtduXutPMDFygjFZnPFHUK4uz4HzH2
gAYnTRubP9IhAV+6a6khfDOZTVR1QT1LCjuzF/deolgvZIbEHzq8j+GdIpKiZBnoQkYKAVpWxFte
ri+dSVU+4y/Fr41Xoh860YCnNxnav64Z2wTATqLRfVR93M2Rctp7kSsiJKBdPogclXMJNobAYtn8
8gAQofIHPixIHnOVg6EK/9r5v1wFn/3V6BBtOQ0Zgay/UwGmfk4xGm1eifxs3u8FNfAvD+lPV8d8
tBH+PSZMxSJs64iNWq6oWwk7exkGFxIUEmGp7dH8oeQ4BP4n7Ge6ZhRxNFprHiXXDIqVApYqTNd8
apFCkMnepK49SBGg5FUt/7/2rfX/64Y7LY3bydZHpt7XzLVl3mjows/ynGb/FzzPjIV8IKDdrLbz
DwWKVqz4nCjmnasUx3ER3/zO+asVxFnbdo3wuwLgBK9ECG2Cq/1W0ADtPfMcGJJlywQ6hMC91qkp
WwRoLWE4jJhnyMPR1fUcwPyFXaExjXQUj/eDbrelLmWioGrFs4YtSQYcmmABW8g0h5O8SO+I5rnG
sUiIThSTop8W6L+niQip/UM/Qr8y7hKFk4mBQ9yeoD1ouhwOeXZHVDRwWlj+MXTJB1CKRuQQf8GU
UhRHL0AyqNYRssmyjc215WPhL0CIrHzY9gzOXdWstl0X0yD/tDWDbBH2I9P16PT+XcuJ/v64vw2K
oaZQm20bcrfrbVo6Fda8JtepKLHKmw2KzhDEemC3WoFM52zdWqMlKaubaoXV6xm4qQlmM8otdLEt
zkv2ZJQUx6AjtZPnjZvgbpvut4LAMmZSMmnOJL0uEpoev976rlcGUys2EsWJT7iGnWu3cAcPCKaJ
XDsX3bZyeVuDt+9yea6duhL6ayvt3ZImtXjEThZYQQP9zDnZFXw5RLGYpHYex6vlMfDkOVy3llVe
wh+DHvWfMJsXHMmUb+MdIZsJ1OBFJofIDrp7w/ZOXOBv/VHF9E62XNznXgnGn5hnhCDnyG64zrs1
tK9FH53l9i1lbFTSTip7/rNT2BSO6NGnwJ6pFDFmHJy6PZMyR8jGamjnUYQW2kcddoGtgXyvctZ2
Ert2atALNUsMaMzdRUFZWl0pjm4ZgfMzTxZulI8tIM+Z5EGTGcViqnPHPOLltLvaT5R9z5FC4aIL
DVN3RgrITnrh3dQSsN1HBWFB/imkOIOmYICdLPJk4fD1XiDPXdVirF0YTVBklTrb4agDSe0RwqdD
+L75R+8L3awa1OXWv1NafJHcUOJJD+FhsRYT0/Crx2oJdxe2IJ8M7eTS0Whu9yRqOOYvs3pvoQFq
tqrFnSvzhsIWP5c3lqmRzLawyeA9w/moIY1CkXkvSAVQPBlTcSEeAUPRVlesAK/88IhVWTtUCbsF
Hq2vi9urGssM8TSEg0bSUo0od6OWufrILFpSqLk2KzCgYUZyVElB4s0LTNFnjMygb3TBue7wW7s7
exYhSNaIPE1We/YJpyVNXTQwloUxCQ2jKkCu3e+sxqUN4IDXi6bQNEANQQxnPpycKd9EqOQp15Rm
8h945r/YVj3bUU0df2v/67jOYw5C8cxq9zw9YEJ7+1WA4mDDk+AxhqYB1i1aEh3YznNTOKQ5s7Yc
6kKNsQbWtrLG5Ak3uq2ogJSP9hWUbFsCVL0pQX0+++T3QoUPCqJGYrJW6+FI2Rrkl3hC+8IwlPF5
jcO/yE124Byp+V8kGCbwiltbzro0sxXtXweCaQ3DmUELsAIbVlNfmomBHTltECa5HkPuNyoiEWAy
BK97C+6aHXJTCdrZVxWDLnZpHb1WsgwCH3pWMTa5QNF4JfX5nGUUmcu2BQnVYfN7luaVkYejFbsg
GisffwFz2ACcCuo9rPEiu7ERu2KhyQ2UUE2+hPgRH+FCEPpxYNsc6riGKUZoqK3X+NH7xKa0U/Rr
WCBUFbYfM/lgK8KGCIUsnWe3X7W+3b8n5u6qy59axPnZk+a2scLg9ZlOUkU7wYl4msyV2OEFYtR2
Fa9F6akXtP3bzwftTClWrolAJjwLd29kwqp50qdz7wtnLf4Le4Sr8WyXYO234Uo1Gd/R55QhQtkE
6dx2rOycPeevSrDFYrN7DzuRgfvWl5kNCjsl3ZovbjPMfz4bvWWLGJbssaXNH4OMLiiOMuQpobqc
sPXYgkhCCzF2o69g1S4Yyy1AKa56+7xGS9nRqy0n3aBTTcY74Ijzqez6VHmfDl+HF/LZ4lS4zjhO
Jvl3y4RGOa1H5x4yAxIkXZFK0K8D0kBTsqe6D9DQU1mGTmCi6xSnBjf4Rv+FanEZFf9otYkia0Op
KSIOUThv9DTqKmYEbSky/yGrzbuTjqCSDR/WvxgBnCH9sqg1HXp9TXoRiDR53qgD2lp3Zs5RVDw2
M7Dw488mtOtDXAaN7yq7tVlOzfGysl3aIZUB+ULMXUI9+3A9FCaIFqkRqGupPK9amxujlrX5QcYo
6kFAEzqGavHK6UUWhDUAqR9EKKxtIkDWdE1orn2ECg1/3gy70lLeyKRPwd0Bl9GlMSLszB5AtVZ0
MxzSQdQjNJsbYznb3uH+99igNSL02NT/TBxCyLi6ytYIGRISGN1e148FuEl9O5Cgthaz6Ze9eDgN
P54T+1t246InmWhQBuAqLnmx/YTvJxKZaj6I9TQX4Py9rWiKi1IZEXJJ7UPQ7v876H75qTcatjEq
2j0Sv+naeCLGviAG0zKpcexxdo9yrBWDIuh/kMEfYdq+Yir01jf0M91xvBBRuRPEF4vU1GmGvLtb
v46uBLMLbvjZQVoWpSKw+pTS+WXPO1etcmvOb3i0NbC8rYQXf3l93PxkKyCpFgFlIybJRjaOdrwy
xKgjXauEe8tDxTFcGGcZ9jBTB6DHx1yVFjgF9WOeUvVea9V3dXlnvOI+3pgqaFCuG41p7GVNxYSL
m/Xq5Nw0j7Xo5SKITO0U0sqa5FFWufHIbLoiDrosrq7APACiGB2ibr1tUuaULd/g7a2Iiry/mWWK
a/0WexuGy50gXxUms2I29NhVGJV4zUidcDUkDB6A/PMFf4tPNe/CLEf2M+QqdKiOSlLytEvRXgmo
vcux82dsVcCHhnHrYTuRZv1O0l3Q0jH3XmGRTI/I6U1cTuBms8bLIRXqBvCy0wnsC2c/WASh9TX2
e+26t5w9gN4QmQnDfu6pY5Mcfv+LOjiTYcliAScFrTXoFw41nOmyr1ICTPZxUotRsiVsIb6z0r9q
RZ1hbNwNWk1m3deKTGlTqAORXAO9WQCgRtVTifXVfWrb2vIYWf7xR1/H97HVk7enwsYbIkZ3uah1
ANagFbYBspdk6YWDPzpeUmIEt60YjI7xDd5gxAC0RVlxEErcXpwuKMHVLDFf6zd7v8j99PwR5ZUf
MjfSgEENexITQik2S0MzbZxJ4g2bfwFrZME+6+WdTvfa73AAuX+M2s2P8/dz8JDvN5Xtg8zw/YQ8
3Rx4E9j0CKFxM0dx7a5EDHIJFY+Wk4yFRQgIK3G83W20+C1avqih4P3Fk9Rg3s2Myz6/hD0KQKop
FoS0yUMw43FWclhmQ9+Lrm29hc1XJgoiE9JTabfKzmCw4iAXFQrI8VB4j5zdq1DWMqLxpdJU0hkj
4yTjesE53MU4UX8KltDbkoBk2V+w37tCQxVLx/Ed9vBNLy556aa+baTSlxK9U/hika1yK35iMrXU
6r1zynJbg6/rNLrxhG3Nj6YL03iS3Ib/kdaLYSVOAiBh3nqF4r9M6IPah3gQSjKAtpg+IRuvu18a
w9VyqDX82LnTTo+JCoYNisd1xRFzRS6SbD2gujYBPrv1y3f82UwUbGPWkComiWUNVDTUT7sHbucv
SUFRp8IcuNxJygYBZvTbwvohCuNjlIiO3DeS/lNKm/UtQZCkY6jKZqkN6Mu5TkcpHTY3OeYNaztR
VmxJgLCbwjoJZ4bEUuJiNm8XBtArL8LgDMzjpVKpCERRkFPnFEuSJE/P0mxnjBlAB7pznlAjpxy/
Q/ZUsKRTrgxRbYJwZzDgx5TSNFAaep/j237wFnJWyS9Iuxxz3S//BCZJvsDxKw63DlxJ+8q6jeqK
y4QknJS6Jsu23UA8Oho472YSXdvOZkC1hslNd5lkmPxen58k0zDAFn/XAbQSB1vOoUdFGSttiVSE
dFVRosrkZyeLh4hzmJ8zU/VIayeV4W3LdEV2FealHaOu4DnFnOKn5YLzVpouiCAL+VOj42UJpQ8+
EqDZQVxgPB0y9liXPySg8sE9aZW4TafJN+T4M8carto1WsLDE72tcPcRIdtlzYWrNSyaEtPmFRf0
+lNnC0G4nMCzSCmdqtDlreZdLQNaAiirxak4VyeLtAbk47jGq8txpq/G/ltcaSZe/ZeOzSXGHOb4
uERzsv9kqWUpRi9VDkwgHHXcfa0GetPjvvackBLOWWVNk50RNb1zz/0kAOgWPEnaJiXLxUDHelej
lGalBs98igOiM/g2WvTXvYJIABxbDmeJ488crGDkabdDewVAzSTttChCrkFnqi8BJ5FfgG4B9OXb
JjvcvmM1q4Co+KVQtBVer0RVoO6rls1ddx3oOKFOd05WuhdoLjSykMGGzeRbMWeApmLRXkwTmKVJ
iosNQEftASJiMd2jpR5S0UGgehUoWeFRbV9cgeOnZ2ifE8pG5z/qhhJTVr57hANYpj/4HAap+CdD
RHW2j4FNhKne9Q6DUWclJ0DN7KK6pgSE68Klwl0NEJNJWAdWdY7pejh+eawF/7+fNTpKLvfekVge
exqnChAcgcM+7RVeO/sWaYf1TAedux09EHZrhiQFMZPphRT3D3BLkKjDhIlM811Bvds9x9NSg7xN
zn1sTJQRZHaEZIhkunX6bmyEE1qiW0a1jkS7tmghcAF2lwdhj3hjlM9XStzJZU3XYYAwi4n0fMfu
lxR1Xga2YiV7F0UjKniASFPeyiv+D+JGTG51n4EgDhXGsLKEEpGer8nu0YMvZwzm+zWQQl8oJRii
6EapbfftU2smwNp6x6x7OPgkY3HkIPZS35d0rsTpdwFoqdH9eIUik0o2bPUtR0GCCfJuaMD7UNz9
cMiPkLOAUMy0bf8IbmH7w5+gIFwf7bE8LcPelk0R3xPL70ihvyznCOr4d5+Rd34XZ1pCWv3e4WJA
/0XzFc0VJn+ysgG82Mg7qwNc8H00aNGxAoVOiFyYhCBlXLziJwHNWNPwpB7vdqUM6ZCpb/5ep+VM
pot+uv00h+hit5vZuBleFRnY6H0KtRAGyF+ABqZCY5O/AB5/aGYb5TnsEqu8PhDBLctVuCFjThX4
Cxmj8+pGDfyDKPnUEIIlTrhbih5IWGLfF72wXgNV1p5ZLIdevYcrt1B/vjcNMMsHmSPS2nbsob8z
RxiH6TiND0naF34kZ2jsPLsQfHVK0gs4jwbBw7g+Y81aIrtfa22IM5hWIFgU9i5IxJw4VM00FhvP
XAfB3sdKmWVoGxe4/gputCAWjlQF0BXTImNZezy2jO28gaT3XP45dO60vSFLtB9H/6OEzTf7U/wK
Suoh7CoH1Jbq06LIS7VvjM2abyLUCdhlTJhvi/PANhMPkG7YtT/Ykqavhopk1zRDlRCn24MI7PfL
efIV8ihN0+HKiklsKfzpoF+0/Tpwlqd2jo+4Vt93UKnF5E2llddyfVZY38Dz4oZy24hyCpOLf+Vq
0UVc6r7iZGB6Dpu/94zs3b8pFx/0d+HqrVYuM1DUTCLTRJFRDa+wOoDArhLcufEDCjng1v3Dmfl/
ZOFGjij1AW+PgXrpDzT8gBbNRMpj52geyrTd6Tqg8lpcoOv5tMGEzHzc/QTHQpR4Q7Y9bQLreeKn
5FOE5JLMZMachxkaewwvpNxbA+f0FwphPwIcvvuzbU2mHC9J6BlZJ814L/EIEsCKXoO1I5GHiuWC
NbyO8PgCUJ43XXf5o00vEcVSTkkD7ezCpD9eFpEtBfgp/hKQ+MIgYFfCOdYN+ucmAFUnuaO2OdiO
VyETu53Ke95yo/P+Eotzv6QVnwa0m/Gh/Uz0GTxxD1DuEjOGD34xWZhGhPXT1/00AuiYFwRVPsui
To8LbhgdZgL3ySEFLVY5SqIsunvs0AZE40ejDo0nBh1i6pgRh/yc6hgYYo/TQvOgN3vqxydDl1GT
I92i7oQTyTqZBHyUlaiaBtsLAZ5N6VnDfpDTyC36IfMFC6Op9Sou/hDRgdHxO95ilWK6x/7Ub5rX
sN/pNG8giS5/TFXJ4Unp77eWvzY2Nzsrzx5k2hVBHnIiY6c/0zc2mf4D8a3RC0Tedh1kQbp/WwRN
PIefLD+jNC/JdFNHkr0ajUHhP1SEsQWpNKADZjoiDKLcGw5hQ+511b0RH3ejwkw7zR9lqyT6x46n
BxXSuwQ027ZvkrQFKzCAgTLbpTXFHA1SonUsDTtPfUhy9BWMKVFX2VwmqdPulryIowWDlF4gLlqN
9z5ddTI+0iBsce1a8kxKD44I8GofBJFTk5LgrjzfnckJsroHxpHsIn+DmCDtuAQmHaGj15pvpcvr
U8nqadwW4VqJ0YUyb8nj4ZvWTw4i4zbU6eNgkg49OTrlqlrPzbFASDAQgPaQ3z90s553+1I2O78b
S2pO58sCU/dxzDK711Ewo5+Vgto8eyDPaIv9JZkTQKknFpDAYEm7lX1HCANhHJHRyoXlm2LZTWV5
tJXAFdbzhFIIRSC7aFLA/TgyrVk9PL4TRMwMFcJ1OTx/tdnV92m+JTDZujkRXstb5dc94xi2+Frd
TnKwZ41regWsFFrRxVfiCADoMo3ndrTOaE8G89z/asVIhNa8xKCBZW8sIxaZgDAYKbz8eTjdv85G
rWPYRyvvgNm5qxgfMgFtsW7o6PiUtQesmnGXEhCW3PhYPoG5ZvuAugEBvtI6IcVYXoLxs2lc38bn
iePDFfFhkuvz8QTyl+SQArZRVKGcb5B9oHFJxYQrGSIx3CC8azxDXqs0ORY11IjcWkXSqEViQffc
FXK+opRzQxwfN2B4WYT5cIo9GO4cn+uAzLvj9/WbMs7wlj81Un26kccbZXUWn6eWUzoNrlNltqXe
wc6Ea7IXtRNbmYUpiByMJ2Aa4h5dfvw1otEVagvXzpODoNi5tHZavJ4wSBiBGn7KF5qEiRc1YJ+h
Y83rv6ZVjuOR39yy1QP+VygAAvsbuOANxSKW0FCBffiZ5umL7LM5T+46vJrrfMjHdR4SjY0DbiZ1
R6fnfE2RF4BPqiFgD37a7+J8f9H/m+mdtkb+uuE80BQ1ev3D9IaTRFNJSBisjOrOZG7sWQmvMxHW
eB3Nd5eQXyzzEeWgOVJdpFH577XskI22RfUY46jXQQP0lDMmwwJgUESPZ4Sgtb89M9Ni42az9pMR
8nMrvsVYt33FbOSJ8Qd8z84pc/Oc9mJ7Zap79g0TQ+i3wWfuAJ2r4HJhFhToBuVNA81u6AlYYvh/
NAwnaClcV8puv8/TY28pmebfxVlBSJ/WaaLfhH/7GPGMhlYkpwtRjmtGzeHgaiNgzom+N+q093SG
EndlA+sOkYsUgAK0Y5tmdFPUVlPMC2BnZwY7aI0zJmKYuQM439+KoldaOqVAxqILhlFEb16MB7Lc
1qcEnoinye4nq25bT/8YpY75UdH44kpC7FXAFbNRsjIdxeFMXRCrMg5bRUSgS8H2BEfDI82q+2aa
tZnRm/c7dZ/FN9OfkzC9Rhw2qXRuUG30ps7o6CZEt9XHQfNjhkSNKgxY4CdVg1+S9hiHXpLSPD2A
4g4QCvzuUQ74C3oXNMpzrRp8s3QmFaU6pzghj8UEX1EdhH39sj0LS3s4u4zsQS4figIvk9rBHt2N
Yf8ljph+FPXBwa9oGi7XN0eGZZNtUENx7UkZAzy0HIgIrzShmLJlwkaW6Twm+ZP/lzxzy7wdaqwo
S1C1DGUALBt4+7z6Sc49QD31V93ztZ2VqOxJUY4sjOayzfT6RDpmxlg4wuHfd2l4baq75fb8Ln9w
Apwnd6OzTD5dsKcm7jz7wnFS9/kjfrIRzrqkNioGIUAt/2fzvJIOVQbYba/Eil+xM7kzgessOqQK
B6P5kO6IiQrZrWRONTYyok4K4VOvhZIzKw1o86axe/5k0SOmp0avhX5OMTTU2bOcC99YoH19wlyB
GzKUd0aDbmuPIUBhMn7XCeefyHx1tu/JepakDSLLkEKlpZb4E2Xm7PxaqpQ+sMjz/K0PEL1oKKX7
uykqeQbQkGK/n9GSi8lbATmJ+7TU9JhFVqgq8sGcdQ2TnQo1sRHY0be+KIYm3s4QNisSt4l7X5e5
2NaLfWeTgPCJBSIfiPkyKGDLy2Xup1f8P1T4O/dQ93kMytpVakUhA+v4qy9LCmjGcCgsKMyfSO+b
Ix+53ok6NxcgQ0bY9yasqwWV6KjsF24/Ln+E8KeIDCTSiSbVUmCTFrIxlIgYN1l7J2n/dh6REgIH
bxGr0N/gwi8SNE+/p7YyEg+O6fzfTTn+sXh2wbv4iiyTVQv+K+D1sOTCHH4fE1Bhq94CL4g1jRqT
aPJJoV97r4KjANv2XmNMAfYgQIzpLdl2NMqLBBG4gAa6Txyh6SInThjf9O+O9oTmtf0+tJ8TIEso
5xF2zFvE510UqOHp/UllV/XsRJHPUWtzU3oCDFX+9RQ9j/EpR4xjfXXOYw4qR8dXfx7XYlA3ybB9
h8O3NZ8J6sTToLdEqbZa8ytnSBgpSqWTbMsaWrCC/qtPWAaruJbwp4IAK8Llm8Jc3jRCMKoZwJ/p
0/BBU1TnYgvpPyFj4bQAuRKN7QxqYKvViKoDuI48gCXNtVj8ne4lSW546qlO1faK6Sxhi58Uwz5f
WfW/xT91V+PtIU2GESTk4DCkNXIT6ChU/OFwnTL81f7iRzG6tVSK2HYIg1a9Uxg9e62+tQddIwap
tPsWllBPWjXeLphjjHjv98KJrsnK0LvY1eDLf6kvi2JqHOL/tde3W4cHWZ1Mm8avrZ1SIvhfmlrW
xYyOmrs52q/XwTO0vQPtuj3DSbBrIpGxzbbr+C5oAE14tJMIaZjmpefwd6IurqwOxRofxUF0ui5x
tMoLmcxNqOrnvi7ceGiFdHPx3UIaV084VimJHnugqiTpudmYhw57uZsSjFCP1cHX7Ucd6nlXwetv
BLYOhfVR+eo0V9Yo3tEMGtsUzK8mV0Qg6pMzyTi8kvT52m7Z5Uu/Wi4GOkYcwfuXx5tykugFy1Wm
acjrOJJ0FgzaXwXyDTQchFzcSf/TZaYYLeJJHEi4xYvMB7+18Thq/zMcD3pPnhiaGkdwmtY70hVP
/aRJ5IsrrRyRwF0ZcmB1waLHmG4Iy4j1JUFYFIf4Gpc7nQZctGC5Q81mvY8HPIesSgPcISdAN911
zTV0ulX9iTgMOd7Pen1WJGz6fAo9bVknTpjEusVB+QSkY4/Iaa6t8MSKjJ1Id7Vcx4EDcSqyB6PT
b1AxIE9OfDW3fP8/jRscgHKQtT7FE2Ehci8jyEnSpju9bqscvKGrXZhiy3OH0dgu4Tid9a+p5eVd
X0ai5xk0m+T+iDFIZl19YCNKuMmN7bS1097TR8KR3LOB8kQI15zR2o531G0dEEtGnLnP1yNYjI4B
BeGJOUvyMCOXQmyquYaOfodJIDzVN4edVW4Z0Lu8c57+xsQR9o5wLkB1Ba29oXbqxOK9glFkh57C
r3S2DE8eFNJBTKG1CyFGOY4m6NxVOUXD3FMaFn0Hpur3u7ujhXmSkbLJVjy3l64oLmV3Qs4WxJXe
iAsMuD2g2vXLolLshAVKEanlpLpSauF/lkPCatYVLP909D4OP070pY7RqOBnwyufrtpynSUZKeq4
2vLxsF/7Flh5RWIOUrFK6Ang6scelWubwP4e6Cf9222ik9VLGWFhREfTocrn6VOHWaGCHxiLU1Ft
0F+4ZKfnBLpt9K5Wv7UV5hISSBCEohWec+LDU2JGimJxryAWtw6lP6jg+pTGuUqeUtDZJAl+gMiw
jvvn/tU+HeW/L8ce5Ac8usvs+jZo48AUJErNMCwsquTNZIytWDz/yPD/4nGYJj0uhpGWe/Mscx47
FhIo1Tx3lUyGcwcn14Gbp+MYkn4YzPI2QZ6eSnrAGF2ff7vypoMzX5ZipGwndL3DDwJW6zbaufvi
jUkLFOhrb6QrSIN3lOXsUzmlzXjojZh4X7maAE3YPBuJtTjSt9ov/V9xr/gvsFcmI28zp6fsqmc2
JXn0Mhmoh/kdXbhYzj9ZVvHAZt1ldD/przqS3bCZLWZFC7LoQoeboOLIwVghmVe7eaYp7a25zoR3
1ZUiw3RF5lpjBItX/J6W66R+gEx+GBooRG2RnzMNLpL6afhSq774PgnrHjgGVjIb8H1pIXETdqdy
D4bJFHabE5SVPrfSjfQzI3/F9A/8k29bhz/vZJ7NWn9wIN/pZtf3I942qyAUzmMz1IpsQdaIBB4Y
XnKeE+MT99m/zF2XcrmefmKEKXV9stl0j8CpkNeoYqxCqD/DNfMvmVVWNOJstuSJUNonGY0mTPCp
qCuBdVENf3zKc7bIYvk2pL6sMvHpp9BMad6oQD8MQzV0mwfo8WkNF61EX3st3Qo7eRJ74a9BGvz7
cldZ82L4UOk+Vup141GTo9FcAj6+JvHDfAk3nqfRE5UsIHkOR4JBHhqNh8TOzhF8DrhjfYhCMUSl
vTfuMB9XJWbvRu+Ucj9lZWTuKJF9rh0uxvAGmg2KtfToybo9pWvGfizWKhQeX3ymUM5PNbYLpuMi
7i40wYKOcQ+sGe8Kti4CXkZv4VL0e4lEwijbMOdqwIVCRF12cQMmmTfALlj0kl7wk4x0tRAVg+cE
FbEohmjJOCCeGO6h/RxQouNtI8UkZNSO5G231ltGBwIyaTad2F2pq9oXrsb7tBXzadY29vKQ+pJE
6PzBxCZgvSuNoTkPFT1Gk5hc4R9QXkTQuOw7agPmcVTPVDZKB7z159ZhGqXMoqa53h6ZUPbicuFS
BLdhmW0hllTTb0/zaXymreFKYcxDq3fcu6qu5AOs2PiNp9RFU7plPxCy/HKCz9tFgKRN2P7Xv5Y8
U+eD/hgQYOUsPH+d2Tk1cPmXiOaHKq09UNaxhcuzImgiP0jml7thh1u1pfWgPV2bw3QVbnxrcrhP
zeg4o4Q49wqqTlkLWGShNeuKu7NVR2J2D5OWGb4/ZTW3w77bx6Qv0GeQgIqdUtTj+nsV9WpLFamj
LT69VrbLKNsUsd0zKm14h57U+Jl+Kctq8pb91qfx2ZastCm6CmwgF39XdVf0rVClRJ4IF5dSPBHv
iACiU0UO9VOUaAsIGYXpvvVl731SZRHLthTF2vjb5Ltbk5LE0bfvOlesmmbksU1iJOIZLnWWcle8
IF7GGM9EA/id9sXJdtIxjAxTeAVLmK9nXMzBy4wkmXyOFIF43Qgcx9iGNttIjwtscMRZZDlO1HXy
2Jlk/4bdoWovbd8cNkOF0+Zz3PrUd+EflMm2TKwddFsxf2JgRnaquPfWf7/jePJaGCt9rYMcxKsE
aJ/CY/FMGcDJDwNiaU8ezq6SoUtt5CE4Eq0mYwZacabfN8L8aUMk8rYi41FuX64owdyDz3vFeJmy
f3ZjMWLSXIIzpQXtsM7/2gKcdoOyU5YTgbxlL9lUpgfD1t7LQi/8wavvBddZCl8ejd3vZmK4ij9l
00HcSZeqHfO0cJ9raXSheuECf5xtlch2a9vrTiA95MbzOqN2WKM+xz3MHe0BPssnEdqrKyKiz+zM
Uf6H+YdBbuz8K8XyOzokyHvXXYdoi8PNNChsl5hKUSwjgvumW2FfzJWh0WeEvNFjwXfd+namv14e
Yn8lmSL604G6lpsliqzpcaYfzmx1AINlcUBlWQ/Otvlm0iQcdamJQnMMKsGm7bJde8gfdZXyMC2D
kYsRmW+OyZ4phaxB+Fbez+nAPfPzoHwsfvfQGjwBNhX1ZnQ/Ahp8Pcm/aGCcKPvUMkNor9ulWXV3
44qXStA6rb6+uS+1v4Odhla4O/mRmOYWiCPjsYuMLXp+crA7kEewC6k8HOl+ohxWt1AeIGO+heKH
vndoKUUuZ8tUNd77wrVnPXq9qBxc9DFNyMLQmoSOVBPEEWyTSI0MvxYS+2J/pKL94gMIaEoBRmlk
TWLp1TD+w496grsfwDdT1zUdIFyRxp0Es3WXwikKgpdQeo+6w6YImmK0n9tDLXWfrXYYATB9nogV
mP+6/BjoHpWPdbjpjm5gJYphHYYJRg3NjFrNjsbha4/fTr23AvyjnfbV+6MOt6LDpxWGP193IwyE
st9R+8hrT+ceKuKROWoKx8R6jAHXzCWymRzxBjZm9Io2xVBsq3PsGoFN+zXZNFqoX+y8pwibQQ/i
EeAKBkxOxJnG7/a69o0puYYF7EmqouzlgQ/dzLXfGh12WpdJUZHUxQgxZlB4UqVAnZbQqiqTt5oh
V5b9OT+TB77ZSgqPiiUR3a7Kxup44q94w+ITAFQc6fIH2CN7qVV+KpUKg676D0nNP8YjngL/YY9z
7IpNHjkldVoIOrEWPHPI6aVoqzwdxrNjrTHMWY+DIrwP+YRcKrkfDz/1z4Q4XV9behJsWrFGptsO
1Crs+alVxTb335wBnYHohGoR5SmEbkgwXxhjqVZl80pP68SYv2IRrgFfLtAEEi+EnfMjiedHZVHP
hzyGtlRL9Rb4+pBOuOFyLmNjoUstHyZ2moK33yQ+faDJr6dWYteSEOeEShCq4BsoJ6EYtQvl3n5J
6fnW5lu4zhR+MrQ3iTi6PC1Em4GT2L7Oy9H2+AXJ4TnTs22EE7ENQBxR9Qgx9GkTsjy26hXRhu00
Ilf30e2/QzKV9zEA1/Ouvl122CQgV/ThGcOfYY5HSuK60JkVFC76FxsiA/FM8K1+ZrSHy9KVQe3z
zyijvOHAqlQ/PrfomdYIUQRtybnpq67+Ea1nIsMigNtIXA4Vbac9igJiNwAmtW8HJA5dz4yMfE8x
8t0q2FQLPuRUgPSvG3/gF2dhS1LSC/tUDFqVlCEtEwjDvgZOYrmgp+dxB7zHO45CBo05yv9jXgln
ESGaKjZFQmsgdVrstiNbrg6+bfNpMaOX+opJVExM/2hAcP5PXKUbALXZcJ0TxW5PgJdBGGMPRf8/
oFqLhVHJqU9MtDoQwvJROYILA91o9KoeDlgrQGVVBMc02QjCz0aMNLU1hqHzMSHwLSSFcn86OkOe
MB9b4W6W9FXF5Ldc4MHVzRmvKGHuKyHXxBFsGlL228JomCid/2N9IxyMRiO07h9qVzDazRJU7uzj
V7vW+JMklgaat/0aidDLLoEufqy36wedU52vyHWRjdFHdZjIWgppOaZdVqdS2GDoTz3ryVuhURPg
MqlmapdikoXvHmPiIM7AE1bZYEFAkGUF4k35fkh7+ornEYy3qle7U7iRyCB7IxoLmK2YkFOt9sF2
ULbrr6wwudKGFitlrjlkuzEn4AoyXruNsMgxEXrtz2ZRRUWr0Kp+Lqb+71+j7xVbYoZ3WyWiIVsA
Wea0UI2qiUV3Mf6o3A18dq+PW6jdsIklsGpEpeO923dOfGXrV4itED2gjfrDpG5z71etz4k81uIz
q76i/wJ7Ek2aM/ToJXLR2TpRKMFcnBXOTIiAu1LgwsuHqbNlMLBflnxpe/ZnLlmgL0DQzFGqvEDd
unGsAFZlG+aBxYUUKbl4jpDtbAD8qispLAufBzT5XPTnoBnVhzpDcNDtyk4lQECVdrl/B/uCcvc+
N15AALvgnWEMkJ6OCOpy51gZHWNeEhBFI91bhPwP5QvYo4wt+C1NDWrmk81HvQOKMpZ9r5xu3sHw
S+b2FfDAxJpb91I6JDoHyBUkLxw/6yy/VBfEsl9bQsN8pA+5Tpn5d7qUMER+tYxcCRCyNphvY/8j
8VbuBiW83sPD5goa9XeBX68MIpBfPfCf7RxUGgw4OaSyUOF9m8QTjLOPcEnme220tylhC5tTzAGE
YWNzJwyhP/X1MgZ9IWIcpa8XwOtF0J9zDc0dONQzw4aS4Tby/0v5cirPDLFo5ipe5PbFnFzPKKHu
N47XD7th7W2/5RpUCxGMQ4J5NcvwFBzxVKAc28UfhChU+gZMAw5gd8WpIzU6trdaZhIY8rEMftSl
1EHdUAKisHAZCucPXjeGUmCQwM9QyjVfuLiT1F3R2zylE/zL4wzqAOmXu8KPh5u4FecewdXlTe+L
tJZF/AbDC10JByOuvZsYuLidiWUqjvwsPjxA1x9cnkfpw3RuRnYJwYgp3avzCnxWhDxwqMHBQuMp
1vxnsGOomPCJ7AZHTpCfp3Mf6DAQzS6PizYcYnATf94nQl6KOwVTMi3px7JCzaXI54HdSAiS593y
7DhopqdvgrXpK31Ed9Ws0KpVLBcUMHARgHlIAR3RwSpqJIZh/hlQ5ElxAnzPo5k/FpvY4YZCXQK4
a5H7ZjjlOsr80T+BH88acn5sdy4aTspgXhBCEyJmGt0Owhpkb2fhfNZBZpVhNKZYte3DD4I4x5PK
lDiEaxZGhDXn6ErQc5i8mrLyqkK0BPq5ScvzJ3ibpMooG6E405hoH7piodBGe/5sJaRF5QVIi/Xu
YwKEoJ2W0TAmhgMifWXxWCuj3kA4V2UoYJvpDwASIJHYeqAQWqWWXdAj3QioJ5OZxSZB/j0HFbPM
ILKIW+4+My1XmVEGsBrXl9nrIH9pqAcTKZ4GtfgeKOahdNmGjjcUl9ARbKzx9zOi8/pMkSFjhnK4
T8XnUSoFmhZ3DPFrxeozcNWReFIp95qj58geXRo9g7aUD52iDq/ieONGXMir/jm4DDv+VxjA8p7I
GG0ijNXmddiOmfNPamW3ROniyHvvukZ+xSN/k6Xxu12M6xMpN3Dw89r7zQX9IpwwzS6QQ3lZn3GV
AkWadtCJRkAWJOUIR5tN9P54JTa5som7f8+BfOc+nbFEHE6aex9N7jzkJ9Hkekq9JuOXvfzKwYfz
M65hlnTQ9jCdcDmZI3uQzuHBk5XjCJQ2DdYWOLhsTkWz1U3TNbSnrX+u9ilEX8jjDqDMbghDEmvp
Xph++tlKH0PlRYKe3+GrTdL6jI+OKWsxrbpKw+O15TYs6GHL9dSILVDhUQbiEulLT03t3ZD3tHZi
3SH2XRVKcw/k4wwVDw4s2Ni+FwhtOYZZv0uQUfrfF8KIHH9MXzkZSTUXWoUTFZG9N/PJrnOwUSsW
+zce+dA1H6bqY+LqvhGnsmVByCVwx8vNSC3AfE34z76FEAQDRnQXCZLMmXW7Qfe8Q0CQr+Raprro
telw9JtmeTVbez1hrieJMXD3764B0VPusF60UohuGxu/l3m8r0CEsORaeGJeLu9EZJB20sx9mH5F
on0wHZ+CVcCWu3sfnjBwOD/m1/QRUWZ5O4A8peFt4i0eS+VSvBijFGhSuDnKWY8HV0gP1OLl0cQM
IRa6USc/o8y8LDiD6MhGQXzA7DQkLKhzGLmvhnQHivwP+hwjK2UPtULIRjub6YsS3nLH8jibk1h3
iUVzyjMWnHplLxW6IXYRCrgqhlr3utwsuZvHJuUaw2oiXmuAXgtRDjoSSiKtYhrUbBO6EWkFzS5f
694JyNv8EBpyWcWT1sLXPio23EO1vCGqKcGvmuRRrKyCdME9+tPZ68b3IQhb8hhEjiKgHBGVTf0+
LkXXVo5aUiCIHOF/M9H16X1rGJztke2Zv9JaR6ltWviXTSHevipLQNpqXTJcf16l9aNolYRnBIww
CRX/7AVs4rZktalfd/nn21Vn0lRmfkUVPvnKv6jJeyS2jFnXce0J4L0qTJWp8jXUrl6AhzxD0ZkN
qZmtfxYFGhLgLR2GioLg9Os1p9o6XyU6z35RGm8YNVXou3W7mOa1BzS3lMzao7wF9ZUevc+tQ8DR
CeDF47Ocbvtq9/LNqnGvOBAheE9G8QxDhMNLSpPBlP8B7PibNJPUIwtsXgY+mYYai8qoCZa1Stap
UPaDstG0iann+W8iplFhdxy8o2TXJ+UPDHvu8uEQBj6byvgy/lw31/Z1PX90g06E6mW7333/nWF1
SVhoCIpoUPSDV3pnmYN5QMl+73vFt4UvjOlz/3sF6dKzh52jZVmM+FGeGKjVbvaDhIe3H06JLDrJ
m6YPbj/+XC5l9YaJgAA2ZewiMxSSonkUAWRbf9By7k0ZfMtBcEU+uxaQXTJJOSVcAgk9bgU4tnVJ
+yVSXBb8TBwslUaTDu7Oz2ayaOikonsjOSmFGIKtauUS1gOkChFILBisMdpVR6WBbfTa/o5Caw/L
SSQ0KZdkx5AORl7RVe9KCoMDT5lBbDn5St7HS5zWDEopFzirnZqiOlojlpEENq+4PQp4wCGUWngx
YS9QUiu6ksL85C5dwDU2Qx3bBwCW5xs987M6eIzbWdz1w+51i1WSkIdDAvawryMeOSku37EXvwfY
+DuZiAXNNcxaPJm40BkUSgjPMABo3BMilQ9Q7URlFHS1FtdF2f563Yb+pM6SUcf0J+Ea4da149YJ
Ahu88vfoCbKQ3C/np7JhRjgHt0z63p2Om4Ite4kXVrxzRLRd0AeyXE4/u64xXGSVwBVR/bj4Mlgx
g5i6eHI71ON2udAscJ5uEeFJNAB6xjivSNVBaFU72stPogIo14n8ph6AG5OrciYsQs62Wrriywo6
7/AQdrr+B83H9Dc75uDFc3pKr4Ou7mzeeCWIgtEcIy6EFppBzaNsKxcSMS0wHLYy3U5pL0f7rSmy
lSbviao02bCBYmZq7/Sc11ndNFybME6yaw217jQcbux7kQPBBFgQ7dmFbp3uxtgCnxfxqHchbIwh
PV8r5MpKqLChjbf2zV9lejhK3rlQmCySrXAfL2A6xzb58ovzlCVO7mwgIL9yNW0afjsxrjUtXHtC
GOHmJd2xyJ5wTstgsvpMkViAxp0EJxGqBNd+gOnl6HZLCCn532s7H4zEZY46vL6SfmiilIN0Y6Do
zRrifHE853rUr9bDunuQWNsRn6sHYBNJAS/8N/0sJKT6A4cFniZISJEO9+LmV70SGzjkxEfM2RZY
XvMXf+O3nzCkDq6Y+qqls1LJhfshaz00XYRDp0hWJb0APSQ7amD4MrN35brRbAtHbFR82FBBdPJR
4oTri2idi5Q774OpWWKkaVSmFYeV5d+Ad8GY+J/QpgP/1OpNIyCgsIVsH72qDTv8fOFfkLUnnzTj
0ZB5lPKBduJwyP0KGmfblQdjigHHZTEfvUepRSAt6/wySjTjBxHwEkRAJmEibUgR0xFZnHCPnQOi
8gTWL2lW0egcUnK9jMtsZWk4SzBR41WIyZwZjAVoqaHvSPgPLx+mEmxXFCnu76bWEN9ojp7tRp09
h/IzYJ7yaAR+JZE3nRmtGBYJsIusY20uEPb4PbFKv+kkLLmQgbPYWbvpUSFjmMjmYjcMpGFsoU5D
I7WaY4gpbhUxoAmXIXtB57JmcXDiR2wIJNwUC250MI8cxof9u9yHzq0eMD0Nfpbge9mYmHRA1tIt
nBL6lJ/Z5QVLArh9DtzOqsz+kjbFMhQozWf/kosIAQn9cQYQWD/2dGNd/3yw1soXahQ97HiV2DTY
9RL220cyP/0G7HrFSQ8jFoE4EnTg5njEXRMc4Sg9OPC6RGMCNj+xnLUdpU1VIJmyqZB5WOnksvoK
mGeZMsuxeMW9EUrCjk4QFicKZZmkG2W2oaEwfw4gmICv70iyVeBeUE5wh7+ptCtgsZfAuFGH6BZ7
H5kUDOljVo9ZHpm8a4iX1+6gTLN3IBpRNl1f837zxrceMCBJObMiSN9pBceiSLH9d5cZWrN305sr
JSn9kqbwRWNQnYKqjnD8oKKD6rCutcUYksoHdOSnSkFGn0EfiWwhszsbNZgKfupjuBFHOnzgpaqF
5jKdg/KkRzBw+rgD2x/tTpaTWWHr75eFTud28BKgR7n+8UUzSDN0IW0unD3rBHfZvrhMTftXa2Wy
3fyQAHe5eM9ZlKqWspunsrLd/D56G7tYs65OlI5kyef45dWMZ8Hmj6Aany2keAyK9mAXLT/+g+j2
/5d+UgNNiJ0EomqkdqnxFXj7+XjtHqhHZz7KWVtg+0FwROr/8XiykyUWNpYl494wpV/ZSJ0zUR3D
gbswg3BfqKHLS6dltSO9r7r7jYTOKzPpxfJgUXx2jSv+USJo5ZiWeoleMxfTGyn8tJqoe5dcZj/8
+hm29c9cL/Z4kJ8jsln7NLR6RK2VAUWzwR6Jx4y4g1RZION4Oc7RgNxVESqfx0W8kiLWkLQz5Lr6
4fLmAiSc/aOccqx8BZTix9TAJUu2LVETilechC46W4/vfKf8ln9Rp/hVO8j5ZAN3M8J2htJoxB96
Ib/QgQw/9WWaKF8qLdDOqYvuHYfhSxKpaplgk+YrIR7FUVWSuu8OM8RsSwmYpDIDGW+JfiHx2iHs
fA2EiIw35k8JS3gmvrVvp5xQ0UL90luWlntY8elFa0DiXFSPHU0mVdWo4KAyBbnTc7mJhL2Fm0GT
WBo4iMZYsVHw3wa7FOQ6AgdkazOSOOjs7QrkgnrF6DWf4j3IHGBksQdpdNweP7/wUdmg0d0NIGMu
IkyNrksx+z3NSmpKquGBKd5VeOAyZqVv38nsrqusET2srezNC94Md70BCta/aqfFZE4INGgcudM7
eGjEY0DqcyOBjumqQteRZ8l7uws2HdXerwCE1bUsB0AtV37TpDDT2yG7RNxUH9qoCQtH40j5fKBM
g8J36yQZNkzYKEnC7VlKBhHgZfS5wuK2xVx0pZEIJN0Mm/mGkPVkTV2epxfMvjECgnhgzFSws6IV
B4HnZg4/5f2+xaGPezpsBPl8J2AsNR3naivf8IBCpmngE182fDCrXjNlfH6kxAScv9tQZyqjfQER
KVPEhg5zv97bcN3qw1Atj8NNkM0HQrqi94+qFPVW5QMirURqXP4RPTyWj1mZc17WwHopOwvEysRh
wgKX7pSrtwcbPkfMVr1INkfRgSlkdP7RAPSMt+jbJRIwcNn2LnqvUOovIfI7uarE2duFGj8Vx/p+
rWETRmVe2WbEf2fke7rImF7rheOGtDO13TVEZjus1O0SEO04rQmvVY31RaAIJ4wIj/DYgD6SXpMl
1a8q+3IGvOHZZfyryuxw20CS60aCLxAM893lG823YL+gan/7Bj48QVN17TCJOFpCDQLJlckxErOO
cIaZ6CaO1zxuaKKaCLKIbml1F55Lvpf0yztI/3B3hbcoEZWouMYOiFH+u+4Vg1DWBmqSzccqWDLq
b9fUpjFk8zyVr/hG+aDN7ZKBPt7sH4ufToHCPgf8S1zx/12FSA3NbttPYjb+uwONmc1td8l8Dsu7
Ajw+zy3ty/ZBB6/naLGfU2fGlKmitf8cSM5LOneAbdun4by+mAztPRvNb1WXSdKNJGqFGdZnyNMa
lfqsx9/qqRWzyerxKYT5Bej9hMQ0Ua0IsuLa2edAq6Kp67w0lsx11COaPzdqP0zH2hqdWFsxNHz9
pArs95vCmDKb+hNEengO2lgT61/zo2g1t675fkzaXtxrG6VlBdQQYHBdo6MFvwyUESajkdBPo9Jq
ig1Lzjhp9bnCLX4GnY15Tgau7NRj3i3rFkl0zXDLzLHau4aM2qPNiDyNUpTdHEIBDj6sDL2m5Mxi
f1lXX4U4n3B+4UgpSfm8ZwpqWeyfqVaCzW2VPyMgeRCqLu8rhfL+C/SjbSybi2zMZ5vkjQYxZyus
qMRD6KK3iT47wTPs8Zy6qQZvTVYBFaijoFx//6LuopeL7GmFJfDOauvZMWfKg/Csh32eUH2MNIaw
5CernJ+5tcaSzLeJXcfTbi0h5mgeQBzKxyVUIoiSHv+pYABlOtlCBaw3GcnqY3bRboLyrrFjdp6o
B4gFtm9kZnuieUztmQNkhBRR2ULjtD2z4MB/AsPvbyeDuz1/6O3hH4BW1I6gx2Krwcs5zw2jT+Ef
0JXkzXS/BPuAkrKsX/VxpGpWqCgBt7ONh9VctL9ZOC8xY0RsxsQnT2u96ktRPWfuiHVOS0gZO2pb
qeOGBe8Q2+hlNsjIw3ZXU4TvxKnhDM2nMLgMSZf8bDarqYX9spWgyOmtaIDBYgZVdvGG+iLwsYEm
ytcTVXlN9LXBNGuVzngB6uznXHugFGjmQrs95GySeprPNSUjpa3VG+BJeY+YjID6bs2Dy58NZ48b
i8h69UnFbJ6WB5OnN9NLlXZfk20tCcY/t0YoXW0ZnwglwjJysLlnlensIhUvG9FSF/jUwe473E5I
oFNfw3NbjW/ngus4tfay/ZI9xFfwt0HNHdesK4wuU3AIlkCyHXVyUHGuP+GEGb00W2LppKdI8J92
ZaaLu4cijGF/vtAsXxNnlvehATvMTSLByUEDpyOiFUCj4GGMKtTQpUP+qNzO5//vgJIKuDt/OfY0
HJGCwSM2k/nJ0p5uwS0PV+Ykr8K0ZwQSMjj9Gn7RWJeDPsp56ZsgtL40isJR60ogXbnQVB1Ce+FX
KF8DvW0kb6kAqn1Awz1rKb3d1j+Mty77Lpk08wpXgf7sSRz++w5Eey7ehfJc9aEdZs+ifSgJI3ml
fXZNkrLK7KPaI21NiZwKVnXDDvGz/I0cIs7xEf2za0jsQHD6WyvFFHHWiWJw7IlpWNihLNJKONNN
JJNzdMfTwjiBZhVx5xwKDXncoFUqs77WIHor6cevJb2s2Rqv0fOheaV987k+fv/ARaKWSDTksvSQ
GDAZ3fJAFivX+72VEH6fm/KvI9QZEN72WfV+3QqsRq7L8Ua5ZJL52RPqJQosL/8zLpyMC3Cbb0LB
ZFxaXg8nMdQZku00bPo6AV2g4Exvm6/1XemPiC+c8BxVMeLnEMSH/0uqeAe7ULsX7BQEYtYR/hwb
uKH+jNUhCqc9AA/32fPIfiUflDpMjojXKXMI88jpF4uon97p65EfwEgOptDOeGYgEDmjUqsdqSeV
FcTTjwaH1J2qK5A0fTfRAbXaJqseO7C8NKLTDnqe6wgBKNyLu2b0NhvJH4c5ZhY8WNRsKp4Xj3ji
3zLdsX+NCOXrM2aX8J+LrAs53rU0Ek8IiBYtDqcJeODeLVgVrkViDS8eFEws95Cd4PKT0iwqyCB7
G7cMysM7C+470EXzbpTC6H1nY4C9EtnOYC+JB07AVNMnEnrwhKOMBDX2TofJfYJj4Ou+Tc0Rbyaz
ZjUk387xuakyNzFi/4Op7sbeI9k+MI0uFiz85ip+Vi/nsqHG7r14wnnAjK41ibAJTQ7ObXPd+4k5
4zTXAzl1amhxinwjuzsOeLn9smGiUEqRWWo2aZsggiKfFM2SwwyGkNevWiULDiCaIJuJag87UpsX
cl5i9jSyavkoTqZzT83Ytw2sLaF26vPE7g7Hr3EKB2b0QWyFmMQmtWX6NbG91HjdvmnrmL/q6Lfe
Cifi/xL5DTfVs9t69B0TH/8XPAsn+1KcMnQj/snH9XPpDf4kxzPgkz3YTSifCaaprbSFfd/fUzRg
Z/kz3ILNgnvMxQDM+q4wsD0RMDK9RIBKvut8vNPu4NsLYql/+sQwi+QsJF+/ixK515WaCxo06+Dh
Szq4aD85KRjBBsjNCOVZL6j/fSNr4/7IQI02K80gKXlGfdoS2D9S1QDa4EPyOE1/iHkc+VGL29Ft
LLDl834cyZbS6IGK1TMCNlZ13UvjJ+QikBmSB8Ed+rMtcKKALJ0Y3OkWAvDNPZyy2VNyKK3bcSey
UDODW/PCfP7+5HeTuAwNIuHbI4iOgxNRXn1Dg+HLMred82BSFoASCx+T9kPCYq7uuqVgFZMeB2pZ
3Uy8iV4ZhnWVMSVHRTt75Ff5Y6in2cu6u1nzLbiASAUMBxB1llfc9cZYAX6xppu8jtnUxj/21vz7
Z2tbKIxjc1APr5rySRF/ikPn/dqTU9QzrIjWgJShpURilRikqvu3dCzPhgHy4qM1JPbsMljOPJCg
fQo8qPFLFBM/82fV/fzR2w5eu8t0ccge0Ouem6fRUktLqR/qy20NAFp+gHsV0kEwpRvpzAMHETCu
isu0GF6T5xtqSj/T2YZGpkTNAYBVz/pFmoKS7uM0XI7qa0yd+o8VGUEhE++nu1p5erdxAWpC4BR6
tg9lAiPw7KK4tueluAGLtUoqmIDG3YmTQw+hkRb8jGWzDmLqGBIxJuCrEiYq02srEf8kSKJAdsp1
NEmeNakIecOwBdBY+rqymA4LmKPews3po6HkZUlVks6LtnbB4oblHtJ4kBFn9jxonRCwUQzf+vru
FbSZE2+Kn5w1niQyZxoN8CJHxqrTphcVnxsKjxJXCmYglk7vU8SHgdK2x/NjIjs/Q9/3/ss+Qscy
wc4/lW0NTfgSBqcSZL+TZA2NfT2hSoto7Vhza6Z8oiXTLclCSH9YnerPZ85sZEXrt+4HI4dPhx8q
T/egAnPKTmyy+9qoBcDgym/WjrY7fa1biUI1VNg5whVu3EO8bSCAt859KTanHdRB5j7IqYVZpl0D
PgOINpjHZydQWsOttf5WhmpiT3EijBC4TXVOE94XbrBAoL0ZIz49irDH2Lsz95yjfIkwXbhRGRIJ
G2yxjCHktMwZ9Yqi97beD3zF1XndVoQx3/qBuSC0HUEJNByvtuHZHyEPaLZjYTOVkWm1ig6YewXI
PQXeq+dbXjT3jL8X5qmuiI5Ov8rYiqE72c+34a7GvtUHxgdGxCTAFykEOZB2/SEq+3w1HayD95fW
9BSf8MbBuSuxGAJo7cNvyn+bXluRTKEW6N2jVZq9UnS6tJdlvOoUi+O1VLqD/SBeMXEV4prU9Vow
IliaZxX97h/Y6Y3/D7kKMaqh4esmF5RpNcetTfZFzrBbbyxBZjm9mZ8DEtjimZ5C0toG+DH0dMfA
I+HbPslONw92eIczKrm9MJ0vZonJyMrhBnQtygnM0uCECVnqOluFXVXQkAk9f56nYHTh3ORRNBNI
RSDR/6zUmIq2T+QKVKYyFJ1IT3W+cJpNKkiLW31aCHLGAlrz/JUUPPCEqIwN34G6RmeBi+Pb6Fn3
EbA1lL2uk0dYBKIFbR36Fn/F5yAj8bKPNetKrde6u/YtVikq/40XsOdoHhDMv5unWBNRO+jgdP3q
iBc5Ei0E//cPbfVDYEyEnPlOnNTu36IRQT8WqnDNlh0BWDpTKi73D/gH4g5lgbzctcvXR0XCdvNu
C/4be3yUskOEk6ThqNs4P7URfoB85Q5B0XPqiLspDWMmg7pwUalXKbxnv4+S1DfWtzlym20RJSy+
zzBgmtSIv/WaVp4pKvUwIB5ttC4Iu7I6eDEnZa/n/dlabUXmygYOBWeLBPkwsI9Gjg8ah8WGnJ1N
FWGb69vYvIhs9a39mhPe1LriMjfxHxIXJc+AgqpemmihbC5YhqXucBpUIYFiARU6bOsDBkQm3ZPB
TuLk1/RzNPplcQoT3Vf1Aw6kmziFYfuCRMfQ6gu9l4rlOCm8MZp02FiEu1W4VQ6ZQFtnex3RIJWF
xJB6v90SGusZlqpiANhyO+I0jykZixZeshpcxIpO7r0eDhVc4bRytPdKkQIpQDjCyCeNxcCtxosL
iJ6GaO+LBMSIucUR1dVx+NlPX6P0Zc6+np2N9GkL9q3pn+ARBT7Y5CEO96+sxn/lJ3LVb3d7rV40
T4f03YjrhcGBJ+fpgXShQdJCff6/Y+yANgd0RxjwGJs/PKmQRCYBK3DfWXHmYTaS0+iSVyKJgami
nQBiWqfGUoti3JGY4JG4uzY8dk4h69fAWaoEvCIA2S8L++KZ71bXE21RCQm3ge5Kekdz14d2+HMn
co8OjH/O5TRAxPlIbONeMOpv487doWN21eWh+5qodFubgUE42QAilj/t2jlYdsqMq/LbbmBe1XnY
Z3FSpUWnX9NeE42QEg4DCmI6E03/mfO5gCOZntxecVt70XwAGypF7n6k3RKcm1yxzYHNRL7pwpon
o+tiSO1qMQYdM9XU/uBj3YbLhDOs5wU5HxQbT3Z0XNoWwHyMMNKkomK7p47W5WZ479Gniwr7BJog
Dh4f+cr5/1gqLEpITg3WQCaUUGjJPJAhKzh5YbZSRwsFxz41VwCTMRrhgLkPLAzMWpgMNIWnZ2Ta
D7u63tyJEivQhBrxcCgfBUxImyJmhKYjpyRqRhsmgyaiLYK6/nkHtajeTI1kWxasdhWPAVQ+s6e4
gd56LBvX39icQo96RZd3Bc7XPO8g6bkYfj1K5NVnIAsMjUFy6dxnE13jgWbPRG7p+thHRXlbcYnm
WB8z4LbEgKxmye+AlY3cx5GYvtBdpSg9LKkV3RSRoSwKgnsuMGtX4S27rIifFvA++HCmcyWUdO8e
ekzxrapRrK/fReGiZTpvB7n89bYrs8bA4jliQl+GeBpzLT0A76UiLKXxem3PBb5IyyH/kKNyxZaH
3QN093w8x16KoXqdEKllNxegOvysKO6Jc4dk0BhtSmAzkbm1wr7n41rWdLswWO/HeeJ+DIKq0mF+
lbVYw5pXOneZU/+ZJiWZlIsOyYiwmyeZJLfFa9ME1oLCVG+QiQCQqvv2qynTvPBRacUf2IMpQgGp
BWb0NQGr4r9fR0WdL0YqoxF5tzjm66LRGxScgXkzCAwEihpGhwUwTMqGkRryjzSA6Veg2IyTbD6n
SSy0dLL4HV+lfNxvjUfYJnpNV/HPegmD1xgjqUnTqfNarTOylRyIfWkkiEZzU0HqnmRq7gS1u5eh
nQcZT8m73/g1FdvHPidY4Il0duZ/pofVAW6ZL1SqUoxW5PDN+gZktCGxtgDAsxS+gMeWYcXj10DI
OyK8O7fdZf7uWEt4svWNo+UyeSZJcTE+cHX1mVfiVJwkHQXLC7e8LgWMyjjwKwdhkExoonBfX0DD
ZhhGoequtbuwQhVmNatDcCh+nny1oOWNiaRgbUtYt9DQsO8Z17CSCIj32H3egdbD76c5D8dZ4D4Y
gAlvjpC/NczS4NAeAbqa7a7K2/L3D+InTuJl1vnMZOa8sFdNbeQoG8jXbN9DiAF8GxUVKCHqmkIg
yZuRETcgucgnhjI2RutqrIEZyxiw8PXZk6Osz8aNJvStGD9v2v9feg4TfGP0uGMUpEcBYEmfgaov
Gc7KVWvQfoOtfbfxeZYVMQM/Dp9TrWyGDcirW4Xd2gjpigUpjjWp8oezbhQJIFej3MAsijXrW1Of
A5j63FmPCg6fWN5eRIhb9ACqWKEM4pdmPIrDTdNGGKOaJrO9B3KubzQmmOsnkFaTjPt/tGXmcy7P
lva4eBuNlb3ROkt2QPKT9ONQ5PSJa7WKiDby/+gtlYrYsECdAR/5JKTe+i2bcYxTYUIQj73UB170
ybTQT+yFm1/ShCUTWTe2BcuU1a9Bc2KGSWq6FYYuy2NRy+WL9EfQXwhemLfV0uF9KnJkRUB80bTp
4KObktBpPSUR95m7u2en2ynzrHni57cjz5SleA94nsVVlPBzg3SoRVxLRP1Vy8j67nStRQIlDdQW
vyx6Xykm58NmWPBAqv1maWApLQ8Jctyswpy16egFlFgo7g9b5WLTuzBIace5DESV5qZXJxjdijL7
C+qr+7Qz56b8+J0PeFuAxhCCvDzh6p8KICK2GP7G+08X+J5KUg39hlXTsrmiXa+7c3M/F53TU6C3
jwW04P4qEOG0cdMcD0Ma5uMIEaq4h2BF7tzzb4EpchTRsqTba6HOcOjA8gyWGvwXui+x+hkO5aKx
wK3smqYQBNkQ8RE+fwoYbOb9gmeXnynHsCn9R2kMuD08cj4BxeLOLreYvfKltl2cJEob+64CtGxc
OS2mSSNcfeux99OxpsesGn53nVbnWLZhUUESoz8EH5BzOee5VoLi2EWuQGCJ7Phks24RfF8IlCK2
UlF/U/snMJ1Ss2d/hIGZnM1lMB4lAv1+vZoxLiFagTr1TEzXKic6l3D++bjBawImPG3hWgB/WYBj
jBJHl1ck8MiUD8OO5rTiTz0F4eVoxigNT2M0Jp+C9D9ebPLban8g6wOSkDzkxy1kzrDc3eU/A6VT
ZPoihCaFV+EsfsUEAcmO7Ba6YZb1HVJ+OhTRQ9YEIz3oz7UEwowrLEU0BKeJ3ek+W4vbcPMIubZO
jN06spR95PdzFzZCl8k1BN7InoBDGh9xjK9sk2LuKzSO5qRbVuaQfcVJsbTIaERzMFGmnJQq4A7f
IPR9KeWsxiLQxhNX/Sakd0NEAY5XPp540a2TbvWOkUgGbk7HCQbORtzq7EezB8HnyIK1WWapeJa7
hr6gOTh+Yj8LfcQbKpIg+KKNo5U7oh0D6Iyi1tz11H0HybJC42ZN6TAGP/EXAl4G8E7Udw62LZgs
3Vg0ICNK+pmDZOCOM46dJt8DYqmRSTHWkSWp3RTzinnAtc1j05IjE8F/UimSFeC7Y/KruPgLvm7h
+iUu7rQraTbIKU4Rq6CplLM5oqZyqHfaIWhMpgBS0khPSPeN3MBbSpWt6RqzRZKDo+vzCQ61DYq5
Tt0n6duTeifxaRQkvq20RnLM0MgWX5TnWRkxhCygO7KBAgml68PMwapxBcFc9vgGPlhTOIk512aw
Ozb0jUtJ65ew8iG0BaaTD/dnlhQMaX7Q8+F8vtEJdQMTlgG1Jf2UDlvOY4y935pMvnK9AB5f382m
ND3MjCDzvp1iWl6r3/vDoa34QHmsVFt1AV/uQ74QvTtKyZ1ZPtwvsfZVMl1nZOcbC6EgWZB3ipSw
4jV3JZoC3p5B8IuS+OE2JbbObfff+inTxs3xf5Y7In9aYiKAN1wIxnfjDG7S76FN0otDxJZyOlaI
kMcEVV2eifigxjUsJNpccUUGAZIKnBQRvOJUJ+PgpwWp/o6TKjpCH4rnSkkU1FhcZ3ZJFe6tPxjs
XQBgbcHYQHpZPb7Tf+yxH/9hUqe3/TxQAMjk2o8Tjmr2v4cyqYPHGOTnGVSqZcqCJ1FjAIWp4xrQ
s61uaYzj5IDauvdPu8fnKwycYEZrf4bbvwk+GBEpCZIfqYG9829PDfwHDqhy83XRMgrWQa/unQD9
ssetay2slsFBI8OT+GplrSqkEic1LryC0VJYwFiTfpGf4c6eK+l2OzGrY06erpAV8ISMxM/1A7UL
j+NHFI0efLQKzO5Ar9ycUVj2MLhQ0aazntjWKMvp+5XtNw3Kg/IufQiIfyvGElmS3/0o9YbvvaM+
lXpQ6O3NhEeE72rWXm5vm8Po+OlCkwEIPqGRO6eqXeb4I7U3n9M23VZYj0WY+tqcpJqdyT03C+hb
HnkZoHG7SkQtJvCYB8witBo2p9GLNR1ZF8lHxe3brWdJ1+5sEwQo+M68PqDoxmvPNRdCgPK8Xj6X
TTH6RqRf89rjWAzn8RqJZP/2CrdgMaH+6sZW7MMj67OLkKzeMW3xF/LhYsVIK41KDDZl+xuSFyIS
9GBu9yKMpq/vpGaet+9WIVTzDbSithPx9bhs/xGRZ8aHdVhnpcOhtMw3AbHCv1i3APeeQg6zOyXN
Y5KcKIG+DfVXa45kCoxH2oFTmKjnd01Kdz77/LosE11gnP5kvjeDsfNvXMzqnZIT4qH2Xec/EbZe
tkqyiay+mretOMIlKX7tEcAj2XIrRZGHuj0+9CvlMtQvVD3oq0W7aWHusBqFqj/Ec6/lcpT0fPaT
4pfD/Qkd8VEgJGu3vVFuZ3ExeMfM1z0jmWAMrIeSE1eYH4rAJ4Cz8KkW/xV6WS3sm031M0C6U6O8
Fg9UEGqEQ9moHs5p9QsckYxon7asL4JmE8PiKY103SzFHVCIOi2T4NmkaLAYaSqS6rRh4yrCvsU6
A72lZ/FTpZjFPMS7LeQuiKNKIUDcpLbzFrWFkdEAeiN4YROELL1923reZdJAx3P1fYBRkBSm16v7
a7lNGbkqcbBI5BJAeGLuKmyGBCPJskd/z42eaKEZsgXq8xxkrZ69pOjfLQKP1VNqeqjALKLRixmR
X8jDO5LC+cIn6VogeEu+Q0tH+WJdOJ3ZCWPYHAXcR9yf6Ha0mdtPczmqohzLRKsxFroyZ5P66P1b
1szh7qCnr4n2xtYhPR+zieZ8ceDfkM1VoHOFUB0ztLxdLiQ35nPmQQNPde+J8i9ig8+v8DQjAOL0
JOP6ETo6lDLBRZwsCsn6mp3N/LM0w4AkzqoZtbg/XmsSuTnTwmj0y4CDmF4x9Q6xBbyEoJk+womA
S33kmfu+bJKeOHn5Y6W2pvKS/IMYYA2kskc9dFDkI8UeNq9osSnlExePr00uhmmw5fK9TQRFfJp0
V3/6W0QmQVxss2N+d38qzWEqcUEEfNVekIihkCgp7sg2LenDAwijR4QqRLSIxOr1HyLl6rFdxo7s
Tn0l6yeBNyzp2D4KOq01EV6a2OrVFdqeIxrviIha8rYaviIEHA67AE/wHhTJ9Cs/eqXDEjVe8YXx
9ToANFfviHIuZFs4a9p2EQK7PmixKOdNGsHBsyc76ysnk/YowJPozu+Jz2u9H97aWNGgpOMH63Vh
RGPHIFk2JVI08uMA+sDFzliX66uizUOfykktTLfaFGqvJCTXWJeGE8cB5VbpF60VcByoTWsSSB1f
YgBEUXXYeGYqOsCronzCBMBuCTlzL19XFABy2H7sFWKsQiM0OJU5DG57RlvCueYVd3+ZuKNfMnG4
FDfnAX9kljMzFxoWQzecCr69UePj7ITKqTWbTR45zXPxqmtR/0ckZQmtQ5zfUUjmiptOvfNJJIIa
2fgUEPE4ai4IJf7VraZ4NsyDZeG70c7VoXo2XZLVNxOX5HUFWmLTlJND+ieJqcAUTC9uEOBL1aXO
9g03QceggJP3Ezsi+qhdyiwfXGwA/p8eT1GOReQhDUtOtEosP7NWW/dEP6aL4J3C8WzkccP7KE3m
vKhSuK4tTvLJLeF2FRjuElpgfrmQY3L8ljZZRih34eUllWQ5pMBpX6dTTaIqx2N/PCdpHSQqt1Dw
skkvHYje7IpB1AkAOREnBn7rOUVQGyopaJRKDV/Ih9O9aMF2CJvxT5eVyFEqUEsAv0bC/dmsZUJZ
VwsYVcYa96YT1jvTQ4GOYMfD5iva1Sl8012cHZnQfiZ9CTu2Okpi6s3cEUeOltWR+AjVcFPP2TsA
4HxcH9l+RuY4FxqhOGA0lRZUJPs07U7PseS2FRCcTEfRNwdU6D2+H0wTw6H4do9Bj8NfLo6nV9WA
QnWrsQ10otqdiX2UFZcuFCzxaxMgLt3IjWcPDhPGjU/SBGxUGBA3RiiBKsvHZX28qZrop7CLns3j
nP8aIOKxatkGLU4PJJJRLPH/7mioJbXu8koL1Q9h+IDLlDp75CPQbZHmtC7G5UHYcyxW5IVa8Su+
+B+UQgZ45tcODFytoxF4bwhShuoJBejf7qfe2QbvCz2cuY4qGcEhjrrb+SKNJkYg5o+PNzAtyVGd
lbjTKFszAb2ld2ZSUSSjB9gG5Suf8Qj+WQhZT57AAKg6I3HGitHtTvHkxgvfk792WawvIY4oPSIw
GLbunfUjlR0+4hDtePxBzf2bkFNEXQ9G4nqXtDyTSQotKR1AIA2GIbPec+xT1IGdy+PgwDTgfpNf
X1UhjqtUSZesggsRO4AFNinPlFMtJcAQ1cTURC0ehSeq7TYT3MWnbIhb3ZGFGkKyr0wSGHgQ/iKg
ERFc9iyafAYuT1Gl+purgj4/xM1gig5XTfhHnINTrFm1EpWLI7YrOypFTujRnZUvwpyhGz2heer5
G3gR6hdi0wNjhnCz4H+scajwUjYK69PyZaCeQ5IlP5kY21WsyUsgKhmCjnk4CbwWRAOpvOlDTNqw
6Nodl+3Iazqn4Wvaffv4VX6aOT59Tt1zLswMcA7aDDjLTiH9B5QwSEdfg6V/R4ZvZhO7hEmWy6/y
MgFhSX0EawHzIrcAGU4EDpU2mHm0ezf5XXi4UO8SGEysfbgjSLpqWcpXfjUCPUuQ0rOJQg/6k5fi
653cnOcHQzIraobMLzrPzOfVFfcEG2I5ETKHBZCs8kwE1xx/RB4oLwWZpnsLKbSmJ0qnellM6FT7
HkubB0Aj4w3Bs6WfXbP3oOwra82TwdHnd95LyhhXZY8Ppogs8EONflVNQB94Br+qOTCd+vVGuHyX
eQ9MUrdslBHjUP6jSZskUrP9GyxvxQH1DKI8DYjG7FcoRr2tMghqQEQvo/Ulp3/5mBVwepeezarI
2O9ssaj082Mx7cDYhYhZDCJNRd33LVauK7B1ld5U9K2ehTAQDifuMB8jhnmIU6p5+8fVLV0rcDVp
h1jvTJ8i8arMIs61TM7KuYRoqQe8rsOauuGVWFmd5pLKOJI2XI5Jj0pbv9zG6ZykKXvjVfZ1yme7
p15ZOL8VTgnN2VeZyop468NpISZGUVkj9MB3m2p5zGyu0cU/Q6SHLcEnHJNMqczrS/MC0gGIbP8O
/gaWiyAkfyNnc9Zk8hJDJlxCAsyDEvas7edeD1EU9MR4zJRgtzq6LK/DV6ZLJ2J2zfY6gOXfAq4M
ibS04a7MiTLG+6TbVnIbPA9m0ejnoXdoCTsWLLwHCVBdGakvR0tRC7d95qEAsJFwtUewvHqBO4U7
GUHCuKFLHXQFKPODKOR3rHd4V9lcEnSy2NUgmBUrq7XxoayiOm2W8Em30pvJ2Z5SEY1epFrp50YR
L+B1Bdi3+XZzJBAx2WY9z9em88/Nx6GmAs79uNnweQ/G62ltNY/HkQPW9+FKvNuGDE71LyqinYFP
wMzVJCtHn7Qunx4h+8phbUgRVjpf8PK7sxqSSdS1xwSfHeCQ/Tex5H95GTBXNuJAwgEkOQfFVBbp
hDDcTCbnaNyrE6TW16Le6gOKn+bb73se2hknIDJyl8tT7+Gvd1N2VFLqo7Rm14NEhGT9SUDjO2T/
fd7yHBmPT+xcCwGUJMoU+tZEm+iSRb4wXSycI9/2sgK+MMNCh8EiSDLsKPA0Z+OUvj7sQxaKutZh
Zx/dV2iIWPj+404s74avyIecmb5kRmZWq0va4iQ85lP/QcNYQSnEO58Z1avrb2MsctH0OAASI3vz
/CPejvRyvka7Uv+zGpnhVpYKHNBmNTAWMgUp3ggt3P0NJjR1Wfejg6xRsnvp5gwyxNPHfc6DTJy+
Y35jNsALNc+Fi2MKyIGIo14cIdUxjnDOj63MfrC/6lJ+8+ZyMr2YkC5kA0f3DENsyWU2ivFF2f2I
KhB1Ro1Bp3IfZ4EGDm7PdqPeP1xxGI132Ki99RYj81Ax4lMzkxP6zB6DkcAOjuyqWkkROimt1uoE
vU4S3a0X24s+W7OA1aj86Tu80ulbC3SwzozfliLelA1ZLOot+njRZi28eDOY+xXTSG7M3UJFb0/T
bNm64bqWB3zIixbdYEj0tRwFdW9m4X0iOA7Sn37biqkbw0mXo+j3UrbS2SwHpzutJaDNRbNNMBql
DWgVeo/UjI8AS/S/sauhoweAKrVeD6YiqL90nJF4/iT8+nMdn5dTXej0F6s5Dz1RVjxee2KdSTDB
hxAIrvzxyGPgELj0KjgjfyDpdhfgQLZ1CUtGRc/KQhvlLhCpYym/51yH2NY5zNvQ11XPkhoaxjvC
vaKmX+Ou/VN2tlhO8sQOhMR6xJdaDtc9JEvEy3VCL2dj26D9lLbD99uHL+hylDdD44B/TFnZcRY2
2YeIN2vlfWsle58NaFRYMueJx62ESLzruplGJVpH5OF9NY1pwraDdUUNEb+ZsD6xn36kllOPifH9
9Dxm8cEZ9kWAjWuBFSIip1MH23WxaDFa/uVisFXRXyKGll1Qx4oVgXqsjEOPvQaf3Xhv4+xpnXPL
62JuEEbl7eU142v7xG/+ngBVzYqDkjYPwlpP8tRlGpYMjBvWbdQazi1wcqBL0E95nam3OC9bEadr
qPvCIh8OVR4gFSKdJmzTevoiEqOSnQbXjV2LE15I45qTrhFQaNVRBC0qHHJ+UAD4OR28WWofBfGc
I/tLunVUHD/g6uHl46aFxRPNV+/jpVZXitZbjOGsICpJ4t7SaW2A1OPAGm4nSUOmxgmDTzdBHMdA
I+CO5PPydqr8ybkFiRD0Sv3orJb8SlgnVU0YT4BpDpLVgV24iBQACjxXOOkAjPDzoFFL/i3+elVX
X2r0YBaFyQU0IFh4Lzlv+WZyuWXTnL5CN3xEq2uhzyZiKvgfOf+AaEZOs4aFbhqAA2FxQgjM9BIC
PqbmV6tu2Kk9djlf/NMt5oXghUbmBcFGXJzP5Qo64ooGreA3DvXX2fl/O9+EQ2LnGEwET6ObzHcO
ETf7Y1kx0MN018yZz5KYNua4pIM1x5tG9+7hRsjc1LkkNBjHm/iZaNLQNQsnooJl1ok7n64mODst
omKnfoBidQipHeT5FxdqVs276tLo5guxs/88DeClwlwemDqT5MTzUWkzbfhwA/JjesvuBUDbfkHl
2o/YZQf9V5r6dYsF4ebNNk830VkrO3ZWlELl8Xq2iQ1xN+WxHfpYAEbp1PbxP/IylMvXYbqRwoxb
1Qgo2iiscvOp5tvL03/Z081gwcuEANul/Jd7qBY0l3DxYsln5p580QmjhtBtqHysVJDdoTrgnVEy
dU8IrRUGx1yBohRtvsddpl+NS9lT4lXaAAwCTq65qpBZkSg8BT18u+IbWmaTU2i+40EFByInyVAH
UXi1IwxD8QoS5gTrlBrqd1KJIdV4yYeVYYZDczChhZcejxv2OQmjzxLFGWT2XaLpQZQnBuhbd00g
NiYmysSG30ifKg/gOrBloXnxh/EMnlJnSiQf1m40AVKVUgjJxfxzDZfO2uAWm68boCBWkYBC4eSe
21dGDBW3vkY+wDX+7S9y12u4aqJyvi2cOVctqJB54s9a7yTya9EXfKOPV5yEqKP7cTqs51RhAcFH
nxOVulQ0EQDU0bztxmnW+FmyXlDysx0ocOj/oCEd2NSpLlOD7YDqLaf7KJ1vOgR5Ld00JuHKVq6y
eSG/iytZ5ra5mcWsCO1QpWqwNbjKZtAzQBYww+G2RXb+us8WGjCJg8aJ59NdU8hur0s6o3gUDzCh
QmrkVr7bEizyB1eiZt++kOD6BhSr/WEnHPklURPHP8Og+s6lkx2K7mHBjPjHTBoVcqojlei4CjKk
w0f6Hbe5t38RwdmUMCO/YZCVtWnylkAdObOP+mXd9GTRunfvQS536uBSRPSzuWhUfQPWOfovvaDF
hx4dAAy1CzXpblTtEQzIeONR0O5H8xyDbIqRZ6UnuHR3NFdjYcMKHZml5/9UFMBsiC0ccL4hWwrR
PtYggRaoyJJi6pFkK2ibfNz96kWb0AER872+BMV6N2e7Pu1qi8XghVb7CTHSWHMGYsPmq28LO6Zj
hiGweTbem4L0KWYWrsI+U4RaIenDQLB3XRJRGi4paHZFWDqUXQOCkvOVY85/m0DFODhVpdrKZmDM
enXMVEcuMP7M5vSaDaUL/PIMVhCKppSnhcw5eIlJm3DPgSYtVTUIg4blPW2QT0jxNno7664D7fK1
ch2T+TE+KnbhtmZXnHQyFqt1r+3Gn04uWtYLzbbhhYYEqRMYKU53nOfBtRea9u6G0VRFKDMvn9ic
x57e35mBmqG8FPXb4ZPFF8OS9r018JevS8qKEWNsMQevm3Pzm9qtOoT7dwBYbpPsUv96WotGBFkj
oFs4osEacjaB7pWWRpg5hePShvCBCv7G59xzpkAngb4O9ryHUZckuyCPCIWUtGTMBqFogihV7Ye1
FbJ2c60s/pCw0rxCD5icgxUYbROnLsRapsji7vxGEXf27+RLpu4WJtUyF5DCE0CfAYMva0WHX1R5
IuOunG9D1wPl+I7Vz5wSZt9DFnTBaXkQpIvykA9NQnsYNgOPmPNtTIVaUbswV1tfJ83zzivv0Tu0
W9J2Jq06/jbylXjqwvKO4uQ4qfhFlabzaXPzEjTEsQILYSrhoAQylI4SCNaqZeQM5x6ii5IFo/B3
pDobtgfUJCKnkZVTVyPcjJx7Bym6cxUi5IlHlKyxRaNhAhsPZkmbOW+M7g0YqEFSexmcDkCOHUhi
a1jHKl9XnnlUwK1JiLLqboroyC/Fx55DQqs6S/FTGhjNU5+LXSmKo5ptqDUkhLDNSosmg9UdYP3N
8JH/aFShrw1YHV5+Qvw1z4f2wp9AvEjZp/a5U7Kvysj7YGQd5QbXweI5D14XNTkidEf2iZh0YcXl
iCT2Y58YggOTaVlURH9LPHJAphwLWGUcbHMIwh3UZwUa6BU43fpQsFCIAITu4h3aAPNGI2kMBWGq
JlV3sTIApHNNsWnowip0PaTPgU2Dtrm/QkPVsskDzTOFdx0UXcNKCBEpLiJ8IOEXTChIkFaUWXWD
u+n5rIzKivqWmiKtY5+LdDLI+BTreOLqaSKp8sL71sFE6/bJBfer/B1YLVaqTicN4b3QpihEgb3L
OTLL0NmT3v478qhZQijPbIIaUuNqfgIcAnFZyVAlJGuZTTYQg8lSkamT9rzBokXxmrNlPJxefpOk
FlGE2J16T4QEv2qzXDehoGp14yJItNl4rgiFMMo5bdMLIRBQDGw+xQgDS3WZ3MDOB/UsN8I9oKdf
TmgFni9G1n0Kv7JQfHh4Hla+ZMJXn7GfSOx0eJMRUFlD8UDCPnGFIssJe3bmsEAYX1SIRd3CDQTA
d7rZLodzaXd6mbF4jzk/5bcm0krpSIsayvtFx5Y45h9GZeN6ieC4OlmVkbq0yR5Lr83VYMH5Y+Wz
z3cR+44BNi6kd5RxaPHjmvm3udH0houYaOqpJlvPmBtam50iLJQt0RcnHVt1bmDTvTN9yBffbJCI
rBCUgBQEbd6yfKULza93Pyb5XtNh0GUw/lpclytoTGOkSPD2fge+Igiw4aFumd1PcgAHtwe83t8S
UEzZOIWtmRVqwIh4ksb90rkW1/ycgUR3i21zk8mY4hHvhXfazHpn4KZhBcPaFXVjgWFuxAv8f8nh
JR5sIUgFAeIS05RvAyKjxFbry41Ki89aRicqk+gdUmfCeWMiQ9q2lpnszgqWUgetwLBYKMwv/ig0
vDaO2UE1hBkjxhlgj6enusR0OHL0wBgHYyuoLOCF6qaq5AthYmpL4NDENrsSTNCpEYQi7ER544LI
R//ynVGnKBsHoQXNmPmLoiPzyUba2Ai5pauApcoB5TyWMKkK7OsSPKbn05u/oDJsqgQHlA9fvx0B
yVUqO9xQLkKr604BrMuZiyfA2rSQjGWL3MlwwFuXwIthbnNtC21lQk1s5GYxrWeTXW9X1uIeblfF
Dmee+Sc7MOwgdVIv9MPL1bsaXanFEjPqZUqZvhOeFhaOlQN0xqGGgwxNWBbLkXa2CSz/qD+WUtgs
aU9CVQHzSmZqQZ9aUVkf3YMzLDB0cJcG+tLlNABA34RoPyo0WiA7/NQgH0cLFnRybx+c52d0q3p+
3cRo7E88BV99Q2oIuhPIj/GxXuRVM2TpVCM+OR/46EpEJtVJ9CafICiCWThJmNw1QQf5FUtkLXRl
m4LLiFkNGPfDga2dQeQ4nNWjqo0hOJwsmoXCTCjDBPDwLjDb6g7z0A9y4w1f7v/iiaXfSiiPW1hB
D677Tu8BwZB4A0Hy9Ni/q9GEWjcLRVwNT+AO2F8VRAodit3SYWd/k6NcnJS4HJYdaVvmnHApVkHx
T5AFyFIGUQennOHCiyDktX6tyjsF1dnVwz2H9ZN7FfrPZRkHL7ShH2EyLFeILjKjTcHDEccmv53B
l7uIVbSy4KfXQ+j2RR2LwpVulzLEG5tmVTbUZQpH5TMVC/IHhweCTqWt6OWcOgW84DEFu/GStPpC
HrH4cNjc8y8EecxzwxBLw8wwLH18ESPoO9EmKX315Hh2hzgx4tiTYI55p9S85XNxp52C5+ei+Nrq
YJ8cMj88YvN8HYSb8rNz9ZksNX1y4Y6Zu53rdg6uHrjIVLGAQM4XNaycpCLkVtVSlOJea3MCAOrg
uDlWY8bmp064au7pKnp9GdXbeGPBFx+5ILEKGoVmnzRd5UGcqF+4EdbhAbMKC6M5jNkAhGF8fiUC
BTJpFqKIGPjSOZVZd4ydl8oqJiRXST9oT2UzQkE2FxsxeylbIb1s0BqtdPIAZhjR+J0NMwxH3gBt
/AqV4tbzyd6+NKyR576+fFKCUaAQOfH/+Lhkl8Dj5xsNm1pF5/sk10EzpIcVbZiNMMpuhbGehhdc
RbXodWMVI+aL4FTIlbncPSb6F8ldw2L+QWFvGrRuSkDmvB5QU58ctirpSlVWWIrTQyf2oPisA2X6
pzwhFWmOcQYh0fTFYuu2gg8SyqbKMZ4GRbUzTAl5xn2r1/O4AvCTIQ9BnoAOjDnI155ptnZtxw8q
7g56HjYBy1ecKR65W3Pbthxr+ffEDynnN+lQHuRK1hzo2h4PZGItx99A/QGropANuME0XPB6sJOV
0m/P7/ADEX8X30QmntNLWGo5EZwKCBpqkV48GqEe6gMQ0nHq6FcNJx8HpVivKPbzbluc3xkVesVH
1fnFjGSd4zq62K5RCWyWJXihrFvIYgfiECe02i9I0s1L8AZh61M6HnJm/i8fZ1eunM3SewjL/7hy
XA0G2z59+RFZ8wHNje0Dx4edXZ0W4xR1Tf5+EVdNRZG7IaiytfFWUCIkEBYc1wLUW+kjlfR3YVsR
NUIsfs6gZf0IONU3pYYfpe/h+rt74mrFiMBQEE4dlhvwS+DyxvteQIFzEJFVLGMjMApHisTa4TV5
+tNYcjR/tsVCkhBFncFxsyRAmtdtbWZxzYhEUQ1AXW1Q5szINf3ZlnHZFvDBzpWI99msmcbxquaH
ja7ayClhkKjU+y9HsBEgaJAfyp6gEJQ2/TOfn8RFlr69pRyz15QXKW+hvK7N/Tc7YtkPxDToqNAy
9w3yT8JECuNO9cNcXFr4NP1Wuk6aZUKIMVc2FJtNV+A690qlUVojXn7FA3BBNIWKYxKSCh+hbKr5
VMWlsf/tHg1V2uYdua8jNR9/mCFaud03Z8wB86dadEcH8Yzi7DBCG2ZpJQCcwX2o+Dk0zRXEGksA
SvO1bE4cERMCNy9ZfXGyyhx0XiHz1VQ732IpEMXIN76Lfc6/ZjNY+nbVmKnl+wXO8i53HwcnNPAX
byt/7A9eAwPmBAGfKOrkefSX4HFDADJSGU+6fd7YA43n/WQkRcUBtYDcffmIVFntr8wdCySFpYFe
wzdDH/gvf2eBO3qIlJLgXNBKvfAT3q14spMfBiXlUsKCfdGknd511ok1bMg8xjcUK48cB4n3wQ5H
AdOwy7O90LaM2S8IaNcCZwv36SJVITc6MwDnUzLdjEj8B6Cwf5WjADcnEyAyNRtovkbTZrDTVElG
8bJAt0z0V9K+MSWNEPf9UiagNqDgDd3T6mnSMiKhhgiM9k7F5kLUjmIdjsddFPYSvmWh25BfNnsA
nGaSbtH5YpAOS9s4i4/inMEtAlDsPze6tNJ69OnSpTxVe/SNPVZ8lAqY1/orJLuCYVJKpUXJJHee
hAST4HCWY35sd8U2nTcir90Bse4xMUOw+b1npL4kOAleedOtT3j9TpeSbRhxSDqNzgcDcyqnaXgr
OdKwo8q4S58zkDHZ+Yn5rzNmKACcX2GQdmcnMhVcwlCHmvZLE2k1XAGdYFQtOajIFT3ucoqoHnBn
k8i6q32zihg8KcYvC3GCJrhmlPpTkvz303LWc+29KRj6nbfZb4SFYhtSmoP9SyY08p5wOj0eAgQL
jjWVa+aY55bnmijd9g3oCacAVQkrdkveyBWyQaevhEkvDCzt5X/4q9qd8a0CQvBAD2giveE1uvPZ
48OlB2fVKl64hPFzNo+AriAfleT1MEt8VBgpabxhgLnmj915IC+U6IBIT/+qE+FYEpQYFX51wQDH
+bHc4rC9bzhMd9lMDVWJGOwa0t3y5oXGciKzJ2OQhioRYeMQE28GUDNsb6etc80IQEGsJSQUJLuD
5JPym7jvg2Dh9ObKuAL46bjdR+ElOPtvu0hqOAXJbF/vtVR4QOhLevyH97aiihY1Dc2SqCJzPH8x
WyZ7A7F4KQs+TCoPeZsJBdK7CRdNPRH797lkCEKY/SuHi5m5BYcE0qHQ8VZ9lP9FZEFiTKqWf3Cm
6tR840nf4lCbK0vvBV6UuJAjCheBdu3vXs0XXK4BiqM0RQq7d67LRD/Dl/tO3fABZsV7k9+5zMDi
3Q8zdkPnhTMZuyu+3Ck94Xwt2khe6KnCAoF9xoSFn+m/YcgeKjXZ2CcJ2uX3VW0dHp//0wQ3U2di
CEt6gTkFYsffC0O0LpJWUNT7ondO4+CNQgMc6ldhfiZAYxHOcJaizYr7RSCj5Rr1sX0FQQrY5h5s
88ax7WoOAP4VLPcIYAGNESsk4ax8WCLmGMdKjaanBmawvqOCR8V0jTJjqDDvwNV7cFpy4ryG1uNu
jAEfi1/npkp9Mt8WVfzC9hlUTz7IEpepw49n2QITYRCF90rGocUTDaMSKtr91ES70vBk+XK/Fjj6
nbqwi2xwNyKBBFGFILTARZHfjyw0j5+Q6WwiZFCBO55dlpDnz7pZplMmNJ216VW4rJt07VduY49w
RvW2EB6RLOrlRa8o9ZguY0yyziKqAQ4w/pWf+FyU3OsEHCYiK4eBBTao9nlh8N2rPM2mbW6d1+y+
eUklaI1vu4WKKgDT3OkxW1/KKB0Ou26vGX5aR1i2t5E61AlcbC6NZQ0GM+tMiWyNtDlZaXxsT7B0
Ye1wlhAlMguffYNztnhhieTfuOazKdtNB6QCcylAkwgpuJ6j+53ncWaHa+iun8jJqCU/gAVXD+8W
7zqxQnt/apEXKipMwnbf+u/hW12kxjydlc3UmBcO5g0PqkWqqPxwemwCGQHnBDklnffWbGf9R/zg
7JEmWNpHkHyVepBtCr32t82J4mqJOQ8IkvdDXHd+wO6ACiKtS8zr3mgPvzf8elhHc7XR2t+mqthk
mWS98ujyyVyinEesDKELD98HUJ/EOk60Iye9XOzxUjfDcbwuyD670ZomVnZ2xbyg8IbiC8WcNGvb
4T8GemAxFoTfMJgha6DrqlbdFmA+jR4yMidJluxPKUWq91xB8aANMOY8rM//EZlvrEsjisozvCNS
77zflkDSqZKMbBzaEne/JRGe6a6VF89WqztFuIMn4MpopaKBaSKnoUA5ZLVqSd4ouChL0C4amsPy
fzDzK4P5TYIbbN+VF53yjM8aDgo8qvF/pJg9VOkX/ENj1CrRRyZd4ZTwHUx7W2YHAgiUGq94VWcR
MVkW79NafQYfuuuSH0Rm/OYaRpnMCQ+foMb7aAKyjCQKViGNkXzTZ2C6fevrkNPetBk/RUUQBxSE
eNDwKlumf+aq99LmT/MN01XGdx6VFwd+E3AP2TaddC4hg24tbcfACHPyW7vqWlugn3HBbEfEu6KX
LSHQ4Ci9oaVE8lDE5tgHJocyUT1OBgNBsEK1cKTgqU1nbvwwlqe76mqyiBSolhit39Lgd0g9aFbz
JSubJF5euGaTBi1wVFso855cQS6DPP3XpbIbHdfCFtDSMQwg/O6EK7enwUgMmsiOh2kWkziTwYdu
D2MElQMm1IUruEX2tL6Ju5jc7QkkqjYHOrRcIHP7Awp9b//BnS/9zXyHTNCRtTA5LOcwHTQ/LLEa
jgax7zSidmE2xEm55/mPmwSZgbkLWx8Wq3wc8396I0rS5udFGtnZLATJhEJdaZ/Aol8a+uBRUSaE
eG7fq6rswwhpK9hcBDxKnbYhSZVnJtba5qndu2t6xJJd4rVlhr5O0dhLkbxV5QoVcNu03jmFd1sw
Hu/5Tve3/n099jEMwm0ja4sjX2aqXFKt8+VrcNwCZBflhIf/ZY9orFX1J9/b2pIhfjb6Sge4eiM6
rfDv177jDTAlUp4v5Uj87EPCcUog7S6F1/9MTQ9rrCVMm/n085tZD1IlABbCdLJdhYDinQylWr7M
irXj1fgxlp59hlW+SKU/j8wje7ZtmBSt9OXOe0SaFWrtZlvXCqlrRcxhc3Z+KzB8ccD16nwkNx/N
QrF3iHIIsJUtxduawJvDTmCGc6fzCyFKcbfXIldgSArhDtp7wJF1ZetUqo5mgNGPaxViSTdfoGzU
jaCG9Rq/Owz6esC7U0yxq+KhxhrDeKO1lUOriO1Q8RIKK95cDzF/0tVsN3ZMiiq6ihqfoYwFkkPN
iAXidkzCxLRsfC56wX0qWGREFdnjH4SW1eDEUtpkE3W1mAaS++tejCMp8+9pbi8aDuYQoMgZdBlr
ABQmGxt3n49FRXuMqltJvrp0gd8Ky/9nenZMSmUDhnlBm3sasEbEUxwJTQ1td7a9a3aGEJoCRE0T
yZFelQ2H+Ya/ZUaKDqrVTXGtLpTRxoO0Xmp48T3Powlyddfxz02aBfWH7Zt0zZmHRpqDIiNm2TmW
JL4ygdinsEOu0chIqzKopIgEU+bukO5Fc1n25uCGJWzc0kHVZiPLG8+jAkZNS5VFEtwUhAAqRP9E
oOd9TbrYKBWM0/2q0R0XTVJGajIqBuaPLegI6l+CfABBfKzFMINpGCoRP9R6V+uai+Y4wKmR3bWN
xBtF9bjyfl3xuzBI5aZRvvNTH8AGX3qW/uO81so5pfnJokWMgF7bzIvBWuwN+JjZ7BaUDDvJX5Hz
9WeXhG8OWIj6mPoEANK4F4CdFmnNowXZ/TC3++wBVa9RyXKotFhZQ76yrzx4CBX5LlfCKWVd1qXv
gBeg/amFtwK0LHOK0goC9nJTIAjEmW78dByOp2JJSq0H2vm2/QXumSx4El9+TytSm5V5slfCDcIT
hpHYOd6or9R+b5NFVhI1tFC2dQFuwWBCTTDKeAdm7SeUm3U3XHw1OqtxK+gLvC7MnMEnPF5r/JKj
FYkUincMIxdD+Sl/he6t9ruJM5r/fLooZM7ogLyj6aHFZkXpjRja/F71OJiml947xw8oPmXSj9D8
meTutO9ecvRcXsse3v8wR8iblr5StFnK9y7uMVh3nG7yRW8oipIaMtK1a/MdQjdeEtlefger3lIM
NvFEwyLw0dCEaP7iLQNuzAhroef3YHWStzVnHXL33iHifCGlcRD7Mrac3CCiGIqTTQDUNsUfNZWD
MqY7l/ZRHBvy2ylOif/LsUw++s2eenrA46zraXrwENMxKVVCHGeg90Erc6UEJLDecfZ9Q8l7JLJo
hb80Bn5EHU4nXKEFVf9KMz5GGF7hvZ+HGEgzZO99Hn9rEecX84CwS8aLjKnQTBxyI+oc+RQOQlZT
lKEnaD7QoqN0qSDOr8J7KH98Zkhep6ltjQ5BfSbnddgelO1QQvt9ljpclu6gXsOQ17rvRBKQqGXE
wu9nd6B4x4FnQH7OEbr7jDYHciCGyPz5lZ3CvmuL3iABKYHEA+Qe5+v4WyfafGekE+BxLMYXbSjm
aQmNdvC4bdLt0CI+7/P4GrZAZOJ61/QMSPdabMC/gU/ChGOch4ptdPgFS4zVIkYcJBGTNncu7b5P
psLXlYDwUYg0SEYwwPfnYfgn8RppnEIftG15zV3lC9Kfju6ZbN+92vK0ATw7dEQXATce0d/n5Wb1
OAA2NGAc7SHBAa9mKrtBqXpO/CJ6cebamcJdypZtnLIQbxfNmBu9fIJtCVLxDIGE+pHlsp/Tn0b6
T9ZFG+apq2z1CiKfIt6BEIsHYl8U+f6Ls8+QZB3ZDshs2MZZmPtOOU0e8SUxoMhIlhc1DyU+BwsM
2ljdFODED8bU4o+HOBWVuyKlh+I3OeyN84c15m5soF6RXeZjNt3Be7mt58Xp4tJlJMWC5wgLat7A
c4deK8mG/cve4KXGDWqoZNaRsNI+pOHbHOMuAVnIImS09d4jh153Y1Ns4tHjkpSrcYgjwH9z/qO1
ghi/H70QgWjJyAK6xLCzbw77vh1eVk5+C4qzgvzMR3hwjnSfmtwE48Bj/IuRZ6WptXWFGPV4e30t
XsghXTMBAEIAW1bsWRm6eYeIX0AB6e2rr0aZkpFpJGU3Bok9NfctDbI82AXdSJrnJWXhbpZNhp9C
xeQiOxTadyENlsESaiW/3PZNVMoCfDkzUIneFIEFfLxzH1BJi9QntAt6k/gugKP2KxXrY+7rIU9S
SibdX3qMHt/Czdyedi9hTIC3ZmzijkOhgJJQNZOW09N4QqC0Tu8UKKmQRCLm2KiwaqIyht3wmn9S
rYO/+GGiVw7G8ZiqnbXkep1W7fMlziffb6zAbY3LzOZb7BXQ0flv2KTo07bhmOZl5C89rjwWDeHl
lHwvh0Ymyr/MKt+rFLfmK73mdFaWLQ3C6o8qcn8mvNrix694UU25T+jvwF4ChSL0Zg1ww43ascjN
y5SF1Vsv6evCNMx/6qJ2HceHmDLCP7d5ka6tBEcZ6TuymUnRJPrVnxlc0Wee2EM/e0j2qEN7k5+N
F4Ni6/b5FWKGXB0O1IfmUXFcQMV9PRlUtG2tyu4IDzv+83FTgyiAUN5WSwn6lqIhCHTF/uwxD7oy
7VS06n3EXfWl0zUrMcDO/6vQnQth5d9a6uLuT+MspmPpFJEpufvpbIZ0f14neeHtGPIGMhRk7bSj
uSknqseI98pYmPg3S/9viJa8aDQ0hDUmRm9jh5mGVbwZ0t6s5/8kN74fD/pN3Wk6d80IQReVCDno
UAa1rTonSp9XKVbpJGBXvATD+ifWiXKxfqbjKemo1zQIJf19tqG4uHWdPLrp6o0Ft6pPSXddEcRR
00tc4+Zg/Pw+aUY1zSGwL6pVTry9invAzn1MkWTw4rzFK8TioMe4yznfOpu/sJGu8tLC9c3b+6Uc
PY8sA91kjth3k3uCrj7HCfz0HRec85fEJDV5WcGLfOBfQUiI5bw+ovmvJh8QUDetB0jzrVqc4fPp
iWC0dWTTDxj0GfcGkfcrR7D7/E5zrT9V6cle36GSKMaekY8lgTJNh27y+kmp8ImrjSN8Ro32YdOR
qRMgSnW6rJ7hTB/jnZURIw8CyxWT+HRAlOFbwXaLzHw/puMIT9ziJPAOc1FSQ0wZC0syOrG4MB8r
jVJuIz3L4uDa8bwrxbjPWKN3coCQ6Yh2vOg37CfEq5rOVc7zt+wCCPsF8mRcQ7+kYYsEWU3aOIRC
8LTCCHKpM5FMfl4oFYkNEyeoQr87kBTsFtVY1Ok34wuEpqlrWu0ot2wmDlVrGInJAOEClXtptbTL
QPr4ELdCFzxj51KTlUu0xzyV2zF6murpyn69FbCyQf5lhW6phxwJlOo/+2dQ2iy9p98JNvaXGYPa
PtvlcjRFir3QzaiQAX1TvU+sZtRE74MrlollqF4Ts+RJ6b14TGJeTxFg1iFcRJkQb9FoCRPDVM3Y
oUkXJZFLmfhvERbBsHJdL0gUQIYx0TJhV2K80N7C7wOYtBH/MdWXSw57LakQuVPd0mgoLK2naowR
eJWvVhYzLrY0ANdgKF9ekbEpO2Svjqt5L2ZQSGAp0auCnq09PUqXo8QOJe5O2Sax1s5LxmnNg4EE
P9gow4OUyYJURLRrrwLDLwlC6cKOB0Aoxg886ax+QKJJS59JFCoABQFkNG3CsYMrjZ6eSgBJjrbF
Fz0UkMH2ZtkgwNsshYLzgaT8VJXhHUQ8XbAojNsyDdkxrLaAj5rkxwN22AEn9JsAOEPwV8XeSkP0
TgypZ8056D1He6rdRb6ADtEKN86m88+ZHonJnA8rfs/1Z+LjJVdOnIN6bWlD/V3zd1z/VWY/iUwT
LWGJzx+FAWbQf2R8iomjJ/KxqzlzXBXnHv5edhMJ3TtRKi6v0Bu/rqHE/xD1yY+xKcyR0bTjug0S
q47886OJP51afuQ//+8kCy7e/gZe+POTiDiBvkG2pRrgug72dLB5ft8sy06mhqo3CgMdnmKlSeTd
UCl/QHOlAj5n7GpafC20JyTvZt9Uju+nXeLWCI+JneCiROmKgkRoFwEvtZTH0cg9ajyKxxV2AFaY
T4sX7xtslVlODs63pF34grqgBMgDw9zOM58ZO+1kIGzB+Kixlba2Oxc65xOzhi5oGiVNy0MnFBrl
4ny/uv7Kv+Bf/wCBF2zMgwFHHYUdpH2qQErWtJlrgWRFNNYQKVK/Fmv4Wg7mtBazuNzv+QJDnqmf
E8BakQnsEGSUCan6tPrXXv6AnBSROrMy9xtNYrPqyGDNZI9s7VkW/L4U1VVMAO+9pGpjhPmQ0FVj
FmB3/8VVBVeRyybRRUtxxvpNFtdUCa67UZPL3IG61MRtfQRuDfhOcY6UKdiyY0K9gy4qUt2iCuNr
OTRbrNsGISfzkTvvqCHBkZ9WUGyWzfcwtTkxOyGy5z65i1hWICIOY+7sa04Dbk2mzFhymyjuGJLv
I+1l65UQhlI0Y52NYHocbQYuiXigkROUylSi21fwc8wRDaA/WxauZ+0bldT5tOzL1g3ffIpfxfcS
dFKXbCMxlABybqRnUP4xjs29PzaTw2MmdMDO3ZMeBthJornYlrBapiQldsUW66RH+8QZq5KO5Hx7
nlREavMaqNfSCgndRkxQYkQlOnPne8zEbuldBshSS6DruWcstjxejrUkob6WUfUbGufYJS+Id+oK
8yT9bhauBc3laKjHPT/OqNUXEIWExYpoNdqQPKhxgKQNx9RHuAFpnPXvk99YSqhoNfeZzPGZoVpe
Og8LweHMlLgxXFNcX5KXW8rwL8AOBY33Q+KpXY6Tvh3LGS+ccaMhOZpav8NngAdCErzf6B7Usx0E
Ir6cKgQWXL6ayUhlBZ46kC1IiKiA8xjLTZj13q43HkJHbzAzNP+nLBhk8h2Ae9nCnvCRqopcmnh2
aBdYW48k7E3OBX7+kZp0FCikuf4aohashJOZfuRJrj+UrAZEXWozurrsyqslJ/eZL7MLmmuOTla/
AGjQr9lvRdmp0+//6rGsISOTT2simicBv7VZhJZiNDdIjrGfZb56L4bIvm5ZGYcG1uYi6WaFyJXL
IN/2REWlAt9nisBp31Z3BaUpgmX968lHd0Tavs7yi1UEyxUCW3BPFnui8i6QJW0yIotfWkuy1Yvy
XDbcNNqsyYse5/tY8hy21VtsROt90zbrYlmBVp+47FDx0oc72cQi07oy27g++gB0H6K/yeQ/2oGf
HkvMdlj4iYek8/wwGW7Om3IT6JZqNyB4DT3j+YfZ+zAA4xn1eQ2VJReQRfHNSFMqS22o/c6w1CNT
gZ6Sy+qIGZfQ4l5d0VAY23Y4C3DssTXglQjJyzFRfJPuQGlMOXcd/1Cid7yULg8ErJ4x+QtUpRNO
g1ebZpbQiqwPBajDNhILQu3kTtZqEo9TeHxT4utE17/d9t940p7Y7R0vQ23C5fN8+Bh5LvoECEKA
vz7gDBvZ3a6/JfU9/5XO7YvodDGUcfmIrkGcj5JRo0+qtj8xr4HB0+LxeqE3fUe+zcKZ5i0RXlR5
hPIz1BAdzZ5tRT6wKQoY4M9WAIiSmQIPf+ax9XUHGwj9lBAVfFooquWGJa/0dY8KrUsuG5CgOsBc
OpM3hztWV1fg8deCMm6TE4+OjN5quqaPSzHJmxmbXru8v4PaqgHZjNNzrVYrNT9swxWrJ5lfm+1y
+NZxik33NGR/BCFrGfRgdzViiv08Jm+UZH7cGaL0BaC/K8tAbXdvoDatZQ035It+WCWLi+8ePb0+
VF5N+7SogEeTgkxFGzDxEHdlugeiXHL0k430w1qurY+a3YZUdfqP1weC4cqOGBNDJGjTnowi3xt3
lBYoG9yqJmyV0p38Rsn5pwTN1u6xpVbWfJq+fGO7FKxlqwHX2/18JoEv7GxBiYoVHjfH04Belq+M
TY0Kwz5KGo7NNf7R3eeW3cPGvTFBAs4+CSlnQU3+BXZcinmlR2Ac3Cpgy6Upyo+X+Mq0U9fM1foS
kXwkYtRZSig8sDBL1fcpaGoh/IbbIbyWEgHJikSNSLoRKjTfNSPK/PA5j4WX2lgP52uYHl0PWwzX
QKZGilb0BzkV7VDKwb07SLYfJcT26AvEyydo4OxaWNKLcbukvtKDgNPXLaHCNGFbi0EAZQuZNqw0
q3/IKOCMFEOJvp625hB1CKM3gGB0L/snlknSWj3lY1WgsuO2p7wrErZMlpBnHQRRUfcjUnHOK6ph
clLbDlD+TsJluDDNxqRP/kRB4r70arza4WNanTY+0zXU7cV/KWAplY9zkWJWaDWZ1zC77Ji0cwnL
x19CwyTkT9lTUrT6r6jLskRwj+0K0K+ZfpG6gun83L9F1oQVJlxVn1os2/oeZjfQSDN8KMjAZvpV
5hEmuIWumeJ+UY2RpbP9Aiyp5OAkNenQwmpzSe/tUx5RRUBkjVvidX/B5HGCit4uiDXX/LhCjPFl
S9sBz21atEmKDidZMd8AcnmlyqY3UwGXXHTK9z2Tgru7rgR0sSxNQXtEchsUCjgwh9EFeH0+BEf7
3dPPitgFrjJ4Gm3J5B7rJPcisrrpftPmICdEPU5senJPrHpQgZWbMYA2yFQ0oovuLNbmtNV+ZWR2
E9t2NHadCS84r0A/VCLaXP6oAlDR8qSeibWijAnfWHMhqaZCy60jpO2U0BdnwwefrF/VWmloKNuo
IuRYmB8afJxUCisKuY5boDtNdLk31sdeObdDjInptM6OEsluF7RIDD9mEUMHwPu9N+l3GsRsSEV7
o5HOCmyfCC/76s9ejXHJZaViRIj8pVwPm88J2pAWc1NGFx73B8TJkNwLfGCyTW9xWTmhUzWdWyE4
sTJDmDyc/01+xLO2uKa8qntiMWQjbEOe8CIu8AapoQorZejN3lyYiPLKp2l9FZFiltVJuUtEc3xl
2IzXZSmoCEznnzzsfI+/b21SCWXciJ6meey/jMzNrcv0HD7C2mcHlxpE5A7iUfOTkKem2sOaDjaG
lY9EjQVjd3W7ZknM76qVfU6Fnfkv0xCYXE3IjPDLu8rx0MhIQQNyY0KmzNYZgQeWyq5MD+hEK6TW
2Z1j1+bMFqVTVd8SMiZqri+gWUHYw8jY/0bbqF/6Q1Ke/XtEzyMhiq8/Mk8w1+x+Upwu5RhfJle4
F6XJvCKw9VpnihHhawNv+httXE331afp71j6nRsrWjjgBdwI3gw1QoGXwUpA8yRTatLuEXiG5L3V
70zpNr/wy8uL7bf5aw5ztYQXHQdhgMXPXB7At3Wng50VNwpm8L49QFa3h2DgwJWEN/V3ysUiby9K
YAP46jRMFUJE0Yn0vwpj/HorkIcBqyau95IRbcpGuuLu/56O4tDZGm3/tHvFVSP6uU/ChNUUz53I
zGF63RjKvUtCgYxAoCBO7C8b9j1SoSc/KNqlK6e1rtVrjfxjoYiMkEGEgPlkInqbYh1v5MLhhS0c
eMcOE2iTFq8HZlCzahQxyLarG2tpjyj/e5EUSzKNmDRkzZvWzLwpPOS5R+BEMBvIArBL0e6XQO3G
uYheSo4J0y16AeTLnv5fpEYOEeUAc0dFqKDsrf6JZTa8mrm1BLQzkZiiSOLG54/Jze/1HAOWI3kZ
7SsqvecKvssyPJgGRH36d4LkSELT0wdjb5XDXHuywN20IGYwrlz7Z7dl/OUt8fThq+6hqdeSjrcM
5JRNPpxSiJYCawbDpjbNed9YG0D0wk2Hz0V40aKieen7LnLrRrnS3/iQAHEFrCzkkzpAAH7Vsm/3
BGZFoWihJ3yErhLJSCESxzqdDpwbB+SDjov25eXKrD/4zVmV3RJHk/sOBYZGPtElUTCdnW1GFyRZ
YsW/SRfdjHWXmbWMSruZgpiqQDd1OnJIIFk2zDRQNknUueFvmd9xRcCToxxtsO/pm0FN4NiKr9O+
o2W9qRn+JSTfgsdzk2pB87cQoB4DgS7cLJoPFdF2cKPPySnWUnr/y5Kd0kqFLhsNGoM5jeMar7d7
4KUJnERKxRzt4mmW6zcyG2SpbTjvG8f1d7GMkOKQ36FV5FzSmCW7ECZ0S3pWKvrh8577EzZLdGfu
cLC01VOEM0jFhZC7I3XfEcb1BdhSyEBu02uAF36MAv6kksq8eo7FoOIcj3vJW9HiCXH0oxbzLqDP
9fHpiY+nOe7V0ZWBkeyxQqGwNxjOZwNpzVeKVkfVuYdt7FamUsC/JGzVx52pYkwX5OgxYNpOWjPH
wyMmc7xkzEDZliDPYcMtvBMHg0sBSsLnH7gM5UPw/0Hd7pfjxUIJuG0yBW4AxY+dJ4eijzjMhPYB
35ko/aiqvVhfueWzmI1tNEBdCU7vvSR/ggpTc4+R9dpMHXHJmqeKhyh3t75/h/+gthMmaPNnLltN
+QtcveGy2Ta7CsOb7vM1env2RH044MSgWYA8UFCYtybNn5kcJQa7H0rNiU2bZOhdSBWG2rTrcHG1
K08p6z5KboCS9Tl4lFnrunw8bsgaQz08Onk9ol6Zq/0U26DKfnrzgin8MbnUzDygdqj9CugmdVqh
Vlx3Bb9589fBxYtHXx+7DCstTP2IXeVgsT/b14JKaBONIg7paPbGiT6vnN272hGWndM19CVwWFcR
iLTVFvWGidqzwEWmQ0QIPvM7+1G6fdw98C+4kWeWSjpncYa+JDBJNJRc+8Yb4oyUGUVb0aN7O/xV
nfygNVXjVfra9loUmqboLY4muySXmIIHERbqO79hTmRsEImq+4GlmNW7U6qAmpTUe6RTndgRs37T
0GcBK5bhHNf3NrjJQ00nbl73yx4aBX/z2Qp8l3usL/ouKPAWgH3PtL/nMs76Ccs0KR/rFTIfvOVO
0OC/6mfV48mMz914bnjMhHOOHbyGy60f+4LldENHESx40p+RvNOV5u1zKka2TkfEPEaccoFtvVYa
uC6AckNgeiC7MItJUdb+1aEfGejQIjkLMHvwTyEGnNe1eLZfrzPQjT7JWC54VXubAdWLJJOawT1h
3C7U+GzspjrYICveLgmcO0ltVIBhvXzwno7JUguSPCxc7hfeFxJr/a+gqcUwes/JPcGr9U1366/2
G31gVHnow6DnucvrLOV1C98ScCZXgyhJ/X5kKpn5CG0YLnxaod6nvHQuRF06aiKOwBx6x5KbZ5fA
3ErFFksCjPDbQ1iVpcZKXPUROPNCaNZuv8eIYRb5unFSBx6KXoGmv12A0gcFKIqbTgcf6HJtt+i5
Aj4UR0K8BozLB4b+kc8KG4lycMKx3PJiukCtjgm5QMdITrxkno6NP9s2eLAYHEs30T+ZAU63TP8y
X3E2XUFlCFXycNbDtKs81iRVlBD1nWQoK/FghlcOoPFfEqGJu1bSLL8Qfj9vn1dSsmNDx7Kgb/92
kF+Uj/3/aNIA5pz/qYLCW+QrwRgSwvXAUyvToXtEfMWkPGmIBvXI2XxY0BeIkhTC5zZzsBMFRwUj
xa/GdTcNp1P2qX5M4yrF9s8lFik9c4zsnDSKwf2KOF4zp0m/Rha31vMIJH1lACBsmQp5Ep6iK+Q1
me2+64LOOO+L4JLM4CFy5jmG8Ql0MT1adSn7A/b3d8sZlit0o7n/E6gx1xxgD3PZD16J1rWAP6ve
WrpRDGrtjuEnTxfzHjj9qoz7HUkj6yneyIzZII3lQVVvPa5owa9HfT/pnODPGhp2MRO7XgxVxwaR
vtr2caY82K0HGTXqOWHjUNZF+FkUDaaS7rYcOspowf7HbS93DmfX/GpxzYSb1fYSgVrQGaNlfUT9
lyzfNcDigaodHNRDe7Hsd08vyNrxJY1oNGlpsYCqVS0YyvNvf08KGFYPmnTqiibFlaw+e3/HRPQ0
WoqoiXzH8YDTwUyicVoylO5ISELzj7WAnTKGubq6w9UFCzds07gY8t256cw8uTODEHu6Qn1miZfL
+5yRr/EJcf0SaOFTWcWw+6VrciwmyA3TcrIHQTg8qigwNXHWhzF5aLViuZWSGrTn4RVUljaKn1uY
rOd/T1sEl92C/Qw0BF4XjVRklzgDDacg17TT7YyB6W04AhjgFdpMX0qHoae3fCGlTjW6Op+dhZgu
oyBCMDtOpjowvNyU/43SAU4XqHbZ9XwhunpipcmaDOPnJLwDRMf9nzUaFWYmj2rOvZu423CZaEZJ
qNQf4srBVPj1czVn07ruXkhwONoCXDIwJJgh2vgHjiJ+9pQMXVvV4t9y5hvj2u0JrOTNohs+Igul
/W0MQJKl1kd6+falCQ2CJOtqUhLM7pVLOM/ORX7Ce2IY+2xdm4jLhif7ug5fKAFOaOnjrsLgxDve
rIWWkfUlIxZJo75On72GqFKxHpMiFwECMWx2Ms6LgjEa8OEP2A3NWtAVwjGDc6ZR7rLV56u6+jOZ
9891F4L1dqts2C/7FK1M2mNqBHJraX7uuYLsAKykKwbJZVG8uQghrwWB/IuMzztV0oiSKJPszYQ9
KS5jVdyYNzpGHCmjKRykJ/InhRWAQX5RNsVn+6n5rBZTDNKoGmN9nLjNFcHzxBZO7C2hGkTpPah/
qlCyuh1Ct9fGaV+5Rr6kfzjj+ESFVduAEJ2YJH/LlaPZzE5qThiPPeFERLH5QSJXA+a+bB8vHvpy
IA5TXJsWLUV6NSRuyQv7fzpLGXLxDuCL1u5QSKOk1YFTJNYaHduSEMBs5ZRy5iM/WAK2HpdyQRwD
ICsAleD760e+Y5ux7cAqJ5znin7m4sb4FMMk+wTh7UUc1Xo58hTU6Jc0e7E05hn2VXA1EwA1WzxO
tah6fiqwK4VvRd79iZsd7OdWY5v0JV/HFsxKr2PoWVvPP7tMaKwjdEjcAgCADOhh0GgZ6nAzOfWr
y2h4PIRJf9gToDapaGs3ovX4uTjG6JSzVbBetvyhj7qrYpCCkpw/imapOnpzX9Fb5B6KxzGPdc/F
LkpnIJ0nWfP+9bxV7Txhkkb/4XHNqox7a5loEbzNMeUeQ/SCh+pbbkIgzZdF4arUmI+aj7iYLEUw
KcyvWNyuATMbHcgUBxKTig8xxe7lvxYzy7+V+zTl+82bsUaVI8/MjkbAFpXJGmhyUycSZrtdRmdp
P2g645DCmqXFW0WWllbaZzlZ2GzF8TVnA8MFK2kCCeRYtbKmHEt/vJSOOfUFpbZ2lJXn+OMKW+/k
z7NjXCYzabeycvAJq8EKGuVgzfGs2XcOEEskdL6j4KyKnNsRv1b9eK6d7g5yDEEN9w5cctmAv9vg
FGwiTVI4uLbLWEIrlhOUsjhmpUstgyxSqGRZwLNa6s8cxBFlwC7sXeApPld1ngW28+55JXW267r7
GVkpAkY3bQlBxo4onWfZYLFN15lWWeMx9b1MbRNL85P8y6ggJvVke+M62cfPPlxba61PMkPrBcWo
aARovlYfbaN5W0JfTpdh54fySbypDNxDo2kqc55PSEJ/QJnKDQ53UogcbojR11b2RINw1AlUpXEn
B//aNHKDG+AWgktd9K4avDyne0IObVWKPBnburTi80rd6YFz+NnButIQFwhbdqVhquHiXJIUPgXv
jwWsJYbFZg++b+Sernh8oM2V6UtkRQz/no5L6G+RhWVQMhz1fvpVv3h6/DHPy298y8e5ZVRi6Qoc
dXRUq6bC+0xTl0MJObyyD1aeN4WQW8t9Z5sdn3bL9KoFHV+cqTc8PDB94cLueJR8zrRArM2lj8Pu
FyWjpGWzG+UNxdOU7iKsg/L/7fM4PU9RjwkWdcICwSX0B6L6sdRit0BzM1mrUIz77mY6ir6hCDb/
JfoDSQukG7kOchL1iZyJbA5yRZWeC41HUUT09TRjl8adJw0atQGwJ4YLCOujIstdMc/QEvfbeZpZ
ZMT2a3t12jTDfUeo9f2tGSCvNCxDcf3qpIpLrwdwxjraqZ+wtcDDQLXmkLktXXCnBuRJCnh6t6da
gH/meXL4PGyqvUKciwx36497gb1NbiarsRq9tY3pZs0ZmUzzmj5t6gBviklw64JAhEPAAhMfP5am
FeeKy8rJUjDzvYyrfgDR5yGcfPI22s8WWQDcjOHwkHvhEzn5Tvil0mLgLMS3v01m9s9bshlpTF8C
8QMdmBlpg7Hhdos6Dby8fzcjEepWwgJ/26FzJwIr28aScniXpnBNQPr8IFAv3EmxIOGWsd/9OPJR
yq2DQk83gmDZhCaTUb4/d6mRjHHuexSwJo2MiAa1SEi1WJCSHnoye7FENOILiK7gfJZffYKmHXss
3hXMo1TCKxvZKDnCNeLMZz1euTpyRmPrtX0Jnaz3NfVdJBeMj7UlbDUl7+zPramWbjGhduROCr+M
knYgEYql88MVmWdMrDMth2ODpyBm0R6/CrcVGdl5O2sL9RpfQB6vo3KKGqXG7hydd6r8EkJdWcPd
Of2h8vM4TbXKj7V2EhliFkX3KufEQfK2p0h/eSaTE5mbb6aoH1Vaf3+I2QufgFJViqhdU/hxmzXl
LZZGk+V0uZFc/081BcOmZ/POTPRrGaxynJqtUXV2DGv6n6ujyvVGhwpdH4PGcBB3Z+nQ0jHwyucD
FdNYuDc8MIuw6k0w70K3eqCAjnUVsC4uDlj5zPQzXBg2B7iHH/OcMYT2jDlF5sGluInSqmLCjeVA
yJ6GIdB487WiYOElDprtRR5zj0OEMwy/RuX4QeiQHSQobmrXNw6uyN46/wCfpPM6i8+iwf3nfdAA
7w118s1z6O4y6W24PDE9JyoQ30BlUtcP5kJ74s7N0hMPa41JdFUS8tXzQAG9NrsKDYiqKAG/QUq0
FN/5aOrXbfQsLOXo8HsA+pNkVvkP/REuo+z8DtYifPrgJHkmyiGFQZUFgm/OAtEJm9Mcaho+FJpN
pphPdLTBz0e/poZp6hO0ot5eR6PA5Pc2mjUL/NfJS89zEtBfmhmAPQrg92ftRpue02YDKZgwsQGu
XFnw9gjXK+oSk9YOxHBVsFFnObR6hsYjtHNVogUHMo9hWn4Ow6pdy1ZkV7Boc9aaFN5mUjcYHaaw
IDwyXzhfQhNksQwNw2E5XII2jKL14phMaDVULVPrOjQEY7VW0NiByMS5tc0afwU6K6igTgGxLMyG
hwykSMzLGQB4RPkV2XBbmKhdi2TNRS8rijOK8NjupaPZqxC+aoh9HvB5vUya7m2LoDsqzc94YOZm
NlmkJMMilciWhRPvF5Fekxf/Myc7D82pT3uDX5c17aaJmo+uVdmrmjSBiFQMg14nFT21y2p/zRr/
3gYY3Rm5Nsh4akHB9Yjuw+oCnlAbWM7GEbM95itFTgHhRhmANiL098g8Sg0R9CaDF09xMZIKK8NT
caDhsPpvGwBVethQr6/w/zVLfyjAeY1bv5V616vn9qX7LIw0poLhN7oZwSMgmFZxDOnXLMt3Kd9j
IZsQ1Nm6jjiMwKoQgIOllABL+duon/GGWXqBTIARcG9Az5WW2v2uSYSRFCDjh53lKd0f4OqKggZp
XmpfjT/jVbh2S+WR7CqH8FDWpbp1rlxhGiRMjDXxdHfSNksSPhooLMsCUlPYRZaa644GnxVn/du4
MLhf/vXYIDrPbSXcn2lyHKTSr2onzIpoe/kuLxp74+xO5M2pZ1gCHM9kvMC4h6DqId74SxtK1kGw
4vZGMuQHr3NloWE32S7kfjzz0Sm5rmv2PdPzCwU30sICjleBMdpxMmbVTcqEIxS/w0axLVuuFZgI
klWA9S8SeeXrSTN+HCjNQwdSEdKVA8t+TGmka1eUKU0+ZPGaG+8ildjsYJhjUh84FDrlbPTlORNs
XJzhc+OQb32EoqaJGE5mjiaU+nAj6K9y78oCN+tTfBa0ZAKfGx0mZFx5weSjVFZHCqCp6nISB51z
m9iIS7IraRKupQen7PGYrXYtlfD+qTkfm1JjbS0tm4ewuw67J0MMBRxC9qMpDHZzyW4nyORRBntA
OTN1F1SYXW60D+QN3sR5O2aX0KvV5xIruka6t6koWihmFQapOeGu6/wCnlAi/CQIpTQibACPVJq/
gOFxC4YK0frxUQdJWXNbcek5QiUuCNAa7wAU2VQT6pd4YTz8azpQFJ5aezoRa7AVnxhJ18s0NAow
MmGUhxUENVcLRcYGar4y0T+i2qc2owVETi7lFe33BOLIq0KVt1601pTMPkasGX74mGzvJw9P3OIU
1xXgumZl5tTrJjKZToCjAW1cPdHW0VXOiVZ7QKBghqilc7gWOz2UzfT1Ha5gmmvLzPK1650KloO1
zX7acLchtLOm8oe5BXrn7Bq6WOkHKsfUhSZerC93cicgnUyS4Yqk2Mobqo3Skvmv253c9gvFT1A7
9qaOCpsuEWtjyfye7JgxB9OcEHpUNxoJKAdn468XFETlc+jFUg3aWki0gHOUl0Li8PZxseYVIaZ5
A711gsjvzc7X7FjpfdvX4RB/aUNL1u9jH15eD8063V44e5s1uC4Hfx5uF/QVEnbBIf7xMLHXGoyB
L73932s1HdsRQ/MqyFAwM1q/+Xrx2aGRjYYKhZwg4d592m/Hr1CpmJHcucX9t+uBwojfHU1GcduQ
5xA9KZw3KOUtf/bJgqJSed8IwkfnGdByPcwEmReS/kFRWv9LyJ6C5N7vjzt1NT1ZZkkM6CjXQ6gm
JXySlD93Hw/s3RDZjFZ9JYcq68EhzIwOZiwmo6cQRlR2y0Zh5taw0+0XiEjZvs+voCa93sex/Q+i
4AZjK54kDvOKm5XDw/ax+RU9B3Sn5f6xi11eMxne9Y5sgU73SfdSx4KlJ/1KlRmpPC2VFg8Eo0KR
r39mjZqbnArAV51zQUKvxI+GTIrpzZyy2V1eDlClakNQ/OaZDhuqG3LJzfwrqIImU0R96peLIWhE
zvElzrUuabxESHw2IqyzH1jRk4D0clssQ3YBAPdBHGgk1IIrn2wWXoW35RK+oK3BjdCV1D3+dS8u
iu3UdMoKTzQJCGw16qPBtq7IOCKVRzIYvYoBOHU3tn7YRNF/tUPMUS1lNPdDQ26UvP5cHpeZTYhO
6/IXrtyrY+PYNHn5FMc+Ozjix/4l2TElVoTDCtbjv+oVt78xmE37a5JK+7/Is9JQgtKFx3O/iORX
vf6Fd7uDw2xq2z8hlPO3aPsURRx7oheBn5ETjqFbKrYOiPYZmCP8yNg2cbp2zQO8JKt1Y7rYkwGf
+tKvt3/vLmTWxKDyBWFf5YhCdpyn++pWKlkjnSPPq2ti018n/9ZAyg/+ukaHjdx8z2Z77Ane9xVJ
WMBNcUrdyTJEkUFwfIw347U3NojvJc7QQTrmhj0rJWUSycV9yPKzz3ipY6wlC9YxSHgrK8XHjbB4
jQ40NZ/MXxO2abyoPx1GfGZj8qmn5p5cj3XnM+3Rwa8wjIyxM+EGAuETRmKxMuxnVQoQtYHWAlCr
Gd6HX6lZkhCi0vOL67+Nj3CizK8SjWjMvJ87U93caNSMReKJvZD0er58VqBBWv2PHbBc72bt0IMV
6pnloq0lKt7UaUOgCus2bNdLIYiLCCZf+bx6DGVVh3EcM1IwkD2DxOmgtPVDQBmL547FXNwjo8dX
IOEt3rt9Zn544h8U322QqUFLuE/CRxOHYxseVUD+uLGdZbjbJbhq9hJCxvUXmr+Xe7jNj+oQP3AC
8H5S4F3+SVQgu4PaZODtNwIfreTaxoiw/mCznqKm0XVe/lqswuMLQwf47tjc3l14QfzcqRITHyvd
Fm4HHAcZWV3Myua/FE35e94yAgcLyUUr7SS0lacDVwwBJmdIvZtURzAwWHewpmhWPwIKn+d4kC8j
5lstjIRkYarsSOp08847RHI1MXeK3D/3KK/Z9aK1svdewDHzXE/p4XCBbGDSK/pLIUvXF6kUp6SQ
SiLwL7NulFHKBrFJI9yYRiX6X/BVPGCoWcV1ueevbVu/tMpiKfVM0p5RPRSq4t1X+SJFr1xLCX1B
dm1ooa27c8bYWshA1LHuG62zYfOik8asI76eil5utYBDdKlADIgTwUgFYeaczYUUi2/8gfwFHbaA
5BXQrKQymS6p/zqQSFswGKuTqR8iRoVYMaMsP3N+DIlOL2smYE+sO/2enNFtiy75qtLh/QfTsoKi
OKYFcB+VJxoHvAkujs/qDWQyLPOikEg85ATf2mHv6fjIZ64yyWZRXxaTlsE2Y4/Q5J3hhPOQTHc1
V+G/E4g1Ee9c8x64V+vsqyr0dPRBobgtGXKETDp1jZSX9RdsgsV/0OtV+/asnYwlJKZRrGwaNlJF
RpycLUdx/DvDhWLls77bsNuZ3Sa4p5uDcsHObQ0agkS4lGoUG/xRHSgBLChM83XFMuLbqyBRFgQ9
6jomQxZbYDwGtf52cEU6c7d2zeguk4i2Qo9WlSsmMioq0on8oFAESXOE4uW4Goimx/6p7/wNUelV
aZSkX+kZa60jKa2cz69gMN710yX88WspUmLse+xPdC+DjNqM9g70/1uC6AUO2vrPm+FD/itj4IGc
4nL3myPARyghC9PWJgpLCLUwHfSyxxqHviHB+OIvVeg2e6U/e/G1POOoZYL9+3dvwL1WoG+20t78
rU71RZL4jVvwjNyAKEDekv2ZHMzRkSemhfDF4HipI7PnSdWldY7RysQu4JsjELoiPGnByINkJQ97
3k9OUzliaVyPBop2YQFzL/mNsOoFPItJQjdys8EkPVXJIgJDKFQgdW7oUDpak4dakenTEyPG/F/j
k3D9YxZwUAwy1tU/7LmqO9sUoAue9CgdsuKGmi10XdTlV4AtiIJDc2exU6UzA1YKSsyNAYaSVI11
FB6H1LkvGgZdgU11QWc0hhVz0xB4r4wQf+9XrIezVvDWdb8g4WATDxlxZTHk/k1gF98ds8TyHNaE
mbSSarOHJfZyUJqiEcBOZLP6zLrCwGHQNAhoXCs7Kd7vi9QoIOXbyBUPofVjywRAatl2q+R4Fjd0
LR5EzGFbEbJolZ+4qUojQOrFrGN6pfCn9xdA69FtOQLKLmYlvva2qbynze9mErin+myy4CSxlI8d
QMIgjHqjoRGOoU2Av8v7qi0o9LYKQV+JyowIJazRoSCTgKpvpxYhO7o67oJZo4pqr+FNJhmZR5sE
qmK9Jc3Ig0a/xjkFx0PQ8lRkRFaMFLUHyr2eWnEnPV/aOILJZklX2YQypT5zYEVG9NKyuFUVZTdX
xe+IvD5DufhdUt3tjiFYYgbHVumsqP9LReyRPfQhmnw86vvsM/DUSqcWYteC+vXGFTV4Ey1Ovs9x
37XDfunZchqq1dEvHC4h8X76IkdRwkp5QFYd+1aCxi81+ClCVvu2WmRE6xu4Xq9AHJJeBntbfWYc
k2v+1uMZeCW1qYOwuuv1Yhip8xSuabX2LbbZLy2+vf7dd+yQmDQNc2Pgs8yLk2XSq5otFBctJjDv
6yRCZdadAyV0oSp31ihZnWGyEtkhNe/qaPnZTh1vVwTFlTC9XOORhU2GnRDWpzWRBwufsdWD8+nZ
1fyFUlIU4sGebHvG3Xme1duqBJnp58edqC6jyq79jTjC6Hb4PrI1phTgMEji5rcH2AddzJFhYotE
XTwaQ9c54sD9wkRBg1wTL+qCXpiSjHiwGn1UCzUhYM/GsaC1Yn0I+nD85LPtABgFV++I0PzinTSK
OKfCBkaOouHMXUwmSWEkquMX2eJw/RpJejTA5eGvJnftSzzecqSm9+C+oH5aiOb9xrGVAheQey0a
kKVW4y0iqSdnuHI9Uo41tYzJdVBIYurivt/4ekkyuDvjOmujT51xNLX38cZEWNJjAkKO6dU0avxQ
5KFW1exuiRHi2rrOZmEY3OhufDEBTab65hZ5VybUB9wTAOJDe2uMri18SRL2kJBWvMcsaO62coWY
hRhrNA9r49kCPxXW/axOpado5QaTRHernxF2iM65Hxdcffj4LkFYyRXptMG74z1AFhY7oFBiX0LG
xGexKcwH5T6sliVJGnaG4unNFbFtBjbyVNLSOs7Li0++n2j1OOpNJcQ3BaIGz2hz9RHsT2NWrgLV
611BzoS9k0599eOnlXZKnkh5c3SB6gMifr7YqTPob+wihL7nyOfUGnNHT+zlxPRBaLsuB+1K0o7N
TwLUM7DOpOHyED/9uJc7TpEI9p3o5E9lMWrMdIaPOzoWlzCUMOZc2d4H7odsFcLmw9XR0rwLmB/a
2kWftqRu2feAOwIJfdEluxP1VWqL86p7vfpVo68Rdy6twMzXk1+xDWPcjtCZbpBaNKfbZVDmSICh
yFJUIGA8lEORgkMPsHJWJGA3CGfI2Ow0b6EIBrZcbCHf3XU241OVuDhcUFRR/6prVFMxKnxTlUGh
/Ttvyq8GlS3yKaDT2lWANdaF90zKLrdWMtdOwWVPerRNRHW7i2PVV1v30E74WjnuKQCMGSoQNvBv
sK6czoN1LB4AbTcKzCD9q1mRck0vBekD3MgXsB17ewPpQHdg4UFGiVjLEkn74RP09MCH0CUd/a4p
6YOAJZ6Fk03VF/jgrN0vDiDHMsogDDfJt/9Trak7xYTdpnTI6wKu/NlOI9DVpkihqPPpCyknvI4g
UUHyOZw9YvvTEm+RQ5M606LGc24bnZpmPHX8gxERhDUu/AHp43P44W695BhXBhN3NFKZaXky7hFH
6aFdmZMWR8Y52fbDTYOeR5C959/w3MZht66AFWJlWkQf6F4OEHY0nieJxGkTY+lW3xoYux7krezn
THencRbl/tm+nySsQ0GKY5Cm4CryZCysxPW+SmR3V1h5X5/eTzyDH84nBp/507nWt2sf7YjzD7sc
6/xob2PYItua5qEsRGPJfC50syKv11DxxGeoIA9sggsm70HzDvvTnbSlrcCvP3HY3W1o2sMLLGEn
hxxyu/BegZUN6NdrWF+zdFR/sX5NgBqTbJvVrs9Q5S8ayqB8Sd1HxRE7y7MreyzSff/hRaFRzc/c
1yRbnBTtIQm/l3E44w+Tb66qTy9Y34V5TvLvYGrxzwsXTMAEw7idPjsZr+cqjTicvzfbpK8sRcFF
N3IAnCmv+ZWhq5mr4nqRtP9wctOt+x4r3baiphNO3CS270oVTFTjdTPAWhJKDiH09u37eRjzbi/X
syAY9c4W54swploy8iPyqAV0Xw8mZG94Q82ZBdtklVAOExbnNVJb0wEKHHiW5pVmCfGmGnhPcIGC
bCRO9TTOM8b0DWT2riMwEP5ArIk+Dlw1Jrs58IVRCp8U1wOordYteuBo4wVAT9jNMyQHqiygu7nV
o0ET8rR9xohc/bfqUwXxBC9tm2h82TW39jx96+jI5zEe18VhWeEujAJSJ9fA+URdUohQ9FA1tX3N
7S+ZE1bNVMQL1vUpEDDMz6+KGS1F0gSwtiEYM8aRlz5f45w+/VcBnuD9i12H3nKAojhiR5oILDyh
yJh7AloVIAGNTT1T3D4ba/fTmqGJWg6qGKtp9vSAJF/Y2FBjZPHYmAbNSUMERi4o+vMRT2P4Esk6
5TcDGHGnnTfDCXT2/5yR3mvQ3CK5wawU+AOOsGgwCf0sJ2nDkkCub+yEeLLKR9jE5XuDoe0KnUvR
8aUpAfGcZ6WkRu7M1b+agHvD9lU7vUIAmk9NBeLT2LFmHz4I8iyywUOeogjCV34vnH1/kHJTBKzY
zsveCwtz6EeHoyTG33fEaJwOD2ioK8m7eqzCxULZeO7nq8Qb/HrEpOeRndXHO7gTcXaa2E281odg
uCRBe5j+hEFu9IfyCEc2VegliKGY3NjFSeiobx7WcIRlkmdrREtlZpzdmEE53G2G+cbwshUxyBCz
9JZGC3wpyvR2mGGKzuxhF4/CLYqgLXh9EDWgw7dy7YCbhdRj24cGuuhfs0TzGNVyBZ7UFXWXeSmx
dcJ5Qqs5/BgAxo47n840hxNUXFabuybvz+BPj3VGJH84wjLYP1L7SCka9hEg8BhvqW6xjqH0IHgI
eX49CMNIUbqNsL5z9neRMK1MsTrjfEJKwSaSjEzsAlWzobqnNWWEkcWrvhHKimVc5Mlk7k0OCkSZ
qVpV0eQjjMCsxWIFNIfqtzphx75WXiD3I+1dCSUI/IT2bcvG2t7amrccTKEJtJ6R+8aOW9QhmlvJ
p0iDUJVh0Tf3/jxNLI1tgHEk5qPuN/ppjHz1dIh5oKMfehrzScRQZhJfOpXSn7JjY16NOk8a8jWl
6y7thU1zxnPBgdo2hwJuDI3EdSo1eAQzCX4k8KLllvpM4ysoEklAHaQnemvDjMsZj4TDZwqDhnu7
SRTrqjQtfr7rTEMw+RKoeLuBcxPL+FZdWTCPzOod3ZkvG1beUF9NJL8N/1uUeTf0+6neE4HgbcSD
dac4+9jC/cFevZktFtVAoHZ1BmRJlAqJmM7RQrWuAYRJNzhAkjS7qebUOEpbmJ5SqfSoBnCU4xak
V8IaIL3HQWnESR90Eehrj5WE2A1Y0a+b0l01D+i8IgoVwFTIImfNCy8n7v2ODv7uK8LHYNA2NLZb
JkT1nHcW1J2WXv/Odt0EOpARN9WNay32KJeQ2zt+WYV/clIm/kWu6Swky3r5ncp+T9vWxq6yixo/
1N4yyDwxrcc+fme1Xr9AJR6z3DRUXZg3tbVF9XD6aMSZPfz32TL/vjK6LpgCXMgP6Wea9c3Njmtg
C4v/GyLblEP157OzIOP1nIeh84czq11r1s0ceBQwGwxr2MJZzAho3l4GUPFUIEAMo6t2BuMzN90e
yy9aFg/XdcFPM4tEj4AEN9lSBrECY3bk7lazTMloFdNSfigaTBry52Bx+XKjlvFgqp26HGTc4anJ
Qu21Tr+tDnapMNoX68YO8Xy/6tavzGmWZy2QqANlqlknAlmN8/SjmiJdBblyZU1g2zM/2twSfCwm
RCLiv9VTujgUlA+UxmAJqBK1kgNRPSvDF7BVIYZrUzy75/aFyiLGAlSNz5nPg4/v9NGZz74C3wei
DVGw71cu96iG603OFxG4ulwbTOnRLHTS87rPqKYHnksoaiVvl87xxLQtTBJJJmhUoKVVAHL0XpbJ
jLrgPZIr8olIIcbdMnmSAMiWwWEd0n9Sokp9fio47dQlAzQA30UrSdsUkIYNp0pov/SKHTxqYfHr
z4eHAU8G+Ug15hqoThsfmXyK0u9BhZIicb2PuVHgljzYYIV4WEmaDcA2aLedWek024a6sN+Ao38R
0fihNnCyRKKS/YXlebKXdkQm9Ip/yDBVSiFFuMBXFNixrCCcNksGZ+cTRA+Ch8hcIH5umW8oJfYI
WicXXQ2Ta3Xx9BZk2zoGloHG7Ox4Ym4M4y6JrGsUsxRhb0SYvJZE8ZSg/qjCdyrd3UuWlRgnQeOE
Tb9m+BxXljgDIhN/9CiV5YXcUstvBXU3K2D8RDYC5XBA3S7aWJ3tYqnZATOb7PTcunQp0Ww8UPSl
5pBz81BNbdLHlGmOBD6ARIx8MfyaNC/0IwQLJAyRGTeHYh8IieI6KerKzhxQpYe4ArRX/BZA54N3
U2IGGsP8+KIjhLsjOZLd1J1lBQCs+ZUYkYPBCkI3f9dxLe3r/MWg3pFS0eWimoEE9tzGxvQlQxuZ
Q1M0h9NA5aIVZQVuIiz7TDz+WwFLmW/DFu2yBvY1HdQxE+fQvMsL3Z0Ar59gRoQnXv3bVBUa+hny
Areg5zHPdyv1lhEs04PZ9s9rx1O/0flnRiOrhBFWCU6poK7e28S5Eo4Yv67VGD5MRv/Ds4EYTHGS
EVqgVRUF04eYrqFj0kvR18k9foK+5R6fTddq2xfeyibjGXc9SocyXeRdSJKJq5kyV/RcP7dg3oyB
YYIbELaw9wO2PTgZL6+WCC7DY3ulcY3s3/LNcnX6PFEnyJgnbH3GC708yEcDjKX4ClDsH8xPpS2t
LZnlBnEoKFXDNJ6JZIFXX5NzbC4VgwHz1aT2ux/eUJthnso7MdEawFYZtpzUHvjkA2DJWTHx+PHh
AyCqKLnETeTrQgVL2ipQdoIEZFp6lRTOoUReowOvzZUhgnF8ATZp46S58UXxzw0/acWHd4JyU/g1
Y/Xaz2RSkizALbUyt9lyUP+5Ro+Rhh25SQrRyx5HeHck3tZ2l3joCJjKvkw4uscPAz68F+YCMn7H
eDdaHnfwhMmWSoy6G7mxoq2swfAHb29bAbS5xODh05uv6PPQLvOtgwmD40M9a4qrkbTrLkTj8mRb
WCkKo3jx/AqyQlRxGIi5Kt86R3quRiD2rpF9OG/bzMYhqhufQlCdNvgM59Soqje0plB2cASJfGD1
lx8hEmuNFJBiGeDNaIYKI537bF5TvhIykuiHrc2myCjz6z8aqbOMrMNfgOnBmZHkzqva+8dU+/nn
n8mhTFlt0VCdTvw+JFPhnAIERAoq5PkxvKzN49gUjpZ9MMzB4C60L4fTxtjkJxknl8iegcrFVze5
E0vzlldsI25wd2G/HHiEeQwtxp/ORyfGYzmcKebuqCu/nMXqqWUZTynKq8DB3bGgOeHzqTivnALp
42n4t8wnSxWQPTCIruqf4iGjD2DupNc5M3LAtSnVjwimltEnYMpEg8BH22A7/BX3UvFfIloZiAtM
WOhzJWLnfpG9znw65C31tmOlSOZAau7kjzLqA+wYOI3W9PiKLOZsWqUKAZGGsgBucn2vxtPBnSpa
K8/j0d3zKxQY7ECMO7/xbQcSboA3hxBft6BLml4IGS31VgXaeZQRk3bekklsXSZInPjNFVFSMUe0
tt4jrqqAsYvvKPB32cPmSwmihqPq2IiowqWeLPu1J2ATo2QknMrglFCV3quwE/8e0hfXmI77j72T
Ko+j5YiI2igWWJzwTpK4jl6VlRpRxc5UUtdl05389yHH3yGHgURHF3RDTBMZkj8wqPDP3/H+BD3p
hCxgHyGAxMDcOeTRuBl/vqMl96raIhGp8xNygv00jUWSeXvoILm0yltkpJCjeMnd3J+7ec1yUU0j
u6/4EjlExAC11bnH7z82YuF8TU3Tbain/6rhdgQDGcQ3T8FNX1R/CRic0cgV0x/iKpFhcE8fnIrA
jzMrNN0Dh6/fW/4XlC+JaBuS7yqqNSdliZNALvxYHG6KTp+Ah2zbbQdgMvq+kqQ+iXRh6yXwUBeG
246dprEnHf7r0CflAiQ4TfY6+6bnCb8gqFKcLhe5NetcFDfveRdVMgKaiMhR0i9anGjvOJIb30+x
t7F5cTJakBL2HsQT7I9Q33D43RRI9NnVDPgVUgdXyVuYdqyTMKUwIMkVBIOLdWFxEnD/TnmnFFlF
89iQjL1GU5vZY+H2z/N5fFgJQJdcBqBROyd6j8sQQ7G6uRM3JIs1Hnoqdp+7DjieL1oN9g4p8lSa
ex6RexraOl820fospKDBEMG1YdiVF04GdTJGS3LlMfhdsMDOEPS56rDx9ZPdc1apWtfrY3V76f/E
Tm5OQ3IOoCSJntGmgmqBAF3hpEUcl0yfdncFS14us8z7rbvUgxiAfJ12CNjAwG0NO3Wtzq/ULZEE
v8c7eflkHiQrGqAOp40oNEUEFp+mlA/D1wVE18Sskyw5ouT0VlbaKGNdrp8oJPYmhYytWySMvphP
GdTilMAw5MXVQHLUvTeGJVSKY//uXg4Jn0a0zaN83ZtA4zwkJjRZ1d//hjHGOS9hT967Z3SUZbk+
d4dAr9WXq7T0bnhxUPnQqQfygTq1msHHmbmwKtcDquPbsWwipwQ5FN8H9uo0v0mLq6ETs7up5r5D
RQ01Stxf0HDKLZXFEqoUb8Hd07pRM71Fb3ojs3PeDEglODyZTyEESqToZJQHN0BsybBbjtev+GiY
6vjgf1gsYjT0X+iEQ4SVjMjY/kj7V9a+6gLJdptwPB97ZMAVd/M3J4YOEV1/M4y3KZLYWqUetTKl
hg4kVN3L0+cv34l38H+9oYeRpktISXaeDbtzrnaBoP3h9u1OScmR7tVRHMhi2jikMLDL2TblXR8d
u4HunUFbbcIQIQDnPosfTYglvkAqgF4FtKahbvRH9zdLt2HAIdShOWCyGQrVkfC2Vztka8d9jSqf
stNBvA9g+k5r1W+fIVfmO8RrDC/9rUjkefw9yhJXqyEvojmXW9Ool6rwDYWF7NiZMNUtLigBVRQ1
qK8n8AeGqMP4xkMnsEiIZr7ZivvBuHJqB2UZF5y8lZXyO668oh+tmYuaLfWIaRLOA9xaAdwly7fd
hK8xgmGmqm2kouENxpacIi9E/TBkTR84MZ8sJaFnbM0pyFaBQSh5MeGJlSg6WHV//ZwXGMfoZm2d
Tvhs69+nAXziGec9qpQ5C3SrW/H8kLt6xVV4U3OzsTGhm6cVMVCWye+DhLxCIYm3lLK72DxlVB78
QLz+9tah/4nvhoDkwu7AHm4sr3YEvQQ/ACsS7RM10LW1MFjJH0UJkd1KOFUCD/n2Ve5Cl4ljzvTa
ITVRtslX3raZt2lZx4h7RB5AvsMZOK/3qZSgS+IvpezBCtLnUy2uoKnJ+gkvJA1wwYw1CaVsmGy9
6yKTw/O/U6aMjBkWAAdLFpXm1JlfSYIQ5b/JvhWuC887ZbWUf3D5lau7hNxWRxDj2zWQQpr5eCJY
CLpiPuFA9OBh272LVMwM5T/uCjNm0QkwpQf0Cd7WPIKh2NBi4ouZu5HJSt2lOKeEdSaDvcwWDGID
RvLwdqokcxR5Xw3Qn2eVRivIYkd7hNdAhL4e/6flJ2wCFcjxN7rkcFY43g+7FTV71A/o1sdf5jiM
Trvj+pSm7HslvDvMF5qRma3vMlM8DVctpjaGvel5Zwwh4EddMay7HeQOTWUL1v8RFgVc1zqA4dDp
8DcZiMj/MpuGD7W+EzCkj5pKUgg844KpKNbf9Yfs7KC36UyqTlmRfqm+J8TuYKtpe8GI0Fm0f5TF
emk/ew6pbELZD9wTVb8F5Gu3mA53e0bs6mfFClWK1u7XU6dKYEkzj09MB6+dtVgfek6GGTXsfew6
E41FFuC0+sWhiRoBGCbBfNAlPHaV1rQErGZ7ruh+Cf16+9XQwNTmAefVJEsHlpzxc0Um79Vf6c7t
QV5PPbiMMCCuqjWYf5gGG1OLH9w+Hth0epxLn/YdfgjH9pmSNR8raG2pcnJCjHzlykdkJcJ/mGg3
Prnp7WPwXU6W9ENcmhY0xlh0yPlW3gB1SKRPgw0ZRwjYD5n4RnlJZ3tKSAKxlu1e+EMwW4dADUrS
+XFY4JvgYYkRVQJbr3KeT7Noc25iSFsldzYVurzG6kN01I3JL95p9Ue4xWc2atznlGsm4W5cHXvs
qdXdVGIBIDq1JBCFIICB8QQXPGQIhRF0grw1wkWPbFe0X5mQlB5A70hbcmymnn2tZe2L2wGDiaRH
ldWcyctyL1nBXz/BskFrHrveFJeJ2JrRefZrDEm7b5bouX5Up7xNsbgdY8sfGO1/qBA1lFRhyyUV
LKWNxh36sgxwmMYxxUEsZfdtTGACoX/GyYTcmh1zivT6hfEhaVWTaKTNudq2yB8AJ6j02xpYDYW/
Csz2poQPFLVB31a1iFvAcp0/sPpUymURy1leRkLT1VEq907j1cfHqOfM27Ty+3qzr8NhxrH7Lavp
ccCnPR5PheYdAlWtLnkyPJ/d6yFRuxAhXLN2D0ae/9HRi85kD47BzDEGTlp6dW20secwvft2UsCQ
+IHtbJratGxDEE93TjGPT3rCa72MF9wf25vQKFK59D/FJgRbBryqMBxTFFx8uEpTlhjxpYfzMnIT
hPi+fn+B6M8IvMRLL2Zh0JKQ2AeMHyi7q2okcQj4apqdn3QtjUvuSqFCIBKChknzBBYUNrRHLTOQ
O7vEN2RDF58Oo1BmemO0cJFUkH6XfX4A1J21h+GFCwpfgB+Utl1ckmd7+9p2N0mXjdW4tHLdbitt
zYfjgA1bE6/LQTQENJp/+7Z/QyDuv/7ogitEJpXqPOpGe4xUOqbGR0aBH4wtyKKdwWqMC/BQN28+
NCyaXGwZcxG9UEuyeMja8FjJ1TTWNZ47fTiwspUiycdmIoOdP2kcUybf2hl8RTB1fdt7llfHlpDM
wtLIeXo1VNhtJDRSrXmsusaCEjcyakQUIRogonU1jl3u1HNqRz6gjcg3p0Q+badPExhpKnGsQwLK
xBsrfFM3ylzCwyXgpx9gfuieGRfNnS+H2T1BJZ0XMqqEjdYcFNgYSOKdo50z078mhMK1vNSLqVHn
6p7e96MR4ejR5T2MdM+xy+2Ce9mHKWWpAPTcZqG8WG8Rysx90yg7QoR+wqf6BzFlgsZdq7kgsb3K
OmqCaP1KXqDPf7qNh+s2YAI147v0AHEeyTSQks6GiBDYN9uoZr2+SjhoccevVffjUFdU6A5C9os6
miYD/hDOjOdSLGzYbgEdYWINy1jGrijoatXFF82pI6RtdSpFHN+31TBrLmcX9tMgGFn61rzp4SCK
Bg5KeLMSLv45tJhWAw1vvM00o0xrJB2b7huSErfmGTj9O3yD+fm8SjGF6In4DFhUQYG+jXJ6clId
Giuhzfyav+VBhpmNG6p82KkCHpx3aB0EMhvaz6n8IHW9dArd+l1AfLsI/7tW3A/hFeU1ZILdQCYd
HkK3ffT2UQhClV35jHW4H23p5ndWr54yPMDLGTtxLqNt6a3dcP3m+29jUGOHjNw5hpsxePES9QXt
fldz1dz2xukgMCNbDBwCEpWJKIAyHOsgxecrsmZv9KQCVFOvwgMIs0xvDGLgRJe8Y+y5+6Gl4KrY
GX6HnKiNT5nlLYdOmiltsqF46Isu2v5FmiH1HWq32X6ZGk/UCkcWM5GklcQrO6XntHMjwnkq8de5
6GWALOdqkEknxtMywXzavrtF9B9/Ex5ds09zeReRkyMLlOFvt+o/NmgFGJdUZKWfLNeqGzsHmXcU
vepaUO2alhUQ7+8sFVRHqEqwU54cHtzTgsC1TCsV8fyfjw86ri7aPUdoyoeblhyyy1NPDe32J82k
nTxtPpU8SMreAPOm3n2Pvv70plwPN0p4E6AWQqFt0gVq7O64i8eprPq+efKVyAxbcT4Tb6bjXwU1
BTpeUgK2SR74WmvG+/N4moR61IMJAwPYnzK0QC18WaxSjFAvwVv4M5YCEYq+FlnC/hYehxSszsHd
cquFPRo3wA2+zISZ/frj+Eh3TRVPBEopk83GDBBVdFTcIl99b+AQcFMrx/9mFmBT3NBpwaiTyPqy
efBVn3tBsOuTN1VIiPLjKta7blPWk4odX2bq7sE35WoHG/6vz8GC/8CPIYUhSDrr3Az8e/KFIwOo
6ipjIQ/scO1MN2twE8tY9lp7E2fpsJExC/wpr6ybAbkCWQLUDOK/N2RgKK3Y42VM0D6rovw9psTL
txphKQMzBnJpALAOyKaGcTysMz9VzzmZCgYYFva5l2NfT0RAavAN67usaaWHIsDWsxIukCNMMtxB
6ps6Tbisn2fpAgM7/n0yFlIMaOMfAowTkR/d8KcDgA71g/aXjxC3e9vQWkNvJScIQxVDgI5s2Lci
s0/ozdhrIJ1fekgM0wIh9QufRUDznrthug+fa64OUhY0XNca3bvSfvryE69UP2aDh2zp11XXBVUq
jALPB1eRn4mcTd6mTdmVZyrL/xWD/SKdoDp0Sto7yCEAM1rxWo4HP03h/yMdelFQliQn9b5k8tsi
+8ks5UGVfqsF7gIzXYV3wrfCByKdhUvCKyQ7A5tP2RiO0CNapOtuMCq39uxQjuZuAPtWq/LWmKK7
oODPMxCVJGAWqxGfxiNhmc3IzDMaETZXh0WJwPww5A425RftRVYFgltTqzX2Fu9Bf8XcQe/b2aE8
NLwG3AbWy9AC6Eb2DqC2BTKbbtmHoIsUNefN7sqALzQOcvr99kYfm9ry+yehgQ5L6asVHII1FdDL
+5Tto5Cct+UKpi1PlR/q2UyPH/aECphMLL1o2pgjTVbEBXGVYg4eJgLMvg8KN6HdukBvhrkaU2Xq
0kw2kqpxKARK8so3/VbQfvNQg/qf0sSo0CIELAXyf1U9xRtT76SgWfZQA8mJga5P14UDcseUDcb5
XpCdkl9UX8NLLGHLJu7TALHRGyQTxp6skJjoyl4KzC8FesDRuJuSKjSrLDkIIWBSvP1HiGZDhk4a
Asah1FEAChuMXNtaGZsz2VdbfJGYyXMgZo098rFYVYwVqPbZWZIHZuS42jbVVScXiY8beplzDryf
WAVxUY2XsgkloKX3Orf/d3YSbwrTbbpL9su9/6bXEBoajiJ0EvI0bpMtSbAdgIrOi6nLfkWeUqSA
A4sq+YuKr6+71MOXikhNNIf9pDL8wq0W/cwaVVyQJHBLWP+W8HjXAnEtgn3fXEKmeYKe0WWFGpin
uToQjP1Z1fBiSfTwPCbGQ33sICFFlqJmZWH5mIntvkMW8xHUH6JKvvZOYf74g9H+szcqDSyLM2nf
1PdynwjXqUHI9oOCLnn8OZf0t7xYrDEyvtcx8zXzgjXIfCky/ORDG0LoLRi4fzQp+k3J6voWCnfH
2yCw8N9FUorR6z0dzqpZaGMvwWo0yB6003kLUiLZKiwsFhuM2t3Cf6rt1zchPGY0Co0y4kwt9Isg
bpBH83e+T/uigYRk94KkrjmebJNU1VCk8EK2vsVk0Q0BmUnPNLr90GipYh4dCSvsWcUT/No4HO5S
SMTLxXGP+XSjGxmI5UuBEai3JTXWOVRO+eZ2DFP0aopsudy3qyi5QFyyoIiSIPi6CniSAShg8Oo5
+WZliCaICq38t51Tfpq4m0HAQrLxYujj7U4lIs0A5SWMYTGzD7QngZNBbBzSQ4betgpp7h9YE+Ii
F8El8dr6+DkTlvPPG7l0TcDRYww0DUG/9V1psQcc4pyz8Ee2wVSIFw1N6mTS2SnDdFIn+j9HrIFT
XrQq74WUbCQk+dCKcYGPgSi0/MWUHw+42i7I6vGgcIVPrnVCHPTyWm+cm703FDV3V5v4tvij6CnR
YljcuEmavvoLYKpADqU8rdbDPRTDktlb5WwFg0mO/7sZ5TB07H3nqDaERMMwEMSolqFckNatyW6O
BvdhLWbmhhbQ4oIiO+oxTO+oc9P3dbitZobMA5U2BANBev4tmMWFc999kD3/uUcRQeoJZSQYSubq
2AGqVXZWFwlvJBj19gtPkOK4ToYZJJEiykKKYnppqfxe770mlarM4PThibiBoxo2OiCh6e26Njlz
lpdDQRg3bHQ+pvG6ohdspyBrOya1eh6OAS1rfIhLidime1ERN5/Sd9WKqVbxmrHRA9FN8iM01bv+
bltxRl//0AzOP1/MVVh4F5TItqQVTEpji9soEj6utTgHj0yoP57/j4mtAKLYgQgVGrMp6+4ynPdj
QfOQkJ4I3Gkpm3KMax8kf3+/RzXAYRiyQq7xT9Rm+VtcQa/GaI8j9xw3nOB4r1j0owlnemLt6Cva
BYh/0ucEFL0pFblpAksYbaaDa5bimfnHGWY19uc2SfexZnfx24aJyLOt1hUpyeCTNMfIZK5ipgRN
1Q7yMxozal3LWm/XxFd3cgvT/40DIuuDy32mKfwsBB2WL2YiT71UJHpAoGCi753xixi0m3gFQqMK
S5o4+JPRXa1BpKNnDBDdTEW5bhmdi8q7+CAimJ/ZbKaRujH9NETVeRw5f3oHy6UAqAfZUt9VU/Xv
9GEuT2voAAYVctFXt3KnpDuD8XTg24q1B21iEsIR0erGYrpLoX/rMwp6ngv1TcXPddi7LjbcN3yS
RTDipTlolKYTK6A/D/oCQptMcvECgDMwuNWXonzIqvp0P05EUQJ8NA3FwKkRUJM3EQi9cRtLmJ+4
BdyqQ9zygSMqDAAXwtZSSbrxCpQPSrU28DMBgsJjre8iTeZEE2PtgcNBjudYwj0svazhiFzRP2Tc
FRQ/qykBCmOIQdjd/yOa0xMtpiQ5rShrCngc2xEqh2d7WmiRNl9kr1ew64zcfvY8SzDI4khYSZ1o
InPMUknGWruudKLazV+NFtdAZZPZBJu26y/yJcChzpi9kbBtptI2BPXgtjadVwpPX5ocGO+YoUOq
QLGIalFeJN6xPnEYF/OgBxWg+D+Zr+SbgbaDoDGBv10o17zN2qxHEXdLOqEwoOQh4eVzv29eCIyB
x2frifXbU3iX1flor1n+Cg+Hl0pWlLrLHWo0bDPSbGge5bZv92W1L2mwQb35A5vIgD7Og05XuPKW
M9PQQ9OEM4mIoBakxlPh+71kcrLfL1LmJcVoAn4IQZL66c5dax65B8ckS83i9ryN4CnR/zAQcwu6
umfwopUmHXAhNmEuVoJmfyKr9puSo3/ZTjrhCWDsWCLWEtpqN8ePqq75Vmn+zyCdQgEUXIXYPFt3
/RivLlSZryWqhiRvdNXhuK6gvIOJQYuNiECjUY3u3yLhFHNUxIobNEKoAnHRInCjSz6pCc71KVHb
N+dX4k2hJbkro3OnSI2xBtVDqWxw+r6NihJeckM0IqdBjg9ifjkwxsud97hqf0SGs0KZuDeva1At
eoYL3B2Og/iZlLqUOgz3tbEdkhtYUT/XaHelGjPnaaqINesF0z/aC4JhxWIECjdQHn/uNMosRSmU
BeXVXcmWBemVap3Rhd7owSNwb4EZGGol+mK1h5dp3dvAzCzX5qnzrofurISOKc69ZTBe3ihnnHI6
X/aS3MMPwgVZO/Md9RFFPwuzpYxqArVUzbY7wBvfStsVVwRn490HTAyzAS/1I0+6yJs21MwwaU0A
LqsqeoiS6DQE34yb0H2xnkq881rPCA6IXdO1SeGH1thzOrjvzJ1NeLQFs6FqbeJGNIeUoi9rvGLx
BMrq2oqD/rEhK5fysqsAPo+xrfoevAwX73BOvBn2oCvIB7sTOpp3UCapKgGxPb640Z22nq2T2ejk
lHM2z4ZNE3YcgVzCDQX/PheE5XpaMuqKUGnivhwUZ6CP+uN8oEyNgJFvvBzxEtff9vnwpRcRvE42
0vgo2shM263M65Khro/0YWPCZUYtGQyMFOix/X5Y+EPkDtKoJ2hN61zr5VeRykdG6BaoqeepBy+3
ux32rZ8jl2GZ7vNFtw+UC8OLwjxYzEzREcwxxQSuW8fJWpgvpuHiw1N/L+JkKqlBOM7Pt0YI649K
gNUvzv9EfUTwYZWuAmk5DHeZB9bT1b0kj4JmG19r33PMuOgg+3Hx2vxnNRDUSlUDX+zcWZO7WLkq
J6JLjV0cG24M6mPl9wqlQJ10u6nKpge/jk1via4FqLHYwJNPZ1fQI0MGkK2+A3cQ3Fdeg8NksupD
7gr2xDX2kjTZPYPY4ZGGYeM8h+S/FWgiLBh7B6AQgRFlKvFs4JZvXkp9KouKj7Q6AHAZ05KRsoc6
uq6AZ+rcgA8nBOqsIHflyWIFlrn5PHwTFXFiq9f9E5AmDRFXi60E0P6/PA0VLZM9iBA3xLVT3q/5
zO0Gyq26Oi/5obzYlr0ymh2N+VXAZ6467j2W/8Rs6ZptB5ogz566JLTIe1F/t8t72YKCyIZBXUfu
7s3mSx/TNLrjtZVjE4hCYifwXSW6iH9za+XL8Mdn/Z7TxJLyj+yBryqevvCwOT8XwidNo2jmEysM
EfoiX51vRyS4My21UqPSsClu43gmKzOpluwiy0f7M6+oIE5ISIE0tKQThY1DOFyxLMAFMqqPbmbT
EoC5bLbga7Ss6OGMOz8WCIP43vILcpN8HsakYWjPOBZ6+Gz22zboeX9LHDJO4/CgfoFmyr0bIrFH
u2NPf5VLRzpJT/rDRfK+w7AAfuzgkRBMLiPrBTxjZvk8yBXnDgiw1yskBj5CXV5J6IdlPeJA03SS
3xSlsFGsZRuNF4vMJt8SM4LzogWsm4k/BI7A7xtlHZWJkeG2vjO5/24/1hVOOyMYLfNONMMDOsWG
DHmhhnv2uSol2haxj/GxfDwHoL0MGcaw12GpjqH3H9te6qdvQ7Biz0zFFCk08fF0Rz2DBoaiYcjC
6G2wFHGd+a20+/pZxYcQavvmiRWSigNJW5tbggwN0myxYV4EzJ6xJmbPdtrcnNSv7sB47Jr/EloR
Ooa5+ZcDeWDrmi7R9Qn1gOXGp/wMEqipfFHrdIGyUFQk9++GOZgNm4+iM/erb7ihVohavttLis/I
p3hI+QZpKUwpVRV3eU2GFZviHvGmzoch73MuoWrFg4Q2KfJQjwnv0wSGD3gSFqtzGoZkzGFkJALq
1BEqsqerMaoBGZ7Em3XcbgVX3iiaRI1Zn8jZIXZAokTIB6cVt5RMqXXfnz5KfMQgKmuPCHEyoDsf
Tb2PoPDwI2Unfqd8Aiu8GvO8NAFDIFu8bJblm0ZgPyXp11odnUNzMgbcKKXPthTISdirhyi3ZOdG
f17XcxoPfdkYRqbBACoqDKx3FwmP8jv7GLboogNcnCbAvOxUmqCHnRFXmKXZGBmhGkfNxpda7Mah
nvzC5h3qn+qHETa1qi5GyjbCSyBfu/tqW1zF6WZPQ1W6FNpuHhyVGzbCuJtzDFwDxQqUnDGVXGkt
vabZqNajlLYm3hZGQkHtUzEJ/oVj6JKJHfRgrvqW+4O1A9hn3rNy73IqIjQWnsmNn7kWSkrdsIes
tZLtzSFoLYzudDzn8ZA+RoaUyQ20mDVA8RYQM3cQu6qaMFCE5Xalbfp/PA5YNDg1cobXU9HunYa2
RKkDPf9Yy7e6ELjfv249UDknsQgD8KfFuosPMLwtxOYjxM+ambAvHzALrYjxlsJnsac7cTY1Eyhp
t36X0ozJeFEYmniVNw7OXqevV7g1jKuExJWScV4m9T7gU9ALslVz5FQnmeDFjXm9DNzHmSewgvsj
INs0bFvUWJiDuvrXue68wA5FE4WttQ0ibZ0GuWRZI2DcLQyTq9um+kPerLeZcignlTXbjAO535ah
JaoYDED2AKJZ//1XFut1EuI3f8S78S4e5/ICUr9VRynJCV+uhKLgm3Fx0y9kiqOaC5rJt+SEZEK5
WwwvjGA77ddUI8hLISIG04loz6JRS/4e/nLnWGrRpa5ftr8QqyEQqd4q0bewwh9O6H75NsSvQUuM
PiFLp/KfaKlI/zPqdwbfizrbmGr33Igrbm1cmDqgCcT26bxc+Kz4bMU6l38sJY5YuehgzFOekKWk
NZZUzVavjG8wQLBxybEELznlvWez7OVRktr2HnHwUJa0mBXJqQWzqAPit80YtqgetDPSQNSSU/l8
H7ByIvSTkIL7yObEeG/Q3evMHRJrxtW/+O3vJKacvSpJx5OqWcTfyjnAchWjztS+2+SD1RgUrPuc
hEvoIWK8go92ZhQf4PsjsrbRIZtA9V8KXXW59wQINY0GEeHbmpSZwkQFYRBdv/GCNEMIJKfa/9Na
lBcFCwKAkmprYqlAQPHwiWlKLce1Fewcz/eCkOLSebdAKImqauszZxUtIwIeljA1E2hhWvNtozyX
jmCZGV+sCFA6tFInuWYEGKrc1hyEgkSnx1F13bUS0zgzKiH0tqbEks3drsj6dmLnX/9NU0GxLCxV
NQASDCvTGGrfvm3Q9jEJlIS0b4+qPvF1Hs5Vuz3/U79ZURS4YQh0/EyDCTSsLR/QdSrd8C46tqIU
KRTUOYKes7ZPC9IzlAGTjRtw1/QepaR2OIy5G1qILRWizBDXdXt+5zXBiPnqhQ4t1x+3rsd0/upB
xLZ8gZZogqs/MOi5r0ix4ycjo919H1z+AKYLwkfiWZ83v78y6gak8IG09KtjbI0BPmByC+90A2Kk
Zq37cKkPEPhVwKjEq7ChqKcFyMSYsJZtRSJCLijxCLwbKBTcvTb9nCW6aZd5ulzpEwY6/lrC/Nzs
ZB0z30g3SN7B/5CP0ltIrRFl2QQ3bR1br350yjO4rS7DD/KO46AhMfCepjnrelNX0ZSQrc5qIM2v
H24EwG+UZ1Lc2LNHcO6gh03+aVrVO2lvTPVW0vgBFuenESFsHb2Eax7vgwXwe/hqvcMBZofNJ2uN
Pmx85C363mK/CeFTEO5AGHqyn88SQI4F6+wzHrvQ7dCBrYAOr01wyIRj+78YNA/NpxY3C2Lc/GuL
ovd7PzxQ0X65hNnyzXYElEgw9kkceBrowqeMJmDWH5BxIRuz12ILxP70ystVM5JeEdGKtVmCmYPv
9LIpzaYyC7WNU/q0if+PalP08M8riUpcGk5Z9/Qrd6lGhHw6r3BGS1gxi8Jp5TGwCaiBapLlKtpp
K18MpOEQCV2Dlc/UkIRtippk+Yc7QiKu6bx5IUVyYEdzxsvZ3LWjfhsCbqESpUk/XRmMTvoN5xwg
UB/vaW9KWl2Use4e+LIQWoN0F7vwgeSx0lO0gXij9HW4/esa4+LjcbCZxfE/wjBgLMmkmXQ5LZgL
0f+IbjMG+Jfdvejyv6rv/La4ghN4T5uVsLrCLKRWqGx0IzE5xRx+yStjkw7k9VYAhkM+WIP5HHeG
ibXxNDy5Nnb4P8JMUq2wIz1okAiT8d5S9TErl8jbMpecPZSxWeIXvw8iEW9qEtw6TR6vb1Lh0+IO
CQ7L56d5EoZotrkgSe+GH33rTI0j7QMNDd0RkX18V8bklcp4YbY8phwOqoIsQ1FeMKKS6IKLD9Fx
hb8NgmS19vaTnaG5Nq2xCYhg2QCDGq3lMX+GcWloo8neDN5MlO+s8b4Wirmgd7E/4EO/VbnReNxB
Sz9pmdiehdpnnf1rqrp03jPRISFpQ5trMWPEuwIYcsy0XMAHFQEOVaO4eI/nkkPNs53loD9Zop3z
IyGUFbFD3WYTZzhp9c0OGLKN/s7VsE80qPZgMxC1hjF6VWCRxU/RgPcfJlIMzmB477hzl4A/DF0W
PONiRvUe2TPtHDeSnM5L8cZvPmDteko5tMW2CKbsPGb38ua0Jz4zhDo5jd3nMS/Hi5rt54yxC7ls
AmjGpgxtA6qJHjgay6E8Nq+Q0qAdH+nCqwU61hiC/ZTat2Ly+yRLxF3HMj1c3IKlpaygHcyxpzfK
imXqnvLlpdoHYNlo/sK2g7VWA3PBeowmbt68VKigvLPZqfpglglgGvbb4MutWkQ9U1dKRzGgufC8
jN4b9gtl6IhRfXIFmchM2ljQ0C+uXHaSYljWm1XGCrbrcQ3fQ/pxsoKMI3FgO0ZWCXq2kSTAynPh
YCum9nHvF9yYt3ajqr8S4Q1qRFvV7S/FyNZBgGFfuH9fraWgjDpa31iQjN+xVlhIAst+S/Uk43rF
FoNl6niItPNmfwrKWK6Y3rNNERAm1swbNUKszksfcN5RhkcXbKrTf3UKSX50rdF8CSsAB42dneeT
zkpalVja7F3/dSEMF1mTwmTN81YYDclYr1JocGlDDRZvyX1AbcOUJucq4dhMXrXwYmDtKopVQynp
hRUVHu0iF9L65LKf7/+h32AAV20ql8MQGngXlGt6CJZx51eHZ5hTPigzGTvnli1QLmy8pC8J5bEZ
BFAeO3rbIIaKR0R9OfqljZCMnENkfzkqdRtDLhc/E4MlSYUXKaGPMj8rWEx41x4syw+PE8LS3ydw
iGVCma3TBmkgE2ZJRvIZGyjJw/DCavd9TE8oRMBqwIJHKVYDK5SSMYpwKiOTwYAfQipWvu6Q9RWZ
SZuhHaLq3V3af4JR3nxCOxGahmM/sOcsyTwIYrrH4aJ7jMOg/+wIjjC5OSofEnd7DelyWTl2G2dE
Yb31no7ExdODGUQABTyl1dmEi9Z3Kh3kpe1zDrllnC2c/7wEmpurIqXVDRrp9Sxw8qwoZ31rFd+b
bBTN1KvJs/NkaqLiRAJjqn9rihhZShIVq7C/1+FIy9IfK+PbNRGCCijf5gBRirZZZMlWxxk0rJSr
YtOFLpwH2qfsUcyvMLFDDI6sBHtBppHfiSCjYJNT0e6asHPh28lkBGwcZoOnElPSDrMCG9PEyB4S
hxLWIhAmQWkjXKggy1kLsTdeaxIjs/2xUtdfq0ajbWJmivJtRhHbw2/9G4QgcW0nQhgBclxkl92h
wMxcyNP36NFZXOQJsw+Yazi+OduotcK7FlQr8+rA67c7kGbszE92u/00xm0nGeF0666dZZ+BN6Hi
zt7Hi3tKwO2zU6SCb1hMHu/DxrTJQd+sryeMfvC5wnAZEbIUVxd4fYTkmQJsyjO7ylVZUD7cE2sx
OkpcTH50q9CmaGWFGhuDEdpu/k/2TOv0VFpnCVRv/qDMr98G+uU3s8YMdMX79AU7GBJncvJx/6WG
D8uY0YmjoV0ig17Ys2NFA81hfxcZnMOurxTHeeAdfMuD6NSkaHwAysQHbvimIyKFsx7oxWcfawhY
JfxpbJza4+OS8dMT53/OB2nqvw8p0VlpF0Tz23icmBZuIbVDv8NfzsmundjzreSRYUFrI2SCuCMf
ZS9xnScSp82hSzOungy2q25cvfxUcXcSRLa5dQngPzMD2eV8mFq2MIhUoxEjqIXdrTvZ6LMsx+7y
RjMfwT9XpxGToMVpwR6OBTpz4hY6yRKliYyiGzQjqU1QbIb3jZEhvl5kAXD1w0V8GDifeX94dNbv
WToZZ/TIqWencAD7nTu57vV2h6P6csbs/VCcrHr/rxAXCx89g7yRClgNwqYsJlxsfiBQf89lIlU1
qLseHxW1tFewKrp71gBiKo8PxB7gpPNikOfDSNdwB3ZG9iMxCVD5fTtF++8/HhkQ963XDFFBsaYr
XHgKDRL2bUK00FQe9gUW5wp7EjMQu06JlDZwJsD6CDZP7aTSc0v+4J8ReV4EwrL2XhDRy0Sf2hVA
BIAFS58uN1Bu5TiBeyHkKB9r1ZsXnu9XGQDotN2LaOYsOhQtx2EemDWK2/wRqX7cIcLddfX8rK/K
TsHGco+YnJn1O6Ecj7JJvSQvR8maOKQEUq7mFhvmKz0KwyvNpHouLLxCIkEc/sAPkDv+RdTstUXi
clRFklqjcPFzZsEVxfVLn1MaAiT863q6XRmhJA7gY9axob+SvRaxG7xmGtT9At815um/t+laTpy4
8p8y0zQpN9ZaTgccqGlzL4scwAynVLX41fjigQYTmgH5hTXCVV2zHS48B5JMfZ3Ul9Yve422tOFD
J4Ql7dhLxKAIq/EGIJDkdQW5erhRMnPkdFl3AdtKs7C8gvbQbEWR2kDNCOOIsGUQWVlHHPTI4Uhh
4amRmw+copZEMv5foP/t1ldfVx11XQh/XhbutZV5AVBwDf5qa7sdO8RvyLr9+JtDO/fSHKATE9Ow
TORy1iqCp2BTXhEwQaSUv1C8nWHdY8wh7gl3ufM8xenP8rXnvar2XeQQDhcHTSaLI5n8XFFQuZnK
sXpo9PBqRdTInlb2xMNcEoNb+FZ8IxMiQMLT0qJS9NGqg9vprGc7dk/bVVaL6OXsNAFmOarJpTOj
611NeHEy2iH6GLr1MexQnO3zekl7KCXEUNR53zqR6RPNPMGZnd3dQjRLX1mLjuFoi3fWN/iL85m+
nJdmH+omkPB5i4S1CjHU1/+jV7nTZ6K+cX8NXXTRFrqd3pcyKYtCMRNbEd4uZ1xWdGq8Y7cL9/XV
yJWGnSlqELnzQTRssdcYAPxZ5rKCiFprxOgtLS4kjYPJKQFg17lf8P6BavJV2ZrwxJYnQqOqfLiN
vjJ9IfjcAhPWi6Ndqe6v+8sxADIFl/TqombDiKh1q/lw45qFd67Imo0vqYd+4wNa0z0wQ7yr+vuG
ukJAInjkw/l+y1+DIQi+HLiiLN0e0/DEIC26VKKGo2o2Rer51LSVxnmi+wU0xVRlaQfBZpFkYAkl
LpDH8eTKIZfsmFFPE7ti7ufVL5d+XPJQk0YZ3z90PSypox+6leTSDt2T3MsmTY3TBqsodV7E/0yQ
DcAJjYYNJl7WXRC8cBHhJo8dERW+ZJyMfFFey6bDreXhWhibIHGicCZV2qCI2pxSExVbMgwGGCdv
LfhGcI+Cs2QlD7gNah93pYUAIkHgZLBdDjdR93Or+J0bDl65eMXPtqY+6iWrg3xAP61QbbN9iIrt
2z3TQFrr8u8JmRzue+kfoRcuw0kon0E1Gvx2uahAtzdXGFUfNWc99Ykz/m1tuAPYhgbNIOU4mfEv
pg2iCHr0/TuNbLedEZCLBQ6H9An6ZL9iACHwQVRDsDr+3MkHCaRMD3GOAByFL2UUkrOodMgvt9M5
hxk9ZBsk+bMZsbSHDvaGn2mFP+jGqGFB6RfpNnwBnG5AxUl/9icRSDSX5KzPfG0XsLJj24hQ2fGv
IWynce+8TEeEdwbdeB64WtBYOCHeGmuf76LJYnJZ9MM7OGWPno9JSRnLh5qDgXCyjynJAfknS682
uFx+JbrpM13kqYYT3eITYbT/v3AUmaNWVVhOT5WDGDgqmskXGmszg7oXDedM55sCQFjb2tcdsP/T
Fd72TG462qiBGcb4G+KHXAK3tzvnKLT9gY8qrdaImo8+wz4AwTcvY1+KL55PjdDBU3aLF6kJdEqS
/OKdQ/1FitcwdLUjXMb2+3oSuYpxCixiqfmhLL7CGS7Q4woiNCWvexYhlGmdEAt3slRGrepyhy4L
01UUh6AHIwhR/fM76LONdqgkstxVrFixAVwX/GdDrSSThz6PhM2wYJs31iqa4de1dDPW2JZHDa6H
sJACh+TVQty6KQsr54qHhnlFi5FcJqrnKdo/bf2IIPAnr5VXD9ACCytEAW4s2fQlCf+WLqUqE3vN
poVRHmdKKAvthFEzD7GghTftURdjKcg2j44I4d9vddUFTSxefI1PtbIe33WvWKIJuc1KwiOQeqLr
RgP4ljg1OvbjF6yKLQtvApsHVlm4UQfixIu2taBBvC+E8TE8n8ESX3eO82H/DlJPx5pZH6dThrTD
XJzZT0H3NJFLRGSepU29CJ6A6fRxAnRTiGK44SsLXqkSUKbgMNSJAvCPwsXGjaVS3ZFcKmyq4snX
X/Es9lYbsfQfnyFNLKrKOpvzwODFRj0CVTkTqplORXmXmUHkJ5tf0WgUUKROwqf95KKPYv+ImF/b
aWp7JZAiNy1cQ3V6Rw36CEhZjGT9dE9kcCigMHm+spNAjQ/48t/kQortt5VJV/bJnBkX/Rwh22Wj
uUELmbJMUfWmhpKM/0t2zLBQPj5pgmTX4dskOyUGaMW7eSLkCTqcrQiO9BzO5MLXgPJMBoHlpM77
NDXXkHk1+DsqYTu1wliDFzpsDIQKS2YDj4lmTzGd5h9fXh1ArtH557Zio45dCEWGj7XOtjtWDDR5
stHyyVpBodDeIsirU2F5V+U8ZK/7xK4spV5KltmPOgphPk4vOwRMvZZ/SxnycNjNBuTBizsyLEM6
H30wkqF46hD1VE0TZJnayq4cxQkkH6NbKIYwd5Ccb5nlijFO3zIr/LcBzNEo5+njHgKUpA1b1/iz
fquwTI0ttehVPIcog2C1AZ7DrB+02MrOAQ1DSBMruV4kUIUpnOTIb4qAiI4uxwF5vidxNZVcYdx9
twMAgq98BPcBoDHX+C8qdSAMNDFYfLCRMRz5Unj+7i1SaQiIF9266PV7ufYQzOWaPPI8tEex3jeS
VHP6eWv684FHaYsUP4yfZlLDyKJL2WVBr1FpT3JML9NAvAWV39aiV9kDnZLlI6VcIFRhjxvoLJeO
hAoG6+n7J77jhBJKyNzqaiuC24a34jf5aVFPBHoanW+HBTVTDvXrGTFj4B1wQojymaNuMlSH+Q5X
QnxDQb2B0qWGsHTDBg1JO6gK34mjoEtP8ChyEH7kh3AfRLkdLtxrv2/7hqyRluYrh1I0KMYk9rLd
LFLfg+GCJI/jR7ajBz66raPfzve1P91vBpbcWHkfzh5+o39uBXpr8NNcrixcOkcW0/425DY9mAbz
F7lsofi/20CLMkbTl7tXdM+IaayFZdkzLPotaRozCqtmYbo3WOL/gHw6rFalCm2LjYxi8QhWwpAa
LKHgtZ4YOHG3g/1fyr6KbzdAQFPIY7GLHxcmwesUVGmUKgAyPoKTp0Did/aa3QggeqHctdpbWIAS
2GgujLlj+4ffYpYRr8dpawh0YrvUPtWDk11yiIFl231kavWOcMeTohdwEOL6nsc4Dn0XmNAGlwUy
kjiWdJpsOaiXHD6/bxVXi19KgEJ48aMiQ3TfKOpHCpCaICi1C64ydc9hUWEZ9GSW9k4dYA1oN2P2
TQFM2BbUsc9wDcMMP/mc6CHCK1pS77aN1djR4YvLPxQrAIY3cTOFaFfgJBX10tggKP/ioDlfER+1
Llkll7E3jqBVHYAsIl4qIZza8mmTICVtVGtNDa5dYQQYTQEpk9QYBnmB6Rkjzq/9A3nuFg7fAgxg
TZz8w/HK/+daHCbNyHQuX+hTlFHeni7KvzhwQ+6g0zmsIAn9wGdkAHboZoxk0ST6Gnr3yt7Pq14I
39q1WN3/w7Cg8jQS22AZY68wuGoFgPxL93sISxtjsStlYq8ZOKVo52cDmQfK7FVhnYcH6SLL2tJJ
VaYQs52afEAcqr/1J3R00uKJWIsmfpaRRnXidIWeANp3IxvVBFzs0ues+q6h88wBXzpStNdZvGTa
79jqgXwBSdNMhhXKM4whX17ZR3WQFwznM6keVCt4qWObr/94Dgcpay37WVzn7NSmUlMobvFHMqJw
2QchPXLMSUeY/sUtxW1xTicGLHTxuSf7Mk2xfHYXqB5LChmPmfZn3FyksV68hIR7LwtZWY6y9fbL
oNiyzCCxuSX74OJDC5zuO5/fNzFrW2qaMcilpsw8ofG++rnAWSaurfvIA5ipSw81HSdj/jzaYVBA
0IQEC8jKKH6jrWVzU54fhVlR4wDuRu3NZxnJaQ2mU77yzknq8IQmMAWf2nUizI1OjOGTai0pDnXp
w1Pv4d+qfM4mfe9Z9klEYTMSb5UEcyzHxOEVNig/m/JWoVZ0Adk9jFpFk9h1t65rOKL2xw1pzKuA
kVV5CDu4KsOn2iVyKKB2VTGo+tRM27y4tWBCwz+5gW+/Sb8Wkt+2+V46qBFbIdpHdhvm4Cf6rq9e
ed9TD0m1bGTGvkRWACbOWYRMduAmKjNgZ9HLUGi7Y/eV/90/de8ibvfiYwoUhYYRtCd4w5WxWo6g
dbSLyB3GaYgSC5NBLF6DiitZpCunifzY3savmb9EtoXNd/2LGGOO7mUpf+U6VOc5ZbeTGClQ3Dsk
03Ukimq8W1EkQewmJ4qNuiD9TEPZRk8gFzhj3ZZ9bGg2NS8a1FueNSe7IK3uTTRzjf3nWshReVCL
GLpNpJ+LYF7flP+rt6NaF/473GAJcZJYNMOziJUzsQnCKPaRuWf3zhRsjZtotP/fPcl3E6o0uvfJ
NCcKqYbkdwHMd+zbQ8ZR2kZBJoNyV1XJX30LJ6370jShQlsl7CXuh0ntDmpVCM0ElmZpew/swfOt
sGIKY8O5gt8zftyA6pSy/v5Ou+ttyn/9+Zs6HqqB6giL6hIOZnQKuyaFWLxwUS0Led8Ce3eLfD20
dNILOq1q4Mb+8jvENaKYxcfL2FVvZr75MpgSc8fKQUp7zirVb8T0tBubu9Ant9h4uHn3YZ3gaTvr
zkGsx14qPD23SwSik6H5oDCrxX7vJ1QaVnPKvH8VLqIuL6B/kxWlHbLY6Mdd43sDVsxSkNW4Q4Jn
HXc76iGm7X4tkUbtTs6mR86pWpROtY+pREmw5g3EZ3sZa90vDrAoHTy/FqfTUtimLf5Q7t8xHEyL
F82XGXyBpS4KQv7o0kA09fukh2DC0iw1JN0T/8gyf4NA+K6VS/T2L4SwLlvbLMS/SxFxLfd0HPG2
aSu/eFmkEIH5hlfXZR5NvJeeyXHW73Arj646ZSEQHGyOaQn1Ob0rcc6dLui6TiDoaujQoZ4Rm2Ps
ImBxsqlh8BAwaCqG//1Wf7dMhjgapB9ggAkBQRfRW8ZY7mGFFG2w+abPtaw106gnoPfHNpg5FGoZ
oYvcKqoWNF+JfYztLqiuH+wZU0Xt18NQBTGU/4Vt4thqvBIAB6e3Xvqaz+YdHzDD4iJmCDC1cMIj
3RgZJgULs+zmcCBquyYfaWZkgF7JThMmM8+kDSM0qGXaRUytxFx++Gj3Fz+YNQDvqwGdLFC7N7ci
M4y4XkYznexMLi1OrUQlZESO7KuNMr9ZQsZgrVUMjFfzJr+lPMPWLqXbzmgW0JNOzjrDNiFKxKaO
DZYdCMblfy3Bflnv/tldNLa+HGAaQR0zkqInIcLgFqeK2iDgPDcQYc7acSIQVI8zFMVSCI2OKZIY
J4C5ClZ8jQDj1t37GgdaDvXeLua/Dg1wFF9ZuFtZs5GOiH8vA3EBbU1/Wig5ym2f6L7aonS4EwAP
1aTCla3ui6tUiU+N5qUi/ZEHr+Jya2281EsOyWaJYwCEyoHAs/fmRx1eqswTdH/MYWfeJyvlj88R
Mk7TVHawcZtX8XLjFMrXrABA6TaJJUWywFq0YqlFqD4QPqXLFauiPH7UhDx3SLRkZK9s+w5LUL1Y
gwuseh067GCKhLyEhe2tSa+JQ8Pj/rVlpw3X3eNCzpTEI5TD0CJ5CJvW0NMwjcU2/lFszdeI9D3a
rht5GY+Lis7AW4KNCpxEj8DxQ1DjalKLGO9GiQKQOmO5IFdyNLkKRcCwl4M0g2+5xlJHWdcKkTNh
xwELtDrbHQ7bPeoqV46RE7/XqPmvA9RL4N0OeNYm5mL1zsyqGzBmb8Igj31GRUoM016uOjnzQn3q
IgIGo38Swy2ELErI9PU6a5TKzHp78ormlsCFwOkxhwXXS6RKtuRmgiMWGqnFAqZ6BMQWRM99tJ3A
CmLVXQqoEJ4tH+0bKrMnnGeqoi5EiNGAPbi9SsnCclQS2Z2REQhB4CmluLggNBb5q6UMoWK2lYvX
IXw7hgHE9sVvlWHatezJja+2Q4ywo2EwVJr5UHS0U0Phhjjf1A6Ux5mevB+kvC1/i0STygVj4tL3
H+DBJUD4T3LmsvHViaFTavGqgO6hbecxlPPDhHzW5bFQIw4685rKxmiJs0qPx7Ip6sUoFY6iwptV
PhVnBFBtPgeKFSM3EypITyPcZyAIfHdxKIognx4wkjny3Yro3egFUL4cV5TaNa7YemnRKHna2Gb/
B4jVdDE1VHy/A5sBNYNfXL4WKwgqGdRDU+wdEV4U13AGNtVgqVss4KRmK/5lwz8vSEhcANhn96Z8
B81ftMQW5JtJcJxyfuGKoh7P1ZC7FyettmXdaIatLRQ4cWuR3P+JmLOpkgvhCwHcFs0yRfiXDSTA
3gyDbBYhLF59Tiuv5pCrBGUNxflKqFCKqIfrudWAh7ihwjjhH+eVbuUvPXV3eQthNovPLmGSFou9
pvbUkd5wYcteNiaJgy51W30TyuweA1mGU6rugFEpsrLN0Wiq+a99OtKp5S43LLAE63rd6CWa39AZ
pT8hN4+vaHWt0bN/rHbpWGpiOYKqiQWeagwtvjDKlQodpJrBT8bt8504ElbU8p4ar5kAIQS+dYNH
kg/OslKapfMq7W/pbELzPKw48s9Uj5dh7aCuoVTvLYPuXUYAhzF+Wo8xIgZlY4ZDkygrb3b/dm8Z
br3O3N1GKRN5DamWaYengyVcXCA5wP+LcKLABm4XKJjVSi1IQemPx1pz7kRe1DSZGEK6Eje002gc
ZV6g4e+O65V1grDXehbuNk6ccJKsx4UlTb+XCIjcCiIbWBE8MzYwbGAWsR6M3gSmYsBKe1xUlvt5
QqvgEHDp/FbRofGm9Y8QoORPGwfAQFUyqwir98t25i/lEkETHV4oVYJTjo6+fdzFe1oITiAbT726
X0BuD8k0OlfsIQ8abD7UV3ma4fNbVoY7/DSjOTd8KrnBE3PF0yari1lTru+/8rNv7Lw137RZWL7t
93UlFv4gRDt/33mru4Q/3QWeUbZGrNYgUmiFYn+BytdJWeUjzUOjaOJPkXSNgnVGClVGjws4Gpmc
BOcMzT4ZZG5M01T+K3aBke4q6WnwPvjgZwtDpkCqGOS5quS/gShgpqsGhP5SiOol0s/nx710FsS4
b9mW05kYHGrAjgHCOGU2m9tvT0TcnD4FXcXcPO9J7RkEdTkASCt8SMCsCZWRIZYCsd5wq5uL94Hh
gxiDeXNQBaMFMhw7tL2Hk6LHtjnhaJ0ejEXJTFZxoq9jP5dI/xzEW51vumNtW4VkKsnO2pNDpl8C
K4GPiSvKzw/K8En5DZ/hmFz1aAf9XSP08dXNTO1Ii5vJbgtV6P1gpDRIrDqMVPMCiOs+guuTVICF
rmHvUFkThh5I5WyD5GWDN6oIdu7yazFs8pNC4IOIlZYdcHSK5oIci5Mag7vIw5MEm5hHo9SgZVTy
zf2vRhGjRp/OBc/GEawgjsztt8x4UwL70XTn1OcMLz+AV54ZWC4klRLOnBnnNasB4o01YIuxMN32
JQcuYG01UAUDdoKCBW4LN1zE4NC6js+XgvQnE523GEHzMfnt9Q5C32Tzqey+voGCmRDuTQNCB3T2
zLqNT+kYZzj8Rul7Aku/gDKyNfmaFhtKvzbCKRjDtw07Hk8hzz+vIqsk5iqEJzN7LfWsec34FaY9
Vue1wMS0uhKDqzEUa+qpts0mV2guo2eQFH2sTLsBlluX1lnGd9e3pIAxcds5lY0quRTEBdBnG8Q8
RzCSn4R4Lc+pNUmgosQ3Z8Twvv/J0qpBCL5n0SsUJVj26ozJ6RAEkLwQLCagKDwizftVduDPe87R
QZz3cLY0iI48P9g8y+Xr7YEnCoRm/G6tCfBJJ5vbIB5QyacfP54s5GX9djFegktwjdC+U5w3WGZI
XF53jRUn4amFSLiFwrynHQDHjSj+RgGSTomRyIN307LxP6WNM196M4UsYZc1BZNA2TZQD+jb28XH
rDB8zoUEQx+2d9OeenWbFMh6CCz+hECb9UlAQHcwdMge8a6UCbB8CLPdF/aoumWqtZ7lvLbFzL72
F5hMOXNSXhAA9wOtfc1W9fYwko0rLlxKK980BzW4z/AKIkjlZYonfotccZeMI4GXcRSCb9+QJu8d
GrFwCd4a38EX1L2R/wFpz+09UYWg4VkxHmpYWVmYE3eI8TtkQAwG9iS/JHrajuFGorvVGUZlJ4op
TMjTFUNk3Y/IZYLAhy+FVrhyx86Hk/CKTOH5Qk5V7hQC4Et8SdMndfkxZ7cUz1OlU6NthwdElNj3
geyEt+P7zrPPm7Xm7C94wKuxrAVw2GWM6qPij7eP2UyKVNI5bl5TouSMnlZ5MSw++QnEvMAJcFJh
Wm+0zwG37cPEtvYMPEwrWE52Hwv60ToKWb9B8N3MfLeNlvj8bBZ5SvgJxHG/4sXZ6tstbSzw5Kwf
I2cFOv0yT8zDAIbPoeQi6OXW/yPBDf2JuEBYbdSiMcrv2nvBfJLS8iMyJXBBRZniC8tB3d4SpRuk
KgF2AEBliQz5bCZhuMS9fINka8ie+mlF9tVMZM/8uwzIGdwh96dOM/NgviCCTOcjLMqRWiNIACmW
V1neCdl0NEgDNd+aZOpTZx0im+yNPE8XPhX9E0wlnHW2zLSnO+A1IbmjisyROvoflIsqidG8frA6
9/X7LchhDKI+1Rt0cEi0J4GH21XB+tdrPZenklbnoUGj5yzKE+vCsnhOt2A5iYHjPq0VgliW/fmN
4NFQFe7hctDy1qNdNE9SRzplkPtDVH0dOKYh6QFfqN5pwCY9iWD2wcPsiIju/mM4o8+O9OK4pUFq
ZtCRpVosSs5Fj6v+oWtVpfmCfdsgYGbYqwS22URESvu60jM134V5ePmU1cNcrpumml+9EukkasSv
oA9+iqFj5Oq9biw+OT21D5lur7CTPNhZVu+IrBajCd+o0YC8Mqarct6GJunW91uum+yiaYyBXYbv
0e+r5AADfqrSdSPhxzkzF4Xr0Rdx+8mBzAUA048s/BJrYAgYmSOVMkpM42aLvva92AWfXh/CNBbK
52TOzDEt3xewze/VzIEDDBJaq5qmDCN2nfYWQgtUXCWmzC2HYNSCFLMP9Zc77asyGefSprNp9Z0c
oEK96xglyZBPqs7HKR0SxuNdCC9wNheP2cx8ovQJvRm0oScbddhEao2jzyeF+MNWImjZffewG66g
EP/hvDIbxY3vEIu4v+6i+krUihdp02lONoYzVL1sdBBPEHITzCgbTp8Q0bp4OZiTm6motPu/Wadn
l0VqWVIlGTlK/cwH7At364pB5m23jmNi541nquJRE+8j20aw+zVoMeGIfca1dkfW3KnTnF5InNLq
w+i9JpbR1DCineVp78U+BJrKYc51wLGpVGe8sDF5yQNF9/KJ5ayHLnGCHiyVxzQwJkUkRCj+qsBq
x/owuTWUySlKZ2Afo7m9blWTtblLdfD00ypNgf7GF9K7pPGHvg0VABlDU1fcGvAEppGinISdF/PC
d4cmLeuO5RtLXFuCVvaKMDTEqIuJ2oVqzMjbNsXuI0Y3Jg4weBlRISrQ0qX38vmLbjCBt2PWrlCj
87qpH/ItQCgdSdUrbvUmeuGOdm4zTqvCElDiAfp6k7lOW2FvaDNvQ9e0D0Get6ZDb3D7JEdvvV0B
bzKqNkX5QD8gTPvFweJt2emxmxwCNUYx73ZZbCbTkXP8bpXUFlvGwLiO//ulQ07oViE1hqztktM5
WSKAGzfAwH8Wu2wOnCVvnVZn4KfdDg6m7dmND4dY7XtGPiBTvK69H+XIRzr5Mu9hQZgaf7HzD/4j
RriuGghgQ0uaFMYI4o0pwp8j7WFA5/wnjvd7nwBwbzfE/1TNmLZV7WiqUi7CcmaANzSgbrFU184D
Z649TWpG36W9m3RfpT+5864PqWQBMUc+m3hDmaqLZjKnoKfo0aDshIMfUgQUiwK3/IGMbZClz/6z
L4DMG/lPJEN/2JSD2BqWkC06WkJ+2I7QecTA5/4lvbcsWXQhDws8a/ufeJl8iLJJ6rv1YwUOKMXK
fUS5VqTh7Q+q6dmOE8DaIZFEQ98iHvoh5w9Vo69T9gxWZP50HO51S4rjOZkN7tkuVA0HtTU3R2Tj
0KBO0WU2mujh8gpdUSOJVxcQb4OvfGwIUiF14P14D9RfLpo6EQvDc3ReU0TQBeEDHuoVGRvMNjaF
Aac1e7a3C0QeWr+IJuZB8RO3OD6y/9NsQLeGD4iCe1LSgoYSmGAhry0WfhCJ7s6tf7HigUSf2Kks
sKQSTBBarN98wEKVCgSaNjL0e5v72LddeYZEEFHNghCyAR7cb8ldNeQkNtsvVzjC1Mv0eUJas0AL
XR8+H0vyuTfOkFkoyKSZ9dGmL2FV8KCAbi3wHPQLzdOex62Vn4u083/BYOuBZbPQkBwoxwOI1q5C
C8I6vlJB5YPVVXIq/+2IRTzcFO1IiDYRKLTStLvDgOPEo/IfutRv/p6rlEfwMt5jCqoezdwYz1s5
xmVFgZKnLD//BRqw6sAsa2rEN0kIjwyQFrMIf5ekm5imq8SfQXV9vQ9R3ih9+rI9dO4E/9/jiX1R
1kGqqFyAhnMNe4CMF3OISzvqd3q+tjqPjrlIEsMVR1DHks0KpdWVtn94tZSytwNqMfsXyMpFulAC
KqyFfvJLHdrnNg1YAaneT7d/JROxYDpdEOsdaiUqUoinNHFU8l9UKUK1uAjWztsbXumBTnp+bxBP
9+N5rZq4FX0NsDS/EA6HAEnkJzKi5yqIk/uUl8oa3XOw7mMoSOsd4wSVW2pgoBnqdiqkUY9kN7ot
1tgF/FAZlhxqdCQL5lLMHpZBIDWsXGTJ/UDxR6nq0kKqq6QWNKNJdpyDfXtZur9OGiJUEkHAMM8g
y6SQXdjBN7tyHV2fyp5iVf+gq3T3ah1IxgsoIy4iZUAq26pG7TxzUkX/+JAn37zIN4uPVmYLYMZa
1NaoZiimtkqL9BUGBjSjKHNlQ5bHmSWiXTCWqzmejSvXGdZohZT/CDaPin40MyHpff5w/Ukn7jZ8
vMAnLl0gymgsaYQCdWfFENK1IG8gcZoBDPovEdjV+QDUbN3vir9+JYy78HhN34odaV6/casm0uiW
cWuH611utqqWmgExKMJgo+ExxgJyhwj636/l6aeR/P5PxHFAzTIhO+AWOPZ0oUuFhBsxR4J/B/19
Ng9XajOlD7FEnTx66iEG3VomW0p/VceOPBrT1eaAL3gdan7yY8di2yqVGPRS2FlR9Xmq1DWF2XEq
LJHe5wz3tZkUCnR83ERDIXHHssgIFlrwwcge99V8MQNkCxWhoIQDLFFFEhVYl8JjWue+PLyyOIHj
Hxt/t5fobR6nuNkf9Rreorohthsmp5U9WoE/fzUh3WLP/1mv+AUhJEGTnmUJ0eeKaNhwqd6o9NBr
97EFHxmAopj8o0SeMFKX0qONfegXxVv837aDgHgXLHFENUFY7EbkXxftGkzLgWjwkA1e2vu79IFH
GTbg7vobdbcHWDWRgrD2mR68x+kTP/hPsltfnZyxXxbAdcBUeSweInd1U7BZLMblQ/ZJ+sATfgQ3
9LT/h8IhD/QX4iIEW7rSjX7okBvM4tdnxvjoVoA6RGNQZRH5dx+IzxaBVwbggTGxdZ5emiWMmBVl
rprLnyIOOXvPwSQl9Fq6r1mfE5Sg2FF14n+O+h/2Qh+thiJalj9tmL8P2QhCcodwEl1p40r0vBqM
/MJ3T+RpYq02AnlrYnFKVw/kZe0UaZUlzqRwPQq/ixVz2eFlu8g6RPp+kqO5HoGTA1NbxvRwvYah
Ttb+ZicgijCvryNeVyEhJZVq8thHif+EcfYPc+rn7oGuUnqLYk1cI2l4pJ6q1CMG10slFBhCIz9Y
mQ5j6F83B+g8TezybAVFLuXI49ErPg6kZQ7uJFdzHm9yBJxdSMfVmhnqV4Tyemu3jkA7VPLRTfqP
CGQnA9MmSNVmEKKC+BlC7dqEukjM7ZX5hi8GzceqkeM8/TaMbmCYJ1agyRjMOHMuH9FUtX6HoccD
05LOucEdPaHAGaBJN3nUthTVPyq8ZiTVo0w0CFStEMgw/sPGGKOIrUP4Czllm8UhNGyYwD/uYJUt
ckcuWEAbDTm5ChcMsr9LxPr5CUrclvCR3kDb6BQN/I8J/bLmNicgn2gqZU/4JvR6jLKgY4rdtE8g
iYBcc0Cl/T8K5aGWcPSopXDcwhX2/DkpdrGCN9cWqkkgEB5t8Ci7Z+tVjgo9Y6TCEeph4IbHvnpD
a+EZJWHsAnFXpN6i6Kn7SnKszzzpuk0soJSUMS7nPXrcLBaZmMSA/e8kuUVl4jCzTPbUT3a0FlQe
G5fZPyLL/TPkD+XBdHTIsul0LWnFB+mWQKnlbpkHvspdPdm/G9F8hNa7TgRf/4p+EZfB8NFAWFjX
FizRhtHLPxAzaDMIG8JM3X9M658LCG/KhOiT5gLCsNBcJhzymaZDID2iI8t+QdDu6XjIHMJufAYL
cUqbpDzOfM+Rav2JOU2NFoDXNMF5aTEZWtmHL3qVgZ5nQvLp+L/iEheSnxX2p4DjjZXDHvAnpBup
nXoWuHRdM2YeXW+vb6V+iCkKEMjBfsX4uQxxFOJIfkbqI3MwsSSdO9PXpKTIg+NQtdK03jzwACRH
jw2VoJiBncYCx28n0lZ1EJwpNFlvRQ2DN/L2L3v8QxwSIgwOfJ59KHkV/wUCY8YzY6+YS2wh7VZt
cyzeiZfTdtc3umcZSbAUTBhDgU6hIBkqIRtdtvABPC3jVi/W9Vb8yd710Im1tdfSiI4oRy4/eCC5
i1XSJvdF+1C5RFTNX0FsqFOTE2XlUk8sj3l3w9A1YNJuGXBWMhIbAhBeZYRBTEOWqgxdbYh5UQzK
gdXb0yzM1IQE2XSQnoaVUmzawlZ2cQfd9EIZTC/vJjOVBiU7vstuDbJnY02uA3rbDcSSmaiDCD6o
Q/Ctda8watj3PBjsQT8jOSTmLj+bAULe//8PkTAcWCGqnMlRM/Z3rUXobjLctk3rgGmzBEaIi7dm
rgYZhYbXg/HLjXBN3uO81JZOfpJFmMBWBIn/9+GX5697A5oDk7fba731d62xXNgsGpxRD8LbxcUD
2QZk5tR9tl6s5L8LaxUzr50WLbgGv9wVuG9h5qVGHVtPIp09obQ8KwSLe7uPyY2q2MYTflnevYLD
g8UmNVOy9+vMEMInCyQFCBwaaf+m1Y5N8S1YkIinfXjGLSDwpjnebyGRfusaKYAtwWPbi85nqqBD
YQTg9diFR6yBX5L2Bvy5tdf1/RsxynJUadZCWg8KfVRcGU/ap3xs+zrsP1Iu2i0gKNRfFRUZWaj3
JlxtUFTwywwkMxoDIg8MS6p6FhhfssAM4So2sWkYFSjDGzZvf745bBlXCGLOJPHqUAUZNAPkYQ15
gkBwS+5Ft9bdcRBDz4Bqf5zeSxpxBK6ZAa33CmClJswG/6fngPIT6iwgVy9Yc/tvHdcDDtnfqlq+
AjoBVR3rP9QqBQkm4WfbkIU9+pvAt5W4uj6eAdTBnA+k8bAkZKdrJYM9cbc/REa0xfOIWQB1lEFa
WjSRtrF8RsncuS9JzYWMD1u1HdID/q3gIuZV6EEB/j30S21dkvNglm4GEwEFZDM8WUEGP7OwnknN
llqIX0gzK5YC9jm6h7xPOdXzhUNWbBiDDwFuNkeWwS7ISQLMx1LPj/bui2Mf4j+DPp2eiF0qoh6P
7JXlP3iqOSK7NfpBs7sXDSjB7DtwejEhZw/2vuRs0bHvv74rNoKWVhw8UiO8fbrXozHMBmJY2B/A
VLo/QRFCD/Qh1807Iv3O9P/daZ7fRsk9L5rFXtdXbb13rX2EuLDhPnOE05eaO89NQTAYfgsQGvz+
b2QHcTHDpVS/W5iTBeNjlnTKzFgwhqKBoSDjVrqvn3ouubKHmYLYvhjUUZhdrzYoRyqmQsoo65gp
pTEfl6KcporlrpljXLbQtj4MfYEngAW4EONU6rvZ3PrUynBWi4ktTlaEyiJVcRLtAIv4Kerp4+Z1
WRx71UiUUvrPuEyrYz1SUpa830toVWPgZOO9E2w8BJhCNreIDdVB4xvGFkyNoTqlsvPhSUAZhwqv
JtLowqIB/7bsGrBgOwE4SZD0Dk4PVxwa9qBHMQZ31/CTr8mAT4jdeGHO6sueBNzSE4Qiuaz2BVBk
BCePseJSBvpWBMAoFVEtmYToxaobyLWvZdhZmeA7J3P1ONUEwi3VDs/PiuujuhNCdhjGMYaP1pwz
h6zroQgpd3bns62UV0nJwGK4B9H/WhGNTsh5oUAnRPXnvUYJBH8bNP2bIhT5wxoA9pbrAbJwIzSn
ObLP0xR3kvtmHBXfiyFm29cX6Xz40ufYazebWR9BIuISqq40xenudhXQFyX7ojFKDCZ5zyxcawrs
4huIx+9krGfZhMEA+vIRz9UZaqIyJMSX7Nqe0qTQ1Ss3eHd9SWb9rMOG7xCJx7rb3E6RFZJ+mdQj
0Ud8rtA+XG2onhhfNWt9BfcaqGUhy/qUyTxe95ezCcY/3Jojw2FNO44NcWAOfkYC8fTI/rt1o6mG
1KuinUG8rOjtM2WEMyvwzKUkJ3tsPyXL5DFtbKmZX+03CWbo0r53ha+ua0p2kNa/Wkkiv1e4LEoH
7lXCFz9Uw346gW1qFezUJKWh+KPoSUZpcQUnNCMooFrHQV3hViGQ55OXcbspO5cFjxYZVrIF+zge
o8Nr1Id0KHu7tFHgaxY/YRoSP2uKTpwzO0rDIypMn7CFHk2a79nZnYIPQfwrkEH7k+HO98iPXU5a
kfrNtlQc13ejxNrihQkqUudSXYCIGZ+fZNlGnXRFz7ZSSep6Fz6N3SxlrzASqawZuh/oremy3YHL
C4nb0MD7H8HzY1GqnQt7ey3LP94G92oUu9SwTt+TNkwqE+VHZHQuVF+dKBkdZ/C4TLQgzSCtToIp
GXlh5iwiFTXi0xs76OVc52+b4pEDPsJLCZgv35cydW8TBlAppEShOiDDPWx+prjUE4XvZbfmt9C8
4zZR8bwYe3eKrhgCeKV3RiEYn/NGHgTf4GqLAx/Ag9bPQktje+vB8yjYy9lKlcNrgrkNj7tRWRSq
3nVVcH4G9F3M/tw74jG4uy5tUmQ1UkP9fveHqgiricvfOX3At479OGuda52eYoaagg0k9eFbZzeI
iPh3Xey+0dknuOC4im2eNtFJ8es5OTbfdNCqSTnkNgrKQQAb6Elh7Lg9AJQ7L/IPcEeXXhJFE/Gf
neuZIS5NX8BuSpEjFmEvbRnKe2JRa5keiYP6aD7c4D5PmKX3+Q2YBO3nf0FnAIF5G4kgXXsZLGFP
9qztdwbrCAqgzWV+A43gCzLuxQqQYnPTM6nyaksWGP2eBF6BJ90Cqc9cmNP2t7kU/JQSeSoZYvDH
+FaxlaL4/LzIjHJ5ZcdPjd6RssPw7f38U56gYiF11cW6x0S9SgG5xsz4VhHMnT4Vk6CHRi5T9nT+
r4Ax+RCrKJPsuPtgEdZLGtaBan/vzR53MrL2uGu+K+uxDsQiCkQHxEL9vTHZJluUSKX51Tt2V1gO
I3pY5zSAfk7eSURB+9AAKH7tJG7mBMPDcSBagmoSfxSZNIbYYr5CMLxPdbWvnyIbFg+J0/lGa+jz
4qI5OPJHt7uuY5p44jjfFBdAW/pEBa/WP6wVy7gVmCXBiIkIkV/9o8bp6bBSjv4hiy/SgdaHyGlD
WSXfUtf8jxeSABSr08HaPfiM4BsHj1ETUrMd6iLhYIcAPkU4xmYwaPDflVCKKMhwB1DYuEFkyuCV
Wm6K8aEPldww4tqmHlyT/vyf6AgXiF5HArdlDjQ2t9klbRGUguhewq49RFCy9GuGefTEBMunjia2
oG3DDHU+6hNo7A/ToM0Sqv8W/ETQf8qYRxnbSXmaza0YLHbbJXG6t+hevhqTDfCc1Sgj4+VBxgRB
9nXgJ/3T3zsmj3mzJaTFx6LS452eUWQ/MnNJzegswEsMUltbPH46kQEE8XDfdddWA8UALjx60ePN
eCkLwMkGiPCaR7y+FDOwLWr4kqO9CUwTKDhQbQ/RU4sRtOSqPQo6xQuv/4q9Gm20tVQXy34xcXsv
Zsizr+Q9G42FkfnMMHSwhnb9lMlp8WrcV4FPQpkIUNqvmqa5yLSvV2aIR69rsr7B3bit0vnJRwcK
t28GQkKQ+ylNPKN+dNXpa90DF8w8MmIER1LlIeNelrNq3iomYEPSq84mBqIreNfMmlaAY5EOwc0a
Quk7B1/+7e1gXuYcrifhUzr9HOZ5MC8uc7Ex95X732lhPjdMeFVkQlzWnYp6Xt0JHCe8DwsqPZXO
OzeMZaHqoktyeeKU31QFFUBt80Td2dJsYwd7bjg7TjwRj1l7aP4gFb4mc6/5+EAMD1du+0+eAUAX
nIh053O9jj36Fb1B0OT3Ga34v82PefoV1D7J9GigM6wNHI9sR8skk3pIgsecbGWbfEJMsk5RRTBc
lYm56gpIruQIXD3Ll0RN8kt5v96cFNLuOmdGCrr+/sMlgGKWqkDLCKozd68U20wbjfShb5Pt6Vv3
v9cvTNtcbN0+Zw7iQTGMALshDY7pFSLpN6EwXw4kOzOhonQ0i5l0J6e66xrlDRxKetraPeNruWOn
VqGa84W+7BKRwzqByPJhaOosKP+UKWhr4VX9YvCq0nXBtrjc44/nh0OiLIzNQ2HwJJEWZtb4tjW4
cEf65ui43I/Mii5IlpSOZ5T2V2xWcTnALKL81bqYo4sFJlYV/rGnt1aXCU4MNMRIwQI1aRcG4nQ0
/BWfA/8Dvm4BBSVZcnwPsOQGXWM+z2U5LDgAYBghN6OYl8KQf8s5bnT/vsmpn5FtJ+IbBJBL/Cth
+8jUmNZfdurYMdI/8zl56ySPnTiiGzYbIuB+ZxbYrTdmpQcTFiAxpMzXpTIxpLKU7RHcWpRwzLBA
rEchDovbe52P2g1HxlF8DK/KiijGhcTsl9q2/mI+d/qr2ev+FvWo6cu8F9doiz1GoepQt6XTV8Xy
tR/x72QWFVhcNNayorokmMlQzYTHh0hrJfsVRrMJ4YZ/ctWIMLnCTe1ym5IwkrJBrEu+d0Ei2f1e
KwfZNiQeX7+q7O8XAjNRROn+GZ3NN/nvv6FgD683ztUK9C4V59igItC4UHE6jwH74aGIu+u6O9Sr
g+gF5aNSzRF5gll79UvNGZ3rReyYiUaFHiHNpbnRpaHBXsd3uGApjRPjQf22btJBLasP9R8vNx+Q
ApN62InGoceuTMkRsyVTytU9ChziKPRZDaVROJ5B6tw/3GbHGMhN1ZjLlTHASclEJVOVwDYkzxfQ
BtE9FJur0L1ErtCbOK9SvkLJrs3s3/+bmmrSUWX6hx8Klg79J3IGiY/MYByUk9byWlBjkwZnVpTa
RCTkw2h2ShnDt0avtLIOZeDFDqW9twuQVkA7/ZkZHNnMbyQysl27toYBVs4RK5K/BzRDA0e/q1dG
kpcD3H51TJx43C3qH0ipkzLZZ5Ka6uyc5Z6lZOEVFRUTfIdCZvX5fj2cD9Kn+h1XYH0UL+ovqmdR
4NuBRF69JOhPGjUa/wfAjsh4hVPzQPrtLXstetwxikFs3bsWCiB/6CuRtDBIneqbUVMmM0rsuCGX
kXnFuPf3wj8+Lh6cBlhOM92f4bALK49lwpjReo9vGA0Ig9BJN9qOhPyTAP8BQpnQVWEJrvAXUOuM
EcEeQKQQmXCRZCih8oXHTeZBwsa7Rj3w4eGMkj6bLb4KhtsqAUm/zDSlBuLTZ/DbbhS7bTPS40eU
/DVFab2XQJhMt0BDi0+j/ryvir066FbxA4j2c9Z/MRCpxrP0vHFGPxnM3dgSChfHb0OoInrdOWKr
u0BFojy/MuRDMNy/Ln0WXgEQjJ7ye2sxoT0N5GfjstyRLONuzqKibFS/+vcgAnh2DHE8UQtFNNL0
PpmBv+kgrqUBO/g2+CWDqft2YXdPNA477W2X/pvYs5DYLQnw6qKzqf9Pmr8lo/1CQD8VIAyJKpy/
4PoqbwNhHatZF0wZGZmDKIzjZ1EVRSlEteOUdDncvtYxmcrCgVgjMfPVfKnoPCXJYu/9PPI1Agbd
IOCR/fMlT7cMWwcw9XlWkjgrtumbkVcJYi/H3134wmXlW5Iooq7gB/h/1c+vQIimq2PiigjEUR33
OQknY2FBj777hMViu9xeRJZIPQmNpCSpNv7YWq4p1//17TjKtvSkeRx7J+xyzcmCcJRdZtG90ZnL
VIadHDJrMlRu6+UX1rQpxAeQjZY9c63y+SVbm4uRDt7h2OdEzmHGJZ7JHtDuNcxGJPrBjgD9TqtS
LJCrUbUwSF319RILWHFkfZXddNX/2sV50sFuCkPH7A2EXTIu5BFcWcskGNZhTnI0uKudh0SGeoOA
c1FVCyqylgN9rHAIsRmZXrXv2+OFI0hJex6wdMA7/JWuu52Mcs3/dB5CyZXlRJdCYHXVkY43SYY5
vSy9jXaqfKwMpociMjBiKfHrDw3RrZ2hOr2FUKWUS0BNf8twQr/gbyc8us5nvLb09G1BiQFkvPJM
r2psNWuB3SULAFbLWa5PpWBTZ9vW7Dr7Ks+DlFYehlm+jMAS76OvAeyzGwshHmvFS3rT8N5ev/g9
PonDZpv2oFqE5KPV23VwJM91Ow1nuOwV4lcibDj0HKWEjGEYwnTCq9gou2eJJISrPxN4DNNV/DlC
xwNh3OtyZg30lZZSyyBYPR+nus53evY91D28OoNmPiEJjVQljjT3ZJ7dWSAqA0qGN2GlA/CR/eOo
OYFA0PZ13rQZkgSN31wem2Q6teeR2uRTKa2m42zoxk9kChZsMOC6F+82fDyI7ABqUsMGtF9KqqZG
4Ig+03vXubiUMw8ioZn6v1LPAp1K+DKpQjguTjImXXuDuARIyUE4OJEUdwwjfHYECMpBAs2z85Pk
ilzBIpNtllitBo2d4JYEW+N2pXCBg2NWksiqRXW9vAPvUk3vr/YjliS3ocy6Bmvu1eKN2NWeN8gD
jR1r6gCPbrzNfD3izlRJaonuR0fb1zbtPZv67MAYVMS6T5wqFbf7uQavfs++6hWXY+NslnFriDbH
PlZYOJoNv6QtHzynG33LQEcMQ614CthXIfuUs6mot3owmhD7RGjC/UJKshG9UYXhgjHsT4aiGEfH
ZLYjqHo+FaDLC4DZRzaBiqMyn+CBrvZJEIbuPiZ1z6ieMst2Quia56QP19zhGU0iGod37WMOpB9g
xhC7pJ+d8ciVsrxx6xYMUEjT/ew+A2urSK3J/iseIRO7MuiM78t2/2uenkQ3Hyne+z4x49oIJo2Q
WOdxrHW1uuWYleXVD/g2wjVgEpUIznZUg3Bdt6nruwGL/+cZkjU6/ZB+XzrCIVBAS1B61k3AZFCW
mra2Zu6sBwMQBelK9smURm1pcIPnOBbV5jk0iQEfh8YP+RLRQq/kzZ3sP3Wh6KbKMnQsIT+svVAe
ltNEHK9w5L1ho//fWfxSePTP8J48fBNg+SM9EuIx+5S0dDTG9zIhersKL0O+zcUrByNZDVcIANyb
aMspyfLOmJ2oi8OxcxvJqL1Ir3xGB5my1XMYJenhkyk6JnetZYQeSKUB350oUABRtJUgGjsQobqW
0qa33Jz2fGHhIfxaszzuepUrLdS2FZuVCXchlo+Ca1Mk101xiWoPVYE1LgQ34a3mX0mCoWxsWONb
W+TTUKlQWHXyaEWEhgTdFvBn5Oy5fO+j3IbgQ7G9Ke1MLjsyy/EAvd5L/a5EgsxQjEELdhn2JMOB
Kio/1R0CwLUfN4AvfPwtHcEQTJU5l3UTGDQs7Wk+/Fjf5/K3W/VrtLNGy3o+3WA73JbIcLbxqod9
5qd9/7dRNiR3d8+xnwcZXt5UyXvBMB2BaNdKNeCkkIOdSiv3/EL17tm9QI9gaZGtSv3w7uQ1uQt1
LfX1AozrHSePayMA2mx2v6RidHQfsG71w8Fh4v5V0swo1hhYjFotv/cHYZO/HyySwAfLwLtlWaQ2
OLmneBOGlMPisRIEAvX+ZAY9Llpnv2vERNBzw9Jbo0wW97A0nhAtbCMcn72iAlVMKNBGKnxZNYt4
z3X4VzymsOAHjBV8zPz54Hd9GUn6Q06+d/o/WQ9ZfwalEXpC4oquM+AmmV9VOjnwlwZHvJtDNUrw
mj+TZPuAn2Yb4VbikVNnoHFnimUbvhHM9gEZl9U+THUuMJB72sBh/arns49l6G/TJCfHbZKU6Xge
DBoPWQjf2+ukY7ChLQ5T7HhpfcOG0IU/kIGNVPHKin81tN2hIJ4GgkQ5jqfdT5cY4UnSnmSLBpVs
7a4MemSUKpT42MQsPigZ3H0z3tlD4uqYOb6VMJ5dfEER779W+q9/zrzYeI1i9EvxDyrYQD1tH/KM
C3U4YME3dIak27t1KANGy6AdF42vy7RrSLzp7FtEcl0a6PRcoViyO3cYbE9a4FdXfroCjVFVzK4J
koNYjYifX1PlAQZ0SF3Qe4hIlElht59jxRB+WxLoQhI7RMjc6Ev+ar4mJ0p18UvfSHUhrg7yj6Gz
iaaZ2fhU6rn06oubF8WPfr5W4dAOz4u3c5vayhpmgfGO63J5VwNL4mMHv63UK5LPGcsq5t/1i/wn
Z8BEC7Fq++AG6flfhsdM04FYweqoADumBr9SB9zCeETlNkUOH4drWleVLG3KQ4sKkX+TUzR0MNFR
IG9jV+ZGKiFVSko/P8P50Q5MkswHaW87tX3tVPOy+XPCPr/X4WU1rCDjYlsTdPa5X2Ncgt8XNplU
BXfHkmrxpmc0FzsjIy9o+T7ohl1pl/idmtAvgeRAgvO7tTvoBnm5k8H5b+AhcWoimPrlCznqo8oN
Bcr2T6q+Xplyh3XIDbi0dj4X6IE0Jte6QOYf1oCCCRt16sG8jN/LnnSgkZ+X0LIRMw38dzf9hsTa
QcRofianCkDIApjYKXR/Y3S/Jpxa0ldivh7kFmVwqNelrSF9k0iBYhDbBUUrC9BexW4lvG2H2383
rn7TpC2y5AAwd2FcPC5333IMrnEGiHybmoCIUeSO0akxLCsuzxpFxND0eUX1TvKpEhqJCPf5Wk2h
1BYqh/Kux7joDtgbUMTenLjJhqDmwAB+o7IrGH9A6HAiqwQVnbVo24bAoJteBrln4oWtCA3k1VyY
FaQ04SJ/kRJRNsz6jT04LAn5ZaXkX+0jqusdflCprdQWks9Y6tBSfDHUZPLxNLIKNGiHL9loE8Il
FZGHyVxiHDD/uOR1yCPi/uNQJ6/I0m4PGn0dwBG1SSt9aKkCLSjq9whVumuLBYLxcy1VdlLoMtWM
b0GURyThYgNVPycAxZjj1uBOzyLivutAHab4xroDwJJbo8u4mppgqMp18IpZNUaEohw1vln+9ebu
54+wIg7ddJOomGs0cO+dMeMNBXtzTQ5E0uw9JYZef1ZuIvNDTKEAGCJfw+6PdIPhvKqdgG4wFRS6
5+lkqyUvlcyHv6UD24mfLNCHWf3wo72xq4f4QMyeySLdjrELpIvXGgOm5z2N43LhDwhlIu57UUjN
geoJlYWkXbRoXwoTn03icfy5F9osVLQTPdyGfumyHTk/3lTBKOvj+ljol2iC7s4GFeu15OBO1D6q
SjNyAwtgbvFloRVmgkTV9hPiufHoolwd3CLMB8n99ShThI/p2hZ5tYCPNSF+8VszqWiadoGtCGag
6fgwj4T14Ip9UV/JluD6PDwdDPBGTe48KQOPw+fvxz2PKrF6EUQJGWlMsxUVKJyPTl1rKjGLSIRc
TFxpWOfgulOM5UeH8dCI9qSywF9LzO5d+zw2ZQOnsr+sqIMNyN35ArqZIlgtTG8Arh+kZtrhPHVt
WLkd8TTH0gSQfiILGp3sLGMyc7oUb1G3crVOSJotauOvCtdKfujpzZxJEhMXfnlf23zm/d9zda5C
2GoASzvAMnJGg5/jb5sY+mgZeBQ7nkmYctMNRVR5DvPie64TymEFSdkYei1FjNC84uX1xVI47FBH
IlJKiPWjMZIKu37PMmSft+NbZfQXe/zQKSQyvTqKeOXu4S3rAmrD02hotMDX5QV8GR4Ko3zUQLNE
fDaUX87cRnwXvjRccMiIWR6YJ+G/nDK+Kocwnftn7LVvCwXWSRzhgHAdaIhYwoeEw/sR6lFZ1y67
eNY8dAwSi62B5ZJHi4QRybQN0F6/Erz3Nv8Fu1PdC6ls2Yzc5rrG4cYVOfmc2b+Li/z1Zl9QNjKu
VdnPG4RgeqSwnEmHUAdNHt3KqFhtctaaVtiS2K9LpgOVoD2HmAhqakAinNv1Y6Zf9i3Jj99fE9Sl
BiLyRiiDf0DBUnIG0Pf/xS3CceiNgrNqy+LtvH0Q4wNEiF3cUQbhsYyoF+BqKbZgiUJLhZkRfvoA
wKaI9X9JAI57rV1IASoPNN+bBYExf+HLN89/EzskFqvm4DhcM1G75ZO4I7FijMxWMGB79JSbIu9p
jhJSfGiXpXDPtpwzgMTs1qFloJ7boH50B8EZhpsdZvsAhFG81kaf4alEYkaxVbSBbUWwTh/FTasD
Tzy8u19I41Cly+n1dfb/Cp1VB+TppplaX/YiieVYgNhcz1A9ZwhjuRu5FE5Y+LGECHG+HHvV2BAx
x3VRp7QnNHYcVwTVFzkhzrBQMTV5u5v4Sl82xo67yFUnIru5oPbN+bT+jxpdlbQIlPJJC6IHUPvw
FE2UJTiRfzVbhmIRZ+carfP0zIt0b2W5ilpem0tO0ZN45gfl95YO7hQzJqcrmOCyFD0dj7NGd0W4
efcbsmO0CJFFxpnaFaP80/q94tY5ZVbyjzg5Po4lsmPMaFpHZHzMhjR/oVGNaZ6zAcO8wGSupd8T
/8f4hlSoJLf2pBV3Vx7ZUA7z0HTZM6Qp68G7074EBNiLByVnaForWZzwaZl9mN6AbXXemTkxcrH/
mtG/CPjO/tfsRk2f7q8qxcdDSOMdjACoj8seu+m2TsoSH3FXVggMAuHNLYvRH667ht5VtUNBO05Q
Nz65nztmAZX821TBs59ZyEo6i1VEHUa91OSje4IKfTaU3uAUSC29J7aEgPvkQ9CxwClXdw1ip0ZT
FPOLYehuUml+dKbkt2NaCW1ZtNtoGP6qtyZY0iA2vtnTiXIksbPp8OQ0qAosXezTmuk+r+ixX7Y+
xBZ/IOt0DZqFbpBlvYj9WGvQ2hDRjvPIecsGIX+SZFFx4mBHWkK660aO/PpG60lyxfCQ8qdr+7Vo
Eh9gkZ/s9hCClxe88V6dEm3lvNFI7wOhIgP1ewYyaMlbTKl/ZCBsG1aPDX5JsJ6X3HvadA/kU1Ox
Oi1gH6XVfaflBXvJ9pedvbqnXb33xiP49ukVlK/j+KMPggoGukD+gV7wFKWQSC/lJtQCQh9HK/2/
VfPl9RFZe+o0v3sx1f/LSk8jrRVSNdzqiYUbaitkP0LLe3S30tS7ykiK0PpF2N22QfTsG2HomuHL
aVJ2iDKRORYgL+Xgy0q+qlDAhWpzAnP3qfvL2W+eVOEBTvcfvp/4eGeu0NNRSD8x4CEtZeYlMbVO
E6CmL7Og2DN8plFkUFKYwg/6ekgPNcP2jOuD4vXMvnUZ+rQ91nf9uJCHfhSy2N4NmhPAZkIceQkk
RboEzHZEmOdfdGa51VSbOr3LyMcDrikAUPvffj20EWw3nE+L+JMTSAKKEvTtSRKN2R1jq9ZQE+qz
LRqlkM9alpdWN80pzI2uOpTS4az5tNTbCfmcf5QwdEFsBd4GLuEKaMyO7cYUZcvnlWVtR28Nr4xP
BT1jfVFfXqbOOtvs68b4gUYQhQTPYibuzalVM/442L5qBw1nOzWmU7PZTHw++Itz/QSw3ameUYuv
eNyK0Obg9ba2yy7sGG+IIH4YORc+rk7Zs31wt+5fF+EVVr1Re+0WzGmubriYvfGup0iREs/Kpy+k
ls1+eKNf87WQT9XS/JesJGBEm4ibJIBaRegT8FcTBMAdsli8aN0JGQFbbk/nG7fJI5xKSWUlMsiF
osGw8w+lhIKPIv3Mn2NQmQTAlGy49S+ygrEDGiRqeyXrKIc8KX/O71e64z0aaaRPkCqeVwlMoJZb
bxL+Fzb4v3R/03RguHW8R82rLwWgoM+emkR7Cwa2gBJn9djazOE6CFSCdTKHSVX5Dzco9ONTrGqr
SioZREyIcCKINqzsHTZfNRrQRwIismbK4MQS4jDfYU3E8EHykl352O8iK6GGFtKjv3XCwnj1cIBO
DuxoJmVm1BCkgyDNEpUvyXFRMnAd8gJugndyH7lKxlIjUG9AQr5KFRBiek0PuKo5D/OtplaYTALg
IpJ1x+H3pHTxG6zvBktm5iAtY3+A0JgOzsEDIA/XAtNWOe1MfLoenPrpp+ucAwVOFWmRduPi2dra
LuUqipeqIsRQbwaMEzq9dAAbCDuufV9LfkyZoCEbZ+LUNcC4twIOemLRHGNwshblH2uOwWJ5QTZV
BemtOEjKO5H/7ONrVLvaesQ2yvBUzsgsF0dohI/GyWC9u6J5WaeJ6pOE6RMEEGzGnozU5d7idQ1e
yEumB1MkcLAdb7/BcFhdt1BnF9/6OhJ6p5PnkgQTxo4HVWO/iWfpl0D7HiAjC7gZL7smqrOy6EgA
LazxyBvyheTeCs8ceRhs2o8jrJ9qphJinlDVsTr8lrAsm/Rt4EqnEbCXu2bBUCxEqx0xJ3fPBPWZ
7YAeZ/OWbDDPf1XfrjK98bzyvWE867hr4/nccUoU3FGrzu2sxaI/+pqnncaaDehKrAZfcB5Hsj12
G43Ggx2DCXUEO+b60GJ7b4Ko9nDGTPg6VIhEpWXsI2+ivgDNDGVFa5NhYZyUePjhnX0Sfelc3ofD
456JZKb+B5RDsCrfdlCWwbTrqf79ZJpdbMnB44oUUnwC4rfdzVTuY5fmbcbyTbp9k9UkEvHR9Ape
HG8IrJQXZi6Led8hjE0Oh4rcHc7ImdTAVeIsssNeXFuYnZnLqgnA0raaTRQzI3cJso4O3nFpWupU
OFBMXb61ioj9vfY0L+2W4tI/8I2sCRfmIgR83GQh450VP79CGiE9NI13CLd7+M/V2xjlbzAPIGdM
yJFMg5+K3tjUZdOpuZ6pc/5lioC/h+3PwQ4y5RuUxaBstSgJ5+CeAmMyEGaCehAysr3/wc+9ukVC
/2S/TQTOo/BSCoM0q4KtFIme2Vna6LiUgWjpZpwvfM8fDmTKdNvx1jPAr+iLb2F59QjnKruBpcfH
WmXh9vOowq7eOsvGSKzgT6k4s6IgjGA1v+CeewrauErzZKoJejyXDE/RnWve08TvuItcvjNDeXh7
MmauzIROl2ntsImTgVFvtH7QAZMBj08pGBz+FlMc+uXhNfew0ra3V/3AczSS90qyltMgVxBDbghI
iW2VZITJLXjy3puTqARkdymtNarBpmlvbo/x6naH0Sa4fI/iUSZBbWxMaMdYQLNjERxjPLSxIgHn
eheKWMgeVajFkAeXr4xsX+Dt2Uj7HzQKiwg9eZv/2mijt/utzB8EHiERce36OlrKQdEooWootaRB
X85wCRvdevsEDK9Y5bDZiEgLjc9e7m1TRPGJq5bo0M0hpP9xHg9AW//uvRG2R9oYP1DEdu+qhi9r
BDc9fzz+BkiEyhnXSgEIpdD9Lj+ZQ1aiMUiUE+ZWAR5CzqcP0VVOBi7KlrK0zZmyJ1CRuBURXWQ9
w7VI4DKgUNzp2+tae5S/ChLEk1GaKnvtSEVLnK18oWT6V9sO1p3IfgLSMUwG+4Mn+K3HJ6TmsXIL
lIOE+p0PpqOmzXe0N+D5H2/Vz6Mp6Z/RvhLmuvihiLAKxxbhSlJDeuS3b/2gQRZAOpfyXRhahwsD
MfMsDQ14+voEq9MeMvhpy0et++ogcJbCeNmXf/oZT1o4uI9h5pQi+B1owlj4dztbA7zqL6kR9yDI
y0ky4qw88vaSOjzoUnkqByDniz6N4EdRiKPzt4sdSus23wgO2b7ty9tZhVb2HrlymUik9Vvqg+8f
VvaVMnoTa3a+Hq5bL981fWR2CjmfuHut4eHk0wHCQt1/um6mOGlRtGPq8UNf+h4PExHNZBMaNnYv
9e+CtsiaXFCa7qzcnpna2Z2Qf+2ms7mlfOHg9m3GqJ43Nfu9p1MLFeIQqK9/YmnHSufFiIba3API
I/rIQ0vsTxvF1qshvMYRgw2Z2/IhFpo20x5Mo8rdSxyMARXdwRCF9qAB1ok28IRw1kpYQIAdoVga
UZM9ue3J0w4pcPYTBU83kRdQtdvWhr4ww3S8q5SGMLwOY9e2sAH5rcKqc6K7Eaz408AZuq63Aco+
R1QYE5BKovpDuGvWh9cB3vkH5BxqUV122a5RzHGCTbykEeeth9YusX70ulNuk57udfBR6rQj2L1Y
BZKEX6tctHkVJUNKavlyt7uBqlz8VY+OTfJvaBmvoPCfjRbDzyvQdINcIK+sc0q3smDTFoyGaYIM
cCNSkv1WStG11wSAyxHrb7tJC6fiy9CSWHpItMTulpVj2yaLMCbOOnuBEaoYw2KTbsGuNKxhrZpC
oiOpwux3KzGIBueGM6i/lty1CFapqjvU3NIdLiI0u8IrGVJ3EYjn/Fso0LyXG06LYPHcG+BmaZhS
UMoCqW21j/gJ4c1zn4bX1UXAeAkdA+dcioMM9xD8tHRpeYxfVCtWVH1sOoOnxJUDhae7azRb225Q
w2qqgGB/5zE/Dv99K9HkquV8wN+CtM9pxuIA2hNE3CfA3S0XhapKiU0/8O4Fitg9DZhLLMysH9h0
uc0YjYMl7JTkTa+97MlxykAT8ZjTcONUUf97XpOVMnu6iVJMI1Z9s75rNV0qxE6z5DJgHDIVdaB+
wJToRviO+L+L08zLno+A1sbnuqPIXBtDDwb7BHFep0y8XL+ICtblVIPtu6NIjqgKTwvBJdY1T/7G
njrA/hLdVzq3hvHZkaBVOuQ3oNGj0XPKE2aZQa9NHrNKStOxFK9T+RoC4WCc2avPFfCPMb/RRu0C
a/bmUF5Q9h1SN9NjwKtj2Qi6Oh6uawlmAafK15YD4Ffv7apyzPvo934wVwb+FY9VMTGq2RtWfcmE
rs8zmwT2w+I4/+c6RCV7H0u5+d4lIhiKhUfgLnDo2/c6M/djKDCTI72F7PeFzRZx3pt21lk9TlXm
T+7AUf8dxgblXs6ypBjsHTxYnkhcOdF7CUIh0nDdduF68/jrm6SkyIFTlxaYniplo/wP1byHt8UK
9RZtexLQb6fRd/SjqAx8vdrNid4ra7nxoqq+dWEkkNcAT1X6enqAVgCnLpZ4EwYYHM451ruqn+px
8hs1bC1z3wyloZAzgdO4KpprHAJUm+1EJGnhU3vYdsY6mD806EXeQHeAlaFqL2DPnbzKQrYvUl4Q
OCf4Ub8OEDHnf/tT64tZ4tbnTYF6onvEFEre0GrIXjzHqPVWYjPNW30NKkiUl/p1DXC8u4wXk2x/
kusn0Y8umLIxuH8/uVDCWByTMbI7hnpOxXviYOi/C3Vh+8yUuU2IY1IPItPNUFou1DoW2hiCoqFm
D4PccrTv9r6fcAiFHUkEsJBpI6DsWFS0/veVMT8pU6fKWdVy4moK0vXHFpa0xR9jJaHAUJJHE/p8
thTV85Ixsc4BFLdT7KlrV2SUVfyy6d1+aaBRVdgG4vcNfKuCTpCQAYq3dS2jXKJ/uci+XZPXqp7j
v79n/HRRWgjO9uzTfP4PArwtcaW2FlWibIFokETWQZbicSZaedZtvW7TNz2h3DCdt1R2E2kmstNH
BlC7+ITQuS/HQECUXgAVEpXuW/Ho1QIug/1wDfGjLJ1/8QEFfSHrfyDnFRJX6qSw01iL0yaxKRqA
dxCyDneVgls7hQT78Q0z+KM5Mf3SHSvxS8IbrXoNBPcbHUho3CnaWhcLkQL1r6ldp6QvZHZG58x4
nqKFHD2ijgKEUJDdf2VmYdB7aGf6RJ1k5AwnH8LenoANEeiiYVYwm7oPY49tRsJfLrzDKH44+2bZ
chMip0nJEgEU1pBg2gaQ5RpiQbGf6VKSN44vRtT9KRTyvJ1FlWGLfkx4ZksfeifdBOsakg12oicM
CjOLjWCoxCNqvnOfJrSjtqQRtuXKJJArNUnF0BXvcNAfMoGyvMx+3CIw6AA0+pZhIZyUhP22TgBE
Xl0MKGFM/Q47AwfcCGzQJZQ0sWP1bj36IPFAxbOANHxPJcKA30EJ7z5zxuyOYB1CWHSC68+PI6+X
xfzrhRU8aJqSBH8xdMuylGyDvSqOB6WNV+e/6LPAMZmV4OT62/UDmlRDRv7VBnhN7sYXNwU/iSEU
MdnAzbBaNMmq6g10NR3xOAz7xgGNUMzsYNJCuxWa9yyXZxT4QlUBDLb//zjTb4vHVy0krECKomHm
tQXTpt0hr/qqukE/tJkOlZ5mjTbVxaPGyX8kld1jI6PHAiwkyNKmgqUL1uYOWiyazykAwULUdn8j
VA5gAjEqoL6n80Z9vcwIPMHk5bBIzbfQViXVh7YM22pNhPnYWIpgaY0IaUtlcza+uKv3WH+579Ap
+xq7OuCvwJBRTV7Qx5MR8LIjADvNHiueLcH2CwUf+cGl69SHWiEtiQvfuIQTR5e6ZQPJzcs2jwN8
rMt3S4A7X3bN4Q8hRd16E7kRRTUF7azdBw7wW6COevmBGQcwpl6nEz0BpgHHLilqvBLv+a5RY5Ql
ebSVzsN2zVWxDynZPaxI2xnNcG4YY4nLLDnQY9b92FOzWjDJmke3cZSyVeexjxvsGdtKbgweTgMo
DdjXu9OdGH1vXtAz5GZ2CrpmeKZfICmHPBs2oqxawsXRwLtel5kLkU9zhh6whiSfSEZD9Pjp1WU5
EFjHAwzmFlaMyEe2Y9SLIOcbQB/w9sSqCybNxs9bABLMQ4TLLy/FGmr1qzKFMnVYWs2cYABnk24V
O88MctDGniis6r5WUkvlyb0Gys8TasIQbMf/DzliYHWhX0sCh4n8FAQGatPMoTE2zGHY8n8AveUZ
XvQ42+0IUPIKIZ99GJS3X/zBdNK0CkdgFPUIPOjCS6V4OriWorplIGU/6e2fEWhhM1ivk9hKTfay
DtjFOg+xQgYz2U8yVsrSBHbMq9W0SmCSll2GsI2rCF8CkRfg9rGUGBMqe9gTH9RSeWmY+1Vg87DA
j0Fx0nv+XM/Nh8BLusDsOmvPJHCzsN5hehmeylUVcy83xlIZHk8LLDAassubcVFi8V3uYYnK2AGG
Gzg0gNcAh3mPpzAu42dXYp1O27/kohgx1KklGA7Dvh6QjoU27js66I1b6/zTc03hCOyS2X74vnEr
wX4Af9SASPocKQAaipeWYu3I+PvmZiGATrRHsU1b9kNIfGMMRoRmNrggzIuGfRUWpNrEU7mt4c36
o0pjebdPvgt77sdzeseCmU8MX/XgEN/S9Z+zDX01/BBq60aqph1BnjWQKxuYMbLg7lguWDiiH29G
fkoPW9G73Wi68aCczuRUMHQMOT3XpKKTTUYVk7RozcpxV+FlFskLURibB8lC5LzKAGih04GNgd6V
mLDlZvSz5Sja/VlrnABqd38KS6QopsmrHB1Dk/2ZCKnYzUkQTkglwlYy1h/ht88ZNKvN3CaDKo0s
IZMQBsbQSQYxaYK5y3v9jbWYIki76nIfSIVtb4E3s7KD1kedIEzT83ppjUG4lTwU5tokwQCAlB+Y
sdWzUQwviCl2ie5DhAOsKAVnllxOdzJGbFG+X6qG0Zq+KchLuE6A27qj+X+vG907lAV1w6JyEp8u
1FR/f9c8S6VB1Rhx6D7cWkDubTXN89KKB9CnYu8+nz+FzCGnvjVMitj1vc7fRXCuz/BKTu6INqn4
AiX3apa+9E5vTX+RPdAfqwvL4cxBGvupM2g/Y0+RyPBFkDgKMCszRPwpT7igFKU1zI5bmYxaJFx/
QBneAzbPn51ifkHsPsSw4aQVvbQ8B19+qLc07aK3CR5nubIl2GRtw8RIdxAWwiFWqHnmtjnHmhNY
+SEFLMV5LmzebiJEYyKw8o3qSTFtQnhYrrLH8ITPGcRM3N/3InT852H9oIQyOhE1qIti8xtslsZD
EK+7khnKY0lNdH0IX/2mQVbfj3aHYM/7K/zPA/eohi3aBNwIqt0vnB7EkNwCyIooTDH6eWbmeRCc
CxDwTRlq0Q0SClXTwXylV+ZjNE2yxHSl2mjc04p/b4B+4PVpxRR2LO6xKu9+UPVW1cWETHsDm90K
bOjoTUA1NYHjokQ1jJpYxeyF+xxChzE35Wx+WwqJ7/G316aTZLyse+DN9ZhIDK2L2l6C43Ni+1YK
mcAaase+MGr0xp+NDBg6lVmGxAsDko4x+9LeJ4DTwrA9DsEXJJHWDjJt44pStuDfDBT0swZE/Zvm
KdJ8fbr1yuu9eAWL8TPfIcmtap2v8mQWOMVLDY3WskUqS4jpK2NuF0W/PYCbABRoXUCQs6DmQitS
BhBnui//0iHDodAhRGmmqPo1K7kUa94v4JBcpQnxf9clOyuUdvgJa1+k9sw+MXNlkxmS140U+ymf
OB9DPTX6FyA1B+Sfb50V6VixCNPi0z+TJajauaDPp9MAAE0UCT0AjNWXyWSn+56QHpTw0NKyFdQ4
GjIoXre7sXpSexgND4c4xeiqTPyLWWMvLNwsFFqc+H8uCkS8K2dEaFOj5cDqNUdUfl5Q2uiO/V8+
fn89IV3NSiyvaF82X6QqP0vQAFaRYCxpc149wfs9GPIrBp1t8yVyraY0nq57bPJfnEL5xDyrv9oK
AkGN8uafAjbAdZVSffOlnROALXXRjpPKdI5TA/BBlSKkyAgbxKrK22XAX94sxb0F3/y0yWZJ87ix
+5Ue0E7YhoFoJyM6iLLD+e7dUm44N+ssaPWtSx77/G/I0weDdDAdVEu63tCbSKYja8vxMP/RDIV7
hTFQTA4zKrQaJhT0pQDXT/chAJQdmOVxH/syihIoZG8cLEoFxZOmWXYkOMgiQVFyUdubexajO3cw
VoQu/TpoPS8bZIbM/R56i19nk24Ha2wggkmbeYDNpf0mJoY4kMI+XWXnhfQVg7d5n7gDP+mB+zK+
W/0e+xSOClDI+T6G15637xQUFm8AFsl0ITD7MQYuwMynfeZQXwtFmDsFrTQs1IUjJ/+AezFV/dMj
Ulx2St6LQTFehfuznTHG9MlprGxhJae4pt51gtgERAMtjZliVFvXVX8QUNLg5ijMls0yYfbhaKpn
w1a8sy6OTMlv0wjl/FTPEIk9AEo7APipqWOKT9h5+nWTfY/AODwdqXhfzLhykKCacBoZoUvoF7ay
CpeojhpK9PFRVqGNTg8QnRUOoWkUGlrxPqvjyq75xBPwzfUQkqsBEt0r/kmNkawqzly0LkMaQUxo
BYEaK27/uelXrmxhSbcPFZqxyyFYYY5czoWNh6Qy/bTjk2la/H5UuMp2NxU/45RhO8bKeOHAqdkh
O8GNk0DYQMAEo6hE6mSCBjpcvx7KpQqMBKoIEFRVbGjrZ+SDuJK676McloxtcRaqv+HeYNRI/fZT
UTZMLjDUPT/P3tn5cGrvV7QAoP5bLvO0wAbmTjyfTQG2oInnZ7GhdSbbEIRQoJv6Htekoi7tzXsu
OHZajIHs1wa0CABYZZdOMWKbMydh9/S1WaTVssQUfdXViZd1qfwKNq4PoX4EEuaUN6y0x/9VqSOA
MuX0r1DBQP3PXGieLab5Ueyfp/VISWpqiyCki1ZdTvfvKITPW5nwfp/nw2+FOH62FtxuDPjw7bDz
rmcd9U7VGprh5ft+hR3YrWrG87VsyGf8l6BTUgq0WjBK3p2IHhIxKQYolY09ambWSnXZZE2BWLpv
xMi88CvnTPJKhGVm94Mv6EfLIkSBxWY9gCFyNxxhH+R1t2jkguqxm/OIDepn6j1NZBHFHdmWsS4I
wfWCNvKCD7RTy1i9R99d/wrAn0Q5NXbKE1HQtAfTK04R2ErWu75tMBu2nY9ENqfp4i3oyjCNJtRm
DGcuG1SiNrqMXrPq0k35eDemP9Jxcjy5UwcyRkXS54vm1P9fYTIgTdA3JwoNLZJo4qKhKiViCAKn
yMwMf4YcUk3wBhSCBNdQUBniYIz0nC3aFiUqGIwUZ1Lwkgyy3QAKXWWAcoChjRFKhNyGPujnv/WN
QZXXyCTYpufTkHGZ9+DGioQ+lK7hf+tPmSIn9TK2kfzenS/0Hu+bQ3b6bhYiyngvxpmsGmGhJvm7
miDiB9TCgtgj5FA4nF2cl4fQZSxxrkm3YQObWJOywPIQMZz+hBIlkKoT33Bhe921pBQDykW8O8sj
6LpUDaYUDIaOAwAa/n7pKy4pmZ6hNEG1Bh98EAuQawbyjQ/sxesw6rcz6YroLyqDnHsFA13G5bZj
uyJb9XB9wAj8jaT8nncjp9Zva24TTj65eUsMLzjvd8FX6IXpj2FosLj1CewixISQlpxjzazU8Y0z
5jtgT9A9BKaHL+4qBvn3hnbQjZrN8UmdkdP9QsshLGa7b/gYjz6z8b5zXSZI+J0juz+Rz5KH7fPE
723HHZMPjoa+UTNqw0qfU8KpAOAYEtTfO63/mMmjZrqz344jkTMt73wLJW3OBiPs8Sd37Ozvo1vB
qQVZT3wc25UaFwLjj4J8WBtqCJVxKgco0kGErmBMzN7dy2SsdWFdhvmCpXuvPSCNeERW2hIy+Z0H
JS+qviJn+uAT/B48nJdfMhlaxA2dT98rPB9BUnm5uvN0dVvFBviqOYng8FTYUMuy/sioLr34vQcm
PPFEK5rnWLSA/HqX6DnYxOxe2Yg917WMMcaJSzlsR7AgapFek95TXuQ8AWGbNU8/iu8XyV7SeDqz
Z3Zh2wxBCKuCtP/4f6/7Az816Eoa6gU33GuHkISKhPlt8RehweTyT4aTvOFbpjZCsin3CK6QUZrz
tCXeIEV/p5Gpx7QwlKZy1EspYnNCKWoRtD/01KMuGOpADSVNvR2iQbiUW5SvDk3fxxJOS5NNom4u
ZjdvBUP2sXo5RkadEBl6orYx9kFKtMoWE+0nxvm5Fcm1Jwdk6EqgdmY8fhKbnbZFXUX9ChY2mFWu
Wkp54JzAyvSU7Z1BnVvHpHQ48msvq61kqkccGUDU0BuS3QtylvWf/HJuc/RU/htnDmCj/7aeVE/0
WBmaF6grFtb9WTBTHG/1pWOQC9clk7AEENjuUG9rsMnUs0ERpnFK5FqXB0nuue79MBf8bo3MXyUf
ozPJDIEKLy1g/mxYqKoqY84Wquuc0AP3GaATmNShDiy668RjUgRICfOoDGjMcHcL3oQw6l6M9jF1
/xaEsSkMjoPtevElTFAr/KPT4mjsi95g1LbJ+mSKzWNlPqbyae7gKy9nmvizWqFYFhEisFbbLdh8
NBft3Y1OBrMf96tf8AfQFaCtdT0rBcWSch8fvjdj12ORWGF7jCJzOGzOmhksbneNWrcnrGUQJTl1
NNU+AbHsDOMEu9GK3AJ4IRBG6ZpwYK2+rnk9XfVyFXWkol30GF0xxWRB8p9GwO97iT4qeyO3lAcm
ByhEgsoDCbmEu/1O1ESkZyrdTUhNQl/AVPmto4azJJ1zg8fLi8HSstugiM83zUsslUXdiUNxsyXW
uiwb2KH7G5QEzhptAcJwz1TTvCGfBHMkq9GBoRmrhXhf6nYq9uIkrQFQ0Rc3ZmmAfkdTkQf7pxH4
FznqCfYwQhpTq9fE0ZDpls2q7oTR2VOLZS3SuHvC8cwGKzHcv3AwtFpqtzckWuQxdLcZM6Cvbgs5
Cft0g5hhIvMx85S+XGIFE5EnUODN7Fl7C9XZnYCTq5DPEoVyUwGdvWggryJa39ANuWtm7VFTBZnc
c6QhhvEdHprSyH873QTaduXz5paD6MDD/skw01LSna5Bt0V85dTNzo7FT8AbO1kdSJRu51MPo+pU
W2U1cCl0ifqCPRcqRR0S0s+QhZDQS6zcrlerKWMTtZBFagmJUNJypbFyGTNaIHzhq2nifsASEclN
3VKuJ/RPgQOUbDqkidy/BLi69p/Q2I8kabX3f0WU4PXFPijKV39ryapUCaqOxaJcPD5EXD4oQ6EC
RCD0EgjlaQANiL3hHY3U+aIEk0fDr4mFC4Rnk02/6zuYfmZnDLVr0zBijGnjRStTRS+nF4Fj82TD
baggtbQ1CoowoQKRfOVgzoa/jBa4YCLxpK/2cuccMksZ9k1+U/L0nRNMBEJSZwTETS93aLgW3oVA
yCZbFs0ZWXL0rP2RkKO+bvxl6dCdC1pUKv82wvjtGjX64wh3dcZHJewx4HaK0tEfyB04OgGjVNFI
j2ugdMm8+3l3p5ZaRAzHaPDThhyliwBUxV0RiiLAQXdOy9oHFP7S9iJ8O7Wx/weP2oc46kYIus9g
MkE3m2/2a4h/dJKzd6rdB+3MLhv7zoN5scdw97h7p1cnqQUiqXhB6oShQWpwBtTlMsB3yZQ28N9g
I+KNA6OCSUqWzKUDPjsIDLiadMN9glBKS8wybY0y/e9qDL9PLuDFzOxDIj7whISH9nIjKYV/5xW0
Az29gjJzDAQh5oMn9C7PUFxNZknT1Tra4XLmoXPhMpqIRNtVHfSVwa2K47+iXX8WEyTmmDfkrYj5
xuOOXddEi+rtCvl7LQBBHmerR5SW/wASS8T6eRmjWUTE/S91YOie37FZN3qIaSoeGyDuhgHlQHVT
TqQNr/uDTIFQ2gpbqH8UZknkKfvdRUZDeLL7QHWy8UvOiR9RqAjDNIXx0oo1kf67m+GL4Yqe1Xhb
gOKDTQ/BGpmzUN4/fzCNc4G8hiiOFPwLfVb9t+0docRVRFo5Hhpmy5mdmIX8gDRUhG8Md0Nziznh
ealRlsUdPTL6Z5Dy6Fx6SB/Y24j5MNhx3ocIwbs+GtCdBFYQbGfwEOpA/1Q8dd+a1Ju9H80gmkuc
i2+K6kSFK3YPOTpFJhflvpKW8F8WEpLqPr4kyDEvF6Pd1guF4R3xKNZ8EnOrz5se+IqFiO/j76sh
kSJ/qPXzoahEVGDrI14Vz6kAPs5RrUdTAkBZQ69e5L8KC8Ul2SvMJsGARKrurSccuLTtfzn2dr4e
eepaXJQ53tKQzZprdU+iFcmoH5uRaePoO5XN9jzGFU/f+HKADYyoeIfKHuBggQjTb/eoFI/PC1+B
68LYl7qDPbRpJPZ2ziM8mm+puHi5XzaeLe3WxuakBOmaeD5orbqPpXRVyT8TsIR95SYWEqM+OsqT
mHVsl6+Om+Yva/RCHbtqIy7Z3Ia1qhPx40fD5O8NC2t8ubHZnlalAhJf7TjEA8MQATpaRDHBJt7w
EywAbT/vYEPhLuDE8CKPqh+s26pIPxTAIf+FQt/ag5GNOvfXyLyeQBHdsEXfm+G74vTm9fzMvtTU
HA1BtSQo3wD0jNpEFTxP98G6IGTK9Sz1Ih8GP01Fr2AwaCv8po1cxBjeNrODdcQdWypkLwK5Vs/x
j53+4xjfrWGOOXfL51nkYZQk/8j6xXO9nTHiQzx9GTNABf/sKDCpK6w+mu/8Av6BfR6hgn/1uE+f
HlWAgT/wzYYbEZwawJkf4WfB4dxUxvRimjz9N7Q8/xTeg1DlzCA24ETqm+ezguPXXLLZ10MVYiwi
1EBhkqbZBB/9kMu5II2fIysn7Y3IPXW2Xj480E0GNKDfyZpQlxLLwcbDN9YPglWt0A/XI3WLO3Xm
29q8hJxIVtZTXZIoRczLbbP5NFzvnkxtYq28hwtXuy+qgoozduQlEMuTFV3Y8b5FVvTl8OsVogfV
H2/t0VjCeIQ6KGpRHAq32bKBUiR/GpqFBjC/5QKTI4JkV8a47LBKWUYi9qA+BBL8cFz2zbJ/QM/G
vgOiYxP3E2Cmk6ON0+hPbnh/XIikTSE1UJepuHfSXuUy2VD3mtITvw2E+mImCvq0Ulvhv1fna5sk
xxSY2heZZr6VCjBFsDmE2qmYpeOgIS53geHwepbxPEP3cs5R/2UL4h1hV/HRXkfy3ooLcLANBqCu
8yDzYmPtzLYLriTA0dvnxm6TUpaBrxCWcK9PU21I1D5+Nu7Swi/xxKe0qDhlEmZWvWTsH6tAstz+
UAu2tWscRWPZvjwPOVwFCst0hW4oCyS/KwKqN1sOL0mJvz+w/uK7CmDLrCNVlTSR91IgufoEIzEO
K6jNKDNJSZQnQ0vV9fDITrisJKmzXy9gJNLoqApKpHD/yUu2X0o9F6iuQrhBabfZNEtrZecd2fBN
8DwLcXFXAXCeACdiq1GfEh/Xss5ywaeqaBf6xXVkx2GKQ9XHl4oBj9dE0ud2DtUmuRqyKAZf51mH
gOwVnpOc8o5BojINzIHIhlbbKqgPu5nEkB/bwyqRGuUSSPAc6fXgtg7K0PIzn6XBglXZlv6MS7vU
CN838lz1DZNyD+xCw+cGCkDaKrODGiiUQVtPz5E3te+GBCR6cbWCjwE0mv8q9Elo8S2vru+vcKE5
sawTjmX/jMt8Q/ABpQ2ZqtZKQ9a0Gd95yHsHWu57X3WiRj/YpKDO6LAtG95CMpITUzR1pGVrmLk0
1sr47KrH6gM4HANp9lIjwNe7hI2JxJoCBm67pT3ZeOHe2GGqZxcqB8NM8/nbXOab6a107xvtmcuk
Ds9irvSaeq6XA6m2wOB90Gzj8FtG1VZy8wDXmddXdBLA9fCyrOcjQtbZHicdK+Ga9niT5ZQC1Ltd
U+i4N6EFGJlSiyyOmcTCBNAylSk9v8l3mAtMMWsxxItd94Z7K+u6b3m4sfXgKqgH5aAyNDcPOfUp
Cg96Cj/GB59YoOAJAuFhxKEmUuyrzJb+0ksv7ycnHrM6EIikflilhx8taYc+i5/L7Of+WU1vwq0L
ITGyBT8+5QAFs7tSzDoErvYhlewaldHMMHwIHvrDmZ/0WUSKldXlpI9vI2RlxfVPzhQwSPXB4Ksf
CiNNv6BYF7RkuMvDqSz0/BW2vRwzHXA36FaznGKfFay6eJvF1CSwBLfWJYI+T4DrOwcCS+2TC7b4
Hdno4fWazqOTEnHLY1rHPiLr/XO7drEeAK8XQQjF5KXm8wuOlcEi7q0mB0GBvztNKF8nNq0CWYnI
6XaoLK0i3DqVZI9rzLwLQ6mGpaJQvLcrZS+kY/7ttkVKelno4GFio7SVIXYdbzmZXQeus1HAflXq
mNCTKVUZrGnxeG8YZS5qZYqhYh24yDpxBiHoQe219zXXLRdu1VrfqFTVyjMHBGIub8UjrnJ+3Cco
rPAZHAJLefYF6kgebspS0L1YjVXQL5y07VGvI9Qjvj8I/56ZI99NyqNk6eiJoa1I/dS5VlH/ACcg
BXBi4CloTqy8HCPRdmHWd8FtPA7ZKmfD1a9a6btFhsuCzOL0Nyp2eQXA3hjOtKWuOQ4gSMQNKR7x
SiTb1g8xIdQPA8r8SPiNPyEz4ErIEsLo8I3cHJlP0FAz1oPiMoTkljWXam7aeoRXuIadW6QCmYJP
vY2jy8gBTfWnyEYHrxTaGQ3NFMeGofPMDnjFw3lylWoXHzli57eh6s98QDO+PVaNhsX6VO7qwOSd
m+fkCWFQ+pydYmdE7K5mtiOZb446wbyoljaVGHTYTjROocRSOkGHOcKApSlSHy6+5VfkoVQPi1aU
Jvfqk1KlDp+Q+N4aFoy/jtZbyzYKrLmKvsVa+PBo7RyF7YIv5t4BBuC7BOCHmeM0hROwRDPtU3Mp
BKNuEIvyvNgcXiRts1KlWWW69JuhUqfjCbQhIim0z7chxqXToCiaKC/pl6SdjGmefJN/A9K3g6l8
6eGNuQESEniUy9Nv2o0QiO1GQkbgGf9TXz23m4MW6Uiyy8wlXkDpVR6kXW38NyRMKFgP66CZqZBV
Hjo4opf+VCNt7bp93fksgUPhvugxMaw0DFS/KYcckAA9kBIvOZO03yXPee6kiDOgCqJItqHzXZx+
J+sObrLHDrxrBkVhDFvAOpc013FDh/ofZSpIPrjLOaahtSn60PFV4S2cOQiG9UL3IJ2Svixb6p8/
IjcmJJ4xKEdI88zHp9n4bFRVPh/BRkuzTU1rla51twC3sUNFFP3efx9dhfl+QBrqha+0dWMvwn5B
qKf6Owo+p1tqHDkFHIEMp1ViiqGE/RIOehSNrXqndvBYWz6chYirwWzukEe8WklUyrpzNQ1yz38r
s464Y1uhr/UzTp+txYCltOzxOQ/ncuDOFV9eA9/AGpgTHvQYlQDAYYIhj/xG98K7xC9sPuv50l9V
TeCOiCglK01IMOmx5yhm03EQKEWkD+NICvdmvfP5HHeKtxsv0PY9iHIhc47OOU3EYYtqEysQUQN+
F5NqJqlFhkj/ZsmTFP6RxuH1cYpTj39pg+qQZaqcm2OdxQFWqROVf/fc960NmaZJEKn9BBHwBL0T
g8pJd5Ck6tXJmdbH080DKf3FpRcOjuvjWIMcIjcGYuyq9eDhdCwfCtP2f5I74ItgIU9rVdd7kr5x
QQkeMm/FN6hKJt4RhcwW/q5mYRKBtzRXTB4PFVGTiAYViJBfhou/ujdSyU3B9YNl3Xe5F3T4xNMc
gcDx1YtTTbXUEQP2peBtiLpc+t4zqh+wc7JaZdneYOGpCkI9BXncaWas6mOlKYV8KhlHUFJhH+S4
Cr8CXRhVAvr+Mu4vohXbsUaseExe1NuGyrj826kvluedZ+Bio3TwNtX+NLGgFv3XZnLroeeczIBH
N7L1qEXFD/g0/k1A4leqoZseXmhA4g0p2HZtE2N604lwS+PhkeZR5qCMqDOSl9tL1lVeP0GPAtLb
lzZu+Mn0GSvm4WJHMPCElWzdRXmR17u6Hvol9GFNa8w2dJJYrKxo8lNa0q5vHXrfuvALVNEitEzr
SUU4yrx4BxZlodhvp+UnDBje9Gr7Cfyeuwu04AH/z3XCPtRU1Cj1kE943t9UH805JoLJcqlUJeDC
7b4tHUKIfLwejUFZeSpKwWtuZZBGB9Y/f/MdfHsJSq039KDeKAkEEaYrx2s/SZZn6qHh1tMEXJbm
XSjkKqh5iXoh89X8qoNe2jisqcDLPmL8OWQhO3IVFbUwgmQvo0A7yIHjOmnsWqLVfpYHTOosiOAk
FZaR37BX5ORKSQvLi7QeXU6yOOx66TgKtMZ95VNyRv81/sxCDiZHH4p17mrTI1062PC8iLUJInHJ
ajECqtWI2mUfLBxAfWSN8b0Pww9O0vJyMrClytssZPtGktwFENqWDC8iDkNLGu8sQav64PB1JY/F
mj6Xt561FBR2Q0pGR6DcGZxQXgKsICM2zDdEj9KnvXjaGZFKcpIZ/VR5vNdCTShJzAlr1c1HKbdi
2T+6lcnpinylNGpx9v/S2MLpSYAfhUheAOCUSyjN3pCkvnNbKcf/x9dg5JKD0+drDmGgtTyK9pw5
JIxrKeniKlwJ4RifwL73Ei38NdsxY/Qs6d/cgtCB4puMKZDILt3TY9eKoGTRaks13iyHTD1NznQo
U+rzmbiwlknfbnV6aInWa/h99w8T5NgKGPJfTTJInhviOmI6IQ43/pZLFCtPPHZ1co8FL1Rxmukq
PSV3Pe+ugfn+zLj2lL3AXrsXsMIhR6OS+l621SQwmaGMkkqdkZlTjSM4hqKtmVW9H4y5iLim971J
IgaGaJ33dmm1E50hslpYM2ERb+WxCqvrOo6K/w1sa9KPnaz20lsw32xvknP60Tg2TZNjlk0+dTdH
aWbWSo/i7TloKd3cX27lOkWAfrmxoGGjMm6UENEvxiUR3arMJk/cuRmbxBNcSCedJHtEceXw+oDt
Iy6f9pEEcVd46By7ZtdHByfurLPgurb5uHwMf0aGvSry4/7kRzG6WzF4q9gUNrri+2YWAj4MwxDF
UrvdoXnP5L9Ed6HZOcE35g+XABfAmZgYlBGgXhg26/Ehvj5FBBlPOowToKxUjBG8BvIuH1FdNLPz
3GRqQCF6UkhS+zM+WoelJ1uy8n8YNUP4q59SswXpRm4TeI0b+yA5jKAWONx2ZqOv10XteSqyVIxf
tmmfqC3V3l2qqgN79WcFbBgLO9y1GLU30B1TK7aIlQrQ0xpTI2fGdr2snU5XDg7chPLFh2VbaTbG
0PC/nWd7tJVLTHLAJQ56aDlnqLEWEq5akNUkst/nVwmRb6wtTkLi3OR3EMKrG3w8F1QPiT2ozrRc
e1AlB27iEr/Y9Fj+lOFB4Jz67NFyt196zfrQToYrpK0aRYahFuWSt5loLBgyrXbcssOLlAGB4fOq
rBfUqgGglPHudexMWPj8WfXqcQQKNwLQukGUp6M1Q8sY8BHvo0vkuGQmkOL6n3X8AWS7lMKEO9ce
PTbhEGwA7na5yT8O6NsOReA2k5+teEluhY9CPalckPKX4THscNeB8Bqkre/r42CK0z6bdwaZLjDB
3dZbr6GFK6JLIYZoBsJDbzm45RVBH405JOVL0HgcQgSpHtK8Btd1xt2yxH5K0hioralffn9AdKiV
r6LeXibxXVzBstKfEunaQJfJUyw44cX9KekOmMaY3toqnJ7J2c1KGCOJhVJBZFIjk8rmNuw5qgzv
uipiGMhWnN6IeTmNYYXwOIphkyarlMB4BELZkueYSpT2cvkYPWINf25dL7MxV5tdPZuk9ZEgQ19J
g8sXERMKAjllfTlgTWs21AvNZffthgCHco+FY4onT9ZycX19tKAyJ3VZ6fxNnWrEc4pMHqT2Ct+j
PKe/RtY5w29I5J527WOwY7oLlJohU3Ar3YJxoETYUxtznNy70Nu/+ghjkkoYdR+n0/c4od4IokxN
t0D1Ozummq7Hf2++eVVus4fbcRdfZJmdUtGEXQgwUAaAUYWn4qcw1zpRKt7jPXMsJL8ttSc2uXz2
brnBMgdUd550Z8Iez7LY9OS1T7W6OvYmlMbjpvEsLoWciBXUeXxNOkNgrgTqXUm0VJccZF7AptLC
AT4r1GaCyPWb7PhlscCRhuflY2aj64wK6sqk2rD/SxlRAJCggAY1Gfmy861bcrXwFOKUBIX1BCYV
6gC3BqXzvdjBCVJ0sNn5o5bX0DObWQs9iDtBOYXwfXXgvzgyyFeWXX0rZ5ZOKCYyccVDLdxqqD/n
BopzTNQlUxk9e1rHeM5P7l8VqZ4sMzjxg1SG+/J8Z0iMDfHiy6Kc5pOmeQEMuOIuxfqFPtJo/J4N
eCctzvg9GgwMYM8g/s8PbY5FjdUuY+PnqgH9Qg/PLBltSy2ldBNMfThC7J1NWuogxLzHA2j870wp
Qdk8ha2lLGU/4jVIRikyjZr/I+m6adeiaqX7nE+B5R7yDHgyTdIhR5MALBMIJqt4J5ueqZ5G3I/6
G+YMZ0It8BZav4RbOypxXSHs00/z4JI15HPUyACbnfnsbJrDgwqyXyxb2tIC3oD0pteSsrH7AzUm
GKlpR+LEbIaZmaeOJ+s05Ef66AKBTmTJQTT+ZQjbgJ38t0PSUqAt+boJhtVsPHiy/vvUvg5zd0Nh
FTeSiLd6+VHroHR1cpi8Qm+lm3RMp1404zHKobK0aL3e0KiXqnxRjtGrCxPmy92Jpb1CMx+uD3JX
hOb8arSj8zLeg9Nmomr8K03KINM9V6Y/hst1BlZEbNO/FQuefvb5QGzi+GPK/XWnU5isu6MhP+lx
5PIYUl8xzTTzdardSewTYJqIb3gIn2P9QoI+lp20WsvT58Tzgwn9UJ1SuOM8q0ng8ldf7JUiVPg3
PspB4K9uz6CI8bLhxNiXCQKyJX7tShEvhcQbPtq2VcQarMYp2VNtytVA8XM1BtbSAhHOLKxPKaH0
ZxlHnZU4n/VFa71xb6UHc2E0MSvx4B7+qdRvLJcpenFloLZ9fUZBaBK3CYcGRoqb9aFJdBKweogC
evMgdjFxyQ6yu5MRykCMVbDSj6mQ/WGL8uV9NfTTGqZPO95So5FJcByStuAk37rDl2eksUS/+Tab
aR7Zot9GnlBM4iEKkfhChcpPeI0NEa8hKTD5LXdXI4wJi/IhIIjUPo7ka29tpTBEL9lHMs0hR8Nx
c5J8Sba5loeFei0nnVCS5JsHCwtJWGJSTfajCWUNriZZQnghYfpduDoWARPSKDqR76odFpOHSKKF
W83IfYIf8Ltd9TarCEZqVS1ykfSv5/vwkXEksfImTMJcsDdfaNpJAjWArJ6FikwlqK8kPQNB4y3d
7WNI4SbgrGleoEDWY1lWlhcX7QZIBfVRQlS4GxbqtYD74siotG+Uo02wE1IVg9haCvW0anBwCh8a
xyksYaONHtZIyIT9Zc7ppKL7ETCx0+5vc51HIfpG0pATg0XY2taiG3h1NJmHg99i+ZzVbx+pn11O
s1vDl/9DWbZ4l4gKGGigObu/zCZfUGx3yi4qKxFHo8rpmSa4x0own4dWKhm8bF00V9eznQ0B6Kwt
tMbz72IgGBR4+qFVzxjykowFeqW+99QTqX9s9hXr7OAlZEl2nuyH+sX7NmIOtPUn3nRrg3SrmX26
8zAOHRzyZL0nWqP3BVTiu8basFUE9OSOFppAOKGP8EGM8SHM37qwXOe8Zbhs28cifPedILw8v3tN
9lT1TAu6I5fY41j6wiMQMFyYYlBvBlfEfzlyVxAR04HSd04qgs2ssAOFBgYa8/awZYLkuhmrmQl7
TX6JmBYJoECGtcFv2++dVVeOI0qYNs/OdGcooARdQ61tUEsiDuwUebjg3wJtlrmeXwWsfMjmWdRA
xu92Op8vWOq+xixcWe98fJNS5X6lfd975pZdAfJu1/FvUDns+EZiVsxPRfE7+afns1C2VE01MpJx
9OJc4ZLRpYQgL9kXqw57GBQdnNp/c1bqWb0JYfHDto29COU1qcKTSYQO+udUShf5dpM8a/u4LedW
IiF67f36K+CcpVVgZERXWrZUPSqeSh/yi8o6sqQ4Vv5Q9B76QZ8Din8nbMsnScx7MVOvDp/rIj/E
mGqBMfK5rnhhaTUICYQ8sgWWnXzYwpnV8v6jG527EGfn6a9sFQlrx8vDYxvTlALoLyo81QJ5eUeq
R7eXbZzN4ojHTfEy8BX/yqhi1vDQMdXegH9aW1l/k/kQuv5Y0KDkk3pr9n/CqxbLs/nGQ/AjQIE/
w2joM+wGKL/Q5VLYfGzQHPVcCD+rZzMnV6h7Mxbl4zvydueHfKEDevZ1btRFTH2vkZhKWKBv68tf
v/l/hNR/uczRjVBp642pmfcY+X7tqra78bWpt8rdy7U4kgHC0PkKw561Shfn9I08IrVs86AFwPxn
MzLqjXXlgB6j10AoDa8D3532LeylX+4wFlB6Uye89uK6/L/gM8853BwrWBpPugbIvCc49NZRirPx
jLHc6FkktufZ4DXZdje4FFPN52zHKhh51SHMcmeHSrcT5BbFaM5tNwbsxwUE2iMcFFS6cO2Q+VXq
Ap6l1efICAFqs6mN7YqDQD2Ko/rhlhvChyGRL2uCI69ic5zoWOhJJc47mldTawS2yFYYwu307gV2
tH0Pbt9QHGdgPvJFFmRSWcGf51N+/xolMgpRPkU9vvfJ5ByMGvpFJV0Fkwx5QfRRGjMHVx/5zi08
AYQlPGKq/aV/kHqRjOx9FwlRwX0PZu6DmYCRira8qtQGn6DUwaLs+WVirf1/Q1EIj2Tk95zFn2U1
+57WHnsTTfXNBsDkz9fFvk/m6LPA6eKKRZ2UTAzGcp9zoI9wQAH79Oo0Drv6r+Rk785cnrzix5yZ
ilaWtZMlzlQpoikgEGHM0JytKEXL0UgoOG4KsDCaPUNXJdVZYkIxCBjN47NYKY1cTQZyDLoqBfcG
8BGl/NSmLxjYGXi6kEd1C/g/ds5tPoTXniDPtEQEsF8MXhNSeonNTV9jPFEFbhihAY52DqvXbC8l
V7rCPiqvP/8DlvxnnPh1x1bGzwMjO2+PJnZfapmYrtaPh0EUQs57RAT63ujRuIQZlLiPtM5rVuWT
98iA/XshHOif4KNvC0UISjJY+PhEtJj1ssf/MJsQKzNCJNuM28goIt066zbGdCWp0Ir7ymoR6PYa
kxTvZRnWMuzH9XDJ2cwv0IZl1IavtweZkEWVwCMC4rHMmCKyvrVXNxMLt0TMUjdInal0WLQ1fc4J
eip73+d2a8R6Cu43bazUeWD3duoaoXdpnn1nV6xxX0a+JBje5gSXUN3bw5ptxXJrW9rKVbzt5Rnw
CslzTC73ezMhrdxHA7KLeSwlbXBFlGiGfkYJ+LAez2neY+FC5yAAIhZdw4b63bUGIENl5cZPiuFn
feypVqlHAacdI7OQ7TfXPKfeEHDLMsuQ3cJPBDA1ZesAdvcm8cP7I/eBQZ/LaT5KWGp1sec0Y5k4
yMlNHMHcdfj9AJxngE4Tah4irX3k98vIGZXb3diLddv2TzzJesm+1OOcHznLUZ8/1xDgLwUUg2u9
xPjyIcEb70l3gXmrDTiijG8QjlXLC3U5jcK/E78Gifwots08DKeRfxyxAiSbxUEdyZd1TdrQYATX
tJod2HA6uajHNOgnEOoAw5Iwyk8c0paJnt57OnxAycjUZy5Byssnids7esJGV3a/J3641Jgn4H77
cZB/M96I/IYB2X9rHQJmWINXk1YjVZihLfUmWooMYbfFK82wZRYY702KvkC/1vRvZdi/LqwTUoC8
I3ljyqLo/lfTQ9CNQdHSAkxSVXFrxYo9UZHrgTHtv4bVxO5YBmS7H++dK2Z5ef9Grt2sxHK/R6CV
nVbGIBWXSRTA/kzITWLF8ghNxwywIyEiFukU9CQurDLKiIs+sby3mGiX4YaFqG5EGHW4bRgmms1g
RsjBT0VrtG3Z2g+009loV1XxQa9TF5nOIFmJTlpMLZL58hBdRxgVfjxuT5azWUXFlWdQ8MP8RPge
FacCAq6KNeH5vAzCIKJO8CR/qD8HoJ+hvF30V1w1VjP+whujpIf0/LIEV1T7/CxtaB3NbVbbk2CK
SU4RUq4pp8gsDSkObkvqun5gAlXfqDyukZxOWxTZC5F6TubupMSEZzw1AieS41HbXmFwPXmtjvr3
MBt3hnHMFavZAFweyEG5mA0aCV6Iv+2mge8i+2MAHLpogzV5b/Vo25KhGPl4K4Bgrw4O9nX/A8nX
CycvpEo6SqN6viL4YE2QzY7JpSIz9RTUt8wpxq2bKvvcNkQOKFt3AE7gxAXuIxx+8BUbFOqQwERe
DFhRg5dAkKfl0hGvEiQiubT/HJixuLMBlG5bxqvpTCqBAlQM+kqmGi5a5w402NIj3raL/Vg0Go0z
7drtUY4mruLyHlcgnzCVJn03T2dztHd63FzV2vBfmIW47D87WZo150J05syqXjfjIAcCQn1Ykv25
KYTvvsnk4aTCXGZcRNl/hMX9QF9H7UNgYk4ykOChlVbd/3rBGBKvC1QpA+B8tLULLYXWmZrLncdW
LgPLVEPYzlNsoi8+E/YteWo/kSC43SNC+tqgACxU/1MuVcNur8WWEO2FBZgQpwxyMXi7NEfI9pDd
rbc2cMzCUzirwkIIo2Mc3gt5TOeHLZ/lsfMhbEX1XmuLp+01qLyU7zYfUle5pqgBEyWWVHBsv1B+
ukFmfUci+CTCdZNzJPWnAzKGzrFyAJFS6MkNj5X+EdxZVaH16m2NB7/tA1rOh1h3JOszAFk/OvAO
Auuzqm0cH8hsFYhDhz09e2kLFuNNa3QF1sEPveLp5g5SSSBfExGpnTZJjhA2ptsPyMtYk49CGYTZ
DNsmk631Tn00frP6Pem33D2tqpNp66hjrU1/pPsAl8Fa98ALvBTWxlhOIsb4zyasnSVV//E+sFRb
qMx2HV/ItZIq/WwXjWASJ1or3sRNaC9ehca4y7POpUTVDTKmClIrlAf1o2IX8uHV/sJxYPEYMcwl
jfhHwcupe2wtm4BzUhZz5a1eZVc2Cy1pf5PYyQ6J5U3X0KJN/jM9bf5LQ5e8Spb6/nSUixJV57KW
EddUG4Fknalb8sb3hP1/G0r70/bWHuAgc0sOwULAuq1DhHRzCQjt4Hir8RvNGDULUIU9asL/kzKF
cyJsBAFOTpItmlqvAh1z82JJAtPOPo3I+lMinteHluGZuIyunTNxrOQqeaAdk5lRVUnS/+D0vKVD
PnBb9IV7d5L3YiIAhafAJjKwffF0Xgxd8SQ+QdZchRuQRrrqocuPHV19ND/1aVWyYhSpxhHzHVAQ
0mBGCra1fY7mb0yH1PEMhozSCyZi0nkHx7fwROpg7tSKZVHoKfu6fzwPuVo7upVswvXIvO6A9Hfa
wyr2rqwLzj0a9uO0z5JZKSRwPjXuMWBZr3ixRWJy0t0l1lguA7x2xzucPtzazdOHYO5JpAz4mZ9m
kP8Ye18qjbnAlhLhclWqRWhLcOEjQvzEo4bSXJqFm1iEUWrB+IQsCVVq/afz0os/D1Nhlgtklf13
iEaLT5N9q5FUkH7f+vXDsyU4Wi33+NUHp6SRvDjMegY4ZC8YboRVddGD6810sERVGtE3UopOX8k0
ECOEKF4X5eAHHak8jk5ZY4dFn+ivbT5LWQsnPE9M/UnOe1iutEfsgtZzxOqjrf58rOCFi/DGwY/x
/aHU7EPJ+vKuVqk47OmSJlJcVj5VpTS3tXFfX1uUF+Qq1WLx4vgAClksawlsjiTAXlvXbZ0K4GKo
JkKzRezHzgPZPDIFhvkZcpziU/jStD2GDNDhQv41Pne/cf9JVaRsdYMQJrwwXonrbsMMw8T/DhUu
X9MiKrfzhNOKZBiUevaHAs3s3/O84fOXnMGvu0EefoY8KTx5xYMtIbExWwL8qx2CQ17UB12UqPjL
/ZoVJHr5RsQ5ULpWuApUdSg99J7sEtRUcKxNz4lbJ2pqkyiNVFEt7eF/WUo7OGi724fySlvJUmuF
vgdvWudzD01OW37nF2/wR+elx4qiTt18UuKJ9NLbzNPtp1q0hLT1Q5rpy0KqIDQB1J/InsfD24jA
MKFrmSJMqlpoKZTal/2+ug9CbeSM8APcB8wGyPKu88rEsgjCTQHwk0vxf9Hu6HlYZ5urJsixopqz
rYFuvD8zB5BDh8rh91gVieLJMFQZVRxr63/WvExhnu+va6oXfxe052KzYaFVFxcVgWYaf27jPxv7
QfeXswxbt7wWodITzWt9qr4nnOADdLhfi+WfeK5XONkxHnTq8Tw5Anfo4iSO6L1FH5L1nlMlkZ2F
dUadfIUXN5garb4fS1l69m8g+QRKociEfjZ4B+Da4FGUjlogISJdOb9MuBcvF7/FjMFFBcWzwOc1
KIGwm85AHDShN3yow+/YDk12zqMOiuMIYhly35LkVPlbBJy4A1zJFovbantMXy8bbO7ZkWb6S5N5
LqWWF9KrWsU7ihU8TkFcOE5s3CVDGkGq01Vg6OEB3VcO+1q+KZLD7t8T2Zl529xzLQ9EyWdNh74O
Ytz5lIFrwyVBuB9s9IoNz5uMV3cX3ukE4lB2HW3MZE8eVkRIBO61rY2L8mTHj97dfnMpfGChhOGu
aOj04ffM+5DbqRsFvO4+MqYTv6MQt3ouUQ3dnGK8qCk5t018cMgyxZjSYfCxuBeGkyxXAKxeKy2B
P0ZcSNrN9FtemsOCr2AhMOdQpT7B5AaIIWzhoHyYXF+BxDtUDT33TBUS/ufciXp98iry6LteB66O
FeR+GWenL7fSNh8SgdFf40mYaFWzdBd66spI4dUD+AIEhmZFK2X3NN6p497rcny8IjXus96wvZdq
XE3OorloVgeaESFEdQKtYoLhc0VO69wp2CJhCDFEdYSecjColEB1CGl7F3n1MmM8S3UaO9a4TxLH
haLbFFssSEz8cfmnQNjxoaHoaonRuauOV4uJTj8MGTzoQRnbpJ8iMkZomQFZq4T6Jrw5BNwAlbze
bFmb8H/SHosExJpDnmkhATt7xvwsSHHsNR+kgWv2UCSGjXHy/QfAg9cR0bsObfUBTdmaAIdEIGdW
jY4K2Gp1FpzstU99JM4aRbdLKKumwiXvmQzONg+3BIQR9Mp8iNRW8twyygq8J7Zi1YjlEq5s/XUf
nfYZ3dNYpiyCP0HJ7D56EpVuGiVShbPpLRSL/7+W6AUSbQ9ri5ioDjf3HahiUtOYBCN2IAhzrtcl
gRAID6fqq4WlnsSlj3Wy21mdUbRuXw/jjrILmtOOP4MOdPtkVBu/k86TTi9l5gg6Btx0Gtp35jZm
9jH6mq9aTiemgxzUIbCI9Q+iY0+Sr+BJQGA4M49oOsrUzwNLXz6KzQGm1uGhChJ0tSXJmESUCsh8
Br7qqM9i91pVgmWrHJ6OselRBrk8Dhyq6gbg/OkOP0UTjJg50r5ZVqkk/2Q/E//GXXH7Fm0QUWU+
GXZQpvPn1uXqUL0hecFdCMIPZiBxjd7b89Cq6X36eQjWnjfYOQUDjlNUT9jYo5TjOftMI6KtYKuf
ud0rD8zKDjc+we71xCN8HfmqYIpZpscGFMVx7vPUVdpzTCbaU2CCAB6/KQnIKn1JVyChvTk4bncQ
8Ym22fe+sTbrnKVz4eqICIakVYjAniHZ8VpZUeJzEPXAwlGTJbx5wy3I2hzEsypT+j2OzTy/fWUi
xa23StVmdwZuBFNRhNFrxZE1VR0WyCAGsHyOpzhpbE8BfPNNMZCiHIJs/cvkZ7mMGEbHEo0mdZ0r
10x9LgrNsYbiYvyOQ6Os+D5vQ4XdQVTFA2yPoGNxgYjZnl7J2k6Zrj/XRIicVY69iK6XEOFeQGte
CDGZ2iznUkJWHzIjGBPPXTE9XIDvuSpIs9XtM3g+R/LATvDGU4E8gFJwLGMbHi8e/wwcDod1Fn+J
0OWfNjVVek9oQSWOi+Y4EYTMa02QjEqlV+2agQaydGXHZCRR1Biml7hLwIK7UUAIWbyAUjE3H+5F
pQB3mN6oQZs/BwGkItyedK4XOLVbRM/WaumQy8e/rxR8fEf+6AcarKaicAfxeZ5IfBUn1x5ZnSQj
jnxWrfKtswsLPsghfY3RNwt4Lqp86TCcWwpVHQX6v5YNwhaebBuVm9HmYYHPR3szUihI5TEUgPZZ
lM0BTPFw6gcI/gy//wr0Slu+3EkyHqGfhJusDS+q4WSyQroGnQkVCYvF9RhxIlrpr6qdAgf9wKz5
MHAUVTUeuevj4ljmMfIB+ske8XDb/VJrI+CVqMVGKRvoR0+9sV2q1soqH4RXZ02WunYVVqvfrBOp
r4hupvE6/eNTJsP255PSAsm32WcsRXBH38HraLs+fEhA1dkNnAfDv8Kxd0a55RJzWvSop+mlLDlp
8u5vjH/Nex+d2LVyrF1pvP4qBL+9wRgFLcY0cx6EDD10zrw+tsfwONoFZAKfv76p3K/q0fs0238r
nYfGehFxklPQOdMAZox1aBtR+Im8N4Nmh6BZmLbNa7oPpL+SmFKUsQ7dztbGure1q7KLdYKUDnIl
v/s+80j+05KF3biuNWVdKcEkZl9UXj/t7O3ax648pkLZkSX6cmdS+AytFAKGW+iKdjqhAJPm+81N
dv0JSX2yjBCGzy4hV74mXtCrJm9do461IFq+ZbdOJC5gXadq7tqzEW6Z9KKyZXEYjR4NcDO9/al5
12egLs8MDWp4JzVgM9QCqYNjUZTbumyJAKq65RVwIsaGYtNBdYN08ATSq6hL5NI8Fk1W/+XZul6W
I42k5ZprazKwdRhULrYS0oILjjjNsAMmhjfegF6PRpx7e3L1ShbYU++9oAsgFPEizlBa7tELUjxk
GpkmAK5mUluujpGWTojJ9NqIFdvvvhJmmI1CH55kzxHlB8xVjrQM4Uv71CvAatF0aH/8nu6i3lG9
BaV+oXPB9M8Et5m7xUl818qAIdza0glHNtoXYv4nLq5H+Iz7xtKRUoE+b9t7M8vJDpzysvnP6tec
VBQp2vonq8b1FcLkC+hkOn4ApMOSZ73tVlQTsH31CoLkhJEASylfCYTxareSpSpUg7iBiiA37Ypu
1H1HDVsklfkZRpepkopRjXnM8aMx/b9kvd69bKSXdz+JviyH7wIINjNoJOKZQV1NGdL452NcqxgI
xByB8q2IMsPfgWPVvtF5lKOjKvnLyksFtYvOfTtB1Aagra9Nl6Xj+hzTVKSXongZxY7R5sDo/ufu
/lwSWq+Ze6Z0MyUPxVU5yXNlrYUeEJqyMUFzA1VWm9bJdvGzt3rst3Y44J+qpdrRNCM+4GKWQOdR
VRvJDGCD5bk0UhNKYmnzG0Q9jfJ55/SAIJxnwWk2meVLGY/hhDk0UPUKHbm71vipkyfmsMnMb9+1
0igqpc730SKf1B9t7XAIDksje1tXdpZJRUDxGghW0uoPO7dbMRG/urrZF3w4YJ2YXCAdAhK9A0G/
MawCntzk83W/OJPvGWS3fK7dBX1Q2Sn56QaTNB3wMSEWFG1KyYR1KjKkrYYGZ9ZI9b7+DtSHUA7p
ljUXBuANkHYS43owOjC/WLN9k677zcryzoMz5cuyA9GzSWkDWUYKgDjK+1t6POIHDZ4SimMDQNZS
4H7VxudFYsVbTrawJRtN2J9ydnm40bofgEcGGXJEVE3stnIc+HyT4+1/sKgiSMWtimT1Of1+PI/p
j3GTp/FScaeMQaIZKaRh659GpgsNqls2O6mua9LFMQqDZHY4va6cctw8luxs5Y/wZmRNoKguH/LV
ShDdDhfMPTXhs58dLO9z4Lx8TuGJi5m2L49et6YtYQnvk7Ag1KfLTvGjlVuMYks/KqxSDkjbdIQ9
napL2iFypTpWrpkS1IdEcCn0ds4NGts5Nok/bY06NwSXBZOpcUhBRC/3Ys4/kQTWeAwoC2O/XCdR
GAOuxXum6IyPsn9DWFPGvlRZW9qhuTlsLJfcgNATNXAq18+g5WZ4n46OkcI6EFRfSJ4K6/bru/d2
F0vpbVR2Nt1s6vcMYGJx8KgIUgWSQctbM+Wdp1yDyM8m4xXp6HxMIvlXtHQJGH+/2xoQthB1vDPa
T/No3XC6Kq2GPCoHp19MnypqwMeqczcuymS87KogS5/P8P2Q/itgJDsnLPns06dlKbKBs7wJ+/Ch
8WfrrKVFNqccisETNWszgRfee2H6WmtLfG7+y+GOhkgF48W/97z6Eijr0MALqK12/LgktbVHHldQ
1sTBkbj1Mfg17+/UurzDaWChzvbkvWa8Cs0G3dppUxetY5j78B8vHhUvrLlfz4RsmS7XzzRSGF0D
AVI61y6kaK6UOrzk8JDMpFhROGZIB7MneX0dmSTFVELFREFYfA+I4jYM9BCusHWq9ojUw6tyvAdM
ONL/K0yIRYQCHN0sKk00LVL/W+FTcNohqkiRpPKQGgZxPIhjYW+dCStlH/xehjFB85ekBqS5oZJX
PLcDL45iTpWwpzFMQln4r82OriOfCtmi2bGA+Yqp8el2Iquwyuupi9MPcXVAaufNB7FKSuHuedUq
ZYLSiyTxB/jxf1KOIp8acuobMw7bigkmf1VBDt54YfV6Z7ABFgo5JDapvcPi3AaQkHuBwG/jGJom
9ZxZtQ/rnJ4+FxyvLJuyUmgxLltN8SEhJqUbqukewVG/HuvfPhMW1/twVjSbxruq+kiDEA6SMSAS
dt8paqEyUcRyLhORzhFG1GsMP1cqrYK1BssxVEpgtMiaBJDn9wjU4KErBTCCqD3XzYy1UUw87M5J
req0lBhsmEuag8FucxYjqNUtp/n72dB37IkHTa3hBNyj3D9b152/nBjhf1DmMQ72WzsxnYCbXnTB
u/rrFuhwDB5rtYEqFKAIQCN32Ka1F1kpCrcgFxB/DM+cSLqTZVXiQQN1YWqQ7aDW2t98tL7PayIN
ukoU2DWsUZ93NSQtTmpgZTI4KQaG2UWtwc9rf9qhT133m7pARoVeEZ2Ql+jZ6onn2H1Zx/Ka9gAA
NjqZ07C3OgnzykwROO/hP5o37cUHiCyLlBCV7zHVgl1YADy61y62vMiCMihlppO1zNqAa8nRipx8
BqHZpMy2M6CthOWSiItNvL7TPa7XuSKUeL4AAEBohSBh+CApMKPurrU6yhw8JUYcUVPT6F2Bq0pO
rUjI8WQP2y6HAN0ucNxIyeLBVSyTfG6XEubPoe0/K+kkwLUcDxaQLYSpw6vh3RjT8PbxwZ4VI2b9
52jhTV8OJqgGEczOp5YPBk7YieJQdgz5AiLtWqQ9+J/NcbMIaoxUxnOL7SCkouVHWXly+SNA15Fz
4zpDxLQrCfcO2/ZbAZb9Rz6ABOZ0GiRuSATxWy13CE/xuv1odIsZ9fqnSE8EwTbs74WPUyfEKDVi
+K/FlMQFOLFoAuhBy9oTjaK6FicYNcoFbOxQsJ7ldoA9j6OLb4GbSdLlU59mJGFrLehreDmaAXCv
ucEVJg4X8kKHhx0b9Zn8q7jFqIGHl796a4XeABGNNCzuqxTyRonlWb30tAmu6s97/8ylwdArT35T
9NC1fxBd6ip/yDU1dluudtgtCRhjZuqAHF3Jq5fG/RHsr2npF97qRLfLdL6vEHctWmzHm/p9VZzK
edaaG21wiR0RlBglKew7KOFP6p8AJl80TQwQrvlJZLBm5vAEVyjOUOK5KOga/S6HqAMNVmFYlNzW
DZKxzzjMJDRa/snHydwOQeZFeqwF7htD+Blzv5nTozor5TdNX4Q0ZpJVdiZl1wD0Qd786Ww0Jmy0
LDKm8gtdIRdo27VRRxHXfMKjlmqsJrUK8ZqmbgW7bYLh/j2s9Bh0Tg7XsSZgcF+3P+cpnpgoZkWb
wt0uHgxPEdsv5npHrhUYweAHSpUfOETiOkY71yyLlwFltD0nuaQ2gQ460oYb/j7A+C2p66ABFSvW
DbEeyS21AbfIXj7s45VTat/5gKi4zD71uZNV/BNvsr96qqT5Me2NBKT8E/AM06H7dv+L10auxDph
KQgcxUAo11f4+KIyaTfucKdtH9I6HteccwYoTE4J2W1bE0sj8b442NnvT/wzX+ZmFyC+pRSrCiWm
RtBuzEN6Ins5/0HxW7IyvnmR1cwdVHV18PdB4ZVLwWpA9YpZo58/Fqb6bED5fdY4DFBhL4msxDHM
tH1dpuKTiQwwYfNuS8E3L9goauJsyyH204OF3q7jyxqLE5zVwbExlzavHkx8ENtDAh085tU2HcDX
cYmGYo0SMxAJC7h6UUVGVsfex6wsHQhI8KvPt/eIkCBwYxF6Z/gcc6A4A1cyqCLv6D93t6C8PIt3
0F8LC6ZHrhIVy3N7HgHoSy98eAo0cmo+yv+3DzxRHECoud25pwxQN4BmNay4kkQktRmnTem4S9dj
meGmA9dJqOHPseYslJO+cQVxdGoZ7cJmG0rxSyCIakq31nKVkRhta6FMijsHqDiHjfB7o8BvrYUz
mWafNEt/974ZmNyQ24yqmrD6PpaIDAYikijlUwavLAfbaVCIaQC5rhdy4rgpp8yt1i4fGTM/eViu
6DqTxJuwEuXB64uLAX90rvn/3qm+pZrCYErO43Sg+oc15SjUC4nDuk7u3fiUYD5scAAE2JwUE3hl
cl2Fg8VCuUJBI/BBUsJncfKblK+qxQn0Dle94UZgVah3nDb1VCxIKDXkOLXEF+nzv3Ez7G0tX+98
7JTaFuWqy0x8vGo27xV+EFAI5mxspoEExsLD7EQizPVe17qznXeFfJgu2G6QUXYPgaUVpv13m1Op
mgM/x+uROJ9l8Ll+8/xQt1JL+ZuR0nAFjajd8vlAEIiK8NEy4eDfBTPT/7bUQFjGVOB2DweJkxdp
pw53tTYBldL7ON3fNDE0t9oj9ZrUlllU2Pa4cjxT+Xoy59NC2WykNtqPDNw3ty69qIjYVz1l8Oq+
MhR5ne+Ycdcn/1M89BfJDzSwS2D9LgEWwYBYpkzc4iGhC3sQ4NX/QhVpAeMurR9U6GD5+InE6pOr
iCIWM73y/LwON3H9n0IWX2EP4c5kO/Kc7+8Ts36QNqitqlzJBUyQD5oCgzvym7/4dwwkpNzkmqCq
61ZrxpMXPC0/vLKQ6DswGe0rrEpT9yZ34AvwsRAWdipt+iAUs8/theUzG3/chFMKH+fpn4lZFpy2
wlTQWjpBYGFFZBZ9nA5osekqyBA6jQpgeDKef/pVv+4us2k0pNxYzIxCe0qrCYoaYqPqogrBDokS
bl4gBvneZBMfHSsr/o8knPdsvxUn7duzNBIpCQX3CMTTO+4A/UVHX78mr0SNtBwfAQMk8t+Zzwfk
T4D5zLnQ+f/+z9VweBkLCSz1aQSYvMx9Xt2/PMjLuaFMkUkb7pqal9j61vLU0EfLiupIdYwEcR4e
NdgExo8PwsK5veeCi2MN3xf7BNPtRCaLAuxhCEpkfIRzqTdnE45KM46PGwpo/CtENgNvxlb9X0Cs
xcu7b4jGGniYQ5ng6ox937KvGM1UaCsl46Ao0SEH4AGeJbrOAd5ThSGKD92lS5skgHuPmPZK+dNq
UGpxwBHviq3drxOgitQeF4Skhqad8dsL21G5tPrHGGVgcKNcy8C5qJwgF6U/B3ndt4Sb8gX+YNEr
A1191CS2TR9EZkNx0AhiWa+LzlLTfAQpr9F06wMOaNxozFVHwFRWjrREAOsV2MYHW18kopDqmTNR
uHSKqoGZ1Jsxf/YwFxM1BvI57ZhRasi32OkyoHW0ZCBz9JQsDC+njWscHce0FDAZAW6P1IQ+Xf1l
qvotV1dJtLiLMw2OSrurYlzE9V+/0yd8s3bwaaotaN8FKncoBRvW4QzW4AYYqFCrhHy1zkZVtRyV
hJX19FkPJiEl9DxoDmt9zpWBDSwTEZ4KDZXGB5bTZH8vJ/ybV/BUJp4YhDkCiIGOFTNB3gK28eJV
EuWrd5tdotB15i0PeWCMJ12PFJPMNsAm/PhqB0PZ1CsCkzlg2uWQvLa+Gnzg0dMrcW0kE8Or8NJO
sxKskPfn9/yFW93hhNznvIFyJHhvqWhcgEtcyObvDpYJNWFsOXPwZPYFvR7rMnNoD5WLWHbUCqbn
REbJL3VsCkN5VL4jCduISOJyPfuygDRynnJEUQAw/Pbc+erlbs6MMS1xtNfFE0dDuXczfmLAFIDZ
YM7XPJFjwrj/ipy2m91Dk17BpAmMJjGO7hjcnFu0B6ZH5hcUpJ+9wpuoRFhdWqaxDwYr42FIo7YV
lyz5v2NfEXMOQ45uQV4xnnSnThcoydltaTRVRQh/y8Sq+vlKsMTZkVbax8wpJsby/s8coNc7RLms
iFQIMud0HuZeX/kv0qAQ6h7iyGVkpt+zXQ+ul6hNy32pxyxoj4m0SNp8IBFuF6XZdBIjgSQMlDek
NJqy7sMy+9FEWaLhotI/Zn1VONp7S2CMXIkA3n9CoC7doXg80/1jmgNUna1S1/roaQzJmEqYCEmM
h/TseOilcbYAlb3iZBfIxLjR59vVGv/TQ6L1Q3fkKGRhlhaEkTzmYoYxAzLr3Dooo93qu8fuaNDh
hvNZfUy+LBNoyBw+A9vIRxB/EN8GyrPUBsvFwK1V3/g+5lKKflnrHdxV0P5be1YIRyw2d5nvAUed
LLu1YUYBfLZwTo9YokedtWvpaWlny9ID3OOa/knmDgAp5mBXFNgrG3T2bRhyggtx8pETmtSFwrm1
ma0zIkBQT5U00dvP/PlPbkSlPREFkQC79fqGSANR188RWZXV4y9GgcgJy5TRkIZEJKoRv2dCdm5U
Iy4w1bdiZ4hOic4CWWMYPD0VrA9ixz5tTb8FE6Vywv4Ye1tFPl9MkctMsocsWlfTuJRSH3/WTKix
zb4jFiW5e+DjGhhg346PGaJR8ddpF4u53hJ/tQhOggRs8UH1O6K8XhQpvTnU6/ufCQ/sUvRgQVYP
X0znh0SlgLRd9X0LtS93pjjQbX5vQV8Yp0DSLRfykiguCvvu5itwVSMlKkdgLDWaZymlP+R3j1Du
hPIc/ui4VmORZ1l5Kd+M/cHp8fxG4WpJHIna+TgmouY/EYtiKfHOBL+hT2yKbgvhfr9pVlwintdh
Gzbq1zNOIPne7yxnB0HSfJloJYF6EeNGGpgGgWj0VLNy375Fal/s+/7MU1VfYYWqHWyP9iWLR/Pf
TOVB1K0PIwrY5PaR65DAdzkrNLi3y/k/eaRtVb2wuxfE85ZKVPsNFE4+cRMAyqo+p2GqoswfYEq2
prrOh0wMads8uo4zafSuvBdld/Qd/5XyM0EwvKAmppqPzWUaXVBj9hk/Lg09Tc7OA5qmXKkIFgqM
qtMq+Swk0xD+ta+YbUjFT8I8ysA06gMmhqJuO9z3CPod2LnCGPzakQsgMck0JSAwaXEkj+w+PJYI
F+JWEUAE9PQk+Uj/I+nyb/qv8m29LaRAhcH5LJe/73FeLfeyz14Xvs65ouKB/maQNuWJ2xy2JCei
/rspRIP7U8ZC7Y5siPyINJUpg2+L+E5eifAsZEJmjFzbImHqqan7yOWFpHvNdCEVq/OU1vvuCetr
5KY+Vz4Z58F9/7pAt2w7DQkTj/SaW2EhHHccwUBw3KsveUDJso7lY7u7AlK3Cf7JYe0Cd8AaOu6M
8kUj2RhWngU0delExLJaCrSxp/rpZFiKGUMs/0QC0xrfRztGjxlE1NI5iBuStxaann2YxtpaUoUy
WladxRZYX//Y1hLY+GBHbpVlL3lQMXC/Fv3nAA1Bn+qS6EcXkRoIenQFlNHdEfUyzDL7Pd9hInM7
FpFyRZrMbaum3bfcRyijWsZ8w+C81El8ygJInh9DWddd3a6VsKcjohGx5bN1o2zfPtfjo+YKvV1r
LSY+cb2++zOBhiqoJh4ywn0e/5xtIofdQSdLbfvdQ2J4lurNa+5fng00lDumiS90KfpinS/fkr/G
CtVFReJS5T7MMjBPEyAZ6PUSUCJ7/Ldpi7mYi7zQ0R3TuFkkbx1DtpzgAo5FEnhgC6bdwWibEB5h
M6p+A6ncdv4BeC3ZVQwzVfd9wExGr7hmctIVrVpT2OBINoMzhJJP3NagM7g2vNtfaVBRv7lRzTW+
2VnFWek6gFJDrrRVmddHWiJNUPB6s9KiMLnhOUTncRehssWaV0AS/j+86XFjeSMYVzQIJcCT7m0n
1mxBKCxPqHG+ROTSmiMa9nlR86Bf55PGe6FCwGGC7E55H2OevSmcwE+awQDf6L3A/2vi8jF5sFxZ
3/oMn6FMCAlAvBsN48m1snoW8I5IISh4/f1RCRFEQwAqkRj3A/apD9iqk/XbLrWVXo3owWeoPHU4
vhmfcsg4NeL/lF8artcnPv4X66jFGhBMMbuTuvNdSkMhZ0eG4JWQ4Azs+BDR6Se1zeSvMzAShAb4
iIw5dSy6n7eQVoavXrUhS8kA4ApBUfc9gw1IIU+khboclu+EiUFX/VD8AqCRU29QnxTWbZt1nPpi
sPXy4pZi9fCHcNgxEQM2/eGgTXInV4Oaj9XjAL4qQwSlMsAbd2MiPXAy2uesNx1fb1Z0Ec14yq0u
uly9vpuQBIVPIuk0S7IKvRVJRfBCQZo6rS2eQdm+Erp3owoTla4tWg/U5FYzBz6pX55gUTsgrxYq
tOhI1InaMTQuj+T+nF8jssnn2HBVZgvwTusY4Qe0i45yuppVkWsUU7i59Atu1Qdii0MxBF9Ew8fT
ffkeZWOCg7+jupIlRY15TTzOJTFHOPphtKTgMlwVI8Ro1HydhZq7nr7sMapZ8WNTcdk2QJNFPYMX
Tm1GtnjzxnMWKIxFEraVyMQrEUlKoR7VUo8o/G85u2C5aAfNofDEYwLYsHv/Ktstpxq70/eXxYWy
JDtArAghJp0KrNInKgOvtVcPn2id6M2lC2TctDL6tzpiVNtvB7aUFDq6slHcqYRrxQC15YWTqpY7
nTqvhfP/uhwB7FhLmYY1iiZYFhKTJKAAbOdEgoSZ7Xna5YYgs+U3CC1ezkcakfxVmwfhwMWJ6nk4
C8lvr47jhRzj9A9uFxgZ8I/d48zIZQhheH3LzHd7b3kqbrUfMgnRhERQshRt5WVH4VaL8CyLetuD
+uPyPc+vASoPc24+5nkNWabv6BVtaTkrhyZQ0j9e5eLwDqw60Ho7kb7tzpCmznhnonNbhzzKu9pf
7Jfn7lGPyLkfIdVGrTMUBPnXHWAtzJomDh58sNTeA8Ofaa++RqYEZ/qoSUp8T+ftnvI7jewIEYFt
3h5P4EFzAYCLaXTNEGmxDeXoDDlLIYsZ1wMmUtFAm4MO6q7LAanPp1wFoRgqP0jp/vCcstXjI9vD
01NIpicsfmOQkzr2KeKhn81aOlxijBZdhXgXV1hZx80fyPjcvTdSg3uPmVYDKzAtNshrBProClhr
oqMLJyIk9DwbA6YfAQ+2LP88I7OB3ZuDnrkF/yPm95r0R8nR3zD7jj3gv+00JJbaBXqzauynJKIu
9lk4vKd2680tAq6JCyEFC0c8VvEB+FaiEmBDYv1UzX2Or8jxPpAMuuFNul7REjb0tuIKW14t/+Da
1BpyAQAH4djUXYnQzLzs7Dj7PnFmZ7WOLMecndqz+D4mghoUokUgihYHEI+Wy/62JVo1vo7ZHJrt
Xy1k8fMoeFxh/9hhcgdxsN5KxsEn0wgRLI9+kXsTXiBDJRtb0JQ0NFofFmchDmp+cotTKn5g5tu9
EPFnCmVnieMD3jx00/LBw1sw9a/Gsantm4SPnOHXGZcfBiulAJx0oEjybzM5MLtw9cwNM1uifARI
b2bwaIvfVUYrGT69VR4y1sI+aRFB4neuRZ+r4uUgtDqyxtnE4FuPXlW6V1qrkbEjy/fEHB+C2uRR
Fpe1qdFhOv/fg2djXPiP2WtnZtZ3N8y6xFMo9HZky539DbJM0VUnDWtRRMI4EIdkd4Bjxhyx6Jpb
MPJbKIddWlbGOiV8DajYeYAuFzS0zP1G6pDMv3cyxuWAOaOyAj817yzlJO41y1iiICJVQmXP+QT/
6SVeGAjsPEHKwz3ac5jVrPrL65YH8sO+zti+6GsfTzkrR8xu77lFg88GI3IBNYrzSz7rvvVRErVA
kozoygKAcwLVJLnnzaOW/a1USCMyV8YZ6JMb2FyubTAuMbL3m4cBBppTqRof16hbbSDI9qAlrv1P
Ukz1nRZq/JkSf/mxGkL3ajXAc6zFKuqgyyKivms0a8LGSs+zxfEBy3fMoh6aSTeCrtX9DI3bVHd1
gaJBttBwtmocc0iOiYefDGsN+2YpER3lU/+axTIqSGN+ePjbcr4lAyUX0ryMrucPzHciB5Xd2lQU
ZzoBd4Z0bShE1Guq/umkvZOZvuAFXCuFHp3pcbM7vVoCB6jrqAIGf4UzgUXFyiukRk4nmpBec5/D
onIG2mvF1jTPP1JL1b6yPNOHdO5AX9CbYT9gvehOQVDyW24euPeEaIREjn4HJIkNL/b5F8+q5Tjk
Id5cPjez5GHQnyXvrRRqJhOB0jBQmc9WYDFheqTG1kNL2VRmsMVQ1JT8jyrPmflZmbUQUPFncPgp
aMQfxIk5osbLkT4XLqAEYYpnZH9Mg9RYj5sy45nPN8PYOZrUZRk8jIN3OsJLojXrHZGX/MI7w/3h
EjuUP73Klww7Zxt1qIQ2NBWPkArFKHQm7KF/Lngay33W6XdkmW/F+3nS6jSkZJgCSsCZI0rvQL+o
u8A4+XI+jbxtDdzg6kVByblpH7Adc1UjO7VGQvXT3NTkYHFJ2Lagb5U09IayzG93JegN1RdsiUDp
tHa6y0OZls+rtf0L/jeYQUgSKHJeBNT0XasBc8RWp/m4VJ/OdZkmrNd56iS35pv5iLY0qxNHK3di
2FiQ1QuzvH/yhJcn7fdPM1j9iSK6y2vxHOC0EGOpRBPAwFrFH6iMUDYoZ6sk50cc8war6ddOekpN
0R8wYJ4QtgGoy5+RCtQBUQAW9D37AxCcIkDhQv/+ul1PpbJ6gEPnUI76ZPNeFQbdj96MLNoAQFow
DSYIiRiCxUUGrkZzxDzqtu9QGzcQmiPGeanl8SeF2o7ictoDkXbhK8UZxHAbC9FkDLcrT6xaIr7v
OeW6j36pB1UTgLFataRi7o/GSn6FJbsl4fZOMm6sdr8YW/eEz2nOxREYtTNSiFjOkHAa2kwLHFWp
EE4S06yHwZ7iX0qsg//4FKDqbatfQAp9TZQMARAUKGzRfqqNIn2f6bJ5xBdosdMRmAO3V8S1Hsg3
oHkO+w9MefWspmaVNp47CJF8SN9bIZWZkRsZpZlbeCCSOutQN0WGKxkhgLaO6LPmA3/xOCqtKqdt
/CRbfo74ojU+dpPwJcW3TpdgDjEd/Weua6ISrocT2JaMSHWcAjDMYThj6yPkr858wMSyobm6y1cJ
E7l1ZESepulfHlrvMaVJ5S9ra3iL6dCE2DaliWfjRamUpF0ozaRZdTiXAKmWbZ5kamp1fYYElX+x
nXCMcieRGu/j8Fe0a6LcKqwmOIqQOSuBEWu/kcPPnpsQgSOZRqvIalkCzp0Pk70LJv+zlctAGbis
Q0ndYpv3w9RpGM+2zp4oK6oyqhLiwyAzzxFbxuqydci+gRD3WgB4nW+mtjCXNsR0ihOE4S0J4cFU
u3nB+H1g+W5LrDrLoDPOWVMShIf4u7I9+GnfwezjxhKOmNs0FEfMDt7DgBEmXdUak2VocRCPfEwO
K6OovZUHDALaRhswtcDrnsNA0h8+4yciR+VEs3WuB1pfcyVQ8u+NOoZBAa1IYA9YAi0ytgXKwOct
8iV2Q8klz8KmEJ1LDt0Zb1co1/4M7qvh2oTCX5GBMYZKKEyGxCFRJvnTX6c6TdELlMHuNsOHfwW8
e0mI1RdmRxIUwuyIy4sNW8zKXGW/sdpyQF3fQn5WCHSDBvFftKPqZx2DNnz+CrVoJ/pXI6EVJ2E3
CsXs4ZQMQphKtByrP+n+TKYSjH7dZOMeLpxxonAZDvoE3ZCv1ncF12HHvWDxD+goglPf/1utImko
suGGR2XH47qr9WgAaM1MvE0fOBM5YBGu33gsDEBv1mdjT/CEp6NSrKF2IWFiSn6woeo8yOh7zOeq
pGhAYoI/zv+qi9RY0lu/QZ7UsXSLjtjks6rs87gykEGxxcNPYbT6mqp1oEOYG3O7RtvB8m5GsqOi
0IGGqcpeMJc9uKyiDSxFxV048hsersh4N5Q/xvPc1nFxwsuAYU6R12mWP/MTpxgqu0LV3HKU47Oy
M6945lZyP3l5mtKVTjbhEb5cYGyrjnCSIqFQ6YecQeHOCwurgPKeP0mn2FNFIkHbTbdhGKDyks16
U0sUZx6tou3kK4tUz5Fqjtd2Nx0wDpK8etdvOpwsRl3Jmn/Aj7u1iRMJ5ALEyFQWzQ0CL8jVSJM1
lVaZFtTpYiCSDUSEruC66C9yEklL6IPMyXV50z63eHTi1/0zIfP6bZUJHwsOO+Km2vAI+58O5v3e
Eqm/eSPAwVUOwC2lVjZFrJsxFAf/F+TFK2xqmV5XdDM5YZAK8uPYlW9zyGzxA6nJetsujWWHBl59
pUYUyHzp44saxzGhtNFWpEYN9oij22+pYlCCRY3S5khm3thwe2oWmlrRRzkVSdvU/afUFmk4u1ti
5fu4gfuri9lCCphpM9U48lC2KUdd0pCSKNASAu6z5yomGk5RuLAuKPreCdgvTCk62PbB+yv8csUc
sIeOQs5RdoHyfioZkT07BUZaXpUQ5V6i9/D+LtogaF7gGvAm48yHnAqHDUG/eyGtVH8QFP5FU2GM
F/tt2fuMneIqU3wAIfjIdB2yZHJQguEB6540JdY/8o692Ujs+rkwzky9IHLjJcm4g4Mswo916Rtp
lNKCNtxbpe0Jh/+DUHbykzQJqi9XyYwjwg6tMwppNYnMyTfbRZfe7Lf/4Un2UrU8Gt/5TExNdRis
YGulrYNRRvSVvuQoCH17jriCK9FwXoLnWgooZRwzNCXDi0Rp2GUNrhbUob0cLcrjsVJfdkUl0ZQi
qjDyBU+KbDM5Yt2MPu+7vmq4khLSkiQQ/QlCuwjKrb7nC/X/AguUMDUU/TXmuAXzGQOhQRjA+XbQ
LCL/Q99xWuv9L9AGkfWSLLDzWoOLNBSeAJzIgZzspqU6V8DDrNJuQ+8kEUSBZdotOyO1+dwKeYvr
PAzS+WrwVqLSE26TxBHikuxVsRdCjvhnPGeAcDcN/5PwuCKiCZcNiBBfN0mmcIbaCgF6dtLkP6qg
OrXHWjt+GSbuYfUOYFzdBHayI5FLq7/CDCZsNtFytgpv6qJnQJGnk1+D2THXdRPpSIvTBsawK5fp
h9ies/KSt1pxmf9X4GNTBM4pqNRXChIelbFZbAtTJ9ocJ7Wz3W1XEV6Mxa40r23krDxZd20e6/yF
bQNfaR2nK5VGw+ijW1vIfimsItkAfTqszOsoFVspFwF/uHjbN/p7jFul5cWx1H+oxUMy5BjBSdzz
jCz9GPo1sosnR+JK5T0LZ1G2z55aE4uIxqj034TKn1xyKstA4YFAPN8AcOdgvDU/X3KcK2q8icRj
zCAAv7Df84IEwvuqDjj3UXQSL7tebHQ6Benpd8R920sT/Bm8AIueMspo1aosniQG3O17KzO0ZiBA
fMc1DJP3SWU1DxY5yLJY1XVohphCjmPvMExlflC2610apXOVllF8c7QS8MVpgJzUI4LbsAP74RKG
GY4aQwqiUNEe75Jty2ZtoUoO3v8WWPQxjBJvc2f8fHhXa9Sqk+lrvPvORD2MRG4eVEdCiBtg2VEW
TMZuEysnI3kcxbYFZRtqDo6EQLPxPGp19+4xkJ1MKYjJsooj7Y2lRNm65I4Rxelf+gH8zRD1j+52
PYJi3EKLcpY8lNS3Ao1qkwTW2w9VnGf+nj0YvIY95ja1AT646CmUZNeENL2wAdW7ACt9Zz4tLAbI
pSyJwu+OLMBN/h4hqL8+2JORn3u2MOryVu885dqBEeYwXnoWS3ERLf7EhB8ikc72cwKbAPJVIJKN
tfIVKe5CGseeXrgjaYZCbwdXRiV1wEDQEy9lxXMuU2S5dP3ic0ySS13j1j5gSkmeVWj4Gsh7rOAH
WsK1pY2Px41cyf88zyMwG61XtSN/+16pFRx6d4Orb0xofaObWIGaWWv5/eVyJ0KvC4mYbmoVETfP
WF2l68SZkulG7Fwtshke/Xfo1fJ+dKXND5qKEFBQRAxeWGE8L45evty5R59lPSbwxxfC1hk2jYdc
GpVYA8G5hq8zZCVF3chO+JsYcintAREOZHzJ43PUcmy5G4ZEv4k8msxknFENGGfr+qPmMSoTLcrR
NBto/IzgEHBLmCtAO+y9EikdEtr+r/qhBVnGFvVlvxZWdccxXub2X/JC6nErqbJ8HfrcBe3mt4z7
kvexqhUe24N5vdl94zbgxqJb3PG1lV1VCWgLwdxG66sxibW6FtrE4dvG75w8HNvHthkrvY9UtN1o
Nvf9GHU+87Jj8Goh7qqQ3fahbJqhkVkQ1EqSxbs5OkSWkAcjNsQGDh0papo61NHCoeCWFNsJqdpx
wZ8y6zw9tZnJt0xIGsogIPHf+gezmxvkHfYfQvsFrpTISzfnCp5oFc4LrZ719tF8ytksbCkK0gWX
QJ7K0+AEiW3pZ0Pt0dqoCOcfQC9ody1m3WtjKlyKX760RE65CcCExDHvRHj4X0N00qNnYXYwXcUI
vS/g90I2pRNs3QP7asMzIFK/XZdG7jBqlydglfH1MydB48tXga3sQ9Ij4W6ZS3O/b6LbcwqAXCo+
pFsWs4GkNldsnYb55typcrM3ox2g9VRvs+ufq7Wujrl3tV1CPG1OIkIzCKIMOTIkq/QooWmsMO1f
vBaJmd+4M1OukTfRxu+mtaRTecAvvLsIoUBWgg7aG37nOdnlvhV12qe5Y9C7p9x+PHW1gNz/k+RK
PqVChfFM6MxF8tWnnOg2M2JqhUIohj0A8zaRxBdFiNzHRVaAH1sFV6jcEMiTMS02UqvTKjVS+6Dv
XmMQoGtRN0e7JFzRKvPmykGmV2V+HiAFeC860qxPCrtBH9OB4D93sA1Ikkt8HlpoCVXNA9n44+T3
16Z0fecmu/WiKjjDPjek2doDYjdRjkylyo7p1ttrBoSTcaw8Nf36p3NQIpQI0RFFbVKKca+LINa6
/WKD1Edhn2STYHapvz3Do9tFuc5A6p0N3HoC6+jO1dztRJCMkv0ijySR13/1Ck8vvybr4kugnjlj
Y5QGLujxEtWfEonHWJsQw9lxtTpcqeDlCV41i0Q95HnZ1e1lDC+bh5pCSTRdZAzr1GziPsaS1Udc
uCqY23eItugZdF6S/BheXzckuV2qINYMbegI5gCCDgpfwTVuwzxrRdMPd21FoknAuzwfFtuW3lmh
FTC955npnhNkL9S6Jsf2JZSXpzlGd6VWmZuHBSJHqHDGIRuwUbwB22eqGCpsbZ5N2MnGwsgTw4li
sNe6BNq4xj+sxt4pQ20LkgzDTWpuIlngsqt2upTwP1agwpJ2g80lGmQMAj7I3oKJgzJYpANAnf46
fPnGytglTQRP4TG0GsItkSY+X+YvCG5yMFxNwU2Cj+pvRBWNsFB+2lg6ENkNeBtf/IJIaBIkb1zA
QvxoiE1ekh0N60BprNS9hzHD4heWyQdO2GCadFJAmC1dXisz6+r6GPhSa4rxPPoAlmkZrJx67sEo
fNKG1qA2khlsNrURCy7QhZH/slioahrlRX8VNP1Hx+DgsS9ivb10Bjl4Xtxwl400xV0Cbk2Jq1Rk
xmvGz5/zxlYJlMJj70YIypBlmRfBQY2kzKZPvo5h51J1sEXd/CG2vUjuXFh54A3Xm9fmFoQwaURU
3xdMRS5s0ctNoe3O0pdmv9I7QSdPf5Rz6QIp5Ox+bo8El2s19zApOiDbxtZTb6fdqCmaToW4PLpX
f++z1SX9ZGE9Rg7iGltZkoRcKDkhI2HuMINH60aEWjM+2fyv5vl1IdI2NUFCYWSm6VzHiyY6Cqac
H7TqCwB3LPZUYsDPR1fb6Nqogd3f/cG7GpjS0G9mEN3XnjImkVjuOmzK4Jd/OyLxAF/OmCsHy/St
oMb8U6SpZa+B4wjPNJP2duK6GnwzSRdU3R4WH//EbbeVxNVPsv+1velyOKD3FWE1SEGe1lOKO+33
evSQbPYQcYwbCSJIk8iwmqB6iK3652I5punye3V+5dI5b3L5QK8eQ5OHMNhS3imiipFEcBl4Xy39
ZgXYUwgBx6CxZ2k7Ke/AI4OxO/zI5B+O4hEkSLVn/9HZE+aGnCvrD2NK3ZQjK9rNhGiFhYsNpp5Q
JlIGEfoXRCKfaXJwv0FHJL+CflPHe0RA+Y9LipWVSs0gRT4EWUQRn6Z2kETtAkyS/ZLBJG5l3T9A
KU0QBW7APmJAqhgVeWYms4QrFWseoysOJdSEFEZTCSHg85X0foooBo/oUILZPcPO8TzEfKyN9cGJ
9i9A7Hpgvrx0ul50SoZcM7E4Nby0wZg2AMI4IuI+CsW5usbVVNGrzG+mcJG7btV1BOxeUFxhDZbv
txTm3S/g4wrnDh6wYnJtduMY69b5jAaw1V7jwWgtAXn1hYseVgheANquaj0SeehoWEZine1U86qm
solAH2dSy4dWEl2VTcbbxV321OGelaMQKGT6S4WRbXS7TnoFtvF1PHmL7IhGirSKny+l6njP91l8
P8vIx+A7Qh6r0ZfdI2uIVyoAOdwsXd6avnc7eeI1sAhILQflK2he6ChsLq4Pe3uyxGc0fhmJ9ZWZ
lISCNf+f1vW9N6YH82iplicn7DasCiMlqMN3uCkFuC4kwo8rluZPpUX69TVk5/GPoSKujgnb73F2
T3IggGkzJlzziPDk0sGQpzSA35D8Z7OsO/liuTRfQaLdwRvm+VGnnzD5BpmwtIQqiC8xn1t8k5qa
13y10ue9ZHyBo5xDcq/NCLsD0MTkWHqOA7anKUtMq1HJJcnYeRCasdjvEUTjs96pvQKIGMwN8ord
lgULyqz08aVggrA+xXn3b743eU5sxgOZXJS8y4XKFsBmIxHesLppi+yOkyjtEef5+0Kmf83z/RLV
i2pg/hkZgDL58Ah1CiTV+GapM8SmitqSNrQyCGZIYCpu+zbSiNUD0v5xfSqhedPuZ5bFtfedSk4b
IWT06KEYH4mcGoQeJEIcFrzek4D9Q+C5xezGcLlgTPpZ4WcA7O6VYKjp5kpftAgpsrNSPlESZwIZ
Xi9yq8VtbPE35MLZhiRqo+0pT6tvQcN+6DbVXydV9VNojAjRlcdfdFvc52FWycG+jgxTfvBXsQ1S
UhlNNBO7GON29a1J0Y1GykghiQTrPCC/QIHnd07qjxHCFmoV8GRT0QXbn5A7a0AuwvEokOrBQpmM
3RmQYc6T9XLlJizVR8ROX3SHj40OjfPYfDgKE9bSupmOwd6ubjGhUPr48ZP/JcpPvK2Bj3DhWAv1
ojEgUrrw4QSQL1aXhhxcCYgsbEhdidTH0tspTPEhP4ZCqi1wz5Ox/WQyIBS7UkWk/Ia6zODlIIRE
mmPpg211CUgi7zZO+HlICvBQYwVR1uqLRpBw+fePf5ANp8UsepKBTHueNE2yKSgJBZSgyOc8KMIE
AB+VoaT0V7eyRMdmo+mWCU/z6N2W23Ehwv4mN26y98JvgwXwRb+ahadgzFUu17ntQ008ZI++u/UM
aVt19JwPi8ly5qQUSI1Y7uY57zgfyz1t5enaS2DfANOzIjM2tjQOkMrOYzKvIJvlRWvS0UwMPAkv
JsqXjGkARaOC1Zkh+UJ8PwMjSmeEmPxQxB1PhlmymsdtlF65k8WNEPK/yhy21A07cWVtOz7Tf3NE
VPb/ePV3QcMRenH4B3xZU8JWB1JkUplKf+1e+u6AXBrlJpKXu11q03VVVqNxdFLaN3n7iVVdCh+P
HESVA/z9lvuVmbbBft/uDrnGchQHGtJoZtfuxHHkoaelpubzpgglMLbUVCx2uHJNPTgQryrXUzJv
BE8vbGyVwPAyN83xiFtC3VpznvartjKBxexRcC0zJYU7fXwOEXGTlSHqcK8mcWuec7oYSN0ch/g7
ezIvMulg9F1hWKWAQskufY/1KRZ0AqEUYUchCTmHerj5Z8RZEtlMKeHYILOTap8gUOEsOpPFvyhD
XtYxeTvmVXDuupPjk9F2d5EG8jMCsMKy6X4uvWs/SKos1k/53WPo1qesdrtDdAqdaH7NY19JAjIQ
pY3dsxLYI6r0zEen2NKD5y6mS6pyDl5z8BlgV9jVXMkjn7zDtrsS20b6+2KKnkCvbXy7L34yEjK3
g/y8cfdqOV/3a4N2HEn+vfEyH+77hYkx4fTx//yZGpGdXIZT1WtehlpB9i9F3M89vjtLDJnaMPS1
THzW8LvR5H5Mc0vBjbHu91f5SQvQGMhd+jesBGpTdmpopgbTHTj5sX4Q9eMJc6nHTu1kWw1nRHgD
Cu5doRwjalDpO9i6z/H2VALbAz+Sr8r7s036lpXCF9uR6S0nipex2ns0bQqE+Rcz5FKxO1eHajrN
GV4EHI/vAWvNgVl2spEw0/AIRnF8m76qR52EPEx5vEpNqJ0kEotexujP0TQOUlIrg+s1Vkll8gnv
Jc27DaDcgNy9Yvcf2qXZZpRAvE0+TJceBf1bhEfY9LsBD8m96HZqdxAQKx2TCojL2t1Lt5srvQ51
zUhTOpLPQjSNRsZLIWDxvrwmRo+0FprIFW7LieuwjopYqnQruTTk+ljnXHyKVtFvNCsESurR1SD7
ikiFcnUcbGmxAQV7ceBneQCaRDRMKmpO/yJXBnztQFNrQnzEBnpqJE9i2/ipkL5rBnRhVj1zBQiR
iRuwavoUqrbSbmY0CoDnfBU6+6OG634htioMz+bwzh+uTCboOQo3tJ2+Z9f6m40bREqsaH2UpcnY
9JP7eKIvNGatsEXe283fNoaBFyWHlVKx85fvnz1ANi0A2WtwhoFGCWOYR3JICUocsWoAV2KQrgU0
x3xwIyZgm+1SdZFPuGw4Dt8tLNvpG+r1L0OS3Ew4VGB3MLEKoG1gQNc9Td6VLsqaGnEVb5XUoIWE
6KgL5StQzbtsCG2qw6SDZ9t6kWiN609bFnUy4alicaPMjlHDfBCPubp9pij//u6FfncNDD6uduSU
Z5vorTfXZRjGN4T8pbIyM1Pv6hkfFjEQs8JHXHg6XrcwWP3/ja/3t2HILpFO8GVstVqeXfgsPl1R
yE1VscCct8wE8HTZDaDL+Oy/fyYmtKO2UgQYKmkarFUG3GeiPDYpTo7su9PGMlv45Tgww+VViozP
22Tdu7NscJmKra6rtjzKpkesFIIFwFaQ8vSxIntNkQqd2lt0MmWaWD6aC2XKPRZ6Qxo6ojKhdr8q
WRcNeSgzBu/5BjC8CAWSSfiYUVP8OFwujWeYXCBU4kWUH5BCtBNDhFJ85WqES6bBTRcnq+X+23M3
HYmiDLWTNs8+M6MbpgjYY/6S3cNsE4+UOESN38k5W+hSj3wcVi5V5/3iC+DIWxiqKjFu3J76JVFk
JVcWMt9z1vv3twUJ+tDzj6R+6gw2dTsvBJVabgMjbpHiqtMLISCX3Wuz7aa3hDcScdDx6pp7pjUp
55CpnTj8VkcN8WQnhdtges0V0V5Oz76ODpGoA1vo3Ad1gv9GR/ou76F9UGIxpvoSkgDZoDrH46fZ
Q3/9nZjm40n4Of8F8QEHbFq1WD3RvWnM0/tkvQ4TRRUHhU6n7DytXjT1ZpyT6yHxwu9hEPntcFa7
GTP6kgV4Zrudz3MkaQDnOQByJyLkrqJmK8RH/05rPgMHeS5GnJarBhqRzpTSMNzQusEDF9dm5YKY
ji0yGXNAm52yIUY+X0zOK/HNplBYDRU7oi/7mLbzNgLoz1uPDDXHaYayl+5xxqszrgSXb7NM2698
q30LgLjAGHWWu24u/mC/ukgh3UnyL+Kjk6dleQAst0GZTfL/SmO/UZ/wl57v5ZVmpk0vFXFAAOcX
T/2o3AP8ZV/SlQWkkE24vf7eQaN1g1Ak6XMRExXiF1O2f+PMfj0sb5OaTe3w6lKPfEDfm97uEFWP
Y9tePtV8SBsqefMd6d34GlgP1aXeg0SeAjHRzOxidibglAeiVL0iQEq3rGuWI4vmjiJD0ahLV0DK
14u9ov30fz1n3ZtrRFcI1vD1H0BrZWTdy61eVZzvURnwQkT4mP5UHUvGnhmMlJQW3KNL6ZtYxwF3
bQPIc4ACXBdYHZwWgXfFHvKLkq4AxGAwKKsik0XimbXKwedfH10TQYacwlMnJj3W4TK7KyZElg/4
OwKISnnIkgYBO1O3fNcp7oKXaJW42csfN5d44Sp9OTRcG84h/UhyNqBLIY7Mo6qGM7y+Z9MquFC8
/J5iqZIG4W2XVBoJ4ug70oVI3ftJs+KQkJm9IkYRFuEq24Q+RX+apr64jZfL6nMcR+g2zlbFz+Eq
kmGeP9XI7PBIVm38yDNK1mAumojPGEPWHtft6ijjySUCKG6JG1hRbLHLAmdSqIAxaFkWnDOq22NP
X/2h37cBiwU8qFl27Vu4IQHai40wedihGw7ATqjrtNm+Qf6wB0sLuW+7Y5pQAQ9Fqnr3bbtkGhm5
HuiL3D5JBkm1oPIvm+Yegmd8B604OKIN5Z/81d7sohZ2SwS0FaW1YFHf9W4Hu8pa0H+r16qfOiGA
NrtSlw1vpagrYBhfpMXrzWGFvhX6UsPcQ51Gwmds068Ujl7+Ud9nfCxK3Bao2rX/bYx6C98TT/eJ
1OOlzEaxLoB0l1cej4M41jG5YDnt8JBrjMbO19QtM2JA2ruinQY3EnHrum0wf2QPt6JC9APXMXD1
QmfhXsflCEA1M/xIJTaS63SjwDfQOuAF3t2MoOgDCV5MU7+aPgMTscVx2qZlNcvEYVw6enP1M8ve
EpvJuTNRovAvEP/XSUsM9zL/+F/teJJMBOVCwKP71CJ0o7IzhhZIL/25rHPsDFY8AXXT8BgTpz8o
lfvMr30TQmtVJLOfzhh++neC3Ga24j1Lqu5BrAKrAu+/V9xVDftAMUYyokHJWo+QPFSltRpkCJSo
bHa/sTOyHha6QH7tc1BAARng/1Dof1AqubPokSTM/B4wNtOq9bQoS9ae+rmIasvdGaWzgQE/PEGC
3KQKO5oVqsO7ftbDiIMgA2WNcMn5v3wAXRj6cc+939WFsKof49pRfdb9qMbzX+wQpW0LdhDCl6rI
MOojR1ui9bzWG+sCXAxXwxZBDKMGmj7Fn8WssGRwvx4rxf884MECYmx6wBsp9XNZlrQkAR0G54pX
QYTWWVyS2CM9GROfSVrN2sgjM79ke3sOW8ExYjakePMOF6/8IbAvfUlFZ36uTmvvmfI6EuJmA70e
K62b+vSSWvBnkq9CXst49QA1Mg2P4lqRb5Oh0eKZqfPV3Pm1wCN4pdqfuN6M2nRdvpMq5YSJZVJi
gPwKsH0KakqaPQzexdtrihyf8kVTaOS6hsA81sDrDa4eV4fTsFOXrniDgG81hTC2gxp4f46KtF9I
K8JumRycP4zyZ3bHECEA6g5yUyQPASXulQN+5L48VNVCfV+nEA2aN1CxWv5KQFhGUrKzUZidpyg/
2DOWieGJAk2q8fx1lh8Jwb6MKSW3WR7IJ+xCjDZYAjyze6awIFMzlVcSgOdzvqJu2eBN+R8So1cB
mYgVvmWmese0Fs30cJHmAH2N8cbdQAOAnV3oD6Xs+w1yb3CME/QVF9XRCNSvhhm4Ptx+9JJ6ApWL
rBndE6DLi6eSPXyYtx9u36WbW/XhMMAB7oU+kTGh7rF+NnVBjs1FU6x0wjBKK+xggv3SH99Ao5fg
gEjcyVjZc6r3ZFsBLWFXZVtmnS4ZcMBsz2BJ2B8o7cGQz9ZPvLdaDUen4hICmmHhf7Kabol3nhR+
XKmnKIBCWZRTjoVaQoGZDh+VpJbi7ZY/9K/M+LB7zDT3RJ0AEIY4H5v/YMYSSzLEfNawH2nbYeJg
lyOR14Bp1+PjHc9kmGexlt//ppetlnO0pW9ClVLqtinqgq3JZdkGfDzC/Rj3yrgEvD6w0co6zOb0
ryf1MedRqHZtmKMxCt3wdMYF1/Zw1zPXkTJv+ywNlhFvIOGYDg4Zj1ZE/39JSZ5D44vNs2cpjvvQ
iCIVOU5Jq9v6ZnWIhfIgzmSmBPulYAwuCgs4T0gUxXMud3HEVMqT+xYrecUPHXU0xMRtgjqoYhkf
aoJbUKk8R8yE6pjAp/pFus31Xx1mEGi4Q+hlXrgy4OCtL0uENrRvM0aA3hXr080JFK4N8WbfPwzc
Io/BsC+iGylfg+wwl/S9PQqUMTEsLlmgmspHKbHaPmf+HKqfkdmTRjWpZQUkDdWiN8bWuPGsS89d
+lnv+nbUwaoEtUHgNlm8ozYOr8h4+5F6MxpZ0Fwxe7jPf1saOByqVjeY6JukWaGpf5RVxGHqF5pV
PuLzUoXbHYV39rf86WE97nVwzmQq0c6kVAuYifsR155BbuvBUluHo67ce0YK+uXBefqafNCVgr4Q
RYC/cyeFUXCAWUnU5wgNFpnUmu5pYzXTnXXBmDglS1Ktw7CQvjFEpv0rY7uDFAMhpbu0gMgtQCZo
iUaxuw2oEIc2bdXopRDDkxaXaqV4LpN/RDCmv9OIa/iURgR5fOMwZuQVc6zztd4rDJqzn/Tof1BP
xlYowk22Q23LzCB76EidHKTeivzMOcNvyxYroijymL9fz0m9yKHQC4ewO8sYk+jrh5M+OSk+Qkpr
SldvaE3u8AoJNLbWtp0FGjH/wUhc+VdhXMSheYdYQHE3/Wh6OI8vjTsP2ZfbfdxM0h6AX369Mvbg
XLQf4XE3tSXA4KKZvZeV/PXm4xvswRGL2Iz7DZFnwx1FV1rla3OpNT5nCrrGDVGeH6U1bXgltxnV
Mz2Vwe2yoJ4xx5dntpBej205cepPA94gG4znZUPyWtmWdRbanCxmO9GiNh6s3+dNk72yVUrH0fZA
/2m/pNqcH1yaBwnH2smnYa9l9MVE0spVxed7VkDrSP9WmTinUGZXQXm8mXM051oC5qvD1lZogES9
fdZb95d/bkG+dSUOwTM6JSprBb0xtZAgzBWeSRC5SI4AvL1/02rkPDo7MshfttuJAMW8MteEsq+o
G1GRPgo4pssE2pVLGgB1RMAI4M/J4gZUhrJPYxtD2dt+6VYkQ1r8KuLQSqLsmczqEjOZGk8r4UD1
lhlKv74S9PjtdtO8In1RpCQUwL2QIrh+UKwbx5NQRQtLEgkU10RggEhO+ti5sr+Gw3hZpDR2Mv5D
8TbolUbJvuVnXFpbeqRITsaBhPzJAi8gXPoo+W3PzqGR9DSnYS1eUY6waKpTqJVxAs7WvIsBqahY
hALkvbUPvTLp1xH5Wy6QjP1+xu6KBtPUNzN4mK9IpNngcWPiQimBnP8xsycaA1PqvfRFjiLIhzNL
2AylBri/YZS2zVeWxPvATtFpxh0Dzb+MwtW2BUa+WukBaqOtkLW0+aw3J1UCXbziIo0QsFZleS59
qcPf8pX3emdTkhnqJQI1BudajDdIR5blKVsmQpavzJdJVjRk0iZ75DlFKtbeB0gS1kjj35Lf3wEP
wTZmsr/eQFixcHTLzaLQ4lQVK3bO8NZftdg6bnYrC0Spuggby78MZakqXDYub250PWxp8fvEIOTS
HWPLjGuIw3XNl9m0JjdbH0aCfthDm1H9KvMP5Aohm07BmaQWYMkSCQFZW7xRbM7SHbUz4EHEqgAy
+ssr4AKyYHwQs/QlHkS3TSF0OISdkEwghrvrdFCuhpmOhksPgQLa13BJK10d4I+xZw/J4Kfa/BC5
kOv6/uwoQ/iwfUzlQth9wOFk4aE3VO/KrGz+NHmxmzhhR0IU9WxQxzXQmj9x7I9hO2YoCQnoZbxv
WDMoalLYZ/yeuZYGRSwp8aKtntGu6guabMhI+pLqOAU1NfnqZpLO30SiDX4ZnqisxcMA0mlv1vxy
9sLAcfBTvPi9vWDHXntkQgvPNi8teHuo8zMHy5/UcsdadfBlnoa80ZcbTILorzfurDj9DfwQJd2u
NrM0yYSczSr3hPOOMvi38JGCdhIiHXWQpByrt7o9lEUkJMDsipS5aQpdOLTMFW3JZ6DVkTQ367wS
zT7c9/02L8g+FhNcCH7D2YaA00dM3eNQqCIWe/5cp2UAl/XBxl2yMocyMkVLOGm22y+AoOedNZmj
Rz6ec1lmKkcEbxcMdKES9qZ4b5s3WciyzeOcFB+YzgMKka3P+L3Pta/okRh2UneIS46Wz0OBXlKr
IZq9GXtMRXtXEpX9m6S2PyTwegeM6tlj+t2hBsbfAXIRRI/H0NH620O1KAwb8MgoUSSmbPU/mlje
XZwXSP9XZmtuBf0TIXUl4mQIgxNDRc/xR2mWVNwhMLhnLMc26V4FUqFcAn4YWbePcmo2Go/ucum3
mn7JJPWuGYTgsdDNf9XU3n3ceMurQ5aVuQOWGe0KeXwVY9cH/bt8KoQD8OTXEkgH8mDbjF8ivnjN
lcglAnH+10szfVw3gwkiA6kAQvhj20L+t9M1tXjTcruuRQTy5hbZvn51D+NWQeNlwHBqTCAdJ11O
HhEIPSC4V7/1grQWYgqavpgWbfh1n4iX0EYd4c7x1fIi6w603R85wNNvv/4qMgAbJ9CRMtXADjS3
/dbwnraJXv1vUTZP5/GCjlD/RZLeM0KZ35h9Bv1m75HDqLa9hdXcBrHc95XOlEGJVEbJh6cjjIDt
2xYYS1pobg1/w/W8DVTI4Hgbm2JUhuhto+Z68AmbaTFI4m4wdJ1sKfvXiuAuoHEOhj5OZ9M52ynl
/2hvDL60AsxjqxC6ehVS6Rb3I2NEVEql9D5JvkvuAGVzxm3Z9ekKgg4qgJv/Zm50ihQI6albWvEW
a3Lm+syFsCAo/twGjkLc74q7Lwstna4tanWrFSSMyvN+69zmIjAFfCYoJ6c5wtPkiUtYo2QYw5Z5
AVX9MusM8bTvq9q9qEMITxwqsf0PUYOrJGC31pGd4czfOurc6ZIpqC4nbZWvLQsmVF4AAAdQFELT
j86r17GIT9rC5t/GvMRWfk5geKSQcsrTgqc5HPFeTsqNIRqzLy9E0Qiu2g1SXypIdktdZ5Fx44xe
PN3ZqTi2ojGo2IThw8kz3Ynq9t7gNyzAJkotN3tAbHLhIZC/WGnR69GqNnEIHlZbK14rEi8/cY2w
rpCcD9m3vpDAbXLM5zOlpvG36agTDJfZQTs0V2r/NQg3k93ziv/xFUqAHUX5P/NtgwhscqycUGTl
fu1WFpPG5gjCtksxxpfy0FwKh207+e00jdgTP7q9iZXLZP/E5pLjccf8ztge2As4PCUsk9ngpqyF
bL8VuNj2MrgYh8Cay/d7qi5e8QchXpHa9pgrStiOTV5faqCxfL+GOZOmBJ67244Co6I1gKuCwSrX
HrKN5yQGIqLb9w8G6dFeHCfXpWnR/pvHXEKONjHNvCJPHsqsfhDtQhImc8PP7jt+TjA7JOQCeQ7k
EZiu67ibDzmioOl4FQfk440sKK4uZwhNvlC0t2Tu1yGQoWLea1LA9K7ygLnIcEFHxzZ26/1DLb5W
qtBKE1ruwz0vxMIPeb4nUKBWwpEk6m4fcsXCqznpTeYd+ZaXTI3EFfh5MLdHBko69Wk7JoSpEE28
MIKtB3XI7PguZZv7aRSoBlxvgZwbOvpc3SbazUs6KtvCksx44d9ZuXq04R4yZA04rVNJ6tdMKQu1
GezRy67rUUDrf1E0aJirt2r5uMdSxhtE/pOKSmolnO4RTcM+M0JL+BKqwVI2yrs65yfYuQQVhhpC
02Ap35y6nUBfHwINzh4/+gX4n4ezugb/b0MSPCo0GUZTnQfiFmQ3ymQKu2aw3VMKAJ+C/IDWQJzT
hRSvX0AI1OMiJolm2l389yHbf7sDGXH3el7L7Vfsrh2i1C+4rV6rSpfVMP1m/cnftRqkd3w3HD+S
5/H8UDNBThvKSrGto9YwtleUq3muD0YRrVwzsXJC5mCvmDLcCHBcQ1xwSL61ZQWCrU7eiy6T0MnD
8F/vCznq5pOxohUb/TYqUK8J2mVCRQN6/ciyW7DS+kLdlKR/EK0tXZUL+3YgQVENYngoGvilUSiw
R9LEEUme/1OoK7XbyV+WrodnZPJjm7uWix6waYNVpd0IuAHdLIY/AXEn8JYGiF+s6OSalimiNtdA
X5OGgG3ky55OHgD928PbUBD4xWNonvHDXkiDFgLax2bs5R+i13HtrZCoRMq4k9nDj84yQ8eTOFXm
aY6XrLp7siUmKEV1PnqFRuF/gn8cq2OHI9GBvXM84nMfZvTFlgmXNKWHaipjO9dZcA2z4BScQW4Z
jpRig6gdfgpfcESp5dRtU5v5Pm2qQs3/T3oR6ZpacPCed3+6fdSDtZwAVA3n7enqjhiVUcODAgbM
JhV2HKLzGa/n2p3Dq9UbE/U45izr3xoo0MN3HXOSztaKrHr0k5ZxM8EubyDB3pe81qh2YQ3syZHQ
/MtQAtacG6uCKQ/M2x/75v0dwe1m5LoA0EJl1G9O8rx6xdyduDOF9moccyE7P4kgbPDcC+oQM02G
wxDteTXNa8nj/jFWrlTA4WILkY3s0+1rNJkm2JaKnawnR2wvXDF0KsXLEKajfHP2lEbi2AaEX3Kv
DuJgls6NIa5NLIYayxtCS0MKzgTgPf/UvasR7+E7Se9R2IcfInP7ZRe7JLbURuYmR36agFTFzaL/
4dj/G7Ea7mBe8Ypm582xk3hNSL1HcSdRw4mM+kh7mjeynXX2JwOJxBOqSt4z6xDCC0dmZYZ0BFAW
+vw024qulOOsQ39rb+hFqVDnWNHTZs9v11gpMP3aGtJFyncZaMq+6VpQK9v+F5Y5sZr1TiYwSsNZ
3LLNkP2FH3MqL67IrO4EZTMODPlH15byOMZAO/S4q7idxU0iZ5c4lvEmWSb4qVDpC/sCVykb60IU
f32mS1M7dsBEf8xjYbKhuWTj38TMoIAQ6hT8v824p19BoDqT3Mo6nQLShOAR/FJ0ImcIRONjwjyJ
0VZCYf96iuOBQS0F7sA+XgzFjwhtaocNIeGDQfNRbq+MxvbYXFg8H6a6BybjEGVVYOpYpZjhQpq1
abDm4Kq5RT/jnVaXfKeFsQcP7q9FdzB3/sxctFpL72jPSO/ssTAlAgP4WdycnMrE1UbNVC7ZqaxE
eodJvqeS9JIV/EA7aYIL6AbkMvx/sG2seKVR7NMuuk+vhtBP3hbwiIq7Pieup+sRXrMFhPDzSjGB
90o4JF+rRtZfmIZCjYgBBDAKOmQg+v8BMFqp/gIQtfNVM076/FDG74gY3uIsLL9WZEGIqjklSnd7
lx9AD8xOOlP9yRq8tTttxgf8RlD6NtzksXZnUKAqCcSJ8Uq6YgsejJnOIxQ9jhwJr0G3jLOhe/u9
wx19fzIVqYn0vfHFqVkIfxzedgeKjrpJqAE1yI3cNMN4S1yBCRdy5wS6kAhOxV9ec49gTLXjzwGZ
5op8WeTXFBuLGaIitJKArHDqdpPDJx2xL2krTUtUCPrn1PZUrfCv2Pq7t6xdrQIwUkepTwplUwWQ
n54sXpcAAL6dXNd9MFo3J3QpmbswwCGP6bJtBJn1G0hPOTiZli+4HPlRaJj9bz06XftJ5pkuFr0A
zmeyFb2FsBImY5tIZRPav7bJ1hcxag/HZklaJteYnAosYijjVKtsV5a5RiT4kDgX6mdQxw78pb0k
mHMn7mhLQ/Izh3OZhHX9j1LY6u1eu1u0LDfReH4/+m5WthLHKgJGRA49SDrFUYZlRpLOvaz2lN62
B/QMYVXwv9wFnR3hSxvNENr6LGOCYzZJ1PXpbX0tsT5MW8X2X3ILWEuf/lllxdRAtp7agQKPv9gM
/HIHlIR7AwLOHK1ccissojrzLMPBWS+BVRcE0Z6xYHaT5Elv8abVNtUpA7UU6afJ1Ct0L6RCYs5L
JGAbiBm3UWxKDKQURtUqvyRlmBuycLwUeajMTud3T2aq3AJty4DtajqPtDfCPpKUrf4YQ/W7HvZI
HhGMb0mTcSD/KyZQE6SsEylFnur+QjEb1mXSxGJp7UZrXNqzbr21QCsRvS5gseA0feZNoZyi1aaz
v2iPHgyC0+K2SB2bQFxrSs/h2pqO9uAM03BcbHfmobOEGO4yc5me7xtGdzRT5NJb6yf4H3OmgLas
fxIrm9FxBf3UBjJz9vnk8/4kL7vzQovTSAXb9ntkCCmUnE7Z8AWb0ZS5CPGAVm8JU/dvQUbMSzKl
uF29Br8TbgjskIQXqwnPTg2H1KoYvBA+2c+jvZpoXc7a9umYeAGrkUPhtxKqTIIij+gyJN5jQere
GNG6womaUiIC/Usg73YS3tVAxGC6P7nO2VV9bJFrGVLjZvZI+Ub+3fljv8jzMBO9DcSQAn1ku8at
Bdf4X21uKgF2MZiJmV1FyhV6N7JNuKm2DbGmjGBZzJTl9iaSmudXETw0gtCO/IqLVf2HaG+0wHkG
O1+xh/NBZ1T0lkYAP5aNaxpBr6hPoLoHFSaZ9lUwO7o97tJXnUtFem0ni/L8FHD2bZhWEMx5gv/T
TMhlx2IscNbe6t7rWsDHCTvkhlS0+y0E7Mld9YIeFC+V+DX3z+LyDhuwcMYCZ/Tn2i/EVIDd4BlS
PVfsc+tI6WHtngGGcFgIeV+MVPQ54fXOS9d/W5Q736pdygp2Cdg153HwSNBHf2D4LZZpS49LlwiJ
gVPKrnDhu+3aS3LEyts/4JA8r80FlJhwF+xrrMnX7FsQ+PW/CwCm5Jypz4zqPB6OhfBuxlCRtcXb
UCoGd74pfHxq9FPAhx54+TsuhA+oiLAwb8uUj0w4b+ZMcryQc5lBtH40LDM1alcIv/iMN1f2TsTf
jX/7O0Bn+vlMc3fIIb5mtPBpHBtyyrAJkR7OW+PRuA5wJyM5Bsa6lzfbVos2pGLuDKKJQbyUNQ/U
6b/tKArPyx9LeiPG/WHMIpAWElnqZ3eTvAsRtsEVKfN49tkvT78NfBZvKZG7VFa2zQpN0yFLX6mU
dc3PJLtW2X2mLzCl4hdAgH18OdTJb7vCZvCD9PiFcToVvou5ts0XLnm+sNb1nu4sXoeGeDuZo+58
hbgZd2/k6oIyG3qiop/DaokvPWK5Lv3Y+v3i9mT1GJkJQII5LEMg4Ky7jY1bAJv+5S5DzlcWo/Do
5r0u52ou1RpkDTIUXwjTn0gpnjPuHSyZnlalgeu7tM/ZvgCIrAROzPyvlnEWVeS4mjGFHMM/zGZ/
u8RMDVPS5SQYZPwfK8zuErkxvueMAd/AquB2+LaZNa3vLQZ6ipaN5M+rYQu7yV3AIK69StAf9jDF
9MUTiyGvgowJWQHHJ25W0GTFHSWBFsSS0b6ZcY/+q1PUNExcKrXsEk3ET3aeby9dOfj1AnBI5LEi
yCX137dbFRe7gd2uGfvJ82m2p8c/JcYzQhABEI/gT0X2z11o61HKJBNdIeLunPHfrPwrteKozJS/
0kOnjpHCh5DmoHUzzZhV6JGKV7daqMkCrKtxxh/5oG/nSld45kFLiOj7cgV4DU2w1F+VnlxyiakK
Y1a0cTVX8EXEkKL3UWAMJIvUe379y4rhgPWeuUCbJ+YaaRSaw+M5dmUF+wnNPG6/UjOSUY3G6t/f
uzKWhaOM78ztGKHvEV1PsjcW1dUaY+ITdaNrfYJbiIqsG61GkJ9ahpscIicRdrbY4R5+VbDs5SfM
BLURhpdEtnhy3gLG2wPVmyBpa4Ovu1i4iYbMh7udSAeUP6znemlGHUsFjS7YtMSRBduwpe1kEzNS
jWhExXvwVnAmN0bWoQqRazCO8bd4iSWpfg+oQ9m3hXe7DDcUcqjDjjJM15o2Abg7MXpl3K4fBlwq
zfDSa7BXDMLbSPKgV0Vh7p/Eu29aVUE4/ZYEzxRNUNvL2NDLTh6exyW5cN26OZvI1gj8eZcWfgjM
c0EyrpLe4qZtkR3Srzoqso1bSWAA4X1NAbH0VgSZfzwaViwBzL4spp1NF1sGAeYf1LUwQlqyr7gx
vpJw8v7+8X8rE1EYv6Y2OukNXX3D/FnP3OpbPISZ4BL5VM/JKfFpqSQAHKHYHgjIDLDrUNInwcy2
FWpRcSsk8RIlsfySmbnbQ8inbX5B7MmNNcQIVhzOBACuTq8k0R2KNHVsBRX0brt0ZhSc9gkQJ6hR
uvksTZ7QIaYI+eajciSNiHzQIIcoa0VtXxLHYZRE5zGKWHufJwIMnkY9eti70lktzqx74Vv3MYVt
49gdSbcg40SihPegseLxDLMolSOBQ7BEN8E34S92pcVFGhGvnswxFIb3PeL22asjt3P9Q5yVb44u
pT5fFj7GkDchIWpTc0ttJDTlpECENaSLgik3mfGp/vdFu0cAXa5AYckN+gSPJyK1yVq2rWRnPxRS
+IYh/N6rwdlbYUY5Z0Z0NdqKl22Syl8fIM8wc6Vj1cQJqD9sa2Aii1OIpYoTKm9uaL78qV7aUMvD
DeibMIaXsUgJSSpfmuvRVT/WPE50u70ZE8pO1VhLTNIxgoEm1XaUF+eVgxQaDyrfGQ169x5YE5Oy
gfP4/WkIN0smgQCMU9PAXQENzPgye5B7xSh++eSR2ms7QX83En2YKQrKRGc4yrsihnsnpZEllR7C
h0iaqOemLKDSmzpqfkht9yLrU5DT2Ip8LbJLX87yUG8FO9vaGJsd+D2kTmOMJrs4bGhuub3rFqQf
e6s0zsTQmdSVOvgKLNevzDZid0/wpojEbhye6YL+fxwYAVU0qxjWAZgReRTh1mfRH3uz696hgMiw
Cg7WDeHjbFPw20xMqswxVuVeZ/M6gq2KmJHGEQXV71YMG4ef8HMXVWLn9hXDYVnTsKZbQU21bZDo
x6Hpq9z7or7gYYdqc0ZwPyQIglOYftCfkQO4EV6v+w6F9JAu6ClDeF4BdOXNkmABsmem7HNRyPIh
75apUAAO4ptAJGCB6UoMLary/Bnb7LihvzaZ5Knbo5YyHto0ek/mQkHV9Ib0FPYgBfO4mNj81fMb
c57kUdOktKTYRjgzA2+iL5npCxVdVjBY9Lp0EIfVOfI+13QGFcnr30IVnQ8YhrMyNzemcry3X0ys
YtFPY9Yt5KFap82u4Ubcc+jAhPeSBZSDhqSX6ngf38B3tbIYkvd1R2cZ81x4Tq999z3ccivQ12Zq
+2rxnzecbzuiBJng1uyMJBBpzhxR2iZwhR6FwVdihwYSnWd6CsE3aszSTqCGvqTiAELTg1Gos/0G
xoEPmJp0VCE0hqhMrZ8715XDRpq13UCYxllz2kYGJr7K0yBjOF+i9HHM3W2ou9mKZ8xEG1n/TNXZ
ScXIMZ+uBmm57+XhMpfL4pz7qej8RpUo1ev0pssZ0FC3pFbVcbrYh0m4dXBMFQSPL8AZAENFN7+i
cEU77UrejmX/5aL/RZq5ms6ecscd2T/Urs3GuZROr1b0Lj0tPsCe9BdmFzDjUqhE8gZU66+GXrpL
sNZ+9kxDxn+G965JPZETOfGvUgRK1zvljEihO0bZ2yEuRXznTB0ko3ByIBoPD10FMYpzx35TccIr
3GoljkYEADaN7dv0AXQen0zpjH52Pa9EZxJHqFahjxZ6C2gcxTCFU0DXUEBriw5oCtsAqkg+zMJy
avwtEJgB4oe6/VPqxKgkEZ4QGO46Bg4/7ijDYOMLAAwHtLQn+a0xnfXvz15d+VS+H9MuZ/5NoRTS
9z0bS3QkzTdKCRYQwJQkFEfPFHUvNtqSfHw8EN4lrMOXq/IyvfhYg2rM+TrKGRpTuQh4dgwzB5OT
T4eJcNvJhgAY16f5Pwods9IuovG/zItqM5FnUr2GiWRzBKl8+ETadED8l8kY02XUViMiWEsAqEu2
16M6+qNBckTCQy6icU5CYm1q4gE3U7ERIZMhL7AX2Bgig9SyuDWnm2mRiq66VKGIwYJGQsf22MiY
K7QSPYHHWNfmfWJEiWdhKLIOYoCGEwZ3SN3CepVIwjNFCNcwGFgJrLZSp7N3rSMLpaN8OCzJfddW
DehvIdwY2Yxk/Vg8UZ80qmnlcMmi0HyQq7uOknT9Q+5WJpgvOu3VcorumXXVLOPR+uAYnmsTLjy+
o8f5VbDNyADyyOtrLWcXchVIRh7hrao+UdWrEeN33CQnBxW/E+RddxkjcwERKQaClVkiD6a3fVKF
RZGADkO5pJTPhWw5cZhnHBLUC8loYPwDvYP1Zql5a1t1MiJ/rJdbBmEWwuioHOYiclm+bwodgw1C
iJbWrSRstmFiW1NP2Ceit1kJg4DuFOxG+kigWAm8LaZOCZ6ToYOcsQSKpZr5HugZZuN/WN7p1Pzf
5I7iu9Yavown22VwhrLsyQE1jfuWbPXKGCqJu/kY/6G4dpzw/2PSsHISfjI294VRMdCavga85QyK
39FnZRLz4o8+Aa3yvvRHe4QMtbGgAzALqmOEB5q/i4yrrmwl7JKLWn2H1e5LqjYMcu325HaL8Ru+
BwMSZCKrsKNPyYlSar9p1iuL87ers4Qg6QXiPlw0tWHIjbSowfQF6J1Lnhqae43BE7o3hwMu8f5W
RUS78NbfdpMYrZODSpRvhk62tLEQmJcW5CcRZ1JXoZSd4jEnVfPHvlubHxdBnHYuIgxlQbk4GnTG
ckWAgYdu0BMM1sGDoDzUmBVnpEiMatm21otOx4yaA6NorhbmUWSd7PZFBUmoXPhMt6GfO+LKwdki
ZHS+NHaunIqjl0uCtdv2yFkuAohnEAMJazhPsL9uRveeVD03pv8P5sWFMT7JFhs5SAyo6I2j1DLz
/6xOmEpWUvv4kL1Y/2xn2kdoR9VarowidRkVXPPtU32ImTKRVVGhtVUulw4tVa3pBI/40tshfuRJ
gko7puZ286gZWej/T1jHzBRazgg1pjPbXLp96H0ED5u+o9L4UCZTSobq/34Oz5/ObGkHWeAXSd3X
kuGhSgjOTIKTS3ROFRrRCK7+CEpHL0mYpAOGWdoSVJL+z3/7T5SBWzoC2BVu9FFbXipeuxL2+qHn
Jjbk/RM3HAM8cn+nSxT0xrbFw9p/7T4v6tu5K8fU7s50HXWL1aiiwNpl1GUUkLKVWTxWmk0Sq+QT
T6GZe6xa9S+MQ33cECZDU+U4dZVLDUsIa677idGXPL4PmFRW4kvjgqaW0VBPcNJfvQkMSJWcTEI5
xqmw3bJ//9s5Lc4QFsylzATdeqgm1pB06TGQm4qFNyLONQX5Il9S88JvDZZdQCAFMBun8xsIDeIM
6g1Q8AzayHrckJRHz57DrXVM9zLb3UMEZQxmfbMrsNmuuJvIScDmcgk0/rdtBsbgzequZYVjzQHE
We7L9y/vJ4DNXM62GvGAftr2R39OPpUJ/UwVZpgLzFE3ht01s1g0iyTAHccgGuaJb1GZCMk1CAUe
oCUlwvy0Aw4tGYa5bHJOZH79ErsUlg+Dd9ODzard8IGH2xD6deQAFLvyF1lOC3LDEiEgXySg0DZM
ps541Om21NnMbzq8OHu3HEpyDdJTIoeoyymIsUgu+4uzp5W+zF+zeS469s5gZ3AYjyWsaROrvxyH
PRNReAT8IsjQNhcKrN4BuCsNJViE6xrmn0HVOdKBKkVj1CGCPilzEHarvNLOFOcXuCZdsbBcOxuI
TLUgD2yuVqUmx91518TN5cymZFsZCar/11sOh5ToT+tLu4K3XEIeaiOfvZkT5EuVXPcuHS+YRZVV
v2umf9KP+NY7Who/QHKkK0oc3km+fgB5ED0GuQTEoTbRK6GTMr95n9UCsFsVkVK/f8wiQQiiGI8i
04qynsrCFDtRHHn086B1iqTg0TXALmrCcNtgFthVudXv2WKxb4lH8V6SsCSsMRQ3m2VSDmxKHivE
TP0S+AViqY6awdVS7nkfgeCQ+V1BdfJGo5vZ8f6XDC3ehjakgiWDI2vckJodJ/XNC7J96xX00Yoj
rYqplxHi1TtxAoYOpiMICQ834FGAdf8fQq9LJNyTzl6vHaOGMjah2iMeiWQiGCqqo9Dv80xO13Qv
bEwHzXggsNj2Byr9TRqRbaa1EuIpU7IuB2Ys7SW3Zf4k9Fo6HczxBSUZ2Nz6TLVHcgtey3FBrpFu
3RBdDDh5BFSRNYNqsVieuDJal7bqowjAkviQk6Zvs1JZhJyN8Xa91/82KvK17t8/QjLPm9mw2cpC
LENZV6VLDgE2TWA46eB9OodZiJf9aV0yxrtmuJyV8oZom7MzqIBU9ixBQPNtt54AoxfIadX5lDVZ
t41jWS5LvWnw5iXSYuYCzz2pI/LQPRFMJKKGFQy9Xh+8iqUlo20XFM79Bm7FIW0pPupNF9v+1N9v
1ZCGsDVfkqCSI+BFpHQc9Pvrl4OmZHWDCmfvFwsgz1tCGyQOnOsv99FIl69YouPwX19QacqbiY5r
p7U4vmZyWuF93OmBy1PbH9WBFvidQtyyaUMWbzChvwuXH5cY+Lrec0cjHPVqUt8SrdZMbuPzbwMb
jejN1h1VacxRx/kP1E6/dfmWGPaGTcbYmpZyV9DoKhDffMusR1itXPJ1C41ZkOahCKX7yvbUqjly
Hen8mEJtk7Oz244+s5iV92+s9brNcvPuE/qnArBBOSVE+qjriuznr0jlNaFd8FqSj8P1zz6bHPbD
DGDHDbTWl9ZVAFbZ4bcTx0lqqCbbHCKdQUEMHb4kk0oUB76vk02f/y8HfKlcglQgR+Qv3TGo5qJg
WHY/3AtWQU86a9Dldh6AlkUhXqotLL6wilWJQNZW/ptjoGBXl8J+Pu8L9oHX3Dt27G8f5bSpt43Q
ynoYu123IOylYboRmBNeQ8eoRAVdjLXLVt0eT71J5C+2MX9DLFFTk2Nnoqe62LtRNY2O3zy/aR/k
JvlUXurHWvv0eh9YbVNa8qPeCnq96HgSa+R3ntU/vjFAod8Nh4pZMcHSEzNegrO6x4hGV1ZBeRXj
uiof8ghaMnKApvA7yI5n8MlVBCPipSfbCIFfhhfDHmTKPRwkTlOqjtMzfIBZ0+Mdp58XuIfqmnCt
LZpwNDHIafcEps7f2KmSRhApPLz8huht+7ppC1JCts30BfXbhtci15/TLF1SqxvREerRZBR2J5il
u49InMlVXuYrvopFiBNUE8SPy2ltjnlpVm4MdmFzLx2njuZuZIj1r3Xk/xBSUZkEhsohokT+IasU
V5OJFroT/FR8NeEyFoz9XatemsYYaUKw1K+DLhVX4VDjnqycDgvpAV7FHN92wWPXvArvIyMiAwtb
dmkjD2O7C6cEXPkkdiN7YY7smIyS6p3hM+xBH5Am4erSZj+PJTljmpN5SinarXG39gKVKxs56gTo
VZYtDDy+mpD0S11Zje1GFAdfF2GDVpPRIIG2uf+2yFngKR241ASU/Oll/cGQkqrSe9dpV78LiZ/B
jPzh+IxheEewX75oZ/85t7RmluB8J3OGbK+pCib0MUB3DMG8ewRfjEnNlZoKcczgVoOPVrzVZN4y
h/h75cKd+YoCp/j23IQq+4k3GS0B+gnNQs0BWwxH81RPIX4XNSG5qgSf8Xjr7h0AxvBh16j6szjf
9YFDPCvmC42OxQw/s31Mw7z34wpdfyjoPO0ILlgIkjsHj1Fs3OWTbIIbWsTVnu8ibjwcRKUbirub
4qnLIvY7rYXjfQaTQTOvR1/LbAkRZL71a1zhK1pk7H7jQQCx94sFQaIVoDeI0VdCs1DcMIl0zrMa
lAq1/NHg7L1cC4tT8cZ2vpttjFEfMRkm8DD9H7BBZBrRouWYGyBdFicmTKINNQ+bBkbPKR/mSo8G
EmgRQuXi7awqYJ+UOstPsqtXn4+Va6qn0FzGsrNfe3FUNyx8l9Cm3liZGEtRKpvyrLsjJnDXmWK0
R2zIk2dTsNVVJMMBRdc74SqolEQpn9JwXnOxfAqNMSGwlh0n1MJm8+Um8Vv8oQ8/hQgShNhydIh3
hPza/ogPWfT5oNv67u7J7Ao9+DXy2kLdAJbeKO7aN8Zymn8Dx3qkSvWHM26Q8T1csKwS5pnLkrIh
FJKRTVi0I8fHIeCxhsDV/TYxH8hMf8Yi9xUgTlGg8AIREaOSCDXRnsDLVVoXk/U/VXB698Z5/dk9
S6kg9pVrHoj0pTwUhqXlbEWiuJ8siskLGwAcbIEAAVJJ7jyz7SF/GuBwDIdjJhayt9wiJNolxqlb
7kPMyx85JpJv/staaxPBW22xmKn2gcbHzxrWnteopuDiIaEer4zdlzFMy7ukAtP60GWtmFUasLXg
rRvZb9aX9nL7d5yQaBSHm/LajoyzQYvlcBi/fA1PWuOGKGHvB7fR792i+wqy9QkBcwOZK7l3MNdo
w5KRAJimioL80uspkZXPwYpl7cfL700fnaOgt2vIJ4Ynxd9L7YeSKYx6LCxlvLV5gpXU3cKe99Ov
VDScQrWItNDh0pVuVOdEBmhY4MaO7rjXnFAEqzhkTGexyT/SvVylTpDPWzukR50uPeWeaO3d4EgR
i8U1YB9B/Kc5wRUYll0oq+TdnKltnb2D6nAD87OiDe8PN3mL6Defd4VhKlRoYh4rVu/hcKq4WhOx
s4KiZMVa8AsjfdmH4EegEM6GfltszojTpyI4CkN3NHU5cvEBHTJHPUmpL/MIG3op2JEce5tzLXlt
elr4kvRJt+K2CYGn/ribPPnj0IzJvsXI2zRCxGiDyUmdGCA+L818fFn29QxEmzpyqjxiX7Bo61dK
NbKb6IHl4XAhP6mEu+WH1etWfkKqM6LZAFfVbkH8SkKFFHMcoM5ebobBsfP4VnM2DNasNHNVGP85
AvnrHA0htt0qk9dMoneb8/whojgxH4tSLv4nSjlXwCoz9lNMhWkymfmBe21hwtTZp/uEcimkl8tk
crZhTWaSjpQBo7HXFBbJmneY0KDekACFdmG+0KD2uYBt44Lz74ks55nI+K2hg9ZzMtzTnnhqnQDQ
BJa5HehDJU+Fik0dDpv+YmK/+yPZYA3ruHTRmlDiCuvsY9O/Y7/O4lFG3p4hQQdzed/de0dQKIiT
b5bCmVJakY9yJKWn2ouJpGoTcAuVnzi51FLWKh6ysCre+B6i1FNXVU461gxXTryB3amtUBeN/Y9a
a+3dOTvMBoqla2NUphphubHy2nJ6avOqK+s7UPhQkdeLq9nZZtYDOm8fphkzmeuNF3VnRyIenmGH
qPqtVlXHrjJy/pI+Ghh0YOwRqf28601XXdUL2CiS5/McnQ2uF00LhKxFpn2Jh59JqhFSiJwDluUS
PjhtW+UYCaTSt2HPdyLQe4tAAFlL8mhY9pPIURgRJ8dzIugzaGuD77By4ya/nPLuQmTgnGT2mEEE
k0yxghUWu5IJntygT1GJ84tjRdVaASzXJJbHDHdgIqYRUo0zPVV90urIWDaLG6WwqAskrIPeDnKj
Lo69nPWVwUpXTVNTTu4/QXZ1/iEUQXznOR37V+tG7oe8jZbp5ZQjycNOkOP8notzDoPX/ABDOGT8
JFCmw2AYLWW2O4ETPditvFKx1L2Zb/lkpt4RHcbP0HRIFsg8OROoORdh7kvF05rX/D1xKZqi15NR
Kt/FTvyqNwFJ8hM84zoYMvekFUK9Y5hG0QPZBs7SCk3MlbsS7HNEJhF/llrx/JT7md+jykOtFUV4
lffYCbLbBrplARkeyR2HEjIJdEeHqF1n+i/fy2QDFUYH7gLeCSnN9VmhRuPYWoUQaXy2h0A8yrbX
JsuOYOy7oYUbFAO/zgcn+JboMRi+/Xeug85FqF1rmdn1e1y9sCYitYxAEqzrKWvd9miGAiQXTaOL
QRGp3dGaBskUacGwdJIABShOh4rRr87jEO7y6j83mawGk/S1NC2rCsFkf2Sw3vnfrqqi+D8LATYo
EFdXrHhkcFdydN1Ofz2ugdjGpBX24/G76DRg0FXTqDfZ7iiVsekIgwqxcfPkfMXH9ekAuBca8A0F
nI5P48giHtaBJPCY9q5pxKCe/B8ZBgyYcBZe0ST4DWTCYw0M7SZDGnRTtEFB3xU/ox2V6w874U+T
SokLXyB4Hiu8ORmPATnWi/EN9QDtpaFII2ZiXjW6XWFgPaLWfKaLbFTWQTxBoLf2h9jCtNn+NA2Z
ASM2dADjd2xJTG5339Uwmn7Ex7hRezLBNQdE4YTSZyMooy3ALS6dQvPIZZwXcfa8fwScsA0SZm7m
R0n1XA4/jk0Gsyn7l3Vxt+LskKi+yPv6xH61XzO0ADxDHhbeGerpYjucFkeimu/mqYLa7XDL4Gna
1KbSkCvjM5iteEDAOhU0HNKY4jOywq4lGk+ynAe3XAsIm6tDkXwjSUAAcC19NYZulmuQY7FI1sgq
d89vxYR3X/h0CwCTvP9BaEbgaY85vMcQVXGBqL/daA5WVR/I/rZ5U/uiFYKz8E6fyj3B8AnstAoq
HQH1PoQZzJ4rujz7hhSyjjcr5BNKs23IC8Kf6fKgxgOiO+fY6DZayyPmzQu2mBGXeuSpLn28Jvle
YPnM3fTYO3B0lD3S/0ROFqk0miF0uPiRga7Ci89Ps8hN/EIMPzpDz87EnYOprH91bPPvGPHJXV+M
TlayDaHhOOhqIn6BQ8UYFKmRZc/628vxXwiR9qIyIBmvdlBXHkqBRuqhqUad9pUSLyAbP0gO4TFu
o7Xk/b1aYw4cOEsbHTKaevdYfHB0/Zf15qNwkaOeOaG/yGtr/mWL45FFcI4NCtMvLCh6+ZHe816v
0ukqtCK8z72Sfw2STGnYs8jZyoR3hpZLekoFmU3xDYal4Ww25GrfhQ3bmPI/8rBJB12D+1rZgrDX
hnqUqBB9jJyhdaEP/iWQxPStXjtarpf+dIFaaMCQJ3dQGyMiYINzL2G4zp9L1vsgTOSg6Hx+//iA
Oeij5qGgsOE14oqTINGQ/pVGulm0wr/Xlv7k51hwyzEtkie/OHJf9MtcsPNG5OdJ4r4g336C1+aJ
V177oXN+5VCgKjSzRDkYAwKrCpW+U1o5w8NyxrpEP6d/UARocEHOezvlyTBlOFVgfDCUphsbLIVE
LfgLzPTtcbadK+hQ65uXnUNop9gpj4GF7BHTvABhZBPcCIy4Oe/m3nlEaEBcuSV2aFQrkMGK77L6
d4PKBp5ZwzQTLteE/153W39LIL+dMV/XZoryMbHJf/Lm/vNnJOs9fvYg2+J6WdIKpbX/20pDJLlq
vPp8tnw7wUlCn4te0h/JqAkuqlEmN8uDMaCIT3Dxw7Kh5qzWyDqutR2WBOlDwLyUOrcHnXuHR/Mu
K3oprd7OxiTleh5uon830jENhHr/cyhn9MgMU+NZ4mwneeQFlFgUBHlBs5cTT6hWi849BxmrydVS
vK2xCNcU1dCf28BgxTO6T8NZl7Nopp/m3a9FEi+3cN2RM8EWGRKkmVqJHrvovwMUY80vq3Ac7wVc
FwRw8s4Wdo0xn7d4vPYMWUZD3n786DJeNGSkx7vONXuviaDQH9MQrpEpKl+PPrQLJ1F9o7mYmeM9
QYnVLA+xxCL5nrlr85LOBn9dApebSupRyLs/8XIpdXfttyXfoDY3hSSmB5goiUStMJBsy8AaqvNe
nF7spV45GO3mShvT/2b6ktcYd2dkiqV/kbXxulmfINU1YjuNjx7ci+7YCeSAeVZLHwb+/4WIxx9S
bdG95KIIo5XlccUKlVZVMD9VK7BxbzO9sKiTnYvBBJBhBDJPh/C16N9Mhgh7HU3SSE1Iu/UQMCIu
I7nsf0SQxO67SBCbHCJeau+8d8uelIObBm5SitjlNJfEyj7h0GdmbEWGwkQSpl+CDAqzt4FoSOBc
wa8sYbzkEMzzAqB7zfetGVlB1CkuGSCvfb2PRWL7Zsjohaq9JSCp81bInk1wKUPYZ/wRsWsaIId6
AtSL80vceWqlJcT/ZKDMcZJ23YIXhVnunYLYmIjKcqYIhnCvPx2ZzAQG5OTDYN2xCTHWYF38VTuS
ziCaqJMhcYvYYV8cmtk/P+fi+ODJHrtcA3mQnVdV77/5Rn5OQOhHpq6ylHpt/3VonLPD8DfllJNe
Vry8iY7JwYhW/b1v1tpM+wDXvP7zW7DTgencZsHJw0+w5pcuHKH3IWGN+9b0moxbIEFKaVrav9E9
dtBKPoyUFC1AnTqtU4GDiIw8q+ioQj9CJXOmLXR+bL6AMbHb73C8RHjJ+TXhMru5ZWd/pVPXF8hz
0Khy56caBcpI29g8P0lW5c0gK2rsWdIUl2HIBepjvYkkxMpEDqt2xlcOT65VJcbZSrego2HCGGX/
itmcY9/xX9jaBzE8CJ59mzR9+5for3dfzV8J3+WKmHF+upgx6aoVp8HjIziqkdY3htZ1Wp9OWYe3
MHfXkO1WNSG+Ci4P1NJAN/oVFEIKTo+WlLE3+B0MQeNd4O1uvhk4XWXyawpR05Fac0rlULnIOgwL
8GlX9X89k9lSo2Xv7EQARjFwX5a7EVt5zZwieeZSP+bNIo/Nk1quiiCfcOCyc7X7Q+RILY1e0hJc
uFX4RS89sYhQYySIjbGZgVQuuuHR1Ny/yhXpqLqS9xBy00/F9qAWCvKoClG7Q8mIw33cmCx6831q
9/E/mZeiZS059ff40D3uwoaZKtRsrqJtcwhbtwf4h+bUcY3aNt8n+mL608H2NXbfVxNlh2FWYe98
0qDctFJlaGOqOC7aO1cIEJ57i0yS3bCkrgVGq1KJhHnVkw6R7enQjzjPkASQyvPWSQX9CVsBaUfd
Gtvdz3WOXq9eSRjv1YgBkTJOzWV3kaHPk3Dt9fQeks3oeDjwPsB4e5PgYuCcMxfODRDEVGOJXy94
C+wW+iGzbPKKnLkjzr9PL6zOLZ8Yos6TjqlzWFXHWd6t1IuSsXms/7ztEqVB+Vu42TAAVv/ak2mm
EneQnVUOSCP9rZKtB3H6xx4PFaDb5UAV6/hXBtFBxqOMrRsVibWtcnz9tn56TqIe+kS0pyiWz6U3
w4V6feXYOFRNfxjF79Bsv2Es7q2mxPROrzFV0MEbt2eDTMzjmL6rUDTj+XhmSVaeGskF95YSitNZ
qhax/bNlRxTRAvh5At9H47MzLCQGSMLP+i+t8lPwGIBQIVNXfNLWdsz8gtWCPjJrg91NEfVkoyRJ
6CKnrV77ey66CC9Gx/tDnFV3e2gyvTfmSjpNad5l+FW3T+UKvjzD9a96U+tgfIC8+lTd2/qmowXX
RdJi2X6/HSD5Hvqo9dnCdpFAgO3NoTnyW7PTK4tnqZkyzxyIyIv/hcqx9aLbRx3rPXZOxfuaLgWh
G7QqTjnhpCMU93FqqR5vK1HlObB0U2+m8Da7WMI6fIxLtFrUW1J7eBkI/4V6O++gGKvyQCH4VADo
4iiuyYdvZdXqq4Z7xrO55NBawnF3ecauiS6pOZ2BWELJng+Gdgm4R4apCQJNsaJ9mEzK26zhCWk7
KWr5mJMfL+RBMADFSOH6cig5UG+Vd1ZgA/5Ni84i/ju1f2YLlrI36dEmPJ6WA/vbuHxpoR4/e6lT
BH87ORdy8V+dguV9Zp0AAyaes9rfSEZNl1aqbIx/uLigWfcAe2CQ98d1YrocKPVGDEttBYO8hIZJ
22NJ8NFImK02H/41LSLrc79/uVojxSxEXpuLk4jOJxLjvYg/DIUjDZ/WnYIvB1Trma4NQgvkNWOS
6zcvqLRGCEhzHa9CBkeiHCqjBOiRMJMVC4Y6ptGkiRuQsnaBKqiqHE9920cMvu0hZxfSq807+1Vy
kLJ/wKBrHOqPC4nRpH4DfMtGEkJCT7docPhcpbblYr4JZFxKrlk+qNdk01uO6ePU8iH25z6mIXBR
PRPHuE9sxxplBQXATLBCY2SFoJRJMXhbU5ZF4hQ/Sj76r05omksuLdxb/7oXffj2jxJRyXaUZ5j1
Up8QvwMiXkFRYCqemn8eX+VcaNU5IK4jDqRlBkWRVeAVMe+40hg4B0SRUEFX7Zuiml4rCJyBCxo9
aWupiINlqEC/Yk99pouomt76kIhf+qBEIVfVklDIyn4dmTrBHqwWtWGOeH5eAe1LBLACLqbXDxWy
2fDU9972cpCuRayIc+WHaLPcWUDw5myKP6qaN321dyIPKxvCSiEhRLEjmBe+3O6/mPw3QwzOGCe6
2xYmJg5aLngCEl8user2kMp3SFxsJEZHmCNEQJFiZs1CrWYZ80gMiKEpfouke7qbcylIaihMBMQp
OPITvwdwWoWOuGf8uId4DKGBIjA//7z25v5lgvT/AQIvVG4s/7vpMksndSBtTRy57GvEyQTrDunJ
RZ+A6X4x83VSougFqBFTLnTGGnJB3sUQnOhZcy2cHxNBgG+/kM7NuGlDKBTz5CG141R6o9s+Ppmv
Az0r+NYLtK58V2eIrDo6fb90FSQdXBnURZHp/z6HbFyBa9Tz6T0bLU8SwbC2C+q3qkAvRYwTTKZb
SwzsAH52CE9VwfiyUlc2R4h39OCdEs3U4SgKQX0WItK40I63wQeFH2kWNbcrNQOjuC7CoXXCodo5
R2R0So1FJX4X+DDxLjDMGptFiu1cVlp4NxtCJkB/Spv7r2RcUzoilLcXToeKKdr2rK9JB+hd6nIB
WKS7PdsqSo1oCVthjPRQLCjkBJt1NKJ+k64eYHl78QdBXEO3YZXAvRme0+1WpLKNTbI8l0jt7Yw6
jFiwSqhw8qZACK8+1q7hSQ/vAqQu/F19zvMrqQRIeEEkheN9spwjVinPeoMVH3ytmJ79DWTy0tyw
HKH/QOaXxn78UwL8gCqUgV+qiiIAiiO4Bu7ZBjb4oqA6LXgHmzcusKAM5MvZHkES6cgn/Wkxb1cW
qXi5knRBfvoLvOZ62FgXO6SXFKbkdSNZh90RDVPw1ohxLcG4pQWtR9ccW1+bDMcyW+L/Euz4wlJQ
B2r3QiP2BpzrhhXWuXbzJvVVc5/awGwbiLpD/9wTTGqiIq+S6g3IGlL8Jo5aczOP4Ta1Ay5ykvRQ
uS8Z7uMrGICzeab9BZGGLnhc4I4xyXyqt2B6jbZxWXt3+POijAj+vWyoUSbfGJlSpmvz7mafkf6x
S8721Mvnb45E4Bh8wtxVwVPI7vqxYxS2G0aLY7qZTMLiRl4Iu7x+A9IehDhrSBDVGZYfAVLHEuPI
T5YlzC7MKZZUqTj0+oZB+A/2zd/YsiObLfzgNhK7XcKC+YYvpHuVVbo4+xJimAKoMuIWWYWyhpO4
rN8f8GhYYWwoMmZZ8swvqqFZrIkaKr9HDph/INFUwshJWtJnpVL83PsEKGPuTE952JNYgB7tAZuo
2E1D6wgj5qrrx3Bn0TiiRqG4RydRuzEnTy5oc5VsWUBsDrFeWeCjHYq+7f5xb7HqMthqWrq+O14G
4+BYTiZ0Af2LNC/TK+FR/Wqu0eombsqmUiLtCVq2TuLV7LlP6LufFodDhJtuWsvuYWUY+EMssuUT
E5or0o6koz8Y1xUK8Kub+QTN8IuO0vcDngYYYqQ6JbtsCcMkOGL15PEVPxzGe54o2jw9hKH5/2uz
EkJdcinsNsWnSOnDXtko8V2A3yVxgdXwBp1w6GLClbvvvuwWz2OCxCDdlu+svJl2Wja5+5djMNEh
iGhLiA/COggqXyr79eSWCksXPc2illEJCOFgzDne+Nvm8bSkYN5zJRJq4QtAbldLvQpG+047xzmo
yPne0NDkTBtPiaVgU/Wu99ajLwrjgbJL4ZaF1Onz+sXhZWa3L8/ULrcfYk4pmfcGvseAYTv8P+Lb
+uB5JR/KkZNEMse9404g3t8tbwgBNCbNU1ZOPdi1EYphKhwhMgUbRe+g86j0rDSOighMgFxEsMhu
9Fq8ncBgYO8wlYlxrn9ZbCbEdnpwo8Gvvk/IZuDfldCKG7JTnIYkBu8TKPeSBLkYuhoalM4ZgmD2
B1VDMkFWjoJxHW/6K801lIECZPDB4xCgDCuNHhECk+Y/byEdzYtzroyFNT1+3fHiUKC56htB40ge
Kr684NacY3Dmvx7fgFZ6RNLk/Bxuz5iYFNqRYoHQHKkPXRUsmQBP795RaC7gYLn2FZxb7hakZ1bH
Oslbq2kymeJqja/xFjPWgmhbXFe9ap+jBJur4bh75fcplweBJhekCSIdnhvJEZuWEOJreipC5t7s
NG2MmjpHYMOdqyg08iXzN+6AkpB8HEjLNIyFNlhndX01zTy+oyutynZ5V/ewTcwW5LbwSYSrAYIr
FVh6pYNrOH9bk8fPAk0ftR8L2A/S9LNYsd2YNES+MO1/++2+o2daFgDqNoA4WQUUVlKaTqb41NzJ
6qgctSx9LbGNIcDDx4l5imCGxGIV0fCRGobw4K7d7V7TyjMjrZ2IzI7mSCDL0SSO/JHMAxSOjGr6
wDbPQUR7pqo98CDoOBET0y3BWafTW9hV9xDbFRTmQPMHkXd3UWZF1ZH+9QGBtsSBzwMPoL+N7Q3N
lY8aWaVil5QbWtMe0CwLGfW8FNz97GNSQ45GQDPH8U4imVilWsRbnUGIlKP31byunZwjm8YJh22w
l6Go9cVCpr9QCBnykxNWLWw0tsy2kwnjMlX1MqG06UtWqwP2WJU5PLatsjLQrGmOedyibzi1J1A5
ciseyLuP3V/SpuCr1G6zuE0CENth0p9ws6zGFSiOU38FnJkCJcideJhHjUgB8z2l6ML06mXLhMgJ
liSMHxjksY6Qs3MntMhpe2trr0xbIceZLXj6kIImWxOjlLCQs3OjURPGrnfJ1svypoNI8TterrJV
vsNhOV5ZA7FYcGjXe4ywNO+POl4+pcRSr2uoWcFTMpJ7T9aphBDdARXqCNzRMWCVEwRdE3xAOE3u
oLM0H7RTDPYQAEPW+s2/xn+yDMGr4EXF2MbNfPWrg5oE+iR0uV3aTcUSlGeyQz34zIIX4TeO1hnO
NGDBOp0sd8h6Tbv6losm62r0eHekE0oMRaXmMEzIgdhJKhtYXWowmvDAbFBxuHrgrv7/BEiBg43c
zBzbcKf3VkWJvjWUbniXEzzet6ojyT7Kk5Ef5E0GD1Q91cw9374m5dDrNYFRDuMdaOXBbdaFufM7
6gd8BDDRruwyQX1U38UZi9GnyIE5t8gSYJX2XAAPUj7ApqbK3MMRfpAj3vgxPtwsVah+qdbFKd5o
mnbDId8oji/k2BkCdrfHhBhBaTc/o+3X9/lxt0aLBT0PtJB/7rxGbZXInsKsVha19XvBd0usIgBL
a9ph+cop2h+p2OOz432IU3nn/n9shNTU/g04YupLC+0U5+dD/KtUCIwDVlMLfRe/ktydr0dO2d6q
Vd1vvyAYOhFH75VCdyjZHhFxAXScNHfH3NjBfbhOb4lCcGsxptr/+pylAd/c9TeLyZ3IZQkL7CIZ
0NduQkm8lFZzq1v+4WsvBdrwvjPeRgsLqg8QRSc2xIOGkJO6rOJMVzNZTOIQVZklM+5Tm2zysoUF
6Ou2GsBoOyfus40kl+9zmRWm2I3ebiIxDX3o+zkLZH2MNcsyaGd2yjDSom7uMrS6kgX2NG6lzWln
JOoNwCeufvLxKYaAuaBkoVygjLE5Celro9ySC+W9ic7RRuxk5rKyOWeGfqpBIdnEVB1czvOiPGeK
kplgKidp7v9DiJeYIoP3Fai4dF7fOk8CCxA1PNYI1V+7B48S34MIg0SeDdgHtoHffvXxqimDqRl2
Jj/1ZuPk/fvk+VR7ms4cZ52c4O0ETZDjO2gC2tLFDG9uxo8e0XlnVc9s4tgGGZzNT17Aosyp82U8
2ziV+ocYn/BMbCezEzzctH/LgaIrIKe7VlpGe4nx6VVHlEelRccUz2vSppv+5Xr6Ru5HD04ZJPwa
bMR6AY125KzrJTPsWmDNw7SX+JOYhJrzgE/kYLYIdMzpXqUi2qWVm7qML1RM1oiJyV0/RoN2gRIt
MDElVAduNFz6B0vWM7krrk8rfETC3CbQCMiipwXUo/8f/UCvQS0HXDfjcZB9yVHm00zOIrZ6w0kZ
A49Hh7CCFodY+XDjwFe/Z34YmsXxpLbwLK8/shK+F9gmRJo/avgvdTQTxYKQH1C9frTvSVbGIssz
ZGLdV4vOUatVNGl3IJjU7PLnE2hWn0WOsAclQF0KKxWSfwksunmHU/fdwiTKIOs873FAJkyIpDHo
VWW8qvsEvR4P6X+zHHbOmxppFhx5Et9c8kP++KjVjyROOPKz5T8JBJM1czMurtn5Wq6Dv8SRvPA1
BWaOOHyFHRuFhLi1r8Dwbw8XxLsE+wq+BPNzAtR6oIKYOo8dxJbtmiAvXZur5uY3nyzCHle3lpWc
Hq1hfu5NE198p/jLoH9rqX/rPdzXFVjqtPpCajpB19r/W9pwPB9Jvciym+PNxKyCepsOaX5V3jbi
KddNzQz/tjwZmiTFayHnvDijFT0UkXuSDmsXTbS3uADyewNyYBrzS12JAtyv04JcRwCA5Todgoe4
Dxdat6DqhaeiFvy0XLt32gSPR2wQk/q5mRO3gzMWddYZlXiXx9J0LPRxBaAfSJKgjKSI2EZwRtGI
peoT4y/1kBi2Npuj4CmP9R6Dr5gGJSop9LnXUliQeE10LhudmMeicgDGovrsIk6z6MqSuvDGRpTw
4PV73RjN2J8/uWa5u0QJaH0dtZbRtioEu78+uPTKMO4m1NAnkWX+ozxSsR3SLoo+pti9J5XYbFQC
SktBOfTjDirhRZnRAuJnXfHBlm8dO9nnpjhJ9UEgxYqgsBwMt3mk/D3gEVmTyp/mQ7uv+GvXEdah
o17yrWubUuP5SLk3nw2AQHosKi4OCKvgIEUYsRbA6jg/iHBvy2kurlhPAwbcrkYU9cbjDmuJTREw
yDmeowtOOWPZiyZKxuIIOjkROWk8kq5TK+1iYTq8RaO3op8rWCLBUyJXV3CcencYsVpmYPt84T2M
OMFjeGAlU3oKP16eNsPvY6H5UE7gX/Hy3+Huom1QC5TmZBOPLA7ITI99Oo5rPFfEJnT6516eG6Sk
W5axFariUwb/+5NzefyTqhaAob7YbAv5qIUizCwueLiPZ6SXhukJ5EcSGo8BwyPSLlEEX335s2bb
9e5qNsTfIxnzN4S0uLYk4XAhasrNG1nnEiwgqaDyXMvCmk3Mc2zGuRkqVG2f0DawuYw9N6X2en75
vwvKJSgSyFkyMj0fHWm2TM1Z89yFy1jfYdsVb1wa8AaAOYAKxqP4GR3NidXHLeA0bpC0eA7kswh1
JJ8jAiU4K+ycqfYyP7CgvMKj7W1oGWd4MutPdaf4gayhfWGWN7csvyjEO3yBk3NMvh18yjgLxjG7
mUYzhcHPW0aIAGSuLAgn5nWJ8Q2x5Zb69ZLahZHGBdlRO/yzhVRV8Xf8XqjJFER06pYYd/LL8lRc
bPjcRket6wnsea5vmav5h6B0vzTkfVKDQEz0jKlFqL5u3WbkOhLCJ0dcR481EN84mtoODanojAzV
j3v9doG3NS5fTcuASAYSaWfIYzeBA4xWzud8T0cSkglYyOSY8/+5LmNL1qO5MBpzDn2HHADs5/nM
4BoD8/hV0oNjAcLQyLFyElonX4gwQYCzjuTsLedkVPctfeb+ODOLIpr++WdYhemsP9sJ7AosaVWT
vId/zISBbhCUn3mMNMmt5Bhl38YDpQBww5VAI2jcwoy8pL6xb4/a6WOGswm6Enn9cDb3NuEaBO0n
YrXKSNoOLz3jl0MYdMX77mAMDIQXXkIIR0ydJu1DTRkvb4o9Hdyr2y8Bua48QdVxN+qCgOJVEAP7
dc/UqhwnzpQARAUrXfdGio2bMoXL/ue8gnebrzcCaeb9V4/2I5ZUkKygGMnnDJ3TFinX284y0zeN
YbZhC/2t0QQ4CCYw+zCp3y/7WaPqzF4KtoJRYYTmekhoIMkog9rdmGnsYcAeSzg/gCPRUoHUWD0H
AgOk34uhGdSK+snhlVQRpv1UWeZLTQ4p1/7Z9Ms1GKJ4UgTsL2HI+4RoYH7w93uXUY2HWphEo/g5
ccbm53KEXZ3qlPzdEAZRSfdItsie67yw9R5ZfP347BruzkJg2OkhTPEVy/son5H6JxsIsrnZjKim
3geVIuJ4pCgFUPJj2ts0i8XwTqMwnJbLc/XP0aNZeBFBSywfJxH1tDTIudYeK00HYNbi4f4iKeyj
GHv2PEsl6XI3Vy+9KdnKUA6gMpitX0wtDri3lxyhjDylK3P0SIMkSgDHchtjPnFVNpdAP7awbfcF
8237VEGHnIlNL1ZFFzH6pjNtjex2XxlyZox3sAAjfNMzssZX4Ff812opH9K9uc140wO1TsyzEa+V
YfxVv3BoCC6hfQiZ7Ok4GdUsrDSEk22sgak2v1HVJ4s21x77q26Od15GVmSN9KiLW3mlcLGI+UFQ
DQgjskMmhbmGNbkyaT9uKeP132h99FoGbguZfUcjF0ePxDV2BQmTszBH2Mjiw/RG9KoPWUXU+QuP
HfV7zREK795PNHVdadkSmcOdieVIlnlqIjsW/ZI75MnCOTfo6laQJEoG52VJP/8gH9p0ldql9Xec
uKN2Oe0XGkuvcHC/AozYsJOFesX0Vkp31KZPkPc4Hh0KmSQhSucXI2N0rH1KHyFwoH7mFhiEZm3I
jH9bCtmg0XLb5yDVFU584y+2+kh91OQ22Pb3wkIoYml4XvEg0lQjCDmjBNkC6CgBju9fZCThujgq
GeTryEjzuXgzp7PGWAbNI/9O1tQnnbrsSyQVFGJ1UPLu2LDJzQAAS6jqbN5nnjeXBOpQnMUXI/cW
x64yxEMl5AYuAwiEZFKhxFLwFi4t10uWeLbeIPZ3BWDRVgsKIi+SIJeN+5mQUNfhnwlNIbq9tzEi
vfQJQ3ViiNa1TKqu9aTdndfGdfDFlaOL4CWNHVWDQzqvzxzzKv3HrzeIbGAvFa+fRMRuclePwrDA
1v84+amrLyjHJcpmbOsMivSANHjOYfBNejaqYm6zNQB5JvXFwMRyIqnEkYUUVO+pMmK/nuPAkCZ8
JvyU9n5lNcqLMJTT/hZVchjg25Ffo3T4xgZwQqW1hXJl5+7g305/N1MZzxuzzPztBIMD/3jI3a6e
ger2sAPppIPFQRE07Kqfq4eURyrAnJZQiLp9YNGM69MlsXjdanJHXTeobH/hQzVXxHV8oZLUTHeQ
k4ia9BqiczieZzN8oR6kY6HEP/7OKer+I2gFQQwB6AoaQIALZ/RehMIAyv5VepAyqphi69ZbGgUf
2qrdW44LrQr8ZESY7IZ7KCfwjeh2Xd5p2dHNacxK2gT7mpKJaBz8LAuJ3K5I03LQZ1sqclM4f7OB
EOn1rHUA7cbolfXHUtzQC8bPoVGu73i5pUligK16BXzSrymPOyi5L+AYuKHQCpRXujw14xN9U6G0
6J0U9zmnq7yKi4G4t/R4iir6DSr2Ac+chjfeu1FTlk4fX+ZUqzpXc7Csq8cziwpgqVYNF1c21yDz
a26xsiLc8gWLexjm5+YtFsGMC6K5zfgN6ofTPlwc89+WTytbST1n9h+XO6PloZUcHi/PUApceM/i
kBdrxDkAiQGnt1O6T3qvsJ4a5fxQ8YEttBDkwTigbZnU1haXZOwYvcmsWfo7EbnRw4PyS0NbMmpJ
s2BrfQR/bZd2CDmXGNM4BSZaxATPU8SHIRdz3C6nm4V7nsOzEL9S9CPYTuEZLd9EeEu+w5xxYnb9
PxhzPd3ddufj51mmDCQFZkOMN18+gTO4Nc5DWg4miP6kGgxJTVFhNiAEyI9I/RVI7JUvpqDClA9P
HDGQXOPH/LkinOue+xreSX5NILaPnu9Z1Mnls5sXWow2dKOHzwiFdY2LXijhoXXYzQMPpPBUdgat
2QgNx2OEb8xAgvQqxMEwK9UzjNkotwtjPMk5KRRyY1Hm7sF0YI7y8hsAF3+7wB+XQ7aYmQ1QSiet
K4KK1McC3egEpluibdwmA1+W06DM+nwqAWg9Petf2ZIBkuTbV2N+xEE0Ule6N++qq3zoHs7XI6T6
qu3VOH0qO9k9DPmsu61ZKHgWCIH9PBJJUJObyuGDryjh6dwIdn58w5jQlT3CGyF3RezDtAWBD19u
aCWioIrp+u+W+HsJP+9nYmUOzp//u5FmX/daeLCk+YTrK3DQZL1tSRGg4aWJFgPnBtfHO+0oHUfR
Dmdgt0WWNysdIkwA8IdFSWEpqgRJZPd/cJaj0433eRw0tte5FIdpJKB8WY3U6WyvMl2H6Cu2FT2v
XlWuMXLmjGhkrLtBovUfW+BFw/d5ddPSuTdNyx1Cop3cGJPs+3i8Dh0z6XeBc4jZUUl2y960j64T
+gmHxaHBB6fNBwzMg2gpUPUW5LffnC91D9yz5JftpbyM1qcUVfjMYTZatEhx8WMapDR2ERRuOVhm
MTgV9C6VuyeY8dPvPqaCJbcT2jfMCrcKllwYsKODhHSmm7eKwedy6jUc/505UptjLuE9i0Xr3+gK
CE+d+2UYFmuNo8Q6GMNlQ+3S8UgCBnlaIi+harByIBXJs+hWthHE+DZBrrW2GlmocT+W6g2kTbSO
2ZP+SV/4wJ0U2HWcBXCv3Sa7mu8lIZp9Lcpzo/+1dl/Mrk/jp/6kwqNgL7UmoAsA7tG51PM6tL1M
ulTlch9srvROAbnzxY5MoTSpShIha4IOVqdB6ZfjU1YjbHzANSeVhUUxFCuEHt9Ka8iv3IS5ro3c
/Ry4DJyZ99r/lVfCIN9GqkTgl7jGHJL6eqbq4StU2TVtUheHR0nPHTGJZi+yaq+V4vnQNXBFyQmR
cfGcIGRepjGRM8QUTTNszHqYcg1RpTwJmIJelAP8/oRxXAc+BivVOWPSavUevJSVlLDtITjjope0
m6fCpSQ/dBg3Ng+M1MQkxGMD8WDNuJZOjaX2oDFQ+oWZbPHkauHToueTiwLDrtFefP+Ndzj9jwJZ
RDgGBc/fFWMJ3BbzOMWF14U6GD34y3qlc1XAt631JWXDOn91chzftSb83XB1zOqqjfOGXSdVyeZH
0Y2SQGSrSdATJepe9SK9F+pjNkzjnkb6eDWf14bUFgF/8XT/tX9Aspohk4n1ApVAKKeePnDI2SwT
e5TJ3CuthgiA1RdS922tr+cPYgILQBR+0mOzlB5Y9DddRR23hHaM45cXjHvRIg82CiQel+CYiyQj
sYyObqQ8j3UHlETF5ppSLutmF8azyonUCrMIUytYcF8iBl32Wltz/LCRo/quAS/wkQ+Kn9F6B4hd
uWCjcIMSc8lG8NrggrjirIt8xrIrhgjXpnJpmE2Fwsp73wBuSI96MnRGK4duAsY88Se24YOUx+GG
j1XtMJdghG3rRPgN8Zbtdm+bWJ/RhflaeVcxZd5YIbGU46Ewm4yaQqGixbx5FmUXnv3GMBUaAf2G
2lTktQ0uyMhGCnC33uDyr8t+YvL4n6M/7K5VZnIBX8smVGn1ku0xDPtCQiLdF/ZCEYfgKDxB46R/
nL4208xU9LI44yVPcS8C+EgLlLjlJCWdjX5iB1h+rqjDZ09C5pMxoG7CiY2LeOqC4Whnl6Phlvv4
GqnO1jjCwuLAolMUR79bvPMk+2h0Rl3lhXKTjR5K20l5JHrbS2BkAcTgJRRp+Q9a06iqNQ++Wq/I
PU3+4FvMRXPwkHWfkR4LyAEx8+k5kQQVWgpM7+OJG5/SiN7F/cZZgZmGdUFduNDUcGYhTGVifBwK
MBLkeSe9riTg8LnG+ICPxixYDGeD9AlZSPR3p5Uya2B35cJDzJF4j+/ldE7KtSYiOUb2J5S+a8Dq
jd8+EwAgEZ9zuaRSgsvzFV/FGselYROPYQGoLO8Q/S0kHmVOPICH7dpBkcctukfuy/3qZ/f93zdX
SBlsuZBuoP0k08I7LY+Z4Avg8fl/y3tN5RRn7aS4Py0N0Vq4rTfSKS9aFmILJkhtMJPYG6azLevX
gDuCIMK6NSj+mMe/Oq1oyfzQp//hnGfxgNexihqG3LjT1sZi+MMLQoi5TtcKNhpX5aZOZZZxRW22
iNihBKkVLAL0JpEDcfQ6FwoD/rSREW4t3qURJsYt67UFn4x23aVZtZVxZxzC81OKjpMipXDNDrxn
1wBRmkE9W9MohtLn2op3NtJf1kNojHn8AN9naul2qBHEB34vkWT55hOTm/QoLmemMhL0nBg7k9vT
kKtxpX1kzw1AftlvUsWvaL1jIvHKllN+EFvFp8QiAB5fLlEM719VlcT5FtqBRTYv0bDOxglcUl+G
5LcOKPILSjxaoenm8yC377osh3hMCG2Q8UsHarraki9DubJKdBKKcUjEvPyGhn7Sv+GuVSlwfaGQ
FkvCgQyVIiF2l+6KJ974XYBylppK/zAkYon174csickoaBKDX/E1p4H+O5WAePHd/sLVRNTDnt6X
X+9I98LuA44U4CbH0oJBjUMUOEA/zFEXde4WaV6e9vJ1/DNpZNEeJZ917/S4RKLo/hqRpas4f3XL
how6W69p/Ajdo5oPvYJBdXCxN875mB9/HW1E5ymU2R4w0FY/YzKAHfKVnbg7ymj5GNibaZPuT4sj
3m/6PW2wqpWFp+xWEmIL9MGoNlovJCR94qrUjxWfMhE7oqwXVt27jpdzQRQMNt2vmB6+V1Q2ADej
bxqSqNwMeZAFSr665GYpB+IAyWfPlKtCaanGfGyCIRbRx1kZ4NioWcf1Vszsc55m+1MbkojKZJbw
+xHjNsC6P1USWSz6HzFS1M4d3SDqcaeHSdCAwPCxdylHXp0sIQ6BpXVsSnPrs4c7LLkQNFmXbB3h
vAc7A+WZUIQinDRVutYE1EHZEzomi7rr2HY+F5//p0WDy7SE08n67Trh9SFAr/i0XSR87v+iOrfN
tOFLKjFJqlGEm41EOqJbXug8NjJVo7tX4FD9vFp69Wit6otqsl/SXPUqM6v4YKS3di196fDNG3iL
2rxFmfuosuX7cGimaW7rxA8sRNhsEg9WXVmcvfnEeXEGzE+kHkcaHPK25jKHNsOTghPO1HzlVrU3
ajjgwwzSWjumEyvmpnp3AVsKA6ZiWM+HDGk3BIvixQW0U8304mPSqOMZS1jN8THutp6QiV9NFsjG
zWVrrK+rllHTaUecUvGoGv5Ghs5pWggz0eDt5yEcnfOiJGQlf1MAYH52Zyj6jYgqXtAI1rYtKPXx
7MPwJxi4j+2dQggzg24sYDht5BLExJfLp56QFaqwQ36yU0aRXIyHHlYNzRBgoa7QYztts2ARZ3N5
ZbVA7O2MCmG+TX9vUxjHkxpcxYqC5xWbX6cDdifCopOb7mxxA8x0T7Jukc5WjCZ18aZ7ABpVbSBu
mn1BuPpdc/knKAR2U82QkEoblLX51JpXBTt0fZCUzQ4noqfoZGz1HxEavZeDR5uFRwA//GsrzI9J
vvk+JTURNbCfB21cNRyL7WCuuvHokAQkqVCtQ5Y9nG9iFXNUCIPtM2EmsDj34h6nU2nsXEfxxFKt
tZykMzLAUT+N9HlP7XKpjaJMf14zcmwNXvScn6bvWtcY4DNnwUbEXw4ZCIICAh2+h7UF2LbxN5aF
4O2yOU3Ez6c+PMdugru2hdE2qP9kfjF4qAjMUCpoRF7yIfOqacsttALr3JER2wSWm0QNa1BT8REC
hCCZA0J4vK7SFr1sqDDAbLu7235Uc4ihk4uYd+6tCjFVCIK9/gJGapm+y3OlZ4/X6cNF3fGVHjAO
zYQGpREGv9f4L0hSYcIhYcBTmGGbldDy+ZHQwSEFyi7UVuqcvh1P9pkEmpuL5Sjdpe5Z+TDlMsw1
3BOliDWZIvJbRg/AAl6gPXuPGTcEk9Di9eMECDh1dnv2YxsDGOndLadx1nobDTANJoSjfaA4AOYd
HCVKO3V07azy/pCGjUHqwpkENtPWYEC0WV0Mt1aNfUeo2WOAfmvclgNCLTrdh9OQ8PshyT0/BZrD
5HOPwVuP8iKFHqKhIMpxu53MzK4oGIKMMVWrcqNze16Ks1a59byWmutUXu8WiYc9N9L8QpyAk4qT
tykwQc1TW9vtAXADtYg7tkSXvCePLjrjIe0wdRjSwnwaIH8i9rd9nO1hFOPf+ggEgnAVqSe4YTxR
NSHqBKMpbCj5Zw9HhyMCkQ3l8nhu1zc+nIanLBK5R8u3VIiWrlihqPOnm0iy1/LFzBitGRUwJkok
Gpu5ghQLg2tlDu4ANa6qHuqJCBdZ08ZYiEhbRtwvZXMQcNYaDSM72LdWu74yCNGKaDldNB5lo9RB
1LlUPq5IpLu1YBWYG8U+/nTyEPn/fAW56HGW+oJR/cAp1bTUwOW1T4LRqxpX3FSC+ytaprgia/dG
hnN7w9iqZKsBiJqEqyhlmJa0zIke2J6tSOkkE+ozntj6Wqdk9zMb/aAhf4EDDBym8clkY+y+/V8m
wx+LWnjQ+nVYO5oYQt8uD8AiTXzVf6RdxKH/cSSawtphgH1Rk8BebV61yESlLcNJ4peznWLhKy5K
ZvgplpDkWmE7QU8cH4BiYl45iypMlgQo9WwZq0X2uXpIUwkgeDUXQ51fpvVue069WmBVZrrN+tWb
0uxoOvdjueC1+1XfOY/kmkRQlHLtKnf6wK1djrfiFtLzP6AL04R0EugocMnKdBeeZcsWZFXv25MU
Qk/Y3+TndL04fF7oroDqq/GDikA0KKYIMQYQKlw8u0n57kCr4ZPhv5Vl5kZRPxo8cRgyrdADv75s
zxUMs+naXCsfE9NGTv8neQzIcFBb+tCUHTeWHftggn7G07GVkO0SJFYUpghf7ZAe6reg/KkdIuc9
rIBxZkb+4MzlLpSKZG9RNDwjXTrb/oq4d6cAC0u+JX7dZAY1BWqmQ3WAlMTspxLnCKVVhUmA3nYA
7ODiiGncWyPVZY53uPWwhR76VeTEUd/Ng3F5nx7+0fMSq99yJ1lGvIAHwp+ybefPGiQGlOfvCEH4
qrxuQ4xolwjJit+L+upKJkiptLelK0pTFfll0UNqcFg3iQaPQwuhvovy71nlp+7qTbWBaAwKh8F2
toiCuNb1YnXcyMkbgBxPz6QW1AMq1rmXa85MPJKqeDFulAqEmdaluKdACnGiLi6NRHfdwsfmZ9qW
T+7GY5avhxjif9uTepXCF1Mnj/u+NyZWxxk6zAYKnjnkuD32NCA/sMS+AFoPjTBzgP+635oX52o+
+3+K60p62/PiF+smTMBfrDGiUBM25lzCcgB26OxtjT/DGWlG3NhNxCojdDB4T1fosYR+9Pd8z5qR
JEnX/QUzmlWsnp9MKYwV+JY+GjDlXSoikzitn6KBpbBezzm05zAEtuBeD5dkc5NsZCcNJhdAlN1K
MPadfefSyQTOfTLKujAFrtgQELBo8EL0wPvZv50sLftRaWHWbeOxHgABBp8A1sDjnZEXJM0qsndV
mJXKCBPXVqaW9UHIz4TTmnYBkPBHlD0KW1X7kf0GVNJVMVafkuwdDcFaggIGH+mBqABmYi1aHNfa
Gn+03D+nK3yfpc1nl95r7F4xDBuxC+9jpFXe5u4Cn1pbYqqwRq60N/yCZS5gajtXLZ7+xujm7BZA
fQYT0bZm8Xyk1QTTus8uuhdtYxbak9OBa0WMgAS/sUCIFwIxpkOb78bVgmhZvZUdVObQGFRQUgHG
x4UokX2n1oa/+YwEnaT2NeQERxipYjsla44vPHnUPvVDi+FIFVLtPIdvk7b88PwXqQyRxARh3voa
eWTMz55YMgZWxd1NS9Sltsdcuioltt6Yik+wUIF7pbtxQCwh5RdM6jlL8H5iTXwAT0GR8+8LcBBf
fUuFhk86twTpTIbyUbq+RXgdiE9OtO9ZhxX3gl5SuSJFH3NfV8SxYAG5nnySJ6Uo6NECcdE+LfY1
mb5fmqCPvkn2K7bsRMa6V6Ux46FaYt0Slpn/5dVh/lpvocWlVqpvASU+Pq9FdArbBSV1ursCQj21
xs9kRZd3DtWmH8kFhqDdGyK1ykoit1xxvH31Tekn9Z+hRKwZVFEH5MjepCcyIy+sxFKixJjDcaHO
t+trhrcXGmgCDdRje5DBqwBzy3HCgJIyq2T1UBKrTzEp8+7rvnqOAa1wGZ2A2Jx5k+nKeTKPjAuM
PLKJBKEwag2uxEeuGXY//u6LH7R7ekGZfBlIeRxRReeyhIZGcLQfIpXkYDBJIUObaAea3gsKcEpB
ZYggpvcb4HrcP8A1I1xPI4Ckl+Gqkp/RUY2kHX0rXU5CltTstKyCPTrDpg1+xIfSZAD9LZat3EMM
I1zRjQzdQ4M/LiRn6zi/X4mhCeSYwo9mvZlTtC5YUTVJR0K3ErNOE0kGFf7UEWF3gQiq2Dsy1tL8
6zDa80Wdxjux9/cpSBX0oFj9XATxz0EGb5jTQycqnHys3SP6UzYPPaVly9cIgY85SWqBtWb776mL
PMLDg2zkU772il04NV8ULi45vIFaP7kL40361HEQPs/4JNPNA4Nxgksr19B6lAQXeyd/1XiU8ts/
yc6loVKkfOgrv411N8JV4feLJMCXWrJpPiJK7jDZ+XWnej83beG/doRCzlhfq9qUkaTclS6Tn2mg
XeOhYUHuuPAC+b0OYRH74bKk0Tu+hEa68yKQur+dPPoCQBSXxwrrKoZCEoBhe4uoXztAHdRFmN+A
+cd2cYixOkUhy+tklAUsPMt3P79SY6C/wTVUPZonl3vyyr/O5fbNm4P+AQlzrOm9YzV12TRvxhU5
rwv06eLzQWAU2dV1KPp3l7jHIFV38guEgDLmGsV4R15ZgunKvSyjjh4UK8bixoLQ6kf3sdQwO9Pm
LZlaMQ7tF/kHVVp34xBitLNtuKYsmW7tsMqkLUlBnB2BPA5wGavuS380ELisKsVRN9HtHIh6qLHY
qKS0vYxu+FSAe2rZsOCcA6UKJGwWXOGuPnWfB0pgnY2puizP3Ouy6WETIi3x6UztLVzep80aG45l
bJ5VTTtuDuak2EQBreM3BUHCwNEthU97F5sZHuqksThf8b3w9QkGlCyZ47Z24axkvUB/v6jjlDUd
oA93DULoVvEs7pYAAvZHTa0ON6e621rJaUFzTyAjTh3MHZqhNiHOk6z58Qq9J05eJiy3UixIcRkM
1w9KG7pCS9NhSB8MWStYmvO0MfO1HMCeno2rvGZ4jHSqaRFbg/RP8geKfvCrKIRWBfCg1s7axKq7
hj+7k187gtORXQfmgQveIueoY/M8hfljTZkcgVGFGN6FSf8xzWBgrIWULpiIevNQNrVwUqOSYbqN
nClFgALtOavqxgSNlUJwkO+ewTpNik0CiCmMFwnDiJnt6jIPbEPG7cTLYPC2bkfBgshWKrhezsd3
/0m6Lm/OMuLGQcKW+158/X8xnq5HFSy+9qOZ7FFnjYP1oet7dp3ImuPCF0NV+3W1IExM5jGnAyz+
sAd1ldQAtdV12jIOxbjUmmXB4K5x9SX/yJuUPez6P+gq4kLnCvFUSyKuqmMR7TTFZ4YJ5QIAoipM
iBasLP2OB5goc5XXs+4pfK2xOvoIJy4osxWXQcxorcgQPk7psgm51/bW/4EJe7dvLt3DgFhmbZAP
j8uOAIRGiSZIIWxX7frsBDL10SGQ7VFGqENZO5DABuXFr8CAbZ54AH59/oLUf4QT81zmd22YKv4B
4AG3a4PHPobjcOQROJSUr7x+ManvME5fOYh5ttDuAkQwqFAfzC/1UhhiKBdu0LcK4QS9lJ1T+a+g
petWDxctAbAPEE30P5c6ZNJj4RPUgugjJ3dSp2M7gNTVKbnZ2q9TgiTEjgpl8SHeB0GXvfPbBkku
l9aev2MZexEWWtpLBWhJLyVcvVV5mRZiYLZrCUt4AdaGlolRZkClC9eYsEuMfjPf+dpTDRC19nj9
QEeYKevmycOQo8DO2HMREYWIv8MC3eZAPK12VSMGqVxm/HDloTR1tGvFBu7zXfipMWiiXjvygsIR
cRniLOnGqRLs3V7ZuVMQGsq5UgTKU7rjItYFZgvXOh9rrIZnN52KPHCVsr0I4Bqc2bCAWB71ZVup
zv3iiNU4bOBEvPrpj+plVmsOfygvE0DcovxjVFEVEoBBRDpIBxTRfFsfOo9PKSNOvbfJbACNQvJ7
PJE5uZtSErqt2j6qwD4D4ZrAVZuonHKtPEJG/a6lJrBiuPTJTg+U920pUSlI6+fRdmURKJ3yN8TP
KCoYkmFYxq7e5cBn/QhPh9c5rFjj0hVeVQrAeJFjTK1DeHYNEOkBns1ucgaafGOfMGMw2bE56irq
mixJt/BtvLde9QpAe9LWi/6UBBk5DKNhHC/tMwytRucWwiW22rbX2xavF4PI4jwGjhF0wv5zMDCA
MnvkY5ty6sRa/rAEEHi+kNs49Z3fPaVFtppdrHEqGCkuiizwrrj1e+rYiHf9UQEJ+tjUqKG18aP+
SAjqKSg4My1Pq56vOhWKeFti7lqyIsIPQCNSMVxgLvREt+4auzQSzigeTkL81Jt7tzWBHournXp6
uyOHY93HQVHCTnNv42T+eq+0GqQjkukwBlzgAfowQzR5CCYeDHnmu1ic8iL7nHscsMAC1isx7+Sn
ZuZIAV3K/DM7CjGi0b3ZuU3sVIiJ+l5dRkQHL3kKkt6ps79dV4OyVhjef/K+liZtkx6S8WvXkUV6
cMJ1rpG0ufBLJuvOk3JqD7FRQk75btQ85LXTMVJY7RjL9s0CwY8NsXuzBQZuU0zLP85p2aZp4x9I
VC2BnbBBuAax0nPlJB+o4CUV62DRQ1nQeoBs2oetM4nPsmRSaox7wO6hIuMU1kiBu2468PcEXIai
uWqoWxGSTUEHMV/pQkn3PUktggD8TVmJzmJQiA1gKnxMS0x+IABD9IAUqBWVM015uZNhpky4fDXV
ytVYbDC6guoyzy52fR0UZr77ufGm2NNn7VnK/HPYSNcLxs3Jm3K2tG52hkDCBhcwYwMSBR7QxXjA
u+abhlBvCvF3cUaoefbdW8v8qeWSj0rrTALzoutCg57YH3MZtRfarAkipwMql2XGYMWHu/scERME
dz6rrXCEelTL0xNELuc7frvRmJpz2qWil5pqkP3pVxKenRH9aJFI8zTXjvJwweV6mRaXooeC4Ru2
j43qYZoXgxUTAdG0dp3cVw7MNugHnym8wzIpisCLwz2og5E1qjnBkJa/WW00eI8w5VniVQwDxOiV
rXezcz5c+AFxMYWShQDM6UtVBB/1FmWFdVNl7SWx/VrK02gAEBD1Ip7NKYBg7oH8tibpgbrO3QWO
ysA5ps+lJx2ysfDvWlPHn3YWKxHFR6VMOFeylX4FVr1AjKFdFJbCLEqtnENhM7oX3HUwmhC9HtZC
RkWcMfy4i1jTqDmD8W6fvC6baTgryuMr89MRwEzgjsPBjUkCg0TSNWhVpxefeovPL5QEIGoUUsLv
H6fAB8jst5Cvvo16ZVZT+7UL4xuwm5LNElHZIgCk2osm99f2tzJpvzzqvbDGMDcZryRbsA3XN8pa
6wY1NpK/vY5ehRpNm3n/S0LCR1GG3v214oSCJpHWPkYWZEidG5X8wA7VOlHsnQlJJU9mGo4YiIvK
iq24nYxT/GNpoS/622KoIZjBDD7TUTlOePISAivPLeeLxI/O2uYzCGwhKh0Xqh6OGp4Etl0aMK9Z
d7c4W8HLZpuhLKdMVtgiPE1eqarAkdF8AOS2J1P8YniQGqvwuF4jizUC0VkiOCYfIMzo0Nd3XHR7
bbVt9E6mvNt0ZhKLOhW+uNDou6WY/6a3rizXz68fqn6/gBPWUAQmj3ILX4xwDU5oMeGUVlaMfmAD
7JPNXZEg2VtcT1h/jM/C08DCLhPpJAVehtzEeg7GPxjZadMaYQxpWY6GYOt44GvbN5vrSCZmNpWn
hZhO5e68LwdaXcUh6QJENaWVdtQ2fycWbcR5Ww2enCeLMcWr9D7FbnXK1g2dFX3fsnUYT5TInmst
91CjS+0QYhyYubaP62Uy5g6VILSuW8ZPPsT1ukaVIzW+6MUy+7bcc6/j+bk13iFEON1c9UYMp4YO
WzkJ8x8lfFdIUWoGRbSHI6X0E9qkJjVri8gq5lG3xASd9KabWUK4keq92odUBYnOz9rb8Sp5/oPi
MYC/Lmf6iwFZiB0oiAyfgvqz2SQWjSN+uQXSrEcrOYWdKgzUTWhvnD6k276l7B6TaJW82m90LQdI
TYMJWkRYTMzEkQEmN7RKMnTdt5EtRXXJfxjbFYXtkX0QDQFOPwIFfwNrvGCyetoyZHuCmG85uMIo
iJcfHo0Z/tzxJWGwPn3cdlwky99/32Z3iCy+T7bh2kz/lcM2rj4MMMnRLc7FAJx129rHTLduWq4h
y1Se/Adb6xvkyyDK+wxps1/NG40DVOo/hHdfk5qfUTyQ5wAu8iarOXr4xZNzMKUXiY6Aqa6LelEv
h8q2s2BOpk5egaY93/hVrqA4erVtA9Q/6+2771V91qegOFN8t5vSUFiocIEpsyOpsef5V6f8c+3a
bS7cP/kbShhTOHmghPHHYfdrsCeVLQokIRudaoaTvH9MHqjPBDBbF+Xw6jYl6OypcFryJeeHqOje
LXuVevPQy0S1HjPkzPE9jP1qvYp6NGnUgAySV6D8+uPI9TkHCvJyC9ydE9suQoih3xYewR78+Ymu
EJaZPHiQaGuITW+2jatIBZmY49/24+CJY3na866Zs6VjKEJHx8nAXJO40paMAZoPdVwkhM+8nhSv
zw5eZMuIpf0MamaPk8ticWMbhJF+B97C8FUXlop19mLMHOGl1SF8yvuewho0fkW4Vslyy5nfRBJa
2eWz0EQZZilowB8skyYzEZe9pyy4Yw1CqT23SuqSP3mjpoHKM4xBXX73s92sBHeQTvxvIypP7NeF
gU2N/ivmIk4H/2+zy0Ty3ZeH0dSzmxIOvNFH8ekoGxovndtfdLVtF2H7jVeLyZhAVfXJaRLLvFX0
WvzZeE70RGzHDD2XxzzCfOePWxv1tudk0Cdk1zJ09R52dTPMw3SU5dqYoDPi38kbeO3eB2Xat99I
JBnK6qgNFRKZtduzC6XBx6cZg6ZEgrYA3n5KgnHeTw28jWzhNFVsBSljH4f6Tqqu4qtkKKE5Dirj
WreNoSp97Jd2yAy2Egydl5gUCMYl76+XoTYnZ9+wGyhARPixIB+S9v587qJ59eGeHEKyVKdxdkCr
8M+pmilaS4BXzJ9zb+NbCyyfoE/A2nBTk+iVQ9WeFI7JE/nxySh+1qwFyTUw94DPqqqHFBCj85u+
dyXFTd5aqPZ2ResMSdTnBLlcFk/xwaPxCjFNWSP03PlCQrW6lUtI2p0wQ6C25KngBdlCgjDSjuD+
XJE76XBq+KY255CrGf3+ScoMtukMWTJPTHmLAcx/c7MSfv6Av79w8nEsraNijOOMMmTGGnsAgMKC
8l335V3xaxxruUEenFr+8GfHhw8FKm0416aY1uxws/e6OH4yBhGXKC1VmhwxhrpGnMDotdeXq+/F
yt1XOpsZpPdFCE8oesiHzUO0ibwtsnGJQsxMfhpcp0DurpcMqQzQR0eeWgDcHvde9NbfJdOHR1dq
LYHkeYVwpJCKjR/3XjkgjVEeoYwNk2+v18Scmt80ImKWTDHTHlHXqCuyeCmkSotnwQNkqfKWAFSY
iwFXxO0Y7vjCAZTL7k2KraxGBRm1y85UTEFacaiROukD5zCt4xmwSoPZxBFW1hZAaRRzddSsAhrH
xMjIGgFMwKtEf+OrOvnr6viUdnKHdkjp6mouvLiWw3yIO4X4m/t5SSK+loqoOHS60HH67Y1+fwGC
R4NOA2O5YYf4pV9aUlpRfzN5QQPBW8WfgPxRXrzeOeQUdaVtFNwmRBRQm/ZG3r7h9E7rkoUc+A/J
jbxZX+HpHNj2U4tRvVw6drgSPSnqgklEr4IKBhddEvHfAj/3vqZ+pyHtz6xLnYckAIiKx+PVJMR/
iMECWuM+ojD70Jbg5LqWVKV+oJaXhm9y+E1mHU+JItJc/YeGm3e3lyT+Fq1fQRFaw4nX7m6ncVav
OjB3T5beivkIDxpZS4WflnxNBe+AdH3lS77RvyV0fDUKPKTbU+MnTeTUbpWF++cCY6VRL8MU5Zc6
yUPSCtD7G30/VSDPLlQ2DYjNfEU8gos8PuJG7rurEKqzX44KOjXuqglignt0M81AN0wL5ZYhTYH1
/pIbUM8BeVYi+qG3089HmFdw6R2IJ58vWJ/dWlblONGKCsr2PvmkWpd2tWKfKV150TQaOWReptrR
tZi5pzlIm21X37m0aA35Wj8oXNDIy3xTWWqv7lLNhxHNi92j8UE9+1KpM9lA+G4Nan4tajeLOBt5
GrSMzsFH/QGpLrU6RIgZQxd18Vivub8ixYzchPEDQBMsYNWMMNrVBFENQBlNMZz2vruxIyaJgLe8
hiepiZUg39zvcjClNvgqwAId3VVDtRasvwUp7ENVyGh690mbmc8nLt8o0x8FCcT00lf34Jxv31l/
MY6cU27tg0zLaiSPKCuuWiIXLx+IVxClVInwgsj6x76vZs2e99wgzeI8luNFtUr2AbKVPl/7VRbe
fABlzUlF4HacwrjblMggTD6Ypgk3NNpCp9rLT9ptd9O8lfJvL/k33RSB5z5f+1lKEUr+Ho/6/LQ0
UOk/5apCTY5FzWEDNz08vrpzFFCbYAU5uNPL6zv2IgLP5pfB8uI3OpzH3rCsiNGaL+mPqbJbig0i
LLfXY6cLd4J+W6swgz2FEYN10d36KszhiMQeGsCopghJwk+CrBqBppYPTQ5uQBIonr4fHIizbY1r
NpMTzdghSihbfNdRnmwkv8unyVcph/cPCCTQ1blqB9Xb3BygKRXbla1qpSY0+eZduIm826LITRPn
hBjVPlQXFx5bglhoD/dgqxowPKZSUuwBTyKzYUiBwmnGye2Vl5o4pgu1zyOXs6ixYVV5gPXoLX0U
TZGvMpEERT1sZS7Bg6etdNmcLp32nl+lNfP1H9MLxuUGjAsf1DIIhG/xoGrXOXRmqeXVmcWf9hrb
jD79MbJgCnUHiY+ohue1bKvyBva19rcdyi3+zk3yAPXXoO6OVnVpvb+eNOx5uGJE+TbQQNwT3QVG
nhNqalfNIe3NAWp9Aoviueq7l2YzfIDfR0ftesQOHmE3BI+EmxxqbkhhCv1HfQ6In9Ik332YY9ej
WT55Ct/LY3/2vlvtPa3UzDleQVCS52k2SuEAj4PcFJAnrxeDBGnWdbT/tflbx3LyxEXeaoyeitSA
9QqSbcSY96idwaxu9dYGy9h8yN9NkKBABO4rtW/WwgZTBE6Nop8pds1n5ESH+MHzGxHOztscFGET
kLg/tbYcff4BJoD5J35oveC3Gd3HNKRiWRTeVzBfjjdTFrdrNOubSCzTvh+CORBeUU4FxuxF2Rlj
gj4i0fJuoiQlSsaBfTVgg9CCDWg/tWb4kof4Hh6EM+h2mLlazbv9QNb6YIpDsEypWyHaGU32AyIY
MMXom6LqsoBkFpN5pbf2Sk69HkEsaD6qNShoDAHhU/VYpUHTaMvdImV/L6GSst+YyKNxYI4XExkh
GLRel73zft1ikDvcoxT6zR+tSmNcvH/B7F8Z9Lx8pWcSo0B6XVWWhngOfDtPEj3sjgVyRONXaSC8
qws/orgLzFsyGqNSdcZN3vbjIiP2eNuss1vKwn/QEz2iKsI/OCY0ZmmAUqRE9sAA9yLsGFIpX7t9
n+kYWI4xI0m5Sn0p61WWTRgm/yLGkICPOfXfhyWOMI4SJoxInyy7gdNqRbWvhCafc1/LKsgKy7C1
MD82cNfd7sauasFb4M/qNKrC6TOw5reVToSgRWrY9teZ04q4SjqR/xJTqsJ4T4Jm2stmHcdcm7G8
SD7Gvkk1LkasDz9C9HQBRZPhrh1i1hHLIx0e9mZazQFC8wWKs8Rrim6O05gE7H6sJVQrd8cGc0gU
1lB15P5i2JcVGG83kAfpHKhfqVBzWnLp61YSUaaBgRRjEg5lgQ59cNLaPekTRfo9bnRljFn4APqt
mKT5xTWQwlaj7035ce7dtI2/2ZSEzDcmIMPV7kG5Jni/NMSCbd1LbAKnRugu6F4keRTCfE5dXDyx
OZLr7NCm3EfdUORkoFy3a0QI0BSXBjEeONGGLEPjIEEk3nwAY6IF9WqZvHKPijcilGUasRnFMb3I
hQs+rxOF4CUb9ha/+E6te/eTPR6SPRl5KvJaWjlTZxwcQ8M3ahDDwFKC7DhxRjs9Zn1dgEaURFjW
D16VLfYq6j5IBISnMVNo7RbtzwhCSCrhn8/a2rkQElPBrHmv/j1Xnwxu1qF5MVjBvszXeurwEB8P
bxKIaSQmyG4MHeuXtnx/GKvmQ1yKvri8I8TvMAwGK+ql2Sglo9doPoGbSQmYRe5N5yumMHrOA86R
3nElTz1O/NTihfH3BLe9pYqC3t9UW5s5emT6op3kiyF43me6PsjFiYBT5R4UMJ4D7JPmN1mbWs7u
MC0q7HGdAIagc2pJVxwrbxGlOeJkbzSKKfIv2YD/X/ydG3KNCGcoZ/z+L8tiHz5PGaa015Imm2xg
SUMIWj/doUfT90YOv7mz7Z00put9HS/1Y3nSj+kJeSIcwrD7jHhs7SG6t/JtYnHy9k1IGZjH+6xW
Yh/w0kVEZITIwz0fvAGPynNSYuSDNvX3cHT0fiZFkWGw/KdWEP2QRoqqXfq4bmIPVaEQDQg1vpKl
BtySNEPKTuZgXXdz41AbmoqRlDcM93VwFn/mBc3ClBhcGyUB/+V1ifFHH+srFVFIXNAEWSyDjPbn
i4hppvZzgAYr3NoUYlOGpQDsFYfdnDN5tal/4TLKzK8v/vorPvWMyphp3k/x60eYPn+fwLTbOxvh
HLWmbj2Kq8MoZBGlYk86/MkDlOTJWB74yuj10WnzL1/WAOBUWrwG5xaoVBsTSxRvuQ5QI6zvaHqY
3pLs3XB+JpK1w7FbTXj1Vm12sQ354n/HVzS5EMkCSF7TKSjidXD7DljeeXZ3UUxO5/ZniGju1sy/
GuoSpuYqd/wsYh4sevMzURMQbwsbBcjgQ/uMn3kHH2Ugx92yM5PLXFYmQNHINwzQavX324kC/xGQ
Rc62WEqWh9H4iKD/6RAkROxZ8QGBR9j+ZdZ2o6MwY8a/GSA/QF7y1o3m4a7+pqjBrgV2lRtiwZYu
F91T8G5SydFjinc3FSg0/6xeAmk6cFnXOlUSmJND3wUQ+Eo76/UJE0/RyZp0WTpWlIU9m71cHCdm
A5iVK8/vyT9Fs1UEawRpbh8iUS/sWIyI9IA6CzgnSjxQu2EFeCBGOjV9WorH9EEK9pEoFmSRoe4i
6CHUnlj5ApwiXC3DQtV55GSlNC74Pzvl34sazrG46zv1RFyAzRoLC/w3AGB2z8O/1EeQLPx+yhFu
BKI7R3ghclmInAJmoI6759rtfVL3oo7TBB0naq9hAgt1zCUSkZI/gHoCiip0C6IiwBXQnmEpeKVD
jt5ydkdcTJMgVzH5s6yYFchr2pYbZGxwNjgilh7SOErbGHSNNN0LRcbBy9M/7M7hfj74gABOFUOt
0V5fyTtN0qoIn3r0GvbzTcTxBKdTRXZZzpuK7H8Gj7Ue07bIOqAdjkNQJ9CCBielIPiqKkV56SqK
8MBw8RXRNp4OFgDTtouE/j+cYNvJdrFkua++r8LMCEqrAzQBH8aCer3C/GQEHT20VRgLcjYLC04T
Df4BU2hszbkP1fGbDB/D2endbvai+oQ9PRcUERgmVz9ACcNpWDqPj0JLAtHJTnxmn6HgVnz3HNjU
n4nDZm76cublaVLr29Is9cjjEcMHb8Tb+hR1/xcmzU1a1wy2YQUsGXspQBSpHrfPdhUcKCLoZxQB
DRpyXVtVr80jtsfjm4nHjrKSpV8W4wT+b8YYrkEds/Zpyd4G2x1nT4pXE1TmZWqWLqiwPPNnG7e8
QBterzAd4J4SgJNFG2/+qW5AvXWNdIc9DGR0l/XqzlzjDlsbs12sx5IoG19Bh8Aydgn4OjEH5mJ4
4U8RcmTLYjCMfAkhn7P62YnTOpdqXy1FTCprveSF6Z9Weh+Xnj/e0G9UdNuMcBiuo+d04N4D2+w4
khYf5G/nU9z/EhGcMVsD1RnmGCbgRipZCkn4lcZOUC5pq629ffrnTK5t1oBrCivb6meoe9NAYPTc
cTTtpKrB7JwyMkPuvHBaCdGUD/7am5RWbGyWkaE8sXQES4d6AFQemm60QPASa7h8atlgGOCQQrPx
myMpmdX6Ej0qwqFrAMtHJxQv+Q7OZRd0GE9a5rSt15FDCMe9UczweE9enkqTTTPwXSzkuIIi9z3J
YF82J3l94Fv3fdc0X0cLPE8PJcR0uT1e+lBgOz6bEHjjN7ZlpW+Zq5RKVbGEW1AVO67CKUtP/yGc
/R2bttCv3Is7rpBqQwoUx9SKVEwN3cKuydG4CieJihSwyKj4ZgFrx1adGBTeEw3g1za/DiHr7ZUD
/nVxehZMxcPGeTYWhROU7gvKJJdnlMXPaoNfrLLexX4uELLD7Gj7Y3jijBziXMHVIP5K1gSB6BU+
viZFq+7RvKJWUTT1TzBJZnjHYI7IEt8LrJKy41K7aoNNGwBQwdRdyBnGtN6FII5OuFHESN4wnl0j
kK7nqmmqgY1WaTtj06sojs7DDRbhTAx2Xwc6i6CVPTcXR9aqea5XzRNxh6XliKkmJ6EdeP7rZZbS
mcc8W007OgU0MAlRHg9YAwnFBHX+NBk/4eXQwd2I1BT1wGD10nm/WqiiIenvgugoTc0rBs6nmCE/
P2syU8PN1KaM9lv08DFH6BEHKuWw4BWT7ydSfMNURyiyduWCTLjQBlzmTgxBqYvFZIbloZ2Yc5Gp
+Jjyjyl5MSkhTYd4ekn3ZYQajPTqK1zm2cPLP7NoKMaNbl1Ft6hVj3jptdb5v0fKTQXRzwDJjOs+
JXTuPetUEmGKkAlBbk75zvkcHDViorh+uJomPe4P78zclPOEnQ7cfFCP+rB+yZ4+2S/1Xkd0mP/2
LWLNZmc9zbOpIBO4AdEAS+zy5nmRe2Nh93YUHrVNCDFzk0lfzrM/Ja2z63t1mktPVdvQIIoni64G
ch3cPj1R/PSDzs5BQAG2j63sb1nneC479MSwRN0s4RWJn/9cBcbqapPxChwvhBgC2jRFpcDyUm8X
sqgvFbEAfNhCrqfP/D9ukfXzc/aE+SiW+ilvNaZ0J+ajptAfZnjGL/VyDthRFC78q8v/MPFzY0q6
as+ff4UWVt4+xQkGnUTBEx+6j/vUi7tQx8mKZzc7HRcJweGkb8uhomUkvZLedP/z/x+enogflHuR
ZbSm2aSJDPh2DjmDStQ8vdf2jSDSqFltB3Ejd6jJdK0Ign5B1faUnpoR1PO//kjpJsCCvZioUx3N
AzPxVvwM+KBQkjL//Zyzgdh3I9RvKJI573XqgxAYUjWZ3QwZdgdo1ftKNNAVtz3/3QIY4LGQd9MR
/f3LfFrgGzZkuv8AXwKkOaNY385BCONjTzAQ8/heUCYVy7hkJXvNwi+rQ7syXIRMsWleZxdYz+Sc
/zQ/3JLHO56nWSdxkEv2fFoFSRCu10DZ3QsrUYTegXhmhkQUTO1CtRdzy9lIDoe7P7ozsGtrwpzm
z8kup01vnJj0HuGh0IVPWS0HCCyDQFiQj9Y2Mw3ESpEg/7TjO/dZKeLsVFGlrhn4Q79vkt0XPDba
LlnkQr/c10NIV98PPhpatbFmlYGbvpgtrOqkeqs9utY7IJRtzypyBA2oX37jHSrL88x7GayF6zBq
vVygbr8vYmvXINEq29jxZlW03rzH6Nj6bg5qu6Osiu3nzHy62TvWXal+2oN5vR1jPHzYLdeP3bAj
tOxPO3fE64LUDv/CCv99/DVzohu3+ns3dgX94xQlDXc3ch8hUziK+OrrG0aR1EtUzWnR12B9VazV
ensRTJlAVdkuXoqYu+1PWS6c6nNF4V6RunueungcQ3LqAn50lqGbWTfJcqqojmcxEvEHQggyQwYL
mzL7DNscrpJsyqhmM7Wz4cNWR6SMg0UA94QsEk1SWuX7kqWSbS57+MDNSIeyPp6Sck5GZaYl1Dfq
ZHl4FXJ6gGzocClpFHuBVLm/WspmiDLjGfxdV51+GzSXNRQmE3ed44imxpxq99YBEHgDpxvMGEER
6nvfxHm/G3kVTx9jxkpsb7a+RUvG4p8mE2lYBJfCbvZsAIaaeBZ6Itf96Or2GizBo9SRX9CSWMvi
8pdBUNn0ashot0bkPyRH09PUb/as73SzItKHQPv1kiP9vkNAIIXREIpuRli15W2fckY2yEErMc7T
mNFXLhBpK5VdXJo8bLritnG/pc7qcqPtJKx/4AXWODQSU2vcEER0hdWoEeh93c2WVn8WrYUV/3th
mpZ+44qhwqfo/SQBYDnoe2qjbJd0xR3LdADGYqB2izSHJhXr0kmO9Z26tj+yjnKYf6daRrNlMXiH
SUX1E3GPsqerqIkYp8r08HyJXTcD9qzFqwF9qclAyUdd1XO0O7+saOL5tEGKeDAylsG8doO1J2yc
wAr1pkrJDtt76j/tC4ZQ8ovk44bQrKQH7sUwqmmxcGudVb+1cA13H35v1wEULYAHE8XoJbQ9JLAz
ZeEQgHaPdqs6qD4/HYLTau+zaleSlyisHipYdVvnon/suGyJegkUUMjY/Izx6DizBF61wdmdNsGX
KEOCF4e0dqmTbJEPDR16h0cvwXu6+zD7YG2blZDNLNVRPqMM7qABO7lkxaxLixhukUuJyfNic/VC
tGjuX3Ds3rAa+F22ZmVG2AB+zCU2hDvx0HFxtM/7jBH5Q/Un/I4Nk83zoGT0RldEB+5+8rZIJT0X
eZ2bRUZTDAqPoApckLeNN1aCdYfiog5tDGv4/fzJjmpr/jMODjEX7C6/7RBZevXILJi5NiwLWQGy
fIcqUmJKFL+Lt9KmMbVsVvI2Q9BpQODUgck6IePuQWmft88H55z60hNvD7UcNag91EnJVN20SdE7
KlLeZH6KlPX9ZRWyofR/R+e30TUSswYImduMAZcG6SGe8CjV4e0MxXRbQO+fRLQ/MiCQBa2h29Jj
iBnOzlP+UmG16/yHOAExIyoAGT7F+o9LPFjndQ431le9vbs3MPB9GWJlheTiMq5L29/wMx/aa4GS
sdH1SjIuhZywGwjkDErALBvGo6xMmqn6AqU0SHa1Y+sTVy8+pXGb6GzgCcgvvWHIDmkcedpN9HIp
q0qy8wHqL2rVifPydFyYXYa9TII0bVbXgmWOveXkqE/AmaKGMfH1l0o4mxcsKQgiOf2cmSrpX9zR
FW8LaMNQxyyou//EDsUfEKIIS7nfniY0vMVpp6MJKUjfUK0EBqkuyYNDSxtsLwrXAbFDkm47RcaI
vaJ682obfbg8ffetAjUypFSX18vx9QzQalHPDpLbB6w3eUT9AzRBLyoAnp4kV3SduygT8CkO3uY6
f77n696olezCyk+HPCfSXf0+TTj5A7lLK1mJ8MIox9fQxABr/9BDvdNQr9EcVe6f/GCGYA84vm5e
fuseLt8h9tsva/Xjh7XJlpNtKbkxBNq+6+AyMUv11ANdv79eCNNYITt6o0Ilrt30hqHj4a3FP8Hr
RXLyvskJrfdCi7/Cie4YADBwnIc8m/5BcpxcFv/2W3t1UxpxoTeolqMha4WjHD65GH0zQbt1uhYw
FV5zF62lLt61q6MJbvm4kRIWI3jBDpnllcOU5N5OgtCwiFeNrTuzm48ZB7bZ9ctelZE6LzfN9neK
aoPIYNV5XWq1fJ/E+VOHeas/Y4gv9q0a00Mj8OxUXxiAl9fbbgbc3qadVIwpbqgURzWBpmgyHY8p
5PlCvH47qHnLdzL0aOEiowjlNuWkHf7AUhhynmqID7kxlRF2+I9tAHQwA+wUD5ag/iv1Uf3VsgJO
BpkMNhCW8NfeEq8fHY74VFNX9w3g1tFbg663bOAFPsW+FtWFZ0znpGV2HWulR+a9P6rLKlBGnLJi
FWcRZqyUN0r6+lYeAbJuXChc9O5Cr5WXkxCh5aOOU8MOihGBp2qns8yEpsyXmcBoAqD70uQQfJwd
ZVt9Y+Z9Xk1+Lgy4crbBqkBQSRcC/C38vjRII3nFjvLIZqM7erBgQqsQ7l1ITVwy3MPTl0+8nTOB
OYDDWPPKZ7IeomOFmY8IYHM8sQ8ZMWBS2n7ann2cjEbG3rzbzucsp4Nvqnpo2fHrn+3GCcaLMOt8
hhRmL6fUpcMqsHuKl+uCFcrhjQArdBct58ik8m4Lkz4BQRsfAnEyOSgw1ocfEPEtwIioRuw0PC2H
PJcCI0N8GDdgs+eOUc8r2oawv9uJeoFDpppcJbnpbyZLy3WoNFFxNv+SXxeZWg6PDSj+Uw9LhIbD
oZxIm2lAFG1YYRLw+ueAgHclGD2jFAExDi3bqy9kbxAa2vmZRW5PXYyQI7iBqwe5+aQGUFJQvNeD
r+Pjs1aWc6Wrtiy/y5hzP5y7a6pZ6e0HX/9QC6OYRR4Hv5FOg/D3J5yXPyuYiJa9CFm2vZthC7uO
GvRsstY46QkH3hwkNDKUT6qnJJVFcPN9payouXocxE0Jz260noxEnUDtXxhKcGhxqXmR5kcU1yw8
ktGrrmeyAk5UAVnkgW1yNdU2p6swiHtDtuvlNTfVaoL43lUSAlId3bbpH4zK2XXo+vMYKgIF9dCH
8fMnteLjrRr4Rp9qFNmEYNjTVCjgzfiXGAiqLYjG0iw4SeYqs5ncrJyfkO+4AS3lXUcOFk6h0G4x
AZuRRCIzA4RPIKLh6yIigPiM2tFuy+zg99D0GtD6tr48LcFgswpI//HAxktpRGd5HeNIMoaeKoE4
nNMr3BRPJDyiluPp4/3dm0Gp7IFK5aShz+kgNFZ6N5X/LmnH0Yl9vltsSMYYmN/vTY62xEF+v3YF
rjTsO4FmqDiuRZYE8FG/gsoK7rSArP5cPkilSlZIL8w8S5qAP1DlFe3Y4ZaZ5CVcPsHqGfF8TYTm
BxQ+mgq3A5CJUOcyGOm8D039A0oz4u35alOXI+LzXDbIUJa79Fj32VnqVcecLZgVbD1S7vTxaWDl
7Q1UwYBoBm6kJqyFHrEgKznuMGTu5REalIFrlsbGhiAhqWomIBpYw/Ae0UC8MXFOYx8hyWw4/u6k
hl3P0xDTAOoXIbd4HAm2Nh2zMXZD88pyqxYt9bM3Ctb6Fo39h7/KeUtGDEGkrpTXtflYR+pt/SFw
65beyuYRdE/fCIu9JfsAaZLqtvrCk6a3tXxjscv73OrPh61WZsWVPeW0N87db1a2SHQyFx7FQzo5
VpbpDnc/SU45glzWZs/DwKZ3tGvhnnOSF5AadJwN/dUsCv5BeMAxseJ0DSzyu6DcOX7lOd4oy/mW
Q/TwX4/xz6AvcxMaNgsGhTX5LUCfGcJ96ZGh5QLXfxn6h0660M1jXYlu1vdCeZsQp4aAalDINLRJ
IU+6/qH/Fn3uKkXcwb0qObCynrcdZyjNB0iqwx5Dli2v+8HLXwmeHvBt/LkCTijDDyQiHubcFVmd
7kiuJvBTtXWKycmuY8cVqXp9+YeC10NEnBvWPzer27DURqOydp1gAoHjoV8BenTqxVbsjNU7R0T9
RvpOawJzemINdJOEJVvaqa6AT4sxVGZa9ZIL9Pig4ZR47oyO//HtNIR4iHW9TzpwvdConzjDCCPt
GqlFEr688DsA7cT2aYtqsm4RsBllxS1neEbj/yXozJP300ESQvWFnjUOKG7Dlo82S7OosDe+FPmc
pMsbh2xeA5cFZlEENiQ8hvnqmWZ2XzDo0m7nBhZ3whhhnbDp64zdSFTW0iRl27PqIr/WE6mHOumM
Q3BNe8nJRCoz8Gq9EaMXTp0DDbkxtVwBYX65EafHf37nXOsaz5J7RF8C3qbtP4VF0uHd6UELzi60
pq/TXmSqZSfr48jC5pnhMCJe4i91QAUlTylVM4UXWYhNIuNzcb+/8ZQY5SaGG64PSKvIdTW8/ydj
e+f4abTUyqSFuvXtIDASRxIopqVoBK+bOV4GG15OCVdu8rf7V9uA0lfF8z73OTeU6ebjpNR5PamZ
Fi+YjM/3ouKY1iRA49DMx2QrswDXWPdJI66ssP/rrlLzx7Hs31eoM5gZJJsMKGGoIUAyRzMQNSEr
TxeNX53KjFe42T+fxcJXKpe7XYSrzVhik80Kj6tekJn8Ui+YQzgvY3MUPy7oURWFPgybTxx1z3GS
F1SeICdcRE4n/B/VdhbA6Gut1Hip3e5RIetok0EpyE1rdswTXaaTfC9XOiKj+M7aQR8APvzGW1be
eSLAVr59Ve6YwkfgJsLfIiECxtGnUOyh9WJpQnRwSHQOf6ZWVnzZlcFlHlS+lIRVxpXVj/BCV/t5
Y/eILlPPQaTp1U+DoNX1T2HVoUdlHXE4vGyYJIYo008Jxt0/WNEVpUJ1ZMHxUgh8x+Zz6qo5zqm8
E1ct4RipiiFq3H6xHaHX7JL8cOzc59t/lgYnFYTMRioqdNHJWSeVmcwmPsfWhDGN3L30j/PWQOXH
4Ba83Fqt8DJew4kEwDwyx5GzA9lTZPFK5zIEIH00ZP3IFEvKjdOoOGTfxUX/BJjf1lDpa9dj3il8
iCnpSjGmQWabuceiVIIbNXNk9Oj7JKFb50QWm9WNPo/9yZi9IuKO4ArnJVYyS1nqmVK4VXkmDgbq
ASltPMgWpmM7pihD2uNde0bpeMa6ggnwFcUBY8gZ477Zf4OB0WlKHowVMB8QP0Lz7FLaInokXa2b
xU7ByVXcceweIefcB1vqJSh2iCExzh7NVixj4Q4jiYLOiuzjxNaUGOjdY5gABF0gLttJfIr1PIeM
l41q8y/NOsV5Hq6TmdOiLWtrgho8/p9o7vzVR7ImQAqCxl9/1OgY71KtmfM3/vLOvMA7NT/fP/9F
HNxXKIZiniwe/trN+8FiAbrPqnI8Nza1zidBRTilrQLuBjpIajjgSkolRyR1pT4mLQhfrqZx3mdf
++FzQdIgl9yiQY0AkylTs3GH/lMK4YtJ24RCKFliKCHHxRvgzuJNjfxoeBqeTNAcM6eXEdOvHOv9
jTqYy4E5qi53NMmqwDB3KbPuw5JshLJi7w7uLLNLUjt9UKC33AmELx8awKxRmkjbmVDeTKkYVAq5
wiCbjeduYpWyufqEj1QO3vnkegOty8iuN+DHG8wIRv2GTInb7+g/iuqx6pmSTd4w3dgjLlgtwhL0
Xg4nUKOPRtvrPAdXHME2e95uPkehgfkUCE5d4w7oG+USAIIkcnTEfQJ5y1Jnt+G2azxguOpQbONH
NVbOiwj9oOz00LYxoNn4//MQmC30mJHbA7JN+UuF8Lxjn259zDlPaP8rp06k4KSBQ1I5BWstf1Td
OLLefTRLbK3q+JsxY6OGyNQjae3wqFqt1xpYAH1dfNv7/ztm1Kp/jOLL/G3KXsEBlzkaG617o5dg
ngRrHWzstWksDMkDaDK6DuaWCELiLqLWWZ8u6RgZkNOu+oeR5D/5Xn+4KEo7zszGBCwxuzDIxVjx
bWjOlUYfVBDsKxoF8CA5U336GHcJdut+/nIU+i8pyZuVcQChxYOtyjAz4GOTuKxOq6e+sBMFj3II
Pv6uVyZmpT0NbknyCz/L60LN2kIaAk+MmEp/V++Eu6nsiH3+EgveqiVnoIhmo6P/+qVZs1qa8NKP
0sOKzTD3hNaM2JVWcaGZD4LsbwcWAamp3C/j7nGQ8Gzsc2Rvv8skfcHrDZpeip0vOfitefzIz6To
t3LctUE5USnBWDKgBndfHfW/CbQEMhwFEE0hIchkhUB1GxVdUgOd6b7Jk8HFtqlkEph3AQfW6hID
SC3sfdpvP6f6tRvOkntZSXOqyPBt9P6EBYiBCBv/u/6EEMZzMVXIrETpxPPpeHXgBu1niCeBa74A
dY9/d5Jz6jbXOqmwuBYafYUik0RF54TIFlEMXe4x5BbME5K++42tKYhQRwIgvK0Ftt3ruMhM1n6O
g9CIb0+vFYrIttTthnxtDt9Uq2DMJ5kIqOHIu/qMwgEdTJCqfOCOhscJRYLqJpS4LOJEmQdXtF7X
Rc2zoGr2PEbR7vJpSfryWFhHQuDMCdm1b/WBThpzj0Cfn4zum9gYyBuEwT+7oLkLmxpRSBMhL4co
TbN71qgpZNfg+vFFapwN8TQNaD/UP1INdB20UbRLHecIFh+lQMzwS2UyojrwCP40sKRXP10xj1q5
9GqSbDfvCPvY656z7cw9gffYuNMo50SPilCmEd0INcJmfqxWncaENneq23lmOH6Lur0Eg9ZY10FU
cRWvMw2CkU67Lda5b5E8TcJ66VZF3kTAvBP6NTIFxf0xU8CAwuqmGx+uNyfAygWfARW2+20WuAxO
sroeQsAGzTp0HYWO1A6ZQEtFIPXgORHthNUb9CT7eSKUejLqni/KOyvUKJqw0rZpCn5EOiwXZdGu
fAHZpFLy4rLAjCdHKIBhyi2MMc5lvoQCCH9mVRXEtkNdifX1jhOLko1OLVgMMPSvnsCW7Q9rj4TC
xQaYW5092rp2sUwL1oKiXGo397Pm3SCalQan9U7UFbCko7+N2iU3gCrZqZR6zJmv4ax5HNAmbGJv
K5N3LrJQeB0K+uFtHe4JeNFaYnhAzbl0sVqRlHr9yW7dnHRMqbryla+XnXRChzyLcyt8RS9em2dm
tiTUsStq8ifNAF9b6oz2q9+H2XdHmDhPKucs/A+lsmc+NAx0nVblPhKSgmMnZj6HJ6st1kh7Y7fd
fYaiYFV3yaxGVkyYQ2H8sSfwx4ZkUoeg97Zplp7kc3DQymb43FpLrg0yC1IceN4YycOoAsQfaof5
DdWEarDNEToNiq+bY6/a6nlrMLbImFXnO9rzQ+bxR0b8Zzsf7Q+9f0ZTpRX9rzeVyzTSBzdhMzNd
vANt3KmzuqKrLmvSBEEMk+IaaDGdctq5216zgxmvRevS+JscIujbjHAR1vt+dR+Kb4MrY0tkBGIq
cG/v57kMb7KXZFC8NXg5Uy5gtPeN/Jd53rqrvk52eE0v9sQIN6LZnEmFH0xjQT/FWgn9BZtnZvIo
+LF7HCHGWQn45SIJ34IPn00dJf2EzmTDoj2SNiYo61xaWEM+x1w60wtcf7fv08YaG6KwngiP0jZh
Rg1WOC7c10k6cFfZlzwekkeCs7uoTDscXuMigybuYKOVVNQLO/hS91gJq0lM5lPgLmh+MJC2Q4M8
7QRUnsLzIC6RVkSbyYuDVUO83dkINxxShnwiscM54672VbNqHUab1av2RTuKTH1pd2Uo51szx5zy
nIaseuMGlKtj7jAr0xSfGEFrISUUOrhY+ZYEwz3bKfzLez9mOZxtfWF1XgWR7sXDIIOYIaHCXOQ2
2MVMiwnh4AwPNpa/5x2UYNcLapbs/pFajSVLXQe4HJQWq3V/iFW/PKOyzxWT8ZIJUARryIvVcqxw
iguWNWIk0YCO5f+DbpUGoC8lKlkrtLaiLEK+w8KEbrtOk++cDOP88+iYUx3RzqG1YN/mKrOMAiLV
gxEBXkqhrkwbb01F+aTKlpyMpUsFT552Nid9sPDFElHOMM7OZosfoPc1plw9MOILvyBT3Ke2VdL+
8qYtarac94XT4JVuuaHxwjvOWK+RDmO4giFg/wbh0qkt5A1osXGIxnVevdS+0QRQOiQiuz2sKKDN
ALNK5eWT6OvmJmOMhZePndNjEkR+pSoK5SCILm0Bl1m6fZvsHoZx1A/m+n1mJ9bGt80tYLzr19KU
oNh4BUl5AAMLGPGojOsiIzJJrTB3sdyl1zx2XGloBLnid0unT1pKjBxnjVo1uzjaJUpL6WuxWRVw
HNagbw/GmT66CsUFVcNvSKp/FA7tWkpdxk2Zv5cQEwAjIV0D6IMaZ1yMjIqb2ZS9YGhGi3dzSyho
OyZBKp4UlbeZ5J7s0RHIufxxfB6CnFpiO+HdzlQxvu3sXiDEc+YwcXOlNCUzChogpl+MHU81DujP
K9EW0HJUbOlYOFK7gmFJFNXPxhAynCaudEGKgyhDAwWJ93Sd3PJvXzxfs57SO+8KTw+/grI2GrCT
+0d2vRg0Pl19NypMDq2Cu8Y+PLRVBF4PyDBxeMHDDcjzrp8nAxmt0ipU6av63TrX3zXIePoExC4W
Bo1ebakiZB5F7GwBpNocYbPirCJdjQL0T5gOwphwg/hoDmPByalZUkxnTzDL8X+IRnRDySL9kKUM
7IK7WwtKX9W5d1Basm+sdSrb03e558iWIaQ0QZudAfjwPiCKhEqydIyOvTH0qGy8MjKXbdGCzy49
Gn/6hz25V85UWlbBFT6Bi/xsyRySkn7n2NAmSxMhRRThmIET+G0GOI3nAvia87ZVRmm5mWFhkEKn
J2viMjMPGwz1/4IFLul6jMZzRlFSCXofmuXyeLyW90q+gOgm6bCamXt4xYekd3D/aE0HpOZ0vLDf
DTMnt6tJYPX40lymmpGK95H9KvfyZz62rwxeDeQ15H2ZCXJFpkxLns1MAPpcDmxPXB2d8rhosNI1
PW74GFZNMc/lWY2diD1/IJ4rJ7ySmP3UVxeAlK5t9y8XFAsF1SDw/DzBhJB3oO0Y2bgfzpXOPxHx
HoTbnNFl0CdAbXZelosmqWRZB8Ypht15n+92aKNkmDkBz8vkPmfflhM4/SL05RM6BlDCFpLjK7IU
VasltxmRk47/7oip/UYUK5/U6RwICsGqyaS/XPzI+jVdM2peTvGorfIAtwbMgJWFNZAepg+KbLf5
0tmpLiUt4yrGOyCdXEbb7cuZPBmvoai05ZR3/W5wx2TvvEU9XXPfQjKF++/7e/s3yDgQvnZwkE+A
tS15f7KlX0g9kUZKZjIxdxkA1Wq8VMU0xyof9T+ii0+N933i9iZjOrfpyrtJG3QcGg2Jiraslzpv
REJhzJ6i/f+00UQMUbleEr6SV62W9juyDgrb4ArsTBJQf2P2zn4yoyG5JeF1aC/5AIYBzOcZZKtH
8+urOXtBPPRfzX2sb/XpdG7YyCGLNhycOEasEDsRsu9qIwdAWRfzP6mCt4p26n5JWtnPHvEil06S
4nfZEocRJIiMPqC6VzJrjjxD7ikdaMdBZb33q8HyChfNFxyghBySrKeR/QziL0vzHeZvaho848Ly
HHPh01cALX407f6NeeCKV9aKfvAzNfIrvHkHB02Mk8xsHOySCzWHYGh59QNAkbAWzE7pZqWMMbpK
hSjInC50lxrcgkfsbF0GlLBJRCpPykdGVB9wy0EKd4F1SFTS/MZ2u2GrDBRPgsdej3oFg3A/Z+AQ
Zj68JuVoRdNE4HlxvHwoqmqmbjV92wpkV4tGGPUIxADG9y78chJWOt+FE9dlI/Sp6D2ZK0s9hLlx
sVTcTrl2Sxf/6UPTJyHCV1N8H06HIyfoIeG3NYbFdy0lu98OdI0eP4SmxumvoKIafBFD3czgSdsU
aBlQ/2/QEHglA0lUtI2kmy60uIVEFODHlVX+411LX27JHmta4ayKTzCwn4uFKqpcnk6NTNPNsZ5R
OV7aYvxDrlYR7PRGUSqraFVB/CHeaPc6nj25SNt/mBDphEhxXsaSSJe3mHW2Xc9HUDWb0jcN+bbL
w6cuv7DFO7qbUOfpD+ni9fkXLzi2XRtKZnlIN8N8vW0BN9FDA7l6RSs14DhPgHRYjTEdvNecMoZv
uVQbzdwfuUuMeqzSyX08DFdUsYhFJrzoPNAyhrhsYanloNHSbssbB46pKKf2782X5GefBGslGHZk
gVNc+hEgm2u71CVcAeT7M6WUljr9yhP0eDIIy8Rxe1YJdZLHGHepfNrQHmyhHPND0xPt4ngnrvs3
jDnZITI9Q52K796JY/P5kV42dOslN1iS0JK6vrMM4lbcVdeEUE6s4OXDLXSp3B2Cii8n9ndSSPYn
wPGo5dDKY+EMZ6nrbJB9RLfJ66j1Dvsl772yTREXgQ/zqV4FblSESOTaS4ZAJrHoP2oCPZzQ9kr2
rID09wrbgomVY6klMzLdx2YIB16kURhV+jjVwK0FZCQvXfoHXsrwYPXjSS65L8K2nSkG1RWi8N78
nGjp8m12BY5S++wbyEhaIXe8/zQWkbQDCWQ3c1QVznO4Wak5oFO19NKrZfk+c0K4QYblV3V1GG/f
mqRG2iPVOLX6/M+OrbPgF3xo48C39+ljYBmaa2evLbPstR0bq18OEmY/zlO/fUO5mTWoYmnfArMb
iprJ4fL1EljDzkKlzFM290gfPFSr4TV8Wzs5E/PWLVnMsRaQdRZwhIxwgWs1uTy7lvU/B5mBnTEt
qiM9GxJPKs3xbCHyQofNmhtThBhC/Fpo/xRCJl1UDeN84DYL6R0NDHF7u3aTZfrivNR5Iv8UFKnQ
mzenCliKxw2oQbeFE+oE6w+DGAKJnofn9O/aKP+A12snw3NZL2dYzM9aEJPZ34X4oQQjIzGvLqEZ
Or+ZsPQYXiLVSUQ1fmDfhCPOMWTVLN92McmkIQ3PrXFgh0U2J7TV7dDqmu2bQRqvrXb8EQq+dDeD
1SWexOjAQcztqOu4hiRK1obScqd3iVrmrvXn43s6EzjbYeezE4NKJElyPFP/QmfC+OcdkbxfZche
5e47A+NyFirr8UbYAIVujQ0DpY96NDD318fmZ09HOsZduoli2Eg/n3o/V7en9gYdkj25Idl0ipw+
jpA67FPu9L+um6tYI+IyXW1JHqHWkuBYs2RGaXu17+chi2KTjc+0zzg6tjgVEQdIFGXrGlgaOu/e
Xu0kpRaQhIbdbuKfxZoxPmo9Op5jjcsjpQvlUx6Km7ilfE1vrm0p6+e0ulZ/Tccz0FdVpoGCNwdx
HYppx7N83iz0YahTn1hpqmukoW0fIVbDirKe0Gi8xgA6XajeIF7O32WeDUi/fqmkoZv+J87Fzd5m
76PqsA0Z/pIMrRuyEWTfe53o9IKGu7eIyRibMdHoif96/iShUZJOjLwblPPKBdGpzW7chQTdcsj7
PGXo5BCzfgHYMJdsva26ZdFTqYLHlSiRVY3Wc6KZQGIxdDfCo1LFQ4ay3X2Zt8zgXx8tdWy+nhh9
SeBY3qPlx7BBAQuIfHLKZZQiSOZIu69bJdmyNgy+skV23jRAeDxL101wT9XPVLLSLjWSJfToSRjD
hOMcQ8z1JZLpcife5POJGCH+aqEsxJyjF7FwEf1gM3JJABXu8z8paQUNvXq4ZntUhCbmaxI4iaMS
ML+tGy95d92hIJxDUrMgIR6PBoPKf8Dg2fqRBj2B4gViYet/l6EgqNEqC4duKAONB+79tk4eybmb
Q7HVUnQgIf9nTsHVUPJAT7N0Cuhwd79ie7lsqZajtrk9BI5X0OnP3zBosvoOMY3vzsGqNp6kxdh4
/vSSHtfH/yDtoAVtKUHse+asAnQr5GAihyElYboxFYVGXLsDWicMxEDSdC9JKhjiJ6wQ/I7XHlOY
LvVqHpQf2VJTCwuRIchJ+LccB6CTGCXZNgiibCyGR9AkMXMO/ka0knYKPgm5GSMX5XVK8Ly5c82X
IqjJEZBOgRcbD/stfDEN3NTKiBRgy+aTZkt3iDiYpLlQ1rcvdXAN3/PPsv+SiUDHLxUen+g7xGnJ
e+BVwxatY+RG5ARzLyB9ItajKNnfqY4sVWWS7/M41WRcYWT+9HQc8jEnEPiL3JbEiWg4aIRyCC3m
+abkAwN00+1lHxtNGfRGWv3QSu0E+ss1hMM8THbl4V0g4BD6Dswy2e9LHKSnzLzendOuCe1Yr8Rw
s0RSPW5ZcRML9dnLIDcr2nlXtmxUvD8khwsKEwKlUWugmLPkepLB5CNKVhoTlrjQnCd4JVFGtDnC
qGiuQyWveRNXu7aVve0Lt4xxfvJamOyZfaE14JvO9iVBJisbPpc7ruIvya8qGWy9vsm006Gu7eu6
tQmt1NRKtjsZbRioDmcAH+LzOXOfAnSfkHp5QewQTkGVPWq2fl05GJMrexzK30pPkJ6cBWhGeuwk
+NphTewwhRmhiVYY58uTqpJ5Nas8CilLQ1JC8AzeCeA89BRkMWIukvRHGQvHOd3n/rdcgYEjC+P7
vYJTK7VC5cnxH1UYn4YDkYnLZKYEdZQ2SDL8E6B3TMvaDAYUoMcZ/xH3WrSZIp1ZFJpnbabNjEPR
Mvl+CO5FbDPh0sudC5LnqKOKKQv8tQnTwLYPQjbxgS+L2ov3tKXaj9TdjcEI8D82zGfxQEIxAzA2
WGEg44hCi9P+M3BShlStcjrOzNHhiQtc2M77Bz2I9BRWQYxPz2jXXGfyYt1ct0JHXs+6azeZDHwK
YAm9KRXZtRmz8+Njmd0Y7mIQYYRft02ooOlOzZUbO2svjcoArYW4uyGnIlV5+vP5s9lXNDwoPhKn
WCegUhLJVYM4BbUBt/l/86b1aWz4pL30//SymrpQ+KCooOqTkLnr6C6MsLtnHMb6JzVd6mmT5a/c
q142rWTNvgj3sT/tygAf0jqM9ciu/EEJqZGUndQau4BVAqcTd/XsZAO8vR4SnHmA1mhbA1okuUC5
T4oHsjfcUgvnWLpzI78GJnCP7YvCpzW1I3639oja3t2h/2Bydx8YaN54vZvURIVDBNivPSEIDv+z
/DwBCSWB7MRU2t9aJ308h1gIaEJ6T3lL9KMtbEBUdikngje/icSReeITz39YLiESU5YLrCkayt9m
PLOcKaEBHUnNu3Mzt+KnrdDmITfLYAUspgVL+SpewZbi6gB8TRgb0xD1vioJ4VoE2JldzGzM3Khr
qJYEN2ZV4iALpFMp6kzDIygxN5V67BSV6p6q6nRVCj/AtLDoXedxhteY6zI/V7JNUgdFCt111qbn
8tjR2l4yZ/bbX8OaERUVhjkGHVzIkmj6zAOmV60YigLae0JebbleOGwT/g/tBi7wf/HTx8gM0FE5
5eN9wcmbZyP8h5eiTQ47zz7OXHW0nyutAWvU9hx5gWNdF4KhmBl2ueWDebp7s8Y5VZg/r3d0MU9k
EXU30d39NPaPEPLB8e3huBiSCFHJ91V2qhEHvl/U1HXpdcxyiKxPrnvVt+Xy49rmmlnlsYOSV6Hw
Tn0PtTJvGUAfLGFhRvfp8JFk91LfVGUjzZJkuFFXfuCwj2FR1vQiCd8xUl/ztY7ia4+3mn7rmDTZ
sYn0rmvCAv80vPu+Mt9u4CfKioYN1+NNgUm1cYP7C4RRdpsRCzws/SxFydvMrFfZbJ7gIX/uMq8/
UXoqCAnh2Ao/RKY018/05q1LDRueR2XU/xD3/l6feU+b5telO8OGAJwi++ouN5Y5tNCtYDrI0BA3
vZn49NqOaI4lUPcHM8TxvigHvT80Dt2/1UMemRToFSJ9C5TWQpNT3iijji+/wRxa3CABK6fJJiZX
nvnOSgf//ooQnBLEz0TEadSWEzwPM8YDA9tR5/v+XcgiTG5j/u1QAnxRs4dqfGwVQiqw0nb0naIS
npzRLxBGeq4VUaiHt1Ffe2YlTGKI9ddQIW4oyR6ZLOD73Fthg484pUX08PYK25WSCRXzhdsOobwX
vTdGqbwucXAB+lfqNTFnlkMkPSw+GlFAMvyKj0b+cOJevd16OkJHzVRKAZAPqU/9IssQVOT+D4Of
wnTVbeDWTMXJhCOqXWuoq0bof5yqylRyWQ3JmrlpxedvKu5gnVHq5tqN+LuBo61qJiPQsRvJoEtJ
xbjBRQzLdO7Zq13cvx3HvjyGjLjssSO8oTQRdZcbu6fsKSi7RQbBMKG78LBPl8/hNHzU5BZMk4il
yEKp4rt2CJmba2W+8/t7m5Yd8w4zDRaeoj8Gz20sloxf/t4haaPvr2S52GSuW+HZM8bXK696QFsk
NR5JnYtpoMTStHmOigljD7YxvsxrbZCcNQ1qBFmv3T7WO4a43wSULy90W+vBUr7M1E1/fA3jfGjv
yJsnYhC2UYb6vl+JkPvk5WuhaWlOTXHcrgQgUUow5nh6TfIojHIZg3ErdJWKJAVBI1Rus8uJdKPN
7hKWpJSeRGhVRgvKe+8zPqzBafRwekraGEFZbW6SDUiHeqIvASiE5i2IUX6TkMOvPQNj66uy1S8q
yf+KbLHv0IhdGkjcIZ3B7ZTQVHUxLpcWJsACNvhFprReSVIfni9Ni4gyTMcjepM8yNI0b57aslpL
7OC3w3EjhPT55FauGzAeOCQYP2jyHk7z2sR+3L4h/qv0Q2JhrOk6MnwOONtOmXITnLXOiapW3pwo
lKf+sw2Grdow0QDKHlQKgvFRaUhqJaR4x9sDBE+EhtGGR5uvsuScjoe4jePO4I9vv2FLsR8NKAog
LJAKrmZUY/G80G1avGX6dn7JDF7vDWxFb3kdp39+S3WGGbUYw9/N4V8401HaqxBs3pGJ1HLcrgzW
rK3FIoK9/73l/xLjvyevTv0gwCe/Dm9M14gWDicZJeXLeEW/1FJfn/ApBmKW2Drlr0uC3tLzgyFp
vS47D8m8yCGONW0+4tobId+85/jh8a9368RW37In2CtDJgIS3hcz9ArAccWAWSOJjkPrWj2Pvqd3
FRetqHQrx5M0SHb0EcsbFiJpy0NGmSS6k556USmoK/ZpYUJJG+tzv2HsElvrq9ZxFsfaSOWb43T/
3KgXnuPCehmB+W8FnzJLdXYn2UaMVljgUBJYa0FVmZy/eXBZcltV+oUShuVvHeoNvLUviypbyNEv
G8evMIoWF6EnCbRSJA+riHG1eqY9Af/8U4DRt7GcOev3n3OiPcAmz0oWGsw2qHpy77jazCCB4UzT
MX+DS2aAPH7TQE1esKqq/EQF8HwEHu1hR6s5VoP5pDs40hRLDmGkIEX24vS/W5nraLhNmj3h4GOM
/YmZtUApZAIXlxy/dHTiGyiRnRtLx8aRuYAGu0vwl4R/mTH00+07iyo2OfCRdbVWV2ja3K9G++6s
XsIj2FQoEgVUePXYhTH/TdQCuM5bwG5XudDcQ+eT7m9a1IVV/q9vGXJM/ml1HmOCJAA+65Gcm27o
SwqkpTcFHNP5rA3eaRictzFok8bjmlygx2b3IX1WMNWaAzsdXxEE/f7RqKgrlx+w2/451QwduFyB
uVtKNNjJ9dzFSw25+zZO/2iyX6JCZ8qB6Npw7TjdjZnr6C0lsjy+jDSc1KFcBC3b3L1h+oN157dJ
DHDt17T3gctR4xXkSqAoHNutoXSOdYsIAFQ3TNjR6UCyj4L+ZkDZHTERR4SUbcQOsmbp3xC0kMUl
1nrtWSsiCXQaa+U4DIVdjgXnWWMBbCQeQ3FxPy84PZ+EwlHqMWRnnq/fW/lFgVbMvHczsjlrVGYK
PnW/a9Ius7A6z67u2FkQFkUHe7m9AnQXNYxbjQGQo+3/Fk3CtvSormAbDLoqwTCzbOzDmLj+5bXT
GuDTfRx1YIIBTvSrDMLpfBMpkqGyrvK7hUcR9JsaLTGEzsJEUIUfM8uFWQwmVSbpAsixKm4xDLlN
nGZuRx6mAU/K8nHOtOkdNqR6zU5iwtkN6QsSVaF3R1YtENyDuU/6YbNH2fhgGDmuGx6Oi0WkIu6q
h3BkSZl1fyrKrWuZuxjBvkEsujyNuuTVhXr44Al82HDS14D9otUUN854KvIZHltcWsaCGE6d3UiE
sLDYdR+/EZ0VNYSOBHxGbah+vkOA+pyzPa12QjZF0SaIMwNiP0toXLHZBTpQaPkQcvTsAtBBhevl
E25bCqurfMF29bwLpfHCmoalhCpNw8MP6xgKo6xbjxVV5glPHqIcpjM0k6oQLG9dLp2S41Dh63WZ
ZD2Xckw/rAzT5sl04rRzSVjZ4DfycZZ7Pa8iCtXHSoRm9rwDrCg/da6UEh1COOmzb5GaUJ2MdUPd
52xS0U2kA3sN47XyYUKsaSnla1+2rhXac1amWJeadR1ixQXWum+qffStAcduboXpVfkZvYjDCawP
+kGmC/bPElKC/9iqvcFJTJFnZb7wpsBjmTgaIw+A89tvU+xVZDYZ7sffMbLAzC597xeQ+65oIYyX
Z8k8XzZN9i9fJ7F/QzUUuyKBfHrnhPu49w7NgyXLO+7zRYBgabmtwmmmvLPOYF3ls26aEWmhBj6t
66lu3NBSDBxuwF5yCURNIFFpffeFhcFxTZEBPwE1n9JyRFmoC5gWgD/1sEY9z8dgyoQvPRADP1Sw
HX2NYGwAC5ESxsb2ovyKFxo4z5+1wzXsuq3gmlr/SHN1h3Y8sTaqgSYCNE+WGiQifmRrsYA2dxnv
q1wtj81fc3u48voDRrfvWkIz0zrmidlr/VxBk0WQl4sAhdBMyvvnV4T4VCxvdltmtGX9uBZ8yInO
IW6qWGOjA81l2KECntnStnoCv5Sz41a8sclBnwTsT6LQitfOqPTVrfxrXk1x40QdguYz4MFkOxwa
RYF6fMebKM2bfsXwIHfgqDdJkA2Vrt94uhqQYEE/3coekRuPz9ftkau978tnH0NoElwHMZNaHggy
zs98/VrNhKD/fq02+KZ5B5eLWRTGWKIVkMWKseQ+uOKV918AVk0xZs2lwzkhf5z5Vjktr+Es+2Jz
GFxMlaKsn5/Pv87bf8VFc3niK8LL+Gg8bLF9ndlTKUMuql/NAMC8ctmTj9uRsQuohZCfsWpV/M6L
iKoysLbAVq9OrAcsM8EA29Nc4O1+irzwgJmQH0BaH5UviJnKMDB87FAU04kam0nPB6MXYERNgOMf
cI/Rvvw9kKheiNaMdkorLe7FlfyV9mqjeLHtGyBu+VoQv5c/zQRlNX3ATRGyobjCaSI2o6gu61qN
pMWVL1gvO9lWWmAqJhVfRHVHt3AKHK2UGmN6X42+dt+sk7s+Mol0uGmYOoL+J2O263zoAvbTUKir
eAKJhQuP85QEeODozu+PNMBkTtKpumxL1TVdvVLPGasfjlelkoHt0AEWgUvpM8jYYgI4qcKkbP9V
uZFPCrTZnquoKmxU3dcr8q2E40bFh8rcpUyZAyPZ21w3Ye3pDFlkPgSWpDHPnDdxEwVzszV08fuy
nFym7/x49UNOwHkacyRsPI34vCoo+EQJTcfmtOcCq7pm0g55lUAGhCOVEck9MhGmuL8C0VLdgSjj
EuH1TUz8dTcGrgEP6099N7tXCdwmrHasq99ga96t0uAliqAK6iWyqOCsZPEJH02Z2+KJyyBaTHr0
oOFsckbdyYXUyQiOl/oV7ztvLxMoOeEAjsrTU5vwOyzyy37vJcx4dleMrE4YSeyDL4/VClC8USQb
GnDxYacJ9T4PtgU76/VdD3ArgT/TmHB4L/3iXiogIKjyxzGaEuQlf1TWY7MaxTO0eZn1MAyiHr9q
C9iM7tZ4W9r4hCwEyhq65BJRlrERRKcK4UzpqupOHb1eSDgH0ncIBZaRDa9UtkP5BJW0wd8dxqMX
6xHV6veI48lcHYD6m7a5JOOT4rszxmm0oSx774KbrpojYyE2DdtYFAV24gCchxJA8Wh5VTZzrsMn
N82FTFhfmArHx1K7o1JanLoDnbx5F4nMAB0fk9vCLrswI1UwUKpNoGTyUJPQWoapEoPNoTNVWP36
oo2H19u+R1wd1uth1e0ygntVA8nbaUZeX2ESFrxrZSWzA1UQPTw5Wg1K839eiMxdVbSzJW7DQK+4
wCKVk+9geEcYntRDMlJsbALxo7nS6PIaTEAp+v02SJS7BxeqJvMOgif/5omWIKsrO3GFRr2Ikx4c
/fjP0/CZLzHXzkuSNMp9LwbVWoP7pyqFOWf6c17tDTr0G4hvJlXYVdS5MwLrCRyLfP7/bO78le2O
XMHYRG8YM39wWoW9oXs/uTEEqIfWitYhxEcM0P6/PrRaxHxnTSLlegH5jXzpGNNG+uLpdW5cByg9
kNidfo0qlu7BCC1Y+qOp9OAAG83dX5K7mOClerP5aFHuHpE5kGuILSRH4U1Axv27OKkrePhND57r
LmLFlCJYuAuhXgfEg/SM2Z6xbhekGb39wJXdQKPk26hvr7Lkho3o9YSGN5ko2Rpi7AX+3SjAylU2
/VYwAEfYVCN7+Ujz2TSUVeR5/hvvCReqxE8mF5Feb9Kqtz6vvk7ukYpnVMopA9VK29Xar7orl/cB
c2xqSdHGTa99nQn1HlNoSEHG2GhNJkhTIp9Wzr4WWXXdYzWjmRxwejygr8Gq346wmizcfoPA+vLc
Fm6hdXnC217YyrPvUDmM7b0eP/Vis5ITkzmCpFPZbZucQdMz1PqLrXQOFfS03oE/o4WmqUdM9T3P
aAR87bVbSSmxBr8pZnhMNXKWvE8o/neid8Co/woGDcCYvjMryLoluwmvG7277G8Xr+WBDxjSPN2d
8aSNx+hDbthXixsQuV3h59DI1V4L87kOzxv8IjUnbKK2XCZTT3tYmNdX/8ZrtfbI9+2goOjTMSPQ
cLQxWRJnoxXiGqVq07ebeieTLw7BpDQ3ZK2+bVw1RujgZBoNqvDtDFwq49b/5FrwFt2ZRtDt/ZN2
ISg+PWXrf3n/4oW1L3g8JxdjfGqDCO3PLa86sFmy4vsPYvAOw4g4+6vwAn7AECeiKkmV3Jtvbn6k
sNYL3+bksfuEwJXDDhWdTO4hYRw8qbR0S/KZIWWYg//d8QNCK1Mhglrz8NhXgXUb8zZLT3ByFWjI
WUYhgAmpsSexkFsj/OT+3R9mBohEZIzz5v9mIC+cHQeAwOjwIARU6jn0T3R+KTcPeBAHfaEKJ1Z2
5okHx3mq/+bEAtwnZR/pCqCcWV8/rKlN+uWnriw0CMupMQhftnKYxGM3wy1shLC3lee+/KVC/AyL
e10OTYqMU8kVvxrLpXbywJLmrtoq4nkduw/ey9sU7Z8pn54dewjB6tarsVzvkz+4960LCFvSGyUG
PFOaDb/BAPIT4cB45ySRqidrHrNndz5ialZFBG4N5wI2yplAvGTl8Yb5s1povNMFxbTvbkLeED73
QUG5iAQqQXz+1H4HwL7NUQm+a5Hy1MwxrIs5JZ6KY9KNPDi0+FdpalUOz4Rf5k/MpuUN1nXN/CNw
0nZ7GbJ4EM4V08cMQ/JGIQNeywb1JhADtCxQ9vni9YHechfgbzgZRh1AGms64OBhxVxtskYFU/5+
hfGLApVF1NPB7XaiixDWnnPlK9uLV4eCS702pj3KdV3ic7mBxRAukmP7LrUpjrJbf9fSGJMnWF4o
nxzSva/PnbIoZPm6miz4TL5RP+aP6A+cLkKaUjk3D0q7dqgXZhXdhjye1+1dfTLuBzy81DT2kuYr
6FiFbNiFt0BGRyYTxiRhHEv6VeS8jrq3EWATUUgqQRzBOrbfk9dTGLae/YTHEUu4m3Xt/Tw5wF/d
BBd8XAko5oh6g8PbBn6iKYyyXvF1RQwM2sY9sO1YCUj3XvA813U2QGhm9Ra1YwJT57nKUx/lTVtS
mKmtfUneXvtFrhtQ8e65Q+L46A7MhxDErgpx0zl+70TIecZ69E8sGulBjsUJh+2G2FyyXyTi7ZHQ
AE4rJg3eRG50GogR1Il9AiKXv6Wt2BEOY9tWc/ixN2YoRPGuHiI1UI+JnN2HBn1OYMbDzfiWlae1
WSC9kKbnGVKPXHMHc0IYGXX/kzoSIyDeio8bP2ZyRlOPK/PMBMVF7LVeFhMD5/XmKFHaOiW+YuHl
5ZeTuZHhTBsYX1Pxt+6fj3fSWdtWqBxqYeeiA9zv8tZubfIuZHCJlw/2uxxyvM+AGQG8fY4nCUox
gy7qDNkfRhtX9f5sberXLQuOACbK5ZVhiEqYMehhTj65pgI5T7IfN+qIqWt4hsJUGssqY3MKDiCp
oT20u/J+peNnOXaJKfpRxZRSmzdHftq0cXBKuzAs476AfcCHhtHYSiH/6Dktw48F+ZSbJkch1yrw
PRNG3Yh1OA+wa+dxiJhSE6FYVqA+Dt2247+9qe1Xky5cvTP2JYoxRdSQUhwod8FIAlkaPpuHoMRc
CksULhKNmhTjwC07d75P92DJY6WfUsQpP3JAGHbfGj5PHnzY8ajjyGXKAdoaOAsnZytnjKu2UyaN
ABSehgaJk6iO5HPnQ+0MRNkD8TObkcXeao3eS9qtLTnC9cd7N7j2fvp4ov8tOY/SeD+B5NLteJgY
Y7QDKznTCG5b+pPtMwJF1z+8s2cYQIb1f4YrJR5jklvppAYuJPBNb/DHbP1WS1W5qeAIpVFeXTDN
8RtDplZPOuKKea9t3gAVcArPgwJGViAAXiD6FFoHUzCDDsGtzonq9Y47ANcc2qCMyw/fgNOSwwPh
a6T4YCREAiXmCrrKDnI+q497hTMNVcepTAmY/zSjpIi/ZiQIS8mwat5k/GZ042XagISvKGad86bT
co/Drh7iAKoYboNgYJluJ8T+1SfqtL6FvgTnN956kQuHvSVERex4KitiC5Go8UoM9QAHOd3V+fU3
PHMv19FcKRCrJI+f1is7SgJ2yQCnToUFl3611Mr8y8h3aPIdQkm3ocjjsdhy7qwspqSAiSGegNqj
XB1r7j4pGU9jkp7xVK0x7U9NEsZt/Pjyg9URGiipAGFVJWu/U7YPMJMabvzU7a+ou6abd4oxQqEG
UrMxPzHPMAeq9FwKA4lLJH9xnc9QXcervymp7ZFOqWre403FJtC7HlLXYP0ksVV7La+Hc1Qycnxd
jL4apNgS+DaJfPIk+1Id54cPyk9ZQcMVn3NNDjT5Oz+V+7v3gdAf+Bhjh7BvqSeOwtoynuYoUe2c
CRTGNlj1eWIFmlYmPdb+R7lUu8abpnc3oEI8u0HlttcgQsqvlNktD2WQbzjHe7qm1kq4qzKaJyOA
RejlDCIT+h5JC/lo2NEfVKwZpXKJLICddeY0t8UBtRwQ/fPXx414Z4s+PBJUrcRz6NEECIhK/C+2
jfejdOlHyqTfQWeRdiM+ZmwALF1jVCJ/S77/0T3/Lgpx0pJ/U/1CSBjkRPspNATUE4TcySYF7/jq
LAdgzivM1XCjRnTrNB/e3iferPnKbh8vRaDRC6WeVMxNNpW/Su88802KdffKU7yDSjUz7T0QWrze
2LKv8jwT+d/s2O6mdDUEx/TbHyOd5yTvqJj3IYbGOZUuVFQEgda9e9o63GynTafT4TrT7igh3Dcg
ZyVBbVs/XlIOIA3T2kGw0e3h18zmmPWjHZNhWJdY5OEDHl7Doec2IhOSfAdwTsAa7gIYeGsLo9Ic
yXrYqGrWtwKGFWSork6RMmYwCptMKODVZId6NVeoDquG01bOlFpqfQ622jrWoXXCsrc7dp4KK38f
2b0bfdUjql2apImYIYpB5VXi8RNRUj1LqiKQXlB0/aPywX5LgByMDXpJdjexJSoRhBwdW4SzQ4C2
iQPbVpxquIBzcXTxJzWtVsGSelb8Mv0GMcWi9dq5u/Da/I4BgbyopKXOkr/jCY18EENQpSDLZ7t7
ICEOuNflkX8wMu4Bx6HmZhHqQ1Kt3HKXbEZjBln9oSD5MbWa3YTZRZelkqA3Mtg/PO543OEtD0sr
6HPruzGS3iBk5SuiJWHe5dpwuJ9gghI1ol6/O/jj/MTjJsRWNFtzfbNofX1MTxbxn9i56lIuYeo9
aiWl4cAOddXY/hQIl5p/eZzn77L9EY5SRFHkc87OxuCObZ3P5AYS1N3KM5I4WlOCFgoRUrjbG/ef
xETvzpXC3wMUdvAdLOrdJABtlcrXUIv6Z6E3mwePdX0HoD7UgDMOqIv/9Xften3MBVxxwbTbQUro
9jZWjW33NoWODLacUzgQte7QpytXZ0A+nxaFHNX90D2n0Kii1IHhJUZjwFcbAn+0PVaRe61dYjXy
cOQoh1RjW0M40KomKIKMt4VZFcApj+hsC6N3vdg8jDd/rIwh4YqPIDJeWziSWexROVxQRBaTVKcH
1dREKFliSSphZkGHR0QtOyeViOIwI3/V3KWpcdrmU5o9u4BxXhsDx5z3n+HrLiAexJuyKOZL8vVD
E9ZGdu/l2xFCgSfKq2ICpYkHCHuladfJ/okRsvwmIMDXPnU5QqO5528GDMhqGMBaiQYk8uYpKWOv
q3BbYlbsUlw73NItjVpAIIXr0qxbgvpxAC8yU476bqjiPEEYIfIEsXKkOinHTwKMLrjawffgXJSO
QMyILPsbQO2feAIe9O+xafS30Rvp0ZLJuu7Pd4CwBR0AmVqQPLFO+7FMg2PVSSEkrWekqJ58Gs+e
ZKLGsxqVmn10MvYKrZHBAScTaYePQVsug5QbHMAcWrd5l6m4zoUTKzwF/Nw1dPPdtBjk3o2IoGP9
gvsmBbsLIe70eD/MHZAb+ID2M11JeyCU8xAp+GNV8NeDXCRDJW9H0ONxPil5eeIgYTP+rix/5sRd
JGywvCi89U8Pdpe6pOihANvT9KqXAmPm1/VgEk0d9LGq7OXiAIrbcT5XFf+wLLPDAO12kx3gMP4R
xxKfJaPUPPLq09ru7jmZ6QFX7AVQT8bY1AolWeE/iWeAn7ecui3gAyC0WpZRkdwEzt0JaPahlpkX
WcnKrgv5ZFh4PdD7dQSxHQ4sLFMGW7B0aBW0vrg4R90O6Hef5SeKRQsE00nMix80N/PtVqipRFlv
qWUjeNYLGi/XwB6C5GY4dB84Fv7Of9uSp5drpHhoaE9qtP/WpWk3j83s2bVCAC8XNFtTxiVEaRgu
S/2NK3PJgTNt9XaIFpX6X5f+zKteqLV+oeN2abRdws1Scoy1+iN+EAFHk0B9BZqP4UwFSscT37fk
eX15MjsvnfKkVGFPviSyJa1kx6NYPJXeQsrIQipBqhMCaTiMKmmbOhicEH1rR0EzVxr64rXzpatW
owwhNWWJxnpMmX1LuVQ+mbHGsDma3dC78udODt+HcrlOLFK6gBUij0CNlxKGyDpvJXLD6zNvkN5T
OIKyfgMvV0zpTvaSNSvNBShx9ocUH2MxGZmzF69gbDYisiyH8BQUAuzeOIsUC/h1N4Agh9SNMIud
KVKDIHEmA0Xmc0Ed03vxSalPY5LFfNdrmCFJbOPPKeNPvGwulJw0enm1HKeROHJD2mrQHZDArowq
W2Df5JaE/L0gegvHDNNTqODHcUSVrPOV2nLPCur4IHsec2wqvKKrtXvg51EoRutj8to/mJYjjKcs
ldZnV8aHtZD8Lq2ZhQSM+fINQPhK7ko+xxXSNVz6XcZ0C42z9wOoTtSgjQAtOC8TL6hRj7O85Fgr
MYQsBjW06SK6x9MrAe+5vGh8+CWAjlZ1tfxPB37ENdA/PRtJEmyydoCRBLgWwTGRregheyzakAmP
kMjTqlqxAZImGvxAvYdwjwsOSre6/1tKZundJCqcYlyWmTunl8aelNA81jzF0FKO0TNSRuQ0g6Eb
AvDGs4+QdnSv/1Lh2BxfszRBUqxBLLInBrNQ1q4UpnoQbeA6UGxyNESwvPlw8/SVpDexYGP3jiqD
3buERhG8mx197fTSyu1LDPJi6cppYekricuJTBmb65qVbHvN+pJLXEl+RlBn4n5WXcAJUnG+pmpZ
Y9sBxIsfPcFdF06SZPKpbgVNoyoVvtLcsMmpuIglaFYxtlKyZvkhRqRpd0i5O17WOq2657TzdQDG
uJC27weqXLUPsfHf835mW7Y26sAE1LpqTIv0Ok6Iu9T5frMMJH5wvANkpqAWlVZT9Xv+eIEXJ9RQ
/cbKzwrAGLO78mQ+QTsowfhdh7GwidiH409Q/4rxPm4jCs0lHavG/a3+2VPn90SEQoZ4FLaRE9hs
tRq3/EmzEFu8/bF7fqRF+QgiHiHF2lBjX/AvWpHPghWUrSmDi0BKGbptKMjEyb5tLAsub1B0MReM
9s/XOAjmdTkHakuhjfygHMm/6pHGqjNZfFpwZWf6SIwPDe+PCAQw1NIyR23X8HoI+O92OmphOX+d
yLxVue42byopDFK6D1AxObJ/wtVGbm5PCxwVr2lv9Ky+FlOk4FH/+3F08x2dYkbjNLlBPwltbOC9
23oxmM7YJkeSod3+USIoI7v78CjJ4ZFWN3Tj1e5HAA7arpxcDQNxaWOlrtR3txvlXy/sRKF60ZGe
V5sBOsFawxPu1VEjBafS+y/4nqiHGNwoBBgk6Kr9skHsuNcctnQtLE8AxrZ7Bq8rVgQqXDwoK0v0
QQotreIVKAabgd4P8txUxxZF/rIvbw55Os8N7G9/g1RER8alXh3eB1jvUyJOSoNI/MzhTUC9QZvv
a15ai97GymsJ7QyKiu/fACCDLq6CUe2wVYIRj3EYkuTghi5uyCuO90OjFogG6O6FXO0jJJubiPyp
ElTBgcI5emwZXQmK2o1ktArdtUV2T/90N3YRextXigD1yy2ZApKw9rQU34jo3OylrobyM2hBDDjA
OuGww0SDJlaXR0NtqLDApQUKWymwgxB/9rxNQYfrv9h4y8qG4cwhKguENKpfY6JtAO9GvPxCvB9h
kqvz5kLXK5K90PtU6bQSIyeQnDPfE9tyPVI48jDsfG/7tPWBwpoV+2pHICreKqPd38Y6jCBqY7jU
IaG7YTc4/8i0JMpRaFVUhEesI1wxq3W+83Olc/dD1Vf8Btz+6QmmvRb0gaE+Gix2//siK3uKMWRz
TcwSYlai5qmni3CnSgi1DPD4zGAr7Ool3zkFfFjjLjnTEyGgx0BPqZfNnJ99aibxDRMVeUNeOJtA
8FHePPVFx4Oc+iIjoETWDOUqjqcHaycoiL+Dxj0L48MSZVBxCAmA/TqlqYSCQSyvEvOtYebdcULK
XqsuDF0ntdt6GpS1pa9qS88gW4/nH52ZiOTGfN68v5nNOmHlVqAdNKYEOwEg+BjOfQhEoUG9dxrP
dRBLyd5lS/Ra+i6xJvrXPCrXSJaUsAv2Sue1oCjeDsePickB9YBh/ePUFzufKu3CCXpLfFV6jd5e
37Nebetqp5THw6MN3IP7trkHzOWh3X7DGF0/+8+sXYLc/AF2tvJkqbcBhPiNTLdrbdoqGkfq/cjC
WtWua9PMOYC1uLr5xTObPC6TQsgwpcyRsZM2aIvKNFZwSf0uISPB3WdAelY5OTnWEQglu1MthMWQ
WwPucOtosvxb8ZGamFARufNWC9ybVSKOfW29mI6rdI2v7VwoSXVFF5b/4lrfFUiXxBWPWFqKCQiM
tz+Xq4H67RCJzRQnz29PT8uvJFtZcemNHtGQs4wXpNQif2ptdU05rESzYXvkGCRI/JfkFkJIXRZ6
HHb5eNAo74qvXnme8VOl+xexXYgfyAvxz0SRRftL9tEDcAR1mGmhshzU3zhcnU6Nd16wtRn2zRql
M3cj5VQGsE8b9LLxMLcAN5nXlM1L36+QJOptyJ95lqxHznU3SB8tNpy89Fc3U8tg2mXRkY8GQ2bJ
RUj8pbcUufM0+2XNmuksng/P/8nFe9TxIs/iQZDvLZL0XUTy7zpzdqJl+fFpFTKIAZQDG2cyXQ1Z
2KeMWgjHe6XziNlhXPTG9D8pHDSZLxj5JU5ofYsVlg9fZJ6Q88K4qKe1o7QKBzD/AGXqjRGdtRaw
NNqh+jsbFT+DJhpVogQuOVK87+aPmPWUO4SuS8vVuW3oEK0EhZQ8rIF7sDWqb5h/F5hRf0cLgZYO
8c92WhfIJP+z9BEFpDycgV10ktFb7cE+nzaEQvA/w6Ra8dL6Am/kzRoRZPC6njWYFqbBFnwI/VZ4
iJidH04iH91/xnIbTbLObeQiKOYhfqCLI5kwANzvMAmHycc7BZO6CGypJsCnyYhXtQ5OS//IA93V
+3x8kXjS61rtxLsXtVp8mYxlA6Y2JYa/aWKi5OnqyfRQjYMww+3nU77g8psm+kQ9bOiRZo3GXfRv
hKM1Z3ppPXlzE2Aoes3nQPGmL5KWT8t/LZgIiofJRylOSa81QnghBVTmbdKKlyzy8218bnh/M2dU
cm0ZQpkHJ1D5D7kS5VN9M+4MFk+a6s5DdDu2OiTmZajUJm1cflKrCPyzi3OXfNeqTAGfKZti4/qg
vC2S0lep/yElDmUO3aBgzo7QvQ0PeHNFy6bZb6BU42SVFcuWVwrPzYv7ZbDYuRgBiY3IZUUO0fwW
3nqeqwDX7MJOMEFtRJZTofGgGMYqWVQOtd2DL1EdP7kNIMav9Vs/jpy3QOU3oAnHklzRYLy8mJKc
eLOUpn6hlrsCXx6I1x4HnZy7HPeLlTWAzyw6R1hCzg262LAQKefGY0GqiowfiWouMcQkQz9NkMbi
ch5+rMcLSbyidB0kv6DWW8FWlbJkQxVSTlAHO6f1ISxkP5Ekasbmy0RzeD2dD4kSzrpbQDjDdkf+
WsBN09OjKdjeSdCOdUb6pshQJ8nqpXqMFnZbA39elTjc+v7Ke2i81aqYjq0VZjqHHnNfLEPKl2Vz
9NlS53H5efdDHYu01XXLZl/qaKSD6xuW88k/rgn5qteWqnbsTCWeZztHI+0DvN0vQ+fBgU8UiRK6
qt9KF//XFOzlVfZv4Gujjg8RmlLZxqXbzBDMNbjVq9dl3PUBUxNVochQwAapd+4CZ3pBNYukF8mB
pCxQkTF93QkBtBlLGtAwR3wlDEmtC507chwd3yJb/kHJNyDmE51eWcevRdOG7qcFOl7bpcxQo0hp
gxof8J2VkDS4OQTyFqv5a0iZLpf9Cqkn4vv2j8c1pikPAiucjWk2zWcrtk0/DvhxeBKAIzI1sgzH
o0K89H9AVP2hXTBqtCN0jvNzJYhpdNAy5QrYtDuZYXAxxYIVbCbuv+jg2Hmv89NeAKXvlse7jtlJ
qJ29Av/C1wzB2os9LjDC3lBcMPRzBTOap2ih7lZ56twpJ/hvpl77jTTVKiBW5d0ABF3rmOt6GwVd
MAUDJS2tHQTCCIBEPF7gGPiKKtirzGpxPnPoO5K3yu3Ve02UgGvQSbhlydK44wy5/5oDqozywQwN
FlLUigl+jjvO0Pds6czLIhrEQHmyYj8214dTDSMcdP0NzlQ+EqPKkI/dT9NpRoYuZGuixBpT5F76
mNq2cLHlnOUVuFkku93eq8HD/elgfOiQCwEMZu9ZU2/WRVUjd8zZ5ucktzYyLC+m9YYX/19kJYxW
xJ62sdP7JCchfdHB9ZtYpklqbSskHlDg9q0/f8o7QXrRzk90QB6gXIZrkRdeZ8b0ohkm30k8+AYi
oSF9OG73Tm7b1Gu+UUXnIOLYSNnYm+hQ8nxSF+V6e6OMrbsLTSW3twrUOR5rUr+o0VKLVknSfE5n
vbbDoxM7PPptnsEICoLkhqWTjv1XH1ngoWJKDfm3Hyerz+Xp+BENtU36gjqR8qCR34wIORWOqenn
01n4t0ihMkvjynUFT6jOUkclyQcGvRkzwLFVrwYRpVEO0FuaeDOCBPTQC1co+o92I011HToKafPk
84nzWxbrzKN9dtEzKzrCqqtPGqciMqh3OYXmDSccjg54B2CmYP8bNFnUm8Y7Qy0MKwCrgDVCnSOk
A3ve8gdUGBx7mkyUNLcAdJd5Smy9dU829VY6qefo27C6BM1vJ5WfXVVhngcOWk0uZZWinXJhcz78
DOgSHsjQoEnmsLwT8R6cgdnvHE4/o4Lt35oh+wa1JzU9hydokkZB4bHzVskhUtnaOE+ZFbUUOBWa
WtLL8U8FrWuHzHa9Hhehpw2Xpsa1UXKgcT3NdPEnXU1MxD2LPeQz1wmsod/ZQSHDHth+27bOVEhn
Om9c3BFedjVQRnwr4T6KayEtFd8L39zzuPF491UzXmcjWbHK/1MyBcakezvP3mLMaZ+KypG8P62k
QcfemT8ZOk7COi4iglrPmaOjw0xjs0LvmM0lb5/tE4MwADjg0oyP/k3qdiRp/IO/vjQ7X5FeHqGm
DEVa8Fay0VGkpD+XQnyrDhqUydDUyvTp+ZsPHkFyhhZad6LzgMFqV+ndlh70MnZIwjoSIZmvBXcU
MGFP2TJ3gQ+YYdG71fX2ynXt5wLqecluT5v6FVXfjNc9hH1fUsBjpjs0VfreJApopGHjovRFxyi3
pRhTSHmx4APnTB2PLsWmfBnnQ7I5EFoL/WwTlSKHydYqayTOvj2Fj+KYgN3zF9n/46RDElQTwify
RRz5BtBqZwCm3azOIZsxyQ0x3zR016W+LFz6fE5D3AF5LE9+56LxDdrJaX8g781M+wpWchGAxBjB
7z5zfdwTDRYraPJT7+Ml+HFDWegd8RnxytPVMPnVKZo/8VcgQB3Oqz1Q+77Z9M7cP3x/PK0h9hXQ
USXMAvWqK5Y5/yub3zABGCs4vvcB6CluZUWKsyB9NcaVyOdpbdeNYzMLBJhAZ0g69gRIvJaff6bA
9w30mzpRBdkcvIQxFjxr948EBqrU22RAZ7W/6Ua0H1wR7d9MxI276Z5GlwibkAsTe1pThc8pI2eS
Myihv0mV/gGCLZmABLBYJs/jQHrwAX/HKcn5weuubkq6Z6sbEPTbmUUAjM0bH9yJ9KmAaguh8jXC
4AAASidMbAxtThK2Ot0QnXkpQkVhOaKtXnq3fAK+mSVnJ+7+6u5YWzlXng216PMKeuAwagN3V0qU
MimnIHhh+86eyh4jQgi2AejIYGoI5o1C2iZeEoZLsKFFIgvModZOBFYHfddJrg3tE6uhfra2ZOjy
5PFN7V5UuJJU75ZpS0+kSJ3ZYB2waios3LIwpTv2EapYDcIZsJWA8eHr+U6oyvpQ+D8v0p8EyVqL
q2KdMCfHNskKgU8hiX03TE8lwF8sWcvfn7zQIX51UxEHyO8dQ9Pj/GzJayt4S0vremFqWGCqb1/J
6ioGBPCXEaXQq58HXwUIPokB94t7b7oxgVwFioxm7sIvW0u0AxlFkFocZ6kanLQyHW5WOty7N/Bo
Cbd562Ty3arQfILlQPv60eC13EwamAK5UJ2i5riDgVBxuK3KvW19fEUBOEkT93bvoIv12MArNb7U
EiJaSWIey/bQ74DyqU3hKRnvLtEXyQlfyBOQiMUkqdeu2ANh0zJox0XL10RHeY7UFvqVQ+GDv1t9
nudZniTO+QvujCImPqZXyizOXZP3FXJgnUd9sAWMKxcEVixB8cJ53d62Fg1zDXO2qaMKqyQEG146
8gKQ428CZO54Lu4qAcTELyd7qyvjftTqxmRQzd1TKbFY6l1fF8bI3ifENaENChnTVI3wZo/SbDS4
bvTmpeceMZfRkuj3evdqBx27Kt2HJCvX8Jzy3K+nLANhW556Hw/jYv+g7apJzITt1R58RB4D+FAn
ad9YKaQwd8Yr2H809xDVdnbz1xsRjXpHRbLOtPxoVkKDmybR6T2Ml6Biycl3vZFuDQAziwwPpbks
Coemi8zpA0pei8c4UmBybJ2wgvFEkdn4KEYj0CZ7iNcpox62xoDLRNC+e54pEsZnn31AiWVzHeNU
HF1tffQGJJHZDYAx58lXfdkEVSa+K0Pfl+i+yV02WYnM4W6oRpAOwr+D1WqTFzvike4jcC8UuYH5
VfzWPW2srEqnMsRwq+B2etCD5bj7jyEl7JsQqebiVicpDYQ45NgR+VQTCS8xVbLc8WW7hl1Tc/rL
GI/ApPOEIRW3EwrRVzfQlNfR3PK/78AO6CSJNwaaiQtogf7GETocRAcVDtJ/REFkvlOd0Pu0tBFF
l/poc72cZip/XS7y9L52J2YPP4Rlm/jdyZrW09QKJKFIxi4TRg4SMofDinlDhRdXkP7qIZDdn379
P4vKM1YciVaItgJpuZU2H6orMbUid/zwlEJ0G8W69o/ws+aEX3g0t5JkAWzVRE9wguYjc8/urgn6
mXR3c0NAZSNS+XgWVfC+rz0yiiNnhBLpE8h6FrBcOVAwpd8wSDf4E5+rtsXQPpbJ00eCkvGIbfP1
Uh9XBx1RlhduKhHHfyYJj24Zdxzr4EF9euFtwUFyF/+v2+4IbERa+FKrFBmr8YYZBD+t1vxCpgD8
vtf213wYR8/cqKW9OTzG5BeI8uO3aCUB7881XXr9Wwzv7EMdtxACZy2Bottf1KWCFMOjreSHYeXm
TSzmVbF636JqOPzlvtMfDqVhsvVTGv5dP4Q2cT3682l4sjc06UcA2ivsI0ATuE5d1ObSZM0fQ10f
UVU4SHgoDt5mYTF6TFQ4+59YUtxGZr0/FQakigmB0oj/RjkeLBP0knDDCJ6lTlTFN/I5FMW+gQYc
bZvMqiDNFuc8vEgvK9tdJ18EHT2bXqie7S6O/hfzycm52dOb9/uDumn5N4KuQklm+XElre1x9pLR
hqrYUBhmfzDCV50f+xeflIUcwve+dUrb16ue1R75/OxTL/zQYujeOqIL80wBCVa7s8rpVb+/9a5L
i0f70SzQmUqEzt189dfjKroG0Zi60UVM0C+FUpXhMxpAZcIWxbhQc2JRpi6PFIq4wc48M+1zZNdG
/fhRlV01CC0gjQtUHpiVl54ehLBF1/udSLfLaBvu38hdLm/BYYwoXmRDfTmryR6kIPYmPTXIHDKf
PtihTbi0OP5YIQoGeHOHDS/h+RIKtUQwD1rs7hyma9BdFwclJeOx3pZkKYPFnqw56jrT5vo07mcP
CH6yzpV8dn5ZV3bb2Jq6XUmF2D2xBqgJR37J6Tmkis/W4cwrAK5fU3q3gj0Kwz6c6VmiX7XVizZx
Xhi4/ZgAyamr07rsl1lr+ty0N9kvY5HaPeNChVA736MICcXIw1RSrn2bIi3698CYFdr5QeysxUY+
JiyC8mOr8eWxLABUJWSg0DazjDUn+QXkbVvl84gKyhH+/iydwSqoSRNazb0GNbwWvk5UPDYW5jRi
OuKx+wVKX6gJX6ku/kI6MEBROAoo5/bbm25INJzLWoEjPSVRJvItBaYcsnPO+fuWhMJNe4DNTpYF
J2UsD1TSv0OOy6qWpc+zLLSzRub8dozHPJ1UeImQWknsxy31w6Qoij74Fi2J7cvtdh4AXD9i7Sw4
BlzkcxsHEnsl9i6y1+f9b3Bc6uVWR1BIAoYboF1qNIXTDVibSUy0xWoAgH8YqrcCDMoRt8fIF1Iw
NRAkybjZiIvqxMeKXkCq599FwEdlNCW12He6b49NvTyz2SJOO3o2yTBOoLPfm4gB1R3RkVPqnluB
3ZK/UirvA+Qh96JN9rN08Ua4fBL/u10lhd4FJ8FzAfmNwYYSFl6SPhG/4TsLhzPT+QR7k96RqVJ7
2YiJxt4VMcZUommyLKptv0Evdo/IhD50+cvodr1P+93ifqnJLmf9wUiCRZ6ZV3bIc8JZLYoyHBa/
/CVRPhNgFDda+mtIBcBV5EyWHJSrDQxRdULf4HgJ2/DXoqYDGsSc00heLK3FO/B/vdSR2UPWkZLG
86hDDiPVkTY83nvCOD/81WFZ4fnx3RPp4mX8CQH3zvcpFU5IeIcJAE1OG5DP7fqMA8J+K96ixKsh
bNu29LVfvqrl81olkf0/oMS0ONwHMUInwR8F/f09A4GWZZi84AIGDBnHihUCEUTNAiE19F3wcU7Q
ZDOVhvsLhNLn2MTOZKNZKnK9WTLiLOPTfCjxpmbnCal/N59q4ytJ0z7zI0y9zgd+5MVZT0fx2LXq
Euvfu19ZjY2Yi2Juf9cIMlKS3ZFgCzNMbnR2S2LUQEhzx5+PtE3SrzCDfDiz55UOzYql+VObFHbX
1+qYlyyyHJvV/ljWrjFGHm3/Rbx+5eSEBHhxSgDDZq/fyuYhwX66MSDKlTZo2At2S+i21IiktHBU
eGGopkm6sn+HO/RFalLsBgy0SpATtMamCq29NkfqDOFgTEie840F4miYsrGQbYDi3xz/hp/ulHFP
Eq7fSFQWg0GSbpFc9Fne8aqFiS6/IRqczQICzr4XxusTudQq+h6wukxZtb4hs0g1Jf0NS+IwAXXg
Xr3JKh9WWAUdqlNHZgk+8IxrZleMQ+Co7Mfkt5GNy0a+WoOMCkxFM5qBb0kDPW2ywf5maCaJy46Q
BBBT1O6wjuGMXBtI0vVdwbfhTHmceNsH6mjFa/LP2SKQUPfCAFKr0LcpZoQsrYqrhJ78wJh/FAIT
MdLvhXkPdHlS5ykyA59kaJM0gtOesx1IXnCaZNZAip665DVWbpEfZpEYgiXAlaUfn9oth0JE/dPt
34h5PybRiMrt+Tu0bkiMaE5N3+B3rnGG/9SQDkGZHVEJhU90nv+xA6ZKBvZxeSUw8JXUA6RNJ3Lx
CyLt6UmNS6YcWgfInmyTaBbfAi8vlIA6FaZ3ollhbHocR+zy74guQnokKLRlZtM1elLS9zkKmDYy
wnKMN3cLOpucsdZOnfreZ1UiC3bowMIPU783q18w4lGQLOOU4K7Ga73SH99fE0xrB399uF0a8GWl
zeqVfMJPvQjM3fEUR0j6Qraqh5p2fFybSrAc8OJmRJuf/FwKIQHmZWmtSeizDtj68kf8I20urZ+f
qE0qNdqykRj0NFAqamqmxgaqrKjJgPh1jqVF9T2bispMqI6UtsnN1zEK+/7aJ8QDbW4iGUtmeCYC
z1XR2BqLpK0mjvLIsKZiRBSRh025Wg609kCkegtW9VeajPvJ0cEX4xfxkgNv2F8T7ofyZH0P0cbC
z0qEmtJ6QGBcNzCtonTmeh2lwZtCbPMhJZctxQWZkfAxS5V9KdMB/lxAWQcLPJqsJWkgj5gvYuCg
jgHcSYI2B4gy1fOe6lIIGNrXufmL5xO9U4KLeDMHebxb3HIVCG2PfGsuTCLzLpJRLgOrhJpX22w1
jcJkKrR5N12ccD1RXxgAY+/K/183llnayNX4VqPkaRGsgnC5cUXbOCjPlwb1GBwGTAfmo1pN5KGk
RD+l9sXP2ZCYs2N2yrhJsmw1SDBYgQMP3aLMi5+oiyJkVtOa3lu0bMp+Cv/5PBWwlr7fa8L/zH3k
zLbtcKdv9BT+TceR8wKDV1xDqP+5nWIkQYq9O9aZc44X9lHUnVU6EbCUxCYudq49zu4dA7wv7IUN
ULgsMW5aYEEo6otQYPGi5GZRc0sFw9sk+Pfn0kbCBvTDX2t/cm6WZYlQC29OlZhS9IDJISQlfYj7
4rOKmpom7dtfWhC3qgBR6b0Jfe7JXKmRTVgXynJ/z/Rmuvb315F0PWPzC1Y8BnVmMORxIA5XEwxS
DelWEEgEJvIoROsCbLnLuvbDnTHysrMltzqFsyADaGmBiKsim7YNhxU0CRm629wbVkz1er18+ptq
JvVE4jehPRCHddyILFTTEXOeQJRn8BJNCsu264KcW4wivkVrQYURMSLvQ73QNtRe0DsQ+OvftfL5
bzESZYI8gRa7CGhBgBmZ4NpWQloUnOaEueKc2ZuHHviCKqxQ26oR5NMDBi3Sy1at6NuwxoHL9DlH
6VaM2AZOQHjfSyuRo817mit9WLIz1CqZRq0P6bntPpgBOOAra/q2mYKxPivP/ypPJw0fEFxALCKO
MFYRhoO25vVYldl+NEioR+oXHFwDVwAxzX1kFpgLR0CqPVAnIkgd+cD0TmKsJ8nsZ7gl2c7xgpLT
ky/uIgGnDzdHBFC+Zj9SobuM07tQkcYyl5JsjUtmFGdh8bOo9LaOd320TYyKlT2l9iEfy779G8zh
dRNyg6lHFritN4vbVPN+PT5L84OYMK5dQMUdIHSjJUn9M0LetXnqaV5f0I3/IMOn5elgB4jpJIdY
QpjR9fTTyiXIOeA00hZmLtddzPdSRf2SLrk3MMW3LEvLTPF5eXrBNBm90Ax0/skYTPSHanWUVnsn
N92xdFvXREHKjDSb+kICIBoPua1kHC+DyXKDXMhv34bImsNCxKRoffo67vg1Ee00uKWL7D+tOI6y
KzJIwY8HljvopF/qc3QGfeJ3pP19KX+6k2bahd0/kTUvQdUcLqb1tk53ozsUDHHDjHKqi1ABgQlP
dOQZDDHNB89Cpj7mMQ8Y1IGsJ74BFhvhJEKtNFQ6g7+EAXn9kqgSLmOCaNmCWdYFE8YhSNDv9/XA
8MRlpsbtknsR1g50gfrxcmGRNcRe7QakaOuJRZRHpk1QLgLfWo/I6hJoJNS7UIcFPBI2CLZE5J+G
snN6uZKVsWhHHJGkTdQaVAWR4UrY9wQwiL95hyiukN3OVm3O7de91Zbo0g7kjeYdkiAhof43Yfus
PB0AlAmndNrHK609ykSF6EAhH5OQOQ38UkPaInLjavddvWDxET1pR5nmun70zh7gf7+7C7XzfVYl
LPmweYn2YkwxRfmqEaLH4d9MVzuCYXULe7r1LAdTcT0T2ijzOZjVz/CMwNoIRDlsP3HM8Z5ryx1E
Ma7mw5h0JiwTk4JZw8Gftmda72SdAEcCgP3dezSDuAq0/7tcY53ZZpLX7muM8CNXqnT1Gf7YWEYo
8ZJfc8FYT8OIJKlzXG5GSlpiIZp01Nwbd9VD1ULC2ugvoG75b6vuM+fO+3p6MJzwztuwbAL0W7zr
aUqDItH90vWLGItWhnrC7ccqbCsJYrvEbLPXifUVa2PhgJ94Kg/E1FM9/MrdhJuJpLHUs5qu6uRB
+IsVWtkOdTtBkrTCBMp/gr/D9wQGpzdQB9ine2XvUAUwBqoGnGjijdHrCjzlIcKp1aDelFJqCJSC
jINah+ArFR+CYZ+JGAXf+mVxUvwIUTxKQk7Y6yoa6D6qp8yzcDd0vnnxft5eqSK3qhGRaUC0c5DJ
uQON2bf4VQMiDKcx/meWbS7p4zsLYSJ0vOZnxiJSv2jaftDnB77Q4plGWWYuVUSt0kdQBNkz+Qrt
fLbH8t5nPbV0sBoCkUtEnWGKEoAe83Y2eFtXa0LN00DitjVuD9rMo2BkdIL5c9Ez1DJ9tlhDX0jM
g+FCGJMvnU8D/hVeqbVTkJfWg6w1qsQGj50BNqkc634m7mf2mG70Yds4ufssLRremVYKarWezf3g
dGzwU8BK6Owx73WetW6mQCRxOTIdpRFKnSZjqtCaw+cmIw+IzjqrSdZHsBsleZmT3Su44NDctxGB
+TgQm1tEWIVTeuJvd46BJJwoALPPbKzzF5V0XMHCWx9S0xAM6HNoROw8uyntNnDMhyJzc2R3MQ+5
77Ntu2HkBxNS2cv3HNZXVv5rjDZhJvXMCq0AslEEtnEe4DSZvhn+IB67YU9TFb8nXnTP/oMyeHF6
xzuRexRg5IzDG3WBbb15P94Z7PodjftQdcpjnOAx4yv2YEZLdrYpTwo4YB3jgb6AQ4ayboIWHS2B
sgPLk23fAr3CDwxtVx5Lqj5WOfTAo3Fmv+JfQQLOH4sYNvu7dj3UZ3ThRAeOyPBlV2+D/c+IJPyg
jk8bH6+AH00PNsH1S/ztIUNo0cey88ZTC/RDil1g+WBW+vBoBYvGrOBrsR7zQ+UdidweaY5MAdVU
rkhxgNosQ1EuGKeuYVMFe3Q4YR75F0HDX7W0/CZP6jyRSb5o5YE1DyNihTxCveU0KqyokagxRJZc
tbOZUgpefDryBGWNUZGrstGmZJXoLI9CGa0Si15ELDYST1HQpdkyerIWM1jBn/PRSnkuOd5oc2Oq
/p/JLTbamy9njYQeDOAdjloBj/0j9fwqOlvovigGF1giMccW9jjNyxXv0TpNKUMAdgNIpOgeAsEY
I5Dr10lsEe0V5INam+O270dITRWXLk7+4djlZgOVEGwfikfDe+CviRbF8sRf9CcmYMqdYb8MYPdr
Uga9pjasiP9kLxLDmo4KL8/uI2alVtVgfbjZK0MyOolxXsN5ejbq+BB/JnLmrwwFaP/gOOzIYwug
EuKDzGU24pXNOIN8pOTLmpDTdBWq4RT3/z4kR+Ctw0aZOxCuPLqXGIQCVNdfwgu9m69+BwbL1gQH
iP/Eo0zEb0JeBSU+eUj7qVT+5GCB5Zmxmoj6pGSsWebzSpnwSNJj1y51UXfnzTmPKzPGepLEuTCj
iU5bSP+HLDxVeUQbCMXnoXSOud5rYOkAc9arkK7SUFX+L8POH/lxcYTvP9VQHmPDHawL+uVvifa2
Nn6bcHa7UrPvfkm9qmEdMswLSMO2kFUtNWy7ncj4GKZNZ/yeGE4oYePQT0uYrJy3fmoOmD548BND
u0iapvfUcX++3BA4Xah40BXpeDSq2ZqHyApIuhTObfyrKjN7GpdBpw0b2jtuDUxPPPfyqMfXEqnn
vvcsMWmAbtXUOYBWGLcAXIrohfp1nA9WGNJcx2CBv+3ccWefS8OFlM1BikGKhAM2vKGkGlHf8N0r
xFZganZdZ5WrvL36L+vREMh42Cu1N9jqzTrpvNLU53mlmxThiNVwdrLiGhyc4KAUZ+59VncvvCIN
qqIyBkE1te5C+1xoOnczk2CHsO1A0eeAMVAzZMa77GBQNnDGKXlDThEu72M+kolbC0QumbdMka9f
D1U0gg++jbqd79ooVcNypYt/DsA7OFt4yXyUoGZiJ2ncXLn7VtiRMsuSJK5fuby3u4TwpPrCwpUQ
aioC/kYgAzmt3iEoLyQJ0ctczn6nizAhonN6c2uKQ3tZQxNk39CQddniqVxcXks4E5iezlxuqfp2
fEvqR1MzzPHQzSfrwJa4tv5gZ9FDETm1VAUR+RqAQrZ79/eMCXvwxsS/o0iMm1MOqKEggU9ElEop
XzdlZAdaa6Fjbfs5FVYJg9mXmCBapkvcrmVyeWS45zjBwlsDhbqPSWMaYQwvdkvCiZcYryWfDgU2
hb8wZ/6ziYEC+F0SU00xIN4e9BPrsnvH2JR7v9rc37itfeLK5iEXyIzNVNediIHwhhjvhH3jb8Oy
c1rzgI8Aelyhh6Evy4YwR1s9wDJYSLN1LQhF5TMS6/w3pxdhiirxVQrVkPYmT27DhSvtXdaQMuMq
yia+94/0wtPDeSqtYQenzIInjhFUzks6/H7/g+s/z/92QL1DmcH5wes3z3cc3YlY8qaFRkWUA+1f
QwrrVSriY3PD9h6LFJXQ/VsRdTSxORr/5vMsGXuNfDfQQrpvk9OKgNyIDQzdVlj+cmbcfSdo79cR
Ozur1eGdmsK5Y0xySyZHp7loZqKxm/v6UK+nxE6QTTXBzsAhLCYoqyf1J5lSHHruM2a0tAsA1iDu
OkjlZFWQ11OAA1Y0DIcb9o7apN4gWJjCmgn+b2GR2/quvYa2VB+nKHafZlI0r3PqJ22wgJhsTtgf
Y+hIsEs952ioRpaU+07L7bKR8DLqIjDXldgbrUjGOxDw8fcupSmN9jyE6BaQFQvFKlj0gTUo+hcs
gEkVx0JSvJzw/WkqkqF5D8xzzLpaX54hNuliqMo21Oi+bSEuKaaOVY6quGUxOHll73/dkJHi01+5
v7txoliW4euyEpbbapXom/PMRI10sIA4Dhd6spUpi+ckFSo6zI/P2ScszFDf5SO4SlSjEEcTWG4z
lOSYhPOtEs0GgplklaLJTYmwxNdNCUT1UjOlWp+RKoZxW4lfY5jwWQEgkMUIW2m3T6hLxcKOxUTb
D2Y5QMmtxGC7EdaM7CLGtqOT1i4RjQCKUdmBjJyT6Dsw8vG9UdFMJ7Fqz2vTe1AdTM+/6kN/tclv
RCzJrKYimOVwtF8Oopkga2u5S1HH/qDLd0iiTIJl9XQSbXZDY/hm5T/xI+X4wqrWHnPbHHKwwG+A
yNGXfCmvyJoSDt+OCJn9+y0fCF9FzcXiBbS7WVQ1oue9lKTYcppL6UXTA6admET7WgPzgZJY4yz1
xmaBzsLITov+OqHdUM0Dv9or9kq18yHzI/p21kvmzxEQsvhUIs7QIiPxAwuaI4o5VarOaWMoYJS+
/exaVXX4Vx/x+khnSCDngl8wCyJt3q2Tm7a6QgboRxH39ozTNggvy5z6VfABHP1iZS35TH4B6PCu
Iky2Pn/fV5Z4pQ4sp4RC4zJ/8TLJDPluqQO3oz2rfj97n/BFT7xjKzdPzYXnNu7sdsLxCyB3ojX+
v0ZuT62/wSyyQpNh0aRg0nU+jGJMlKE+ms48z5L5QirH7wM/d6PATAgZ3NXUEAgvpphL8kuO8LEC
YdJr2BluRCW5YBIErxA+PpwLLr0i27y+99H3qR6qWg92VYyACLEUiKos1FJHxOjRO3wTGSyOYpWd
/OVKZiSoR204wG2QJ0XG9wana//7vPw/qCs5y5iVdxFKYQf3BQc5oEL/TWwKephOZY5GAoT4ZtLj
rZSt3zq64LYuOltJ41W8Xu+1u/ISoYfcyGRClUxc7sSDQuhlbYynL2hvjaNvttqRDpM7BGWmN0oc
fH8gE2/TCUS2LYH6d/Jwar1+qMIfiSFYEmamdBwUm3ZfUDGBhRmfyF3MkK+CP5uHW5cv/4FmNhUH
NPI3y0yMWyhqAfmwIJ6TnLqaXwc6vRndoouAExlxeUb/77u9kiNWSRSYcgXbKLoVZpL9WOnI+Mnj
Ue54okOf88Yp4/Tt5VWEOsyvfpYRViNyLgfWt+RQk1RZqgtOF59WUTLaGf5J6AI9Bmi6om0ZpO/K
l4JwqLmckciNfhSMrEdEXtGjWMqeQAANfrJ4ZH7YFE7n4p6N+kzwbbK9kTit9PZBpao5jX5RGvxz
77GTngltTxPKXue6o0NAHY3Fpyy45g7G9waRcCvvWTd7Je3tIf5FDbq+sWWN6S5vd/dRv61nDhNt
5iRAKQ4pv5faJN+V1YktIBCufkFdt+hZbwnK5B5bpaNOM2fyB/+6MdPy1n/rHrmSQPfePnyEE4Fu
UyRQGnNpk+IaD6idPJV5iRMBpmF/cSvDP6A/2QAeEuK4Z3Uk/l/7BJ8nWEnfnGQbzrsZwP7jaM9H
tVj6FPjXWIvTShKyHxCHM6Ams8sUdOcBVyfdZuj5yJYV8j6XtT/qCJZPpIAEaLtwzmEe3RXx++N4
AiiXm9W2grD/XJcd+qCe/H3co08pvLODew9fR0HOPpwRcdSHaWTWOkKRP2Uowy1QIFeMmIvJGu/N
4f/vX6BrUSqLvi2YD6m6YI+Z9/mMSxHBNx9En/c63Hae1PjhIbOa4GqjJpy611tS6Hm/QvrQm+qV
Bc1zcbjTDdnEklnWILp1XgOE7B5GUT6DzScLptGRgyDmvxo4oxr10sCrkdlOEljuzIHTAd3yVMn/
gk0I1hzYif8L0QngwS2/Sm42hd8KwzEKVsXzu6ZpMxDXpuTrnQr9YEiXBDigoj4iPH6tmQUCvPTT
fn/4bxLkhnUCszk57+zYdJSn/1rI1pq2mh9R3tLb7H2fxITd6bVxpJWTOXvQ5MH3vjlV3omZdbzg
LZEBmJpbDnRmISG+kq0Nk71uoyTwn/qs1aIwF0HYj5+LpP+L8HQV98AMxoaG1PrO9Ja6UUHlqtpE
oHLw+IfX9rVkipBhws7QNIVB3Q8XCTFTbMe2ql0pICcnLTC+wTBysF2wNnGdQ68Ps+yhvUfQbU1z
Xz1CWS01jqfHWkb5E5llzENdiRNDs+Rzs4wU1bHGUQAaylKxUVCOJmalflViTo7/r5mvb5zaNYm/
QQN2nsgjlDek72vyu9LPpJDT2heM4E3C0fBdWc9e3SjQ/OiIzurlffD0Os7v3SFONgjB0SjR48aO
76XCbogh6+W2uGW4+1dhwbFMIyV7I67CguHeg2VrOPEfDtQJ7XRyFZen3H2HijMBpkV3TF7Q+I0S
8i3sezS586zjKdavvnyqI4e91eyB7bbFSOU0mgLjfZm62owf1k+dEa26DzNly2IQM9u8ohazrN8f
ubXctnH8Z8PSZBvy/9lZ+U/Y+RjfcTJCNI5q7UOxiGew8UkNiADfhWlxo2zbR5bLLtug1s7nOgj+
reZk9h4P57kvI274x8lSLte9/bbZhphNjzjc1xAZn0RUf7tkICTNn8kS1WJlTXqrTTv3zxJW+PG/
rk4bzRSMWn8K3ZR1CsGuWRQI93pa6YuSzpQY8wwWpPu/7h4cf8GUXhz6maqP9514est9YMOI91EC
C5Jbrw/v5LxDmGJC6vZkuzU89TQ04w/CxQ8unFQGpyWQbPqb56jIU76RX1RgNALZ7gNvuFK3Ncad
Ct/lirz114ePdCZlgRMC0uffnTnwJt8OmVoriQqrPE+X6K2WqlJs5H9gCCuYDE4oVsAfBzC560mG
a5iKV+12Zn9JfTPbQXHl4i2NHxp3N1dBI1OMoQiS4eKgqGHWufaR+9wnYVFEU9OBsPD4hEJDPE3z
wP7sR83rbDJfc9yIImYbG4XT18LZNbOS28whorAS3k9BrYiO7mkq4ZEzyy+W6lzFHvFAWkn9sDD4
gImQLcgiqXFXA/5ZIy+98P/IY+Vq2KOf85eG+fZgIrijvMmHXl2umJdo6nhi8RV0s0PpA3FJK8hG
gd56TgM2K6IlpiO9qM2jX88tbqqonj2AjQL+8t9t+VqOYUtLfbpPsZb53q/AnK/BcriX+PWrqel2
7iv5roicwXzVriL8UsTOBubbaglXxCMF+qWV0PPY7M/7xv66jaXMdTUjTqHjQVSty5JWRCgIuiH6
3O7mx/rcPTOdvdS/11/FCiifuXlsW3560D6w9GoJLCQAG+FjOUaOqPhtRB2DizriaKfswLRPtpXd
ld/ILRmjUMImL5PfBMlgN6EYG56aHch5kf+wFCUbgWzwrMRdLkxmG34rsOVR/3lKekwxMMBzCfo1
bX32tUixpDF+rag9DrlmLR7AkSxxi79HaP6Uy8Qf45iZIuPjF3r+pfKxGTBetKX7zxKBVLWaEpt+
aZouYayCkqPK8qe+IylxO6xcYUXlgKNedxeMMGifURJ1Fmi0gXt1B7yEiwz4dmRxUJd1OPX+TsTl
EDgcsbLEoPUqqeMXIbfvnfiD16W5pgMocdE9U/46JiVR51Rem7QW+AaHTHamKIIvMybm/kpZJEnX
oBNjAbvC04U3Iu8B0h6uD4IliAxIzw+GUZ0omkjPI+Mt0+i+XaQ1D+5ghq09D9aKU1Wwbh0s7A0h
9FITyxC5R7hIX6emiRfvs2MXMEBdxgy+v/VtPEasySYOrPsUQZwNTZoGzsDr9Le84V9uumFtblK+
Y3N7EWzPBxfSX9MwiP3QqnURJNVc9A0ML+nfV9MJ+nPkqydyhcYMLWmiPz99Eb3dtbvxEKDqzQ1f
VYl+UTFdry2b/qcZJpPhG6oCJFJybmpZUtGboHY60bDmPr5+/bnFtPdm4qTHXrLbVbHlrhRUvCnu
EDmMtChvKEnCrtMHjqaEmUopj6u6ymQZj9UhO4bjiDFDpwOo5cwO+Ga8Ub1JdwWnSpu89P2ptKjB
FF/zBHTkwk6jXp2EQ1sTexn+KeoAF8ciibNkiKrcvO3d6qD+U82tOhPCNU9M55OrffM2PqxXYIBX
OGGmhtnur9WZQXmZRE+NhnG4YMROdzvSD3F0lmsJ7tNtbrYUIhCgOxCOYg/dMvYO5Bsuv8TSOEjX
BbOHCe5yG2k6kCme5DUPBr/a4UhVr3O/mEUN3pyRH57VKk4iPSXW/E+TDVSp6Hcnd90nozLUYAw8
zVdsfWYrdkP9tPimhogtVHDsG2E/IFKQHPHYSC2yJuUOL5y974DhXMNtYn4wKoUf9SMBEa6+8LzH
Gy6J2s0iu2fETzkAADWIsMi2HEaIBp6bvMazpj6QjamFzzXN+Bncw12hbNtHhjX3VsF7637Prht9
ejgAxdEcc03sxZcqf+8NJ1nIs35Tyk0mdKHDqNIaTrVrwu/8m7VbFdKCT89Ka4+jG6MjSMX7O+VA
A9KdfLrUqJXNl+YdlU8/UCqhWLxnUOQwAa+i0H3tYLziqDG8GEJ//e5FuyjaBGikD18TVLw1B8wG
3MLvVA1GjuQ8l2ZkqXL1v9gHDnYyWeABQiUef+2u5h6oQPXx/0Uw2s7Sd+B2TwKTYeuTAnIWoEdu
2cXGTgh7Xr8Edhwe7AzSStaAMvhq8LIXR1V2uQ43r5q5NRyod0SVGletvOA/A/CWH4862y2IuNcj
3l5Au9JgEx38Y9wALS6XMGYgn0AqjOvuzdtHnPptBDrRHg13yqZyFEPbMVTDXAwQYpgNwN028aLE
OYV87kNpIErtRFOeFTeWwo9VssN4yhbXBP2F1E0O0gYy03UdgDIk8qg7Hj1aoRMBSobWP+IVoT4F
ZYxKjD9iJLDezwh1J44WgZ/Lg3WqOIj8doRzBG646+88Yqz8EL2YTL1Tg+gjYgTzeZIp0+5X79Ca
JWyIqWhRYHBuDfNpCi6S3j29q/Y+Jpbx9hOaOgXBMZB3459xB7ixHTWp2nzvAQKSUvKduvtFqaaY
A1YKkWRYXvyISpw1aUwT7YapFKwtwjgzb9l1KYOpS5iZLCMa6VGIEOMKFW586AZwgP3WeBG1EG/e
9QAfMwuTPsyYulCEGKiqroEv878f4BrhuB90kJYYmQ0phFW47yb/o/jtYvFMzG9v0mJMBD3C6ilV
OeVXUrpC//dzqM6b3NYF6GP0mtU29x0TyfLba37BmoNyVgKJJ7Gdsr9P5Od2tSg/hwrVJmN26ZiJ
sfwXa08mtrDH1y8LPgG9ltOjX0SvFhSWE3LOgjJm59rCJS32J3fgUpyY6a4qV6zfmLeOp1xlrlzz
cYx9RvVp5qyRk7LWPBuyCgZ89EcpkCcZfNqafap0c7U63kUvm6yGA7KQCF0w81aWndt7jNLNRcpZ
zuXgXB8Ww0GBSEbYio/BKYyvSAb4SifD29VKoSpSHr7PhfnVZ6SBFh8l+qjcfCfLl//BzXrtoeO8
dTIkyFk8N0j6VgUlEZtxQMNLgwGNKBaMp1f91rNk721qkm9OXp2jlnMNTb/ESDa6MxBsQ1Q4qYBP
z6sa/NMnaChLayUlbW/Tm3FZNxS1VY1NudTKDA564eKhk1Zvnram8WrYXoiCw7nUrtnN9Bfmm6tL
c9FApOsHVU9cSoln2sb/NEP7LVtWqq+z/fBtd3QgL7DCrBI8smNyH26cY4VtmoOhf/E3rIsCwj0d
WaIISHIPmJnz+YxPiBgJGzZO731Dcpa8bKNGrCOFFTRv38uJdMf+BLW0/8Sj4Hjp6YYadkRoDt/x
A7bUVhQuWGa4v4Q/79Hjp07tTX8t66RGFZdvbnzsoVqFFvy20omIweRo4NQ5CCH5F9vmM5MYT7cB
cr+DfCned1aqSBoxpFGJDMCCs9M6wggGbEWVOjABnKEZ2Vg9qREzYAsnbxKAtJJOo6eTl9IrU+VW
zCyHfkrnEbDRyVN2wkYNJ5mm9PaYhBJFXvkkDlIfsF5NLzy0M6ZymL+0HWk2+vcREkeQzVQ7drnP
C7dS4MXuy+KvyQNpQTaG7uJjN0p4TqLdPutt4vHcqIPQ7jBY0oQWN6rBiL/SBJztjp0OZYF7gWdh
wbq6w4UXHbQQ9ZZBY9jfg3l264MLp+rioRg6w/kHCC30crK0LCF2emicChVlURv9cyZ6Ip4cWcPT
v/BvHlbG8QUWD6rRzXc4jRdnk509q7J01+gISX3r0cCnoUkZeAfOB7X+RhS+38jTuTup2KXxriBK
JExD3bIIs8ow6r1anhHaM5yh+w+s0O+HLjwLhomtO0j4fC44Iv5/iD42SxVsH+JzfE4WLQ3kd2/T
HzM1bzCRWa5UZ3nfZv6tIBk+0xXN0h9Sgl4hbyUJvKPTFb1o4NwtsAq6577hqrQ3PKJRieyzuoFz
yE4DMSoU9zYY4EjYSZpX6poPgezrQlnvSx6IkX1cE+aksuUPvrh6IZVNDpIW6DlcmXez264CmHgw
SV4jD0RgifkVEY4JVKi2xZbxs8IB7vuxLK732bypWzSsTK3cZiqut+/OfBbkp3xImTSgleRA1qYR
Dcj9l9YxQSBZmLQDlxtQZtKcEu61WMZXnembSr7T71VWT52Wv14PFtSqbu4tnR48shmWvXXtkaM+
p+ieqWfywGBlBYuDDAVxRtFwrpy7x0sCQ1JEyU4f0TVY341Y+c/pcJQSuLWDbaattACunK/MT0Fx
UzKxVyoITiQ99m9uPefniAkdObKvjKKUT1uFabr+1GYnwDTw8FS2FVfSkNvX9umwKsBpyyYM9Jzk
cs/q1fCCPvjP+8z8BpF7Ju5+96rJzGXJMV3G1EwEcz4uBaaLfjXzoiOHTimxJjthXJ0FT2N2wPYP
Pg7gPTjy+ryAJb2za32BUTnBpVbaKLDf+yuiKvzrmNAu4/VhBvj9TiTOf/7P9uzUHqizFcLhdUav
cAgSBjU4SaeJvDspiIBi/l9H3GdYUTNv9fzWTCOd55HsVAuwy/ZFA7GZ5tGpKIurW4ukMHjCp9TZ
JM54H20rtpkYLaAomNCWuVT0sXz+g4K2l5w16a0Wo/vO542Malx+AVo9u/hyi9p+ZS20FLVySfeA
EN2UYLCGIQmHBRjOiL6q/TlC/kQBuLalbGAJqWkEGOu18eokwj+uCGig4pTOJZ3kuMFnSxEE7YsU
9STg/sGASX2GhPpgNpm/T8bb0IY0YzZ9bDgE5jXZ2RLFXe0tXsw+bpWECuDQg9UeYmW3m5a/QNcN
MP9ee6IXUGWuM+AuAo8ZZtU9ZGQ2ChaDLxHvOxZM0L3ip06DnUOp3FqSKe3tVqprxp7+n5CSaEer
uBMpFehtfpepqrGQexxX6ii0/JuHDVQomVSgnjn+xtJBfqjS4J6Y8NeBZEkzUzsFh/kCBrvrtkXr
dsqSQ80+G1Mpr33MKBbdlzCyEaPn8X87FvfKzRcKmNKfZFuW3NJD78Krg4kQIKSy5ioldDEAZ8Wx
rWYcgwlE3SUKbAAtWNO9npYUHtxkQRWKrN0ari6TclgODJqeZzd57fjy4uh4/k5QEVi87b7mIMqM
zJxMUlC18xO3dVeRFT0Il9uEcz5mBQiE9ihWzF6UmOj5/FolXJZttrMyI+tIDD4ZNUFjEfQfiEwV
zKkxbDI+CGCa9tCN/UyIUqi06ji6s1vK76Jvh1T0bSqEi/91iMQJ/+r2R8HsSlhxvXz8wfByXWz0
rffZViAWab25XwVrH4p6bYpL7tf8XCV0q0jHqb1aey9Atdq3Wy7Y4sV2cq4NByY0GRij1CgjlpL7
yGEzEoA+CkGOA5RDVhgdiMbiFrJVqqDo/p9cDh5ubVUr2Ejnp7wxzlawGYufITfXEdju446kHwGC
LpmYjEuoFiTogI6hV8OKZFGMEDZ6KitbFW59hSr3zkPXsj6irpTWOHvIG+9SLthCzyoO8dRkIEP+
jF83rAKbFrpzH+DGoMg9ozSNjF2xjiaVN2m3ZXv4nr+NpWZhHDJMp4N+7InXZmvcpMv7NQkutlnB
+ziRJwG21BlGTxNXxYuc4UuywsmR7Nyfg3Dbq9iCqIIXmKOkn6XvgGm/8M8H2ZAO82rA0lKzHkm/
2d+kUEVO/NKXfC1LbYKy9371y0iZ0NfFMPZWVKnxY02Wz0RtNJ1MkN7SifefUwjwE8kSUpp248l4
IRbSUqJ7LJNE6SuvbBWyLpLfc+c2kWmsPZkB+z5NAnlAY5WX46VSKWVR/n49Y1omtwYs38MDLKj/
jLT74d26qydT43uanS1e99OzwjeCtp1qT26IvpjXXKtM8V0eM/dRuVZzgsJ5GVbhFjYBRhvC3Rx1
Fam1PdRG9ts7U/9rOIaHwDkZNlqYaK+aQwHWd/hT89aSL9OYT+YWH3fkd/ohpdtCneivjPYAr7+i
4/ZQhAia5s+JpHwiQqmHqtgsJxXJomIYHh77Cd7SbWLze+SEixsL93vuRsxpS9GG4tFaaiR7nnlM
Vkhpl9k2FKMKPFxsPs+v1pbMVqSdUD31E/JttWHrkCAjp/F8LW9XXHFq7HN4+2VsGVF+zOteLrDc
cEHc3VxrSX1KKSWZdASJNp2YjMX5TSzDQ/FKjdrKitemRJdz/muIpnmkhjKaVZwhHJYkSTpyEoe2
hvizjeCAi5TWcPSDr4P5paTgTjnh32ayigvNAO3DTPXjtZ3/gaqF/0LthSrz4n8ukxvGV/Wk3dGa
UpJB+2QFGhsjct9P5VG5bVHJ/jIvK68fX52+VvfuJyzLCZsAu2pCmMfNXIJXlHqq598hn/veSsgz
1yXeY4KIPC8B0O3wSM/Tp0FaNrT7FF40KEsbi6xEAQTGZlwQVGpzisATZS6056uO38z7c2FN+LJw
nouKpORq3T9xwG0uSUewueDC/WiK4svq13ZywZnxjWPcMPpiw8a4BD0gp6KzHbZ5DXmn3F5LYAbX
9X1WCoJxP/UaLGPT49rFgkvI/M8OXT5X7fNaNt56LIGBG3p1WBY6kyuLzJFCDxqa5zVbebcu6kJG
Wucpgrc9HKIqbJPYqQ479svknf3HE8zob1dDaPDW3DsRywFFFXjy0Ixgkngy1uEYJgDgJAGCX7CP
h8zK/bvl0xD5ol0HYdQ+MTzvrIqltY7ZZKFrO2k25NbVl1FOu/4+2FUdQcoHxkJ/ARbp4x7gJs3W
ZjXs98r+ve8lbpdxBl+LrP9KrPbOgm+GbQCifeS//FqyU8b5SVtHn9AKJ3+LCZcSa8UOhiTX4jy3
jz1tJZLpDZlkWO6KhV4eeEDC1FywUVWBHIdO0G6RR2UrKSrHmq7XwR1JkT5loBYgvi9Mui6hrlCl
fxMB+xumrXgV/j0Dt7uPNPEOW0A1jIRV7pJjdtdcG7bU9lXLuYOVDCVUKrM9T2WhnQsjK+r5VzHF
pwovTXuad7wFx7pbhX8G92Il2sqG/hZOII0V4r1Uhr4PF9Nuo9rkqat/v1PC6JQjnAPSm8MsZFLT
uztvcyTu0s9mHFOeD8SVB1USkbfY+pcZ8CSWpZNobk21yvocanPqheQQtYogWIIFdS1OWx8tfoun
ZaA+TBxp0mPwKZBJgfl/ZVtjrzMwc1uGfIVfdF7Zfmd432y8m+46aSOrhkMoVfB6uqKZfkn/bgJX
yC9bR1FYwB5HM6G5tPwTjGan06Mvg27GaYeSP63IKdWQjWMw26QrYa3Scz64nTigZeC73R2U97Zj
ySQeO0Wbu/rx79T8oNnVrIHcZpb10UqkXdzoRceSi4+zZVxYQ57KsfP0QHVYBsENhASYxggkvBxK
v4SXbZNlO714j1AAMQr0n9sWfMkEDP+DpLeevD8sPEMxXkXuYz4rZzBQddhsEwKjabANAbaXyfPI
gqm4wjNd9ovgG83Nus3rQOZMjQtv4EE+zIcFWZo2L88f9V2/9r4qWrVfK5tE9qIsk6hdMxOaqJ6t
NNuDIaxtwwOoO9hM+HYt6RKIKJYpHN3K5rdhZKZ+Fi7gKMPc0iEUzak5QBlT/OdURMQxv0W6rYsi
m0J7zqGmi3gD9zLlu0UO3Q4oGZ7x2gdzyW1jrtjtCaODau3zi8AhNOSwzVdh9ulLFMTTOjUKKogg
XkovjZvaw9KxbzbXxulJ1qxBxB3CcD73CzLZRq1CPaDcb3Xu71PWxpiMmIXFmfzO1260d8HOr0sh
Oz62oiduglR/XOvnxPTXZ1Bk/EZqIaVzekrkJ2CKdYN+8kRLV7dOQ2/u/uQLW5jL0aT0TvmxMZ5I
Lp9IMpw9h0N6s6CeAPK8nnJDXsv51wjMED4sOeKsgfTlXF1IgyR0fC7CTd9g+0dsWUQzBAh0DtM/
FW41+lFiW2ncqPoFKvoWTrlUk5N5LsoGTlkpVaubbHpHdsFR2ipIKKctFAL2XDX4Dgzito7oho12
xc2DXRRGEq5Ilx2wkcVotZZ6bfOdcCh//3QAzlG1B+lF1ra0My4qC1ACsfd4rGZzwEEYDJjmuIev
1NWFEqMK9YR2pl4NlniAu3/g4NdsHO5sC6oo0PwFoYHypiMbLQJrLiTXEcKFK0k4v/9UZcpFg79f
ONspr0nLnLSTukouK7jvpadtjWx0kN0zdAridHTCA8pZwjx1JEZ6CegvCyCL9McPXv8WLzpAI521
jweMan0x0fUo60e4OW8VDbJOjfM6MaOhIlJINcWL/wEWFvXY42q59Qhyuz2DdYNm+uVptM93ioVg
aO21uHWYFFYORZ1PAemuqGcE6q+pwJP945vtzivsI7aeE6t/5TeE/y1F8kZIuN7nI8o597KlNTLi
CmEUp5j0OVbg4wCkoqMN/o4+NBFVMBn1F3SRVCIvkUGCezj3T+L8BamcuVhAlg9fxe9cZ+HSIG7G
UMx2IzlCERS1x5Z0f1S+iDVoIpH39UjDxO+/HQ78LT5l4W9lsUCwyvVToJNzJYBLFEXz71+janzI
kArlUBKzzYwGJXpmd33fRX5WIMB4wev+DAO9ySmsysKOdKKtMP98wXo8AAxfG+Wkbd3dNcmHepSq
D9fkJA4G1tRiQx3Gr2/LxevRjE/V31j2mNDbmphFbXcEwr23nmDqtUew7oXIR/LlZpOGMBnymdAy
dm0ZIdGCj0QPBpX8kwGLJyxTkRgIS0aUfu2yy+dfk+IHfEIZFdrrWnEgp7Q4K629eHjVt3IRLDGG
5jb4W2KakrAhM8nEIyu3qyo0ASXvfwFovpn2Z5XdcrRIJGHxIxrvm4NlBV9IHfkDMjow6g3neX/J
7VvHLrrA77ovhiHyFxzHdknqpzpFStpseZqPk4By9F2DCCwpSnVmAeWNn97O54w722G0sL3kV/WS
swaTB3m9+ynKCRZRhmJPjKth8nN0q27ohKAJ9CHH+6kMRTAoez0YB3AFHPLiEXXHmMZraLg1b58i
NjKuMZ+As4ybJckFyDSaU9xwbfXBJnxAVqkWOtNgl898w/Y4K5LtGGgVsVgtX9hUAN22PlccMwv2
SpqMrenaqLy6mYySGec+nAbpEVl/xt7LDWuxOzxV15bDT2vrhKfGS10FNfXHxf/f+8K02n0TC1Ov
nzEEcuHpqeN35GFpLwQqrTqfiwSxTUtuNmJY75lD7x2Eh8oMnGdZm4QknBVxVQpzot9AQJAPzMUQ
R9qv9qv4GDDhG9033iOuia6i5rWkwxKSh/5QiwzWAgJeKHCb5eoh2ZPBeBRwrRe3d46ednUcbsPc
mx/+fXMJrWRBCKvP/AB7yIar0y3zSOEX+67y+DEUHUj9EDbroOyZ3wuOkVTv3LgsjLc+kOsICA8u
HpWaYh2sc7476Y6J0xPHk9mPMTmlresSWNTLvKhE3ZevlGx8iAhVqGdoOPyooPLb5ROg1w1pAqWQ
9dWJ1vcXa94JqqVBsPhLeWmlt9zTappy/u9baCE+ajYgEspZ6jIifg9TC3q2/8YhBcoUuwA60VMG
tm54jA94ZTiOyI1FzrROBLrfxx3wakVeBuWrhoMaTM0j0bqWx7sS/0kM0gTyFetQ7H+emsxoLYom
lscm0d/66h1rg5o7Zv1lqIi/JlN62DAomygV8l/vdw4L6/poq+JG04d+SCdNb3bgf0N2cO+yz9GT
JMXlq4I5RcsyFP716neQuCAH6vZsQnKVNCTlGUANlqp4Rnh8mgqyPzXRxkt++q5MG+TthNpr61yW
AKbN9uNCU9phBsJoNxVkaofTTrahjFXgbFdoStfwsdFen9ocZWmg52vfQ0mCpxAieIEA5BSbyk17
RTLPOR+3P1gCg69YoN6+03Xo1GpJCj5/+nZNcDaIdyKNAGwVH6NfvYQDMC1TT0mGuCwlvSOfJl/c
iLWdb0OGLQjGAj59/pB1BoqmJEEyS9upq7AwR/BSmurqN3g/y5mmjRUrFWFy8mqd8vYMoyU4t6us
e4HC/2sAhsUYLhG3QbjrmZ6DMGTc/4bEN8RBaOy/bY8oC6EVVpVyMu7GuLSaXdxcz22G0s37dMLc
rb6GP8iODa9dh+BfOO2hXhuWhkYqLM/DuiIYyKdA8Gx89uZTvYLjjIcpyZVUtSa7WrT60Bt7f0NC
try55d92l2RwN+st7Bu3+qIuyNZFDXQR38dXzbteXy0uY+fzdXkkhYjfEyjTKdn65NmIM/ZwFwa9
upD4JUtW+SE4lJL9Mb3CtbXUIBG3895rYPsqRdiLSBoONCM/GArKGScKeRBA0JDxjZhO82yATCuw
hkLClU04CRa6AJEO/QgC/q8rL3uiR5qmUwyKuCUvan8d3g4vjwIrmPNS/O7gKiwMl8FdacW4RFg2
2FTB6jMRj8MPkSqKvgeCwLHNsQZoCT/5lG6g+OR/gekgW2DtRoj2KteF4W/XsfeUIpiXfwAWVr7m
yr6eaA+BzxMTFdvdC2LIeoXE94aNjh94vllRHT5PAgMRZC1EH+lhtoL9Bd30Sear6wCWBXZlECVr
4X3IhnFaehSMz4484ZLrIYWtmW01ftAmFvm6PWAale1T7DaGJ+N/RsT4ErAhYmDBIAhxikuBD6XG
DQyMMSEsycQEBHDUHEMpFNmbGJYvxvNNqWEKnXtAClKF5On4DzpXToaG93M9ITePLTKQc+240E1X
fSmHXtNzM8YNMUqtFtBrCRpF9TQGVppJZGSMuL4r+VZowPo84JvRFWoPLwU8JIcNFjLfWYhiT/bK
EVukJtQ4+pvFC9R42XbJ62vgZaE5MTfrWX71LdD7G0Rd7HzmZOico9MTcIwE/Hcm2Mrc/cpbgXE4
uOhwVkDE3rPIEAuZ0wUcIjcCLLC6+vyZelR5WUj10ogsteV+2W0eXc4K8mXjmhV+bZ8xYTa8x175
88WY1Onu1BylkKJwdRVwNyq4a7DtN6Htoz+8iOtP/+mZEC+NsnS4ASE60EbRXMNfJVKKuQxphyZo
Ki/B+2WK/qQo9A5O1QZxK8M84+y55hUgjx+IyWl7Bxbs+sVTItqzGb7yAh2vJGcPYwE2vl7o3ecD
c/HiMd2vB1Sk1U8AcrUCar7U0rdzBQNaPD9/KkTPmBQeGYYmFS+EPWuCtuhnmwLwGJ+ZPRQD4YlY
ztvceXke9AaJuYn6yS7qEHesiOUCOrGbIUu2GykmWM3IPRfE8ZZYnnjfxaYOeAr55eOuy+iUhTFX
5ufayVr6+IGFi5f9qB/BmvpJuz6ykdlcVFrnAIK/ELwv2ijurwfglqHvUxfoM6EThEzTir6ozHfv
9m7zUGddzfGkwJ+9bsa4sQiJLatslKKf5rDJa2oVQt0olHRe3E5GRBt2mYbtXBssTqMH/Mi8g3IT
H4xOp7RftdCxqFwHENDkwsWl2PGQC0JdXu90MJkZliNLXoFhIqr4woBjvF2cvf/eVlL+K74b1uE3
tGIf6eo6oGILH8lZaXem9n54vbFJfsJVtACFkSYJtG7SIPvA5gwhr9R+a3WiIMBvPpMTIBOubnDT
Mrr9TJWxttu+Jedc6jJximLX0C2h9AkkYKp/ngrU1WcHhEb4RPyI/APL3VDtgnltNK8A5E5Sqmar
t+APiMSnRK6ZcO0jQcAorUPLLdSDQPUNhAlTAoEVKRGHZvQVvU453iXBju3SrErFzLvGkB/chXvM
dzO4sCFMxkENHWqUAA73pZbKiJv3agNeZ7VK0paYWQBjKMeeatEzh9rPToEMjmfWJ6pYCGnfPHI1
H9b8gfSBZECUi83i1NMIlIXd46Wzn1BFyZse04hNuCQHCudQ5cO42B69OWsxhFAWfcRk/l8aSkR9
CKuwpUhtJM/dLCScw8WQ85UDO5Gq9qefWzPjdYHkzIzdpr1EcdJrwqQjr0qDiux7ByUM8glKH/rZ
oSSMTC3IPow27uz+uXUiajrzCLViw2Ysur6/RdEbJmEUT1ecRddrcPUGNXeeYLk5kwqrRANtKCFJ
m8IUpM+UhQxp/KT7v3DqJyMrNyDkPCat8NOB7EfGvpywv88gIXithit0oNHp9c3x5oOcHqg3xtUJ
sS9KmMKNbTVQcMlxXEg39K6m6cBHsZ4cDtQpzC/VoYTB0rlySoHmgQqvAgnvl8RFRn9f60WmspG2
DuGJzygl0eWS7pl/ziuYBzopQHm2FxpsqcQYeatnpVhfXZ7G68W/7OPZIkz0ZtJbyt8EkB9jpHGR
vF5u3lgL4+FVcZ3dbnQhmrNN7hejuENHAz9+ktw6FUzP8PtCXroaGyumFil4zCzciVkSt7rZe3K/
KSkMzGcD73SDWyU5Ax1pn7yGrH1jn67MiHcjYTDREVZT7EBxalyR73RyBDU9lE62e26UmtYvraDr
ytUU+tNYCLAvnjxAdqcgZZZRjhJiTlek6R1k3ThuEuCFUIaLIibKsBZEk1prWQmpN1AMybPqKie7
arlfj8w2M1FNnltO2C8ir6PLKSVNh5hWYfOTehl88WVa7ryis3OdW1g6RlGSCCmeDEQBpCin5W4x
1u3GlqHUCdgbiCEBXAYhibPfiBA9bABPN+hFhfPRZPoQljd/n4zg/q8CsqOD3BPQKTY37uhkPeC3
zDACbu0ShTzzTZWpP6EEvBI/di1bySX3ieccATXwFSkYQ5gkQdEuC9ZFdmC8MPI1n3gnuEVXDTHg
P+8+4RdAgz3gwH9inPGtdnOwwwXmL5dfCBGlZl/kAMz/dQQE813yyH7hEBUdz1c5dASy1y87iI6n
bdpISZXz8yUUsxUXF14J9HAMpFqN3YjN8+oSMR7VccOA7e2fEeB8zdLGt5RhoqbgUPpmcYpMucY9
rKjRQvw08SoAXx8dWlRGswENM3R/pZ49ntDY0YTA5vyfMroxgA9L48fFeqLsyUb0fjYYGfcn/+Yo
EE0k/gF6Xpet3kOIQ+N6P/Dy0fIBaxDgnVRmjqEvBHDSx2U4Alp4W2L6giIcSv3du5Rh2mZeVZKz
7yw/khXw+PVPBcZv+DrHgzVz/eOmEPn7ZjQcMAK06KUUnzNbC6A7WkmMsoZYplABLc94EEgdcCMJ
rbYNqqswkaS8y9iFU4LMOphmCJVCTAbc3xHWxX2bCIIBz3H+PNX8dvP0yR59qb5C5RAicx0erXKd
4/L/7cWNAY8TK83JAsNBVt3tfU1NzumyniwK/bOu/uOdLPhje+YSWkFoFEmhF/UCU8tTW6WgcInN
NHp0zDOZny0NxxFQM3FnOIXrcmKhHXH0nQVp7pS5uN/l+BL8H4vOmKfJTLZwnpQeoeWksi3xuiTX
3rHh/tMao9UO//IzIzYfxTnKfp8InZkPg/3aIPI7BNItrqbaRUgoWFdJJWbe6V4xxNsuYEtBe8mX
39+/kV1m++ASlAVMfwMkVvZKXzQdxiJbUjCe/lTZSYnFyP1YpYYSZAJyc8g/i/FW7db1hQU+GhAg
DV9RtRyW9Wkbw2zVcKcrc2mmBzwRzA4CExcF1BT4Ehg867V1wVG3xJlU+qzZ8u7tsiVCDjg6NR+f
vSJ3eezduqQyzxenK86qvIziKHwoJqJNZt+8J37c0DUTvx0dDqWn1AifDxKgtQpsf/v+8M6OSc5m
UQIJb8Gp3XmM7lPXYlGefwB1Uej9KhNnt5ZlFlhK4A2gceEKwKrTF4784n7woLMmqjbFMRsw2BDX
B8d72VV5g641QAhbbhwc/vElLIUH8phyVx1OjvQAfupSB2tXatHKbGMJTssiXnAsenSOVAmctLtn
n5HLweHVX6aJwn8mWjA2Lp1i4m6Z3qUomw1RYMSpsirZujyudiVNpjJAv7csHgfi//Ry4gmMObp5
VaiARproxNn5T2GAtw/6FiyhzY5HR1LRwr6zUhJgHyij19TtbPOYdGVd48wodmkOhIC6y72CGeql
vfnFf1xCKaVf+phIcqsrP+uXQmMC/c/Ga1cZEp1Db2e8yNWxj/ztKLgfFtVnnoQ4PE8pLVWjVlFO
eemMbJC/e47KuUV0uMRO3dUoTXCYFMHMKka2/L3tKsV0+JNWnCrswl7m7/fu0mAP3dRZQgXXcubP
5g37hFSK7UXphydBC70C9ymp2M8mxKJeQKcCSLw0PEzhcl0J2TqbaMewdbJz6Jn027M1OKvePp2n
Wa6spx7QxlSAvRWBoLKMnBbTmPNfyJJ6evn3RH5A+SKG0V/SZEOSCImR1rPvVZCfON/+WjM8BenH
KdVjLdvGiW5xMXguaQ0spfflj9oPOVHNI7TCqdENSbaTtRfYnfc7TCqVRA8/d6fXQ9DIFhFDjmeA
8n/98Qkwha5l3DGz/16OT5ZB8irPEizVfWznl6tg6L8gQg/mDVAJPL+lJ34YzML9u8aJWU+uUTeJ
bOJ+2h74+3j+uFS4FEZsZCWc6Q2p4t7+Ofb+2RuILa15AzWtQ+zBu90X85P7bedVEYKY8lfGCYPN
SSqDRvD436V4yE6TImPDAfyMTPe0NRGKVWNdaCrLSzqM+1e5NTisD4eFxCi6obAtJ79G+iA+pqU8
cmbsTMLPLCKnpaMaP1abasI+AZXG63o9N1ha8SQGvKGiStm+YbljYM2SbRNzj0XyDtZB9hTuvWlz
+f4xwXbHqoH5zuLDhCKpwapt3QteCbW7J+qMvey5LYGcXF6VSl9jbkZIQeGiWtkKfouH1xEAal3T
N7czJI3EPi/GhfQmMp2/3JA6fs53WiJQNDgWnWCiesjri3sO3UKhu0F62IHbxW4cFR7zZWoYGhDE
1S7bz6Z+UvcAd9G9UBzgKISuU4SGW67SZAhdEXsN/c8lqRICX0nDt4Ai0YxR3eItiUKCVI8TKny+
21sljvJulCLW8K/S9hPKnfgwR08HTKXoS7fNPfq23A/E+E1IUQo/rMZMpCi/sydzXZcccDKTUbAq
XAfFhU40HiZFNS1fesvf+BjrpI5dFjV5fwPlzMUNjHHquFl0liYBMQjgWOdL+C4hUBBxlCeVCIAq
P02+iDFCnaVbQA6mTAmdkHayATmonB40U+JXg4Jsj2Mv/shXX5zLVAckvBghLTr/ONRXwMEa8HUw
oWAm/61j0CdjkYFzGm/vloAhVC6m4QS/6a1mh5fbahr8tIWJFKcah0V5F6AdfL1s51V7c4uqhHzE
ns+vz6yi7Q7GtUsP9cne5QZ1kLXh73U0opfYBjKfPgNUx/Bh4IuqpujEq5YgeCcDR3UkFeqGVSsk
XyBDZtFL1non3GiK9ZYJe/yn/w1dcEmTNGg7e5EGgTWp2SVa7Uri8JlO5939sbJE7WRL/2rJNgf6
2SB9HrLLSTp7i8+hiFiZrXuq0y1f6L4fc7czPWWZK6ad2BhJzCbRbo5IhbxFLL92JEsqPqJSjvdn
Qsk3m+GNbFUAWmZ0j+oayAE62NoeOjIJX7sG03XagqDJTU5OJU4tsBwTybe/02DDlwzXieXFmiAg
dUrU52hdTl8MTvSzOVek+qPPooVI1bDdEQYSJqcXsdIArlHRDToL7PoMCeOg1B8gQyLW7blqccQC
pPNB13z2Qmape1PwJAiOB0gjhHdsxruCUJrEzT9MqrurSsySWiC5SpaHM9vF2GEYq9q7YVQuKq/b
6NDQYiSM+U5x/9xV2JNyeHg82S5ajzRx/DD4Vwaeo9rrT4zxEOhkDt+vHT59EhaqjtAsNeLL0VLe
8TLnx7h1IucKIIxKWjNOC9g6YTUlvIXlIOd2Q83hlPTqSW+m13nkxLal8u2/QBkHFph0inErllyV
Hm/h1EbDDpd65otU/wFhg/Zopy3R0OTGa1hkJ1zo9VEOw9DOpAehEqNDlnnvqwYm1LAhCM6gDyRm
PXLUs05VryFgltuOySbuvg+EUjVjb7kalH2J8ORS7WuomZtRKn3f+sLOp9lX1DYKdeY1wsCK7KG2
pKYKT8pJhaHWU9HMhcXnxulXvD7QtLWswsbMpg5VBFoOqMk+rgxcdZ86OJiXF6ngJfrnX6Tw4qKe
vLubsCkqWjREyHkPSBIb/VC3XbabYGTlBn+RGfY7ekG0QbUhWJFEJ//9kcuqM63e8FdIdXrLy1f6
5t7MdztH7cVe4TUQo0JSTtb/Vv9ZuLHmTXrLYYXajHE3hMfG8aOMuSEooQPXF08RbYdN83l2Mnr0
LbSOBtToQ0VIqTzPau36Oc1gAmKvacYCn+2IR5sJUE4FkOpbrunRcy+/4G45cpEkzVUddPvfqNsg
JsGubkESN+mtoxcX5ncO4oxE+flJujqP3h8uWqzNH6KKDwAUWaqMXKTgWHv3gZe9t7cqtFhFJTo1
Hm3x0JRKjhQDI3PBpM33XS/D44ikv88LxXS14P1OO5rkIYVuEnAdWsA/IYQMXnr5/SO/b9+WGdsS
FFfcr3KJ8oQc0CBl7N6D53/ql9pxP7BuYWzYegh+XGY2yC0mL1O7UN4ES1RFLSGHGWG/s68NX0fv
CFMwEprYGKGi8ZKjq/r45Gl/1vMca6U1AVHV7KDFZcSk2naaIsOxdtXAeOhZLv2C+7vUxj3aDr0H
aEDK47bFxyjCLtsoCh8KX+TF1bFlTV2wfJ3MHXvwnMqk9BBciH2VaIVW2iTgHRMLt6zAEeThFaWy
K19fSMvzMoO4QNRikSZCbMO5t24HIvMMHBEN/yG2wRF1jsnwjro849qEbkiHoj9X7T2B28FIb0tD
eq9OXVyVzQtjtSyOKf7y5T050C+5LDg9i18mCuDOoop/BUwKKHPreL4+Xs+msGS7ZW9lxTZ9z8vD
YulbLR3OBMoUQ55VE8iGxJDbcLknlSL80os9sDIMX69bWsVKWglULPaR8/O23FZt8etNIEyRFtAb
fPj1FgJg65Uqqj5fBO8gqXE7hrTWdlT4gGYnkMq5NeHjVQ2R9ub92wXBGoro30gXgpiBNDZlCmUv
+OiC5wIDJmT0ScxsBGTLR1jz9Vg5R42PF2rdj/KxTAuSG5k3TYmM6aNhva5Pm6zQ9PHASvTI3wmn
wrJE1GK6rwS/LCSOWiGA245WL0i+KumBBKAJECoJ5zM12ZgWK32ZZRBhujpM+cM8Gdofq6RGM/ny
HEQ8Klx0MlbPRHwWbTCNTZwnfIM1prsF/3ZIeVZOHl/eUIwFijq7VDve/MnVpQLtPuKnZcMnriOK
Rj+tqIHBS3WeiDPWQRvrT75j1ilZ1Hd0lvdklJQa8OfI/MokjwP1IDKF8o4pcuRrebWereYh5wOp
dewxFh7BsZiPr80s19wkYZKLb7r7JCBm9PWBpJqK4A1Qi8mUdg/Jm+uJi2gxuy0JGux6u1Z397NB
kptPdtqI5l6XEahgrIu9G7Yx1J1efv8bheDaV9Ea9Cio0wpmGkU/rbXdYAfvM4Ee39psWv61l6dA
6jLDJk/6gU2Fylg11UvFkv4Cy3W+a9WjtCAOc8ieqMr7Lav+unHHaqOl1pRhKF7riNVpY+4i63WD
3x2plx3H8IY8EGbWR347wim32tk4oMPPMvJTjOlZfWAwu8aiav31MlA6vzPEt/HVMVa1CM/XRJ2T
sbR+ETOgVYb4A/Ocm0FoOhFATNQuEJ0nd2xl10Ys5A68pWNaZvX2qULcalvo14QpYeH/fY56FCoJ
Q+1RdFhzbq8m7aVkUwf6x1aSgd+MbwxJiboMLLMvcZj+InJbv6zx2EdXIu1U31m7i/m46qB0iIOh
mFzIey1+zcUDmkN7SupkMpf0odfvb/KX2nF3Zhye27n4VKCadtPBBjkM4JzEes+I/wK+Tvo4ciKd
9GZb2D46URaIxsoNIOmn9Dxx4+m8gWqMke/wGT/TH0YpEWFviAH7xdxAfGzlNw+XK0zFT7Rccu7r
WijDZDaxTmNPHyi74bieujDtvKoGohijrMgwIc8W1beQg9bitt/GAOt2isFnn92liCs+fKtPT07L
9K+yrHxpP/C0HP8fcO/1hlo4mUGr50KkeBvpeN3RjJJOsyy7PtV1kwXjI0Dwh/4vGF0aU/ArPRUk
tkLbeKBnvPlQXJgjwE2stgE5C/eK/ixk9+6ge+YVNJLnFhZEXwlNyatWha4z8ST2SUjWuiBvFXvC
bnzqaJlHvm0GsEGXnpPjtgyBJSI9gYzfo2+dnXUYQIap6Xc73a3J/iQTU2Q+uWAZ8NIhaZpKHzdj
qORgHm4AYsLEioNYq8gyAittnCDWc4mF26pS8sythHoXhPGui+nez0OJ+5acljhywsWO3V7l2fpP
aSOpl1851k5/Yul33oKVYkdcvqDUlp/bIXyrrpaZjVEPHH0mh1gWRsau8NJF2S4/fi0ziwWaLLdg
GNrVF6V4pA4SfAxKwDuPS0+XxgyHPHp39qZ09Fsz9Q+POZaXY+8hRDHuVjKRwNMikzpG2pWYxhP6
ZGsED/9lsu/hLHls2mdVm7M+gvHBQWnGxwUJMDbPRDaloEMzFNW8C5hJhGvs2JnKNPY8DF0EC3FU
wLNaRXWJFVnYGY3beWdOgdrZ9pQXeSLpbEmYdn9qYgTcxrGNnu9jNoXYa72uLrdfrq+ETd+4Ovbq
F7XzheVBqEI9/QB8jnTUqIkvkVCMogbhVGftmPLs4glqLElSRw/06v0tR2/lFINcy9eTj9qpEiXd
Up7q+mKDlX1iPLfepwLHR+xNzqOS0kOIYHKNpRuntw/yoQGZi3K3mst4OkBSQtLWoEChYjqen7rf
lA5Pcv+v0mLAx4Z94qPtdBh1C62uF5YPYqXgQdK/VZ6PIwBKS3pePMmLxdnhz9U8eUAJmRVnqLQb
AVFH9FQrjFT4Qy0V3RQk5uLUouZL59BIjubJycShalInrlumj3tg+RUjpr74gMKMO0GyfvlDdMwh
YvW5CpzEChoXtq6RZzYJtPvfqq8SILcqVc/gHW6P2smRON1MNhjy9trXDAv2an1dYB2/JGt+NUp0
SlpdUDb4JP5jDguU09F0Mh8e3tgan97ruYHj32W67baQQcwWmMleOei9u4LnFs7HciKPRFw00TH2
2iNovF4ZL8ymd+77NUfuiuNxMOGgCmx7KnauT/MB73XpeEZESw7M26G7Y9jYZbOJk+6kelZ4GXnb
6ST6H8+UbEUggWhnqMo6af9UNU/Mt2+epjPEeXi0qStSluIT7WcrteVwwlRtRJaw7INXs+pxhIWe
UEAcqXspXcxOhFr8AzHtVKtfqSrHGKexHIhX2wZ6DJgn6C+AyKjvElYgLrJ4CWNMsxaN4vh6I5ES
r0dkTKxkOdzfUce/Zx/AzQXCJLVG4eNcg/7imACmaHjgtwnpqLYj2VgDZVsjV20CT4ROkwt6phME
rvhc/o4UrznqTCQHe3Nnme+jtTjxbmP09U2e6vtlh+s+bSp1Z9kb6WDNyOTI+iSoiAGh9ETKa74e
4FjkHbVF5aunUxSeepS5nqIOotFM058NcN7pq+V0lnFIzHqjaBcwinhg53I0neEyJweLDzx+059r
4ALG4GiF9/D3AUwtobbJ+vX6Rnng2JcGMkFRr9ftxhS0BF9dawdUK5Ypxi/1GsqtAXHa/NaQ16Fj
043/0kQV3u5R+1BGmvH2NYXAAFWgER1bn73uxclq7oU0cxjhf2wCU5li+sDeA9l7RXlv4dclvyeq
L5MyX1Spf9QDeWDOIpgzRFJ8WA3jotDRllwyumsnPP1qJS9OjbWIJKjzBYgW5gOeiCbQP2MPbS/I
XZFKto3NOYX6wKXJfSVSScAKQYCHT0RH0XpIXnpj8KseioEiMMR0mHxD9H3RzC9nckdNyPya83Gz
LTWOuxhtfrPc3VDZLD2017gimex0DccpU0FpG7xv9laOzG3NmjjWtAgSeqLdU+n4KiR5ewUtr6Yj
3fCA8+GGomT0Sen/S+IRh7rS9rvBnxn7gUgY/RV3aYiPeEPqozpRs1VpEf2BLO91YnWwPY9Vi+Cf
yuTDAYLYZwGWoGEdpkui5cbanqECEjlvk08NeFWEyXRDNy1ECDaXsKsJLeE0H9I37/IAFE9mhrpU
z/90RNFtxT4c6mi+nhzBxyMAhy4l9r73BNm2uoQkBAF8x4ZSuXNUlB7C+X8ovC7NyPbtUUfOHtK2
kDhrNnEpZPjhSB4onDhk7GUBksZT8mEAADGJk8EYGYpsJEnLP+2YxYlljvcRJr5MW5mVp+QKlGuh
6YivWjA5wLshDPV8bicFK+C8A39lQlRXXVlWKgc90DSzSCBDq8ETJgoMnl30ILfa6Zz3Z263FkMO
vvMrpVjnA7UinOz6+ORQ3oEycj/CSB7rF7Ua7sZrqA8RQST3yssztxtegqf7N1aSvKg+kCN+l61o
+QQjnSpOCCr7KROs4Mmmh2PtaECLxx81lHeQIe1FA3adpoZNRYaKPltdc1feYOmu8wJUiEFehUDU
YUd1KyC+t8r/U+mndPFxVKPgDovBl6QZESaO1VNcwZ4wa+rixIxBJVKvpeEGq70dFZkPNCX61ozw
kcSRPJtY16cUszGPq7IhnicR7IadmB9bHwurEVW8ff1O9MgkpmlafK7y1z0/miFtfbTpWgJINSOL
ciHW2q+VNp3Rj5wTxpLju53QnpKhBqHNp5WPQOQCPuX8LZdakiZyKa+qOScnQiBg0z5SRPtTpnEm
CyiPt98YiYIn+7c/5m1dRir+tlH7Y5FMBej5oiQdVXAf2j1HACKc1JGWUnY9gIioZvtlCWo2l99d
0ORoYeGgTgbgdaxEXI2aYuJQWisR4sHJz80/7gD6fMcW6Pc2xrdiPGnUPwHWdxAxnM+yvWAQpkWS
bLyuaD8GHJS0hZyOIoDL0FgdFmA0a3/f/amFt5aV625vkEpRwjUgI4kkKuRUVNd3WL1Gl7ZYf8nD
TpVU2AXbdHcj5k9OkgVxSnzLNVehw2aU0/wOfCENmnJ9Tc3bXsQtbLYrQz/TTgtfa93rxxhiF6tQ
vCDtCNswOl7ZcbECiDneOgi4lOJk7bKWWe1Zrn9fnTu1axg0LYrn1P6/g2js+JW9g9G9y+rClL0d
Z76XlbxW7RS24irwv6rtCkhwL8gXMuPJBQSL7dA80n8AJyHvfrckjUDrxSoMm3hmc6xEXLP732wL
94CnhKxn6RBXpBSsBQh+CLt3ePtRYaQTOce5EcN1BLy7w+oEsam8mgu/GudyW3WUuz8RWFYgNYsp
7cLD+K4hnleRFFkwwOWgB8ls8C0ofmxNYKVLzk077rVXSOaXCbLk4DhwdqXSJq1XGp1zNE361oyT
RNsYbjyGDf1pY0t+lo0b1+UZfV2sWUcwyMQie+33ZFCicLBIOd78IbSW+/EwPFoN+Y5DM4UQta1m
v4X/ICq6BUWmAcxApWKhjEAok5lDD+C7kOeClceqSBOGcP3vkOs96ts1cx052iQtOuqzKBznxPPm
jK3rBK2AfQwJv3hzRjfBkMdj8obq/Kme8/7mi3o0fT9wNs69bVW7A2uMWqzHvTbi4gJ1D2ZJEMjK
4oufvkCNxPxGOztTeGkyHlR/eRxGibJLGZstYCksfMPbYV4fFJ62bJQTD/1+PGGjhYJiUFCfZqhD
FB5Mkkq9iZMM/5NfJwZ5SEC39WSC3rynRaoV+6e2q7dMbbmjrJ2h3jl8YJ8o5x/y61Ofhu9z+0OK
NtFTIpFkrsLRvDAt1A0fsBK5W7BTARAKSeYFIpq34DIdafQdPsvkdN69ZyELbAf2ldKMQb15zdUJ
kcPq4dw5fgYZuo8gfTkQ2JqlVgViMOtzvcEZUYha/tI4q28lVIaF2YQGM1bI1V27sHy6RFO1eDRl
eDHxrR0Xa1qWbifxdqKh0+zsadFXMJB772LynauItpB8fQvMlvtazT+1pHnvnFCaB0bhS7yrRNok
vZCK5u3HphyRuxNrgTISSaB9y4QAABbAZcHyXoeMcwVPOPiPg5gz1nH0U2PhsHAF6bvQ+ZdFvkOD
iZonNDqEm8NMHizOBfcLrEuwR1N5Oe2+3Y52km6uyJAFZ94rXxnDSOr03vLKnhYTwIhbNTH/jbSS
P8V0cc2MdgCEHyVkjh5tFrlZ3LZ/wbAepNi6W9DB59uD1M9w7mmfLB9KAiri1yH11G/dR4VRes8X
ZYkHYsMoQTFqygn7LG7tTpdZhuNIh6gnutpaFMfIPx1Sht69DH5ZSWdT9NfiCIdyxyn+VeU/RJ8H
21lwniRtCLM/T+3Z0Xo00cLG4G5ZtdrOmoXpCYd4iGvNEoCVMGcVjSxzyDvL8WYLEXogmK8R4hkN
3tkU1pOYLxwSvYwxBX3EpRq4t//3jvZnqyTNt+xgoWnEtbADUKZsKKw8QjVnpvVPehe4GYqrmzxs
KG1X9hMJ9wsAj3KD8FNRmUPXiNZdPMxjA7414r1V5Qe0onC4IQviPjHeErpfyMV2Ah6yyyoQvwlN
A5P6pUhGkQkba4JjAWzrKJCmcmlH90oL3czCOYSy9Wr9Nc8i4FZN47Tcc16ybVDcNHg2oc6wrZd4
ySBzYsqvlimQn/9uIaboT1IMt8lSfjMX0mMrQnglrY/JcYoZq7ymhOWP7jMyT1xIAbXFbu991Z0F
RYze/cOr26anUx7KXB9zeI3mhu+20jq2IS4RkL3/Bjjlnr6YyKQhZ+cGfPPjx8N6csMmYJwiwZEx
xHH8hTVS8nl0o8ylEZeJUIXJ97UyoQanIxEw7GYR2weF3IqMhgIdgDS1kIgghxY5srOyMJdLobIY
rpeU71aeeBvoGta79qhr88SD/VUyvLfOSQh0/pfHizY/jNxRoFu5G9iC/rFV7vculwCWOJEE3zxM
djt83fgvB0BWXq77K1lpmOQ2SBzylSYIwkzrGWlrqDmP01UoIi7UT9i5Z9fftxENpPRM5E7T7snZ
WYEM5VLlAUcMeWlNRWyBQL4URQCq5RL6KfELyB+9cS3ijU+PDMDu4/O6tsHgRQh4aRV3/zQeJrBK
ML4PO2N5WJGNJMuYHMwHPaT3NPUSMuXY+Wzg8cAyF9iOFFZnG1cdyeNsHw5eDc5bgLBMBOyZe+/F
/1pFL3mXBDik+WB6i5uHHDBgcK1lwvwKySq6mwRsC+DGT6khWh4LHJrRecO93AmuEg+3+x1p3w7B
OqUrpn69kz9XnIUy5j/7xu9jO0N1UEp3I8iOE4n3KLSA1jKMFb93IsLO8RCTWJWy/p8XGVs0j7/j
k2K7UC/t9bZ1IPVlLCq/6cSijknhcL7DmznudZbWi16ECtSMiGFq+g0b2+1ENQR7fz6XgnXF/PTE
9R9Qo7KmeuUG4UCtRcnNZfW2fTRdm3lzRCoCrVVX7HHOVREk4Avd22LtkaARd1e6AJf4DbKLjQnT
6WhiG4zMmYFY5X0+s/1U+WTeY1rdaeZlr3ijfgI38hcXFQ77MFClotSJK1bF5eXJeGCU/JrLvVGb
ooMht3yWXEyCNaqRhIFxuqKnmpc3j+omhi/f9/utNS8xTNg/ZaoVFuKGWVFffa5kjWGnImq+Bxrb
QArsgJ5ZDZjxGYJ6rxjZ+ilL3SJzJjSPZz8OZcPhzSONCHUi2l2lJBF7J86/HcZyCC37Neuuss5F
cSJa5NKtlN3GTH8mHxBy6ccj3rAPSLzdoSYDNby6Kl1ku8PNAPP2jCuCjMpjlmjS6kYuri7bA5fu
xga3To5kJyow8gtlFEc8U1W6oKVfzdTA4F4s/00zoHgqs4BxJkTLRctE/peywbu4zsu8f8Oh+C/P
N3TTodSppr4N99gszt2epBXo665fldiml5KacCI1KwEulDUif2NH3TFHfWUtz/muzG6DZ4GZvZSl
pt9DyGLr8Jn9yGKVUgVUqbaEfeJr0tqbkMJuR4tinSlEH0WmnnSTpCtTM2v9/65ZD72BLq69wYSj
kJl1UtVuIeNsjgfQ5VOKAsceDxMbPF15zWlHGBy6e7WjyQJAv+8/YOj1/jnDpQ/gpyxsbRA+qks8
HgiKapPRx6cUXMJtnvsrou5AgrHvYlls4nCg5Dlesc0D8voMmnc6RK6XhHDocBJj5bZjEv0+sh7m
vbYqvJ9VQDj1LX061AIm1ECP8XI2405AvvqjLzfoN5L75e/bY7DQMbG7x0OSrB6rAeofTHNPLykE
rMt81ln/8Aw2cZPHSnoxegq24fbZqRqFv9Xu2JuLQcXiPSBrQItRPJXbHNXDnQmGhtT3fIX6N25I
AkVD1Lox8RvN89ElVJ791eaaYiarSWpWQPYk+dXsUePftqYMEq1rCa82jYedSqfd3ZL4hcO+nt9B
2BrCSXrZbZuS/4qXP8v7KHaiaHVparFU96edPreBMKi6MxtSe+UwAO44X9ORMYCbjwPmdXGRWbPe
Sw1zNTps39vH/8ZUnb82MjNKVEJyyGa4OaI+FSJvP+O64qHtUE8Nc8KIOYOjBXI2GePdxRQAogeS
eQFdJb+Ykg4J/Q6eIt6BifCxO7SYS/FKeig0uMeRmDZ2p2ANFbG7lRGw5W1ysK34I7B4hR5gYzdA
78oB0ml7a1id8t/6G3QZCpYq1mSEqo4gcyxcAGbzQDlNPROwkzR0ap/73Ew3uK5ukA9hj3QaWtGw
52QU9EeHdBr7UixqpuTvZgZ49G0m2r0HLs9buToRKO4MP9Y4N1Y1yRuu712cSDB1S9euCuY0xmjM
9obh7G8S+giDuVt5e+D/0YVDGQyKSRTN4QNVw2SrL3tkjVUMk3Hm8O8dS2jK+U00qZC4cSgyE+o0
ddmYiW260ZMIzkn6TUrEiGpIj/BxGC5ijDkj7/QRNefaKyCbaTxS7P2SbniF9lAW/eZGn+cP2XWp
kkYZ3Ro0IcyCl1vk3vIHWtaAVGDmMTqgal2mXIqJ6NSM2aSCesZxapD1m02J2w4gbuNYfBY0ss1B
IEDVTY3mZCTzMJ9WO8hybS5tML+A3VHpdIvlzzRHWCzHXONNoPf41RMEORpd6d3OSRoCOQMNO15o
bLyw3yYxMvLOigkLAelXh8w7Sy/ivxgdrO70Ix0rbFc2kl4sibgLp7ccm+H8+CbljAj3j9StySXa
TE+5bB3N1pa0V+6YbNeIwRS/0sMd382bawhkj79L8B1F40515CXShwcMYCscDzUnPjd2vlHZYP7M
MXlu6+7v/+SDlmophxPIRT990bUMyGFLfhq47qgMFf6UnhTogoBoCK1ILeNWsNCYkBSL5J63DWq+
Qy806OeaR6liLmPxHYt/N8JeF3P9sZvaimXK/jwN4n241NtMW1ueOOXB4VsbX1VOvnPy0lMrxU0Z
1MO1sI8BIF9KDTP3TuTKjlRorHjzQDhLQufVCdxAaUBlfgQE+YM2FsFfhuz6TRvhXwf7ZpFFjyVf
VCuLPi5/LdE+m41XYLlxFQTt9b0t9Czjs42tXcXBINpRJWusGr/lMAOl7dsZIE1CoVrsClUiuEN5
+YGwg1RMgVVbqjx8auBOzWEjIE3OHs/RqAGZUlnv5OB8KmAnC7zUrF2xqKbN0xvlAQllyMw26pBh
xcT/2+i24A33X/FM+RwDAEx011eJ/SAhOevRwkGCzWlLGCIb02BCwjiEqitTrg5umKiqP3BWC4px
TAGkvJPdSitGc5DBWHR4x/bXR8Ry/+j/2DCjqylyQhNJphf36E6aIQFqEHLsof00cNQ6HJoKc8bh
TvV/KS1K/Cw3lXsD93fSvHk/Wju99MVIRmX5HoUD5BxpI+UGZBag8tcnKeNVFrZoQlu4wRpC+dcP
ArOYSrEP4PHE+V4p3vDrDwZ4glH9/j+z2m+Gd75Rjx4VCx0DlUNddgQ6nprFQHRDq8A7eBIBYM06
uNMrmkELfo8ZH34tzZjvHZl1zS84FlQGdORC/Vq/VAm3pzeyGpjV0YnESAJ6hckyZwpxMEBxLBFw
wBCvkz5nqpfrbSb9kGUctS7QfDGY9+CvcwirDgImz6dOUp19kJB21sXDpxZ7LyJLilO++k9eePOk
4QYEzkGP9ZhJ7y7WMiA3GQmk4ntqjd4itaApfDWQyLUny9w7SfflwdQgoh0gSjrmR1bT9rzvDj3b
h7K9fdp/T5xLyNdvDqbCVhIwC+bm7hHIBadHPXBGgvuBeoIOwfXsNkQjAkHY61652I7etDG3DRye
rzhP7EYCqDW5pdvoxhw2Fth2aTKI1T6T5wDSQXRNf17S2Gb6KGjSI/drMT/qn0V8JQlbDv00/2oA
qNVnZnRoAwpkhwatfJMIePKtGQV7MppFP2bmG9XKhyFTxBNXCoZ/r8rA8UUtXfraey+u0MvqxEcN
8YN3YrzRpsSnO3X8YZ0JC3QeoEPGUmIBv/OM/ckEaJmXOzGXzmcr14M1ZLLynsO+p2ULEqLVUcpu
z5A+pchQuztvYZ8W7Rm2tu7Oowde9I/Dd3Shzen43FPxhM/N9JVmVfatbNBu8oNa7/DTiTUR1E42
MJ66RiJogV3Sl7zNO1UyCp+HX5P4/M9alq1zafTM0xTBFzDbK5q9FwJtl7OQ4+poG+Xv4ci2MvYQ
LzVl1bqJRAWN+LFFq5nzta8K9obYhGeTI9gAhL+yp3sdIIW9uWif/1uTnOSct5WO9KIzVT8EN/iB
uCSrYkNvA/HPqxMbIWty9Ue4LSho5cntRWozr+yGk/Dtq3bU9pas4r5OO8lt9QY3YGChty53gAOz
3qyeBNTset/Rl3JA7JXJeev954MFbgI1lHWLy501PmesZ4JUpgLL4cUHzNist/CN0wxs/FdnFMMh
TjPBSwAPon2do93HdSEHgycelBjfJiW2SV8jI+WunpIZmVN5Si388j2C33Bl2uk5styCYMhA6mQw
YjBBj4qD4dQAjYc3HnEu7jTBABYAcjb9HCkd+vNS8n6nz3GXtDkPP1KNEwhvn+Bp9F6V1VrlN8kM
fXirTcjbIKiygd+ETT9pOQqhvsS+CmB36w6m586HED0ou9JLLnVxZ6TWbAN1F1Ab7HQseAghTsfp
+nuOHdYTpffvAwno/Q9wo7cAHOBPcWOc3dQ/KJIbKs9Ua5DAuWwtxXgLlCD5L9skJDPihWItt4J9
2ROdzu3fNDKpjgD4NE/KlrCjXeHIkBgQRfCP2l5OoXaapAEICy/SSKIN8R0QuEUeDnQmLr12dH2L
uIDCTubFwkY3sbXqabNyuBs+SCydUlZx79Zjhm1zUwByGD55dIfJOzIZOXVQYU83JT45MdElykD2
mrkc7j7aTmbjJ1wqk1F0fyEV9/80R9kJ5aQe0+G/UAnvibJ9ssA6VPKpsvrC/sVTVEEL5u01BC30
LQgEbKVjstj9nQ8e4x2/Eqe7FZHB74GOtFDMBITk8iOj5Xm+b9qsa7ZMqzkEc6E8kZorLePoIxdj
nM70W3pnNe9VKHJ26PF9zliB8a7XoYOdqVY+F0OkyMKpq6PibQPvVDn7cAoEfnZpdTRCSOFWfh4/
o3+rDyiqCyy8Hhju3OdA0VReKA3v3tvQFfotBYKmK91sZaQR7w6n4oamWwnCyR4axA9g2L8ph/ep
kyyvZEJaC0C33VjvjkghbODFaDteOt3Cdo+NPssiOQUf2CqiHYf1PHuEb3u2e3Ynb76iOna47EhX
QRB8nTlCmfziEZOOCasV0ItaQLqKPFLPzp1bLudFA3gCMwmtWVnWojqELumsDgU0aQ5zYp2Fjb2z
y1t98A4VDFldftdN/0i6uMRn89Ri6COjB756lYioIv29RlX2Rv+J97BXmW8FQUt3f5Mjk2MRjD1X
ExmsGAwVOLh1dhTvE2cxJHtTqxeYh/QPx9pYS32XbobU+DCDRsdijZJ3SD/qR5M8p65zB4FhKKKs
gCF+FLJ1MsOgr2Kw8kO4Vg0g7KFi3E6ijayf5DzwW45raaI7EIAguYNwtVHu0ClI0dA5GOshYhH5
kx4ZvNI8dFicgjTL1z8vQW4hPXQEYZ0rgCEWTmrnVlhVW+IvvLxT0RBhPVuyCu7yTaeF2sixxrd7
y4Wz3FrpBuHkKIdGVB2czUh4P0D72jkr5qOpRKJGQklOph0kWRRkmFiz5PDAODnIzziW2i4yDrFH
ZuT70qOPOnnR+gi2smjsYJe4jTEMiPshYpMtiAcxzSznL9ahJXB6oKap6H8F1MtkPZziektHERXE
GX4/MuLiLIORvhsPMh0vsPFGLcLwLvcUtyb0nfA4n2/kRQYMWEShz6bvIB+bk7T6eJF/5fX8djuT
iOC65UJVwCm66yOcq8gic8QEBLbmLs0hCWOjUZrhp7+SYxFYfJIuLDmAuxUb5/i0b6KjLt9QxvmL
Mm3Lp0Y1KSt3RC7fnM7aYboqnPRGclF71E9sKQi2wI786jQ5+F2g3xep5mHJYLRUZIM9fE+sKzQg
Y9p9uB/Vesp361XA5O4+TgdzwNQi2cMgXbM4wMQMWXao9yAZuzvA+APiM5/vyA5tylUy6JG55nGn
q0QVDpw3cXHz74WDJDAzO053C02hspkpi2Cqmol1bHt4JngCSXZcqSs4KiWtJW0RUeKWcyih7Z2o
FfRZ4hTLHt9RKYniBZd0jB6Ou0OpZfvAp342hWs7YSQ6vrRHKnqAPk8ZmdtCLisQHdWFKKvHgSsV
hmMgHHk5PFDfVgH0A9WL8KPy89sW/+OSDhM406sQUx2//uBa84i8P2DKpJTyT38AhCk4Oj3ZHtVK
LmN2a7q/qPWgDyLnYzpnQlTKttyL4aKc1manf/cGEObjUrA8gMHD+gSrmywxb5i+Uy034Li8CdMk
POcDCKxHkpHTUqMVWax94qNLc8LrSN91UhCj7uOlILOxG2RdjAX4q0cIkhNUXlSwiksM6jsYAfYt
dbRWgSJKMZIPNa/Da6pU3lG1V6k2OylTsmoPhGdSuaibbCGpDQHlLzzRkvNzhVnkSkUKzNTyk7Gh
J/QNjjG4nW7mFLbzyLndz+S49x5OEbb2eF+zKxgVhl4kjmrYfxMg0pZLfwsqoXwU94s7CduvLK6a
mSM+yb7yfFNuK9eu1PDaRqddhk2+Y9waTGaqsoMYGb0Ngrr9eLmjti4qltT7uvnLzVk4dpfkyLQ5
7PeIIJ6rJ0Pew/FTKcpEIxfun1VAhbFHdQHkEPFC3CZkAuofu+Y5h/XJ2X31CuT5ygJzs3D9ns4O
D2dGE9qTLLsKHLt7ldZAqW4OXeP35ROP1FNlDP+y2+UMpu9HHqc6W08dXBwhLwT7zvnh8TgNX8GW
h8EQbLLyRRPsSgt6uFANMZfd3nVnMtKwoYx71qLHbK6kQB6uceCqUw4R0gylJFWws79MzlIjhxHT
mkrSBz6YoPSuPH9rg+F0oeo1sxZfcQf1jTEfNBjvidSxR887Hm42y2jIxkXDN9qSc5F8VUgC4BtA
PtQPgoU3rnyf3My/ZGDioD4U3hYr68u4tXil/AZ+NHWkY/UD0BcTgEK+EYU9aJyqH6ekZJ6rnn25
P4+vywJuz/STmTcsXJFUzmdQX6qVhxsiKy6ZK7DCCbYzwu2pYsJ/zmCo1q1blkUFK4pFhB/kccKk
xYCQX0m09K7gcLTNWwHOimPibiZvf9JYtUJFWkF+NxMXqjGGF/wErMyr5OvOZ2xet11yKaFVsyx5
vQ4iuSrP0I3osouxyDyux1Y83XkJRNv1DJ0MyqkUTmJZVFRe3lwJXANYrGUrF/RPuEM0Zgp6T85q
mSeBrQzCY+2t5pM+zURQMMA+gnbBnCej2GBPd26I2Yw8BVUI/AtVVWyVVF7jymjNZObIAwqEqbfB
bfaHEt2QdZDLSubMQXMhbK8WKQZ+4jOdfCfZnFSnVsajJda3yQVl540XXuod4ZWzLCYjd0/fokrU
6uZigoKzIIZYpTEtOrzZqTw+MGUQEO9qFWAnhHVRDktq3lxrzCOAl31nGbFWYtaBqOg0ukjPFjBG
ijg1Xe6CdzdkY6fKEci8SYDWfWvdpdEMOPOrP7zR0xYG+3BHJE4tNo1rx513flEuX/Ic7s21EDdQ
aTYgSATOT/8Y4xGTSzzA3BSMfnd9LCBUCz7mIurKEKyVTDoBTNPc3elcHSiF7ONa0lfEa6tqOZLK
bu1yNsmSI3dZCVjV3kYLQtFWivBML6m+a2Us0b5bbaP4JuFb8ogGXbblX1RjjUgBfswsvEkQlVY7
1TXEC2dCAHW2yWyux7npGgKMF4G9huEzYs1rgFo2CQXSgevwPltCps20GgddmmZfIuxXVx0p8f+i
ax4WB/C6C+pnobE7ciYqldiiWeRvlfcTBGfOHBdcsbf0p/iwT4RtXjksaJ4vCQ+XO8Unyk2UrelW
0ScOgwZ9a11GOfUmCWDiviyCVgLcKWNwPihDnebLKAHK+rLHZIlVp9jqBG4/ghNvNPAj5W6uuf0V
P8W97qxRBEAlG6ut9djOL0IMZ2w3f2HtwEt1Su/dvv/IdNaWmMTAz6Xt9oEEwS/36NeR3Ana/rCa
HUG6uzhSzgWJRDx0BRG7dtFLpb1+QqO5rMfoE9EOzlmR1IrgXmiQYkqbiKKE/z6vWIIU84Zpt4pD
/Pty/xSvoE+Mhl2sBZTNVCwXS0W7emabI104IgAIqZePVrpFGNxhEqtSmhC738v3yEAK98MxIImt
Kif3sZqro8M1xguVA7tp/HCAz0iIta3sl5SCFJx/IMSohCCVz/w7dRcJpR6+fvHM7TnGNBXs+fjf
ckzpN5x9f7jj4yIIREO19E5doBfILVzQ+EXkDKZz76PckqN4sTtit9aPcLoUsVdLBvoWoSxf/byN
hKu+/37WxowSJipaLy4Nb16ibPimMvQ962Ov/F5kLNjE+cxLwPDFc7AWfK0BP8AT4cQO3KaWYlXe
SFBE/Zo4c1YXeyfVTR7zVuQHU+QiRBlkezPerqZNTFl+ptkYP3N/VbH75DMZ/I+jqwE6/qOIvvpW
ZQdUn/C28MlDiruEZYq3xp8zdhQeFUs5Bw688n4Ep1nGOSaBX1DRU9ykG5sAfu8jS9R1iglI6n7D
g2+ImGlm/MwUZRhk5P+pjW+sAK96Ym2wFQh1MG5cgkIf9umP07B+LcUEOBL2c66Mi0eDe6FSD5jm
Jax2NKPDJi6c7ttapjCqnzdRCGzGfRKPobj5efQzbf++cuYYh4qByqz551gF7MfT6nK0jDA4GWFM
1Ul3d9lbtbQEmdTtTlP+hQxvmSMQ5T/3qnMLi1FxKX0jdsLR1zR9kye9E/MLTfGCEFkrKkt7hLOb
Yy+yesnQKtasSnBUsifgT2bSzaXv6sUumWsFLmqQPFmaUGH2VffLsaetPE2rO9cUheAIlbIjE7ud
lUQ34yfn3wE+lrJxzCGVurT1Pxof9VU36bZNk5T+2SI94McGaDmvmg3QZx/UMO+SlAJQT0LGz8cy
Kt2F/cuc/YQfl12JeFiicrTJ8PwZBgxLYRiIIVX7HSmfBVWWq+YwBbNnREX1yc0le6FwHMkFCI6s
97AMCj47G75ENS1dkZN6gzHd0cIFADAPNDfndyJo8rUyhkDAjReZ+dQWF4pgLtlmmrnMkABundAV
94QBk6Lf2aJkV7OyONw0QwLkPMhvWY+YpqwrBtFFvL5zQh9bZVDTiZnNqqKecZh2NSBtPEZDVWPI
BDpVObYWHEx3cjWP0Bz1VDNh15tvpej4xlM/44nlTSn4Va9QFwqZuI9egDBXEyUSak7uj7+E02Rl
ql5xLga/vPXeXRh7bs2CXnCyQy+OVxTAaSWIzANOAvZRFQA+GouvY5dQ9XS+lPEUSXzE7TJScoan
0OiJXhegSRSb6z0hNzcb08bEucrkKo0L7mMmTSH5AnOmshTkeVVQYgwwNrGKZqs96RDSsYHZXThn
leP79PHviKh4gPtPAUcrC76QChBQrBP2SU1icHf7KEc6DXsgUgkCUY+BNy0nb2wpkEt/bucFzDUc
6prM4WvIbo/tiqWjOxyB/GM0hQhyfQmbodXEypIat5g3Fx9MN9Osnu3sClNkdH0Kv1lKbM52edq4
d7K2PZltV0Vbn36zeTTw9pQbKPbUhHF9KOrcAGZoml9JlPdgHBD/70AEE068oXBgC53EsrFL8QYg
7B/Wam8TNuG4StB62Dy6n0dNWYOJlkT+Cz41lpffRaXUGprUaoZFPqH4Q6VPYV5RBf4K2NjsCaDH
JMs9ZDOS5x51kgtqfwhF/YJidG1sWitkuVY07i/pMuqHE8qfRlBeLvv0PvORZPuxtu0om7HWMeUa
tQmVZ4L8m3vytG3Qvi165TuymFakI/0Jyki02Ary/7KbEXoEmFXzxHjdwfvkWOKqEfpEhtvsGh5X
ajIsaE5MK1jRGtOvliH9Ca5p708mAMFhtrguvRf/u6611vx/nvlHxNTa7gI7JtQbPCtHMQHr+HGK
L/FeacNtpBISsRRg3GxUis7Shyv38w+fl2Iscfse1Cxc9F5i/9UgZ1a6ujsGf9wIeUNOGZGUaPgG
ztyI3vljmpdkRFnhlqURgkBbq79WXQOziVEidp6ZY7fPnj6vfTe3ivWebcv29QlOd1V/XOTO3YgN
t59ZZwDfmuzrNas4FbvlLYuYZh64JuGFAMjj0HywskLJam+0MYwJbrPo7IC3no+QsS4TVLhO1i6c
lkaAthriBlHUJ7XEC0/bTEMvrUsrCIao98b54MziJfRwyM8CUtinfzARpolNJeZ/vhhO0qM4t5Zd
01lrbsjWaENvC0s0TVyMs1SKS9jK1rk9+OtHY+jP7bkdzcoSaVrN2RfPEUfS9EUy1UMFnL1Mem1+
w7DDGfgV+3y2QWjJxHr7Shri044jkx6ke5LsjdIe/5ARxiA5l18R4nRKLua5gssfVu4Dmg2aPkSK
DLLdRRB7riW9IQSr6JntT1Ky3bwjHQLfPwTLcxjnnVWAezhUwaPRxZ7L02kDmWbBHh7ONKfkBxAm
DxFnjJapxlH5lXawHWlqUCeJ2QCpOAb5OiiwPXEuqXkgNTar6EFNXr7sHRbA5U3uvqYbkuxyISP2
6znMhCjLdP9bZhloCpUFXFO6YmmOIEucnn0R+gOmAjgYG53hinxZf5bl3/3k9cF8M3bmY9Edr2mJ
2w9/knAvG/MhltGXoGs8V66q9eiRv1RUIspREjMKGwL7d7XYwS/sm+CpDKliFiCqtJhFqJGy1oZe
IHC59kqfZeZZ+7LzVOpmzCQzpPgX6f4nDtTUN0vEiH6ayElq5v9OCCGffMbXprZxLENEtNhj6ckZ
w7G4E/08Rv9XOL5P7xw5VPQ5Pq77386ETodlvEaVIBADIyiKM/znH9X1NoAguxhYAkUtIlIGksEH
038N38RticTbAeTAZzqcqAi8tS0HVPfnzpXl0zN1SE6/w6XUk1NAgt466bdBeokP6VtvA51oRmev
Bhk/Xp9I1Shc4tZJMMO/rZJ5101JGGI//BLxkIqkKQ+FSNNqO4k1BF5XbwB3JMH2sw15EBL3Is1o
l1kR1TYr1nCPKNhbY7r5EYMKvCKw0Bhn+OOLm8pnbtfJYjo40/e1Q7BjQHxVAkbzY54fNwwu0Pg9
679uBi042qfNwtPpcRZsDcPG3z0cyJEb3lipf1lcuAuoIrX+b78TZ821Jz327IYZqmZ2YVtX79AZ
4REwcTWWMfV4I7ncx4frRyVfFHo3B+CbzG8vakP3TayAxSDMp2TGq8OcDJsFkWvkF599GdYFb6ti
EgnaPSRr7PN1UzCm6Si+PtVSr4iRl+6M93GiwEmXZzd1MnUaUvaTDH/D6+cCBzS6qmtY6gpMM7qz
OtgSJcuQy5aBsQXr7m44kOC8/C64tTFOk15eBSIW5kGB4aXh42ZvTzMdhE664quKcgph1mPrtyQl
IYOMjmct2mZhQAyuKi5B6L+5DHvlLohUsp7BkrdZzuJemIPUJNbxjTCNagv5SAaTz7p2CRT2gAK+
yPdndSsXmFbBp6zSEfiHqv8rTspoNSmUfvLKps5IXKMF5Gh/n1Sj3Ho7mibNSLYQsdS52KNYDP/W
IWuADw9j/BGnKn88f9zzNHu6OPvXXeliFaOtnxZNvzoAlUiIsSqTxqFkRc7al3oOMl9dUpPKdnjt
cDxYYZDkqG+2tKoSLm+H0flhNV5YTGMazQKCwZf20lECKqZTG7LwBvaC8yH2lkAnlMyHiydEiRM0
odbT6eEhPcZEAEtJMsfRgmjWBG5AWsZK5L/Fru/w2nCgKdl/uKLQ2DSXrEO/bntfEoljk7kwyxgj
/14c8wiV+1vKnD+HBSFaDnqODt9M+85V6Ys4OuwjZZYEZy/GlzdYRJqCR35UEUw8BTn1Ok0IThsh
+VqEKmb5H/2UUC5lTE2m+B+uKdYV4xBowx4/k4qG5VykN99BneMzRgRVVVgbCLthbrbLoBcG3LGZ
O8lqVIbZdSU9v4UQVA+S7rd7uEh/KAwEm028coREopQfXZdWMxCvtkO/ad6MDJzeDeJ434gTRqEV
FxFozdEwC0bGUVx3MQMF63/813vQa6WH7Iudpmgi6YyQNWrLKEj7AQolQGsjzboTJyUivGo0Ycl+
r8J0TRXYLdurYCuMvbcdMYTEiwj7cpaAcc0yrTt5LnNm7/wTIzt1WAQmTHxxS6LQ1dYXJ4x64mzY
Jzt9uDbO18SJ8UEAgcibngyskNmH7gWjPzdeKudP73AiOVUD0vx4FcmPWnGWFyAm1OpuD4p2Kf/9
i9lyAD05ujmFu4d5JiPyiElG23TAtTIHh0aLpmIBmNQT/Mu/JvPXhsEU+3TjUvovCCwO9ywb7sb8
3XLfgt1qqrpYmO/GO0c3bc8zI4A/87AGVLs5Zi7Q0bHoki3AdQhK0Dqc+5aho3epunNlVjP0yuPj
I3BsHEpSycG2UmXIz3eOsbiM+oAcv0VVj5/5kD7qn5Ff64E3Es7NDA2S+59gmhJb2qratCjNn1KQ
J1Tj1S8TK4rBlq9V9fu0JiBvPjh+fngqJQ8IA19rXMyv+/4aZZGIaJY5atSBkckIO/S2f+1YXDfJ
0tETwTLUPt0cdCZQ3kwHRzEPmWGxC3VCGdRk5POfUMzQFSSvqiIfxNlVy4YUxhoqlB8IbwAEK1oQ
J5QO+qCPJmNAxEmdnYlycSRLTyPas2hYWfvJzzgWFwe/fYlonmNT+kHYZWAIQopjSFR1ucyK/Akj
O/3VYm+ww8+aX5AnSdc17qYIMWjpOgidUiwaV36B9RoP3v3iNjnUz7Ne6mb7GS9buIFTI8RKA1c3
BxPG6hBiCQ8fdV97aNaVmKQ6zmvUjDsYt1ltkV0NKhrVIUA24Aq5slGyDIBhXFzblVmG0HHyfrjq
oHAdLNir+ki8WMnzzkAUCI8lYtutiBVmomd1Wm0DR2RhntpeCvN0wfHaK6hNAo4UNwbWOcFdjk6K
PSaM1Qf3aA0SOz8roeT3zyoekSQjGswTjieGgMJp47KFCRHGA4L4iiZREx2ucwnxUcXo1FFGwYVy
mP1pXzCXo+Csvp580dBHkEDsJ2gfUV0A6ymOQOaRuQTQbLdMnLO3H47Pvi50DIUL3gItFW+fp2xD
35yRaTf5+S/aiB+bnYFX5YRZ2qe5vWEhJ5HCfgn6n8iuTURyTReQU8yvxQ/DGmbcDST8/2jZaK4u
jh3mW4Q0XyPZ1EYTqhwL6o1S6fR32TmGL48s8bJYlsj+Xu3fNctmliqzPr9lqmZlE6gd62I3sEkU
Tw9Otw1GEoGwfJK/y1/sQtnDIaW3d1z13uTxoXXEHDF2CvXXocgxfNqVsGHcfR5GQYVXoIvu6Wsw
UCM+MHCJzRJ+ahj8SaxwW1kndSBXD73RWymeF49jMcuvp1huMr7iLKBjWSstckUn0BzOpEc1YRNR
VqLQFyS6YPR79wXSNnYrO2iCifQGadcs2WHOz87+0FvWpr2T5gqZ4cWZ5FY32pzckbNeoaReAiKP
bpo6A85aBp4u5fcGpDuPQV8l5VLQhp0O/CgbaduMzfy4wZlAHrJtNVU0XdC+SEvbf1wdLXrgFQvO
N0OfzBR1XtP/rHC6dgZHl5rALQGP56PJOfilOiLgNFhAv18dahgSjHK6LMRM8dqu5gXN3xtyvaCq
pjXHe9xk2r0C/LTf4E/MgJ8+ZxoyXsWmkorLlg0p9eBhi960mRhcY9Hcub4kJIVROZ7cHuhHVzYI
zqaZeT4K6MjBAecknG6xEyV0s8t1ffSDsP0QKUgEj1BMYcXSIU1u6thU9SxYhys3gvCIraepK1Qr
FDIzPjR82fJ3plPT9vocT72n+zCWxK8qn1uT2XCz6waPTLh57SL9iv8kQBA6A9ZlteCJRv4Tby6I
UfK30/JvgJFXC8Zubuklw5c3ZVFGF0sV1Drs6kg7zLweVqAHLipjUUiDM5W6Bjh5+FCoBGfIyxpY
WmuvTkFMmxZ66c6Li2i7zpAiHaa5JMv6d+sy+ujXxSNOCoD9EW97EShcQ6JGYnIFU/M1DoNyBbny
UVmN+b6ByKLk8J8C9KSNg9R4IKsV1U0wXTXtaGAn2JxVrWG/IR9s/grlRAojdMQ+SPCH3b6yyjTi
EZ4/bdngnh2NQwDDlY2G7pPn1FpI3RMlfbOKobjn+fsSZah7GgcF/FZedcYVN11iVzIhc2LG4EE8
tW1vIZt7+HB43l+XQsVAlWg0hfaL2MKrAGuW/JKrRHmlSJUofCe1lWlp9YxG9rNFFOCeCSO04o2c
BlU8nk26odB7BSkNDpZxB4parSEHBW+nYB6+vggdRyfmtD5amwZSbWCd11ktLRWmsdTBFVSumK3I
0fN0EcETkAwV59kf2AjuNTWoijpNMXFc+eVoClVDrcGbfskDrXLM3bOnM9WxCccKyyW3R2GOVrhO
T7XKI5n4MI9GQmOFOtrLpVQLjCPrM04XgxQyMeXu+RcvTJS/ezLYobBSTOW3HWy7St64G6XIaKvR
SMWL0UXhdKDLxooFHpBziaTn27mNFLihH8p7xjgKMQ1rYrC+1Y3t0NBBO8aKbKUyZE56c9XfSEqq
0pJQuFZT0qhiX9cx8LIf1MWHaE+ah0/Fmtaqo7EwqleuikmZqj162X/KYzEW4omIWlWCfGtklN5a
G0raCQpJZr9mTs/GwZ7ZJD7T/3W5mrkSIwFC3riKJ7CsjLnnXe5Fm/YaFN0WjR5Li+e6wA9vN0QA
BCbpBkpkvbfW3vGIpHxHHPJs4ohUCja1TzsEkRTTCAcMNabbMLcXr8jmobeC8J5nyptz+kPJU5Bl
/xnAdLkovM2X2yYLoWXTfH9p3/ln6Gsmo6dNpT9dCyPx2pTwwQsoPaTDK73y0ZKrEziANo9y1077
mWF9/h0ulfxGi3mgFG/KgtM628cvVeJFXFK7eujXbYDJhr2mksHbjTVupP0ny5j2u12nA7iko2u/
0qnfClFgp4fRRl6ROugcg6bUdjDwE7UZidMWMR2v/STj5mRKtTlGedn6BuSrzEXgnavg8IWclRUR
suoJsPPEZvgyRc0Inu9SH1RGHPQtNDGbV3XlpmMM8mC0ocZ5g9VgLnaUDf7S6WAjtHOKjVAfHoEn
DjcGeMv3P8IPRLWdrlcHquYDnSb6ripBjigJXh4umdALIVRGXvEFTRV98xPamSWp103Y0tFYKhkf
gZV21r+/4b8yuVbHXvuCaWPhITCeG9Jke1S/AcGNNa8HV5nc3RplGx/tT3dehqj0e0DK3lhuPTnk
XsQz4uqCjr5FctzbaFN0M57bYWDFOGlOXd9PgZKOr6WMv6e2v6vejNZgsCoNV3GOugPUejidwlLE
FMQbNWA1Zfi95gARe/KyecRq4pDenI0dOGX8nf3mRqY4w8a+9PBh8KLsaiPDA8ObNHth75mtuS6j
DVin5xM+dOBzjxTkjPfKTxP+rQ11GMg5QBUVvsRbbXjaJhFhaEudmU1dQvOlfSz68Q7uLVFvp+1e
mxrHb2yzbtiGNTUTr2e436Wl1nD6JiReP4z+i7vaMCnsgUQsQZy6EPppvDdBncQ8Jo0LuiZWpCmk
OXW514AQJCRi66mnC6K0iaQAgww+K06FpUKiFCjWunajAZHvC05dhRX1DoU5Nvmuburp8go/8VVB
SF7O+2NX6La2T0lQ/u3a8ZGpYfiJs0cXT4Hd+k5K3WKqwG40G33HUDCnsD0TlvJF2LJqo9FcAmlw
I6l1gOOwsj707nkrzGwk5KdW/IXcAxlMVbDe+3/rbO1Xasj/R/X6dMw7w5X/AGStoz6kUvD0uqm1
KEElBfYEnglSSTCzbVpAF0DIBcgqy6NZlsnR+gEn6K3sMwjMYC88yRfrbFsBGW/r3rbKMbEEYjQ1
fkY7sB9Ls8Fise6GcgIgpP4AFUGBl1LrDg4jK73UsICYnIn68dnb+W/lsYUIXmmSmcn+B8W+m0h1
ifxw4RUzEuM6nnzkYmFnfeuCLDFi3+KE9D4ppEPvC1umsKBqiCfEd1zcHmQZ9YvSjRwTVx+QZVoZ
+/NdytqKyynd+4VPfSUc4Mxb8r2bR9JDbn2Nf1s/7tUPSkkyEfBPNELfFf0p3SnVPDZsx5ZlD9CM
z99b+kgrn1yfMpGsb/FS6VFfKqqPyt7WFM78sRDNtY4WoX3mLJ+fKRm3rweg9qofZwzFeM++L4SV
dK6edJcukbNB4aoPU2alGzmbM+bzoIWs81oB6hf06g9Nz+9kCav91k/3BpgwTUQfwgQRlMwaNW5l
6Tw84bjXLbQktDVFV7XMHR6H3xYLu5WYt42MtZsfy8ZoFtNlMO8n57t9RilMF5Hj3a4Xk2gcb32v
GvxPRf47bt1Cxt7U06O8t2kyqDzOmMvvFfDsrH+Npexjf5HOY+GQrtrC2KS9vdN4xPRrzfr+3bOP
zx1mlO1FD0buUCH3JQwbTSycD+3Rtci35eMTEq+0iBUkGztzNskwDf2cb5mBPrLnQpUcSPFEnmzB
Juv7hMY1fWudFyohTYfhRuJZlBM0CNHMipjK0UXCHnXPOJwcnWDeBKlvr85KJDFXwSgovuE/sFMA
/fekh7jGMu1h5uH8sq9BpGmUCJlutayOCZqHB+2Hf4BJ+jSiOPB05A1xApfMUSJ5Tw7hIddyMZoY
s9LDM/qQ6bgoOYq7gKi7dEl2ezOgCw1L7srJ2E7wIFQjQRz9k2rOasKPGvHkcKZwCPQ9R1bGxQ9y
AntPVtiOn2l5x3ZPgSuXWmkDulfz4dwBRP/1ygEWSHPejvLfCFQpifJenpcmUj1fNBQvffCgu+hH
aYrnuiGINMVzci3rjqixYc94dTUb0SavvX6XLXtAGKjoseAK6BDMYIZn5bUR/SVEIWP/e3jT9uqL
vZmRwP4dPzxY8Onupos0FgE0MOJTjs4SH4DaVB2Pb/qtT08CLRTTpqZZ6RkPPQ0D5/746HhN14ZT
9QtrQYYWgLUEI+9xiI6mDw0cIJM78LalHBT8q5TRhLeQ9SKqx27dVe1LSblCZzOtAgeyS47jLDyF
rtBS3xOkVLVUd2paRQr9Xsihc+KcDQme5dTFj9CYwDF2jYtAbgo4t49nSwL2evbORG8KqPD91axr
i6MCCL4JRL/UvmdORbPdoV00qqGLcljL3OtbuAKzSo3D8Cn6LWz6KtwRAQQ8WUiglRyp1wLKAWVk
iDei/bqOS05HoLtBvh3FOUDGonPNZ1Gw1JbE5bwBO/gKvI50GUhb27ro1i4QvUO8jyorCT7cl8g2
2lo0s5q9i4RmNfd6906EUDaNEar0F7nzWyyuj4jjPDjCWKj6zkuY+YbHQGMQdtre/A4GGGpYFLKy
r3vMhiDtYQJq5lRFMgygID6Hm59Ax+8zAa/Y49CWi/YBk/6kQQ62rdpwHk08l6KXGmYJSvBop3lL
RndKo547/pNW+ow83hs1sB1XKefSbK7pSJR8qYWWyKbOik8J4oMgIsBPzAmnMlgLRkW3LOjHZczn
5LR+UZqBU33RcXHnxXqeuQafRa/CQlWRk5b6sljXlamsO3Dxz64cLuDG/pzI3WGquNt9Obin/hNe
FfKE2AIjkpTZHj5TLEstzNCegib7i+U9xXFJrNKV3tZBTRkT+vjSYw+bJhbVc3BI30HIGIUG3azX
bvgXQgBEAXdEs/KKdGnIwDyLFIlUV/bgTpmSoogFcGMFDaB1UrI35clZ8OMON2z+mglPOAfcg3rA
JKYVuFMBbkOCzJM5bNKpZeIuQfRg/juhoAv2reTp3UwPYJ5gsifqPEhyQ6UGCj/IvcSJkHCrSEAc
eJxzKbwegQHLvcoaQh4nLqwM7h4vm5dd1Q5Y5oQkWYUPxRwQ21qI9pDSTyw0uZhYtIkJuyQ1Meo+
H0YcnWVsRMQzkZV4dmrb5xz4loVgkEs2JXRFqlJU40qtVtx28SPHYL4LLHHOteTPvRR9ygydtYn3
4FFqpbd6DJ4YMAS+HyCxYtC4LNrQDbY3QblpskNvsUQ8YvXqd7dq8flBVCEPdTcueOoTOmibvHnk
N3VxWFIExcFJqKeeRoFUv2MWU1qAaRZnqmRfLDxcXQBJGTWJhLbXu6wAq7hQXnVQC5l8naFH8qB3
KSldhHyhznFwo0eqalOaf4pAF0EhzojWKeRy+qW/eo63HSOGYFrpx2pn4yGOZLhK9zlWlgZ6Sd+8
J1cCdPUgyukTqHWXJOu7rMSE6lcYI7wwQWA1ub/1+lK2pJyyyIrOyYJddmJvvf0QrtxvwBQnQ8i/
x/jM3CRVRWT4KeWdP+eiuL0qNy8OJAg1QRvlp4KOrhmgDAiinzGnWEaJQuqhriyxEa01BgtG3R15
bQ7U/tO68WB4FXycZYmkGfOGA8NQn1VurQpT7Gw7SIac6dmVpIlAMJYuKLqMkLCeg+KBjryK5wJA
JLhWN4x3rmID4+l34UwtQN34Ezb+uDr1rRf+PL47WHEQtQZDKyAY8/NINguW2Q1yb3p5mO9J0B+U
fqxlNAQrZGy5+JRrgJXStq5/X53GvYl/gn3F0iT1AU2ebhoIKWFVfnr0OTyPFwhAB+7aFsPMXnZ7
PE8qnGMAOVksDvb1iLicERkncQHEvYnWDUa1XLV5E7Yq7I9lcWXAy9b0i0R22CGL+LRDMzZsbgRx
EkPpfsSGTPa8FoSDbIDgQX+vA9BV5eEDGNr+xTCbgYdQtPTUitBwlSeyQlmiemE1jp/+K2HXZsFO
C8MlTy/rVtIQFf2h0fBIDTQi+b2uP3blW9v6OVNdyWBGJ+L3W0FLLWQHGm3ppvL5N5NAzCsKZ9PG
wHiiUBomsCX979vpeu33rfmuVbkj5G13tr10cyvf0ghMQqDV5e9W1o8f//4xXhsYC4GrChgOP01l
dD1wisP5R4NDHgoLs6S6mA49iEgksItyPW8d1F5Ok5Lep1QxPFquDSJhSeRZfEAB9k24LQJeigwt
0K4mPQnNZeZ2zzh2EHrb8hF6XdAwGP4ciZn+LxSe0ApLbKrVC0FaGPFHlRaXWODKna89D4LiiG4B
ffITXIiS3FO8rd4267ezk/YbrW9ELquXPnDncEoO2EzqLDmWVtXM6Gnpbks28p/aiJ/pAUTm/uAz
hLZ/U6+sa9eVGwrb5gJFmK8S4lA56gtAfknxfH09rUmMjtO9qYPuWWpdK7bR5+9h5RUxT6WGZa+B
2ysdaJBzurKBSGfGzBHxBjf19MywpuSOGDECJV8Zoc+HzWxwzqQqP6Tne37PPnxqEebSvGsGOSQx
joKTPlNW1CLx16adDLF/q9hy0z69YtPqmieRCn1UDJVdMbitwzMhSzJBMEevq77fCwSu5ZFvOzln
XndOM8payDZPvqCNYfhlQ3AYmvVp9fjC+b6N571N/TEZ7CZ1sB31k3zzhqLRts0Neqw7gaZSwb6/
vYZkXpTVY78sULyEnpe5X9MW0M983n3cPTX6dHibwNHMUDkD1gav/fFtyVF0kmxMHviK7Tw87jcK
OinsY4Qqp+LObDBFNZmYLdp3jLUDEAFBtT7CW1cebnl0103frrm0vXWZQDfvojPPL8KALisgNVLz
PVMoaizrcvjfASf6lp5Mmk9voebNDI7LVe/kGbfBBUcngBKsA5bApMYAaq4ZuHibbRaJLEn4q6Ko
WasmAcau67HfMPs8cW6JySZ+9EVLvq4ZWMsyF0ADbPi/YOe+xFabYTKE49kyo97mju/NKpAWGTCo
XHe0yZh+JhKj0kHGeb6O5kOYB4Q65Ae2B5uhaQtxsOVr6va5vE4EXNkAyOvth8d3oh8PeB/A03XB
/nF03dDGZ32/oZpORVLi2iX840wnU0XL8KgslTXLxD6rIfJ0gfvqLsU2cbOe7Ci3oDmU53hylpgH
aqxMYHJFB0bCmwBKI1x6GwqfTiaMDKbBGpchx+dLRSWzQYdQBmdi3FU00IXeJc4RI+SDjtSfjdTV
K/6wyJSqrTcKLCas8aZJtBk7eli7H+kkAznSO4g7N/M0G5sNE8Ljy4EWVOLMp4dbE696QohjyYnu
LRbqZWW/4BfnNS0EwTjQN4BjjJzVEnCs1ldnpltMMP2YgCbUDbj0yWNwjdv5LvHXC7HsoYe8YnFN
PzMgBH5IQckDLCfhEC/Of5DHsuqzplsixxbnjzHRWAIPjyWTrCIxJfChu6k3MAEvtxyO80oIozPU
0ftY/YqWnRci93/QzklK5kFMn+tbmw8Tvt8/6GnVIdgMQ4+qQOKVEk1wvwOzXt7OklQS78xKWbZN
bFtjrcBtX4j9Y+KtdNc0/wL/zXuW2f+mVCuji7fzIGnfLNHo47ELKqXzGd7+wHy8ueNLI+nfswVX
+nHhaXp6HUbJLzASbPB7W0SwhFDK6q99zpconiX4WL3dN1aYQL9M0dXgdDazQhpOZjumyHZp8v2l
dTAmlfTJSynxie+IbYkHnrEm4THcn2sLOVX98qdZr8L8xMvfOagQIkbReHn8cUwx3t6z3VJMuB16
mugBSGOlJWG216+zv0pct01D018FXEh2HJOjONMELLH4qfxkIdGwLSc+py/f3c9KsCE8M+Wlfo3h
81Da7qwnxNOlsFW6hC0fPkcU99yYp8K/I+3lsWhwBT8ZW6QwZYilIdRsNvWRaiyruPVeq7pieJy/
2fvODb099QIDKDUEAbSafhsZF2gcW453xuNYgos6nulf8OFaJZpMv4gtn8GaEGr6VUIkwbYQJlgc
bKLLhXuqshvReJ9JLELQbxFlmANqXRjP77Me3mqMvxpjY8yC+5GvJnfyuU2lXAQ3fwlcMHvy/Kvy
L836mtllcBtmyZcJx/Os9M6SseqaqqmjidRw+702uGsl6hNgR/dSKzlZfBcYYR9LkOSzjKhM3BPL
Eb2Tvt8E8zd+11pir1ORsPTRYj1LyhXWgs01DxPvzrnuaPSoiX/A0r9kWkqlRRV2nmPkas5N/xXs
gksA/i2zGmN2e/D8Jz+Zo1sdvsL7ecarUS35XKQCVSJ7evf6yWXBVDm/tqyrQ+k2rJvjUpDAqT4O
bz+ai+WIIU2W/ihkelmBck5mxGvL0OuU0PP99uj4nqtII3n2PHdDQJC5w+60UpGgCA2xXNad3MTU
Lo+ogIMdlyd2t62ykl84R5UzA7DveaYiTaSga5CM13B02D7Wx+2UdXVezj2s2RlfYLGMxBwpa9EJ
cOFgvpNAsoA1X8F2Ot7YeCMBlkyMUmbVEWnHpzhlJbhcda5oNBDjJZ/33hEa07GRnrmDgZeCZ0Jt
XsrwSVBAa+dIfYplt/eZStoo059LgfNxz/uB8ONJ6XccNAJ8DVM/SoiGZyNZjpapZ1Lm+dYGiCev
BsPoAfkh5K92BK49rdPBWI4UQys7bHV/EgMQmXJk70pJUsShGTGaRyevk7ogpwZcLuqUTC+S0PdT
WKuybMKvfaI1BNgIpEgfapLX1IubgiZRf2AM3/3IERc/MBddyYl/QSp6LN1af52Ya6aN1sguS6Xh
ExYxqewoRTO7wFMUh/Q0p+XDr3sk7c0fHIQGg+uxvg468popSMNUPWELUjjnS8NF1oA1+0RrjQ2c
afqDRnHSC5SToUcB1qEEJ/OYlAYq8xGyTWwsR0icd+4wg/QqcsNuhhIh26P2wty+jD9jHnzMkKT7
GvCU989Ch4mx+mCOyiz5Ph8qPdJRJTGoQBsBEIXUJCwOvvT0BmtU+Sk/ad52VFK+XqKPYc75Psrz
MyiHxxR5fCLkqna0UrMmVNLxN3AFh9YRcPowRH5ldfX8kojuqopg4Qok8J+7+5jRecrxS7BJguFK
2mwpy2biX5Cy/NzfG5eve1pAL2Qbs3QjW3LpFUoq20rct+IPXVbVeYr5Z1TI7qH5/2q1U4gZwgZx
E8ejvB/MKFX0lYJEKYSsgQG0Gd3M/Uhsx2dwVRxMHZsyZRPsLEOTQk9Jl+3ByVNxAZk2W1g7yYca
uf7yZV4zKUf1TEPYb+pOuHRJpf6oEupvDT0TPDcjaLyBT3sVIsADp0Xwb2HoUcxENejp3aAr0+dh
Nf4tKezklriRgPwGotu0ue3mPQZLEkpxmY6BRu9bqOcrcRys8yDDEdFvIAK+YvLiYaKwWmPPpAPl
YzOOKwIkFfpIovF2d0DhwwrivjSR83NPFNzVr/yvFRJ7if4u2AFbwXRcoKmA9JSCUGEFWd8fbuNI
TUHaIEcSnNgm6m5l19lw6gFrvyC0dTfM3YvebrjrNaH4eGpmKd4PkzpJyodDKPeN3k8bp1sth5qX
UFywMmc4qB6itVn4x8KqCOddPCiRBjxUC94Pit8jlVYC9MfTlsYf9XTo6bpLBiuX3nCgqTuZ1Li9
37F/3q2lqDarVtHmqiLwrxVVmWbOVobVwVwk7tOnmFU9DhLW0Hw2DOLk8RwtomcyahnWfcyzZ4uD
Bvtv55W72Zs3A5S8Y/WWHykqiAhnAOLYu+JRMT2sm8KrU2zxHhCYI/XaXyH4EBdVbuMdoPg9V3B4
jpdTv271AsDL7a1FyrjSxHxm7qPNssvwyF0whEgjRUDqFUGAYvXrbXzp3iNniV6DrRMrXa2wKh+3
zbcoDcYZ4f5nOtOuZswTc82MPatueJV69IaeOdxEHcIKRyJgbgRaypQ4S1KW6spu14Wa+BBjJzYm
gRDCgfTKB9/qdC8EvdhdUN4GUUInv/1+DDvP9ccyHXpXf6WO2BAuX+PHfzvrrsRVqD9e/4Z3NK3Z
R2wQVml+J1wldz5qvzKPElmPva9TZaogU1xHYRJwhzvVfTssBfC7TYoJ2lwrMwxP1ASGisb7yNQL
N/OQuCGI6fssp4sUNWvweA7OHWS1Wvb/cgRufALTMHVHhhyZrgpVix6iKyOvBdOt4ve8wFXWKWjo
zgou281ti2JBmjbH7LXm5Ib/tEPtx71ao+Ggjok2A60eRFwGmOcXSZMSlmbPg8sgBSuV/EoPUxUC
k2P9wiCqS+qdamsXZ8b9PMVtHCQCV+L4I071JHF5msJ4qXkYNcs7ygkn4KNDdYJedVMwghk0Et3h
QwYFFC7OaqaBH754v79H6v72tEQDK+ycylH0HaBeniaYQ0u8dJwKvekhS6ENsCQYYN9SZUmhMQMA
gQS7mG28ton5Dwqlzln6TunuYaLocRiJQ2ITj8HaS1BvHbqOefKjRMD70BhgVL/1woQavMteSo65
KXBTAUshHbSL0eb9Ceo0vQCGM1zWkclQwHbQFtuqCF9PmnqM2/lczblW+PsL03Tz2JatbjjHWwfd
gcHOQ1CzfLFvyQOHQ7QYkNc7u5snuKGEB11oFGneVUJUh0AKsu0r6BP+EqcM0ODZH5eTmzDOFMz0
fq3+7enyQPJyR8L1xcEQ2geaiju6Sbb59g/ksl4oW6B9lZEtg6Wyhf8Ai3lymwr6oFxSv3RRZYLM
jk785n5PkAEtClwoVGlN7k34O+xQ6464mcn6ZQF/Bar6Uda3kDuFvi/u0b99FERBBJ9hdH4JC8/L
SYfwTZVClwT2ALfoeoVd9Oe6Muuqug7CKRrbtfdAakGJnnNtoqMuT3U6TYrD41Yek61mFFrdfxKl
0ztOX9GCnmzW88VlJ4VRzbqAON3BN91fIjjPa4nZ8iRPAleq75ZB8EKJ1BmZHiv3CqAprQNU7+Yp
hQzKnL7thfgM33NEUV3xUYluc9vBMAuoW6z3dP2T4cmggwjdekP1Vmx7n1uneZCXQhFSrfdM1rC7
kjMqrEicAMWlR/92Zn0ueAHyeFphQv39WvUnfl0MGt+P8TWc0xDEOkgSV0kE/zf2Ah2VT8/z5gZS
tkWuOwNxS3tzngAQp3QluSD/s3oTLumYqdF2g4glpltM0mUY6h2+2GDj/xpxZ8T15LNC5994u7rY
R3WIRXwvk5G7vJfJK04sL3Ta8nBzj9uH5tkrp42k/ghdTGAU46/oxIwfgq8yd7D2n/h/Orzv9bgb
XMpz0nDDe8c4IjnRGu73fGA+DH6n0DuWa9//pdgHvW9SAn/+5ZbCcA3JgKHxlNCaCwvYpjX8KJdt
hSx5ysYnZojLxCmwgzFf3VEA9DdQrIIK+UkrzmmKYELLRly4BJjQqqZQM1g6rpRaYeKwUbhDjjuP
mCJMxfs97R6GulIZXzmBWXBCMslwM761KX+i7ugaXcqjgSmfw0C+aBlZ/GkGS3ZiFs1BfJWBdJ5W
ISP+Wpe2gwTLrtPEa0TITxmqn0Q5tqh8J9gUtkliiu9EDtaPTpfssQ1IeIyAnnpeNyvS4fxxKhY7
JJEmdUsaDEs0ifbT2iON9lTXHj85Qwt9RC9KOc/RfyQm12QLniw4uY4GWM+EB34+gWWvkceCsO/u
qi7P8et84Tv6CslYdCPST8iZCD1kpuRiNd3KTMaKROlCfilAWEGrDawptNSXxam5mzD9vdAmvN6A
Xv7dPxvxYSYxl2+aLeaAjCtt1AqTWY6wBzN2cpiSjWptIxQVZk7uGyda8QMYJ4332e7ulFTWJHPB
Q5qyBvt7TEEN4yK84rHzL2RRY1ZmXAv+2HrTy9fVwDOyI54sajxGk2qDRCpdB6SuSJ7fRLKvmUUm
PfaAO6V+erMJniNZa4q/E0b3whS4to5hLG2Oa+QUiaS1x405VvINpFlaZ+B7o7xveScdxWTu+O9O
3hXhWQ3W54D8Bm4Qj8DNEmWzh7m9/GIAf6piKXw0g6zZ9aI/BK4zeWN9EvrpSn3fVUlIAwYZKZUj
RKy5KWFIJSQnOU1wXGwQpomoO5PJMQ28PfjQLN4/1Uf+v80bHjs/JitrriMgpRV4vQH+uPh99N2g
N18QYF7GHv5HAi23gBcjC89r5hhNsyDq86dba9m6lzCDJ9SP2S5J21Ywxf//kFpI3B0FJGCj+s0s
6AzG0S0R2brtm3jTSeLKlxMVaeSkZXxxBTLQUvyVJnJy2BrYWFpg5F8fLZFG5RY5/VTXihYXEp5Y
o5DeHXUyUeM1vakGEv/xj6lFAfJJaydN2vmBAgePK69LjyHgrBLu+EIaNlHW13n3CDyeHZEnzRjK
rMNoYrW1uNrzijiHh4bthhS78Jg7xjyUE9UiX4ujwecGKin+rZcpAxgK3XGpWG3EDo7SlVwkXmR1
Ijoa68Qoj8VWbJLD4Buj65FtSJ5yKC03KXIKpGXG7Xf3lPPuApk+Ryd7V8JksNhnjnlLuuKhva3U
aua1fhpEJ0hkcbyqaOX3zUzckWO9wRATViRarNIA6jOPy0TUP/EPSXuOTeeD8OEe26SJwyp7Ukko
w8VE4+oKZxin4heIiSSJ+KsUMD0bF39IMGJ7PUny0wsWtfXEEKV8CDf7/F4ZURbfFsvGdZa5hd1Z
CpN3tQhjt0HXlljj1a1FiZg0PorVKIL4apqEBlmWMFi5pbVuKrOkF8V4UZPEMl05+2FbU6TLEovC
XgY2Q1dAxiJvhGz+rnJM/4QP140gQDNgXr1a18mNJ9tNVU6GlVwcOI1LSWzB5pQF7Ocp4PJBgV1L
g7mkuW8d/U/LN3cfi3TngXsEInwlR0AoK14F4bOleA9+S00R34u1+rmyWWE1aJfjXedNVYtE0Me8
0dRutooN0oO6QSUbctbWTi/nghPTAjP4B0nm0gwO6Sgw4wcAQOXzRMZRp9xH2MX0VB5b1N3Zn31D
15KSbGKrzkr2Vxui/tqsczjn/EaudWudwgieT4xqeNWyzshRU/jr0nxNO0/1njnhqxN37miCRhbV
T+JaGlqLIcH78IxpbxdoANaytUyu4yVstLeGCZSOHoHCQ45TqRfXnZwyO01WKrcjbkfGC2cS0PAC
MUTWMa371KMc+qn/uEBQX+ALFjqEZ62BswlxpjkYLyoHBtjv3aNNF+7DTM9Y2JqGRb8/8UIojmCt
yxGBBFNMCuJzTTYMHq54DzPETe2/RDvrTvs7XeATE1AlzmVbuAjOGN0/zqg8qgLDgDXszwQzt4P7
bTTVJs+Nw6vgOZak9wQYICheGM4PdOPVYfTqQHQI33LhC4o3YRhzkmMemft1vLLaqWZOyGfCdHce
rOOuNDVvOy55AIK/kGV9gMvvqCS1LsBzJBcAy60Fzb5HSieWcNIQy+cskEvF1R2yQjSHppWeiZct
pOKamFtBjF5RDeKqY5xCrgZL9sEaboaVNEoxpebj6OA7Ooi2XbCJmSoLHl3ceZ6RD/yasSMkwYVi
6vNz/x8qCrLa+zYOQIL+qjXctgbviohLkLeW0v54ACsaeTYqdpYf2KEnUhbuB43y/S9zglvY41qZ
gGRXkZb7jjjUV68KP94knOLQr1TgIi4PnYJLcmRN4MLv0Z6ka69kdps8zB+NqXHqXnjyJUE5KXw4
ZyE+oh4mJGUpdekt2VyriWcmo0KmvGunZKXB9bICtjDy20r63zOhOmE1ZD1c/qGk1VeM+Q/z0gR4
8GJfuWblFxpn5tHquUiC7u4iBINFMbUodGK0Dl6fheBUdMG6RurQYwGtsxLyoAL011gtXpVsaQMK
tc0iBe3A48LANHGsU/Kl6ILqXVqnOLnuF9o+BOTNLwH8gncaiFX04spK80i5J75gPRS6thnJ/lYg
Dmcq3q4YkBOSSPZFRswlLwwxBMwsQPKn1bTPorUYBm9c4LSTZCw1ZjiVPZty8M8J6MoYgje6LBrJ
cmsg1yMI6/CimgGsv4RvRNC9oIHA0D9pK98GbIvd0h5o2D4aMiZEMMSzjXA8RMy7LtY9mzcYDnbJ
GkekpXEEiCJFSzuIMThSqC9s2ML0HZadO5I69kFq3+H/ALI/lGtnDAZhUWXUMcLOQ49G70pxOyYZ
vyTMpLjBpfqfGqZoYSPTyNGE6yK9cu3nXe9VQmZkF2QFNenVsoVnDN5lp9Z9wmjKRpWDDsdF/cCZ
1P1tMkYDGuu2QX+SPtOuJ7f/WEM4j27+r/RyXzYxVMSKs5n2nUv7ZLrR6WP4dwJDRF795yDYONzy
llW2raIK3l4cft6sxhkePbYpbivaIgSq48dk6zmVfHDmqSW8C52TMwkDI75HmQ+Sy43Nbk6r8gOm
p891uE3XFQLkeqzMlOSmMeQHGjBwODDKAYXvJeGieTMn58T/bHnmuMRLqAhGYSnPYt6TfKwWe5XG
lULfYplYs9rIHgQLxe/ydzqTZ2jGuTxexUzLuVfuQLth3HndHwKi/MeLgAyL60qjp+H9zKpIlUWB
/S7YbS6Ry5y426aoPEJ0FM5NkJpIZRghIaLtCKNyZoqMEVUY4aAhJCLow73WID9E9B/VB/T1fqaC
fP1Nt7mjPSXEH6CkdMcFIqBxavihqbygg75XFPCUptUfVzG5lfj0qI+YyNB7djMNr6p3f4XsgIHO
lT1kefJa1g4reWCv/Zuvq/tfipkye62i09G2uY6LCKyHlBEtvfMNH4MrY5+Jc6grtG7Dnjd5YX7i
tY1tUfVOear5yBGm8DhOFpiuWXJPzfrACEke7jQ1h2jxmvofSjs6WQZ5TVc6JIdHrwib3NJ62GpE
HNXTvvPRdeRwe3t41q28C9huuMgUcT6OrrRAHBziu4wFeur3K2QE8yqBWLcJBkFzEm82/gn9LnlE
YzftNnPv28oS+SEZa6ehBevmTybBpxl2+y3y1oYhuIz8nOdPKR/NoToXrS3qzJzOPVI54m5JZ0oY
0m+U6H4agi48StmF3PUy8dwnuLVvXSgzarAkXrShFr83VLemlbQd1vgU00iq78cRbLRsFquUWjQZ
hXLu1ZbN02Ty6WvjRBaieBb55s6Ic1oQw/Bt+0j3tbp3M95gUStV10IIhJ9EDcKAKuf7JfCLvroK
HKa1Lyluug58UrWv6FXXcJNTGuSWPvXz97egaGHsXXt17CANb6bAz0wwnw10YKD8QUD8CwdrfJQr
wdafhTLMzZk7kEL+kOp2vMT29wzukBgJzyj3nXeY9M7SrqSmUSIsx1CuokXPXnPNWKmE8G/or6vL
LQV6uM58WRIvdM9xmnx9iW5DvmyQ6cXJjz+1qa3aan3vMXrv6yVMZ8MzmD11i9RvZRXAqltb6pft
PfN/wgmqmt5avbjhxS8FDsjO47jc8uTLOVAkoytDvfUtHy0YlZ+9Q52+Za/ZGpYR5djWl54YinNA
kK+QwpXVBirYwvWRJG27qjtHCAZjNnAvEeKpKIpDIB8W/2BAJR4LegDeP2kk/Ek2V1eW89KMPK/6
DVXhdGGy7UD0H3M6I6zvDa3/szZJS5dbbzbnze3Cs/d2fLiSGPVXhVqs3RdhXS/2HbesM/O8mIjw
yRyoIcaeyTQjTaM2RI5cm2mQtVgrG3IHe/3z3SVJZTYjdudWRpfVbWnNHUgTRrNHFm4owvCJ4eB+
wKJTegPCXAYGfvwEuoDwEfHj94dP8UhKvZWSJ0LyoeWhCQ/mZZoFj1ALeJG39d7Irc9RXtwrk3bo
FrIKkK20XPQvV2K9xnJVkxu2p4HfS3jR1WD+PPeKNkE86A5cNe9i4Q0Cbp/SFeukFJWQl+0BdelM
ierRBfyYARYlBhfk7O1kuJui217Q1epYougT9u3Ua+V9jwxtyDsbvIhifBFlkf5okhLIaj4PG1pe
kcWPQS808ZwmBamJSzukiPc5LvYW80uSFfGSGvN7QioG3JOswGQycCmVXuTVdjwsAgIIsU254xNB
FWqHyMlCZnu4KejS/4HlgxAE+k8zGW1ADVhf7OXALJe6MUlNlhfCkyPjSYPWCGWahEOXqqkPmSIU
36YUK4waCE990tJQ5n8c4504FxP+M5TuSYICzb03XsbSGdPf/F2LQfTDrSEUBj3eatJSEIaJ7fEl
e5MpJrrk39/zaGPKhY5dgHyh6T1yVPs+s+jPsSWE8fmunQA4bHmJ7Dxu4lioOuMTm1LcvsMNvxCG
MGk9R8zw7ft3l1+e1NTSJLWcMb10IHqouBw7crMUUQv2WqX7qb3oIpf0X1CIbUSiGyej/NFM0zzS
UWEEIcwGVhVo8+7lqLYCgmfRcXDuWG6jr5a3mpzfv6P2jJss8GG08LRgYNvuc0GBeTBUPt1SujOI
L9RwuWrat7WUgCUOhLxCEwDvKs+57e3sfYP3Fdnsp7zhJr4qojtNJb3WmN/fQ0cQ+dpR+vpH34BP
B0J5qHbRJM6HuC3LSAKTaCAbr/U2/bLnxmhtBYVRcU4+CRsVzGCdM9e0DZf3P9Ox9Rf0gB6LrmUG
+j3Oq2csyYnAk2UvVlJGwgR8WJAretcH8fuVmrb4gd12Qdfl3AxhYTkdWAzzL16m9VAZ0PsXhB8R
lo40qYkAxro+QUhGd961Ekb53pB4xMUW7WKLdZKkHzUhXNFKZB9ogRff0rODdtrV8t7aPPSEyl4o
Y97x5oAJYYi1LnDQ4WDtO01IqhLcTodnD3PZ+Jj+wDeefS+/7BBqfPZMISiTvDO+sC1mRIqxxPgo
pMl0hPvsWalSWlCJJkgSgSTofcmpdkpE3zU0mFAVqApU/J1zxzYdAdFm3vwV+qbcal2sBbC0nZJj
dIjsMwPJQOLrBnySKSxpVqSmbFt1gyjdzrifVYny/dhEl9XtVrPOME9s3duekRjd7MUJvSaUJkrl
GHCX8xvrZ+v5K7aQKMLD32oWbyHGKbIoKi43pmcRAgDc938nHu44Yt6VTJK8H+oNaUW33PUAXBe9
Jl03QuRnaMXliEVpGfN8nEXeqbpyl5EQC4zIPZxIuXM4VDXn6bLHrb+x1F9xj9m9wK5Ge+deaDGB
brKFLWMRtMoF20a5Vy8u03C0JOVI6uhu0pC/VbcjKtQygGffAjpFi6KTw+0b5tNblwfEvClDiVGZ
ElYxtyvpxWJVJWipZwWP9HpQiuNQX7/ntrQhzx8laQXMYCkmNZQAAObfS6VMXUg4SJhxdO1uyMRJ
WqqSp3UskUzdRThWarJueXOFDwPnx0lwIycoUp/h2GdOBPnD0RYMu8oM1SjyIdJybIK36PvSngHY
yaVrg0gsweeIN6lz29Hpz9XA3facpGMXqug9wKpICw73q/cT+hfvy0C4+0blNsRWL74XqYVPztRJ
WrAtqeVnOVQdBBtkZzRDV2GQ4Merfm0mGNz9OLy3LxoO2dLuv8Yh6pZFtPXdlRHMwqSsH4JZsXal
/pBDWrwvTfCoSf5TU2wn+QJW3aTvJ1jjxjPvAoQwX0Xh4+OCzxc1NEn+ecaQYqI3LC31wkWnzhH4
2Me3NnI1Me3BabdG2dailj+3sO0SjsZtDtRTICsRHMrZxZqFRlowaxOno95czncdB46aIWFSYL4E
dKfiX4mW2l4vFbGlM7pQwsGEHvwnmUA4AbMft1wgjsYAL7laxEaxNKVvnJpnR/BNjDb7++6jYkUC
s9/bQxWywbCDxyQRPnSfyjTF1x33TjMYUwDxao+kAnGUCVdV0ltT4xSdjGhlGfOCc42CB0iGoGG5
ME15OtppACWWWCzbStxV8x0sdAcfbamVEDCLDV/wHl+f24Re6ydG5X4LZNjhgMBX+E30YPzEgO5p
hNmXofx1On2mroYLf8Aba7yChZXSDgEPEZUdrkApvlHswKl+3ik1F6vu+ImWmcuu6D697oMSJX1Q
QSoQGerF+7wQTZdotcSqCE0Ri8EUUVQ0S4Q8AmzE3x/BAC4dUwmNwS0DgA8pYkcJEL9ufY3vuQLF
sXm8Eo2CalO0LbenSnI/ynleo5sK5YN7U/Gsiw/y47JUCZtW5uYrDnMUV5Nl/6/pMJdNZuzpJC9I
kkG7Bwx5pM2piP1Sh1v0nKLynamumiB9FTkZZ8chi6Yx9qy7xTro6IRsbhDezXyBIDOgDlP085Ei
7qN0XgX2Ve/+66o2SBp1irlACLNr1Gpy+OreJlV5qKemNMkh/Qzcsly1o7ekCDbKGpfWwNnnklPw
xPk75pCTcLkrkEw6Sd3CfgwdKbrDb+ywSrAzRg8Lcw3WF/amzTRdmmf+vpSFwUkFGg4yDT7qAICA
egqgBthqH2YOAIt1MQ3Ecgx82CQIZyg3LELOtzlTJEJ5AgXqwzD6UfxGOPdfG9tyIkPUC3f7KsZ+
+1kx6dlasW0l/orc7FPt9ERMrzS7B0BD6/NA/mV3cfR40danEFNQslndhNtGN7kerU0L+0zsO+T9
TzJkVTSzTQkxrThypi9hWJqK9BdK1dfDOUKYU3OfvNabSemluofSw46sPpSmeTUUeEZAUrMVCAPr
um4wwssrS4/pkzcH8LULJgAWQ36M3fwkjjUdf5+0yOgMIDowntuyizn++h+M9GtA88ja7jxk5rEr
E1rGUs/Hz3LWNbJUktPR6HUZFGVv9SrmcpeOwxhraIgpZ9f5Ceqiw2q9sWP3IqcMC6wSUj8NUVuO
saCMmFMctK6vp8m2NPBQ3LaaPyGf6GVKVW3aArpq7taG93lpI7hMK1NwfbEhECmtZmXZQVNJ4xwQ
eULYashQridjf7cBXUGB6zWWLoCceSNKmMUeQWmHPcDIN/IO0YYunSVgjJm90mHYHaWdLQRMveqs
lyE47IkMuPZdI+sALnH3NfjZpKs563uZTAbn08jUgSPzKjrSo/y1EvPlnzbzCAc15JfqOctpVSLG
fW8Gvg2gYGJv72V9qyw8GNRzmKfipf4y55Cu6eTSL7WjklvkDnzh/lddxZAsws+M/RSHPnWlKaZB
VquV6BoTq+BYW+HfUct4v5tdR9kItA2bA9yTjUXmqeNy+ctTxhQNDIcuMSq5+WHwvrR1GX49Dlti
g1YjelanlGWPv446qSW8tHEIo6oekWm1lgfowCVqkZeiPu8R3lKxKiuKTsOIyA84ngSOP1gh3+tg
0eK4f3lKNuRgNmuBccTh8IvIWDso5aq8Nk7syx8mosi6xgFa+0IQGIK6N+cSGmq7rxsB6MsH1IH4
ZPgX06j5QX5hmFMZ0kIMwaDzyX6QMkDI8ZX6RH+/jq4C1/mT/dCIKbdvhdfdQNi60mVWOIzzMi8t
PpiBTyurSSxDgX4bcxriuAjzaFICcek1/JaPmcQhG+JKjcga8zLvBe+K5gmPijCUksxZtEq/bmDb
FnXsd4rBqiMIt7oaQIOruWJfKpi9HibdKLFfT5gI9M54Z/gTTGu2MBlmafe4QL4Pwmb2SlyMKpGj
ahI+79jqjlRJ7SVRNw71j40f0EmtWmZCodwQrXkBxhF7dE89HaPKbXhEvszL1nqqbcxlxaVWTppR
E16lt5nSfP6bsQv2oHXaT4tR0yuGXNbStHYesy/FZmkdcr7qdNQ/9MyQSqlUal2mLdez0EX1JESW
vSl+7ndB0LYDDFzEVbzBxoKbAEwekmByLQ7lMqQePnvojF/Wm5kK2C059F0CQgEMlv5udgwC0TMv
waiSOiv04Fn7q1MccFleeodZu2RghALkW+HxQj9+/6b/V/Egq0NjLPOResXlq0+4pq9tI8BAk5wK
St9FtKapAdgzqLDPTe6UddCUGF0hkBZu7lxdV7oSc3bXQeSR2p7+J6I+odu8Z0s+OeYxkfy3h1mw
0ZZdiHZl3OyixdS6oqQZ+Nve3usek3C7JnqF0ObYhe1hJSozROGNh75WXoYERCw5HdL+y4Kq6hi1
q8/Q2o4fdgDWQL4Zw5rBkn+s6QoJaDqCM/gcHzQTnUj/CvQrpcCRgH2RWNTubKcHjSpa6cyNEZPH
pRWJPLXS7XO1RhwZMAOUmFcNOsUMrkqvjEm12RcP8h/eHqOT3xYsRFgDGsvkaJBtn26+6ix/2YZ4
tWXvExxiJjyweAwFVwXJJsBv4oRDo022ZjDNT6tsLtzRI3htJZZ9zyHtZMBqzbahWD1si/j8wOfZ
xl6ncyHuZhJRXQxleC3+CdE93PpPXRSOJvvim/s+mZDre243Bt7B+pe+If8dZuKm3iGYt+kZo8Uz
Oe3C58x8moKrprRdiuCY53cQ1VnLSfcUGi4jSopa88HfU/HCwjDdafNiy7W3cox46pI8ppvp66wl
953nXMARUo/LTbyQY0Kbj4tSE/op44nq6bH2+CmNZ6SmFjuFJNjAk1V0VD+55Vkn2x5UXndsgm3s
9jCnnHPge+VOj3BTs7nCE0cPVDFdDZMC5u3EzPdVvogLzXEptMxEezy4HWhvWxztBQsT50ulqDL8
DnB1D4PHFQOblGKNCxaBfo8saIxc/mtYL+h3oQeqaVcsTQS1RxPp3HPIZAZ6uxQEF6sDoMcuEx4G
7U80puUyX0AXT6ejA7dvfHaUocilDWcTdTaySw37Vtq5qT5k/WqkwORD+0Sx0aw/y6nXHcjEpqEE
GftJ5vU4WXIQCCna8Ia3BwQkvbDeNGUux72SIr18dl5c5Z20MZeVVIsVPVkTgcXtcZlyYtrljivc
p5NnkEyItEexkV9FKYWpE9SUCXncGe2gR2beE4NJthwMe23l14GgbhfJuvN1zFgtqZ2i9LuDKovP
vRiucllqMXqD7rZyznCd3TxjAJ6bhPiIobHTH4hbg45HHsc4yg6YyaSxMIj4bm/Qfz0EnEv5Lzq8
hPdLUULvDX+XgcCbyFpdc9cex2WF8sBu4gNiSWLWT/1ncfTgYkWOLdr6tiv6l0f5sovlf1KHhy9f
C6j3pVIcBL7E3A0/mv4JZcUccKZdeksLtg8MPVH6GDQoqSzgc52j/fM7str911aF4FTJgC0p7X/T
K66+nnqQYpVxxXWRs91Kn6Pa5Dfc/ep4LAkBb3g3xBC16h7R84+fcvY32mMfPLLEo1TdNieDbb27
qLopuC6mlKbO6P/8LEHGRqTEOrloUfL2YlndO6IJdkcDRSuKgZPFH8YYpiPFfn7tip+QDlonbq75
YbQd2FZUXdasshdRBekzGziGONf68Ie+EU+OT3VeFOwltb3aaeRD4G+NOSiNJ7JpNgK7ykMEK+dd
c9lpr3YqJLzJqwq/eIJbglnxV7UecdmmkZPO9n6ncRrY3TZyTK71plUIC72aj9iXXh0Ka+Nl62Vr
tqAmVQH+g343o7cCvVfK0S2+iGMHv9qhCEuryVssNWzLZTpJEK6A/DzlBuIFfed4T+YoWc/ovhaV
o6WfCKRcnlmCESYYW3RjvjSgJ+w87I8YV81uDsIfydpQG8tgq/Ki0zEddsKjH/9YF5Rfsa+Ho2Z4
pSBKpdp2JVQAE7VK6cDj/jmsA8XoVyxrsOiaybLLrdm9OxEXtgU+Tb6SLwCddewvGDsMwdL0CtN/
HkMI8sAU4t1FBbRAC9LWaOSzyb3DPOYt8K/kYN9d6gumWwYMcsXBSYIYdakqTHbae/Hx3M+sXQSq
xbZznXZbMCAAG9IXwv4hRypeuM7vaQowe2FX6VRFhYma5yVxjmXlXQ2vrkeffpA/JW3aYcBeG1IG
eQsCdKvIFx2dhZPDB4x5mahWrzg5MzdWvyLzaEbVGIpUA2d0ZCyLeog5F25sExMPvUkJe6d9qi79
5Hlfb2LrusG8u6hTfFho1iwy6G9pLPHudmCmKoHIxZCHcU1h2lJY3sYPesX/H/R9uIXKJCOuGCr+
NEtVzCTL49u2H3FpwN6o7saL+xpNqwphBi+thzWrtx7HPrPX1o0urPWJg3VLjs682TyJIsiThKEK
obK/cpkdoAHYLQwXHynCnbN/PHstekdd2KuMx/0vWw/eAgmrk5SFqQssKGWCGVHIwfL6c8CZdGVU
9xB5BHYCMLvS08+e1wBGnp+VZxEbagdHLW8aU7k1rPNffhUg3HV6mhzNuRelKyRNretfQ+rsen29
fqkTvA+GwiqUpgfHEe+61aG8IddevZMpTKlBrQQ3E8QT529mooP/U10eptMiZHJxIQWZkk0c1Kyy
+3jrr5RMdllgzB6D472us2a4CMZqgo/ruB6EOZlK3Rp/Zct1LzCkifHzNOUpvLN+Mc6ljS8si+Pg
AbGySM9HFVysNKQY7TAk8wS3KoVxBkmFEm8mHyKX8j0DuGVY1FoYqYhT8/yKplT7D2cJSGdWWFWn
STbaQM52SgfIXTofSmP9DxP7KS7N97JqXMG5+N+YfCaN/p0jhhUDVeijjvooTDHMNr0Uj6/5UT80
nL1uQ31F3HVjyEAaiDUa3YQneB1l+uLCUuLR6Xrc3Re0eU3wS/cd7Jsow8Ikpu+gHesPut2g2iYS
/2TFw+nVQ37JfuN6HwqkIH9JR0wzacv/+dZwXUEAnPYDattGZJW/cjaHhnfuIMgPSeInPXj3f+Xn
kDR3E4jyUe3CIs+8EekdmBC8yhudfHiZ+odENyHQgcHoU3IQPATv5zijIYXkaynNf09R9JtVHa6Q
/re4JpyRZpjraVZBVd28tZwQAdYYzxhI9GGKoypmGedjgQun3epANiefox8TprmI5pY3xvjl7/af
1/kSibhZHn2Gu/wCeLB9uVaHvMBuLcHOzokHZw1XLgxytx2g5sQf2Isjga86KTBDnVjp/MnQY+j6
/7+JVVhgVj6MGvEqc2P/GWy7y+wsf+EumKuuBNLEruaNavq46dkwUNcVDItWSddl/+jQbrdb4zZz
/jrC+Oo1IP8Kx4Vs/JjaWBumRuefKwAye02QdFp5udeAkwB+Qqg3OjBPVRSSXDF+ZfOy/AMFfhnS
2bS2KwAB170/lhajUkAU+TCRIPdIQBg2qrVwNMJ5IdcflbnBest+Wqy9ehmoQvUtkg3V4fp/ooa7
lmeXjnEKdoMhZKSkvpXRzAXyXhWn8UiARW0CcGSTosyPaNCLI2FwEZr81uDmRj6JUu1L5kR/V4g9
wrbhWfLE49d3Szsu2HrNO8LTZQsQpLMpTTzlIbGINV4fw1QWAeExNfM9J+qnD+zw6zmVf/T1g+ap
OWBFDyvZH1O4p1OFb4Gs1xsPQdJVz+fndzp82YY8NNEi4NUdwLSkDOd92TcaFJl8yIUzB6N0h+Xd
csDPzKPe0OeJBMLZyBs5+VYO6nzdakRl575oCRWd8EcKayNwU6xZ+Ys5+YWGsFxWci0r8sHHREzD
/haW91X9KkIdlDVeuMQ7M0gagrqgi6KS+oh3kZs01N2m1wr1gY72Jih+FXNig88215vRyDcF16cG
KM3SvZ73v+wwBRfpjDJsDzgMyv/h4Zrr4wQllyxvregnoy4d7LktX5IVjvmbbegMv7VcIZ/0lVOY
TCbs0PnU98CAJ8MO1RyG/v0ES/BVk/YEZhk2iBqbnExKEegCd8wWG8omLhASv8TxvSpKM+rPjaf2
dqKyGnbMmk7OS68mj6/0Lq38GvdDzLL70yJGTu4joB+OrdR5tNh5JP8XlrwXAJzAqnZXEJ24DzLQ
lH0h2mjQg6iJ9hCef5WMMzdQU6zBG4t3oGC/7oxwVAxwokqf2JPr7lnE6AohHS0jdS+mnwuOEPp1
x2skAbEShDJxFbhEAawIPiiCHaeUc3KP2ulN4DfGPMh+iAoqhRy6i2/oMCWU+ZsxTLoauaoL3ebx
xxBj7FBk6QzBcQObDK9XvJPsK86Fyngx2OkYeVocRjF5eoRgvtpNl0aT83UmjhpJNH97C3SPDTru
Zzr6Z94A4YsKRdDmgIrLJi+UI/U9jzzciin8+Ey/1y6uSzXtvaPqpud3j8ZMI2kAYZT9vS0Ry8YC
DGN7vt+1L/KiqN8gLG+Ti39FqU0SVdU9ROancGNbNSoOCZxGvWMY3vsvAiWtRt0k47AqpPUrGX0y
0Em+t29jeCP5+7JuTADfbQL1tiwFalwrsBQyEqT4KrQFUT5gL5U1zVPrj1HzCssrwAkvuACpcIb2
FsTXuZ8UX1kFUOFmyzaAmzZ60/Dpu9uNVcG35FDP5ZZLrPLDO5cUts2t8wmcVKeqMTPSVWlPTFFe
b+hIO2SIOqZCc+gJJQpTdXaMAWhSpz0xQolg1x9xS6uQMi4EyqfEzKClMT792I5eeJOqCYoDzGI4
1O2Oxdh8LfmO2njXQ1Dp3Vgr1Nf6/FQHpd2kzyEzo5Nd3JQIU6gMicTngwIoallqESf9DxDlt+pe
SBB4QESfNy2nelvYbFwbRGeMdi1+1pMaKvjQ4+EhuNuFq1KD3kU17OG/jjIFktAR31fYy3G8laba
1sTan0q0QruslXaSnVYF7Asemgm8MuNqaEUI8k5910VBMxSq1NLzu0fbhggZ3Pp80IiK9TCbOxxZ
xpXed5zVeV+U3Wln410S6qAhQu4DxxzS+psqhWMv7wmyJdCQcnCkNAfaM7ZlIWS9afIZmnacYW3k
ryUDMmpoi6axgB4fEk8i3OeyHRt9HWBdTRL3oYknfIEV34xQqFLX4t5IJ0tAXflI7TF7MGNAdsot
4vz7ZugSyU9RZYw55BFnVvI/k8MqeVifDsILQKFYuFZpfJNx3VWShAYgvIZxovFeTFcu680C3Kri
zz1yaNIs087/JRzguEcQPbdJZikRuYE7ruFUaGysSAODcwrDj7A5TzxN14xcDjmGltNNe141zh03
iaZvTOPcl6Ww6hdP3eRfqblSEDgCOZqUK+EzM+xD3mahwV2pHHAhuqGjTorw0orRxJY8yC4H+hJZ
OoSYKyFxc6uSkITrsWiaVdBFZoV8QXvXxiyyJ+bM7turiXhmFI6jk6lPOdi6PcQ1Txc5NPmvWpgp
b2/Ie+xuZ7qOJjsq2hmCO8MnWIUm8t6MveD9hW5xcR2u7pyNYnsBq1a/2CtRkoIn2UNHrYnRGq8/
DHj9+eddCs6w7jvBEHx6HScDtGEMNjiDGVIlQcaU7u8577XtE18ywdE3ljxlzDi1lUhmYnlDbGMr
+Nt5GHzsvsZg8iol+/AJSQMoL5WU8L42e6IrJL1MS1ZLm/u3MFsZM5nybwZfU6svUwpqLv6mS0fS
rIEBPd0t11f/j6+CG5rOwJsrAzU6XY3ZgpL0NjvCl77uC9PTX8lJU7VMdyGRcz54Tv1h1f4aMO97
j2XELRQ1agZ1uwy1OI2yo5IrPpGL0y9nH/1S1uZhd5bBKZgirmX1ks2NK/FZ3jseXzMWaCMGg0rN
4jVa4urtTVJsErB/lwNUCvqeSK4JC/Xm+WON2yrI7/tjWQWJu73+JKU9yCfKpia7rsbVtCKn9Ctt
nvDa5LeePtata9Otc5InnuJaD1BgpTTSDLqTRQjf0yd/hmBtyGA8xyz5G8wJEUFzoPP3Uh5/ByOM
9qw2NTWFiMSLhg/OM0RA5YsJ93E65iZGD4cEfZ7zNzAPr+Wuo8w8zVIDszhNaDpxgu8nxQCluopt
0LH4IX4D1jTUh2TE/qJd4se4oxv6yUoPSjcO/trixUZ0EdNmmLwjG3RlIFDYZJFz2hD2kaKQhzhr
S835Db0Fcu0j9HPqdvlCYuyzDVLwOkQeYTfXjUkOO8S19oUis2RW/PqVZLlF5h74vzaRsCZSO0Qz
NvLrC7CKUHAZfBiNtnJBOzEbTCMEpJypiX2G8CrUKLKfJ3YQik8fz87nneshA+ZZidnY6QZtkEL9
xXkZjFhpQVi3ukDjuPw310gXbzKbKnpTj8Aml6fvZfmFTM5SJPAyNvZaFVMa+PUaN7ADNkPSV+sd
kR/6vyd8suvcn5AThOqASH/RID3vRlFldwAyjFNjKz9E7zgLE8wC+ULBMWSL3Azo8vsUzuxSv6Bi
U56B0Kx3JndpSSOttoFzPWCqg6AKOYFzgkmPhR0e/q0zvxaOgdGsAx6imRVCqdSHkjLupBgrIWHN
bNcJdcz+NaN1UnjEBZkS3r/rIIdfGBsHvQ0g/IwKP4z/cXgPoLtEJs81WANq4Gr0hvD9EJcePMmi
ipiyD3t7GUBpsrfIazBb7U/9qOkbUQ1EsHKDbjL4B1bsm9+riYvKNh75mW+4dpscdexigO45fleq
MyeZAEv+5rGEdgofQl7Ms36rVckKEIAmYs9VN/TgA4a4y0c7BIOiCQ4T8+9nl6erJ+W8U4a9FfAB
t4npFyImnNrSizWDg0PxTPjblx9T1JMt5IuTsdijxQSsLHk/kxvOO9fl9oCf7CZhy1BkQjLlunw3
Pm95vJKopIPojjagJpruDTM9VA02Z4WMHuFNqTImlBxwawJ3Rrigc1WJ4HDO8dblTPHyMy7NwP5b
O5yi8UeI15g9z9tWTlts+DycII/uecZAgPjOjkR7jfPOPYzIkgkczkwrMcV0VLbMg4bISH0GSLxV
JDTSbPqHVSWFdnSf/P2NNnuWpQqZFx5fIfrU4CpZiMbX9+UvBfDaI4FtTaG6vSfrZUXebbOYlcex
4Pn+/yUtAvjXzLZ1nsNGpu/OVN30zvPes6hi+Dx2W2pP+ExOwAvrqqXNJGuHBPakuxV5yjo3zW4M
Z3/Yd2SoXbXaTZYsdj17eE2hn1tVIi0D1JMQ8iD5Srs8bR3i7J0QcyQI3Eo1hBtaruuZrvitvIcD
XkL56THELl3BTCZihWWbBLK4HrFKUGxmYiTo0kUiW5eVO5cxrulZnwPJkhT3U870vMCca9VFuiU8
zy6wGxjNaQUkvhBGiiK5WkEmcH/zA5aDKJGekGVy2B0mqGYO5y9kpez+4YKcF46v426OvHVtABAG
RLlSFKf6urskCShhe2POyrKMxoh0hsOxiEg2UoC8hmeMu+WtOOdg6INjs036sfoWpAS7+6LMnczd
MiR/5+OFvx5e4edSgr6ijSD2ULeapbneJQYTpZROj7dRDZehfHSPkcLL8UFjomtRy6H9GPOsyhqi
1OJfY7l3ya4Ekp0Dzj8O/6TgQWi02C7FOajW1c/ToM3Zp1zTWu6anr7KC0gkfJuZocH2TSF1nkmr
NZG8gFHL5ZeAkZRJexPi3yVfIyVNxA1eWUMi/4p9s9i7vgzx2HBWfdCtc3CP5vKOrCuEQImFAh9A
oA5hvoHV944vDwOlhAG1nHUuankky9/RrW9l5rz/D6TckySIMu/uFElTHFxREXT5SGYdqzOhaKmi
s1SmPGOduwVl2hMSxiGGXT4QRpzC06hVJbVdnnpWGpCK6r4JlBmW7qBZxnx7piD0AhT0QWDwLth6
+dy6IbUNRHE0yeykwY3MNaKdLRGJnGV5Ksjoy5kUK4W6I8bP0bVY1zs8YDooB6OdJS6FeJ8L3DvW
o2AAJroh3qlFduRADpIFoyISTBjxo6gvNzHdba0eWv3XaKkRM/6VE66XRiSEsNgI5i+OgwW5BNbe
YPJyHZsiqwKPg3SyZ38J2OhtU8LsZpz8O/Jc0fgNAa2B6mWk8u80cI1OEG1SlJ8LDQ+NoIpUUUVP
LNZQDfBDTXk3TgsIylfL0klPWFJZ0yT7LwpacEIqOYBX+T4QlLyjpvc19EuIQF2TxzGTCmKRt4wj
clxOXYirdA9jo5ZM6X1GBdRhuGXAEzNrQDC2AkD+sVSq7RZ0GMJsJIW6LdMF2HtNLYzjUUiqHKaZ
xDLKF5TXGoGNzzN7gHGwkY9RJilEuKQl3+YzcwujachJPghfzgqcRcE71gdABlNDVtWjaNZH+eBJ
txBrV7v61HHVHmWXpwSzXlvI0whLoJJkRwI1qKkY/k8nAA6WxV6rrHcjrHmv2zgeu9y1Y3eSQk6f
TCF1b0eqwfpovQO14lbf+lrflQGh5CqOexJheClXB+pvd6GGmGpl39v8R67qo5VZX1SVyQe2FcMu
RZN1nkgHAKpnSGLafiQ1Dsn3hw9a31DVBqQmP5QAOqd893vMhOt69ber9W0w3fr1YVhMN8nzDkTe
kDHuRpiGgfIRz4LF9HcXDGzZNMPBsI6/x7g2aFfeO1kAqxap5ZYSgE4reb7XQeuMSGRYwzD7Pj6k
tdKie6IYf6dcXty/600FUjr7qiroqgtHvjKg6Nu3BHs17QInvm2ch7quEoqD0DCfHnKLL8TtVm1R
c854s0tDSzqqkSz0IYef7aHLe/GgmBeo7hud5S2XT++g719AmScW7/yoLNqAM3NJkT80qWd8XHyc
PyIf6n0fjtOh0cTBtHYE2aXmPILoV3HJxfVKk5cI/L8j7kQq107GrEWy87m8fvg0UhzQKBP84amT
60AYlUhdAterop4cn2htLwDAgVvVx7+7j1X3tvfAq1wk+A+dZBan19L/oIS4ZcOyRY2R0xji1XEv
QxlOFYkMvYPdyVLZqwutpJbDKxrG4Xnd/V2JPK5gfaLWWhVv0xCpdAX8n+c/tJIgNmxImTzkrsNY
ZudkGDuOXFg8gBy5rmXDiNUxhsZkumpQfgXbLQF2366jpGmjgW7B73za5aDL9xaSqll/REa4C4q8
I1kWMsCSn9vhTCoCDuSPTN0b1JF/qsEAtq+ooxvfwZVmzQ/t1MN2KvG2ISGhkrCIGKwhUGhAuTdI
cFXlDShOPQKJNGnzeVEcI6cWYSbJo9CDrjGsnmn8J4DT2uxqmV1s+QMx+o9mbX7vJneYr23d53AQ
+bYohT2XZb5r3HD2Amiyl/DO8FbX3q0FO4yqNG0euXZ/iqsgJirRL1d/NSELcfcy2rhL2Cbj+GCY
AV7Kl9I6CL+zBin0zk3tecoFI/FuL2YpPSQDy19pJJ7ZHXMO+Q8aFF9wG832aVST2izhRysioWQe
M1cr4wVn+qJs66kLZxMxr4AoPMT5uFlnXxioadfuRH0GkgT6rNLhA7snCciuOr1ZIdGMVacQUlmT
A4oOC5Ox9iHWfL81YSuZDgQJdacAE5YPKZ9xB6FbbzD/h0gi0q4a1hYtpi5sAYvFLfC6+0V/ZfJa
3Pzp9NOH8m3KnlJdx68X8LAKBrykoRh5ME5G8/vlN09AI5POk14meWwT9mJIZekMpZErOr1y8ggy
wKR1Viber42pBlWX15XdDGBzyMfZF2UzquT+8P6AfslbjuKPaxH1fiJ19T+fIlT9ydJuFIVNsdpF
Uio6wHDzbKDgd1JnqMhRlUPm+0zd+CDOcG/EfyFQYd2pGZsMqvFgnu5Pv1aJkOyi3jCUxRKVAxk1
HaCDARxqDhihwCguf+BrRHplyqtTR7RTHeD4XVF6Bt4yJvO9e04l8jlfSx4Ol/wYVN7XTKXSoSiF
/nLRn7Z3SqaTKeLz1bhzld7rVeVJ1t9cbcDvacb+cNwwMzSz8qAKlu+froTOQVGuWK50LvajuBZ0
rG/yjWzBUwdHrIvvulk8Or7+y2ecp2p4mUFAI1qEfN+qUF9tYkbp4mChS2QvsbmwlwWbXhzT/9cr
0WyRaVGv64DrSVJaEQofMP5T+vU1S1zOeDxgGj/4FGUhclXTkK5NfsuQaJfy9qImbtC0sS1aSXJO
LhsEfEFFUHBqWPrZmz+Ece3qSEYcFkvcE1fq4XZrad18V4/AABifK1EWHYMzbICjsP+i9YSNx+zB
3VrxMDZsNcpTbX/GG1hjKkbEEIojXX7jajBD9M36PyggQT4K/5huATW4Mf5j08bTmF9rqzrxRoJI
NtnTEIS+63sXrOTiGQWzsWbSZDeHbTy9W1mJxbyfjYTww/t674iHx9nE3QwxjP4E/aDgrGjsqGQL
/ODhHfrNkgUjpm6pTE++FAJZsfbL4hQcULBk81AC/sy+TFJfXNNPri7t0EcfEAptrC3nxsKIpq+W
Gy/giNBjbXSXPA6nq5lOicEGXhmi5RFTiFe8IgxLR1uySes3dhnUeF0bqi41+3NAEuwNDzdc6jZn
vzOE0syE5vSG1q092ocvnJ3pdeE0PeWel6MQsa1N8E/4Gpi9BDWU5lLKZFf3XwWOG6ywOSgYaO1T
Os93lNg0GzpE5JbkIqMSdXBiFxmKTreCl4VdyUxvpZ2KIDAukaJMgNvB4UhiXyrg2G2lRC1xOvzf
DQdvf3fnwx6QpfxX7JyZE5jQQJYiGuQxNF55IegoAFVNIz8HIvJ9Gzc6XhBGzp8C3JMIXJTmbSJc
bpFi0DpfXSg9KR/f1B7Z8WH/CMUndgw0KrZlIaZq46GSmd+LeYW3fv5SZJ35KyUj36c4AuAJDK/3
XW4DSK3VaNl09NIyzX5mbG9Gr4nwh+W/ZOvU1ZH5WHP0peMLPGKnPboyYpjmB8n2SpUgNlGknojY
7ZaVErG61FglRTQjU7hU9E1erm3S8dZ/wy0y7yd30VysFjc/qkmomha/NEGWQGp5Yl1VflPHhVRw
qPB2ymPoyW3uhk06n9+tIbOSEaYdxId880JeMKwVag0loUjD++ZWgBTy8PHlCyfpSaUokp4JU4le
HfnqhVeFJKGwSfESSsasWA2RuFEeHzl1l4VRCcOLvzimItJzuMVsZrymS9tubH3LbUE/lSE+uhnW
snYe9BUlJFcl+9kBsQoRQNL9cDbDYfERrlMz8Bjm/+mKWddR83TyhBaXAilNyzIZLIIiDSAIOY9F
1UaBR6peBXJq0JVdr+c7T7eGQ7TWRDG+sFLkDsBDnguQ1XGgK9MIVE0iPPvcxH55U0RqEuDHsb9I
YDYspQfIFrWeZ8uMx5B/dlt2jDshr7YBukOgiasW5NeQVlhPbgNV5tOiq6V+sEQVjCy2sRIUWEkt
Hr8A4E52f9I+X+FQhkZifThombh022IKZJ1O+Bn4SFnYVkLbh5tcXmrtJPPskST3d9Ij+16Voojr
wOpwKBeH6o+sQ8S6QZvWJokYnJwP4LTEqX7API/BlHxE9z7pDc8iWgROTyn3M327m62Ry7JCAVAi
ic+ZtoSoj74UDdsdwiBPuns4814RILtzC93VkbqOemrCwpyYhIMPNoOqv5wZOQKoL0AH0IK6FR/j
fVVLqYwqM1tOtiV67FTDgWbR2ADIfGjNndvv88S23eTEX8daIXhPzhG5thLTjScR5ZWxmmgI8Vmw
fk0NN9+2a/X8HDMc1OX7sjLge2KSHnUd+6vs+LYhrVPG2xZis3I7nxWZbHpZL5bnFDSPAyNSQcjH
eFH2tOvgoamsHHE28MD+SXs/xG6F+DHDbkoarHn4rf3zeNiapnML+qEioOP4Zt19KcIM2UMAclru
kKAdhVIcHYarE+uyTQGTRY7bDbEW+MJRQpXdder9NNH/2ORtHqPsB9A69ZRJCQH1ncT/KQ0BYB4C
nKCEX50mUS4qXunXDHHfSpo8i8hfLqmEb4u2xiDT0UTDKMAWcCAFf6TgDbfPDa1+I38m4J1o8zd8
RRLeX9+f2Ny6tAgtlPsJEimcTXbW3cHCn37XdqgMYOU2J5H9UMJ8oKTkMV8va+gSE1XfHkVtLTf3
He0sbn4wt1ePf2pze6Q9AokdIFE/ca0etHZjgXwZm9+DPDi16FZcWXwso6XfZwGg7uw5O9ciRlrM
wPpz8h+BWOqxdEpJF3Z1Xb2HwpUKYBl9L5xgyyuGGGgBSOOHRLuQE2oeecunpuc0MPzlJIyJEgHb
JHyNXhplRuQ0+g7ZVcC/pCWlB8xpCfYRzQxvBsh1lUAtj6s95VgfkwBdQJUsX7n4y3xELDfZbKfp
DMPL02ctIn/HB7H3VmEqombWh9+sbUQxLJDqWq95fT6sp+l7bvPsc+bnqoQe/EVU9WXrScHzkQGT
W64fFCMC6215/oS7SwzYxlSb2NcelnGk2LnwSwfYOXj4gTQckuz+dHcArBHArRjzCoN9L5GuPDmp
Yrmu9ngVuchPE6C7RsfduXhhzZ/2OHsjYyXfrYGvLIOnzRp4g4kw/9j4SkB/QtKi62E+EZ8dHt3M
KFk1diJIRAVG7zKGfQAKapf4LV75ioGsauG+KvrRDbEPs7LIbKrDY3/oNkUJm6CDOo9uW6C6lT9r
ZDZ8HfOSD/SRIo3p+/xFasbHl2uEZQj7hkXgucocLS3y3UPfZ/MZO7gYba5fKa3o4NfZQu1dbY52
Ximd1kPGheHKfnb9CjquM/5xCDFIThbwYsMgoWPnObAsYlHuaqoGSZo/0Ss691+UtAOA2QINkxna
nS32AAWh6qqgO8K0nGuVIwp2nQUETpLz3s1sKChcRgZabNHm6VAvvuN8+fTzgSrauugLxhOhtRBA
I1MKdXyQDmgtst4iFtS57YjPoVGEtq47ppu4vz29hS9DdWBFf8zu39lUraiPck/DsPPyY7TFEvQr
7UsVVmKqtbbINtMQlkKgjiET8e/Twmk3Xt2+5fnPCps8Ff9ldnCK+SMo6E8jY6RQ5SGobG0nfbJ2
XuJux5pT/JsawxO///NE28R3+HgyMxa/vD4Zw6D7DT7j0p4Z/FcZrTn7GPvE3gNklA1wXVKvfEro
YRkaSMD7SAzIy92TrDTl1ta2Z6fFx8eAhhlC2SYbnt5ZdcUz7AM+U1047KSBZkpKezfuQexbvTh5
Ea2kIEg9zv2vdytBmjLgxgMGp/MF7U7ja6YKnuJu07YXCU6XEGKqZKArP2QlRh1NULpAq3wOYPMW
Z2hEvMs3ahHgAmTEGuxgUhWsU4XS2CyXqz4DeQqzdbYKi1nClldze56B2gbt5C+aoaovuoxY8UnN
ad8zWGKDToCORXEzdV4oMTBUoMcw2yoBo7L/CH4nBB47w8nk2UtAl6Q9GcRxcWmVq2No2v7rVNGA
zk2CbOpHxHhRS6jRQy++ynqJqConruVcX9ctJKPnYxkOEEul7l/ZiqF2EO3sXaST6M6L7SLcd3HH
evZrijLFgMts3xZUyQrfZj3NJ906kCi/W+kl35dWoU8IEoRTiZwsQiiz2UTrKzqFnFexhRiaiP1+
nlOl8EFDnqu6zNMwWoxZSMAquyYXAXLQn1b2Q+T4/0Yz0GgBpDavqXUfmdcq9lP4QiHzTzac+BWn
yZu5jiom8nzDy0fcYh0f7Gx1NWBQhM4VC4UNHTWVY/B8uXBiqE+Yzyy20Qu2JTKZZF4aWMt4dZ8M
0NilpNZX5Ek7o/XFWDvBSMBNuDtJZVxNZ2Y3yi2a1VmExUg4I4Tsr6u4VjMQeBHTSCDuDemckimB
Xxgc+Q7qE6BFsxh8SYiD/fWM1mHoefYoGjFJvCD5Ey2VGt1PHKFNOXA/LEBZqZWR4wrzaiuunq5z
8rNMFuUvJBdlpVmvRtR2OtIWd0ws5QCCadA4EkZ2yfSXpBSQhdsTFzBWxxC5hLRyelLQEFrcyRNG
zd7y7s+kQGFGYHBAHlLVUsT+kRq9yvyJMP1nsUAp2tH6Q2COALcagQlEOegbeBoYMCS6WeFw/0ib
v0wbVvi7zKsY18FLwZYGSJl3oltrEQuNofuXOWc/17WSS43M4sSdPXm5aHUpvk4Fggo3Z9xFJIxs
nwnDQpz78oEJb3ey+DP4EQrPRYeVuJhu6RcmIAnGTtH2UmJG39qsPx849MlFeelzesr/Bo5AIr31
P4Ypl8qhf4+iDkkI/S8ACRRV4LmuHqLMuGTzU5RaOUMik1+a9wzme/Rp03vJymx7IsrJLe5cJ/YR
VFJ09vk/RLNicld+DvQrXTEaiyk/KE2ZXKnzio19FN1+m42VSDLu8ZIdMUSa4swYZThjqnz8LbcJ
+AMiADhg8FJ/5A5bLNdebefe467LUC9Oyd0VfTfSYXCjw5gGi65iUnngHfF1FwK1Wc5CrjQMDWrp
tBtMc+4IO2zXVAl/NcQ1Luq5hXtcTbRE0EYb54KBqWtoJx23YY60EAGb84wm4VW1ksHjJqR52R0C
OFIAXUZSinz4cc8mYCoJ7pf/5F/4tpS2OV9GFLyqU9T+QhxlorjMXWQD5eS9F1HjhIooRYwk/QgL
3WY0blhQheL2n0hnOg8xrbUGYZw6vl2zRSbQzdNheCBK+18k60KcNlNI2PwapRZuxf3NUHLPi7mK
iYsc0tGDJpYgjJQDRWhwG1Es7Iot3lk8r5W0lfX4J6/2bOezjflF8A8dfp2jcuM5tvU21cAezstp
B9uuDEUf3W1kEGH+8arscCnXvn2j5MhcY/aaUCBkI9q5hE94XB9h/ozAu1UiQ68pPa5UAWmghnee
g9ZsmuAzWtmE7q7rvU06cMEudYh1Y/m2ws0qesD5s+MgS3/3ymqQqFpYTGNNjNlgQvvid73fn6ms
lfThyk5WU7l5ZoaRNkfqfwMTJ/z9ai9t9C9Fvg568qevDYlLwGCf1aYuQHMUWDRhmEu+kUUeDSWH
WrazAY+nrYjT61ADEaJf/LRz1unQEzcSigzTQcgu6KuPZiqKLUZaDXIvxun4xod5nAhgEVilk9Sa
EENiOjIRy82CB5AkjgtqYcMIP/G98ECWEF1ylWjyXTHkBGXwUxjvIOeG24D+0jtC7Ei5udI4Vj0u
3e7UhhKikRJacEEqMmtoD/irp+1orVUSdbvFoZ8xM+F19bNUTK+QF3Rxo5eLWkQ/pXlJGKiMhrkR
ssHkZuMDKnuGRq2105KtAml5a9LuJsSID44XGA5+uVhvw/Ik+8z+rgBXFoAZfG7kgLUIDG2xCz6K
nU//rwGrUE7Q5jFuEjkfBEOuTbOX37YYrPY0HTG539BK1B2fo2DR9uNaa4ZlVcbP9hqT+AUt3Fyu
smPR0q4OCbrlKYAxKQcdybnCk5Jni2T469OtdqTpjdUhKRVh4nU0o6s/VshkHJZipGaeLhcZgjar
t85b0LF8Np+0QfKLNvnubu/yezFgImhyblf3j2TD90B56UKSKbfIATuAOuNqmTbtk7JF7HJoBqEt
zisDziucPHAJYLIw+4KntkCw1XG7F15/DOnIU3DIZzprTDkhfv2eKBLNhOQwRWVnHSwql13K0EMJ
aFxbqHl7Lul1Z90pOqdRVYTzFa6mlsP7KtFPHCAAHW64yLzz827fVQV91aO9F8QMOK7JyAh4JZ3x
wKHyV3W9AnsArLxUaHdzjXRv5BGgjA6tBNqDEHUOnkMesYyihnyZaSudMfRV4ZBy7fu2enoh9mvT
UAorGUDUxxiogGgDjxwutx19ntLL37Uh9xl3GRJm7kn7vpI6esxpwp4yrIq/QIsB77TMYnlwVBrZ
vg+w1A4FiAb2tMpaV/jliawqdtqjJYXUZ8Yo8fXmBXZDYi0LHSjJ+13I12Ew9ymX9mvtdZlhSYfK
3EEy3u0DUZeNcjyqc6yqpOw4hGruHpNS0j8G0zQLSfWqt7WVv4zgrpYmHA/Ij9dHkqCScIZPO99k
JCEwja7rspKKdv14go3U2IhZsp3EuXTPhbPvK0HBAAOeZqhd0+mi6+fv8FTVNPf0CUQUfUEFDD7U
Zep68LY7PU5UICo1+7gALoU5bviE4a7ykT3ID4BxWmBTPPiD3OOq3Fvrq746fEDQXhPoVCyxT1sw
QE3Dubcr4ADNdL/+H+/v07FfGmM1QkOumUyQgxDRsjOFFNI0v8X17caFrlifo8I8ZPHWxbM+oJUq
5QMj48sS3uixLUNyWJNhJI31wQrBpZeXWilbkRjZdKhzIv2F3lMuhSMIJmkypw/Z8n2b6h5go2h/
8vcBabc+JFfVZ3s4+5Cxr3rX9SjVkSI9K69wM10pWfU7Q3Z4oheSdkfU4oX3Hj7UJgIFRp5Xp88y
4PAuvGEvaFxUYFiloRKrIkuZBe/RtulJ9gXnRrL4PTmsuhmtFc58NPDFrD1lIBeJXumMeMt1uSuX
0HbzsoIXzeNXjCaM8h3p1AXpXk+Ce3UNLx08M0/VbwrgPrWKdf02BOUVHIC5pMEgdnvFMdiIRx59
tBHnjXyQT8Xhci70nKm6QqbNaP85HIVxW8L5y4fGb5P6r8LstBQsF1ITcGbrEfznVh2Wv1627Znx
fgfrVkNnLpt7I64V8ESYMiB2NkXO44upI3NEASDQ607hjGjTHFdUikEcIzjDtsCawOIZT620AHok
JSX9+JMap05oT4DKqKKehUTLaWeE9D3wDoKmagci1ZUdpHkbznuOT48KLUB0VMVnKbacAkaMpjwu
30t9UUr0OBSK2e9mj/pt3eVauo7kenCUahr4S4FLYWN/X78wJ+7mim0qlMlpd0zdHa/a/Zc3KdnQ
/i0u3qkb+zWVI9x8GOsSYxIw0pzA4BjSzla1bLqT8jmhiUPJskR0MCql5AAXsuqGlRRGCp4M8EjN
wZMmFu5qnF49NFN8XGWj7q12ETkJo2OQziMKn6PoaU1LeEOmlqdf1+RAHyMD+PdBq2ib+hZs5bkl
ro3be6ZsPandGBktnnqvVvVfdgOQim/fZ65+lVyZEXbbZUaEfgXTbduKLxL+nd/Q4cveypde412N
rGovwz9MYU02684Mk/JZd1LsM+EljEY1my1196BKWFOtMh+21xrnT6Fjor9NwDIGUNHhyQpW7EuX
+SRKYTZ0j1OlGYCXag1fTf9ppIfAmaUhF+U7aXs94aU3/fbdBp97sbsvRLbzZmKExNnuOP2CHkTY
4c16gsvQ3vlIXsqEjpJqnw+m2vO8+2W5eBzmcZC1ImIDpQJJAu4IqB+CM/4LMLwWi509i/pX9mPi
VaRTuOQt2CrsF6qje2zlYSRTj2gnUWbxcnEgwIDHLHtTRlrCYTLuYbeIj4em3fRlevGYw/LJbbt3
cQ25nYCSgNc1DD7DhGSazWMPMNGqDE2xVlqoZgEgCImjoQELjLqRs40TUhtDLKJvB6iglvCCg/2d
nkw9201M8LG28zBVg+vqQvnF2HxJ0Yyt2V6FmVh80u6THRuWN1oTH9ZWq+Sg3USUDBhrps9uM1tD
IrOJiN46Z7JIMgZF2fXwnUpdg6Es/SjXad5Hij5nP4Klc3KQQU8ZwAN4v7inSsEhfikc75xFBHBC
aZyjEnCsqZdnDHUPRlJyZiJh+fjVAlPXgMcyktynF7awVKqqhXC8Fk6nCWWQsCHj8CATSbMuHZRs
qIDOsqz24iTS3hSnNAiH9LhE2CUHTO7VmPIVwmb2ofH5vGZY4fnrgB3zCClMVOGCkhzsRj/yePCe
nM0fC7rd99dVusBPcFCfmlbZUjtZNW/SeotVEyxUi58in0eyg7J2C9WbiiTB51NMAfxE/vsF12Yz
ONldBGpeS1vvHIYv3l+zf9VhadOQ18Rre+gCB8cOS9POQojOYEn+bzNv/bA1KCh7lBFEg7XnyP/G
m3JTAdtK/tsSDY0llsKVlr0ugErks8XfesFGotefJupZIkzMRVzUHw/PcXTFXb8Q4hvlFyctSJ8v
c+B8OxEriaryBmvaWqilJZk/r9uurZtB3I7Fh8UepsSJhUFStZXOlgvIAd0Snx0TZ4GzBrqU466y
yZLmlvegYlkpK4PmrEWQogoLOqnw2y7PrRH5hYTDsVCudpCgZciNmuG3HGv2R5JxFMqpvRO9dccA
B1YJJHI/h2Bnv4SCdhBqLFOKRt95xdNk6nvPHCGhN5VlInnVfvGTmsDxQSVWxyCOAkWRHuKqFrdi
flYM4LKqARMtjL2ybS5SfmDRgJaKinsT8v1Zl+/4nePC77p7qKMe7vzK6pSjilfbvELkNiSt3Ed0
Xj8/GMkF5K67uKi7Ta2UmouOTUsc7W1ahhtPc6LMnKzBFUMQjGTPjp/VQBzRb5tr8TqzOqqiZ1jl
QiX2j8+7mK5k64wrGGMRumr8IJyHRvd2GT/7xUCqDfgzSdrR4Ejx47AaGdTsMbJcuZVtvO+Vgp3u
N6LcPyvf8RnPAHkvw3HrSjJspZqy7ziyOjm1CknQ5W+NYfgcF1+QHxE42u0RJ3GNU6uCWKVNyAd5
D0zzZbFbQtF98EBA2yoK6jgm725zvHk2Y3q9ZSaQg8MtFVozOkvHj/8+3P9F5u7CoNr5ZyH8D1d1
Cz9oJuvlCvHdbKgakpTZUP2T4AMShfvYrD1cYcw60MG0qduXnFYsmYSqxpeNJFkow3f1oUJRcAZB
FaO2oLQoBsn7PDh0PHF2Uotz4Y0vbDm/4WucFt+XjO6B2RgxeVXyov5pTrRyDfUoVk5977WW1AoL
iUxdQL30wEHO7hBxWTG2lXi/5HQoFw2bCHgnU5fZCC+fufsEPVjMdqxyiwN2VfBuILDLbN8oC/bS
isuApWKw/OFElgteCNcvqpj/VaEgFDMcONGOv5Nj3Dxapd2VAm1chG6eepioMqMYP6kqprSC9n3Q
d78IV+7gQaQYAoPmi5de1iTSikluQ07lWlLRwGlMsv0eCVoNhQopwgcm9mmExm8KwDDx3MrrsBL5
M8URyJa8/IklP8o3zV03s5TMQP1izyFJSn7BCXyeYN+EDADGe8GlMmJxCmXngQTqVYcxsoqhCenz
JJzT7BI03kcXxg9TYKhmb9OiSZzGR8BPtLra7gme0XqwqsCXbabwAOHraKDDn1roAkvWWY8k70EH
1/1XpuTh9HNSe+HK3NlaAIr9lFG4FvYwSfaqIlFZP9Op0f8ml1Oev4a6w3A0B8MFCvju0r+aunEc
IBT+1Tn5kAV1JEPKbZR+UZo3ajHfL7OilOmJzS1RfcReEw6/xP1C0G+0ssq6jXsr96G1KpEO0f8s
5t13AaLs9erGCcB1HbVvFWMpRbMOqiEvbl3Cu7ND672oURzZ3YZ8kqZm6iYWsnuVnPsk1vJ+O/Bh
3XEb6l0wm0ajyEa7QWjIH7VEIiXw+gkv9jgiByxgBt31aVbvNW70hZCbCCdSXVG7q9d9jZuNCEAk
+t8rAAyy7XRlUv/FzBqimTe9Sw1cEzYEH8SrrG+DK2RyPwiesOrNm8b7/4lle2fbxud+yJSTpB+y
6ng0ZRG/AJp5NO5my2ArmYZR7JAaU5G8plJ+4eaD27sEBC/41NNYC4YQNtV/Sb2zkHAZjZ36euMA
eZqumrziXJypudbxcbxFEgTn175Bi4DsG9pvGOXCjSxLDZCSUAeLQlgM+BTi7b8Vc0TDckTBQM7w
neGSW4v4k6HSRIlNOYYpT/qwy8TbfVQTShxDDzgAP2oqRWvDTFH045a7xC/NdhrJeH6rhP2H65SY
Oh6CiMFGs/Ku+wz29W0uruVCxeSGyuRpm3+hsTUZvqTl8hwMK1KbrkJ8zpacJMOjXHmTkc/QDpke
48sWmqhP3JdeZ3stp3DvlwmawqmmiUwkIcCES1cjeB6WE9v4+9tfOM0NuFDLE/3yAfCrQyagdWIT
Avyu/EHJcUIxyD8hkrCqOrYli5vTG2052xVVfGCXOgDEyBsHLPVgOUeK9WuZXP8cbB/WDcBF81eT
Mie+0v6m3852RB6mVoUDBz9FBfRs1JKPYi1cZ801i2OT6WICJ6fWKkQzZ04G4WPvb+OFk9ekkhiH
M6hu/NliwlDX0V+lSaoRrNFEwSxHsliAqAdVsp57Y+/hSYn8+fMYwhh8mnXiXlQU1B8G7ewzznGx
kjlzaZR6rYEFz+VrPhES9JD0eBdMOwYGDYzmiilESS0CIDPoNlKzi/2GUmgIwyZJwoN3bc83O3QR
DNLfcjyoHiGq5gpD29jO+HaKGDgFnebiN7p11wu7ek48C47s9jD4DtDKI9CzdTWu4ha2gVqr5EGP
IbrkzTmcVq+DHxw8aKpmk36Cj/Dk1bm4IJtIu3B1BV/MK1PlOP+PeD6IiIH0Rq3HAggLR6xEM/Vm
mf43hdlZQmLuBP1jVEeRFFDoRrZ6tdS91yGVF08dtrlHm8Y/okBv4ee73/0iKpnbUuxoTm3NE4yD
EF7c0dMXahVviT/lyR86k8MuGU0H2drbsaKGiA09XlbcaGoB8XqkiCxAnGPu7sv8+ykFX2uNmbzi
rmjwNd9oP5dmLS+r0EELHxM4z9dQ1p3F+I/KusalBgRcW3ze/ExlbDYtAK2VgOiaoY8Vvv8yY8AG
k02L8haRKseoQjCHl/NOsAakhst1rHVpT1B7Npixa5q45JxlUg4FADuiRE6Y22auPb1swetaGGLD
usima3Bxi4DFtUg1oCxWW92zYXiaIWrwazF8YTlo+ZFSt0YNfv4yFIqtN0ya1Mm7XLijMeOEATQm
4fCLNETL6xRcIO4c/US4EVsELoXKIdAo4FZuAWShS8R5vWPug022bFg0HbWAzB+/t7Cahj1ARzhX
jNzdmiL08bcHqM+wt7nKxQATMRGU4vETZ1ZRF/vhPhI8Qh5V1Xh8pLRMyeFABFMpJHySXaiTLLsI
Zl5KFtF3L2KfIJoeF1MLCmHjyFieMXqpdQ+9oFH3uun724yOTFdl9HPrDfXB5uG+AWZGKf3T0QaX
O/wlXd6ZMImjtnMt+rNw4FdXescHsPsad2lU8/3JUbECs2ZLDvla05UOrmsUYrybPZ14X/fvZZCD
F818Z8XlYgPZ9gOf1jTZSlAG03X/xBFmXciv0bi+vQpwd+gkWcn6UgxYrlJ+gUOGzJolAdgVdU5L
+SfIR8ftXnaRoQMG9sfASKSQUKY3MBQDABsogy9yqWUUG6UJIaD/bAmlHtsQnkHuvliTg+ICUTk/
PtMio+UZzUcyHoRV7Ibw//TMpOePLqSoCXVd4cO631Jl90V0Z9IGjLODzXTxVOTK5Ob1KiEbb4ie
BOIpRiBolOmAcn4wTJNSTJGeFbGfW/oSRvfx3bO+fY+NdFXSct3gDWcn29sNvvBx1Rpeoy28d+sH
tv1AGtQWdAkWgnCo7v3lbKyy92/8XzN4ItF+No2tIlVQcfWlJknA7HfFVjdxXgPoWwrp6vUD2gdY
RA5Dtth17DdPgBpnbqmInBoJx3CX3GqdyCTFVh/+VV3sHwmJNoEkSYUF6VYuVaZf0KFZfVXA7jkD
taIBw9a+CLJUrJEbFU6eU/YxwdnOWll5Bw8VtkdH3hRQDLXxtJcGrPEuGfOCCSnpIioIy2tZSpOf
A8whIPArDBQcsYF/E9WLXUNOJdOzNpxNnNSWqWn3xNc+Q3ccEM4UwEvqswhLFRZtagyyybazL5tB
DDFf1Yy6F2cZnbGCwovskPBUQsd10xPf+8eHX5q7gDqAt1cHUJMBc54SyV0nZHYC4FU9fNwtnz/j
FvnH07bxOoyB2equ9+ZhiPcRSYW+gntSZwiIiM1PTBBD9c9ALbr47KDRC2dxH7YEO+AR9BsaxqG+
FU0gsqPYDexohoyDqwjMGjBR7f2HBtOBnscFMYxqFS53hSqERDLdTUKu9U8C2I39dTQrE2Pr+A7K
uQurUToZPOPPvTJTFlgPy3ajxLsClq1bIWLaKJ7bRW0/2686BriiAUieGN/gZtC0EFeYag1OgMDJ
/LoOeWtm6cO7mNG42WzCq+VOEXemZ5T5DoGURajYoYxP8fwdBmnY21UPM747B2roODjU46tkk+ED
Of5JssUw3COUkT2IwkQTqgHq1jKv3lnBigPsDNSyBZ0i/JqB5EzT78DnSHbVa+493gJTcQRCIsMG
1EXDhUFmwWpPmF5Xdk+diogeTq2wotJVDJ+EHLOU8u2FiLJJqWNzPHaA+qD13wVraxAxVeg0lvYJ
IXqU3LIhoa/geWUMglzZCEEX4oHMixC3T66TIVm114lwTR2uoHogLZcNf5qFE42SbczfJZOtVXJB
K1LC7WZDBWZQs5Qi4EKvBxYssLytJSGSWXzAlURMCDpISUhcPQGHbhNox/ULH76n+TXj0NauOZbR
nMifWmnq26m5c2agUR76LxLR0YCpHXsmpnKcDEW6SGBkbhReirGoCj2odhqEOlyq9z9Buztb4kWr
dQjwEhd2JywQMCobuRYTJ5EO3UN5szOLTy1BRLZUl5wYwwMKLbRWVI4YviQkX9cLt6hKZxcpQmuF
qEBROq3UUpKSUNEtlSLoIY3TThqf9PsW93PM8kaKaLpfLk4RULPkALCPr9B64Sj35sNne+n5vPu+
/Br6HS3uqChQKduWh97bs+7pcMv9YywyFhupR/Yu0XmJLAap7n3UrHz24enaBZ8lFAkSw68ex/Vc
cQ71nYZiUaCPRuH50YLAZUh8jjFCvDykK/8ZWLlP9Zqx54iR13Mu186rT9UhC2zfqrIEqXSyKVTd
zDCOz7BrHVYV26WtempqSuE45Vi84Uz+e6dLc/UPkoKh1ApRDvQ+YYW9hSbkwHNxmTnTjU8f8ILO
6EtHYkKEfqAqYPo6CVZ2LeCE0w/2RZBpA4ZOvsCk/RYRTa+YGihR6DDN1yklsiM4ReYej9c8LIyK
cai+lmlpVnfgyf5KeAJD8iKKEuk1A0oi3B/m1hO4I7mrCEwUXyk8RQAHQzSE1Qz8bXCSqsAe9D94
wAPEm0nzqZOjGPu7EXp/l3i0N08d5/dIGcZQzHl2EKpxShex4F1mXWsVyDZ4ubWLrbqjIDECSXDQ
g3EDIdIpdqi0P9txjC+BPwMMDQWBn3kPHgvh3G2mq/iDVEPIBbpdiR5e93rgupP6qUNFeH+IQAM1
2loYpBl0vbLTzakiyTwwjUfpIA0L5hUlcsgJybboSj4lC4mqs+gYanmDiDpKfidLS+8EScTnTNVa
qcwqCfhlQ+ZRRy4c2tiqSJ66LCgFy6/xQ4XFGQXHzZ6yjTnVgHWe6dWFlFnBj8pWt5sedSZ7MqnZ
j/xfml+NaeqCqzUj3VJGySGdvkZCv+swUz7KICWYDu1tS2pahS+ZirOp+A9mc4PcJkd4TpIkFcq/
SPIk76GICdwa1DiIN+jsEnKQ3y1uq/JNRvyJ5eG5LzCyXKCiBqCIdEYILAeGWvAvLgmVpGuTaG/2
LNvr8fV4N+YSF9lzFIiqp+lt21Iu8HV3pnNHDDcEjDzBHPh+eYKTv2cWLJwfR1rQhutxppNYPgCb
xGmM5P0VABNscHhrIqInWivBIehQWBxFJ2aB3qu4oyVPclr5/Di675UJDsoHCwCdXbshY8AwA0q2
vo3XzdMMN9QObPaIJCXyy91duat0u9InRhgRsbg9uUwahJEtTwY4snL8Wowj50TSolH6+xPo01E+
LCJNIXUP753mVuInkoriju/kFtt9GQLoJyP0VoMzbxyQJNYkRVyloP20AJsv3VZ3t1zBkA4XGr5N
W4p4+KemnwiM0Li0GB2DDN+iKBXolIuQgM5BHxPThpeX9R9ib6BijoAh0fN2Fpj6ZpJZ9XVaPvhs
FoavvEzABf73CQWxVrxGjkqx0HiryuaaPv24rwz8ULU8XYPQqHF/XatDiqZSyth8lwUtZLrzm0Fw
txQUM9cX2ZmeJk417tYcoSLNG1w19JzbQ0lOsPlvf18dbajBarf5FpksesmyjcwsiYlR8hCG+Olq
2p5j9H4qJSnDhh0DdHjV6apClFUleP5Dzh8xg/C4sySXesMdiBgoQMuxdLxFfNeorMUsi3BhrywI
33StenJjNGyZWq+InT12rnVoBO7UzlyPfTjbwUxFzc48CQdUnHz3QnBOST9UkMUZ8UkJ7FwWMLt9
DYRtGIChm9/3BgKIxJuTJGCxWQJ6Yj36WSF9Cz9CxB4gNXUzSxAniajvRXA8H28wBfPezy8lU/5R
pqDPAFUwZyjQI7t7Bve2W5FrnwVxFL52z20muadjRHzVo+jRFS4pPawwnAeDb1QleqJLv2Ev6HEj
pjWVrNz76Y/Le6Lg8jim84Z6xZJnBVAKjOx1IqHnFt2w7K7WdG9RD4DOPP3LYS2/wDPpziYIaEMe
pQupfIHuRNwzcK+Ri+4jyfojkk5JOy11YdsaAtjrDCRUfIuAi+ZED5yS/mxgIDpG2of13LvsnCXV
NXjygAJqdWCekziNXaPWyQfsAPuaBP4zCYj/BRGVervudoBPzEastdh1QPLioIpI2cwru8QA/xiu
4qVyEFQbRDQgwfeJ9aPxAjFTd96NlfdwgOwXY4wNKKjdvViWxZMH/ssYw0zC+eMpCYVBEclophqd
XfmfQ/Ug9517b2YlmTDjD1RqPcgQjcdp8Bp6/guSvmeKa3EaYIsH6WJcCJ7saJdPHvGXczy2odB7
pwUnjbv0ubMooMfRz/ZFxB20CXHm61Lxlbnu09sO4I6IRD4k2F8diYmEdkI7sGdhvCeQPuzUa6jo
C2Xuiuxj+dbwShT48EZgI5pjuXLpWYZRX6lv7rZJkn/gb39xRHQcaFAzHZZdiX7Z7CVClDE5GUdZ
PEyKcYGVDXK+L4kUhYeQqkjYIjyk9Vp0z13D7Y+SJR+MNp5jEBl10yMva8q7zxZZtR+peZh0Uyjw
zVHD/G6nZ8DW1NueqJmRrs/HHPygqo2ClvnEbYp+Oq0499657/o3oGTDkhXS81wAGW80nHp/wdWX
nqTSwAXQsWhTPAUG4xnri12//VTkGqwCRsGWDi5zlSGvawc2m97+w/Xhvy3p/2fTAENoZ7qY1ySd
l/uRwbiQ0xMqG96W8TJ216NOs1WalN7yTzMpq8AHiU5BwTWMB1+YVq/1ozNERq0Ic+ChO9Z+tgEX
oQxOmfzgxS0Or+jGZKtA7snrE9CRrEb9RmMcoghruTZAnBOAcydNOis1i7JGoT9E16BYLZJd2moP
DTno8V4SDiZZbIDs/n1F1kdRtsbSoH77xTRsCjiUVsnm6b2DPx2kWen7N6XeE0C5WbkFVZNLF983
yAlz++Daa/io1PjV1s+pwBMNJLkQ4qH+xn8aAqLr4WmitOs3QTk85yNV7OzB7QaSDeT9MIiflei7
yJf/GaCGBycDiuDPeHd5TeWF8gc2DaUnM8kev00Gf7hkUKWCJnYRAO2V1vQf1kk+UAMbaYPzL3mO
nMiAn4GwTj+NgzVtPLszv9gFjKXmJE4S/buz2soyg/wu/8q5QB6AOZNEqTTORur/vGkHzSLhbbHQ
79uY49CN1gkH+gEX1Op82j4qgMEOGLTVNpxlaaf1l0btMNWtmH4kts/z92SutAuqrLTT73PH0sYB
dUvoAzc3fY7maqHFHm3+32R5LsvDPXW88GOx1FbxfRw4/mQ/u/XyFHknCWGZn2DgdUGDFuqnnqpu
c/UPK/y64ov8yAfZtPxqawFjYEMzBRHuAtOEeJ3DuS8SyddTfcZZlpxsneH7F+KXqQR5XYRyUThM
T1O0YpQjiqn/eyiBMnAYl23o5B+JlNkjkLswXTrqcGKZMAyqoo7HVsZpmwthD1Oo1OFm3b/X3CZu
5xow7pGYysTW/UdorxeOSelU4/n7Tx749ICDXrYQUXvQCf94Hgn1T8O41solHPVRq3Kyahz4Ip9v
v6y58Vghkf1ph2/AK0McUh5g8qU55KA5FEGRswtqRDYmE69PorGZvIg6y+DLZ7XIZRgsYK3fbVdl
NDp7MuR7aWfx2J6SKZ4akrNajsycPWvKVarNd/6n3SxrDHZbVX/rIGKzrZtyAlbYUw1hEgj8wRHR
W/ZCsb0CYvoTBui3ySzMev+EaG8w0UUx6y2cF8h3HSdbYhWXMRHz90aRNoItlHKWTBFhyUe5Cffz
xbglFFd1/il9QGwZxPzqlza0pbupeNvSckhodu/Z7V6jIMYbbWugPVBiTCk1poXKExfUUGExoqsN
LlTyG2iFrSRuLpJKoi7ADb6veV5AQGSTrzsezyUU0AChBQ3sUn+D/TIxdrLyjJTLNcJhzyE/X/Rl
Bibxh8RKed63QZAyiNjOArkQdIg2aOEz81f/JnS3SOXMk28hx3a9MzdR5qFCOtwbm6XMpSY0kaf4
xM+1ZUYRdvHel190B6hKSXmOBiWB3WSz3uoq5bqaI3cb9KGb65XT4+QkoghSYk6X/H2soU3qVX2G
224n+DilfcAXU6R6z1Co4Fj/x8rQFOG9yXiPeGQVAQFzW7JTOyfo1OTGQYtS1ixDrpAsKKN6yR7f
l5+HcerGhcRBssnaXBkHkMdHeDdJJEcNEm8g7pbyOtL2sfmK8EYlsSekpPOW/N/vsyt100kFIQ9J
KaJBOkus4nq1alooZ/uB6zEYLLFMmOGNYJuKAx9+OmffLG8mmO3ZApM4Zt19ErS5p8tJp4ziUCFQ
RMcN7UdYTwkCqWwaFAebx3WTJtzyeYjnJyu4JcMP0IBJGMotE2AfYV7E5EzYfZ3h38132yK5w19M
bgASGCu5O49rTl1B58eaIftha0FWlFPZHbDYwzfphcieOxmt1SR6BnF8eYcI765PZ0SetNv/miSR
5TCUJv/K2hTmpKy50fCI8Mos64M+JOglzCvedLAo6LCeaemnhotu801nnVUGJ3gg9VNYEiaeDwKs
KlGNcQMOjWECYzkbJR3uqcVHzHGxJxOtzI3jToWd3FdYH22V7eEuMVo2QcK0IAQoLJ/Rw/UcBhUo
Xwhe1AsQtFBoE5lYvawLN4kyxNykS1VsYEI1BTMkaXdUORMDxsOQRgjg1GudOEy8IuAgLeV5S/T1
4M4F0W/OngU8r+QcTdL2H8ifxl7Gu23H5txUogoUmy5UDhoVqmOiWWlhP8MHY4dsLXlMKObRohIn
zke056E2FM7wh/p8CZSzrnQscWR8gTEHxnaOm2n/7e9e2DB5HD8VlpegLGsxNtHfzMCQXfAvmkxm
Fg6owSiliS2q6PaKW8yhE687p/yRkxw1R68LujCuD2Fi+DrklkHWlAxunzAXJP6OO1aOijc5rtA8
fx0dn9QpastJdx8v6gS+OqfQec1YUWo2v5qYi4tA8jR5nwi6azjaNImoq3qku0Q8LPaSMVsBfaiL
Nlbtp2gF1VJOWMTanTEDnsqWKYRvdghuEXG9BKbdmS7NDNkRzQ+jFcMjmdSWrx108I9GWn6P+0ht
cVhlLgxozceosaz5A/SeLUt0Xsv0qcG+e5LNv0FNjLUuc11/zIkwlf8CfTuk1v3DhKp9zPKRVdoQ
B80DOCXv162wdB1o7i25hanh6oC4HB0S7okYbBuoGL+zFjmg8mgWhO68MJwvryDLaY3V9aTyTFV9
W+gfqd0ul2FmPBoMRFiUFEsWkmBv7/f5eygcFSn/rEzY4KjKJ1Ekf8ISewcdupRJXaws63U4dC4q
i3+bty5jiypcebP0mqoGtofmXe+K9jzg6468qiSh3cH/SfNHnzRjyRvs8ZZxZtB8QfJFGaqQb9L3
g30HU/V9EFqIvC9672Vb8dv1glI+4a7BH6Hqbjl4EpWojXglSmk9pRCLaPGuaTLUtWT4Yz1SiO96
0GISwUkKlEJsrsiWoiico3CwW3yx6m6qN15s0TZosQFbUCKNEUA1GaYv4u17OqHjWc32B0SKaJyt
qyVA1Wyrtjr7OiZwSunX1uqpnZ2WLKAwOc3G9Ki8vuqnYtK9I4Rr0Mlzds9iecK4W1c7m+i6ph/6
R2nBZJe8AqMcPv3yU7FTBp2RU4+8bE5RctHd/R4Ft8rTofUSN/IHp+q+S9XTycrfK9PzmFA2LYvO
Xb5r1hP/+sXXgfcjU1WtR0eT/OjYdfSMSrb353scA4I7OVYynIaebutGp7bBqc9ce7M37uVM1EIw
7iaZbgx1JjSYN7NuQUH+FVkkS0wsiTa+KlarU5KVMQE9nX7e6HZy+qPC1Km3Vs8yOfERsWAoFJvO
WHDCDRV/sZrYJNNIvCEQ6GpY5ziC/0/CYBhXADCy0y3WjjRvzV1aS25fCzcyYLmOUOPArQDnwngv
XjYsWJUZcUQsF2qEJ1YJ1/I2pKosFipxKncydQ9jEROhPbMgEKlqTOrbb85Do55XrrZwY4qUEP9I
DHJETmG0z1aVbWqqkfa4tsuoCzAyZt2Rmv/z9D8+22/wU1i/sKU1p+g6o+LzhsHoy+yEVH4jmuiw
JGNI19G1QjsstMhhv3Jm2gQm/UALzWP//51qn27X+gZaVVnaOe4bmYNO4bMwQuOkgMihojwPD23r
un5ShlIVBdzE65yVAF2uFviqbOa0zlqzDrGoNTN1A/RcKpHlLNWpnQjGlrfyXyPD82sq+B9n21+2
yJtgYa+XthJL9Lc6Ic2WMTMwCzSjf+7etETPE5Y5rH0KWzHR9JYkpX1fPOUTD+6k3d6ic2oiZnFl
7h5qCHrKrdgGJoxgw7y6wjdDg15jYaTd2iSrQnjBdk86w2nifN2EZfySBRA5aNSM/2a34Or8FHhQ
Lnv4DFHCPdWz9sOElHOaH+LzIdV0RgPF8ZrAZM8jj1PEQBmYpQpKwgnV6AsG85a70rhZP19zdQgr
9EubuhrWJSOKdjlmbGjuntxHzcbLVQn/e/lnyx54qQ9SYCwMtUU8oSm6s91Cbvwq7VH1hYbaYQdg
KCEquxpcs6g/7MngI6atfWgv8cPoskmtphBwG8mYogW2N6e7qhoFnbb6sU3F8xTZe/PWdDyNb75g
iCR9c7FQQEoAP6M4zECKQICbdKVSiwvHYZn7so9q0fbB+9k3NT4RxsFCjpsb7pcGTr2vWJZ2bTNL
MKwXSrh2t7koaBhRl7/YWip7Zhp83q8IAytOml1jyGYf0oGufSeZILQx0IePPRmPO64Vv8/fvpja
7kN/K8USNGOl9/yKso7Eg3AArzopNCE1lbYDDEvuU3VgbV8cNIXqB7qu5LgYGlah0w3oQH0TCT+S
Uk3boGrCiVZ6CnEpQ3Wv+RUCMqyCz1bEL4RUdDoyfIE5UauqFQNkzQeahphgF/4Y8IN8SF9alvl2
Bvk5irrq8CgU2DZYTZw+qFLPZ1lCucAal2t4I6hl7jMAS6ssPBGZdzgnq/zc96nj7byKv12hoTPX
hSiGgNq4yqN5Jm/ykhKHhfzlrg4g1kw+zmBr+MNdUvLfMe+441+0+cinK6kDU/g8zItQX8rPKhDc
267JCuX5kNHjVuw9WplsZ4qNZ1XoRfizcfAcX8N8TR/NotG9vfTJSPWF5DLFm22+QVhFZ1rgZmhQ
xJN4rLUL5T+s9EDjf7OwWUIOPUZpIieKJum4k8549WtOR7finxEw4yCAg69VK7ceQarW5Dxj885H
DKNXMvL/PbcyAxYXOltzKj7+jFunG7BkelWl2OtZPqnmIcZ+uErNao2jtnqB9BHCFfrd1UgKRUal
EcohAE6DOlSTwHxEzLzfDNBb+mLOnIXYWmjz822tCbLrgsStizO0M3nLRVwmEgWKscgwQVB13EdJ
kPqEH7RbGhKRr3AL7DZDE1fjaHENpAXHZxw0anxPnrl6Jd2at6g33iMatO5v9zKp1BNg5aehqF3u
hW3E7HxbG3YtWwayqr3J7NUB/IVubo8jGMcM6dUxVPupBm+gMyEx6sp6041M/B2Rys1lY2/RaLkL
FJP9JEaznO0adUci5VWMTWsqbKNsaPkE3lzwraZP++yGuI4B0RFqc7xM5S89BMqM5CkamoOknH8g
4LLHEZKynOiHQlrmp3L6+NiLkocXoYlkL2CVIxLfj+n0XAiKTX4JUadCPxTro4/TbaSDcbXyVWTz
SRM3jjvIinzkWoYkNSjwxz9BKkPlBub/SS0xSc7PWROWRbKytfYlzdn7hmk4zfXckmgAK/48H+Um
Hhb7hh23jw5IoiRvK30lK8NCnX3CESCEskgyr80ezPBYXVA6RLmT/vshROwb0ryt5BdvxERPeTnh
5Bz8EvrM415HsO7KejyVeByIMOQ5/RvB5+kXipe8JFVoeLtzZx7kujqQHW7SGn7l3oAG1Dwo85zY
2w+bpuPbxkNOFE+gTZzsR8ivp1WSuombhkZlfJxRjcF++9hFp/q+wwND4Plon+Zcntc5WL0Jxi86
eXJKDRnYxnu28Zu9HIH0ptTqRgapTvAwmY9TwK1aGcSPzTPWXV/KmPt7gsQuTFsVi4pUQUtaj5/G
ZiA5BKQSXYBcP4T4WTymjtpr6WyvDLfJdkC/euc9oPVIbY+zBbx9kO9yjewQIfJpCLd8rU1KXBeX
4gg+s9ArFmofmmIqljKcaITAxmja/kTv9n5XDeCog2O+v17FdO90SIY8XKVJnus7mMOf2PTLtvX/
/3HxKK60T9DAxvtzgR374W6B3xqMguHiDDwhvBu+25In/pt5CWq8BckZIAKcTCx90cmpsXzqD5GD
AwO6iSBjQNMNFHBudX8teJ6pz9i4x7e83vz1Hw0HFpq95qUDqH2QYg9ETGjLrEeeIDfKF7l/5X1P
dN/k6jqWySH96MGLB9BT0ejXCfPB189hw57LyuuBiUaW9JfWtf/+KeoX143QOGwIyxwiUEJeZSeo
gvdLWQ/kDFRzW4TQlq7WjXSPLZ8CD7IEeuxr7iln/uCu9RcQuu1Fzadl/0bavw6r4cwgNwjDp+JG
Wj/yjP/wox9Rv1kpKsG7+zeJ6gt4G9FeQVwwpjN5ng9aiMcNMXuWLmNCoyQK9Vja0TXkXWP7yYF6
Xh9ZcG6gCWwUw9Rid3ntlnIPNaz2exjQSnKrPmqNJWCeNSIcEbQIBHa8cIlVzjNPCho+gqWdDbI0
y6TEqEqYH7CEvjTQa7UZMU/XnWV+vfL3MC8JpxETO/ywSVI+nj/jDsZlo3RZyBbo8Z5DIIqhqM44
aq4hn0tHr9oJ4N5FpLU3C8tOWuQ/eP+Aec8PmeBRSAQ23MXIDD0eHWvmLEJO832KeIqsb8Kyq7hs
GUeWe+aRVF8YZcJe9HwZvfE+oJdPvh5Od72mEzt3VzFLZOBBGoXb+FONI1iP6TheSF1dmJRlJ+wT
l6s++CAL16a0xcXFSOS9g9DfaT9+1OS84Yksnbf+qR42C9YKPcVJUk2mbVGaP3uz6iaHdcagMIPg
VkbysN17e1710o7HkRsa0ZjZ2HApHlANcgKwutRlqpmN5AgLHhqdfRCe6FcASlUEribo44LZcinM
FMq7IpugrhIlPJO1tDaUmPFmM+X9GMThoad96u+GRMvnhXphMOdp0Gf/meQ1foN7laxxlAjOtlAL
9spEruA2mCCoufa5dBz7E27TTyWtFM4BlcYoQFUAbJpEWlPOAB4qezatPjZ5uUCayYn5mkaziOQW
tqcrwP2HnShsj+a+IfO0Hsxe+wQ2hMw7SoX/lkgUr+jTaIAtiz2bSS3YvrVGG+EXFfRz+5TYa2l8
wZNaAwwncqjWMIc80RD4jIOpKCZYl2ACEDBaVZCbJn5I7yZBI7V0HHZWFqWH6WcvehtAP22fP4Ye
VDXzYJbrh8pYIEtmZHaqM+h8HhjrB3fgYYVA6gDHNJKBJ7DRoI6gwxSG7P/ehNaJNluYV6lfP/ul
bC9wIBP7+5fSvcSjkMy8HLqen3pBH3YKFW9OxqJ5e9ei8Q9/2Lt7Mh8+gCpJlQeRPJOYBStBsi0k
K/V2NnBVS9bqu6q+O1i4yyTJ/VRrWWohpG7VBrocOomUGIDKp0eS48k6AJN6P0xBxBwu4+uHj6nA
3ok3a4DnIfDn2b/AabjYm9mvrDy+N6ctrxtyWRSP0vJyYkPJDDEWTJlflbul+iaMnmhDq5EpsYQ8
gE+P09SknPSqsYMJ5HZRg9Q3W3RsH4BDwTw+/h3BlQ2f1ski7JLDK9AwMTF2Y6CQDsJ4GeNiibV2
vYijxO6GonIJOmT+pJ5748du2Ne3iGXF83wA9tncDSpbsXpzqhZpYpH251ZKs7rghg1y+MoEN1LO
WHXipfHtlqs26n1nX0EiBKbL8TwZGDMy4mJzuw2Gnb8DmQh5sj+JOOHJp35WCw/6jEWhhJh9bJ6q
wjTXx6Mdf4Xz6RTaN79tDYA+PNIvclV7+oEAUOd7kkuASCt8yQW9QOrMgQF4NRWoCT2JAw5/5nfl
J4SDGkVyvWgqUyr0PNlQn3ydcRL/UgTDoW1AESHnqYbuvHorHofpeJgbQodFtaXSok0KzLMJ46Sx
+cMezR1rIW+QzCmz9oajHb3ejmpYJEY68lx7gyfyys4E5cdsGBBCcnDNpvzvcKhcXvP9JYwiSq0H
DhsBhXb5KAgQ/zMx1N0TEly5HuPEICp2DvwEgaM2r6BddnK0GkTxvpm9cfed2akvRx5jD0rdLGS7
tRL9cutlnAl2F3+HkFewtoRq1DPnWOki1gN8FWf7PaK0ZZfeaICYq1amKnVS9/QJT7lvtbsyji+A
qvPM417a6c8jzFla7R78kj5IL9hINEin/uVi8t80ww/Zvo6ER0+hXgxtMti7Tw8u3/mhrN45WIWT
kVYCW1Qz8itYXvveLL+xBW4VPhsJsVSBdr8rBXhMYwQTiz8eCv+XKXZjLu7S3CVxK3kW7LU3OcNL
DO7lojVwU6PekM0e2SqIN9O/h2iYIjbv/wT27TvkpaFxrBKEl5j4vvmrysRZ3V5Edg5d15e1c+w3
URIeysks47CpGJgGZfO4Y4Xnb7vZjM07NQry02XzoH4qRoZXy97r5dIt8klEJNwgHt2nqXqGeh++
wmlLxwJmRXPKSnZ851qK7RO6Vw+e/DMef7JVKnfBliDgwByNUjJci6JJPyccRu6ngqOkYzALZdOC
5eNU8YBhoyAlg3NhlpLawqu18pZt+PmFgpai/J/UUB1hpn1hR2SWk3JdL3Sb6RTnvk8krZNhz5MI
ZuMtPL45KIur/B1bcjnMsz+nXjMhYah+ZAoqhI2z/Sf/uN0TAVbRj4Zd1JM9jxivnT6+x26Vz32j
OGmwdDn5GUlmjtS6kkpzZTWT8+6nWRr3kJcqKp8JQmBwxQZCnsN/K62GAvjM2LElQdzja5zcN9If
UF6yeF774YUV8j+q7g114qRNOLmxCxiiIyYiA32n4uEPh0oxPAyt8cDeDk1i2NwEejW4zBLhO1I6
pjw7j8SsN0T+qrkzIV3Nt+hif+yZ7m8vRROp3IjLkiuWHZzNXP8XT7NL5TYP9WQvDglg9LJHEB4Y
WGiri+j8fOW9C9QA8OtKP8e8qYd8y3Wnp4wUZjYy8EWZNoO2Z001PKwfKC3Ou+aEShJgsZwdbdY2
PvfafWNySjLQhN9mAr/hcn/ysVwr0rvDlE/zzCV29Twr4VpQrqznLPiB+Ogzkhe0JB/N7K48WATO
bAu2ulv1AUl0ypi1NsTfV33vDGjrCrjvd6t45qaJMyUD2Mkmjn9JNkm7iCLOzMQ0g04jQ1b/6ups
jGOuxaSE2UEwkJy9MNJaexNynmmH6bk8+BsjeahfixXs1zoCN19HSl8YRdZ+rzKQLYT3t3Q6UoUz
+lOTemFK7917q8Bp9Z/hJqTI1FWYTKljLl3VZ3Frwf7A3YN/2oYUooS9we/y+uU/1J8CC9RG+tAW
BOl0N6dZXq5yRriN3q9GdZBV+NjEOPEjSaVZdZgc/mmuBYouDvxDKgGSGLk7XcTxDHasUn1FlvTk
R1l+fVnWS+tS4ou/YRPv/kXoVhUiLmVmOPrhGzncGeAUxIl4QiRKkzmlEXWOyspF+mQxDr3Ghgka
wGEqJZx10lI+22Y0creSwVMwl3h49IaU6GitoKCa5NRUQGGnXwxCuZBrhzTLsMQ0HrvxIDFkSf6+
jbhtizU65ztMwOotptV7jewyyrpeIcyTXb8rDWywGTmACJn5hGk26uDygm2sQIIs/hrQYmWTvE0B
BoQl+JFiOjTraBOH7IxHBiaE5BLDPcery5g4sepSvmFF4MHvNnPBrLt2+NfNFuI8c3Xed+5mzoT4
Cc/mDhGrw5Khsx15RJD86UGOY57izsg5dqWusTsoTjPOHKfOhThN4IBeA4NzbMsU1EDqXbfD0wCY
Vhi3BergqncCoY3HbZwdac5wcj5k3S/+bS7bglOCum58d3sQH7QK1MfmoMvjk+/QxeCKF3Y3I4Cu
hSaaJZaxTL9EaW0HUW/YN8ILPqXLy5kkMMU44T7PS1/x7OHhctSAUtbuO50Fw80O2KMsgSvErhmO
Y4pywQ/sJBjAjZBxrYFxqp0/z9sYKjxyCBCu3OWAeg9YmOF7aW/N0inzOwXOZoeB14nsthSBQYIF
oGKcW4R0xuRv1QmLUTAR6fy1QzAkBafi/fk9xFPY7tqczatYn5TaV76MUUHn3yD6Kv44W+H94Z2D
xyVy3JtI2IVVzE6qaflXLgqqLLRVL6HlW0aqSPYB+ErEIh9c3WNY7vTyfXF07iOMdaYIqYV1Z694
dTcFmSXKjGfkWKa7F6d1cczKGBwYqYzdj7K/+aA5xrtZ20kWpFqH4pW2zQROz1wLXnQFfIpc+KUw
oSb5KAGufnkQq4YhmhLqGKIt1rYADimpaWxM8c/bggW4DwQW3OlsuHeEOMUPrlY9nAfKqXTsWHcs
kUApo8MrK+9jYF/L42x7GtdC0rzqSWXYTPZYi7tLNrBWdg+KGL79JXC9HTee28JvRbuXs5fNDbvf
EldxASFMcwGYkHnQbip5hRzTuN7diavpNJbNHZ7+XQNqbDG3vfknjg34vLi/MXJ9kSyZlftudVdE
wgPIacdGUD+sHhXTTXU1em5/a/LAk4ozY8evvP9ZeBbl6p9WWYkKf5LpvxLxM3NFz9o8hL/pOizA
nGZXYPOWvkDwHtfzbJ2/nQDRULM6jmXcLmyZiJzGzw2Tlwg+BBzpJHoJtQ20mEB3LB690TJKpy2g
NniQ1tksYbSidsirfQW5PbTYSTpPtNyZ+IkpBl6yX7xzj3oKd9SZtMr0QiuMjHu2YxHmcEpry4uu
cee1Wy7bn5lUUF8S9y6JEA7Bdo3zxP297Nwln+ZnObA9HhmWEcOr7JH6vJhbdp/PssoZSXH3lNnw
ZSdq/Pvm/hBg+PrZOyv00/S54F99Aquh5X3uq+3nZPXu1XxzhehlFtsZThl8jCDCD7KLdccnCnoN
rWC4Wvt04k7DsbzTjelErANEOP9BsUYYQ0uo/kuHfE9euDDT5ZEY+0bav74OmUpoSQV6nKV+JiY1
Xtle+6EIMve2vLV+Hguhj2M8K6DgoPaojS7aMXIcfEyLcRa4HkFay7zSv/QLLQZtwqyZfqUip4Pp
ALj5L0pn9n7YigyT5OZdVlAmfHTJmTMwbhMWljzWsxkreuflYYOb6QwjXQ6z1Nd0SRm92WEEFw5q
v8vhUK6HaIX+lTL/kO4UjBCV1anrVC2K0FnbhRvsTzWlaqaJX5NqnLH4zpwEinmM4PgKu+yGZ7Zr
0pWRvGNnJj9xMGqySxIdzcrUY3NtGEvALyW/oregQq9Ke14Kod1mn4KEn+Q7eWS8i/fzZ9ElB2xF
pStazhbbjMCnVq6kZswMVVoIWGz7N6fG2jmUVaAFOMTpdqggpNtt2gQQWTdJE3h4cBp802KEBdca
aQUyVkjLnWGYZweca4syEZS62sOXzBDj6llmasSFdtj3sV89mFb1DuwzPzjGvx2sNtfcFB5JrB3y
5MviEZeGhUNYfPeUz76PML9WyrJLlCOddSIrXhDIoVIJctudIZMx6hELenYIhS4AFKRMPrjS1S7K
GHPNpJn871gXhtxiySGxgnap4e7OjdI1cjF90a/6B6Ewv0Py9GZ4OKBwoljoJWkYDfkqZiOKjdAM
OSzy3yHGeUd3BHqJRxr3dX1qCObPYgsf4Mw4oPcK85VvGUglcKE7JFtF6JcJ3iYjExI4a5aHgxj3
fWfQX/Oi1vLVnYUE7J7wf83NcaFD8wlLX47NiyHyzpUBDmEDT/YOcxgdAoE3AlDTe+BLzxj5etJ4
5xDwnZ96Yp7y2R5e5dL3eMMhx3Ynr1pZNOolwxxSzSWPMqmQeERarcJbhp5t6rc1yNJgN23CShnZ
C5YQtOIx1KqwmuGRWqIqs0/VmoJfo53s8AFbaVluEUQXg7A1xKX1q+QZq3E7XlGZDU0b7WX98NRS
AcwMgu0lAznGjRPL9bzAz7i2ZIljdGRUxyLQCecFQdFNPPJ5xW1u7bX6RyVbb+TUZHp5pgGZ3I8w
YlgYpk06FV6vwuApur1P+jbMmEWA42sMK+ovDu0PxFgNc+S+ZbKWSpr77QjKGhnLio6qYE/fd6zj
uIYHZm4tejFX9hDcNuTPujS+iPgbro8Kcg/ObBcvsJmX3V0Sw0wZUdDoVxgZCZSkjfr6OH7eKq7q
dDj8GxSgHKUSbz0VwoSx56nss/+agpADgU0SOAorFehkFzH+LLqo0sWqLW3B51EkNd8Uo5lq5lJt
FnZ7Y7b2LkNiEhbXSybJzGJo5lhl/+vePZ1LhjKTmD77El4VzUmAbYDGVDHFSvgKHc67wkbXWg6U
8bdlaZ3Gihf0xcxjg0Bp+hmztfUz5gfEaFMX9cQdj733ZrLKLJ2zhC50sBUpiuv3yg7GhQmoDpOZ
/Nmb1+1UAVG4VjQsWAZzpbfEqIVr+ZsphPpewh7+FNJOdLyn886aM961OroBO2NHWxp1EVZQs3Er
BkygtK3CaYVHDLmgLJMgH+O/l7tK2mYJbwB5rV2CaflhV7tBht28m4eAF3Xp3GrAVkAdaLc5Paig
xKXapGn4wuvG1shZHmScB1C+fboyEDtV5t+PZKZMWboVCj/ig2tZhOGNSP38CNuXeg/H17J8opt+
3NNXQEuoApHAqunSX2X8K1YSoGF98oB11UyYhdF/JP1PhKjpJMYFYSbr2n8hL3uLMjasFVWdRoYY
ynATXJI5gYg+2o3a0iXsL+NHA81oB0WBdI/Vld0ouosDWXW8+/QViTUbKNhdYUi5hmd55fqV1nVT
IRrVDZh+NwoQAbsjdGkrNg6PB/2QVGL1QkMrJUZSynI+8++175fOve3K5HST/grYhtoIdRbEWA7+
cL+PU28HeDA0VPrLuy5ztzs6sRkf1spZbeOzru5IVcyaLeYSTPMRKQq//St5J1uzXa1/i0zrPRVq
jz9zC/oaP+Yj1V6TFUDfSEnf5Mp1b+/+1kyp/+vmvZ+/HcLjBCqSINSNLxZbITv5LGBQjI4lMQJ8
fa9BrFMn66KqRm3fLM/xNrSfKBwa7ThJv+dXfot04FtjM52DYGjpBuXgRLykF2wsge45iWdJ1LXL
0PjAktXnSe81BPbhGJJUjcReJgHgNphImyJyUw03l1VP34aBiy0DkEK/3mHnyV3wGM2vvKQ5XRrP
w2qjNkp2lRoXjS6xG7VXEOabhccPDgmVH7Z0mjWe9Bemml9wTB2ish83iWU8rrAOA9Ax7E+UQYBi
L3QLvWOr1Tk3G9pV0Q4rW3iL/B2E77AAWcvwrH/p5sjZyuFQtBaqHmSaDd9GQpqpjqMej98lHZLn
mcdCyjFfcVizMWJeDtIunRKdQzE71B2SCAxtxpHoTFwgxhl4jqz0CQd7OCk9CyOYNtT4qtHilOmf
aQbMHbYRICRE2E9GRbnjO7ekrP6qNGL00+CTGcFDikhT6pgyp35eKKCCZ9o9iEH7+eG94G0H5cQE
5fhC1W2aAwHWjm5Y8mKotLlDtGc1HPHPKM2+ktu5QWxf0moC66iEb+80pR+FSM0chFDVJq4KUynr
SlZY0+uyZ0ZMMeeBVJwN+UPbFad5fjspEkSXTbQf3joZv5B7k+r+AP2ChvVsrsuBc+b5+Dbm+lLJ
9Jb6JWEZzALzfOPvssNpfxTHAqwKFJ+SwgOICyPPIxJdRb4f+oM1hQukZidJxcEVVtyWns8mzHdW
tHWINc+NDxDnA8Af2yVj+GAAu6dxXIs/RF8A2kbTon9PFOr4DoAgBPAuUrYWojqqoghhDCexwv+a
xfaQ0setJd+kmJVKAVFwKBzAcFIEyCQpwa3sLWlJLAKHMRXZ+3owcuD+3wtoxJbZEYj8KOz11zkL
/jgVJ+Q7r5QqtZAHp/sPWJBI0aVWjq13V3yTt181drzkIXVaTvfw4h71yFjue8FdDUPVtNSZLxWh
ni5ur9VIwX0bf4GHrMcKB1R/4qFH943sgethZ4idjV8t+fwCCS8zvB0FxUAY8rRLm4YwTIclQXJa
ushSSBD8PJn9tM5RLheoJXH8Sk7xqTJbin6unYxwYIr27awCCuZCqZqk52Tgpiogap3VRpkzHYed
qy3pKsr+KQJgsY2EOCpBfE1bC8lKAJBjqzYISsk+fUaLV9mgEtkK3f4hhP4Ze9AFhXVt9N6xw5Gl
sjjr4KqrbX/ezzmSKoDS8ZIzR/r5ocjHs65dx2lXq3KRR9ktrCOJMORyIIQqPP+1TTu2MYFjNP/P
A/C2d8GTMAKC942s7a/9JBldP5btODVLp0juAYkNUr2ibq2cRm1fERE20oLWdI4BNf8n2OON4loH
QbX3K/vPlLO8G0Pt9srJ1xANdBDhh9f0QqZewMksEpad4FRhxtel3dZbvCCJPNIfFw1l8BaeM889
JKcpQ9odLDnaZshZ3iPoppGo7hAbCel4cTM8ElmW5vPFXaTTvAcTL+xbl34WgLP3CFb3caavhqUS
PB8I9pCBhbRRqvl0bT5DGdK1XBpFQOv9g1lexV00K5BJVBxB2Nqs2Yl/ZGK/MauNLrnpUkyAfGPX
0ywg2DxBeYzCG/V0JQVLTifYCei/l+FQxj31EQxT8IrIe8wFA/yGfYhMfKk/zQ1jww6hkfS2oVaB
3ABWuIE3z6AnpfLRPCbpXKJg45Wgh3ZPfR5YYNLxDlPcDC11zjxq48HqUg94CWo1vB1FiRFnyV+U
NS5akYCDg7Ac7ebNC44ZANN+FzH1u3mk3DchFj6f8cABUsM3aHbDquGBZ1tOAuXG7/yfk5rKavYO
mwBw7ZcvifjgIJbAaQcroRcn13Vge4hT6f+DgTmBa7Rd0lM6rIQGqrE2ePC9d6WitlyLohDmpi2e
aZEU6KlQHhvpVSiGVBQXFykPEiaCOE0EjJoL/O59Lo0QQTqkyVEB+M7HKIFYXBkkfyOLTu+62Q+7
Nk8VsFPIrLDnEdDxKDn442IZRg7lUWIE4q84SIn9uqbjBZ8XiXweNrKJrE2LI54l0WGHsdWKnFKo
AajvnSTrpZFlrkDK/KtMOA7ywupqvXfiNZJS7x/xSVrgc02rYAqw86WkGSQubKy8xmu38PiC2lml
/UK+rsiYak/shDCg4v3mi16JviHi1u8XlFQrlZQ8b7uUi9hDkmUKjfsqGQaZkEwU2fcb5155aRmG
EUW/fF/H4n4Fi8ATFNT0qE5aRCCnWFejgKSfGA4e+583S/bqwzmqEmkuja/KdB0x+aMPHD3V8Kcf
AuBTwYl1brEXaM68a2o0zKB22hJQM33+6OX5TVOW8i7IkQ3C4Ej3VYbiFA5bD9V+hu8I8qpfIU6j
yGMxRuZsqxuZprOkMUbQqDa/hCDxZOIn+UWX7438k7T/n2LN0J5VvlD6Z5nagwWV6BARtVAIgytx
xHLdvBINyT0xzbjuyTvvKLWhg34cOnWZuiLl/VarW2taGnlUj6XGZ8NhhsZeP3BHk7rIE0QNZ963
xmVhZJ8wQK+gpfoMLfGRKDtu9u5hfLavjjLjQw1/RYaZW0i0AshlE5QoeW5d5npnY+d6h7x/hsxB
3//+FAd3ny7od2QTPqj+euclTiHPklrXzUJ/OlommiG9dnusJ7SADWlgqjYPd0N4BNwcqWFF2bL6
/0rYG/LrTLIgiSTm3qcM/NCMO6lRbX3XHmh6Ssi8BZV/kzVDMnzf+TkyyHfSHhPsmLb5Dd1zxQWq
1SYgNstghekhDbuuPQ+XLrwNJmlJEKIAfzvQ8wkNhbimxAumCOd/ywhjYOTLRGr9HqrkFkm/XiaB
qBaw4neWCJ+tz9dBMSR/JTDYsmd5mfOQpkkTVh4ohwM+7gW3EmyJHD0TSFXNogzoPbhVUGCgZ6HG
2+y+XSAR+yR3nK2SuGjqCJwL20cR4BxkC9RkJlXm+ITnVk0DOUW1oQMtzUFPFiG2hgH3Ou5uQENw
ASuuN5TW+zrrCrwz+ZWWmfGCQg2wDttgEg3R5W2ruP2/VtPKUMJVSV600yKcAfi71EzjS5GwMSjO
i2Psff6Rf+VQT0kj9c0T4SX6r84MRug/u3NPiOs4NYAlnQJ932ToxnIauGalbyGDOo/Sc/iNaJDB
vEy9sdEDfCrXGj7DFZLL6Mbq+aMa1G3m1UNIt7YYgzDVS9SkKtoSEhZlw/urd579k4+Wcn2SoHzc
cb90ffqrRjB4BpMpFzGJSeiv5L+e4IqGT3f64yJVQ3GtPCe5mi3F47R4kZksYO6UvhU/SmYnl4vR
m9vfKXNx6Sidiuf8nIrHvtaysrJc42HjAu+Ng3FGebci33crGbMhaJGIhsqOcJcrtlm6GFTDKLfj
z0IVMxb/ukpKm2Cgidul9ImVae+XhD3pkJ7ptEUpFfTzYozBZqgnVTu88IEv4ERiSjSCIpg2P34C
BiQiZ/OaqfBSyf4NJ3bZcYp6VTAzYnW7U+w9skdPYQmxMILWAAHYsz/Xcft2dWGHLY6RAV8HUC55
6oXwh9FRvKPUeJ3cOZx+PeQvayIa2xS9plEvp1MnNAlkyM53eTtGGQU6njmy4WyOaRyTTGTYyZuJ
dcWuj+6mGkEfg0VQ8kXddvuhELMsvCChcaNghBQdGMvgg1nsPs+GxmDUKbpfXBGe2Mahu4xndzS4
Oynm++JhnfIO1cHRmICqyQyZ8aGeTYd8z8S6j9RspxblRz3E1WlkaQO8Oia59yZVFNTyyow1oih/
gNtJ8uCR2QGxBV+g11rA+d0Xh6JxjmGc1dTYod3M4pmP00y4eud9m/AEt20nO6raWZ9O7AAMaIzz
TgduniBGZVf9LEa7oqnVgg0T4d+bvnsghSdvlP7jJWR4ydNAemc29ZZi0vcqog+tC5dxxNRqnYnb
BiQebU/ZiFDsikg19oCMzP9M5OuC7JM7ls6p2WV9bmBRyMXaMo2/HppD2DCtdlFiei4Zxpos+LBM
TQEUpU+Jb6wt+sMWZrrMgHC8Nb+QzJZfw9A+OAbxAapTSND81brnvy90hlhKrC6Y1aptN7DJWSc5
aEChr3qD35jh+plo0xGRs7t5UAckZVx46Lz9tFM6wfnRkOA3wTakz/YAD84e2oBHvPvLgWlUVMAu
Ceaj+LSRGRszjxv1/+DwFlRtxrIzSWLLkQMDSsRlB5M44cVFV9WN4sUHizXMXQA6Nm3O9AsjIE00
uqOPeo/ixyf2iUzrzka9EFIC9yWl9kYjjyaXrpF/DvD5E2UH4+GLiXyF7d6+5XDCZzck/d0r7hBz
AkfQq0R0mx+k6esp4/eFRXF0NZV5mRWRyjqc+Lq6HMC3EEAwNikGDo00SYHcwmsk5HzK/Lk2Ep1n
NU72fZyUbJqMnvBJJY1wACl/zq7q/rQLypJAnF5LFQXN0zN19X83Y61RP7UeGmi0cLx+W1XzoTim
Ue4OOwBChgGtpEMNponoApWwniGgDG+NBxF9Phwd6wVefne4DkrO/5HR5eMfCdsGfR/hk10OPbSy
CoRS/b751LRKBr6cMb/fKCtkyZmKxPAJVav3fBn5fceHtKsZYVl3nY+zFU0HR/97ADwdMUmyyQ1R
RQWXhJ6kqVBvPjvnpYigaBMqS8LuTN/TkJRCYCE0N7uAozJ/uxsddbn1EurJxb2hMd1JWHjIYMAz
B+i3Ve79dST5npDnhxw0BDFAaHHN4m+tqjq10Dx85AzCpUI04p5fAbaqJsFPnSrPDbxDVfsRnkN6
c5jqo6me1VLkKHNobArxxELNcYAGiQslak0D+CeIXfl2Zc69cM5LPpPe6a6u31RXlOKAxhE5GzhS
7FLKrWK6jyCY/U86hLPEDAUTYdaBonlL+roB551h534Zaeys6Ub4N5fudrApWYdJ8pKxCJ2gIgNd
dZlWudsB13u3t3Zn401ypckDsXN2B1N7ZI/B6cpcLaXA4DU7JkwsISBFV+/iSNi2/DBmx8kuy/g2
TH3RyMpwvODl54wmTcpX1PbsGdLtw5F8U/Mo/96VGOJ75AakblwB6LPUbBOrqv1305y+Hvy6wkzg
ZqHDt4cXK+sQZ1TLlT39mFVohZ/BhGEeP9KIlb2RiGZssTR4IGJqStKenUH5pmJodGV2XVuUZwdR
JrJC0p7xI+qUnpf7WEjLVVJLyzoBA+KNAqXBcra3Z+kpaCFlnj9KoRM1N9aYiM7dbTtFfDvqFBLs
UYVj7wsI5KIBuHZIggs1sqeJbI4EzE/OUUrhMcGQcmMUcKUexG12BrlOhrBc8BmnBdWzPR1oTKLn
NUHjTLqO6XixdFolERp4lpE7yjZNSvVzC9rmkVvtUE1vqH7qzF6cAdhUCj/PvucLiTfznX6sJPsN
YdCy3QQMkM6zQw+HZkTDzJWaRE9DySuLOy9uD1TWdewHivl9rd7nlGhfgqjxHX+U8RgM2TTMPnrN
Xr1MjclcXTcbGHcK3XkBpwnLVBcoQEtCpH3CHFFBaPPuUN3BUZAvXwWON2imy9SAHJuD0UMfdCvt
qQADzWWt+ZFPqwUs6Aj9oR/5WgojJFNENIrMT3qKE8uGWGJx3rG4AS2VfY0h2oO2MOdYilAB53+d
mI4WUYKCi9qlCCmBTxddOApea72bSkQeFFw3v2/njYeakOxw8BBZU2q8j9jd2G/Qef4kDcNxIQM4
NaiU2YY08jiWd2eGzJgVdx7+7C/c0hXpqhittGnIPXlOvcx9MrAdiQWEqiT4ZA8o1YBKRQCddMD3
pB8DKFtdwHkDOhYRX+X/lWdV3Bm9A0RFCHsdWezR+/dSvJChOK3QPiGxIrErm/py5RKCSZdzxbYZ
pyAY6++YYJyIMtnmUpP5AFexEIdBmsus8z6Otk5adN+SBDwVRDZyJ7jG1Knj9bsBULr16cif81m6
utcJNgYRfdVQuVhHbK6mZbaRf2qbeM4aim+Cdbz4DwPB0vSkSWyOSeGfB2POnM1e1bd+wxJbCRMI
rqmYf9+UJRS3sJUaRne4cLstFOlbVB79bCHS2ZyZMJSZ8d8a3ktHPkElURQVjKhk5itcjBA4t8DS
TucRrf9SZeZSh0R0NFMJWfEfBMF+StZtrnlzXhSnk4ht0ZIq6GPMv3Bt1Di5tYA5hVYx1R+v+CAr
AXmYFq6vDdAiViBMDMIgxbMRvQvnbU9SxWVDibjkqH4XrmLKIJ9XZ7w59njT6gPgQCcmbGJYEImN
jcWQoCTyj/GHzOIUkCDFkHas3hcNL3rlRDxppMjT/ogPUDjU++dMaADNCPEzQw5lrqonbIhtd7sp
wlmdDZKgAenvnN6YNaiw2tL8n5jEMSnOuClBiBXDt4dYiKmyEsqyJAB8mqS4Zk1k4y9pwbm9BVCS
Uf8bTiHLyVLhblPisurMCj0wpvjVwU1fhnHCpVJQSL5Fb/EOaheKLDOAPA4ocmQZD7jYT3egtzp/
/MCw4BIMpXCGY2ifQgNG7uT5v+LC6LFDz1SyW3dYUqar4YJkfClu3Hs8gqz1dYkSn8YCqbqB+cop
udNpUonxRcfQRAorLMKXBxs0syjhiqJJvp/zmjrvp3QHvFNH6fTsLA1gnqa3l0wvo2Sf/U8Nnm0x
I1HRk1+XuEzmXRRgMVRGtWZMkKi0MSsDIrE45df2sf6elK19SbuoUmR/z0+lQLk7XvSwFlp1zZMa
BXuuL90hwcj918CjNvsHwHmI4/RSK2SzCi4OvzRDHxd0+mWG6zSLByM/3KBdjHoUnqOjuPB5ZTrD
+uYyQ51ra9cgjTyaKURqjsY4CCqSQYdju937vpK3FuDukW00FyqBjWO6hEZPjAxGOP7eg8wpLV2V
Ix+YmydMfsKOAXMwtfyASGo8VKMlB+W7ooT7XzObTsHUE0dR6/BklQpqkQb37u3WkgWs0Pnm7uDv
U2eVzJ81iTqRehoRxnV8DG47mSrhXq3B2gWQtmBEvqG3n32uSDz1UOD27WUk5QFSAN17i0Gf5MYk
f/v2kE1w2YrmroEKEMc9zLUS76JuR+v6R+yzDGhrEUt/oDjpmpTa2HFXSgHUvY+qdy3Q8dEy2BI6
pwfb6qVbRyBYgbGMBtg4RFbzXEN9cItBQDjWiAP3d7dB1Cc48voACnUzUT4nblfeCQlzv1aEhAXM
ompdL2/uN0iVnysJzoPzUyRwOIksgz53hUOdUmie/ZgGTryu7dETgEtWFPQglvfzdNPW5sDq8eYv
/R027iv2lQkM4dqRNdgPyz9DxgAWTNHyLIqrOT77sCD2bknARmRJ6y+FkTU2oh6KIRfu0rWQATzc
4qMUZuZklxG8DsVyv/nk9cY0tL7Aj7ggZqJ2IHs9NC8z/Ux+p+fAl9ng6ebFy3uN8Ygq58j1WCeD
RDeu98kCy2P5jea7mS1xbcBI+2/bZ//YwhKCc3vVf2mPcvbAJeySyeScFp2YS2q3ViaM9SDlWu+5
ke6lqUCIvPgQGNKQOW2tfrL2os/LbC7OChaAg/EEj3AJS2+RwvzGArIInibJjgMiyL/wXkLg9uWL
0doT8zGPNqab3T/BnpFQNbG7CN8rzARE9UzytWhYxyEjb7aO0HWGSn/PLIWhzlhJ+be7m80E+BDz
CEvKl/IKx7hvxFtb/J2QhR19w76Xr1OVVtO+Rc6mf2TzpvkYRDlObsUQTqCaoBh7ZeB2HMErEsMA
eu2PenuGV8l5dzfdg6Cp/gqvvbJhvgDk0VIfLCD/YBF84oAom0iNsulWwDGt9+RT1zXxxrjJH65N
E82wr2R4ULZS2a3CRII1b1U7ALzXjv0JFlTvsi+bMZma3LZfv2S/Ggw/7PPRbWrskG6nKiZCRKLA
+yYURzhww6bdfx1Z5KL3j2ZqBRkAf6OrK2FKyGST2PqG9kRrdYKPBb6Nr6YDfc7jQ66MFDFZZB7p
PZjZs3hcA4Rn9fB6WqXvDCzD18YlDKg4Iq3vlZJL/xXVdk6of4wwix74CBwN42LeVKvYlX+S5On8
azKd/Pqaesi7O5BXx054G984IRp2GMqoBysUujvzyM1+hvDp5TAtG+7trebKLrc7ObX+nlgGz2Ko
V9sAWJkkjKPKiwiBgtF7ptlkUVoYNKoB8LVwNPMuCcoMkx9nOR6IlL4KHw8G20PlkF65WgA65IXr
6Bv6VT08pIe0A1zQZxFORzi9/0++wuwC2o+AGgTtJM+VwRWfP4eKDcE/lsZGX+8CEr5pHQLY14qj
JxS1AtcmNwtgiJcICqs6O+mviZ4D0+WWGsPt0IFQokCzAVdXsjhjzts74NM/myfwL3K5IWruTkag
/7PG1krryP1oqiquihPslecmRKbuECpLad3dXS2Nq5aH5iRGOkA5nOjSKBIehM/qVcsVMlULrL1a
Xh+1D+TDCFOvLhAyyZ5c29uYuIcCoo0M3/R5LfnptUY31LoUaOzEkaJrJ9CCaB9QAy+CfZTdC4Wh
Dq/qtnh1H1wB0MuFRY3uR+qoxvAgr5n0P5cIGTfojPNvVdBoNCg0zW6nuewMk2YX91nHQ3EnmjSI
0syUErxkm7TGiYtYYOqvCydvn49S4WZv+TxUI4ssYYarfGPZklO4rCQkp9rfUVg6B7FCkeLn2qRd
A7IXAK9p5UFSJtt8OFu1Kkje9U/JsXvnmFmEfJbWQDKlYyP1fjsHqIRGFXJNtTLUuve3d0pZHhY+
dGn6wNUtC85Awt9C7WAPT2Jyyrk15U/C1aSksrMEe+wQj79OmmoPL9ZmEvZQq1VJbJmD/EMONxmz
LTwTGzvwJdJQPiTH65TriCMOG9CSBHoY0yJEN9EIp30SdK+jSriLsk2VQ2wxe/GhzTwVsSfTOB0x
dqE8ONGJgTWPU8of5rZqjEtz6DZLepltShkZKL6hSMBd9Lf44j8MM3F5GrEI9Xahh2hDqqPG1BZj
e/8F9dYgux4Gv8FnAt15JlQ4ZaHwVYYmiQ4EbLhiDSmxDFntAcLZmaBJmoVIjhv2r8QfqXyl/WN0
qC6MtcQ3BpQwgFxgKhb8Rm2rIa1FJ1sCGKVNhMR+7O2FqEP/qfLdoviQew6BXOKO5eyRQkK4iv9K
ilmiyaOdW59X8OOVSSx/OPrmqS6NAE+8wwNEie1M1Yom60/Lmu9jxWSZ5rN9Pv/5H1nwl8QE20ES
/wudongDAY5+Rbm+pnegukzVtuew0Z5RTmNbwBwFaFBcE4QekaXyt+HbWeirMRop8RKO04ZRb3Zf
ZwTRgkUxKpb4M0WrcB6g5DrNSM/MiZ0elLuhYDlGWcXfZC9HyyBhk/F6PyEjl5acnafzBp9RBjxx
DUUlinUuzaQWSiV83E+gtFaiSfehbu9JoTOcVHuZQhJfCmPCURddEFj/tel06miZmHfjlLhEHkw9
LT3nPyGjZKPDSgGaBrlwts9wOXjj7iAIO4BJZ8HViOn3Wtpw6Mm1LlDhgNipB5cset40C9QmTpkH
GGANLS98n/eaZB8AofE8JiTUv3ZPJYZMVQDTR+rJC64p5VZbu7ZHKHCVxSFxVlmv9E2XenRaMaS3
NlBrxtD7PiCaJ6M9Lx5EgByARDaRYflZDxRxb1FlQPYYLZejXeqrUwb4Lpe0w6s5u0+QQlGs8N0R
A+LRkp3DJpbNjp0JEt7zaCPjXF7zAEFXzym7jhprnKjDcba4oh4nNAvbFz8FDNjehViYE7COLv7x
hQP6V6XdbClW8GRdMMoc1oZL3fnxZ7gjabW3IXdqpfNH9V70kcOmnRb4y5eDBptAgL48EwMLllU5
hCvrZpoK0YO3OKIu6OCWv9R7YJOTFwJMR+gBhhh677jBQ3bDt9Z6YkZ4I+tNX+I6uVlKGsYG2q91
RXx1wtKek2yZpUA/32jIk441h967LBSgHKGCwfVAxHDCTpTVRaVC9zPmvm2K7zFyY6VXTALAMV+L
Whq8LZZaXrMHdgMJh06mM1ovaNeuBeU/elsqpPXxzPFjYqXEv0r/cgWR/evvXmuTTDn0BvPwK2rQ
1fM68tXDym2SReN9kSG6Gmr1CaoMSlA+SZJ5RbSoKw1WmF6p3uKHpoSqgJ+cshD7u4Go32dGuTi+
AK7EPz1RHcCpeBEF9FrC7T33Y1KpZQ17T5HaeOI7iWzKO/nSOAokJQvyuFtDh7t5WoqSPWp7dp+I
NHSw9UYZc0kf+wSOr1YgtbQzb/9P5h6ayOSwhy1w4y3KoqFSInI5UOKxPjnULF75XRNeTScl7GBm
fDAA4u5qtQJfTF1x6INsemLq5+MAgLm8kIEf+r5AtNHGz0D6tiMylQMezY67qZbGNDgIZKamODl6
8tXhuKoZIJVQ/XD5wkbjkdf226Q1bvMvYpx20QfO3esNaZki1sG9WJFC48QDk8/UBgHfMriyBvHb
g+bEKHfpq1S5eVqrbXuJHJrxSI1/4L5zw8YHk1Yxg21yLXMUg90rALuBz7zY6FrdLh/3Fi7XKPOD
F2JNxeRDAYV9/44L2EzP/TvjTcZB397W2DBjnbDveObJ2lCAm9yUzojlycvTDllleWSvzm8wDFgk
u5/o9lddHkpN2AsDbwB5Ok6gyqDkCjlTz2iJVgEndv3YqsN9cXwd/5+a0qLTeu7AKmUC8Ow1CF7p
Wju4XDH6AJUyV5Rx9+KHJAl1p/rGsWpXJSzCgxnIb64uMI0KfbUMEae2AbOnL6eB8owidXlaZkoW
FDm9KannLA4RBH5zet083yhr/cpVcu4ipsL54E6bwisbV/68S75fhrHlhLX+tDIQifC0+m8XB47t
HUTkhdMCzp8+HKu+/z9V8bUkUIsiIUkA2/9VwfpE0elKHQGvqLhnLQ0wlf2bLuhz8o75Un76bm4I
zAajU6mc4XugfPDC6Pv/+fqonzWd84K66+2uxJ3NcQI1y6AHuArbEwV35zsA/7rcJUk698KlVZ4q
aNMz3VYGFziyk9txQ6MWRpdkFKAWGl9Jf9TsOOJKL21hFnPOHyz4dG9qjeY4QLji2al9A8u7SpRk
U+Sgbuo7dfkP4bOMIE4KXB5dMgBoGhMtBZcyDaPTdbJzsBcz+LjCluLwQ4jl2kc9uhZjj5pMD26p
8+vcjtVHK0w2f0oPD+MwOdxs4OfmV5MSSzJlVJNUZ0EkoYqYpArmqigepXT2ERmAbcz8P6CAnMyc
Lr27S4UyP6RAqnNw7eMebkpH3xG/c50nl/rZygtkJRCNccci+YYrycLJbXYfSBf2jZqgAdRQTdB1
uU3KR+4gJQKH29zjELQT/HR8WR27behDu3yI9OpmfXGNLH3zBJB0qeXvNIDLrYhK1s40pYdH8oSy
Q0y4pioIGWkE8YSBCc2L1RIGk5iLto3WydPF7XqsOQsSBqJxVaEzQW5tvv9viW6kFl5uwSW8v7ao
iNuuUxoRXsG619frOUvjQt0tl7hQt735DpsxEMJevcO8X7jPOqexE630rtLnTbaY/L5GpYgbNCjz
uKdg9cDIYeTpnBvwht7odcuUWu2SvCHSVGj8X63L/XpS4eIx/REuKE9uqIDP6ZVPrho8vmbI1Q4n
v/QUCvxL1kGRzuqfZJKPnViUbRZSCDd+4p6bmLm2fli26WRdmT25ZCfxLw8LOKDxt2uOywhpewl1
hQ/NSU6vz/rtXbOsKrVZXly7xbcUT36+CvxQXBh+qj/qHWBcWgFlcvliibFPQ9KqXyvSeaX3YmCk
C7EeY3Pyb5N1eJ/qgokv/IRztM1wgta0KocjuQe/QBu0TYkVLyr4rYOmjgY1QaRllPk679kvWRta
PJCTxgyoBYH92Gyvq0WcPiioMFGwCTztCv8pYIrC7NbwXRS1q5NzN4cal8vGXwYDby2rndtr6TxB
+kgmP8OPq38IMKu15gpg71uMa2i5r9PklXU8dTnP3gi88hOEpRoLxhQQL4bcDsoYCwxTnYKsw1LZ
YQUq9qlOXilIMKBxNi3XnE//gpFeWo8D0fCxId52wrojhvrmpR6YCY9YJF6TDT3ACi+PRJrshcQ1
EsJ8UDcOxdQszjgRLsUNbmDoDuiMPu8DKeBah2j8Po2s2q3d8hk9cwC898UhTZdDqywGTFxjaLrb
x1wLMusSSX/g0tlGoRU6gMYuEnwJKWgSKl/Mt3JZYGPFJrvQg4u29tZEtk0IP9xWu8qZHIjncBaX
S8ozi6+vPO3sUS8YWTm2uddOydfdNDun0oSqlqkhzBYCK0L4FE7gSD9FhnGkwIx3K9/yFcc2LMM1
Q7NhugoIrvq2GaTEaZEJ6NXBRrWV5SWUJjj/bPlgAsNQN7rZ/V0VNlj857Cyni2ylk3cHkPKwfhC
8FtmfWrHwPNGkaNUOxJ70ShLnJVzZOv2V6+B3iqjwPYc1bKATJQpXbdaov42I0kJ+72WnJ24OFax
mAKF3mitAU1pDPX+zB5yBtgB4c8I/NMjcssyMADJefnYFUdTWS92dzwHP+uT60IiHHxJ1i00YBY6
t+JF2BCHpBgbYSHmwxlgC+N5QhdTsvyR7+KLXnMrw0iCwjYswZHzxeuGeYg4YRFuIoPmgaFUTYr+
j00+r7ERyxFhje2opsgOlwVLWhOBTicRp/OtOO9ud05qMKBWRtog7kBkv25JYiP27TvpK4eIzDiS
jxu3ikTFUR7vUX/GKKBjZs9SnC3mpvthbYEKfZ0Kg5uC2+gRzmFAuFQn4bxc8x+Eyo2n+1EfoUeM
njYcWCOEfNrBFnPPexT1V7Ys7EXfe0QTY3Wpg8HNtLAeOATEnxYeaEZhpMx8L4z7ddfVkXY8VEoD
LGJndiJ37xSKjT4akp8AqfbFPutSJbSddtXk6pmohfq5u8m2BqMISJPywiPCK0gvC182j9kuamYD
2qZUatIOpZIJdYa41XE/DHzgCHqYoAMAwk6zg1gOWKjEHmn+yzqNjCcs6asqD3ww/W8nBMihWDsf
oBPI4CAaGlwyt9STVaKNCYz+NYJtOe0VbPW+KoQXqDRGT6ieKsTIrTtbRvoN6H+U/z1FPj+E7W1r
Z+9fXlWTb2jGQ6s48uo63FxrUiXfog40/FsCDC75zZGRbeE9YDpY6Ea4l/TG+w4fcQDKJHThYrfY
uV0ZM7rwJB0+EmhmUUq703zA/CTL99FH+yAjN+BWlP8fr4UfNNIYCN4S1UyD0r/NQf6j3WzEPi3T
OodBiXPiXF3Wptew75gtxZLGURqs8i/INS0nQBFRh+XL0p8mq4cE337L0+JE71aIcIyqmGCyzR+5
WgCclOZ2kaCPNrdCqwnei5yctjNlekFZf1sCh0Vl+j+heW7hfhNt5U2beE7TSE3iMHgqeaXWH0NE
rJgVBp8eYcPGsEyjpuQdoLcXSwdsIBzUb51WrefB6BWItebax6qd7wgZjzwlK6C1XO3WqNssohiM
JwFUjqwA8zyqqd7BWDNVmRejtCb2HHuUHbtQUratiItBAfQECNvC/u7j0jLyuZB7qVo0QRhTDMSy
d6W3rCTF422l1yqMp36tQC4uhc5qcvEWTsB8nD6VJ1BPuBSrFgN9fF1WJTgF/2J4S3gpS/819deQ
PPka82a+uQRIVTQ3/i8h+qgrGU5yuH5S+YiMRTC/Id+UVouLsa64NwZCmQblFocXmegOPV8gmjiH
zRqd+EYaKgIMIrQ+rVhrzO1XxLIWZOt9+MeL7qbco+jsjYcsWPlZKKvYnysS1v3cbiMOmHeqIork
sWL3LqNckBsF2uVDE8hZASlnlCmBj4uYpYO3wgu2RKDCcbVi0iChxf2wHqp8ZLkc0UI5czlrPz5m
JHmi6gnlaY0SYmXrA2tanDkwkDHjIhvy9FRWD5iEdwnD20fwxov3RtK0ZN8IABHA7W8vgJL7SVNL
xDIYnQCK8Lpk+Sgw5znWABtCj/Q4DK0RnBQuMQTOMHlUoP8AlJHL+vMWhgXbxJisKEvmk+hN8PM2
oodxF5WYWfrQdXUHQqOVKgSHstE7m5ETm9w77BnimJ5j4+7Vwg4vXdLYbdU6Hv4DgFFamvo11tiw
0LpYrPGoeShQv7IwUOzb5f/Nm1wOdBSYiZ+iSuIOwDT3s1D9lMNGshvY9qDfq/tJ/0rEla68DS7N
7paW8SYKopcKRREcyNS/pTVwLh62LSLj1uXJw1aAIAC6AVlJQ5zNMvssIMCvfBeqnIirhsKl1F3s
i/fmNhd7/S/wCnKhOXvljw+ZJCtj9ttPau9kBpfB12kLuEZSFhusis5EMpv2Go7EoawoklntP8Sn
NLDsTeyGLhufs0g4hUt1sv0BwIQguv/9UIMiYdIICBY5FNkzGhUpgkbNSMnxC2pW7u6REmFSzKrG
UrbocaSWQbP4aelP38DhWS3nNutm0mtPN+L4rMbGEHUoo9MCkgWA4kwwrozyro7u3FIGZUiFq+M8
+fr4zIuJiJhZ1NUajouFLMgEc1kqgv7BYBn6ERPZ/3gQbfLVp8BZEAspGR9hLF8pfv4dywM9W2vJ
Dg5IjDTg5w0NbTd0v5RUGeAsS/C0OTvD76ClsC9XceSzOORQqKUciWTQYkrvacFGJSxlBrDz5/in
1bdNOu+KXOgjHjC1m0S1Lw9hTdH04MtAd9fRiDmzpbUgZNqKwfkXqmxGE5Y9hBJJ3c4lBExlMKOC
K3DwqkBz4gxxDt39h1KKmrO2YEmxan9I5MJOAuJ+5Y93si6f2xU96UxrrRwMQB6eM0ZLN6ATyyeo
BgwrQbwpNikjcbCa1VLx5dSI2bvnBES6I+qVMA0r0nKeVxEqjNMLC4EGY+JKNVm5DubGMjFLwKx9
8L0MNyKk/K/OarzQkxTMEIdCxtqpw7NxUhm0kkeTUU5OT+ZXDeIwE9su1/Fwp8Cti23janEXRdqP
5FRTrxwhzybHeeKjLJSmsxY88zjlo61E/uu6BdhSquJWVWWwVCFQ0RzQ/YA5UFzu5ioCH8bwxt6s
cnvmglNyhL7ur7+Jb8zUS5X06GU6glzxSoXRvn8yzuHbhiTtBtnXOCWtwJUyJRgKkfaLMUcaiWSa
e+t570xMc/KtN8DKiXlahzP7Ddq7x/5eb70zxX44u0aQMaNW7k1jHbCAA9iDxIvBetfiXgdKZR3E
MJY1ojPd4Y6KC1MVB3BWgwl0Mt9HiJhtLmkfCevH6RIUPglyErt0EVUju0+8hDPcKgd1BHzpeVpr
VD6SGM5H7ojUfF7YVfvNZM8Kd0l80zt/TOx7tA2FOZ2RvCulChwIxWnjDXIira3O6Z/B6Y5WZcDU
9tY9Bflva7We9fG/98sk0h6EhpoK6MtK6e60/amho07Gc3YU/7Y6kYsJLXsX7pxfLeTD6O08JLNA
tQ+JcGHSnV6nBftE6FEBV5XeebPVDiiogADXzse7BumaQEA3okvPrb67yTC9TGFt+PdVNildJz5T
/uG6wSO69SaOvYXbhmP3hZopLZB1zEoYvQWJ6hNEd+vz6qcbZO/RkiROfmt4qJtXAz9P6JRsjQOF
75p8vxTYojOyrdq3eDScdmiQdtJOq+O9lMaX4qtktfvryhZRvBtk2s9OiJ3q43t4Za/NuREtjfwM
vjLA7xCY0U4kJA73dudQpHPWiQwMtuoXWpagvfrP3OwLdCHB5A9bPwAk7we0fIAm7CL9blOSOUvG
Y5UfHu178rplaCaRTk/H/bfqAsVh+YbJL60jpQHyuAQYMia2sUNCq1KFvkMvMwyymEfK4h8JGkcc
1TCLP1miwCTeX2XGrk8FqCnpiX+DqHPGLQyZBqrpHRen68Ow998qm/mM2DLEZH3LVkGu38+HzOQ5
SjRB7smOrqNgyG4M7aqVyGSzQ9PHoOIBFbLoeEQlThItwHYBRRvrsRpz8XDMHAW0iYPUdEP3zD+2
m9ahsMQJAM44YvD/XHRS/SC0lU6tzOjTyHiboMcixPEKhP7Gbbh9itgUvz1yaOMxT54dLuGhhdfO
G03epq+zdUArqe/X9Di/b66ymW6mC600tfa8Z9uVThzBGr7fLQH8HVeXQQl1Dp2BQjyho1IYxoIm
XaDPEdrLRlUIA3Y1ZLb6d6cEk3Vwe42c1GFvpiN8S7axk9d28p/3UZSQZTtPiYkIIBLZdMjbqzNz
pgscvj1Gnd/gTFxEWgTV1TQ3o68T3XvPgRbCdDq89/EHG74PpFDc6ZB4QgiCZJmPGem0A0n1nWrt
NIRwr77w+WpO9ZVLt3e+Vha/1YA5nmscLDW8ISXpfFOfsn2lJNxan1IgPJ84yVVT/eQZYTPG0qpx
uX1f+Ac0It9dyUPpL++lmED0qH5VsYbo7tiyPOwRWqdq6ovyS+udNjz1ilLJKu9N5ntHhB4Ch9jR
6M9qDKvEC9V4UKgIEnGYinjJftBikfdsLKEXfPbjwSPh1X0FXi1wpjVdT0gVy5vSp6TyhvIqwJ8p
RFW4asXwCuwzPQJ12itKxykI6941SwdBP+tMJqnvkF1pFKxFzg1htLm/EWNu+GRHyBn/CV0QiAmU
eTmj2R8yPMRq90uCQa1vRIqDSQ1MkeFWRClAIK5UiHHRwsQtrXSvPE4hAaueCkP+pZ9CB3x3fFG2
Ti6Qvvf/0SHLlG9CqKGqcAuLPa3fY7A6co0/nPqfPe2USkuV6o2+QEccTirn+6q7Q0i4QwxhyZvk
9N3pAOZvlYxC8b61epjVNd2Q4ABP2oUVEp5HX7kVUhI9IETSnSWrwrSGm2yl+DIPkKhiD/1m+Woa
30sNsrzUIEC4SaiG732gahH/COm1KNeWhZAubT6TihZjlXo3aFGqsl2usyG580cxy9JBqydtYmS2
aUrpvcxhJLTaXBYY/pT/hrrQh8tGUdHLfaTRNSagJafR5H4SrICjOJlWFVOeE8jJcAkSODmzUIdh
m27JRQV+jz1G42B4Ijb1y9cwN2c+XQWGLJJBgME9565u6BmJ2Sqr97AHI20OnotuI2EagPx5BTYz
HmmttSOgwKCHFb4VxLM78XMd7/nJ2mSETn+1UpJ+tx0LqW0QECGjcUVJV7iRILWeTn7Qsm6wu1oI
xsW/pWgOtEa30rq0ZQ6t/41ELJsRWKniLNcr6h+OadCCLijZV1JdfBq4SVDgMNhDvYCpiSKMyU+8
UHdNyvi9mr2lQPOeBpTIfyLIEyXUwTZwCFbq2t7A9PqKxz6Q2BfPqQ4ReDuPRn6D/F88eOAGOMxt
BJr9WUSJUqG3PgUYIRlGCOevGPViD99xJTHKtQ4P+9xXZvYzBz13C5x5PEMjj8//jhO1lMYbCLXE
ieKqpG56bGbWgYEWSgYQId3UAlsgD/3pv2e3vf4H1SbiiVIpqYSW8T4UUeca8sUQT++6qxeUpMpE
z2+TIt6fQfgzWJ2pcWcE2UxbqQWsmcKOtaB6ee7ei0brct/C28S6Q2C7gHHMtZ66A2x9lr4uk1yV
sTUvQcRaSNV7WvSR1FuRJS0HW0yirFxfkK7PGVDy7s+rJzmQYFGMaJy7MW8Pi0EMRmi3lbsWwvQr
tD5bhN0ZMKJA2CER8yxlr832UOSqQ/bhnB2sjcxUP2hprvs0V1+c8jRmyQGNvD/CYndelPDMbF1n
2clKjfi4X5yMlS8c3K7AXyUEvwqSqK/1mmd/gNTPbF6dcZu4lMAdm1ZGKuYVSycLx7NquNTIujXI
M03mjyPmdCHcYxAhHv6QPaH790JucVlcwraXzSBH1JebbnxPsiipMIJnXRYL5y6eSIde8LPwOSU1
9uJwxL4Jahdkksj3zdvQcdTPXwXfpvsi7AEXEnG9VMbdfXcfCs++epxSUCIzs2XSfTQSw/1LU9li
m6nOYsmc1uqwuvLQkm+aRajtQny5czaaR7jB3YNBDInhoKpO5ChI9H3PAVP+iTSvAwZRu58Ro+yY
DzGfv4izf4RApH8S7OuMvDEZEbhhasCCXidujbIugI/qZxZEJ0RRQQQiUfEBchFA9Pj9pNpXNl9R
5FW2Y2PY5YH2OpAl8QjPh80LQ6mxbQUxoXPGcoJMdKcayFVkERfM8ASGq1eoWPp2VtDUNztdCaBO
Al995fUBwuQhefM9Ao3JVsl/KR2umuziceYBlYfjGXr+xDBUxhcHLVUEPSg9L6FnQ6OVXgJy/GRX
rKLrKp89ty1uEzO6ii49b43VzYUQleyl3ne+zUPsCg9FAVEHhTgmOpyptiISzYXUXH/Gi1du+cgM
A3C3tku4o4Jfarxb8LxjTd/PgT2ySuRHITDotImkAP8zPi64gKV0cp6bMr8QSBMp7aKZ5IjH4KIX
R14oEsRwoY9+cu5qxkIhdhr1qnnFpI4m9UrhJp1ug9cLKsZG5qhCYaUeeNsc6xLWHX2c2W4p0HqU
rCkUp22F0mCI95TNS5aPobYGRLWI5cyT4QFwXnEA9dFcy5IUUSk/X93os2mkxQz/uYuAmsobdCY0
XSLvbCCGO8Hm79hlx0NzP7/Kjk6v/wp20bXCQsDnjuyp8hDMmSxUqa8/AOv2AOo5JI5LDxWlyJYq
o9LiT8sCH9ukxNVhAwhrgbkfMmvYWDt9y94hpdWwu9WdeYL29Aa4REwZsBHVrFr40uxyxyYcv77a
uM0vqMFL3ofbrPkAawXJJa5+457gyY5ozTxaUoXiD3NcOSKYLV26izLihT4sWq2lybwvZZE3/w/j
rWfEJbEMPX5ZjpeD69AaiFhz7ARm6gGNNKtNXQhM1RqFis3MaSkqQ2A1v40n+BVTMDRIKmNe/78F
mg4k3K7PCCEIlQBLCADXtN3ut1XA6S1nRT03sK6uQjE/L1KK9GAGgLArL2NLAIwlKP+MkhFEGk7x
87vDoCmiBt3sFVLSQ2KR4uEzW5vjm3OChCS2rHAMcP6gNd8D+pN13nfFrza1l9mmopoldXXdEj9d
sTrzbUrN5Qz2nQPjaLD6UkWFnxyqmGORHsU1Y7EoYkTJSndSiove3gfuoV41TV8S93be/jWGIH9g
5K+/Dy5R8PPUGkDe7DU+jOpjBRpV1s2SOl3w8bIFCOOubgJ24DviEgunvDFclCuptC2AaRTt7XLW
fv71h6pPBB0SeBoYHkSSAQ7NlC4iZLfSdmYLKJ+yJVdtjtd/+9SaDb6tBGoVf24+Qb7NZ+WtmSMV
9QGLz+yhpM6I3wgwLo1U8/GC5j5UwafAAqE216GiaLpk6LBiJxbwoaTIwC22rZ+tFdQajB85qJJZ
dqYZer7JSmY1G2uCK/uNcFI/NTvIkEPND6g+LtzvQicIUHbGZ430KxGlgunBVcHigorxyraRXIFg
lPnJdS3QFM/MafP3PFBPOu2n+DjKPfMUlirpvm+oWn4tL7HbPSgwomWIvkKtfmlkg8px2xmgn8Ky
GXqQAjacngD72JsFzLvKXqvL/zG7hFT3D/wqWA7NViVJuTdEyh2pxhePz3XYEv0ajIvVOeg4tUMz
SWXD9C5hqZDt9MxmczrsNtpv9kVFhgxy4gPot9arKNXzsDEPknkw/XzMbmyPoaLDmQgv0t+W6IdH
xX1ab99afM6Wh3q2jKQP81l/vmoIIn27N8SNurRx/f85mBMIxmeQJDPh5ftqBRmDBWlPV84qcXLv
+Kxw35Akkvq3KV1Ca/3nErcHNlU7SXGO2ktk+gWkSqVx3uIvfXgVDxZvX9rjSnG/fWRCFbTP3UZm
kCdVQzPexZQtaHY82KB/6pAgTNM6aSOLpCJuuneXCcsGx28Yjl4lLwXoyR28GuY/fv8cW83/K09i
2LzhCsqf5qiLpOpSMFvxygTDy/zR28HgHymTvft0wiL6C4PMXfj+5xtuiF8KP+EggfKKABrbzAxn
BzMUJyKf3H+8qC64uL2ZC/VHxlsSyXoXwhxOIOViHbYRNYmN4nsuYHba74SxEETDBfohPW2IOpcR
vv+YXjR83A8fxlBqUxIYi3uGdC00kvR7m4DYF3sQ8YgD2APqv6mU4MGBW9xm7f9GZ5HdK0LtY9Ez
1mv0nbNq/j5JcBXYKW6IWja3mrYMEKnArySTBzldS05PAKlNMHux898BQOHW1+3meFdX7nbBB6bL
kj+KwtkZUknJojh5fOSOQxKBqi0XuAleyClQUzTvo3x8wNHqa9votCxoxGXLgH0DLNX69CiDJeoQ
7RV2SG0UN7Bhl/5AiXlhm6QWYt/PsaDz743hUiN77dpgZflnFxJ9zm6zXvvsgPmQU5EpJWivnXCz
uduKJAfwmnQiwKYu9hhHEvF5V4fl4q16ENL3Od5rqaHnz4X6ApmKgsx6RJDfulWz70hVQU4PS6qd
qHim1RrbJAr451Ev85eLmNfwPFE6PduqnQDorIuNQl2D1M6yiOvcFEvipgqgTfK0ievCLcd4o+AY
qQYN805xNAHZNDkKEpCkSaB9h3WWPbgeo/gsKDccfupxIiJRLL/ljn5b6UqGo3rQwXp8rYyQOc6L
mb8jg0uDfUQ7NJwtBM+2R1cTPdFQ92G0C5y1DkUdXliQDWGPBTdMajFrst8ajMYOuOc+aujZc5EP
sUS3NadvgAcz3laT2sahczz2wDLfsfEGEbeyUzdhYsYtJNWuU/u3kZR13ULfHQ80hWYFN1a1/Nmn
EsQ3DK1e95jXehNb69P/kHr9ZCpOwhmUL0MkTGW2mwalNNzjSPdyJvau68diPGUyvmEVYm3RD/dr
IDd/cdE14rcE4HPArRozzsjOM+eo/ympJ/s3ZzYRBhPl52GklknDL4wkSyR6B1jFeS08ycQ5pd2j
znvfe5WDVuRoyeKr8BVlTExA1R6ykky/DpkdDYc6rXwAYlAGr+QPHz5/9UBZ7y9HAk0Q0ApPYLZW
pqPitgcd0F5FkGKjPb9YKTwWVPIm0AaYmmnetQOuG14ATTv2C8g+yms2TxlCbxkA4gchji42Z7++
BR03DT6KT6OIS6APTujNg81jS20NcXX3h9R/O+2yCRCI2sElUbxBDGMoD2dUQjbaVKBuJIn+A91A
ar7H6ma47/EprU76e29uEL3c6YKCbeuolK7RzlYazds2wuN22rlJvnEgJmjqoocYuEqHtZbCBhhN
Z0shTSe1wSfotLfd5u7s5drv4+QaG1Fejtx082zeRNG/ULrKl9bwFpzqrfxfi7mrCohKaXbtckJd
GbWm8wHeztqg2CiDQApdL41SCI1VuQ6/1qCI2SSgOpiAbukc681FU+/n4FI4AdQLHSRolXLXh7a1
Gh4noIb5Xgng3sT965oWufK8/HrVvQPWSqoG6p/nc4/IAAwGZd+7uktNVcJlAuQMGaKPLzdEqTPs
uABwTdvWCgcIzJcVtBYuyLNd/UhDeA231u0z1NeTclL5YFg+Tpidno7bI0pCmymijH+p3GUf48cP
2Q8iLEl+oLURWSJWI8AlNoknNRhFi4keplloNVON/bBcw9KqYKhFqAe10m0WHLeZriqVyAiXLXzL
8t4LcYZ9yYFJwd1tnDepT/9gX7nIv1MYK9SCmReA3k4m23SqE6Y4GXWVMEi5+5Tnz8SP4ISN4JN1
jzcoMhcG3MQfPJbLTOMXVxt983mzQqX8wChylmjNm9VRLQpiB8QUwsyFjvKc7TlqS0r0TkDc4blU
XZTwFrwJCsEuwG2g4UpuRtoxq6l2RJAU/i1YfeufbkyWvzIeQ71FnlVpt0kmuoKfxDkYKuLNxxvs
WHC4gcEodB7IopWywoskO5q0sZ7OL8nzBWDeEO99AnmB0sSoRay53L6ivwFm5OUL/JNKhISOa1Iv
xCPJGS4OBTeO2f4PYc9YpXLyM6ZK7zFuhyYgEuvroD68WsD+RWe8NGz/duFiK0tch+b3ImFD5aJh
F767p5RtUsEX/JCPnlc5pnbNI4jZYlJ7OUSlmxgCl8k7Wpe9tOLOiklHnRUdiCM9wwzhtk0HL4YW
c35nDOy+J9ZA8YkxA8Bu2r9JhI95EA1pVPfikzVPy7iqsLTf5E7zII7V4KIL0GXJ+AG/JnC+IOu8
JUGCgVfPLqgx7nHNWMusgjgWwNWkI5WGbLtFqP9PzaTMUXz6y+AaGffNqSOc4uK98l3JsHiPsiJ3
nXqYzhgAn2THwyJ36vC0hdFThNvFXmRK+RbTWLmicT9d/TEWXZW0zxEFytiQdYi1JFv1T4F3lwXK
Gnn+D3GTFdNQqmKR2ypy8n7f4nGKjvmxqVxP2kQw9HOOMAlKIN3RDkdUIKcDes8uoUwWpNQMj/CK
E6Vh/M5nctWZOTO/Zkxc8qHduVcFsDLaVwNI3+keq0JKS0blSbz26ClVbZqWyFSkctdFMZMVuvRk
yypfuDf0xn85MIb+J4V9ySl+FfjRvxP+PLFjERSt8i9bSGq0JrNVUSDzHzxX9zPbs2NynI9mL9cd
bDLHYz9E2kj+vCQCb0qkgaANWQpA9eRFyYjYRi0/9+zdFTDDSISmvkmugjffgq53UY/mM/W8OOAA
5ahaNR9EqwJI1hF4xACsGwPUfSj9HyHGL80dwhJRXJNJOXF9HQ0QTubENdzN59IQF0D1L/gkNOU8
ZgtKhr2uxIJ9RrTwxQLsBbWSIJxwo8gRlpxI2697G74AoGihHdH8xV5TaI4CJA67ltAhG8I0PdTS
oB8UN7nEwdNg/32K3bKdi5ksCkSFJ24yWC/QWVVx3+R1PCnPqgvV7oi8yZaxb8Oq98RndfsuXIQ9
ETv6iO0mBwGU3liuKkKSCsSLXkeBL0gYkWKPzGH7oQcpHeazXcLpouH31CDrdIx0xhWe3eEph/n1
7RdgwzvsA5TFL2snGRTdHmYOqCr9pTpdDveLKkRXKPv3csZxgMDawRfDZ6e1lIVsJuNaIbvwGsQu
3zLQaHUbPLFkuN+cWLfjEDKjQMH1SNg5tXoeN7E8cuz4TZIs4wDi6iLCVDsj1/5u5roVJlw79R6e
vnra3vmCs+RqrnMTp/A3WetdfMvBWsoqmTalgzSl5sIuBz4z8is1TiGWWTVAHm6OGtGIwmGGnrh6
5Fw58Ia/aHTFSLqvmpG8M5lo8dxhezqHhN0OXwl8OPkZVrV8y+Nsw5dyezfhWthA3YggEGJQJG2H
k5hKqvVZTqIJN7Z3DRHnGrxkHtEqqkqEdioFimzYlBESvH5S0d3Q569A3Qkm2NBgDpEL5ag3MVCl
fUl96ygcIuaPSiSr63VAthBiW/9/vwgayA2lLm9pnIaZVDQ2tMrAqzvNXjPiaOsRKBDxGipHEDtq
myzyN23YSzZeQyoe9/SWHlbN6tqeaOGqGb73PS9JMkDNJluDq1g5ZhAwu1f3oE0YfeZMLDL/qQ4D
Q5OsOxP/wXk2SQHB8T2puK+TUnUxGjrXrhy3/HWr+J4v6aKVyJgl1iyXFh7UdOoPScRnxmcWpFDd
FYevFD5BTCFZUxo126cdOSqEeYhFcAHLUQKi+KHdO06w1+7yWOLZF0mO5E7VjQvjgJ98uL4JHlsv
52xa7DEocC27MxvjhOzewFQavXghKlFaNalq6CZ/nYIrwFboireAUvP1aWxhnvaKRRfzin/38X3j
+QqXMDOvaviwdyOpQgTQFn0Dvs3v9ZfDS0nzzDmRharaU6NSf8bVV8oYatEa/FhNclFypBO11oPF
DFDe30BaMcWzwVTivFUi2yQhhKYUAZrtKpSNJ7yqFhwbAOhPS8sZ55YZ6bZB6XSyT+90nbgx80To
WSv2h25LPaonsGV0kIAY+Js2fnfwKOfpK8sQeMtxlGNdyYWA7naWr5luQNm3GWIV38cLBfz87d92
9a80JCniWAIeYv69vt2urJrTgTFQ8x5XOnDBHqFmo2X8HBKy+JC9o/nVK/MLwhLQIyNTJza5gKd1
Hu751xtE34lBTOWKcV6rGW0Asr4obmniVbLqQeW8BvfvzzHzvs4zkB0JKf5kQCGY0uj7OkFP7ZRz
vAg2GzqxtgmO6W7v56cj44h/zmGdCgl4D8GtM9d8iqpGHkwm7ZXgQafXcmT1S7aYQ2a8aoE8NPm9
2SthsV9T2TjgWytjaD6vLmYufaWgQsvAzqOTol85kEALqCemCO9TNTDd9VZPas9te4ojSpBw8wjm
tFN0GRKP28YY4LAN+9bdzCFZioKBQoYP1RSMa2LajXczPmx4EZjABDAUtl8A8MvaYzy4T2RKg9MA
0iAB3efnbN2b2h27w9RpAjWdCnKzvPVvXyc6g89h1hEm7vHr449xxkUcWUNjY6sz0hjbk8Wl1bW0
e8kN6JAmocGWNjs1HX1gIYrYlqTDzEXjUuNCL0bGcY9NZR/pZ1PlhYI7UprboyUtOjrHihXAJ6U1
/+61Tl2CTGLekr5Wssb7wwo8C47Zeo9WlBNZo+ThCx5Ay3LqYugbapz5LUrYIzCW08Iyx1CV1NDx
1AmnG+SN8ZtWMKy1GbGyzVeAqkxPub7TPjdlRsepmTt1FVkMEPJ6+x2yWi5HkZD9FTG/5o6E2umh
BlnhYdZ90T7LOOsKA9PcoHrxWWN1w7mmyDbuuK/nqnf+uUUERV8gdKsLqAMXubKcI56s2Ky/BDM5
WgSGHFPep1ePydx5+X4P2Z10z2nGg0H3DI8oondBUjtUVija2Wh1Dd96QQoH10R5TMDNxfUg8C4Y
RTFVsSmH7JgFUOqdXhpucFZIwWJcqsZVBlfjwy7Ba6SObNRbNRY6gk0aGEeX+dSWo/njm0CrRHiz
SV5G/J23ERu4Jsbk8Ca4/od/03AqvHY/AKwbpzwMtKg0cRdccsAOHTxbN6xn3zj8XeJlDb4Egiw+
KYWodEeDiiQVdeCe7h4vLrRMhRDNaRtmqvTk+31wR7MZF6m/wi9ZR/2+21z7AV4g5j+iMTdQabIN
NdfknR/a8lVfaiBu2WtCQ485BBrovzYMWTX7E/nwRhNjuDFxyeF/Fj8+PDMpLwdOuXRfzIwDb/pd
2PA4B5ywxZ6PyTsBnfS7vk7yeB9LAtn5jM9igtJ7UGui998Q0dxe/6RZBcvvPUcMxlVB/df8XDAL
+qqCmxitmmCgx3QIfLoJHSMADzekWEqiOWVq3oRnFMF3/2ihkhwGCFZ6SLOeTmf98XnY8U7Uk0sp
9VWrivlwh2EtmrknHrCAVkkjy8fBfDkqK4dFK+1C42ij8Pv/GAkiG9YbzsD5ZJ4rsyL82RnYrzFJ
u5LA3fGHGB15j5zO1mkBf2HN+1vwF1S4C+1Z+AW45LFu0E41gTk/RH9IJ+bZ5XmpXr73egoHJnau
llkaIcmNSHLdN9d9dmrEDTTf2te0IZXmJF7ZJffzcyj4S+5Rb3lMdnOSc+KhETjUFT1ArnRLhzCJ
A0hiWv4yyu5KsujPSAHOmyAed8l1/xduUTXEYSOpkCb0tr8scM8hPEQOFgPw8R+uEHepHK0kOtUU
tGUw2kurZxySuJWxTmuctj7uko8PoZ05aXzKpkh3AoFvkBtwQUeZLerQR/1qwFbJyO/4HWy7NZhS
ah/BKNyqCQY9M9gxx9VIkm3witw0j98eiQfGtX8oBzrLhPM5P0GVaLSmCESBpQWWpwmfnu2M62s9
vyyPk6Mh/Y1Z9a+ejNkrzwm0NhOGyzewsSTwtKa7FBo7FDOCmR1yU9/dIz+/te3b1sWP6NMM9nHJ
LzQBkblXYTAYB1zQz96IvMfzS+fH7wdbotBqYc5f8BSlAeprY5JSDGWxGkVN1OexKoWGU3IFGKGr
iI9dQdkX1CaVg0gBIZDkArVEhRazMw3f5kthZsA4/gkuU+CuB2224zrSWNvjkML+c6UuwlSyKRf4
lNItA/A6DvdyyePppyYCeCbb2NfuvIpA8nIlRz06/sgTBE4Jznu6+9wJoe0wfEpvfJT8pK9IaUCQ
LC1bzfR3TVN7nHE+XFah2I0zCUubfVkP0l66ehRYl+dLSn6qHyxh4fqyH75DUnCNHmXqtwml/Lil
CLylyJBoQoNjOnZGPhx0Ck7hQCc6P9FOmpk0Zec3FL4w93rEYdXw27o2Tt4DMhZiZqrtFOwXxdsi
ALZrjXLVYLIGFL00VD91yeCyeGZqBPNkdvN982S7qaviQIYbjlWti8WxyDq1ylXTUYXbgj927F9A
PMSp/5S4CKOxFQKw5dBjkEJnV8e6RRJyjGL2FMEeZW0SWlhCjA5TWXXRL1i5xrnpV36rjNDO0pcW
G4FICnBGmMu4T5pnqXFWoXRE3+ksxJaQn2//X25XdYisiDqQRCCVsQi0Xokx5jSxIWEmLKL+fXsH
5BpIPMgrWbhkDPPMYtdAPX9pCGabThlF51lQziARtniEZhRDAid/zIgOJbIrM7c+xtzIyIlwOljR
0LfgcpjVgZjAKESRkdxtpPjW7Yplnu+cfHwHvhIZPkU4nevUfGQ8SXzqCJ6L2BbhPLt7ne52PMOl
R+ZYJf/MlmXmck8G0MW+BbT9osRWljVkKaBgUCdYTqpFJRu+f/ANzcGo52wDQfQ03fL9B1WRGLm4
VWVc/y4vSxZG5+CPCYM1WQ7vCuyZ3hQwoAEIJwgBkZVby6fdqQcJV/NXK10qOTltAH+nuVpQb9WM
wKi5jcgr7X3/AYAZMi/ITKJ3EXUN6eq+Qw29UaW8ku/B5gumjCRb7q4Nfm4LaOYSanyD9IHuWQJl
PYrDy+24AuBeM+wlehDlHBZjVGHqvEfA5bugTFc4itH3zjz9Rtvztv/BQzLUCfH5KqJLiA1rnWhV
uDKjo0bjVETAYeXnh9KyLGgff1C5VG9iSFR8DLdye6joEWRaFLXsnXrok2ZnRUnhNOqshdKxo1xu
ZMb/Ar3x/A7m9m/LDBCcODr4UWBd1biHRvbJvWqjncu0d46dQKyuZeAInoByZpIc9m8nfLEEiDMY
iglHxYFQ4iMqCUxceSnPktEMySi/5dxE+kwSBqhZb84XOW3gsYN7L6x8+rNacWJ/5qOYE0KdFxGt
4jg4Ev2ftwtXwqNoOHtX8GHw2gvio/S0PTJCvM4UqKFgWyEd0jdhrqpM3XmCD/4gwMDmHecaPCXQ
XuXZtro5iuZp32ZNssuqfpKLcT+Oi1WOUAX1oGnwIIvEHBalH6ZKSYcTYa9yz3JWtDEQZnhNU24J
U9v1pqKFiy59Gn5OWtLmQwLUIaQpgFu0RPO03cuBtnaIgq1bBhfFgD8frn032BuwCzpKdVb/iqv1
auUv7FWEc/v8g7+zigs5tdl33bJhL6stElZJ8fJgMAI3gisKaJvEZsVA1inIhMZZ1+DrkDRWW1bp
h7k2G3RdvqlX9FtpuzgbEtqndvZTmUtQj0gRjnZ2LG/1vK2HolldSXpR731nZDNiLFmWkR3QSP7G
8tjRXcUeMNgjSPD30kwYVJ1/sk2niSFLyZMEksRFXaz/OQ3uVP0J3c9glYQ+tBzw//ZkhHGjNsdb
en7o6YMa5zjTRuW61ydJWcWkx78d4TbYlzVWcLDSJlGOGHwqc9wz12VK+agC3q+2BGDuZHUNZXnX
SsQWpMnTCgY7pJlYYMguEQdn8v5VPeeEhSjaFamo5J53e9n/e7rOXEtqxrjRSFQX5B4T4aUh3KMB
NQQci3Cre9RD549no3WzAKs2SOEQ2JoLeygbGP+YJCb2IRYbtO2utshLHiGJq3CGKAJFJvSdT5A3
95nQLq0N61aL9uURKeoB4zZ9nntWCtlHiJhUH4TU+HXSl2L2IC+58JVMePcuq1Gq8DWSVZ/ciArm
vJAeiAWAKMaHoaUvbT+8f0+aQS18rItzCGzSOHSDdn5o0DUZb3h6l9rLA+lzxSwZaqdRkUKa/qZJ
b19oJk1KLOATU6IO+p98ylLB8wyWApVOMIbZ2yTiMJPNvYu0vmXUtDBZAOxeCYTs+uAka6j2bCt2
Y8r4oXAqImOVDjIJwvt3igWoHkafUCMSdKeEnKB5EgDaTcH+FQtDOHxJQrLLzFzqHhubF+XR2Myr
70vWgrNQEpIEq/if48vv8uF2iAdX1Z4Mw6gn+cU+eAAYH1Ogy3tKivTdQUXpppvhaVlXes6ECyZW
zZwY0VZfg9a+8ufu0kg1QBfPrJbqrdTBZJFW/sYd02NG22XAMZsK1NW6Y2JdxsZyygH6rA4UTqof
2yx4OdsGTS9NeYYuKbjESo8zT9lyYmHAFB9iAO8rK5YJqWZb3YjpXBR0Tx2a13ijdGYSeHxEl5zk
aFffxHWrhDmpsn4APGGNG5ATDl5e5m1lwiArnpU8DJ/qHMBdVzjT6e0EDtcj8RLXawZDxBVsl1+O
yK5OJ3ICq9PWislGL790G/JjARKtMk7VsON3BwvGwCg8f7csaOlqa/QWSayz1okX3yesUrtJZ0hj
9s4k3qExcp8vIBFkvTo2YbibVADxwZonscHdmukFNuRBnmIF6piFpU9AbU8KpJZye/vJ60zVvLPF
+nT8yyVI5YyBhyk365JCxU5QyHkSkvR2Zmc+pqz4wB8o73aZi6HXPWeUyNcVIB/9n0b2nBXRcTe3
0HUG1megSXOCxK/R8wtBgolSeGkFy0CSU6uZetZgvFDVQUg2MqTLnmdUwEK11wQYdi+wG2dN5xlc
2GeaI3CUfuZeuJ/jufLK4m75BJpnIXp8A95U0dvy0G+rJ19EhGBaiIacXQ2G2wXlqUrA5xLjj+Pf
9rWAoKH/k66YczDxDVU0UldGJnkHxlzng+Q1I7TY9sX9u+OmC593s9zPr3Cb8LZa2ZP6n0bZ/qD/
uN9mQRo0UM8B4fkE5pT/h3TfJFgEFeqdusdWu0cF0S6AnoYYyECcVSO+Zi4dMroUSKypdhJMYC+P
dQQiSZlfnx/4rpVE1CLsYmOFptkmZEYpe0Q2RHvBmlG4h5T+M2O7qP9J74O2+qg20WzWfUfNQ4Jd
Fls+SXKfMMwtGxrxSn1sNxZMwCscUbnzo+ytjIonEtuZFw9ESMGq0u8p/3ZrfSFkSgHT3w59btRH
UsVmNqrGbr01n8113gsGj3mGFCnNt6XNFez5DHFeqPuLbkfSpOMlicwYTbfqhEDBVx9hgYTrxA46
pnKcBdKVmfRP7X+rdQTuLWNQZ/OibG+427AGuTffqXE6Yo7/u34Bvl9xpbNZO4C7cs2dD9yoKn3c
gQX8YwzRfClfUl0SdtUmMvtqkhlHXSgEgF8DnfCHSn4X/0Os6ohj3liFZSy84llZTQwXpARYOdqD
McmAVyJ6sC1ZNRpVVT46y2HXyO3sfedZOEd2zfcD+lRYzwJN7ivx3tdi1EXseDwxPc0BHqd1Wofs
WdFsb9g2IIq27sJnIMkGTO5PD8wVfrFD7cEBdk50rqa/pR6VEVssrYxGQXmagnH91raTlzaWj2qV
ZQ3VpFfPoh6sCllCdV5UUjT8fW23LuubXqZL4fhBVNwpiuqG8w+ohCVjSMpNMNo85BEKtcWevFhb
HHhFqutgAGsnNjntw3/Bk9FpvGUu/hJUdg+SekW3mHPjC+g55ilDWgnIHCHaCXZtS6A5qjiwSYRY
pjudO1XaBEyyOj2lbLvN4EYyx7efrqgXR7hzdgn/K6Nsgh3lN/RAK83rUWP6XutNCtKGkcf8fSAT
vFFEXUkNRM12okshWH5qncJ864zA7oVGB3+9LDIqQ5MS60D8lnIjIRwaBtFGnuzjb9MDr2OX7Xxf
W3FndRqIdc9Aq8wBKPLxt4Pco81ITuI1jM+v4Pz5YEL6a09Cm2aX+DGjBXwLxBXlDftLLZrKkOLk
CyoEY0ac9NlWD86HMWMYh1Hw5U+6EN++yPJat1LlYHglu8FilrcA4R4CNWJ1nBmzT20gaKaPe6wE
QMuINMF6PLK9+prCy2gkUGr4GEUv1Ry0wbuKTVx/usaU8fuyKpu1E01syE5BxSbpKMDuKdiHvLeV
ba/AeiPudrI9OQV4QMqTwtOJdk0gmA5vPIFoK7LR3a4CpxFDvSHLuVVC/9o7l4UzkY3i2ncL5BU8
mNwVg7gUpOJupgWdb4EJCViPJUuSxnjASUEjdMr4lL6WCgWGEaDJpHBNslvwC+43IdcfbOBUf96g
5/6JwCX2fBrv4kToF43o5+eRPT8BTDcNr486A5TZ4zD0mTKv5YfMjrbSCcuFyx80lBjT0coJ0Ln+
78LoOx+CHph7tPkvsmqJADDEp+kwWoUfL37Y4nYb/xuXt76VVyDmM0BBjmKYMyUwPq6bIxMSMTZC
kVD8r8MEmKuaOEVBwDYEqPTNpZa0J3qG7VwOtZzUoymPphotBFGRtkixRLYQGRAXDJswNwPktp8J
ilQKyIm+T3r/Nq1fg7iqjrTbNTG1K+M042GHID1nHmTspRQ24e/76NqUkMk66OQ7wR1FxfojSmf2
TIdIZcnwqTUSif5/vqcoaJYRSc1yAzaF6Ajff1Ol1UputguN7XFfG0zppv6RPPZOvKZQoAIKPxFg
Gu2TB/1P88CYmYgx8XWizF9Wi3wZp8fzkyvvAYPJ22jlj1t6igakDdgNr5JtlYC19a6madTdhJQx
sjUkm0vAg7bt22xSg/3pL2caf5DCVt1vdGofZ7QLiLpnR5oueTu5hlPPB/AX34qY9Slv9X85egiD
io//5G1VuS2T0z4n88FInJfmhcjQ29eM0FQa+RvkBsy89ltP05XOAid8lTNfsaqdHe4rPKyZS3y1
5QQQWITLSvH/mFrMTS4jTRWrgvMEu3MJeQ7CjSBD8hd1rLKP7eAVK/4JXCJIulfh07nNwB6f7gUK
kk8nXMsw+bq2I6X3uhaQ/YdRlcBRIkeSHKAsu//HuueKg8piMOEKX4ZzjuNcfHtQo+vAck7T0e9V
+2i/knR5Vs1zFccOJP2HgvpFH/fKXVXlgq69/L+DZNlaB7sJIPOm78kTnN6OuNDYy0tO2GnIVJrI
Bm6H2L6SiTOI11HT668LOG4HO1yoFHPMfUYmMa7LJRjLXYfDctoQefyRQxAXtT0w+2aNQg7X3v2B
X4Jlrc1AGU4gvqSzrl12pJ4oQ0PA79k9LPEkJwX11NsmKpIPOIV0rAiDSBUSO1O6ZQ5ZgVwFr+Qt
Kb9Rqckr1qkZyquO5YzIdKQLvV0CQk+H2BkW1TYZy9FpZDQSdguUrs/MGj+K3CnEBTkasKraXD2b
1YJjfZAz9zsghHl9xbm7VeOX2rVnBMc2cIvuOHRj9xXeBtr5WsRTILMCoj2RLcOJ8E0CBrns5Hyo
du9CQnCF3Py07uX+quIapXkdoZNb3iVEEt2ahArpHKeEFMRXk/t4ENst2Tc9D8I8YUkNf6g/6GXG
tD5buc16Xbc8VH0vaHa4cpPwK4ujR5ZLNASLdueQ2ydJtqfznXNDXw2+Vc3mKM3p9dQmx0ZH3XTI
maxVx/5z6j9Zg6lwYTPvKnpSvkZx5UPhwZI0FVGodJVIYQqKNFwFdrg8wbLv1CW/6QgGKJcSRze2
tXIoevfykSsYNrPZrtmg6tLRrFQJRurAwyLtSPNfQnlhNewUjMwY6O1V5dBe4c65eachksy+V34g
UArCZaHMAGvdc4Of4vEKKR6gc6ONpdebQVbNac/CF/84qjCQsO/UIHeiwOa4znS4TceGtiUpsSNU
j+AEvdZbGY/xAkVTghsePhe5ddFrWzrjLTxzoS84qKb8R/5Z3N342QgCV26JoQhtZBko6XGKlBAp
UAXKVhLu+LcKZDmKCZuvHyiK7QpOx5RW0QEPfEctf4XLGdcHQ4rNLiIovdj+t9uZEXuqUPhQkKc1
4+8Rw/dzXpSiE18ejg6C5PSrTGElp8qiabFx8t70vwam5+QYhtkanHVyikaMTG8CyjOpC8gwLS0E
kehOY2zuompJ4yQG8eRddjWhKbbwa3rHdmY+Le06a2ivJ5uqUT+EP8cyL4C8O/giDboEm+X6m9qr
y99eGxsxWrYt5V3c/HNDBmwi1XwQu0Y/aSOSnbmNNuOm1mQZo4nxGPtQgTMiMFoeR/FYd6oOiLrx
SvxyTwjxK2xSbAgsEnDHASt8fakXEhVp82jkwFHItWq9LfvQzYNgVfsoGxiqaz5BWsIOCesjh8L/
b8xKcFe5RRLdWBfNLKjmHlJEZ3jFsmggbyLVF5L6wBnaWaalRmltgiZ3jRVpMrZBVCNzg2mwgu0u
s9SeKxfxpTkem/xX896iu8e3QugJ0Hc/IM2F6OtKkbK+X2IeZtHEejKwTy14Bcr5mPO6RNqif7uM
xG766nEIHzpEYQnyRXocVexLFqyOjdjePKIt3uokieHAtyWjYlRZ6NWjRBhO+Q4h6ZnMtwu4EE7f
7r7ysdyNn3CDGdoBAP+1AYBnyR+5UElDIbAeiA23Rk8l2b7gAV/oltJcmjTGuMIOKzs+5gpd+CM6
6JoYVWBiRDl28rFzBZFNOW1tq9bPgQgSTbIqGV7Y6AJAxOdK7vujLyTBblK5FMEsqknB+LRULzYW
OYDwUYXMGazOuRmehVeQ/oJLUg8d/7eAcrf8Oyp3UtGhl7SNJZX4FeH+F/dQeItj4jo0pCQ45bhJ
9PQJ6WlvIo32ro8lGSMr11J0vjhzU475dSrlUXtuc6ryJammale6BuYIqH2/2ezy1mn9uLd2vPcH
dETEH3zxVZBD7KvauyOnR0i9jNV3EbB4VM/fkda2oQvr2AglGxhd8ErouMMfxq35OU/zrCCYF1+9
MZyqcGgLk4rwoho9l+JMbnumBoyAVeGuyzYWBFLfdbkSnBKLdCVv+0K627Ie0vmbO5s4ML9zSa2F
pbW+KuIJjIqHOqKG843frBg1ll/aX8hk0SLKZDUuI5fkOy+eNtUWYWp8m9SyiN2Wvuqo1AoJjgy9
Gmg42dRK1fVZXBC6JtGJ//03O0ELISoUHwkiF8LkreuFZlJgPNuiWmYorv2RLfTkFU1RFDZeOa/5
Y/ZM3vK59cBa2w671ShDAVNsTPOZ4P1m8JwyZKheH+ZbRtnH4oerTUtNX8Wwdw5qV+xo2dvcHq82
5ek1N49FWVfQ45gLnuu5Nc9wkBLmlBUPfmU9ywBtYz5lZA4rrLbu++dTcwtCCOUaOWIVJh2US9yi
m8SZX4Xb3AKp8QACCRhd37OuVfq0o54e3ZEJVTDlRavcjO8AtYK/UfwdrarC9n+m9LmfUsD+V6p7
LwyDWf9M8Jll+6LNQ7IbgYwhmfX3EtWg0os7QYkqa4PBQHTXcShfNQ2LDyCUDlgwfKJ82UTbKIB1
H3h4ZuiAOYZnyhBiljClWau1zl1H5GT3Uu8TdoU2eDuA3ZvDoVzXFc2+ALR2rwUuiaVBK/pxvHts
/2f10XffIoKnOV5ym8wttn7qcD9Mqxm11yjbv4WnHs4PZDCOxH4TiRjJhrAD1YPyNgSpBs7V9xkz
Nxrum3Jg5yKpxuGeiPRuZnIe3PwjiGCNtUYlx+hnN7cXPbhteIaxC9f/aTlDpXgLAso+FYmcTDI6
SkUVFIdGZnbYCMMOlVfdBTIhb8hG9NGFAKXDF53oGPyaT1lF0Kge0lPaPGexz0yIElOf3jkeAW9+
43ynJJtlPoJ0u/Bo17AMh0znJXsk7aSWxe4Aono7fLy9hLOPyVLp4OlTeowaj6aD03q1S9cSFxxw
3gig9l0yjliZ+PwU5wpR63u3vYC0noJCrpnQ279KxfiUcS11UXD7jjJIhOAGyP5J55flGASzmRYF
4yEw50ag04GfxXlIS2eRbWXojp3kFoKItWn3kXHlTXk1BnvDVCXatCttv0BTLOzuIVg7CKlSA2C0
hZuI8FkBedvtLl6nwPiKG6g7DR4lIN6VlSXvf5z1TCwyOsiZBqbzgDj3zVKAHcN6BrajVWSgYjto
373+yafcOWvLqkMUEvcSnVLZ28fuMraCn4bBTyaiJ7Nc1zbViLwFmdzJu6g9OltucVY38EGoY6Ug
pDy9nyPr9WWfuVsW+yLIc4NXqpy1gpxixA3brhgUEEe9JX8svTYwhw/JIdgj+XBUxWk1GHDxHOLI
uDu6fN5BK+65yMFrBhJ02zodGA4dg9fkstQgVdfMqztFDAZ+fH5JtsdjuBwvWCp+6vuliHwVs9Cs
/veKVoqJKajRfp3nVrOOZfoJeouk1rTQkwLQWi1ZDaNwlEBKZ7US6iPinIQ89ZIXYcuVDC5MrghM
n0MwAXJNwYF28LiAWNcXwXbKO1El3dOhAz8dswCUu9UOqqEUHHdVUtinlyIuzmxDrQo8r7PECZ7W
UEvRZl+rrgPpiWVuKdvh45ZIpo5v/YJMKlRx1U604Vr+bOscoPiHg/IBA7ekIXKRWFPLYlVB1s0R
sxUYdJBVFujDrdqhdhmK1BNoX3N+KDlzhJ28d/4FAgUfUxREBveqNzFzW18n6zKCovsDE7xlA6sJ
gKhHj+xX88vCJcU9i/cfglv7cPPbUvpJ6HYCK+dNrw0S3frW9TK/nznC5iO/S8HYC6pF421QlOqK
Y06DoLb3NqGuDwnXTgAT2VBC0iXKJ75nteSoRJUnb/KwZNoBR2IR1LlZeUdUWRaMk7lG3Oui1y7y
YXJ45d9LXWOhMaq1o4H6Mc51jPIxq2uN4UEDj7mvKhZUBACdATIMeld3xLI7+lao4mOh6T6bZuaD
u4f4BX2EiwtMISuSUOQoDEN/xEh620ZsUbwleBnXRd1p/0ouoKzpsZbdE8dyTnPzQNHyfX6gNpBe
GzRlxNF4wvgennlQNabziPwPzxvebaC2RWLy4EG+WX6mJ5TeunNvjoZuPRXi3IXq1c/dmlG1G/vX
CUDDhldwz8OVBVTjJzGfINAksyB2GSZl4NBM4EZWKlfIGXagP4YyJXLY6VbhLEsgho8aiorCs0uK
y+Wb6yNFQa+pOkk/ueSJxh7xS7UZCdgwxJqQrrb9Pcti8c807Ypqb+Oa4mlUplqQFQA9gihYt37j
nsh9NJ5l2zCERBZRg40Kd3VRM7mDDZmsj1Gc9km+RcHCe2wSW/e+Yn1X/Fyo3Gaym23YP+La8gRY
vosIhndV0AKchXMaW8ZsOVdM0RpR686ON6RkpXs51fv44rdkzQl9UxlERF3qCHC9bpt3lChnvLNG
YFvk++f9MKF4euUw+PTNBtfr6PRobEvfKkXCL8ttZG+CxemieAqT84HyEkc0UUApdG+EMdlIyC9U
V2u/oUS5k3DL337aJrjaPO5V6YxZqdcxpG3OOalQeJwi0bQ2siofSGNvngmpOIbv7zUKVnS8mKnS
4CHdQQtBNftXNtQTPJwCADwrYIHx08dTbq4RcFcmshJ/MYBcFBkqojB6idhGIhLfxEO3y9AvxSfo
JtLvKla+dT432/wUxv/mfA7CWuL63r6eHAod3ttnPcTwnz0nao/vvj88DSBVb786Khx3fNmub5Qc
G7gs65Gs3a4jAanwCW5zYYIS3i153wFRqyYgzV96znwAjSvgrmN41nGJQS+PrviPi3U9iTdxOdfX
Zhc+n/35U5ftvLjPVYEErUpsEWoNsaimtkD9SvrmRVzXiM3LXgcI9Q98wzVy0k2H7FtlJXGuzE/h
yjZ8f8Y5Xsp/395EmLrNlsrWWq8uPg2U9X/FKAo31wbTz2oEco1g6rbkCmuk0JboVjFAu7ynW352
FnwZgYpU9sk+McYA2Eh3xbcNcB5bYDf2r4tI6Yl6aQYnHKNTTfWwUL9qSMYrpM7bXcsb3ZFinf5U
gnIstOoHZRCjoRouL6fw0PWGZxduNX3FP9xE7+dyFM2ci7OaSxAHKsE+trKX8bwQqQ0AAHd72KlF
5pUUweXiYGIoysHcH3GUuAIGNpVFFQCWiEU0pgwiC2hiRDNijPpHPd9i4/9rdJEVgm17/9yM/HFx
LnuyLw0YOQb/ralUD/WzzSdJSWUkRqNnQWOW7YQQfvHyTi8Jy2+7pEPvW5eYpJ/+ke340saZwysr
iNV52nHE1ptw48gjv1wmA3CtBQT0wsDPUK3Aqx8/C+lbTvpGaHlpGEV9EuIi/hSfgJL74CNF0oqk
HJU/vYQ7qJUAZ9zxndpiZIn04PTdjljeIh6oIpkBb0sJTCKPZhpr1JizRZ0LlPbDAzTWsIBbTuMv
L2xTbxOa3uuZ9aq97lCot5LdL39nq8aLsJ8OWtleytjg5pJZBmdaX4F6PwoIr7gLAg35rnhTk2BW
dJnUSJZ//p16ONtiQnKxtPDZbadHBhiyrsONkOsJWs1VdFUcAJxDbuXu1sN/1sVYjIBb6m6pwv3Y
8jnxykSgPnaFAIjzp8tJ18wsF6RjcMfMRKFHnBHcgem3D3K8gqzMuXeNkBsQYcFKZtqOhBaJZ7LW
tqVe0cdEHk8eTlinJNIu+KTl+ghZF3ILrsKUEbTTtT1oNNHNEW7lFO6lmU9Hy9iZL1UkqH0a0cEf
NdIn31VXtw6GUBVxzgioxjTHYSWP/Pr/FTls8e1z0/awBtz8eTn9CcucZ7DRONzwtAmfMNCFiE7q
M/eTtLQd/tGfQ4zyg7HTWedDqeAghgEHZSOE+dVh01WQiYtplciBgKCYsXBlwZphJ8th8gy5llW4
1p6xc6w2QOrXEv8n6seDdYuubLwZHZx1boq/ZMeb1bEPumSM2mjBItcKkuggCDMBq4n2DL1LeyDp
YizfyZy+uDDjdOgFWdHzhhYPzdmxRTBdvNvGcXBSbLiUk8ldrEkZg9P6E8gmHYD7QFd65jQwUAok
JK1GtViOAGq78U4I1Yc6EmpxFzPFlfZIPDOx8fl2m2+8fINpW9gO7/eP/5UywST4TGsvAxUMJuyR
lVE600Abltp36t/4TnbFNZorUGxvGZyzHAM6gKduOP29ibH7mLSSXhOXOBTRQ6npAopLJl3x5eDl
qr/L/SqMLvfyx0V9PbSVjVnlzjVHOYYNhgZPUADUuKh4UnbSphHtkrYQV5v7Uwpb+CXc0VXjTOur
AOjS1LP8RRKCMQnDuVWenZTiB4Ype3yMo5BBR0KsEvV54B4gDQH1KmQn0eGcCVl102BX6Iz/z9RP
h2pzvt5uM4Rqbsx6D9y5SNBe2kliDg8MxjC5jTX4/uHHY3ZScRa/6It0WSgGrJg9m8gdzfJw41Oq
Sf+KZBY1jiTdqWW908Ser7mYIgSYF94iEgGI2JxVBDp+1CecaggQyHU5isXo4Kmw6UcwZfI6XX4E
t2F3eKibp1DqR5Y5HcIPpJJDd7cmhVV0m7wvRDmrFU4cJTeIADiTvkMUkmw0X4Lr2yMPddU2g/xJ
GezQYxVWWRQHSlDmqsLREsGzP0QYUcX/iz7rXHE732A5P9VQuEdMpYdGmV/od7VHgMXVBu/f+svV
eA4BYGxWoyv9hkpXXS8YziM5/I/rokS62myyI74za2troB5i+XBMH+216z10JDntCU8AIEmh+c84
nsnxaVJJ/GELFgF4NP/wgJb1OxBLX8OlHPNZDz7lHS9FMiGjs2EFN47jJvZu+G8sPN/gN1Ph7jN1
DNHgMwYlWLYnF1PRsRpWQzFNqiD6QiKBNaE65j5PRJ+we0zh1ePImur5gSRVbMSlDJvT7sx4YcBw
skG9r+KXYksvbJuz2BApRddqeQesqocOU7cuZEZcb5HwvdtvoFykY48K87wrUBb3LdywtivotRmf
2fj444MclgU7nCSootsgv7X9HMHhUmWBG9mvXzLypIkHGTpbh9/NRVBFn/8lHrGi68eRpRs3sSHj
vjeNaq3HWgh60dxwp5+fdjlSzD6CkuKHuzRcipBWkq/oVI41sZDSNKXk2ZRnmJzMZBVZJcP3gB3Z
y1I0L5QrAhg/ogfRoorWdFYb1MpBN1NB1BE6z9dRDShAqrv65sEqXGS45IA0WjSjl3qcqPZG5jNL
GQRRbZsVa5XS5s5ZSP0CQSG3+/KVZaHwL2qvC7e8+4d0sul3gj0Lr74wPYx3vV9kcYG6cMRapUQQ
KRItId/2RZH+nTNu22TcpiefPOIbOj2Ya3f+wP97K8zVxGn+eS+Q4wR4FsjKQhqQkZWPzcAhsgyj
5HCyJX8gvKt+Nv3FE156C6TkhHEEnz04L5KdM/JnNJYFaDMkJyliMSrQIvbxezCXgBwy1LfFZGTy
1CmeZdQQiLSne9w82K370SOrM8yYGui6apBNUcx/HBmwFpv3XH5js3wWTMy4q4ptrHjuxft73Ipu
MpuAUKKg42FWL4JSh6gMiAYvqwv3hOpkNMFQnIRyolbJKTwtljwasBzbbZqhYj4diHhKcDRpi3AZ
rdBKYhMipGAsXZIcpLdtZESg5kt+7CH3zMwLsHXgHO0v6mHRJ846vfCAhu0ednJ3TgikTIi3149g
tjUeIgdLwskBff+usviYCY6jOgX0h9lxxQsp77s1wbiGS36YQ2gCRz8zynhi3OHXIlwS+dkJGew9
k6nqbkvScq1EGMb0x3d+U/a01JqGBuMbTE+fguKTbv7hYQON5Kj6HX06Oh1YolxuugbjRkzWTg2K
khKXy5N8RnUOTbb/E338T4VF8FUQWX/pPEKimv+i3nCH5S6/GmCgIO0eiXHOpLeLrQl8KCtqy3B2
N7JxOQajyLaKPS4N34pkgEF912MXiC80rjhX2knkcMUiVjK74fXjMRMYgDQIyWBZNbexw3tM+g9z
8wGi1yn7soHCG2DRJR7xwHKWeykm0OUfelDJIRV4CiF/iaf9uCursb6ZQld6+Ggf97vqQudbOcrE
BMYdutOR/Nbqa7M58Bot9ESAIspfvxe/aj8hN0tfqMu+pAbCECB23/NcpPtmn8kBmiOXBosDKPwN
GywUjWqteAt2ikVVlLBCLiVlPVg9lh2iXmjVoReNoADadzWQfqcAQQwPC1vD3q9VisdXirESY3Av
aOJ2Yix1b6/6x+Ojf2ntG9wteejnhsIOcVUPpj0o5+LjkeTYdQd5SGRXYNWAG5cmWFl5qBmmjDBE
DjbNQG2NcmpFjCqyBgkngw7vlboktpzLTTe2CC5am1FZfpc7Nd16PzUz06EqhImQ6twEaa3u8USv
Y4gWonPfsZgFZEIvPCLMeW0umHdtnDBK3+ALG/Tr2kaCntxhMaT8q6ke7hk9o0HbcR5WpCOajvdT
kqcMZ5Yd6ztPF5j/oF+addxHxDdg6IcyG3zkbkiuBpKgp/dAkXsdZNbI0qRJEnXPAlefV6Xezo5A
Q444RmtfcrexEFUomHFPhUUSKEdef3AhvlmC/J0fDhu0QQmJExtD3eLDpdRkoBX/qowbJ5r7ZOwo
3R20Lb399xsk5KxKzlNchJjz6tgfF7C5IfJwVyPolwcKa3JEPwvE1tBU1GSH/PO2SfbK9sdRWXcA
UaeoXYUlymbMiNiHjHtm6VcWysM/Ex39qwUA4ZAMw3ZL6r9KJ1vhpYyBlKNd7R4LLRCQNjRkDXYZ
KoBziqYYxR+SbSm+VM9BujhhKWwkpxSKJCOLbOzwB+7jdsXMpshf42RwwLK/12pE71iSwZM9kgXm
MTakB+051YqCM/AepZ9iSu1f0vU2kXxaiMwkXUhn9uU9cWMsOg5V3cH3BjcbbOwjcAbU94CmPouw
oBPa/cWYyVDizea358rRccIc4wA7UbnvitBpTjeYaRE2Nxa2AYJHC1n9cLps0LCr1fNHMpNNdiaZ
V/rcYp3T/916h9VX9EWtRN6y3y/s18aVn6k6aN3tsXuQzaD/Ok5VWWBAWLCR8qUdFFIqgpdxft5Q
+F8MySovnnWvV1JE9bsYpeNopKramnfSeQsnNanlD+2o7ZpsWFo0qjgayXdYcaBqRHitkgeiB+FN
rfiX46mwqV1qsHPzf7WEyKZbPNbmg5asQ+O05xN7HO5+heXqOev8zU+qjHkGwRpj9ShOu2OJqcZa
iKaHFUjQ+hFgkOzubpJUoqoy/UeCmSvRGLcFC2xUS57S6lhCjJjzxclSQ2JJh7cpQXP3XOoYVryp
mCbIRPKj67acbZj74VQenKK1ULFs60w54nfKH1qL33LvbirUcCI/3fHhJji2NNlyyc9jkZWGve1q
yjJjfIcvTIpI0W8aqxBiUprq6PkIXC/SFxYEzv04WZZZwIkw4JB6zzMRYQnZ+CtEQzPX5lx54TJr
dWXNCQ00uoX1Ymcqiqs8iG914hLPDcCZ6yZ3VXPndL94uisgdmg7ovjPmMRjjXv1GeYex4CcIhjQ
Qppr2k2np3v7hpuycKt8fRD1XNbTaYwlQOrAMy6V8f+mkzwNCHpqOpN0mdc6vySzyugKuxb3yoct
SRP49F0kJmekwum7R+5ovWAQmhtG7phqV/P/T9Y2QMhEE2dug5JS5GnP8XTmQnB+tbChxWs0g7CG
MuYZnwfxKXV9zVj8deXrZuEeZbCQzNGKpmh73nZed+W9HeLgFnBLIzxgHMjxvJ1RChP8/Um3ynLj
H7wkyuYDmRvOfj053MvZrLO/pXPnpokbPbSSk0Fgdhx5bIqVtZ6Wlz03sXDEm5Uou3ms717W77FB
vt617Y3ThPAw7qzQF25ZFxROkVviZLm4dcqCdgCIDH6QxaXqyF+nR1Zyms/A8SHsn91UgaxarL3k
YtYlYsvXwMP5Tulezgdd9ui9RT8x/yMOje4Ke6lecekGjpiWvcNLOGgm7eWSwD5dXZHqmyWFx9pz
Ir6uGoAZD6PB4x9z5hIEoKTNSyGxn7wjEwFmYdrrgDL6V1StJsQE892QYi4FoLjzmFQJs7L5r9UG
U1esT3SayoSY8patqQYCbE9iSiw+hcFWQrAnuYCFz7nLP6HhWp+/Lw8IxEKtgZLPjX2RxlSs/WUf
6OkQo5PoopyquTBG26IwR6+G43rrtovWbeu2EyK+K5LYgvrj71Z8yQqnWbopiMdy/XU8FCMOHxIP
rpgm6UqiTUlPvjCvAdv3Z1IXmp+8fJgz2onI8Yuuu7Pm+xNoQ2rZFsz2uuYD/+gkXUr5uUBRS0IQ
ak4Wr/3b/+E2XTfiG2il1/pC0o3pkwQtfKUt/0hNvbQPPVaMcEi58CsBcts1yCpm37m/K1GWl06S
iWbhRkXwSAUgM/2U00ARi7lYkaxdl8UrG/xQdfLJ9C2O+8Wi3wH083p1f/1dY8TwpsibwiG2ZsUe
t68SnNSEbYaQ7QT/UoNtDW1tPZzzRol/KDCAgcHmZEP6UwCZlgySOBr7s4MNNhHkbOSMFxGvcZjz
zb+ivoRCFX32hWtNImYKX+oOoQq+jTsMr5owHyp0uEzgpXWYMTg2bIsbGRQfOha8GL2M6cXAnrwp
fzww1hRCHge+NuuEzVKXDzcNNgWccSGenML/mFlihy0mGhsk00E2sMYxfwc534IJUCY8ap0KMeJE
27OQzOkHQZlIVSjSRs6SeyaoMOu5R8oh+0zgn+lXCjj//fXXpJLncwtL6xSnsItvFL/W+9bQhp2O
7vsY+bAxblWtmCody/k8K5VleDijp1g/ldWFXuHLcWRd6uBSG882udHkH5W6RsA502K8gpG8wVuG
5eJ8Abmz73eJ8zxssFM+2aGG+K6uFEBY4r1Pb2p/04xO/Tn+bqnlqpdr0nnfJrB0HTYlhgvmbtAW
q2S2EpkjPwZ0xlJs1Q1R5DKxFcltUE2waB04aVL8pnF1HaNyQMaB5MhmExdccPOO7qA21yFSsvYL
A568REKtmAm1Mhaof/2dgYX2KkOB44RAFELB0dyJoDfKNTuhKsaZ0W3zBlPabRd4Jq+zeCx2Dhia
tm+/i+9eYFKjEJc36dDkO+ACLQNo8DXmR4NeHylbFlPqVf3YnMkIprd/C6sejJsVlRDgumakIntR
3nXP+xlyYmMVnOmbOa6y2nplPjolkz+U/T7MjyNb48uZgFVNqxBfLA5/A+kSw94Bm9qwaDI1LQbZ
INDcBa1iIrSSqTbhN7hZ2qTeOb5EA60RFCj+VTSK1V9L6tGJb0w9t6l2AvVQDGe+ZTJdwF8AniX7
uSnfOdNorh8VyDvYkaexuN8bcJJcqV6hPicNn5mIGj0OzwR9fx/Dntw+2g4Jo3S0trdBLX/pNnur
0H0Pa/lvt+MUiK6MF7kkf9st9CQNzQ5w7brWoL2Zs9A06h1R5hqXf07kHAWosnfj75xbWTFnXvnQ
x2a7IferS3K6hSSPwEUgEPfPkMLLgerQCzjZ+rYzVfXZ0a4GpTKouXS3vlmsPVWiK8H3920k2tX+
tqO18CDYGh+07lwSu1IovCaJc983byaH8pXtXt2SonhiKSWWt7EG0zMnJeJ/aodCd9S5fABrxOrE
zInDb867dSi6nMo0CJnq2FdasRdsl3yFn2NQxhxXtdnw0Y5BzN5N8qivy7TgIf2Spwn7ZDov4eoa
UdkGeKjFrRZaBJyPO0dOkHyYynYdaYpHQI/fhejUBPnYwBhEXK5Ha2ENhLvD/R4/yxMMW8+9vnh4
BH3SkR2Y1MK/BEagpr+PDn66/JOYMcKrX8HJS3DHyVAskXhuSIJ9Cjk8NngLDR8uiK19lG1DDFE4
MUOKnBQxfMOKFty1uxaHM161o9fPIRMAdxSNuo8m8tbcPHBuCTBaWpTLXF7xJwQbOJgH63g0RlTJ
uRJHoibUoBPP+uN+S7YJR0CK5RjVMy+qt9DqqCBff9zEvXkOakmUAJBpkNz/65SVQ3COr4UJyyQo
EaEwxWM7V0Gs4Q+s7/KyCUk7DSawpvEUUTzavYiRer8DLqWldCavNrJ18JnGo/39mu3AVsUUhNxJ
SpSfyN0gb6OEOVH4BSeSL2eNSPgKQs9JNMeZjD34PZ1nZ7iGxBT8PTPzQZldcZCba9WHhFg0+8f0
ZPugCsflPNqep60/GG2Sbbq7wW0eWrl7fOmKqUf1wFb5Le2DKjwU9JeC32L7yS1YCqmjXKt5YPyS
nBiit0IRw6/eqtZakF4Eg4o6FBDE14KwwQxKmdUoKy+r/3oYYfQ/VwmTOGD8RlrITyzuQ6qOtvLw
Y3STEf6mtkTsTQqyKW6OurRiOWY+0rwK+wpFCTkC8E54Mvzu9rQrRLAUlHPFw26y17/FuGy7eSFM
Y9nkCeINK6yiu6YgrgFKw47Gq+fgddVF0E0NgiIK36nXF2Nbveac6b5RUPFomWclPomY2ZlNe3P4
VBoAK7FvN3pdpL4E1S035q5+Wyho1AxjPJomip9VxZZhYPB0gORoZgtluzUYhjxHlVqdGEsSsXLD
m12C6VYdY7qiwyxC5G290r3vKF+ZxSRbOPEqfY2HeAM9zlFIFrJ5c+9JgloFc946X7SIjAMEUSdf
nwxQyBjClmTBX+5SyrGGwy4Eii/b/vugktkMn5ksdc6NARhzJF5xa7TOox9m3D8RwFQaaNgXOayN
bpvFS4oZgHSOgWnOuRK3pAQH/QPLMttvpfVulUKtvIz2fvF+H4F6LVTL8JawmoAL1wGWEaejD6In
u491/oPgAcOEqdRV44z1WHaZrQbjbkSQNlx61c1fCbc0jTwd/A9ManvXhP2gW0pJXrHf3zEeSp8/
6koWLd0oBQz/x71GRFX/wuz+bKpe1AedVaWXtxDKZemB/qtsG9CRJd42gm7372mSyr0VCFTP6Y/Y
m+R75AMI/NbHX9iHMfCE4o+ZUm2oK0oyMhcKf0M83FzcsWjnNxm06tRkhhStZeXKwZnySCoUK0Rp
WcsMP1FolR03LHcG3usbzvc10JmkcSLLsb1U4Y6T5EEfUJ+kUFDXxiKSo2krovcFKWNU3VH6MHf3
QiDmIjfjHoJQS/xEerVU5LOv0aF6jWtx6GrdnlLFTAdbxyWQ5/XhTbUjTQz+5IBV9SjJwTVBvjlB
CInnK4GzVhvF9Iq6wyWMyOKQLw54trtVb42dGDIJFIyQe3FMYydYfOFVzBBotWAjQYCmZ/bKjpRF
ppZPM06Pi2bQXCtnzQG9C0wOrA5Lvn212M4ElEW6TJjfijLT6IH3dKY7TCNU0e1PVAsQ4Yd950s3
3T62cYSZjcpAgKipVXSQBqpi/g9rCmtsyYtJkhigefsfHbqxlwEVO1moHjgHU23rmY0T4ZELBbjY
MpazHZlqRi/auxnj5omDg0lKFIk7Sg+mlpkJFyiHjHBnqdglIaWFTR/OzK0Na2qDALdXu2lwmsgI
tmxRaY5w5PkwcSobRi40xF+lCM+OSR9sETtstx5oBrBS18d0PNpolICeWk6JHatTHaPmCb60S6hU
KE1LTjDd3rrqn9f3cmP6ZPcnRhoe8Rgtym4qFmWe0dPeTlZILPO9I0/IoS7pUKwAlOMLfiBve+a6
bF5iIk8BtSLSbpO1B1jUAsZfJAyhrkK9sdtu4XrWghOWONcKhbOkcwlkjfeKbKkxfFU3VJl0ymFk
HWN3+OM9mjdFUGqE34ym6U/lfwx7SiCjcP23rttGTyLhh1sf5qVr/0RmGa5VpbA5vPB6tvv+DpWZ
3w02SFWgH1PMSkokcH/8LEBfs8+e0XzNaQVpD+zJpmgfBvBjf4Dxp8VI6aRX4csHfjmEu0r1Pg84
rNYWQAjygWHQDu2BEYdzPrOHn+zL+sWg1CdmozzyuyZ/Leo7BK2JFkknjW/5EQO7ALnIPBKoQt6/
byssyvpLGLkSwCPHt17LuJ2z4wGi06dIR3g5WG2qKGs6jEkIBjbUIBRJAdIqaHjJVcswjjDeX9Iu
rZg9YyvMx03Sfvjak9rDhSekifv1JAPk7JcouOU7483NdbCv52/V8r+5rlJ1bAhKSp11KyX0rQDR
Ck2pB796LZIFpVrZcHl1sPlGSeDr2XjxyvB2gjP63gU7QZcSNIctaF3YsIT9q56c+D/DCKYIGfYG
CA+eC/oIVGhHGvelwSIiZkjojDQBw0JoFA34knQaVz5hJo5LKCBTrCGnhNCjbTRRq2AxnVk46qNo
PsOnlntunwnand7aUtc48SyH1ecf0Ec9qGANwOUefA7byjMpZo3xmiZkOvXq0BU1usZt/pCGmfqf
b5jAjRv8ajIkizkTc2V/iWMtpAdse6gxzGw6ECL36GN+3Qg6TtV6g8HX+q25gyF3qCwAH6Fc26xD
ipVo/rvwHjowgliziKSJF9yinyqFym0rdWRmv883w5Fzlqh+FdUYmp7U+b5aLXfo1ylP3prib8I7
X+uLirUezsh9t2AI+uO/Q0+kYP02Equ1da8uwrYwZrgTD4qv8XWHnyAMoTCRzt4pXg5pPF2sgYSg
4H7a+esIiJJ+45FLVk4x4wiwHQVUAbE9bcBnMwcd88HyfO06cpUdTISC3QfrKqusY9QZFfc/myc3
IdUi5zSCqBu/kssMH86MjdCi1TAKV67P+CpD6GywewpWFnYEY86PbaWPCx/wG8AkuNyQ4qFI0wM0
vSStTXqREdIxYKijwjO/THZr5IkP3rO3fFITrSeBJeuaLoreH/2N+LgEIE7tRCUiQEDCNBEbOkK9
0s60NjiFY6zypBYFt0gNaSkJjBx4ZMqMSC9ftc4rzYNXyz3CCL/TZEvkNF66mtqO+0C1Afplp38i
tN3BAyiEOOGiD05/W2yzg86mtb7MOnrTpSwvrpjBCLIyWW4jbTnnETZrHe/i3piBO+twPxYRFZ8X
+YzAxADBM9h9lpaMHACzX97WH1fg9LBHTGNQTd66o9G1uwb0kAoG0ZduyLz6Qwqr+KUkqhLptqdB
ZzcFzGXA27xYfxuw3NjcaYEX23fz4xP/rs2qU+3kS30MLGnlfzBJRLIDIfDXlXJ2VctinZLUkcEX
I/ViGL9rc8VDk5fme3OBXUDwX/y6m3tdSjlhNE21Sb/E/buaO2XBxRqjYNlB31ennhtl4LygLnT6
xAoKhfBpYRY/HH6DDFI0g5G6UAvVga+MvSU7xTMaGYZMmpN15c/O9NA38qkXgxB1Zxizk9S4T4q0
TEhCOu+QmFRE8+elp/Nty4FczXUQUGqoExxlriH3R+bq2OLFjHQiaR/mTUimFY+hJo4jGuoEPnff
pH8EJRA7gx1Hsv5k/MJTDNtonpSHbf/g/GPFRz63nZGKgXar5fUPFDPoJe0WdIyd1qNKSbEt7EPA
fRnGg+1BZpS6dheT6oOY/RA7mE5t2VRhr3IB5AkBrNvX87ehEIwxtv7WIOd6pn1gZPO482Brrb7e
beHi5Rfg12RusuiEL4jjfjMYZ71tHfAf+NpblZwJixTcSv7zCRcD+woqXsun1ZidXFsVTq5CqPZV
BwkQbSBaK8HTJrrcNuTwAp0i9RGKX1EGHjwS4lbLPnxv4CxKCX9xm1BPdUm2xt4jY8SBI5wXAq+R
khI6VueRaVkRBQSIMi8uuWqy7lBZ9jIOHH1IkdeGwKv98UGxuawokng8RvbSOSGRrVL6vw0Zy5K0
11G4oBtsSR6472IM+DXoGB+T2kl/O/pHRIfn3+uzWLoZBftVdgjW8/oOui98APIBSD895Mvr9h+z
q/AK72J+gt+bOByNKjC0dm6ULbRpHD4ezcvoKKH5p8Joil19NDmAS4k9XtJnEUaa9shS0DzYSpXl
8oNLBs4p1bpOU0Kc6Nsg8r7W5buRvYF+gELa7OW9WQ7UVTLnkjsoqY+ILk0mWG2Tbln8EyFMgWWL
gU6FgUzrHs+F8CI4ALLXcDldonQ9+9aMBQ3JVXYMeGpdAGq7FltLDkqiZ8ylGRqfhDI8HnCJTtE8
v0B+TdexGFrOIFdKzuy8F85ICAKkXPVhg1MfVCgDkOjcEUyzH52oxFBpvLlMhqhq3Zux3tLQGSIz
f7gKw0UfJvkOc0qqALeb6mCzkIlVfYVpJfKPprl6CmoPoJ/h4zeL84PLFM+wjeJwqr02fIvmPRrD
Hx9GLPwe8jOjrObpJylgQftRyBYxTnXuKT6XM8GDLuum7lQLVDw+3GL/VU9gCByeGLFb7f7tFPKz
8XS0AldKqSOGRO0FbGDW1Uy7lIM4gO5hGmOS7pEb/5gvXEjN9pC5g4cSxGyZ2FmAdDLPVKKwypgV
3bu7PfIKbj/2jxZ5gDj1dDEltiTd7kT0tIY3RBerVAWCh+PH7BVuoOTHfgJ/CFKijJVRomi+35JP
izN/aR51Z43Rr21xpBw/wxtqMtclmlN9PaNtS7Q0+N1h7rgCe9WPNO0nffdzyvh9H8qSfD9EajF1
NBxV+ei7UH/FVxU2BvL/4nlP8GNsVIz59h9BTUBeK4bv8qLBufH112UdrV3fmMwjKbzHoRQNnW0P
EmORJZ+kQ2H14XZ4YhHAiNWDj5gzy061QmZLZAlZHKge4TFZ6+RK2fRQ6RbVN/60Mp0Z4qwbpZpC
HEBy8xS+DABjt8QpNKjLbu1wi5OhtQIACv3wJsTTEfrG+exr7DR8gwG+Dw85aFhHSdrQm5+ZSzjo
6TCjFQN8BKHMSaEkX2f/7B+eCOtjX2i2AF8JqoSoyV/VBDZPxCkApAADYHpcb8AnJhZfnB60QXto
LkJnrVPRh9sp7NGnqm1DDTRWa6aq+iBO/wqbKFamUR4AQDXRb1+skzRzytnHT+xbKgKUGPspqbBl
SHwPMug6tsbRdqrdyvEoGbuhQgHn87uO0DDNKnO89ThXEytnogLb4ABaqe6W/bacHne0lMeyLJw5
8ByWHgC3qJ/QNRHfiOx77EqTTsJq8otxQDDqbQZ0MvDQNrgPQ3beKyr+555qGpmSa+Hm3X7j3n0X
dDYI3reiF4q41QMaPoiEEUu0/cnv2+LRp+ZU2CbKbFEXegO5tLdb4dK6uStkKrnN9nZsVv+fAVsD
K0ftViFmHxurMpq/SdU8vLsA7VfoisJeCyygchwv0vZWLqX2q0uMCxY4wPt7rWLMBSaQq54hDcPm
f5SCUyPAxoEQWqIG7o7RPuI4ExDOX4MOfFOnyOTrgQXJjAKcmnGYWa0oX0Qbcx15bnKwPG+Z+1xO
0uLFErjoTudfSvmd6hTamQufKcZJOofjOs4I86aK7VYT+yKmeV4fDpjtaIr/Q69mNURx8gjLVjwq
tq6bcTI/lNsNk4ygcbt5oWcvGQyHXk+WN3TtbY3bPi8PvSSK99HicZEmV/51fFBxujPy5U8WyUTm
eWgw59GcQtaNbcoqSC9uJHGdMBaKTI+ynCtJ39KWPRSlB6dz6m6KHew4CvqqB8m815GpV9R6MAWf
yaPka75XulwJbE//Isa2lzEQbpmaDc787XipYLuZgdGRFSYFCO3xSVx1GW5iSPCpJi5wDVcrPzd+
CZHBeCn3mJI0rLaEqWvmPUflGxKJeZ33J+chpteO4CPchJld2Bq34iYY9M7zWUFLIOD/z4en+0po
KQbLPewLCqe3BwiK7s+U/QbIjLmuMPHCfv3oVEFLwNSfKEc89t0jMEZN03mGrEVCHn6UEAd4yUJO
R5/MIzVnjUSPbGg+/UEsG0axJjUBvMQlx6X8a7bxxORQa3VsqmXeztdp4mD6V4hbs1UFhxA2Ih73
nKNLpvpE/E6XlwWWUmbnDkL6Zwji/omT0s8WNO9d8l2QpnAiIaOtEiyobUCGM7gvSOVajA/A2JSE
/EctoO/vVYTcoCTuyoBAOjBx3FMas52x6w1BTPgtYYhZBigKAyvXbYo0/KN/S1m4IuPG7GWCdSoA
tMYQwOSGQzbL9KewLdbvKKbe727qBFAR9sCRNAH4P3usj2sJ5n4pXRzGIc8pqsmfUXvx/CgUKx18
t438DqqQ6M2XvnFbz3h59hy+0yK52oOxaQneckN90V6Iy5qf7ZlG5VzJYLUaTIrH3O4Odi/ncFkX
4wmLCf4NK73FIv1y9VBk17tJ71USz/5SL7NO/dppwxG7/Kpt/hurtlm+9ReFPBX3biVUEje1oVGa
MU0p15n4yINiO1iN/cfKFrWTnWZO7vJbw1hcgI/WV+5nEjn4Ztmyf7rLqT7LZ9nIje3mi3zRJ5Uj
lbpTLdq2AkcKiCavOIgnfV5RbcSqENEmagjE+Q0ZV5ZHMBRColaM+5ex1T8NvMJkuOJ3KQTjyPi4
56VGcz6M2wMnOBEjsdFgGVEKyEVI6tH4/VIoJRKHET/LPDgLrOiJq6vzPsq2EOfsGdV7wEVp/m83
eazeepJDUDC0IsgwYMpd7iN0YycFeP6HDMMQuMRtd26kjdmE3aXM+DgDNTySv0p0mKpaEv67U9aU
qGUbskQsS0QqshRomGKHvmW/uwiimQs7xklrx8uGO6rxAaHUhMwEynPELIFwaR/X/dqkr2G9JY98
E85gli3p2bV60SfeC3slBC8GcAetoUuemXsmk9HUfb+K2Yrm6xKOTC5pAUGLLlR3Ub3luD2F7XHr
OqBsJTFmBCSzxo/qQZK8cobtsH2upTscjv9RfzhJmeozdEHscLnOWA55OZ9lL4KelzI5KRNNUzRM
b5z3FhtQkwPynFgjlrouJ5KCrMCDcb2kgbfrIyCS6BDc5NrIho9f4wHF5XkPk0WURq5aE4bOAPrW
PCEgDv+8FL5zZnMTDZmRyLfluvu/9EBJjmj+yL8V0PFh+t7L0GUURgSfbNpYlZ9kSnI3QN1CWbuD
+cCUTawdlVnpRgA51RGhtZBCvrAv+GdFSkkwS9JjcCZczB+uSv3XQizQJ5uyW0cHfmV1VQnJHUF2
2XHSzcYNOaWnrj1X9UQq8CbQlOOuNh4Ax+LUjZNyDXK9/o0vgi2tz2Kp844KnczIUn43WPsy0vWM
XHTAjFUYHDE8tkE37f9KWXBvIutAG9yjwMX1mZWqcu42bICnAmxwgEp4vjr5pMhEf52gXI80bkAU
R+MCSd3JPiwbf96iq6Gtv1CvPvIWLRuPotRtOWMMWGom/ctUuZlgNG1JfOy5DTJGhFGwCE7fUy00
pXQfYyzGwVyrMe/nbnAfVgNT6Ky3iczpEFYdXNxt9cYClVxK/y3s5fFl+093rKk8eOGcARL2eN8Y
fU/O2Q/Ste69S80oP4/jkcrTF0fpiYTFFgaW7Na/wCmVg8GCYHiKQ/njD026tCXOKiCFU+cBUqGo
CEabeI1PYtXGPjRjP/27oIH6fvIgasd0WINl9W0OJLoVIfcdUJEszF3+TS3+8f7hFg7SjHQaPqVN
EgmtwwXxRPx0ZXKcOgWUknmH0S4gCyxQoy/81B4toFy47R60itQz8vAYbNsArSx7oUXGPilXnjZh
LWtoDaKzgorNY7j6qZpGkFMSOGm3ImAuOibYjmhA4GbaGARd1trP+cEX5K+5LfD+yZEexJ7VC+y/
TXnVjDYI1QAvTnMaY9IEzIeKkfz/SfOT62ffPX6AgRl83rchz8UhiIHoUqwnI+uxMiNt3oxYHxdY
7PBHYgrxaiRaP2JMgyzvvyQlam9MLLTuWUdlfVcbxgpB2SCDevxoceMxDpNJWcaXL0PDX0H9rDK2
BzfxnHyvkdky1MhCD4pWtH+B1vHp4KSjUhIrJ8KiObU2RSdjZEMeiY9VYseX++fwG2MdZztpAyMU
ArJkJcGQjDUhmmGo9Bo12CPc+lxGw9bzRZdrHRrHQTx1x7REWYJ7ZcQleBwjMZi94OoG29C788t6
I3h5Pey9MJNk6EYSxdzt/PZ9/1bjynHy1p1YFS4GB6cqyjLtEq98PqEmpimPUYFCLK/gDjqhEsGX
m8gjtw19SFuPrU5+HdiPG6K+TUhon4+Z+0V72dzEJkoHC3gzF1e8CA4DFb2SjqDj4KunbW5gFMmt
IpyRY8MgCQGrLrq+ahdswZxq8/GxckvskNu9YVGSihRQblzPqyfzGdyUPg6hmPi8tKoBaG9qtkVE
B4PFIQsJ5ggSwlbrgmXCsHpsYA8v+1kXfkAxvfzHxUQWPwsjGsUo5+vwiyw/6fbG8w6m7uzg0HrT
VSJ00ADRCsFr1F/6ySoXeTpgKKxxX6yc/wuSs9bbfpglpT12R0xVCT9XTF3+dV633OFTt3dIPwhs
0DOcjAfpcWjAv/vV5de35/H94BsRSmqFJjh0n54FzIIT3A4L6ec7b9jGCL2DII5o53OXt2BF+yec
4EdBqh+YgpWhxLv1ozrYP1KPABMZ+2rP9mVxoW3emTlZROIT+Nqv6n9OP7VZRBgqu9v1I0SjnhRt
q8sxWhVlQEPRsJC/RR1rpasnOwkrNAaLymvdEMGhV6AziRV1Kd5bZ3odIT2oaXKu/I695d5JFekM
0vyKFD27G1n+FAAZvhQASef8rjciuN7HrfjZO4owIswUDqKnz9UFD0ng3uERzH0vfIKof37Ko/GY
W0vFe9uU5fSQgvbFB9cupa2JGagYarTTSNzfGud6CFC3Q4wmTClRhDNMvsjcruGANNRGVwiOVDlw
SUcQBlHbefWlKme5nUlzh7UhJXfPYlYf2mKKpAmySgxT9NdZSd3176S6e49MNos3UimCkDEA1wFd
Fi9OYttxUKDpg5suDrZ5hu1HUm9aXc/IFSEZn/m5BwWdWRcC4VNdIozq1GX1sG9I+ivvoCq9v8yA
7HF7rbhrK7XonvX5AhVBOdM53Lcia6IF+qUNOuyPZxxtdcmxbBbuXqP97/YlwPKttKC9Z/9sW2fz
fjrmDsTzOS3eeSMiOUNLhE4smlwuDSutlhWrxSeq8YG1Jp+DYIu/mE8AHKXSdb1WvPz4GTeA/iHK
EWDKqrl7HA2HMnFhIq/VWg+tFIRBzxrNwRlN6ZR5EYsVzHnEKbtGVIwId4UyqZb+v6QESyYnOkZP
CVgkhArxp4FVbQZlbq9KqH1xpO8oDg2Bflo4YJ0rSTeJq3tldJKjfhvMon4l7yVM5HzxCMYOySY5
wpnHab1fXNd2AyXz0VPgVdIg+UZqYkNb08cZFifMQJBksCrhYWhlDt1/7Pt0jISLF9JsVpci7HFa
0yW5bAoeaA6Wsu41rUDyHbFcGMYv1d1zoNiXU04/IXnI2kXDD9NMCN5/asCSDOSEFW+w/KX+AxMu
YOgM6RKYEhEqDxEyg6+pgLq+Yoxio4Z9Tfb/yVKLGbllfmHsxaBTYOwJ2tKCfDE+bX3B1qlTYZn6
avB/zc6iLhObzqASoCCZy4DLC22QH3zh6HMc8RHBg3W/LzN6KV8X+0/NTVw55gFH7QhzGH2PSTy0
bNJlXwhpX+SUT7Q7BRA0+1c5N9wUFSXzNCUuV4S6h7aBwD9YnXxbCNLO+6czDIgzPg1FCl6cdPlc
jh3QS4HOWHP2fM9ev3VYbO7YaUpB957aTJGPvkzDVv++tbg7jRANhUWjoXWAkhVsdIODnguG4/3v
ixZUzIagT6Stz4RH+LnRI8WyQUCIHiMjkElllBqDZTNu6pRB76jYYVufiHfwAVFSLQ0nl8M7+HZJ
nWLAT50u9B8w1h9lvn4mRNPlAbvQ/gwbhVNX0Xd7Bqc/LB/amqY8SvYO+ksGW9FdsljklCQg7vts
XNsaS+mlOE7iyCBJhzjLGAxyBYqVrXvUCj7tTjWKIFf/1Y7fo0T7kBr7EpgtX+8Njo6XYmad58f/
F5wrDwc4VTlt/9WMtUilZh7xWGZWTKI3vRghEqc5ev6ldj0z/aHly1Fil7A0Axn6vx+FYBZSOidL
e/C68Oo006KhZ0vAQZgms7M2sL20O755Ey7DSl/a3ZNIN5ffDB0c8IK/gLAnIxsdnpr++3zjvBFV
jUdxRVqSWYqqh9P4pBI0pOihV32ktJo05ufmBlAtc6V/S1oZS0AaYplxAqJzaq6Jm8cGNAgWILFQ
SxNTCd//QmrpK9npzq7v7eHaiJshqmCTpIuWYiGpAkAvk2PXMDGcZAR1zhV+a+hY6TNL3h0hi7Cw
0z+b26WBfYE2WZaAT5gfDFL4UUsCd53OKO6Gq/MeLSIkifPIuQW5Uh+w5NDNh+J+j3wdrRRuh0/7
P8CqI69D5CKKCbPl4BlwzK5fPX5ue5w250CGjn9QgHHBAia/j6JMtwFa7ilUrLPWFiiP6/SHhsQl
b1j7f83sanUijxJ7/lmtSQuTQA04TaIKEmTEspU75FC2YnkGxkWCD1RxWyZKb+RNRRP2xU7qRqgF
f1/+5WGm6+sAv3hr6zgQz57wHuWVQr+uvIGaqOnQcQw520p2matyjU91HhAx0nBlHj2yFSHC0Xrs
oDmazD+sEq/9TI0hXEPBLgmXCE+nxWvngFBb2dyjo3G9kfxhFjM8B5ELk7AUD/Wb+AJzufA6ZzVY
rl7Oe7agRIlsfLxM6T1ZaRrE9coBL4SQCS8yG6TFke3xVcFNecviBRnzmPPZ1kuMq+wV6eFDeoWq
H2Bq4wSvBoNdF2P3qxZZIA9rd9GqD0x1usxQsgyC2vjKD0y0cYETVpylolk7YR8HinReBgOBPnR1
Hzbne6VWMIEIcdA6qXIwZHOvbQS/SxGzmqdoBgMKcX/Qw2HVQYV0cAIbM0l86He4cRsXCbg0PjSi
7IHsSujZzDEJYlyOkOgXbJ1Ca382etv70CLAuHct8lzHkKNu2DwehRZl82tt/i/rDtQRRSJn6XJW
HeMIhyy7gyqua0VUwKeVg5R6yVMkGWMgy/ItOUYhNTrXjU7Nd0R9uziVPGm8G1MtT1kQu+un5X3P
I6A3WciOhdlnjMXr+u3dAMhsQjgzIU7IYudPJ3+kMYfeecRDkfASg2WmyFK1w3And3eIlrG9MuPe
CLCTYXQygsehppI0rUFyOZypwjFy603pOS2ReuCAqWch0Jcty52FbVMlMG7J3VoN9jP4aCLpljWV
SBAIYLFWx+WFGXHLbI50AZ8t0nHUZynHsBc45RsLs2oX4GWSfK3/J4MN69BQTBfFtw+FMmG85Jyt
1c9og4gEJRB0PcbRnK53x18jNSoDCTiRu+0LZYu97uV+AMkVwO3f6IrchFBb2Fy3e/QJ3N7gK9gx
sUOJX+SmXX6lMu3SyltJH0Ajq5zYHqMeLp6RCal5BiTad1HAM/IlBbqIDSudKecnTCf1waMMqhZG
r3wClBYyY3ysuvGdB0jordsuVe43zSQsIuv39PKSsKKqyp/Ncl34UHVgj8Qo46fPNM624rPMufXw
BBdgwDt5DFfoZ78Rc1uBERpyoHfdknB7oHhHzRiJoSiZU1vweNY4YqFvu5W09vzZnOcGrnO/CMYj
Cg8ilAW5ZP/ld9p7JFwxbEZRVQJtcB73NEcj7ACQfmpY1/KYwXlDprAq83lWsCZw+dBE+59tSMTn
BNmaSZr61kThLaSMu4f3UAmK93LKcGVetvJqcx9oJjsl57rEsgjXPQJa7e+yOec0hrUx1EuGA6d2
CgXhZgIlI+occZoyYZy/pmPvSSrZkpFi5pa4z0qZn83RlBxScmmb7HBMmOokwt3Qz9Fc+89pnb/i
8+Tn3hlk3tCU3m3OOgJT38cIPUvsX42kFiqS1HI0XgWi7AGulv3Nnc3VHmSLLhDA+TEN2ThyKUyi
qhh4DR+y0aJmQTllF4tnXPlGl+m8PX3T+JBVRY7OHezdGko/AC9F9wW8D8TaD5DRAd7m0d07aoRq
n1w9WGAsAqHGVbpRzwJs6FYt6UCr8VUe6irnZt8ySsYIBzz+WZvac3OhhvuRXchtrqjbiP/Blnte
VnF/wSyigelYmM+8jXouH1TI4KTzLRm6nozxzi4nXQgrfuh99osDSWPXWdoxcdvrleHtZaioAtWy
ihR9a7bNiZvUZYK8gSMIe3VrTCHf0Ejg2zGjGCe63Uoq7V49wMrQ9qiAkNijUMToXTIyO2/XfEdw
BW3nHVPQnThjzp4YYckHdYGQEXna/4sdU3KdgYUXHD6YUFgxBP8OwUykN3FFTmZqInFR+9VYtiSD
e2WKX9iCZ6lybIKNmkqfZFjUrE6QKjIBLdh6QAtqBTj2AihNBnnK9NwBh3JlNfHxFdO2+TAwvKFF
u0eoAA+Mzo2Sw9AF3cD/6rmLsTb2STkN3Qqoc4cwrj3jBhwAib/Pxj4PK+Y9UB84gf4b8x+P9e0I
W9q5uMBOwbi9vYMC1vSdlZ9VbkTvAKSePaEWMCynWEwEzQTTDhF5XTCTLz7xBCgzTl+R3kp0YIXJ
fKZiflrm+BEC9LswNCPh94erMud7iNML95a0IaHpVTEH0NI7ljZ68il5hDjeRCI0Y1XT0RGeeMeQ
tMxHMdcvjUbnumv5XPnrCEEwuGktgqRIiPe6VvykOhtsI5+iCph3er5JEiLX7VRJFyDIj7zu8bUv
U78jCQm75xOzsTqHxF04xkBYpeOv9qtHXPL/wztTkgDuiqrUxLPTW43uwLztzXxSktCG0mmpze46
8cOLCYmxbH2rprTfxarYDpsfYdEiZElxcLmukrvxS01yNMDDm0wDb5QK5TeTzAOVDSPAbui0JkpI
Ld5FXgxrVDueHv7XW998mttH0I4VWaBYwJJn8CxloryU2qh9sOoCraetlIvSR0RjbuQO2enZ9aSE
opW2A8PH4xNGdYQbxeteBUXlGxGSqOHxP0NwyXrUkeN80oUyCPHFMZX2QfOYNA7yq1hlTVXMcf22
D+pyUHhZmua7g5ahbP6r40g+k8ucgfi4rAXg0rA7vHy0y5KEJiHiT189Ggxn66arwH98Izq/KC+g
KbERa8YhCj6oZA1xbfDOAhIbI/GaUaYyCTvsCCz8rOJg+a+mC8/Clvyj80ohQdZzZT4o0kIMDOz8
w+HJqI+YHxvGsRvLA4DA00+7d6/rh2wzU3cAs1H0ZFoG8di+CGdNIgqVyZDfDaYEJpBLebooNFtQ
UQQvQdHuDwKYj5b7+ijc5S4OWvRdZN/VjEPe8vswBO3Hr26L7p3wU0Uv5aB+DEbisVHUlURXGmpm
nnh0+kzFEOnNvdT0ABzA9HAsZ/cKdfXVlE0K6wZOPsnuOPN7rwWq48ZQ9M1HeFbne28Y9PAyKzF/
7K9cRT92b0LhzV+HYLgh6VwaBdD6oldjChZnPn2EJ/F+3GtL7RPgkBs+w3UiX36HRuU+HhNvQtiP
5QGgpK8hNlqwEJqBBpxGZwp2+wSRC62kjep9vlPNxMiAMK6PL4Y/XhS3nqsWfzCemDkP55Gci1sf
RF2qQiX+DVO2+K1vZg8LdYi4UPuiWOKXmv/RvgkuQCvtWRDUhAx9tihXzm+qaXO/Kf3g28MVmU72
b/s75vHRlHUuHWCFVtQln51QYBVNTKL9GD1uT5Xy5tJKgY82AiRIkYGolYLR9O6zKZvVW8fXaApx
pml288Sb5/o9NfpWMkLsZwaeZvxWNdcYgMRDoizte5A+80EE2BY9bnRfqDQRqjGOgYeyBfhvtd0I
VblijA2cauKHdAP2DtB1nB2x583r76QgiICS35oTuFn7DK5A8xLWBnm8V51Int36zzTZhl0yhSEf
PPicsnqeJ5ozAMn026al0Z62evsWnUhEnmizFdCcM2JGEKz8mtqa9enndQbS6s5jWN9ixkZcy15L
BHO3CPS6ozCM3iH7kFUZH3E6XZRo5tLXs4Io9PEa+n3FV5ctJY+LhPdNZlLM1RbhHcgSfz5OvoEl
8nNaj62CVfUc+CUquQv/RrZttXA7ALeKCmqFehuQtTJ+gQa9kdGUK8tFB36jW+IOqcEM1BdiH8bZ
vxUUqrk0wMmsdmuD/6rsMkri5Wg4EShuD7t/ukkTAT/iNKmGM8UKAtltrCCtGPkGQajKXmbQNPYn
rBjhls4bmtqLlT3yt6g3FTFC2k0/cE3018v7PRDfYfdIznBQBgQq3auYaB2wle5wjO1FfoLVAvec
X6b3Q3dbsZJ7GqMpny/cKndY1wMWLInJiHPDXb1XdIFcGkloq0z5ffuN3/N4QuSAFCBV3k/pFFvV
wypKY7t5oi268uQ8QO34c79wdGRxr8Gy5Ayak+qWYhaBoLatazvJrZnsAkgVc+XEzzm5CgtK9WVj
NI/vupnxvigWrhqxOxM3MNk9gurL0W9RTqhjwE7M93ReT+sx59R7lLXS8JmUx0LcK7fnCFd5e1Eq
SgOGAFmSJTpOjN8yA3wWtDArvHBuk14GkhGFIv3tRzZboAVVZhm5ATUkY5KvATtpJ1VZT4KwhBic
tymt7e+GbHBhqJWJFRq4p6aPUqwIL1HGzsUNaigtCU4w44HjYjhVJrNyaHwOZDTs3kRz7PwPVyQD
phGrnBMQxjnckATfoWb7KmYylVNN5BovrK8B0rv6Q+vLIqVJdbJ0LynpFgHFTPfLvzuEJ7a0GR7O
jbfUYLFVZBNaFy7d5CzIEYU0lSuhK39OpZfIy+yGaNVOWdiMTQf2kPAawYTmM6N1FWfPsmXOmLTp
Spqogap2eig9C3AyHbvX/Km6FfL0wzNWWSyKDgLJS7m+etKVZbD9y3v46o4kcob23Gd2FZmE3RhR
E6r4Wlcdll0hBdH07WptJc9k0SgijE/ZAUOksqBYFGXbe3NBGyFCECs8cQekXVrvAQl20Ov8RfmZ
RdKBuvku4wU6xMIrISAEPYYFftjpZUmgLN8URGVZwQnL9KDn5PA+1pc9iIh0HOeke1kA/8DhvVqa
vCaD4NtNuD4Al91lYUaM5h/EDCDtc/Tt1sXJIBUsn87qlKSxZXZGNJ8AjFx4FF6nEoGkMXyvMZdw
YvzxzXlbIGqTVum1kT4RuQTCSXYT2dUTKjaqld+hwWzgTkfgxsyb6E3vu6JbMNSL42WDInf9Ovu4
XJGzS9X4T06kRA14qmxQPxzcr3pu5MEFKQ7DQzDySkE7ywhQygBBaoo7Gq1kZSLp9SkIqcIMLk/y
o4+1KemC2p54eLV3w5GYzSYXz0P58SwYEC8Jpf6/lrDqLpuNS4cR4tjimAFYu8JVGqcZ8yg0rqxx
QLHxXvgfPoilxgNj6WbMpKSI8Upeupg37510Vg00OKku9wLmF2WPfShflf6YPlhbkyYcVDPaJwfU
ZUeUuq1naE9ZwhozpsWHgmkW+Ah/TIyfhKT4NDCe4A1IpJOnc9PI9rOITZBy2D672K+669QYKsxT
Gzi2GsvxPKGSu7CN3c3wB6SD3roSzwnJk3x7F8KNkPWPWiczhVqbuI1WhZCOXHmJHx7zOXu9qH+S
kii2Q7+YgBz3nHfoZWeYm3Q+PVhXUYQVa1QB3bHQasVhn065kOLioWmpopukKagjcWEpJh6m+kVg
Zcxr+da1VM+sNaRjTZuudFRbJeChosDf+/9im8WRIBZyZYUhUx+7FZVjpbrTWbrbiwL1SkHBn1if
JsKc3Hoy6vN/hF8ZcF0d5JqiSzOMVqbPy0eCIezE4QSw1dJ2pFsAsjL7FDd4YvrOV5Zn5W0LHOFx
WUs8/+Zv4zjn3dUbjx7Ly+AQpA9zxNtHeLQAqa3HDgGxiV8lGXm41EtXAvPsi1Pu9tzu4rDjJQEN
w6at4C0OdVBBMyePb5+gTVIzaEed1N9QvSGm7/iZiqw8tEhNaQ/GAPj8hHgO7aMy3AyU1QeNkNtg
a5/F2NuLOYwNdaRf7EO+C4H1KG0GuDEOupvrq6y4bvs4EDoVj2f+0nwc7l9SSrjsWlUssvJmPyDE
K/feXopw+ouZZJRprzPOczs0yrAK2gNgvQrmsMW9n8JoiOw5wbWVCfjffQWyLdfbreft+74XALkF
kAxRs2M6H5W6MZ/NOsf5WIR/83RGQLTYps84IIGKYqLFxph/EIrabrqNNcxMZmU8k4GX1fNzjY9R
RCNp9xnhNBlfbHdozdhj0uRRVe76geZfdg7nUqemYY2elcUG6N3Sb1xrMLmeUT2iHDIrUBq7Pyij
9AALNP6X7x9cPMSUsOyD4N/mVL53Y6hWTbF2uB24Z+XevAri32kvftUbakEizUrmQhMrcxGbPbZL
ErPQcZ17TEdP9jxz9tZDGUShCpDJBwjHvij8d2ycODgx6ToougbSmh9JlP0JHqGwxWtPnwSu744h
oJTuhUVrLv+bK2pZRyzvskFeb0cuweglrlNIPtlhP9JbKbssdM3BLeaqhlPIn7htelOg3W4qNS1l
qrqHZtYgVDplnoi0mFKqnz1tUb6PXPG9n8cqH4fsixS/J8OSluO0eHnY/TpRUY+XZk1bJ+drT16Z
zh6H1s4/sp/OEy4P69KamQH67xHKDSYiLv5sdoqz/AoEkkqC5l+4VtQPMvmQYotinbkWSqoO+TJU
ZqYq6/J+K5SuqPmpYIpsIfn1Esfx1Gk5eVagzHoodHGW22HRvdmgn6tXOaiGrz4jDU9qFrV+JOk5
6RLoxBFEugd/H5avCS/46UfM4pwkU69IHqaxlCTRtAOixufVWCSqbfrusIUai70bUfFHoEv4ZyCV
W+iaXUU7uEStwJzbvPa116GO2ucsm0RvA8KXDjyIdkWil0ENociKSP9erHAxHLMU88QcDu0OjOwd
upl8cW+/41HK9EkGfNiA2PoH48qADwsc1BnHF8+eocwOeQ9IytfNpTJJJ6xPMA4T16tywjpdEgfQ
IaTeFMmltV2Q4kk6Vx0p+Q9EoZEDIVfWcgERWJT1VuBueOX/IeIVcyfXFeq73DJmPlZR0MPu09Yw
DQzmKzoE4W7j3f6g1EppeoUlq4kqeN2Ja+fLOzvY6GQ23FlNTjPCYBYamBcA6Rj5yiZuj7dYFXJu
2QJ0a75RG8OvVVM9XWlytXD1SGFIIUuifp/lu5DKg+Dnzmjh9puNLqc7hKVqv64Kfw3f5M+xIauz
dA35yzCOv4p1bFDZShX/CwrO9bn5Dpsl6h+Z0h7iaygYD+eWEcmq2n8eKA1t11FGZB1b//A0CdaE
a5FdpMyrbigpSjpTAXGviDltuwKPxouhQlhOrM43muaGWne9TVYJ/aO+n1bHoibl0UxvtvXVpNcf
t9tsi8A17Vg5Nez6V7g9FzjxDEbPwBQOg6U9IN3kP4WK8jkw0O281TvVPDP+NTnpcUTu6ceeZvGS
WR9T+AF0j3wcr89/4IZGc4dyRRLuB4qe42CwKImBRclyL1htIoJ5BP6YGLmR+DUEKlCgw26DIVHE
zvhx0Ihb2Npwtu2NYAF7MK6alNwT2uYckWlQZVbqD0K6GLdB3J9o5ylplBNotQMr9uUflGp5oM+i
h+WOBZbrYVa3VWAyBaBpR6OGgBYhnhcj07lPIph5IYXLPo7cIv+72AE8BKApptlFTAKt/hm7uWgA
GWmMJzd1Y0jYmjEigx8T2gdCvuAtKE5/zM/mA3CIvTvcuAiIOFLItqvKmU9hxOA8M0HNXGYrU7+K
d7vz/3S9mu6Clo9RLz0N75eaaCmoHKOaEb15at3sdVv+f6V69DHGyPU6msaXkuaJ/gMMXvJmzvfn
ymA9h3+x+DgfRg/gUpKcpJ+pRgNRVW88jrn607qlBSX3wvJiHrvuMEiwXhPNl7GnS87DfqkdLRJk
XaY4nrzO5OiVG+UcEOi/dLq4Pj0FifSJj/P164yeWl4WNY8MhBZFCGQ0lVYhcv0IiEREp7jc8Cqm
JQsvNFyGP0bTRSwTpQgvP7FPVySx9k9i0GYabCnZItTaZiixrB0/iriK+8wTu8A8Gz3mqnbr4vYI
ycwT+V2ZtMVbR6XTrWKtOvv/RZX480WeVNK51pZK6J7mBz116LzrmtrfGTSw1EvhTNwq4XEm8uzA
RpZCcPPpAa+qn0iAlmLUP63ciVY0fVeLUm7vBUrK9FJ1lW4PfRaIBnABRLHBbCv0chTGLwI85iFg
OHEuJ1Kx/CzoReVbhixoUrZxcTaFNNawgghTR+eGx7ITze484coqeyZ3qb94M9WMufRJxvet8Khu
8w7KPKza1W6WHCrFwOpy5I1noGllhADbpNQxwKldiJ674CAaQ5qGg2EALeytOwvqOJ18DSOThPAj
o0r370pDmzwY1jHN/YQUu7W4ZhU2aKODoNlo7sK13PmniVvlLPJIYcCusxc9xmOXKTWjhQ/n3ulc
Jvf5DAVctIY0SOsQ9XSvQULCRsKZsnxBvQpr/Lm3pfnetn+qdPXzzjCe4elCHFBmhdANcIfNSPIB
EurF+tGuVvd2lD1mw7E3TUZNe0X9DPxQ0hMAVm2DAnB/0loFPcPRhVkFW0+AxJiGyJzCSqa5DwBS
ICDPddLhpK2571kS+fdFK1zd/0kLF0jzhyE6HhNYay+YB4+3QOjCdMZp2FBEfwQ+ia7+WGS2Up/M
H+6F+qpRUbIN3w66Qv2ZmH7RqejiEuhSSd6ZqU8xbswy8LnPjS8bd0ftkYWk3TBX1uRyW9OePQ/H
vmnUH9jtEuoOLegpRR1S9JuPtCKOFXpatXcZO9BW6+vbPaWSHPvbnezXg2jmyUU5ILsDtlAtjoJl
fGqBO1PPlSUGk/u8Oq8dSx/zomFUk08nhFi3AJO+KvlBMQsGdsInRHP2UjzTxmd3EY3N/LF+hY4f
dh4gUyOavSZoggK/1WHOPjEwqAZIIntw537k9OtWxVPo5iGJ5FTPWefH2wYZ6TjREPHcABRQDs09
B4E04xwRtlCPXdFBtNkj/YbrUI18ad8XXk97akhuGnRrqeakjp4haKRGnvAhBgUjdREZc8WbYaa5
9UaRM5pbTusoRjZtcMiPeL2oVDDWVRAhPPp0TTWUwqirszk4WxF0jtTqfFc4N1g9D6KHGIIxKWyk
Wg6Eop9FpN11S693M1oPqxF/T6oM8hKJnI47O30zIu5E85aiZRVZo/i7GG80IVO+ZQ41SUTbR0K7
rgYZSWPyCgfnvW6bdaa2sVy392Jr6v/4mKKu0eDH2WJVFs3xmeJARgUbvcjs3dcVG5a/lcBMoATg
KERaqEU4IQpgF5WLgFaIXeEHr9kOY/eng8XUbtKYlSAA98kQ0Qf7xMrUvkNaoi8yewgzSL4xdhcu
vj+KbmfMyU9KKhSXjuXsODyhNxl00Ng02H3u/hDa6LOy5ltX7tYG+a3SaM2GhkGBb5HefpzdyTZc
IxXIEMQrekcR821doCilYD+IKlyZVnDjSnDdj9Ud4WQCqaKe3KkfEesXIWwWey93pjM4DyoOlywA
RxhkBIc0YT5NLMvfJMKhBwZZDWQb+7a9Fv5Lm9NZIIyajk6/T6cn27XFyB2R2jdKjkRs+pJhWayA
C90LFMJ1bh7ETbF2i0vY0+9mum9Ocnb7ME8a5yzKmSujgJVeyLXvh1JOUK/pl5rK9RbpFx9MWus6
bQJlI2bSWIjJcFMTaQmm8EKXTkM7OLBnZ98m0zg7xveEvZErnQN9oBex4l5IM0AYz/sK4xiVR9kH
uW2DicvDa6tc6Z+3uFgKrHKKZedrX5FkGv76vTVq6A9M742I4y+dPSFzwcHy3stHRZ2EG/RwIfM/
Iqgy03vbcw84fZkFKBCmPJmBctY9ODVO9qee7cwvPP052C8853D4MWBRiH7KWfLjDIahpXO32Ier
oCQ4aADHl1FBEuDe3Hh+7outtiPVeR6pvLp/T/2WAYZ7NLPgw+tQPt34spWh5DQmuU3dn/AlKw3a
x6mfPXtsLjQ65w93GfdkJYJxdG8nGtuenwFf10KbYSooN2ILKHk9lueRUDyBPYlCmhDKcKapy1WV
O0h6TRbA9620voQbfXQXn74v29vT0wGtIOSbwXLREYfEeYgKWR5X6W4DWBlBhwAKz4QdsXY/BYNw
4JQ05HYiiGB39+vdgDv2p+idRU0gdp8bMacN6cDKSYwjz2accXgFq5stQuwd0B0Z4BMVWuFsCF3Q
lcYXluJ5zVwW5MEOwg6jTGP+UnT8q9V9EWMfrnN369/T2rjOlRdvZypKPFhMDblfgPqk9jjhkUGG
sEp2S010Pcg3MJrGaS5dXMFxJTnaNldc9Bpj5GFz2JzK2skyhHsafRWlCli2lWuRAutgLUpNBpSj
eDdxwv1fmvyCziDdgd7Dk/irvNvDlTccXvgcquwnUNUnNsDw34gdw5jpP6Vj1afXXADjQLRbytPw
RyU0lrAQc+YqqNqIlYwFtXs/UVHI+AQroL2ilaBjWKWEral8RLkM9+foCXBS9KeLByrDe4Mojio8
cTiyM+JnzJzTxHgpz/59RXAMQyO++0gtG6aPaTs7lLAqStH7zdyyS2QMuO1N9IJUb0FZlLBZhv+U
OmoqTIsmM8JBPGLANOItx8WPKSVq4AfN6aDmM2RXWCuonyYoYMvkSF8yT3c3hV7NjAhWnz76dyC3
DyLQThdHx7JFyI8WtaLq1DvLInHTnrGtRgKPzTFrEJEMOisukkGjbUeokG1o871g/wqruijxU5l5
QP9ST0/IBgwcg/elW6XisKu1mb1fQGElgtoAi6fRL2ZgDfsvjJeyWMe101nU4hRkS4SrMuFfQ53z
glkRuxiTTqT7FAK5URjT4Nx6wOY6jTTxuEIbkYr8XtsO+MYVxsap2sn9qIcVEOCsw7O61r5FDmuX
LJKkS0lffFnr4obSCkZHvqEB1USbX4YdK9k+nfhzuWBe+VGNalgB0+sb/8UPsYp6kKS3aCCiTj/e
g/bjGsl+2nT4PjhOM5Jp34iKG9WuCSpWC+7TL4neaI/o80nsR3hCJxdTOUpben5x2stgIYxSuGRm
pOYAMAY0z1Bb91nQTBja7iGGeBDxxeZx5MjdzP1DZ4QnMwfGdQHWRsR9YOzWiJKNBznTapPOed3e
07QBQt4TpASvym+r2Tat4WQ/0I9SjvkLNlpwh9mWUrMAUa7uTWU2WRrMKsOEsFsVHTltFPFVeAh1
csac1fw5ajSXYZAbrJVpHtL6oeihdChgc4ETcBCNSq27ye37m4rESNtqO8FKyiO7b1f5Rd41BbYU
EHAtpGLXAsam+uDGOqFty4BkRzW337hdaTHu/4ULumPfDam551xjvyd6pgULKhh+WFOadK4EAaeT
DJA1jvhITQyuS+7SoGnCsfjJrZrXOYJvL3oqAGSBYsdrjHAhWcWASfF4s+kJVCnGPH4bSHAhGER1
EYMfBk/KQBaCleOmqD9r5SD4tUD/9aUlSOvbDwGugiFHUnI5NO7oZrP+PMwhs/tBFz1w3Bprij2f
mMxpsCLSffgNiz3H2NbZu7SigxDyUS7w/rSB0U17hjTgSmPv4AY9Ise1ckqTIW4+Xzu61z9jW4BA
C3W4E/YjVSiAAzfb1A50cuWhqF9hGMftmRXqRmaI0IYgLGX+8NasRiSh5fo8/Fh1Ar99Ye8VxAeT
UN5LK1mUBiue1uQCesbBrBhZV2WtEz9qwZkyVo+2RRgmrKejKW4EKYuQrvwk0ENsBE/ylpQxyAjj
bw2V93aSIdoZGjr4vOzA6DbLKBTYak8fRPJMKZOg7HpG3pwkTYh7VREBoTHFtBHSNR5S69SXoGEJ
BGkJ7Iim7HL0BQZkyKjHEIiCkmB82KOAP4Sas0wTRs1ISB3E36Yea+DVfygajpG7jeQ/YdwEi9zq
XJ4F4yWEYvhmgR6kvDqTM8kRMyzZvnLiqOCxgdvkgRMKQU+rFMhagfJdPMAvmJR10Rn3c+5JtWQY
DC4MEJQQ6ajFTu1WkcHZK8FnhmQPlPm9lpxNqgW63LiUigNbdoqRlwEujap1+5nyFp6c82L5S8/R
UdorGN2H3QjaL8TpGsxpM/cyZB+Dzbt0PHYTha2l66qh8m1h81jb99TW9qasNnk+ihUnL+iFQe3v
Y3qa4NYTqYuTHotRms0sZCy8TZKyl3nzg2y4VjrtwDldoB5EiHqRQYr95VsxiFxkisQRv4EjoJIK
EbN9Psh4aZ2xor/qp+SoblWleexXBUfaOwEm3gy3YxIJUPD2b19LeXdzK7wYU25szLEU11yOEJu6
/9io8udb9kSw19H9Z/PhjLPkRcRQ7EQ9x2aoSCFJDTuK/4VJ0FsGdOGFRM+WhqdJy3wNqh1rmJDu
aJy7top5gJCvMpLUOEgEu2rwaTdps32GKEvWSbHAtxKztV8zYNk7hwCtyBYaC9uJuKV63gGK6Ur5
h9vRoi3aN1ziVTAr0OWauzmg7x5lDpry+yB5Mp384zxVPLA6xGWZDvSwIdK34pngtb+9NNrfKrS4
OuXaJrMHPozheM0tUDAEwTlqFBzziwQDcOBbFguRVYkZil0yBnJuqayAa6gSnn37VDEaHByfgeKO
DqgbpOk4fbHmK1dKxFyK1lv5rBQNH38VeKtlPXesHDQ5N0NBAtxdTtRVEqiTJj46nuAH2cPJNgyK
1f8frdCHY5Q/MnBTxo0MXD/RvZgrt01rKg7VYLZ5oxQRKtkaKdQaPvUVaqLKJzdJCdmcYEqP8IFM
mT3i5WJOfOOSCo3k1pd/3VfXEJDHiuIWv90zCKkUelKugCfZAN5B0jjwZdX2wfjjWXc6wlZAqslY
5L9GwM1x89fnuaW2+MbVhlCBbhddF53LCt0WzoayC6P+yRm+jN4U2kuMJ6TVuT9HV52OUQitiO44
2FLeuyha7IklLfVgKIpGwJDOjJkETM/N9lFpi63UZ+CRvJGDWC6uZ0kSNVv8+Pq1V1BFM/REjt/z
IyQIlidwVoWgzpcXNO/igzDXyB92MlYkKrbWw0mIfkyuiCTFwUT+2Mg6iRxOV0/6UgaCxQ6f9HRq
FsdhSlREQGNwmF5qgpohpiRB6GvtNG30RiofsZ/gxJfuo5Ps0aGlCatuiB4IG6U53rYGmVYsOEq8
78UNQU0JuIAVbMWCU/wGjPJLLhmMamrEYjpQRhqR+gIgNgS3ITUMbFodFezBCGxklqH4OvtCBQxj
er1D3OKn6rDxYR3EH8QuDwHugZEEAOvQqhBW4srDwSHHqhPiN85oMmWTfeP3b6YbLUflJtDEiMib
2P75S9AI1xjgu13QHbqe1JxFOGRVB9U5RW2ipJmNju0NVUOAFLC+XS9WxZiZHwghsIlq5w+vsYPR
j9MAXdaOQ9COQQZtAWcWl32BogOTgp63zppuvK1cJavel4H3TzqLDWkDno9B0FldIl/5ao4g+T0F
uHGt3HqlIsowesRo6jR9DeFopmX9/JgUzrWWto7nkG2rNiOwlC1M6EgE4OvhGG1sPwLkH7DszI7Y
6kLiUYj6gbvBVwzl/4qyNOWm/5MQ72EGPF3zDFi10XfBAJ0MTsd+LeUFocz+7XOwKd7rPZ0N9cVW
NM7HzAC3sI0TgusvBQID6hW9oTCNeor9j5RX36ktd0nQkq4kbzYeCvnTbDLnS62eF9NH2C1+ZeID
6a8Kp7Vy5zeukrb8Es8ObiyGUVRe+CL4wvqq2lq5dH2ufDftyT+mQ/Joi6DwKH8ptCgd2vHSnHg5
MyakSBd4jOMus9ZBbzsk2lEoZ65NwP39GDnZtctqLLvzceHnUibR5lrK6OdntFOfTngicIf+tTGb
1j3qtcAId0pmloBTqbXpUnZR49ofdJmcuHEUx5kOkpItHqJU/MeEVFLU0ufEGIFBhHHhWl/NV07W
fqVZaSFHoc6Xce9wAh8YML/P19i4B8Rvyf8VfCYh3uqIrILx/a0w6PnfLjwqFuwZDZJyxHjMUrGi
cLN29v9u5JbgliTdblSp7rxyaS5IHhga+c3C8zz2idAkYb3Vz4t5hee/T8lRa12vuLLceK65UtCY
qmn/efES1MyM3HkWdxcxS8OHXhPzWseeCjtEXRfFtDXa8jIWJXnNOXBtid35RGjmYlZX/9CY6rZf
SNZbmrmp+sbnV3dVbKrssW/am5tleUhnWYQ15Y5o3z93QWLMJAUpsUkdNrfiS8zFH0xaXytY7UrG
v8RiIbHdDQuvGxTDT8+Aha5SaroFoPR4ahukqEk2keiFUcM6VAQ47w2taMKzXBNVY/LzvqwdNwnG
+BDD/hIhhNmGpvBUSycZZqQCwZGGEDFAlv84kTG6qJuTgoTwIuPfUNL6KBJ/3fbjEIjwDc1GT/Lf
Y8u4VBqdPnVIUjfR/56Pbc9ozv2qK69vNm6AtgHgaaZiJjBqgTQoJ6YUSqNeTVsr4u0eqbvO6Qnm
WcMMS9/wcXGTFDzhZViZLYmA+KF70PLLyYC8YNbOJBmgTmwvWmbzLlBmf5F3PJqphiNSUAEP/V5V
LLyju011EHcO+wKdWAYHFBW4YuO3m+Z6pNpFbJRaL79DeL2l7kf8SE5WX5MD1VuxYLMm1ZT/gYs2
DNdGYbrlH5ha3TCCJQ4nzruWO/2HdjY+b7tMouw2hxeXOYwp3/0GMtdA4JppRYdEtAs/a7+9rmmW
nbS522xYdriZ62CGJLSdAHV4XLNhZY3ndYIuxrc8SAyokbNP3Bj36301tT6vQ66RowiloNyrI+EN
zwIbh8+5mwiAcV3WG14vO05iGcx9a786JflnhhD5N8E36BCknZ6tH4hiZGIBfojIEPHuszhmJmkO
nncFF2zS22zs4/QtwzNbgTmAbm2SWnaIaB6TZ6Y4jSzNU7l/1CBxT7crs7gLejbyJs2j19lky4xF
YFOb+RGZfWY2kx7SdalGqCWQCy49S3ydIZuWHyskxk73Lim5aKdVAE7XzLJGfhJpmM34LETuFTtv
T8Iy69y96uqpGLto1Sdlxr5KeUhFRUOoIqIv2H/pusIfDTsWn6JCpGF5FHGrbfeu9nOeu1oym2NI
Chmh9hwJkpw1gLfRipBI63eZvzYugOiILjT5b5A2VxNwR/mCQGldiQDnrntuNyEtoLufvAGz4rWH
MXodcaKtkZoH7GqH4exELbl2yQTqfqJBvqdKhKqXxkpqBhL7SDXLloSlyak0Zv2QZgtpmR86a3I4
5OhH7ZZzUIy5+5zgOI1/93B5TSVINwRU7FW747HxnZlLePTrD0hnJNeHw+HrnOGJRff6Y15tZF5c
xuloZbGupZhBB9XRgYrVy5jKuLP3CIwNY3Zgo9VyCj6jAvlkU8lYRR9efmWhCYZEj2eUhNi8KNK4
oJ+UR9R7tT6xSh8mrXS+nAbS3nhxfNC8Wk0ZBjfRF1b4fcsRQ5IKa7yCbTRls6oJTgYec/+qaBYD
M4re3ngJ8eBnzJ5+k112S/HgX0EsPZ8KqnLWSmoVOWF+pnGolBK7Exzc9acF02NQ+wyNgc1K11Fg
taByFX/vyH8J9sObo+KsWnvCQPLltrF10AY5xan8fFzlQxUDGRhdemJt64Nbv5lC8zLItOmaHmp2
Fd8zrnUeqzkyDsZcVQh+7/67QtBbITSLl6B6hOtkMZiLs/zhKWXEfIBlIQl1sm668ITWU+H+KZtd
YUySuSslxUeDQwOigzulnihDkBkeUeBSTFsuMtB5xHWv+1eFbwTTqEWFmCNfYS4UJdPIPhsTuXJ5
miQckmMFhdGc1pm/P/RAzDyVG9rpxjo7oftZbq+pZDaMZ410XHWJ+rWlzvjjB2+1mUbqgYXm+JZw
Brq5I/qiDldTeVZhTAkrKTBul6Kq5LJhIzHrjUGRQ0rC0mJqk2KqAvoaprvLDf+O+lSdtWbyq4Sp
KviT72yAvw2UUUFWHv6+dG5cVFBgOXomRTqUtYq6MI4qNjq36Efsx5rFCuNxb6iqPa8FOpSto433
pMGuAhEzEqATgM5AbBDJZRk/puGUZU85PVbfVfF9VZH3Ph19wgvX2ksfMh8WL7Pzo9Pr/KUJJCPs
WjNZlWDQg/7/RddqBSpKmBbJCbD7HT4o7OJn1iJCSLLgx+vHO2pV9Zh6pzxMx8HIY0527ZuX15ul
GNAkUn2tCj6xz6LkofX5H0blfHntaNUaVxlFSR6dYkP/nxJnBayEm0sdXueXKONgdYv1WU+uNTuu
+U0kibhQVqG/PvxTXSeg9OHmEunkM/5JzENER9ZBBKIXjXyHiWOfa1g2UemeQDN8XTW7y0JqnfrC
VnfTEkEh9OxsBpa/BVdi5d2KGEzPnLkyr5TGZRjwdpQU0U8tCUAuKNWGc7DqOHiInhj/f2GzuvgL
/+PU6At8/UtPhqVyPRUQFYuFxFvhQ4+XLmfuTLQU6HMcEu9QPCG/EDAChurfGMHHBvE6Rf20ENR6
PlgqDCALJnl2UqD2RGKoGLjV9pkFtkjWS0sDj+j77lbMSLJBj9UUckqE0zWkyYpBVUk4B6ikbCO7
gY27EolA6rllEk5gLdh0NtFcfgV2rbDLZ1yXNZsUUrVgaIQCwplAKCTkePkuiTmMrsJhVP8sWKDD
ipw7yZcgzrTndLEHG+94rLeFWJymt0dGw+CMOuUC9NdFqo5ZPkSFs4lHyNfue+MwnPV57AKmqdPA
UAclIIZ1OIrUSpRsy9ai2gKu9PDCCajfe/rIixInwGNS/i27YvRE1RYVp8FMbLmjWOrIixheYJFw
Z3JFd8/STHhB/P5Ij1e2g58nglNmzkgAJ1ZgR9OEJ6FKoE5uCTgKZqhO33zlgtqLE9rznQOoBTLv
gjryML452uh3McTWVebNoSvwrCBibJy4NmpAG7LlRU8AcyvwZeguf8258CIECheYGJpcKoNseSnx
h95uHsIFY+IF221Xs/+iiDJbBJdBLqhnnLJUC80uaHIA/zpbVQBAQGjHV0oOwpOWUp05l8LguLwO
fu3UfKoznsXDDcPOGgvTQYJd/2SNNHT4Od69KmbBOdaKJyTaUwxpJdxGjkI7KDGdgRndJ13qUbL4
AvH21exdXqveJED8zWM0IJz5LUlQ22ReySnKwBdSJDbYxgAndjZOUWFxmnPviEDBSlcJwqFC0gvE
jNSkdQQ04idiNveRJrWIzQnSx+Felt9fpjG0CtzFmOx6/SqVQNtqWQhepklgfGY19niaf300QxmO
PPijm3aDf5EQiiYloDunCgO2kHWZpbXdTeEl3G+XzRDHyNK4Am0Ky4LVotnbqg+3uPJ5gpv1WhFv
opdIxABwjk521qEKiXi7msm7ev6Kq745kcpY7EexxUNAlmGnNgF8bnLRBhI2lMxziXjqcnw6PXhk
l2E9TWzLYBqaFz+wu15FjEG3a8D4I+cLrqZtW4o62nGkr9ar5S1ihjYEd7DO3mrdhZ/w2TVvRH69
CoHm761iviAx5MoysCBj+vgU5+Wz7gyhQHB7xBMJKZwQVRkZ717/CszVqS/NBbHuc0haj/u/XjeR
Sx347EosXTznFLQaeywKYWsWd98CqHvQqGuOkL1AgHylK/0CIkFpzwM6LG6lgc5U8y54VwGXN7WK
BGPxoe6uKn9Yfzo0nngi8a+ZnjJXTCtio1CVcIjFL6BiqwV+5uQ/RzVRJODxe7oH+tVIZAswqSdd
VxLAhbb25+pORqEpTLAONAib+q1LGKYL5EVWuSh2i7DiZaYk8vgCbc7e8ZcLMPPdaVaxnIQ5pnjm
0cq1zJVAua2XWdrTxQJjUtyCL8klNsJAzdbmEsKuvExz8qYRsAfHk17sbaYJfuJil19Z/Iaa26oW
b9+zXYvElZqint2wdBxtTMWT1FPn9kPnzMhj7FeFlxRUpC2hxqYfka07Y2pYuCu+wy6E42p1PiYA
LFMMjx24+HC3yl9TsKAsytgT6p9wcLpwR3h7GM830VIItoBmjXB/pZRzbUJbXvZtxIK5DgevJPTK
U5GpWkF+bzFiGdPNDW39MfQJaGZrSm83fxW/IyocddrCdqs3m2qNbGVRfrOzXWXi7tf/xmXyH3kF
XjfNjl2NbwATz+ufrS6+B9MhNRMQ3t2DxcNzKv5onqeX+PKIt7dv4HWUMNKIN0OcFyR43K+kPV7z
Fi122a36ZrTpxMhIKrngnJkjdYuqn7KSmtGFLwTTV4c0neriwQN19Vo8q+02tbZhl6z6CnGf/oFE
Wi4SjytBvn1keWBDFd1X0O6D5dKxRvo4mIF8PMn+2sGRsw159uAyVEn4nEou43j/HXRHZUa0wSb/
y8Mz9orpiKekU+fikof9VugXBaJagkVBff0ef9COE+e7OIua2Cm4YCRxwMe8KJsLf0Z8Y0zVpTCb
SjOSd/UYYZsL/CAxSVBace5A9C0hN5BfTQZIkT3ndc43C9X04eUkckK+UFRJO/vb3bYTK7myxLJJ
0AW6GJthmVv2MY4jWT1RAKWB3MqYIUVbpvq67NVHKCHIs2UryP9aMu2RGCjOgzgGKH3DOw8D6PF6
HgjMzKQ9eKNSMDji8IhjsO9c4VCOG8Wml1hytoxGrVDbpSas+skdC7/+SQbYmxs/A2G8mGxcgznk
Jzp1ISR5LCbfR5WhaOIwbff07Qx9jFOoEK+SS/+umChPB21c4iuaDhLfXGBTOkR0AZ8qHUWjA4yS
D+ZpHrQZdo7P4KHUJG0oZV9PkJzwvO/hlNZC0n14BQV7+KA5wgd2grlxPEdQ7CxpWoJkIU5vEv6V
Xcjt9cP+2bpPa4p7ghgDZJdxUjUqwilh7d7zDyv/M4o+O4vO0VHq6bdXuoPIsUtoK1uRnlWJwLdK
8uyBYscL3/tWLyCwRSLcXGomNbSqfeURlf+JCRIGJImX86/Uwz0AUSe01W2ksPl51SgiHmiOLuQF
SiuXtSGMPKELtXZzy3LDzpiQbN1oWYJ5x3/gTl3XpGC8ooOnnyQi0xu51Ws2Kw0ggfma9/QS5hmb
2uy77Xcy+b4l0hCzF120JsoOKeGxhHCvoOPA0jfaCSndNnnBXBdWTIWQmGG78ncZv0M04BYl/Z8D
3WpSNQ+yd5RseOO4myZ+m6MDpDRq4OOpLZXdw4nMA9DF19meWX6rHb7yoJuxC/8/fCE+x5tLBoFi
npjuSVQQ/KwjuRxV0yfnJZBh/P6U+xNkvHvF3ax75wcLfU8AEh4Hhcfog369MJ7ViXuC5geBb6hc
Jw9bFi/sgUuTZqQJyeVxdw0wYT/rNWqyYhyKRrhuPnzVBUPsucqL+/9znq53TFkBRYrMQEli61RE
azC/42o1Yo7NvmbXldlxWxNpPffX6lc5c4R2IrWQXOo9DBF+Ui+m6EidN1Y29VNKebkfSHRWlMW2
3zeU6vI0x9l44UCda+x6o2J96HdhcuD2Co5G04T87rVK7luzcyTCsjpvQD8syOCBjYAYYZ+wdi2G
WSw9Drr4pMQE2ytPafw6FyMXQfua2A+iXR3tNcpTEpBUpewImbc7SD62pJvfy87WSrFtxxqTZUup
scy4EZU4PSpedETwIVfo7tbQItx/v5erSYRkiCxyDtsr64bflKQ5Qx556OSTiT/fFs7isSfDqmq+
VxY+orbsPFP+BMzkQ7cBDdOLjpjNM5w3+QClm+F3D+3q4zqRKUfIDC0ueTEIehSsDySV/laKx5Hn
6wWjb5l+ft82eSCcOQZ7LE74xVOdVryu8sOIsaYe7XyNJxZKkVnTsGuUM1VhaeQjLXOotF9hROZ2
Nwvo2ZhVzhhJAYcI2lg43bIVKfZIuKSRD8aH5oKCI3yK2t9LXg+WAd263E+GJe8pMtsqVOpKoiuM
PCd2DwIoqA9lK5B7dVw/GOfxGWDDK41my9Xh3VqyKOBERe/k83BoMxBFMUJlrYWvxEa1uHGNftir
XQ68UpvKylhuJ2ZVdXCiFPKWc8i/cCoaJP0PSYsDg2gSbVhsH3WhhlIvEArZaXWy9hr44Kv8MXUf
jXQ9B+NvypDWY11HZhfN2s+QLInyCDqflwgyB4zn9mBHtldXAf8EHyj5rNUZILKWglnvD3rpWyM7
i46qVpzi55WtMrprr5EZg+HlSw3ZkAdiJWwiZzs4luUhGIMqrHNetC2mizNY5AbLjYaIUJ53LRQ3
RqSQk8LQI3BauEMwbqJnpQ0btNPhYOgAvdcEmRfbXdRCMciUC+kxZegljHtoRkJUD8pLfo+sHL8Z
yUaJEZcpp0tjtGjyqTzAQK3is3hklFGzNN0A4CycbYdW9NUfHr6B2+J+hoSqZv6nGPCLc40MXTIp
TZSYJKnErYnAOJT+C928hR1u4+IsdNf1y5HGHr7NlHJMu98IZyQNvEOTo19scFo94UqJWDPP8H5T
WuI260QYqQUY19PZy85bD7HQtKOMFlTcvCwx2MTDdiCpjG0wWWCt8jlUJhLQKx2fnZ0nFTZ49bu6
skkxpBg0HN6Gb8DzwTM4OhFlmhmSf5jatl05K73DNUMZeErEaMoPKRCfGx7r68XQxrJeTe8jnhCc
LfBwIrS95cskRP6PFGS+pIoHBZaz43yYTAUFL68jnfrUPL3dCEpCa706RrFtSCsEYOLDaBj+tLM2
gf8ODMJyTsQb4adqXfFgzcnbxQWgr/bggoFtA0nTTQdXLbyM5caGMKR/MOtDNuIPoMXK2Ru9o2ZK
Z1afBNLldwthjJqu1w1cqLyPLkkQPGAbgLUNhzdrfp+CKdtPIlGBksAQ1rz2y61Ts2ChZeMKTnDF
hPZsjrnYLKVdpiCujUq4lESzgF9mI0dd8Cb7vYw9CyhrZDUOMHxM1Xs9ur9+15ZdMZ4V7AhtVM3h
SkXg1hW8BZShO5rVxI6qwWkEt+Io0Ika8JjXg5RnvqgRwgSzQdIoHmYt/SSjIVx6aSACqlLcgbgA
iO6qr9dAdiL9dMGe7t5vcMpDX9tFuIkJXLjmg6hrDqMTPNSs4xMs8VXOQm/0jtQDgQQOxEa6Vcpf
87wTr17gJMTnxRa5f2JrtFhrWdbPi5funL1wjeOzrd1/elMWUMVK6FzzoKdjC3RKMgXCrigBto9e
4+Vb3bHGNzF+jkkGIULjlMAdTn+Zq0unSq5Gv2Mr5Dt3v2uxK7x3YOgUW+XqxnxW0iRi8sRq+Hpd
UiE5FcP9Xv7PeWX5GWXWUhcVONhD1jPVbLKXUu9zbynUkqlruTicMngBdcB4KZfmiu17u0xtgccK
2AXlvW8IvZsBFxSG7L+kMUe7zJtNe7qUmDY/iLablxZTQzvVLYoBc1lhjMccmDS1uWDT8hZVF105
3nPf1FxoW9NW0Hg4e4h9g8c0Ypl1aQf4A6nPyC/HqDqd9xuxuLhLcqKrD2JhZAm4Oh/spjPWeHGu
2P0xHRB6A4K08eipnCE4AtSYytY1P6tNA2RRAq4oQl3AqDhjONuuSrpKu83m9aIv8NMS6Q9y5O+N
M5m7r/oE2kD3MOj4gJvGHhBzQUqQ7CP9q5nq4NhCUVbdXZU/7xpMqk+EGzg6nADyqaCz38aq5Zar
8LfT5ZK2y33/cfZIJr+Vudt0Ft3IerhHYhYHggmPZwVyoltC3Rs9ni+ijtMR7mr5wdV09qt+IwzE
SAMbU5psW9g0hF3rMJ2DmBVlm2YQSiqrg3vccpvwR0mnXVkjHVlwRJjoFEe82vpBAGFTKflkZDX0
4j7udFV5YqVi1ib209ezmUgPQF6kwFxdG422J1uj6f1vncuczMi9T3EBx7XbBs6pAd77NL4iYvYb
yDG6okb09BLfHrdfJIyXm7H3TkSjomVnY3tot98hwBi2sfHDzb3Ub5Qm8duEIiBUNK67v/7ELdpu
F231EhkAzWXnRGjzOsrNhTV94/V9vVCGROEFAyyu6Yanq9EM/7Kdoc+EwEoSZAngSX/0eiHjHNjS
mjFchoLkfpKRk9TIMX2pLmvAyi2mfp99Kbpdu7v8hPM+uAE3JoB/6wKsk8bMnWAhMrAgpayXyQYU
KIb8SKhxM2TtnEyUELHINAnjdOrWH7PnkiIWhHNNMFqRvsjrAH4yb6mSjgULgo8RQmX6exb9YvjF
bS1azgljD2e2OEhKho7htV9PR5QScGCRymuvRg9IANCOMWQepMPDn+7x0TV57G09rB6fRSm8RQ+s
s8nLTowJEKEjXuCL4fcODK4wIcUmAaQUVdbGB71keRRDUMx/BUoWtfFJNg7vpxoV2nr6sUr7/hi1
k44JC4SPIz7/MaxDOfXd0SohiNm7N5Oxl8Nkn6z+tZOfl2xqSivRDXNyc45yAp5X33h7I057f21y
T52naM7TprGQUStD7ony6ivx80G+MtaQenykIymji940yzqPhqPcybr/lMqLYCu51bT+snPC8i/T
nr7ZPP9hpfR7L3wd4PWIY1aZC89QChWFKcSf0jUvm83pQBCzPTEGoZsGyfgIjxLDJ/ua2Wj6e2wU
/QCrIN2qma0PDBVMAHs7Ust5eMTO2C+PEK7DdM6zmE00DC7yYzegRGRC+mh8KAa3Z3zPmXl/T4VX
yb6eE3+BJyv4GPV0a0uWBSvFPLP+wxrV3IgSzI8maF/c/Otq2DYQbkjowQ5DOZ2lCkhE31hBLsWj
NwzJqsrK0tBPbH5uzPgByzPgXk2FtwR5hGDLr2PyJmA2Xyn+W+XPNTOAWU7NTzelyAyuQ1Dz6P9f
aPPjhWVtIIV19fBBGqjSErF7WxDOVFP2sjNFgKGyCiPwXyp1YruYqVVoLoG+aXXEbz2trrfPGuhV
LcqizC5hHtiijWL3izmShWjOAvCjBWyvULkbwvP1Jjow36JCSesdWNXEM3UlETOov4haGCfXPaY4
xBHMA0CQUvZT0lTMhtn0nDEsQUdAPZvoyELThQpUcSQvvG26LgKikmrOTlgAcL3AiVRp3C4UC4Xo
DKbuMvl788skogHjx9NY6FV2jemoVQcBvSGVmZIm9yqxy3geS+P/MAFTiw2hCC/NGrKaxEjmN+Jr
ZQt8oEtO57WOzIr/DoTV5Cwp2VbpH1G1ZEZjuwAuZClyOjcnYatOveHajWFGD2izIty9oBaVtUex
hcDXoBD+VWyvefa6tmeRHgNjzcXG5GOBn7encNlgKZopOWViu2URFzILGjgbWcL0Q5yD/bcUjjSF
TC8nK1H9NxBabrm5DuhAOTsPKvQSf7/RlBiELH6fbmkTxA3BWoMjtHYloEo60q1W2o+38xPdy+6z
PpLrKAJpG9PT4oeeEDEVpNB6OXdF8Kp8OES7zOpnpzcAQqFZ6I4yosurdlIFxOGOsdXc/SkOrIV9
KI49i/X0z2V0jbiH8gzyHJ1bHOUm8akzwfqdmSAO70UtnWqpqxMiXXJTdZrIjnibmCeB55biIxRX
ptBqiy/5Mu/F3TuQBgN3aymJNUxhdl/sQUBscL8atpuhe1ufWf1ucQ7ZGWJr94gmzFQe6+OPWSFg
QZMK43NgIF17SQCyKOiFgsFR/G+t138QopB4qSqFFKF1kgJrg37OwiPFvJi9z7degQ3Go6KdkvCn
XyTkHw4ofsiVTxntkN0yQT9FTfRpizxzvZOsaqIst7cljujWBZanP4646kv04kZ/FqGUHb1Lc88U
PVkenJaaQUbqyi4duGj83vxoLBelSr0ZJkaTiFcnZKBp63VGLcUtMSAYZIZgHDSH1baQpCwXV6e6
Msy34hmer4kgEHITM6hKmhBHo3E7aC/iGnR5SokUFUnoZpBzqzxVgy93h5LbB8zlbm9e0D7ETk7+
YFy6Befxqh54R4RrGRNpIYwcywOPZvPyHQkrGn6c58S7pmtMk/Jw6xN/IrCjwYkO6ypgZ/5ArXI6
shyL2bnDC4ernZGkpyqT8vENPO3DWjPxbCBLeYZbBiBKz/v+/9e+mzcV+lPD0S+RUmA3IKjwuUeS
9RlEguoJwF7xWFayVEnbQ7L1Se7MKcFTR43Dmt+8Jmw4bxhg3DkYv7oCZ0Xmu6K9E+gcKDP6cZ5v
oM+/d85X0Bf6SjhAlXf0QLLon3POjcTm0BjO6GIwHtT8pPc4YAlvG44mpHyLzIw9DCnBYxP2SMfH
YtEK3ZDmqo5/nUntpn1BZ9csCJHdSeN3XlBCUk0ROybH2V4vnWKL/41q/Bxl4vqBnCdMTpUIDARd
D6KtH4mIUMagyCZz7ltvJwMGiHBb/BVx2rkPXnyJrenjp3jjUvIE319DIxhhUMbvgJyc83pVxAxA
u0AOL8DUk5G6mdJHrxx5VVv7qMAm7dmuHNvBQtdzIvbmf11WLMhRgnkR0bBrrKf3RLgSKQnqd09f
SDoMfPQbbMJ7R9qF4S3nz912RWSfafJmDmAR+l3qCQ6MFXKCD7RwdM1ykucOb3NhckBH1Cu+hZ0z
32G124jnbXxxfyRqYwNwjU2TqZSdFkT+IaZ1vluH27hBmsBE7WcLJBmJQm4wpO4F+ym/f3LOAUqs
bTTciL2nUsc7uakbthhCljzptVhVWbGp945kpLSeknWYt/aObeD3RXkoEJpxERQZ13NHttRAEMKR
6JPbDcdvsyCe1CQtp4PAf84OHXfTLLiQ1kwmlNB5BlpOXFA5FcKe3nqTwdhWguBxRMox47qF76M7
RdEZ62kBbty8fER0Ukui3cXgXeeYpNVx2p4GFSyRtaHP3YPwdQc6BbX2AHdcE4qQURe5t9IXARmx
3Z1fJEd4EZdwTZj0A5W92p7jiehUuok1B/dSNCZRNgqKCIjRvDARjQAhWlwuYYt+SFNOn3eg5u/k
aXUbst/x54evlvnkpPlaX49LdZjpAYGf9HzUqhqOddAI6UlHSCHNDZMbHzNlhYbra59f0LVldLpq
Qq7AE6Bvn1lglHcXlGIE/w/gXHZ5ue78D+mZtlBrKkDAwS4lDvRpyhUtGsHNhril1xcURH8cqc4O
BUyim263Seg/XpnaAKz/rD+67Rx0oGwyx7ESkaf5/7zLaJNGFCUHrpGYla+tjdLOI9ONUtIf5/LV
+MpExBNCoVbVLztieNLDB7nCni6we9hss5rNafHBFFO7AllQolhhRLV/ELiKVrv3Dfemx6h2QP17
eDLnljU8ib9lE8fgJxgt/0il//S0I3Tp31cIKN6GUu2hTxe0DzVIc6BnogVWMKHdGJG881a51yW2
ekWu+S3SJeW76PV1Fomk1V1HQ+8zvc47L32jLqa5MRZbBr326AvQf4td2Hf1z3NnbzkC1/AVuhi9
CNEw6SG5irgYdCABl2qamhjAAd+GNFsz3ZG7eiGZFLot1bBuRU1LYpdWaGyCGmt9ePXzcJCNOL2L
CnObFh13Jo8OKGt18P2mbYYoAnbtgjrgVbUZfMJQay49wu2qzGyObx20scvpA+xTR/HoDt68Y3re
luUH+kyZwmjzyBMHk9b+W2zteemorFjp8XKZVpERaERK2lLKtn+AyoK84B+465EBstzJwlPP3yo1
Go9nJ0As444J3Yc4/LRLQUBGRev7dl5o6/u/NDPRuF2kFCVGMlkHxgYKp8MA8fNxCUfMgYWZWgg4
bSeOyCtHMdDOcKRIbdfpSORlKvFbqW7sr5kvwCoC3aotd/WvQ5lz3fb9nzuyMhT8QGP1pSaMGZtC
4nShxvSMIszCYgRgkD7F7HQUCzIs6gt4GKisSFOfVdFLmbEoRr6fyTgUvIYQdUK5pvku6tqt/Tt0
5cySzcvrhs+2WCJr3nRcbCz3Y6vjwyqr15YWvdvqI0JddlqRiu9+JGklab0Hpd3IV+vSGdZV6PRK
jo2Xy7h+rkUrwwO4EL2cTzzO54VHjjUxqKWMY1Mm8EEO41WeyT/nN+phM3IKk5/cQXoeCGinLyrA
bOXW3xqZjjGim15EWsFsIRRQJcQV4JewJ3zR/urAkRV6olZOg4bDZV1yrI98CsLBWW5FCS1aErmw
exmJbnt2uB92S4+9MReJroca/uTXDQAzZtskCIw/hSPIrIHPXWGZw2n+R3krdT2YpTbWGq6fH7cJ
UpYeB0aMIf1Fqi6sW1w+rsQTESH7WLfqFoGMMH9t/rsHMlSQb+yiIfSPVjKV/XooO8cPamJOFgkl
lKkZjAz39Jz2o3EUCZ1FkTqJuTJVcU4/U1wybYeiOaXy2552TDfT6lmWKChPnqLeC9YP8Nf7n+fP
C+n/rLPCcTUahbxyoyas2l45TWh3lA2Y2Qtlr2gEypQNlXwyOpYkcibz8UKUNqSxIDELPofMjULN
RPy9YhllkHCbPQqP+Oo6qKPHeAXkSfVk4UBLITPDOoZnyJPpPDFPKfK9jupkGzhL9DOCbsm3pyHH
aSxgXrJyeukrKrYTXNeb/SJ1heKfIErwYAn5Jm02klCeqAZEOtWgqFaIYUQCTRo9Aplwa5iYmpEG
eIw3j5tkUoD9AE+Pxeqqaln8RLAStAddZmfJO5vrzGEdnrjL7+SKtzhj2fY425bY1KrjcY9QotbD
lJEFIYYRngSdXlGXAVNMpKCaHp6H53Z3UqnaG3mmbcnijGntVykBMjjZr/osG5CvzdjTzi2jhWFn
oAd1lwhR7n2hUiZJuql46vZdF7NTxFAYv10IWgxxb1ee2yF71a/zFEO8H86DoNE9oeGDX/xBtYOO
Z60KGKg5/p7XOpwFcs811bomzTDmrNlNnr4TGAyOJ5PZv9uSFdYUSiulGOeX45dvEB2SxHaFGyTt
BpryNd8/w6m1bYH8N91ctKRx8MTOH3K+C+q+N1LIJKwnvJTHCKRCcoWV4YjTztw6PEx5Aj+gofax
7TFTQZGot09xwZskMDmIyJx4weL4Smz6+RiXj8GryNaTA6RCxilQhwi45jzI/O5iyRml5/QvS8wi
brBzprxRx0nLMh6U4nAHsQfB1ER/LoTLVAWovSqv7/ZtMg49anIR0yR1eqLaz6OZQTcGqq8wXhlY
uUiSrIn9sByJ+tOxdTCczGE57fXLiwI4YgH7swhcUmWc/doXCZzuJVeq/OwvJRykaRkJ5YDNjesU
ClJM4qw3gY9Uca7Pl8q+fq5V7WjIC+mkfskfh4mwmH+47yDo/d9EnBXUXkSFi+cg8FJcUFDRGgte
vizNIi3U3n/YIQeBRFMm7yUFVp7Xv9Y39PjLuUgmRFDFJr0xRObnoXYuRsx6MgIszMmPwxrml9nO
dxIV6GzGz5ogl8gBnXrTXhVGadSyr3DFKGX24kvSJrQMeThmox62XAI1wdsz6bIulsRYMUJGqygQ
10Y7bWELe+jDv3kOgXJ0TiqJ8W9lBdGXkbqnvdoBiINzNrVX9ay73BvYyWPJZIeCXz6IgKJsYEqR
7j+n1Rp6+aIl378TKFH1PLNfCnElCrVrIy5ibsaqhqB8TG8ZjcHxckWDPvGSPjHkfo/8mShrHUq/
tOQ5+1XeAD95Lpndzf1caOmh1+FwksdAVVEvKBn2HiSEdS1IKZ/LJbt0YAbBiiPbIEcVsOLt0PIf
iAYc9uu9UrVrvLhFPsNZwxSa3IwW+gmSEiAx6aeSVJqGzUJNiu4NsbfbO3MY4UsJwCNLYqnDoYnF
2wAylsTg/DdpXJf3mSs9qW5e1000Pr/Y38xthD8jsbow408svL/enFQSHtLD0O2dP/FoaEDyEQwW
VhI+7OaFN2RYs6j1IC3Nx62eZPIXcjLxM/FFU3LI7NVfXnpw8S3LVzG8cOTQMObpssTajRXzVXad
IXDsDFdaDKOOeBX6xZFvwLZj/5bWMOsMA7n9cu/Ksj3UqLj/TnXkSL2OCi8a5bpfaZ5wzzxqvCi0
cpRTt+CrNqeAHLP1L3+qOIbbEgkIAUERooU9KUjzRI05dN1l9BzvUeRg7AbDOuZzk699jeP4zGdn
DCZBwXZMd+Oq4MsADz6R0jGLo/WCOPAIjmzILNKsUNWBKamBpXHIQYa6eXP0PonJbzFibg7vGgoV
IM8Npg8Kkhkn4l9rdn0T1B+vNF4awbWPeI+kz3J1ppHrHYwurt2/m7AwqNc6W5vD2MJ8Yr+HFvas
TvvOTbU5HvI5NOtjGGwqMrI7RA0PC/euvo6KXhHVmufo8tZUau+gDTSUnipEGUAhOLa+5fDUfaYV
VQH2K6/l38KYgXSWDJ7xt86ZJQHVeq3X53bup/xOroQRaUQPQBeH0jDGiKS7L0bDkBbfUwHznzkQ
jn4ptfeR9kgB+EwODlCQoXlgMOuoCGiILWBiPmMZ5f3z05iSaLn9+iZMwYkfNcLbJKAFVgBCFvYH
tFUl5mEpBu8FVx5QOe9lUxW25D/pjjXdtRo2fltccSzt0TxksP/fv36mRplyyMTm4EC0y+0mBypN
UMFn6FD2SR5NrtK8/RRowO2XGuLpLFu6G90hqNHY4hOKmSNWwDyIBsXLAdQeps/dr741xmBVUanZ
OdrwdYJYPcFVWul06/kGBeFbi/Ba5g+foqw5oXwfKcb1MO+Lh/OtAtWffHk9HhW9vcg3o6AQBxT7
Tp58l5LjNSSLCoPjR7PGlssjC2h7LU5rr99zzFcLEjcEWpZ3FnSSGRuQfQCnVlBlG301lE9nHRx1
M/A5pTuyDsl6MG3IIMIBgs6b6A5WWPiijwxRF8rcMsUxuiKGYRhePruYW/93mpE8v1i+tvee1sz+
I6l9rg40InkafM5S3SeA0U08/uPfRt5K/JekJ+WBJYojZFK3agHV0b/b4WwSIlKLRsVUxfnJrp45
nY68han5BPFDO9bR2PMekCjFi3b26zH6sVpkps3QylRZyatDBNLVhgT9J5IYAZmWbv0aADpdDf6O
7gEGGz9ONEW4F0qyeVup/YROVLpqRoNwdSJReAZBDMYSRoOYO6iqyKQhm6FixJI2I8W1nmWw10pC
bU9SrRZlKZ7+BfzdAwK5kTWTGIQj+X3n7Qudv9Hjv84PPh0mX1BlnhTgEP13Ve8wumIN0oBKkgXL
NxNOCGH3Fa1zMJzAX3Qy51K27xkugtwbUbvctmpNLpxXpGEynT/cqcicoR+q2lvjANMTqnAAvMB3
cu1pIeYUn1bGBuviLTaQwKG3ivcAM4sUymB9JLzWHFz0p+YQp9H5U8D8H32FnZPW5Rw7DaRGk5PR
yV3u+7Q2H3I/LYtDpPuNXZg4KEstShXAF/cMZSfsSBLG1S0DepEHbOGF2YixtofVipjvt+8ZyT2T
t37Hh0gSmLNRLfV2pXClU1zuXpJMulZkATq6kJ2D+G4yEfC1Zqw3pO+SJS7zm7kOy5+xe3vBk5E/
vNHMAnH0t1yR2/eoLiDVLG8iMIVg4UHr4ONbQykCvgf8rbNHVW8S+ECrSwjgM7aqXBOqvUgcDxRJ
asj13AYLpdmWeVmkvEw+zT97s4nf5oVbU8TDlQjND+A2/sjE+hra//vWTufb9vAG8oyKayYh5BUn
aidrZLunLAPaLrnhIYlABcDEQQeRwQyGBqP7T26h1NxfpOLv6rlr76crMO7AgjWVL4ORzln8/CWh
GeXn4M4e9n8ax5ZcI18qJ0IOT6s0n8DWerYRlpbjs3kgijBrFCNIVhCwW6Yv8Sz/2XIMR6TBtxGd
8ht4L4Hlb+0BuWT42sYcFRDgRsIQcmYQerkreqDnwXoseX7LQyzWZiprLlS3JMQdlORegIJfXAQC
Ujc5tLOsNXQYSWituNhmHEqEQzlxYE71+PI6IqxahF9xBq6u7jAFyGjoaOqPV64FJ7f9fKde26uq
7vjecH2fW8sEridTxsuhORFjq858oQ3z1hHs7MbhveInaaNWTtpBNhX4KtKJOLmwblySwT/Q+Y1N
wVOWpLnxshAWj+iCdPTkM4U510Xyk5V5Ddh7d3bH8UUIasqJDwzYN/wmDfPvcvQyiHwP7ltms0xf
NnkYVyJFyJuvpd7YghOlMS47eRHntTSUTwEzutSinuFy3c6zIIGPcWQVH4V7gik9yyMyTNTIV+mx
Pp1784JbBpPvm0ZzVisqd5NqinyagG6mgJ+Ajwy2QGKrKe9mb+1cTQ+IS5Mm6G98mBAgA99Klza+
jzz3qc2hk0OeVrzTYXumgZVgUp/dINEN/eKw+Mlx3DLb7put0xqzDhCSiWwaVVoDsxrkhvpCrBej
OHOCRJd7+USSrZ4WF3QyZvwBeDpFyC1L6qkWm1DoUmvS5OKpcqbCC7zOCI2x9nrG2gn8tFm4e++L
VZcGAEyPylZuw//fACskTGOdW0KosmlVXKJOz6sNQa9bocDlYJ8HnKy9iz6pY+U1TRlAUQE51g9c
1h/gpNemntMniwA+Iv6j469U/OEiig4lH9gBleyD1xZIN5CPQ4Ee8kS/6lb5LmYVtVRGcup/8UEo
eXpLiLRJDCxuaczlyjxQe0E+GpIvWw4TQ0eAe/B7JQT72YR+RZ+DMktagT0yOIxxEKqVVynylwdL
k88NxXJFLwGAxGTrLG/5m4Z5W96aB0nUXN5+6GXyAEctsFl1boKs/Vj3RAM37BjaTkGg3o46+xZl
en2AY0sRAV/cxgOp/JSmq08KHZ5AUV2MEyKpKb6+Tb+YUnoFhF8HymBQTUlKuFw6iVNRCdA7xq3N
sOCic1HsX9k+AITqdJwuSSZ4jsGheq5gMaT52qq7IZ+us9mcZRbey8VgOEPmMPlYZJ74j+eKCGrU
yBmf3rILYAFavW/v13mODyqgxwlZF2n+QBgXGaqk3+PaqtXrsEdd3WAKuP4YStrXgrkd/FwgTqv8
g55bnD7BQAxHIVvAojLwe9Jz+NI6R9P77t/n5JdYCUznUSaxYM4q/L+ovF64rjdmGMwbqdOIz/ci
nUaklgF1NOO7XLEikNR2xcoT+Hdhl9UHkfvGg6lvTbdt2GXxqF8YCoQORsGvfbK4U/6lo2YnIsuO
jWeZRg8OLxuQxSEbKiJN2BcKZU0IJ/A7PAsgeM662EnOUz4w2M4tYyOVcdjMshE/MLQr19x26evQ
7rajIgwAyxDzROki+eBzlJQQnMifl2wCRW6xnsaFori3vwdWzOws+ETjn3vNLmOSDtVNsPNLEVBu
T+Ub9RfvX63x+WTjEgVWsIUVpL9LGUtEjaJTXFS1AMcorQv2EEQQYG5cN2020ovbKwO8Oke3Nzrb
HuQkDVhfuZNkkIW8Gul1Ky51q+dJV3TXKY5eseMc4UtXBmnyeCv8L1v3hEVXbhvSheBYPNNAtyuU
naoxAQRDfcVFK7zNnbCjRams11dWxggoXjAH14AAkrKgqjo9ONzos/Tv03NU8HIz+WKd1GsZL1L4
Tvd/hPNAy7aUBAzapaw7arWkgh4Pqh9BjeS2ZYKhVknu5RDa/s5KfW2KdN4whJhZO0EuBPR7qr+b
5CNMOP3X34IXLYoaX55rDaYp6NQknlX6aFWLxf4na83NOjzU7q02CwxqFnsDFVtwkkYt4Nch0jsI
w+N+wJubUgLii5i9Auwz35YSafnpS2gsS6Qiz0D7VkSk/8lUYgTseRMVx3XXlyOQ1bs7jo/IxYYP
OM38mgBdVt9FXd8Lay84hbPn5Fj8iIXnNYH4e9xhxiPcSFI+gZi7dhpH8oPF/NnhnV+uTcMzYNAw
OV1HXcDPZxL1C7pPtq5LTzJ6WgZA55LMLJny9PsdCEOKYND04mjQ60Gi7U6DGZPCUCaMCbxmSSE/
Ybl/cCjiiWZN/D/cllOp5pnc0fidaN16UtGjaswdtUk6KLLTxinwqhTPy+INPdYZsJzXcCM5ZIBB
NNQ9tB3PSmn/hE8zCoe/tpumNnF4JsLJf870OuLMN0VY3alKD683nRJJfpwMVXvCvP+c6e8+QY5s
AnoJzJAf3C4Q6Cdv/m5FhDrWx0017R4REX2vytGFhvMWoeJB+NmiasFU3fcwkDQ0sEdRSPBf9kL7
r++tHmqWZ5TFXTRDQjST0amyKWTkafE6FOnS1DliCovEJxX03WLZPe4KJk1V/dKSIIUMnlV+pwq8
OY5GCRKl3J7/YaB7lNJWfyc+WIVIlAqhF/bGUzsFonaeNNc2JUR2+TObFgHZ2AAXo723Hxu9PmlQ
AVExiiMGyzSzSnDqqiWg+7HpzC0mkny4Lc/ANru1BBbTzCsDhK2aNsA3BgN1i54DV0d7sRVEVVZj
gRYh27vu/deGkjGzXMk7K/rJv98OafJhhlyvegXYGN/wpUMU7VuoD4vboktlY29CNNSQJlY0XH7j
nGBwwQHUjngvpF/LfT9Ejc/uuOhaObPJ1oSRh2gu3vGIOndG1kiO2CaCZd95VvQeHpuhYwnn66vk
Q/7dVHyI3Fk3eCXX3ZRI/bmIgPX2An6fVHrqjztgMn7n1t+sMPCzPtdQYDebB+M9wsP1e/XaAvjD
TMwru9wOKxDBYE3eKMZLMl5AtDNnkPwi2il55pTJ0+Qea3SwPntX8KJSckQguQQqVyxWbzErg55m
1GnH7HHjAZ13umPBwSon7SmlziHk4pXG5CV3HAruFPxznIMmTzaAjo0xQm2wKkqLJSoO+OE61E4x
x2JxDNEW5gk+mJ39qfCTVJUPnNKIgwP/oyFpblDSBsFEkduXGukmYoEhVBar1KfaK7Zp1M8IxLAn
E3fSThdrkxSpj6CYKoY0kV6su6isiOaT7ym1+pd1cZTxz7X2bUyb2T5lHGYHEh4yY3UaWTMJlT/4
MgD6ZOk2+INmL/kbFk+1SBDEeFrGE1QEmogQmZkLZHE0KFCK0A4T54lbmpEX6K0nyYMc28d2Qusc
1gMHJCYV41t/zztStB0LXzquSMC1EA1SLQZMcgFkjkRkAqOjqUs0NfPYBf+A5DPdfQyZvpoTIeer
7JrR8j4GScsQ030xX+Rl3A8AfVpZdSiGyzbc5PvZxvW8NViaP0GNS3NUF48qLzIgj+79TTs/5nJK
YdfdCHVdNbT9SeR6Ym4UZExlWi8d94RQGQeIE1CGD13WZr2O5igX2KcIYKYxPxo2Cvui0/kJ9vCU
WL4L2x5cH647HXticvuZQB7XYaRR76hgVg+PwiTHi4WW+liaqmZTwfnxqA1fYbLSZebOrXPqtCda
lBavqgQ+iZw3rZEEIN4zM0ika3rPr5J7B6ET3VaXoyW9G8G6PrZJr6mc4/tVUcPbxOWggzc2zuVA
RN4xjL+MfGvHrDiApY0cAuhwAVwJ9GE8a/Gx898uGwYoJLO3B09bkDLu56KewaA8DZokjezUEFxg
QrzxuxrMoQanEsLHxtW0hAMy0V4C8x6EEns4wDefQnMS2b2IKlnC9MEs8RBj7ThInOKaSTz1MnWQ
TJhSxG1h16GpngFi4wHeBDwa5rqX8K70g1TaHHEDy1kwTP5c79RDVnzRr/DWrdrgxoglFArORJEV
NKBD2OnB8yXbPKXkUwilyqWfy31Y1AIz1giH4oTBQTnU1XwKbhhJHpbLjF7NiHdWLnh1GcV7ppgf
+B5m+yjbHytD+leiQYtopqly7CH2CyiBJQQTBk71PccxX7N4Fu+MALZypZaZuA2JeFOUiFpGJjsH
EhgTv3jzR+l1JzadIKek5GF5C+OWYNq8g0qZmyp+RILYqD5nsXpsDOoLVCPwkFectJWChlj1T2Qc
ueJvfPqmDifSs3BMqZRikbOlA/cqsPoi8srahAFwqWQgYcWYEnmiv2SGq3YzA7v4gvQIBjuLCWwM
43XZeUH4b/yPGzPdAyw6DIU82BJTyGHqW4WU3a0CZ1ZU++bm3yA+NDzD2mB+9AU/r5hqZrignlXS
fepIGxuYY4kK3vmtUchZuyq5oIjzpHN9AS50gs0R7nT/veq+nb+QEwkKRxoHUc0QycOJ+vHvBnuz
gb64zxUZOcmIX/3HA5PB8X63kWH0G8MrMppgk/waUMgPB5/UBdZFwCMBkvjQq1eHzdEoffx1NU0t
EGGkD3dnBJLEiE5YmPZPLpg/8SnsMJZOyllUczE6RS+p2aK+2TkwzY+t9jzAJGpBpmeOW+3anpN2
2iG6XKX9063i+Z55k+aqZ+8gL3fdtTaeaYAQF5qZjDW6JhHPe1T4rWgJsNJtm+hbAmapPiFw1M9f
IJP4Ws5kL6GoLZAg1dqhO0WvjobCJwCcuM+Um+5iIT8XbGWKSbpjWAQUqKD3OXkVmaxPxY+ZGkMg
LdRUoMuGlKXOzO3Qgosutp9hCbUzCQm9iV8mYFX5MemsIaqEjAwTgsBl9993OdHo3cdKjhDQAUEQ
hm0YvA6+7/nfrGbf1fl0HMHmipwWkcqhcG5g43p1V2XpNBGXIm6clTxHb/4O+Mtqx+itGjqzy1CR
5cwvUvbEqDNIHtcL9IhoJWAY1F/lbqizQ4bRlwIn+npH8boQTSYtTL/sB6dI9wAEc83GlDDB8oPd
PdIMjNSRKX2OTfndXBmn62CVKBKCv+zezr4bJeMeFf1quHUnlrO5l9WORADF6rcVPgk3N9YAPEg7
nBMz7u4s2IaQ+W9RBResHUs/51wGDXl5CuiX64fRNgNWEdEjQk3Mzj/gID4AMGFq2Zw/YiaoVB5a
scrkdwqG0i0oRgTetjfdnmLGS/ukmkpdrI8+qmeZcTntX+9GvyWWfYZxmdb7YnTAMEZJuiGH1m93
lFwCDu8PkyR1j1KJxw1N3YzgAe7JX8zmP8eKN+okWVLIDnUkkJfTYRUULUNxotLsbt5Jo82cbm5N
MzHlNNdHZ7eHPl1yc19RtcXCcU3X37oRuvjP1liQ9QMmhYJh3Zrt42O9oZQewOEPowGfBR2X5LlN
i7efugxSUlSnFa/d65lVGGoUGuqcgopKfJOD4HRB/atoC+zvFByWnpeAg/nr5c57XHz3xVq7tgnw
8IJhzbJ6tOPkza+fa9/fT+9PutvGQ1MKrX3jDl2BFqK0oPMDJoQlDc6j9JJVZYZ+gBnypVNSn2VJ
giLU7m3q7iGU52AVx6BrtMn11EFjDQaCWJx20ITIIAg6dLIumxVCCqEe0zIjcKOYDTHQt47/o9UD
9ZEx/yPRSRcyEL606yisNqzb2TDGWqDG06LA9/dg/5LFpwWjBJFWODDVUq3jMMqliwQgVZvgoSzC
HgTkOQVkc4CKhZGpTr9Hq1Vvs2tFBJ9sCvBO+JQzvuYF2jYjD9qqnvlec/7IFem9gGBWr/B75QI9
LkSO1gqnIQq1bAhCLOSfBxCgcTejuwFuu+Ng3nStW8zo4APZY9y4gklNyW5XutUMSk6pteTHXkMb
J754wEkOknG94pfsDV3gWyvAEQTKvIN8vuktPErMD6HuMjx2Xo1MKsDONCekZBshA+psyfz/RNpL
r+R9epUa3Lvxt1SBq+3uKSf+PFuFj9cbVeeIDNRkI6ZFE0avo0NlegcRC9JB7mo38ngIyRve2A8j
XAxzIiZdu4OgHhNsZ+WF9xQaNxVvWiUwOpZyGGQQY24W3/rqR9h9DPj3fW852F7Zj5JFT+LMOqIh
S9Dd1odeKpvrhYdmipV/AKxlirruHRjroRd/MC8At01lOxTrsaiJL+EYzFStmNv7qbvVdnBsuOFB
N4yea+wzj4knUZuNT2Gf+dDMDTtc4vte4OJcrSVu2GTLnKlmmzSbVQ/LtmkTo3nJ/X/l/FeNXcEJ
Z+lLZPdwgHa5UY3lBu5xu7xIAczemLZnlAurCSz0bZ9QOsbJCBz+selPGi3lQBbom3wonKi0VooP
6cvfmHIxKjMCXWjInIdp27G8QIfuZDqhQAPCRORiso+6cXPlSzuQ5j/fGoAaazvlcc41ZXRREdX8
8ueTkQoamvYuu4UlY0UGZ2dEWb7VkF+UvSqu4L2hLt2Q8dRqNj6CpvE8YjAcjW1u05E++BLvxMqq
rQdgqNDQVHNdMJfiOrnBlzPRqTc/wz05e8UqODaWy2rwjnbzNBPd+JsyRFegIC6meL2L/IjfecmI
Pa9g0k/2gotYLpTsOl8Rkh0Z8tdfdWCR0wV6r7KtUBwWtVWeyRPfGt5TD9y0cNJWd8WLep0bHExT
Emkgyo8qF6SvxrwSrV4/DuQlbRyXjCS3tfPi5vwMu+vaa9d+bV9PKgKXwT2KajTA4u+39ny19kam
Sw01sGsZ9yguUHgFfhsUFW/ptRuhUV1wMbKOUk5G3Rp0zHxEjR8Fu4Zi2Wy+0nxAOgoeGvveh/F0
vPXQRFmoLg+/ji1VHMIzEqqwU4TlJMYFn3gBWuExx4EuGIM9+8RL602a0hWxAl+LPzbJF+ybDiMC
ei+Wb00EBq14mEo+BmmC/Ky24OrVYR4S9DMbpinTha9KVvFZVYHGSlAznprI42VrvsloRaDYjOfq
A3oSVczgoHfvAwGxT5vLpCz3XoyD2OXT7bqgTrNlvm8YDbkOgwMewQHXcq2kkm9yYWc9LrHeYrkF
M1CT8KJfuiSUDpawbGQwPHt4VfF2i2M7gPzsUdsi8BsKXR6IrytzhfpRHTQ0rrhX10XvBiud5NHu
5qdVSCNJ5XvmvVjd/jrYhmR8xjjY8YjdixnA0EZD8KadLGtmmqq8qwf2c4T5tiVWm66Oo+NHicg9
ghvhm1XRj6r4/3j95nWAv7QiJe7mcR6iynyxe17O49/X0BWxEgrl8B0nDzI2u4pEY1qbX4rM90cn
ABd5R+014E63oFeH/wvx59JSODtFa5oI07KrrKpSfSo24IzYFKaIgFnDZKnQspzXst59tD5hgYTD
2DQ/iClEFUw6d6iBMrSyJllZOGbfDV6/Uz+7njilpkIsdZMKX/qZQUJhQXnA/hHzcqAyAQOYpPSc
hdsMablEXVDJ/Zpsz0YnazEdpvxh1aIuNbehEKqpNnor0mjLqnQAIDlfMmoYyVfh6sa5bR903nxf
wvVQGpgTlZ2A+csnj/FV2e7O5Ff5/i/7tGtjQBkvMu/a3TWvnQ23GWBUKIfQ0osUo5IT3LVYdnLY
gfeP2/fGThMGRoMM6xZ6lOpdMce07OvJmE5lXKdGiv2oBBapRL2jdOhH+KWGJGROlGqWEDeP1Ew1
EfUI1PvGNWVbgrJJ+2QYrSPzyPKNtWufyQGpjW0aaVRPGl3glzPESDkupAjZpRNZZ0BVcdGnYWgG
W3o7+lc3BzTmUzptxhvPPVFwAr6Y5tlgWSCJm5KGdgOlageNOvNb8YJNJ2Jzm5FxS1IKUqhdK/4n
/8X2lSBv14tqdGZ6gxtAyEvv1TUkVziu+nXvU76Lt0m6ck3vnDZSibSWNfMOjk7D7AJKYlEkkh73
/zcotwUkK7Ssy6zN0bRBODW9z0tkTUoNDD0UN3AUL0rwCZT9bLFLIARarpSWKbcAzFDbrRhMv30N
d+gfNJ3srQft9GwHimUiUnq1E/1l9jrepT0PBT9ETp2sXyZFeY8S+bFu4bxLDWg1t7nM8wKDhVMx
rEeJ2qPCYFEF3REQ+LLpNPxYGcYk4eV7W8vXAPYdjppc1uxvGrPuxZodtcqc8F4m0doe5EkmbfPi
rkaCZ+LJ4Jk2DmdgSB/ykdWytA1khoHfgTfDieqKHv2XhM47KIfbPyVjaB3eA58iJU10cOn+q9uJ
Kttd0EKTLATHbPVM3lKBFs+vjXf5WYd69Pbuja3lYsbQHorZIBeqrPpWdnXgX9NGn0gOML7bCPhA
CM4rUKMhthi8Y+xZV/7Nt7aMDWzZrRmVjFQj/7GelQnXOBfhcQejrr2BwHHB2reCgNHsF9JGiToT
G9Wi7RmGPUgWIVW3c68nS/XRzugUjhTw9P+58fogyrZcRButZ4wVwdlCiCnalEOO/eBf3/WU1NAb
8/zDkM8EWk0naB4Z+HvalhY7IH00woW4z25FQOuXkJXxkMj5ke71NhztJR+vCiUZhicMGIc1IVWJ
kSPxNcQOT960sY2h3EJpugAWVtIEWW6Bf3jkC4KahrqRRkpD9lGLqvqB697kpn2zuooO76PU2oFd
Fot3GK9/qSU0ty9ZWNXrGfsfx/lxGHLZVU4IYK+gDNVR6FRdSXY9UF+dt+X6LnJ4jF4OFR8xznWL
JnQgi574EM2hDzd4JTjrec5S6gpRA8RpasRpiT+h96J5jgFitKuRy/mvRwd2JX+Hz760yqZ+Q2YA
GD4/bhnar9dqThjOa9efmz840LnZ7WNNvrdNIRvZWOoQ2RQM5O0H3VGNxj/ki7teJII0eF3Sx3Xj
NmJp673r74KNHtUwssolzYHeHCXUKOjTBnLiyyNmXIkv9gjzH2mQdzzq9LNG2VymvNM3DKXiheFM
nTwzGt1McA3ySuCE52Imueg5FaSlCUCaC+p+InesBeYDosUxSlAPHcTWhy/u5Dzwe6t9sjgRePIw
co33S7pSCApiAOwO1jWFON4xHTb1+Fi+//IWzvSPmcBuuk9CU/skTiv3yk5J+69x1uN9HApQWEQd
v1zcDVVdoDese/vjKC9tGrxeXYRKiCXvhGivZBJMnE7HrSAGVWzGoI7UYiVKUHOe3IazNJ+Id6YX
Ftxph0ZN3On0LFWKwVFI3FRZRAwBelvG4j5XxnvNWVPtBK88AbC+sEmI3gnJTkEg3oubZEWIEsuD
gG8bIU8crJI/eaLCISs+3aUBUVKNEZUMgBDE6x2UzOD35rSu+uJ+2hAXuEqevingazcoXdrf5Jqz
/Jl/pQKy9OaJnUAcldRP7KFXooB8SZxVhnAHrYeloxGs3t9kZrY4cManlQ76pug86Aw01gVvft8e
f1HpzFVwx6lAgndw/4u2wasvk2wQho2vEDi5kalhbp5pMeYIpR4+MxQsVVr8027BOZdOrHJ49a9P
DI/3zKOPGoK2PDamvoNxv1/xUA3iqAllE0zsOE/HHCLL74DHZbQEpl0ThtNV62hZLG/WxWFm5ul7
21EoCFgE3acXLn2wy884IgRRL9IH1sSz+7UPaPi1eMbgv+FnHKqkUf+Q+UfPMwvVr9qS8Ljf8TEn
/lmIvIJ/qccLEj70mv+KrdgbFmNfjkvmif1l+7DkvZ4ykvALm2FJRkOawgCxfRxnRvT4J7Ljap1n
1impweQpRtGGQ59R6/dz+oUYDL9+RKKG1XHIYsOh/CJZSfptybOgjZBWdtmXUqCAglt1yj+01LiZ
aCo11l5MGlhLJaZ3L3a42QiWT/9pYqSWsMZN+bAldZVo+CThh4qy5ZrZLTBrvb8v2Ea3Rr4SYB6p
/ax2ESiJSyyNOnBjzTwEtvO7VS5oXRrgXFwJRCtNB5Uy5C6s0jVZcUfrU3V4Y8Qbbx5U4xowFMqF
OPkSEBK9pIyG9Lj1UvjfKT2BzsYAtHTOweE5/5m1IxL8KagfICIJBhQ1MPYtEz93CmGFZQFzto47
lLJQYW7V+35a+1qZij48IpIAje/fRlzmjv85N+NSpTT7+4wgiNr/RWFBhQjq3vyyAwVpldxxHMyI
ARXZKN2yDoVRaTpl0QxPQpSpePlLMQPkohrtVa49DO4VywubaNa5DnpI/Mq10v6TT77dRDarh/7V
CryLa3cq3XY/JEAoxM1PcFcZRVp7JI2KJkbjlij5+Pq+9tJWHcqrbd1RKv89/vmQ/BmbhUzKT70T
SpStlAxLQuIFH244/UdYpEI7pUJ0YOTvqMcXn6hVwnk8mD6qf4NL7TxUSFrNBtzdBJJJFF04kbOv
hSs5aHzz1Usk9R0S81GwynOq5CKWNqAT88iPsvinLaoa2iVE60WfMQRxlxD7Og0wmmFL0Pm13xfi
GfvMOzwFJL1QbOVaR9hlC+/rFkYmLpm8YyfziiMrjs4OLGSIgtnj9SiNUXvY7CaNKt6TJOG2BPtK
DXvGFCAwqA2Zhg979ZC3Id3Rrw1Mk79dPzqc+/jfJF5BryVb7wwKAI06LGTyMtJqAt1UNyRyK1Zh
rNgDVdPDvoOHhzEoMBxksY/AH7MCXBkI6PNedh/h7xCNaHcPJpour8iraQs1+qeCaNs9fuW0/MIp
gRU6rbnzPMGtxSAFJx4MavFxx7Etll8HZdSwEbvE0a57xsEWGwmozyFjWQNSkTjm4ip7W03T2u1y
/q6gfPUkDJTZ5DS8uqXlmp0BdeLXmF56Te1zjWHpt3x/Il+oEkkweq4X8ZLHkTlaAoO9ODxM2B9b
mwOPoePvque7crpAAe0PcrNjvVnXwGIVCrEpRV2agXHcxQQzDqWOpV+M1u7Ns3WymGDm7nnHrpXh
bpXy0kim8N5vDfUZ6eODqt18G356gdaDA+BkTUF9AzbAa1MviU7UGGpFtvYsQ4d1N5TBvf8CRr8y
zD62REEhw8iWGjrp9IkBwJy4uy+LSXWnE3L4q2njhboIf822W613t7028I7Z6hmNQfGR337x2JBj
dyoYfj0DfuDdrBwK+HRuVJqkEL77kn1Z8qLokXY9bG21liyg3yxnCZhK2gfq7jfG8dPT/Gtrp2jc
BS8/jWqsz8XN+Gv3UOub8NLQb4AHO3+Ba347BrkMn8HfcVtdEITTWEtpx7Iw8FPyT5QL8CmgCW1k
nWeJqy+aF4NarqQo28r7kUZtSyYA1cVB/1DCQoITqrSTkcIlgOb+Qs+e/8Djx2tQ2DZwewvGwjs5
fG++jb8BT+3Y9Vwfxl6aIvhWk/8V/IJXupakKc47Hn2shMpKBogME54fFp/d7N+pKvjQxmbQjgYA
HQl+WCgSC8cAjvfk5puMvGGCYTavg93HzbY9KPE//aaooFZM3GuVCmWLo/x5IMs36z3AQL+KXBV9
t06qtYAvIuUjwWOSCVNgHBtin6WLbI9QLqI6OZaR1Qfa3KS1hBo3I3tkW2eSe5c4/ohKHWr1gBgM
V8c/z4iGV0nCA3e00G/5tZIxhkxRHN42eUpvNhDGwFp+9ShXGfQ47KvDNSP/yi8pazQVA5duHktH
o/tXNKBXqXm8jQRa1iY8oSY4OJqmPJEQxBRY7T7+kc+aDkUfL+OFNYoqYNJkaWLgrCBcS3gc3qmB
y4S9uBgIEfDSo4+VJXvWofC68vnwQGiaY6rzb6D5rCNKZ5mgNLOgwdcYFnXcI52QJmqj5qH+iQuV
7GvhXBuBHoQ1R6sxToUNpGx2hAwyu3aEkckQGU452nLBHGvykL8lq7rq4vaPl2vWEyPDigqKw4RU
dmBupyvwF7MFPTp6NR/Bju1Zrkj/DQK2X/+ybifzI7SitfJvOhRI6zAs8R87KUuyczlGbeQ+pLhN
qdd2RH39+4g8y13PL4sH0TkrsYBcA8IsFNKHXWAYtHRno4uBnif8N2JIXVz0QTiSPz0dcp6vxGSy
XwlazCLUA1wnelENKp0BH22vJb5+F4GML8w+AO+1mZmsvQLbi4q9PqR0O/o4N87RbxXzBUiSc4lX
X1ZpMm1lazy8TtalydTgAA8PbOk/h1Q4zLQ5AcCvw+KVvc2rHarLcafbwLmTR/1Pnmg3MPMIRCOe
uYZfP/Gn/x1OUGqmKX6jq1vY7QBgGRPd/4+GFPtFDBogkA6od+MvKAXzpvdNLXgDnbDjME2/16dp
WGLH4oFR9ylkhNBSeH/pTH2+DIreANekB8a5VYrYbPmGBO8H86IHySJuKYWu93qXJTspUWyCstGQ
4APSqTlw6YmKddteRMuE4fM4DK6FsF0AcYx6jHTBW31SbtYQETFI21frtPdQEY/tiEMe66ja7ENX
b8xF+dP7SpLFLIB7XQ+wYR0+Sp7kbec87l/F8egGAH2DvqQzg2KyD9RpybwkGbB+Wsox0RIS1s0V
WJqiS/LvH3MRPxaDtXNV+Mexy9WbP5thAQM470fCWW8khrjvQVSr5vTQGjBUaBN6vnoThxKFR/dJ
FsFKWq/R1XYjjP9qbO2YI0YgQrfqlxMARCTa2HYmeDB6euH0vE/50SO7pvP4n79PwjNI1Xbmgfa9
7/EOjTC9y0C1GtZFdzOUpbNnrn/9CkwwRvaBvrHbTSdCQVw1tqGSJAQg6bmKvQ1X4P+Arp3u2r5N
bsasviDAd6fMRXQD9AELTrkUAdWKz/eeREppkUFb3N6/A8uBctC08dcKBABimviiaiOzcUhRO+Xx
UW04v/2bWP4Lx3Yh6RJmr94KCm1Cd+WiHDH6QZDjQk4HqZNZsna9MGH96eWEtnoU3UX5TKs+aPKy
Pb2zvoAG8mWL1ChsgNhd5hgw33gyp6bPHluChwvMBpwiH+bHjALQ6BqxuKZWQ6uawacxlhF2Hgjf
Fkdo3c2sN0EFJqwBuGOXcqgz7gC9/JNqgyZzIzwcRjCOmoLPA8YT1jy5DBlZAFcGpTpFmD4BYush
/hZIO1I1pWQo0yGvILYgT96sHpOmyMumEQSEbmSoVX3QGYBE1e3n3Dfw25XYT0qBE5zNpCD1gAeN
IQC4cpVQzI0pyv+1cs42C47vcx+6+pL2c16Z1oi0+9s2onav2b84eh1Bnfe/+W+hUPFBPx5pseoO
kYq3I/2u1H0af0+kxk00wQ30ujI1dgNQpPE8w4qisRSw4h7nHR44LQ5+7cemT37LSH7mKcDBgz38
UN5hbPQHMPFXhjTU2HBAWjc/VyyN2K+5Lmgtq7XztOj8JB0OVLPQj9C5kW9vDiisVqidhYj9QSyZ
i+41ZrVmyEUVvvypKnKr2QRv9SJ3mdVtJFFQRqNA7N/uJOJbD7OUmiYhmQFDbjR9LInglbRmTYaV
buvsmd2bgePzV9szJ8TnFPawUerainaDu/vwUSd7h2G3S8UlEqkX+cy1LbaCTVEXaJwB7LIsGwxi
dUcwjn2K1GQ7jIAZIifevCNA1YHV4dOenz2DB/i7rZJOqpm+nU47eE9hDyBgIuvJ3bj1IW2JlueN
BEzNcqVjGO87S9b4EZKDwtZAeuCK7ALSQvVK1kkJ0uhuaXtO2rPQNhrDfjwinIYWAeSfXyoMAW5R
6Go8lKfbEzEd1zQtvRhv0f7bpu931IsqA0D4mpJCMB11bbraex7ZVrM/e9mtIQmXIxLeUIMCKlIy
SEOz6C0XE50Q2DcoGro0VCIcOmSdb0o+mrMjGvN1vbUz/7AcOelcIz7qAfzK1TuspnMg1ozZZo0L
WuSZyquRffzDm+jvNfaDUC6VeWuiD+wV4LkdITkedq8w1FYDLpTqz9zKF0TPh8NymDU/NgqLf4dY
zWId5Nc0vBEAEZPjeDqlh4kVdxPu8jFPDD/rR7qUiKtyu0014q7AYIlfYr42oLc/g+OFGhMAHMqV
vqJw5HT5vLe4P3UVmsi3A+T+JMFNFBGBDvgo5aS8Bqt0MPosjMcqr4NURM7I3MfLs0rlj/TJOUMN
hqdVfFU6Zfgqcl20LFEzswAV9mQ57RVzaT1CNPFhVQDoCIsMDvT/suhbbcjVWWbO+oTAPIdAkLXG
IWRo/k4O9VIC/AAk97DcQTo6yoTnGRR3QhXqva8egfHrwTCvVcMQXc68accZ0yW2zHEopvMZST+T
evtvSslqnZues5sySc6o7Y51UZHKVs860UAOxE1aMA8KZPQDFSQmMWQ4mzd65FkwsuloaOwctjgP
SZ69+55M61t1MhhMnOFo+3qb4UV/YuxS059qsn6q3R5xfAfg+vGa72169tLNLjj83OB9kMgjExFP
BLSfFu2cuz+tMW9qgBKfHbB9z64JWxyJdYz4v2ew/kV5k0s+ka8uBk/VuBxFnHtya9Lz8wvQGKxg
QiVrwj2SdQ+yve1t9nK+9kXBgVsYQT2s6acjOYCrf4TN6mwhdSNDGoyUcT+v7ek6GLvnts3wX+Hx
KqJcWSTZCgTL063UifrtFHhZ60S3Jmpn7+BEzfmDBK0FlUZgKm5gYFsvtpLvdAil37nAW2/QvcMW
BLyyqwBHTGqroycM54OLtJJYH/rhIAcaFDBpr4Nufd8wgoJU4SAN51J5xK5ogb0iS438alx7JDkL
Y6AaHIuQI+BLb411VCmzXrbsBDvEiUovp4clreewUqixF75ag5v9XBj49JsGuHhjHyILCLk1XeMH
rCQysm+8VSCQhivD1RyIP5Mjc/p9AR6E3YCaKl1Tc3Qd6lX3L5lnKdbdg4QUz4VLzu4WavoGt0WZ
e2FqTcIWUtyrMRGbUdV8U15BGXBr57ZTqU11dcrI72fE2fa7AoajO/2hlTPJhsXwoTpGb0hona0u
z9/kU5i0n7KOE7GNZOmSZuckiU9iMC6VMap4AgAZTD1uzBITLGcMQlj9W0MRNtsCo0oE0Xnal6La
m04r9y/ZPrK8vWfJuYbxQPyzeROaPuL7UD+qBbbwpAFcGorAJK77fanryu1rxPOsXZJVuTJqZXU6
mYejWYY3XcjSij0qi9YJZcIMO/Entp2IfPxQdWad2dByYd7p4kXEJ/jxHit2W3MZhdOdGs9uKfyk
J5geezREpviK8F2/3RbZi1xZSFivgmV4seCRm3ehd78oUccRz1t67k27plbgNjtIib8IbEj+x3DH
/GjZqXdqLX94G1HXr1skWuqWVmxHWy4QNrhjs6BXBMGNpmk/aT/TX6RZNqymujPdZufGoyKTesMo
2j7nCZXrDImANoGoJTOSNt7FL3zsUdosG6Oq5duehoJdjIvi7IguOI1l0zdIxCCnICBy73e0rYKE
Gcbn7WSrhnrgCcC7dJbok/viP//4q1UvLY6dz9XJ+YzJgFGdM5IJ0WllV15Iv+6uGHAPV3vpbLz1
KqY3wX0QYSMGwxXY/dwotxiASqc1i1otbtDAuHwT5SGyhfhAt+j5dqjsY12KR5T0ux7XtAZGK82+
4x3TqR3RyAQzKfaFSwdwGU+kwqfGcZQFveux1erUy2v1zyiJBYizs9Ij8IUVBm5S6abLEUlAKQU3
HQBydcblRw0sGxI2OrilYhySnSLysU6npQ+HxItc0lNkTmDnG1qixpJpq+JSKOe+sMcSN+B6BSAR
t4VbLj0Xq2dAijGCMA3wwbwXnLldGAV1Nw79+dKYwtZ/P4odgPl263WtVmwLBJ5LCd5dcVSPh9M4
2pQQstCtgRtxA3Y8jU5FsHf2pKQL+ujrZb6sO0lV77ER1ovyP1HaGwuyKcIldZCbUyI25fF9J1Xo
uFXePRhR+OL3MBzZ93VbAC8MssJX0YZt5RbavM7ssrt134n8PKpG9maQx7V8GMoHHOUuDrF0tSJq
Wx10+y1tpKyKRahErKaON6Q02DrG3XI7XNDH6hR3mByCctnF4AsbOdUyOw+fFIJR3tGKeAnfRgAR
0Rfv8BP8zwLJEdO2yb9kmYnOVR5SZHqJv5e8BeTJkLTSshQyAAGzuuaNNsNjuhcCXFxPetSUdj8m
aDrPXO0D/y8iiLfY1T161hdk2EV25UQ68nZqZ331xP4vXS25lQ/S3pCRSJIOWU19VagYd93cmHkU
nSrSRxosdgad+t5VKKdGUsjj6Jl3MwhbSesznPy0Pid3nkIKr3Q3p9I2CVd4vGZj4iCgvil25EB3
GfFz+BB9Iq/Ep4ZMJEYoTbmlUf5SR9T3CmugDxr91LscFFzZD3b19ONYONF0XzHxenxLeP8NNlAp
fFTcmudzRLKShEHJ0doCV8JtjORGgafsjLwGy1RrBlHA6IowgMzgNCn/Oz3FUhem+PrAWfFK2YAM
jrabHGJ6MpX3WfJnV6DPCjz+dJADUZKHscHJKDffZv+xaYBdXsX8aSZYgfQlLMUqVGEAw7TCps8W
w1H8RyMhq4nbnCvW496slqAVzM5ZpGzNCMy9d8qqwo6In9FLFScjd4jOVk0PcamGl1xVJDIRfO8w
GNQX6/JKejQhh4lDYszYQW5BPAkvbTePx0UwBbN0JMmn0c9AL/XfDwI+QG8SXavui0EIcclnSq9f
sSOLEyeeifSn5T+WC+MhXHytVpudU/1JM8ieCJLat1Uj0xvl1BW2FFbruEEE2Wb+0e4JCgVQvl8+
dQaBWBAuGV8xsoAEoycMLtLutb4AGScainxeTAqSSajCViveev1Grli1ZMaWvamRLeYDqF32kwkn
2Kep//yF/9oe/rBZtk6eeWAd1T+cdlgD2bRaaa04LSZk07o+P42LOhQh2OGVUZ7G1+Oq7FLf4SbR
1/0cY6IWAESsRAqfxcs2UQE37Akfy9THU6xQ0BipHynZjqoLf/GPe7B+UuOcqcGZHQg6IqvALSMN
D23WdvTvPd48diKgScYWseSnxEd24bpDXSEVoYe5ZNmepySDgQdWfACvZMddpRsvme9WpQPVhwu0
TRKLbiwZP/TqUiM52rnlzVrpCoM07lB+Zf70fVYOrO/W1Zl3MP/zIb6Fc2ttSjlAm2DJd7CN1b1x
447Nw9sdLvDhM353rwodmw7HNhllPoQLBwL2dz9h+9hUx92Bl/r/kU9mu9+1TySi9GqEmCTsnxO7
LzXkxXJacrExw6+NCRnEetAEPLkugGMIB4NIJ/v8ZBAyfRv5DPkE6JmQZzQ5I4AczCqNPlXFakGg
9S14fIRkZ4QnfttsiNpFiaLMvtQh+MR438GOSmXQzSXlG/8342B52ng21qCLk2cKbNYAormCcceB
DyNLhxDWAx1ikb+fe9r3sOIDBnZewwrYiol09cuqqf2phENAnxQtvs7KmHwSWBrRyeG07MG1y0Yc
zOk3cT001YiAgT2Y+AZ/6jnwnY06JyRJAvb3nTeaEtX3hdOVAc587KqTpw+LGwTh1Sx2a6gMbD7L
er1N4vWZ4D8hgAhIPN3vxNm8ukZPlQH9mN92JJeXPDtwSb/AI5nccW3rsMhkr9SPwNe8Kji+4Rgq
kuppfTd3Y8iEADzchBQWoVidDcIOyOfcjeUPT2ZV5vEoKRf1Kl8yzErYmpRwknEGN2xuZ5WqM3YD
OJFSEUMfs6XB2ALaX8xmGtPz6nOQH9i4NZKhLRIq92TeGl00oBewwfoxL0MYg+BRQaMtijZciCE3
EE2wO3GgMt8pxGZB70k6VKgsz8OMpWm7xsRcmm+gB2mTibEIxGv2JGX9MhisAbiiRjfU0PPxkaFo
Wd/Bvm4Y3NJvbkG8XNvA2uTh3DWn0CV6XMvoC31Go6Ma0eUVw5KL5O5TN/lXnIqKxlVKSbzuz8RN
sjDmF2uF4TMETRNAiEH/OA4EP/ZbvyVPo8pvohTZSk0yVvtSmGwI4aDRg8CdYEKBAy0x/Y0qE8Tg
ikEQlIGXtl5a4kthFhmCps5WFln2NKedDgdH/3zwFEfTMkytPA9hh/DVGDl+pMXeYyqaROJVCPBz
+0YgwhDBhxzzk6zEMJzYlqcQLCYzqpFGwR5iuMhV9heilenN0y1aGzT1Y4roz8POr0xcqxH3m1sz
qPY1dWYMPOzd9rrymPOCopW1iSyhV0IJtDT4KcSEpZ22Iml+RZow3maU2nbyFa6Qj03IUYidqD+l
5hCgeSaatWX+q4MnDkve0uA2S03zMXvkpKByWn1jXq37UJwEzUM4dEeytT89MUGkZGYas4ylFTGT
NvLBPTHsRctkt0fBTVzTz/9g+nJVDyCcnnf5Xq1w49CGIti0Vf6aSOTTRi8Fzqe5PXOdnqDHe0b1
OsU3uhGqGh9VhhYuiOIjniL7oZwgfEANNYpSF/CXv/MKCEW8dRw4GjD/Y5iUtMDjftBVhS4aZoog
9rcmyQPLSaty7N8e+VBGDLunC0wPqI2OESF2afiRAjceXCsKvQkJWRpJol1UgTaJeHCyDsdJ+3Om
HfWlJIEDLBb+vBqjWXgMX9JGbkFxgS8g0RjgmFjq9sWdde64D+7b45NJpGi6bFcwLEyAPzpYMN39
nCO3WQd57+gcsgSMdUBuC0zlghUIJP0VZUkyti3GgjhyQKuKA5H7vdE8nFZshHfVJylFDgHgaaSf
3SYTGkEoF553BreOhMcR74WioE2hDUbrfonyv77huVgZ7BdOBxyntkK/Mwc7C6AO5aN7hwWONKLN
8Y0xGs3I3df6yWBNvnq34JE336imsbmXHaXs+dr0eJ/hwOD6qPChlthWvOx/ys31Mzd9ikL/pMZw
fWRNrIP4/eITMOhXUSBCvC1j4Z1mc14kLVJx8vcL/gYmznTTD3njMlulD174zn9ygcq5J38HgJ4V
o9BcEQDoWUq+y1MWcWPQl83EUvX29izR4JQyY+/hRqdWai6iQb6fvUUNGa+BpKP5tCPPtmdAagWI
6r/IeAzHBD/K1+b0nSJPzKOW670Y5kWe19IXFNPCpvBm8W6KbO5iDUqBeZ0MoejHY7gUwWjf385B
SUGKwNrdPTut7VJQVwPYdkvMw8aHMPW2Uaf11egzk1Vw/u87ysdFFerkv1m4fPZt+WrjHEDaZ1NH
QSQQNvXp0Qy1iaDsmt+DfkhDUAaPwak2KCrVUJAb49BirGetVKQALEzbKzHi2aDNiIbihIw/PlWJ
MfnqrvGIZn1fGBZH8L88+OuKk2Anl9YJ55bR12ZtZLaBErcuOeocGZ8ZKezwatNOkriz4i3Ac1Tg
ikVczwBhXY/d/cBxhx7IF9Ka80HT4L0CzFk5rVrgFFT+pjHcqn9Z12SmAiTH4V7RTKNL4tzS7I9l
7vqdE9LXNXTHjmwKFQGdEG6R3I4L6V7DBfYVrrzgrLB4FWkfqirQt4M4Yc0KThdXbfgPpASfUPHU
8maR20WOgnAXdb//FX76p4GKmlI7/qatT+K7oOCktyKeIEkiPB5XZw97aCn5lfp1W1OfCZUKQI2d
jIz3+PO+8yQ+g6s9DzYIVz1hONsg+yVHZA0WOGugsW3/Ks1bDeMWZ9otCzz/61gCLR/g075Zplrl
Go94pCgWCIBldlyEZbez/kFo9YX2TleeBkHxgoSKI7Q7vWdxNTxKlFILYSAeM4Cx+OdgV0DShoEY
UReoZs1axRUFREMWfj1hGSP8s2uekPLRCv23hD2rsRUV0SF373qBgS6Dflr83X41ZQddm/VJw73v
Lhj6Hurfuy+B/SngX5lIwZsGLS8LGwJ/YyDJposQOqJMgON5EE84TBwc30+bakRVpqqwDliLFS4O
Vdh05OoIOhh1QDwvgkoWhOvcRNQuISLw62O3CbPAJW+0IYGdhZIxtMZPA0n+lZVYp65V4qEbO9VT
rbazUqbSUAIyaPYj3eGjPVASXdScIT5KHW9PZG2YqM0Ag7eAPoTsPIZkY5pJ/+R8P01ZGXOo7OXI
tVxfcNiD/v15KIOPEJ8115AsNph5/HCW2AvqPkcRXGE0nTAqPEtRoNSalmmJbKg6ke3oPi1DbrK+
WbCdvcznbwmmWWvBSVEAesUvrnv/yM6jC/NkebCrhSHWSnWdCCtqlVXTECTvfW1DQLgesIe31Gvt
sfODjYJTNirwTpd8gcyUSmxE4E8adWVdpX5Z3OOCweP77mhn4QoHLtAPbdUUUCL4HtRM7RGBntRB
FhtBAy6O8+NoiK1Exwfth1QTsZOPyJkfrlJJ1NeXvF4eVnGbvRGfHn39WhELfyvUJb4Bi9/isLxK
o03+6kdXgVm1D/MkApjx45Y1PvMsJsYxVdGqJ403Vw6MSEJHzByvm7MkXY5qo2+HYKi0x3qO4c8X
O2JnU8Ye/uoA6t2Rytb7koeIqJWvCi5epUoDj/e1wIzjI4r632DSO8JZUXuBSyC1vWzcz8/e4Xm1
u2FjhpcwaAMCZ1iHiJF/ftVI4CA31EQ4a2FAYjJFv77yTUDFIuvcJe+gRxWAjb2JLqIgDZtp/c2X
mEKcQTHPGVTquq+1I/2GC68TNW19nkUEeNMWMdsurigRtywZaNxDNQA6ShtqX3LKN4lL4KA01UuD
g+u+5blULSiV3RVCNUQA79CXQHsYwAzrGoB0WHp/o0TbYaAHITo3u6BSvjpukZWmHZUooHys6shM
gOLfR6KYTkHqXcAK9bUindNsfZiMZQvxp6zgyoREj2iTFdN/g0rnnEHL2ITzlLEYgMuFMeaR8PJa
qsi91ZGHcS4/s675aELxSEBgtVD7BulslF32JuoVkLVyQi1xFX2wx7ZCJZ6+5ALVWJLGkIQAEzTK
7JjkJohWHDxobzORJ8rcC1FfK01sdOM4AcknAE5F3JSR3K6kdd90t9hxLESs7jeRmUYFvphtSmch
uKq/nnwhUlkcQEN7dXasnvbRAAXYEjD1KCfBOFy7Gvl80RzquK4kQt2JiG40twAJm/tdrFBOMA0d
LFCmYBL0fUnzPplWHVklkSuqAPUCYkp5X2SWNqZV6irMUgQa2T11RBDsaY468wzTEzD5WyF9vyoG
Jx1pitjTu6DXV3Wy2NYjtENBkEnkjxsplJt1musz+8Gs8JmE1Kre1dvQvx3aEkHeaSdVTlQuHcHk
/3wcs6P5vDSN6NRz7z5GNAlJjk7fo/SUMmj4+6PNbc5Smz/egKF5TJPiR6Br1GOYQPivZfudf5uL
VsIdlN5SZ0oK3pmWyAmOKzE4iHWIgwYfsA3bK52xoIBS+yxaOnjxP3MIVcYKb7yjLAkWCrBfOYxQ
fT40uxQPFh2DHyxyQtXzPoj5nIKfeC76G3DRWpozUJ0g11jR2fChyUvJV/O0GcLDE6CcO7IEqbBv
Ld9arYiUS9Xk5w+EDReVpfGaAddT28PovXpApLcXEE65MQ2aJC7BgPoTstCisbuyyg6Z4DHDbwH/
MyJhh8fIfapA2qpHMj10F4FYGRHTCPe7C7Wl607o5vBxk8yRSIu2LRBgCpFhBGM3MYc7C1zafBCF
vvXc3n9jNIADTeEm8nSPtV3IMg/L6Gd7LwDAiLAuexWNv+mJaKiIZ55xDbptNMFHQJ8o6Ggqu+Tc
aI/c58RTEeX3CO4vMNeAspBDoleLjLihnI8FpgANhT67ZlsY5Pd6G0YAIOVK1qZKqumX67mqN9IC
+RVPgiFrFsJLWB4U0AUDC4daLss92Rw2c15rVSL9EK4p4tH3hHE4Y1dyZU/q8y8mqerbYc/2ue6q
6N9/BBnXbiL/ZTyZ2vtVfhHPkVLbvOpc4ZdBo3cC1D56LH1Zca6BntdIUjKvd0ylvnGYJLxQlc3k
LqXNrvgSmW66u1TUNWxIXkPfxtreG3pwjXzCQkDvxKkE68lRA1nmEINFf4zBl61N7XEwKqLv/NBL
mqQbeFTvaHRgOvUWHuolMIheNVsT5LzLXQMJOJm/u2WYJxeaWhein7hg2RW2Ek4NgmTSCNUUTp82
UaMuPbHZID/IxJMEjS47O91CDryX29hpdJG5Vc7ZYIXb7ElAyFosw8/Z5+bEqk9IEmkpxVsxFjfe
/NqDv/mlnrXGdjnEMTA82qZFv0zgCMOkiP8bWBCwOxXSfp6NJhGE/TaOB1vz0IqzX8Btfc/eG2nU
vjUNK2sm1NfyHqkD6AQoU1jhxE/DTedAXCAHK2U0Y9A7C/rMcHU6Mg92OS54Robnt0Iiz3X7wqYS
vBWH3JqR1qy3oAgHhIZk9/qGn5aZDw3ZkWhTUPEGQCiP274SEPQhL85OeBXyk6YrdehpscZtUDCD
mHlZMiSi2G5pP1lYtWZuX3TeJbCftv4giVY47VKBW8SPfb7ynWsjbFj1TJxoWUksKeUsW+bCkJhx
Tj9QsN4r+fziTIFKFWtgBXCQV57XBNaxA9r2+cCGLufmyks8LHCirpSxY317+5I4iEftmQWNabAW
lvQwloyQrFUO/t6HqosOIDvI4gZ3EX6Q0Rs5KiR6IG9qQPBtPw6Q8tv2lsDnU+Fe2SLq/SKVoR/F
GazIIjfLBRdc3QiSyYmsfPCKgvmMuoWFolgX7xrMJTqaCL/OPK1kgDxZVrPjXiOKFit7OEXseGDP
bxemc814vg6FqDL3VJYvIfhD51kzFMSuNCzBKmc1B92ZBKzSt4zLC2zIf00oQxDfWrRcdxdz98oO
InKuP3MkYWcP0eYE1owGuKPazck81R+gin5LKZtu1A8F32s+1/g4kwzTPleVMerXi2iAI/xMl5R2
Soio3/SpHDn3/QlmMAuw5L3NI6ZhLq5tdnz/KYQTqtpifjAV2nx2u0okivgadNYeHDN1D892/VPp
okyB/7E4zIdQULTn9wQhqkbJ2aoLSdThlGz+w9iyw33QMtLFRiv2MqoVdk/PX41NQkyLpmKhhzDp
JN8u2KT0iwj5+Oe8b8+xgEwcUFV9SY1B3+GSKIxO9Pkqztncldl7PxiiKvKjAwaJjYgzEhUDlstm
HfQJHkESsIytVW0lZyEx/Uv6PzKufp8jQukivM+1iOa+yuFjsscwqKritw3SeCA5pncbonfs7xX9
J2lb16FNJfZweMzd3DaJwCWimJk3tiOsqMf1mMjK1BkfcjDrnwJWs6/Xgb+5b948VbsTy5BFEDmA
+mh48GMwM1ZSq8x17OKofWltd5CmCD31NdHBKubgdgcI2cXK6WBkV60MhRqNtbbPC4u3BkL/cDzC
+Ju2bcVcRUhI9k4cVT+RuTtys6a0a9O81IgjQlEXGMfW1idDpxS7mex5Xa0lPSAthsaMWXjvqxu4
+EWTgG46RybE5i6/xPkLeMUrdlMr1URUOSn7OE8qWiB1W1a7e2GfbuMROwGPw56FYMa6AuqVNG3h
Ey0/DJ7o/ddXraqg4Bc5juRhIQbSVuz8Q9GSiUA6mifn/RhN4sT1FZFeDEl0MfW3N7GPTclfWtuY
36FqJIKC1OSnjgItS2eoc7fHuP8V0NRJBm+H/m9++dZ6imW7bjD5XwjtsUZ0LNJnN70geUHhPSVK
Za1sVWBbeO8e7Eydy7wn/xIt1cNfAkQ3ohX6h0dvd/cZ1DUgD0RGXk8rilGnor8wpmFH5cJ1LR8p
qVEYYfaOW9A3naQ9/YDo60VprLyodsJOP1g2tze25Dl1sPe2iN6ZRvbbRfCF31ynOAtay/xU2alB
UznPpD10b9l95dB8MvAaNUavKNgJmKAN3Ot7St9QadUf5CSW3X1+Y+kvm2rUY+xanOyZEa1zx8d3
YMX+jbN+7T8bNMjtzEebAoUhyFRBme2Z6r7KbByfkERkv7LS7dKVr8eMt+xDnqYG4pac3xp5un6G
HBas+Lq3Ccl7c25lmCoSsIvr7xOFLmO3gYGbl4109/mpefSGjCSQOqBUYzVKnVgdn41k6VzTf7/s
o7+t4lONlEmJnC0GQSo1G2wQHshDwYSWi9Q4ZsbfEO9rjFYJWbcOzW6FFV+FXe5PLouig4A34jXu
GMJmAJ0Hmd+OYB0Wwq5HHKNtQig3LfP9zxsEtdU9zBs/7qaqZJY5IxBNV0GM1NgFZ5ihlf47O7KV
YfzhUw0oZ5H+EzrpPKNFlu36GVa63zzyyc4gyHkKUA+NiVDCSu7FGoiN/V94h+dpmYv79XraL99Q
VDW2SHnoEm1qgoNj+Vo/bE3Yef5MJFr+ImJ+bSc2KnhwPLTRzMtUhvZICQGfNBeoLIwblL127a4P
6mwgWWpJk6aNK4n74WZNZwPumMhgteDZz3SgPH7MrzmSrCcPZnjVhAWmfaBbLjMH+MroBU83Egbk
nl0ve/SSd1aIxise5Oh0VDE8nKRzmi95XrJwC44MGfv/g61IaRuc9N9OD1Q2UlpmaEK+30yAn2O2
KOH3/075s0F9h5yPj9QhgyPkmxDFxYItjqJZNIAlk9DTtjcqTWO4XVNzCxgSVtIlt6y9b8K+GQ1q
K0b3k2Y2WeA0To3NYs6IpiVpCognDvwP0GchZ49olhyYOncguoAXbcnLLiTEdqsBPDnVgYnQMYu7
4mQWII6dhTY+3nywZmlmVASSCobwr5Zxxb/MIRtZZiIpS2G76YcLswN5d8ZCRazjHATtD08di4TL
GuwxtrcwY/mwBAAJfCIX/qKBcl2eXqCj6wK3+FZgGFVY4i6k0ZJ1TBwMD5glHi9jXc/MhDLitqDl
69iqQYt9+NYRNMtT5OMhkHIIWAEIuGPURBfJ4TxvH6FPjcbxujp8Jguz2bbFZrO1ItQ/lR3jHS4x
I40xmpMuWRK/LSuU0SVUWSTaHqQK/ulD90VKb54D63Pl2lnUYbaCM5MH6OrbMn1IvBqsnGJ6Di6N
nE0cVa026PyAa5FA+FZCNsYxFokJMHEWbz/mALjZIISyV1sldoCKQZNSNsZdWDx78HvSDCWDY6yo
AkHqFUh7+0jZ2xXawPGI0XuSHgtn13AoDe+wQe7H5JNK+KgmRRRbW7frkkWbRadItAF0Sq8g7CL+
VtCd9cMjr/ODtyUH0qpVM9RPgdcBm1sY2hjZRUz5y4uMaXokmSZNjPFVIB4QG85iUG8XPubG4ZcS
sgnlxgrDYIPTgH/Y5E8Ko1P0g8e6gk8unGbm1cuCvrnhy3fc1EOydsDz2YykfONLIGuf8cC3W0Jc
j98HKb3m8ohANpCkrQv2uhjxb16mxbI+mwxKo0ouXfIw5wVBgTGvdSGVIkaQDeuoXHHkxdgfVkxh
f6egjw+E3lb1yQuchnDK8mdZ5eWSnhRZB4BRz/y3jrm+MCVVdJXtTppRrduweTbJpdEvAU4xru33
b1bhTKZkVDG6ZKtEMu1X3i665dHFd/ynnk57P1aG5gvL9nunaNh+LFv9Ro2qmtEH2LDmVMkyzYDx
IftOv3C4v10Cio7dX03hxQEc4kZxrW3LylWvUAzllKIXEufG2E7ef5psjPFZ5pUFKGNuNCn70y7G
FYV6ZtCMHVYKlX3Rp9ZCc47oETonkgeE8f+mfAV795pyZo5flmTqSjpkgI9deTsNjnllXaQ/RcXZ
Ss+WlvgEAg7MIbZjP4T7Tcg+/lc8+x47Ya+LbMBlbODbH8+6BjokjAUqdtGlPqtX9l5+jXO9NGYd
CYzAcF8T8VZz9IOJypy/5fA2onQi55LeRVBsfMthNrNFILFkGtVqyDxKCNq+S44hbenwUi/lRa7n
hw99O8Mc5pPUEFSznyjmzGm+Zo3GHRvqU+01+QB9gPbbyRfPFrmuBhroyuGYMl5Xfw7jL9K+uCws
7mvhy6ejT4sSn1hFDY9ViMINDIhgwnB7trnm5sOtjvPllbud7ltAw80k5AD8SI3+C1wvnKTjD/Ye
R7uI/vS1QyhpBYN3ByQmEcp3zGT3OmT0pkk5Kya6YYXim4K56Nv7zcjdk6Hn2eiTtYEpmdI4jHuO
+6EJMWyaMDV7ak9PTq+pdy7ddbiwVVPA9RcGjZjpn7+v3n0VkoY0LFrmPOjWQdx5/YmIy5VqR8mC
rGUXYWbokeX/7NjRn/47SdpIdftH6vQc3DmBry+Vu8PigfVp6M+yNSVdEjAlOMbSkUuUpTIPTTHR
h/TiFmZRRIUIDzvkqXzTfDIkjUvikz9rxeq68QA337RwVupiXat7DgwZrrR6Wb0HxYgzbCZxSLf1
t8UfeXrKyt9vAiiDsoh+ybBmgxoZjQQDlSsBsss6ojRUhnCH/M7M+Wj0Stn5TcdhZDlTmh8hviYq
H7Go5NH3eDc4KoEgR7evUvkLXjOodpWpndzAAoK+64sBcO7WoRW6TkSwiaj3Rfdmex4dwo7RrfEf
ZtVHrEmXGloZH5LA8UFY25495SDpZ4hVHz7MkADHWHTN6SdoJVZsZOiJYAL1k4OSkFv1NiO8iR4x
7omhSVoPB9yPgbUA2xjFmlwFcLoKYCXSexK4xRcSgvW6VlSGw9TUMZ9MemLwXV0P3E50H+dlcOAW
fb3Gnou7YZ0J8xSuma8jbnRqntvevNx9sb7ejHc3WO0XXEQ7LDwfKUaUyCLDjU2w98uL8q6qANx6
U1Y/ea2vQMxXesKZOkkbrt1HCf9Z7gVUyRy6wyePCvFmNbzows7BgAqMSTbQb6E7VcZ9WmQ6W2bu
CeoRpmUHLMXo9MeHk8BTnTsJ68sUEun9vKJRRePiT56cz9wNzk/ILH4Isy89hZ6nglxCJR0c/7V2
TLXrLlPM//vmeXSFGnE6pk+hA99VcuwbtjUT1VYR9LEl6Lhcxenk5Zuf4jEjMZzmkVnZoUxhxCD3
FGbXbXOcC8yZTm6DWFM9jy7/ElGIhyVwa1eK8Q9yZ2HDYglupgLxsNBvoGEL2nyb+UrWdsD1BSTu
eFDdVu9HR/96h77El5koiquEknJrZOTOuOAR1Ds975MUiN3d1ihd0sqFiwiqjY/ZDK1Gw0I7vX5P
BieERAg9na9nEnjZhwlylvz8KIJRtZtQWN1cyN2CLPAKhK65epJq/czIm4W/uo86CsUXRKacC7Su
qEbktnLfKZQ+lorziCd+BTowmyFVOquLYn/adRMcFWN7mCq2IFhi1wL5A79FxXo4qmXtqGpYMqtU
hYgS1krzrcc+RuaZRmVjiGmkSf4c0FsZuGytxYsfiqAhe7ZYwqHGIh/641tnUn1m/g+cY2gs5fR4
5cSlHIocnLc+VGvbzcDKiLAj6XRNgtrngWB3Ay7SiwCUATJi2GQ8+4Ce6IFUH8zmUUHHVXsm2rve
hDHe088F9swNkSJMh4qK2cpR20qcrwTl6Z9/5G5p3hZ/BBcfYnXV9mBvHpwnnK88FCXmrgxw2bb2
+QLDAB8FHdz93L0RhgXvRwuv4wuN/nvy1slV0RkzM/evZsahhlrvuQsyhcqqUgznYQbNMcQEDzxK
WU22MjLAeXJOEAcWtctcKwr5pIf/qdJB9ssc2kP7oAZvLl53w06+gkuiH7QaEyaclzX6LT2v+bL2
p+ndinYVFmDg5e5cH+D/ueJUsshXDiuKOTF9Hip0UwomTTQqa6bMTY2zeqYPlgHfIwQYfKaR28uh
Kc88VdvbXbtdtwpgS67LxJStUY23otF9tuNLFZNasQVYgmW8x1MZk2I6x3rTu4yRiDUOllC4cKuL
3vziIy49PHNuBw0ztOr5FTvcfMRra4XPgZgkAQNthOx6P3oBbq+QVBzhjMHlNu2wXEU1xaPHj0EM
SRLTKQvSepI14tIO6ZNQhmivuTAT/blJael1Gg4Cs1mGPUWxO99Sg9eiFSsrDGbAockpfxJflswC
XP0i50/zY/yFTDDXFpog7LGfR7wIxrOWsS6i+9vuEzGLcFldfFBLHBI3E/RBpIG6C9Oz63stuPVx
SN8yR+W4jUmxF2pFR2DLX/oZYjxYUcpnKujTfslzIX845jln5IDmwLvpXoR+NFNDMFm1QwRuzDyv
TAq/QrP4k1Qt3f0ivDbJ3wAo+vQGoO54rCIkGOF3IUA6+3/aE/gzdivGQPcQGbGE20kFplDlTKpK
ldNCFg/X5k/rUNqEWYGzO/ARvvPcMaXqb/GEznZ0Sb4470o9s/ZaDS3/hngBSJabqUoYpXbjiIYO
/zoK+rTOrNGjTeoBSXMNqDeOYOA3vVUQDYKyPgy8sL77/MZwsOoTuApItXzjSTsDsrMM8MZneZAM
0902084GCvb23f5GPJWd7BnP51QzriHFw4/txN/8oAtNGVqsV/Iz7kYVpqn/oOYTqg0tAslQSk7L
VIl9+sMexUyiAMtPOCy39JJw1rRq5YGpf5lfSWibtBn9HbHjah0wSHXz23sHuHasrx2KAWMehRUt
FJ907mSCD9gopRGsDEzCg43cVY1ZB+GQhXZcaVFS7dypcG7WprfdYa+5NQQ5YWsBwuvQUtSGfiAk
lmcI0kn4A0/t4pPlD3mcsKc2rIH/siI3Ur4aw7zHlhU6gKcG3NcD0/0+h1pR6nR1/CQSb96q5GUR
tSDa2soxKKkFAHaNCtwgIB69aPvLvziyFeOGmgX7P6GXKF4y6o29vV8sTwXSKDyi+lnVJO+Pz+7g
iExorcTiXCD/eFRtw8Cx1VTWQA0q2uDnZ6EscDwklsIVLTv08eE09vCHFVIjxLuoVRB3+TgNpwIs
wdEoJM54DXHvXRUxQOXmiBPEzkiU1csZYjfvNWqcNOAv0gYgLuCw7vy9WrD18/4jRZuJUC29Hk+b
qNbsXXMd8sl3ooAiO4Wy90YJ61nOuIE+iOliFb+E8vcd/pwdtOpeQPlD3fxzMeSRTd2JVsoJfkKZ
5qnWAN1avlGe1Wt+leab8fxvlXqfbvXw5pBrI7SyhG+j7QbuEL5tKeN3QfEUCurPrUWjrVIw5eES
xMHAwjnFtZFsD3rc/GIKN5DzfzkyE/tw5r2OcgBfL4oQDUtLtL2hqZnyd2O14UMK9ru57q/65Tps
zmW+DBNlkEVkbjbsg2tWl3b5vrkzzp6Wzhk76xyuffR1leieQpP3CscNikmg3wXlF+Av9xBrixWO
dPV60ukLwCe9CbNrt50GhvCGLbkxyvkMwLNot3g7YGcXVSOYx7lj7q7lNLUgsU0eqLI/eJvbkGlo
qmHd6invuqunB/0iPc4suZ8mV4tsArl1lV1MnvnLeQmTOyTAyjs5rOVlr2FL2gro2+OBKVVUVjnK
m1fSVzG9vRZu760R8fJoDU05Sc0c6dh4avVMM+gI5y7pnQ1NbVYOaABIuvEwYqLIu1YCv8iwhmKg
JDY7Xx9skH4lIupwoLVWEzFmcJNuWfrtDl+1+aRKy9EWRB2W8VvKtEFYM0vIUwWURiz3Yd2I3XK1
5n5Jz19SJz+FbHyuRspCKMkL5tlREhxduQbAUTyhHSB2JVywBxehoUcQGXDVS9XLSF/urWy/CvgX
Zgs+i9s0YungcwCIpbRtW5L1bly4tn/S2wEZJGD4n4oMDkfIF7ju6SPjYo8n+YQk3tLj7ctlb9pD
v5dx0sveQFqTqW1VbTAYBkYpsWbGpkAtH8ACHF/VLUqkl4m4KzuJwgbov629bcLvgFaJBYRkbRgi
qujEuT5bD9j/g/+8fzo1fJhu/vCztqWni0FeouTyaQycXXQKFkFVk4HY1/OSpK1GrFlRPURYhhtx
EhB5DdiuzRXvdK3/te5aHqk57aL/KgaTByLHA1nN4oAE3aLPW6oWkD7NEvIOADjJv3X7fcXjqQGg
4TZIpyIOuyOk6OJZDvQjogeQtVv9JDHaL7KLTcL3pvjJ3not20nDM6u4MrJpg0pOm85wWRZ4T0mL
yqbZEUQAHwGrc+cYLown7fB7lamY4/9dj0GzghmMnzdRkBq877PsbFI6HA414i8bOvbGzQrNaAbd
IjUYNinVFR8sHY3nR+A//83xuS+2QtN9SyLZLaFMKTpwVziYqKYizKg2ChrUBqscGx/yce9TCyNY
OsWoWICpz6W07WH+BpkN3B9IfpRhw8OfooZJXS6IYjhY/1Z3glAyDvXjtUkfWRYzR6v+HxQY+iok
qcGjOUbOLRbONjWN+QaD/Bt1a+3L0i2oxUFTnCt6Z9c2v0K+bFE8GdAb0jvLEUVhZKP7ief+nM+e
NLQ7a23GJSvaswz2Oi8RrZ2BsZBjnV3vBuomqRrC5JFLAhI07sv3Uw2v4cPyhEtaP9OwwxuKApfQ
bvcTnXomFQI3nr4T3zfeCAOVFRe75W4LGSVNbOgixyAIQ4Cy2lbw9Pp/lKN1OJ7kp6zHhpIgpBpA
wRPI94CWLleyLLfi/yu2MFDm4U5fKlr8cO0EDW5wB+lGTt2jPTNHOsKIuFrGIUn7/u7tJPoDs5UA
BJqgxxGOPJQWpJcC3p3nUrjPkn9nYrHSYNrL43FvS0yrhL7L9dgesQqIMYFoWCqjlAQHON8OfWmR
dEAeGVxiIYcNnRiP8r3eX7SvQ2iS8WITIZxT2P1ke+ZXnAnhUxc8tC6x41JSVRfRp8CjqZT857nq
JnaGRNp8OkZJ8gcXi5hAjtE3naUOmgK0g4CnixCQGjGvl+jISjpWQBXSnoTF9LsGS5unKySOCEeG
MenEzWk5atxvDX2YvigjWRIHfTYYY5yZ4UBVjR+ZGEzslqOH0Eq+YlxFsWu4vT3TbKVYpjLrXEMy
DulU9KoM5HvvB+y88W12tDYRmZHdl+pw3NqhY1qIx9oFEQVFeJO3MMRhnFsd+GNEyliXUzwzEBJH
tnZiQwjx5Bn90jEM1u8pk71FDKqyh31LyPIKI/+o8+KVf3SJuQPVNUIRpaXRukeVXw9OBDJhYSms
L9RcX3pR+5CcKF58tBRJ/jhPq1bzd/qsd4f88FQrX/XzAp+d1Tj4lave4qKHf/ZB9KjxiLaX68w/
FF8HvyGuBbP0Zfv7hbnNBfUTJvFaa7eLA6WEKvZBofjr5Tu4OxhpIUfZtVJIEEeaAVLa8uPzmpEW
BVy0e8XzMiismem6z0UDDFkvBIVpPO+HO++6so8Uti01QuAAQGAE1y0+gpi0eWg0pyfqMlsB9gck
Aai3efMw25ndrZ3G4Zy3a6yTkeqfjjgFo99vvut2EdbBGLKfrXP0UoKo+Q5I2u7F05Cp/e2iISr5
jnr9K3c80nNxwsABL8vSEo8H8wTqk1vSwGSEoEiXFUiaCMpkWNFFKrSyJgl8lvMTN8F69UAZ5m2i
whXt1YavuKNxxo2kILtLY3MZ5O7GKiIrxOsvFiDgxkVXYNEfdeHbyzhFw0uP2LCjU0DufXUBOfdT
/3tGXgiMvsdA37D1pK4jbA+GsuFZg/r+00IwvVNXsWtdm5dHXSTXxNSWPhipWJywBiYd3I4rl+4C
RC2nGTpTssoaOELj+n1h7dL5IMmufYBEHyVkCuITDaEE/wTPJDaxMB1u5H3jvAEMo1gO31jVsGyl
T6gq3i/mAqMANXVld97M47c9rAVu4+srrMfZZy1ani0IiDqV64jCRI2m22RPobarFaiOxOsz6lzA
UuuZbKZZOg7FasbHzOGRvBtxIbguP33E89dJAlM5B2gMrZOzRbrjfR+LNj74PUp3JSzihxHzfOXy
vhjR8NFuTeYUxPLTyEAT/fEmxcsIi5OCbeJAlFDwrewcJzoDUt1xTs6kOpc1gnQeW9MkONZdswfw
KvAOdejTFIDS3ipHUMGFReK1nuGKvO0+f7EzEnO07pfnhiCmu8RsU3U9z5rjyauKFt+PaNovUfd9
wUIoSBKJeSqJoztwzN8Kp2tIe1KVDrIXQyXIZhVGK4u5t9cxsiR9DfgGHp7NfL/dqkvfADtlqj1f
INU+/mU9lN6VQd9i7i6WAE6Yinbv8eSjJ3W4aiumnAqKloke9JnGoJsexz59zkeKW7TWXYmyBEQD
eZ10K7oJ5Ri1ozk6wi/5SPm8TpGCKFjicdTAB4UI9RH59VnA9d+78Wd2hWWaV5unq675xQFq99FL
tN7M3l/PCZciVOHXXazL+5pDBn2yEfbxeElrzzunG5TZ7Tpe9CQWXvsEjLRmWwxYLkFCZZr/v23T
wGRbKZd9ssF5O5qbfe7M4AlAnO1DCvBKaHK0BuJzY7Ew08pCKoyAutz7pPNzpi6mCPZclVSlU9cn
dUKLrXhhjnzWRBQJtvAUGdKCVTe/KS2lvepX8eIf+klNIe14PbWLP01iJwR5s37Pf8TwyrUh2vMR
yJ2Ba046Lqg3d7F37OVYNPDAGOvvoboD5epQW+0/gZ0xX2MwsSHoBvj0mrI4XI2WtJj5eBkr+9C3
DNNUJun1e338TN9644fJbYuiqB9F1wIRNbvIN8gFdCsof3y3Phzy2g5zlwlryiUmLnFAzpv7q7yQ
9Blkv9Yq7ReSjCnG4GPkuEeiR+YIsW1ryYFvMUq+whTJDQFY1yuU5dizQFEVYtl6dmNviD2MbzCi
z/lNrpMhzxm4yopz5BiA23Km4MQFkp5WNaJuY/HSn1XZhZ/jCarmKhVwWi7o+KgVUoQnx+Ar6TBp
LN3A8Qr3Hv18rn8UPZmlNojAddiw+wOjlAm0o1mqfbcSVKGmjO291/6M76boGfqotjsT0pK+VG7T
ZJbPC7OEC83VUj/dRNEWfrxE2uVYui5v7omd4oUluNypYExkSuMM8WSHEReL0QbXff9rWzC9vXBU
Salk5WmZOKvJK9LrMNmiIke0K/QiQsFewElUYgbxSjrjxjyVOX+os+2GS0G+PMfrcQKDGvoxJq3B
mtbs+XTNKU0GpxB6bgLRD/EuNyOy0rVGrDrMQJT6w/MwaV9ePGz57OWgvRCD91K10b5LWZgIu3DS
nN7C+PTjvDdlTdokXdOb/3X3cC2xRuvCthwTl7+qCsP8HxNZZB6bt0/BCybawqtV80H3SkNvCNkT
exdAfjRBw8VVrUtSQJJQh3Sqk7TmcUbg+9nubCZPyrGuQbg090qHfcCOXRRU7poW46HEHb+IDlXk
pKGGWxQKep8pPmg0V0q19dA8WWt94VB3YicbEHxqEOp2vF411IrFb+TdAX1Eux247ZSeDezhAPlO
plARmJm+Sx//B33vPjkttDo2kuYrEJoVC3UUYlOaKucAWnXJsiN5rzeiHb5yT2/Ul1CZoq//3hE6
AB+1bpM/bbETiMib5y6s7wFcC/3qG/+MpbmuGOHZpluZRcKHUbkSpvN5TzYFLErYMhyxjAfDgu/j
9PVFlsLNc8KLuUkNIOhHgDCRQJAVjEuF+u2001+sDlOgBIecjmavFOdezpYexuw+gN/Lh+jvDiYX
MHoJ/pOhEiP/NYOJncJqRC0rVMa27FFGoXSjceJrCdYbL3eM3JcH3sa3XWDH79CD0VUL62sL4GND
W6Sgro+yDDKcDDB6HXvObhRQoAIG17Te+mamUVdBuqYFiV9G30ljajiaSFaRNwC5xfEFr8mNzEDx
y0o1UwTnOh/8rwlfKj4oIT48ng8nTJRsqgPDfZfEoE2wKh0fZtKuQHRlI30aTDM6XRkUFHrR10hC
Bf7ZwGF/QFJHqUsAGPfhUePcbBknVop6EkenUx8UCEPt4U8h7bA7fC5UpTWAGfTVlnVuRrer4Yvw
qrq3E4i1ZVp68fGV0o2k9T7Lsl6D1qJP0/8rNv6vX1B8PTc3al/h+20ziKpqVSceICL4wu3dFHji
lE5LFhPzE1fWABcjaCx2R7DIHOjNjJ9Bve5yCpQk7vzxTyrR+ArpPEc/loklLtyhpjdNevp0UME4
p+G9OcGvJtgr3Ff0TVCLT+d4OjuSHPWNFm3Jju7plVY0Z+x3nfHnJ9a0IspNR0PQjqdim2oUcXLC
kTV0EHyTEPlv9n+bgsCGSxZ4cvB7soG0zjGJptw3JmQYqfVOIX08NzJ/TWXhQPy12kR7BCEuE8DZ
sXzSa3wgSDP2A++tFBQH1RvgR//xK0vxTVUDeL1BSapwum6f++iNCPBErlYCI+guQzqxHprkNdnB
4FHGTRu+7Ce0mpZSRRzE70ly46gavjnmKTrf2C365hRSkq/4x3Cv927xBXo5T66EcvdULTbBWx5g
NPyjKWU9FqufGVakps/E6pkT/n5mIYZv7fRO2fnY8qbZwgxsGrQQsS7BUUWfaSKVPVbAyJ0zd9j0
2tiVp6C1LBUtBmnB0r7gSV4XYDLIJSwdn7LUPaq2bdNEFhDEEWzqwXjPXXhV8jvzwkEXMcAKLZzu
VctVA5iVICg1vXWQ9P8UC8Zs8mywFZQn7tr7x6sGpwYJGlblbAwL5EsCBBiULAEcxCX8D1ZHhVxK
NdkQIVdcRFf9BZIctIUwuVUkytI8D+5xIWk981E8No1ndyizy4AOB+EvbGYnakOeK2t3HR3SJc2J
thuQUzgzUSfzonazQZGZI+U6ZI8Ep9mRNijmq035o5OSi+ONg/exZAqc0KFXs7CR5jKdFs3Hz643
yKnOjMg/GborJOzVcZ1tv7V6s9efoGG2/JL72g9OoWg9UQCNdwrF/xptT67zcziy8kKI8D8U1TXZ
EASJJRCSIQGsP8/K1ip5K9U90DD2WP7tHbX1DGrYxcW4VvLjIdC7azp7TWQICO0PXxzxbzIdakY6
6094P1B0qvziryVIQ0/7+g+WWgN+Y3xr5WJ3d0P7yqB4BDwjFPRW55Nx7Mc2S8TkVrJaIw1d4Y5P
jjbp6WW9GCs91Sxc2Gl5zgRZc50dv7mw+XLqkyku2e7F1K5aRyB7kj6L6XHfS5f9dLOW5VVnC7vo
e84i+x4Qerq+s6egCJHJ/JFG0vPXWlH8yT2ER+AscMVIy45sLE09xvSrECD9HACRS/3UNAobpWvv
bwfooDHkGT+0x9d7q3NiKMoZj+uJGeRDbLrtO0Ambhg0QnaeUxkMNB8hCNNvQCFH9p+eXpC+wmA1
ycPFNDsornPIVc+Dvlb3xjeoHFUTn3kGot9TLIUK/OYeoaGWgaqcYq6jNY0lWCZhLEBCtTYvQCT0
BJLIZIT2m2Q+awB8dM5mBSSgyvOEMbHdLzaHp9URd+5iaeZIo6YFG7Kpu3BkmB5o2eHoPkInhX7v
GkEAlwrKuxpkllbhwFGTEMCjvBiyVkRHO8IFbinjhuAuG71oljAc/AtyYgTaOYC8EbSQQE84EPO6
rjcnp1whtZBjjPMhULQgxqIDcUe39TKjCGNtbi/duY17aeM/mR7Brc37oDh+BSu1X3arTG+RYurA
MHQP6WC0OEO150QDZIpaAq/Z2G72EK7oqk9UvAbmDbMp0nHum7DkONo0aXUohiLv0S6Ijony2HKr
x8vo7LOv5KvmCkjS9NiupIlQleAGXccBgN6rvdGaQLOybW6RWob7o8QVK9exxVLQi4lQiRn55LfC
xDCdfPAsOn1pDGMNF5JDAoPhk4aqxV71JQAlEinuoIT4E8j6E5ohkWx5j2zKiGRp+TwvkdCzLn/R
fWxi1UB2t5vTZXkdENr+X3dos2X2Wp9vKX3x0pCDUnBRZjpC2ipVx1gLk5s6Ivzsn1uIcysdHcvH
VMD0TsBPrJ4moLcGh+RpGXGnMeXhrrbue3t9PplplITzqz/5dGvBr/5YASzBYwa+ESlMWPHCLRfY
k9saJB8NbDB4DubcKq8lDrExevbjSvQsv3RNUQaLWTfnXcAz+nJfUYWW27FaFxUaaebc8VuOd7JW
mQ8bIo0yjDADZmqIR9giwvWje59WyloG53LdQmaWq1Q0dsim9t/W6NL+Dfqkk58oTbjKguwK9ggz
OqeiB6upiuiPZpkqORJnOm+gVxIlpIWVl3dGryGpUYBVfBClZIfaL8rMc5RSkh1wnWF+abUG7h7/
/19PJnz2Qq+/N+EDOLao6h2KB/sipHWOQc5FN8UK3eCCKoossS0P+wQoeOWKfvIS68+xAIK7J+kt
s2kjFnEYq71id0oEvIQj0P9MX5SIwuSPAKKwWaF6ROQ1DbuUPj0sEaJQA9BNntz4iHxwmSbkkloP
H2hbsUJeBLl6vd3pX1OIwxZwG6J54k7CjMl1/fOC51pb6lbUAp7HHcjlBkA9OGzHHhgScdxLHtyk
lRnn7/N6+Wos2EGKhQa89QaEUkx2G+j+KDdRZnBrpw4xjtX8ebuRWKEuzlTkPV+zQ2LlRMEnVLQ5
Dg6khUswEVGaPzrvtZMA7t5qgTpGDy39ZXvcik3LqvHuXlYsrw8A/ULk40QQ0F0ECD6bn/Ixhroi
j12LpWvklOcBFBoGr2x5T+J3/s3aJ7JDNvCZcaL+hJB2J55dtrBrurcAUJCk8BK9PGLHXrnFTqvO
WwK3dkn8RG0nWicQkEAnLyXC6ApY2E4iemMTsgAdrXvOeJUJPl57wtRldQyjEj9aKq+qcbbWnhvu
h79ZdtlhVCiCo5CNrWhrlTWdlmWwuVQBks4BRQMq5b6Y6C5xVTRb5tpw9qet2D2tUMrrqiQZv60E
kvFMmu7UZJ4BSJi/QUD3lwVlWh3+LXfjpH7TkLlWu/0xbwCDB0xsw3tPCRQwE2qUoyLRCnWPZDEQ
oPclDRSXFoy1qTalqS9Qko+dQcqiXaKTFfB4AnsHjmOvbu66RJGCGa6Y5lVHJ9GVZzUCY2MkkN54
mXmUt6i+6fEaowucGL34+Duvuva3fcviv21nlub0m0ZIJhg2vAEy8E6GMUulfcskTQWHbSwOZXYz
DLUsHUAQyUPEcGKsWGo366JzyNJRSum2XHUfna8NhdK51xs5iIvxfNajdOtG1vYSCvw3VBYjZrQR
gFA7bhfB/bhCXVlFzwXgAIVs7akF0jsX5R8PIQQk3EbYqgy9O+axevVcD6580UHxBSyqUgpQ/eUS
wEcpBfb0yDXx/SuUVWTbs0G9ZHofCbuvOSBKnG1ERytNYdV4HIFkdAiESDEL+Tt+liWLpqVqUMQu
H4FK8A6qBiqW+ViL70vPqABJAdeO8zP3ouA+JyB7EJzwVjbllgrfd4Bt91dl+RctEPsArbAw1bUq
hwnUuZ6ttXJ+e92nNT+SOvrn4C/nGICHISR+x1xR9uquiPY5cpH2a4d6iEN0UKtjLHnbY8JgAypU
otCXmWuljs4dxZFusiC3uekIetpCdTkhf7iq08cx6Fs4i9aq2dKwlZiClrb9wfeXJXUIH6chAxz8
lvj9hzskTNGcWkV60eXQyXByEUE4iXzTbky+iN9lzI5oZNUEkSHpG5vZAQNTSnXEumZvhcWkywuu
bxIjDL3ZtW/5/RSokQs0pRUF4LUJixMA/V9XLlauaNyk3jBxVJERaLIwwOfVRv+euzx4EscdXVsF
UtbmrdUhXmJoZLB58qWRi4aaGsGcdCRlxtGsf4eUkFD8J7EujrCcNlz0iKRZK2ROTJJ5aqWwBWtN
H2ymeU9scjizbcawq5QLiT2xdQi86YA2C7qg0Ir+fHY5TQhP15Hthj9kQZUSVXtK9B2OB4DQcVtL
iI0t7fhq/eZCWx1tcWk3j+OhSdNDyQKob66bgSxHJDz7mpAErMTXVUamYQN7WJ/gdOuBIS5bjPqI
nDF/jNRFx2VFoerbnD9MoF51HJKuNtSSuzoWOYWemSTu3dSAfOBqNtRRqtE1m/sQQ9+XqwcIC+kH
RHPeyrzHGkKe6y5pKdxjl1CDHpk1iKotJYlEFyrOZBweGm4f1YVJIY16e5mkLzr37oe1JASa0ci6
l0UUe9eaTOUkZNK8CC3fcK27PxNhSL1m0Ev1QS6PITC583GMMu1PKki7huqIPlJwsrMfnc7Jh0x7
AAgODCme/CBAPnVhyBvDCdH0dENebtqTue4cE0ovDPmQTpllaFWlM7aPdIG51WFaCZY/D7KkxagL
d6aYJA+w+FP4UOCCFbX/j+diGq1OpIprPzGlx6/AIXUimFK1l8xUa+hn9BSF0ELfDqEpLkZ6VEfP
b7y7aNQaVJMizA+RIh7kQwoubw+cg1gjE1cXZ1WSt0lqIrp1B3hwxq7Klr31/5XiJm5DycHNjXr4
/p2k4JjvkNVYMqE++Vxs4+YlZZ/AYJNTxTkDaDOOjjq15WSaPB/vSB8T8Iy21VK7AKYkM3pR17Rj
qzaLaQSbwkFfN8rOcaIhLj3Tr7wT55TFuBGMTuAP+nsNiEhhnm4j6wQLaZ9LLQ8HA/ycmslwSIaK
BFRUMEpvNWqoyzYKiYzofB66cuqxPCL63xEISs3HDotdJaVoqOdeQiXfdDkQTUMAr/h0QaX8Zwx4
Zd4XQQ8IPuOr2ZepIPyBCYzgtuDIW/q+9zQVRrVXrLfsVQ54tfGJYYwmRRtCgD7KKo6muiMn2Xvp
9seep0AUVgBvkEgeDLlyPqTE+tzS/Tb3XMzwO1ZOxp0T6ufxVnOEjfhCylYFREnYGMM5geepg0FS
NdvBT49u2xBYTJw6mFC03dgG2bYwKCeKM9H4Jn8EYR36lPxRYk+RlAG3Pt+uNNGkPEvxBoFgk9wz
2/rr6Sg+WkK1tgleGuAHtBBZ5ejbMgm+WEaDyYtl5G9iy58xe72/fRVf5BcbsG1opQan7lXeLLbi
7o/L1/kSou+IUsvgpWj00C7w+YnHJc2Bw01vvqK2oDAZyprhKUbJs/BY2J/0y2ssmm+YBF5uQrhg
Suh2qS/Z/zI9bBzm5uJnZBGsrVL8IVPoC0Cmd8zpB4+YdW+FM8oOc3du8r2VzaIYg9mxMjYonrJ8
7tSNsdotSHsGRMqqiKNi5R9fTTd3mPFu6GCfet4IudcVSNRMoCLpqWNrxLYrwWorzd7sXrVmEeQZ
UFc0KO4sFNUVlBEyW62fRWLO7hJI1+HN/NuY1bWo7iVJQFTWtMVO4NIfhl1NxSOdmQU6n7nP/ByU
wW9jrQeUXV8r3VMV3F0V64OyR3uBayjRzQTnDRcGMgu2PiYPeY/EM4zL9tQDEN41KsWKHtXqTx2L
ldgW+eTsUGe/x8PPmY7MmCD70d/rNuV3qnxtKd4r4buDPFtgAvPFB14EoLUbvj2J/fUZv/AdLBpX
F8L62cKkxCKXjapr+7g3e8bj70yUnrhVzEatKl8H4E9huR6sbbBk1TxkT+wzlIvYto15dYo8scl2
tm1T9+GHHgpVmhSVP7LQ01GiPV/hY+zXmRm9W7gZASPGQr/+y9yFRF2HXpC6M7OdXcSD0DEcbbWz
1DPwyhOez+mSVvW/jCBJt7wInA4KL7dMoeLOGdQgOROX210ukY3SPcHrx5wfmMJd41pG1Rt34qd5
ZrdRjBUiHml/P+lNfl94A+oiPAh5RqIkuUbufj/zBt82401MB5wm4YuE/ge4Jo8wHNGhztsrdosx
8zcKq6BA+zk3L2+90V6bPaK/RG2gjZFTBo7LOFomqUBqa4wxyi54ltnCDWbv/+mY73f5S227bMNM
doVvJH+c1Dg3CyCn47JYFvXYuSLAzTJu3q+UjsrxxtaAL5D4vtoM8ih+BJBGKxeXJq7GQLr3slRc
3SBjXs1xBeCzernAKuXOvI+eNR6Bs2uS8RiXBTycxBzos6uRqDcNVlhP2gBLng98ooELMXpgSuvh
FD+e5I//Esd1wfpipAEW96p5YYY2dkPgI0E7Hh5ssWEFx1j/fVdy3QAcWXtTBZpRv8YHe2G2p6av
VVylE4bJxjW2FfP2zP13ww6KMVG3W5I37SIOxGCZvbHkQHgQ/l1kJ3ydax5SyeArSeplnJ9vxw1r
KCrbwWgOOm94AGWgAfb06wUyTeOpugfQWr9jvig3j7QPElpjFutM9oGZp2I0nm8LZkmXTYgJn6tT
oLjfnE/kCbW0yKp+JhpACin3L0ntEL7WtHeOcokrkE73UrvOtuUrUnSv9cPlyeNsLh4wrHgAX5oy
GGKjOLi86HI5Z9uuXRXOpY5mNiIUd5R/IoNNutdpOCYa95EKR33synt+tCWF+bQhYkX9XK7EjnuL
ahgLL3bC90boSHLlNUvmWriGnJ611oaNbNwrOuQlwKterIcAN4nZ943RypLleygFEEDLOA2tCLFz
slNLL+hy4dECoCoTbOkF8TNiU5tRWQPvbwV4LXGzwtygoGVMa3w+Re6M2oT8r7XrXu5vdstQVP5J
6AxqL29MolTNBH0TKEwVDU0VKYHvno1QLHq+pvAoFJbFMQVYOhaLr7V2tWezOL2pFRnZMSGAeSep
3WP1JZR3GjHRJlhHGPbAhtVxYoKDXHvpdSy1j9T+52VqlihDxOGsQjDCZYvpqm0XM8siZrwJfQA5
khSmDqQ8Ys7ZFPOCPnKgr+QvPy9t/ohn/Qih9ul0Udb6OQSea/YhsEvgTHdTH6MIedBxEpPdM2IK
yxnxZ1iEPs0Rzg6pibtK3PFsINNzBwq3PW9wUBMEMP+8BVRwncrEIw1ONL5LDANCnLYDCGLPzjJj
bh6CbmGUDzejyt+ENTLdvSjcwMljsL/xQCDpoqNFaCxYKT5lJZK6kPnNYLGjpL37hycTFYRiPrOZ
0HEm2BLw8f/rS90q3nqtbCKB2G8IRplm02rvBBAcqa/CwNI1JlJ4vybEl8Jv5nmotTG+ISpYKo7R
Q5v0bdjoTDiVEo/VS1ePIXNsWY23XkAk7+dMsQfpdDRhWBATT2g0awhDTY+/bM6x2pSwIOgpKurE
B2fOtksBjWLwDpKyI/MVM/iYGWVusqrH2/VEmDy3ezv4Kdb+tJlEUDiRYXyGvbAjHCAk5NP3r4bw
yoYfC1BdIohCFgPYEsDguVX8A0p5/4nk4b2rJzXZwT7qYxhpG/O01flHqPV+mWh9gg3y63pKiXSB
Fxkp5vltW+Z+6AZTcqDGOsswdFt3XOX5Ohh3LGnP8NvOPqXp4xNP30H5Jt7Gy50i0pu0g7+h06As
Ehd0yax7VDNIcGt5Jop6n8dBjyzKtqJB/tT9YNG9KlDzx6svz4gXsiWhiiSLNk4kZwe1IDYPb9wh
WAgg02XcV+kVzpFKN/v8scM/k00vuug8lM98UpTEH+AqUcL/6XCeWF9uAsu3vlX1UZHE4Ht5iEEV
dZIQ1sjIsv51C2hP/nEPjruMZSM49NjtsRjOqZ5SP74V2JqcAEhUX4sKxw28DO4KI3Q8a8zxeELJ
ymsvtx5NMlG/lGBFaQM1hIETLwIX9kq+Z3WuB+NdKbtI9kD817xiY8YDeecBG5Ag25RvaEoFNGrV
7zp6QuPA3nh2T5df0FAK8O5ee6Sue72VlGRfYFEBENoX9ZCRB5LerrDwyGKdvA7kJk6lDGCxleTM
6eo84tURZi30A4dmE9ycqB4E9yF781HXkibGp6SFRafBPyDjZ4iH8xVc64ctWCU3/1dIjoMwrY5g
UdsMHjSU5/1HXQlyCqQbOXrNgSQWY6MDD03G8xrbzm0bv9DJgQ6/WiHPcbJu0XqM01WaacXXZSt0
HeF4y6QbIOxXpdfrkctxRnXEUlcRy1M7o8N1kYyoWT1QidY5hJi9ZD1bmQ3d3oKzJRysNg6a1s3i
VPF3L6AZFFrN9mzCmb6RarpaFllFIEY4+rNEr7yRhpImbT81bD8A5XHtAOyklG7L5oxwPLK+C5Eo
anOi5QZQ1s3nrlL8+oDA80ULFVtR/ujwvgSWewyOzvtJMMRSt036DnUFGel59DDHNsx6x/ZZD2G1
Sx4yREsvwhnJkTs/68TYA/USCHVIQaS1sHdgfEwYUNmko9yO8ELhJaiDiBUxN+L3ZcdcpVjxvUZL
z5+xAhuHLw6puRSXZZ5LZW+Ew5QJE1YVdZl3nHWJJzSQxszMgJCIkacgIBeWKL4y/sWM9TKYVrLK
RkACUHFuOZEHnXeXIyNJxt7O2pq5gQ4uL3q9X2e7O6DggZCvpeHFi8HzpfGYRtK7A8F11aUyBlaQ
imFaMHgDUN6NZXaiRgtsCec5TIRevftf144uN/r5E6X7XNLGCSgRSU/siq8/2nJSIj7vauTS8zft
AzXjTvQ1hSia/C+xHqa9fL9ZgivTiDf1AZ60utVmSrul7atFnWAdl6seetyjMaqxCzbkmStsSGKp
ibTjnbQ88qHb2Z6pGWbrCN37Si61NmuAtJVBeaQWRDmrX/zayuYQGt0Vt6lLHpEJ513JG2myKAsC
+ZLz28evBQJvl4CFH6WQX+y/Vy+HQ33d3V2DQhkNLWloOFKcxdgYRDnK+3hMjkh4S+pok6I10mWD
je66p8yv3wcEOvZjEAkoW4kkpXV42QHbC7cxXcjNsr1KqSFctv7be43v+SJdjhr6Ad9c48h3bBTs
PF86nezK7xbwsYEGN/Z14p5NArIMKkEXBM09QwhCGa1hySeAxrg33NkPeOWs0hmst3QTx5RhMvss
3NH4fJ+TvzHHkeALqFxe99LbLNQUc0idcHKEvNMH9ovr578vjJnwzEwKGoBPgcx65eouWdEvoFOM
nMUowG3DsEXwOeaNTXbxm6EOK5NWPbtGtIQY9LpUHWh7oyOuyxQsItvs221T11hVZgbLV3Uv+3DE
hUzOpY0HQ9/JxhRIhPA9PHhWsh1F/OyKbxQBpyoQoeJLRDdD7cmXEcOhW65ChJACr44m5HI+Uu8+
fUm6TpRYQPzOOEcE7EKoTwEvI+qw264fD3rFLcoCjpSFD6JX7CK9SpK81u+zR83cSumujNnfONRV
HQhFZWaYhAk+/G7TD1loBDUg8NRPAqo8NUExZuNxVFJOiBQFfBYo10cwARG92GIC9gnrMgOvV73r
toT0xnMSAmKris7hKXdT6fjwiJ9XTPcvwwTH/16HXeCllHI6S3DXmRWYo/HMQnijR1tIQcmYqQ7Q
ZkKSMrox7mbnNCA9GYWBXp7RNv51xBW68VWSZ7j4UpmtlV3a4zY8WuS8+v4DF1BmtXMYFZAJkf9V
9N/bB6UtioMp9rjrX4nR2FunFqPe6RpNM0Ccgti5d3OY2uqmM9ZCwgpOSPprH9u/b4W4MS592tkN
D64A40XYfcx5YhBKJAY0Jd9rZgZm5Ddt20v7ZlduPuEAgW1gpRdKHlS/KH1a9gKxVzp0We+xPp4P
nvupcIzYJ/Jpb1np4WCBgEh3hZLB6DY5LCVWWB9bjXVOoK8Z/oKWBscbHsi3rdvMaCmNH2htMi0F
ceM3ldpQwG0wGDTflZyTYVv64pbxt39R+/sC1EEj+smsDF7WOv8zPbAoILudGYthsYPJK1mO2Ypz
MPm6qAdqs6IiuQReVawRQ1ebsMGUkI4JW+u6mpgah1rP1/XSe6hsk6nJt4Xvc8d+jZX9GvDq6hZT
OQTX3mP9s1UjuVhpCrH/Hnm619aJBlkSHiFMIeR5TZkURqTDaLq5PoeV9eywjnAaxPpEyGN71mqX
+dkWztJESt2cRxXAfy6KvAFYiracovjtl0MxKk7HdCYZ3VaEpjWf3wYjz+oH+dx7i+QNtlT3j/OB
uHfzGS1h+dRYIngfW8RRfMzxDTcGGqFfsonxkinLsFlYBakGeN2k2UldyH70jngjvPLOfzgLpKns
XQHS6dQxPKmLPcJEfI0eMhI5HYX+v3eBbevbsaV/gEOcxIci0qx9UgeNYcHaEO+pBpePrvDHTO1d
IX2OWi08o7lJzrHECx+vnXO7XrWpI7cUjYqxG3yw9rHOvJJ+1gQWVGMMunoUXKQxoECUJQuuabsR
eAwv2FEwYOSqXh9djNmWed8NomE6oGZ2m6XhZtaJ9CqiwRwpk973EcJLyu9Ms9O0avO4/K458jCW
oa7AjrnmMobCJ9pPqDtTO7FUeduviroDsHz8HxdGhHnO/7bmi7xxwNQv00/XTVdLMjdZG3AgZdXa
YZfeR4hCTlw5OmsPb25wR2bWB6zxCVoWUE89JaqUeU0+2HCCPxBN84eGuzUq+DP6AxALJI6dfT/J
Dd0Epx/nvojjAjHmhJmvha9nB1+XrsolQEet4fS34I4Vdx8RzwrQ7f883h28hoLxKh6OtPnnHBiL
gMgyMmim5G6YEX2rfYKvl8f2ANpTryaLKufYELlRTCWvKEGilg6RBLIIMIQzp3XA5D0j0aPJCUQK
zl2e7RFWjWTruAtrgkvJxsF6Pn50sNggqiTb5zzMLeNATY1sHq82vCpafNXuaChi/uB1Gy93OIoI
LTFRuuhzAo66XIbsGZ++L24g3BScngej3NedDEFYqupmBSajAbSTFZQU8neX/Jjsa/5ASb90LQQs
U5MO6sfhH9FufvvaYk7COXJapjgfMcE67qMcgv9SsKw9juP2Zg2CJJUsfmnWlkzpOad6lsW8fqu6
jvWltLcjM5xqkJrM05YcTZ0mmwGoS7iO2Ff22EeX6Rg8DN4Mj+gp4iuwAghVnaYBOg1XkcJArx1k
tGnEfUPnj8J8K5DDcCV5lyEwim+UK2Rzy524UD+hEz+aDJcpegdgWJWdY0DRNt+xHsW+hhVF1uDD
LtH7gx0h84anv0nu6R5yJGk65XvGyIocVnXAe1Maz3iR9KyGFZ63IU8Gmf3ylu3yfEyf4gdybTcG
yDXzQcWwWKrODL3bfTR4po98cUWcNkxqGjRl2o/9ifH37QHnEp3clMZqyrayLaCUYv5FLrPRqLdN
t6r/eg1Azg4U7dBfvuz0ZDO3Kz+HM54TumzMJifQG0EtWMSqssilLKvFPENWoEK36KKPUqPK76u+
oOorIjtg+szW57u83fb6/qUbQ1CHy/2lq+4L4CQadW/WyMuj5vxI8hlD89z/Nf9cgknx9EMmrXkS
H7IUNHqujXV1TWBnCVTBQcDRvBSYpVrqDGnrsOeo5GmszFgTdY69n9Pb6ibwZDiLDX50WOLM6DGO
WGB7Y95gvOAWD5iBwoMR8/FQC7hbwUDExWU6E+437931VjqIfXwbOAzVOU/XqklHhTgtN/TrtH3W
nNJrMI69Fr0AlEhVr9i1p/dABULb7rh4fA7q7UTSUTwzaJKACws4yvuxIXW+TTSFqplaARAvTF4F
9O68W0Dg0SnVZD75loE03P3AJ9oRNLgVhJbODVrQxvJmaZB4m42XXs0pkzKGWLsfxQXhBRgTJ9CB
Ex1UXr1lgPU5v9InzDoy12+uQRs1bAFpfiVHjoz/Mh4gz7SQcPHgEsvjJDABByZBXEgxq2tGNPEV
aTbcHeSmL4L5jXLvYTqBX9Jbx3WUWINbs6J2RpuO94D5CKKgKtjtJ2cdwcWCYmta6A9HYyVyFC2s
Ib3yV8O/XQjjYUUgHN8KvsnJiah6mclW/5mcTPiSv49LzGC69Hlndu+bvCF/WqqcAv/JtujIi++C
4hdLryHnA2G7uR5K8Sx3TpfocchIcIhqlCnI+NqJvmZZSv4eqe5/HIUWCojzlUdQN+a2PaeeloF/
ol3McxAfMqxTyxxkyMgg172Cp8f1CyhS101Jf0GmTKX05ZAxpO6c68Jfs93Gf0oyex0vPpry1hna
YIaMZZNZf899Sr0NJyMUua8q3HB91linXo742uETshOFd9Bam/Ey/fXl3vFalIWXxBW2Tgo1bezL
NOtu/8MVOa1ggINIFIRdGKUFRFNgvOdLlIgrFtW2cobEtJK0iTFINuG2YdyQRSRhFcwv8qXhB/I4
TIe0h/9MPCEBJwQEq5Kt2HlRTNuuV6aKNdmqn1xGwq+Za+fLTnB6njaT/JROxBBW/EA9Pb7IhAPf
xuxV4Y5Etk7DBl0NliVIORy/MOAb/4vmpbdqtdXoKTPLj2loKNf6HPpYMsrVId5NRT341WrBL1qf
UHLnFBtPpgBPUzzG1uIxqrRMfKZU4UXy1GPhGxQ8u6+whevh8PG8oLmkB9gd6xoeB5NFf8Ngk07Q
gCYFBp+ovVMoszzrnzDyMNAYtWPKGW8WYzC1xAjCZaSJs2qbrQWwc8mfSkq1qsBoBbNfXUihL+Vo
c05s0K9HWyv/GtGzKTVVZ41TU8JEFpyNqOSdFsnnL6OdD/L6RZkYlcmq5GcHzDxxq7jZFjxYRcaX
p8wdoGsq9f4FO2zj6ZTN64sAEVhHvLCg6ZnNNb6LJ0zp5B6imfS9Qr8XIOI7zTmi/EhxSc4yKLMr
Uer8tP3gRhAbXKG5bIIO1yo/fZAwcTiyI5DdOokQlsmcvIlrHIfp0r7Y15JF6AsG3b49icwDHJWf
wkwiJ0S1cB0J3QDFfsH6tVtRbb6xUigBoXwDeAKspBN438Q/09/i3rCt/gPC3XczOG6mI6ri0DAD
rVP0WUbgQCenJ1H9ATa+o1YZ6AwsD93pcq7SKmYBkvWOuQX3AiBzEEIvnXDfOuiWfFQpHAGh43cP
dYwhQQXQYdq05KxwXRqPv42vvkRgyZvixRXkX/4r1/dGUt7Wzc30n8kEN2AIsEQtt3SI5ForlvFS
kKfwwHYtHDTBhZVZKyrxUVgaG5tlTEDiKdAb0VEyUzxWsEf6aoLtH6j5sMmts5ffNn0Vftqohjso
mYDTiDJySBoe2vsJp1mCuUYgBlhH0BXEbAKq4cyXeUZOo5nWyxjT7VBOS3LkrFsdnew72eYGqLIk
aPix/PiNB16A425PzkZCeTWna0qOKij0sZz7CP2diatNCddUdroC9NmHALtnuqs2OxvLZtGfxcDh
8PYJZOOEKlcYClRNNXB9v5KxYll/qCpndgbyW+HCOduE+CNYA7nZrxCVD1yjFtJjmmOCxcxb+J7f
PeJtQ6cs8HOvwdzA6aiRGcfaPi5dv2BKAwnsS7AzN/zhQMNTKDZkhQq8MCqwiZ5oCpyiFw8STJVR
2B95hHeD0dyF4ym8r1ueqXQi19q9GKgTTDGZMtVROxm7CM6UJFHKE4eAG5Qssjtve2QTuwbb9GuU
sEo7L6glQSnRSrPqjCZ0P9qik1ygSwKvwUg5Es3mlC+tuc86dQIoolbUni+1cX2a6x++YfpEb15v
U4aHUiLy4pjWGcyI/gmInom8+rX6cqZEQfTRapgyCWMY9iH+uLjwftIR6A6bUfCRwHYmravH29hU
Ns8ZtCuC3zqi1o7vEh6gm2RW4liEm2X+n/yHN8BSTgsnN1QxFgxeIBa83DZUfrO3FqEX8n2imMq3
CyiH3J80qvxbfl1k/jv0Oe+RGvZ20g362MmjvszzWJshiYHpQNovTzwvzwW8io+vvGf9/ml0md4O
lWYkQdhkQnp1Yl12DF8394QSTeu/Ja1SAiDgiJdlQLLPOZCr0t3o5zv7ws3TngVI2/yPJLWUK5WQ
Hk3yCx+NouwXiLdMqnkUNTcf3YsNy/gscw/QsMmBTZoluGR+CVbr3icBcz6SMi+wbg3Oyxd++7uQ
JzJfwwrwMnHVVl1OM+V+f8uBqK0snOHll00mz7mI9ZpZdOWL+9OYHvga1Iph0UoqHRsdTvBT4M8Y
VhDCgsgdf3hVJbHn5uGaja8pNbusJ07YqXRaaV0b7lpE/Mf/6srBahTmXy7uOn7XRKFkOBPvLL8T
d3lekoI8xZajN71ErMGDFcLBy5+rZf3jQQDs2vkFY13QzLyS/84TSs88qUXRL2/6B+79aH/PLSP3
Bh/7rs0cp8TetI6a4GsNYHP79dJuilwbEvLH/7ds17mGn65wuTnkVcD1UmXm4zSwBPof1w1sDdFO
9WJKbKz9xMyO2xd6yGZAXMA7rWXXlWoGfb0b+Hn7rqiPtpmhRgWN5SYJJQTayZeoLFn7KrHR3Kye
6/lFyP1dAQswecp6njXVZ/89BD6WxQv9DWzSEyJ3gd21qjTdA38giMhsqZ/NoPMK6k1y+g0IeWnJ
ImmuvqpuNQ4p2T6/kZ163Uv4tfdWIXs2ZrBDO+HP5YI1u2xXIHeinapm7nfXF2RzaGCpWhgxPKal
VzcBspextw3ZrVc66+J9O+UsA2YT42p/nhhpoi1IHNXOc6PX+5sV7pIjvjiyQYbAdesPLtInsJED
SErmKce1kF64VDGTd2EYy05BJA2cZT4VSfll2Lox1EJZkWZzvd9nRO0/ncTACGHkYrV17EGMxwq2
3XaAmZRiRnPJYfUpezTofwn0uNW6RRNN1bZfdtxxqQkWMc0brMWvXazZoU2MsXtxl+p5AEC8MA01
L+nZDaOWyQ4SYMxu+btflfjwXsL8E8wIxmg5XGNa63EMizqSWkJgX5CE8Po4rOIlTADzSUPQWcki
C1dBUfiFocuQ9y9oXegBUvnrcirSN/Dq491LGTv277pn619Xv0gfa2P9rGySXmN74LTOlRwH2iJe
lCaHg7ChGOBjFHwe0KxDInjh7SM3l2KGPCYQw93biHKaXf13PjAMK6OOxMbKw1DFvMxnhOlyopVU
CPP0cOn/buDQA4BnNAlGdtGpnyf6ssYJBxtKZaWxBOiXnQlZz30AEQWDLrIg0DNVlNUvqHnWHqk2
UN+ElHmLXSi9EX8/84EHDuWkBUMV6UoD/v2aRhvbH2ltQAowyAFFWZOKaivHY0kk6ZERL2pXuVY9
VT4zlKjOqzHOinriOOZwddVo7tUvW+mTygJW/Ccr4FsqXaLXz4OXjdS7lbIaMjf8xDYPm4T64mE0
QO1Sm1LAHRiZR8mrefD45ENzQ7j45hC+nE09RJAdNBJyAhM5v2Je6AJZb+cR37i2UItFkM2dwmrX
WeCpTuteTtC8X2AWa4kkRJI9iLEv3TyuDFBnR4+PWuseXWqOQzGXAHd0EHYPGZ9+uId6W5RiyKF0
p/sjnRXvgC2oBWjY+xKioL+bqT9ERvrjYoDReGuBqoFIXGeWBKn3ezwngNuP1srHDUueIbamWKcF
dIAsvlzQssipHWk+IJinl5fN8ibVwJ5UEMUMpafvJuAU3gj68cycRJR7XpZidYbWWGP4b3w+uPhI
8/k6bpPUNe4kXYr4mssTebQELgzmt34FxKpv7VF50XVuj5QAmS/kMV8gBSRWrCwF/9wQxH2eV6e2
aH7kzM2zlM8tmgBtg5gGmDKE9Jd5AZAtgTjpdCRpSiPTu4iPUKp9OT8I7VGMFCNnfX13tAQ2YNgc
AByRY0DGmMn+34NvwCFXG2PxG5nW1KC7mJLJCpX/7B+af7de8sGWVWWd5idJDpJSQhyw2T9pKSOW
yIqZksb16Um92HXvXOfuIiWT59N9E9JKvlP97d61zfuPmMAwktSSNu1nRaiJHbraFq65M3Xbp1Tt
r5eL22bbJu1/wA4yt5ny3gbBq8wDWEXSRXKmuRer7nYf277lYIqmzFxCIj4f/V5BuqrN5vhq82dZ
eeFq5e+CIgk4bVuSM+ri/YwOw9I/rbrBq3pl1utqbwCu3zdzijLIX7iLqVSmORwP4d7xGjjIDWGR
yJPKJ41SC8oy+yGK2Lf6yqxtnApUz4x1TV/vqZsVV6yyB0d/ukri/y5klTqRBVRgvIMG3yCxDjdP
rE13RF0R6GpMS5E1W64IBqxlsGX7h3nyPs9HOMtci4PXb6S4dF/JI8lz+xlvjMD6Begs+x58xcAo
8kx4sJn3jxduyIYXiNtKldLFrpRDWFbXVVBrfkP0EVpSrBoCvTdTPVS2Jcq3Y+3XHhYJ2qydLLDe
8zhHDnxK5hgnAEA+EmwUIpcUo14fMaffUnMLZhZkXpnwex4yWqxOSTPTxAgWYVdEHtpUa9f02z/N
MhLas4hG6edTuxgI/U1n8LblXSQPSmUfUvwN3u8JEFrh88UNTBMxSgu/eWN33kG76YBPs6yG3BNT
JPHuMOwJhmuQujPzo5FRejxHsFbkwOjNo3CLyjZ4gnEg/T4VejGCEsrbtGxPJItu05DUBUTS98UW
v75S/QjKb92DHUvqf3xXWFxaHyl4vj3Ifv3j6GYOA+T5GpUrP6iX8R+SFIf1PZ6pd+I/HguMSkEe
PKj03TBqtBjen1kOEzstJOiO3lerUmS5qJUpayPvlsd0RZujV2fuGf6YDlteWCGisnyURkIetKyA
0idbgGJDkobnd3gtTqrxPdN29Iqm5cviXuwflmsYE37K3z8UxJGVx7t83EY+gLWZUJkxVc/ybzfN
RYi/3jgiEGvT3D2++zQAKQBu8KoGwviytZE7U0qDpma+Hsc8zhVwCMMfo4XBxfH+CGe5IitvPRjr
pLP9fqEIDX4xITqhJODDx/WfalF0SPn9ZAbKdHJQvgoGjMaMYQUz3hDIyo+I0BNJcxGW46UYiTkW
k3B7LZS2R8Lp/l82KXmtg4D4wiilKI3fTF5qTsKnXiU+IF25228AYqswQ+B4nyZx+BqFBGK1L4f8
mfi5PaxH9zRb90Gu07CFSYDXNfxqwIIB1jRI7q2XliH+Uny6QzjeA9iHZHDInbfSCf/iFHMbH2fF
bRvvudCoMy3DHHaimgjJzNo8mHifIVg2TyMxSV8eM8Ewg5lIFXHb7JctbV5XiHReLSxLh/4MNuFC
kr3Hq8FfNa+ZqYJmwnYda8n7f9quDNBC0Rde1RD2v5bm5wUrvY2GI2zXEdkLiFo1yNNDp8mSI7ID
jfhiRCd/Uh5YENzq0OMkQBQoMKeOXtW5Tbt3KglqK64ENi28r6apGoI9vcmCsYgwBM0srZBNxq8W
SAOQT38PWVMy3fxJfh//9JcITcrdQp6gekLxFF1Zo6TvXvqGZDtIH/WiiW06jcv8SQVDM2yz4YeU
aJ00twU38Zz5Dbb3ubksUPsz467Ilm9TaTqfHBZC24QHZTeOMjvB3dziTpJjI6zq8vExpd4u9Ju7
pU0FoRBSbjt8EU8KWlx7X/YEhBBz9rHGFU46lBVFaeWrURSJUxmRlvGpsZRqvSzRxznsvQ24mhk/
ycfEEkpmAioxu924AUaOIDWM/1rQzcsbj/Hz/qXuazUS0FXwRgom8mbb9Fpn+8hkXVp089GdBZwF
EslC52WQrfDaX12+ramE2nPpw04maLLJLSwZQnqkCxvUnKSS60jCUJ61eSThmVQPQWTSFWxC2DC6
YhHeD2qifvJn06E16eU9VukR3FTp0JVA4k7M1aPa8X+GQZcWhmrhrQfUcjjDwFM+2owgba/+Bd9c
YDtso/uSptTydh4L8EqrwX62JY/MA+iR1GdCThwsKPEjCpf4bzFvaMNZknLzTllYPvG5Wzi/qpOW
aPTUq0S7mGx+6BuUP2VaXrxbHOybxl1nKdUkcAL8hB87Ts0VH1iUogsSbAG/Vc6iT9Ir4wXT6HPj
a8pcWCGBY3aSroIlh09EqlEbtvIHSvGCTjo2EMcMrCSRvcooASO+bOpnw45PdQZs/ucYwKmCUk01
OjJUinOeq55wsRdoaPFSZEjgwnTP/zfAkLkzK2KkUJJi+riHvhTDQmEkXUuIcDIqs/crHsOw0lrU
ekL5EXEaq2/2ZZ919j/CCPaFc7eGAvOY2I023YsD/qhWa2IuWO6WvDVg3AnxdYVbbguUllzsply5
W/DKGfSs1/AQLfo00qzctyalQxKUULhQNflvbMVw3wp4tzKMgl78ym9KiGpa19iftXSNFuHi6JYy
LKFe2tzcwMH7rz9ZA2vIKifA9sPcl7+uJ2U04fA89xqXsA1SwePIgTasbC6TnbBRCcPsrZa4l84y
KZiFzRc7E1qHl6M8EkCQr/5pO6Lyx1DabMaQQ4V67JHOCePirme7An4FQss8Pn2QdQ7viAz2yX0J
eVIohnICKbIstDQ+TVqOwHKo3HAVhOkXwQoO3//iD+WYBjPZzKlkn7Hlz5WoclgmJ1/h7Cr+UPbT
T391BWyUmbS1FosTK1ubdk5VupgOvLKOdVjsfcquZJFXFvMFVByYgpJxjBlLzq02xf/a9C6dJHiw
2EQpJyAKgQrrR9eYXHWGJaBMfvKBiZetTz/Q11VfppefCHpEhRlqqWiebMpzrOtT7eDpisDh1++/
fZO3bMxhc7no2YJR/B+uRb52YlQCSm8N8OfNMWTQATmp3P/6MJJlroGFa65RySD4rUv2HTTnjWfG
5uOwuuxgzeqCY4zdtr86zjB2dYJTf4LCo+wgSvuWRt6+3ko4QcEaRBdelXLbvhXTnfJnITss54D3
hPEZY4UjWffnMydBCOkjz8SsmZE+OJbHYgzunTPEwMv+QJ2bSngEwxcRXwQwnuExuNRkhSjLhrR+
D0terDLnPhnYUaGKBbto6Z2m2d9b7QytOYdOwjzqtriWJpypSzoi8DbT1pnM2Eqt5JFsnPx9sozK
H3ERy90SxmtUMzzLs5AWbaCh/IAIzqV/Z4zl0aC0kz5VlyeeSQpZQC63vwrtlTGq/cd5YcElSBCr
ktzl55olmCqSe027jpTOInGG+qKsCJq3XELk4OHlsYZEe+hELgc8377jLSwWtnI5lrFaWzfIriNL
tz3cYE06VZ3kBy58jqyocU05W+Zjjx/hLpt20yGeU8p0cIQJJ59O/KjWyehOjQNOELOkcrERTfqj
tM6VLUVOBa+qZgmJOXc3XS6b51WrcUezY8XvJdg4wFeX/1Q2/WbSQHstW3dAExiha+kVLveHFA60
A9Gy9GxroTCALhVKqVZt9tiySApk0+sdQJw1Kg075k3p0SgUjX0aYkSZZtgzKSteUD3dL3u65oxm
YbGYnjNpDUeuPqCShEpBdCS80DugMhI6d4te4k16ISlyfu1KVlwKDqgAFmmvnTkUJYeIW1MREFE9
9us3FrDEgG37x72rN4nXB7OPqlvLQIY8bZmUz4OwkOKVCSIWH3fYqiJwO6QcqOawynoTsn4bt9SC
U2y9bDQ616uxdXPbRWbgIoISIsK/MZSi/FJCHqkUZsNX5AFZ7ktAJBGfhiWbmjd6VmddnoLPxsnq
yk5G5NVR6sdBkEhMFwggb4PoB8U0j2pzrzbcrKlb5RQqLjX9Fuo/c8rTYRl4b3DjKuioi0gqj6SH
SNHp82XvVkpoF+RRB5fceA3vm02rAN3Lhil6fLIvtqis6lFKQbcio5DsJDslyenHcsGU3VjGuXNN
eLAYWpoYpYk1/2U3D8bpXfhnPt7OymHX2wl3ODCmoMNZqTphcu3FQUtM+sIv7kvo+fclfQCj/6pF
Dm4n9NRPx3ImQf+uMlu+JuAwStJzGmJ1sTJ6lI1KvQ5tZfqzv68FTiX5H+ZBTpdBHvYW89hLImWP
SqqpjHOdCdL9EH8NyReWzWWHX7o/LSV7hLJRzcs+cOSnxdNKbOZDzcI/oO7rbvV/M30fzu2EEgeF
RjXDNwk3wgofYq2xfJvRMHXOVf9dYcmuLJpzS7L7v2Tsy5ej7Yv+XC9PRIYSAkZZ9DhfEbjAmvQ0
FxHcUlp0i12Xj8L+OQ44v10lA2ZP51zuMpgBZDsO4qfyNm65S1jfMTHKqLB8BP/61HpFZq6cgWCe
BMMjKq+ADxugj7cPhxWf6FI0wiloUSn0twxnL/Gz/9PeyGeVVHOJZPLpEOMJOLLO5+s8jtft6wbl
CrmBS+6FqDLVJbC6k2oxVYcWU3Fn9vbVuy6wDShH+iSmKPH+rrdZ5Xe0PANgMC97V51vg7vopS+b
fa43GT1TDG0OOb6vSKQN7SdyCKcfxUCVXsnxWhFsYghoYA4yLgE7shYqHRUEuHNwyJ6emLF8v4PA
rV9TaWf5l5p7FkirCFkcpEvGRjj9w0GTflS6mvH0osJWEPZiWLo0JUBr9R+9pGulH831O7ViDJE3
KV9zXUWjYXRvOBF6mrpuECeydEwm95j+Fj8IOMYh3J+OebpkwKF+3gP31El8BAGfGqtMT3l4Rcff
l+4D9IHNHzMkakrxQQc7FiHT1oTXlHjhMxZC8I2uY10TUhSY5Hund2gP9mfmalfPTS1TdW6F8w3Z
fuwVJcFi6xrfaMTWhxZ97o7yYHw4fpTTl5q/w8/nX4JeSzDThvrDOPQP8jrhdvGoKhTlOlJmwqgm
0IyO20LbUC5DHsKuyvZC6wUD9qzXHsbO7rlIzFXZS0MOU8W9GnA/L1leLGyKCoYBngCu7gimeSWy
tEiI0tU5zap4cMdV4rrK8n+lem/T6ue9W00w2DPRVBLDZHQ5Ac3OBUoZ8ASQfET/laCGObjNq/Kh
t+rId7r8fl8YXLU+nyrswYBEze21SQJacqxJV/OVKc/noGYnDh807IrQCodURNlAXrT/zid03zQn
yyKrhrgf9rnaDdHfoLbOiK0FTWgLk72Aec0Yd9AXSWFBDN4RQPH/moBPQ3E8HV+Kke4eGZwOv7C7
VSk4Ktgch23o2tAmZ81YOrqEmswtiISup/73g3rNKZ3nLayL2RSSFE6bTC/+TBSRlsXyF2LVnh8v
ANdnnWKzMHnnc67LNU+9/OEgOQjiX+So0M4ZpkxKeL/hwuGPcUB7Z0R6TdNqkX/6y9vQkCfMyScO
UxTAoFV84INScYHS1x5MmxnCd4gwQB7E7xpItKJIQfJ+gedOLV5cb81llESwtHxr2u4B8PNsTnud
JM9mQa6nrhcpHO+zcvLsIptGwPLf2o3ErIRG/vzF0QK5Vu9Ro0VLbNPathrU/Do17qc+Af3l76QX
IXuQI04mdYh5lpWALg3tTL7U6+GGNfe5N8Jtl++BKnOx6Qo63yq+ldB7c2IICNApJl89G2WDPzqZ
Id26d53G1adhTo9XCtgGD7jf8ACSfy1hlXTkPS9njovE1orhfxMHBob/GHRNtFSqnuCK66UdL9X4
YBaYitq9PhPhzDX1rg3tmc03oSKuQFaKJydUTnmhKsrWKJDCyag9XNS/QnvmH1eDvoP/Au+xmqJq
CDEKVAhUKIsy6ruL/oHUktdVGnF3y3xGrWwHfQgd+kB5TIkrA/FuCUUChrm18Jr16/1wPGMRJbEv
EOgPv3Iq5vNXyzBk4Naic/MFXzeS7VTnS4GMgENQlae8bcA2QmAOO0lByrkVrTECLRBVAVissMgX
TrZ9oMx8xmGPk6rRnh5lqLMVKfxFv8NbGsUWIPAD0stP5BBOoyfhGDEzIY6h+SztIlLX4jstgTH+
OEQ959wRsJCws0VncsCNY6JGfAUTz2OicYGNLm7xSSU7zhZCVhj41fehXsPPf2a/2lhHkcYKyQXH
oC/W7pnwgAQyyMVsw9xCwrb6TvSxllpEnkxkbHIMzwV/+ViiB2iCp9ybV8h94GJbhdtp8oN9JcT8
0hVXs2huGafaXYArVwJEzlkqmzH8KjwEEx0F/4aqtLKfCR3geyJMwy7WuiB6QTTWObDKOzuKQBaK
uYRHdT52wIelitD/iwbKlv/JXnEnWWwcee3VbdUBl8ESt7drLuz8HvttMzQwzX334OKNi8H9HtFw
aX+06GY7Zq4LflP5oFBzoGudfOtIcNPQ8RH5zY0njBa7Bx/mLFJv5CAIJxXMRMRTzl3mPR3EFKAq
Et/FaQ7Hut3eUHBFrZyW8spFIOkqrqRIxFAvRAsCb8GC9mXK2lZHIPK4M31nmi5dynp5kxS6Gs5t
px0u7cOI3qOPEIFvgWBYJQeyZjSR1/mEnRxjEY+QKDQ343SXGGlGPW6n8SjzYgxbTcZj0xaO/bvu
eZOJY2uSPVczGAo0LD6OPEYajsw+qElr8bPqHmqq7H32VrWSOfw7Y1C7pXGfLNZdVuRdPGZiUyaQ
RF7dDFAWZmEuifbRmfhK9oR6LVS9885iDPIyNPVyKjJoek/n0JbmKP2Ar/8XJu+sROhp0J+F/zj3
ixIByqGtuOeGGMXVviJ2URlczQZvNmwkJW+9V4dD5PrgduVv0RMQlINAnjCxkRBkNFBWM6zhmiwS
6o9XnZKLKa01Una87HQX/VYRwVYxPPYuqL03PDQpE83e7EfbuXFrkU31g2E1IQvNe4sp8BFpUkTA
9MVRZ7qF3kgCbiwAp0pcLL/XQdvT9e2z6DMO4SuH4QOdhUDMiAxpLV2Nds7TUWkOo2/E4agJ9zRp
6Br7ZRiuSBZRcOvy+9FFk9e9dH6Y3cMj6PecezeX5j0H7gnA/0YIpOnukaRs/d/lxmUT98sjv/5/
X0GHq4nMde1tQxAffOfTdsHh605oNODhUBaGdBYVJ3n76iZemI4hRw6LRJfz7wJvg7QJX44/uU3D
mcpN52kyepE2laAPPXnjq5gmf4XMyysDQzF/GI4Cp8V0RZPnZ3GKUivnKCWBObQBZgSrmQS+k3tZ
XrXQJDsu+cyjElEzJakGyfFYFDwwcyfunrNA7hdk/zY7hZQ0ofIvLNuQT0CZRFecS/1/0J/CI5UI
V//CEUuBNqaE6vmm4q5/TPGGjOJjCV3d0zmWceTpwH83i+6KChNCd8cm0R2NThN5YVmoCCLqQSEC
N3cj5wOVMrWyAFg/3aKWsQcD1wVIrUg6VxJmXmZ3Y5ZghaLYFb2tKH0pwWmGbxhP7ceL+bG2jLEK
atnu+run+L415sCDHyHey3CWaw/XKzTPhvQIZWJVZRsxJhphy66NL3afA/udSN6sitD8/FuAA9Io
QFtABVyj2XigNG+KczBwRbHOCn+xyc/HSTD4OW+S2W8LZ/0HADUv5j6UPn3tdeogmH2+fHOBNbR/
w5xdi4Youcocpc7R8NTIB/jSCSbrq836vDWcSjKktsof4TMPKXRftMGmESNi6mu+UzV6CTYJAR3A
YywfxIIKQ5DOpHudrAPExdSICTos81j/kX0YYewJHITWPxaaGtcEeJ2st6Bx4azjxw+x06X9vJvt
NNfspeKiayQ+GiPkiSXSNZCFoTFtpiXoDHKNs1+RjU7GAuOMkk1KHGZuj40QDpDnJkleDVmFPHgo
sgOTFo3H1ien9mrZzvyxAXOAl8JZrUpWzmgrQXDXpnbR4twvzRDSu8EB3BZ+RRgMNcQt0EAkNnvJ
fTetvtEpebpLovzA3cljoRe+dwxCNd+eKrJhY6U/+LfJdtC6rfzDXPiVsmqQYDDLOcruJ28WhfCh
Zu4BUDytGSmAfRVc7p3QbBKYHSCaYoAWb3EuzUi2ChgH/ELZl54axyxjkeinUdgJL9Ddsj8tb3da
Xsh1/KuigaOzsvzhR9a2MybA5Bo01MrSd5PpwFOmLAr6Y80VqR1xSJScSKjMnKmfrJBd2Pd3jwE2
zyqKgUTp3aXC2dF8fzPHTX5lMrWHBpkNtLLcLV1sX8ZhNqIVm04BvTfQczKSFByyJktH6NDNetPZ
Vz1y86/W9NF9YuxUybLorHqtXDtnqNVwunDxqbL9LV9GjAtb/1o/hBC75wCxF/+mIZVycB20JKdm
PGCiXf65DW/IlPG7mrN8sfz1hyPNAJS84CpCj/+WHkaT8sCJaDf5gfNrOOuao6707J0bGNTHBn2j
sccJnGMqSo6zo7/+ljSHuX0WLWVHJnU1njXz/ZvE6DSWSKyf+zDkOep2RXGQ9cdXhYEmXvvTAKK9
oNd5zYVDmSkxTks0LEqDXxYTIFOKPxiP3bKT0hYxyVArz320NTRCEg298TLKCsPIvbmjj/4WnuYS
cDu0ITPqh3IYXJ6lJOEbbA6WStvK/9QI2phEOFrbi6CHSFnT6V9GvvIF+/OwB5CKlxdnn/ld9Vkg
n2cOZdKoFwofXynJaN9bvVGxSVkOcIbtaPkooUdwlTrIQMydf1RPDU+6i/t4zwM+CJhqGnyY6MSy
P/HH4WLdnN0LWiLMmKTLUmPds+1HFXSwz5StAwibsW4RowqPEHIzzKyKS+AvncZDaKc0GXYaa/z9
cF+eOqT9ulaya6gQPEJEnLDgmzVIaZLVmzcdFKvE4JjFJuETLz97Au4mdeBeO9dSYGVoxArSlLNE
bfIawsM4+DU0D49YEKlUIY9CVa89eEHMf69cs4WbXaV/VQhv5D9sfCjaGGb9FyX95nFa7HMGZwlI
/aZTPSDN50Giv1C9wHjSmfx1eNwWkYNXJrtUnCuvWoCtDRSAYjcsOJePdgXK7jrUTU1HYXgNizL5
OpSi3PAGDLYZCEa6X4H8B3eVHDblTb6nWnDN+uAHNKFA+pynldL1k1tNxy4CZ8SXA9zHvL2a9ltY
2PQnVDHW58Wj58SSSnBmbN43KW0u36P8zyN8rQkJ/BHzGJx7jBq4yIA6UT261w6WHoBlXQZt5p0J
0X9AVi5cqXQuHp2qwUD3VxT6R40MunJphxNS1Mlom+dtSaU4SdACjb1b5DILCqGXjx+RlvdA0VbW
Iwy2rwwte/QVgKRm2QkHce4wNuL7E6nIQr3m6CNYuSPEKIQuVDfyiDA1eYumSpUojJ3TmF+yDcZX
1s/vlduvWlE3dA5KoJZlW60sIoU7bZrZCxKiVvY/jmertKvq9yDcZl24bebGhP9hDkolq0a9sYvu
D7Tfds0SAJGbQ6UpSFW6lQ+ACqkScSV0OJd9CmIDjZLuE1/R7g8oVS64ZslnAUaBtlpNK9I3f/EC
VKIk2VE9mZ6PROUgK2927e32WtNVreboQftcBfPxu2msj33eEyapXrFfXA65dmiwpoMRouydFN1t
xw011fYAdVrKskXUmm7I+O+r8bqUvQgkg9cVnPkIrZiPZ3paILIMXT8pRD1Ah7xh4/EXX4nzgPiZ
pC4vBXuBwnNBRzEDsW3L6k8dyxD//mMeLhS2UAxto8bEq7bS/FNKBPOl0hb0Q3aIy1cro7ErlwFL
liE1+/IDu+6LBWpOJaJrWl68IaIa6vh7PWtzodlOZmRzsS6OkFhdPAyU/1JNQYhzZwf4nEeCAOWc
r0pqCUNEa8j0Hr7+lYRbkBAttGSP1cyFKWs+k1bY0uvySFOzqBIBhlcrCmMlad35lOAOl4ETxU5+
BDcvrVowfc4A24aufETEvOxeg2R/AmUCXiHSOQK3XOqtCrdDWhJr4Oju3Hw7MjuY2uVGg1e7ufhu
x8yFqDbmcFmoeqLHjbfHDnvaLZtIJKniUVik45qlfgbGQOhK09zL5C3CdVk9uDkJStU4FPGyvWiV
PWfgrfF+LthdkkD2BxuXhGylh7UNYDVK4ccKiQ0MAWZNqN+FI87oPdTlW9EAuGtOhA3zGbO5PapT
FRRn2JyyVCP5+/idNAWN0EdeImCwPBx+4dTas9dBbmYcUFoRvyw5Hqx42BrJ4nU7fnUMYS/LFU4t
DmpzCWRIdRdZYI3+YqmpUuuoHs+21uCheuQu+d9vkY+EcYmNNm+kTHcuqc24xXAbCQ0mVbdbYUei
H0SPjTTq5n8ck/n4HnD2MXYFUeXzSN9xSMhTFvFhRgQF5zlksphDwsEzx7vAbNt+WZ74T3OpPPKQ
0oZHIhBx0XCkSyFx3h4ezQyIdXh1ehmKjFDZt8zQqtb7Vbuq1No5NPIYa7ZyS9WIqJRTez8VoUpT
tdBaL/WGbLVE7xZgVNKTfW0aUKbcuX880f5L/LQfQ6yHKQ5hK+j+NUMZAkHj8MNU7O2zmUpQcPz7
x11wQLhkNTBKo3awCCrhyL2E3XybFD4ddWbYDpZMhMhXXP2JEnKMzgNV7MH5VWnu/yVYiPCDJCJT
eaoFwB77np0eNDc0gkUaWDQHD5RzJQiGvdyw+7ZqZptM6/ITMgocdkGIzS8HRjZui9xhRHxjyDOc
oHKLmsHjRcHzra/ovfB3QT64XBGT3RRC503iI0RkdSNpTWf9m9PBahlcTS9BRx6xXEpAPufM838E
Kqr8HGPusOJxUKz/GNNf1uu+1uVHDiQhfK6UE3SHL8BUdUgWzasxFMOYxDah2NlJ2x9z4fD1YwDZ
bqHxVemLZIhjr5Mjv0abOu8DZHbXtpldXMSSxAr7+Bk+5iqN+CLAOZUbGqFzXgUuA7iDY/5Mx1Pf
e9rzN2xArs822a1KXChuw9HnAYDUM13SN8OFlA82aW93jPRdc95HTL/y4AJuXnXq84VGTSWovamC
RaCkAiYU5D6r6n6O1enpBeYKsTz245mnS5ZXWhWdhUMdXCClO/4OXKFaZMNLkNwpkHKgmC0EcwvH
fiDIx78f5z4tmppqPM+3nTRbZ2oD/6dUteJOvztOhVKW5P4hKAOMyAwimoKDeVjzcz4WygL1fyZ5
923kbx7NpCRVl+2aE0IaBCCT9BUYWWzVOZT4qvTgA4tATt8qBGmnX2dI9TqHV9FfTUYfxu+znYWt
VAxM0B3cLfMIadYecmpMNXzufXf84hdwShM4Th61h12nr/EePKGDuZE8JRIFgO/tElyTvhFrlvS5
ekqno3U0qW9/4ySIAkEUtF7DS5uoLvS2cEkygQgivmjpK3M9OigYPxv1UpvPA93FKj3riI8Vwv3F
/dWF+iXy2suhsqUD480MnSeFeRp876LE1yw6MQ2MUH3V2URdxZ3+wKeJHr/70EDbFpXDgV4LoU4g
VKKQAivRV8rK6HApGcZaJ1GTVpfXA4pEsMogsrqrRFF69Q4Hz74fmt5VHXbfct1VQhYr0iPEUllI
FsWXsi1gJ3pDIpUnI7xPr/rZebo/cVS7AX0ZotTO1fsg5OTVsK1A/IOZxSS8tfyjhPXqIPsHu6Zd
c3ShKQu5kK+MZHiaUkyUBHgjLWEgjCKrW4m+qSLAzGHfTh+SnlKyvVf3Rp9GNuNAj0PHxnmqnrYJ
nq5VePPSX3aRweZqTJe35+SpxV6QGuoTukGTClsYI28cc+imzgYHvH01HxDzjXFnlCctYPFe1iux
UV3Lx2tVTM9ZqdXFFIf5MQZNFGNEmjs5sOicbALQljh0UoZAf2ZQxYXZFoM0KJ3k33yhuIhyp6ey
ky8RBwTK91bP0U+SEOGsmQCHGi1DxzLvgQ4x8bZt4I2u9uqfQ0rQQH/ftLiFhYCSsZsz8Pq8Ppg3
PVIDYQFROlImyZj5S3zJe8fpX73i28IAhRH3NjNSYVb78l/zjm9R4gFteL3X4gMdMU2tNT2+d52q
13Lph3toMn+FRgM6EKR1Yr6Hv8v4pj4YJ4czls1qcIWond3u5UxL9Zuo/TUSWQLATJOxxsQorAiY
ixPA1fCHidBFU/a5HvOavAIb1TFtn+6z59JYhpAyLR3lJGfCO2fpz68PiNMo5FseBSesFRuVpZSI
umfszPX9ERdsGOWF6dFAgo2q8D4dLicr8DVFlXGeZjkDqF6nJguAGvHSVvTbIceD65dWqzs56XEj
RmApzVtqB1JPa8Po921vq2ZhzbqvohCRJZ3XfMnox32eZpSM7NALz9WwraE1VEhczLiKc7J0iTwP
x2B1VIeZzP7K5tZh4ex7t+7yCUtX4RnGbCy4swMojr9qOmGgGCHsxynCgpNi7pbMXPrnDCFleRRv
im0dDS+P8VUrSInzNRNWSEVZOfqB3kboMjHa7D8xJAAbvjad7Uz7AU/4CCL+w2vmL4t6LynjnfdL
B7sL9s4y4N78rLyxDlFa8AvM06ciMeDv3XVTrxvlnKsGDbCGWUQ00u+72JVL05m/bNKqcLOWU7mi
E702q+QEifszRW+pCKy1wf7zV/JmcqEKSflzegq4jQFQN25GuG5wdDF10D/pvH/pPSqFGvo2b5Fa
2cNyqi8SQvEO5VhH6mDWIX7NGtBkpXWNrnJdcNYRJSBw2CyFd9y9JYozp5cFHreEWJEeA47UHonf
rp9HR8YUCSnVT3B2Yl484RpTJGHHDlNMDHYyxxIhDA+LggSuEgxftlirTCV6VNC8QVK/DTV/kbk0
nJYroDl5g0R0M7lZ0eVMn2b5B7kZgDtrjqidMERziYoeRlLFd30HYRPrNq7Xmffu/V5yGIN98YwJ
5XFEUYyrpgCpZuc88bMPBbnk7Ks149MefiqWqmPtx3oJY1FZlaHXk6RAExYPUU3vWnD9jxkahs1T
OUfNrlIBEWFUeGGcRFLBiqHKAERFzeG74V4IpKyQgLxKOeeCqlBkdGRMRxKy5IhnUEyis/mQqLWu
xrCpLng60zq8CYn0XkjBwA/AL7R14IuzGa4zdSFSgxQNvQR6KwEfE6FD52tNsMJY5dGAJrHE9aln
e3EDa/VuaoGSng7769DhKEHOb1FFjW8YmZsELlCX13QAlAhShirTk+4vrxO/SYHwEWdc/XJRMD64
gicrK6aczLT+aTuDjtKSA9Ti5ff8U4IM+DG+EAIKqdBSV/KVqV0JrCBReGU7YWAizAHszhCID2Om
znS/BaOQlZTSYZF/lHFwZ+T3zP81y+Hin0eNUEg9kzrFOQu/FJyiwlPyVwHEIkQacbEYmxcsSTGR
537A4If7JiMmzaikgwXBIxMJo//pD3I2A77skzdo7503YSCz3UYk4/EUNAsnNVvyWQuFSig3A7Hs
l0kcCPpSU6iftVD0afckDO64buR66bMu7agfR4lYeWPIGI4+E24ITKbKkNUC2gQx6jKdyBH9eCFu
0zH3SNRFfj3HHG+TTFIfk25iHSDA+PzLwf3V7QAVncQomS5FFgPhVu1zx7+zUmJQVOXkgKr7CWko
PPwC72TmzBAUiSVV9XuqMoUVsxlmk40SKqw2PFgXVBH5sUUXxQ7GCagUyRBZbtKcMScuQh0RhptM
D1QhH037SmAUXoi6+OG7kWJ7FZKI8BphTY1Z+SlVxK1ITkAA33jgSQQQTX3SF+S2NkXvl9kwa7vp
yF4QS16ppfAsA4H0+KEZNaYdwp67aevhcEapEQTAHfsBtea3MWzeA99Bzg/FSzA4J3/pblAgOPF0
QtnmEdABIqnVE6r/yDoSs2se5hgmGN24EPuo5sqLsNHXlb7mtslyWpDfIVtGyJo6lQeclx/q5Kj1
vs0QCLbjsy5Nw/AUQM5zqALR2usUncahRN35z5NsNYl+tTeC/skr6oPyMeZmj9RkjpN9I6sDz0eb
fYEdjMx7EZe9Yj+Ozvs0nyaY53e41Vhppghj9bGI42q/7NYMqafLld69OjCVNKduGPtK+ooAJuhG
CZ2ut9jLRNDcFLVOaoeTEbOctK8t78SuwZ1nK0O6pBhWsHy/SmbxS5GK6HJiPehZgCDga8Er7i6w
EZOjpQ3AFVkSM25bUWTaTs9DSLXrMA+sk5u6/4vVALAtVrVO40kw2PesmeaDRs3qsOWpQ8Qlu6y8
gRxPyhKV2+DlOWQGaDpGZnRrJlbeEyvfE8ES3H6CaHkeh4FuZV/ejwsCG+8uKQGRKEjLg0IIff5V
ZDN33wrqG02mw24vxOdgcE7HrheGLEMKI0eif/NuPmkVvYlPWcw8tbUXMUCX4jtLcnRM8DzoLNdY
Dg0S7VTQp0l0vJBi1VhpfC/aF4dHYcMP0uThavGCXoFGNolZfdlmvFS48yRt+MwXAPBYEDHENxpx
4UvYUuyviC8XIbKdLf5j6LiajwaCWoN6KyHHvokI8dj/R6aTKuDGHitMmByI9WUmqmPMu6yio80U
Sek54RCwZq4JVAdeys+KCE/+StjgwM/fugL+6Zwepjc0f2GWMFCcrezqJJLmjKtEHre6XZ9dpMjX
1riTqEHf5Cw6/yw+3p56m+N1+daopkakjYv8L0jl6X+oyAKSnRzobeba73ZR0aQgy21y4qhbFx12
iqZrn/2DtXsyDclptqp+8WIky9hbEh/r4JR2iS2Bsp0osmX91xFd+Tpb1zWapoekdITpHPy6vCfg
KE0xctj1tykTBgZ0dqeifgms+M8ui49g5o4xNA6iFtpS9HuQ/6fFlLvr9E1hJWcXcTRBfa41rf2w
PEnEqTmuoZXOkoPX6yQDORmAxei7j7ii4E/usPnOwoJSxKu9zFthZE18Vz/lJjC+Z0UdtdmfdVyv
P2E5HUODxJSZqVkSJ9vRWureR+h+uPrFEV2d7IvYYCR2oiJZBmbq0o6hgURh0uQc0n4VVgc7eOtm
WmdZxeiLpc7ilqu9zPsoktcDxbhnXsuSG8F4u29nq7zRQW3HRkMGacgj1szvK5ztZCkzATQy8edt
txycPpxUuNTRSjt6OVdDLxXl5TRYUaU7oK3ub2FxSYbEtheyHHF6yvXYwIx5gkA3e9Du9A44FHWt
cdjPkcM1QgA/Np9jNhwTdr6/LtdLLFqFXZAunFr/9SacCgsgAHt0w2sAabGuhUMSEak3L5Quc6Iu
/OuHWaTCy7Q4k1p7xhkWcbl6fsh8e+zJdFtqkOsL17arr6rlWV0mc7J50vxLN4UBaINtzyLNuEf/
g22NDrl3TFQp5a57FYDwuglE+6t4K6zBiu1HY59xtms9xe6CyGnOgLAjRI716YtxVET7ywLTKTFd
N8Y4PlDq76Vv8DrtVMYU/qjOLtIpmRkT+0e3ZzX4neSITupJhrbGwLvt3Vg9KmuJk95K4Plg/68G
bjfacIMimBZ9PZsVDaeNb9DFehmCaYnxV83lT1uzsKBggdmv0epc+3yDOr8hVyETREwjMLWIHIPD
g43hS255U0ng3g0YEmk6zzGD8Lja5Qw8xrRbkDmJzoigQABv3S6Ynu5dp426Px6fpEPrW9NFZbNN
BHHR13f/oesyipecSdHdh5dY7Uo4YWZQimuKZKBXOgyvnJxRSSp8n+bC5rWciz6HxhwkJiAEPntM
CwZF3nwcN3pTvOy53hUnwTeIPcnJBfBUvAroQsYAagKJw2o2qeHmGq1qbGbMNYtdeAoD8i4FcjiT
EFEJ0dy/lirT7bjzL3DD9TEdX9x4ah6GNc742+NkUGTGFkI1KhpZph01L4fndkKysYWU8mGdYzKc
capvF+a0/Zg0NPqhQ76MUZs/at3meo7+gwdcQkyNWT/LY4PuyyNQTSD68d5WddM4FikV+nvc/KL6
77OqIFKEOdYUkk5O9sa0m8z99+5oknrC+degk+JHNjKMg2liT4Btwy6ryyrlrmcgIpVeiDgFUqVG
oqGt/abuU5pIrsiZfITUkqBqsZicnv1RTDxERV4yKofFqUIhbQo7okvvH/bo1XZhtJjAzJu42hU7
IrK1SvZNF6dbfIsmb3mG+dyUv/geKO/uSiTLHbuscMNaDIJmohvU+fjasG0wev6Xm9i+FwLNkR/Z
Gr7fsAK8vegGvz/jsHdFBwICYYbnmZVPHVw8vMXBNUe5riKn4bRy05qw6uhv2DJPCXROgcyISsIi
LdoSzezzTXuAxduwLJ9mlt05zhHck3M4YgF7fC/GxVKV16YlheKDPJwTcdrbUlWxurOOycGeka52
vkWeCOZVnxDf/EEGLsnf/mKHtAdVpIlOCkd5SaiJbJH/UcfOM66MhGex1nnybv9Kyi9uXP4c+Tjd
OwqxqrQ0taX1IJ8FEVLjmzkNi4QWSrTkOaHzdm5tO8BPSoDxVlhazTQOFdz7uoPkxWXH/m0JZkIT
YNvLimglgGLZKBYYBqieT9SlNE8Dw2fpDvUD8Ire2/TwX25XwJ5g7W5oeiQb/O3a8ZU1V8jyTpmT
PO+PHKoXHb1qapzB4ez6mbI1vOWHDKpFsPh0EXPoogYF7MrIbgUN0aw5m9t4w5qM9mOMwljDr849
Z1n5ILfJsWaLyCBbUDv19CLlvm7W82suKg+WLPaOi8wNnt63r9Sjszg0ukJcJw+h8SS8ibcFV2ub
QI8SQJWKK5tjSIKjmJlkuQwXzpPGaHVJ8Oxuzcim4NazN0msMGUj891GofjewGCjHU2mSa2N/XFg
QoHMd18Sh4bcx/847Ks3lK7v5KHbLS+aiTwE5DcBpYxNtnD/QYRnwLtE6aKZS1AAjrEvFcvvYEL6
MtCjeY6RV9CcoA4tEvzUAemULo5f8hZdYuY1AaSrnGSFBQtmc3UNjNialdl+OaLb4mXbHLBqNo0d
Np5WbJGFzePf/xiVmn8zIGx2h4zVQyxKE3fsFxDAvHn20Cq8/C0DS0E9qt6GwoXSSwpv6nfQZDbk
ng7EpIDDspApD6o8zNCQMTaUKJF51YCyBR/WHd4psoiezvgdP3/1uarywRCb+CvgRhYPhPdyv/x6
Esi68Ua5fGkWrNDzQcDo0kHoEcOXAK8Ncb4H1ueElP0K7R/SpqcPoHiHLJNoLG1MI8csopv2OQX2
PsRlGDI0UCRPOVs5ocpckN63snXUfHKSu03+Z/0sFUUXMJOc8/R6+S4yUAygUThv3YLyYB55zY/k
TPl1CL71rLRPuqczqSBoIdlLV/kHMAX9AWqGQgtBBLQ3R8N0S7m+IXXX6omFl0llBzwHAMlTGl+9
vinBzckxLvpaUDnj46NhLfQNNrnLLmTSammKO/7H7uD0UTID++XK4h2qgju/JJxKxIoOJ2FR923b
nNGPb9VYtZ8TreAWMqxnKDKrWIsumtNVM3ExVVKohRD4p3QqAex4i/KLMHpMIPKZsv3BtSmclIOb
gMQ72L12+/lu4Ce9zU0lx4jUvvWBo51O/1lqaUbic4BmOPx03z/liNoTjo0MsJKCCP0p17zDs+d7
1bPUpODYN1ShP3XGHAIUVWbsasC7R1SSBKesyUpwRSv8X0qFWUGgURyzWL5GVsbLp5gNTVPD43It
Oas0eMTk8vSVlOtJRQyev6bUgBv/hZo72HBgTQl1Hmwm7FjKv3ynJpOXLLg0i640xkzcZ/GJq1bS
RbtwNOV0Vj5PdH2FAhLS1oM7Q689iesGy7FpcfG7R+LLTbohkGAxliITosjPcRVrJUicnwXqudBy
Ni8+lOc6oSQZSdcZrS0z9/sKaZyg9tRUkmpxTn4FG4pCmNCfq9OgvYSSsbcA8GH9KeMmyGmuQTpM
WauzIzpLg8CBnj2jtRHF7UG7m06XEZJT9Xa55bwmPP3USLHpmUVN8gw9HcosbR5zI7mKUGpxQdSI
4h4uDLSN+m0dKF4qJVJbQCgCXbeBqbFnvcWDEQGt29VyORn6HngB3NacEoB8uAphXgG5N3I0n4v4
pQduBU4r/NhBirn6EsJGYBS7aCgHKNDMmbOiLO0kbh+YVsOUIF9dYatjFOQmtgMGyr3jhvaobIh/
FEa/kY4dXvVrMiPXPygA20k1HUvqZxosDWXBfNxsDHpzrabns8ilnuwwmmpZrL7rCeO+QwtmKN5w
5e0ypguLAJ5ncvPQEIkz8/ioZVRYUTzc/l699hcT1sQYjczFvatN/+1d0Sm9zLtf0C1o1Adh9y2w
uSra9OscC7YW54x753XQIjIP+fCedCQDW+o2WOb6sPsB2u7muUBxgVluqsFAyZeBG5phxLJYBZMi
6tDSkUAdeqDmrVybKhd/M97MA1hPrGohgavv3dgSzYFav5woKo4jyNfQusseNFvQqWRv8i8O4Fwa
6DUzj92HOFgmAokVd/NR5mLlgZhX7BJfEqmuepP0uzgu1ipvjDbylnm010u2k6Pz/pfTi5ERdXPX
jCDF72m20JBq//EUk2JOIYQrrJ0bU+goffyKnDyE+qsEQ8MMWCR0cCx2XCMptri3QlkST5+A+IYP
SNhmi5CCAqfvSyVlQHyw4Zi+8SZOUSlwQMwNutnpzH2OaAKeb4KFIR04j1zcZ2kZj8IbXfM8VDfH
tp4ibL5OkR76fChdK1AkTGBc0YihB8TrriSALRisQ4a0hT+H3Vy9pVDuHgdHpfLSwg2VuZpdehWm
flBFeXgXDklOmBd9zoLxNSmGTb5/MqUp3RNFOoT8r66QigcBxe4BdfA4Wu26wejlkb5lOVRgEtfu
eOYiUVAnoRNFVbI3yaJSwmLGWdiUmh50uxJXkqENMtEwnil/G0Ec1sTJGWhEgKGxyUdxA9vplZ+I
nJNFIP/zlcHFXdts3oZAaBkTX+RnneKtCvL9py0nvLV/tAdwFs8m3i6w8xJ8e6/BSSDBrq47cdAs
wW3DBYUwdvHAQQOj5Ql2Of83Z+32Rz+ceHn78LkaCfYRg/PJAc1OqZYsI9AWnujMMKZwF5fM7sLo
Xc2kjE6xmZ0x5X/qeakvGdDdCT9Z9f62f7H5mD1ge8L6L75IlPoqUELBhqYmVG9BsCA6phCYyX+a
Se4dhXaajoMlEGBE24LkR4Jyw+q/Nxn581qOl/nSnD4DCmOPvPD19HF+4qScS5ajsa5LIC+S/y/E
2GClTz/JBlBgJ/U2zU1iM5pBODvkkLRyiRzuJMRG/HC06yvJBn+RM0XT+tW/8hanASATQUfWTyg7
HBvrF/3mVmtQrP+17qY1xZAai3mOc92m4tmKKRwhudlzHNGh4Qh3PzLe0r3h/PugbilCkHRVpI86
LVTuruJfNp9yOx9Kr86mrgNhR+ASzi+MOuYqYcT538YtSE8lLgx7ugxBF82XC5zfVbkzQ5we0wFC
hHyymzm9Zrr8qjNuNkoFmvUf+JPkhB/K3+yK2tARJy+rH743o4n4GckAP/Yjjp4SEC0iXxSg24nw
Mi86F80CqvNFsEQo02cfO/EkIDaVCC2fP3E4nvPh8o7etMuFAuwFlqesxa1yT3dgfdhPB8amxsIs
13y48bc95yyrKHwP+TzY2IBkFmUlMW+gCC5us7q3v2djgAjr+QBkhgyJNX4edOYW9zJHJ3NERS1G
hHBley41rwFG2lFCuX7rZ1bMoYX7YJvF8cnKe7ygvdPXtBzwd/MqeB5WJuV3U1BJEy3glAcgdiMs
JmTgV4Ze46swr65dTM94durmXxevPc7T2JliDK09YwGx8bf5dxEbvuq8VWmr5xU0GmanTKaJjTGk
PMT0wneLzqv0Yutocpe5kyO+5f0K3Kjwdqk+md7fp/h7plZd40vjnmb9q4gAz1CbOlRZ1dQ/RPz6
yuTx8oEErFh48LiDAOudyXlJhKJM2RwJ1/ouD3KuGjggFxYENyDltCexNKOyXJ9+rZoIlpaDUOt7
dka5zq2tL3EvQVLTRD1YT9lQnedgXhCnu4THuh2B1khIkJ7NRl939rDM8lVfceF26ZanJrRACvuf
3E1SzdPGLGiaXs/jTr0uFMh9fTgjAiaSIVy7qtGaLvvnYxvCUdEJOFXtWjNJvb3GB4g+IcOccDNw
GnGc6fvju3IHRz+ovNfxwRilyg/4Neof8IV+RhIekukRmi+dNU7CczZrxB2eNCWP5fs/EWgehErX
npeqkgSNzuLc8gX11cjElA+imMnvX2bz+P2DKV5QCZA44glU/JPKPnCh4k75eXa7DZnq4WxF5cea
avfblex1Z7VHo+mW+FRm1N1IFTtJtBn8j3bxApjL+UxiiuQnQe2NpKFECVcGOMjBuzIDxJq6LQu/
uIKgH7YdQ27skyn+O4B7pYmQxHjtyWbYk4LCVw410JokKRFyqtlNA81lp01P6XVJnSyKi9d5uf/T
cmKlwkR+XcAMJ2LPkvcg5DnDEtVAzjqHsrUTTIiVZm+cgkCDteW8VePbS/6wkcOzHY7iqdpw6Di/
z5+AxXWBlXKiXf6ANUNUozZONuBiz7+sJvSjrbx/mFnsj+L7nlwZjOEOP+KIWZatUu/71sc+HA0x
lSmaB/TV5Q/4vPV/YjvMHcIdFsyg+aZCedarxzws6Qt5Zt+wAw4q1Hxx8mdq91H0PL5bnGpf5lWG
7w7HOihCmErDCxhjOWRQBGSMb8iIqoRlvUKXFFPYZb1PT86s/j1ZhK/hfrBrIbHcTNPJKgBuuMzO
ehOAkyLzF4ZUopHFiB7clan8wvNG13tmFprw4Y97jBrj4gTtkHjgtFrRNduUW795OIuvy4QBn0g4
oae2syHV01R3aBlY2HOVHcet2YGsOXRxqc2hSpxuWrorPkv/J4cG1HjJjvqSoKpjlSqqTxXg2Doo
0CFIBaN7cFcRwbNXySAMs1zNMxk6P+gsA/2rIpc7hOJlRdSP/735THSlABjABzkzQBQ3WuboiTHK
F6+UO5P225vt8wTBBzD5pLhvCG42034eQXQQLG+E4vt63GVXNA0TT4CBk300gPh8jx47bHtDacyz
HymHF0EdprUpBYj19Qi8v6GJ164YeVa39AveoCQTYdEoyDDsA7YCje/UP1h8eaPvrnKQ74C6D9ZJ
zmIHi0pXKXa+igqlhaVg+luIRwK3/DFAL3yFGWh123jPIoV25muL/b12JuLp/24qN8CIDAdsFx7c
ql6J8BYBopJTmYB/fd2lNdDNcB3PvSjFAE1lb1x1jMKZDVR40VW1VVHcbbe40Wmr6SporaIHmNs3
o4cUit6kqMH4UTL18il3pnLlynftrzHlFmCvegeM3IZuSIEeto9mitj4eDzL6DxjFTkhjpnkYhwK
2NXJle6DkYdJesbK3doO+o5VdLG4fONz43/bljfEvqNa1NMF5ShYJXsIMAOjqN+ClLYh3yuTFtv1
/kDnqRjAxz6nKZZ8giMqcsRXnbgHj5fa9Jfe6rW1V+XpwAtom0yOjv+YrLPHavw0umSYU8mSv9sd
FSxAxmtadC1n72vTVwAzUjslG/Ve+PjpmjBOLgbmTz2PeQ1xBFjnAHyyRFYJvsYtv1PGx7rBy/ke
zxhxfhGGKDVtuw6a/DmYb1ESCvLbAoS6Qt7B7ysVk8PmCgvVmGm08riPHj5hFp8EWCLCLYEORUSQ
wNVlYQ3TRgJnt7BWEAdu2X+uecOnXo+WtGyItRrNYX3nfv2Bq6X0UEPxVS56JY02MOTlPiXDaZeS
KLw7ydK2UQzWhEYDJgs2rIxrMqhXRYRTapR/R6JKTouR9Pg7THuPQW7+nuQz47fmpmbIJmdXFh55
ELHd4xWxncOJCpdYjkV/X6n1jMPOU8OO0oqWEtizzot+i37YAlTkZicY/WMdyRvI3P3XnIfyzfZy
HC3Nv7g6KY2uigyEjSZE9ewaHf0+RaD0RvrdtHh5raE2+mqFWzDvCzE8V0A3hXG/3qEIsJB18+JU
Mvf3dtAzTEQQNQbgcZ35KWGjo2q6oM0TU5+moNAPtFmrIl5OKufbW71PkSNi2P5k+PJ4kJp/j8MA
fo/LKoWDmQwfPvTRNeFp+dxbr5GeyxmJHmqnXCk4882+GJVjkR7sh7AG1CW2Trp5Kl/j0J0XihJR
DLgvh2R+DBaoAu7PWehDhJKWHyzhbdD6YKdg2wxmhy9CcbteAdI4yf3BjQ+B4gVzqdSufZ4WOgX8
3svl2DyAyr6WrUDxUMC+PgaN2JcmGOWkSxsIoklzNaI3ahbsINt2VxzjqneqYwwzHiMxeq/la/Xo
Cf4Cjp8nYPOI1IlBEfY7yFRZ1KnVJ0FnkQeba42rkz+XUnWN3b8EEkAvmjzBoqpJCiduwwU7Ei26
wUYdOrsEx9OjkzmvKSSbSWKuXD6ldGixnn7hljohVizX13K0jYF5KGDgmTlTypIiiMCBuUC08w3w
2+2ntiB7xREAhzuigtLJMRNFVB2bJxxq1r3dsK0KMTwWeSLZiCN6XKTAC01DYKPLk9n+A7SzBXv3
wj460x4F91ASYdsdQ/fACO1VtByHk8o63nvYagZDitihFWBwTXbLks34RgA3yKym/E4IVATTgAdL
/HyzyNeIrJEJUi0BdtmCL1WiPdxW30bGM3xR3tMGurp7mgZ3JXMSPeNZjATMRnqYBiengyoPnTpr
R3a7ShZfPloCJotEFogKVuNRBMPZC5FIa9AsNO4AX8pUjv0yRLF4qcWHXCVF8sT4fObIDgaB/MOt
8BOLXPzqHcqRKY0t8OnYeIKG1ntUelvxtiGlWBT5POZj8pqgew3mdYeexDoMXBDAdzWrbSEAV24/
rgb2bQsI0DaDAwVxXfkOC2mvYX74BNfIvLr0uwzgYr4xFXEOYwioG+EV9Zr/KZaqW6KveUtTz9EJ
VdnpHLrcoLcYcXq9pmJhyp+nnb9i/QN/aaio7/57b5CHcCXVzFiiC+DIwFldDlsmTcMNMbXOj7NF
6Pak/1M2RS2f+6Tdz5HLNkXolcWMiAEukjstq8BF+8UhMK18K3ilQ/gsgM+K2GYkpZ4lPaSyqrpz
bLQ3LTKdLwZarOoj9KO2BYcC7OiqvFhLYjGffluWYRPyjA+tcpL4vxZERF11BZfBa7Zq030d9Z93
eWBY1GvXN0RQVIhGpPdPUXjjIHgmBSMycrau0EIRp+mbfQcbB6p5O32GlBOmBUrcWu9Or3hxpsx4
sWXneXtnE3VcsuLGcTUJ0Ay8wLxOi1NV+E92Qov9tK834MQKgarAcY9M3ZrnZerFl8LaKwliVOnx
1zz0K4t6PFx5Op9WRKV9z45xLrhpe7w++hk1PYD4KlcSftKTKaqaCgg50OQ7/WKNJv68uXd3yhuh
siScvPJCil4TWl2QD85TEsVgw5FjeWgFehxMpiWFsXZca4+x7hqH7UU0cot3M8II2VleHBVwlWn5
1CSqBEKxtcT5nRrfqJQwiKM2UFwOA/EWbIwVNpnUIkVIdm7VTFbXPDtWP8K6TA5A4Ea+fsDa5ztc
VZI8L+Upho75tlvHzZDnagFTxabXrClwal1V3YRYf3wKVOXqkEIkhWzyjrjYhJYxuSYrk++dw/oA
aWiS7BbEvlO6YEWQ8b4reMw2f8xg0Jl/l8W5IUeiJR+ZDgV9t8U4bdieIvTASclTMljyNEvGmPm9
AXQFuSjp/buGbItuyplyUwjqB5XjJj7PIBuU3LivOl10OE41N5NKF1Ghi4ivr4MFST1SXgLhm0tz
sn6/MdszqhoWsOdT2CnNdsALE52xWVFNe07CVAWpoNAW/MT0cDLOCTBbIEY/11rtIsXImdbodhkh
fPyg1oJKL3yt1m2zLel2BCsLTdZ/ttY/4dgvWbNcZMMsEqdEAMZni9EQF/RluFoOT3NDdFOEEFv4
ETZEJJD68Bzj9yJHhoSRvQLs5/RLLPjlsOmZk6+rXlcaV/eVYJHAzb/LLIO8SPlg0Sv+K6SH6+4S
q06sOQb+5JpSxOHkaH+ZvOObOxqjcMl5BGmTa6GKLynYEMFbozmCpcmx4v6VXhBsf5utMm9mBsdU
El0/yI38z5YDOxFg+RqNh3lkoLxvL2br2zv1AaPtE4lXige4gJ3hEZJwaqF7Vakbuvo+gEXK1KEI
7KYopmvx3pVyEFxXK0DgaTLlztkn2uEU8MAJmD7ph55MFpQNdL3ASXAksdCgiXxD9yq1l8C5hr75
UEnc64lAbjQ+XCxtObzb44ppwUYxPNgXQTBUvvgiqCdrdR1xIm2Wtw8yg+M27gJyEsFG8RMDEogB
AKMFCuqdxLNheYtxE7GLMkOeToPvqw+Y94gI8gZIF247lxWr+mrlZxJSD/YcGjfA/oC7eSvxzSjo
oW+X4mqsNkeRL2R0Zs+SmoZv6M0xqQ2Rx4G+IcgR2ZzX+IBgvrgMuz9WB1nsGkPvymxFudbDmely
XYWVUMBiQiuiFrECyus9UBwvzTTHKoEllfm8YXWA8u9UNcWKsgx42BQqycKjn+cuyPbX9MjN1Ll2
unZZ0EORhyznpL8AAU+3wFuu5YG1HW8kRNYIz8M9Vr/TtEdhSqPt1y61ndSp80A6lTM8tMxSS6g3
dl21mc4AcPwaG3PtxYEMLpMJcE40LTKpeJ9rAPc3vqJAKscyf+V6mjxpbaUh2zwT+pKJRVvK6sLI
9KIcZIPDG9wrZebkZ6GgAzf24XoIUHCH0LvczXNjwyORG8RPZruDmu0Jy164zR+xS4nbZdIQfoC1
DOCrYrIm3Dp9pCCn3NMPKBVdnf/rxrbEntbHU9RsMy4GMeJCdfgoStq48/oQsp2uzszWtMmdmH2h
SZZdYjiSDa7WQd98zKwGLLTdYoKFdX/GG2LZjfwLeZl7K9Kx5zk3XSAHKS3WG+IWwbnJ3jVrnUpj
jQOTlapjP7ThyqXOH44tSsKsxufKodLRmDNxmxTeHoqJLf12nmLQGtoBXgzF7RK77hZ6+bEgKQdb
qZgqERQiOecV9KVxe53SaejGPxwyvFW03hHEdU7BkxsGjgLdPePxRh6IFL/GDSS/RulfiIZiPT84
iP0V636N8Tx8PrFeCxmW+VgPnXZIeBevEYCUBnMUU+QmPd4i70AHsCql9/grYwRvZB/JTa8QyUKu
K0plNCc8+/UI8WdI9zjDu7gWRI1LpcNdau4FhpveBEhMU7MHKwrog7UWfkusr5Q8LyLEFJ83HaYd
WlqzCpVYwwmjEku0i1fcbcvT8FW3oTyUgEzjLx6dTEr/oCbtQOkaHfAc4buU00PQNuYm/DdTAk1/
5uNZUq9gFkA+ouK0MelDsmiP+5fF55d1+iIajfJ7EiuAZU7Du3h3A9Ay5W7GDK5JTfGJ4B8vk95m
kGYKr+bJtTJPzXEQZXBSQXh4jiehq6CjSGtPMoMedsKL6SC4Cp0ikBZQwx/G/xAXXA41tIiToMDq
fD4wNgYDKnHFYgjx+E0Cf/XlH9MOI95i9icxHp0rVXLkLqR5dnVrnHAeMkZTXWYCZoEFpCqVqk8d
GwyVHpOoKKsCUdnz2XTUIZvxRLMPlccfxSKvdxCu6wuxyI+UfNbeHk3xRXDMBvor36roI2BlQGbG
7g/8Vy48DYiaIwO+8tV8cX3c45AJ0BC6yEDbiTHTknTuN16y+ql4PXwhtCsWmbXDk9ZzVNM4QVCR
X4ZM1fMsVUdS3ha2Dub9iZ7CLdWAy8H8RLAR9mQh0m3XMr9LU8ToPsddFCaCEsFLt9C3R1IofsEb
R/pyFK0yU+M+EXo/UHS2Slyj7YXRNCFqhIA9+qeFCYfYZSjnbiyWwFEG0mSEuDX1cq9e6QQnInSz
BtSv+CRcrOArg8lUPE/HuHFvi7bD9KFMOuziYEA3eUzzmsrpzY1ym97Ixjj7vI5txCqnGErex4gg
RlX6Ab8qGge4kWxOoEKeHdrJkKO+raEDalY4xRZIJ6thEXAMMIyhisnbyeNj1qqdZKo3Y2AXJ5tZ
JOyJb2ZlomJSuGcL9+zhyTISDCG7wdulKJPqh8nRYrMhON1L2l6lsYBQWkF5eUOicGdfzwlbcJBM
Eu0SYag0XYlV+RooMLBszP8ROfa4FbSHKoDutXBevUmVqTJxdNki+P4MktNPyKc2yBYKgcSZzZkT
m/oM5ocgM3der/DUIJ4FJDFGe4vE/Fcz4Pqx+vMmzsuV3KFEcbyNG0SJvlPuWe3341pg51o19AH4
zPVrKY1W5K2ZvjYQFqUnX6reGP14g1yX1iafAkODuEBIqeDhiSgdcE+3L0aCI6GqQ11IydBc7tXA
7OcM6ugRarQSpA6alF6XOtd38+SA7Qj9lBrz6dKYc4LonBbBXJZGwU6QIoPcHMWYFOH8YDb7DyKC
oPr+3CyuVa/jx5JawdkR6XzT0LCQlr2kHSl/9wyzf2SgyzNG9YSQVJwjN68xlDSpY4uDQxKq2vCT
/ZbrMRaNa2QEXnVLVPm3vgzWGBZbkJrcDXMfkQZpigD7Z2elRnyqytE4FjzWCOLiQ56qHc/NYcky
peGWIcx8B62Q+jYYDVmwaE29VWvBSkx7PdV7D5TJ+ViSet1j0Fj2x5G9aRW3oQH+HtzC9F9DwLJk
0rnqOTUZpcKNzjcnOODwTI90pV7xo3RX8rDstSsGbBIsGulpT3EMipDUqn3HEwNrj6vh6JTvieYr
Oao+VIXYMPQXw4CdFkqhAgiUGdCcLgcOinZNG7sKeXwall7tPH7cevzyABaYWNOiSCpQGisWgvmd
nemquEhPlKJ+DDmUc4xp+lBWtQrjgd3YvwCGdvyVILqSSnShWQJtY+ACOM8sOM1xzVqhjnCcfdVj
ZT2OsIr1eQoOYfrAZyx6n0NRpIvjdz78GMpEnDzddHYk3WXl7jt8rXgoxQlLWebnJLPWeujx2pqh
VVNqewxioQ1Qc+G0nw4BC+flqMY3/D8lR9kKLwGPFXjHi7gqlLs7yZL43OSpMi36Br1tYfHhxhcw
a707kJsDiUBqgdaJlWTNT1kGsQVdk5CUlZF4Nzl6i4OImvt5w+vfMP54Iqgzc6QFyA667Wa7sWHa
oFeXCSv0EOGm5TXP2i05IfltfQvsT5t69G9eBbLLiatuQloCF0qONzcU2+iX8KzT5qzrZ+ap0sSA
FTUqmOvnmVCxOnGeULN0WECQmUQMNxkgfkUAjETM9/R4bpZSkavsbbO85hUfsxzcStcjn5egScnU
u/svKwh8pMiS5ORndUhvkfTQ893l7s4gFmvEEsdYou1v4czUPIA1bPbBK81giVFN+ZXQRxKzC5Zs
mFOaGY/Fw/xfPMA/aYoleDaVsnlveXYhLlI4zysTOpJGUVZBWk87eDkcEx0wfmhd0rT/BZ0iH1z/
W6CJJaKBptmkVQlIRR4qIl0LkmRE6uxe8adPfNlFIzqy0mxCDxaAg1gjQOSqUgGpCzXr2x7a2/Zw
2/jdjNgA7tZk5pXQr9jTwKX0ce/YIFGrWcdwq+pyNG0ty2+5aVnCln6w9kXCKknGotM7NO2rt8rj
wUrXc7LPDu9d2lB0z+vfKLbROTMeNiwgMTgHvlqZvMhs6vUan7wi99nqHyOEQj+g5LagHsz48LRm
f/lpkNxqL2i4nlbgDlXgCb4wKusmzZLWDtRCokhXnaqUMZRgfUk7p9n0bs/ICHnTeStm69lNKT/6
39t9JrFayRVb2eQRcUS0fxfiFXgvh19Ga7bHYB6KgW7uJr3EPokHPThQRG2HwIQTAxO/R5p4ocsW
kOlzERvAdSlKAeMwnA2ODgauNyX4OYWpY8vACGYxpAd/he4/YHs+5nKnknafzAe5Deskt61pvf3l
ej/tROz80tSRMyWaZh8swG3L04lqZf3AXdzlV41mbhVQx2UZQMjyRKEYMX3arzENS1Z078n0mPEB
Rv5e5ERdruzlIjY1y60XBDngy5wnjdnAp//006jXx6Qhh+s2RPYEgTie3GW8OVP2vabQ2ATKPtMx
sudqnsVbCMhHoQzqO6n/WpusWQPCqLanekoeI4e8ScqrP59nxLIcO/5j7x06RnExUQcl1d3w7Zqs
ERo/I7td72xI47xKJokiqrl7bl8NAblzBW6OBKP/HRbiBbWQRz2bKz26bY1odTbHLwmtl8muEpEW
swqZEnBnSTU8rcZ1uSUJPZTUAl7PrUA9buTN+L987ww3Znq4afPAwYPkc8qx9SRyMN7AEUBZZgQP
f6zVkxoI+Ca05k4mQmmbCgAUdnX83D4msPrXee6lKfdSZAMbZfCIYyMC8eZSAa0gd+nAaH13MMw1
tz9AmHfuAohC8qSUo2kO/5XMZy/uZbBYNNvxBudV4A98zJBQiR98UKDApDxd25i1XENRgMQI9hUS
+wmqueYtQGe4NXXlel8uUVHS5aZ09Fw+vh4eeGSP5K/zu2/poUgkTnbQfGYczdbE9jJtaehhEEZt
kmjqQvgBWmy3+j8oWqazhwpJBhGHbQ/sR0kkisf4JYS48MGTAKaRZUgRB44YY7BmDx+5HpOBMPPW
biQZhLENmP20lTMlgay0rgFpHzpFeEAINmYcIHqOdH39b2qLra3kWBMC9GjJsY5u/2caPfxEvM2t
McHsmvLXbkLeGv6BlXqhfUrnqFAPqHBdcfChMxsA8U16MJBPn1hVIPGVdvak2SrQuNPFszpifR2e
XRDmjj4tuZ+lkCfE9OBr4DgAwaYdHlQ3Gpxg0F4RuLYKON/Dev4w4er7inj09qsIqC5509Y42bsu
XQRbxFxsuNigE5j6l/DpjuuHxeK6b9rJycImYikCTLPDBUmcuQ/9iX25IpcXjzVtoPOkod7a8gK5
Zv7vMvAljzTwmPYnkErt5fIuyvYaqVpaKju/YciXW+GEf95/N8o+WX6GizXYV94dupWYrbyFzTOK
vyRVYWRX7vyivL81naZLr0pApi4z2yx6ZTqJIjo8RNoG9QZNEOcbe1+67+N9CuH8Wu0T4FD4lL94
H6uwd8HAahwPAo/1x7IT6zhQrXyxHER2GgFb6vx8CfjLPuenDD5Eawllc4GUiqRJNlJs+KFvmjYZ
BbscJEJx728FmU8HCOL/I+FMQNnzHGdHhVaGbK/DeFpOWxVlE8kV78XDCCBJltHxqh7/EASzy4nB
vB6xPqK8JXBafcB38Y2FUbzHAu0Crbs04XzXFmIYY0nUXLwSEx0Ap8xgxkROh2r5q0l6H3PqM+sH
r/StA7yBw3y9OVrTvzTqr42UPmtnSsSiBQUGpmPMb/nJWPYWWUUIBJbdWu2Sf/8g0aIsOeE+ZIAj
JLxezyDKgRMJcnwG3zbGqhcvevjs/NSV+imR+z9wq8b2Nh0EgEUyocwxHiZtffQ2zKrx+72vKc0o
TohXzLRv+Yx5/1PJkJwknJapGeL40TxrYWR2o4BvS4Gw9n4nT/oFhFiVDtXjjXQ3902b9a3AiJKE
hzMjnLceG3gV4IWIooRqfAGDuf4GmS4vJEnL+fiX3VGz/1vLOHrYGNiW5s/+YCYUSrFTwv6jIW+v
w9asF+9lAz2lZm6Z8/QwHIdOg9wXPfuPSNA4oImY8vNuXi49W1CqtliRaqO16+OfuJGcJYRHROOf
qHs+wb/YgPN65atM75M0H0Jj/A4EGYtqGtPPfggU+zWvKxt2ZS6/34AActIPgXRbam1bssVUo4La
TqS3AmH9RP+jTgWC28dX+89asfSQiMuFPV6xC08GPxBjPTNBOj31yCUN0JktFE43ZigXC0sbCDmn
OeOUT/ZzJzl+elU8KuOHGU/Ahesgj0qPg8HX/sfGKMGJWLvWUb61S/QRlmWGgI14VbZjBsZam+Gq
s/KIdcEbOv8fIHh4A7CAIGzAnLuYY5vL2E2IgGnzCkCdVCv9eNFAf5F16JxY0FmNdPFfZsLmk3Hg
xLexjgd6Fx0gEf6ZRS0+eukmMIr38qm1oe3/Y2s+bV6vuezGbz5m7aqDkKFptDmc7h/Uiu9h8vs/
+JdSU+oy9PPuNSWhVjPWn60E/tNEg0cCJXNoxGEbUzt/hRx57gbgLyzY7cei+oiocq+dwmgEQags
R5/nrL8cUDfMEUHRio4rkSCX0yH/H4zx3LW/D0wPSSor4LEKKVTTzqvxae/0eFsIlP4q/rUWNqLg
doPutvkOpuibM6Q2k9vghS7uJeHvwapVwftx7+lxCfyOaiGI09kxgASg7bb3/hfREmPym/t5OKxX
DsxRz1rvSbd9ujnx6dNZPqjTfRDRoQ4bVjaUyHGDdjzCjPFXlujVUHE5piWZqrP0zuDBOHQLmfai
Km4SKUVTweCe4AZU9n7xEl+7eIw8QmNl67G4W06PnLrQkolj38pTclvZu08bhwuhJukcQ1x4aNR2
m9vXbl03nqYVOOq0Xf3D6rVv23P2dl3lMGQKMWPZu+UbcjfFFOtlE5j2SDnknpiF0toU4E6E9wZx
iBNzhFUWTs8ueuA96oCENuVC26xq764tiaPeVc+XgMzVzmewoznYpfo1EgWbePDhl1env0KhqhKp
WyCo/e/dQFIYuvZgEVjkiDrg9eNWOE4f77qk845uN3R0iayYoTOab/AlKA2jrj88/Foig6msgd9j
GmXtDpRrvO4Xji9zu6/ExVPql0kzr3zLX+DFMs6RpQvRI/5+vvb77zhk2jmpu/PHEo4HBHglBhaK
83ghYXE4xzeq1+R7dG6XnbMkCRhnLAZMwQ2aX5no7amOVkR7ILN73ef938mzx1ALVPGvueKkUzcA
bqAEaMIwtw5A2bJ55jiJb95y7FsUkWD0WGLwEYEwEf+os+jym0e5sA9Iow34dlR3a1F2HJvh3kSd
5ZM2/gxrDlhTABI8ZvAPweAgKIoDQsZ2xrcm6zHNIBWjjqcEKQu776KBVopH66daFWB3UybHtRuE
f9oTDUZL+sFI+3rUB4jpaWrSrdqz7Jnwtvk6AyEZZEWOFrxE4ExjKZQ7M/EcpKrsmrIZDyABE6+a
g3NzD2Fspx6ETuRtO755I4MOJnvnYKxFAD/LY6ur1zQPVB4ZsMvuVhRaOGoMU2XASmjjX1Io2tKi
lsmL6CTx6dLIiB7q3PYqSUqXGtSkSQkQu7xows4+tlTLJuEaPhOADhuSOY5jZcPlJUcFD5YNC9pC
7rYQNtc2ECdxetTiXidmw/t4mIXvdzEobVgCDFFPlrIX4fZFSYEfFeD6hemVkLwFseohMIL1NWaB
fdiIRW2eYOddX6elAHIIrpMF8tbQJaezLqEILzfp0yim7sk6Fn6H8M4Baa89PpXPGionuXXqicsN
cKqWcR+siH/xldwBIPc6f8dXP5x5+mNmx9WnJHvaz13DoK1Tu7kidxmV8Iuvw94WNOpjwqqdPCWv
pF/CzzN6xPR0Xs9+En2HUNgPFRTFHnNgdVy6JOktloJSmoZ/WO1lhZpHrN42dDlTQA/j2gPtoZt7
2FoKX5nyA43W6pQWCFpdst3K0467wF/inyKByBpHaqVWhjoxkBE5jD8kTTPu+14DL57n6YCL/C9Y
v6JNPbcJpi5gIl8+7HJcNtzgxWwXnF1w7gUxue4XLeUkkTJEy/Zps7Q9bEOICMXwCZ/85q7Mw3Hk
FoCqEpKUBQve3utLQgDXJ5ubx2/7jBk65XEnde4dvs3rlGQUaoASsa2II2MraRgn8588JpripYCF
4eu+fRbZcxnaFOlvq0ckmulRsZcNnr2MjaKkmaRCBTcWCUqerWgc+eUgxUSF9+zJEe8VcTPeYX3f
8z/kpDsPC/ha8OR8vdcsrHD2QwcKkrfavu2oY2l7YpX4YSznrTBQJ3KwVIYx4+eNMTOEfuvTTduA
ggPrgp1lhQ0+a2It6Tr1Sjr/rx0AeycjuwBsUx7dKS50YE46+7vwpEjeFs2OnTmr45C/zyxfFJ6B
kLGmQMFDF0uiC/N8I3OcciK/EeY+He2aXMJpQrProQz7ccxMczf64yfWU6xIOtSuDkoIXS6lJzTb
xiEGEgg/YeqDRQdh/ugNi2IlDID2Jm4vzqbciQghQ7baD0TGmIaZDgfQ3KDyKxJp78ODuPCG5JYy
OyEr0EQ0LBGQSe4gYuGIxPqU8dr04l4tUTvUkNcHrBvUrbV+slj89MaRsS6z0NNXgCk4XepmfRny
wiSOaeqZVWArFsqwyqBV/1JrEUFOao+iGIaeqcQ+4CE1UIeWYCEmq0rC+qf26rnMHz1J5CBhkFJv
KT07rCi8jFdhh8cFP+fcF/TJ9Eo40dhkfZ1j4Kw0p1yINziSUit3UAJY/G1blj5kf9is5AbvIJ+q
9Us45eVrIM7Bf+4HkNA4c6Nw1HhM4bzjvjl/rxUB5g1T2RUnuDBDQ7o/vrQdHyoN5ERsXHxqVLWk
PDpkVGt8G43dGHJbAgMO5EIvIttpAb+gBKr0cQsMh4BWyPHfwCxCvqbO8+UOiDkdPU4mi/iiclWr
VMqq/UzF5sAcVCemZwubcYpz0UCffBa0oPPM9pM/DwybZXwPCvvItzQOLZhoeQoLuj34nuLh2pZU
5E9S1fgz1VTeVwnoIscLv2PunNtbaWwDY49JbdV6o1afuxbvaOZWACK48oPyRRkKoeA3swxPGBCC
w0boylOmLShy61gQIrPTdeXBRlEX2XXmfDggzsWnoFvH5L9jmwheVmOwE48PwziwoDGH7X0RghQ8
azpgzFknfdD24aLSBz0DtgSvse91QxYFKanwPZ9W2cIkO8yR9k/3d64rpGoFylR7zrAHQ3PERqkZ
5wXkWlyvolWW2LyVq+fNqxJAgd8jD3zihyjOe9nWWeAk/BSxtrB0Iwpip+a/Q4DFJ6wixlG69gV5
u55R/5YT+RWzEqQ0Cv13kiu2JF7RwbRUPGvCin2lkP/Wk+T2r6Z9P0O+svvNmsMIOnRT7ulPL8WC
dBT1AFwd36bUz5ydLGL7I4l5AYzhojanTYkuXNHOaOEqxqRAD32X0bpfdkhxa47gascjr2Je+wYk
qByHBxLuH4JHBrQn/R2LMZJwlcmZ1ACuwufI3wLLCWh9ZOGcfWxt0Js+Yx+qsfTEgmYXJjgd0Q2Q
AolbLAvJgdgZBJsqvS/c6Cqc728WYDSFuGlhkusf8jFByUlIgYypmoKbPCo7J1JPNOMiNntM1Nx4
M6RV9flm0Sk/mp5AH7dwfqRW4V5BS6vh4qsUDYSGcmOuKPfTPqLlalPctSlYcNCMZR/MhTDherhA
51q5IX5GCDcABMs/gIWgx8mEqHHqDkVAQT/AQ4bCDwLioPuymWhII81jbU5dNof9jb+jQLoVGioi
uonWwt6i2KlHysGlCsLzT2nE9pL7YS72dgXW+OOUDuO3cMWxFZqzbD06bYlgVrkJNHzOiZ+hQ/S5
+O+Qn/qK7uPwQ608nJDhO30kB+EvpE5bAsdrVjV0Yb3uRBASGAKk10/Bts4hUgdehTyZvRU+sxeT
iUz5BMX2b08dVDFJyW2ntZhx7pV5+D2PKnpAumxR8frezJpiN7/SV70XU3zUBfSYl+Sw3dPz3Dxc
vE7jkFP61AJPnPfDL5ke3MBr66PyvnXwvb35ccm1/BQqIVU3C7oLpEfDk8StIcCVAvmzxVjBv3bw
t4tcX3lLm6DbNa0GxelCEJizO79IgxjZC4H7s9W9uSH9KyfxblbOyjLhkeEFXG3H1Z6n8SJHrW0a
y9L0+xTNI7ZyQyIe/QQfsGbkFw4V6qQpSBlDhTUIvei5xDWMsqAJRYYUQpJpnOnT4mQSU6NQT321
qQl25C1rMkZx17O3cBMEArFZ5FRJ7t1VBcmlOfUZgscoqwnbQevf7CK/b6HIa6w3DOgG/JzIlN8P
N91fAhOnvRPhm4HDzz0NG0Wmji4hj/AquFyQA6zlNqTkiQKl9X7n8HTrz8ZwENsWfwI/xVQSpMhO
eCPN/lxUDaopX+kweBa8HjWdULw3DZKHVtDaS1T7QEdeqRxhWaZ1U4hWSR50T1qhlUgIvgscMO4Q
6WMmvPXoQfBg7s+jmGSk5BFCeMkGr+zv3YseNZez04Fz+lf3x6GzN3eHeaFdFV0eLACsz9OdVdDk
ZQ53x8nPGpS7jVlYtpNw2xNoc2f54g4613ercbIUZDDNhse7HD17AChDokiXRDjd1aEaREEKvssq
NRohMZrvtx+Z40sd1Uq+D6N8SBC8HqUYPPi05poM0l1iwwkkZf2sKPD3BClzU6Uf/V9gQAnxP3e6
Ay20dOjoRC8URzA4um/zjM888ENYSricdtH+pDu7GU2BgPFVFs4DP01K5hpUbLydJ5w/fN9BDfZ1
HzleK2Y+F2Ikt0qL3Lj2Md0FrYcdvZK1Fg7badfOwvf/ehidJ0pMCtxkiLM66sqUhy+UKibCSa5a
Yc3Y/vOoU2hRnDLbCWmiCxBuQBQbgiQWQeAPj0TYdpbwOZ3FVp/Sk8/Fny/MMoi9wG5u1ghRHKAV
pW8MfwPHKd6ht04ahqMgnF8ZS3qvUGtXlVjW5KfpecLj5Pp247d5PuiVA4S2GECxcAe/n70E+kJL
0Mcku/rsc+M3DaAaEFlueRXZF4sswnCoBYH7mDA1geclwOan0C1vYGfbCNh4f5s0SXPvjtjN5VgY
oNBz5FwjdzChxhZ50Gao8N+KwoLPmwRL9TdRNZFDqGfiEYTf57Hxd6vYnXtEzY/qRhT3e74woAvP
vk55YIPZsOLe9rrZqZmRv5pa2qv+9H7Nz8v/cjSXsmGxYziCRHgrBgheHK1RofQU9LeZsn8m5spB
+0AQtrFLQCNd9QNCjae75vThXzb7J6m/CDbqBp/jjZCJ/hlxubzuadSmJnXc2hm9TVVPdxyw3xTy
b/MTHEZ7ZD/fsg5OPPehEal29dwgLdxLyK9lX7bRpxdWs2KP3bCmIF8VBmidlYh4seinLqjmd41N
78TDYLKtAuWOgMSLHHIvJguEJT/uNPyYW6gvIMt+n0dyr/wdiqAoxNsG8k1Lk2A/Q8SInSRozSCT
vjlpkOrQ7EYuCCv9KZsYEO85kJr61D+xrTtBWTv22NweRNTdqcGZ/hrjMja1baSyGY4AKKAh3vaT
tXn9dy8meS9Q+bpVzNuzu/0v2WUC/B5Q3sbqUFWxxQYqRKpMILeUhq0dgzw04rK1mukHwoaDzwxo
yoFSIQoM/7Xsbw/f5oI1FhYcEV9IOf5TDvUEfO4PNvqejfTnwDZji4mTTT0sfQUQeFmBEBDvXUXJ
yqzck7bLGonzO/f7qqz92+IgiD0sUp3qJo95Ciql3x2GNQ1hhfAJAz7ksFoLLok6lEAkKlX0MY7l
kvnJkfqYTITqeqylPQD1k65YTd56IzWYmvyT/wiN/oLLUCeOlKEr38hsrIl/7jkau6ZWWvf1hV7u
T0JDJz6v0og8I+1CjLCB9zj/lKJcH4QbhyOtfIvCpP2XTJdKtK+Rq+cQHHEUNiZbaRmc9W+Whiiy
xLzBxLf0Z+fzKr1hRrzMbqUva3ixkNdbiAl2+27bgkj9zomokY+gOM/i/OUAOGhgFYFXQlLONf/j
kn5B26Ve54kwQPx94QjyYnN1OWytgHtAg8LkojTInpSRcNWdMqToKZR0oGnekLeTzVvIkEcrF0FA
vJ8BtRS3uOdGMIV4vjt2hfyXNegFzYyJa7xEybdpAYZ/Sj/6H1RkKBnvQ4HX8bWYhtWBjvzqxamQ
ZK+oet5n4HwxgZMMcBs1ZBL6G3Cph5uoose7/tL36P62CLU6ooNqgErZSc5h1hAG+fsh5uLt2yB0
9uleGvfuO2iE8tc9e+sa+Bv0mMRgGRYgKhUAkWU1qTAG+sucO/twn9R+I3AJnKqrCgYZPqlJKWkR
aHJlcGIIr8Ek/d4lHi/7D7KvbOvR2hynNEsIwnOheHRQ5O8ceTFbReTIgIKq6893LoquwdK1829e
/Ckzsc/iKPG3tiYnSl5B3NIRCpZMGrxW1aENYFMv5uM28vMMFYI9PtO2gc73VnOrnq2wjuyaJg6G
tdi4dMtPQl/jyhIDlgpAX/2LMU70nT5EUpp4/6T2pEM3bm1j21PyZnaxeFw8p11SciP+7Zb3ecmr
qC+FMb6vDzMu3tyH3yLDLAbTVR5sgPkPaCjOugQPRRKXJhELmmPouZsuOj8WuHEjmPK3OqaTOKAm
WviWqUp0QwOAJepiQWjuHXAXN9GS7EGcPcYpmN7r+rBWr+cexMctEDX8mLCoS0h+IyjK4xY9DfGf
wfbhT/sn+YdpH5cWy0QIqitpg7dOJftBelZBAryiJ5U24lewNbBpZCy2vGAaxprgLPHbtImYU21/
IzCyTe3j56wkg3b7kC7HhhNqhkwHeJYPAgbSniuPbZr+f/9sNqf+ynijP93X26WgAT+mPAHWkygH
TCaSlbPYfDhLhwwgQJgh8nbDZR6A+Hlchkpfo28WWkVTYzjF3p9/RYMkUvxf2UMsKQi5eUzvnA7M
IrKBLjY6pE5FxKSUWyOsI1VM3a4RwRJXdM/K+cnJgmG7MsHqFQavNwvc6iij8u9NVh78DKvj7Ypa
E+dXpVY+OcIGYCzsT1m9erwHmaotysKdBXv2A6/6cIcO8ctMZFP1SsDHHm4uOFTMNgjEfcZ0X+6t
a4c/oHcckR0nd4DH/r7Ni/qq2/pMfhU7hgH/ohe3VTTyhyBOhExtVfSr7uxfaUBMv4xfS4dKqK1t
Y9c8528ddXBnkEIAdngFz785umviYFhpoPrpkTJtuA58f50lJhQnMl0BYy4zI3A55VUw4DF+NQsu
9Ewysq0IJubV8dPHNVHtJ6GBPY1+opwSL8fsmTqSEp/1Hp24uTVhZWrFZ3Cw02/ZnTdl1nKoZA17
nzvhJktGw5Z+QKoWlwgHSPfW8cDuhvzdA9FfywB8kg0FLRXuSNKL6EOVlFGsbFYPCKMDhY1TEbos
cBoWfgjDZIdZNYjimajA4KXliiQxxihl1O82SwMvTf6nzCi11sq6pYQgOCg6VocRNv4xG5UC0Kcr
UeT8KldPIu9L43w4SJHZ3cDsThCbo8fUTl8bsF/khCFDAkqu5MK8u4E2QlJtfS0EZo8HqVqrGjFA
AwGI07zLE2nd07R0s57YaMLqNvjF/fHh+oOlH5PlYtyYFhG8c0WCefgYjIs/x/cl4Pv6JZhzroKL
xh+iyjYwvDN/fh9HxkGxRPMuv7XrZr1Sp1P8K2BmxTqeZ9Fcyi9RNkiK3cTPiN/L9i8h9H8bkXGD
mak83hOsYMx2uFk1oKl8Ju0P0sQuBMnjRbNQBEyY1z38I+rLxJuX9LotqWNl6HfscThfigW3jPvG
469z1aq+3HW20ROl/V56DFkhcSId0DlD0m4fXo3HbwCPeEuzs0JR8VZH8p7BAgC29bQHjmL2pIj4
S3gdPjLZFMwaQq1ll55Ovaunf8EgmcqZG8zBJeyG9aP+Gp50d8fMowJdss3AxeLJydoHlXzi9X3G
3gbEGzAzpPiZWlH/aikd8MeMmQCWsVe8pyQU+qEQOWxXgOAwefrVWuuE30I2OgiQV0njOuX0i5Je
ynU2t1BvmPl27FsR7W6Gzchh8qlA73L0WzNyHhexW25tH8r4oXtJAdQhk21XwHk51+MIW+P3wkMt
3kR2EN6qJ7m8rd4y8ynwQ79qI1I3N47p/E6+TmYQevQTYuzuyrqAOHFz6ie4i+HCw0/LfTGGNSyU
l7EZBsy+ZE4ofWxjzUVPQib/xws1Z6XgoMuiTNQen4QVdQ+jCgxDvxzGHNrYrlCrK9o8SecE6w/B
sJC/Eh6U7U2u0B+fD5ycwXjec1Cb43nAiJ6KBpOqL+4eCg+zUzTAp6f8TlRRSfaFdQrV4PPSPuJU
JGsjTluIm+dS3KvWtTTjSTiWTmXxM0y3rP0n6+3pVbveQj/dcHZgny7/giG1fCnGXnCIHOaldAe9
l4RbYtdLJzkDfsAh+nzMvsMQQfWBVg6/CfYPGIfg/aBTCNnAuvvOsQWbhi4KYP5NZN/xz1Sd05Rz
nhkZoj+VX+xWtxvU2fmz4vW3bh5JApUjHQ7cjbld3QZFqi0yJyvE7dE6J4vcKmYf6LIa+lUXAHt6
ey79ZrTsjpLRognUJEnxvitgMJEn8dLihyrzWNaSqR9KwkWv1lzrS2L55HTVufwtvM8BvhfuaCYl
LHTjZeqTRIc8DesvTgzsBuKTbRRz1yT4ZFruJGsCxIVTYe9zzwiRHFWJ0XkqN33rUxCqS6Nu41TM
OTHn/It38KZ4k/h9Cg3lFmBlpfag7vH0e7/tzBe2INeylaMbBLFNy0vYzHfQd3CWZWlUGXE08io7
mHstQnqBQuS+YLooEtEA83NxaUZUU1AjjMQa23JQIRLQoGSYT02B7rgfjQC21FbimB1tvVJB/Qvj
zofTEF+CvPNs/kzERCSS/gUv2pWfusbhbVKjoOZVZn+rpGKxnor9/9QY8kcz6WXAn5N/06gaKI8d
MSfHDVCf6g38+6DKOZjKt5RTsoRNygqWx2TxQgQJtiqrFaaoTY3SIlBoMINyIWuI9GSLCyeuhpds
IzoYBLIGSDU5/iZH3qxde9LyeCNEe/Dzgl9E8aTv9tr19OayijC0aAKhDeJskx/4jOW3eXqpjq1a
08nXQ6P8ImpNQhHJYldVrVqoyqfWaT/hUtT8fxSuGqS4lYs4LRTZhvYQ3PBzlbqFdpXEecFtLDQl
UlzAmmGe2E8BysHrsgTl9O9UDhkfeHXWiImvFUUIgzlc/exsH46cGY7jKkvbY4wGVe0a0A6/wEPd
/nHezcc6yRtRyu+HvgABgSwEgK158UWlLw4F2Bmjo2RVgQIaJLdVUi+eewOkBBHZTrszi9ip2CHJ
KK+9P5j+IP76MXU8Rs+VSrijEadFmZhNNcPNz0/vmgzg+HgFLorLzg3Ruwfzyvkpftw1vOuJrv6S
0VV87ZHXOBHBs2Cr/V+sQAtgtVIxnZtX60qXirIuk8EoNxBgcUHmUMTU3vvWU7Dc4HgiBFFBh5zm
nTcgnXhDVApY8coYGYr9u7l0jwuJAJteBmFz+GOLLyPNRqTNlmZTAOYPo1UIrZfJXPa+8wX81/4h
erscZ++4sUzkrSD76mEm9DaezIK0dSoVPnALlskD5qRhLwTU7ixfIZTl6EsiteemIwb6PaVXbO8W
c8eeC1dXrmrKFFvo8wMwMtyic16lUDK6CtJdNc9yYt2gYRlkzWIMiUIEiW1vvZ1MYeVg+lFppJ/E
DQYInphhWJFO9MAVxtq1WJFT8iKuRQBsKqFxHwvNfNYQ1hTvNrW/lWktPz5ybITY3im+UzShlol2
+3uINeYWyZS+UIOMXH8OgxuQ9/mpJGKivhtp4vgheq2VijBbyWKfVzzEJMowBEKF6FEFvOcr93Nl
zwpmFKIPeGfjgt5mUfw50TPyoCDmuVWpnJDb2NBIUaA2dBA9Rfn/kMkeuF0WpD1FRLymUpEDf5S3
CWoMSJl8s5QHNr7g29EeNlBmGP0BSZrCewtFT3tIdVtMkFH2w63wHbDY6mGCaKH//xMHSVJVCvNG
Gd+3naftVhMl1YobnxvJDObQ9t2z/w+goWQvgXe7kgPX2df3o+yfA/MFztIUPCc6e6mvZ3v5z6EA
FMEm1MiOf6ZwI9WcAcYGZBrlshU5K3A+mrxO9emJcrfZTaiy6+quib/wlX2nSbybrX7fFgYkyzCt
wjYeCuqV4MD1/ei87NJhVoex03CyaHB4UsslBW2vaLsDkWkxGqNQKGwGXwiSUEg1Tg5zebhx8hQB
LuKlNMfls7tA+c3/5/gqZmJcv9cHIT5aWNqAPVpHzOVHY+hC0WW3kQY1VaZNYviqHiJMwGFjZxPE
/ffADIP1lCnirJIH2IzF+shuFEtdD7qg+FFw8rN0y0+WkB8pFvuSzydQ3UbpQp9W3myN0ULHgBnv
vwA5AsIhU4VfzUYKAslLx3L/C3Nt8P2pHxJqgz7HsRUBxA9DA+NBuh6zauQYjlevDJJ+68wPzE/y
ob87z/e0CDul3lF2IyR850E9bT9OJ0WqrbVzV+7KrGp6o+5dnvvMAa4i76JxQPdrUjgNHU7kRVhD
PIhmo1op0wFV97nqeBljf742bcOfzGOKH54e4JIFr5th7f7ObFKiDHoJHY2YEKHnqhQZH8BhFnZ5
eLRqNqDm3LJXGp/jEoiD+Uf4FaaRAHX75v3q1YwzvqVeMf+49IhyjjJ0qjr2dzUdLrusEEk7d+x1
LTMDfeUsyA6qEI1Vk9sPUfeigjECxQNZkJj+nQJQwfLxk9zNIubrgxDXBLLo0Lyf/Z37VQGyKcQa
bBPMG2ohL4kfsc51Z+w3nv8rVIZnVKsdDTeUD4yxBjXVmhVLoOKYrOZxvXJplBPzWyPyiF1K1aTy
BE6l2NG+f3x7pXclXNV3OhWYodYj+zd5bt7zkoJOGA0Yaa3xPYQe5ZPA8zkqchT0PShjcls2ECyI
GoD9OtMQHKB1EO1l/cYgd+9dOCvStY+n/qXip7802LPzXQhJHcgew0mrTHcmNAfG76C2d2ewBWcB
cv33/pGMMOd3qBBbGD0jHiKaAvZfEI02142rbX376q7zMC8ooavr9QFbBRF29/PeVk0ef6GID4H9
F+AFViHKSUUkrbG8NbUr9A7DcZ472igX1YO3Lb+qcpI8HQ8Q3xw84GDeaF1Wj+2wrn2VI+wJ8+rl
FxsQT/86HcxHuY0A1ERYxcTJg0Ab9Kd+sBYyD79BCOkO/0kI5s4MFChtit5U5UOoVHL8yH5vRJSx
LBz9MkTc8vHeXYlbj1Ht4JCT7e2RW64+cQlN+gPDqG1pbJY2oL9hBBb+l9LyDXjbvuRJAia9Ug1l
PfsclO7paczi74p+LsM6MnNaQRBZz3zS7d22Z/qX/aenC/kKSJ5RREc+XYbKHuqvUVQOfOgVrPpG
mmgnvQUxLRqVaKoSnv+KdxQiCIDVMbOMOUOo/jlWhlX1jRLk+S4hUzj1h39Is6OCCs6GW6STn+rE
kOWIdNQTkzuxL4EnwxV01SUuUx9DhMA9/7tsE2vTyh+WLRuehFg11xTpkmF4CHIOAWH2OJuGGNM+
iMhnUrGIhgjwc6ogAPdLIK73JDv61d3zZdvSk6YboVKVQUBCglQV4Kl/g9rVmDTw/vahXIOZfZqu
V+miFO1SV3fdIsFFF0xBI33mV0V47uhZSpbem7xupIWqxx5EEzBV+zOgXPOsJOuDdkwSwcCDvIvj
RFBT2N56DmNqlkx/ZR8QQOW/ujUmjI5yU1JgKUP6ytltanzN7pXYDK/3GzrfvG90qGyNE60Q8mAx
KdaTxiZuemL4qzYu2lZvhXqwPIxX0OOFcSVIb7q1ss+4M8sTccTR2PQ+hpskpMFEwSvniGgSg16u
7r0oMAHV4Pi1Iz3+n6ZMyedSnxdJvqVqUc8alIYXdU7QsQxu6JY2M6ZjYdlbDLku+MDZTYialDe0
60tNjbde02N8nr8L1mohSt+Sb3ly56GU9r+c7wlp5KJYRpJvZwmzbw2YIIPY+Fxji0MKlqOKYdvX
rqoRI/9VhIIUt97vO8p9eyvYUkjsrQ8H6oTpqAoOW2iqATMzZ3Zuo+8iWS/AF8qv2a4bwQ5ft2tr
iNf03fJz4USqHB2iizlllTPEwZ61iHQBLwXFAK8yDcI1RBmBa5oqFEw0Dd/AFUZS4/3IA6NJBunP
Aof85CgaUwstn7yqBcP9BtNNgzfVM65hWpnmfwMSMqNL2VNFN/MFBK+7JENq60yrY/AgAvVk/RG2
aeVf6TH6ercNq5KQg6N5fmlTXw8SLT2ZdsxsV+h7FHP4TUprk84tzletoeEq+j3/QA+85DuHSUIW
xvMC/s4bxSIn4BHJ97fqBOLbzkH+L9YZxHOY7AkrXW1GAuqAnh3o5jIjzgIGbu4EQG0tKwtgeDin
WqK+7lWzE+zTnaOVyk5AeHO0jSN9nfUxueCcPegdiJv3fs6BtHyX1TSOleVA6KGFBxzIvhMsGaU5
TEkta2KKI/z5UViEl74ficshGqn4BMW7LxG/MlZIITtcceYyZcumPeCGnDVoKyHrWpH7luDDykVv
eJ/ejDU5sLnwdpUaoFfMECELCf/hpRp3ykXfMKQIM82TcLg3ig+/B5Jd5rmE50JBRT4KfdUvOD5H
U08fGHDv2hVhSFzgo0PLwr4Bv9fD6q/YlfeG/HqazBovBDY52y2OCKmys+Z2KSh5AXvGkhQzjrct
UOI81184GBE9OBZgRUl5pRJKSMbIC53sSFLaGgLRo8QpUNNL4vyrM8I926sI+Tu6bNXUoNz7atDy
XNxGu568oDmUmTIcIEds8g0K3v+BW6OigZNUtHkLwsAmqHtRXZdo6oz5GD4RBmsrwhQ7ndPxoMeb
ga4ULnJuBsA0sqPhRBXBJIMm069X66YgmaCeSjhmnQIsevUURk6q5I9uK/UDG8ZkuAy7uMFXyea4
jgbFWZJt/lNSJcJrh5sGXpBCgmVlTxbuDIfjCz6/rt5ZEvsL9/zteJb+65+InPKWi9Ut424yJB0N
SzqbxYn6wyWwSI1ABrx7eLueLcljJLVL7zdyR9KEgGvdH9tBSApeDF7UqRv9pb2e/hy29KN32vf0
LEyZ4XYCO3s94LSBXj1qTq10cCBA5Pe3JWlrTsF6xXGfLK05ab2L9FTBg7jz+apDy/O45qS9aog0
n53s7yNBZbghH6hjL5MLm/t/7wgr+MZsm1+mSMMXWNNy5UPdeqeXCu5mIVc4+b07jqHsxQTl567K
Wlq719zZZ3TZuiKviSqyWokKEZaUupYc3aIGD1G75oRjyNaDbxbMqj9XaKjYsG+c8yNpuPxEtums
nzm3d1TTTxr7FBK9x30JHN96RQEUD+cY0JQaFIZbOvi4nyXwKiacewwzFqjLRLoqnA2yEFxflB4w
Wkrm+N9vIF4R/Ifienxim6wvWlJ/mcaja5J/hNRAK4MIhh6PGL0KA3TpUPhjeX3B/77duIkct6d4
NTfLjl08tjNspdQMsd4RXCgBomz8H8UvWwkS6Sa3GwQsyZsf1A6bMbQvKV4VCepP7n/yHR6f9mmu
3A4ol5ezV3XAZ5yErAgeGkxVgwjdo4G1GNn7QaEbTJ20qk6+k78vAQSHf8DlVNOlQkv91Q+r9Fk8
TLCVl1CEtvsqMRasC5ECm6YlXV6JaDyAOZXdaKviUWfG4JwP0wCCJ8L5GCulCggo3n/9GexGJOib
Tfj6jNeeSHz5ZGLou7oqeKOaswoUd08Nbjb0xFpH2vaBrW0zlgLGcY4JsAcGQZzPrVAZT3/tK2e9
ux7SIJNPJFVnJ6vwpImvTgSZfW/dYDKWR86DKy+ipU8RcCsMoyaGTT+y6y2c/s8BuN9BaMtshVA2
CPb5W1HcAM2NyD4zdByqmTA5T2oFYvSZPzR42x6BcYCX2vAkbIdA4eJjokZxPBdVQEDCu0X6IqFC
ewYHvcWXcoUkXCdsvMxZ8kc4AnOrxemIEGv6QiFUVxdY8bEU66uWiLkBQ0fFP22al3TuIpUmTUkg
OJhaShAZDJNyEKTD8gG0uDuQGluhc5+rGmfMF2JFVUQyLG15mRa0/km9Q14ZyLsXRONqH/xExu6E
EdcJHuKs976dghFnrjYw2AplBkUzLjnhu1SnsT9ZpYrGOnCc9H5LiK6HIvLPtmZXMqUdWdA6NIco
JvipbYealCbawQHswpp7t95Lwe7ZA2t+lur1rEicHYLdSEvXkilM7YQWHfFLwDntUlOXW1DZSL9G
+Fed8qgIdwNTICejXEA6gSNM+G7WNpnx+7Zgfjfmp3MaBqN1JDSMwoQn5yyCb96aYtTmqGzwoLq9
UaXph0i+KVrj6fHVsx0gwOydp9KbJA4WTIOlFokncfGAWonmVgYti9KUMNcMuTqVCkytT88qf01Z
ArlqKAEo5ZZkBaf7Io8J+nb4kyTA8aB75b/NelfdYzlqY0Z7RPT71Z53LVzXdvMCsI0wqsTl3z51
ZvqiNXoXJsoaLho94fCUiNuleolkdEQUShFL8/Qcj7LH9kCriKVX+urAGt/0wSfMzKK0YWSH9Hbj
gC46VSR9GqC+7d7fGi9pXIbbQ6/3HfC0FpK+jX2P6fiB1gR+lmkgQOm+HP2xWemODy3FzKU7hvb5
jo95jWrzKYi2hzTE8Fyv7kv7iYbEBlvFFUaA7duz61B5d2Y3abq7udbEaHVlHd2+Gx1sjOWKa5nc
ClRwh9m/aygd3oElUt40Ob8jEcU/TX4G9TaRVis/0jFgH7sOC6LfLnPFGPZzgYp6UQ8BAWpEx5+3
9ueP3f4gZ0sS3YllSkRbyO3bHlAosmiDhCor+wktCf2qco1EN2rMS5d6fc7CzIt9KdWI5rTStkfX
zBlW711vl+FuAAnzzWlAgasm3GyOJzGfA/i3b9BfHkL3GkWqWH10nxVd4+3DgnW4TawTVTsUtKoE
9UQmTwXXDYYx+YpVlrks0i/dxDNzd48bIX8g7FJpOTFIcZBGQZfgbRFAJLjx9TNM5x7JTQtpd9Ci
u0ujBjQvm4WjPmJBuYUUBFXRl6lb0e895R4Ryk7gkQdAvq1G4MtnYEaSRS8vBhTlnG7YbF/z1v3z
PCCCOQ71uV4QwwoYwYEjIPmj7i7YUAvbEwZRocfSQM1BfKungxKYDTVWWyB54spvcyOXZGnk0Sf5
kJfVg7Qmq2UZyklel2uu2Ir8Ir6reEK6x/hBvgsKXNstaqiFzxbG/P9oP+ViicbwgkSgrH6PHmB4
uYWe9LqD36H1ZIysSWZyE7Bm6IANtAL6WFFmh8iq1gK1wM5aGl0Jw6NAl/SKwdfGeWko8e1Gr9Wv
zZQUC8Wn566KiDCaLHVmLknK6DhR53ZFQuQFP5MYeJ/SBy/CkQJGRqZjqmLYYSsZR6WT7Src3Bcb
XSzKdJ6KHUCoIwSwt4Ox4PZfwRTymkrGSMmokQ5MrYf5L7ODW78S/j78T9mABj6+a7Ew9tadfALz
LkmzgTB0J+pvAoNt8YXb7Zz7S90jOr8R/QFv2E7YVuy5GokfPyX5lpSZN/kZ0VnpGJSDzg2RgZMt
3lfkipTK9GrZBhSYO91of8mcHyLmOvd1UccO8ypLTvVBz/VYS81pEI8MNw9fSjwmIbskCHjdyB0o
O87Z6CdaZhlEPPFdQzH00C6qpZ3TDCUaZdPa2xOQYwhxHIww9g2aHRwvs4BoxORsRw0j96zFVWxi
+DFQKsO19rPZDVWGUlUGqbL4AkG6uo6BkU2nnRyyrSxv//NEUTrXwt3UTvGB0SSYAENtdQ9/lfGt
lsA84wAV3i6fmJ04z10Z8Zn4k2+ogyqbvZ4w6J6hLxb2TLQ2AolmApVYH4Fwv1lVT8NgplXyl+s3
wat334SDuXWe+P+7WvQsJseGIlGcicFuhpaqlSBt+BqEQhsAzq5gxMzIqrv1g42QoO5Bvwcd2Ikq
BUmXPWv43EwQ6y3UKBQjBOlY0yf2p1O93KN8TEsNkWxENEgdb5WLJhadbjrsvv8NGi1glUPMisdC
QF1ECUTBlhIXkJ4L6l5R+6AXknJBLQ6kbx6wlf0xxLrvSBJPzPtcIEO6T+MT2tnvJZBGEL934pQj
MVifpe45T0K2XPeYa+kge0LCBRIsX3CSh9ZNvbnctNnuNXiGq0dcFELrBSv/iiAx+zq03uKoGsxz
LJt6v1i5k+OuRdMnR88nkl++leO8XXXU3ZmG/hLgz/20dIQFcqjFSBoOSzCI6IfrnNXUp6uLrQ5X
J2PYhbZdsFCIxSW8mBM9P8i20O3od2s0vf4mZ8sji/6Ac4Ze2zHn3CM9txjVkwEduYIbmhhK1m4S
wjyJHLUfc/iEgDts35y7nmQK4M21IZwupxSLIGcKcfKTOLHPcc6ninnC88L0jtV6P2JpAibo7gNx
nwqvj3bdmoJWMPNw++lo7JGFtah9xPm+OalLOchnmSh1YcwIB1BhnqDVjazi9Wy7AdLRt1CKtYxP
YFYJMLSy/hyOFN7PC9AYXiLfG+6IwZz5ZTtc/UXqlj/38Q161t81s3ue3f3VhM1/0ttQlle+IhTR
2y4cpCIQrJM//opxCZRS3D+w35WqzQzOdG6Yk1MEYFlhwLU5q0yoHBdrk5/NnkgaZTaAMvV8ECs6
O2F0tFI8W8+m1Fzll4f4SqHmGHJdUrRtWgGNPUcLxPYpMZzVdtsaf4bluMkzu+JXpDyYb4UmSL7K
pNM5AmlyWTKrlkXqIhc4L58sYpyTfmfC4AKqui0qzai7vxiBxnhbHq5o4OeI/Zpu9YzCC+qErFga
kiOaEZXcC9Cn5rFHKm97P6E9FdgYazyYP5pZD545P0gpD73/EFSogYrmdX2a+WIiFtAwwfUk3CTl
lwsOPf30X+nMDZgbwcQM/HUXjtHFH2XQJXu69/0Il/1+DsdwXTX1JUAnzApUvPs2600oOwDz4nYH
NACTW0fmZCFJM+v4bXiBLh5NXbX0PXMHqrbcaFHK2NAa4sP5hJn4a4h9C6bPptfn4jY71Zb/sr9y
Act7mDKUfMTplOnKUh5j2MR0BW663ucS1dzYxiIgaKNKz0PLJlTJzrcvz5o2lNYdL86Ib4rgSKyX
hAAHrFCa63krEkE4zppmK/qzeJvZOKnerSn96lhOeI6BCMQGDRFIBgaEI+/7ejIqfhkSMD40hATT
M19SiKW4HUhI1dXmqqlAunuWdwoeygiAWLQFWYSK11fYH9LpGseJNzeOgRxb8zB1exCzyiBGH7l7
uR74BIeDD0+LKYMu/Job9bfqHst9zyAhLEJrEKZymnBLLSSXmX4FbuGyXmTpEZWAZEAjNNPwlE11
RWPFvgRxfImna+UmdroAbwcXLbYbPeNiJx/y/ZccfzEER6PJKVckqaJxjxysUe7Q+tQire4fkca+
uH22AegDvS3+A7uLxQOnPjB7hL+5IigSajyjUwH/m/iFcrbuwb6/s5NgQQxEvQCcqZ25FSrHATu9
GRI5cCAmEdVnPib1dqYb9zzqSZEQPH6fbh3gadi8n/J58rZYPCdioXjBSTKMymEojWuYuuR+94kF
WaX1j4f1TSbmRgwC16U6KwXfhSkDM7vwP7GxBkJvSIE5Xu5ED+Q5ar/eIOQrWhuun235/noLf6k+
W547VZbnhE3kveSrcmKfvQfK7/m0cIdzGwyTagoX4gxf3dvMYNo0cLMIUZ1VrXYghBNoCeyliV+B
fnKYFjeZJhmYoIPKsAxgAnCbrZgzJCc8krfs0Z/3YFvnB6f3LMlvzp54KvnMkKcXBXiePZPuF01g
c971raQ9wfS0iADyLggff55bE+cZRH9dpweQm5T0uNxVyE1BwS1w/oY+/w6OOQaha0vor5cKNS13
BvDtPC2I31xvsy0xEJz48C6+tqUXBTlcP27+paSvR2oStZQKQatiFPIGo3xIIw+gUZo1KezD6PSX
8eVTwISAlNxkvSeZk4lKDESfXDmfwaZ7R7K5UF6HMACiIjuZIJQO5tRrGNm4rywpZmeQjr4WkH3T
9rseG3Bi8Dp0y2BPGysn/4KoMFWpXgCAs4avSdSAG7k1BpULn0FGT5Qdcp2RSs9TXSdQZVLGQgPi
dogfTByw+/Ntx7AuOrTm2DoTvonsuGUiLFZ17gee/hr5OAPKFNgEq05y+P25AlbnvjS/5ERmqAQ+
N3z7eNxUro+9wfQKD6xtfYI+2PoTLEG60upL7piSAnv8I6DK4ujWOnd1NIVnspDSzl6BZW7vPQNp
yEA0jajgbqC8hdghdZbzDuOZ1crMBl4hxUvAfcKIsK1nZWzAqRFTH/HmL2mD4ZSWgYGWO2hoKjrW
poygR31gx+/RWoB7Z/3rqDiccu540JWkMrLg1jumWrD8SmAOi9RR1NYRBZfxPYIGcqut4yavjBv7
Hnl8ucUBOcjNA94WpuyFcpDngH8+Wkivq7axdbsdDdC0HmZYnuZezMvudU+lFS5HTuAv0fgCizbQ
4hbKeCF8dS4vwnkkzP5ZDG3MC+sxSpu8YofNy3/3d9m8cwlEUMP0TV4mcR+gvYLYazqwbBcF6B+D
5wDVVPP9ASxeAb4hOMzd82kAvCQkiZGliJyrBB0b4qwkfZ9lYcSS25qhIhmQ/3MzSk1NV0JZA6dc
7K612X6xqfZg6wGtuXxTE3mM1d7ct+vSacvjurtqtIdxKxOcTTxXwUQuuBRYFEcZapOjT1SealM7
8QP/+8V++uBGO4H1DjmOGSzUtE9gejArcXHP2+2SLDj3OBbJ5kaLJpVUv7By7t+P7J43+frGkk98
2PUNuy22efepzQHA+RBC/t5qQCKsNux0Kwq1/tdl+hAe1D4MINbCl3on8ElEV885YltlP9ovo7Dh
wxhePvWiBb77J3lpD5T1bLI5o4tP7XvMnC9GZUQmsCCp59wYzrakWYmc4Ya1XDowcWoGRNVF1q/C
z+JukqkjZ8l2u1SkvTw4wgx9CcnDOxQoyF4NDtS0szz4tAB8z2++JE2i2lSAYkopXYUY1yUN4jun
rZkRn06FTL8NsWGtzvEykpRmxBRSYHJi8z9r8wSrOKO1hzWY+QKZ8ZbBXXdXkBgtXT1RZ3cu5Jtw
sydVas8SFp+RfkjqFbkxW9sIxptoKTRXW0JclVvbmtXy+E974c91+QzDtTDdAh4ITSP7ikQ4dwm9
XLA+9TQM30xy611cSD9FAmlvCBSaN7AC6mfrQI2OIXjjg3VUp/xr26hsN703WBqu59ohgqqTKwvb
JOYH1Jjt69syaNCNwjjDU2nnBX/adzJfKFwVo5SH5eXHDBfKkKmMh8vowshs0U1RQmie2zKH4LKv
l4bVYZZWHB663ETt7iSoR/nf1zoi7hNMDdLwT+/p6wy9C3HTwgtWl2anHh+LfhV4CElUkjaBJolc
B63E0pBZR6nH1nIPEqRGbkgfsVLxRYxPpx6Xa34SPnixpBIRSUxNSMMOCX7dbbXBsAx2WIgU2LsX
8bNilf96L8KsDsT3MABTLm8UAvRyFF6zRHAbdN2ceTY5FPdnJ1rEZRbN66xStgJuoOVFoGDMAdDZ
cCQyxb3AkPrkBoDKuNgIDh2difCRl0PTfcoMjLYEbJ0bfmN3ZwqqX+3iFhKPaxoFbGgiezatvAwU
LLShWLU807EWxx8PJRHtqmRPx2kd/+lZbZVIfB82Xn0r+SUZdbQf8JFXY6iat1tlAwvSQr3jYs8E
njQX6ab/F7IQrR6/vjT9is2d8usEwAIgVPO6Us2lTDxqw7w6ucuY2c7qVC1HuVYLpk/aaLcGNScq
vyJFLqSrLGN2iib+LG3CGkThT9RaAh6JdmM8LvwA87Y8MUxfjcD0ULcrBvpCAtAkcOLukDC3jGl6
ffHUw/LQPyiejC4LLW/43N/ZcXUMtGD51Hpm4CL8rJ2HjCakBFT08vQkNAUo3bY6dhPCdqaWYJCp
lkaVW9W0sGiHEjDZEHruxndDT/6Ohh0voYf5agZflsGnu5P/KGdN5geJ4QryWZ1NYbVchAHBmIsl
qWAJ1TjYjsnunBpmLt19MHu3pOfxUnm4u2NoQ8gsFt5vKHxCBAwcSnkRINzRhfWipwpm0HEiO50h
Iq9AEb+MYwGddffAetymEL7FW8Wu+ywx68eAAyg0coctCVxfSzLq5EvVQ89dDGr3Y2me4MpTLMfR
jhoPmYcVQ+BecANbV2rK+S3T1nwc3UPBHLbZTF2xgmPLXXItpYc3k8/B+bz4I6u8V62QDTZkXHz0
N1mZOCw++H/HtpQn3/PuRDD96JD356DhoOUd90Hj1sryWEv5EyCf3aXjl3fk7977zR692qw2HVvI
BNNg/HsHMftwdI3ZqfaQdCurCsjij4wDR9XGvD+h4ERceNZbKbg9QqDIphuMmDFyCaqvR7U7gvoY
RxlNFqYrIh02gKWvDRxQTCHAinVi+yPeR4+svW/6E/T/cxfwne3ZIfaLOrUE8SNhkHpNsshJAzjL
eyuzbDl6zhGreNnV+S2ta/Uu8wmIoK0XkBse2jesPFRfdCo2dg4Wmpt+pDGdlOEcPOhzsHMGkdjb
SLT2F3uf+5aaWRw+LNzehjt7xtRtKzrIq8JyXYRAFqX8RSarg2hbLG5eAojviZh1YA5ri6Y8uEbf
npsfH0u62bBb2afbqb4QH0G5PMPXUUouXueuTLtcTeK6qLeZIHn17FznwEV7yFk/+xG7jva7A4p/
Rm8B4Nx4hW2khL2UXa+NsU/c9bsdgMKG1vw2O8Geoi7qjuKk8h3s0zjH48nIVtLGUo1RO9pOnpV0
TQfS+/dy5wWZGKNF7TkN48edMNopQQqJlITIT4iTd9a2yzMEE6hG3wrLrs/oDxoMXi6DWfgoxYvI
LgwROU2IFlztV6xT+2tjxR3QbyNIGnHAKJAgaUOuve9TgBDjD+pQNxGd7dNYMzAF7xBpXH/dfCtT
W7SVDmZBJAtaU0U54G5c/GFMEwofm2pt24ibIE+65WHD/xYgPVvZyWAnO33jswU41v2Pa9qoDgOI
e6p2/q8ICVR1CfDXVk+qvy8eObV15nbOblQLWjnEIyg90emVjdTlA2jySrMGs9LCwlLt4rDfNliq
FANmnstFtLNspnzJLIC2kE5Jb6gD/kGuqFimU9WyCE2YRwbQt6j64J53FrO+QlmAD4qoHZuOWGuK
Vmulr6qq3nA+ymJnYDaNkfOosKxYKid+MsiOvuHS8HidoeG3K8rYGpfPPSWLrjsaaYRvUM5eiqXN
xhMylhoxeqb88BblERFNMU/PjJQRlVDwmsyxIlagsH6ddEfpJ16dhp4PU9rPueMd9Mr743c98b2U
EnoDC5sbOYa21JFHRn1AA1GpCRvELFRIpQRh6kTBSfxHonkc2OgSLgZOqg5Gy5dZmG/1uQlEkvaS
Nn2GYkbfGPk30N2GZ1FMcAZ/TX2UZOyTzJaswYdeb4D34nEYj4r00mfDVDT52s1GD1FPz016goCc
kaAtSXl8tSusJzyXuPz42LckcKsQ61F447iIqhQIUqZs2Sx1zaoOInXsy76BAzDjMq+Z14qU5hHz
y05WvlyCo4aor72BKaoyNr+ii0+98cbkMzBgxy62Kwaw+nNpM6FG5GuHsL+WFAqCo5/FNmWQ39IY
wf/yhQSqfOktR3tb6dMcdTR8y4NaIWKYo9KasuCyTe4wVHeAdJOeOCCCopbpKtgu4JBcecVqRNZV
+4zxSOIJJQOs5vz605Gm5OjMNJblgU6wLT4NnmcIghfGorZCCYrPsdJXrSjfWyG2aWNTVfqo7aYi
0LguCtgVqpLVZJSYAJYL5ymSLrMnoxQe2GS1GrrZ2PPRNYrrtVbEcOv/DUCQV3KIIciUy+5sG7i9
byWQezSU0olG5rHqH38kMHW7OmiIAbrkFSC7cE3RefQbTu1xJeqCvCbxz6vr7Brwk1gLsnEAydxH
Zc2EQo4lONj+1+i/9KG84Sugaf0k1TFBrlPuVONbh1NnPcIBHiOcGKtELHccHru7gxr4ToFIsrZJ
Y+dXHW2HRS6msjtr4EftUB/Q++E2Jy/YVrSlzeKftbkpUvCUOjXr5gYenMLOF+cGuPumTomiReXv
Oxw/Bftbs6Wa9U+TEMH3o2Pf6eJIxGKWjsh9EsU/Lq8i+Bzrw0x+M+b+muuZoMePgsgk4pUm441C
4IqiZMEB1x+bC7IGOnqxEx1lHQiIeKUVd/mtRMJt3WapFj+Ygt6757SnHfb8NxqqaTEdmZ6bqpAQ
TZZ4dvT5xPc5TOcZXOERs3zJ04n+bgLFoJSceMD+zoVxE4GdhyUZ6ELu2aBndAWiarQhLWU7OorJ
HGDl+eeTgjbvDv2WJw1LUbb/lzRM03fTlPKD4OEgzqrLFnUmIUQ982gOzzELSzyLigfMX9Z/qN53
Ap18jRU3n0el9l9dDT0D5jPYZ8USdKSCJi0CVrS/4FndzkWXcXniBsgGH83KNNOCLj70QZxMvO2Q
myQTvpNJXwS3PAV9WX4OOepxLdnmTtcJLpfMSLZDJUoTor2pe/2i1cIPEIU53L32/AU96CiGIYTl
RxCsTgUcl+ghCJspVmOqw4QH4hIlxPT5xpmxzR0JBI03TpRLnJdsbGFsJWqpl76Z0IJviMyeVitH
IEs3sofJ2DAOvvNuJQe9ilHb/mPmEP8hgT8SjIu4jcyMl0SFzYIManc5cZfy4mf6DGPbEx24u72I
umenoCTcbKcct6wIQv097LwLQn04/Njuu+SFE6FPiuGNbYq7puZmwrhHFcC4/Z/dN5fE65J27MoT
20H/Tiwjg6X/TykBMVAxIvOdQCuZ9/pH8iFQozjA1krE3QNDk8//UfSFbqbXttmGOGpPQuG+GIMH
YLSKeQ4sJ74RGwSrgrMP6VDMsqIfRfrYtBItIDx1qwl04Ot+/SfzcfAoBpdCDFIUEsT3lSLq28up
6cj2OmcmNBpDHOapEBeufa3NpwjINoCFLCTN7OemqItPLpAHcPG14m8YNNNzLGn8P0wjWz4BOxcP
C2Zfj+fpWRyUXfcNFe3h+4P26m76tTDC8AzRjlXY9r5ZMDzBaintaSzBjNEq2WPf2M62o0TOKA1y
5W5y6E9MY6M+UL1INiKdb2Hkpmkt0uDUxlVhoU8dLnC7LR1Ec/nm0zYHaAKuj+Ym0wneHy+iuW7y
KJtK4QxqRCjrYoYPKCFoWMRZp03HRDStxglgNgXOmlaHDNBleKKFcgY/aI49q7nEKuUrsI0LZL2R
78LI1sYS12PngWnEB7kY0xbsbPk/xmFxoPNEIGAhOsb7Dx6Tfxgl9mAaDlLiuD4iRsiWpnH11Tw/
Vpc94lRdpxhiMSQ9erxKYUmojVfqbFtL376qXkivT1RrUT0A09NZb5QKuzfsrzXvpPoam1V8wOct
mfBm/SCKO0EIjts2QO9NwWCKuN1xeKVYrU1i6a2HMs6LfohxjbP963gjROgW8KZqM8a93jFQhGmm
r/Qn+SWzSFinQ+MsAsvVXDFfld8NnFXTFo1BDdyHXnidcTnOogJdDlWH9XpY3QcgQsEP8zCrrtj4
p9UG6DcgaCvGXVeir2RA/IHlWyjw+T9Lk+zmzzZMVXwV6YcHqmtgmI4+y7a1Mgorac/qgII1ggv0
VTbuLH/98ddoo2+OFssf7JTOHHnMnX6kdexnJkLOJLIfMOKNqFUlWSd3xfmULotFo++JieHa2oio
IA/IwfR5Nw5CLy8YKtb3hFsO5W29zhoajmIhQAxQzP4xcm3JOu++v6LSyPXl8izSRzMTlgyTMTzD
x1TxkFIcfhM+eFNo0BhRisWRzqfpkTkJrGpWs4tKmPwjCPQdLh7rET2o2NNMI6FTXhrns25V/xNQ
M15pzTx8ydwwMSCLo2kCEn31fo3akkAqhFL3EP4K7B35Spw7QNm9a7uA0jENQlq4DHML36qvIkbj
F+RjCLSlozG3T10XcPOWvGDLow268oNA3E9v84jAVNRV9RqzRTuk/K2rDtpxIYbXwDLxWcV6dLtT
xBsSbpIo0I+fXkRSfL6sQxEcqaQv8OH4/5c0cawFgKv/eQvbkk36Ws0Z5IvhRb11n+HsDEGGmZN5
u3bfFalnGI+jDi3G6OeZAuF5Qh7vI5qxnXnh7d0sORtzE07TPfWUQksUoVXtAA5f1aWhaJiti2Aa
4iFjcCQjCr+9DqF4NP1TWkm65Ap+fBQX7F4MPJvnwgfZG1H6wRI61N+VH87ZyyM3xoP6mufMIbKl
nCfEAI/7Z6ONSIXqd/+C3h2gditiaIoEkk5Emrz+eCE4WhfFWOV11z5r8yiCJnIvKr6qA1svigic
hYw1OJVcPvrkYVcXNqLr0gz3q5h+m7NszU4usvietChHIM0jQ3ZaIWwUy4WQTJn7SDLi9AlJ7u/o
drFyzMTuFziNTlx4GVtmMqkS9bFZKJVsTHmZuC8YwLliQJgkJD18u0tlMPdYXdt39H5nYE9GZMs2
Tx9ulArO35cswXgd9F2K7kcyXgceS9LL3eMVFAHvKmiHswfwXr7XAc82wzMYmgnD83NUQkNpPiTf
/rzFgcN7lNSTFzlCw2VRZniQZRFGxQDznbos8zvi7SY12e3eXSsB4cEdhdCTG13QVVpQr+8c5wdS
jkBZLrqSua0uVw4LrfsqpuYNxz0dP1YuuC+yUdS/2r8BKpMcujP0emXPEiSe+EidFFvELsyad4QV
b80VE+42rCoNVnAB1eNmgmpWKFwt/1OrMoXXSE+YItCXdh++02RgY0pu33Xg0SObNzsl6XYruBZC
RGX3QtfNZnbrsqMyML3eFkZln5lkZdswmoN2eph06j4frK0lSWTLANwsk49H4gl+3xgwdOSYMdpB
TroY0JCJr3m+o3qyHksQrFWnLy1i56dBePMU3XF7HSVnpsS7YktOhR/Uy+258QFleSjGIeTIWJ/n
f8A6CjSRXx/r/XJV/PxqTAF8DLOIOmu6WvtaM5Kp/ZBz2l2B0BsNkpIE4Aw/UyqxoPO3aiH4ZLhr
XS6i9Uw3Pj0PqEXfoaaGao87UDAqJuH9zXZFDeLesjT45DhcDsvrsBfwHYHg4Si2GjOVjAfvir16
NVZMwkQE8YukTBst4QExtUSD4tUAYOmLt2zdbiTkCxnTwPut9ngO+5Sxr4hM3Hj/dxxhYrGhdfmq
CzaXCo2nMShWsneyho6xcMwoR5NWXVTWezV6dbj4E0As49WoS2Q4Q0Xq/95La0eZM7NHDBVJuY/8
vRL/PJrzyezHuW4xV/ZUcUcNM0UHIoSe5A1oq1cnP/MTIU3MkOIaO30KxMocOqLzb4LVyCHTjhMt
xqPAXhlLT190Phc4Baizgg+MR8+AlnRDSwxaePbQ2aeBwJyfb+dORuEpzI1gQxaAU4x+QC1HIIvn
ioFTFCDQ1C2SGCGCltuz5I7ktRQxmYY2sbLsvzhTZOZTkQtfk8IIDjNcTBTP+9HXTq5UAg0h9O3B
MDMC17XlUZrPymcLZGI3TFrhIyCm2x5QBWWKbTFtJwnw85OKPit8D/Nki7hYifhzaWbwGBd8mR6L
Yqk9YMvqXncrkx+rlfaOEGSmINgm+ojlUbyyWgGqrxBOMsJe7BEf/zzfrFSRtX9O4so96Jzo7wUK
TbQf9Uw4gZtB8B+73NMp9qDi/KEr1BV+MYXJEFVGtbsXXdp5mYPzWWt10ALTsHhbRUsSKRHAm85g
8PIrmvnlY22PxyX1aytUlId9CJKtQfiJmWdVnc1WZP95sH36ubXHx+cQzg9AgCDsA7IiiScCr/GR
h2MMKYPY9uITrwHACZpQHNmMw2ztzJRHmXhje2iPiEJ6WTU2V/G/LodyOZlLV4zX2VQOap/jBhv2
NxF0bQTOciHzPuLeI3upHNTPvb8A7dfeuldmkS8AJJhGGIAR3hSYq1RmInxBgDeDPKgUGV4aIgCk
33DskkS7tKfACSArm5PhO1oNcWQApnyU5kya9nnYuuquFLTMOKybjE0GMFTNAFcCi+dGWgVnuW/A
lU/UqexLOjV7OslZU+iZQ5R5/Xph0viPfZi6Rda87hNMkjggT8UmUixnpKISghPOHTRplXmKuyj6
MbW3EA8hXNr4mma/IxQ3FYPY1cIIrRdJ8rgosG3fTuvjbMuCtFYLO7CSopvj+11vmaFZ4ibrNn7p
b5sBclftB3dzfb9hjHPojla2bW1C1u4CkngU9xsQOgbWI1I4DhSYjlI1y3ZPi/Z482cdUvRis40L
TpXvdH3VmlBFkjGZ2RqpY5jKiC3qK4/moAZ/oer1dWBMiR9l/UeESWWIy0J9u5G3ESE+37juQK1V
UdgOPodysGCvW8dd0xZVSnvORSp2Gp7CrJXXSSgZcFA5Vae+QEjZc8QAiGY+0fLEAdx7QcWg7B76
LRVLsDPG1UrRTx2e5xaZ/wOjY0vzRHhSysVpHQxE1Q9eZQ1tuZW3c/VLPx7divSjl1jNi2gyaRQB
QcSIJTZnn9XobTegIq/4oCgZlJik1VwqcWobAJof0wV3hICfjc5uAkbizEGiyYtJKq32hRc2pTp2
ef0m0jQVbLm8NLw3hEO7DENGbVQwl+mbnlk1+UsyGjiLPjd0c6gNjc7uGpgs3s0B5x7r6EdhjSm1
NJ5rSDIxvm4G7v2qyL5+i0Oi+RmtZ7ZcWKdY1IOi1w9oZ66DNUJaNXQymCdm9+gAH5CL/QVjf9z0
0T+SP9lOl6051AKhXuBTNSQAJKbofeWO5JUiIrqPwzlPCrOhylcLk+CPOu4fEcnc8nLGW0ZTUyJm
mTgFcO9F9j4OFiXY45Gt2xheGMQwBnMwZcVFAbx4H77T4mpILEKAm8Ynewd7inDcH3JAA+d/fwFe
F04dWFN3IpSOeWtzXo8HkM9MBW9sBm+mupW2Fq/8zMEMhL3+qEuCWienrHeWhLca/QTwptGJEswg
ifEIV4Y+yuSKeasdBbwSiXRmXwTaowitkuwbJ508xT3GXsPONCnIKA8F1CikiHY69Bz0VLF5Ve4P
w98cuq7DkSswu4YFhMDmI496EMolptqnj27ksxZFCO7uBuyeOaYyaeNpifPUAluImFOFziCfpZaE
jgbAAJcfxv3a2/S5HYK2WPlacqfO1Bug0TWsBWITPAX2DpFd2Nrg3K6VVEdEJh8QpkUmK5JWaW4/
0PCKnsEwdyx/8Qqpl45njofWDtk00uCmHSb6N+SEgFj0Cq1FTRImtUfHVzx6FbRFEQOHdtN8TlBR
PIfYks/uilwZ1XpV7CdhIv1i/n0h6B8CiFBvDGUeW+Et3IscjLhl66BiTeof0momgsDnukgea2aY
qA9NLF9SrkBkzf0FE2B6+lVPoS2NRfi5K/JmS55L7MigtreORitA4b5l8vAL+oA/nimxipuph+pS
057NBl2YvsYn/TMVjNgAtkCwUU6BEi30lxGfxLO3cRQecuInd6JIWqobx0Aip3Qgmh8+sNM7mPQ1
93WdOEG0mNzxBqG/3cCPMC24oj83H/b0r3+TzW1uLkjSGspe2BFcwS3bHvSy+HRJxhL6XT2n/jtq
Fgnp2d1Au8TubyU0NBWkYv5cuFFItFuz2EwtsDeTDvZslIkViKIESiTTfvoliYa0m3raZ30yqb4q
sVbidBZCZqEavv1tmLCkBqmqvf4yOhGBY6Sp9m6jRuWpw5bdq3ii4wPKGiJSDJjOMkDxk5MlO/14
ufw+TPMS5/sSHwoHEykFX+MQQc0DVILYuY4vbxY8jDKv0TSa3wIhggaKL639+03LpwBzTx+vMBjt
FR+TsVpmwEzwfhyZ9OU8VAqe99RzpeFgpw6DoJdXPQVTYis4TNrN8zkXSwOzBWH3xFM/yT2g5cQi
s10pwRkQRAxo/gpRMoJQxACTIr2QdPrE1u4/eBHUeIEOyphk8bx/sGKTxVciX6BuHBHdiPQRPSv8
vQrOb/o4ogo8bUsTDAFhAuIuP5AUCiCpvmakteQWlKRPjXx5aUE5Yoz0INKDX50y0YoBBCF3u2fB
MIyLFkQheOTme9SCRpU0uYQMfq0pt9+E+gHmlvKUejZ/Ed5D/qRLOvFMEXgQYaL8/JLuh8SSOw5P
E8H3r7/hYc+zILesQvH6lryZQQjAcBHyMcQSotneUdP/H+0I3GjaQk1tEUUEL4n+BZOji+ucNdM6
88McXXJi/xG1TyaW24S6NGMZL1od+7xc5NftRclpRI+JY38zR7mW+Akw0fyDNmEU+e/5xEE6LxH7
z3vuCKjfAwMJd3QmJN4I4V/BUPaTK8mxoJOqbT076p4qQ6gFKIgSa8qDFevowh8O9JbQGdZJvAju
p9VJHkFAV9XzeU3koajRIbZoqxrPWOzkp2IeM+US0Jk+FjXCcx+gehz95son4epL4tRamu9+EaFn
E0oPp/wmn03Kn6BIJ2D0Cjfw5S/2b6muMJ65qZ8aAcBHNhhbH7gBRtFsNgeRdeXWh5dl+nnYfj9a
ZLBdKQJM8M+bc3ZCkngUvdHDV0jfR0TpDnujVmiM74PzXmGNQGS1KT3baNDtOf5JNG0InyIb5RWm
C5Rv27TOdbO5cxmYA3pojqW4KCll+UFC1K2CyJphIGUje0HU6DMfhEfkkoYdj2jBnTNKrnseYLF3
S0vfcaI6J4JiOWg/RAvrW1B+p9/25G1BmsZnzhw6HNbeKQ/HN7F7fFIpQqYVUCUSORtJFyIQHw3m
YJwLXcO6MD39aryoe/q56yrXH+Kv6nrOlnMbtTkH3erUdGOX3RWTx3R85HlzUES9ZfOc/xLgZ6ma
89B/K8V2AJUA3a+HgmE9OqD5Txy0YlpqJEHIvhGfbjKyJPq5fHDTCqD1HDd28YdnomfWjqjvkjUL
XTebL9ttzFqVoUAJtzBXoLkYtEKYQXKLUGQQXJ6nI4d60TSOl68yKBEST3nV6Vr9IyunBRyGVxsa
Zh7X7JIdMCuPTltuB80X4QD/2zuKF25Bw5qMrXxc3LmB7wmg1u3Xy9+MJibNxC8i1d8nEKBbkHeU
oH0cdfuVgGbkFvRHeEFoXpxc5Ms4tRCSOF5lBi1cG+yvUGsxoNfHj1GuAvH3234LBIAtMJAxJe7L
lmqieYn22FfQIPJMLJJ5kx5+8Mw2KibuS8cJveGGrixfVo3NhYqzDuehdG6OrFj5arR2hoLDM1+R
SwJ03NVBDgTaeRWzqTIUAqmLPYmlnFQCZiNWWciZblYbdbLuP6tzK+PlHeB42hYBvC5uOK0y7iJ8
K+oJJsSSxukTv1aEjon5p///+jwM7nujjpRv1hXagjo5aOGtJTUr3FNmfMiiPR1hwayY5RC3ep7Q
s3n1YWaena5tAFqyx2iAqIicwl0jfXJaIyiOaNsPpPHwIbyBncmCDNIs1gpz4xDvl1Sp0cxKpkcO
xVoo9tkGB4X/4JXjwjPitWV9JYewygLcwbQxcI2WRZrOR/wlwZa/3uOHqCYXeq9+xpW4KZ96MzbY
3QtFDrXEck/ghsbKH00Y/6xMdBoEPodV/cLmWNDxzoDgFsDz+LTFbq67t+8KoEQfwN5DZO/3RL9s
PCIM7/orkSGR6Z+3tyjqqGbB2E/YSE+dBtI4mYIYfkEK8gya9ymojPr4n0n0rIy4HoI5+m0qtCb6
BKkcZdnrXZaRBsevEBEZ44LGC2FcE6V/sCTWUdDISOE2fgYr3Mkz8Rj/wjI18qP7EGwG5odixK5U
Xyl0xatPjcpaDaZF4TlexNKTem3mDNWEjwRvFM7/rE0SoaGNjotVTJhAUiu/+VXBLiu+nX8tvUB3
FRrUFbRGWzXnPBZqb9yHGBCZ4bt9Qhr9vjjxhPWmND8rgAF4+RazQWUStj3kHNglMcnQ0oC7Pq/6
FIka0Rm5cqh4aolPz9ZaRLlPLxkvKuGX6DnHlyAuMdz5D+TQLtK4X3pXpjLZIXsBKRtVKtUurekA
JxKTzZEw0HrxOmG/AgxhGNEmsaVdeKCBF46rML+mc3LtPwpCs5LU7rA0/U/EV3sWBfOMn1u+cO9U
pmhZlvcG/0dnJrsFmyl3C1ZpBR/qBGvkP7fTTGoiEQXakM0kXD4g/2PRI6SpGFdCXhm8Om/Txp/t
Pxe4pmATDgu2P05RqX5mUWdNeMpZUfziGBvn8J6HDN1CAaFhRIvK5IBXHxa9pPBSC8m456C+l3Pc
GuXlbLAuffd42lmLu1H+HKoMcHe5QwgAMhKZqdzac77bQZHmG27U1TSaREOPD5cn6CaZt1TbzsLH
8hKcLcdv9Efd1OykxCRmeKmiPXwkadFlTUCZ05x8YHEFSJcEOcUv4kwcaW0OSZSxPoAsbDLWTX4+
HPVSU6b5pCtHXr0O2K0Lp3lPX8KvP2OWAyYQQ13qjjvHW8COih0TAT/MUW8PsUztC91+PKJmVJEZ
H3trXDlGlceW/UV1VdOA5fKh7c8PryjZnOc73yzgBQaS1LdHaT5AcJJ6xbNzdYxWJB7i/jFrPKIv
cqxPhCEAIbkQOmoKXJAgL47CCIpUTjwUe29mBv1MXTRvlbasT18Ib3Iw440cbb2Wn49ClUHhbH2P
KfXw6BmkGSQ7q5uvR6fOej400H3gkaEg1YOi2JBiW3iPiyA+ObZPRN4ELE7CyHujzOEql2G3Zmaw
qESBh7/MiO3G6FLO1T+zpYFzqh/NAPykMwWBalAdQdBsuK7r8vRXLDXclTEf1fcjz8bo8NpUYSCy
Z5SXMFpZZaD0TNLSb2g4jWQ0in+v8mo9uyur4NQTc1cJCx7LPoctnDymI45q4xz9sqdYTkWJqLmG
26TeF/2zJwBV4hL+WsIDokzUONG//quwXs3zmmHMaUI9M8iL5nwOfRkG9SXfJGW7/84/gFj/XFOL
HrZ3M/dlmaucrRyu2suOuYL2nBajYvb+HQLQjgVtFvjLvMFgRWNQYWhn9XLmMlj/ojDfimQ7JBkU
BEybZ8PaH+siQCOIZpVlRDoN2FYdC79oNnjalsh6XjDDo/5ECPwS1vnwFozmqm+a2QXXQLUFWCgB
PDMNTd8+/wSLc3rr+xD63rhVpUygj2zSFnc8C3pxKnLgPfrTgiKzUseAnDLiKNm8Odjnf2uMetnd
SU42b/zkOaTDX17b+VIpINEd8TPjCnjR45WwgPNYCMB59jvx12ZWwTzR8kZqgDEBH/zg0wXoVULv
ln4Q22b1Ac4hgDEnchLCDRWCJXnCkGgXbiLqUoR/o/bTLMlNxnbIU9Hdq6EgMEuafvYghS8SmeRI
U598k92ABbr2CbqM2k6hi14WW27p15gErriCwQl+PwvXx+aaafKSptXpfZYsa4AoyC8S5+MulmmY
modYuHIvs7vzFfbS/J5qfsjUcZVH+NcMCNJBeaDmUPCt9BifsXIgR+/2Kg6NdfjuSyNIVVQAv9nS
rMOXqhwN3gSbzKEV94AfpbwrbosmLLOSLjQ783Obql1y7XhTXorFSJCCQkACOi9Hl/66fH1KAkgf
nDYIjZVOutyXllaBs5cGN41XDZzOZ5ZaLY8fWltIwXE6VcXKnBWyotdbxl0B1Boaf/JrQU3dZM5G
AuSbxPdohQcX5TKXhqsweu4WXiNvIdrIuzE0ohddY+jJjmju9d4a6lYx85Pk9ql3Y71Nt/vrW5qd
LtgDZipU3TivMblxt6C7VdcK6VWRapnxyW/h5UUx4F54WdUluoZHzQjSB8F9sD6MoVPtMVau7UZT
LdMvo4OXM8y9bMVPLRu8c6fHDghTsNOodqWbMQPAoK+qJ/ob/YMnfCN5so7Dfas5gwnHB3i1H3dw
k5YPaRNm839zpZaYYhBW2vilKvHao9su1aBJJqALpSiEfPaQoYwvKPpnydmyW//Akp23rcS1YbB8
JOjkLY9I8oAB3ULFIrSCqqsF7z9hM5IWCceUnx0Ks0zTEkS0TiUmb6J9g5HIupYUb/l9HLZm1sin
KP0cqOdxhH0BimecFcTNaYl+gdVrSUAAdxUkPLjreDcdw5Jh4a4hbqBLs/wkcPc17ksckFRypVuW
pJLN3BhRMlDlPOIciLvS6ho8f/PpAIWPd0NlFiD4Q2vXhRmQGspXxzsffrBxz2UIiM5SM6jeAgmI
vqvo5nEUji4ztDUPJvkPYnndsp+3kXQ96AAvl6ecUURNdffO718OOP9xiIlF8LM2T0rhiqcs4Qnv
ZqP1V+9dv6sdginp40/v2R4tmYJXUY8CfJXaFNN7nzRsw6UaDQ1aIVGId9nQB139ep9Ip2Qp/Xk2
NA9LXpa4JQfou0jp75FQwVVXp50QEsADUIXqvQuJ8L/d2A2MuWfNxS6BN/6y/n9teV+Vq+HU31nz
WtTIIgJDvr8fJrN/xwV6cyXbIZFulVjPbFF67jjvxKi7wzVDzdTuouNuyjLV4EAM9IwLU8MATgxG
2bcSEKBFKq3zBJ2rHb7LpeDN+CbILXyEqX42B1Ji17hw+5qIuu2Z1ECrQ5ij+mvdJQScPTGV5tW7
UMTRFStWghqOAwxHMSMf4N1yLi4FZjCaDEHzgvspiKU9K9nANvVeonZVuD5a6hhsbCkTGb2sbyea
yNT5j6NbWTH0h/1xNErLLAzv27V4ec16wrUN44uAf5J+fUQit6xAlzNWnU4VJJl2YCobERbZcdjL
x3co7cJaPB6RlPTAiVQkg6VVxz5evp8Zj9adj3XbTQfugCHNhmhw8WjDVlldrLqjXIsOMD+Vj8HA
GuSbY0Y5N9VAsnLeWmtLdofgXxoSyy9PhE9N4eYcQ2+D/rbFoa1o/3c3mQTrXTbaTyeKrw0s+sgx
nt2Wl3qHcDAxJTXhAlFoyr1d84GVFZ9GBhscz8WQ8xuXLTzcn5gHe43iA8qbkzC5xKwVjrYQDx5h
n7C3xwKMu2GJhMo88rsADwNUPmQT7TwghlgQ83bkb+TJApHX/DYat0cgDxdApD9+fAGQb2rEVDOx
Coqph4Nk30IH1gdzE8KAhkNGo9oauMKNYcZXgUAvrRn53XBv/EBC1we/GoF5ORt7TyOwwXnznLZA
L4/8/qio8s4P8+R9XCJ/sGPurJUfUSTDxppVaKgG7dZMt98OqdvmoGV1GLa572zNAoXxZpcm5TP6
TkL2UeG0EZQfwji/2bcZzcew3vqBHqBSzIxsRPuB/YktPvWwyzCurLc3AhjITPMhJ9ctTuiJb+xP
E0mUwqoWqF4e5O7N9Pm/Pva0Ybmw3XJd50+t+5Ori6JVov5fFDSuo8z4XCnnqfCb9Z1e0oaXGkHr
EGTKlP37yNmmsU2XzvmndPgHHxeqGQ6wF5HUVAgvXmryLruMTIJs1Cv8WIAtWJSGa38HI7Vm/yAA
2HeU+F/FBGUhhsC4YpoaXx0erXdF0jo6BxoU2JwuJP7xv5FqXwi3N48WnRwLAwDaTwM+SLNTGTLC
efnEfIbBpQ+6Pz6zIJHk/Zk//PmbdneFmMjHjyysGLEiiPWROtrhh3uK7iZ/kS3Vup/OP8K8L7Xp
Grga30S1378i1YFEyKUMT2/pC7PadsXYDc6PqmhCV90H0EQZqdn8ByWTZ5SpvBaQ3bVE7/iVAdIF
QwkIPo7JDvIX/SKMdufqZm5Tw7nEy1R7DY0zcB2sYCyN/ptfyLVdlC0aanQ9Q+gYe+tjS+dNUJ2l
s5S1ghmW0qbMdJqMvGmUSFyZEGZjyIyU4xVmKzlTnB0n9H3RpUvIXeTRb9zUaFUonSb+5dx2srMr
KPjOY0q+LVyS+3wfRSYssFQmZd4hR28oqH+GzDQvXoGpkFhaZUu2RRRqzzFHmnpZXZsMjRoMm8TH
ZVUAO5XrpcXxRWrcBHRvWOZb7/3n1oADqJotqLCtX28JE2igF2hh3EYVcxk58PP+vPA0jvrkVMct
O4qpGhY03Cq0AXw28aB/Ifiw0PO9SIYKIJzV0X8rF/jAsRu7u7eZbo9cKhGrHwrxGbuB0SqSRFTa
xXK74Ws2MEPPCP52NXiGRzQPJ0yN1NFhSPUbkZbNdnvUjzlolPZTXGLiQbLr2mQGd8cwOdl8XToW
ugbOFmeszqzfG16/Qz+qT8lq05NHjBrqUdmGZxlbQfeHQSjagD3Dy1bpcyWfKUqAewqkWfBS2D1n
m3zGwf0qdSaVx6f3OMwuXjrZDF8GXa9cuIjGdv8W+pML6rvneB3Y2IJLT1ZxZ211L++tPUD1Wj7m
5SijzEaJQ9BVLElK5AN73V6eaiRz+5qiRNVyddYYmpWgpmNslhlu1fGYNyi5WMOuoTJrvUr0e10l
WE96o0YFDnWgQfgJ60gBry+MwLOsKeEr5fJYDOYHAlfbPZTxKaaR4sGHT7+kscXstvkCbznxicDE
ZfpuGRqUgf0JPVgzWBjsIP5YlM56Uhnxsu1aFT/GED7Ie0bJdfD7cP7/PkweTKw72CJWR6996CK0
Na94Uw0U2SthveNZ1OvL//RfM10GbjHOO/UhnWukxTn5sKmAkcmaJdBkzLrOk8n95FAu5nhGYjPv
P6AT/TRR0yDUA6IWbL30KuBLlXP6GN8hzTW3c08GGdGWtAvxP+tqYawDepq8H5O94R8PjIycA7NG
NGBecoi/Nq7RRHB0+6nZZfmkZZBqoQ0jgtWUd2iNFw/nD5t4Aj+vl7UU+J82l3akccUJ9VeU+z6i
ZHpP7kDxKQGuI4OC7pOdRGYMSTQ9vqvH+aAuhjRYrIdToWmcZ+tHqnDg0C9SXUQHvyWyYInpw7T2
bEOysgS40BU4S9E2KRllJAioJZhfbyjlEu//F5PLuyuDp2K/4OSLatlJz7tXaoHYnZG4j8uqpDhI
pIqj5taVzLUrc3uS4PNltjy8ypraY5A7vSjTWS1jeeuR+XoFhI0WSYPlsYdFDnRcG/R5DYUxFeYY
oAaHztOLBbyhK1JyfV/Y6QUGJV1IBhCqSljp1EchBnhJboWyTNFCTYeLTn+FWU4yEnc7jgLedbhr
xAP3OyNT2TB82ptxUAmhben55TohMwjzwGWIJ2izHXHXRuCkseLULmQDKW+SCGw5tt657I8nvC0i
w04TbvvNWWTiZCTNusPnpJq/wRRiPLZVNRLbpQXXFhWuW0RfzDdo8OdEXS+I7ylwyA/ncNQ/7st/
l1kfm4T72JYcPGl3+rMSTk5kl+K5l6jgjrr6LwDfF/bPBViA092f7QVUp+raGcU1SnEDSwN50oIF
Rt7n8acyc6vHrxq0ezkQLW9jySvuqFBFn+dUIZVIkAh/XN/CNDyNIL0MrQ2F0jG7+8gVne6IVsSl
rBvU/gbexUlaB+JJSMX7TB1JWtGUreYZWSquJJB24GNlstPzN8csM+6ipPwt6ex4nCURpNo2xSoH
Hs31VbBGKJgp4hOO534v2YzXyshxTlk7E62owJ9B2YpWqvD3+HOARJ+aWkeouk8He8yB3CelqaKn
b0gPkDL6xuxlmUmwQK22qQiifYE2q3YrBNfPXmo7XlCnRzjxeUpsIIErEeEIkQAwMIKCISfKimvc
1NN+O2T+E5ITVppGy5e5NP9Qptvh+a7Q94MjCwgW3Av07WTtKvKU0gjJPnlGR8XGL3BFP9hE+6vh
4dtj2reD1o1WMiYg70amjRmr1uUqdgXJY44hbHHSq4c46YIGYaGEwuVDHIrDzMJu7OYZ+E8Wvck3
qvSTmp4uGzKKTJCCmlDs1CKHRS9YaF7k3QDl4i+tbg84DIgEQ3cOKAIC+DS9Bq+oz7W1Hv2xFpTF
LGPh1SZC5Agl+HbOo2cRDk2O1+nHGsKFfQtnMsKT6YZK0i8lzsTE0q/vz5UcHh25yycffAqHMWzB
bNsNjYXJ0UPobVl2Wp0VBn1rFBLknhH5a3w6OJzbABaEAa7v+B9sX4KCQiJrn3l2m5a/59CrJDrI
7nYpHa7cruL/k2UADRH7eyCUuuyrGZxdMNXNFozdCtM+lJaNq7b7EdyFizgIayYor1ee5hemPNWz
AMsvTozlm3t5Ji66A9qK2xXVgOxEcnahqGzDIJg/FZXW69Jualh5dGwIuR+Y4z/Im86qvFY5FWEm
puj2Vx1luesOXtJ2N+RdpRbf1No/ah1BCFqCEmdikZIXUwQtupNdFoH9wJEOPhDjJ3qKqNsIQbwf
tw0WBnk2naJLgUGnVJr1KTwkHF3GtiDophAkNBf2fTE8IvY0rYVmVEbMjMAc0M9j0+4U3NETBpEQ
sokdubv9i6Wj/vw4FTwyufBTptiQDUUuIEO4VPnuiC8jGqBqK47OHafSuH9OcDMDn8QD3zlhyhmY
Op8Uuw8nsBf4f0U1Jly0XiRy1IjRFsQxlnk1NWLAEafkXBCNO8k89kRduSph6psMmBzmHneiMzPa
4hGPzhyR4RL48dDPLwZqlUHmr5mmZBUx68kornrLEjN0J1qAVfD/AMk2Pw5EZLnUEFWPnBySihbP
+SeVMiZKNDwkiUtJiB2twBqZ7nZ3e1NYo3JWgJ2ZyNWgMfYAOX7m4yWgjjiQrMeCKk23GgpvZRVJ
53JnqSUfatAz2fi/AxKbGnUbyjQtRxHW0/djKKTzivgKRJnH35KjRtRn8aw06xVSP/v+itMxS7k3
Fz7e2LWHXVrJGAxTwLtxwd9bn4/xdvfr/q4BHage0UlyW7+OCRDNtHB0ANsDgLbe6h+zmEoUUiqW
b0vJ8eyl5RqIpoUWUCTROd6ml0IEcqa7OIJ49HYoE1Wa8nXI+jpDjw3qzpbsJlcypTjTaxaeMsNF
SFZlLdH9Bho2laqyotMaxDibRk6zluQdizT1PpiZUmNWyi68U0iQ35qgurHqE86HGQQOOiuyL7WD
AYQj9mLe0jBsvzKpNpPzdrkyLMbVTypivZCCWVrJLPkrWm9cTRzQ46QbGmysNcWadhnJt8CRjGbK
VmiwGbA4RPBovfmCxcieJIsjh+IKJjoDS9dLnQPKj8y6zHApzZ+MQ3F2t3gBBYqoq/UfwzZ9oi/O
QM6bQYYIzJLbXAClKkKBghOkIxCADMlauD9768/WHpghVy/VzyZoRpurTL7SytF18EEaO2CpoXl+
nZjqsZAbQyyrPB97Im4ypBuTC1gB2RqPi8YQQlZLumdNAVu2hCBLXzXj+LUQ83Z7EkpQ7zWEsOlW
uc/YEtrLvkvn9syyIak07TCO6O2j5FSW8V/RCctvaFvXZcRuUM9EXqxLDieY1GrepsLxfkr1XC5S
Pig+9uYdsmhwe368AJMXr0DKWuca4FoPvV6+/YDUD9capC88iKzSe/7aHxWsLZCb7YviYdVUcJw7
gCnnJcOZKfz6rIGX1QpOpF7Y995tYkDckG4NurN2dPH4leZ0gY6Ewu8hGGpXRCmFbpfERGEc1IJk
uKaS0MN+C3J+br56ZRGM+6DVnzLMs6ZbHFjLughPx5WqA1BLyx761hMBdwk4QtPh7fpzng89vaD4
NMKmPGIJRYz/ai2naU3lqRZ4a6xuELPPKvHRK1VKjnh2OBNH9n2a47Se8Pyop7ZJGZBYFDxW3YmG
hL3xcQXOUkXjUAMq2eRWk41b4w6cKZS8vxiZPkp4OKMDJW/BrrNAWgoh05CsFXw6S+sqVCY4KKG0
6sAiLgwJx6Fm+7B06MrL/O5ThM+yiDzwnKS9Z5W7bnBEkygXz+sGpwYrw8GxJMvbALg7oIkYuF7V
c5UkZZ7KrP0jRIWAtYWyi05NOIcAn95p+Rhpvb5Hr10WP2as0PHY0NB5pxDUIckf61DSPlp0ZT2e
J93DgCURnv7C7ls4lYyqgeiIt7B2p48HZ8IIBE/x7Wfwhm7cmZDqG8yAmSZWeurGMPfmXH/LuVIz
hSiSeO252PgoOT3r3id+jH1c6wbVtXvO0sjceDEmJtGAHT8k7CZnZRRcmIaIUTm23ebZoa1TB1Ym
UUVihBAsPRcmg0eaCbrUT4HLeibAfdZ4BJLH0+SWxzkL1dh+OKVwjRzVhHrXIWVv4N/HNRsNupyj
vfOVbC/e7ffMJczfpeGiHdGGoobZ5EHNdE5mmnoEF4rBU+0Is5GFmtJ67yFvDVBmmncMCQ2HLTcA
psnixT0UAvaEKifR/mzHAZrXQ9wc0EnMVlTOVDkYs8gEQONbbmiAVltcNf4B2ttIrPmiat/d4XUg
hHvDTGQSPLLJzU/yXflKUkOVhb7NUqi2RJlnU139aql82geDfw+WDYh9vEWzECduRewpyGiPjSF6
0K48o6Xr8j7jGAJFaXhFIYo+J8qk/lk63rnAOdnxdau+1Zqx42O357PQKprvR4CvGFCPSTT/soVa
4nCpeApGubtSEgkJ3j8QYWvKpnOMg39t9PULcl3PUJ1T7ZxBVFTobxgZJdFFYhByTHfRSnwFBLMt
FTeEYLWLXKPK66YsiHtSO4aG8+aM1+9g0bjeFbBzU8uaSv0QuunknagJ3b1yliUxPSsdXi7ESWjI
rODBDMLCXmXqYhRHcnvfac+eRUoG2vLmJN+7GkEjg09fUdD+/BsdB/Aps/HCpi+VgauYjP2ZGCWV
DpeP0RzuZde/sEpzvi4PC+gPty3K7KqUqRavNEuYXw10zrikwEZKZ+dNrTJ/0JJywC2CCF+yrHEs
RGmvvWFKa+ZrzC4E9YzOs/R013ZjX6YgUmxkyl11pO+6e6mxzGVFQQwovnog5gn7s7hLy3FYCRfg
8wcEIKsPf+958CtqpmI8SoqSpL6BY787LOp1nbrn2t/UAMIUxm7tc9zmQubRXcSW1eJbYIsPQqV0
8RpbYBCWPBMUGnwErEHOmyUXIjPWB8UiIw2kLCr1IAmg9pgw8FepUSTI0aAQYLqUi/2fYQeAWZRs
DNpSaRluYZXQrtbtnd20SrRB2jTz27Rg5lvs0PXM7FWwwtSelLyUYfSTmtTDOQ7fmolUwvnBpghx
8oiBXGmWA/13nU1/XUekgn31Qhs3sCcTh4QQQkALLozq0BhufOhlHCWoQYeIj6oQwsZhNQVtXzJE
/Cid0FdFxVbOJFwmd9nrYvnIjLHl4WwRubniMrzWYvfBXev1emijv16Iq5a2avRp5acoMDo2Oy9V
IThzSP+1p3+VqyP1xAWY6ezv5IvEbm6dTdnosrQKHVqOHaDctOk6/omgyqAvkcTHUm3dEDOGEja9
WCjEOVVjK/sovllbcZ0mKRVg3RUwxikrkKByAEFkmmnVHgWppKAJlJ9CQJ7XdcWCZq5+XDP+PBVE
9JuaK2VezbkTJwn+0nBnAuAkUTxIXg+tji9R7bD/MkzukyViZmaG3HrUXmb5wz52stjW7Lilkosu
LyTKfT4sQEG9knnOy8O48tQjMuXQ8y8TMGgwJmm+zDjuNIDwaUBf1Vhe2bfaeyJKAYYWyI4iIaIm
DZsBRljbl/2XquVdVFiAN5akrNNPduDJY0kyqGq5s8muw/eGHcfYViPXgogOK4Ggg9+R7OGRNDPH
s9FOk8iF5M/IvnkeZi6qPx3heKDBLa4FwbVUKJHCA3ewdgylHKHdOW+KI+Fc9MVGlnXzS8eXlGW/
ahtOtoV22JGQlkFyg9o/dFPCoHz9J9WZVPOVEYScdfL2Jr/fD6F0w63D/wxmjoIPMBiY+3zGAgHW
a7envO/HW2cym2GYNGA01CvXMjAMK4cSWwD+9tHsk8ZUgaZPlJe5Dcz2jJmsKJD9uLGshtWoijqM
4O29e16TqsECMIR6LIYIIBk0BLOwyY68QWkOp3RvMGXa7QRvgST191YRogPTHpcyU4rBYe2qIxP7
i2uC4O6q9sJR35JcvdyYREKdlTAXYoxv0FP3QnmVMPzkkol9d82uGmUzSYd4YZCq5IUbaLjNXZ+N
lVhWf/i64U6iOWWDnl4Yvbuv5G3S91vj7fT2ZtVg/g3iKx2FRPNx76Oy2p+L70pbEEeLQi7y7sq2
gZ4qCXAhM60oFwr0R6HL15ddxWdx572TyqZsIhupr5qgq0XoMrl+hoPNrgEW9fSCoScS+YJF2hOk
Eow4cF8brDfLlp6rk2l1XNsGkNBg0hB6s2hlUENJlD09HAxAoIcZd8mZHEgJ59qLdlDHQguJwW5P
JZ+Ny7PWzhfygh1Cn27QikZYQKGzhhk6tg/a5D6YJjcEiomqgEXhtmun1ePhSwtJCUrOKXs84s3l
25BT3lJM9XIL4UzaEcz1JEZiwz1+z2Fi3qjGpebFyioKtHMI41cq12YDLjqpCSJzqlgx/9dLGSBG
qB+VCphSy/Wot/lI2yhpprhxSdGRWwOwYVlMk64G6NK7aTvhbsg6laoZBXSDhgEw7/AMrv3V+66U
x3hGqkL/LqFVYRCKfzat4Jszk0dwcLbq8zOfUXJrv2ky06Oq5y+9XFsc1/m3lH4qaK3FrGzoC0io
7MgVnVkTE2SWXG84BFbiMcAoQOyu4PyEHxBJp5mWUH5gLWXWouozPBU8dHNAnCt07m4Hyg3ePN/0
pJxBO9tVXiMBZt4sD7GMD1qbByRx62Jex3/k7XaQrl87SFUtXTj7Fy4l3lSTosvpU5miQxA+m298
62oVrGEBsg0cOpnXLGcAwOwbcw/KA+fizi3AEh16phwlvvo5Hb/sGmyU8YzJVf3u7zg+CeO2HJ6b
vNGDqvsV86P8N8YM/XDoDPAwzb3KTIF3fYgPk3F+QymqyAOfn9+G2DPcUe/Uc2LWrhsa45pAAEK9
kxGwIGQ14JHUZq+kws405G28nV5qNHlQliof+iS5y/AK2bV4E80O1eAMQgNQnrpoL4628bNlN/+O
mrsdC/4+udHuUdH9OewF4jZg4sLiGrR/gPzK+RZ/iyGh54qwkEzJnh5bIshxPDW1DNzq/BGn5hEG
PrHO1Wj5I5Oiw+ksTgEE5MlvAjYoXQePgLLejHvz3bGihMbHZC4ouCD1bVi9ffaixziZCVkrzgra
rs5vqTkDfY3G37nM1tcFPtNY9q5TvAcWJY4XbuoPjZGxNy+DLyfwMHCk/5D6TrZtpS5ggdR3xfsS
fx4Myr0wvTI5ajLa460LgkZbMsk2m7VfHkXw/bfDbQi2sSxgnlDl60LyRGCgwShC28VChr67OEYh
j6dj3caRMaFNE5n5QtcNXMulTRuNS6gTPfrIZPf/GTHx59wncv+k2/67gM8WTdZuqbiE/gu7oyJ6
rl4Aqc+xiHE6V3RR6DGtcifOfHavFIOixxKORISlIBVLHaxb6mGy4dIMUgyYq4ZaRgBvaRjBLRe/
VvdXyJ6n/Ow02RrM4VLJAus0FqD+TpHY6eaVAakcugGpxKFYq3zdjZC4fcibI+tLFgBc5+7Nwt6L
LUEA/yqz4Hr3HVuI9lRQuoUa5P7tnlI3AOfPKsSsQ+uIxt5/+UQPmzhavO9t37Fz9ysXkRtZIKij
zDulUHJLGq+/xxPPTYi0j7G7fqzCd8xl+RDu9PzAy9VBZ1reLWCUTV90woUXBJ3rCH849I4VB1y5
yWV36Od1dR6jkzANA1G2S339Tv+Z/IJDNKkChYpzNMWvVjOKURCLKOiJEMzLoSemnKyFG/nYJorw
7KTUqs7JjehtFfYf4F/SZmzMhOLmPj9bcRcjjjezI6j8oZhxsOfJMXPDHzSy9XQZu6omuhsBEJzQ
WSqUrqwT2BpCUVGnsa67MfB1snO2YZ2aelH/De9uLWscEqna4ZaRLLynEizu6QUd8mte6Rs16bKc
j4I8zO1YiW9hjkc+PL1YHvAw1/yOg9P5y/wQCSLPYrTX9F03eFCY7Gb+/4YNjFNFUx9xMC+CAM4V
E1YDQP6DHxvyIj/HKm1+BwffKRA9CS8/6AncktrJG34lfTc7cH475f68hQkpcEWpD0jQX3uTkWIo
5UJDUxH15xYuzeOw3Ns3/IlP5hxMNex4CBm3nlV+cXfDN8UN989nuTpWKUzRX0TK58oFldE9md5p
9LPGdtPu0t2msMehBKsDmOGs0SGe0JwuEx+9gevX/j8AWJNM8+HYHfqThpjszI+TcrDj+QYPvZDe
99d70YXyAL8cuplSdmzW/TDehqaqZKRLCrXKWgZz8braPC6P/0hjH3tvqo08Jw4UR5miToPdUSLQ
CkTTnp3XDdiOJe6sJUEUQHJmTSXP/iev2uolV3oDEkcdASYDLQcf6f7zjmF4/ljT73+Hc2z+yaxn
l4P5EdAQfYfhwuCtbYiu6U36yUtcgRRisJkNhnwflAk00Ze60UVHb9+kwhRGFpHFYYUSU57fLkt0
YwF4yKd2l5VvdETpePhJzZ8m2wU9BZe3l9AUORtEIXNAF1zgWfVxxKMul2WQElFVJsil9Z9d4qBJ
8IxFkcxVDLiGPmeE+IjeKBqBmFbfJwOMj9RNi7dl+PvsIH8+RjzYtE6NXsScoh391nKgjYWCmaI/
8LRHtK9CkSRx8qVcOEfkNjifeD2RF6QL6TNgl/BBRnYMv5SKL//qxsHORGXorMWusXwLcxhUjVe0
ytcFy1vnVQ3OlmWXu1GwebIZGtNaiL+SZWsN2V08i8fLIRvyKZ6+hF0zbaLkOp/xg64VHNfhedAs
vPdtO1aAnNMyky9DZMhb2E5bLTzqI/3B2SpTkr9yvxdWQnVFas5xG2/6NF30aFY0hUH0m8StY9Cq
8h0tp1EgzaeUEx/vRwV2Psf5k8dV0KjNfmAtPVHhkfCyJ4g0FysyjCvdUfnmRkfu72QMUMtPN5Hc
YbLEZlNRewvtqD6ze75cza/eyXY0vtpi38TXFuiuzi1MLLiiQ5cdB0vBC1QSovG89pi4nqRNpQ/S
Ce984b0YlC+lHT+hucgTVhCqsY2JncK4tOt/Ai53WRV1N2Wgn6oTIuiIjbW96c1AWdc55ZhS/BRB
gFteUaxpNv2ddh7HTD/RqSuWSI3Tfoux/1NQ0dLE+/DDVNy2/kzGQ71+lxm4f7i2YWE7tEzeMZLn
9Wv7HMgla0aCExslo32MeZU6KOHI1+nIV8KaZfpYN6O2M2Ow6I7jN9TQJRU3jigeGIShe/oDUX9m
S/zMD0Cp3IwtIU/dU6TkaN3682e3wwMgkcscdRK/7SR8kD+wWSZtzbSTLtZnc3ICpYbwUHc4iq/Z
9Y21SjZPi7qDFiaItrqb2t776ix/JDKEMu5J05GARSfdXZ/joAmlLKwUs1yUnse2/hrCEkPNHuwb
Keo7cu75yg7P33MU7w5gnCz1NwgA/MJuOJjGdjXuiCcC6XLe87WHCi6nIQS+n9ZY2AEoUgtDyk6m
rhHLrI/1tQRqq469whFlzL1wFndERJLbkaVTy0HFBbK6YvZ07vTBBNPwEgO3lfdqMv7TlC3jZWjz
8knNUDAfJ+dXBujkOhL2lCJwfa9aKeg9kilxh/ACgTkSFoRTulOT0oOoSB7xEmMa7l00+VE/AR/9
/dFMoaTx4Slp8iFH04Y6/DVyEaTsVdXOe7OA2RXa/qLG17A2nXr19RZiLP+NN6PXDiSG7WsPNWZ3
gx360Id9S4FqJ7Rr7goXIzfqhMRZviIJl5G+IO21KjHf8djg+Jo98urHiawVXvp0401gYnOCrySS
43TGfRXO1dqruBj+R2h4TdNxkl9Ot6XFfx71ELwAyAUOSLvCvoSjaQrIb1+1KhYK+pKCn0VoG+Q2
9GL+M2AbhL2cVA6rca4wX90AkiSGos3hbJe1cgIIHYztY/b3m4Be8mf4CM5py1MnfMSLuns9flLL
Vj4tWEGLP/t7T/TVFuhUb8H9qq92h1yQHN0ZGP4xwCembMDjrig9bnqHHBzi26uxC68tAottlSMa
5RgDV3fMRY4f3XD4ds3BvXBawalMq6I7gc03gSVNdDLJd78cQHHPFColuAbtdhcjSRHFJcv37ect
a/W8fzqeBLu2o4H6w/y5uMhfT23gU9zuXqB3a1liKtNeiAbfyU2Eeg8JTSP8UPXXpRBhROp+P4nM
wEyfyZN82thvCV6bq/rL4wqnkZrxp2vOtHnSgzcB9XFfn5AeTIgALF40F+hQ63N/0a2DbXpoYbOc
OSQgmqTFihPlQdSumUbT29LKx3V96tx1C5lDiCAbz4WfTdX2tluK7qb2cHquv+PguL4WrQH8MnBv
owSQDpDt3Mbsgr2nyETAOZQOVr0s2BNclLYC6osr9g276d2PMBzi2T2VLFKnQLmeYmtIXP0334H+
Lf6uHdJ8D8FnpfjXjyT2hqZkJPfvRk81Dkag650C8sBgMP/46Wv6rbQFkcv5CaAmNlwfebhnzmpe
ws/193Z0mjJXbensrrFsXYNMISl4jTU7aK0CuHpAntyLCRpbh97nwRiNoGKY80pherv2AKoyythO
W1HizY5l+mSiCXyrrLWZsn602z3QIz4FZM8cWnQe3/vjEOSqrBQk8gWjvMGR5iyArByyMCLTn6dw
JB8OGpG9s9QnbLPRxRbWRMSKaA7MeZA0FVP5FE/1GKI7OE6NxnbWhp1okQqGe3b2W/w1YQYk64Vj
BYhEBE1z0olEsEOcBmpL+EBunwnGQGA+q32VN2TXNqMCdF+owOIlfWYruQt0PsfUWB/mEjS77WrS
m2lQhY+NDCTuLOUsM7MY8mkI9oL5Ji7l0vv7hTaPsuZ8WxJTMkHpGIvmzn5W2RjRkTp1zG4b8mMp
eooWYrqO4DrRDjAgBlkaLWh17rFNqdxwbShd4W575mOVz/2JqjCMOrGQDwv6Ff+D71lZIdy47JmX
hydtjKz0UB47pgF7F5qIqq9ivlUMtQVDqbi4IcBT/B7XWWkdUJrCZFrDoFidqCrXtfMsfYfOzyt+
T4Jo3WrWc7RHmoxJGb+P32CpatMecSgmNqTvWEpDKFBmC4jurVe1wKNdpNs58nNYJFt0c7FH1Ka1
Xm5z3nOpItISgVmeGL767IzxSsn49qSNtAhFJI2Og9ynJlW77bVqsfPeFeHEgAGV9WajpUUqibE7
AJdLzeAwiJ+FQdZF2KdYsZYyRvXnlnYzJqSr3t3gKflFSGZShKRfKVgbrwl9WzVSSq/z2tUY3hXN
WFa8mcHLAUU9w59rU8GYEVkZRdGedn9M3mbxDm+VHJk1NvF75hMAngwswx+Aunt8FXkd5Yp9GfyL
wELDmwKQeQA7xVlhmtVxJ/pLXtIeolY0NbOQvLp6ddTG1e77hlKrN2c9C//UmH92xRuRhJ2OTy3R
gjznqlZQg8X5lyvtZzCMRoQR/lhxMal0YjUfZMFR2289a8aPhLiEVu2jQOJJ+yxF1kDGyi12lqDq
NcLvp10GW5Th3gquVMmNAEkfVZhUax6HNGB0CwnzktfV/gk4BmK5XbPb292TzyjcevpqEjZte++f
ljHNZQ+OhtjToXbEqnvX1N2dHS2p2fDqmBHpsf/Um/Ql3NQvNK9WiFBOcAtW3WCt23S5VNxUee2B
XA+VcauC+yGJUNsExe6ow91PMN2m0MI4T3l2CkL1eR2XzK+6SONhfVg9YLJw29YS9Y7Ws4v9gTe/
XrKmx/MfcpAOVVQHmS/+cqWntyUYl0jXpIhAShyNIYYtAfanw0uRmibK4NgkaHZbVTqWKX1EkHNR
sRKzERf5h5CVS8LM0FiWEzHCml9GSkWA3rtB6QJ64cIovsGMHvxyeJbKqnc3iD1Jr653rmx/NP9+
PNyzpQRJk7ydrC6ynWuRBnlIMICW4+yTGEqcy+aCVPdqsHeuYYYpy6ZFytcDQU4p5cgj2IWVuLLM
DT3aLjR+BkaJMEUGgFHeWHV0lgi9YozyIYmCfE4VVV3KHcNrdjojbaEuVKtvkYn3MEAQaoJtFdX6
Zkw/UQI+MCc8tAmo0QhL/jJnrPPXFwJBt+DsfrxsdARsUAxfM8gvpRZMXs3XtZlvqClXQu00I6wu
Xi3+4oyPzBIm9guZsAj98ILWQTCLeIYyIqSjj1T3IBZZEKeq1xdfTIQzHIIeqoyDhEHTc98VOANu
ftwpL5zQM1NsuaHHnHxrWkCbkfifQ2af7WFKz+u05KmkSDW569AI+QbUt+w52youoxwa6Vynf5IB
s682EfNnmWtWxCrss49ji19bWYskKlPSNaHWQ7tjs7KtVi4IXsNou0J7pItPIT1AkDJASPvjAN8j
leMjpPTJ0GjZV465Z7GKL+n9lZodd+TwE0JFSCcoeIU7ae/SiF96vVpwe41nmOuF73lu7YRsuYt3
JIBi4MFuAbx36y1/Z6xunazUS6iwZ0ePyUPhN+4Aqp07VumGVDvJhbWT30vT/8Wp2+pOS+hE2Vpp
f2JRub5Px8VEt0bm3iiD661pMLq8Fy5OQnhbg4RYXwWBi777NChx81UpaoLDZsf1WI8hx4ZQjVEy
V1FrDNshxRQj28A9dnETR47f68j57QoTT73dKwfU5i5fPRHJxLYy3EQ7gD7lvwWR7nDEds+N0fKo
DHATT3iVjgU/q1iEFpF+BsaIlqDHa+d3yLlZkh8J+yoTrU7REB83I9EMHT5rBXq8El3J6ruLXys0
Ofk9RUtjqjIoXfatOXFFX7rvn5cBSxueQaV1Sgm/+LMIzTphTIDiz3OUkefjEq4ZZK2rk08GA8Iy
JzRDxsa6SYjwCfs1htAIgdh1+/7gjlMvc4kzaoCc+ZS7cu707kS/sfQa3mbIqiJKBjQXJ3/Y0NCx
tHGs1g2TR0mWVanisMH4l7PGKAaMKIeBQnBa4is17wbDY8Wqgmban3ZnokmhBTRmT1v6JhuEuobC
xSvPt0KGQrtGvQ/q1PSnUX44SD+yng0kYatmZBnyJBqccvETbKg7fPFXyrkQUraEH4NILS8V0uHC
6cJx+pITPJWjY0DKz1oAxU2CHH7qNRjffRpGgdR8J7lfYfS9tbQiHVfh82GrUQA/DMUVZz0YKTE+
6qs64D/1ealozObU+eJAIwJSoLiJ29Oesl3MRC4vYJOE4RJjupJ6iYSuF52Qe/A9FaL/JjEd1o23
r1nnZl0BOUuTzrx4baDtZr8+z7K/9NEqpC68EPcUDkP76LFxvhNs6/h6hnMp5GjL9Uz2lSAnbaeS
QocIyc6SIFywcGJhoJO6AsxAtXYy3ecwXGJk5e/u97Y5GzaBExxIvKUmCZ32SBepgncMr+XquM25
5RqD+8LoRvuemEBGBLzNu36muvWfeNhofgdy0h4Bw0HElLSSXaqDhK0Y6Pf41y9q3mv9lRpYq6yZ
KElQG4Tp3er+V02NdrCYOffjDf5OCExP4TNbyq+pmdOO6c0QPBR1iZbhkVK+fVmN7UphTYxh8HDB
KhRPFlqmp5t/Jezbp9N0W8h3rB2xT8I0n8VZylJ8HfnHd49PSVr/V7IQsDDp8plBzBPyt5UoIsaA
o9CSgSUGWaJIG4mlLqLahOeJuwfmeTh0PL5fUHZkzJklB1tBweUIgSj6z1M/OO31xkaDEFnFxzbe
QqzlWG2DKD2QnzNHdy5yy8hAOJ+FmxP4k39+e4pOR7wAO0GZKec2JxusIp/eSdcvWUDKeMVHKYBK
8mmuaUqUwANGE75JtcdkRndiU5pyIHB/ucJnmNPxm2VkqOlc63TgTHlulX2In4vUWMwreWPf7L4k
iZ49ChlqYipEL6sPQqoEZCLcGvPMKa4TC82XsN7e3lgf1Ktans0DZuhqbD4dwH/E9yS4yo1d4stz
uERc5ePoaqskJL1vwiy6YvgZFNslwaPDbivNAe1w7hfnA6uIiDssbm9SDg6W/jUWyZUAxug3XvAl
JW5VA4I8/ngIFfX5gO3WXUSDGLelnLlak3aAiplK3FS3552T/wnVhW9zo2i8MHfAnHVcFVpqZpnU
lTmhI+pGHvc2ZtFntciZnjQYa846vjr2C4CKYov1ZXnKjSfhF8G6JwbcAjBK0dEqEx3MNFEhhhjy
1nJVrOx/vtYMXaS5rkf+dkcEhDB9TX6Heybck2aoQZfH4ZthA358jiWLb/DovpGTuIHOK3v1P6nj
nXLoaRVHVTlprOQfagNcKv68Z/cL/OUyYE/6nH4okIuBoxgzo1IcAOVn9u7j6OXCcahQukhibKv7
0tH++87VhJaEtUfzY0YfCACGrhXTgP2B6qvhkMYbxuz8a7Xg+Ty1IeKcBjeJBOSdx9NuSxx1DmUK
H9uOULywri30NYLcY3VTOl5S5WwKwxw+6jizVo5Xq7JWfpVD0p9OWdnZzzwPheJ0WcU6+ceecQD0
a9pR4FglehijLTJx5F+ezUpDS3noHqTR1L8O1CdLAu1rZ7qErRqrJfTpEX//wbIFKdTy43QuELYy
BSDsqWENLYv/Mq9pwrwh0czZ7Ylwrws2yzI+8V6n6aVVYVoBkgjwLdc+7hIN0V74Bm09wZ5k5Ayv
UqZtKFw2R+KrfrpZTBdoXq8L78b6A7u7gw0vh0ju+Z7S47yscX2dFdhw7PqHgdplbsDhKLJDSiy6
q0av84Ffdvh9Y3J8ZL9JUTaK9IBbZJ0FMgSRhTcC8hdpykaj6JGTXXcoLARdx40iW0K4BOWMGrS0
PmN58L/lzfaMXY5bbMe2+k9ynzA44fn2C2I5QSLxUInjePh0JWYUVZMQ2wKgaiNIePzusXd14OCf
bLof82aou0sZqBJXqppgTczHWDi14GYJd14NnufV55e3kjZr1mb4gHoAje6ztZ715WblX8JSEVgK
wK0YQRSQ9dExxhFrhtfxEQOyLv1dAMQY3qY3taDDVds084e1jrZGzWIjgdDKX5+v9EsVlvpTXVBD
vwgYdNKhnUwMEq/iu483g+fr4b1ia7Qjgwxj5SJ4HUELfAo5txCqi4NxGROKoDg9LpdMQE2ubOxO
B4r7bjGkWjfD0UfbuyA6DRFT0U4AUNUZwtwcE3uIpvdgf6ThxPnizhR9F6Ub+GqKLKiNc5KSK43G
+8l2sCSW+OvNT/nEPvzYJOBfPfyaHOpf2dAc3veaufci26iO5vSkOkwDzBpsh3Rg6PVS8Bc9OXri
onoK0tpp1Uejegn7RFWzjl3uyhdRCkOkZVAJ4PwwrWiSchpMD1ewwijn0us/i0jXlFIsP1HV9d6P
KxyzDhUf3TMc4b41XREYJDbXdX6WxvbFIPZ5zD57uYNnA4YQv3AX0O4Iw8Iu0OP+1wFpbcOSxZK8
LL7v/4d3UbtrrfxTYafQn+RUFHFwyjlCOgKTzslSyiRr3UreX5J2CA/R4MVTsHaPVFTYkrx25xay
8Y3C1qpDK3NaYqsU7jucBafKaIftWikma4dQoHXs5sXcdqPgY65dn6KIxJH9/yiJXbGi2pCpeL1d
Y6+CwoUTHP/cmFxr72B0E9x7dCpIYfjU1xysO0GHnzTmNdTo29bybo1UnavW90ihBd3EHSctEIdZ
SyiAA+MJdY1/5CEF1cxpxebCCYoHoGJsVeJxOiB3qvRpCPFMonUxf8xr/oAdLba0FghjJXIRZNLa
NWbQOUDUI8R43JEVxBtxx9Ym3LoFr+Qwp6HTlPUokY9IaZhAsLAqXzYldnMofwSDllKMMFlYiwqJ
Muiu9iNJJltF6+NhHt9MGGOmScTmdkjNoy1EYQjpszkVIUUlPnMxLuV+AQ+IGEJ5zJ3cpUXW+kKl
XrxvwnTZkQf1A8Ci2vq+i84DBkaGhSpkfeIL38R/purr+fKjgg6tXPz49OTuE8UgOeW0jPAPE5EP
XCtl//rRZPEHsFGWC7KpLRCY4lqudsrd+TohmqrzoEynUMiSC4O7LpWY0gIZ4e605LDOaTKb8zSd
cZpPvsKsYUQ/snaGNfgvCHMahFUXKrgfC/h9onW+aGJcjio9kR5clNe55D1tEpqla8wKZlPoClU1
YYypThDXLcRUnd7bIZwONBAJWmCfih5h3Ovkk+urjiNRFo/5924FPg7+mVqFHnkVwxm89eolCirJ
LycPubR0HNY6f8jCemOQl8HFQCEVR3HilE+DZCJGg4WxJ92xxBOo6tSlGteGJv9PWr262yB81qE2
eaK1gIczGKCdEhq1dMM+6ilCAanOYLNHS6tnyzmuBLc7z+d1phmjYv0BrD6whQdkscbYZSdydkf0
Qs7CbJkwHggsuA9pahG++CTgIojXkd+MBcGF5w4zvGNPz/+dd6oMcRYLVZZgNECEsxJwOgSZpkbp
Cna9YN8+xLQYyVN5elnv8+7aZDnK/EN1VK3je0aKHMNAGRXgAlXFCcwkxB4ZLZRPX51SZ24WWjqx
piHr/kVrojEh/NHpQzb9eQqQS1WhQlDxRm8JVSk0qACR+qPzC4Mm+hSHfeCQ9BDYVjDIvFW79krS
ob6/S3kFe/D6DZPdVoqI4x7L92MLBPOTlXdPIeSPsuMMjV8pb8y0vnXZsxhBJFhk1GDS1L1dMFhJ
qBdhQKeowvzyQ1mIgZ6BBsm+qAKwZJRMwvYwxSfrg0yugp2RbVJgIdwxd/sv0Spv5hoG5qok9HRo
K17Xvz+8cywiw2Y6HbfThj5eJ7gTC2WZ6C1WRAXX+TH2SvhaU7UilqCofkIHJxH44w1Ow0iwOZYl
3JOuNcQqn+2GAVyHnFDTv5b/Lfyy9VXhZVx0uJK7ZZ9JvTOX8f9/Ggf/KMI7UVI21pw8YuA2v4s/
qJIRKwZ+dwrITwf+ZV/hJreFO1zK9UEF2UYUmLsnMdzFTGf3cTGKtAgRN1PUK7hNUGoN1nveqXGK
YY5Nja7fi7aJrQWpULk1YVT1EIVk9wGP9k1kJvALCs8adJNRw+9lFiZh7H+HBYtV57iOorUeGSWo
1fJr/KNkTXQbK2Rebt+Qqni9NrDk1cF20espp7F3+L6tslG1oyw2+TKRqncVfemakS9vnRw56w79
D8oX5om3zAZ3/MlzVJ7v5vIGfSa4N6f2C8l4yREDmSk12cUNzIwCL1GUZhy7LDv+nkLM8WWoXcGS
UqeWlzeAGhX8zSX754jJgreL3Y2mDVzy0R/nUp6JNeJW+YlJv2KfFHQFaf+TFCj3gvySljXNbcJ0
YfUOk0Kbtkrmw7u0gNck3DBQID7Ic6i+gHfAwfPT1y9Dx7eMsaHHj8fP4EnoI4kYmzbJ6Z5OMoWD
4a7YvGYaV8g+TL2p/2d3ec0VHNwB8zl2dcGGzGNrA3Gp8rlqAWXDQ3zAATsYkdlbDufYjy7lm4av
/ukUTCWCwqiB67T7wzffcwTdnksIXFENxCBdZ0PZlhGgGmeRhtN0mMZn4hcyq8Nl1SNg84ckYPz6
CmFR2QtLCfXNJsV4xlJ4HtbH5SGEGVZIlGuRLV77E33ZRb8yrgqfWKiMkc+d7kKBT7G7p6lEMnH6
2ZxsglyPwfodEWaa0GUqaAtlfqb9t4+sUUk9F+WSd0NM9O9OfYbigvsQDnlfweS/z1PHb0+e8Ym1
EBWxaBTue/04AVGghjY8yW2RkMqjYG7H7z7WQYiMOsUyXfFgKn5NdLZwlJt+NevxRivHtp7+4h3k
Qcg+ZOGQW5Jvll6kkx8hVAXclNIsLnYomd8Y5jKJfTOkQeHnDjpGqKISGCwd1PRuBykEFzuVvR0Y
zlOkCyvfGiuFu2GQisSj0pl0xWSrRgGRELnamo3mNHBA4+PKW6EObfzsxFKn+CdZYHqCLWnW1tjO
6+vAOGo/WFb0vnx8jtiyHewqq5QpWzFIJnuFZL9Ul7czqzHigNdU/NSEIWX5NfayMUVcd8XtcTnG
9u0T0UXbo0xyx8H588AbsP71Wm6zYXq4Hv84CTS5NSjqDnfp9sJLySGTArhsNSzGfFYLn6vsrQPq
NeTW7cew2ao3Roa1G0wgwKeKxDzv9qB45+PMdKc7f8AkNmBuNzkBpVYtk4o9HA85BWZxKSUfipql
tJjMZXCQEtyqUfSVBdmoHBbpwoDt6TzlaQBBphs5zdUmcDrVvQM+TZSFhLjk/3DbQg3jZwftTJnP
ErAgEEMG+KeV92jRgWWqS00K5dglZBxv6G5MzdWO8SVzGCZ+Qd4kcs3tqLgDF81RQj7xhFLjMY09
jkfKLoOu1evl9/lLY5ddzaXR311j7OTULiBptt2Lp2mjwGzDgGWkA9GfQfDrAH9BrAxAPHtcbIRi
RAFI8ZYabzLfTCXf6e4ZTI1kdssqZYFGzGAc0qUXtATfhL/WdUsnYhE51tWlm70hQoT/V9cx1f+K
Pi4xt5XlXI3Dne85EnNFTofc3mLOvdDkd9J8gsZnVRP9D2X+wr3RPbAdKNS+zKmIEQBmVqzDzlVJ
NxUgeYfuUgioELICBigHNm0j90nDJoBefY5QGR9h6err/UehKGj3NK4xmySn20t6eghaDMXTt59O
eTNQxIwSiTd+/Sn1FONRiq4nKMN8iv1ZSsIOLI4nfKmWqwOFxtfVZkhUl2O4rXXs2sgXlajd2VQp
4lqLSHVT+LjiM8n0tEFsWYBh9qwfzJIJNQ1bPm6hCIrbMqvAUUz27j/79QR5bLRuO1HclvNTGGVy
EMJNwfV1wNyus4izT6TyeeVKQaKXhZwDtc+WqXscUI6ayryPbZK78SuN0T7RIDXM6D+s9ro8tEiN
7sAWyNfA6kxl7lP+Ufs+jfxDfzyaumkaqiFGLaNG8o2yE/PyS+/BIzgltSL3HXlCVI2BAUn/3i2z
a0Gn3kCg2wTx2hAaAqemixlgwFojAODisPTDgEg8uCTba5FpXiZXrw21gxHLGrPZqG3BHdKO1cij
gPJFLHyxFWcMtIRx8djEc67c8JGRxtzdIkYIuB42v1WPUAHO2v99or9aXBab1G2NUHzJslU5YuIg
l1SLHz7zSJ2ZIzRh4qmGO11VMM2xalkiEKzPLR51eUvLwivm+iH7HRD4jOyfPxoDo0dCciWpG1EF
pkHUavtbwfdSMaFWi2pqrTWsgEqBZ0ah6NalFDyoyMNxtigELQ9iJ1cieK/uqg7KmBVEKzH2y2Wp
K3gBJZw1pFPFRpnOxJ5q/PCowqOUVj9SJeF0KG0CrncV6NTocFUJqVf6FPNqp0ISaaIspVRKnx66
i+qJcycj7V/6h3luIz3PKfKt8nMR2dxCazbqA0GlJgw/3xj1c3+eAhH3SZWA9FSsLaOKMyOOd/aH
qAoKp/sLCI6zsrBbNbYaY/PZ2/cpakvkPPNofWgJkznTatNcSU+b/XOlTPMGqa0eHj8Rj3VVCVXT
zEcl9L0YEDW7XgT3NuG9kEQIiPVisDMc9CQsScJ6MzBN1ovra8Yf85PWhevU93V4UsQ+z8lPey19
IQJe3jaqHgyZmDg8iKIg+978M891rtXw0t8tkkHRNVMs1mn83iltFZTtuMHx3Ui+6+FlxtidDxZn
D3OhC8j00UezeBdPsDzxzJap8FYHebYKDWQvHzWNUZGyIP9SFZBTd3eh97uyarXHxp0kiDteYlF/
i5ptCQBl0IfYzEniqAc3fsxg2C4CcT+oswKU4bei8hP55AXkeJ2/jx0wcvkHtPT52yZtp3tNVh5C
1Ekkw3f9dLDfFSfNqs/cTWTXWZOX3n4mXc2+YxEeHRTh4s8ZJrZwi03KH8wO7oya+XECQWfI+O60
XjFirtGGQuVoWsu2QkOrb1k+F2reIG6ItPW+Oe4NaqfZVKXbquoF44ssAt+a7cWHYswy+piCkJwf
btrk9CJ1jpajQ03M2CO5unSZb2Hlcu3hQcDxo5MqHkAxFKnGZdiIBOBsfxZyfuTxwQdrI4gJ5Xwz
5Zs7hyoZrflt7PhIQ6zH24rPa0Ov+5yJZO20iVmfSlB1w/MItBtrERot+fkShCRmcHZig9z8e13I
G2ebpnYQjlW9HI0z6Ab+fPWbUgcBwQ8f96zZXIpaVTlgQ/iwljCmUHonA4dT8mdCopMLxq+jwq2e
ouhN9aShbLSnq3aSB8tT7lHQ216hn5bY+zja2mXZtXAfFMTRR4sa0ztBRN72hncXM/HCEaF13ppZ
45Ana0/nFtZsa3rxywZEBM7OTuzsbEza1k2Iv11KpBBNLitW332mQGt9y1pCn1N3G7NZRStM08Yi
9NTDYpdz301Jcsp5cJIlFd364QGDUPNrlTsrIfweDXOPBonbpzU6Z/gAj1aj2LtCU71kMLJLWLWx
Pq2dGcMpuW/UfE1Z59A0Ff3EIrOIAprWDWaOkXXSyjtMOggikm5ZxackCOmBgJDhgJS+4YF02z7a
atHKI2b3VRa/QtE+dsGjz8byRTZSiqt0LatiyUHUdEHpN8vRFenms26aKHV59B2kQZSAYMMbKzQe
b6BfWnShAilZh5E0nfPe4mFkKidC83gyFRe+OCCJNA84xSQrbtzT9i6FqsjqcYwGtOWVKlpxjbE9
D/ADXnOxGdCHf+WYAhVeUPKbX2Cyi8sDiZYheMjb3cPa8LQBxROImSJhTWttRbQaJp59n0TBY8q0
tCwQKOMtdIIafMYhhvqf2RR4uQtcdkFoCleylWFypoGAYX3eEgJC+TXGnE2VEKnMkbv99OEhGU1r
mJnnXOFYbQ+mX2fNdPZQ0TgosXz0uwSNGhfSCckdgqO0kEGWxvZD8a8DdlvZewucoUxjV+EkAu2z
VuPq9C2D2J/QD/iAmMsL4RZYx64/8MboYo4XU36L8qi+hkwoEHeowF3MXVC+SweCVZ+Kat2wuxeo
h9UryfVgq6nFk0XKm0HDsFbUweiLUGfiCIFPaz0HwCfkuDAuK1NKlzJYGggKlb1xdeTxzTQgxtyN
2RuYmsTUYxBwX+aWiMSd/BrFRbZWCg3OrRsOeaE0GkZgBHzwkj/8cwnvMeZZOZaKtxAGakkVHR6W
70bDlWg0hDCnQCQv3BVnq0ckUpS9DJe2/oBL3whQILiewVn3QzpSOMuuyqm5V8y7eIc6QGvYk47D
gmnlVEqQNZQSZPw6RSTR2WyD4KCb3O8t1y/wfV8Vep5XVhj4o6y4bcwUH66a7dNzE3NJMR38eluA
jOqOBPCn79gevs3b2OqI8Oo1VvMVc6sy+2qdk6ex1o0oGWdSzjY5RUp5RQJPX9RtgXkSgBKn+XiK
mCEh2XOLP5+CvraV5XhvRlyjjng4KayqDbTS7fv66hg62kVZjXL1TWbO5M9e4bJUjUpfBvJCDTbL
ysMZ57EvVXMdfEA1v1OP04D2tR3XBJlz9p4IpuLzfbI1DquJDlgAEosNp/9e/IDzIYicPwbE2Bne
bY/JMGaKVoPxU455pIqy2vXYTumiNMwK/xEdgeHDTOZDSCdlJxMQVhEJduWP8VzNRQBgoE58Xa9w
MPSKaetkVWI5e0PSaKn4o/PtGapdBW0JLPympnCHHNWQ/kyucRwg2iKq2mbsFWvdtuz3/egunV/x
hLCT4ZIUk4AWWVc6ASyOJgZxUmvMq2fduLBt7Zrns6txjvQDYhhxQ2n0yHj6f/So1GmgJaT0hDsU
xWS9AyiqtbrOWIdwS00AWgJqmo/u7S22T9YEj5egrfuFE9wQn25Qn9k3U+BjvI2PXUWizflOOuHD
ENKHgpw9Ln8JwJTJ20qbupa+Otmqjx0k5sY2KXAL904JLj9RDW8FbGKwCMBJWz277z5bizBYKyvZ
JQ1PF/C/OPGQIqv0WbgY9m/CldpjHrQ1wxQhzefCkm9bGtn55zbFGhWlWwXfzRDPBNcUZ/rmiSn/
6yMn2yMf8pKFDD307rqEh3fjTfx6tCME3g9RAcQbTCXw9+5JZmouctsbnQSYkyvR9TL8RWTv4/Vs
nhzNuQUFvveNj49AZrh011x00M+dSh/JJjWcmxKYyh3ZpFQMY/yFDMeE4wa7ExXNyGiyKxBG2LwW
v51A3Pq80i2H/MXlXovzn+PBT73sBR5iY+1ZdNfWY0H20nOJGhnD3zB7BpqpQ++9fP6mptbPfqOk
BrGZO5UehIkJpzyLIJL3/komCvMjdu2CVDqW4xFlRu/xjz7n6w4uIC4BggoF0R5uyNoRx7867Fbn
qPme2q5P9LPLOJe2q9QzAcYGKL4VCp3gNb/ILuHqdQ/bCIiOLNpjKEJVqx0ErOFS5lI7nFatCrt8
ihAQE8GraJqVshNcDGpAKaNJdP7qC8Bsai5OPdv04x7fpLpLo9ic/pVn56TV6yia5HRMc47xvnTj
cDyp03gIloVCERPQ6ZBpKuyjqyT8dHzL/ms/ewKaCp20OOg3mLtUk3cMuWKU/QDLyIJ1H92diDDa
Aj+Dg6sn+WQlJIb8vz5HKH/hHfkiZ9KMeXOU7sA1N+HHdI4HHRXN9IMYo0goh3WKeZk+0w7r88Gq
Bb8QU+/gujiCgNSrgZK6jim9U7eC1KdQMm+YaYf8TO6UVOob6TBFuNT7NuYyXNQ2HpYzlP1sqTWt
oQHg6oVNs6bRWRetANWEo0fiiygLApWuEcH7VJ5OrpDCm88hTEnWZgn7irItSTNa9NmZF7xkDQo/
36p/N/7OOc52T9kuc7X3HtRtNbPhjuP6/tubmEs04WeLAbCgbud20uyRx3nsSGMv8Ltus+yNI9DZ
zMD8hmWRupyiUqZ8Z07Lg1bz9S0pBSjQZODffVIVcpSMYSFcsqX9QydsKjAaPH4aUpS5lWv5mJ2T
T8xjWntJLejsA8+Mcqu3jKo/JOfDUXrsJdADGSwXpG5Zjl9/KgTkydlncuukCXoAiaEpEja9Zo6+
iNfdA+DaKsqqT5FUpxIbksOKJGsJiRqDhcRZSoBQuwKCL+PZ4mtL49qrmdsaDr0xUAfUYabrBNAD
yfk2MYta/rddTCIWVl36w2Sm+chDpZO4MH6ui86hlOPkvv1lCXTeaMZlyVyAmCl78FNIQGOtVpBv
jQtknEqplzNoewKN7C8LKfk50z/aJghbv8LD2uZr3WJ/C6XjDK1pA0kMxhBoUTaU7PNp1CvHDz5P
fsZYvPSz9oE10DSZSmyYzu629863pPV4L1mttCTeAct5Ffjrp9ESIRXsdxu+HAPZFQdDykZ7//Tn
AKde2/AHne7R/veWS1t6r8v5RSI1iZJRjnHWc+EqrhV4tqroX0yYba1/fP0Fm4jhUVrS35bFARoW
H19b+JwnmqKDG3hmNHlp6OqIF2Grn/wZyzOC85kurRcisJ+TeBT087LDYA7u/22H2EaiTmO04p4P
lO/voYShpZGkTEgqnHtoByK9oGbHtJkVQV66UkSnb7IuHFpHcZ06EHdooy5T2POBzRtQVscItOq/
GQIDLp6JcBDBpuqG3+Gj+tKfg7lBJFhe0/MUISOzIsFi/ViLeV/Xq85W+MXQbuhle5W6ipU3bMrv
H0KdZvbH+XCTdOk+f36Lm9PkUNZ8+0iKmL+X1qEhekEy66+PWzzLqTkoeNKq9dkloP76al9ACUTy
q8G+ma5xMC+eJ1N3WEeJ7OrzJMGKkKl+3mHVsscOdh8GDtrv2hGLcG+miL/gluyEKDH+6va/tzdI
XcIktrqM1romgo6NbNF96Oi0AOEFhhJNu1UGdnHT9xKoK5hODN6/NAVmhdW1S6oBm1U8KgdjELsh
97zj6JRSRhxVCJ8tnIAEO+eKfhuUPJSPFoLQQcmk0QpJO58jCGwydJroV5iagN+Dy8TrmgGG/rcs
C7p0XSK5A6VJ/GVehhmvMM4J7RhYhOGjQ/xJTvpRTS+pF+74NBCOxOnmdBHMOeNEgMWnPeQrNiUS
0pTtGK/BoLScxbkcgH53Un/T6oLnCwsCUVHtC45BnWV5oQNWS6KSOxDMeJad+yBG0227SHjbo1he
6zsqJb48Rlw0MQfkG7AKDK9FFrYU1Xxfgw3HcWq+VHFL74Tzr8ipRy/VwS1aXBoHCAtlt0d9D+NQ
P4GHKyu/xd0j5GzBSjB2DpQNsjehceHCXNo3aYsDMzzqdhAI0tbbX4PNi/HSeK9KV65M8nHCgMPT
a8TQyjdiYcjbjMUk6y4xLe6LUt0sllUUQnBLqX2IZLU7o2YxAZXb7Yg67SWU0Y5KXD0Nf9sDM1RH
IdYSy4DI1Zs6hfvkbqp+VERKDwO1l09SoE5ByZwqlj+PlWHQFVJyOZQ7s4fkGymtoRsXgu8aQW0L
DhpkSX3MLZjO/Yl1VuJRNX0aN0TcZLXi/v32HuqrlpMCDKtJsMrxT8eNwLIeQxfa4MpbUfDsFjbV
HCDc0WzePk0f5NIWcx1OSNgGcu+AajIT2BcgRCMJua0vcG71RRO44CgPkdxiEDO7FhHAqhqDXCkz
igoH1YewiOFWRxGoS/2hO5ape5gfD+5uf5bhsQifPgK+naSkq4Iz7xpiSsJKjGgplnqJMdYpyEYm
WVCzwW2NehJrIFGWQOvmNm8TNZmX/pR74f7c6x2ct6a7cVXPP85V5Gub+at1r+lnLeA/ozLFL/PQ
j3joNlxRhotl3L2Kwe4T2W1LdtFVKGWonfGqMfexiHZZ3wBnkKQoFaj3xfeYr53HKqa0hfqY/ZhA
r+LRm5g6U2kC3x+yXHtelQcMkjPlZPJg40PsJZbwECPA6eyYv5rsHAjRAVLDOAf8RPmrx3boMPzl
Q9gN1ukZp8SqYSU14a6ij2itW7QlGNTZ6VjqX+foWJ+p8qY2knSa9Kt4V+3bmeXePBboN/kXcYqk
zPMdkU/mulp1Q7OBZXrLJSmkjMfv3l87ybHA5D2jj8AHjZdsrsRpM2idP35QYJQLSLXAwQXK75mX
ea4BI1fejpwyt01XdhCGZMke3WrEpvEKmsg1/Yp74Kc9477nPqr6S+lZX/qfRT8u9wJCkQiPQRHt
xILMJkb2G7VoImf7+z7fC1rk0ZXeSvH9L9ozCOAQKkVun6BTd3EYnKUjYviRkeHt0dHed78+uaPn
Cj5WQhXebNXQSA/lhJJWrFKpkJP4Q6VBvpgJWuvJxfpSpQIoHBxmAD9bOqytIVLcJ84WTPw/qHp+
TH475ALpTbKlSUxdCxVkOfaQil+XAx4vpOqKTyhick/4NOryLPDSBLZbqKF+Kp6KxGllN16FbohB
BvG3bJV6sc1WFd2bDexM8Y5sppobIe+SRG3mG0V0op3DN165sTCzchzknqnCLwBy/UmfpmbpsQA+
mxcMncZJSouBtrkuOhhzmDGEJkmZ1UiPiKHcRlj68sliEnZHRCLnSZ71dZUZetj7a0Cs1ceMgBVc
beWNmzLU3xGVT+shKeMEQ5Df7m0/Pa16ds7Q2UNJEIzE1qPvhcb5cM5QHoUJrFnTEZj76I5I02mf
ObH1RwrRr+s/nV2eTBPrUwF7Rkybfgs12OKi3JTmVwjjojIlv2af6SOFL+Tyd0/4yhon9NW8CmEV
X0d+gpUhuDUONzGzVQy5nV1cbduqLAfsidqrlltlzM45XgxJSE8ZE1jrbI7DUqox9Y+iAFK8Qq5t
Vmyn81Z3x88xSk4+5XRlsSOkuguPk5/mEyGZMXe5uNxftCDZvOrkQbDkgB14LLTUbmU4afisQ6Zc
M9X6o48mrv/xJRWyXKK0haocvbHXRGfghGyEIb0mN41uf6sTVxth/tm12n+TsFsEPITirgG0VTfo
H1vy+059aK0AC9ko5r7TAaIAOMMNLMT5wLMSA2F/vx1+byY1qiYi+bfKtRAOG1RObehdHdg2XaUO
CXhfLDM3B+yAYmb5NUURT1LD5uR6hEELFyGpa4uH/QTpZlZtVkGG/wVXx6zdXdXD5bPPeeNdziap
xOCimmcTJAYqhkD8/CkJ+X9TUuebHCk8IbDNZM3zBQ0VUcZrHv3fWuwS33EsF3XJ65hmMem38K8S
iOsiTA+4xPe99zP5JKx2aweVDbX+E07Tf45H31uHFLTs3kMZVcprBIuIi4IgdMTPc9W3S9fVizQZ
KCuWCf0IcIMxpNz1FvB2VfcfCmpN5iPOkZZHz9wtDxnq+rhXlDeTipD9jyFzCunnvU4WlFycJDNU
YCB7P4v4LMnJe3NoSpGbRHA55ZcPV4CcieZiDLJAGezi35CdDwlovThHeQebpC96FsoVatLoUBiU
gLTuO63KgU+OV629nCndovYAd9JC65pieUxkNs3QCP7NB6hrxzc7HRgMuRTfi0NkJfvWUgbJYWz4
RhF4d7CLxC6LsbaOC3USYpx2jYC7EDa0JafFmy7iNBfYImGizDSb/8K70gNP4tuJFlF1LvVUBXo2
iRgOJq9yWDD55VX3O9IhSQlXJ3FKIqP8TukXMKoWMTAi66E0NYtAMjeGdqeQOCapRpIdNkIJJvfI
kmulqsEdpt8nnC97WQ75qHfmJPLTXAPR83UI24agYcDZSm9/OFMybzaUz0V7OKaoK1TpRRys4sNq
n/bNDTulzU+PESpYYqAV5+qtVCXniRWJ/Xp5JC0Sy/k0+aVvpCWXGVq223ABXEbTLkjfsY3ScJcM
NRxt/v3SLyk3NpMeZ/5D6VVb05sH5iVDRVUImTtASaHDMMPDFCnWAMcKCGjcdMgSneye8CmOEjBL
7czC01gcXwcgSjpwzvOGKEivR3mfWyeUWwF7QjyX5Kf7YI5KLgcD23rYD/pQBJ3oELveJPTIRVup
omnUrZYBLr8xokPYuq/ZHgmPmdCG8HtpV3OYlSh1N8oAXIlru/gRFzl3cGqrzOMYs6O44vDkUyw9
cG7ldZvTF6atKPglfrEgPgD584Ql4U/gf90ZkhNTaut3544eQVUldn1nWfVNgegAWXLHCso/6NKl
ISkjZZ6N68fXLVT1P/rWUYWV8LJf5ctv3lLEjWykZc6raB1Y59/OgX4fQxXgTgTtdcqVDCvp1nji
rE+cNRNzuI/0t1WARrjgR0/eaLnoApqTErvD0y+QYeAAmAFPH/0C5xHRRVa8GMkEyw50WObSiQee
eYG7WH85pOCB111XONkLp4VB1S5MbXYujbwaAZsWSceH1iynF+HlzWrZHPrWiBkGL3L6E2AuLX6s
5S7l9vkbrGanG8GqmK9fgk9nlsCimMd1Zwuzlg1lak5XUjqh5DNW9A0q7f7dbUNYYiEN3Wn6oHQd
Brk2EWq8ftxi/Srtm06BFlu7Xtr/Vw/HjT8tzZrKJxnJsbgetDjro0Zqp7jBu+2+9gpgjbd28ewt
oFlrqkSSq7kPWgCSTggMrlvRM0ZSS8TOyx+0a/cD5qK0KcH+TicJgYUO7itUva6L0zkRzWsu/6GN
tYv0vUmn2UaxjPUAz/1AznRhsp86irU3sJnsjkuXs0u/n4vR1U4mAcUs6QdKcFCjMw//KKxY8WkJ
QP1Wu0x5HKLbWY5zdY5JqK7Dp/VX3GGRzZl+Ty2h/oL9o4JIIxKO5ETxd25PwjGfiskRJvlItspG
ZcTbAZdyyT+NnBWjzzC4NiW3d2pB1Rw0pqCT0r0zXirZV4pOSwr+u/YtScVooFk+wmUppNo3Y3X7
OdCC0PxYBe0nLme0hNbE1f7CMmIqTrOAKlVkeo8UJ8quw4/gUUJ6hBTn/qGAJelMQHCdCX4yIuF+
VECn55OAAGwvR8KIILyNcUe+CeolCuCkCkmz2gEYvNHmXCxTvqQEsD5UkA6e1AfEPt1gohHcdppd
OvdOjZv9VbY5NHRcmkh4uKYrJiB9U04zXKePdH8MrmLHJHbA5u5CRChVOc8ikvG/FLAx/lNsZ+7i
JaI4I+uXsAXQIRjGZV/UVC9AijJ/mBWYmbnSq0SNsFqtUkEUjpC68WwX9Dn99dw/dbbEv/bRN78t
u5wodKnfrrVk77QOk1rnokwnyA9lsDj+mDIONtqcEiaU4rJPcfREzkryVEMIkEGJCY71CYfQCV7I
nV673jlsgAK+/auzW09YuFUwi1ofIHGGKZwd1BJ2YIXorZI2hsc5F5Cj7m9SIgUrVYpvv/GM2oFa
b4wHN9NhVjzfg7/N/xsU1CvFjcFwUe4KwRbb9VqxNnJYEVKQMnClLRN4vq832p1+Guk+rnu4+PMv
RexJTFRcSE9qhQEWgv5gAX8HVByuSSa3yYMPHlZud1EcGRUgPyQcyafmeDCwSoszyR1EorvAErl2
lqzUX2RdwBgQqtD9/k/plMUG4Oih+nxADMTfq1vCoqG9La5s5UqjuYxQ54O/VEZtppANpmk8JkE0
Qf+IDPvpo95Z+zSLWoc4Gz/ux/pc5MrswdoDthAVIWzyrMSfeyMqfq+wjeG9XvOAsDfFrNoUkAe1
kEdMv+Ay6y8LykgFvUx//sKU+C/zF++U41hVU7Lzmps10UDsSXDdWpEYODE3qZC3udW4YibLcSJZ
M58lQdv2JKkeOclLILjuvfXakyTu+w1fbJGOVDHqT3XB7nvh1023bwv74RoAQgIvXeP0MHMfRfvM
GsgIU3v/3i78chuioNduq1eNCg0kioBVVPpre5AAmpkVmqzAEOh9kQlQ8aultS3nCidDQJLmHxnP
zqxNWM2tt29kDPO8BR1vK0lmW0ssx378R7fcFugaz5qQaLiNxBz7fGPZ7IwYkcSWHeduq5Cid5AT
yP2vpD0BTBXpaGCoOB3KyS/X3i6uSKjNX4ggzSXQG0Bu6K5H3xZWHwXi9s1gHsz1gNsNKvglQX8W
sUHrLHqBFR88OR/6H/909v68wVBBlvoiBO8Ou4VGwKj1KldPhBtN86OkwnN08stS3ZIRlRHBJjFA
ReuH3xRJjfzUcI93EH25qYT60+qCj6Myv6zFO1GM4+mQyuWKYHCYB2zub77p+hRy+JNyL4oyWvrZ
GzpYf4TBbmLDUBtx8wrfD6o1u8WbhuA3KE8GUIx/jN1hfOC0zE1tzKQZrdia0ESQA5rkRF0/2wdt
gPBafZjgT977zQ+qphYaDCiRMp+Y8NsAKBmMbjULHyhwbWNYHpGPuP0h0gAhn45Z44ef++oM0nqK
0qVdkNvtVi6BiLgMF/i8Bkbe39b//1RESCQm39JmpZFOFsBIBWGVFlauPWfRrkP41nN0SeBNckTI
W7MUCYaKIAjJJPtKh11k9gZVO5GYUD6G3VLcrHQcscISVMh79f6/j9OYMBAKoRFHSVy9MayGe7G6
TI7LUew6T4hFexVlU3R0Jalj/WEh1fjnWxOwV9BwbSHPNfHtmD5+ugt4zPb/LFPueqC7n8fa7ALQ
Klrs6zaw+vaoDWT9ctZfxa6gcP99uEkF5+NrKucwPQqzG/sSz7U1nhjf4/d1/GKPQj09boqJWF2k
Zv3nGiMYDGPF/8lJKBzM4+f+qhlH8HzZ0lbaGz+5PwtO7Pq1dkb/TuQlAF83y5vlCku0ziqKAm9N
fZjGqguK6kubBcH+X9ygNXAHabnPz0ANnesqLY0AofqZAM1BUD9vcJ7/E11u82aCm8MZHouSyIzX
K+TuIE8T93n/zNxqejW5QNo8yMW4ChniMek9rQ9VAeOt50l4GlV2Js8aAEx1A1YWm2X74f4vnin4
ALB3bLZRVpnRWZcigQ7C/tC6PMgkR9SUlJNMtez7X6LtL4+s1FclNNk7WJJ4/q6IcpRjlnbQq8sF
km851RFosQApRrKK8BjhqJknJOz4Dl1FuQ63g7U3+J2uyGh7wuOSKxcQD/Rveo57uVyIa9VYJ3Ym
pFs1clFsqp0ZoHeam7tqPoD2plPnqH3ULkDmKCKLhCO7O66XjsTaHm+o3/xNDKU/gtWev9lqqYwN
Ujhh+hTAW5LqhVkr5mAxgXHuEDrhUBj5gz2qtCUJnj2In/nZBGk2r7A+h9IYBcejwTke8ko9gOGG
cI1sBwz8MLH7YooSORkT+95i4LjUyyALn4/2RSr+0xv9ZVO2bkaABmaG8b1VmyHEkdOfKwDJordN
pFB8b8d3bdd274/wLi1ut8ny/V2nRMLoRRdzroOEEHjiGsLszDLuKvXHERaPqRsipVzPuho/Uuo/
D68sfyNtdT+DX7Sm+Ku6j80rN9uamiCgO72iO0k+x5IdDiG9qa8g9fDRz+1VuyVwm6GwviLa0WeZ
NyTn9FUh8PObNEDxsbeDX3oWod//DRAAt/DiQHDHQ89WNvXvk5lVEFx/qwjLVXhlh1+U5DHhkMl6
0Uc6vRTxKAB6oM8wOgCU8nbc5fucPlHuO9ySGuhu9vncqI4lrItzQVze25tJ1eEgLFoXUMgZQ3y9
W59+9YH67qJbz66tdKymx1S6SEd2Q7GvA+iQ+g2sfFDZJiGLKrSmNHUGdul3svLIKyGhwFpvpXw+
5AcAogdxfYKATTrzqt/gA5Q55Gkq2xAsW0OGYVCD8VvqtSniA+AL7L9GIfT2VCxsE9tnl6lo4WdA
QDyymsNwkp1mRgXUkbnJfM4FyZttbOf5l0wLFdWrkvuww1IXzO0oXJOKyY8Xc02pcc9X2L21iqYq
RNqajXwGCDlNhOEEq2TmtT2ZXluY/KG6Thh6a4rnoAzEnT+hq44qzRqk+5lzzPwHFot8AOdf6637
njcBnRTPuOzDJXPo+e8EwBk6PAow5v8wMBklmShDrersbNOr2AGj9aXzn7MyOPsncsVv0PNKAgIK
fTCdDJ/BWrjWw/2awsvmfl1IIcsfntD/DpEjFwx/zQJzV57yYybThTnWYf4xbOCdJ5dRYnHx2iAS
r4fzdtV6gxIMfD3xgFFuoSDBbHyuMbwexDR8NCfHGNdlpYyDxrsI26Cgpsd4F5E2fAxXC0uH5EXf
rIh3DCZ6ZhPYp1brFeDVyNgOz9bWnwx4YhY4tPieBtZGAdRMwrvy9g82bvJ2QdRQBdW00tXUDiRn
ZdC6bxJSRh/VOeR1Mew1GFiboGcWQhhbZd11zc69YtTu7buU01PXswqG1NWbto19dkarwPvqtDug
g1qVhJ1O7yRU3KWFSmKkiCXHThRG0Mf3TwUIYO9iONzCJL3Fr4iMwU9UASB+pztKP5QV4j11bw73
8v3Ik+d7P+zJZDRcXKT1SJ2xbKBwtxCWYn8uaUDLNaViKNY7lywTyFlue7/GDMIIQdgRCbXcKjXz
69CfLJKtnsFgNwpNp98thAkBo69sFYYhjpJTxmlApqiMXA330dJDyvwlzWO9DtkJpAP+Io817LRw
MTfqBdox78Rc0HRnlgsiFr3WLOLxoAsCzrftfzLP+sWuovNS9f2ijePzkK7GASOkvSSxa/W3p2Hy
NvHNzBxOj7Zr/Iu8/ZwRxwxQ8DlFOqlnkYCfDW6maxrhGlGFvVKUGm6Q+LygNxFTx+l3j8gKRKKk
+4pw8BcUolPiYMn+VmZhC1WMQomr8K4VuHJJDYRCsgcs8MVP8uy2T0zkruUTMgWyCc6/SFKFQPxp
CYYcOYCqyggJ1Zt5+R7aKH38cXQKIeWCdJNdoP9nqQmfy3Gxp1flgMAseZAEvBMmO46UBOEcPahB
2He5wkNjtghr/e7LC4pWlvYF/uQlddn+oyJYv5ZAPRVDKXsSiZMi/RW421kL00pNXvyBGNphwCRw
jyR07udukQWonVMfAFwhl6XTNWgKJp6eOO+2pBDAJ730zr0mBMkhayDtJQ0OP6UzWqsHkBOHG3NP
g9Pcz4Tat3NFxMcdKZxUSCeO1Ogbq61ZFlLGEqQQFAEvrajQ8d0k8UBK6l1Wg8zGXVj0Dk/pmuJZ
TTCH46vAk3dUYSWqVCqHJPRw49OpCuNczAzsa9mX4xdd86TCbYBeyqoZc2JhTJ3aprQNHRe5koqG
A9rMQCfDfWJCLEtSvfZ6A8GM6dfnu91OZheYt7rQ1QrzMmMZpzm2y1pQeMfz53tCvZgrobZdZp+D
oTzVYuuI+4BxBPUf4r6+oXf5piJSOZBG00NL5JEvKrekTr36o3WwoA3cIeAFW8JYI2G5Zb/5UvZ6
ZjvTdJMXJ08aXqW3xlt03jaaSjnq7+lWchs6YAPVGB0GXqJBACqCj/3i2a4QEdLy4Y4l5kpyReUa
EDV7+X6D3UZLiSIu89Tku3xsyQiOoufcxJuWftMIyntiyNeE37wnof/dUG00c0ZTQpLOk8bZU9aq
5BB7pklKfg4Htr5aTUxglH6GIto56hsin6hPHWkowfvqnC0qbjg4enOMBap7Uk1+nlWwxxDRWvHC
JRBajfQb84U5bDSEIcPXUiLNiiZXzrNNr+g0c9L/g1B0bFfrvwhzHyWuLTWnrHgGqLJGY06LA0zZ
dYJlvnEQAXErbGlq+si1gAC7YdOIdY/O9URE1jMiFuj5ObpgWeHVGvec170AQE5p2ZnT2Cgp8HpP
c2R12qUxWNmLIBz/8/kc1saK1QHlNvlbCq8RTfeVPPvVt6Z81GjdHRF48R2Ao4PrV8WVSTBWXKId
nkRUJ2TmBHL6Vh1Vmu5PQKIdiqIBa9PgnreECP9diDKLFRBGDTm+0iBl4tLsFCjFlMOXI9V0Lvox
5G2LHzzPHTXai2NRnxIk3k1a94bNtV5nIprfZ/n/rddNcwYsyMZOT/J5oltPaR+WYe0LqVw6YI6j
yvVlS4PtIxBgfEfuZWKAC0cSbrEnmHyD6SL3aQiBbaKfRYRJiDEyj7CnciVe0VKtMM2AjZjq0ON7
0W4/t3C77oIMpz9AnhKwCIm41G9fM3emCY+Q76RCE6ejArIVxrQWdD23RonKbCaMhX0WTyCHTEW0
TGKsgcPvwEGdLgbW9wIIULVBFr+KNqhamydjqiMIBJefYme6zpkVk44iFzGbwfz2fZzrkuUAXzSq
Jpzxqq0zlmDVwtMEWL1Ao2jSV5RGzNoSbht2mYXiNVkGfPtklxXowQQxkn3YqyLMk2f6cN3Sf4Wf
zp2Y79+sVjRhRp1TYWgYVqam8D/S2P6I/ztUXos4X9e/cNDuYBgr/3nIgWfV5ATrKCTvXW57ZSPw
CJtMvYMRwbe+6Hx9KyJmRFr2EOM21jARR3Fu9j/7AJFx00A/BtXpyV9MXBiJFYMIEjU+BsXHLMlU
ihqEDmAwoCtvR6CeGLYZXXkNSD4Tv70LmnlNKvPy1PHTvou6j7ij64W4blbjwZzvMfWq8y5fh40S
UcfSKUn4axem4ww9F27hM0S9uECf/zHYjdo+xiUY6b3iqNILf4CrB0wqIKu+H4AF647WEKvitPDQ
A9/SQrx0eSzqtr4kgKP64Rvk68vAPEqb9hq0SSjvq5fshqknl/nay9oljBJ6i6ogdljk6Z0CzSV4
dkLsfRL4XfUd/pflCqtNxHc2q9CYEgxATVhOji5W6riNR+zVzETgN/b/B+XsOs8ECcANINb8gwH7
s0J61Mw3wwjVgam5s2FeDnSHyCZQwqjboshquOklAT+QZoFFG4moU0zZSISrNDaykZ0DxPRiOI/i
wvto/TCTm7lVZAyZSx3Tg0zX/iT7qdHz4EF1fRYAElzYew05INAu/Vz2x/tUgDTDQyd2I7Z0lkIE
sbvMdJDsppffhpNp+VETXxIe1WT0VYK5mComGiCogP7lHobI8WkRRcsPrdAkcjODOstFnwzl9fvt
meeLwInFxZSvX5P2iQ4wcfFVeI4Tk6zC/sfgBjHt3Fjn66oqAykcLIHkNVaVQifasFE8Iwtmh82L
wzxNuTGmVdMf45mSKBTGF+3KJVwsvUG7J0MxtL1fk6Vqg1ecwEAaqsWdy2D+ci7ADWHFQh584hgz
VdneXyfAOAAmWpLboEoAUDAexsyautQaKmv6U76j69PnbBONIxBI9SHdaKGn37Ma0B5h/LzRPhq0
2/MDuLJo1N3JGFiODcOz7Ht/kT8uZ/aQrdKA6mU0IZ3LUFcO2ngeFdlhwhzOCw05mAl53e1+LEd7
YxdypauFqSod7H9ckpoGYrUDu6m1Z1dfUTauhpZ/F7rxErJ7Inn5HO1RBspiRnJ9L24yLxuBVQh9
3/i48d+9tP/6UsPOcGYy/zhoVY4bnIQfTJxPmr/bpyo/3FGyFEi5yZfg7MK7Aa5OR49zO2vbElIn
KHZsafFJ4mE/LWTWZ7HWHmqLorSps7ofDsZJ5wf8lVJXp5tvbCOITpw/XfxlMO1E0HLEV/xnlLzf
SsoW7mqc0D+ke3skLZKYCgdD5BlXogxH/yGks1BnvKUcxGmGgDAUb/iqlQIXuZ7DlS6+VW4CL7HI
vV+3MgIus7KF2UdOWY/BA55dLQf90hpt4koVN9zUAdPeQP9v1oM6tBUSbYoih5R8XZwhL/lZ5Jgc
fZDPGvMg0ZOEwdDCUFfEzluh95q0C0isFgQ7ANvONoTH3zh2D02oXWJ/WkIMxaYVNuFqZURQnGKa
ykXBri9DpHedvR9lVjJmMAXsPbzwfD2IysQL902QwrTohyIuPW40evdQKYpyxH0ywUCjIL5HdYMw
BiHfKmTIjsXxambVF27C8KkHKzEgHXuG/PzIqm65vthVSFhv72pLmrUzdgZAMxfXZP7hqzSGjzMl
ldLHBk7gNYtFapGy7Pch3595BLSOnQchgeBjfkHdsMCBU+FFeMFQdVCbj+W6hdwZJ4LjEkjNEh4B
xH6SqoEhqp2jO1q/049huZ1gBvZDKz367iJR9E6Zjzrc/srIqqA0uGN8vsvVs2FwIPibB09zGWIi
h9CGYHC8E20rmRJhBpmD1PbI+IE0UkRxJBOec84IzS2jJ4N3JmtKXMy9z3mTFr71Jkr19czzE4eB
sIqrZiqY/KnSy4POZJgmv32wslZrvkdp+/2TZLlOvgTGnAJJHi9daCNwZcGyf3CghGY07KYohlTv
3qol2ZNG8hOAT7IW3UprALIaRkXvqofkE4p6IdZHtMOohQS5py4XwThTKvVLBbp31EGKeGCSSFgq
x0i9Br64el8OzYtBq8hy83Kk9fpYQAU+41P+sq/oJ0k+tH4fils9juQQkX86frBFylGstut3nmHH
F4MMrHWN73NzLKgvAOXAl9umOOqOqIbxVTLyF3AwP9/sM+kceh+BWCTCuKgKoHVGR12Rr9IgVXXG
5b6DqBV5el2aYEZI74V6rVITujhj7yQbtsfTJ0KSHDdFhSMkBoNTzCMTaZUTQqtEGX+Hq+wkg/CP
n6JFEAavsHSz6w51c5Ez0/RM3Drq88PuyrCcnLcQbYDHP80dPSCNzkFANSW8fp4WrViuJJV+ny9H
RBQgTCf5Uu+UcSxoO+z4UmkmlDSiZ14j0rVhsA4g0uESGmMhuCpHYimnltwwlEf7akyNz/btE/Ss
Utnd8tJSBEqdCBV2zWqnbiNFYKWsXSrHs4vWuX2PGRkkFrQ3q9Hex/lpaXI+aUxfUrQQYu71jHYJ
lgPJMpnPTBHX6nCLHQFmMOLyL8kAT+i0nCUpYhafw2SfpLJ6Ggd/j2qdOcZC6fSbeMKROFMel+He
W4Km2yqdu0dY1EnrLxtZnkfifuEyQg3oD3W3CYeuVnaZCeQuy/9H1vGTQ4b5sLUtlB3rhI9/3MNn
HA1uh0tqXqGySp2xiejQhLnaTta/I5/B9rsoEKVDkFHatmVxF82ay/zqUlu0LLdzTYL1z/FvApGp
ioVhFRQwmgpbSZQNf6E1v9T3080HF8G4KjErKvCzvdUeLVLROhrxP28fZhN1+A3qyLA4SnoUBeMP
2YSYssZs+GO/VFtA2/apmpzQIZtSOQ5J2t2RpVYOF+V6JzpzlmzWiJSwJLm9TGU5QH3dKvfTK3fd
HQZIzuLvhr8LozbtH3n3pT1aQoUE776lt4HT3dmOtUsypaMQpzl5z6reOhefbFYzsRLl2dj0sFU0
Znslnh2uVUdoNVI5HcIj7rPm7aO4CK4ffgG3UezHQAfnqa2NHhgaiG5TEMlowaOGrdq001TEeKG2
M4Z5zHYIdNObP5H8/7F9ZJNHSoGboh9cJUZkXadIQNGNuz43NT6yi5F4ipvQMOf5SOtRGhzl2bKR
2vprq+7fR64fppQegrtsbxp+ZrcQUxwX9NBVj/3ADOZI4CRuCp7MARnEikAx+ZXSGJiVGPn+LzQA
SOWtHZlmmkWczwSa6E05k3koBUJHAawhsI+91BMAeW1NEbLeP/w1+Um+UUJkqxxs3EvJ8QiSxi5A
961ImhmfKn2e6fSJDM9/SuOjMRu8dHpI7HLu2/V28XWSnMrU6qz5jMQdDPjq2ofefH+rk+Kebbzj
IC1nL2oE1dGftnbUXO1XtFx20ISg3RvurHv/3ZjYxMClXKp0S085/95c1pEVtEbHyP4h3v94x/fz
Wo90ah2BUMBmGZb/U3nU5aAlBKe/nCBUH/pQDWmnEuvyly04G+xRQT7+voYAKcNpTka9qX7HdxIR
UI1wY4bPDVk5WOQNPVQrjkgs5WxrJ95r2YtvuYu4iCXfnynKlcjdAGXIIlXlXsyn9jJr5jrde3Gk
c0WoxEsPvMMhmNkj6DAdyz0mAR8l6x+JA3se6Mb1qAwfdh/K77QoXWLd4XpamTuPmEljPXVGUMrt
KB1whKiLspGcOpgZYCLnnNL7NAKCATB3SbRL2qDChbobGtYDUhR+XgwcOI6L7jzrlF1rUvtlA54p
lL48e+5fB44sWXkKYmXM6Wo+vLR1gcEwBoFwvi1iWTJ63FgeMQ7iFTfUwKvypC0LkS5WBrJvCDhA
V0quH8cHZhs4tMEKPvC6pnLKjDqFyo0vB/wn9vT96Se/DJGHUgIdYrklag9Gxkf0f0HUQlKKILpv
isUF/j00khMSGPtVw57IyUnmfT7wN2JIKYVWkAf7NJKnSw5SMdjbq4w7bDW45z7gFGzyAIk6EJYM
pzzSmm+whsCgOp048fx5pZJt+U6v61oLrtGf54rIT1+VXFWdxAspweJlV4L3qNfd4LuPva/AIWnD
ScErusIYzGgHX4Hrn+ZuHBlJtaUexRN6BNl+XxGla1RsZQUSqdH9HIQtE7ZF5lJPxmaVx00z5bgh
8aZytE5fJ1cXOBR+SJ6RKwYsaQ+0TBkIeeF8OVe6i1VuwCwvYuRoRWtrh0MKjh8zeLFhxZ9uCoxf
CvuMIuogtAhA7Zvdrdq9GDCl+QYNoH5SRiQ4bsoNXtUjF4q+og8eG97XC1h3DdaovIYf1qkFOd4c
goSJmtNDqDWQkKb2BOsnehTLxOzE1vzSaPgfgqCI6dQrKVw9kpT/lyD1eSPS09yta+eMRZMfR3Nn
XTVZgkRnwqMLWOzPuVwRzZxTL6+a5EvzrUEebodxGRTyv16lbSxW7SuviVjwpIEEE4YWxKqLo9Ij
ka9ypI6MlWi2v5kKlMTzI2JNJWWSoPD5L8UbRS2X9RBr0EaNw6bHt4rXFu84jKuxwrITRqJ/jBap
qSZxp855oFbn+OtlG7TcDGW8uTDV+wxzmYIRygkPJfs3guWDFRJxwcLjsNbqnF/o2iBvR09zPc6Z
oaY9l8hQk9yYb43FKUYH1PVr53KQqdueZ35khBsF1u7nYhsSO30qAhAMp7e7wMIdFonGVwTza4ls
+buYkyD0VBJMccApekKZgPcf5C/piar3yeixKepy0Ln3cHjuQBNd6Eskqtc191SlZJH94TZ+fXvV
OfewXMM8v62hS+vVr2wOCzfI6jwnU866l10Sm3yiaWgLucQptpYAgSZEaQE4d3nQn61pzGJ1M4/W
WVChatEpF0JkOflwdiPdVm13eJR+VndYWjCemphXLaMOHrMBUdIXRCbwESvaL080m3IHG1QLnCxN
oboc/YkShlLdBUhYbK0D1hPhunMQF6+qgCCU4IN5CqNZhAPe8GiFNRNpCcx8awNFRvofGO65ouDz
xgbktaMH65aq8ihEsVgSWlKTIRgWRwlPtZzD1dPzKMBWyQCo/Qy4fe6AgO7fQxgH0GVerC4WJLVP
nfqJAHttNWaAXbKFsaII6xZExcXJXGYI3CKqJEyo4GwuEC8CzV5DSqeC6kE1ORWd0dAVdnRJR3W2
vjc62c27FVa6IXPwyUQlfQJ9nR7MSRmFGf1jqZ/c9bLpvWEt1/jJ8joBDR/XP8R9QSJVZhWRmQHF
AS8EAhiH4wz4m5UG+zdElaOg2Ttd/MjEQKb0FU5+6gZQ7uVUp1Yniwrguh4jvNkgrBM72f6FdJfW
co3eaSKBjevTJPaF1xrpzP3MsTy9Wbu0qTx/jGUrK1nMDMOhiffAMm0zUaaP+8NcSz+lUABnsxNT
z3/5pktsbIs4YE2/bvpInX85Tonxvfox/zQ70YPxqKLWRh7JE24OoYZOvSzX5hwhPMPAlvY6EYXO
lCd7kCij4Xa96ft72bg0jZAJRKscbhV6Fll3bFN/Oi6akuu8JaBezIyBdXC/j1lbDDH8UqOD8fFd
6JDe/+H+D0PjcL7x0La+rKzgyxK5rNNX5+//pXozC7Em1dQrTJzU5meaBHnl97o+ZVY7Qm9VpkaW
ruyyO3kkhQIleFX6r1PpwgYT7t3QyDWCt3xB30jL6cDjw8nW8Plr0iAbbzYPW6HQMwrSqPToaNQ4
Fa8kCtdmcWxC5kUZJDp7rxGfl+dPicjCek2A0S/sEWIYqb+D4Zgq4ALpHqkjx511+kZfVti2nPeY
SNouhYx5wvjk77O3eCsy4jWc3Hy7lVLWRbUyCD+CrE9YL8vuA5NqpC1UC3Z3llrS623ssqbMytDD
0FqOsRI8HWDyTGAV69SZnALXLyJLZJyrUKKuFKVGy9umUuDz8crfiH4vHm/HdfahrOWWtBCmUZT5
re/yt7LFXjCopKtEhsuU7StTql3PVF9wGHmbtVJxeirq87tZeKs3PcX+b9Vg/TFM/e8SZm2Wkkwm
uIVuDD/wKXFT1WH2f625FMCDPyuvydnQ0exQDlwsiDxsMa66rRh8+3CnRPEM60FNsfEJ9W35p1KY
W+HcIa6JzKif3TiztVEHAKS3YsnL21tisWqXoWzV/p5kgPmI36boa5uuKWqWLzJA62uiCuMuHyGG
v/udIfZNAo4axyax5B3MVI0mkbVjmyZN4sT4gxKhVbuY/HjqhA7bgOrH5fY3ApRri9PmG/jZC1Av
fJkGa1bnLSlU2IHxVUNBNNXz4iBvDPrnoglJzBqAPc0sqejv1x498QpEzGlB85lVtRN+pMMTwJfM
A5KMT3I3xmuJ+7r84yerlCFf7N+iqPzdNhtS3DxgMk8CuuGqg/IvF5LKah7meb4J0G/eVHf0XVDZ
Mi/SSrbLyyCFpiRXoOWGhphhzya7tJaTHObmjVxvHIpzlRTzYhMn3wy6kPXKykaRKUJFloHNi+HP
DbnXCmPqX4YV7DBarYWgsXeb9rOsnX03k7vame9hp1t1pmFKwHKjuX2KpnvxIvuU3s+eY0yqtkkU
Wvc4Ag+p8VIMlqsN2PaLMhlJLQQxKe21VvyDiQ7eGVPF/HnMIBjwDE9H0/EmY7boM2IFee5XE1CO
rQ/jzXjkUEwpdlnn1NKCYJUsmmO57v1VyOTAPG4L9dYVlcWpvosfdBFsfRrCXdKeYGhuofaOuEsW
HB2GR39xSKW+tZZBHi13LQWSUNOdYg11YFbYRn9scuMPshP1nhyiU5TM6sRJaoOB2jgr4EdK2k0Y
ncS8pV19WoQPBZTJUnpJ6Knb8F/I93z9LsCXCd/EvlHlHyr15LjC7+nxD5rf//fLQ4BZQGeRsaVb
R6+25DgkDV3WvIwRz9lFmTbPxJ5yD2DDfnssK6vFOuJBjrLGvZ2XkcdGjdXvWgizzRjrJLujb5rH
lSMQTOpde/gl554W5jVw9EMTl3dWI8Z1DF2+UK2q5zKVJ4SsR4m3Eo/VqSOqri8CyKtENLia34ir
QrkDYYAGYXks+4ztLZaR7xAmZJYwo59cPJ9HCvg2e4/lBCL0f2X/Gi+0hhb0T0FaRYAWMxO9DKrj
DCX1O+j5IU8QSBLrtbwgveIWGzL1ep+E32Bm/4Jz9VNpJPVUK03smtHbqbSvnRmPncSbgQO9l2x1
g2Xg9yjELCdsjqwMkQ8tyZdMcQpSE5TsbhmDxYlmxTiV4H5q9pDAs658eb73wHqV2ad/BkhX5Mgy
t7bjPXhjdfR1W4bWXVTzYKq+7aEomcacTMET3XocvWTCOyyvN00+CCUwSb3etAgG4kpjHBhJs9Rj
jGZ6A/oK0gCHacHU6UjaRflN4ZXIzE+sAdB3WYvTrm5+3sgysRHHBxk5qCBETkatZg89tYIabZcY
dDQ2LTNTwkWfdnV8kiw66uvp9ngga7IPoPFpg/+4VpLImrZc6Yl4fXNs05vdzBwGUnFh+wSljAmK
O6+i0gQ6+NIL79ycGFFPxnUsA7wwJOj5X+DvyKEI2uBgZr0fW3p5+PMqnCDD2L3aaA7QzlLKQmkZ
IpivHYqvVGWIcTn9ZCQBpNlFEin8wirFTDk1lJWkzjvDVaBJs3y9kGMoZH7FSEtXTzlMnjgDvpxf
Mmj6uprNE9pFQJwUAaJ/VsffftX7TKYvlT2gTafuSOXdPwTViUoSPZgJfP5U4ngHpTVZEBIX8SFj
Se/XFxJqeSCA0zDhHP9QBKNreFQCQC5l6TvVBMMIE8CK+1WVYiJaTeRX1uIkhqDrJbkU2qjb7LvS
dY+644wmHEfRAXFDzDhvkt7/XdYnjJpqPZOefm+ZNO8q/5huKKOseCGMAwcAB0d30297h+ny97Ll
KbK2u0RE6wiXGdwwA/Co9HR0TpLYJ4c9W1HmPAZMJ/WlCjzgaCya9HOKHaPR/0GLq95W5KZA6odo
92tSgf0QRfGZ3J/RTAA53HGXLjEEfy4pOPH3BpPOh8MOgypNyK39veAIf+NcqhSXVKiAEFv1fvOX
8I/tlQcYaL4fFxxrMZt/eaUW9tNBBp9hTR99zbQ6wqg/GC4unRqctjty0tvWPG+LimKVpDQVSxoP
NPr3hWcfQ0jlKQp+qBzunezwqeMGNtmGi+7KYSDYriifxdxkGogu9kfkBjkLBYs8bv3O0Qn2yedI
/zkxEHPLOExpJlUg9O7hIrXmOuaXJTobt9VOJUZDJ5Mdk2/NLmjGhPZT0dZRqfdgLfOPixcQ4ALU
L9hEZdNVE+Cm7L5QyP6zppXtib06e38F9bCt7If0lqdZqzkVbBwGi0TWZJtkOmQzddud57iv9bxl
ygw0XXrfPPzVfQaKSmlHhLEMA3dAfqv12dYNySgXutKHO7nXJV4fjT9jaTWuvk63tOWJI0WkuZU8
eTpxDZpLZcFpAo+F+yxYcIfRGEIZkSxzC29EjYNASX2BcV97ILzh9vM0/rx4uuWjaXVoaDXc/L19
QEQv9SNPlCNVgT0fqFR6cBwzOYHgWy1bUZ/s7/zeN0jWpvnHnC7uvAkIRz81Qbj0ICUNci5e/DZX
4Ra0otE6CXGGeEM1tq0DlLgKQzAKtd+NP8hwRU0uuXjHaeALGXlekCbvirAy+UjFqvmviWngNLkp
WBzjInazJ4EUTsOuWh1UE9xA9gZG/wMtDgfNH6VV6crRTbJgqgNsRHeUMGPl0GOA8aZ6yCe3gYDz
dxu5dOaQelm20VTFNhjwDQy6b+yg3lDmAzyap0K4lLj4CRS1gUwBo3Z1TLvUwnUWeSQp7mzkEK8c
nVnxSu4JxrLbUWo5oOEBBEUs0pU+DF421kp9t17a6vPzvjxsi9c5ibhcEGFFcGFTjjesTzyG3NWf
fIbJRoqRDMPWMgNAqV8oJOtQUocfB9FyVf4qMu/+KSuRjF72RyjVG26k+HuF1+Zp3Q3kpnSttlKY
mFpOJMQcDNbmseirLA9LmmpkSpenoQkTRCdMq35zLZZXE7pdyXy8tHd5TdwtLAAXlBfTU2ifN2y1
M7BzMs16xWoPpeqbUVQQHKEwNu7O39N6q3QOzcFZAiVtzFz+HpN/fqSY6X8h3fhlMttZahpsZ+I/
3k6U0BSMN6o48SfFj09kqeiYKuKBUmnQEmRhZ1sl1WtHK8RXQd7T6VKWqf5Bj8VhfSGGSC7naqd7
Z7qhGMhA0giAznbmgRvNsks+pV6SRuElPaA1KJNk+vgwNrbWO2QCh2zzIkQ7qcvUHbGuk+1Y56bn
ClmyLq88mwgsCOQa3HSZTCaKbhjWLRv+efPQtIi6/V/J/nbUDj+GE858qjcX5rtqwSKNB4vqKsoN
2NuBHIGZfkCPMNZXJpPcx0a80APD4VyGzbrGZefG2KkggODS4Cj0veQIy8Vao27biQd71VRi9KKs
yan5jajJlbF3j4zsg6HtsloaSDIPuD5yWtEYqFjs04VQo7ZD5qC0r8JFbXG6Pb8krO5JICLaBsBi
OM4V77VCH/OlcY986muCxhFJIGu7iWZh0qHXl02ixNO+vCnDuFQrV6pQZPdLm+I5Q+y5Pq6u94AL
w7Ejs4Qy5OnDV3Mw1pW/WhasSmT66wGpGG2RguL2A+9auYMe3vOE/jGva46HAGbuB0qkKgcAuWaA
bt/qLULh9oeGJpo2ek/0IFMbFLPnxlTze2hXTTcnA5wcYwWnwl6hUqskbAAvDHlq0yhb8ur/aVvu
aejlJB81JhWt8bnThz+7yf/PF6o5xQtTyWMAzTigCQt4LBvK32ReU4bMEHVLuf62rxQ9zBS5KxrD
sZ0Hk+zFty2Tv53p2I52F05z3Seat54TIcBVnXwIbezq4AB9aPbn5y8eJca6a/W3XFJk8LLwj+3a
aiAPGI6uAOBmK4zTtY95TFoIeJde3ofxIb9yaQ/lNGgE1kG17OsGJGRSN5olvZfK0PLD1bwPmH1S
o/S6PPf1+Mz965O4bu4IvemSQKwZrFXx1TRv8/xOnk1Fz8T55MsSS+CalvjxHcQABx4x87sKVMKk
pWUlK0AZjyHNkHYqTAfAiqXlko3NpAKzLIIQorzkvmbf1ItNC1KRduoLQlWHaotRKOB11qpV+Q5M
PBo6q0lEV66+tF84NG52Y9p+Dt9yJcVQ+mCCLE9uCAg2LP9XD46dOCk+VlomZVKIY8wk4iQ8VLmI
OVMHah4kN36/laDNb/3/hHg2NTj7ROGoNZ4BduPnnMt8zX4sWgAm8+zc10I/PHC+vwMBF/8yDL4n
kNFYAU5VJALE10tVLwCIZW7OjMgZDEJX9aY26FHAugJuYwhLoOidZC2Xgmtq/0MdqWRN2FTlEbFa
AEA17K66XazyS9csni5qd4RoRjrwMLkqAbElpC50i4pirFzA8L7rczJPE7c5UBa8t4jm8G+5gCEI
YnI6zeV8YHjLfWqTuB0Uqc3aJz0Yj63lQlt4IaGxCgGuvkjuU3ZZK4jVB+P6EJI6Vg6bMmsXecFX
EGPWzUthbmaj76RgdOA12fLi8DWD0qbiNgf9uqRO8UunJfwPRdIXrCA24b71mvYHvxjKNld9XSnm
AlePga6Y+Pyc0pK9ZacX2CtqShYN9zUe4hYFCLCoiIUJ4Bs0ZtM1NDwfDEPmrRGt54MwkvmchKnJ
NKAwK/CW6OOkbWZHpwC7m3IxrUqhEyi/VNsrt1BDZ2FVZV+d3Qlwo0BA0exItafUnUw+RZu3vmWe
18nc3peosGaDftBO6/cnypvMwswkg5A3NLgt6ajvlZL2uemRGe+g9U+UC3gY4hoJoxDjU/RmQ9FV
tZlHsR3HnNlMZjfYTKErAx6keGKu/ovTI/Mm2h5cxXPYqwmsO/yotQXewDBKWUAeAStfHWYKiPtH
vE8VIWpWlmYXmri9V9DrTEenI0g/vm2oS4qxdgD8K0B6CuTxtKRkwS7aTrpU5nD6QdZojA9eeFuq
buYxem2eS2kt3OQ+R2hDo3NXFuyCAIhwPSwZ6u8uRc4ecIuDVPIsvCv1FuJ/A2llu4wHgr2ZQXM6
5ZwZN3C3z8kpReM9xpM5aiP7gsrlB4OHWRKehl/ZMFi1WO7/vRH3TUPSxK25QznjCmtkQaB0lARq
c2aN+p454jR31GgwUS3B+YyloGvPaSOOozeCJ+OZ0VpmXKfg+IUoilI2dgZNNVRSc47YTaNXGmso
w2UZFNIIY4C6ctqZ5IQCskZzl4EALfcjZTgeL5rEn3kV9h0vC7csQVg8KSLnecBMCoCGKth9gQBl
rtPgTuiSH3zo/ctVRw3wHCvYLLv3U4giq8UTYZLf9n1L+abqM3MtHl0BZBZY4KVRRM23AMo/QflQ
X0U7qywIaIpIhOtiw0vqpN5k/HYVtIKYqgYlABWpLDEi5eJpgHOp7woK2syoJTz45C2gZuGIPz4u
H9TTdNaX9VekKhrOBUry6Mmk6su0V4RQDF7dLPsoYsRH4rf65at80UlHu22QCXzsmgW1d/vFDB7P
vx3R+0UmkE5OmqvZybQ2FjWo/rFbfEPpzVzfuigDi6yJzsA43KeB7V6rimHrrthq5gptBj8lhv+u
/Yins3pGe3Q7tvqNb/zRULrO28a5Getxxh+11l6Sl5Cr+Ap6eeZZCw9zblPr8IKK32K/ikbna4Ty
VLspvrIXns+LJqAgjoGtIwPx4yNYXyoMzpWfBvbR7rkHl9B7J5rNKw7xAoz5Lmnd9c4MnGHQvKmq
TJ6A7A5lVGyFJXVOUMyPiAKV6QbK76b7VXlJko07P3HCjW4i8Mq2b8kxajakN7hMefaHs7LrS/Ov
M5tId7RYhd4K5UEY+GBCp9cVnv4Crd4mZDRELQcLxFj2L6Ff3HlxZmI2mZVu713ic22nXeck/5HU
oJy+T6TOz/cJupZapsHzxDkFMNgLhlzxLPmuECTJaSpn+1PlJcEmYAaab1p9lesYZ9Ax+v/9ruEx
RwKO7OiN20PmSJA5gge9ywaqsqTKuT9eKutmwmN5bOu4TQroFcGInWN8dbOWFrLU/LJSg6N72T2h
a9hpnrUzo/bfdwSJy8F3a0qrVdf5AsYxKYeOq2IJVltLPgDMHUn4vwvvp5NI+UJ3amanCKPDQTi3
9qpYqRg0uHhrYu0yFZoDkAquvRiSI7MJeoMZt5b/KlWqtXoIuGS00gKPGxp4qVk3a4g9b+D40m0B
jPxZ1y8U0syQwpjH6lhsolu8aQZNAg/GJqtlQWlZohzDF8bMpiKBFRaC5UJYpTKSsjDankMGdBgc
D7D9xkrxStCdYFlTvHILYG5TzfsjuIVbB1BZB+rcbg9yudPCbOWXflzmP/jX8RLEo9TcFuqkB4F8
Sd9xbJ5X2sfIShhEHqUJEebf/sDBeGf9NCL1tUCqMc2/cphYkCWsnq1HxCLHgMOQyI7vdv1wM0tD
6XWbPZKXLezpBjjTHrE6HGv0EZAH9tOYDSWEMOu75ZJCePWJWkMMJBHB8Xq2C8W73q5UxQfsVTyY
lNdbdGcK/+f7H/QpPjALLPUEUaP8PKxahseRgaCXgLyUeCYtfLwpCnY/kRPFqUtXwFwE0ulUHiHb
QXpUuPpwDg6D4MmlgRO+7AKqt31CDNcklFpudKRzHBc8n9shK56u2WeGKGJDW3QmQmYVuNhkKNX5
3iXtpHhr0/756fQPWtEj3ctuhIOeQeOw3yKABbQcyPqJnCefNvnUCqa+cuw+lQc/TYQ0lc9YFgOg
MdUP+LGEqO0m1Of5WWnWbVaZ9ypl3FA8RZH6sMtTm60OPYI0TSkESPBfoH84XsRCrisrYuI2YdGn
znBOBfBMF59qAXgVV4JGLmRz8GZgr4ee+0Rm0kIivhCvVXyJIVBpNCt8f0BwatUpBFBkcsftXMoZ
sW4aagkGMFQu8JmHktZlzgTANReJWFuq2YG/VYIwlOtMH6Dbq3qU+lSZVc5JXInQ3an16BQfBrzS
+uQrAwg0U4IcEqeL+GozvT1nZnwAHMMso9DZwb7zOG3FJ0FNgljzdZ+Ig5F1iyvbW214zEhhxleP
Q7/ctqOtbsx0AhFcbhk5ZT5rX+hChPEBY8TnVXaphsOaRGtZF5glv1AneH7WN1zkwHKmi0AgTapb
wx4R1Lz2fNfw9RGR+Z5B3V4H4Xo3rmpi2OImRiDnMdMYbBKZ4lu9B56y4aERnY+CfAWmwsCU/TMI
mreOpKUjvXhMEOX10uNsUNDyhJqARfzkHF52bhaVBNAvLepVh0uHspVcR1sc/7tXP95w3245hFlZ
S83Cnf/RQpVSjfZHd5K4OdFp8YM1gIw6Krw51KL+8BeocSDEoPjRx8eaKKniSr4jWvzLB5Cwa55H
YMFl5DiAVZDJduA0Zy9yo8I41QSZlol/4kQDEnDEy4DkAyA1GlC8c158kuHNwyPTTU9AeRKQfjPA
czCCBwlwVxUd4DBbWDVAeAd4KR9nj/h/+aqernn0HNQOONNfURT7z9hR+vZ1Gd/+huWlpxERi8yn
31yw4u4+gRuTPp0wuOpC2kUaWGZbG0eaUKno64OCXyIhF380aGv1C/hmtiR/TOsLj8ptrnDyxVdB
u15rLDh8PoulW0W1EF+4Dnr5h3TnU5vspVrbIZnTV4mXp+1f+WeUo2hlcuv9mwFxWRBmuGehXuRI
+Q6/NNrbpSIiFpn5HLTC/6MADm830bsI4LmGNjHJB/TCbmO312+YRDXm01gSjqo1PAIhP82BSoxK
Pd3Rz798Qz4eyXtMEC2/jLui/u+ALAauOsFGoSNlApFyiRvcwkcv1In9ZV8E+N0hFtNspm7LcgcY
2aasqXO63qFbWTgwgOQH0k/5gtmADYICC5341qlUmpukwXCC6v4sYtri8uzugNbg+qzlXgYzu7Vn
OMf6pGrcfV7FQH2Q5Lo/vIQNtdmNGLlaECUvZcioQwSUEoY/O36KC3bEi+S5hcR27WjMfdoWpWJT
BiRIBuOValtk3wi9UQZGDopIVdC9BT1oJSEBs7NeQAXg371vvPTaeQE5SEfm28AettxiTajhS9fJ
lZcb8sLFo9y0TmkUHxQiUED0UqeaKRQAIOz5DzjRjQ+ryWs8FEFti/jMuxJD7Uiv1jHc5IvAgbaN
WAWOlCuPeCRT6tyZJO2uQs9Hre8zvGgTKN0x6mN3nq+iW9wOE7MGeZk4NzHUOwoxOk/ax7UJmfAp
u4W9RVJWUum/5ml0e2EK5+8ssKNzRB1H2ZBWi1zYMTn9DLslMCPP/i+J4Sq8noDsFDYllzLjJu9H
mkxvafK+8wGzH7PvKIsWUQ5QwS9AH0mzskGsGHDVhAkZxqj3/gBrQvaRK2tybxMk+cdDxdDW8rNL
Pg4v/UU53YzTUyUyu0sIY+CWKKvBt71G4IdxjFm9O1J15acSIge0uVOMw2tmB+DVcwqsc2DESvmt
K4irLB1jvzsHOu+k5NSH2sLwNnBPtsi/inMNHk8PCnFMbVIcqNECNqQZItAzVAYKd5jt4XT9KuDF
esz9hWS/wdKKbBgOOMej6neWP0i8Tzjszb4Df8T1b+CN41qVEDqteCPvgzFYlIzj2nJ43tBGW6p+
0IR7sgyYBSq3FiXzhO4Ncn7AbWG0yiZ4uy6EaCTKiFbEdR3bb0sztzo+RfWdiOhqfjjfyCD35Oju
i4lMcqFtEwR4ZvExBT6N7i0ZoFZB9HBx4GGpcTybqEtMBn1e1FNIKsbLy4qtJbKXVkBTy2FJOYu+
XoHg33tHlq3jztYD7Lysf+aa41vhzrN9itwBBvaAVfT7aEfgst5UHTkcaXArf6JhilVqV+ts/Xgr
9SFtGvXcPhC50rJNWB0oZz/vzY7OjxVEFnUXAJZDZxrtS6AZfHQd6Jlh9B4HFdlJHKPkR0eP4H3B
DsxS2o6aHbWGNui5iaYhdcSmFjIDVLC+T9tfUPkB7R9ueSZ4ymWSg+cUn6tcRO+tk2mAuOBqeigp
7Tmf5EeqCUJma02Veds7QT1y0onaV0zw/nxoU6oWtKPMudGwYNReA48XwOahO3Q5I1OEW4RpBm9h
RtVZLCYYVC6rCScWBf9ok6Dt/+KpX6Hz+gcnx2+bMW03KazP54FtCoyj0+4Z1UdPy2bkAD/uGZWR
fwD6UGmcp5UQbyIWc0W56ujwKefz4O/nCMTTM8XhcnshZ+3VVnLmiveQYNgqxGuYIj7h2+e2om0S
Es/WYXx1P2EH86vpkSahBTLslnIWWTh0weHoUipkYbgXpOo7z2xmAorh/2Xc8pYKYfIKdQFMz6xe
drJKmqJskxEZr78X0aXR2XbufxAEfDUlUJ72tLsjzsOxABbl0dWfXzaCD41rUc4PM1g0o2YIyvBc
9eBopdVQKeNs09A8uHTPI5msU4s6mi7cXZjVHte5lDuxPQGWlqAVPsqq/BXwHETPcrvgOx57oSWo
3abHzAsL1qfcMh4TQ6mFAzNv6LbdjiJwQMqEgYDvIQIn5dXl5GTjiBdJAi9syb3hdSn7VeeTpFmC
j80wgtmktPurUcEYu+mOIcslxg0yCkGkPDeTBv6T8A3LwqFhHkxDn5SPctqi5nXicfHFC/W0nJrw
bq1IzgwVI671F8RyDKeuspiDAVtVfghT268iMT4Zwp/QvTwMjns5XsKlLwz+NWBUp3MKpxwHcbKx
hjE8l1vCwZJQy62C3MNyg5BoSmRvxKxmml0EDTyrvdxGVbUr5Vv3DhywxOoKJP+7WlK/ltwYhKRT
7CIBBrmnSVAEJDChV4n6QI5fWWCf67v+3QmRjqP45nGXUqOmxYk8iADKE2qj5fLT1NjWwEdcALM1
HReZZa0kAN/PLaN4fkkGahJf53qIhGf++sTSNEzwleEhz9931uVQOisNa/70CBhpv7awWgcONikB
ULmMqHpRVaDuHwOyU6/IJnEEHfLJRzCyocXGXZq55DNdFHYWWYUdh0t3KOZyI7KMhsVrsQUYT4DS
EIWwKESG/R2mIizyZ/gjWLZJ17dM/Y87lXODTuKGKCmYJNywRI09JjfR/WfGyd2IQdTdzAPrsBCa
v1oulY0tS3+W4XSIrNQ+nfXI4RXEz0Rb7q6ORPd4n71Y5wOSEjje0Cp8/WQz9AjWpkqPrVDy/iPC
dYbdhK3bB/rGwtecxlCYTTz3rIoAvJoVi+tOV5EAcfhyOaZbNS+6p3cRwu5tvF4w40Ahsrnb5fDD
EgIM+vSt747du6i0xSyyMKzjd8XlbCYzkPlswd9z7ExoPEuGxJAJ/V+qmQE0lLop6mHsM03RjQkH
rhJvNX6TigVEeIGtspa2Wk6uUfpj3ztgBfrMX2VWxeBXjO5a9PFrrF0+1WbpNTfMEPk4FwDaPbpk
lAneYTUJHBk3dckVv/P2R/XpspU0EV8pxbma2ND4xkYdKRAJ6pD+FVVxWl0WSn7oAtTGwtWXUbzb
4ERShsfgD6x3c6mLhcvpx/pxrjhanGVXvTpz1JEQHGFDTUGU19xOigAOlhWgL8j8oZ7pdjopexSR
RrjJ6avS85b+UOreYyaas4OXxrBq1hfAzIOfRPrOEbJMpL5wU3Pscz/NOI/XWjJ0F8XEUtMplKhw
g4gV4giUXX4mFMzf8C/pbMu2+JkeZuxMz//kS7caykjxe46psrJNWU/ORXghCLsjZODgnj51dLTu
BBubUvjyhXCB+wdtV4kQHPJkr0c5o9CktyXmBl4g4lhLum5QoGqXs7v0aqrcTLuXKd0TjvL6VeG2
6dBE9CRGNl2VJ3qxWRJY/m4yeyMQoRLjIRm0P/rKypj+PRtEjz1qeLzgC1eL6Cu47PioOR2RtSRr
9Nf3d+XFvFPH5NOM+8ngZCS/0TyDVDX1rdG0YfZsCixuV9R+n5HhtAi8nn8kWUNQi0xHknSPHGhY
nvKn38Iipb/2KK8XR17NtQuUG6no7zO+piR1P1E36rScXTMRguUWi2I/fxNSvMvJAeMeI5NjORLR
Gl28z3kOnYodRhlNxdtB75wjDNNfuW6fInv3icRF99ZfoxGsPot03zl4Ns1kPWDT8MP2NPtKRafU
PPgSaHbTXjpmYmcEGjAIRkf1IbmkTdvlcwXBpjqFq5kknJMVdFp36uEyR1JjslPuh8UlW83Hhr71
PFiFKry39bocktLDbbLeJYPbQwiblEyfnCRseWB94ewA8pOf6HHLib6Rx0TWM+klsWOAQElBT8PA
zP5UEUQGlU3O1uMMJhkLWzMOU16wgUZXh0eY+g+VZ+hk9NdNOTgAfwVmCSMqGchHmFd5lA6POvTn
nsbBG/adMtyaYmfLbnJSnuuoy+ZQIMw3laYLchmwUHlngI3Nzo3K1h6KORvG+kU8KcPgThVLa2g5
fdzjDwydIxT6TwrDQEZNiKPAI3WdWPAQ4w2OL4xceeAST4zLm26DHB5rDuK55JEN6+dPFh5nDmFM
RmFOw3sgacub5RvRHbQYqNoqxx0QxO6m9CHNrtG8Q7Gowv2dJrVbZ5EaVC9zDdUSSrtL799lUB01
Qpkn3UN6E5IOgJcqpC8muke5sgaW2r3D1pdlkzQPsKZVSSdL9GjhMS2iRoSfAmqZxMmC8JfKb5Xm
UN03sXovHutxTbxrBvOihQ2nYalg+fr3832dZSFyDy4qkqFSCOvbVJnvkCsoW/b1K125HkscW2rp
RlkNm2q0Fv7eU7RIsXxWPEpLLXS49ld1h5YgnO6sp15gZ3HTcgUH+BKGvQnRO+nnDRg/eNcv5P4f
xqapOLmCSJQijrYki0lLjr12JU06z79xk+adOgAsBRfLVfixrIDXgsmcz0cI2NDICicYrVF2ggpK
CXCFV3E6/4re3b8W26532j2XKay+Y0k9/8QqwaQROR75KrjvSCyYz6Q0AD+BeqZqI6XAm/TIk1wX
1SRjXgMzWLDQDq8lGDM6FaDZbsT5Xc5txywbC/LMXSmeZppeBPW7hq+rJzT18NW5hp5mIqYZctk/
2EvXrrnsb8UAcaiLt2Q0ikAXDVxRRDY6FB19hSmN1YDNdKbzRW5LY0FER7j8auvsqP8Vrau3ZTVV
M60RufhG2BxUqoZayr0nMSDWpbuIOMlSqq6viB4Z9tZUO6a9Vl/A5CBhveFpLrfe/MwMdoDhgy5F
flGQKnhQfzIUgSe1tNpfBBB9RB9RTRw7GcDF+Pp92Qt3XvvxlzobSSMDUd86EFVZpv44pwAw4enU
LGVcHwTiGfk8/5SUOwjSG+lBMzRFQd/Ms7xq8zMtVEw0MuWGny4nJVBp6SMK0TXb2oG5OLCPTbey
YK8/1iMFODeWYsmxkcWiJ1Wkn2Ru0dcMAPziSwL+tN8NMAPJyY2W4z9ysozGh0hUrrrVk3zw1aRM
1IU53sXCc9Ih6UzCUfj1wy5d/AUesV04O5Sw1RTe6VpgRD9YWa4XWuPTct4gnjrusduWb/jGXcWk
6fGZ+7lDFQfYu+rB2QywxsGHDWFNvPyUh/J5cDhgT+5TDX4w5+0SuAKX9qdHoOAniAyN3MVKrBYi
Z0+AeqojPrTIet28CpLUmQzyQ74UWcO9rygbCz1cjR92XJ9UxGKBZYlc93FJ72gIbIelBfWa085M
YEhei5Lv/O+oMbou9KUJPixTq1+uwOFzaxxjlPqMQCDMxKa3eKYrJ4GL1z9prWW6+d/TAS4m9qrc
K0slLC63VP94daIDebM48VN8DUxc1JBvBkzroj+cp7vOlK98X8AvkXEVHcRDh4581E/U+q5lE8BJ
rGkWC5XCsfbawPQp0+oeEcXA5SPgCuXYhEYQ3Yk4INYhsyC8wFETXrHijbUUlWKBWKJurFv1kZE9
X4tuJ2AmwdAkcWqeDedMjGcCEbcAWtFsI8CwZf7jTjgVneYu/wBoJDzI1UwuyQOAYNrQjc6lxnhF
7OB8trZ9Gu60DPcJBUELPOq/ANUByK5Pj0rcmg+kMhdYgZR5YVjb93goWC4JAZn3d5fAvvqu24hz
INanYyDKN64/w9B6gB78KUmbfHfevg+d59wLHWcOnyZWBNLh+pebRk5ZccNe2JMwrl3i7RUGc8z4
kJGC1yun9n/fItNJ6wwEDVZ32YW39J4pRIRPKVFkJqH5BQUfcOlPHFLG/1OSFGu4zjV5EdfKeC0Y
56jvQI7mMD7VFghcOpBrdLs7P2s8bQAGwarD7gQlrIY/jQ/R1nQe3jDtVLVLlvj6ngIu3KuIGndS
Ws08aBe6q36yUzRhGLS1fXzqhcHPiVlpAhqcDLbof7d0JqttPshigxy4Ftlzeos+AKVe14jEcLk5
zFFCwjvDJjaR4o5nPHnTYwpG/+mH/tQeoDsP/5ZFJfvCFnmxTVkNTKlMRVXFIJu7+OKFewcv8JhY
9Y2Ad2qJYsOTM/3r+7L2Cg6XREmhk4zZgtlTqD4jGiGt0uwWWQ1DDrOhFtd+ie++Q00k7dA9Db2W
VLHod7QpJ+ClC1yKVHvEbeZ1jA8hwHw9HEJTX8IrEuLPo1aoc7ChgcIpHtaPhXvxg3JvFbmJlONj
XT1hyXRs5NitNpPubWw8Gatr6xgPqMjkbW53IGbHwSzLi2319cKG3qUl+k5pzod8plogXLcwRdFI
91kD9f5MuFRgXy7iohkYJhEH9/HChBUX+VQ6/iHgUtd6X0DBNTRoQUs5l4s1wDjT4NV0F4jVglt1
M5dr4kIvG21fQqUWeUSHPy3cGCoX1Scs2BkKsXo5VPsRHbd09wkL4Taz2erbPG0NzBQc6jEcwCPg
u+yElxqMsyM0pQNI+HuD45kq0T4FX9g+JdKiCu5EAJ0PHVq7P8tiqYthsPopDTwntfIGLCyjp54f
QNu9GStls+IjfI3m7ePqlkvHKVpm0WKekNwwykJRhrkQUGduczy99IvK4HzrHKIWuLZdw6NMjUhT
Nr/lGQZ18ua3lD4FE6H7Y9knqPnUT5HTBy0rzvJZUu6jsguAiwyN4hJKQ7735hFEgA60JMCIJP0w
D7o0Igw8enhrVCthnY5ybxIKguZoswltPdzet/8dZ89JzgiQFvRgu84v8cxXxPy/SC5s3lG6QRj0
HZefMClfpd02IDplY1AgDC571t3hG5mdRC35HCcveX6XuQAinO1jj3lmzX1j2ig89uQTgDt9lrSr
MYhpAFzqxvQmZFiPfQItRdr3/ehY6ZMLDhc9mTI2WROTN+cs4vBJf6pvPC8LE9Lz3TjrWrKJ0Qnb
N29YP/m2BNAhIAKNURaEzW1drkL3+L46zlhPbFTBoAkfEsjIOnN1e4YAnPiWv9clrQQKmdN7XTKi
tYpLpHq00OLirfMuuuirfoM2GQffx95jM9tHJw1rwzpf+YoJ2/H0UfVU+hUuHztsRzF4PG/djlPk
0ZdH8TPuRdP1Cr6p8/gELrpaZKW/Ss1G5p2CuEBX9EzcBB6VG3CTY4onXiVrnOF+fKY2VAH2y2o5
1/3QiCtQgCqTTKN5b3B2JWC3o1WImUlctVjLQS8g00KcZDT7NvQwhL3cs8jgWVc2TiWTF8j+BzM4
gvpfxhmlb2kond26bqDxeh9GL+n0IIzjppmj9k4uWRqxX/2eq9xknzCpDK1su7JDyU1ViDQ7l/pn
dTgGRG4DNakoQxFaJh3wvHn0ZWPKHjy95z83wgb9xUYXPaFm1EwaKKUqa4/ubeYdk6p+To4vqHwB
girAWfsrr7NtFn9JSYVXv/8bz9nDYhdI7eiPrlLv1vb5D/xTy9MjSRonvT7C2pZ408t9mP1GtcIh
XLAh0yhwO1R98BU4ypbVjulbnSxjFVZhF0XLqNwBf5zZxT/68u1+rH1YE6rJ0XADbtHaZTcCzku4
9OEUxMEQrjOp8gm4do2xJ3O577NKqgGtz5h1ftDUZA3x+kfPIbhBiwfUIGjKSUtqVeEHl1oHHvu5
FNXtXgSU0SaAwbDOp9fhIpCqqGYuY5+sZdneFIxGxbHVP03H/QRICAOKaggFjOKRgrjnxsajN4a8
1q1dvaAI0UbaspFkERft4OkBuzitY0v9c1Mjulsfq3FEllhiFJNvHN1iYEiebaEuvsPX1PyLreC/
6Ycec6l1/AquCa/dx4E0miEUdQn+p6hxz7Yb/PDWDSEV24uw+SNhs9n0Hq8OIjPy1HXAcGSnDggm
cxVrc+QbO14Wj6Fo+1wYP0IdecpnDV8uK2FiubI81x5xhDVG654RfqjlaosAU4yoobWhT4Al3Ybd
LDdu9skHiR5mWGGKCJZeSvsgaAzqE7UkvykpO733ngGUMLAf5gj6y212uX+37QAIQwaxhOr5L8Mi
0RewlyXzfSflbYRY3RV5YxUStmUhrjDDYe7qknQCb4KGuyZtFUrxzdtNQRL34KNbrteCExBR4msb
1usc4wVd2tTHPpMaCkKJLo8DVjKVfu3fiEC1TP3q9tTS9/Pp7sBPjKv6kGThL96ni7wYyTbHqG/X
Bpuj5OzbnLtP4HzpcXT+x5y7Y4zWMl0gDWZHqMOOSU7xPEA0ICI7f85aVPy5JDmRvBkX9U8FwRS9
8rZTrIaMZ/5Y3+YFuoKgYJKcpbhBV291nK9p+vQBn13HJjP2B7DYJSabzgatNl2/ylKtDKASQFzr
fgkrYStC4Wn9XiNweLYNO5Y0+3nHN0eGUcQo6pyiAeXPZpuH/+8aiMQ7LowTcB/HA+Bl44PSa0uS
0EMhoLysyBxd1tdrusU6i/3k02MXXdDXGR4vSZ9U5gAhwCd8CRzNCLBPsBm0Ig1//wTuZMlAS61x
W8joeGwEEKcLTWHjG9Erxw2PawP13g1YTlF70O09oFiVMcjb0o7Vd+5UEyRkO6y2ApzLhRDP34XG
DNoCkTktMj8T0cL3VU+EmxnGdyyyhujRDOCw/hFIYGAY71iRZPWRGF24mIrzRp37DJs5s01cPuXs
eO4nUcagrwCRj30vUYySvoMjROG1+nAVulS36cI1WFkAjf7eX5DWjjD3Z9HLGS0DVvmd/cleejTb
ofZIMEdbjh/Xt0/4Zd7aIwTWhXZa7hZZEO9i9oAJyhS0JQBB0xyf/H7zc/NmH6gSqoA4Ia4L6qWj
oGwLPeRl7fjGtdGPV5zcmOpl3TtSZPz7RZpuPcrv8Ui3GH+TYaR2tE79LfOwoOCYNubUQCeL4rQT
czNsYdAUKYdX0m/lfxHz2i3L6x9vcssAtIC7y4Eu7QJ5QZgZHqVlRJcY2SnSMwdgmQ5hks350eN2
6dNniueSD/DPwvhmiBtsa6QQUAZ3A57VS4CPBN5qTEYFZpoBZj9yJIzWQ5gIXINKzcvkst1lW2vu
c141rAWE5EwlBCXJkC9RqN9E7lXiVgcFNDMSoP4x3wObXU2xCmOavIIzFBl0cYNmpbXsvuowqQur
aOOfw/pFQPIO7+2HkE/1WdcvjWg9UMfWrEUSoQoIPFLTqfJvr6TUCRZUFovEutEOVfjCzcQk2w4Z
m6/Al+GPlJ/ywwx6S6Jx6xPbspr5/pF5VC+m6dnYK2ad0R8T1yEyl0E5rged0OuH7d3G2QGFzdEm
RdJKT7vtKxlGggB60TGSwTHR56e92WLsFacpS1+jIoJOTif6+6L5ipqGjfCP2BdlKZqR/+fjtPS/
w+/FbGm2cKz1W6JfZ87SWMvZmG4XsN0oe1ZTYQDXZe0Cl5TcXoLDwk27r3QnZyS+xdqkOlfHqu1+
yLBM2vNFPQ/LJOsfaTT2oGR0kfakP+dLRyvTsKCD1ODauTQc2g9E4u92vKVS1yIyIveNnoCMZvaj
88wn/YeRdbuZN3JayPbqlorNIluNWTD0ZdDcq2x2sUFOUCok90A/HwwEI01zhBEDq8Gue3ffzvCr
morIGDd02YKeQyrxweCJ74L8RJ6T6cvIjbPR3TXqK8KCz+qLl2oLLyt55jxjeclNJ3vLeY2kWSpq
Py8Io5gE2AuwGSbi/XxINKwWPi7MZfhSszwRKnezZP66UXH0YgnO2AVerTGFOTCqlIVQjJamnXLU
HcriTJbwBwbtadXHGDtePBNVZTNPExR1cx8ekDEsyZmin1d3tAcUBbKfLFXnNHub1/yaUN680u2D
gHEPZ8QyCRcKnmJUZvrQDk6MafDTvMqG+hEd1vGSOjffh2+wSqIScq8m2aCRNfH6ppkQ5Fvx/9aI
suC01uDgCdhXxLRCOim0cX5uhBqG+xPcl7w73ZvNvCA6+75E+njl+bHtLJqOxjtLL4C/IHuS35FO
qBYf1cnfYRLUaumZ+tQXhVAwIX8HlCmvnWQtMMfN8sQuvA/ih3gpr1HOmE3izgWFaKGJaw/oxbwR
eesKX4vK3eHR2aopvYyruGPxQKJUMl9hp/2rahXoMLdfOPTY9gCyuuogW2jHwkM1WlWDZZffwp8/
fgXMpfKIRsuEEmU4aKPDFAkJBQnJbk+w0foypm3nwkb2t54lccslQHW/2D8tOlqAhGH2aovCdY4d
AK82hYO8A4wH8v0LmyYEqNhnrwU7H5AcL5NUAtzyX6+HEn/xRO06pIRABLdQ9ekTCzWkhpo4r+Cc
lYQiLdoz8i1+3+pUEqTEU6qoy9J1lH+5NJOeVQAQMwHXdFdEXoDR3Likx9mHQRxvLC5UifrGkBf0
wnLmKTMoKzLjVe4hp0Ddznae3B7BOZySLPOuqnoYrDLYhxWNC4hkvmvti0QnNyO0hmvBm7iMnFdL
TzwPrdnpAdxJiojclD3IUcr/sC5aprRLEXbK2m43J8mfqWKE/qIRMcci92ssc+nKP8QU65bK6SZi
P6UgH7K7SCRgjo2ZvR10yYEMeeIeNOtpyMViss8EVS0AXg+1yavmxxLS1YFhoasiHFZEeRce56c5
0ASzVT2Fq3MPQvvSN9oUTbI7lyxHJw8j4UvNSXvsy7HmMXTNwpDGnIaV/xJRXg/vynLBXNjPQzFq
RW2idaXJaVpWZ7LIO8k0g1pTADDTmP5dCnHiHcwft1cCkrtsFpmjuVHujJ3+V4+G6n6AhU5BNHQ+
ki4sT4v0s3QlhUfWK9E3G/P/PPej8lPuwnN/F2AigvKapZKgXW9zT9etceLnZ50NjPZSAVSR671H
g5gMyfD2cibwD6cZKjgaxiUmIMzDvhvpo0E+U0saldP5J7I/IpsN44YPaZnW2Iau2Q6FRaTFodaZ
gGiI6CsL6b3vygZYIOHkHHLDZK7xflSm4JaYGQ5bXj6QXun5hpT0jKeCfCatqMs6xSWhDqeFbC4i
OLHtoI7umKs4UFqEFZg0NNhZv5jT15Xk1QoOCgPDJqnCXVim7Wo4Y4aZcFfbCUbLIfQkkRZefeqI
9Ykrk0wDk9vuIpUwtL061GODUzScYo+DDD/0H22BW/W6VTlb5ynY8zBb2rhr/dFnHClhes9dbm8g
5vynborX39Xii/5sl1TEXkyGcAQgngXMePLZQ1TgKAtTt5cU4pNDcB7pCzMb22KOxeVVkelzoCbo
srK0vLjHZlL/6nQ4090h9Cp8lQG4ZHqi4AYbZdW6Pd3iKGXDom/YHhfb9f5nNrbpGx/yjaTx+zWb
xWG5Y2a5fpruHE6FCtHmhMUd52mlt3ZRxNII8sBy9f7oHfhkCUFz+Fq4TYsqItDxYel9zMHRZlui
ac64RMf96cJEhvxOJ/NkTsVIGkDla3f5OfHavmpRGDcRTzyESXymauwdV8uJHfZ5mBGIQdiMzqdJ
rn0dSRY9A0zpUaFmwyXJpeiGGWFbyRNwN4aIWYIbZbexXFCoCxdS9iw5vnhRVJY0wLO1rq4MrqNl
rzNXvt0IYDba224OYh0jp9ml9eN1Hzdl8CzzGNekFgCxS6uk/LkSUNv7V4+RddZCrLtIiPyITnlE
NZ6Qbac1BpMnDibTgHI02tmIq1HVwgaHe0GyjK2CIPitDf8j9DgaZobdWUbzoKJtIi4UcML+eMqk
HSFS0+f69ix+eNw/X2Y9oW9qYltm32XdZhMD/uuupRgizt9RDh+FF8St1ZpNAyL32PltGGKGF1Qw
oGF11e7yW2Hp3HD5HOchO77JuPCw/BqM2yPEoClx6BOXw8FMv8DGo8Z4xmPybOcZIt4sCh0kO00f
JotFXETZjijw9AO8nz0TOT9PncqDbLinagE5WfKFBnX7fw6JBWJ8XQ9QijKhy/Pcvjki3it9MYgx
tH4YOsg+r11JbSjD7aLN8FuyR5vBXXp9dXVeFOOYXDScf2QFHjMaglJc4TCfunTi0Zh7V4rNSyso
+Sw9oHTACjLCZIUm2mKW6QzRT1EvtYD8N3bj9o2C8ssz3W5UMraOJmV8Dz9X6nEzSz2gzduQRZEh
ARmCV+cp1XAiDYEoj/pUak7frNSzdeq0z4EvzTUqjMxzsxkEY2FJu12IPrC84Ehaq3ayb4E+byUk
zuqX3jpPxPNwxSVx2Kik+DtUpAPh9xAWmgDC1nJ4nQ4TvR4WsPmHCTUf1oEZpc+mdK2lnBXO5a3Y
6SdV6d8Z+kYmJ0osqJx/l33oClSuzHKAMExUsqmPexod8Ql3lOF8I4QavpbhEtH9Du3XDEB+oJDA
9Tt2pfF8t1H7o35us1PDYlXwYCTHxtApfwb3VTaiGpiEfKcrlbdVO6UxQloOZl+ZmMi50bZjZAJ2
dTTxTDN/gdHftATye29kl9j94A4MqxB4aEeEf1SIkTtXLwatFlrRQiQjzGJ3jrXo70J2UCLO8Wbn
3OsdkrD/++GKj3ng+CYtjVXHEg2SSdyUcLNwSjf6lhBofaf/0KGJbDa0KaZdvt+JOUEZf3+bjFrW
IyXhKYQZGLdR5DxE0fDW+0qwTJjPa8/7Fxq6qNSguuueY9opAwm24EOx79KepvVUqkBK5Gybfrfy
uni9stE/WG2C6AnxYnDWv8IgoydMO7pZE6tS2/Ja/ZbEROcThZ58zG73nivjiPM6fDiYzfP/jWuM
DLFbpzpmUgvt9tgKa19oJKz3xkCKbXkQfJTQ10MdMgj/EPp3dhhKJGJ5y+ufGovdIhHa6bojIEGP
FsXInLGwg7x3E+CyOZYannzCtqmsCrfO+jY2Ic7I9mTacSR+FUiDeLD4ms/a5v7sp2FYztRM+SMO
vGrLAJa1U/+SyOhn5oQpOA8o+r3+FM2cjzXEBbQatqQPrTyzrE7IX9EiOg6K9mOLsPInxHYfhxwr
HETimNCezB3YBEVH6cDxPPGW9fQ+IgVWFYdjQqmN6QePkFw+2C9EwweNLF7Tg51H1u/WDbudDjmA
RoIvVB9djUnoVBY32TJ6QGyZGidYngryu+S+0q2FXogEQgfpl7RUk6zV3jsK1QjFgaXwXljovlU6
MNQqoc9jEQMTZ/8CvwGL84i5Uj/RgyEJlf0AKGclUqB/6dBDraOgByiLxiVmkxVjbqHkEV965x4K
cdklcHV6sDqbgp6saBLng5Bx4lbK2E3ecadsrtt2ab1IQpf5LkFSPkOe90pKJ1xi/QSWKIpbcHqv
5TciTTC+VDLjuJrKkLAc0aRh9wYIaC66kRXLW9Se3a3bhkr+4Y3pv6LAoQcRAweH7zVipm0UlL3H
S+mD2sgOsETQugLriVowCNkDPMkEErSjaumm9SwC4ADCfaTGjIe+0tDUK8qcYLrJzqspp+mMYdhT
74sDR8cW1PV1/MCfy6yhetDDgrvxQzXbXLMXViaGZx7IChSwK6cXVnwBCw1h/vi+8bVvvPgwyrQR
rc5mgEt4/dWoPMFWEf3WLPZi78hixGfucx/DWtWQzRiZ5vk5MBCnza02JuL0pqCk5vJN2z6pvRAB
aoZopCcft3aJcQLRJoWYjwh3/867fCtqwfbk7zbizdVspxoJnBcTwQ0ikhbDkJ1XYqtcuboQnxlQ
iyB0g8qoCm4NZsShaDvc73xbScc1vEhpYXXhhoifExW1SXTebuWRzK55wVT7v6BW1nYO6fdmENzO
b7fS3mQsi2qK8+UdQH4t2onnn/HG0YgfAVebgu9KVOExK3pID4v1w2SnBicxLjCFBZ+EOYnmYI7T
pdrHJIU8aEMEY64/vfTbhwhanPpgl8u9Nfmfq80hRImoIJ0tkHJI5LnuHwQm2Z7NLYrPqwPdjJQn
dsQZvZSkAvK8ZIzeHOxQpSGf+BU85qxIyunEQVJ7rqJtZsLr2WOmh/EAw3O8vdlNh3qUaLhRm4ZK
rlxyE6GIDLKZPKZngDRAzXWelJyBTGaXRsRGVDEA9/8aGIQByeI0D64XuBnpzXteuGz1sbH3wCYw
mEn/Cg/MsHG6/MzMe4EbBGWXeg4gdhGl32lZIIEzVCW+D8keZ9484j8Wiin2l9N3S6a8Z0bJudqn
Hm/i2R3MrqAxfgBe3GYb1A/aMOozwCMzyPlQrW6GfcZ0JNzJyvp5keISfOMvC1cKsZd304EJOSRl
jl8sL3R0COr+6m3hzyIeI1X2goZolQPhIhsN+G2hKB581NySDvjzFy0NLGAWErjSjSmLK+Ae9PY/
8Y83xjku9UAVwzzdodY4TX2juNZn2OGvCeGX9u5X5AwOg6Anrmqayer4Qm773lgyokEtIv44v6WO
7BJLcBFVGbQQQO6RACRPQ/lsbJKquDgFKyjMCRTtGQZQo5YQPom4S7cpekgdmBMYNPHPFT/xIBx6
RqrjOEeX0G4Nfa19Ht8hkfL9CcWMepSWc98O5wBw32ERYAY+5KrCEbT2RY46jbtF9XEGKZbRzPJG
/TAUdQZCAWh+BNdUMF0eXWdDKuruAzPfcbnlOasfeGsYPxG9fI0R5yYqPS4L9qVFexMheuOW2MyP
yNMDo2rWpS/cCaDn5BJ6L+a5AwYrPAN0XUPm0N403n+Ct8gCGVhcLxaM1DJ0ZaxI71yqOdYfM3No
1NKXk22mjvxsCeJ3gdJP/kLYzVw9hltvwmLqXKm7/htLad5SAe97BcxTnMPQZZwDSBzocpIWHEQQ
T/h0s1yDCmYDsIJn7RAwu6KxLyo0FcvLwgZMX25172fImR6q5P7dfZyPiL/uEjRUTDh7ENJlpFJb
tIIYSWvoUYZ0Lf6NpxF2hDc6sIQSi7AUxiy5ozgXdVnONeXK7ZiPOieIYPz4d21kyACC5lyDgWyr
tk0H4dfDVEL50uiOTFtbR+aWwl5CJJ+puzZ0qdzKaK+nD1/fk8uA0MwDurc0qSgj3K/HyPXikQWh
K6L7y1eui4YPDb+CcbAp0lwqUu9EbeDCbk1Ns1TVribH3J27ntzzZqz7UI2pcUi8srDnq/G/6SDj
7Oku51yvVMv1Z/jhrFh1+fvBU3uF65i30Ctpe9uco2wdqMRVi5xEKWYwsHH2Oa5/DHt5S4iOaT88
SYbvGwUkjgj53Jf07uLfx7t/BgxxWsbBLhrcCULN12oQO8K6Bd2+1fhzaymgeTZXK5FE4+49sgmx
HZetEOQhHg6eJB+6F00dBqZ/3JigvjQlimws4BkGOyp/j7sB/XP9geP6cbZ2pOc5gN2yj9kz0REE
3GDtEMHM3Z3KCrHlmyQNE9mTCexpx1Y+c1DB0qP0lKDHt8+5vkep+9anW2IsXzAaROSaFEm6RDJ2
nZKxQDMN1CsTrih1D6qSQzY3k29FwqEfVufpeZHP+2x7wW+mq1lUKtRGETCCNHTtM91TfzQe9DpK
j4ka9N3cQhrYJy4R/uWXObigeVWUymVBee5yREId1F0Yb73ci7Vg40Bo+vUlkvW6PdbYBaxflBKk
Ym6O80GhBvVXzhEUB45wZjxt9sXz/cSCx1mlMAq5L9k6Ksy4qJZQ7TTp1QnlW7oLI9y62AnFTozT
F1THc/R2BuEiVTN9ZUMMp3a9VYW2PI5rd9Am7fTFwId6Az87H34Bg94fzWSJ3hrtfJ76LPI238hb
lqQzuUtvJCwnJUluBcSXsMGJNSsdjvpPQMWOah2sZ115LTZn37S1PZK0Ai60uNr86i9wyylHMAnb
aQ2M6u+D+nxhdeI/y5oWoQDu02zKx7x6gUEhDozrhZ7dXvhYQMWofr9gek3sbylFw8QiLCiSjWUT
F8WD5SP4JWIt6BijpQbj2j7s1PZT7TP+VNil2vFfPYaxrejIQYjMUPGTUn/HzuaPJyKgo5P5nm+R
daj39cYMOK0erOO/Y4LKxqKgPiijYXSEp20ckjo5qL7FWIAWOuVoxLEPKGXwRI41ox/V+Igrm3Et
Zle4h4fTIVisdt4EoxTnPRzYBUNiTGStI2Mzavfvy5nxKzTCUGbQ9uRiqaqGQY+jjg9JoG9LXQYU
zD181b3+7nfBnDCZpEmjh6hw4mTiA7RO2AZGYNuXhoD9fT0GDqVOsphpKylwu8h3ucVcErMU8vhm
KcqpusQRG7ULvnGPWpqvc9Mkz/LY469ibsR3DuASxTepQ/pJG3NUxvtqRfAvAM1rhT2l4065IopL
NF55w6hWzgoj2rMBYhliCStEUTCtH9UGYLgcfLG813gvaLDbbBgfWcjaP1fSOYB6BGZN14uig68l
YNZ3jZrTFnh4A/k9aE7gub5W6hJ4iu8tRRUs7HvdszoJOfWMEpkYdGX1px3LRqlJmYnK2Mj+6XGS
Oy/LdA/NAzaQ9a1GTxaxYTXBMYCud02gbnQE5zwxbc5dHTf6rxfKtlLQxugxl6sFOJDME9A3CqrG
F1uyuc8USs3VEcnRSIehkxUcStFK9TuHQLYwtRRnkdAScuKpqIkbHbCjg5RTd77LMQJOjxvOEMuB
EJ364qylezx31wdocfGsOPaZJ4kNMvGStfCPvtCARNf0McZifeH2BDx7As65JBhPShCgeVx/Re5W
H5Us7SwVTZ3Vgw9ObuQlg77vSYEnCfDAmIgVj12mmgPPYY3sYVmtm4uQiXfudBkwJswVRdC9X6gq
G/0D67430hX/DII6mXj4jK2m/RuuBcyuhmbAnxaQh1mWqKi8ga3fga9XJCvzUq3ZjOUqYho5Escw
N6bu561hVrSc9RHgofRtf5lBT0LmUP00yllxqxHEUycHyRCiGBwebHYVORXofGqaSvsducuidQUL
fBY9/X4iLooyx659luZ635qha4FlK/VbGFzw0B1vn+kYEEfA5s8Tj3GGMerPhMat9+M353a8lFok
xY1SKsG8JBVQAiRuQ5XB9FU1E9Qm+7Ri9Sc5g0VwlvlIIK6DXcSJfjwNNmnAFxlgOYL5Nwvo0pxg
LriGVOKhU6zVoz29jeJwa8tZVSSBkXJXX5RybzQnpqij3yWZYT2Jx2BYQFmgSPw22TrBjzq7zQkV
pKCqJXOYyjeONVkTITzCtUhgai6Od0DriqO8Nj0Cb3iw5UB8bPFckKKDrlhn1bwjrrgPbWY0idB6
AMrnFjzWvdkh7Fkkok9XgiyaCRXSIqQOx2j7R7k+EgJ8R8hK7vWcEMBCm64JLKmyykfRgVNdXdOn
/H1FpWo6+3xw2QeqAt8HfhCgszq27BIJSaFkGwAedQZXLCoVDs4UvI3GsWFm/yx3iQPvF014Xvye
FxLgCLWc9cFMONZc3urZQtkX02PzxfTYJ/LoBmgLxQEHiulcg6iRtOyNCgLqeJF7yUwI0rkVdu6U
1MaZwoAFL25CBtxi4ezF9yZoya9gRNn5hUr8+A396E/Maf3J2yze3wtt2KAQatw0Hl+A0lS8wO7t
uF5yajEh40DgOR+HdDsq13NY+RkbCk/rQfocaZwcKweVLBnpuVx5lML+vwpZrMd7VkZo9sT1NgjT
dJgCZXjoVbKEfWG3lR0eQIyK3ubbgpc3ss2P5LwHfbxplurygCCjTe6WrrDAzc5HGr3i1Y5W0IZC
v0Y5FKpcf5GgoL18CyivG3FlQfMp90vUiF6ZN4/OaXbt2aPI+yM7MUxauLXTSkwdqCGmyP/v+xdz
0hxe3fz0xcjEd+QIVMhVdc5uV8ZegiN5dtFITSib/mXa4KitPbOnz82j6aKd1vLnFU+5BJqOTm1B
+3LUGrLGogJ+lbKTeE9S+QpgGri4dJoUaBN4kz5h5/kJHC/XlUDQT+IS7y6nC5+LbdAiBoIInnxj
dbV+QbKzUwcCWCCarsesgfkBfq3lDEN9rfB2hWvE6UNrOODLp/HTwFWBSaDyA9ffit9CgY8PsCJb
8RBO4sb+qIU2DeZL4lAhTvbKL0uUr8IofHv6R9PSXVW8dcmpdPY44vExS6BZ8NI7a1v3ES6kvpXd
ERRxA0b8TPbFveYwXcQgILUNnyC3qVLvqB3lNHDY5MUPHZ3U/OtgBaHKfWspQV1r7DE00PvcqlxA
wINz4KdaoQX8JKPFceekKVyRpx+5deQ+Fek1b0DoZXIknfyawKh7p6VsPx6Nzqms+AgoA28KSpYt
jL5vi8xRSKWaLzO6wflxjIGcEl3s1dgu4RtkY0JignIjBxMSv9NHX9kyyzukz8fyIbffK8vfEyKT
9RHlYprf4kJG8cXKfzJblBCD3Hez/KTX69PMWULzm3zy+T8LAX85yehZ/Wj3DRWCnsEPMF6uFUtZ
qUnojCyEJ+jXOmr59Cmf30oJvwmNr0FrAcVRq5Zsgo6RHcf2xixi7Wsyw1ddLudpZtmsli11ACGK
IFU76w8QQ46tst2m24DPAr8gARyOHbKg46VBQoNbLTTA7HGbbLuScMmoMkoWd15N3o/rnGHDlcil
AgR1GBHUdETRENYA4iis5A0fEpH+VfBzeRIOQ+45eWBMgi83YmwomPyOhLK8S+vWerEmS+GzNoa0
7/xMVsza7kHA9q8/78LbnPODLWFLQGmUrplaevM/zRSxZ4zpzJzchEso3nhNdIMg0VDernBdKZuI
a/n7SZ/Wg38T3gTlsIUl6O1FcSf7hqj8FMcy0ZGNnpk6Mbc7KPmSQhkfTJlkhg6P+sCweY+P+w1+
P/QSAD0in8+VWccKhGh/uSyE+Db29FfawWFIIKA9bcjNfKeplc/xCHGnrHmGV9ySYC9NPDlJ2nyA
F++jYak9oCCsvxNu+SZWh+Kz1CXJhrr/Z8I330kQb8exNAjfGUySlg0J1+wizTRG9FJMck4qbLDO
biV2Kq4F87aTspYszCCivX2r3Upz4FL5LLfAS0Oki7ezXDskop1MDbCngo+HDd7Y+iPtK4nGCWEH
rDphrS46adkqQtZo8/OvfD2H2JR8tmxM3jipVrpKAm5r2uzqhZELTmFMVWxYXuv5oXO5xf6TGp6T
pNg7TgwJT+SDgK7ucW5orO4Koqy0EUIk8yT2Y8hHuo5XBItbJy2GV9R+sWbKGouHzICUEGGdDYA7
5NNNqiXysnY5ngZSAGqY0IHpxqnatQ78gGGCTW9AdbRrHZGg5zr1FTwgwOgHSm6w1/tqb3Ft9zFv
bhEdtX2oeyQdUkkfeYofXojxgfraEbJaGE8NIyqHEvoffsFFZSN/lj43Mm6pEbAmqcdiMNNQ1tir
U+6+cq2I9sr1y4bKtJutcvTpifALNHsoLS6JJClAvZaTGfbbKPfalUAK/IWWIcQ+fizEumfh7QTK
EeMPWybqKkmY+ydODjig+AtjmRYbS+P+l0r3N3wZlb/hkdbvcs+Io61Ee5hZvRPoFcRY72jxi+hu
INF9xykEWfkH9O742tjWthpTLdoIA7xuETjijjuHuhUIzwqN5sUL+Yef3lCRH1tJJP3Mk6BPmbO/
7z0aXdfTZgCFvs09Zv7Sw4zhnVbnLFS99Avj4qV5BLNSGaHnql2ubfTjQS8GFfvllA2kWGXCpCZg
Z7o7rRXxbs0Pr1y/w0usK/CBaQ9XYKC7FidAemD3dWr7+dTcCS7DFwyv8ixUn0pSj3P/MHlsuxXC
zjzCJVwtZzGsCAL2dKu1oNwNiBISJwqGCHL4/Ie798tkphIubcc7JbbodI+KP8ocwa4n+lHr8W/u
awmRv5x2tPKdIUnUPJAZx0Ayrk/jeoSZYgWReVP9oMSAimpB3ZTLS+U3yJCkSZRa+IDOanAmnJvS
ItRex1Sqt1blqwGN+gcUfPqkl35ngcYmHfiBmT+dut+myTvVpbNq/JvySUCHO3MzojW7Omz/UzbN
haBiP025cPHYk142RHEMhFGFLkb0U4aK2rbosilQh4uQQsMm+/K67+fmAF2bWfIPco5u9N09bgpH
AEOB5E9pwCSj9UcNZqrct9sxwyKXAcu1zT1HarX3UOOgXAYgYk4NffYagvupTZSK2jT9HzInrD9H
ekW4/3vPONZftNdAGrn9LEJ6Fwuwhm7dhJ2i9wp9j2Ek5awVJNSM3FaTvx3cTnvDLlW5mSpBMeY5
FdC30phQ5OKx6JeaF5myxUwuCHN4VUTnagMiVsF2PgDhKYe4ufpSFxy2qLc2a4a9kALmWCxtS4Un
CbC+6Cv9j3Rws1+LMMYLNSmboLChYY9u+gnayJe6MDnuKKXWmas/a1ikUNxUYwFidAw/GiOJO3iy
KdwQdWG0aHvXWU7yESaWfidbSMT4aQPjUU69x2ZXspuYWzskLkrYcnb9icjsQLz1fJ5aQzjE/s95
tDpqHcyNUTlc/g+vHsGf9O31LuWWbo7bKqYfxEAWawE54JZl4jrCcW3Ts+DwWyL4ahD1Vb4Tvb/t
KSpDpyLTI4BrYUoY18PsOtTOr7V4KbHnnhB2K/Uizo6444CnxVGROdqU5Wop+xrmFjbu7bPPdYYS
UpcYQuZsYvBMLKQZhw3T9CUrJbrzMrIxnWPgw+S4Gl7IXcYuAwu1qQXgQRcELuBeua2NYlnxDeQ+
Jm5kdx5aXQ7eOiuJ475mWGoIRWJNAummUTWWXJMp3g8MNhMMpV7ouawF7pv7QcQv4Z4Kmmqu3x0c
c+vQCz3Tihru/+2JWVrHyFfxFmbc9SobcgM8Umt7U5uEA+kNxi61EZdKqnpma/d7VRnp8VdPPZTP
Q9pQwIXzG2hdyPnu0EJEZJWpOMk7F6AGesAL9ovw/pQ3HOD+uSggZtvIFd9k63645g/IWVjPBTPY
geT/oFWvD2XstlYHq+2wXInNOWCrbmdHve1ebiRw+4K/p6F66EbBIeYqb8RwkREvgpyrl9UWxfug
QZ5bmO613Aiqh9xjouDArhm60zA7bnsCDrHU+MTMpK1kZ34aSLlAoIjuRA51ykMVKdLeABB9x1/r
rELuVQq7NtdnYJ2dvhxpfkURSzT6PSNfTS6J2Ox53k2teXZMoWpELNzakp9ltjVXSAjYhqfA0QOW
raYparp1FsvFvbGaPZcnj1M1yTcjZXLNOSLMn+tMh+YAuDcfrfiYQULFA/DtjCAMo/0Xq8KheGrP
WvfpEy9joINl6a6A64QpxtkiszUAtOtXlGK1h1QSQZexc2sVwiBAd3HCxYfqmBt3Pof3hSzvRRfN
huHD7fgzlhoG8irJhZkvC3WvSLVSSVodOyRi8JJfv/0GWhTP8g84HsRrZ6gMOObC8s9h41fHru/Q
DeMXHyFqqftidCe1SwgkKB8cXtmMOMzLN2ucapCUM5llg6sninZEiAyrmwUDoF9LkxDODhKAlxZt
nzirGqLLcwWxnLQoZRHX1b96y6afWBr005ILaCOYPTsk2BYB8IHyGZ9qKp4+lYEjPyX61hQqC01h
cyY0PlB0b1aKenY1+d9/DVmvgwIA/YArKamUgUZV4OVuARi3rJ/3C2jTUa31BYE2yG8pslbUDBPb
fLxaNR8I7qhRUxnyoqcEssl/5MomIcSPD1UEDt1sXHq/0xjiv/8TLAOphRz0KgMPyAgJ5p4PyBha
6MkHmmhq/B/aN42qmRRix6jC5M5oo0djYPNA2ZLA9+if/EM021SBAM4+Cskn7oG3Aa+TcIcCF13T
m0LkXlbV4KL+Kixtd6mgmoCxNvKVxe2rOmPHeCtFRdR86g1WM0UoILVLSnYDUK6IeKv0yO0Jk7s2
64St/DKloPc0DOz1bpLSZRSxPpgG/bNUPX6Tv6jgwnyzHB2UlNC0b3Yfa/JnSDEz6H/UcSDLeH1p
CtF8/gzVRxiQcjVan90mZdozmChpqW8jvIx2U7p3KxfGJwCUYB+Z+PRvoGgMsLMotXeQzw/MsVCV
drYsAFIOBweAfSNc+Nd5evQZgwjuEPRIXkyflJejF+vpThVwkis8A53MBCsqVfuiYq6udi8VVpm1
pr5ME0botH7WmhNmdWm6Rk4/N8SnLD7HWYpRQ3d8F4+E+gZhWcnzcGvgcFALak6k7CCJ1a0g9Vl/
+0zNb+0hoywRBj754Dqx2s+xrrdHdfhdh5xExpENVxe116EhMnrurQFbwNU+klH76zjvObrbrgyW
ipzsWdq2rz+pwX+hY4YWy2gYKoBsqNYS9ijchw6Z0EIVqI9R7Ekl0p8X75ioxzVdwSF/7HBTh+KY
tFeN0xuomBeRFdNRMQWxM9WzY4n7DXAAQVClE2XfCEOS+aGIAN20OiO3Md4tQtywmninkhE4bSad
m68wGVFFpy3fSLKlkNOczj6gVfs/oKkc4zBK49/SEa2A2tmaTUs8bluKZM27D03knItZmCew5BB0
iCYN4/pq5R7kQ5sZj8KrVuPzKKGTgfBVO0UrXToGaTZFORGzQBeV4xHlju1MHP5VICqPvELq8Wcd
CApA9wXomr1pWHPOepXhWnmfTUOmYnfPZtz21QnmVaZki2knH0rWV5YcdRF336GUnwFtfZSlatUA
8e5BZd25OujCUphq8kEJAGkNYQwEvVdBHqbeTRoBCq164oE+lgAeYM2Cz8Ai7fL77KYOE1LdUOVr
nwEgaCw+H91EiRqS/2Y177HKZS3/HRnhljDu/WR4UqOl0VTDxsslQlG47D0WsWi+fVUKcH4Ne3KU
IgVZIl9kl+9ktDeejDl8bua4dVVU1v/j3mT+RjZTBNvBsTDuj2MFiBC1nVczQFt8lCSQI5tuSmIg
S/hYPI+U0XxLFvTQhxqnSKfhmG9cNKcAoNQBunnzViSmOHFU/4KYcArVCo0fEAt993bjXBaAEuHd
tEb4HMF/qy4sFtNGdJNkVkOG613jlj8iobDjUkAoyB4KsYrxZ6SruDmwdKNCUX0NVuvZJb6ETIax
azshKI78UIdjDKwUk33AsKyFZ56FlOh208MJ1eOBAYLGR+1Zt9J+QoeYveC8pv0sTbzWXQ5U54N9
88HQfB1uCvI0OkiSHDfcbAeOGGyKg2winISXKarHPq01b9ruS08s92rjy7FdzjG7Ygmb0VE0/ICh
TE/Pbo1VntUaubOd4LqSGSfVxPTuVofaylcFJ9ME6Xa6rt4g6K0Uuj/fPs3kun/KYAuy/rV8bkva
6J5JgdEH/45zk5UwmROXHfhXPdWy5ZJ+O8eccp0Pyi18HgsOX58GqQF5VdjZcagaqT5M1vMcssoQ
iJLbmNsqoTju6Z9fqleLJK1bsJc2rZuUdCYn+O54cm06Ci8vmxSvMBb4bYMsqsnH0fzPUP4WvWWI
2RAKy4IpcEeemtvL4xPI5VfTtV3Kp1ZHyxM+lbids20w0/WCkoS33G4evlB8KWD990nbMenAXTU1
wYwsHzq1vPmJgZUttO7W3vZAYc2+ZK3B9HkDfEBd2PfDOr5Qb1Uj/NgoSgCSvMwYrkEWSoNmTNtG
SJpCR7YG9Q4AhxCXyV+z6atZb/Vv1LvciWStwKaC8ioWxhKBHE3HA1HIbnxWvzhp9b/+Ejt/dkmN
ZgDlNwWXrGHQPD34h8lzzD6YrUICEZyGbQA/a/4CnXaqrCX1acJE+qa8+C/mOhYqN0+uyjrAMgHu
Q6QbWZ4rmmDr3wuK5kg0pJALnlTRCSSs4Ebbcvar9p6HEAQy08rLGP8SvFEZlqewoEjhllD7Fe7h
5Db+DhsWjm6Aj/ywJgdmAOcr+TBdVfGUXh5UKpmdJ1vzW9b7wag9AZ0cYlL8PQmpU7HNa7uJub5W
oDiFlhfN/wESMhWjqViMSgqivgvysuTSW35/xPyyvjzeSUHxfP+XrRibbPtqMcec5VPvT6eRPRTV
GE2yt8/myvOKcMu9id+7gUPpKRfjy66/Hc2JZycvUz5gYIkeUa5bk9A2gcc9zoF0+Ty0NGsM1mZH
hidbyEpaCoXlYpWddaOdPUQGQhpE+Co+/lfjCUomeVISjBIvNJPVIIQjXqE2Mc8wO39juAiDxGOu
31X7/k0KUhF+hm2q49S+XPP18Xt7t8NsTZOMixOOcVpVH+hudNfQzwmiUWNydg2VyNxTBZQKQcbW
xrb0tVQsBD0Y90UispXgH7t0FK9valVevaeVHehTrY9A2dxz5BiQQJH7JBou3h5Kp3Ic9z2Dnc9M
f7559nGo0y5XAB5A4qjpQiB+50IB3ul0+pQxyyFAl5TXxwdq8yul6V1fhXttG65t59al79Xm/0YX
7R4Rt1APwKfahRcSJYmOzp5m6Ms4gBDBlmwOqPWnIQsYHeHU9Fduv/DpEXNwqvC78ZTyIfMyNBPN
FDGmwUytuLU69rGKRtUUpmPU1wOBaBCoUjqz8e/poQJiwCOG7j9ey0KR8jdhgKaEZxbWQgDiRAus
wmReZJV7AZqKunXmyb4z8vC3lDw+JbZoSr3H4vxG8LWFuHap4NVZt8TOqy5xnhdzyEB+d+IMc1Sk
QESdXVxKMFBu611rUXv0TosXGcg9jQ4dJJ/fhPCl+6cx3eDAgFTZ/2pXUohowBAps/GVAoYouE4/
ZJz0hAhor4sQkpVxqm2ZwMzU5oPB1TJZ8Sy3nHWDKTuLUiateeELIfMmLNyS7XPRTMPf/juzh85Q
vugfiClXcxDKS4qA5Asffpk++tUFEcw2qSQAoTLS2Y3tctKz3sGVMgbm9S/+WtmSRbyzivGEVSbm
GrWB6YMFL70vWjWKRtks6hmVi8zA2Jx5aosTEDRMZKZiowCmHZfoeCuWTkEt3z8G/2ZTWFCOTXVV
Q/3AA2G2qYfPhWmPX8rS0/8oguJuspdovhs+LM7gufblSC2YHCvTGnhIaoD9GIagxN8AJacwaT5x
gOJbngW9Ts+Id6RKgLR70GbmAhsRFL3GMg9S/0N8nIINKZeoCKcLsuSwrWHYC/63B91L+MjZWDhI
ItMDYm5zXp2bBYWjw5ZaVnqOS7zDcsRONEOQkwIHZUC97zDBrW04kVOYKn4zTYzde7v5tu5pHDnH
Lg+NA19NIFDG1N2iaWzGsT7AsPfNyJVRrGemtFccjmAkiy+wfu76AcyDmDkCiP7oiWBuC7nSmC/4
RwQqDTOumPvfzDsF5IWqPr6dLCt+33gIuzkE4n7VJTZNshoKwgU7WlUwMq2/H/8tb7f1L/XI2EDJ
enQOKgrGbroCdNBuvnBeQraLTfAJGg+LlP/zFi/BmDn3UPzCn4C/vzQOfWFp/TnIr9+tORlqxkUo
SWFtq231KdmkdaWf5aILB41XWbWuC6e81K+liYZkEmZHy+VrTq+KRXJvVXVb3QBFK+hoYLXKiEBX
GV9pnxsku4Q9bDrduVzFdZqdS8TE3m29sg4HzBaJEg0ctwOeupNn/1yoEzqiR46hbFzpMrSs7FW0
pgpxmFGxn/Bac9gfR6XgLQ/C23GB9ENW/QN/akQhfIZhuMr9elUncWErBHJnOxzXizOEC0bKtcfL
oKXhknd92QdS7Fdop8DcapmoyR1u/tVPJFny16JnlHC6Y1MjKoKnsNK53I6AGZNqYILp/Y7zCxjt
k8H1ms5pI8s2TwfhjhNB+ZEsA89ZkOc4ZPUjS4KPTz1iYLHDBTKkurOMeNTfDMBEaESRWId2+TWc
Dcw8HJQbOID1x0zYiJVd9H/byVeNrc27D8e5cTmLbjJjmqKHRZJradIdtQu3bQ9nross04Icyfoq
0za/KNnNF8EtEvGHu1xi9/FylRvUee6KpILoP/ZlnwdQUqkzjRrCDrJzPPPJg3bLrj670TpbAFI/
TpnGyhD4okgvCJVbDp+enTwQZ5vnB/4nogGU9lwoPm2QL/dlUh8b+UeP3sfgM9QXgbxNk6pje9Ve
4k524JsChu68smCi7nI95Hi3x1QDEWE7FSKzFLIfnGHuwHlJf1d2UKK4RGzgx1yA59Ot52Ds0axM
045Qdl2lvDgQRI53u9X+MeQrbDHwsFRoBrxYQN+3KF/Y3326YNPgmmsFwvnv7ltrmS7RvUQ4fy9C
qf5hw3+BIZvQAEvJT6NHtFBeg/jNTt2OfoYGG+li/97PnYslDOC+Gnns43oSLmMTXVcgX2CpmkMp
FYGpZGRVQzGNBEeUUv/PnKyr8OVbppxhuvg9bEOD6WMpRFkR/VSFqR/SkbAeCmuwufmlF7UpKN+J
ec0i88K8vA39ZLPezOQHSxJwng/CMpOeGCD2CzyIrDdxj3W2xj8rBeSDkg0ooEf9a4LvMAO/ag/V
PnR8Dv+vUTisOM5GbpEXNi6Nf9Gnk8ad+nmuhcXvXoEv9iztRnoDNHoTNRnX13YyxOdOsPGi+h50
WeFQoIQ77psL9YAJf2e6gZqOuykT3Y1OFAQuKKMoC0/cFWC9QICh0oEUYzyNHrkw6BPM+GnNPCsO
RIh4jifmXuEmINHad5TrPH16Oah6puElWGu185fY7YZ086NK0lT1qh+xfvYGCUMfRvS0t2aPuZY9
wGwhU9RCE3fQvbwxkgG6+UUsdk+ZpjWLFYnk3MMM+4cqBBFmuQRcamJNBUu1tENvrshjL7sHEzMt
YmM7rquI8lEkwfd2dZtx781+h49mZ5Ey78EEiCUcUMeQWbOxvDZKLeju22kcpkhlbEU+zkynNZMv
oOd4GyytaDNuXJyYcwME4sNBgpI/Tv1DM+qcZHPkEdSL+Bnluiae3kwlxnJd0MJ/Mlos5BWm0D2a
ijToXDFZJe+/i+TywbzvCiM3SWS8v/s8lVDboOLs8UTYK45Fz4iTL3RiUVSX9Qwh//bIrzvRZ+p5
FTAlGrxsKl+IqjDLydJYhqOsJSFZVmivsmzkNDwRAjva5BMfPINWB07gcvI5MlPSJxpuIsKjjslq
rOdM0JvPXNZONRGLONnGxlpeSimJ0z2QYtkI89UV5mUA5BqFX93ECxp1zUJ5B3HSZY3KcGWILU1P
DPLw3QIKakH5ydxKAgIVEHKksqp/S8s1lVr39+fKIVb9/HWSCdca3l6zG7nYxCveiCn1/dDhpu7D
kceR7+8v/xDrI7pdFXCohrJEbgdFmWUrsWk5DzcSQydR5LQz8OnSiwphBds5Q8Pci7c+b3tr7pA7
qGFKxiaEgaRuRA+3yksvIQ08kB6Ut2UJsPOxZubJO+OEEAC8A5YJL/hK9X5NKRfIYso4x0dlZGkn
neAXiR7nLN0CU0nf4XxtR4RqfJoFEO6iMosGn0OlxUhD4bkR3ivXghU91/Djq9zhRELBHD9Jzy73
x26pkUxtMbhOUv+pz+fQ8HCsMuowd+oykZXph0qBPUu//NdgDGsgQBf+hrIAeiPeUPQVW646+Ozb
MqY7jh19V5bsnrJ46TRHXxap6RxAhhe+dvor6vgGnFNMGypBFBe3EaOY07YOKrrac1wQW2rS02wN
O3QuCB1IeuRK9TCXbOZgn3+qki39WG0NQGyU+r8+JFKaUoPb26vEpE5Pk1k7VQkHLKn02nSUDhob
bIvge61WelVgqA5/IIOVSc7TtgucmGUVGZZFw/729ihDLTthAvNerAxFTGSyrXXZaI6WFcYEwzzl
RYH3xrrYHf3ddJJaqbj2t1ra1Qh5KiGIVxNgLod4AaDOQkRZFY8KGSedby2Tf/90QpIhiP7N3w/L
05KHCJQbnXe2+8FfLmb6PWjVvjNOwAFwd8hYcz1h/Fv8VJf7t7xWajeXYaeXGdAa44VtEutymlGP
anmu+WBSalA2uPx63NjCRcvx7Ecij1TpiAq6h51JEgcS2kFabvZ5oLUaRm/PbLSQjDdhY1qtnJ+q
4COQ/vnZ0qazBP1t8HLnSCQjk9NanebNRU7nPyYPB6DC8NHo5dbk0SF1Bwbn0pD1Z89+aAt6zzlH
jxkgR6HidTW4+bCKUNUzhpX8t2AfFH9+nEprRRAJHWJ/yMkSOq2oqDBiytpBBiNRxeQFCJoA9iUF
cQWI3UoMwFzyJk0hJGtRA0VSHRyXO6fkLpI3Grwzlu4jOnNTCmqpc+gzvAeu4E9UstodXgBR0jG7
l0s1F4EZyVcfmpxLL1XG20gjB4ZYML/X3pNn7DL/CkB8TgKhmZYkedQz3WgZ16NhLdFYHLqtzgUV
fPmOPqJaK0OoKLfxQ77sWdeE581dbH0crBwp7UHIIdu3XI/K0qgYRqBfElmaqbARSTBPfa2+ArCh
0HQtoOoeC+h5fPeQ7yyLCk8AGSzdmcSnytruSLwm3QK6cj108kZwuGzLlNcUAKxw5tu4fB03pWP2
AuSsuJOWh1asnizR5L8fzGIx0wbqD+qG8uhylCH6XVRFeZDUv1VOD9KhM5tXJjyAE50uMRs0R0dL
zqRvDUYDbD4OE+U3V8cA/mdrNnzoElLzy8zDb1hf7al8D3q73q04RJLrB5pGU0HnTXFnEh0Af6UJ
gX1X3QyChUR1pIazI9+dUs62/GEoIe77SYC+AUJNaMSW1mWml5sECR0y5x4f/0gdNUfJDv5EKO6Z
GA6N5eN8pHCMhqCJDmtqHbaYaRNebRXl1nrE9INO4nrIWaqBx51KKnshPnfcg+7RkwOop99fw2UE
x6ettidtA0SQv95nKHVMAu1Z+Mn3W2o13iv2TIx9QAUfqJ6M8IqmdmaYzCPRn5o3nKueWKkmJWTF
drN0BpdF/1x1IiSY49M2NElRfVXFZOXktymapFzjq+uGs9e127qcLhS+e+HvRZKPaHps653VOprJ
a3HGt7KL3IyK381b/UeHvdOVzJS08WjF8izACcWrYFB6I1YRQFsv9kjnP8nnm2XzpXSB+YyjoWGg
gars2SAuQIlKfgx/jss5UDRnar97freDx4j2FAo/K5ViOHASRO5WXRTOTPYN03YompV0+oqygYa9
A5ZZs8p3yMjPdV/+i9gtgkNJU8lXCtpEayCZ1MNT2gJ67g2anANJoX5D76LxY8pLRbZ4hccy9xtt
+pnA026N9jYF73ubVmOevTczal4En074kEuyBn9SIKMMJ2R9ydcUx6tIobg12s5IoXfPh5M5q//m
pAQneq4zbj37jDdNPfgjryIY1zDcdDSBHxAq9UroIZBTv2VIlZFkBecNRmXsAbfEnlRcit52eH3f
0VTodVZVJ4NUSGJMLkJMmUn8JtzN6PxkGKf0xoTRXEWlSkpDCdCjMa1W7Yw0/kBjxlLcwntdp/CM
+JVOBHTVEKBxVCa8/fT+/kN8MD/uUug9re+EaLkmFDyhMWhk3gUaZ3IUIQcMtJqjz7Zxc+/Psh5J
t9gitA57zUjenrX1LiRo1eZI1bDA2Hi5BrWGbIgGsmFWGqDHnNgKhKsdTWEw4LKx4umgtdgLrrwr
l/4geO3aBKZxZsj215C2LVYmQAXE3wOG4cUjnDJX6WYJupC3HMPlFfGcerNwO69Ht7QC1fnMnRyd
KG3ZGXfF0/CDgXIywN7ACy8f0cXad5zswqNQ8k3r4P4CMHWQrSpj2QME1KlPdOXNSnPFh0T/ARoT
u59XN0g2RANwQgBq0M4zXVkJare2TD1cyCQ4pnkPTUzsRf0u50gsWNvlkuWrJSvyGh/crda1qYM7
OFtRjxoz895okvJXLSUJVHATDMao3/Q5/qFmZGN1/SXe03zRMCSqNwnqFTZjJ5NlXGpw0cmLrzmS
hq1gGNh2C2w7LAd0pRCUBCN9oN0cT+t8JFINhd+5n83GIKv4cKWaf2rBu2JfcJrqyUcgiHnGFWla
NpWr0hyAuiEgDGkbE4qD0JPgfXVHqjuTD8cnaD3fh5tHMGLc0gKTwmrasyQ8aOWBGtKdRpT/Xgvz
cEi1II1wrz1UeTFjJ95gYmzIHhV8Gz4j6U3rUb0lV3JA1xXwQL3b+uGydA8rbll3pv9ieQJcNa1u
c2JgPJ8tt6uP+OAbPgHODd35XRByax0hkkmQX9m6Y6zQ3RUyT+ITAZBFhGmbWfjm2V/nZvxqh0/e
pvU61sGtLA1CrOMv6BDmmLwqtYuYlAr+8rfUPxRdJ9pSuOpjp8c41mrmFObpzAfTJfYY9yq5qRt8
CuzamLW7+8A8F+pTBmTiBCdkZzy0ZYLYQ7ZRdO4J/j7c75EuxeYvwGXv7vmdXVk3o7X9hvwujG9L
VCvzpyZjckm/dkY6eiSnwXYAY5NDep2f3NV6c43vU7aGh0JnalGIcS/vJHPkwLfZMjdL+7n32EGu
amsfjv3hLv9ehmxh8yzlaxI83TOztZkDdr6w6oz3awoZ/trWnOyrepy1XW/1TiTSiYgwI3wGmtBt
+KZEbskAAo3MAddkxeHfcoyLG2RcKOPC/ONZyeaozat5TwmVYEEcN/ZNYZtjEUJav2P9O69Gjuka
qrA/hoNaQLHqaJLN4y5VMfExC5kGE6Dt1ZoiEiZzBQ7PA136KDrwkTS3eJmmKE+O6lJIJItIn5MB
JrUc2l4KYWCPse1o+AgSlLTsZWQSi0So//tOO3oNnDH28e9bV/r6vfYPfQXTgXHV+FGEvtG7fQSE
ErOCFYqy4T8C18myPf7eiBcCW+O1HZeKQA2okivoHqZNY6fWL9B72vuYtjUP9Z1MFqdUJVcQzLhU
GGYN1RmOP51dsGlurQcAlH7wWUPQdj8qcanKXaB1Wvk1MDyZpYCIdTrpVOeOxiBXHscXpwd2POrX
+0BA+NlN3mPG2q75gDoEq9YZ7BvTzguZldWTne3wi52O694Bjj+UP5a5Qqaq5FZJuxXyiYDRPKLa
pNkI7TBJ2fRya0KT44ddUfcUX4p6edTzke39cTgR9QpvV66pGD5ip7/NkJZOEo2I2r7l8VvW3092
pDiyD3WH5P+z11YpBhtvm/47edK7WsYo4Nm57TWvcAk1oqv3fG56jIcLbPQEIBQPvx/ahFzGiT1F
dq0ZeiQY56+xCcZKYX/Jy5hKBp5wM6KY9l1OR/lBJJpxtXtaKj8tWeepNlKpPMt5/fdPT2yjWsW3
gCgGNcJkupHkUqWMwa9lpkPM6wrXVPn4SQi1vibag9rRdIlEPnJwYN8B4ArFoWNXB16In8ydy9qj
zMrry2A9IN2yRewp6JPUf24qrwybtcNXG3Per4R1di2S1wYdJLccrshHyX2eIC8lOTeXAWkTx/cm
QOd6JK67YtoGJCeyTOyYh1ccX6dzCer1QptK2GCp+rm0saFlllJmw1GUgV4Un1qpUxvm0uUT3gxV
gqLy167dnDyTIlEYXKQQ544pv9rsiaXSYQp/EgXHzHNo9QSBQu8uQ7Q/NngkeI7uzrDcttD8lWcL
ggTA3KzowzXqpBGKkoJlXKXERkb41QzengHAagg3qUqlXZDTUBP2ue9eWivfCOn+a5Ipb8hI9uty
iTsBn/10G0qF49ORBNl8KAoJhwY92SOjI7NyhwE+hg/72RFUtbALcUjtXJjEj57/TTXxPtIANMXA
COFl/zizXcYTEXMqj6a5nFYp8sv0ePuRtHzdqxcfPjs/6vow8GOOPrA2ZlAm+pC2KMwXU/rdbw4M
pabvNdwT0uzvqTnl+g51B4UtDC7n/pJeAc91F0JPr94gTNj5zTSWurSZMmHtAzv4b39KZUGerVcb
euGi6+buOWxsUjHAprRHYSX1BgSb4V3r90Ek/uQTsKmc7MY+XStGT5DQS+4Lqhft8n7ptH4TyxsH
QSCBxxtqVxm8Hl7EwKSFOsUrz6bU02wDULkYrH46FoFcB1Sj7xYAVmWX08dTt2n0zLLZXDJR+HMW
RRH84N82VKFKteFl38qIOvMeIdIqndqMYuAiVuF4wijoad8iAPvJnd8Szee1U1MiibaX+11NsFWo
uO5RVYrBVtjHT6HcG87aqflbvtgV6M/zlHrKN/75sGEHn44JYTAaOoonW3d5ZIGZtwBdYm1Hosv8
30oThmbpucmTeYHLvkINghClY1N0m2gOfSNSVpOOToekdwaTm+jV6KCq6aPGxYHzF+Fh5geQEBLU
301mIH2KGBsx6egkDBWjmxSRfCDhDvFC3NKy5ypqFlY3/RC9QtA5k8TjCvQSbU84RjvT0gO3v81q
aWh+tYNSS2PjMyjZ6inYwjiNuwhHUShX22VLO0b33b+mWHcEWDIacYGa3JspFSqi5wkIR2NEGUCV
Oo3GAM/3MUtVQ4+hvqA4G5FqQRMz+YZVxyQAdFsF2h2psz1HdRBCqDtu2W/jVodygfn1J7hax4/O
1Mq2so08+PiEQ8c6VNFjXT4xm5PVygdLgej8+WDp9zBMchq/L7K5VJd8I8GqpJeRKPvZPswQ3Azy
d2nIKm89p2ZZ6axXumvb3VOykj6QcVhldITGNAJiHZ6fKEUoIWoE2bjN+wN07j9nUHs+H826zKeB
GIla5XXp54wiAFC/bKTba3FFamn8E/s9fuCFm0jyqOmrY1Zske6HvhcGNHsAy3DSMTPLdmZfv00N
PJuTNxHtMqAi743OFGdr91sMiPkeA7fsAJO7SE3+pudJn1cIGbELWWBzCFUbwAbtPU0zvFIpkIj9
Jhw0xY7cAXsAbtCrhLHGrSZvfOruwqNs/tbAbn/esuB+FYt8F0s7oHyez+w85c0xk2Db6zIusaP7
oq4JGmWs+56G0+ZPnboDQtllon47u/MXb00PjjzbatzRNBNaqveQibRaRhgWXy+s/MN80rac8/Ac
E4XgTFr4sHrkUmTFbx9HWPeEf6d0d/I8lW53iEAJlpeHmR33/8+CblDzEuLakKXAmMOaXxmMbSgP
7zWWAUlsxwSna85FKn+kcZglbWOTPTGCa11Cl+pj7V52OWGLLMc2EZZoCgOMc9oHUNA6oac+Qunr
4zDTCa+tFMbZrcYEO4kZ98UlMCdeZeRlVnazOGkDAFohwtkwmaK+J8oFxjlmzV81Z4IxvZmpp3Ir
94TOxf47dZ8H8/bJvWNj88bzrYebpmT9gounqWaxv1FkwlYrAip9jEddHdXCArFYg2ujXuIA0LnA
njn/FnZvym6afblM9tHk/mrurwC09SWT/AF0L/vUYpdVWNOCXLDZTWMBooteUMovzlASF91zL/gu
s+7RXd9O80OEoAIIT9Wf8NXimP+62ZkE2IPVhDbc0QvX0hHQhMtMynXxL6xrRDkhP2sFXL4lyefS
Q+JiVRm7PvJa/3bAMscPVSlfFGNxxLZUd+9/p/ZDjxxWVEKCrcPxJnRHqRfUKWGZvQVs0IVurbpD
/7ClGJFl23ndx7rFxVYEIFv0dSfyrmbcND6r4wMvYu4/XDXT/jxRrezfD3QFxuWAvk6EFXuXsMWk
R+WfHrMUZr/o4k1Tu1oLBKdMgLj2HL9vzmu3ZiJXXUqSgXNjWQxz5H7aoRqK7zogfct+4Yss2quD
wFqWYvLEnEkMyLoooxTpLiDpM/8Z7GlsQmq/RVRmpSuEd1A9cFY0wUpDhWEJGkOINRkjwYty4Jte
UbySmJ72eUdNY7K4D08IEI2DQnQLcuNI/SubMQV1G4gk4VX6YHj0kj5Lm7MylK09B9jTMjBRlUNd
NkkK2yN5s2PrwSKsOKJPpu2YYVWQtvUJ7QLvZZoC2JYgOMcObouC4iXLLy1+aSZJwNTF6m89REch
S+l4TFA03lBEBBuDvAJ8hAj2PuTSx9EWgcjhGzzy61NfYkq3ICg7+NeVCn4ezdUzvF9wcNdfnt05
uoKNVhGGZOoF+kAz8SLn1WQKqsAywAxVFdovONiCRiui6h8EqDPebYaZnTHkBphAboiaqkmioXPY
tNfzDl3RNzuQkE2SpReJDo/5roGKuoVOZo0jrLENhHuh45VeHg7fJF8wtOTNBGum4837R0Pee2OP
5y7FqEcPv62Ux1OZLbRkBaa5BgRWqRijflYmbI8kPtQ1SOsI+OnGDLntFze8RUmF4n87kKf9vHit
ta2Y4oWh5iElzhH1XJnlkrfYlf9hAOkdT7ruHGnpn9kdK3IHHWo/TlNreBBAwPvHUppn+IGnYAN0
VPY0aZNXMOFHzHDzc+fAlq6cOlAshj83i4utVP1QJOY4gJNoyzqGWyVZ1RamiB9YJ1usW1zsRpv4
cwB8lrHkg2ii7Y25aZXTaWxwwpF/dql1kqofW59AYzhDpbXm4Yfoz86jZAfaLxfnoQUO5Fg1UpSV
UCRrm0/MqjTx6HfWhUX47hufV9ykrnhyNfdom46Eunh8idouX5GrgKRoXtrTjK+M7qQJ1/zt9iyS
B2VhcdWfv1xBrD5wNEUlfE2yyv2t3O9gxsBjY4lys7IxJ8WNUeC9FtaYpYi6+ruTx+8MBnOJhlF2
4YwCt4rE1Yzc5Xk33pixkGkQFk4Gb1mOJVhgFAx8KypUa69xnB2P4Y7+81hpQvtLC538CIfd2pQ/
X5oBsc437dCRFKIZiGoEhoJ8eaYNYD/zvkUr1l+v6i5DILFmhvot2JhNbyGRxpYlano/kgemLc6I
qYcbxLyAXHwnuQXg8yskigFmN8V9VvtVMsj8pDj6TLXg2ZPs1S6gF3k1sWa9Naii49XJGYiOntfQ
pO8d+q1RQ/ZJxpszTf/jexXeGpKI6aSidFJsUsgIYnH/rlS9P+zbNolxe4ty66T/mJqOfE8XA8Lw
yuw6r4Im8UchNeQaOWDwQl3xp0KywyMZnj0wkjSzfFtUxicqqAYCSs1n5QJOq4G4Ax3wU5hARkNZ
h8pdNp3tG+ovNufWTmkA2sIg4vD52J4Ffof/WaTEkNc+FUI0r+RsRO2zCljqR+TgrMrDLtkM+X3Q
X27YaEXbtiaEbSRHJakvEjiEbZ2ZZ7RLmG3aQB/gsjjBPWvNcZp3a87nW5dWTQmOV1409whLbkAc
SsIDRNLBfcAD68Uvl/JaGPKSxpu3qUIJbuoVi+UXwJ97iozB+ROa6KuUSgAp+uJq3WgRBhSx5cTS
tc5GtYQohIQvCoQCZa6f1rN066f4O7xDoHwJde3+xKcQ8vrICbFLVXDVvB6wO+9O2qk+GvPiofgQ
3jiE6Iq9sE5o8loKKR3vMb6yIwzFkMz+VBnRHcfoiIEmFxJF4jEAIJWM9dg6mnmLAj4ks2QNnoe5
fAd7pn1GT5NqFGBNGmz8CT1GY1jxYY2idocU8bduoCCCVsiRLdCI+SF7AbdsFNXxzJhDdKLNFJHB
N50meKRRyYc1eHycAUJ1DysAH19Uj6RRqiQ7YacQbGA8Z3wvT8BT2eSrTxnC52VidMnEIvDAiO+X
rG0ZOLEOd04XhvrncGxmjImzWETu1WQyIkiDqq/1qpwxHk2LNeUf5XHQveRu17rkJH0asEwbTSxn
YV4pHneWkWxjgBdq5WwqSCdquon2VuOhNw0q/gLDlq44vDKL+jQOyn+OVrLXVx1yzn2qIlcJ1qB3
HkSnul8YslZLLJtCuKvaQbg+UB6eOdmEFNEfskqlQSpaMvN6DSNOPB5QKl/PdK5cEf0SYmS6mYRF
z3Nefhq8F9sdsi9TeXYAmDrqrCnr3a6Z4RaifvlpIehTIKgpVPHVQEnFfw2hcxP/A+5KKNo9zmWf
Q4CSBSiRxYE5ol1WEZBFGqB8HoquYKbYU2+2T/I939UeJd34YTaB3SIS/jriob8ODiszvRH/h0bS
3+nUjPKdtcPboxWS6fw65Rbj5uV1WLsB3PW1JiNobEBTS+DfdDb3qJrd4HNuydP1dlEuRcOQeHez
jLyMujoG6/ytnPwNXKbe2SQpEoyLNjXm0jRLaAuRAVPOvoB60cnz5aa3nu1Sx0oWwY67s1P3356z
7J/L+hCkziBpafMLHEUWWZn8A+UPerJA7gzfbUyFS/6Ze/CPhml3WT8ZJ9aB0xAt7ZsaiEAvCbhM
NQ6zFXsLU7jLDhqwLCrlCb7IQb0PWrzVIus5kIuWBQgnXhLQZj0ejVwTMsPbwkinHfCxSzMImBGw
WVV2LDbfz3Ga70CwrguDjq1HfofjJFhmOVS0HnXD095oyS+TUqktddCZ2HZu+xCSmyDCxTUn65ir
7Rn55Nd0KzYqlxGiVT3cE/G30bYPAd4NEKsxiLwaxFekxMTNNn75QeNa3iIS0EgAtsqkXqj4YV8t
DLn0ZIwq52k+P1ijLdH5GuQXCB7lOwlgiErqi7UIFhcxUIcVJZ3+GDYqa+PPTK7DkTzoWCJ4Bqnt
8T1nrFxlppTO1XAZocUm4MuaYE+cGv4AEzFfwZ2cRty+B9tfaR+w0NHw5QwWBAih8hqYCLxkXALs
hTTzQsJfVYKjb5e8QqcDH19x8rHaCqee/Sx8YX5fgz2UmlBl8/Kn7xMm0ADKdhLWKe534jpomTv0
aX8epCFeOOZ6cicvSnYb6KE6MgcvNzIbpEWIEkXADZ7Q3aH/zHYfiPWYtpBopEOt2WOW3bTBpt6D
HiiLfHBVXW7W6gZP550YWproCMnNJyNvugJ4N/cW6DUy+NYCLap/b98mc7C07qjlim40ctbdZ7fn
Ysj+UfYrbT1IGS8AC+9HiRTzQ4HkuwOmPH0T/L6k4mTBfK63oyNsFKojtcLGynqiQ6ZUG+y6zzOd
BvkFsEV9LdUynYC+ufT2/wOX9Jg5hNGZoIk0oN71YkUc+gh8igzWmyKUQ2owidkIBQxcB8d2QSEd
T84xsR4bYKdNTbJa+HJY8GrZgx8pbo4zspjuiCmhxwe6Kbv3Wlna0d++nELpPP+suY1UthNkCELm
DWDH1XtpHm4qLqvpQ9Xg1wqJTQPuhxCPaXnPSjtXj4cwySw6vW5yH135aH+70/pMw4HEd5PL45l9
nERGMAdP91R44lwWktA9RV+Vkx6O7oNw0NHtuDjHCCxnR+p3GSmsrrhK3+JKotiSPnEEy6wjX2rB
R2uIzntzv8JudFW8Bl4TMlVGvzMR4bGEHTe6bmrc9wJFXo9qj8dThxal5BKQh738zM6xrgYfiF73
gq9lFdni+/QDVJxxXFc7cZadUmV6Eq9snhvNQ8GmuvohGQfFf5E0G5lx7WHEavuHdACuzB4wGo07
i2yD4gWE3Cn0vozuFXpvy0/mJNzk6Y47SkmgyR7sMp9oKLRoYxlm7uHuS4BGJ8d97n7HBAuev3vW
WltT6IGXF62xzrg7inMUUuJGRQZg+fvHq6qIeBKHt+0WcU5M6cGBA6DM/OdAcs5H8r7y17aPSR2L
uSwcqcd5vD3Lue5ng6De4vhA2QVtB/r8cR4REfW1FwIV88tIIhKMCFrte58q34vgJOY0ulqPWCZD
7LWeMtkkS3Q2XAUxUNlf1kf7xw8Hh/8k4IDDwSPOHYXXeQTGWx4jhzcsWaevCaJrp/rzjkkHBV3q
LQwqH0sKL/i2Y8SR6OIBYPGuvW7O2GXDc2EpOAjg9JgoFOMF/ozMhnFSoZ0nbxOz4aneQ3z76B1p
BKhKnifG9EyUAc3tul2+oEqnHFb1GzJHANK5cJCr0edYjDbqp5Dc4j5CafxTbQvt0qbLXBpbkHR0
II4+cwOfuoMi0Qv5oSJHPX8Liv9YYCLe8Tqhop3XvXf7hHEp/13qjSJ0INVvArJXl6P5amrB21rl
f80XwtldlxtSgZLFZACiiePt2WoTDm38/aFSccKqr0YQbgL37NOh3ssqbbdg/YfYC8UIsegPUR6J
9ACw1WGO7VyIeKCUiiSM/Ve0KaX4taE2QHcXpFPunfWq2tFFhPWmaoJZ7LDwMhVmP50scxhI7FmQ
OeGvnhqa8WHPleYNg1PVnV1CWnWt7aX3rynFdlRx/7x/TH+rr+WDB6K5vhb4AHo03WEl5whOUXwr
Vh+QIQM1OsrelpjFtx3G1sVEs7LLS0XUK02UyM86xMhLodiYMHJfXvgZnTwdj8URMv/kSD9hOY7/
A5S6pVU93ULGn++P9qVRPoFfViNNhyvP+PUGRWKt1GYd+imuIIGAXhZwPfz3YJNrk0zSwSzIBgNp
fYuzFgAV+ow7rBppx2LrdjD5/ZD5A8usm/bMy2Uu3q3TzxseC5p+rjC8B7UXbh8tfTCcophBTG4I
9tv+ZhW8e2a3VfxgcQGKgPsPO7cAJMPq6N4u60xf2dzc+dWHJu5qdvVPofzPOM0hT8oKMCR3l2+S
AeQQQ2EHnq+5e8bVa55gTetm7dTK5Kub3sqVCFehmXAY0BAruasFQ93EUn8CBBscXkm5HpYEVPkh
YRGUREWJAsbeqXlVLuBxLj+GOHfV/D3/wtZvYIO3Poqwt2smpw6SXTUP6k6JRNbxk9JXc0gzFQ++
W29AsE6XFxtt43M9oTbBRWxhSuEuaWtcXPUzcJpVpFB+09R4lNua5qWgMb9eh7c88qlXXOGvJY+L
jhYvTsVUd+9dj3yD835RCh3Hb5FLH63hDFH8eJZpOLSGO79Jxwpo8ThRl5Uc3rYE277t/7aGogaB
eEeeXxmR19vYCBWQze/2VVVOVRqWYyC2Iw2MuimxvPewA6q7/qIQoKerHDgNqkqINMZ8Whr/JpID
qT7AaHtj40V9OEPpQghdv/3MOhiZ2Oc+5PvlJUQPfWWzm3wGvmA63BASb1oupPa7JBG1T/o72svP
9W76VyG9yT4q+R9p6pCy2clZxhZ8o5NcdjG+uGlsx0BN+X8tF6df0vhjJNEt8bMuxexzz2yDhhy/
N4jxs1Fb3+GJxKSUQqae6e6CXcMurhcc3HeSIxYK13w+f4j+c/VQmyIb55jIfnjtdyr7hKeXuJwH
EZP4wRoq8eCQu8m7WK0uRHcrxfMCIBU1o8kZzKBLD1JQOIX9LAy0aFhQPfRBa2gNfAVvx68o+rb6
TgcuZFxzAkHcY80i7z98rRGK7hQ4/ohrDEfhDUz7wEWlwqHb2jHYeak4NrOhKcYkPwm/CUOJzH4e
tIYYl+K+qXNHYmc+gI1wG+qtO5MirqDAJ2yJokji8YxUIyrYJVBU/O7o8VxnLrUQ4zPHV/YN6TGL
TmTJulm+7LC5XztsoIQCwAq9HWqDIUdRFG0XTvK152uI2RsXllz6QeBSZOEZUTPpKBLhiWQNO/dZ
QSOUmUVb6VdU4IS+wdpTFFB5yqmNkQLNlrnbn7nMR5JSrfhhvsTwUBP+syDj4OD4ssQELeGx6qgE
c6hLZtSz6TO35cSdiSPJ7lPf3ntCAPXzWf0v+8eWMuzAkL5v8UiaqgjrO/IdrVkU5DRaOAOTVQh+
vfJcmoCgHfrZ6xagbBjyfmpTFxH3dxmRvXBgKvehPaXnWYPilAKdhA8Ngvz+D25LjEXYuIgtk9lL
+n3QVcGNEzoUBFw/qi2C9M/oIzoklLINx81Jbeij7nHiAO9Vop/3En5q93MDdrdzGWITWJ0JXfV8
0GwhWmrZYQl7W2wcF0gPTLMx0UNvIrgD5raK9LWHwUKDWDMSW3ZNtCHVhLXkAw8iFd7spQBsU445
3BFAhp1HWEJ64WV15KYSZtoNFgJ91Ya6yxw/UzgfbdmidOB6f73nDLogHgssaxwv66NU6zV1li7a
VIp99Ipfy86C5c8D+dygmemo5VoAJ2kqwReuWPB0D6eUzuiUZka601NeZKs3uDQq3by7a15TA8tc
0sH30ag9WYNWohOEG+BRGQL6GNZuctpdB/CWKvBcqjldoREIKgjWcUrEhiFqUxjvkbuwEB2uzdpP
aNckcuXEUFaNphV+RnB4uc9g/Be1GQWI7VlK+PiIAlXvMQQhAldeeqV9qVvFwG9JGqkgPSRzWXFa
zl++Wxq++tDQkxwgCcFsWJ9WJjY1MgXsMpZXcwN3ZEm3thYqteU4f5RKtmOaJf38DzWCv0XHznew
oG7pGfKp6I5Ep6ibXXoEqHzt3oqN+k4i94RGFfTp1NPauD37hoXkh6waH7TSclQrRIsDQyqLn3/n
EPc2yDKckK0K99bb//LLrgdrcCuviq/CCCdeJO/FoWirheWCCvXMlahbwIKBj90Z3zgqlxdgQsqA
hOikHq+GWoRcirAYukd65KiWAmm5Ww5e5gwIsg7clvorkice1l7bBVtZlLhxy78HT467i4z7nJJm
UdmPokH/AOEKe8TAiLku4NJWniGCuBhGLF1zb/BD0RftU17fF963C8IEtrzWFNKphchJyZ7r4Lr2
NLpYnzwyDeW3rbwy6rW5fQGsLJ1PZLHoFmE027TMmvqZVlHbUFwzhq0I/rNXSUroc6FpN3nYpT89
SqoPbFGdgH65RPt8D0l0RVIM4PUQ4VCnGA7UN440Xo0ubeBFBMH2JAHxcwj8PIA32sQ4oUYySbNh
eQ1PbCLcJG04u9YdB/wJfTuMT+Y7XRdgnyZFOpjxRhfgKbt6T/AgSiqzFsHFbriKwT2MDga/xtqt
H8SYF6jdMQMPEl3V6WHfoQzZYpWsvHGG4n4C2ZeJxlFAK65PQfn2RshGa3+sbLP+nhjpHYhwr2mG
ZCP2ztIHhnDxdOfwPgIFLd3Yxq3x0gS5oPXH9f+VqAedUt7K187M/d95nYBEQ8TY/X5iz9f63nrn
QrQD7ajcHGxpjhn+QNhM7tDq5XR0LrjLq9egJapi7sIBc7F8ALme5vntkaQaxxLt/4+bHyHLyUF6
2slkeltPTed52mtRnjR8Dz2NnpwfzWgCVdv/guYwtGijXpG1D/b13+3GcMzlks2VRLNAy+FBJ639
51nuT9ALstWGjMCxFuewW/g7TDQPh228dExTE3i2CDimrhkCoFMDDY6ofxyPMNAAASiV38EGxpi0
FzAXDcwt5r0XIMmmcdzAEHK8Hpuah6Q061Kezmzilx20xWJ4focztPnSsXUz7RKuUFi80x294kt4
T878bPwRPunPaAUySoq2+aEf2jM9jP+2swSxJEVKbVBu+gF3hgN7+Pw6WCgM/CMWQkEk5Q21sVGT
yCabZ3obGQQusBuq5LR4ij+mM11y3d4mcdUgJJtd/hNvmqgaAmbzI5w53MMoEkEkfX1CavXDCxJg
dL7FYG+QRSS5m00dFz0ZMGLxAHvQ++oyvyOBZLFJaavzZzk/mC7v7bDlqEIE7axEkslqOM25ulhO
2I4KZvGv3tj8lASVCxiIlaVTW46IwES71dG5+gF4UaOYFvurpYBNS+YHcjMRbE6IhhFzKlzg+ltt
Cksu37XRkFw5a+q/fKHFL01BLC9SGmBCbsZbavC/6cX5gXU6FxgGKAO72S820rBvHrRcGkta8QaS
bLEus31kr1DcYmlojntvKsuiLdwLsY3cYCg8FTAYKzBAgQ+K6/ivnmrFeFST1uGKGdpiptwInmrE
Cp+1qbpxKQ6nGvstoQ12FfFjd8Pre/5VrpqoZdqecniMbRB+qwTur7RGyNJuvJNftulnP9MFac4y
tDERlFz9r6zC1ezpUGk/fpR5jtC1AgDhnFRlCKq4ArHFBcxhJ9CHDntmtrtIXluaT08d3YiDmNtF
HE17f/s3O4j8LRg25Xep9gf7RUTMfugWG7/HxRTE0E+xRr/H7dQfnj3o60WasX3U7gsfKtP3Y3Bq
DSZ1ZxDplejKgLJVuY+ekynycX3OvF1d6HO163te8nMHXyQRzzS4UlJrW+VekN3bmWSF8JY3a7oy
DkZ0a0o4QqOhTg/O93W45eUoV4ed3vzl1sJZ5S3gzjZJIg2itoJZV/hahP2W+k9px7FONn1wJxaT
XWWv8BV1f1HIx6RkgDEM6AjxY/KGR+kSQCtmKeu4Ivls6RPZ5e/Kr+WYHzT6H9gmgnek9IozLxDX
SpLfUPORDK52uybWAOeSBXkz33/F07gCkpdtxXeYjoUr25IJrimSLC1uHi2xeFUCaPvUfyraNa8t
DQdR8/6C4e5qU1iq3lR3kT9F9a9bCbh9ZoOV4iO1sOOHWzodpyeaq5/iY3B7Walh5QWhff28yeSS
1vYMbzickZuM/srHC2Kmtql46EHB0BADrgmEbLEDn9KQA+kyGOsep3s+QhPAU2V+zyhKmRJxxyuZ
8uwdTYHYh2sHI793+Xoc7pEy4gYNhVmGpCCekWCHt9dXIv0+f9zf+/nsNPYBoICpGGudKY0Nr5ax
c5pmtg1B/bXE1Z8R80jf54K/8w808mpeyujQBLEuF552qA2gckOH+3MPwEyWYjWsLLElXivBeW+1
7V/G20LElfZY9koLXnZT7BtRN49uwnaMFl7iXt+nQ9Q2c+8eNAO2DFD7Ajhk8B3FUoEFZ9btZ5Kc
Md8n4fy5t6nUCfwAH+nZuOn8pwci9JDQolwjeQhKAayMCz0myORQfG0ocYhclfkJIgoHaKRwrMOO
OJqjwBvhiZ0Iot9jxUy8SQljjEMAdENS1D4Zi5e7JEBG+E1E2J3v4FjGXe2E1q8i3qHytdsoIJbk
dys5Ltr7fQN9t8OvWOLrSCPBiWB8xZm7FEY1Hdq8FK7aYmmGF37HAG0FFm2BSRtS/X9b7QWb2qNC
WonhNvN9kPYXVCa0CYCBWyvpwcjiSGCvnd7xCpn1VWhbibvSloVrMD//vRjcnEnzlugiDx+coM7y
e/JaB8iZLwBkt275AJ2TINjQIoae6GHjiMCWvKvtwnin6IRjHrQlQ7HYUXdxNZLjryITokmp69hQ
CSHRzqDSHfp16koUpyXjfz21FNbwLJtshl3v/iOOYlQ4YFg7zyXRi7Xp7qzatXdeREkS3DydZgxy
XghC9sm2KLE+cD176pzNQSamB4ip+JH0MeiWPNSBkk+Jv0SzxO/dAZUn5sjycV2A8UhVEWrPF9cW
1q8sXTnQtU+jYd/VKW97bjvE2RvQOmnfx5DDmAq66CwjZTqtxCDIb9Yss7zNl90axLhZLX9HmSZO
elFcW6lcquVlJopjrRaMLk71i26ywXelNmdr8StnpHuONThUBUIODaEthkdUzWUY8KAIPtAT6gY0
NjdJjXNaXtaS6F1yeVyjjj+bFKCdD1KYsuKlLL7+2hhDMlMP8xcOtMWN71bVg8aw3OkQT79Bd6JR
olvJKLDMBdoHr2iHO+rQbCZnok01uNEv6CqEykLDb3zXzFADzATYNIliLH/Q/ut6afHOP3Xi9xa6
wFMcac8jFmjeWKZdG+GYdok0TKxvhOs/KtxrCGUswmX4gFtLfQgpn2CWYjbwR/sgUK4zLb6+GRkv
oW32Ms/9vk456hgorqZuMH7LtswC6RoKJT4DKFsmAVQ9ccDcwtmbmj4elhm9NWOn8D9ae797XKYe
4tMENfEn+JLa3lTSG2cLWH4CfMpqporf6ESXnwj7yDPrrmES2ejhm6omQihd8Mk2MBgGudM2ORyH
2Kltze3vjFEcK5MsZV7785hjok1ZUadYUGZGGyat4GN53+l7WFFmU2skXnYSd6GuuHRcHJ5BHM83
Yt8zBN8ptNWTCKbqI0KaMmInkstnJIHjSYli5UG3W7GB8Isl0g7ntqq4lDByvNXdI/HPDGsUstFp
+DkFOqF+BWkiQaWl9qCNKcCTQAmnPzaXVRSyDhXjzRc6uYwbjmuoORJ7REI4eZ9Fxe5zKQH9Uxva
TZyhYhTHk2kmqo7PBqoUmMaStTF7aboC5cyre2oT1gbx3syNXDox0Vr/YCthVMsU6/RhOyISN+RV
fYRobD4Ts5k87zl3pOkp2UNRNUAG7IidH3l8QszOWZgYppmMQhbq+QlN6i3AM4mBwN+i+mAx2Yuo
QI1x3kNAZIKMPw/cZ5wfOABDJ6Z7IinG8W5iaTmNAfLZj9yJnS+KK+dcyoeMJcNMJ6CHROIV9MEG
zPZTzhenP7i/DJL9cYEy+5FGDHsBRlkEa4xycMwdyEyUNV9G966f9qL+o28OaSTSv3sxbFeDbKQw
pAjnN8nVg4o4vJJw2DMRRxbOHBqU5Eg7q8fqRH/hCZVShZGEHok6Xwf9c7q9vxCLWS8QwrokfXsa
5UKQ4QyF2jxacBrsdwSrRjuMXkbXuC1w/wtGkvfeIiKYo4RtJBb1GelOke1Kg2SUDzKzO+S+Sf9i
MEYVKCVUz7MaD2adUuP7H3Ud9sJY1RckMOCK8MCTb3py+9ZcsCVZl3sIVRNo6gbRTyfdzs+qPv3g
ZqCQnmv6YDnu3ke7jeizxe65rWqIQPvv3GyV2G6FBKhvxaZb2ptykyT1+DQaNwpdl4hKS1/sdUtZ
QP6Nvi7d0TEz75GY0uQVcRmP+lyonupIUvh8FJ2L3W55QhcuESA/6h41rtq4Ceht0W22o+u5f4xv
DzW+nGipnbuGjjUDm9HW32SRhHlqAbEEgH75Ok89omH3W6Ps8hn1IQPpQ0S5C+UzO7j6rqtn29Jz
3z4haT/66HlxqO9RmX1nQ7/WgzvBUUNFw+IUedT0eRerLvBxbWDXiX8myyuRBBMXjmQhhRtg7hfn
oGbFgwDlTYwnk1d9kPxge5J8UnXp3SlVyjU4E15wpyCVphvpr5sUQVBY5iGy0MYChp901BWVd3ra
59uXVkbzfrEfhGlIUXW9GeAldMePhxrdCkQ1CQKJBmlgwMvuUBCjNSd/Wb1Rhck62WiRrQn6dgri
JKr28xbNLlsymgxdo4d+8DpwrUQics3Wu9H/NHJZ1XXFVLVe+T6FMcNqf2q2ejFV738PDj/Xghff
UbgrOMJOdjNy1FRRh8U5B42WH9EREow7bTsC6ytKQwdb48McLmQvyCKEvJ/f5FJzGV38ck7spXKj
VrB8L4mhJq+1D/xCS8MG7oQvQuVe/nu8/isTBZq8ohpXVkTkSV/ZMRzAOa9I4H+4pqCdOSTOQcvK
1VejrRW9cDAaACg18u3SNkqGir8G/uOCKCiWXpCLF16OGJ9DKwI0HNPRlhTolBhTD0k3+RAO0YAS
NRAMg1+LRqiJapIBrx7wPhrdBBifxMUCNnM0A77Qe5nxFjHYUimEgy78tLSPSqsVGZ0T3eJe/RIA
DGJGmCASbEgovo/6jv3/aPu8c8fT1QzlGB2WFHX9bdS0+ajmXBmg5oYP6HexrnjSUjlOzS+Tah/x
yVXOXrDZLb2jxrJFtqDiW2q/6AGMdpbbRYuZMnSVxF3eirDG6G1AMrrsbjjbTMdxqOLr2/1lowCB
9pN9PT0o1Z/y2J7q1e1+b9w2Q6J+tVTV03pN5Yd9IsQnkDRSpJmL3S8NjtDURHyzvLxhwcXGvtt9
5Th/OHR8gqMMS+dxE6ikDqT+k7u7pxvBHYIPX1McDudDWL39CwVDU4oxmDRi9uP6v/lr8NnOkiAz
ew0wuaolOi56WcROe2gWJkq3PkHQHvNbiw4fNJQJqmMEUkejvRvnkotXcj2YaK9aBUZJI24JC1i4
yQJXCdohiz1lvHfz7Bxt5EkJeqhiClCOztgpGDEPTLrX0l/VewAA6rlEEeyYNBrzbfhjMTjJ5N7n
2fa3LuYG6YgPDylhDli2+nTVJfKC3beOGHulPYXWNihuCMujMgawenjXKBv1k/7JCaGj1aWYNOTl
n8U3B22UZ7YKtAZ6AM9Xm6aMvTzaj+rZD2S7Gn0LvjySqStwfnTcSIbb4YkQvCbw5j2zmQla9ovn
Od0My90BNM/ztcHDgRLOedHQ97X2epM0Bv+r0+FcveVJr2alWkTJ5oCLNwe2y57qds4HOfy9vljm
hYWXpCDTOBCv8jyNTlusH0cfq2XmlcXkdwMgfWAt81mMp9003ObhedQhXaYmh/561vNhr0gR12ya
VC49d5XXL/MoX4FSvehQh272USxwDCtTII3Qz5WEwTVZlylcbGTIzVG5M9L6PnniJ57bJB6pyhjb
hW7RKD+Bb3+JBrYMhExeDyFSc3iwae+sNoLiH5wAGl9Q3/jhJB09SiijBLgOW6/IKKxrPGYE8+XI
fCz8Q3iA+fZxekvQDlSVR8H04LG768LX+eXZ9DJ5xSBjxvJr3toh2RwdfcH20hb4kDJmWt43DQjw
DrG9BgeR9osZe8Bp/kOsm1KwCZwhRz1IEb+DDV087+gnnPOBcEUjf79xD2ITdYiOF+/5p7uomBFM
knP3QvVJB0Czbw+du8NIYajxNKvE9ghOHGA6S5bJms3SgskDWizYDCQ6sr0Wz5IrpL1jt7qinCVk
79LdkiqKaxQLHCaQ7roQCLiVkeVdX7wRB53JspO2amZvHby/eySp7qpK+qj4bVM+9b9jVPz5jK2e
+3zpyIviznaNZM1fL733wc2xjDs25jS38EANtUB/uKKGKS7SezGinwRnTo66LLjWx8/IrYvqb1PJ
b3j+PRk0YZ3su+wmMg3/QJvdiVapKgkoHGhkQEUqekmtoNY3D8omIEX2thZUuSkuNxF449Ppkm4m
WWgCdVORU9+EE5V3DLHwEzznFLOvuUgajNeaghUmEtF9T9GnNAxUJb7GfV397ZTzhcq31wairKmP
sq0nXH3K227+9e7WHS7zD4PDZwiiyv/YkTZ0GDoWYhoyu0xXKe/e4DYd7aeMr2/by/6sjZp3hb8l
IA2GXZPelkPH3kPTkU58BLea16m4FFWpWFUr/fHu97ceUTEOcwwejKrf9XqvPO3IGKUgXOb+/DX8
N84S/kcWABQ0nn2noOmyf9U/uQKUwwEQaojLg4fAq1kwHPgyzJtpaaHwRTb4+OxDBtRnoyCZwS21
DldP73DAZIx4NUzKUT7vIcqYdfvAouKH1NRdeMDoCgM6akdT6ioRVmwBnUnfbiJAReYb/RQTdm94
bq5O2w8mSIcjqxlpqxSAiYQQmW3gieGs74hsgbSv3vvzYTYXOUk9/YvLHjmNO7wdXYIFjEcN/YjH
MX49dLLkRYxcSKOa/hP4nJh3cykRnH/eoY9fLFSU2rEBGow6B1VYwaz4F1TC4/RFVwnPr+/szW0L
QQaK/d+obCi3Xd/3DkRENoeESVWA1JNwBTzVVDSf0Vx7iE7aC9WA/jkoOKqLZIx31vA1t9A4g962
r0wzG9xGtIsGouVMaTluTPjH9v9HKZnDRP40/Xk8dzehqwoIIT7YK6pqHKTt2TYeJ1O4OHIHsKXH
FKMuQpn11KD+IKAV6/sleq651jcjAjTZiWc9dUdMS1SVPnXE0+18hGrl4YTZcwMsTzTpW0dS7Ej6
EaQgozTHKN6HqitQvmu6DtvVnvwZFjyw2G3AWh19AeAXKwctoV5nRdA4W3WZHgTf/HX6fxTtLAyi
50F9H/ng9pAWDj+u8GX9fzhlVDJdl6ttOOtXZmArcpl72vkcjkpK8jMwIvLv/eW1W6CMgFdRaLzT
884k9i/Gig4oVhLdIRVzJAYNEHU9E5AMBr9zgxJjvDxxBlJNtR36F8upjs4fEZtv7+HId8xXyy8B
LdKKWiQsy0dpY184Em6C+ZfXxKkkFg0q7UsZPV9m2Mn2XkO8WYxcoh6iKQkGWF3Do9EdVmI65UCi
nfN+CRmavYWfqhwkdshQWaGX7bit+YVnfg1Yw1QXjnp5Y+c4FCWWGGwxUYKF1a2ynyQ6u42IU1lC
87JyWuOkMvz7TcTdZbri2/y2cjbe7gedM+i+kR/RjsAU+z6iDh0XuxYPZe+Kr02x3CKnd8bLtxVO
zIA4Dy7FlouN+BlYml0iX7hXvtjiXk/fcFu2TcwEns+ekTYTFUt5pBeXiZuV4J2mdzhCz8817Fq/
Dy+S8J+cWRj5s1PCquqenS2zqg7eGC0r7HS+gn7uBkoA9BIvfuiSQKM3PnqwRC/3KK0mkRymVECM
GLaBNWUoms8u/d2XFg9NDbi9nziwhuPy3atjVyX5KKey7679jZGXzTZ1Pz9NoBpi5fZ7Bh1eNCtk
96OmdM+aesLZZRPxbGHtQVi6cmckMEtQgXdwn+0Em3tqfXH+J/so2wgCpNvCgi+SCjkpLwu5Ns69
Pf9UKRAMUFGTH2/8S6//7tVYLPaSjqCdqtlEzKxt1UHqm5v659VfeCxrUmjXPXNG4W1sWYQop7vq
AD7KoAxk4UHibAHzwGg4KcIGhW3o1zPw4XwYGI8pceG9p+8CHKpPPeGj/g1RHV74GXys6j5mU0sE
IANYXvY0b8q5YYAnkvp6JTLYp+VoK+yLIDVmNHB/irQCMNm6RpoFfolDve02Asje9tEDdV4TG2i4
5Unj+9RRRWtuqB2dgO/KL+S9o0jxZtTmjtz4cVkjHULXXFIYbqGUbuvxyD+Dhe/INFFpFpvwlX0f
e+anMP/XO1642N7JSCBTf1rWl9IhnHKDhHAqlNzaJq/frbc65wO+UFDfD3yfmlVLde62I2RM8O0J
Vx2UUk3hJOYZ7CtNEYeOCIM/B6Okpm62w9TRf1psOMNO9mKC04g7h7iuc3BRCJtOHWa2ld8YQ8ox
2ME1VIVNunz2Dl65shhnaziqsFejFgWu6T+oyFuS6uk11Q06QDEueuJ4cqGTV44Jl4koBBlIPMF0
CtIFGGq6NY1vv00rRE76abX23tQSfDKWfCPOaOm8/AgHIozGyPC3OLjVUXWMmbxrvQ9IZT022ZoR
BxAofZjqSKCspGrrWDutatExAaUAeLCKYCtoYWLaTvhxJrpbCbFy8M7EGTKb3chRl2PP13GkWhwi
isQTi0DmhxlH3VeGVk0yGAGQ2SwIwVrjUzrUiBhkTUeVDpdpIm/NhfAaCMdLxT+8MkzYOGtNGK2M
imL8l/jGtnN8a7LGvpDKy0eCbwrIWZ3gSVTHFXyz3JRl+2ihUoVyKP+iPzDBT1uE3TeyK8hQu9yO
9FGe69r5+4dJnKKdZ925eeLvvyF2ErG57XkKPf9M7Y2uxImqedNmLZfUq0X9gFVfji181qiHmsIz
bJj0SDi5X+1a+Myf+uLDNTdjK/yCwtYUH3CPjjXaB+oXHs84mLgtCfCwx9zWaFGZtX2n9mPzI8ni
NrDTFWVimACMH8C6UtCEMWfXWPEDSZ6733kwkLafe5ku/hmRTTDC2NjMvSPVzI37tdFCL90Zm9Go
LQ005DRcj6TsabnO+I+rwrnsxUOtHsDTRZs0nw8AUdGz1Rp7wC841XZtpjtwsOCZbHp6UJPQTKbJ
tINUWzcW3Lit6/kWhUlRcEuE3deH/oLxJ1nIkUDjtryuwhqHa+klNNQrabLvyhfCotiw4Kj4Dwk1
C0siqfC3T852wra3GBpT3o8mTEq5HkxFN8f63iB7jtMW1tX+BuqC9qwYaUFYj9wZzAGouRRH5VFe
R57n79v4pZBCzweCIafTfomNSelPn6tysPHuV98fh8ZZOjrDhkcgmDuq+aBxKype/Jnf66LMzzhg
h0+JHH/O4RaibtfWpNLz3ok2GNRm8KDCUJSiKREqbOkTcrJxh4aO2iqqbQOp8WORbFPO/GMzjDas
4oFQcP9yz7O9U4l5IM0JriiFa9brpEtI8OuJTj7QnVKtVKDlw/QM8WbPlyvZccIeRaDVmH1oFVlv
E9MaRsWfS0/3rFq3zS2xitS1LhfbsdQy8o3oTxjL6Eoa5XfKFjYslsymjWisYEpMqJAzbwlNzJJr
0qLZ0gfxv2Q5dJPHfsb0k/6+wlNZBIwV7wp1JTz6fZK9qERH4xCc8b4WYyjRAl+uR8JbL5DdYznv
Co8XdCapk9Y2xglZA34XTWoxCiAfQX9j0K6CV0D1cOgiYScwQ6+JLaoK5orJsTUGKGy+9ESQAmCN
Bavsb43uMFglKT0HzebNYf59ZL1nxGvQ2RpwET4f4fVtcj4tC1hmE+6YOwpZByurDYLNlyEh08yT
z+no0cE7XNkBpuP3uAZbCKKpw5m/EFXIE2oVPBZwhCFqu5FOlCaHDUhvsDt8EUnqCQHAAb7VsQaf
EuxquWDEynhdW+HBevnQHL6bNHbbiEnxnOMfbQTiBNJECcUEi1ZwFVc/ymcgGR+NPShNkQbwGhEB
uIe59+Y42fCpo33gWOTO4xp5l4P1NG5GDK41f03TYNx5ix+D28y31GcF2uEfDVs0NONv/dEzTkTv
LWf5D69PloJFCfuRNILdndTK2O0fUXivxXjA5T2E/0C7mNB81OQPE9cb8RP9v7MpOqNyuxjgeXTC
wKko6tRgbwDcswJ+5G6nmLP3BSIJV5QBcPSuLJ/U5TkEHTKs7TyX3hm/KKL3nyrl13BGKjHbKaeG
D9AvFsqCez9kRsfqRArbg2p0MjBtjF4wYJeVQMSfIGSYPIUzCPQx5FEiqOmiVAw/bvpNAiiOqFTV
e9u42CRw/XaFXWyNiR/wfTHjslgY9Q/ip3mTZm40tg33YbridJsu/DZohkV32TfNCEFNXNcuWB59
38Pus2ynr7Z3I6BWrEqLfdwG3J8DVz0Hb8eLoA/5tj6JBub+ExO5zLGxNMxxjjrA5VFjDd3rW4ty
Bs5tXDyfvANw0YkzrmbzVKX88cT4wLfNOgRW7mQIkgj6Ydl2hKEVTToML3LJ1rxGome8PP0K91ZH
tAog+0eCfaGorAmxzRM4116MvGogsEfix///D5c+Dz76S4EfkEXQ6vxK2DWgNi23DKo9C4AVEr3G
vmP2GzWzHZpmqRQV+fx4mI8YMRYnbRLatFnKb9j0yHn85y8FXD3Aoi7YsVkIShSX40O7TapOEpBh
Z2AhssxNfTO/FDbQ1MtW3aTnojLPTK1Qk79ZUuKupJ1lHfZDHBAFgLW1SuxZa7AvRCqYgcXh3pz7
yeoJ1mw976uK5zqOL7m6V8ZFcJhKOr/rcs9S4nuvAdzON3XCVmeof33CO0Ypgwf2nkxrS+jvZ9et
aXQMsax3NDyooTP3KBVVpuReXjL2pT1taAArnAUBX6DKccysG8pgBqf86v5TS1R/uQsUcaZ1Siub
BJtGAj9h3oAYXVUisp1FHT6dcWFotjVSapNkhesiIBG8Q4SiQVC93AFoG76nYr2AfonkH4rBzecY
rvwaCb339rLUs8OBz2i5605VOme3YvE+yC6CF1mNVfi5WUUYoq1sHtjjSOegkjYZ3JWyh/ywPSFI
a8KbwmGUjXahLEIC79CQP69Bh4RSayyMdK6yaPodSzjvFelU+u4sUUq4P0to0lQVfAP987dHI7uS
dPU/zdhaxf+WsUoxslKq6UKV/90UHX+0wE5GF92Y/1Yw0M7lzGvvYmswZqNAbpNMwr9WNEXsM3QX
+G1i5xNAS4p3TEE9cBSliDuS2ehyVV6YnwPt939ozK9PhAZLaZrwKjob2JbL+56kxjBlaygFuNuD
NL/caw34YdEFeZNRKfD4Avxt4J4Zq/3X0MfZIikcMg1ilOSfYE96wrDq/J3Aqv/zgyfFmHshSWyY
z7HSIk81n8+ia75O/AW24NqCj2VHE9TvCAwBLjcMc9bdNBS5eQ+DXFOfjDvDZnHXg0gRokTYNBff
3cp15unH3BW2e90nfIXxJk01tHdveI8+k6Esq71oD0+IbN1jc4s8Bmhydsk7/uPa3WT7xQswZYqS
IrK7gP7VcsKRYVjZ2g256t68g61KRql+As1W3z5C8L5f//hHg9PNg5ArWBNh9EEQk19XfGndaYE5
nQ7qHqbIffUTpL9jZR9OJbYidEnDJI5CdojQ3+8ojS1IqBQ1fRJLiIdMhjOKej6SE/5wRlyEwqU2
PPgiJi+0twiBefLkzoseBpEZbh0rUgrd2lJSORz9Cyb7O7lP89atxxXT8jt3zZrnNdVuXdrdtSiA
unpRVpm1rQOCdwP7YlBpARC8gNX8DM+WJ1rgHS9HPCA5C3OonluHoleiNE9ZMEyS9XZ0uyEJYEzn
9gTg7BxU/Ax7D/mBKNImTy81G2Sds+XAudOV95cUzho5UE4CNksEeJSLz1GlLgposunJWoLtj5Do
wcZ9/svLsmozimZ2yOetkh7kyx23IQIsmfkjahOl8NxHUphBXd3IuqVNFLcqXmXUMjm/zj86H2BH
iNvblVeEBVZDdRUrPVOehPgxd7CHgPFoY4dir+R2/95UHMG7wmhAszj0hkUQwnoKWfD5KlDd5PKR
3lUDZydvtt47r6BTWqQB1ordNA2lBii+xOmJbtHlEgck8ziyf7jEkUzkzTd1VeIdsmEEZA8cIhMp
ifyESSAu7oBdziIOOiAyeTKTwHyo10v+ZovQyjTe5G8czmuQ4IXjnCs0Z+c7gj6UFXIWBeVdseYA
HTB7mEXqcKpcim+Qt+7+MRElZLnzCoNFhF7q8WCQG5N51cHbZjdMtKk1YGYCNYbIl+CcL+hF6+YN
3Mlth6VGXHYqwBgKSRrB4JrOQ2CBkIsK3rcs9Fu/PFrFn/xREK77Yi5++PlOPXzvvhfOTaWMeS0S
ekiEgyrM+NQtaKQtaTdS6FTWRm6qyrhr4hgxFP5PWsLqq8rgdJUd+Ttbwd89WB7yhpNXgyVa5hOL
aaI+5qYWGdrY5S6cFOHzM/JM+Ecx46wxLPsaSmKBkszVxYchiralqZuLTMwULtOQMoMK5I/Ynn/F
EZMM3gYMRRmvR7MMYPJPm8Moqr9RKOqqfqO+S5xX9K3yYLsAELJItN3ssgae26Hocr8Gy5zXZvZa
5rISOUuVXyYW62ZxNzUXcsE9tcYWNk9oPu5veTp0GMbgMEPJyf78NN73EWqPGgPFDsZOE10ivpxs
a99RyRIXcTdWtTllpjK9L2PSVhfMgttqJNn9KnX1gUYQExo2NF57MORpxGxtlm8PVwPZZqEYodpk
BDDy0/xYeitFSZ1OcYkn547AkTPWBYbNsN5J+DJ/roEVMDfvZu4AKTgj0lAX4aYfeWTrsa9myQHn
j6I1dHViQYUSWdD2lHUSfSDJsHCjgizWsKC8ZRDdM/JgwoLova7AOv5raUW3pCqf5YgcI5YhYgJg
ErjieLoEtvreY/0enkcFavujYd2QDXrTmYk6v6BuqoEgriSfn7xsJsHC9m/ovu9DM90eotj1iPyA
BM+kaon6uFNXQsSven47DNwt3CwKPVXUAtO0HjkoJR62CS7vyYgqNLRFjau+6XcCUUFd4v0CoJJs
+nHzZE697wvQo31l1lR3vmBkbyvJoTWOHkIMkVkt1ythrYfQLZgr8EdhRqZJr5nO3fZe6prhKhlT
paowYltrRYpI3BAfltHk8flWQQOb+WP+xc3teuLgyYVDXRAhYocPdg5y9Kp6fqZtIK2Dfabzzx86
q85V+5rg3RvHG4W899iiJm1jnykqlqXks8WywvW7eEA2prv+xI7YwoF31PJPnmWQBQVN+PHia4Lj
QqvG+XnWA5Es5tusw5UMo4XbCDeRpMB6t5NsBw8qZJ0f2MYjM+Qkq8Izk6hWKWU75lxagHD8yq38
cH7N4aGhC6BZ6bSzWIBaxEEjZtTmM+IgoUYCCAR3XP4SKHNF15zaRdiV8z8sQ+dVvZMZFNchfZEs
fF+RpourRlKuYjhdFoD5LIZgkiUelVrjVfajLQ4wokWBhDfRoFH3wxTV98QS+vVZEGktFeQJm4SZ
B57UccEOWgAdn0YjY9XU4p2soD1TSENV+pxDufoDeH4VG0+E6Sf6EPlSJ14s36LBAJtUMJPE5Sl/
/S0d6z6dTa3b+6WmmahQXvj690eNfUn4VmIRDUJmN3zk5iIGOvK2VGNjkd2oOGfgl1QH1tvLyysN
oMX9dySsIkhPfvtp6crRtsf8guIE1jMhFTzajMY5/VMh88TYRpaI8C2Zt2G+R6lA7lNy8kBZtCBG
r0v0unpA3sn03PtI4aRhsanT6tOuh6HYmHgi5G5CPZ9lgCpAazY4zV19S9LXGkVrvBqyIoeIVNdj
+wRVX9PrXK+YZ0k1XM4VRNm2wLkRTunZGf+ciOoG5ZqGiUL6FndjYBh80IS7mWkJsgBcJZUDee8E
oEFnDwk6ikyUaG8BhuPdYn6c1jH/6x1pW/ntTNlZxpZxmZuFHXg1rSlXAj7QDzFNTepBwlgJnTz+
pBt0JECK8n8bJk71lPzCy/8YhRf18b3wmmf4X9JE7PUVjglcorPzARYMAVjkp4Kzup76kOF3fFwS
jfQ02j/1zHsdfhd4s+ASYMyaqrgMJW0OPTsNeuVnXGnDXyiWyYPmqAzbdzeMdqQo4Jzj9FH/Bn/x
oX9inr4qxceOqM5pjhicKXNBAQnxfRXP6DDBJ6AaJLHxAOoumP+HuDbSpfnohFhuEQ2T76bZBgwc
iubZG7pmvw58DfnAya22LxbfpHhwX+KRVrnEcFpm7pqa6TxR/LYuqvHZir6HF/3qh5XT8mUgE7Ew
QIdjrUTfbKBclDXyNqL9rZSjtqH4XrkynAis154bdH9aDRg73kaBJPpRgqRLv3dVcbiWrnxmM2c1
MLE2swF7rMfb1LG6kuarLZSy5+elS0IRKbABOVpRlDd5ic9eWSvbVMyAFYtcb6Sniob75IXQu4PV
GU9b8abgJm/aJvLX1Q3lqKJN+IC23JWZltyVgp9UZF2Zx55EzgGZYvrQKJ857Vm2WgR1N/8NWJUM
VwET9ZG0sGTSZ6fMnzwXv/T6nV6Ex2Fmb947/Zsz036uKpunBDXlzpRh8KTl1LHCHod8xeUaQLk0
TdI7Jq/2fekbr9O23jeV5vuGQxfj13NMJ2WwQVosAUN9MEXcDne35aOf33SG4rT+RoDdRKeH3inb
LXlqBE6xmTB6MGeIqA0fM0qrJ+feNA+/nEOLCFUvCdf+lj3BnC0ethhwKpr66OvC/SSOd0Ij+lPd
kVbbOpEj9gi5bucZNa5iGgke0hOjV7+q92IH2gE/2gqEKkmQ81kBJJA3Vs/OPiWxgU3smT3SoT7x
gqVAhP+5mwzLDHnR37Qud+qwonuY7uiCkjN771iGMEFhBz9gruW2U85KVK+ZteYB9yd1kds0P58k
iWysjumoC/B7icvz8Q8Y7NkIauV1/pHlqQeOF6CjCBTQex52AeRMMV3+1b1aN7RXaB6deZQMwBxe
2bM7S8bqo4SiwSm+jxFOM/CwjG2T5Dwfar3qEee9fgPfw+qX+5gkL5sYoKgF1Zug7iX7A+mPgxiq
5H7v3QWNV062pb/sURVrJEzymFELlFePGUoMxooQJoMaV6uWQ+2KFzZvqW3l6YfmDd4LtZSTKc2A
hfn9qXcx8owt96/AHtL9CAu07LW5+JmIiIPVdI/Gmx3a6kLct73GXdFV+CCkQJC2uBZtqvOjXaHC
UCTqTgTypKaAnxS8y2oVBDKThFzF0Tsl7J3vXP6topiZIQ58ui9e6BvjB+v9dV8zKnlVI/Wr+trk
MmZkYo4ZKK2NK//P5x71XBEKDn/WyPSHad+V5IRt9gx8wkLJdRLlBA2TY6PiZAYEsL7aFi14c7vQ
MI58gjZaqeGA/l54dC0QbgNj8oaD7Q6kUaw1lUGyb1J6+X7LtJhgUPbYI5FXvQ5Btw5fMxTF3vE7
rXwzY4hfQ2k9YRZsB59bHjfxcwlK9G3PGcjIfNDvVyxhQXvaOJuBEs46oCJ00XedWbHVY4s5Q6Uc
eBw/S64R8hog4/dK72Po3zwAoZh0YODCEtNI/+ak3xBeUnG3dBeczNc43gZTHF2sa07W9WunTaIN
L6aIKzQcqowYNVT1WSwPzakA9r3HoHulZ1MMc1/xoJ1ln7E4YGprPu81YquhLLcY78rdE8t0xMFu
PRymW//MdJoBXvjupw2nk9FJG3VpZ1HLqO2gvbf7uhu2OFA8M+QTfz2JRgDXHJg+9/BNjK6FdQL6
oKTdI6zwVG7jVMlyL8XIWeTqajoEkaHlwBBHKq8mIl/gvmmJPjdJBNpTceS1aI1Xt//bOI72cjCJ
oCb/qR6sf50zKUfSDIIJlos79qbTJi4kgtbGENA+b+8iG/Tmv7QMZh/+9JngH0D1hVyOSBZw3cLV
ZKefHcYQLsC4SCHua/UhfCUgDAI86dzOPPWNFj/sA4McoAdPfRV0FAWO1eHat/ULYIisGo42AEmZ
uPY24lzuKLlPzVZTvwcQhV+zZsIbaZ3l1rP3E4JiLnQM0ROwV3RDN/sgtDrn2MfS65CQg7vWlEGI
Zzow6qTSIM+J6IvfDI03xkZU7LHkMj2+v1vQTy9MpByKFMFWmiVbMhOou84fVL4cHkqe9URHbUFF
IxDd0WbNltbuEfZphQl/TeL6i7kIOs9CSA3A/Vz6501keaC7VBsq1jbSSNMV6tcuLKOnBi2N56C1
hz8F4RahRMgzyX5MncJiIKghc6oQBKrhKkRt706pjRZ1iadSFaY3cGPFF9i948yOnaB+8pnACpzq
OnpA8nBdCMLtL7eHtxkP5G/OT9dOi4Ar7e8BFRTFoU5uBRCjtMTJrZJatV1b6ymaLFnCvb6cGoQ6
pztr6/dc6IkdW4G/VnUh4diYAFAoYUh+TnrQzR4UnpCzuh16kpAf4/edSgJYQaL/VqbNTV3UkQxK
odw/oWSd9YlZMw6Yl5HJpT9bcJA8IPcT7lI4AMITPW3ttO2J17kqUfe5XA96hhNsEbzsSB7YmzXO
uX7J++ZANhcdy6pqyoECLy67D8z/H6BL2V+LEQaevukH3yLx3PGF/mh2Zz+XKVOxULRRzHtNz2a6
sXLxfpZ6jl+B9vxvYZZH9tBpS5qM1pddiKxwL+L2x3Po2uWWzKH/I5eptEjiBOooJclDg0I6nnlO
rjZUb+XuyZb+KBmosHH0u0CY++1GaPCKRBzHXC+U/gtmrdXlsdoLHLVtyG/ArQKmNzKw25w/zzNG
lIjQo9jy9gITSArTaT4GBc7YqDGAs4REzhPhK3v3nEL4fP07tM90aQcq+ZxwZoe1gJOeOp+vY4R6
k3qL94ihVS9dWKb0j717pLpCmKe0hJ8WB+PShLf0DXUBrkz9n9uy39ZP9qbtQHdiX2+CygCu6Fah
VuvYoPlIWkWGoxvR52m9oygSozuGITeNWp0xZ2CrlVGwKXhXHz5sGcO9P54whXB7kYfybA9W9u5G
0nx+uALuUUWbJv8JzXl0JsMPG6VAFZ7g/aTEG3q+trdUgqsEAq5xM8cVf/onTi7jLkpMYVFQXmHF
LUw8ZlzkZM79r1HbSOeaugAR0guxFSH9OjRRiBEwhFiC1O+6RE1+2xXtPmP3PSCMD6Tpab6SwNL9
Tpm01Qm4QrbAqn5plLZbwf6JBG+NFXmseKOdn2X7ACA7rg9lSriVf5XRUh1lZvVTRG/mMuhwFaNz
a6CcnlpY5upjXzQYaJIQGfahtPVrSjTjlpgWQPOuscmG/KB8okQi0YE4WAL55Ifo5++KjZoel/wg
mHp2+FaXc5mUX+F/7nY8nRiuYxb6ag49Xo4zjV6lyCk22TNrGqEn83Cz7AGV2NEYPXyo//Bm0ofQ
S2NkdPTNnuHbOwXammWoBAsvgTZyIoAE2Y9Y48MugFg09As22P1fED2WdCP2o7sco6nCJkujsqa/
sJdJk733G+GyJ3Sumgg2VZ9hODMUal3iJ6zgoseOiKBHbfME4rz8u41p1tgDLM/85ZfXRJ9PuU8Y
aoEOgSWsAiRvZbb0XKh7+7okuRo5cxecXthevyM99TdeEkFOvvrk9G0YnljeYryINfIxezxh1WjZ
hQKal+SVFnspJdcqDixW7mQXu0WPWQHtXMu8tRlUDkz6NJNMHKG+kyoOq9oluV/wckHnwHyNCwaS
Q1KKMHTAgfpB4DctBfvVSduiLhoOdvMJWCIA8J8Ydqw72Vtzf4Hu+jjO64uBFw9JjS7Qk+1970Le
lWq55eZTJxKsoNsUChqdXvaucRZaHFXe3xXVuGFWnm0ibBekcUaTWabtSvkjJXMOCwhdG5U92YDq
OfvcVpONJAs986uEaoI3PiDNeSpsz/uMgz8FkiCKgsqh8w/hovE0hzKB/4uYHX0mB9INvZ1Y84uF
IActYWaOmGCbnND+xPLTTb8PotyqZ8U8L46BWrSsWUsbc8ybr+F6ORSdvXyj47rZWRuPvUfvwYEf
x29r1Y5EPRvQNBwRXxej8N/DHI2Wk1xN/J04UQ/czLwIT1GUuFqa7b02j/Isn0SRlPP967tvIzW6
chSwRB2E8p49q6fEJzU5xZBvpNTaeBkheK/9hos3RPq3uOKwDLwUqOdIeWTbUmZaxU/qLhsxBcbi
Puq0zZEPmWfApvCiZWFQzK+Wfo3q0knCn7OUEDiFSZtz9PVRxXejKB57Z74liAa6kjgbdwvBLPfC
cJy+8ZEPBDGFIiJWXUAJISAvpi10Va6VCaI+WubCVFpgaFr9C9wCKXoiXnrvHKYR5d+qabonZu7r
sYbres3rHWIBWq0jyjH2fC7DbZlVi/BNeJG+2tXgggy3MQ0Q3z9BFIL3mF5F7paBPKGIGtn5CUj3
e2ItMDqEXUdhEpuk25wA7sIJlc9kxwFHraqb7ZB2g34u2kMWOm1mTT6pg7mdTSdqRQL51zqsBxgJ
1f/QlpKgUT4+QRevNRayT5mB/czRAY0kGhHhc3WL7/VwhldKn5grzozaDKDKS0IAMW2vkuQ+F85f
CuejRDN89YiplXWZnY2+GYVUAs9VRhsw3ZsB/t5Y4NuZdr522+7dfFC1WM5IePfDCeuZJ5XARwgW
EUH8G5BtXXU7rdzAl3G5w5ryH0yzjhF2GIJRvDJ6bsgyfHiz8VVZ06/xCEHaldp0N4zaNXU6gKFd
w5knoD3zBq+PYxHa5lpkBlrCAE+Np1E9MVTm8UEp44R+oC/FNIiRtYG0FLjsBXG0CsJo7ztzlfy5
1OKdGgH2jzs2QXosfuaMLsU5sGax4yZyWiQXNQYhRZBo34mm+dKb+zzERXjQpxB8Ft7BblKywtYR
4TLcxjDx1L8EdJNP6JTeIA/k3/1oy7eViNfni4QM78t4YBTSXoekTt3JJcKfsojSgpuXkTx1gPIH
A/PqTcbacjRna5pGDhAhzCYU6LL7+rPAn1D7onYobhAQmEj+abzpx53ojpq2JnfLn/FZxSUEKrrb
bQrFXOX58QyT5DTUD4vf2TE406TDcuwSNPzU7hecN0RIRKVdMzq3dm9LXvdz6u+FJ3rRB043VrQo
NbRdY7ADSxTJl/LEH692Q4N5Ybim7BnBNTDzZiGgJxgwFPk9zWvDDlgdD3vZXHmotQ/D9iwPVjGC
30w73RW8t7AwN3tfiUmVnOZDyy+j/GyGouaKzXskkSMtBu73WwRaJHb+aLKi3YNXoRNf1ma24UX1
3V8Ks0+qjY9H5traAK36GHiXaWe7sL1f9lCbQD/rKPzAVkfqPoKZrVviH8SscdH7cAGIR93e+Nt/
+dmp/k7gmGtYjBTwAQySWO5bWzqPn4RBkNkI0OqKeGH1ysTxQB2qd3lDGdm4KORiK68CmoTlOFwn
JeuxxPkwU4kuCeY+34T02pg9wbf/sjRIUPM2k2jCSDe1jpvGs+T98/U39m7vNyeqi8gz17nD9g7F
rUFtA0vzQQo4NUliv87FYWBUGxZHj/6lR8vmY4KGXcW3rCSUyng3cONshnaHxYgdQqvK/TWYGnlg
BGO5oKfMokGatP+phXHIa5d9DSVHHlWRDtSOsz3exKfcEocopu99d4A1+uWlma5MDgYqMubzFsy/
zhsArMyjQxeTDZKCMDgPnk0xxLay3WRSgrAcHOG1gd6Xk+W/MZJQMts7w6Wydpztq8oT+K8ZyUk7
jlUv7kH7mg8RDS5W7IohRJyyt7AqP3UPJ4WCv9YjpQuk1/KjVf7Cw1Xbv8MTW3T/TXfE1oWZi0c3
84iGg6BiZdKIW/qWVmm7hL4jE/6gHJFpr7U9E1vof/ZsB0lqpBXRNJE1dzOFSS45/bDk+mEsyx1u
vzJoftkZKxWiTXC8DWyRRfMoJ8mEACv78YR4xXFryPX/SjXPFX/CD9O4VLDuDyMggHzSMsdxmeY1
CBRnP4kBPazHVIDZLkZljWnZIou3Ip8Q+A6iigwQlpncqn+fTdGHHrwqOpktvisd4YLU3SGXQ817
IErsTtWw7diH7URWWqnpMv043w8QL//MmzQSlf6UvHocaXsSdqCtRNfm2p3c91D3ArFC4uaT4Kbp
tFotiuLNDw2SPE6e7aJt2zlYwJzyelfUIiQSvRonQe/4S8rGkujXTA6VLBB8B6BXFE6WmC9hesSu
aeYhHNB4Z10KMPfATmthIXFVHsp2Dg5zM5ZkFeDm1ofmAnYtWhdx1AvtGiUm5wMjGa5H91/5kOf0
KSItVsr48ElR9lWBEqmHyNUL03QwUv8mPT0A0ymiU4c9yFX9eCsEhaeNykkay4d9moY7oqy2WfxZ
zvzj60BIw6CA9OYjjS4Ofm7IeXKijFj2GV1RJXg2qpTz/FalGuYFCPEAYfaTgQs1yau2eO3GtZ1r
lfVkmRzR3SJgPz8oaygqMX1JvDfX/OBOURG9fk4qre1NbE5oVs37C8e/LzJ+Ak6QAlJqCB9rHWiX
Rqd93TeJZ1YXln5gzreSv294dCoqp476L4Y7xVMSVVh1pS4HOoUB8jd0gopmLxQEo08OYbKqY3kF
f57azLRSdrGoYeX07mON87eP8xv0/ArSCvRqHIB6V6ybPT0B85epDV2dw9IwxM+BRF5sDHRpcfSl
FiBZLl263braZLhZrnv5SneS6GhvwuEr1vLnViryLnUYMpPnhlWkkFOBtoRyzqDZI0mVO0DO9Jv9
CiZwEXTbw6JdbEGFoG17BAW3rc13ktMWUq6Mv6ntTzpfl8PWTJdl/1hA753lwaTXXGbzsRCJZtBb
l0ZF/Zi4k4ik3SrwKktyDKQ3p3W/XHFBbDjfzWLTWun5wYSpb0/i6WXiwjCFj/gDu9EWGV5CzVul
YsGDvMtFrmBd4Mzaz29d2T12jOZAkhEpuwOHW28PaLnmBkPAX2B4T8yU69hCH/8oWJb2N3SAc7Xg
FXbxAPJZrdENsZuWXIwglXVImvWN++YskEFB7qAFLd2RtsKU9xiJhcQb5/tUzkGJYqZNsAi+GpkW
JbndkRsJ+5prm1cz/ThQ9ciRhWcD4Z7imckpybPxhSWDiZL1z1oU7QgXGXukWkfEG9/be6NSwwCd
YRhZfQbL/ypLKmmkAC4QDhJ1a8QVGlJZ3zRNKxLT69OB+WjxyYmqM16li2EcG+pr4wKyvBPB0tQF
cT6lYzhq4HsEurIlDFLRj40DhvX6Dd306uim3vxjCAW0E6HhnODEuC7pMKgLZ1anIA5TDCX9jIOY
uh8CchZhQr0fo8WCVBG3ylJeyVXGu8x1Evdsl0UKqIXLSHmMN9WefZTHIcL3VJYJJ/KEQ74En3pJ
TPzDl1b9hvSG5K0jParnjpvir/hi5diaQbLeSYCxM4XixWaJVDCTmQx0xUtvpAwmhaLShOWV8zl6
Kc+OKGmboBNX34039WREKKGJuhZc7d0c2WCnasM9JsHpVtXaj2AR1oGgv+tEpWuXSd9Q4p1D2Xm2
gtrlAuJTqWz5U6H+qjUgKQiFEn1jeGE2921xsgduAs7DtINE+tXpkZFuxoWnYOOiojvp9+ii2YA+
LdngrBbXR06AGhO8P7FNNgXSpzG2SJR26mR0vhmE2KYrOIt7Q+8hV+Niha13XqzeVWBSin6KwlSN
8YPxQneOOs5Fk1BAs+zWWJRrqdu/UJvgL43hAN2eZ4z7bjAOTD0TXrlJmou3JlumC2uMgka8ma7L
Ndp7Jjp8ksKxn3HPkwjl070dr9/xWsQCzHKLKmK87zZYOSLv6HDt1eO3scBZTUBMmFX18Mk2J2Hd
W+ChIqJOQklNFCuFWkt+JNLmqMM22I6InUTj5xztwQMrTWt9+6WG77/kV5NUnazuKziulVJmOZVe
atUNu1QYYS7RwiSddSzYPfsxSph8ptJyt8aepcpOq3YeDPzfRzuGUUndIXlZBDN4HX2+Un0sfnHP
RW4+vmXAPeoGOZ5S+5LtIrxw34RCq2xXyijHkxFqksZgyYA+Mi81r0dUr7EOX/AdKOqnSGm1R2iU
D6vHPC5+n1Vt58P7vLv1BJKNiwrtufV6ZtxidlP9dO8gRO+l8iToNnVb9xNG1TQxwLtZ4ipPHP/Z
Oy1z9lAspU+uxjqyufovhI+tsbzMBn9c3nkPpqOiy5RVtWZwvdJvi5l5lub98e/XyrAImqdjSh72
XMF51Y0dEXvWaFS/lymmQ9TCjBn2ay5tQkMFk/RJVqy8yfvlGkE38dujrJ/HHKYmvn1LDRuosw0g
PkLrSh7FHcvM88Lyn624ZHwz7Owa2zB8NW/ok9SEGSvpB/LG6G6uxrq7RljdnZxkCS8Gxi41ymJA
kWWje7GYGKLIN+4eULIgjojnmlYYlzHXBYpJft142gpT42gzR+kJT6WbJrUHO63NCGmfrisGc5AG
C48uPg8VGca91eamW4xeB1XyEo2IHqhA+9TYkeP/VGqJMlzqD7KIzw4hWmGYNsR9+TekZVNAB2uW
HF/2W1xg8cZ4nDvlgYqmDrZtkph9QZmS5Xgm1iIfvvPLIrVRXqKxC21QdmWvAfhQicPisDacRs0S
Pl4nC2CzCYO2vrHONWunCtCF/9z4xWBa/flTiXGB/ybLmPaRSN0dozamu1GAB71mRL9a6mYA4TBh
gAUrtJpdel78BP2UD7nQOhRjqkWLM9WT+RGANOwI3cT/3xy+LgfsQDr8b0Pm55N7kySYTIgVHGud
hjFzq8s4b5Z7of5/80tPZbMmo62l4fpVvyITDLZ993zYGLpcufjGbdGBOVRWrgbuti27ZO8++e+D
9Ybb0dRPjE0UKbhm7Z5Am2iABUv6IHEs2s5niACd/FFSy/P4FQtcfOF3dPfBg9Jx60aQhkbQkLGp
PjPrrIm1TReJWjQmwJRyeRAWQmvcPttZ+eoLeOyxF92AJrRZgnrwMuOwzoDDl9bCkje3PMq9MwMK
HSNeWU1sZV1YuxFouKUejw/9FipciCwTMs1f+kWKZIZvATxehViqGfeKQ4CuWeBcqExfiYKbeEdO
LE1PyNlq4GZfcnVd9B05VkfXMcgGYxx9xo8L4HluiNluiWIyBd/mV5ZeC5NX9vxMlmO5aKaosH+z
amhr3DeZf8Z7C5dfbIMFvHtfuUB9xt9aWVuw3aOyEWODomqJ30GPf0JUCwZ/eNf/7WR84mMH4Tc9
XGb4syzXdy0dcu80zo0Hsf5HDhnESDgO7SSPSrym7e+nf7KGvHb6dciCBfmPbnvU/VxapT1VaFvU
ec54ZhR96AYLuSm8LEieUJ3pxSoOL39vUw3+PHSEs5KmBi5T55ZGFsHNxfqQbYmOb8NDzZ40brKR
u0pJLvUskbbQThxlHl2lny3cT/eBh80uhVbaf5lwLIO+r8DqSwoLecGHCIKvqaMKzuf9XHVjM691
8xn2stU4QnaaWe9KqLtl4LI0cK+IGJt2TCB8rme5qFXT84cN2FiQdTerxW3k0kB6o3ejWY2Oqy0a
F4pmt+fix2hH9I1oioO1zccaERzIPaeVGWVnMOi7kTdTpDbjuN3U+sm1xOFLmgVAZ/Ysar6Kx1T4
2pMELrXTGPYVctfzBjsiaS0tvsOn/94Id/MsB2XW7Gc4P/gamSUDNrCur7rUvpiP8s0cAbNQJDtQ
1dVstgLlRFLiXkJdSaMRkYsR4SryT7goTjY+Lu4W5eHbsx2ZNbD87wJqIAIMHdsAsAjTnK3LGn94
dNs+RmbhYwHYUzKVEGPt9xcQlRYDHfFzCmkc7q6YLbrCprJuevnrZOYtV3vNJArg+R6eBJd7ec0o
+gpOzAHo9zP2u1KKW0rhoC8XeL22mSGyVyY8NWqqBGp/fBI9j9ne3wNt8IlxCAVmlV9frUrbwWm0
mKBwMthar36b1q7SK/tUM1ccdccsg3R9w3xCHKjiLE7smG6p5THbQMhc0IbTLCgpXDi6mBBQFe4j
T6DqjJu68oe591Q1eMMsog9dDIMetUrw6G20QU0oXVMLAj52fwvvfQpd/0SjjOUgvwzDjFHf12Gg
dmBSKl+kt+sNe9tabrB1qu6jSO7ksgL3E38BDg+AQkU4TVLg/Nk9HMbVHI8497m12BhqhDNno6L8
duLSLohzSwER6jopr1azA4eAP5F72hLbJvlbnNjXUuwSdiQKx7i3XYmMsZsERArnJIhrxbq8sgAy
FxrLgqWszexDrGLNJNd9W6fsTaijLVeJW5QssnKTj6EIf/lZULrYMI3LxkYwoUvt1kY8X4hvuURq
bVi0pV+6PBTryjKPk20xOUasRDpbGCFuvDKyEU0mj8SmToGHoxUxeSpLwOfyZ7KJrpPDr8RNUqtO
me1QGwL8kLAbpEvXeOs1qkezASLntT8xDDYu9z2NtBgyREhYfkNWp38hygQHwjuePXP/LKppOedz
oVSyT2nCjep4ZlZqS4Keh6Nt7SqJa0f4yaac/XkY2/6OAO5KAI4rNrcwfqJdYyx+7HhF1hN2Kop6
E1XGgYZOWpFy9E5Ro834XqS0OkzwSRE+vtHIOQwmC0Ft9mmXnFHXZdwDeK7VSeNbuDzfIZ69Y0Bg
BczrASEPId2qyYFYCGk/EonNrI153oM0wfVciEzx3MK89CZdCGS3SYYpEWJbXbmwdQujGU59pDsh
++3sREQnXu8QzJUUSMBTdirvyAmnMsP1slcHZ7dUwIH49Wn1BKFpPRoVStVIxoWnAwIJQHL5CfAv
foD1KNn8JXsiMVXXTngB+28WJvEnRoOTPgoypvcrZl6Y9dAGigMJCY2YuhS+HSbW9b5uujUJ9745
syEHkcXHvZUwfPb/bNL4U+PHb1XcR/XhdtKAFy/NFn7rD5slS6kXF6oEz6RWK0xjB6A1qsuXmhKs
G52noUltBBHOo8HpeoyygzlGt8jmHZWLmZRxz5D/DtVZ+qxZ50LHXWCA2FhDZEuN4mwS7IoTZ9C/
uEFEEvJ1iNTwHDa3AHHmSRHfhh/3ZI0BZR+zRH44hzUzWuTpWV7nyJ5KVMfclLadgacVwx911hgc
7aib6IcULaCrlr7YG9356Dk6bo2fsnxvpGRR1z+kFasQ6JtfxKxGC3BpjliMQzr6ijWiU7mw8fMU
GyD4UMUy1UGdQiIvvNkd+AvKerM5I3JdzII/xeFkHL6JGwRHU/WW3oaX7/+crflrXNjCdYy+2J31
/XEq/ECpbOSmQrRprvNpciN/H1JT1iC04IochmPgUCI15IyX3tIuU18Aaxa2jPBghXfpBtsiNV42
Z39fGa8h9F8bRE5VwP9pp4U5J6PSy87j5/kpUavu9qNqyh1bN4z/9K0iP86PB6TTQt/8NJQ87Pqh
7TOWfbJp04YJKpy+Lc5tRVj2hBAO9M5cFGXScTY0rML0dIUu/JQ4gi8G89+8wbvRkBiq7Tr/rt7J
bQ7cNGbDOM/DSYsA/YrEyAMbUmv3LZq1pLy6/ko84WdMoRJ/qvrcvGYu9CZEZO0e2Upnuxq3Yzl1
KXDy0AbmQKQi/g6pksDsLN71sIVZ9Pw/GiOoN4NGjSreeO4o98pDq22ocZ+pivhLguu+yhNrUZs2
Bd71nZf5v/Y1hZt833ZmxIbDML7tqCIrRjVBCglp3IHnwdRSjNzZD4B38GnRSgptz2iF7I8OueBl
kOLiGKzOJyr/Zd1oPi9zSKT4BPhmzzLeQf0hMLZXsTBvpoDFx0F3syvSSahS6ylE7vhs21KacAWN
qB9zpaB8O4nlkeewYLmShMU9wBHBS5jbeqba5PYn2xBfWNVNmuqZHAQ8rDO/DnbcblWI2KlBCEJi
k6WNqNK1DCFF4daQs/zPDwD/U0eKHG8RAVZbJ+rtWOBQt0I9WuYsvCyai/RB6t6mKctT79YEHx5Y
kv4DpZOaybFUBmfUnqcDDEDiiMh1gBnoBWYVbhTfNmYhR3Haj8Bm7TluEj6Cy1HqkLa3RsegAUS1
Vids/JbsgiiWoPBHS4pLJWuSjUdXOPQ0YyOMIYYtBjy2cLxtfDLEGY85tC0RMxL1IN7l8968H9LF
TiOw77reIkggxtsa1DKgzlM9g4H1hZXQcYCCb1MgbQDyuTvU4Xq0mOTqXYBEV3I7JGwzn1udqtfL
ZgaJ/cKBJ/MZaDN7KQoxLCE8bgxI6BfG8WG3nIcKtuZz0LBSLuIJ5Pekg8uVjgUCn5Yewf1oIrxw
01rs0ChEfybCzETwQXp1nwKpIHfdv4tUK1vlTzFqpmotqvd4+mAntbgytnyMC+XDT2UlguuTd6a3
B0df7u7nId+K8nf/lZ2zxilN3WDSCW/QjbU+c6tUOjuwiA0/vew2kfrem3rggH4dXpHba+B/JZEd
70GU6ANKMxlj50GPkhy06zK4HM1LIe0ZIBqnIyvU27j8hLY9SO+wK58yJl9GWMeSB4E6F24IXBN1
vJ0aVa/SzKh7i6QfVgathwHj/gAZ4OFc83lLcwIjmreQmaLer/G9D11BXAcQkfdKumhZkeuvZguo
YvUGmEzO6hfivL6CIC6a8xcZT7TCm/nD0VSQa8XfKG91ygwDgDBfPxiWAc4FLhozGVEN2ostL8Sx
cmAqY8AcWvD8J1cgZpWHN7NcO/rSPI+lU1JRk/ymJxCvXh87eK9/vSCcDu+m4W73mkeUkOMzre6K
Yj9vFEC822b62uVRse/S3a92cyb1WJzq8PzeyB9aqj4Z7os4FA9/4kpO3vgSX5Ixejl6mpiZRoyY
COBwYm8o0M3QN9FeJF9uFaihVyEJfjMbYuhJmW5uDQYiK/yYM00t4NqqSq2wh4195DDlqHzt8lUL
/JDWhaZnCwMfV+izwsVikr7lpEzBpwgvzrs435MPK5NrODXpUISSdUSpkARj8uFe8XUR0666nn/t
QKHcvWULqbTN7KewnfRuV8SuuvwpDoC+MJmkoN7bRdh1t3lQLKMwnBIGVhClPqeoLsgvLq21tqs+
g2SVmN25sClN9hV7BnxtxXaPzQguugG5xElW2ibZtf/ENveMu9CC0G22Au/m69woTDIpJHtApa3V
yr7PhkSpeBE6GXiAqRIKCVu+eVK6H7uUcM/oRzB3v2qjUseCFn3DaFndwLKra2sjm0tobPxlIYNn
rV0j9Nf3qX3ylDRX6yu4HtadKLqRCImQPrJjWGCGrOefhC6ehaiCPCMnJG17avAxchzhohvX2dxl
pTmElT8cYofIKop9gQz7N8QAlcwp+R9+HbDje5vpCBeoQPOhIsZuLVFyYmw8zkuwR3KjTrR725uw
/ScQyyiI0LJpYsx1/hXmgL6LnQkQzos1iofFa04XgywoQziVeIETfAe88Xbzhkr9Sw5BsEU340in
CRLZzW/1YAW2Ljaoq6B0SouHkYgnQxF/TqofA1a/cqG8foAgL2zQC67KXPcY9/i681TBW/EsjDge
xlslueBRzEcIouqP3uH5mkp8dB+orOLQko4fnMbpvgHAsX6EYY8stOwin5UQYWtU2QxHaN45EJkQ
8aPccCVXsAfMH6+lkYgnDfZdbm9S1Dwj6Wj9Em4VCNiX7UeaHAIXrDbLlpBx9F1cVCBI5nEKU+wM
5Wb1BUG8WKYpiZuqpE+5h/JOWCvGGYxPosVcDmC6VGionwoZZjkdPoB7Ni0qZ/RoupI4E1ouytVm
C6Nc5gd6HQEthteiWDr5mlVFMchVzvEjEZF7SyxTjpgRxVh7E4+cSCPi9iBaXBlJU1EfMRzBduC2
Eh4zZK4Telr4pDsXVHtNxBIxgcwfjg4DBQQXJ03vr4b70oRTv8VCt/h4/2HyPyO7Wm7xknIqoosZ
jw+RUvpPvRNV1Suq8Yza42OwEUS69oSBQlNzgypvt/s2l2W8XyTRrwMsC6CuVyV0JY6EV0YQ1Hmp
wGft19kU12KG1oaKUBhPgxCb0SbcCSabD0ocphXwVP7+SEgAJE9N2becJYAP7aSy0APyIknrnGmM
PJNnU1h03MoAJqXUkl+g8bFkUQtqwAI2Sx8yd1kzU/FvygZCQfw758/1CyVOi1S6u4fwWxOHIN9+
ppBX3q0z42dmQxkvU49CY7m5aJJInvx8TILi1EWBwWZxk+bK35n8kO4+iHf/k3caZbPZgMuCNQGG
UPN9M6+nWqryqjRxXcookI3Ckx28GmRjQVD0yhSb80IBofIzgdjiSO3IMtJDjKmHpLXi6BirwWY8
HYvmBIXt/CLIlgVOuL9GdJWeOG0YLnyEeS3pLQdf+GfmgLDPJABd8md4pYCYdP5O8Eaa2gCjenqv
lLY+56bIbkAsatVV3CzXY3ptO02htzVdb+M355URKSCcvkKiO63kwE58YNvegQLWtckkUm9JYc0g
00Hx6e9mzjWFo8DfyuqyzFjk88ydIO/dOY6tbdqUAGjv/Pt7tQgjYQ13SCgYMlG5N3VysRULgvk4
amgoP2zB+k9NKeEQ+QxrvKRY+Qr2hIv6ggVuqaCIwFDJXp7nkn50jfZPLPgf17V4x4EXwxaNHIJr
DcQOKL1wug2pvxtM5fuAGTToEM2zwP7aez9OXwnAyfJNk9L3qtsdCN2gJuEb9guF/BjgevrGYvh1
UFPh832GqoXpJOjo6PG/FFYJpNt5OfHUz778Hyt2ix2u+PdEcpq8fMR58S9PiC3ZNn6jsJH4CFgN
q5E/iOG/PzQ+97AKJPWodk9H+Q4JX0oKGVTg4H+ozc5no/WCYRBe7U53CXE9DfFvLOBGv0BYmRgh
IY07pr4WGEYHWAH2mlf66YTXoNB46qHsemr/taLWU6IukNC6G8c3rYmAO5Frh2GfSf7VFqMOlpWk
LTGceXjP7gW9jLmomFocx04dhpoFRp3n5fW4DZ2ouXndpr23rNhGzJ6sRuoTy90/EEngBUs7Th5F
QVyrf3K6ugg4xOZqokaFx4cFiPPwQnOWBX3cB24HhlJ1reIET4UudYVn9UbjkEH6lVsSjU8Q49sT
LCpqhdA794JkJoSktp7bhh1Q6wImqCt+MpMkqn/659yWoNjwuYkOxOGIDa4rj54QuRiUqkKGBAu3
cEZj3wcOM6b0ar4OcObYNEqk8lft2rZHSbYmNOT+vdCfi6YR6acZwndGKhqsN4MOzTSroYvGAbH+
YczslW85rFFygjLVm0Q5T87fmQ1xo2OLboOc/r09JWw+i244M1ghiR2Kh3+yfunfjzIrI6KWcQiI
l7RL0+gMvGdOV99YaURV8Zvl83LwDkI2CEAauQsR1zZUAr/oZRwrIHYdcp3NWpnio80NVY/F0hc8
8FmPJeZC2moBBaDzsZN+DARw3s+5aw8LfwO4wHYuT7JGGfOF7oSYk0z50v1n12GJOqliRlKvN+9Q
yDslrpvN1rPfpnhoYPTQ6M35H8MvyDIWsopk0661DlPO3/662cHxrWZvF7VgvNRZvggIl4vD1T6Z
5gp2ICMtsLAbhRF9aPKYmY9BUjT9hK4l6t27sAsFSZ6l0biih5mjeFPy9VPA+sVnk49SFMyzsyAn
LTA0Rdz6sUFzRz4GOXEQohRghLUPyKzMH/7pz6muA1bvhYRAIyLpt0BqRcPBbAuseJCraq++mPln
ER+myYzZ9CoH+IqVH9xcHmTixkwgmWBucV1iSysn+Qlr9ijDAVYc31EWdpKA7aKaXoMMyWKo8/MO
0sropBHR3NCidtsM9wi5nODPzbjrtwMIXN5OSN3j04Lc+3ndDVBiso9yKzyacqz/A/ob0TY+Y1iq
oDA5VR8Iqr/cliUj0zfKw0t5IK7k0xqMnVTfHuWYX5FgVVwfDPls5GueZJJAhPHbP2/YMNuakOiK
GX3Org2jg/ZQ0/poYkPaknwuf8pTj34JGyifOyvkl5e3cTlA/+vjgTXgoieFcl8S2uh9JSa0yafh
loh2R9UfbJdS0y5I5kNH73rzUebSHlzGyFyb/zemMjXwP+LOUk+gJ8rcDNK4snN2CI1SuLgDhJga
A+nYj3pbyBFs9HdCmBMBrcbFsEgedkHf1jfpuWeEVFNjUFWlOfS8/2HeCQa8BIQ31fEyTZQ/z/qL
nvkW763ON1+MMvdtMyel43HU2Kd54mKN2+q7XLlYlxoNP7The4+8akX5wDNonzknbLw0zvX2MVw+
EmWikE8L1m9q6dtufwbVdOhzyN3ivszkFJ3nilHCUIXajmMgOot5zSvqWC0unkGolgHODGEahYXn
cVYElBfyC6HeFPaULTqJjwB++lPURU46kHLoV6GK0qxfGIiCVLP9s7rjmwiGdSk/tE7ZokIZWpfR
HLuZbDVe+6HKMR16AXQH8tEq1pd4nbMq3EORnz7jlPt06HMyUyaR3re8bxjdTr5oRKVx2bucRv9j
Zm2rPQBvsa/ughpODjhJsqdF7CUSwjq5gtTNRWn0qQMlKUEe8pFMXoeHJPKpHF4I5dLkiM/442Wx
zKexR0jVevbuYqMQDi/82dT+4wTpnW06hzNQXZV5bZsV6qDxm3JFzucpf4fqzWMuOCjJub7EBUKW
ZMqQ2b+6mhlwqX2BywLtdIk+xWVocZrsQHhmp8ffftI0ZSmXEwA8/I3s+mYTVPCxt68mu3iqRQDz
6O4/OYZFTqEQ8WatVeGiTC9sNOD/9ux4swju1R1xATMo87mDO9CaCdB1oLzdklIQEqNu5UjKDOMf
8NoFR6b0Mv/FssVa3ORC9Dsk2HxQ3tAEjlo5skHKNDyJInsocyyxfNhRpAIGMGc1bYDKsgfl+QCP
CBXXLUZ3BMQSQNcU8e3s6S2S99COKr+MpuZpGYc/TznvMIGhY4LjmJnnJwlkUn6Z4PNWhLLemzrb
bQEOV5iRpA83AuQswEXWye1gB8nZpdtoik1XrgfoBIt1yML5z99fAxvxQXB7eXVCqH8jM3wTDzVa
DnhKFjm2a2lnL7o5vckEI2KHJjGSF5871dWnHTefzaL7gXBhz+dva2xdL1EtUDpZ1wXXgfq/MTX2
Hr5b8FmpwbK5Stfj1Q/Lm0/5vlYjcns7W6QeAFgPp2iUc6x5RLNKPEjcouK3zthZ2gBtNRQK0AD1
+44Xq8Q3Er2PoWBDY9Afjkh2kzxH7WNbhIAbWm7sQGRrOxjW64rxZtP3lHkhXBJQPOOnQ9j1f6cx
au0FZ5PaFdvurODPs6BEIUxqJUoy2S1fw98KpHwyiGw8+RczZjaVrXglMkqJDAuBR/l+74v8wbxb
27BKcbHQAHxG29RJbTn1fjIj2b/qXffcecmHaKyVObgiL0enEqPOuLQV/TiJOVe+KRb0qOQv08Dz
9S9C3ydi366F78BQWmIK/iskcn5HipgYtOznNpJkO95Ow1x0H5BiLUzHUCjIHRmoq4ujKRZwPJGI
GWE5HHGuWSBw+N56qgCd3QVjFuucsD1Bpn0pOo6MZtra3jy9uJZf66z0IHBUfC8bW9Qdl6jOwSls
k/yR4FEGSlujQ6JB4ozSeGjP/OphSe8s/H+DVQupAGlL9coHAVU+cHOWLSyDuzhM/UZ/2VdYXI1/
d5n3o0gqhzicp7d4sAgW1+ad8P8IXNCsg2wWVJcePNvpHI5yUnca0aEhTn0YhQi7CmJYLIkctLeC
aj/dAFaeJZ1L9HMRf/KHHQp/NGNKRZcP9eqUsIrVC1MXeKBFKYePkbcyaK4o4b+4jwciPboXK4px
al2RzzAGogWPrzA0tVjCC+Tsrcp1Zl4hu8WHzG4diLmNb4g1QtqykDJ5Yr+LboFLerYWS/W6qdYM
Kn4tab8jNKAPJsSgvmR0Ys4vJFu0yoNh7c1bJ/BVfDWtHft6l7UCLnK1dQZsthNYLCyf+Q58voKU
s4yd+cLflGqAILZbsZ9A7S0FlC31aUCDiVuRrdhZGc0BkKxM0ONnhceczW+XqER0DqTLtLcmtUIn
Zy62SUjuaStmqXveldGetljvOeOCUpFpz0DoV+eV4sWQcoGQOvKyafD+bx3CyI6WhzllSaelTXZV
WD3/gf5QLo1PIdwX0Gc8JNX5LAHLSfsFROo8GxzFYNzj4vd5WoY3oSTd29AkUyuHKe98kbhyk6MK
ZxSljt1lupc7EdsO0rPttx3G95RUsLmhrphb3zickwpEXXMlk5/f+TaDOszXxRVBW6ylNZRKi3uE
41WVnhTuCTApWZlZ0FBfJZafIFjL7jr6hem9c87FbuEZduLZHo8xufgXKkMKm4WpMEnJoCEFlV6D
lUczWaxYdqfTmD3jNnEZcrYA344JI5TcZXM3m5Cwbhh0DUYWkEvy/0N9celDOUVh+dwH7gGKRSag
2BB8Re1KDtmPHRfUXwbw5Ocn/gCjTNXTNfXr7TfFRfU7LMOykZqNZpm8mzGh0NCibC5lAq+45Ks7
yMUu2rxlImJAj85MepISWYF9Z7SGBY1l3mWNxrGdKr6Y/NU0vICBCZVdy6Su5MFiuXhNWiGGOQ3X
QVBkYRxGStiQsxPZsKy5pDMGPdfAOKvB0unMXgbJAcBgO5gT4qgrulxiH+v4vzl1QqoMPzMFGDqD
oGca2KKct4Mtrl3WT/xtJ4Q3DN5F006KpspeiV6+p5Wkyaw4eFUDgI31dfiCzpDRZkV1dzzxskCn
Bgo0gZTzNtMPPmIrAzhSyN8Sv+BwwKSCMGkfakP5yjOxPGM9OpK3482dheyfGgKl+8DF51N5BCIJ
31ZzdYGeHcDj124yPCD+9KS7vneFvaBG0PbEHemtZn0Ati5a1RBT7QYk5SGcb6E88vbpD1UZdmEt
we4qStgwIPiDgr8Sy0Y9aVrYjxZGXioslGTul0SzcHLRCOrll9205HhpJ3+6SmmPgraRRbzbcZ5i
FtdlmC4AW9BRBBfEmd3GWtRsGkBQJ/2kQ//rm43D/tgiqW03G+e0UHi5wRHj5JnVMsrdAfiUKyUp
7rJYWDivydSe8eVrSB98ahn8jzL8JjuVcJ714WmLkTsx6konRJkLsd/cFIaqvjYYO/eMoNn8ivSK
aYEF0A+wu3KnpStRJc0plztAQL3hB2I9/VdVhi3Xf7Byud7eNQfV5/StKbOLOQy/kNoYGf/ZxpWL
7+LSIoIUu5cuQ0eSI1Dtc80zqGNgtbLGzfAwjx2rV5guFDDKKEaUkw55WCefrhOIl3D2aAQhhPJF
zL1Kymy+lXJDAWFJjI4RYLOn1WNIJC2v8ouVc1nblwQHdIYJePvY/W0CUqOc6ZJZSPo9NhoIOqXP
ffS+yZ00vrcqGIWJekprFu6FT8RG6+tC0+GrhvQGGRq1TuKzSJqT2QzX8J7GvJ5OI92fsyDpP8SL
P6VuVyrBNzmKT24W/Ob4r+i7v/D9ZUXTBlOIkj7u3HelckilFF8WSPEqZZ7RX1dSmHo/jY6wA2nz
X/s3TrCo3UJztpe2blnLSoHmi55zbpA471AGHcKzczauQ8as4Z6Gclbv+WGkRX1+5SBDzfcaoh74
j9gVug+TSCW/M5tx96dSzZQwuLvRUvotAv+02z7nJ/p6eVulxKU1ESmK/Y8YtvWSkprQxTQjsMEE
H/7zPocnTBzQ19mFr3vM+Z6NOs0F5CeBS3iIdH6LJOEjB69x9bswYQPhVSc8abJjBMx3yrz/WRrX
10dDYElGSJKhtNbUEwCo8R+uSoW31ZomdlNAV4AlRY0WxETgXDEoSmOd2zK4n1CyX7UIdHNTAOzu
4kvHmLwJGVL1C+K1BAmgpuO9CpXDu48I7HIP9c0PVAGDKVtkOlIITdVSBYoszT4z2XrUmstP3Jom
b55pKw5bcZk40Ar/wB8uvP7sZDSNJ0D4nwLTYu0PWu7gjs7aqUQnv/3TZhU9cuS5MiwZcRiNC8Go
UMKm8hr+Z7jHAGqp9RwkuUyFSXMbEszx/Gk0H+gioB+5wmjrC5oZ9OaK30dNLoPd6NzVnvrGID/h
/DXCUz8zOTWadbazUBoGVQASib1T4Mxt4ZBzb/4+L47Ixhy//L34R1syzkHRAlqVrNxYBs2kd7XS
aZxrw6iLIfWy2MZCmEU8XJRB2bdtmc6RAPobDKa4mHHiPDcM4PRXTHIcbaM2F3xXP5ErgkmpzBw5
xYZm/rBgRwQV2idtnQqmP5DpiyUP1Or56jVh5CLg+v6VxoGAipZXmq4gkA4hGQDRa9B2gnD3Qayc
gHZAhRG6bGjKTZCmatZ1gJPJLLPTtVe2ISkelQqVfK08BurWhxmaUVKLSj9Js1VifE+j5C2fhY0l
UyKFvhScxcu1vfuh5eqDFPmuq+wRpgb6MAa4qaJ5cEUwRX+4wlGg29w2SloXYvcp1nE22Ps0DUdN
nkFdJrT+Ftj/+OAjV/kn510qEmvrMzrMMIwYroKYihn5AQ0QjUa7PQoyGCdah46g01mwRZZ1Mrsr
7WNE4g2Y3mLMEuL50gEmWjZhXQr5CbmDvQhAn4cF88QoA7XgHf82Xme2CoDuvcnLq6GaALAPLa9t
6VUUz2Ej4Q0UKTar/6em+xH/ajw0RnjBI6zgRYlJV+fGDtQdDBgp66xrX+YRtgkPMRUR16wn+cdK
IuEns+J/23c4BHNcRe4yUAVi4OMX4KPZYr++nliyBav1PvWd+Rvv8WMzy/nW3krKc26HiDXzvDH/
L9bbiWTNxCwxDfPvuC1P+KL413c9bsqVmLanYKL5EFaW5txk0ZNOYLjhcQeTcIzuAgMdBVYrc95q
BaUuKHUFtyiReaBJ38VL6Cx1ksKx8kVkImfEsrYU4xbs5oAnjZ/95F/OrFRy0MxdWCjt+e/kF/Fj
pjxxuhqyZobqDY2l1EDI6OAlL+jUBdS0OODhSnBaHeDb+WQRibHqDCFFxCEblSqnBLTLofs5q8Cf
jQE2iE6+3PHsxax2qjoxv5glMD0GsjQ2CKjO/LdA6LveBWdlkAFGu5tQAUAOWF4JI/nYM9P7B5nh
8LBKW8Y0nuTDTQbUt6z7ClUQmbPaLseQFezJM8aHuhZhgypGK4QH0jMFhPgcU4WbQSKN8DUGbA/C
+DlPa4DTUB5BQAm19LxPV6qPM5MfgmCIDlj0sA3zcr1TKiDyD4I1fVUczIyK70wEubf6ZeGqXl9e
tcRdsTGKthjJKomBWcCrI0vLu3aeKhMJPNkKIoLEOvEBdzltddYyeITOBpwwfzOsSTu5VzYPgyq+
s7STZU3MxWuUxK/exFRsVrppd1u5riTS2v2RaAZ6DMUNUVVkQ4RxwIZtJ7S9Cufkm/7cSmCPv2Nr
+Of04kAvqGNeQJFSj7SAY9uVFbhODZCMPtkuB7rcExI9i5lNcpuWnA1VTaplVfwYZNeQntJawjFs
HnnCl5oxxRhHV+jnP4iLRY9R+UUFAccz0gun01fFSFFb9OlKkSRhiS1h7zYLZ886uMQiwrhog7z8
Mj50Yjb9yKIwv0yac/8PJIK6JzbtWzBwiLp3SWUn+P5wcPH2qSYje/pA0AINcxkd4Ii2rpHIkWy3
iug8V70AGIDnHfvTUgmoBaoOf14P3OsUlKKNewgQJdddseoZi/HKCgwL+WDgHo2CLxBeo7YZjvzM
C7a/ViLy1Z5TuFhVV3e/1qJbVEVkjuR+HdfkG1VaFh54QZghRPuGwac1oRNlQkqhFlw8YpfnVR2s
BiQRO7qjIf7/ksGfE24cuPXXgdyIucP4KlpV5i5HWF+J97RBEigOcwWJcCw3HIQG7vPsNpcT1Uit
HhGh1pXbG7hrZ5RajkWAmVB/cViM99xvY060AlZ62WQskOlXHi40w4H0PM+hFBp7b9o8RvuCJndL
OXR55H3ksZxlMkoeNodwLSjeGWRWmMApyhkCILHtGttZ7LbjtIwgEYJY1vVuCxt4tdm84iafqudi
Uqn9Yc+t11zmfW/vG/ej8j/FS4TGXE7B6SgUYkAh4Clj9nMjRqrwLs5Dt6rF9TFN517+R0qHDIja
eRj8UOK6aw44DDrL6hBuM7rVwikjZddO23TVW0DiUKLZvd25JJy2PDg/Wahn/dmgoRWjH6uA+a6p
uOoF82s1aYvpshXFHMvds5RGvy4vgJM8S21x2SfSPgMLLlnbqnQ8D5soOc7k0ns68KNFFeybCiUU
l/LYDU3rvGr+t+xRAoUxxMCxQqIA+jh/aNc1AG3qa0WqazFPBLmR7ngeHwpWv7K/aLPl2bm2gqhd
m7bv3oPh93Z3q8qWQMQ0klxf7DsWusRAxLTK6hTRhA19FRwqeMg1OWDXDIcF4BEkmlfXaN1eU07G
qq+x+kAb4YLFoX0RtDxapab+R8r2cpjX1VEgnE0Jo7aVan8L+WVr60UALqFXA8Q1QFwGckYaxGkH
Nv+Wn+pBoijfJhPeH7PVYZz52mPm8iVcPJil/w8R1tuHWWs0IdFC2g+VbDIH35vT3MX6iO+KmdVr
SpIBuCr78wAIrTPsuADEiz0HMdRKWdaKJd/xO7djB1PFRb0cTJ1srpS2XxUfQBc3brkw4QodFHcW
Mg9yBquOkmSlPTb5fnZRwMqZN55EOMmUHkGZkOTA4Wvb3UTalRmOeT+f5uPjLgaXH4kxGlbuTCrg
ECf+fg9wqQUn6ioZQTZAVWSb1oBhRPXi9MKIVmTcXmldjv85EXq0bJ/4eHjMA5FUBNNWeMHzmxVm
xi7npE5nCqGBBPhEyJC6mXNOF62mva1aYAH2EX4Ra1pF7d6LictKo1oPA2pEOYS0UxKGDyqQuQg9
+EJ0E9eeRqJOplR4YYKMmPULbuAESMMfceksYE8bGciAqJ87tlm0b8VUECKnslpApx5D9kE0qbmQ
+ThVGjqAzZkLO8dxtvXorgytego1zPpQkKcfj71Ao62QOh6FDdZR1i85t3jgWkfa2+OL7IZfR5Xi
Sa1g/K34nfe4iE0OVEOurvJmAbaemEx/VLoEprZ6q2fnGUKU7pRQEKqGABQTi8B8xmBLoBfd3wPK
KSFTESHDwxq9NTpNtHK5o4WkGfK6r9DnW3mSn5HnZKI/uLE9+worUccz9bVfgo/Ukn/jacKYyebJ
JjP3NhuzvfPqnaV2yE8GiZqxvycy+qtqtkubHYufako72XD83qXDhRBp9518pcJ6At0rrxjmSXEL
xGA6RBVtt4nNgF8kLLDeNNVy0t+rSsEw73tTV8jWVHAeXSx+LLnFZQb/5xWsZWvjHqzAtgb392h2
uNPaiRKC2FPOD5Bp9KBSKejr7D2BjIJ8/joUlqTAMrLrChLNRNwAkFQptnNFZduNsIEhJ2Xckc4B
c6fGIQFsi59vhu36w8oGuDVYWrBIwOSmXiVJNJGfLDEcyZTxkjnTNJtIX2Sehwa8jdb5Tk22Njcv
5r39dyZvMKMzc1taCAlnvnrAxTT1I9KFooYQo6Q0BXIXceyZVl9PZLcl8Dvq2LD6j9bn7hZi4yUE
MCRz3+33/CK+WEFHpvm0OG3AzG2Pv7FaEORnnx+p0q09d1Ha6DBIlQ1Uij9xo9dRZz2yt8fFFRwR
CpMZU9WekmKjbzDRasBi9/XBR4qyGVZ1zVFQye/v7vR5Wu/L49YBAbTsE/VyLUPS7soQcQ1Kyngo
UtZkyBi62g238RNnGsWHeXASnz7rLAHKsGAmbqet929w7+BiV0iphCkZ0Zmo4d+QIeKw3Ss8VuiI
q7taqNNdv9dBqGH7yh8PQEpaEhsx7rpgdyoejLbmcnN0vkOEYIbxxvgYxGedRL4LSgNiPUPazZXl
msvkFrv2xkr4cAUFew0lJKGsbNMaGVl6/CtL9e6+wGz8DWX3uaTZoi7VHAUFCs3rnE5jA3U1Sc01
DOhXkoOcTk7Qnxg52dO/r6GKHF7KXAFsaZvytZmPE9SYBCw/3BWIg1xnenAbVVhoVYYwPBDZqcLO
j463XR0ijMCLjmE0L7Yl9dcFReh/aABHjamUgXp1WQkokUkHVVDZ2lnhZVHgy4TI58vI+W49dH4E
rO93nJr412QFO/dZXLuMc/fwe7j1DJ6JfYehBZoODN5TD9PJj1uvATIu5bOdHoNd1zezPCmv6VgS
73VSLyWzV54smnq1ouTS/qHaOcSaLHqo39xVJM5WOeo44vf0iLjJodLlVae3UJL1TWxb5/UVmiVN
hqQJ78PKUR87GiCpNJaarI6Oid1E3hlSVEioUPRkAjG7fOMyCw46MvtSiUNSDGWDENUGDsrWahux
RQpJtcgpKkTSYCOjZPu1Ll9/gRlT5uqzrTQUoKf4PCxgoMkJ9FFZhffTd3QjOk0B9bWDLV15fR/C
DZ0rFcBfx+QMj30w2Uzh8GeWJZbDBxmblkZtftMB+YM5VlV6nOvnNIZamXbwoNArKSWv2Go9TGst
tLHt5Hs7CwV5YxKbWHsDF3gLYFcLS8HU7BgG7ccLEKmFmlySG1pr/DjIsLVVyF2BUSi0zYtVhYRT
tdOeHVJDfXZcSWwYLxNVTTxf8j91VhLSvqI/sM0kKJoOxfrxqLjoSmj2488n7pFqO3zJau02t7ql
obSyvgf/w8kaGLfF6uZlsj8I4tQ9Fd8DuqRikUDBQR80FZRfpwIznu5nJ5nLH0Vg5/AfXBS4TXiV
UZGPBgDRJKzVSHdlF0Yv1s18HcuRpIDd5/jT/L/XxRXGf55xMDtsXqnvRFJ7S15LBwuKqof6lvrb
uAQvDrqpvC1acTI50QZJiP3k1BQl7g3hwYdpLrBiSixASwJBMIIl8HR4mSTlBZABBmULkZWMgVb3
ZBblOnF/srGLO0kFE58AHlwz7cKVhYH7QZKPXXUkEcbsIBoaamd3ob9cy9HGguqsWkjU8goR5dJL
NumG+kcdJOgtuM4UqcjP4bFqYHSfcqt4kSEj2JcmINUGmFFaVT9PzgkASfladFxbUGeuEOfNn/SX
Cf3Wf9DnsTT//+pDZMGiXHeD9mIFs8CN69i1f08dVl9Y+QpXeKk/mepM0BxHjSDbLlTSlGIuCb/X
n4OBvFmV9jOX5KwiBY6u4H6N3lWJS1xukUvAxoeIBV5iNNjQMpoNcwPXLTj/CabESJUz8R9C5Ja+
orU+y9vNb5apoFclNe3m9EpucPaMDZ8jW8sEm2fZ4o/LBjubPFXjq89G9r8rqpa5DDONfW1fETc2
9nAc+3cVzayqh4NLdBbmWJK9cZ1+dk+ZGXkfPIrVz4gYJiNRuuzfQJrHS197GSA6ELyYkhOiYm7v
sLB0yydBazhaZy+732cPEIoS3QBW/Fi1+fVy2+VwqPF+EVp3hf35/tN1dFp09XjJkjCfkCybIch5
a9nm70x7DfYmsaQYIicUX8tiogOHaYxSiHx7XyjYub2u1dM/wLm/qBl04nOYt68BuyBelte1x7Yy
HxajeYqQONUjMcjBnoFVgYPl1OUnc5YBh9EzLCuYrMKWHCT/95zRR2LqtQchspWvFWKIwhqAmHcm
JVa7ub3I4s4V6Nh3ZPsQGTVW0JANIPnEyRn9JhoqBx8YMD1LpJpyaQHWDs3jcnxhfzh/VYzT3RvR
t2qX/65RFz4glzDCHdrPJgpQuxmzwGJqe8Pceh+1Cp8GHw2MClr0DicHWMSsZktvBorU802qdD6p
o42u8SKOP8T8SRZWw8qT2RDzJZkLso6CnVwE+piLQ6kMzwvyJOlEqIx1njaK29PP1lHeE/71LFg4
yCV5UPZLWQ5DKBwhNNpU3/KyTPEIQ+NItA8kjukWYwbph9QKyZue6ESNE6IZq7VyYRgW75gLPOFL
w8HcTnEExSZsSpCFNhAyGUy943TF3pM4UmMQ/eEBelPpGwQy0tX+GYstyXEVLLs0MASyw7wuaF4J
3hppE21VNN9zNhHjp8/rtj1v3QFizJexwvVhYDpuuSMXkdafnJS3n/8s2JVsqXeWCnYDn1edaKks
RxSNjFrNRNxbwQIRs4DZEicmPYTFb32FAbZcS/IzBFZn//8rmD8bL7EYuFz58qOiKT0/tgv44kCU
beIY/wJcV1OA7wvVHMOtTyVSbsrvj8W2pqbDZJpsxLg22jBDmDeAYxVHmBJy4BJnoO3cSBMTUu1v
0RZyhk03lfXPeubGcloEAHZDDK0/jPdR7sq2nTVWugSHIeVCxcyulTGxWYlgdS5oQBAYE9k2cPuA
4N3/XrtL+oljmpVAYtHy1qmBmC2Ab9z2suEoSNdbNREjauiGZAWCpm8Qjwhtem1bFYeVh+euDgBT
wf9+kTiMz0tKZK5mhZnFz9GGRe8wl9a4eZNu0uIQNpxDCFgKRllNcSjBksTDOiNNCyoFsxckw0FX
muy3iSf1EQqbgKWQC3CeSe6ApBShrShXveQSCZCCpffj+1GuvUQp3choO3HJTJJb8g1+9XxCvbhy
4h6we5nh5EOZdCsoOup7I/7A60jb+VOOj9YkHnv+MLWDYOGryZDXAh98hnGBvsj7FSmr7/YSZzri
eVerEprp188Jv5YYkVB1YRJkuv+pcz6f2KbOG22s0De7ptr02FxeUp2NvMD084/ys4JrcFEezFit
lNBS6qsZDTHFkDInQ5ti/KiSDbWr+7EHk/RD/SlTeW6E8Ubfky4v+NrcYWYmy03qWmzilPUyHX9b
pj3WgfDVm9RVFcMvvC5yGy4qZJ4QfbzvuwmhBFx43s1XeJF42Hc1QFATY0rjewvgNj/Yne3oGF3/
+Vju3wFkqhrj7BqYB4hoQdbvzQIy8OOS7MLBYU6laHVkiYhOPNes2gmHCRe5iMGaX8JV3vKMAXiM
wAd8oXwKlvpUv+bKmuvztRzAYG8iDzYXAx8rbMObpzT9O+f5HewjWK/qzQYvnCbcucAEqu+CtC8y
2Y/m4IlFBfESz9qVrg9h29vhQGUsSA1lDUvBSMk/L+ibybPNj/CVferuGFZrD3NWOHTGjyKa4/k2
8LuGMNxwKS/PkUqNVWcTOoeCcgS8GbW4oyHEVaj5PVq7cCEO4Lt5DW0wAksppIMzdwN8prkuVgdV
QNtGrqptLejeKngNiXKS7KKrlxLAbrlADH1VdrNCSrwgm6mK3132yccAlr71wOJ1orQmPxHFT0+i
u8z1LBNcIra1dw9lOsESp73x+JcN+4VFob0VqtSAEuRNw7ixbzw2WjTL1MBVU886U7I64zewNCI2
K/t0GbkRH6JeR2dTHezWDa3XKOuHoKJ+V8LkBMUOUbeSc8j8dbIMnkXXNOtAQYrMLd/5wgpDezZy
Inuobd1GZMj6rhKxRMqZvwu4Fo01Oc8kCttYhdXf6APu410PU8rQ/M89MLwiI4U4LDe3JkFbKc/t
WMBOgwEaNY9t8wUQqmFM5BW/c5RD+geyYFt30dnQ5F57ncVRzgO7fgtyj88Q/tqU+L09aTKY0qlR
vqKSolCVL82nea5UzQAAIMk/pupRQCBwpljevlEjo0qDEU5kVuyQXoHLhw7hGj355kM10aeJJXUV
lp/hN3t3CdNBapSmRJkIpkZGNye3YYyO9d/NFo22sMQUpJs6ABGlCT2ZOyElEizVSGRgVr5ljKIn
/iBnOQpyjWC07DhHdFzcbjzttvwb8LxPI75CX83oHIbuLfFkIKdO2WeFPG3iKFr/iRqNuAQnYKGw
9nHemKTKpLmrcKd3yAnmxNN4aNqASF90H0I/kaOcRtN2wfWDhy1eOTE3dCAEFOt+Vts1QpaJndRI
euzvWThgvOsPKSMvlCK1NQJTf8wjVGbEKgXu/0qVnzo2UjTIyN3V9GcCRQzNnYglFc/Sa64xYO+Y
s4BE/+7BMwR59fEyVISfEN8HhOjRs5JYnjNQu0MiAb6HphooQ8Zuak6yAnOCay4ZcC4QaqSXCNt7
XSpCQWhh8vb3h1PXBLAbCCzvwv5gQMlHW90itmMk5Vjq/PpA9Heo4jOGpo0FkAJSBsKZ+OjlgSzR
aDdcX6kZLGOixnbEum2bTti6g3E7JL4+Ulaz/rLxuMGbv0LFEKhCUwBdogu3ze6AOX8sCdtogHMr
iztluIOtqfWcMwMvOergad9lEbcHHg4wIcgqkERGeE/6e26b/sZ94/9QH4FzzY9MxnyZ0BGHTS24
i3hQX++brcXyrn8bpnfb4tz7UUAq3ljVhA19XXvR7VgfZc1/iVD+LDiox2ndF/72H9jIbNVrLmNf
9ihA5VxtNyW8QmGMbp33Y1W35nvf+4E7icGPOQz82KSHmoAOzgYUJGUQNWQBfGbD3z/ekj2a0u8O
sIqIbKBuBisyeo8SgfuPDQi0HLRjggVc/0m2H4/yXZNdY24oumCyuNBwJ8Vda3MN4iUDF9SEhau5
ikjsR3Qx7vn9YGBy1xxUIr71U8CbLiEqGJx9yVCx/hWNMLUiNoqIK5HtgiK4IjNGWKgG2WrFbUld
wz0Ij3JimKRoWc/yPcPDVdvGJ9PWdLPb9C/rDgb4fZmcZ//3K1f8NSZvFjwdCO1pPEPKAv03RDRx
TnjcFGHcelOz5zsbHc1vaPHtfHyNiIeZD0C3MVuTeP2+cBoOrMsHFqlfLj6vFKJ8dtzPvPlUOput
Xr+n2N8kMbaBQgDpY0mgq21L7es/XXJnlqDXRLLNX05jr/maRRPCh00xeRwap25nO2dgY59KCnnn
NjWqGTWabUv3tHWPHRi310fsgOwvjJ2mvhKRK8aig/15aUHaWlwRmB+WEQj8ngCJJQKGO+3mUnND
Xx5y0Pv9XfFkgtLX1RIMcG1yL3AH+p9pEq0gBdFu5tyuAAe+0whO0MBe3vmmY+KhVDbOCJZ8cOAa
hO859PgdTyj4Vl4TU68WN9SjjebcOo7O6fwwCkQrjfyG3tOnj+eWvkwhCIYSGzJRL0GvsUEhTOvY
Lu62hqz6D+Ux8i6niSYpwhSoxS7DlTu4LftQLiQMWPIDHR3xWmcVBwyoYphi7TW7XfGd9TOyDRVu
kGqMuRl8T4xLU10y8PPpE21HgH9mYzSFfHeaPEN2ntdGcCMteYznJ/O8Z/utyrAyRnJam7nALzTh
CkgUmZqX/6V1M5wh0FJm1cGk4J1Pq8yQy8Qmx3KOQ4KvwAxIl/tElxzNqJhsQ3X5Zs5ReqEgFX28
0LPPj7FqR7lFiNkx2lr6TXY5OAihnADfWpFSP2RdBTyBwZoPD6xRKC+aqmwHwXT5KGAuMN/Icu4X
MyZoO8gHVJfNWvCNk6k+z+mmiqBFwZAICeREyat/ijXpzEpJWwE0xjvnTmba+D/JwsZzDsRQz8mU
XR2CPBiJsq8DXp85nF51bH3dwUjmyBOZkpP9UCPPjae2FyW4NmP02gAk20VVNzAIiQmLeGemFpFi
vOexwXXy5JHjX14SPt63a4cxjPMhCQYqx7I5FnTi1sRIOb7XowuSo+9uzaYvj5j1AZ9vVxgLU1aq
8go0bfVxLPdBvg5by4hIGH3OkZwKNmvgt5JALAgKK8qSD7to78foJyvgVdjgI1RYGPtYjIMlWy0U
65GTR8tp/HSCandhHsWRVk1crApa8yjO+PXkGC+ypaCaGaDaXroA3J0LO3XjYcpZF2U8ApcrnQYl
zzWJ79T/8xYzSnzbQANS/+lFS6NJ4/i0eyxhFO0pVi813V0rBp4gzgUmyAaDsz9/VLUGawVT27dH
EHd8f/IPM+jAAjSoDXnI3axwzUsMsuXKFXNkIxuavwZjGU5tp7OL53Crik7woJM+rH4iRCxQt0Ae
jAQDOQ0sx8cEfK0Cfly+js4nQleeTSMEAEPoYHZQd9ufqrBXVriL1+w8a47VKEML0QCp3F+eOikK
ZSnxrmF0zvsjJx0fQxLrTpR+ybVvUKHoSCQa01TSXaWvV8S9+a+o2cBvQbylYe1Rx99F/bS/FTfW
falBrXnjLnZOq/rJi5QXe1ITJiDBugxRtyFf2vWvTtK8gRg6YINvlSC4B4qUlj8WLOJy5XIAPiUu
uRVOTqnxxqiQCnSP5ic+EuGMF6Xqk5YLD85Lu8GGNSMIiZfyxDIkbOhA8VZNe21O1eQT4sDlfzei
gmfHP9O4G2svOvLkLuUppDJliSqQOOp8iaQTd0IX7aKe/SXv5FvQHAYfsdvdDE34LzWBhpiZs2M+
Iqns7y4E4PJP6HxwbcuxBiboBRaVlVMHhxh4UWAyUvMWyXqXFTjY9HiyOTNjfBvpgkIGEvGJfkcZ
JDAATe5xkxp++DMOKhc8u4Ky6rvCNPrUSFLqraSLPhvF4DVklJu2Uzt5sJ4CD3mCYxPPkzqmmf/n
mPuipGTXn/zuDNNyOykadydeCOwKOdS5xSY+gwCVX9EyXta42wzn8ADp8TluXTr0UUXqshnfLCRC
A6qzeFsuHKfIucpD9SbuMCKS3YbPS5NupZG7TWYWyAlqeP4IJlUKgT1S4NkH6SPaqsIXnV8ydB7d
PPhmZDj1tYphwX/whQGfwVemxRJaxfQ8HwqWPzRH7paoSXm5bJk0/rcT7ciiL7sZ+zms2C/H8iSZ
t5o79j+9WThRozXEZ+rSPs/KRvOYFuxpK7O2fYMO9NfTMhk+flPxdT7rxJf38qVl219Hv412EDvL
z5A7/bTnqnuWjmFJr/9hcSZ0r/UImN3r9AuTS1ncMgqXzPIzzy+idy+uOiPvJrVdh95kfX0i/v3K
kMuiNP+LVXcbQPileufmSG4B+4X67OyMxk/n7R6dZ0kPeTfvvzYNl2plAwGguJR8JXXEBoDgIFfT
4G/Y/43HaskLA2Gx2RN2+8DAgHiNeFn07orxKSpTjVEoaTWALV5qscthVEb3gBMpvgXsvP1l88lv
JfHTT4ge80zNsiRMOzVpHHYDJPKz1CpJL8xYi9GSzUrI0kLhgfiVMCCku6xTzQWtmY5f0RIiXFO+
BcqASuVSp5MxzfiB6eNRy7uik1G/CTUi9EX5G6IF8/jEDTI1B0DVilXwsmxjBwykStglNLWwTUN7
fYx+cRdubDZBjwAq9aw4pbXSrpdJDdah4xZa7y2peXRvvfEXWZMpSLsDs197mihhUqChPOWDAn+6
THDpA9+QhWa18QQAoCuRmXjBOJDGDY0kEgewZg0kaGp9Rt5A/h4TrrqHitWeayTWWAB9TVRorqb5
yyMEO9Z1ydcPGZPdstIWCANu1eiYBytTskThX7YOUKKzco6VXoaIvr5qB2Njdfp7mINDgjGlik35
sZZpvtBQwJuFihJa0SPgEEhXO6F0GjS+ABWJYrfwyTBjdnqQyJ6GMNJNqTQDjxJYd1la4PyYZ439
g4p8xdap4NKZ9muD968EZAJiOH1LlVprP1vAmz0QFpCl931E8VEOXiDwGw+x1oTNFXgLvxQZTzzS
p1B0/m82zNk0Xj+HN5bjS6k7Q3hCgEaQciV/m32GaNO6Pk/KzNW2dl4r6NX2HCMLBZtLkmXuCIFi
Y+HBm1cJQX+Fbji2tLyguB252Ht1Cda45ppY8cs3HdIbiNrMNcXiUfDqVuWl1rMbdF7WTzer66ef
jC5cgd1zb9rAfGJERHs0Y1fVjdMAlTu3aHQ7hFaFsdDjD0yzmCTmTeFy0gqIUU3FrMQuyOb+ai1h
DkgZUbfOtlJTCUqvAqVNeXZyJeP7rjutefOob4LpkCYo8mysQvDu35v3/epfuh7JF0qnJhp5PiXm
BwiV5FNZ1/ILa9wNB59VyDokmJrAHEtqvpvReJxIqF7/JMetjWMu9H67UHc6sKxit551RGJ1KCop
S+7AvS+9g1Djzj7O36ObIlUt3ZU5VrODtp2islGuN0t1naBUle5q2siE3sPioLyeQy8Y2Gn5Y3F3
YgJp4ogYdo2K/ta8VnvHnM95yMal/7fN4UzdPIMJMTb1he11vrBzw403ozswwksT15hUB1x/9H+I
k9UUmGRc78IiShK9j5kQPuLVUwmXeViyIGYv5Lg9EM8Txm+uZm+k2QCNpwnzi3QmU8+lH0iY9rC8
35h29xkzKx8DkmQuR2sn+KA9xUcYYmH4Grhtu3e26D3fCyelQSPShcvDm8RvAt8C4+xVFVLS50zG
NEbjBABor+oSWrlqqqHnz9MzRGf3Uu65mkl2xond1OAy20cz81N1Phq+EE6O5im27k+rMneqogGD
jIu3wFY76J91Ma4tgS3SYlXHukXm9hgS+SuOo76PbCcrvrbju98eX4NeKh2OsjQ8BJMy0UnZT1YC
P3HCAA1iZFA+kWRikQrLI9y50VPJVoQgskq3FM2v9FCkMOutpDABXylUfT29xw8Rl/QWOWg04Jbx
FvR8NjqABqW5p/bsAXXKuCT8RHI1kDNLymiwme+8lsQNEOI/M2UWmqVNDNxu6Husub3OB4S18nwQ
DtnDvuJW7RL1CYpNav854PGGF9U7ZXTMa772QIT67c6o74JGX21jf0Ppd6oM+8Q+afRAtv2+DQYn
Gj5xTt+dinYjinr1t89VCNNSO9etWLGSQtO71VcB4vnAAvAyo5+VB5alvbnQmiGi1jRQfvghqBew
8nG6b+nxXwPYKz2sma5yHHBJaLvvTb2iRoRTdBoZbTR+OBCiX/ha6/UrrPaxY/E8PdtPQV6kSqXC
y37xDtRBLyReWEBL6Az6NgoFBXlSQ9otnyWvc1pAQOc7t/rZD+bixcfdT5YTf1qdKvsuHI822utM
gPfBlI1G7hZq/tlX24eYv49bi8/7bg6hJpdJ+woCQQqc/kyM+JeVRbX9z3iKZodlFdbYzi9TEQAI
gDdZt3ieBPwwagSBpJmvlo871h4k52Q1VVZ5olK352TJH2jsuOOBa98KVkNu+xEVRiOcHj5pZdYF
hRvm8RBUR7F9qTEqkQcc7wCH+mBWqaEr4p3/xVWFpAf4AcuyJM7iKVdHk4dnAwqQxt/GNsc5VigP
bsZbHGeGb3E1vIrlEZ1jDsTnio1dIGCp/EeOae5KzPZKGRPrKQ9bg8Cx0nc1oAO+VDX6ewJrYJm6
ND6Lyl2md2G9HpYuUJVemefN29pwZFaCa2Kkb0lKl8lfTMDkXK+jFYmE7C16bgzhc1Y7Q96RbzYa
taOAB2jCWfJfqiM4DE/GdEVSr3arAx0ac5ObNxvfzNJ4cluSaslUM+DO2OjUywkJPURd6Zt4ShCq
1bx1BCDqlK46zDSvLnaESDfObpBce3JW4eVUZDyEAqZzlzZO5y2fYW+cnyEnQqGabaw+c+DbAYcp
TEs48YZw9V7O6eMhY1szWpxWHNPTceTJXqaWzLavXFKiRbHFeXjzkodf0LFRQCrkAgcEq7zrWGyS
YUr3qqAIGEUVcV8sgha47mL/AT0YQP47462CtZSYkD0VFobl831cxs0WAiCwfLQM7L4F69DuHi4q
Y+3IRqkl7BUzorzccdwmp7YU8dSVbfkaQSyARFz+uI9Z80asrQBH2T4OYZj+29A1Bh+z9Zhvjh/H
wgUFkAdzun1mvhsKF1fVnkSm3uVRNo3juSRTNZ8kVVeTYvcpZ4pbQYade79r89aqj69QSdla+tjp
TU5HELAF17/+Fh4666hKF7d3KMx0VcgHicO+A4FYKOF7Y4uwva2dHmESh0HK+zhurJ+QSM/PLEbe
RkzdxsuZcj0uIYVzCwDFGvHwCSMvCpRUu2IO1+HcO+79KYHXwyX4MHCVVwFoMKd739wqOkOxBXYy
58dWiZBa0NuMEv4NrE9+FDe756d29AdsIwiXnVwihyxy+4SqwxFq09gB5gKNqtK2uL0Nc8tCZbgP
7HfZcjaL1IyXl0JGrzD0CY5NEd94xAzdElWzO1yb4ghfpSSKAmpLITx4HKg0Aoxul7UGDvFapEP6
7Nu6yCt4kDUkLdrwjouNT8PKM7c0jhoQBU9iVNoUoyoZo1qfJxoJID3zBXDTY6MvI6ypkVGk3hKB
iZNlazV0PT5fHIoejPcaj3iydEF0QFbbuMC1gX0peb2/IzIP+Fj/BcyY1903T/liYqFWh3T7qHAy
KR2K0KDJA0wHoJTZczVfwKQ1oJUKxjIjVlJMGepFrkcb7f9AzY9J89PpZ3CM/MICDdgAhHfoEV0d
EK89/duJgFDEtZrbosR3jKQXoOQC8CzPVdlM+wSBcYstCf4k6U3MM70bHuvw0r64WWCUxGQTQLyJ
HoDAP+31y8ZiVY7a8bkEbOCXMh6R11NECxgOmkAg3TG87ydjXKgy8FjK+DCajwAy1Cq1nTN9eVbP
X75hkGZx3chMa2p6GOAltrims06br8X+pdJSnGlXqhpX3EHav0twEVk0YIdI3EMRNlmSS+IzLMtI
K+M9Q3rboFZnVF66R5nSLgR7tlJQ7zwl2HDoqGDP2dv2szKnRmPfeJvcv+A1ngxm082zuENeo23T
swPSyASsAm6jm+GTMj+vTjmf8wcWisU4yEG1H1QE5nILQ2ApmfFlwAgAhtDlXuYlxMZklcC1dzkj
9sqsRYGI+lcWFGVbeCR5A2glb6CKdt+SOzPSX3xFPUySf6sgF89655/3O7DGJKce1fBuwNuEH8Kl
HZ1mvvQkssOP5a+ITK64bZAfpbgzfzO+3jtF0gMr3AX7k6U0/f/3bcr0M+gMY2igv6uWEfn3We/9
VvOwOnKIqt3fNtw+fEWnhnzlm055j6XVr4mgXjOpgopaiiqm1D1oSQwUaVsGeyOtHybfO/NjurS7
V0UcpyKctxtDLKxo8gSlf8AN17elGNCohp/eWSVbA534OKcgncGtJ1nBhZsfBYIcCvLP+K0D4M0D
qFiOMU5iDwpq3rrBOtvp6oglivbV+j+oVDQ+XL42sTyfaTetOfxD2CtO0NP2eavOXIKSFtlFQEaJ
FtN3cEY1LTnb8NzVnxVpDPoCd6cZvPlvCZ5WW+K+M3Ww55AQZ2eH0WJXqIizkKiEv5R5yqN4F7u1
U3XOw2sT4KiAa7VWJTkSm/5QraZXNXZ4tp6Uv4EcFHYCeZyqvg4qopakC14VZ1fP7bYUr80ehAT2
ApXEFjL2NscMIXjhYAdQ+jcPYAZ0f2hsnZrhCTMkYXkKdMWYyW/M9LYZcRW4KRWG11Yse6GBZc9W
+ijJiGlReBp3LsjK5MSN4b2plV8InDxzRmN59N7LqwB6YvOZoVO0tsMHpFRnWMZ97/dN6vOcbBnq
Pg4opLEc4cojdZLwURoC4PLTTDXKnRVzL9MpMmcmDdvGwj907MHYFyOvZqu8vt4vhzMb3+thFR5H
wEzdTMrNE7UPpVsSsxlAsyUQJKxlZCNTr3Mg/DbTCLc8dCbjI7SJ1ifIx1PICXZT2hKiFVZ1KkEV
8K7/pFY5NwfJg/bOG5JtCyy/+uYxvW9WkgcNCJo9Lw0j5lU3//7U0LO+1n+1nMaDC2kRGwrZPI5O
73SxoDAD08pkvbx6qHjzC1INxZi8dw4zyX34D9lB/9eFHYw1GlhlAUCmbmII7isY4aVTzE8+bjhK
sUPqK441Bpxqg5blpnU/wMWVikxGPt31bDkjVjEVi+QEQvuRuRbsYWt2zIOn1WCNm+VZoEk85+gy
f/BC3Qwb22Ss/1psQfZy67EibZ3hX3BTbA5XwoOn7a8ycsQIzdLPSz5XMG7h1g04LzoOWqw9FiZ6
lwMhmlcafcRvPFyUZ3m279tBHjSQoNNHhrTuAjOFdFrOFgB48xE8O9eYxXAWgVIFBb9id3E8Z+/o
N8EhyTf/RsKY7Ojnfc2D2vFylU2Zyy4Ywg64AarRFOZ3ecao50QgvYmIjqAKWo9uoLTtgB0bD9kX
8DCtwdbRTjGnflYRQVx4gTNstI7iU7EU1tSZaNeOsej8BGGEcJrpIZDL3TLJMJ6dOFF0WwJ0W//D
zX4sTYKfE29prmvUrWYkx5hktUO6HnIODm8doS4waBnbl1lOka+smtkEHgtFH5Pba3Oj3xhfSUJl
KjjSOxZvJRQU7N42zuAMG+J3cqsa/j66ZXTMNeBTN+/JifGUkGP+VWhL3ZaNElyxBGybBEOSgfLy
kIUl5PXG6ukWw3rkvxs/TXmaptaEb+4cjLGz4GdrnWCewLt/7rbgvNOLQNHhCAL/ztcVh/blUv7F
9lf7IepxpzGhU31rz2KD0ADR7/2F1trpQ9fHVi3YexgEwumuLEAE5u3f6DyA2c4rPnkqyVj17BVA
clqpEBhsVe201QmOgZ0EJTkj7rLejmexaOvAojan+a4R2hEAuFKU3GNraweV/V4KZadakSEQGNme
59ALhGFeD9LemQ+QtrLpdxjj8MZoScK6+LwtGnrJfqROnZTSlp/UpzRTn28vyz1DSTgcRnUhl12k
OJCIVJdUXlYU0/AnsskG0LbVQeFINv+V8iwxRqR2TslFup9fQB8qb970hH4LnA0l/xMKKgpCy0E9
vak8ABC2cAeWjV9GUs60YB7sjbucMDAW6wsrqb+6/6VR3jetdB1fR2yaWZJkivJCwNsk8OONfEdT
I2MpwE1zb6PQaB3bPy6P1QHRGbm7ME+GazG4pvov/9yaLxeaLa5uBtGqbxLte+UnjhGSDG4VGaCY
G7+ivm5GXlznIbY1x9li5u5graVVfsq//sy8F7dhKE3v6ZqWBixJylBKmMXJwU/nUcdTGoPqZwx3
jGUH2WJGhbI+fUDEE8sF65dhHhLzZZdWnfuiJ9itL1m7p97DJYbjipMMdese2WzViryz+Eqo57+O
VLg2V4FxImWO9dbebQNrQ4+D62lmO19ppKs5R70dgT8qnd2cTawQVdO69QnrJW7fU4h1891Q8RwL
iFEXijxhurzT8jb25zqKkh56i2T9EdrrrD3+b1TD7H17lH5u2tTXko5dypnUQOyjjj9+uhJrdCrs
wCfikpIAJlxDnG1O4I/8kBACCuUOG1V9Asz6BtEYeaIHG3HfDNw+yGFh5N2DF9j40Rti+aoH8ZDT
bFfhS+M1UiDGE3qQVX/SZlE/Z/MCiS0ZbNmQkxz4QNWs4OJoW5nXi7Z9MoM1YXfLZy+GtNTgc8Sh
3cS9iTdYUEWyC2P8OjqYCinheKltpVl17pBW6xQANBmxeU1TfuMOTBfi54U+tShlv2+ZQz0tINif
6DHT8Et+3w3zM8fEDSbqy4xQc32DpLdbIMQq2sFRAElolAzID5DAkKshMSZ7Xg3EUaGbfXiIBLz0
zOh97DMeKBPYAP3Jza5vo3m2g7Phe2bsC2NO0jZnDa/VQr7wLoS31z03oivDdssfa9U3U0J4uHam
K1ZmWwPhD38auUVum/F5FEDDz41m6kuEUuPyd7Kj2tEtXPyGQ9JfRI2oxzZKWoHQwBs1MkT8sUNw
ZgmpQvVwq6JPk/MYVNc5p80d/w1OZXzJKtlnyctlEUjnZvBkfxMHJ5ePrQzAFVfWrYCetIleiudC
BRJbMm4+e44uP2C8bVJxVeuTdS8Vcg+SxI2ZKKug0nsONkMVNr6qXQIkEXGRYATJwEyJAgD+zI+/
2kuPrvPbcJTxWLeTC/TuxmDwrExv8AQehDV/nKZ+0VY8rO/WfeAZ1AA/Jq39OngAjb/ywTx2/4BF
72qBw9oOD8T/Z5F2qqaYhL39d21fkHihtRQCjV4i7rQNK76U+CA+3qDAifoCpWuLd1hbbic7qaml
Vbxt6HOyRbxAn7GFrAXl9iUQuZfJBoMsml3N+mloZKcOrAzOGserVbv95nbWhf+DZxQdEaLxhceq
9tw/Mu8TLMW201xAH7bewce4pc7qTHdGjMVDP67letcxpgdKoUxgFO+pprK27ggA/MaqH7RTwGhu
/zzDx0lYRfRXpmqKVe07FaG8GaTBGMyWYxaF255yzsnCP8q1wsUVOHZcacNUBBE62VhlOAWQbhMO
guMbl4l72sfXiMrhcw0qlH42I/vMw8em5lyhuz3hraejUSt4bnJTXDOh/fQ68Yya+awKlkAm174Q
l8nizY+0NBdjI3bSwxYOkiR0mNTkfojOwEbGEeI0ABFaWUZsx2GPCaC/iWcjiTme/HWoFmDkFTmK
SKk6uIw3hTZAPu0+SEI4qTEfUn7uSrVO269keJutnc4pnZwUsLblebVyZJzE21KAySS7NHAeCMzU
dB7hZDVfwObV2uJzei9zqtLMrmRApPaPnieGeqqfrKEfPOVdEArZTq6bOEcRScPm4w+P4qALci53
YPkfOC/RwMfTA0tL8h6EsCcFI+A5RgXFMZ1dSkN8a5AW+IB9Bxe6LBs4PQKbm88Nf+fAAGickUbw
5ypAcp+upFVW1zdj83nfhCqbTBvLU8bjY8O+Lw4am+40ipMilK4f6l7NiWWFZPJdo+SRrJvo3gAa
80mW1+5nsQmYqI6+tA1+cJ5ulWOXehgg6mb0t7IlNqDHW8qi8+DcXklpeAxa+CjH2tMXZ82GtGyy
kldQIINluH96Go0Lvxt7a/bhQGAYdrTL1Xg2gb3/B+S+DssJ0I6TN8c7/nI+XJlR/Wl6LYPc+TNO
Cy30FiE4X85HGxEq1hMKjJ8C5B5tvwjQ0iyqNSR5eKa+okiaHPRqkxHIJ556c5RFZPPfiMOIwjqz
AY9uu7fQcr/yBmPNCvqgHUKBAg+XHF76IkmYm9lMBpY+Lm58O6+edS5tp3KBoIHyoX4OXelfYfvB
0yTDRgt2GOJLyISbq5YHZU49jgkGqteZxg4Q0++s2+5oog5oviaI9O72XNSzH4Im185nBkeuJa2O
ScHpCnuHCfVaj4yehZvDMnmE0GkiByXkMjHx1Fj25rR2cPFSbe994mpAOYMcLfIRCMiEWaGv1x7U
h8pareuH1GYDRYV75stJ/G/qcLtE/fvC5LhpVk8jV+zyITeiScFf383t2Tb1zeU7E2snnIphrHy7
Yill7HPGzQs2nvJLe15GpO3e4kN/60xZtgJdg4+nnyvsQTBQJEZuev+cqsVhCZqXHaoF4y3ONc1C
EqycWHFLMgDwLoEDAUZAYyfFhSORL74M5nlAWxAWix0TVCz2GuwiUcfUkPgMb1DnS+UWNFq4iblz
Yjo+836ba5TrwAHFVwGkzGRnNKgUarYK9Gh7RzBKAhAR0IVZqENQHS8jeTdi5AA+PHOGz3ywLSZi
pWPzNHuV3g9F4YsdYKyuTQ8ZXdL4ahhZ3wID7EsLtMHhAWdqPg0Q7ZYxgZJmQefJEaYha4XPIy2/
x23tP4ZjOE2hE/tedOC1CibxAd1YuHMkDsJaBnx1tqfwx2pr/0U5T43FcQ4UkcCl1X/AEza/bedh
JHizDL3Pq0m3uhO/AodMEiNaupv5+Pv//0OyOnzKBk3FgY/fUNpRk3LUCMY5tXShNLD9mHXn5mtn
5QJwkJZHPnV3De8soxYvZTs1CoI2YP0zUX+ePC9Mm141a5KDgTMCGLBxeqJFuxxMFwAWI/wwuK0Y
H0DWLPWTfjSaFSyDEJK8ZuxEhwOkTIT9HOXNVZheRQviFEAo9KKdt3KHObi3a7dL3R+7dVp+QhT6
OkjASV3Q3dKTB0GCdcImFo500MpnGD/4Ko11/tQXo6jj3ajAV4mTMsbZf/ZthAW6LpQ9W0aPeC+k
ofLshqt7ksZEwKyGsjt17r0SuftW9waDMUYRxh8dVEEr0KpZnYlBl8JpcdISHOYJWsGvPj+DHKWY
04G+BUQdVNQS87RtVWPfeOs7CPFIak0fvTxhrzPy61cxZeM6VzR/dGv+iAm+BeHxlMvzdU9ySkQp
9NN1zU+9t2X/NZcbfgVhRK/A/3mxCLElZkyNUjRtlMSNdpoNrZqD7630PH2zRPQ39aXWWXGg7bTc
JFDlGxVyp77VrCJIR1vzspdQeQ8x2yFHShwEkIwrBMZisRJ4aL+NBbdbz0eCLrPWIRe866APUHgp
FxQ+xp7HR57DsVyRpQgiDNcqoRkDslhGfz0UEGNoVIbDtOLTejp1rYdS7DRH8MawTpEPjCIJLoQ+
iAr2BAF03wrLPIHzdwt9k91RfodobvTCF2YgxO58IVoMYEqpf7KIUtzR3NNXwxNpHBRVkFf0s0Sb
bplIvihiDr9xI1wFze6+cmvZsTELgnZnP0CgD6T46EaguzhtyJvN59MJjcuMiw5rFiW4sDQyxx46
qBq2041sWIBRl6+/OB2+NxSgrv/0P3IVf1Jv2gDUKXmNOiITcvm7oRQEe+gtOSPsyiyNnIDYmeOD
+1sQlS6/AZOHv5rhiJsNj+OwVFUuP3bbbycj3bVkKECJrajDO6oRZyCAKqmQEGsXfwDor63651Ln
puzYDzygkjXGAvOtAUppmY3v9arStHwgNghuFe9e0VpgpGu8Cq3Gn277Yy3k9rPXWU3gwrJ8Phyq
MogcnczkUjxQHCCGp4mF5c+4IesGkyPxEGvTtzY082TOBtVaAPyTpUKK7OR2kaFfH1yfta64vVe5
WB9gMJAG/duY5gnxVGzW461gqEdGcmpV5jY+8wb350SVpUk/zaRnWVZRjwKD+xo8lD7k8dYmG3bM
FXrscETnzuYdgOILcTaowcwWtbkDRK9tTlJ8k0cY5dxSeKWkMOQtxpZ5HpTbHVSrTYOQu2wJ9pMm
WfHDFuSzWc040w2DtwjoU5FqhpQuPtCzbu7EZtu+xYqtFtK6tJcqrl0a7oXFRzK6kczBHHpB/Xcb
u7w55iQVrDSAsdBLLhPShSZS7pfPhS1FoaUarK7OXV4kzCuWMv3CKX/0Zk7rNUoESnmiPvWcnm8e
achn68nwmCu1igA2Icj4mT4FZ/lcaZdcPqYp0bgWsCsvDwPGFu+S/8ihL18p69zFwDBo5Ed/Tfek
P4LFt/vur1+wWdKk5jFJkhZXSqdBG3itINch1EindTc6j5ZLyFC0ieIflEr1fauSEpgr5bIS8SFf
TojqnJx1vqO01wlsfuoRs/wVMQLm4dX6chZr6YlVPOKV1CA2XBvKrb/HUF0F+eXuJQWe1lyg2V8W
7H0lB4VF+TuqqSUA7PxylURxjGfGftO3Dn+fbJhWEBnHYahnHBlMLLzLaGHAHa67mLA+zSy9LLwb
n1cIDv2beoOcu+k0sfX6+62C1DxWUMGy3llhEqUkjwotOWxHzNt/UL59uLRjGMikdMFo4E+CCeRn
WNRJVxxzIzRG89+36Ojh/TWTSIxOlWLN5cAJ+ZWdTXg/4GXyXkrcRumjuf5tj5dZv6w+4eEF4Avp
p87LAY6xxC8Q3MSDwxjMe0lzL0wn4L2MHosvArbkCk1K0wa6r52rohBmZg1ksb+VTguFuFN6Dj4a
ZhffZGLRnD3XW+VaMzp6X9SGprone+vG47mHipyhZkRoMQyxvwNfPS0QqhcB+8XAbeRG0uck29nG
diyRxE7WnGYXRMO16uaM/eEVaifbJNW2NYDzyvSeXk9GBJEhA5wQm7DmxWluzOhqR+ZYloazwxkb
P1chsAXoNXdVjBuhiU8Olrx4HIg7eSUw3FrNE116SXmDYW+qP4l39O5fpEt5ANeBqJe6j8JwrFeR
rsslsxsxTj37z3JsT2iztM1aKHCuqI8NuraUbycSkQkZVBBa+VGXcDoAO4lptWy2bzHYe6TeTmbr
pxwy10CNpzMFuZtUxZsv30auAnJEGQ59E2ieSLizMs70yMub1WqgjjWmHFowcX8OaeigVhFgrqOc
H0sSLP24wHpJtwmEjBcgWQDFQqPeI0J1UcX+jfPueKozN7A3HP9uco9u3NnBYCuvORjnMHCG/R01
gWyZJu4GTPVujedie9RluqW750pKFpmtkIze+h2u4p28uJ2rWmrFvzHAXsJyEbVUG+iEXLn548Jo
01AC2QgS5LqzRO4U3N7d0yX1UCpSR4h53tZvG3RzosPB7umIzwbLcCX8r+lbHn3On3l4cLDcotFW
H1gV8OSqFXFkhBh/iqSdtjwWsIaNC0AGtwMje8MbLXqS5H6P6aPlrNWd4e6940VTEyDB9KltXTTU
Q/dL1CBMns0PfZoNLAwNzPVng9LTuL0e5gurZ82kCAwJ7tonrVV5Z6cAsWnGYMyzLbCRkZdnWDc7
4sycw3R5Kpot0sZHb2y2kg7sKyiHE9vtTBI0eLW1oPirVtQ+1zCnDrMefPS53Fr6+m9rKEP+eFX2
94Bl6IpjVMgJZvc0yO5pX/q1JU1qmecKcCtmrR3Cjyvo8IYe6whqZmlzxXX0CFoM3/74JAkGXCPV
t+YEFw6sDUyFZwIEtr1XGUIJ24eWYW0M0SN7apDuXNUUV8CV3XQBHkbP2hCoFFpCt6QkF8Yc01Zy
JdVSr+Nva6CxDdqN0w/0YYAStR+O+qPboZ4u3eXw8EWL9uj9BM/9FAifACp+Q+I/etKR3Rn0epBb
3YZ/ZVQKMUnPeRmt+vxEgZKnjekkmIBtILt1Auo1aLh8CxosDqpF9bNsEJ0HmfKOuMMFwklcHxPM
SqvNiIwZ9HvPKlTvLGT9GV7JnlmRzlDRFYzuILPcJ/83Qz0UvwqZRAdQaRWSriFq1WuJm0+VDcgx
IsCqRF9H0gopEQ7uKcMSjS/V/6cCiR0617Yzo3o8CraXJFHBsc8DHdJMnV2XrxSFcfyZ36S9sMu1
n25aFkf5R2gmYA4gYoC+qYK8LxNd9INrUObVcX5nopCqpqGKENSrdHCJ/ACZiagEsL29TwTSAygh
zCCmdQaPd3ie9bLZesBENUo7xuM/U0jf7YZKgQetoFwj0GMJx5Jpr9HWn6kP1at3evtqSbaX0fN2
U0pcxyhNtV1HM2u9S8kPG3ElKJvAEi+f8xSQ7M4wTb2NLxFQeRb7r9cl1PJoaZR0A6+S8gqfBW1L
G33S1ZuQm9eRXjN6QOOqULOuQVgjpGB3hLafI4APJdJwHbc9xL12JWJUNFY61eRO+gPGvUKRffW3
Eyyf7Lw2Lbez4Z/O3UTcqV1upefYKFONwya9VMLfkSDfkD47OG2kHOyJblHuGMS3c7xB14kYcqvD
z4M0hlyWaxENFgB2FM3Uh5ldCH/KqN58yDQNpiptXec6gMsnOVyhKaufdZcFQo3CW9ib/w5tWIpE
yGdIWBEiN7c5t/imi675zDU90Oi9bdimeAwR3tfV/8N0uYuPo8o+80bg0XCq6sh0h8cEiu9BcKpC
mDw/ZIIuA8yZ1kxtkWpwEPJqlkcaL4yD4u/s2OK1lMoG/yVGN4AUBfdiE3pzohMM0SyIz/mfhItE
/W5uTjbGZYR3VONNzBsozJM0141OjrHuAZaBf7QdD/I/hwFw7aQ6o5ZlQ45wh/Jwx5Kuks2VjThO
wt0eHMVVK5fINAHIflkv9trY5dq4EwmyuJOEFbRIzN2xkQEML5hM9a/Jo/neqe0eEoMkj3rMgQD6
uzIKfwBEhm9LDQZi3kt1f4Sf0jwiuXloPZAog5gdAEOWhGZmclSnRPXbapipyILiOAMd+SCYg4W4
l8Z1qs8ZmNnpFSoVK/GQfLxRmSTDE65gL/yS7yXpImArt04UfpxAxmpWzS7EwrEiQTGwcFBkVHVI
Anzs72ZwnGIqOpD77pTr/2bZIcQRndhfSqXpljnnmS+CnA2q4cNSW44XrTRz1rUxg10aL2nf+zjH
L0ZTiM8082I8Se8BcZTpVc8h+7r2r4lSvAmK4AHZTKTxKTk+DzMBmS9m4kOShF4/odCde1nK7aN8
0QcyWjL0EWlBN65mfFz9to9r11HQSfU1EVbtcivkpX5bJIrjl4F+5upBh9LgP+x4l6DqtQVCHV5p
6stzhXX3yVWhg5C/gnOHj+GPqKD9HMyQaJhr7dvX6I3gR5TkQdM6lkgnjy6xTRoWHl21pwlreGU8
J6tAspBQV/zrax2vYquTtWGb231RkGFbi53+JlS9AUO5h3+X/iXC8OWsdKRu8WSim0ljSHlaETCo
TxFMoFHHi8hqpBtMm958lahhFApX7bL7dYQzjatjBz172jWFWqmOtoXpYbtlSObklXFvK0/96Bje
bINKFkhaM8eVIxl/fjZwXLL7AZE7cTEhQRGP7dRqyZR2CQ95DoGYJe6+fno+Iyji9miA/Iptfeo7
24+RvNNKjPU4uT1tCC+bcE1nEmXcSVavzouai3Md8Qj8pdIUkvyMEhiFZAggdZJ4/DkbggIXInwy
gQkSko+Jc34wYKEqzhdKQT56ux4Vr5FzR5IXubs8OaadHmRFahiC9BU7UlsxSdMy1Hf3wYePD98q
mYy6IdzWJFlnkcWGQc9blvum9AY7Z6NwC9bHopPzcGfIV2ngGxnQd4kjd1ja5myuThklqLpb2vi8
uPBtvIvepe/7jbYib5wY9QTZLnekitMtuOHcGVpsCqOnQjPqvUVxLZmZDyu5TJMaLklRJc+00GdW
s7Z8qSSWcanrudRUy+3zZnc8+sDIKR78O7uou1aN59IyYOT9LSPAwt7IXxAc2D567BtnqlBZYavx
7/QXSFHXoyhOpyhmB0yguWZ8ElwrrP9VT8fpidIapvYdGiK9X2jbu3SgAguS+XsxvdDSsTdrX0oJ
Kth02VFXIe//DMCWwkWSmaghS96ZTDWFWK2A7LtFujW1WVq+aLoL5/oHD/6qf6/4XchYCKwBhxOL
HVRZVEeYG6jTIo898YB1y/US/4mUup/TTTc+Iwq7PE9Xenjfw5bbKt0EPPuFWFAa64qOWxSpvu3i
0sXq9Btu62qO1KrsghqysM/gBPQStLqVuhMHQYXPspTxp87azpSsAiQ923Kh8yRy0HqPBunWvHeX
SAGMn0sTKVC4WNsdKzSYmTrFPsL5uQZSeksItO8x1mR9+s+5dcmW33DuxSvnyQDYK8eE8bQZ18eu
b5Kd4M6VM5oItB+TQVTRjtjyFIVFwt44x0f3WAESiWe1gkTjnwtnK/sEKLtRLwEztFco1p9XVqjh
l2fRXs4pihsk55xTwcL98Iiwlf8qTunnna0kLNjAiTslrQ8F7t40oiV/vqW3dEGJzGc6fY15u+Rf
0Qs6xt1WJZ6sac0bFM5ixoqO/tMhP0A20q0grVA6B6HhVqpTUvWbLbRi6oBKU+rsRfgjEBQZ37oD
8s0vFusqd9LUSpyDQiVQ/VjpxjSbAgC73pzvj8lSZ5iyt9cMDsUWOQdvYeJcsP7S2pq2CRcpWwiW
8tVF9RLd1qtWt+LksWge9BtJhAZKRLr93nsa1NHpEWk8mNonwMEgYTtiw/pwQiBSDluUpluber6I
KgPEHNKYU44XuayLu63T3mtHc1RQbhGNKKsgo3Med4NqZimAPWxM5v2o68vkGm6eMGdV4P17/K2M
eJS4jW9/XJvkyOxHsZoTQJWmI0pV+x2pozQAEJrUhc9kdxomyYNVMqxoF0qBJhwDdIxUFYquABek
viIkXV8ZllyhKm9DohumSLkRkDBgUkZpOhTVFa0heSclMCEMfZgTXhaQtmASRePXH46V6HcQEcbV
Hj+UNwaLvTmmvRjPJpjHbm0d1uKJTJibvjtvu3PpqzaRAxS09KNCEdBrDEPY4L2zoYMjngTjRAWn
KQSfY+QYoL3v8sIxzG2J+4e/6wohnlYDe6HifBnWNE+Dm7EKpi2hbPfQgb0HitFXS1tzYgMQXA8I
HVJUA8LTLaJV7Ox884PfeiqesycUvw578A3/q2wrMrU5aVjyalizF3/+pj78QPoelQaMYsGdn1Gr
ZBRfQZ2ugbGpKLP5B6OAc3yUt1DxMCTQqKe7kbTbEsTOzvr2lU0iHZSgrPBsZOBHDyf30JJneCX1
mMZfidmSue36lubTUjYIy0enB+Nd5353l7v0Ua3MixG0Hk1HxhquUFSbu9ITETV5UWU/WfPXb5sp
0RGK1zU2MVrYtBBiZWt9OlmQGFJIsmPhFpyyIx7vPz05swpc91c4YOO4xPAx2WUkWtoiZkVcettG
0VYovxN5Pa3s8ovcBKJltBQ8UGSLcjt6FY8lQHqp1HRS4wxNNEcIWnmefMZ9MD6iEnY7EDI0ICRs
GaT/FEwOzbg+bs8+VfpMZfJdXPTGo+b73fV8H2cjv/4qTuShJHbIlsgxD+N3a7aFPw1AjV6ttJ+W
NUiDvZdsQPzWG8P5/g5kZ8mdZffRGODhSiqHsc9Y41ZOuF+hi1kl02uHC9Nrqacaz/zHfwGOvXnK
c/FpENdyDdIAOj3FXj27JUX03/JIQhRJ8It9M55Fhad/68oiopN3yCixcZ3L6ZqbKQpHe3hOzkUw
axjBMSZAq8IVH8LM8gQqJywGZWGRvr/asakjJkXJ/vkJThUsWhiF63BSeZRNG/LZUSpZYT60d2QT
x8oxJE7VdDOFOGsMQzSCimpgEhptst8cTt8TDJrySBBaXe3IOHHvdgocOfQ+ZVE5SaJoZu/Sd+Hi
06eoXcdf1ULVGz1B5ggo9LqqNa2nbSpwaRva2nslgKWAsIGHfLMBC0mEBNEM6/ziVlWw12eBtEm3
jF+g6K1IqTqKXilUz/WJmGBKaYEEsPDK9TjHSX5Fz9/mDBI0BYqpug+U83BqxabmE7WkOVyfyrQ2
kUt6fYkQsge6xev6NfFCridK8syxlZZLeBDfWP3cyi/449Y+uxC1KaGWBGRoUHnwPnyRUFaSUubd
kBct1PIs/yP9+uQSZns0COaJm6yjAVndBn0+EKAWa1lduMIZcBxS1vd7hYc6Y8hv03GaS7sbVY1+
DPX/ts0o9Q2lp88cmHuWEWeB/TTRKx9QPCJaXXsgqCsX12iw0tWivghWCC5sKMSQaQXalLs5bhoG
UlqpchqbahdMdL2AytBYwBu2bCSm024hTkJ2bsa5l2a/WKL7E1qaZxedk2CPXtrmB7i/FWmslaoq
GUKG7K+xawNAFtEzni4GVLmkqHfd/z+ZTVoIYysGzVg70UwegDX2bW7QkUI04asH5AUw1gQDrUpy
6VabcnJEJ+2O3lp5u3ajd8GkwLuuwxAbzrBdz5ld0Zrtw/GK46SM9ZX1RLwIN4S4eZBWl0X6E2VC
F36EQ74dgok1qR/zWHlFe07HAj/B0fWuT9t2cdFZEG5fZ9yCbiv2eK6XXfmvn26Mi5nfy/WBofzp
66c2mwqNJ8/b+GRhqWeG+BLI89H50Nho8sTSoAARqsK/aBmoO486LwoR/81mEvNJp2QwDnOL9uF4
Hu8i6b0xSkQS7/VNkVoPOL4gmubualExJPXduETejYmVud7ypiHWyCFUrJfF3ILNybl0IxRcDhHx
OEP5NBvp1issKOwRPi6hrwBfa6Aa9Eoa0/388bU0a4sEFw4kUnwNMb6sXNfHhns54+am4sTGaDiK
INKc8upxjZ/Z3q7hI7lyq0m2yb+LAC26RSscuI8iEj7HN4HYfrVgokT3chQl6zrlPJ0Rdfho7e83
joWqhVnRtaBCpDLElsVvxkDaQp2oJXPjpHj/zeQYcp55fFTGbc0EkXnZpDKfsnN9k7I2nUqP/ALW
4y0qwb8bzlAo2pSqsKBu7nCQ1FfkJNG4mMHO5sk95V4LrHozAs9rUJurx+HyBVsGnymu7DB6A6yg
gnDof3h3Bd7H6PcD2nRVATctu1aW+bM4Gt3O0pcO9bfoh98Yc8AmVzcVasNOB/UOMx+lK08cX4XR
1hpbvhdmK+Iy943Kh8aqE7I/AFcmJKWQegudQ5QKobCPZMVdo0TTNSEPHz/64loV7Cr+4xMDy6Ei
emwfySkT5v64cLGiymA4A+PKsvhh+GvChknaqBlCyz/gjaeokSG3qcRqEYy44J1l3AUWQUBI1aQ7
29XMNxDubpNHxZCmcpyiDAgCIIXM2wzGmbEJDZvzgErxdh9LninXbtHxe1nznPlVBOUoEKDXtd4E
RxyZaAeUIrG4/q+FNoj/IeeZXFwcyMO8AVxumvmqiATuhOn63diaNSq15e0REJ13po4wCRk31No8
Fl0lvz1qzd9pN53oa1f055aEg0q+YZ5lmoiSgjEUiAh7QnoLLxPo5fuxQ1NOs7+2KBQG0ieHWRLh
PT4mYiAtApp2UHPmw2iZcOvTIwDTqTDpe7zumRcTEfBJbTGpAfMVirNcHSfylSmyTQA32b9TayUH
Dw1ksai8Os//jvnOUzsUvqkR38jL8RJzcCUxIhXwmInRH9pnk6Uau4UrS6CVrHCYh/kfcYtnPMMh
r/g5dIZNtBop4ZRssXXwrrrI6agLyfXMNRBLJgKkONpvlSOL4gnATtP21GTUKLVuxyjNnq0IWkMG
xjZCokK1IIZ1j0sAsrB7/ZX0yD0Q633qnmd+rEQVbcedCLoyPShTDmMXmNAMdI06wa4vnj16bwj6
xmi3353xc5SCBZyV7ZYDcF+AyHX85SsIrs/6GOuQ6sFXpOTc92snojmz6w3Mkv/I7jdhavHV9gyn
cVU2UFICuw64hNeCcl+UB8KmjAkmOvmHcoePj0797nMZFMbdKo2vMHVYDNK1i0XBlVV4sgiEIN2r
wNCe6Vpk+zQxgjFBfwX/kz/A86nvOcnqSJ004FS9fVrA7yiyRNNYNEG+yeqOUowI70cqpn4lqnAe
+ajur0XE4LQxQuhsCiMY59LEWr2nWLtWuDIVXnbmrH9ehocmuBxI3PSd7lt3vZ9O1plT3oYTg2c6
XogGND/TNdDlXWxv6ubA4CGnGuXYAxVZzl56Vqle4P0tF8FyOZ1J47RGsLZDttxzO+R6RaOzKcWE
s/YxfQfyAZv/f5nXiH4sOZMaIBs9Wrcdf3K5L9xBVXgBt86Rj+Y0Ms0CP4SUlrOfBtTe14AAfvBR
owDHzL+e7ttpVuzfR0se+N9G3mLwrLyKoEA1OEVaA7Yill34boXWQLchpgBZKSESJLLF8f8Ox5HR
0ddYVuTblxzuHFNntRGcRmeHm3mad/SdU8xHI4a6dfaoKn9sE/Pw0xeV30kM6Y792oqja5zyZqln
P+5gucx7aIQkAfX9yXMF+W6UrzQykuKtWX7mpAv5qr3JQxkMvW9wjTUsXisCGrw6GOqg8W/GQhop
bjekv4Seo+3Rmeu+Bm7tW6R7jAcEqAT6ryNJsYVk5VGmwfXciDAhGMRlpdcn9nm6lnvfkCYl0N4J
sEP60bOJARb8NqB7Qv/gyFQU98vabAJcMHVLfUFjju8CYpGLg91dvEZy0u8Mge+q+7k1qODozKYH
BnmWkmltkK3W6XNC3J41yInVFEZJJSqJn5YzLyOptzjI5pk8lpSoEHMtPOgAuOCLcrDbHykmtW37
EQqUQ1yXjyFdVAUE592+nrvOkyhZakaIjmIsYOR0ptEls2Fk74zmGQpCSiKYZCsGmy1PsiuZmJQT
Cf4DkKNlClmexIGjwjf2d7qtw2ZHt1TRTRHsXr0QUzEobiew0L2+EzA82vLHK9IymrC+JRPFf5to
0i2DIdhy2Uai9BEgZi8rR9olr4NMN96v5rj6KoRQDx6oXVPtY1G1OmgSWoLdj2PWbstF4SFHZ3mJ
4iMziuyr+GaUDu8N85duJM6b1+pEVBXM4oIrghUkR57iu2gZNDi8l4L8O0dstUk2Wd1paVywo+JZ
3QZaVQUr7FYqiHt6npkB2L+VZ4IrqtOSdxL3uGCHG68m94zuJJOtpV67Uo+TI22MnTBLbMqsS/MN
CrQDF2/VNSuZUbDtT4GOiNtcgp2/C0EYnpD8DE6gaPowZt5WAUaylqjCKWctURosHs5jsml2xK0T
IWVfSb36kz88sFSQFdLyqzu2BzVJ0PnZEBhhvmABnL+7ZuoURnWxGAInxkg1tTaQt1D7kNHN7xjt
GEbkGQBRFaH2ljK4rjJi70+p2tVWDOvyy+AmflEdRxglDnjNzVrBhspr9ZKXr18KNKuXz98HtsIS
XMoK4Ygv5WMu/uhIt1sk+pwoO3k68bGHFuJfITSDKqpkCfHGDPzHWpE72HzMSIz/ufpFdrhoQFuH
+6S0+Z9uNkvvAuj6Ib37erK9VxM4Vn72p4xk8QUFfFZTpTRKIXkNBxpQWrLVgpugdTj5Gd0cewCK
rpY+D9+RlVJqqypbiHv6QvBVUV6FzEu5ujNX/OJ9I07i98GztEteEAoAj63a3JB77EwOmY1DkgEr
Zu9fYLb2hwMMpUfv/oGD0cAuicke4z6VyC7QktjIPgM+gw739N5moclXZbmuU23azy8OkHsFDSUd
hlnHXEs6/HZUphpCEQQWZSXlzsiZ7vxAlBX2QdhXSW7hokZRO41wOREqGUuVfM9JxVtH6jxVv9jC
lS9DqjrCjh9ZNi3t7BQUdHxuOnRZjMEirMSBFs5q/dC6ULLYOv29hmil4xgdQMxxHiH3fHfFPgs+
I5Q/EiPiN2+ET7eTzHAJMNRrjqk5aLddCaWSGLlaHhoJQinfcXWSouTQmtlak21i7jcsILdiIh0W
PCZXfpM+m7+aPQg5Wtu4CoPxKfMZc+aj70dbrVktqFfYBfiq+krHvctP7MWkOYxTqpTAy6t52Zbv
NqzrBBnCVx1CyZ5l3YtjvtDB1pXsJ9WXOTfhivvvMKkTyxEz6NfqNA52iueEOdNciWTBMjMlO1/V
vwjs/8n0dT+rRS/FhNQyL2PsOUN1RZF6aw4BO9nd155PYUVgYZMtQteSYqs4HZk7SXzHZIMRatcU
rn8Ky+25F91TGnaP92cmSmPropqWz2GbLN7Te35a6OVuRaA4L5kLB2AljDu6jus3YOe47Ml+4uHP
LU2Jd6tZ3M3+YpDLRKxEywE/k1mOa39xolKT3kyBtqK3E7h0TzpCGtJ2VO5k311AiJKYVYVPrL8A
iyVKp5PBYiTFVe01T7arK9Hh6YG5BN8wKmAGo6f97vJNvOHk+MW8CwJ6+SN1rLttx6yBPuoC7dHV
M++r4J1kieNgsuPYtQlCoFvv8hnlPoagbZidc8pHzCduuH45UxbqO3nrYIuyzLKUfqMTgtJLy5mT
Bg5edwmumOgk9u7oMIFVEqr/B3MX/ckxZchOl6ICqtI9snqXhtMiLGgkvP9rdr/3GtdCUl8/se8K
BDNYwcl+nT8PcYVHuNVklEFFC34aWnQIn6Km/5HxCTEpMRJOliWmI7cNPvb920wG0/qAIVa6XGU9
a8MyhsTOygUfzSDn8U38SRKBbyAjB6KhXRQezEcDFWf49sniCKmQTzRUQLwd4N99bjA1nYVCroqr
+tktONQbviQT9piFrMXRj2EbIOHMvsz6tkILnaVM74PTEjAY4t271fvgeJeFN2X3t6eormSpOJTQ
vguTTgASJqAF+BmGZwJwlGjTN10rOIxHXXvyHLsV9f/4yfLj4+yCpL5RcmB2YD9qKwKp01fdM+Ty
U1VnDBl115AS2CoRysIPVyqfE6NvR+F7zFWGcF0hecrGgcOKJe3fcPBf+I/XzqfYP697Wb5rR7k5
iUCTXFrwaaA4aODV297dFvYjxfcwd38xK0/xinmKy/HWY4yDF4htPmgW2TPVb9KQBdpsZ5fjDB6W
A9zaVbgfAjCsGPcAlQWYtj/3Oihta4bu2p/cYZQ/6wWkGjW/0bFD9AGIGtsM9nStZL5crak37rb7
fD6z9kvfQuMNMfyGx1P6mrCw1BCig6GK0bsWDVNMuRV+8KaGctk7X7j3uhbUDqadpNCBmaGidKbh
sUG7T4HNpaXeCvP98J24GuqnbDt+mHZDpVjoaPxfuDO3Pm8yoKkbaw/tT0GMz0uoZt5jxVmZ4Mdq
R4+CH8nfseK6TAq/rBi49eL9gJXfOTKEFO0PqNXrVmpzrLcd0KAkcriS+HtoWbSjSqYdgxzZSTCj
vAQB9PwqIXCWHg6MW4PzAX+NT2RMcLc62QHQgGIImwQn8XcB/7LDS4NRbkOVv4lvRJDd+sX5z1sC
SQmvoWEuoV9topMnU30S1K09pLtJ46CBa/b1fRBO/Ex54RIB/MlJ3oxkXV61ruo2M5R1Lgu9UEk+
0+OmgQLTzUj1FR110qjuOyW5cvtHveS0QPi8rjwRSc8IXO6G8uNUl/4XM8tD3oGQBbdJtK4e8A0c
gItc4w++1+TIxLXAuubOOeL/Z6NZUA9jdeMWo00IFt4LOZSN5PsZi1algv2SvWO9G6c8KI/0yFL1
ySkkTEyAqN+Q5cI3OBojkN1GJtsYwmeWyCp1gtOYQ42mIqvFPNYC/NRTXMbL6h41xl8iMHyJMcG5
qMzyJ5HrK2LVzPHnjzOCeSgNLI3u1RuJrC5afho6yhE9H4adSzP3SNBmb9LrOYWKwgJJbWbh31wT
iGcDcQEjuYbWAO2ky3DCL7UaD6oRZod/VEsXAftsGmoUSDzhkYd7CsvRbHzpBvNWnRwo3Z9baEXZ
d27qIpJw8g/lCVlN5KVmdPhtPg1D1iHYmSeLCoF7Z2ZoT9T0Y0RTf6pieZTUlzIEk7eUHU/DvND3
cGsTUvmr7ShZEAJEmJORbNiVCo82F0hrQo5mm2/wPSv1KIEJL68U8fdT3dhWao7ooo6PmzbZgGkG
FCD9b27AoOz1LtkBf915kLw69VEKQbskpcejy3CUTTujzGdmWavlDvCcMWR3bfw2wmkas4lPubiz
sVd76BpoogIl6LRdGok4pRtQe3YvrhBJgDh3LCCGTSxGdkZ1Pf0yj11Kx0NKRDphVHd7VXRIygXI
hwucdWe/I4OkIcj6Hx529N2j7MtAiUu3lfZ6PVXJFkCKuQrDJHih1BD3F2TjtdM79j74SxVcp8aj
98raHd13GPEca8UVtcmgHlJKoflL5dq5GW09UYzgCtKygCc9eHwLhrc/fdp69Ir5KIJsv0gD2jFJ
3BB8Ci41bjsRA9HC0oCarTKXqVZ9ZAgxkJZ1lPwy9TNfI/OJM672qvaAXGEyZHzM3RMizPJVJwbm
1wdouyno5zwXVrz9YfPDRSw3zdaQv+JHTFh6M2S1PP+TKkoNwXsZ4Gt2DQCY7bIZ3ysddzDZzy5w
vnachDJNmTHTOGYoiMNotOC46j1UuCcJz4A72hXvG5wNB2sSDVAh5e4vVVuJhguWW7JsKjArhVWi
8hlvqakvKXNDV8qjYhuF2eW5b4OOyy0m+l4Q9hnj5cIdUpEKvOF2vFxLAYrOAl4bZhb0St1fTkFO
RDVYWwnAgZOrJ7qPpMFH+WqoHhJhlW0otpfzfPnhwtecMInDlw4LEAVR+blDqzA6qPPV6lKk0AZ4
R+CgL4v6uEoEA68pGD4cXw64cMht4WXin6J+xXpLkm6MIy2TsY+cNj4a+enklAFzcLKTuV9rG2KN
dxy3fMn6UGSJ6q95GxstLRR7mmKqDww07c8cghHPhPV2SWODyUaAAYFBZnXlHMIKdRwaE1TfIhO1
CGV+kI2i8cFA5jlA6pFdZIfFWFQ7H1swAygUXHZtkSS5ySDlxjHgdTdDTd4FLr5sHmLVoLRiqcvt
fDtOJwX6PPbcVKQQRtAQAAZLfL+Su+ik8qRbMljR/4oc0ywSM/lKVHO4JC+sQQeG049mNJ0f26y3
jDlaM0sXVp74DIj7nMX2DTYiZ5lkgwUlRTn6CirVLi5s6i9TTX/MIJlcC0lOgvEVnxCtTrX+hI0Y
jw/GPLOQHbC+S9TpwUcNUp8BZwtnz1snAUV5TPmLC50QRe9xUHEjeeCg/BXrQTWVCOjuEICjhl9U
1b9LJVKn+l7KTx2qm0N30frCkdEjZvqjs4A6YK4jX2n9LqnVoDyFNPWmhPBz7Th1tZhB3UOv3T94
ANpCeS5gfRvQh+gZK431ehyNfQ4rGMdJsSc7SafK8P4ouzFmlB3bktC26JdORceiEIJls25qv1LN
AJ8bqNJpLfJvA+VTppnY2tLTK4xRPmth1Y511JDvzgtAQNHMo78V1JUzsjudfYgoqt0nPcRFOwAg
gcOYTo04+3Se3bZBdne4X9NSxDrAc9SWXtL0BsMG8noLgjMM/hfDHMnBtZuhiKxHmGUdSbD2Yf1A
hEq3F558ZYSPLOe8ly89kb9p/mzcRJglw8bRlpUJb60nmNbm5eLGdLSUe9VAGyIdn0+1cCxS5dv9
I3NzuBMKI/cLEhZNuj+xXO3GwOfgpZupxOmlCvFImSvLdb1eOMTrECWzjv5Dk/+VEhs8E0yGPoMd
COfpfehmFXfTNoSIt1rwVVOQXZaU3jArFgRcePiWL86Rc+/iVNyFYn5OCKTjvoegPlhtvtuPb1iU
mXzuqUQ+H5s7w1wF/acUu9O618vNJMxVABfynd2eEQdkkgwqPduoXgP6OWNA4xbSBxtePLNHytZO
slQgvq68vdkOtAi/jvxCtSqTI/tksB4XKQX6ZqKdM0/mf+ZRAuF6Dw9QP0yoISlNVDXpr+0u1tSU
M+RwzswESZ3zH7UkzJMU0Poa1MTdDQ+UBNXrLKBgpsHR1pr59FmYo+2yTQPY142ad6LLzbcl6mNd
zaPhqTpZDzhNnUmbkdUcy1MYP2dk/JRa/slhfzSOcsduHR9LFcYKeInGrM7zoOa54cQos65L5FxU
a51KsvTyxqxuoxCEKZZiootVg60edLTLJ+aj5ywjkVFf+dzDnrp5qddrPGqUcpRKCrhUJWtntXNN
U3jZnqoARmFqexs+BW4enIaL3Ok8ObUlJiCgRuwRWq3M3Nbk2AuA5Nei8gem8k1zPJsM/6cMEPZr
qwYBjXRM+D3Mr2+MVG/TuKdSNOT4kcWjXzb8v6X+uIIeFdtde/Qj0ZgQevYbhLGs5L7ADW/1BPhY
7/o1eHoOiGDYGuRccZi/6pp3JNh/jMR+i/nz+mOhkph1fqM4KxxMklG/Y6Nv/4mn3+9jxsZTrHjy
59V8/D8B7eUJqP3nJsp4rYkkwRi33Msu4/eB84zEJarwkfDNBf7sqH5Ny36CIkdPiUoUOKQM/ada
lVpMzDg+5nYXwqAxzMQ0sHEir4UvPw0kaDsYCn9Tb6Stf6k9oQGjIpxc6z0bhqkTMeE4Msrxz0Sr
Y4MmbZMcWdqHN0REfiBhJJImWlju8rm7aFKhMPo2fheQ7AxghayTbl2oMRCEXp2ci4ua5YNFjc15
ZUkS4U1r6pu7Tieyo2vROcUJfke938pKi5kBibS0xcG9g7S8cv355dt8L7dpYFe69czffao3eNDA
ytL/Tyanu1i6n0IQ14W3p0dEg1UFoLWQ+2MdxfD8hkoEI9QYhBkM9/YDmfQh1XLz9Xs8ndAgXZ1h
hjILzlm6/syO3XK0e8/NA3ejZaphYXO4puMtWN2Dx/7i8iWcBq6FZnXHXcyZ0T+obTeC/SM4yOGG
w+TCx2qzYJNknB4o6jiSWpAOjfFWTlsTCIQQGzDok+Z3LnJ7t2aLzw7igHYxukZcI2fFTlnLZ92e
RnLyRnEU/8L0rhzKGonFs5lvjyglzT3Z1wrqaN+vLRbO9V6jT0lctfCl+Mhz4yaLg9dgnf7YwL9g
elU0R4b1r371/wM8FcPHRgtTFqwYiI5TblhN8AKsUvF6Em38IMJj/15XotfRKgaO3pc5pINB/KqR
VSjW5QT3C3RDsp6JGNpuja4wYQEJmFtPDpaaUsGgnNqFYA3CtmuYDVV/BtH97MJOwhirgDwtw+aO
fPfZC0llgAMtNvADVbGbMeWnkp0ikbZdrBZvtQ3wNmA8y71hC+5asu0wLYQLQyjDKOH/WQqyq+PP
zTpPvxJW3eOhXC1wJ30a0xWQsc8NNvUKzyzbNN+xDcUrxZH9NL4KaAyrYFeQB0P20RUpVQL45YSk
6L1yswDaJjx1YXjDNcJo5qtzlWvU2mWaOxG2eXMByLLah89AhbWUzgaxfDaeK0pacgKJkkP4t5bT
N4Ej5SrC9CZJh/dB7qcKya/0RbbiD6kaqqSJe5+8+wV3yZAb2QgPJsV6zDlf0Y6EnnwsH3ZzCLL9
GEcjfxKycSq2ubOZHqnAqo0CaEk4nrpTW47ftTzAKKlBqnXwTEq6KpXV5wIKKnnDLZhxG3TDd+LI
s9vcwaTKFeFHd7KNk8njiadxJZ2rq2DgthYveqgs1bi6y/cuPpbB/70bJtJofJ1zMN7Jqn6jqlrc
hOOloV5GYJPxUZObZYtxYIJcV0sWrdC8qXPCVgxaloxB6Yp6h+89/5nNXKIq6P0J/p68J/mDfZ0S
qMDmqH+NFwAvtA2+HlFeAf/7JOBSGfNSvEKhiyr0oalMnrQFwnlxkgznCEJ7nwWTjtP3XdjCfhnI
sy1pY5Re/1qiwovjRWvuJ5binkfe3VIXnv7hnbBeCyGjSZboXma2DuizPDQMC3DDFfoxW4VfWUCh
k4tReWHeqDJwiz1xtg4kNxSUQq6HJpCcUpFpE/BkKpfqowcmNb42xOtODR3UVbUXMH4uS20Jkcrd
bSTYJ8kIqysSHL/HqvT0aoubN4T4sZ+bs+OUFrck6LHgRN6O6zj85yrA84gUex615eG47PY9Xcy5
WbGSCywSEeEgXVm6n2Ki4iJFM/KziP4poiy9QPSGRSpPH+dZx8YfUctFAwvw0/7Exo3Uv4dMygNf
WPiSCKFcesFRsC6ZLVpBKPqHy1gv+uT8+y17reqoYr4Bex/2KeN34GcLueT7ShyLt3VGAatyfqIy
T+XA0Gf66IIZZGveS67IfgPL0Gj83n++puU2NM2yle2OpnjVM1huD7Wx3ziL9AGSzY+7aHtbnca4
RYsQGHqLOOvoFA8wh6J/DgcFhF7VIHLI8bSzhZgIzrRMzqkZTLYfdm2rDlgjl9i6pHzwsIKKUD+t
BZaABJ3PYDDdyAyUFe6D7FSbnZiMfzwOkkYrWBZZMz9WNcwovUNfQPutPuvmJ6gt0bAcl5Fe4ut8
gKzInsaSP6DUwjQOW59HaN64RBX9JNrqmUQsxKTOTlAnt5v+b/I9T3A8NN1GcE2/rvxcpqiaAic0
W8PMpdInODbsZ6ytetZuvetOh0PthoLKKjRJjx+7DCGjFj6EI8q/HFEdy4x78jsAslxbTRpS5H62
cEidxZAEkQLADFWX2bJQV76funlDprtUhQR4bMP2Q4iXM1TlLgEuko7h6UQsfN63Wd6Z7cKH42Jd
8LHqH6g8QEIue/3QgME1jnvY0gBJpLBffIp1bY/miB2lEeh1oXna7pA1HeP/Oas6qejWrxHsrnho
uBdfPSDW8hUDhhk4L4H2TSRY6it+ElvB32t4Dq5lxE8kASq/dd3ZD0f/w0CebuV0LHco6S/Cutv6
e/5KDPWZEaVvyDdyMz42T2YSPOsvmXMvp8FnYlutRXrzlqShQqTfMig7KOUEdf9YdBI7g+B4tsf/
CmsvkpQPi8BTEgNQGaqC19ZyfrPhTy4n+tCPB/pFy7YL0qT9YO14x7O5oHN5fR6q+lOdo2rVUKx6
fpCa9GUm0wDhPSsIO58v9gTbqHAV7lhSl7Vsk2r3hxdm6uznG7YBSUR4VWjdzLhulV7EVjfZpP/x
Wcc2rWriI4aGgN4qaIhY9edivleY1HnLjAihaYG0yHnS3y3c588P8RswiSwNIcAtEj1YGVNIXqDV
lPvySbQI2V4Cex/F04hfPHPtOywqd/i40H3GrO5h8BmqX0W7FgKFVl5SmmuvR+Lk8Zokm5h77hnW
mbFnZEFBnnXlwMo1/Fqp/AP/J2fNRP4hWECwRkBZ4Qv4wpkVeMR9NBfKA4HTPDE1iEd0c39H1taI
VAwVEgeJRlkkPbga2GlEp8b239Wb5jagN+zN6YdAYPHUAQf4/DY6112kAYk8Mg5U2HVt6LNjncgD
H1uNFN1nLZSuIsu0sE2khxSX6tWFy8n7tGyv4SRhcMaO66YQmAvHDLTVR62biYnQZis6GI8cYVvJ
08uO0MAoZdqZ6yLtc5J3IRZnTaperprnid4lm8iMCiF857eiBME+R7iepvjslkoE63DgIdabChvW
mU/mg9oMLEuo/+sxQ6FBeAlIBj8KPpMhsH0SDBkJ+cVytBz4DEclO2KGbvpgtux9CtW+IBhWNdHr
oTsDlWVhYYrCC5GgzR8WBd96sf003FZobBbscHvGdzEuUhdxQPZhoagKToRBbrDD2e+jFvIUmXWM
pfrfJPgFJO5x22EDlWrDiQJx+HtOcoFn0Xdx9WeZCBoBr9u+aQvD+8F72MwGSGwd7IRDVYSyxmub
k9VRBg5bjyK7CfcK+GzR9xRK4thU/eNPn7O8isnF1pqNnpMApK1shgEg03z40j1QoyrghB7+sfHS
jWqbhbgZ6f/LH1ODM85N/TAjKBwekEaL8tvx25tXFP1o4PMk5L88vnFKjvXXAfOnEzQhIdE+PXtb
Fsbkg5LoYUiVlqTNy8k2sqzXas9Fotp2PNp/XNu0U9WjB7QSj6izbgSXEqaj4EvqVEku2YMZA5jW
n88nRhmJDSdmevofJVPVTb7H7NHNIYPtF0hz4zLDgIXOND1UoSJWtF3D5UbaLIHWWTgmgKJaXOZA
e9fjGH7dORLGd0d2CtIpvcNQtRr5SkxMvQlRNTnNB4t2G2s31WeS4xsZiqbQWRILEITFO/qnd8dC
96QNH2gjsvyQo6RryI5cUxeis7oT82p9mLShhBRWVb4O1/QxkWURht0hpz7/KkG+eQjLrcxstP0R
ofv90QX3/qZFCbs4WIsC7bNbPyfcIiyqRjwFVtCEhHGqcY7XKwPmdYyeD4yEDcqBab4wxH4FWYJ+
ERMr7WBZyUgqW9lI9Ws/Upsr83x6N3/rWz+V3w1q9sSgu0cmCHLjZq3ymRKDGP7XHhqfX4GXALDl
sbAaabxuzKbXvp0BLT3Zs+Ozx/C0ycdRpkfcrIAS3ORclWN+j9COHesGAa1lUWHrbUHKjJlxWqKF
8WWKdUPnwH4JB4zD5FUlvm8S+WtD36eYPt3nQ99tNKVLLHX6VMxAtICYoiSaaRyXRvxOy2kBaFOF
4tWEn3oJFOD5/wTsUDSmzlSJ2chDs1Z/UtnpN3V8woGUEfQ2u1IDKydrXsiDvQ7HsUfs+KFGGSZ+
mKiBpI3epHUQqeroJStXRRZkYekeCGz4DSLgza65uDiocRSU8rdWfepIOScwN4GS2oZBHtvvXUwW
tNX3ho3QaPFvdnGtWliksalzwBhECswSRJzJDN1M/Sp0NvPdamB4u1YGHPVQP92fKwv46yLWxeck
TWboyQEZC4UUkMtCxfxwVry8HUXZ6RFmJrjnVuBAsm0TWH/+91dPKNqESbHzjxK6nI4mpyLuKIVq
sFLsDmtP/LIehKbaGiM/0F3AcFl/MgTt6YK4+5r9LVJewe+nvb4o+puKa3z5WYlNV/q9iz+kZIWc
rU7+5OotAPUDZx7KvWOmxgmFQhDcBZ39+RFrgEyWxdW1mdxfgCJgpTz+QyuMa5woZ0hbyjOKneAN
3ZD3i5zoS/YPxSMTujZFUeqd9nCm2o9omDleJMr5J5mnCLG/LfzVc2bNP3qA90r9zr5v9uKY9yif
PlSx+Fc/V2tiWiLGku+qMJctTSPCqcj0bIVfFvjb20Lxt3UsW+1/EAnRqXaZE8Pyzk/BtfIQvRb2
zINI/794+ytzAgn/37kwd/ZvDcovbso+Sctzg4EeW6LLY8dxs7MLyp8r/9Oyja0+R0uxwcNI4IiD
c3eLAjFEAgAbuLFOKDSnwn1toLrQSIIBfkvq039o/NDSq4nBAojXK47udxxtZdCDTPp9BzEAoMNF
LY5FDiFAlBrCPNqgzkHywcLwkkbju3w24qW0fgyxvTW+Jy/QeOL6QPJFp4HSAYcQh8pOOIlcASZd
M4gP7FphF0GcyKkMxRqjHRH+QwcB6M7jKtvVQq32D3jH6voIbFUq13LNxyNP4NuosicQxis+aId5
JIFY5aP53wMHdOmBYJLdnaHWdPvmnVbWuwX03vltPBTbB/jOtjMBpf8U0uryKhpDBr5LBVbEEp5X
Revj7jCDSo3xO2YbqciujNVj8AI0DSRwnIxmbY7scS845rfRBreYZ8C7eODVtsokcIpqszwT7iq0
dvI8/d5v6OSxDMneqi/ijpOVVhgct+hD2ecUmXQNmMr8j//vY0mEknR94f0bRt/CurDHye9h+Iy3
heMJcKBiqcxRGICwXiC2733t4QZwt9EAv7dEqsPTk78TLMKvuoBbMZpR+4aZTYiBrEOoL8CAzxfS
0g1cER2MoZ+zqnPjhTe7k6XbYRA9YJG/P1vLyLP6J02q2bHZXr83cjrCF120k5X7n5iyci01gzVG
pVrkpKa/Gm0T4m1uxuw0Fwh/Zg4g++PrJ65NxWrej9P9piuOVNVHlaZiNHIeIRM2wKUPup/jC0hw
zZhqnKJFlvE2AL5xTw3E0vW0gorvyGTzZY8NfYWulBBvG3N7SyGwIqj1PtbJ1XD8yx3y5ecbuTFS
w40/95isRpS3dAmv5mwo7XFqJ1XyBXVZvvS1UFLz2mhay8IF+rzpKYfdmHDECZRkyu2gg+6iJDGp
v+t95SzUuT+LoVzMFVP08Ffj6E5ijHLffHIOrinwlhxhiCIor7rhxfe6lJXuPLYyK4dUUaEhyeew
uduF/rECMJsFfZmnvUgbC3HCIumb5ciV8UoonMkbrrvvawKulQEG8GDyQiOx3NWJSTpxzobfeEj5
5r0eZCeKkZ7+hXJ/0i3DEkX1N25BXdf+nGoNC2/LR6VSQBAJWOpeGTHYCd6AeTb70EaaX0tGgur3
rkAYw87WDomK+4VBDV6FK7QPsQoEU/28NSH2MpffkxlmUE+THxUGO4U2wILK96vXzMJaHEqjzJwP
6DLmj8Vwh4Sp39fMbrpH88DVEKKi9YGec0Cz2ofZvl7179s++LcS2TLq5aMPce4mwQ7uJH2IO5OA
v8s2yd+aQD/GWf4TguwR1qxN/IGZmEkDsd2bbDBAuC1Ed1ftr/kgm4rSWHzMCxbcVTBLPGOQ+ngI
qB3wvL9G2cLCS+P3AbxtI5kJ58zZnoWmRa3YzT7XuAD1yoGtmEJD0w21UZ0sWCM1gCMSYilC2mQU
0sR3/4avsRr7SVnSNjgsXtA7Llew6h8Aiqxc1MV9MFVShGCaVKVIiUNQiPnuC4+kXlCJJ5AsYya7
fDnTDAI8vmpVUszuFCtlEMmEv8RpzC2NsgQDj/b3rIZDelS6nIW4341W/u8zuSeM7YS98uVMi1Vw
bTNeZGrqypoXBk8KWciadlYkI1GX/CJXoq5Y57742+dL/cPQAXnGU8WOtosY+DJTgsqwQI7P+sxU
mi5Wm1qRQ07C9UWMfinj4ybeNseDzeAY0RuZ0hSNXpfMUKiFMWnpl/q73dxMZxu7hn4smyjF/IPH
FGTsVT3+YTG+znWm5tzzra4kuOi+cdZ7RTciOhx4NVxZBtW2ytl1vllNBUGpMm+v29m3QMUl3h1/
YCEyAhLV2DK1Eh688OfqDT3jUtgbtAX7SdFnAFI3jKLsbi+OayhtNP/0ZkG3JwaE1Guf29TkZz4f
VvHoKaF7OVRHE9VTzHV/sidRlTptwCIv7gJINk2q8KgTBOKPXMVM+5Ji12i6PZVp3URzYjuXELum
Q6oN7qvMG+wXNbSDVLA7h/93t5iClevuoB7MJ9QKl4gSlaXqwK268nZVlvOIi1N/Mjc0AJa+CFtQ
+64SCpdMfoYiu5lcV9yF48szSkaryrnTRvCI0LOxkKVSK74hGEIjc5QmQ+JrYkv1tGX0KDFkq1Ez
etEagcgSKVYsadKXz/qZGA1MlLlYgq12mVc1dX7yFTB0C4W8co3tjHAi5T/VIHxssNorpMs5f4tZ
2cTbuHAFxJEGbuFn/ccLiov6hCSDKF1ZVbZmRY03nbaVRGpHK9GzYxdOcvj1wfom7ShrnBONaais
5K0XA5Q2a8Ybqj5l0153MUQ6CeU03xsn2Otk5NBR44dvJfpHJAXGlUJUcpMOiT7nhtaQdtwqBROo
9r+7AU0cv5MTGGaclKG7Jk73tTSpC6jjAyFcOojv5ozGjdtVx3NqzZJo2Ufe5IjY1ypKRIx254wg
pdnJ+sC0y4xnbFwzTihPxvTXDejln3Y2kWlVq9MwHgtU3dO1P2lW9s6dgk59eETeLLMUYT6mNYM1
SCTAkyfHE2ckM28E/vr0fszHYvzOXlnMdfTN2F3D7E/G7/5AjULQEZe3sfgd6LroGTrd+rDf+eJd
CJoripcxhEEeht4Vx3f/yvxoB4tQFJuC/NrZkh01oKVEObaj7/rkVDj00+dU+akm/E1LH/xbMp4v
U5xljruY4BC140fCj/ORP+HCacSMAxeWtAe3wNwtaZ8K6xxeN8zvhOjMXjMyA8v+0OP6o3hlUwEj
dpQ6clBvL9F+SHHEOzQaSJdr8UAWd8NuIiYwLitnMF6sIuxLYYLDXzONDD9GvMxMJG3CdRSbgENG
T2jrJDIZUgmDFhACYr8gwpjqgzFlA7ZOB5yvXzmBAAN5FJ00vi8pVm+N9eeFkMfA5vq2dqAHwdX7
0bQBp/fNCVGhSTRiuTkrO1i2MgAgLEKAoy/5zzNYgupZW3pPb+58LFtpgwPLQulHy7Ig4Po+2hbW
2TGC2B9xQatwy2+vn3EPRxbYQFnyqqwt0Vn6MHY8hlIcGNbOkQz1knC1gqu11Y+iSHmopnsWdvXQ
z+xIM64J8Qrqce/EaXLxnDzJKtxJPiW1W/a6+6EyBXAn5zKhpXlj66Wa87C4GZN+be4nCDzHzSXd
giISYQKplvwk6PZZvc/Ql6ba0wXcy99cozfb1jKOOwyaF+kM7Ad3uoNG3VLcZGbxFPO0PyvbOpef
xBoSZOBhbOMPBJd5Nr9B7UiIVIHgp34frj+MHGU1scl0SQR1V81BFm1RW1WhF5p/0lcuisCcJPQT
hXCHW0XfloDsj9EPzjbWXl7c7Iy0jXkDHLpj/hVmD1oUnkW/XuI37nMtQDQ2qKR9CyMtZJaMRpDb
ieP/J2iN6hBr6pCdXSybMfH1kVt7dbeHiFn2JqYDHq1xd4uaS9Z4forbnEf9xKDCbmnPI8mhvQk5
O62lPafAFqUoktP8WDJbXt+FrxSbUliBY7OHjtm8uZ5tIA/8b9UjWCviGS8uMQREaL0iflem+LFA
tVzJbgvxyvdxL+haxta0vza6CcnQMdsBYqcpJ5JXCKW+vhdqRqlgHIHc8e4ykxdOlUVEMvSeoCiT
J0wEVRpHN0i65FJQqKeV8j+9kAlRx9mztIGQPFevFlW5bC9Q2+nvhqxYljPOLcS8xyNRe6WS0jJK
sPdKVpPg8zhomUZqUABlsNCgqTQACAL3JeZSddi/Dce3yp0w1Y8PsVxSaJUO43wZ6uvgFA3yv5iz
mOwAQN6ZcHRkmV6RIis3QhLWFeJJYEAFWCldRrjMF+XqVUE+i/O72OJzd124J+yBqpkm9tnv9Ocy
Xtb5H5LNSBOa1xnt2MmR40pfNkUoe414eoGrn+enI+FqvM2wRvl7nCbPXg3VFUZ+AOYN1Cpnne4r
o5c+ojHTXvHpo55jgnrQm+6jdjjqVHVl4srvjkO94viXbvzzfkJLT/PQHTMyjOHZBstwsg/gsHLY
KgWZXO6dZRdam8qGCz66fe3cOZHgo+nsfTWTaj2W1OK6JQorVkrokOYoeY3QFc5pVWq4w2By4FRW
l08BQB8KIaVOZNnIUNKZHfJqGC4qNS/RnXPJfYu5ipmiscJbj/beFfexC/HYwr9y8kf1rukFEsye
CjagS4mKUSXI8XogCrfjjysFKcSnXMWb9Swle5JUve43hJa5l/H/PqEG0nULlAbAt1HqQuDN9XYG
+A4q6dVQlSxW9M3IOzGTN3FEC7Ly0XGP7wErKmX9sVpwdmOw9xhhni3EoVyKfNd1qb1Pg6sGie00
CJHdGI/OjhlC8qqQqMc1O4pW/4hW9wQ1nyITEXMDwgWtdrJrZlPqQDd2f3VYoQkg4fueLMHDuFTs
xjfqTMx29kP+E+8glpjDEpMvQkfbYe4z4Hp6xKLgTs3aAz+iWXPW+LMQv4EXXVnZl81B2GyUFGLX
1a9rTJOxQJlKawjClo8bfdkHNdCWn9mKu3IxoLRbtPZ//kjtm5tgfSuh/zkDTCM922ol2Iu0qkBJ
P+pGGx4Q7BOxXa29Jcg1UM9dXUHWZ+2mRQz3fFxCDaUfFFcH1PxVTOWJa84xY+pX4LpSVhZav3PB
a+UfAXpBhDMhNVd4EvD8yvPMUAht7PLdrARZu80Qr+FsW+y48sji7XTMsv7aPEwbkmWEEPKVNlVL
U9z1L17GPzyHRl0xvCIxxXDrCLjD78q63Ci3DY4zNEtf3oKmqw0Jr+ku+VF5TyWYCQ3Q3wXyx2nX
cQeoBdua1ahjskdMyXMCOB2UsIupRqFtn5KgYR/x1xLw+G/QIkKEqqLMrkR/GVgy5RH4EndyelMM
jEsGWWreWgwDLFL4jKQD9KDCdPdEs/w5fpIozVe+Z9kZ9MispfcyAA4r5u5W51z0iN9UFcvQJ27A
vJk/lZFRb2r9Jm0YT3ltAHdgieZMlDXiR9Xhgpp1kk9z3q95GZBuO8wKwGZpExxKrp0XN8zDCS2F
7U4FLi9p+sxAa8IdBPNyd6B3CHDF6nFEqV5QedhcGDTnM04jRySL5IqoZ+QKZNmOGng9JFEooUpz
bOooBlY/tCeRjGLz3GsMif0Ctm/+lAejtaJsRKXyrNZzmxUU9lxlxDLIrpfIdpjjfGRFel/q8RPi
yb8HQ7wav1uT7Jzx8kQj7yr74mDRhbUfwK4xLit9/TpHbDwVpMp0VJsakK1SHjgtALCM4dslkCVW
xlCRJ5GKVoK/8UP1uJRe1ki+DP0vMBCW/MDY2qMQLaFESU5uuRV+vYww3xAt00SxmyBUl/uYbuvs
7LSAdN630oukH2oTQYqEN6r8cDNR8Bbtvp7PRV+Q1ucQjo7D7ybhcB7t6fDNd70uZFs1DexWCO6G
4MtudCgn8y//hIARLiYOaADxj2SnG/wgo92C6sp2G+4WMm1szQu5sfW/1YPGrg+LiXxqqHU9h8lf
2Z6RjiDpSP4U7v/g8kvLc3v41AXKY2gfVSPXtVNyuHrwvl2RGDkYcirMDvFRLOB9AaW2FSj0fAxK
HG3QyVIUCRYOb4gOmvlF89wRCxhPMHWBh2exNwflQDHgzx/xlB55QG1w0r0tYtXQ8ufCyg+6JXPj
1Al33Ka2eJzcOqsxHMyh8MAQ440vtCXO7yMadTnuNkLZpshNm7ccDwelal/lXz6L73JmLOUzvm6r
yxszQuLBBrc2aW64S+nDZtifsK5IN7AGXABsYONxryi1yua2a2HQ/lOwXp755k/Huv0pUKIOblzx
rB/iSNRfvO02rQX4bFDgK0tiCORL/jCDzSWKepI+sqclDMxLVUhPCx9UUqwOSOTOjl3itBaskFe+
C3LRhsxmUio4lIww+WHspdMReHsL4HR/sy7trE4cOwDD6Bkex1pG6fZGi1ZNXvE0URIIf+x8KIcq
8G4SShJfS5iJVoIvi7sXS8TK7touNYFgqAOTIAoF1mPplvnHP6/XlcTJHE90G+KuiRc97y2VMFgo
WATm0iB271oZVnl1Eooigzzolpe5EHyP6Oyw4Awwu3WohTmCAcQn3IVnTCw6w82VASzFgiji8705
c6DlLKQntyIFWIXhO2Dk8O3/tjc+NJzm9DM9HpevkzepbipVjkqYQRVIY79JKE0Qv8NDs8COB4Vk
YxabKtGijWcxkgIkALTYQZTYGE4PYvnXUBEpV2m0Ij2Xvn0t/r3fYjHAoesKP3N1dldBZDqcwesn
DHIt6+ts/4b0QsLq0IV1XL2/Q9ZF3p7em216jQaUhX7o6/XBKVBqALI1ER7ru6cfGMfuAUti+dKa
9QaXL2VCWdxAZ8KoOCNhTEM9O0O7Z0V1duJJBTYyZ0pLsQirITjf3QXaPtTsIW5fzCU5YWp1WDyu
G+ztVks7q1bdUkX+pfFYF5arsgLHjip/tRLlm4OFjX1RGnEAvd97ZIlvXm0cZtDufrf0ZzAyicNF
9n+iLl04WVoF9gjTwn6HVkzrXeslT71MWxs5+eMIB+kCvCpiH1ONUdvZIfXzEGi8tg7z9KR/g7Kz
pGp3MXh7+px3JluB3tFTIxjRDLrtPsalJH6yE0URueB4mDwtgUARpmtEkY3Irtm6aGxcbnKAHqnq
wOh9fe4WtVwTIm0hyTmlVt4sxAuSNiu+HqrxeA9lk/s7Es+OYLJ05mZ/YzF38qfe/lSjaLnfn76N
RUPSwKlQJEzwlTApoT6KoiHUj02Y0V173FeiMsQN0TriYdAtNmdtTNPsz6AnO/oLaH5KynAqgmtW
1Z0tjndKHc5AlK40VKn8U+N3bOkvnqpiB5SMAj+CwX9HemB8l5ahEHdW8AodbHleYIQRO2YfTYmb
V8z1cFEgMjqe9hAz7Leb3lbqNUnRrGw3Ag+mnlzsXv6RYv6eg3W6FVJNu4UqUGrW4C/OpE4lmvst
i28n88uaMiTjwxIWuQ5XYa68MGr1FUh0a7gxvpYZDET/HgfSs0VsTMedqsBqe0t5AwSoCt/xYYM8
HTuX8mRnm5u9kFzOVmLwQBI8gy9tetAk7ED+urFldGDKuF4cxjZAr/gVP13BpJmL+v+rpJ6bhbQ1
M0TWngMz9pOWOnkHHjiQzqvXfykaqGuaxpAe0h21vNhBD6q8LbR7EpSz+bFv7oXId73qOKynerBk
YxbprdjgbIiZd3T9jbmfhD3aPY37mKeGCXdpoi8OfWm98el8e8vgdJxu/mhBcF043kE8WFJM9FFR
8uRQ8CGVTumCTvWUVovWlrReiE9L+TFHZP1IZcouS33Q0bMboY6BMGi3wXWeBktHzwAshjlblSw4
JWxPnhgDJONQOOgJGTDzThY5qJe9KFd15NJ7Z539SWMZQwoA+9R73owins1Rk2FooYapUV3Zhx8h
F31qC/DZzQtb73Wm4Fpx/qX0qVIhKdKH8QIc/O3MbXdThYhh3FKXi98361cSObB08GvQoLZmJSdd
I0DDGKPp9wROrKkuOqQ+s2GI4kJAxYU8H4AhiYpdJkaB1fb+r6P4lzgHaQP0hsRB0NKfks+l4QAB
wgos868c5Md8run9oR2n5UVhxnQIFpKRC7SyfrqDISSnm8s7Rd6hOt8DrED59+qriikxNH4aAw3J
dZBfQIYYRcxAiKzvZTwxcgl0l4YiL35wPvlmOi/QMW7WO5kjyqCJ/bLiFBHW4FY/ovc6Zz/auA0f
T2wON46DwJ/m3MMkWGDpImtpiB9woJKgeZmoghyuj7sgGTFrh3awvpNaSBujuudMbY7vvcYWSyQR
3+rVQwWl9P0XoHZ3zw8t+3FvhtqQKDzXRmuYEs6fXHgTWudxpSrCinld2s10aHvMCEjjIGeJ/UjW
a+6TCAWtb1pJ51bs9ihezc7v3W/qOssCHAGS81H/Wt7m0KHiy1wRfx277Pj5BQBxDTkfblhWQB8r
//RyXV1N/4oIASNCv0pEWGf2VmtJSLZMyFhMMnnf812NRGKcQjQsf4lY4VUCT884ltTe0YfduOJ3
XY5E4e48ccRIT2ppmFEN8i/CRnGk7v2uSRRFtrnz7moH1X5WLKcUHaJNkwwC0O8NM1YICfTs8+Uk
Il+3pBwa4tmc72O5/rjrHOLllRS9WYhWb5e4o2+0gBrL25KMIWMMlwuWlGhhCJyk7F62gY+AJqLq
fN+mxUar+CN8K0v7n0rFv7DNd978ILIu0TU8wTZJS1vjIhZD9zPu4+/UBP6W3Ozd2FkhLLYB6GPU
3pWZXUaORrObLTAWECKAka+bzfl+P6mUDVIIxgX0VR0ZnBvMbDqNvQUoy44sGyJogbXMpKmT6yjc
cUAUn1uWcO3jMZv+MeLfC6MV57ZEgUkgtzZH07a2U4IwYu4Tn8ro6mPXTphMM+bC0KGSVtAk0sIt
YK+kqmF2NY9HUW9zyyYflEOe3uol66SJD3+5088g/XVCBlpoUZIU0osYpq3AGmjWJ3G7637w3k8a
+Ot9hqNPLHVxQ3oAZhNCKHILulloWNICBiz8L+kEyX17xuorts8xqh4Yi6mIWRAEECtPNQMrsaXs
VT1LoNlk0oTjqZ25lTegpCJEzWKHVjV64SazKWm6fHceJZkMYsDyN0RAP9gLP+3eDCgfuQ99oFO2
jZXgNNO/StoSLdCLC6VZ08ZB6ZoWBVLZCW8XjYl++tauGhaJb1Ux5WTtZc90Fawqs7Lx/SFNDxFL
WNrjGu3c6iHZcqsZ7FUlLkEZ8CCoyzdwv53pJpJjIcbCi4QWlVntqRg3gG5btWVAhVMvYM60LrKA
dUBHWJedKpkL8tifMVY9QauAHsyaRKycd33DyMWa8FMh7zhTeqWjHK/7L62Mc/s8VGyD4ne9YI5+
gFIQ6kPUPPTx6dMT+ip1oOa7LV1H/zkfa2FlM95VW/C+LkA6g2VblzDPOcQnvsHN0scDK7KWJRX4
tEnHeAn7abvMvbp+ULjD1mnIy5rOv0V1/ReuoWzlOiWqCOHQoyOl/1wSUwseyKt/HZkiAJY6iDMf
TePmpxk4lgkyQctLBvNGLM7bJ5J0+GP+tFZf3KKMSsAXagF0CX6miWr9QxnIPGdA2vJAfIxP492H
QyEgVp+eVXDeNXrqfaoGeH4w1EudEQOnl5EWZMgRJpKW8J8jVbkoFu8eGSseziacJU1rhiMlqH3w
84dYxVazb8nMK5gBQ7FrEKs2hLrnnx4tTfT8pKGNd4+IVS/vqEOcKYyoOtiJ0fOA2Vlu8m4AFYwK
E7vpzjzgWzgq/A9PcoayGf8rPEzF4/UY1FOH5gSxDagcInjB8+eJmdRFrSrE+ih8wkZY4ifs4Doz
Y+1VvMTWEGZqe09XA/ZW9Eh82G0Qn+kHwDczKh2vIxtHoqSsaOug2oCdpUZ2l8QiSqxJStfuleAL
Yk3nZpV8XLhjit/Je1lrmCT7tkqkgdtdn0mhhTCSVyCHSUWZwY4DIfEW1P8Chv0HjS+tHy7ydI+m
LLppxCWcd6coaLhzakOpyVpoNw8zacSIqK2WcUu/z7VN/xdBL7HjyGdM3dos4Rx0qbXnFCOFiyex
4m+NQJR2UjscXW2nEc0Pmtzo+NGffQ1i9ZwtL7CRv6p6Wloy9ffZ4/XkoyBFzQw6gh3vqYxTZYPY
f7EaOGewt86t6gLLdXoMRPty4gV45ag1PVM090wpR2pxClNHx5WZOxDa401iYIlJRsObZPig0yBe
btqOydJyjQgDoWenQ0LBSCIikVdVuIbD9SnbbLhsgHhrEY8My0pClMasW1Ly5tRgggYbbE0/pjsZ
TpRJ0I17a4O/xghkBLbxN/RQJR77zrlZCH+DEQnF9TLWgqPA3VJ4cdtOU/oKBkaepZJ2yLpbQze+
mZzQFaldEO2O1KguLF5zG4oKQJCjFUL+HfeWopGP63905c5dbDxZhtd5ok6P0z4oGh4bpzSrSKs3
XFsqIm0YWpP295aNsOnGssuPSWtOwHQNmqNrFLtlakNwBuRMZjYSO1KIbr41LaEiQQQgmsnAxPJx
HxPLoOjX614fLL3P6z4+9klHKJVvXhiEFuqKs5ejpx6HOdPsUNbNRbrMY95BQz+aQD1v5cG5A92H
oGp8fJCHJ2gEWNT/TQaSdiS90fKbMLHx5CeGV0Bc8+o+iNbOCWXDqUfJTjPtDwg+orb3QLmDoWPd
0xU7w9GeL/RAXMBd233wx1rZSS2tQZSCEE1+Q9LiyjGwnyjhzINwi+Jhg8KlJN2M5y/B/dr8Al/1
AtzSTg2WJDsnX/AyFxNMG7532pqeRR9urxqx/dpuy2BFdxmJ2Bdt4jXk3qWZ+OF3mt+LTH0PwqLz
b9ESvf86b1cwNXm2/eJqXS9BB3DuQ1Q+/DUREIPuF0w76A2q/B4oUzzOZ5FEY/3qyIpBTC6UTpEo
4VDJZ+llNGUw0FSyRRUZC5Drvq+v5p1hrDhTim4lGnThrqYAjrOSIk8kkF/OnCx3zntzEs9Hl71t
WomRQEfJTJwfsdKAFWkiAzIXz1LCLQ9SSpuTmOlejzhv553c0Fvhf2cL0m+HXoJsrjP9yTAaUrYl
K3L3wd8UzrMlX5ByQ7sjFXvokELG7VaKGdhGuDyvccUZDL+3WgLLbaT+Hz0GH7cGHvWegVO+5LAT
rBCyA0LDtDeVm4F4Cv2Iyk4Pn7BVPz1sWHdKD8Bw1r1ZYi2/xW5jH3rJQwF7Yts3JrsWLdrYyo14
1pU1oTKnisb9cFky1Iy7nfjt7xoBZ1a/foKkSdn1qEDy0UeXtV93uTnneVcDJZW1r3aAO3cGqYB2
yu5U+l2RVqswM5ipkAvji9Nf0o2ve+4nbXZu4Wk7gVgaUmgmnhEPBEPXh0we0L5r9O2D9/VAQZMC
eB3VBLwez2xC11JWHQZUTvh5fC8b/P0ub6GL4NwnqEmc/UsGgfa33SqNo7hFdGCAfAi1+hzk0gtV
YQCqpUtOpNdtcM4SO79AI46maE9eKLv3TW815c/NzkkfVEupLgfsBACcx5lIR+H5DuQzk+caN/Nf
7AJ0JzDw+9iBJMoxPYge6CyttjtlWvOlLf2uBBxfJGO53r6CuOVp3HDYbBTPxCJwgLfG7H4+f0EZ
aNQIFyJsipYEly1sbFDvPYMqrsB6hgcIk7YkLLv0TsR5L5UcPcjjSDDtCRgCMulHQD873GZdOQ9A
X1LelvS/PufMJ/BbprkSfzlPsaEQdvy4bHd0a0SRIolLyAKjfDd82AqWOHqByw4BPKbntJ2JHSxV
nVVCdp9yDEMDwrR7oMjWf5+n2ObwWOcHG8WlYRMqw0W5dwQCUCW7NLT7TM/MjGMRijFY6Q+ozefA
uA/xLDjP1cEYPLO9W6oO3DEKxHizym0hkzd4vhznTeiiji7czNhpaeZaUzMiHR4PZHQjtIckpQwG
aoydUF8JGqfX0YKFl07bH8MXxElO265x6HTlXeLParNTxpTUWMNVJok50h0zpudKKyMj3gvY83zA
HSctDKDe/JtfdA2AudqU1t8LiceTg3Q+D/r0USKutWcLhes4a/lDMjfK3/cBnYKac/rO9tVN5D0B
mOs7DZsjuCUTPfLGwhr5ZrbvNNOw2lu2ngezE+uddpDXA3cDt5zhvDK8dEYNmuWi7wyBTZpf7+ow
GJmRf7chYp/5lQk+d1Kf0Z9lACOvLsIU4fhJq7xNNqUPnRqGcVPC5jEiEdMQQx345CqCBaVupGRT
ZZ/rlFD4bymDxbJfO/P5UX+OrvCGxlnISbDACTis2x3u44mQH9bAHUvemhu9CT/pKx5DpCQz5bYk
EQIicR+QE/jdAH6tQFP63fXn66raNxaqTVlKKQb8Tutw0oz5MMaTYqO432CGvjPGQGkbVPuUX+y0
jazCuES5dy+S5G35hUulp2MCTHzsd44TknFJA7luZ/8rSmG8vkRXH60fe6hcdNXSkTstnr1qZRps
MvCXGiTXdeJDjmjX0F0bTpkFIRXV2syht2kRbcKDzrvgWmArHbKlwXOjt3DC0YWtcXah1iew5X9/
g+pMfTRD6DS4/+6vEdWE3lnaJaep0Wb8saMwJUeDWONVVqeh5cnk+KiUwJCBn7F7w4ITIDBKQxe7
b122a6sVVIhhifxXo2TYcnWh1k580/bSC+Gk28n4y4q4xjgt3Ye0njVg4FtF+ODthCaG+8fJsOXV
sGiWf59pMDEjImZLQEq5Rc0M/uECWGKuOP3Epkp7tsuSLdicwnKbo8QZVCWfeDIg0/cIsRtTIC0v
iWD+wWYdRbKq25R43ZKZ9MvynRTxCWvjanZxDkTEprig7joKOI72e/P3cDAJnxNFHjNO2JJBhL+5
F8NnOe4xFTCqaT3f4xKHb/JP+/TjfJoQwlc6n2J2OLh/Q3EBY26rQDFNzwxH+MH+OOqHOV5KtWh/
PxXP8dC9UtnugX5USxNxSH3Ur3xVWTxK270advanR5dRylpib+JtjtfbiWQmxs27sD6uq+7eiO9/
NNJaYUaHTxc8dwINjCuS0mIR7658UPDir5uaw5O+F2J1P+cuko9tLkzxRdRAunJkHSvCtMQ2EqKc
yJAEgYLfgDV0r6BCywhysvQ8PyxHpwy9AwzXSUhxynz048nqOkQZSGpTtPm0K4c2eZ2RqIRLCcmd
Qa56PUxPV2gCp+elOnEo9tFYrTH6NFCxi7r72/0xuWi4HuCyuwTEP+0rZ8wnfDdTDrdG9dxK27Aa
8DlT2Jhsn9Cnp0utC4/1I85jP0wGT7hx7JC+WnMXAvQGILkVZhPzAm9/u/BSjkPN6Tx+d1/CDa6F
SqJpISFB6QNBqf8hvqKaCLgolIwExCUUF7j1XxtuR72iDcKEthv6JDjhoaCI6AwOUw7exJOlVoCs
Sq2De60xmN2RJxBzgkBLDRp/wDskS7CaXgc4ExFRup62oX6rG92hyrPv6uMbTjOX9nPX2BJblgGN
B0ItT652akIG1HyeQhmARmuH+iohZVmntlaMyHe4NPO+oJL4AIObPnrwkCCbL4CWpWVKz+jm9HFC
MQUlprH6Q3tXrbwTiXHN7D9HciiDTZp+EmyBZn41Sp326j7pRnUrPsxK/n+WMQ1fTXwopf9t+/uf
zGsFFgsRZioMCDSam/rkAgDvafx1YoUOjjdn3sjSClQhyzVNTybdh2cUrUizISiNgUUz4O4c7ikl
LX35ugf3xYpTB0hHlUWw2XBjn3i1MUT0xz+BjOanJS12SSXDJzp0yC54pEnojS/EvhRomQjEjdYt
VoLkm51eR645wqv4iX/TOA0gZ6/7Ln/cVeKSOIzj9AlhgCmzci5Zgytrhd4f8lUPjcHot07y+YSJ
4duGkAi2ytYIj4lNg4wRVMzmmiSAfKkothTZV0QaSVUsclgg2sQWXVez5PGNd5WWGPW65JXq8HI9
YyxPPfGOJ79IibuAlc+9RlBT+hF5rynb/m4j1zZMMeze2NlDR0RlGXmn8WCOU+6KKCc3t5UDrcUy
Qdb7gcu11krViMk2v0KwRYqCPDSuMFO+hJm/CcNpREngwUgj7VSwNYTzjQDepqQrj2BJzX9hclKA
6f25YiyiKmvFXRoBO9OoVEX3GbJYT1TtYni69uShdp6P4BDGR8HyKkp4pqF1IA+W+tqqXbqRvRz6
XEJoQ+CucoQJvrivvz/Vr6tTcmSf3JDI5TWQnQjx/dPdBuOjLu6jDbt9z89gRl4piB74TC9k65yw
tMLQ609SDzyy6f+ME7p1pdjO6gpgblkP3kVIG2P0GDYkXgHMVHPuGZwnaGKLEpgRW32RnjSsFCSB
1yWKWdki2wSxWCKWBbEU8Ff8HYSvId7Bh5tz6VmzvMiCU/Jg8OtJ0PclAtIbSv262yUGYaFjnv93
gH3mWy8pGGUgMQ/y2jmreYO+dhe5aZOkArzgf3s3hBM+3XSav88/o2663zI5M5hGVluSJv5lXXf3
CsSNbJpBOybLt2ePxpVUhgQuYFF8RO+iGZTrm9iVLkMEMl1Ka0ZEhGw/xi9ibqeaZaZXx77Mt46s
OCTI1rsCb9cvMRwKf72rcau+dQgPcXwqZ3ybfHROHnBBusjb0Tg9pt0kmryFygsUpZf/f7s9W+wL
hMgBy+f+FUrU8o27bDJQp+p6ghlLoKAs9ZWtr1WdGgBpcnkSpdgxkfi6Wm+fn0k1qcDKer8FRpRX
VTA3T//A2B2TJ4CwVnCxNoHty8njBowz7i3lWKN+fEURwy9dQ9PAt6R2KE5X2yT52xl/IqFUkUDU
xVfw+b3J2GnkS0XBALtMz55GwcqWS9kI8ssdhvlpA9/h+tYtAhJeoRY3noAvxHDKkLcICRgJvt/v
4aozRNNq0vJ9mHmy2ka6HHnBQupVDzn+hMWbJz1iOP0M7lE0HRY9eHV2fFne4jlbjA3PmufqADNM
jLaOv/3anKEeQN2V3zm+1+tO31TZOSCtfaG1lDOD92w02OXSr6VVfJhlagdpZWjNoGAjhmxEOgFc
ZK1h5c7rjfrqrbZMBkgZgDim9+yETJfPQuTQwEVBoKHguvQ3Fka9Bc8doG5YO8KnyhR7r/yQalOX
+KQIi+fuTC8GklSK4gwkIqxVvFZgQcy2fSlCoZoMSw5q/JRCrMhVCY2CMJvCJS02M1HhKLxkUP5s
rmC6aYveLQqmDBHfrhF0VcLIa/GJH9CxJLXkwWvYKlrtci5FghnDyCvqskoZbenib0yeuf66yYCU
f0XBThLSy3o03UEQ0MudEWhlsumnxswpRluh5jSyCkHRzO42O3TaEFMpS3CXR/t2OVc1Xx+d7II2
icKTDTTFdLc9H7/dJ2KSfZN+smqRBdlbEpx4VdIV97LUWdbCPJCjOcvqQuVDmAL7sBmUdSVysvHa
/HBT1pY1TE8kLeEAspXkTWrrv4NIgNlwUD+woVMvplcA3ATcKDZzC4qGJ77wtW2gSiTs61r7iXMQ
0amxqjhAnlwRvS81E/edZJ9y9CSLwIzq/lLcelotB1gY6Hd0c4PfSp6w58Swd+9XbuMDzAeZ08U5
ESA1PB+n2lm4P9BLZW6IWjZSeWhn3yZU6LJC/dwJsNd60qPyqTh+Yp/aGewzK4QxyBKB7J8AQFwj
i1TsHsKrCxljN7VhzmtVeWnBD3oZIsqok5DL2EJyqd4CPulhDNnt07OL0j2vs3oV/xEVZc3B+ZgJ
SxCsTNXRE4uheJZ3zHDb6JwF+bWb2zvfq8yOabXJHurJksonX/df9XhB8b4SbTRf2qzXTBGg/YTN
YLDq37Ij0tAiuiPEB4dniNcLZXeqPpButoVPIuExoeBMUMPQQrZB+bafmnByksaMOLlz7YtSM/j0
p1OugN23mLGExKAA9flANwegdEs9r6wLXzGrKr/MWsUOHSJRt+740TcqSUpDwyGFVuoHcy35NCzw
1elMpO7p4KK7vJFn+5T/WOPQafrHcsT+C7JL9aqfmPo00P/AHG92+KezggIfU2/X6sz96fT28B/z
sijt7yxVdmA0InEEieBQb9rL8bEE6VWpeYfO+YHD8EikAbAyRi+GfRVP08s/i4JUmBfngaWBHEul
cJfgBWCsfNplkoT3o+/aLZ1avmzFjv0bAvhYLGmaUrzQr89GjrDvp9kFCvZUDPvkjPqhUYsUpgYc
540hydxStpc8tG33Vum9umLDAvrY5E7lQReza4TWyJNwl72MAhx2Ca7sXjguu2wnkjxytAD13lg+
pCDL6MIIg2TWElAEtM4oIU1jQyUgEb8G4eIrY2WdBsHvaGlFE4i0OAiF/eZahYbiVn1Y3XAzeSoJ
n6k+Q5mE7qB3jVkMdMSlSIQZh1UgFAaSgGn3BXviryCUaVkRha126Z51R9yPiBI4+/4PgyEucaTx
0xud1kwc5gSLVx/ICxJ6vte/BZRm5lkMohhz+ePRnTeQAeqOQG4dCAlyeaRYMbSLWp9K5jTzu9nq
r90PfR9xZeAhJi2LzAJGqjUldkOuR8Uh18bXZgyrhxMbG5ut3bYFMDENtKNp2gMI34ac9Ts6XJ2v
KzbWBim7AQH1FEUX9GgzfOlx7qy6eFE4vpCPvxp+80rj1uSI643vpiOHih1H7WqGI5WnxMayFxI0
9fOxnwBt7YOVPwB5uX0KH5StQBweb3wAk8ByrHVcO/7YtFv4QclJ6Sk6Rmejy2wlL75BoRh5sXEp
azxaJikYYfilUKyilWlpT18ctYgvl/6XPJbhQKnZCfxVh3YqImVLFyAgF5F/5/4t3TE2+1AJuc30
5xz7GsRBEJYeTNUeMV9mVlslz7+IlxI85FWjlt9ZumaCUNZyp4ZmlI0BVwPtVZWq92mVMpk0SnVh
CCAXyH/R/1gur0k0nda/Te0Bj7JYuagBxtiXhR/1+Y3LfMMPhm/qQX5vQGHHSzxMJYFb0dd1neo0
+WvxlrgDCxayr8r98HvbPh0m8FvdP23khDV66SSYf1c4veHB/5TteX6HqhwgUtsSdTI/a7uaasIy
rSn1tOOZlecgJ26DwmZgflOKn1EsyNZQ9tE7PWnX3bEgN7UVRLt2ZK9jhgJydWYIzorHXM4hwclA
1fKXG1j1DEpyyT5yJOZR1kgH4EbwgVisPItMIxJcGaPMoCu/oBw6CAf/jA4s28rxLm5K8BKkNKn2
7TFv9GPVolxoH+wiCVarmYPbY+HY9hgflQYBtN8n+V5dR0OT/0JrObP71wQVnTA10u3xfDFn7S7J
3wRs44F4aqASs+cO1QFAhsrIsosa32KxQ8McJVY28gWXycSXy+wqDh39nADB91WJh/ohyMo03y9M
Fzs9ncHComiUHrmMZuuYz0ApZf4MBdOCT806Aqhl/mEjU556F/MmsGf75KfaTb99tkoabeP5mOrA
31/HUS3nhLbbbLyWHFnFhf39K8HEj1LkHqJ5LSj9LGh/9i5NCHvtRL3CE61wHLWXfsF7U/uuhxTi
pEQgCh+uDrqpUDisoHgkor1ddJA/DvMm/jcs7kQFM//3/pL2bJ3g0EGGHPCMU+KJRJtKOZVK9PMa
8Jh6hwhCNyIf52IWPdzbNV8sAaZIhRT6r+wm8iY5eae/6bfjhf9LkyNC5mHQAhm0okS9/OnDEHoK
AbRwltQtYJ6ZTouoPjJTk1KNzv2NAWxCjeJdLq1hH6udwhWZhYBYfoW/j1XzwzREnRZvZxW1iQZk
oqbPQ9knspf3ApffudRUz0HsY9PAYITEMox49MTRokIDoFy7sue+Z9gGZ4md50bYB05hRMJUq6+c
/X1zc8sXzwlCTiTSkA2qTIkl7PbWaH/y8kTniL5ij6b/ZMXIdomGReQET/wE2IUH7e+IKRFpmcsA
4oSFxWHfR+pJAYkHkYZhCcJGYsJvew1lRApKPm145XY9NZKlH2ro/TVQgWNC9hAVZwMPCGIlqqKW
8gpJ4MSHUPIbk63Io/9aLY1pW6V5xN6pZ/qY2yn1OTA+YgAJ1Bvuem1mj3up1dqok7idK7XWwsU5
BCXY70wVV03cArk6S7aVzjxOSEOpTPyGtImtW7Qiu5CViAEWYGf/98PWv/uNIMDVCLUIwACXiXrg
g5P+iiJmhYKknD3sZkVaCWbcU2MceNgDb8g7rDUpvgFMfnUf/aWUmwOkkHdJuc3T9SThLMleTJnL
nM+zWt3SAu6dTNBYyfUHNWi8pVEVvlkRgnnPireLNDcTMw1k2+9xv3T/Bz2etBX1pb5m4iZfudZI
07W/k4VzXPSiRRyGodonJmsBY1R/FcXNnMRGjtYLgwWORmq8AuzesEZuIUA7fT+PrGSCCbZwT7ZE
zSQguDcQsUiKIPv/h8zbdvYLOPMnfnwSBl1dah0xzg8rovgHNv0T7XPcAyIBMb6YpdHhJaah38n5
GT/6vJ5VS99olOXy/iAX7jt5zS65CIJx1FSPRzo5PAbs+i8b2X7TJSU2okdV5rXE1x1K1KBxnqWC
MF/zWOWDaV0/+E0A3smxUQySyHuOy3qrP6pac6Ttb3ejmKsJXvvTE6KP+VBA0DkdQF7CQgslCv4w
JjB1wV7XTnxG+mBtIMweXvrnUE2N/FlbLq1iS13LGzERtbTkepLm6+TnFAAnUERQJx/7dMv1BHpT
0dQkO9J7SU/j+QnWGBUf3XvKCSHhUogeKBapul1NWSJfzNiydCq3gJyhYgVEqAZi56151/DMATI9
6dbXvDXMtEg+VYjFwReEorvHq8f6jOq+bepPIeLTB9GIX3p4icMy6gnsk7ovzfG1QiyXfj8kq/Jr
JXfp7LV84IutKNVpd+658g7nrruZMVgwOMv+eQjVG1ojGx8hIvb743VyXX1lm3B9t5o4Fi+82s4i
u8H9kGYF83C/bYrWZJolpRNFZ8HPPBFKowtg2zU179x67OH7tetHQdr4N1oX9QqMj+Ixk2cdJ88L
W1BtEkmew2XiLmM/LXlZyfLEI9JIGMLCpgSl6aX6MUHlc1wXgQ0VkspLTy9/j6FXUBhd3KqyQPYA
imMt6gU0etxAfxCvTByiE7ek2893uOZMOECdMLgkhspd2EJMcg4psB0Gp/7rD+ZmVOb9B2yoXImx
k/wZoExWziAuFdVxWYoV+a+koKstT7/uEx5B4oqs7ws9On9Cj4ZVfIbY+J7wZjaosGeIbtJrxXgU
9VCW7ze01rJdrDI90qc05lvdlRvfJq0bGCtJWph7w07VjhwSjrQfHZ43PFARZQorH5dAeK/KsYuR
XRj9BD7vcVsfqoZcE1rObYx+ivA9//ep22Tpby43yw0HT/EbfUBHgUKeEIMopoeStg+XMo8jUDIL
vAKCakrmT6IF2Q8blwm9C5TgqQwKgu7coE6ngL7Be0hqRsDCwELH9xkJic5AkTzTU4EEEgOyKk+h
uAA5gqTNXirMe+gu9rbtWLAT+98MWSQitvu+sbiM5MfGnlrqi80PB7aLby+AlA/Tejgwe7sTcMMZ
xwIWhT1IzLlJbsgLbmiCRwCfmf4Un2gZcPpqtfsU8PPpJREfGUlRoYnExCsKU2O/tbZYndA/w0Ya
r9fK8OjgsFU1ms/4QGIjKo8dNgnwUUX8F0/0jkpNT0aZPPJ3HKp7uEPoOAkBDmBDGTR7XBF/c5cg
NHYRk0HTU7ocGopcF0s3cF+/y1ANUmdxP81PXaakjSHFtioHgm4lD8FfOwPOt087ZaJWPt6+Jy48
kQ6p2UeIGPMoP+azfJzHuhnBXgyt/Dob4y0e4XFXtpxycPVAabnVjN3TRZx/KVxC755s9VqnT784
0IDmFDGdUdyti0IbNwvoW4P2SO5DWr7/6kN7D9mVz4mykNRr9T4rKkAC8eMPrOC/KkRY8/d24REU
v7UMw+gwAtyWlnYSdHJzifv53QUwN+8s+LvoLxVubmuAkYZKTuzPAUcLr+auCcbh4Gh/pRMdZCJg
XV9i6JjlLn/DDprAJ2MeLumHQfhHYkj3iZkLsAfqC5ZLJo74lvSMa8Wiz4Jjqii39RpHoD8o2v9g
CaPpjAVb9BljrlO2oQBsFyBbkfMlKw2jftWK2IY45uZpH8ggTDu7WRMsIjVqhbmqX00GmHEXmWVS
KrvsG955GEWKonPPp7CcmV5N2u4GJ4T9KziPjtspgQMqj56vcXD8E+IvumgWsrScrFWboBeLd5xw
PyxmMhITYsH1zeeYYmZJojRoEaby7WDTfdU/Lr2m5RlZKhaZJp211FtFmtkhXhxUpuvkrRJqdN+M
eUGDRLS+REQsIo4vvwgeJxp3I5xi/GMIh1qEoj6L2xEpzIkGO32jRpZEWTSRMMnmEc9StmHdetid
LiF+0ELcE9kfxp5OFptIDZrRKKiuFqJeR9MMFMUNgSRCKUpaTD8egJwcgeKsl+GxiiCrNsFpbvEx
bNc51aINd3jO6nzTcnTQHU9gbkH5TLlxrLXjhI+vFHzmtNmdjvOyx3BpImRVT7AH5RuiYTnOECki
muIlpO+YDwb2IUCUkDonAy1bTVjESFv1Y/p8d+xkh2dju2j7a5pFVC/Tu6nfMNAhSNqoxjhrVFXo
ckBEF6Qa32vbhrRiXAcj4/FlOk8E74JDStj6JTach7OQphhQpIc3GMkmG9npXXv/JbBBbrpuAl8e
sJq450xYv1tPdc5bSsbaCsCTFnYulBAFn0xp6JdEKkb0WwybQudz+ELjopUQKLtaT/EfpFCOmdeJ
eqASdUzzLtRH0MaA3HevRJlgHltMoIhKdlpvn1G4+Nza9HYMwhugkIssceugvjysaHgvvOOxjUnR
xH4OuB8gcuKlJSLnaTqOb3D92EQb0HRRp5vjxGaLTgSqUjBcT5CiNC04vDvzyLo+EpJI+ejeR2ss
wc2+CI16pOBlcRpRNrCHloTohMQYokb0PUqpR3TJnXn2pyYAiSThsrTbVx67DQyplaLyylx7XA1a
S1J2xgmiWZ45OtFHnD7AUdqy9nMTppjjdEGnev0sH7Nu9lfLgMD5UUdEAdFwEuLZKh/Nz3IX8Ex5
fdQHntEwcMcvGQEdm+xNjB7j3DmokJyYqqCOg2Gi4qvSQ0/yUKrv9OF4twkL1wbD3NO1SN+lSvff
eWBlPrtgJ3rgGrKhPKvbkl4hRCmTzp8Y8wcfAZbQYc2hVQ1pAtp78pHHD9NVFYrgdaJh2U451e+C
WutoR2SjeYE6PBvf9109yYo7PtC+P10msM0Ne3yHVg+jomwswxgrW17xvZIL1zlfYGkiJD14CWp3
BdD5ODgr2s+YcvVFpGMUwudVimNlvjc7emKxIAoWJBsPOwIaE+QEW86m7hYhOJw5TVFTbuoMepJd
mltDVbOKaCb0vhQ5JGxLIkM93iS4yhgua2CDTJsZzqRJKtGwPUE6rEiizc/9Iojw62xvXYETzOM+
3oIDXsL4WixDiexmh6MeTaQgTb7olXEfasqmzyYXiw9gC/ymGZtqU1SWukz5o+7uELJPh2XLKyfc
hNjpZaX3dDTsBBKbhMwWIFX7DA7+rEXB4qrQg1DVZzHfhB4xgsc7I6PZR3NE6lB9/rAXHgSzIBuZ
ysj/Y2YAhRKp/qTj4OA+xK6vPEHLO36xh+FMo8Df0fO7fmrEAMZuZZcDz55NjSCYbGCOit+qrzJs
A4tUWKBIxrkia+KrUz9Iovi6v3AfbR+GUpToa3skvEEMNf8KKgP0sugywILrIUUUR4ZHgmEJXr98
SGEehAsiICEfPAAwIyfSD4ghJKZZLJfsByjG5N+KuS1HTTH5jQnWwUweKAK7Y1eqT8Micd9qqe0m
xNjiPmUahqrZ5SkfYHd5thWbdwyZyy66VfwhdSAf2YSXMX34Sxm16aYO1YgR0Y5LSHzj7VIIkHaw
v009mlx/FLLJIrGjPy7vWnRONvYsV7AvDe9yzfuVyVjKfcNUl59xO7lFTTdtE61+3ZHohtk0Qtnz
pXfJKLJg7gc1aOPrvOO/WJcmmYaQunZjL6v18dxuxwPSi8Oo2rTl37rS7CraHPSoLuTRSjwqe/Y8
S8klm2Gdu257peoTw+gM3ySsp99c6A+bVdz88rl0QIuiL4hfEIXCsp/PLcBpngYdkdPuxlbrgHTQ
2HVWfXPSqJ2uPAhAWNhoFGZn4lpMTbp5nRAPVjrkydHQ1JYU/Ew7A9jB2akgmQUEIO2K9X9QoP2b
GgzYU1Q6uBN0Iq3DiUZwdBRmTcbN+bkYUvrQy0MOwwXeiiyXN0y/3XJ2cHD/ag2UR6E8sriIKG3i
eyDI1gqd4tz7XUpNyKkZ7Pb3rEV16963Ml4odskCdEUshJKYd0hBVfgx7t4tTiLUEWSAtphbJJ5y
iOKwfrF2LEpqZdHlZFxl4zEw/44zFcurrOz5Rdim0zLP5PktEgL5PuTRNf+u+xsj3DRvKAUxmw2U
zSBLyEef//OLcvg/jiaRfgk3FHfFzc8NxrByFTfct7uFZhc9ukz7q37PVx4cCSyAuiRPMvdMz+Qe
sE69GDR0UJtk/MBq4zqShmKnVgEhRIUrxrE/wsYfqPFu9O3+6zHjFhleW0peFxP+NahvRzFKrS+m
jjmsdOpYw13A6xSY1gguFdaU6AXnB5vx8MF98RuZldfed6zQqR+PVPX+PvEohNC2YieDRMdp4GAV
xRD1JicbvoWYLBireb+ifdtPrIBVIX7uWsVNHDSlYcSHeClDYIQ+EznkRmvqNDZvNFLUOvMMWiFN
acHckt7gRGIZFANw4Y6bSDysJ3Fl7MebJU1ytaxop8Cg8woW6fkaQLbggyOPaDcGBSK59skac2wX
C6f99lmt6EuGF3Auid8JNo4IEMqYgHT4rqmSuEGfBG71i2HtGxyDFRVmkjIR4v6pIgFMWzcvrhLy
0K2puNDopKCZq1/xbVYGj+gDOZxO+m6fIY3P+zOeQvZS+L7LAF18Sc8tXBsXyY5m52RQtMMlYb63
wdAJ+vS86UABsV4TnXqZmYj7Adj5SpgPUObLYZxR+z1AMIfarP35FfZ1hZvA2AzDhQdqqPd9KAO/
hMNHNrH8was5vQoWJI1ZlD3OyQaFXdTn0TDfzhMS6CIluiXmEZTA7jh2JfiOBqt3m2TV2cSOhHak
tG5nkVczHDlMT8f4ZNhigq8jFh8ftMb9Cqm9yz977XGsRUnUVnfbgH0IVKYhzhxx9AVd5FUd6yFB
LXZb5I/DT5CkhGpY0c/c6daJwLKmM9JMUmgDZb32LPpFKqAzaLQ8Ilay5rZu5AjQJSsP9Zdm4Wyi
A8xvLhk8RjFeoq/STaJjE1dLRKz8db8zxJ7TId25Kib+HUKS+rhdlOnqgZCHPMZu4WZrt0ef5BtV
IK2WOufikj4aVdoE7pmdl35GTbCyCH+ggdAHY9TUzRzUiUxt8brTLMm2N+Y3IdV3ZRg0RzY90LoN
cu7mKg78ZgU6pWvVP6md05/TtX5h6rr3lzGZyv1beDNCwn0ucono7kHWUnBEA+VrSPFELcTj4UIp
/EauPqcguTwRw8A5VMlp3JsHTLTVYUiNXExhvA0nR5CBtet9VNQXedY699TuJEp7MMs/WIaaXXn1
tAurPj7QlAjtA9N0vlapicXIm/hozbX8+C35GTJ551pQAA4Q5vpO5chm5wbLza/rXWyPiT2QxpPC
LgoPgQmtFyXhypEcqO5q9CKpn5U/AemOb6rdegoML1RIUdsjkiEydT8mO0ta+fD74OMJn+8017fk
T/tDzTYKEpA4thaBDeHJXiRVYdD4YZIMmFNZ0kAECd9fxcpYusrE2Ang03gIw9sgWR55O8Imvy+1
MzLNbW2NqA8mJZjd+tbKi9xWLwF7HbeqSegGAbjWBYd14JrqZJxx6EL2FUcKmQ7cUMqFaj1Me5vp
EWwE7H2PfcZgaOT+ordGRLmfNwUEWt1UeqHfXQUrLLr1ZrsTbFShe1WCy89svhYAQwM0ikaGxAE9
1+r5VWdI8Sc50gzj96eRLk4Dd+vn4JSWZ8ot4zAwrBkevasgW9gKkDTXDsxEQB6gj/lRq1wWzLAh
Po/Uqaa2olbolE98z7rzEMv2sg2LnzMGmxhZA0GiaOu9jj815e2zqEcG841QsUWrnA3ZfdghF7b/
NrpGQcy7tcsRu5BmVxyh9Yd3UeV5T/wIEZ31aUAJBO6ENX9oAtTZLz5bwcdQYxQGEa4+88RUSaGe
3/BPVW7hn5BLjp8IZLgUtDvgUulAfQ8vwg7Wc2yMyP8odamXMqYzLDvNi9vCruT4NjifznzAoth9
iYvunZRcIgX2txHFO1cJARC8wT0Xm/U74n+WP5uG6zIbyi0fb1oAAtxElVBulqSppY9PWnxHI5wU
sZChOQnVlr7nJNI78D8lxT3PvJBTGDunAEYQ/9moB6ADxBoyN62wX8+w3nugNwOxe4/4iE++LZFB
xSPByEIQMpv62p5jfklj8YvjT6QfGNF9pAaP5Tk64pvYszGBZAi/dtmtmDWD3SazZI9uR6HvgEyF
pHZYM3hf/GX8y5LJncvIxtKB51+gDkvoFax+PVSuppucTtqwqjDRgdRuQTKxSw55bDeiRw9aOfW0
eNT0noI0f14KIb8Gv+bvnAF0eRGLzqr7gdp/FkwxIfrDvIooNdnNxVd/1OV/lzo8GuvWK7KoN+2i
fToXlL0NjHKYsdq1EKkfojX5zO6Kx2rpCQybj07IxA8GmuQ3VORDgP8ieSaYz4K+wIMJbtBvKFhf
oVggOUxDVy8R2TNhtliJ+vijatVVrksmHkaDkYxOVl0xV7E9ZR9RnhdrwpGGBh6Rhd7cAVgVvUiI
VHBlc4EGI8YdSJyXrtSvSKcVLpSOHek9ma9cmJVJyznEatZ/G90jR7Ys+ypmW3sYao/G+HHzf+U8
/iIC8jAgPms8CWkH8I83CKUWUjMERwiJG50JCsT3PEZ/W/e6VjDTzLDe88x+ornSWe7sQGRshWNX
wuGYDh2Q6hKSbQ/CX3BDba3goCjhQxkmDysfy0sSOODuM45JcYVPxagKuQvHMfb3DZShkDMv9rnj
PzG8QrgbQvASv425Tp4wtnG66CwCGK+OB9LYmOg7FBs+7RFfxv5OlbnrkIRA3aFA6bXNrjS4ohrt
uNYaP578WUK0DCAXDyLO/4nOtPcc8097KrfNk9bDVM54rsjUuQTNhublt8SnBf9CCLyboR6qSFe4
QNm9mIz5NzbvUxVdXWUqRf2IHlp5Vq3QFISAgwo7InpDN0XGFHsy14ULZ2CLJK3nAShxXIRhTKXv
wAknrt5JztjgHMX/X8DrnsU437C8RXni7kC3D+Hr/kBMyEWVo+DCfOvFSasKvYXt5K+VL/KWcurO
YQOSo/sGAQrOq0P0edSWtr+7ViQhogzwmKcQmquR3RZUpQzUWtyGif4m9j5UsCVgNW4IyZdb22sx
MQVoch7BFUPcU3kdLwf6wC6yRyr1GjpDanrNvA5TEHL+skzwWyVldSdQnIFyNmwOZK+WahvPoN2A
jVpvKG03aRR4bA5TVV0G3InokxMjyfDB+JVkLwltkVp8SStYEDqM98H+ScWqi/9LFMbow3dFNlDL
7Vlw5ouYvVHKfsz9si1vBFO4GIyl7+IQUz4NhIjFpMDZZm1gXc7dHSO8YoEE++kfrnOF4RhPSVbw
Q4wMcc2fBrx5Xr5U53cHbbwzBfKVHl++v0ztHEV0TkMbpKdd3gLqW3A0GlmhrdDSIM+cE/VJhmca
KgqqyJdHkDtg95Hq3afSBnVWec6KStvvpZbPfaGuNicjHv/4pNb1bL9WFvFrZWyZU07DUTlO95/B
h3ArAcMRs+uebsc0cGEDuYa3IwUhu/4eRKz+jRU5CKQ9Lb0S7LvyIKRxxrwWLeA5F2opjFHWj+jM
C7U+di/NkaX6x625Py3putQHFjAm4/j9mvPioVBrIO8JTBmsuHX6afku8LXkhP4Quc/OPwwueOxE
ipOdqMIBbi04RH1hKnHPOcMnS5YNXkLhsKBIHGRlWZjPs91PtBREVM3Pm7btCBeV/J3jiOE4nukr
iXCtKKonmafbR08W4Ox7mSal60YLnYvdNFgqzOST0sAfOWXIby1uk6UOBahbhVKqNvzfu4TbdyYV
y37fmF1pDsubVgC0hltCwY/C3Hp06kea79IxLJJwWSA2VPw5PYt1SMDvXbVl0eixNkukBaKnI8iE
Q1jjaIFAw/PUQDq1f8Khtbylwz2TagVfM00bR8H3owVwRVQtc1N+EIp3cl+OqeRkRXfRnbZIMgj1
+UjZN8hRsCkkRKqoGdOmpFXv2opUMc4q4YOzEnW4uyBHbihF9QmO9MW8cVB+w9Yez4S6BKnpCeJQ
LnN1VqlWhYb+sgVzhNyw/EXNHKPivwEuLEBfoOcYi2LIsWQMm+yT7z+f7+WBrPoUuThd0kPTngMp
P96VRkAMW0ScTYBhfPqd3CbUU3Xg8fYs+qegPU813P2ztEkjVOlfmPjNlSu1QcrQZL101PG4ZMb4
XL9qdt6gCK+x9giUaYbJYSicBuDL+mJDMqil+bhqSnXbj6cu0e4Cg8hdxpU54deTk9Z3GpVbvSV7
Bf8HyOobXACZy9Kh8XjednyzLs8XwPCOGqqHdgiSrpSb6N4agthTiiaFl2+0bKl7eMNrvQ7QWjui
vZ4Fk0ybQi1WW5L3zVD+60j62Z2lJ4exh+WfL2u8JOGyViiMIV5LIzZvdh8LP+aJsQ7YOYbULeyr
Yd4hJICH0c8O7hJ2VjVK63pYQquJkP//v/+BHkqUeujA7c2V+leqv5jzwKeW2yVlEgdocvaOPb6Y
wLAJwYTlkka/O8FnnXenPFdhJH93qsIiid2GzSlxRQAlyT3rU/I/oBrEcL/+J5aRiwYauoMQxZi1
YrMHhg2Py1UJtLfiWX7427mumgvoFri56y0ARsKFp9k12KuBtcZZSzhgS735zmw0ERUO4nJA5LEq
FmWOdR6MpIwCkY9gt6EcZNlW2zBWk+/Wroyj1R246XyfZcOJufOB/3dkn7gBUaMGJTMqz4Qcfknb
3XoNLgincoEyOFBADmFdIOCfYXgFrrn52yP+UDVLoU820VQP0A7LjmlHlOZpYkpRppIBZ7HY6k9w
wSfy25S1Fv111K0QsHTOyVWu8BzGAQ+nwzRp2m68uPwCxosFCAcy8ZFijD9F9rHp0lEMy7BTZ6m6
Z+aQk6ovluBTgSuRJq6j5SST0tLHs7EP5CFwxqAth5GcAjvavLabq+c8RI8RnBYQsaTM5crLE7wd
A8NDSSrJKl2f82bLQV/I8D+n+MYEOw2XZAnnT0fFmSNt3PlZfSexbyoY2bELdsh4rzad/YcbifCv
ES9QiYC0npZF8QgsMDxNmfxZ/Z+4tjNOszVpbPRHgX9qIiBPZY+HF2Q8b79n0KaHGiw/8P1O/kQs
7NJoxhcpG30mRiY5fEXN4rdd63w4uaCqxm/1h3hzu+kt5Yn/F/iR5o3GK29Mh8sHuCZbuf4ZR5FA
b8kD/qHWevoRCRw05K8wEdvbJSHKi/U4k5l2uB/JdmMm9BygAJn8GHU6AsfH9cKucX1g/4evvP+8
HGXI+UlU7aJVItUyJWrbwCNPTPBwoyMGGO3emD7sZqLvzvI8fEcG3qzNz+X23mhcAhX8ooM2sVGw
PuQJ2kcuy2PJMVi4c0UJQCct5G5/ZxdCV/u1h41cGZrx6wIZ9C6ctJLoP6CAJ5w9RrGejwJb2go+
iL+6P9jFeqnG8vmOEOqiu8umA3/RtYyoA0qvnTUAP801tBoDpc6JYkNb7KdjYKFYzr0XzsMxzNGQ
ZRrG55qbeCNa+BEU9sSQ8bk+maTii7kTKX5ppDZ+pLN4d+baDR85D+Ejnmffg8ycM/ch9RP0lCJ6
pQuzhq9bYU/d/MUPITJQ0wnnhRNvHDt81AUDq3xXBXWtd9RBJXGlJbVnA6hqCUP92yulQOBF6fNE
HkB+zAK+jNp9IlLZSYK8VwOk3VHdBx4f+8whPBiS7+eZbWEjqqLEzC1/scpg7KA3KEjf60wxpVTr
h4D6m46+SU5iovDcAKdyzmTVkDraL7gWv+KUWS4QaK0aIlzU4u1a0o8dpNRLzTu2OWPh8Cy4RXtm
EQqHQI9dKixVp/twI8/YRp+zpiboUFPnAxZVGCxIJM+Rnz6/IdbDwbiI/yQrUCiskmGWDiyOIkqf
2pEH+vrH+wP3fuzEcjgJdimo3QmerCcoT1WSskgVpsE9NICFyKNpR5QSPFvVIr/556kt9hoLOWCt
MEaeVYO/aijdt5lMH36odsB7MkvULExnbriNVwf9yDW6A91OPS0sN6NANlcvsyf6SdAS7+m8PisS
oS9XybjwgaPiyfZN2OAKcsQ/0AGgXqrt9p2o9B2alvAwf1HrBmbEu7nlFVlxe9SZHQ/zaSloJ9yb
6Nlj7uaIC09D3fGIt2SlqqZ95TLdt0IPBs1usDo43ue7O9ImU2p0ful2UB79BjDHh8f2NfhBT/fl
LYErKU3b4ENUX+SOvQEz52I5XAAK1MALWCJUiCurDB3LPOR/+A42K8Hxv03HUNhoxHuUKjnCdzZL
uBgEYGPKQeBTVKOH64J6BVriJtqngGhxH0rYcBlrK9VgBUmYSSn94JOyKj4kuYtsn67IUJjoJRF/
AMliuWwUqaD3H3p9wggZ9ln/pv+uv9GAOQufg/heSnh6zomjOKAHskw0uPFTol6gewbbOknoCflo
IgaeS81bmo2Sfxrn1IRVNxAgIlSphFoaE61PCu0iY6dygV3Qc39mFoT1ofkLXuSn3i44cVnbkkN2
YnObdLW08wW3odQtr6BV6hpG6Be+jSQ/TFsecK4m2cbWp+fiHF07CgUmdnxASzkg7V9hPk9vjuju
A9u3PAb4jKFzSihP4Z0/mN0BZOC9Kp7vH8QKhV16tkZAG208LbWDZNIcCulQ7uRALDGQnsqjvNxj
cfmFz4MQN1NcTNd2luQxQcPZ1lMw/X9QtCsG94mkI/91wMcRocYZ13Zpt6fDIcy3q5KdNIv1RLEH
ApyGbi1FWiH2Uwb4T39LhjGFpi+Nm7ZV70q7HyljuL/xWqZLGoY2/iowEimbkoclutO465HGc3Xg
Cl2/EmtHXeT4eUxEUpTfLmt5YyXn3ImG5SdyKjULgmzkOCcVaGG08Rw5N+26CuGuymyFIaA9PL2E
5XIlOLnrmfiTav+ks2/ACXscfWziccCSHbL1G8O8nbJRNANiw0uOMBcU6BH66r1hsyB0IOoH5fbC
Op6XzZuZmzFMtoqyUay2KJwaN4rpfhEeoJ6Wxx/MZpVokD6OWTM/4o6yVpl2TDyAmotpKQGkx5j6
j9o9nxR9rTs4v/yE/ce/KKwvSxrAmNVG78LB5i8R4h87WySzE/vAFOHEsqfXYzzeRZa23erTi+qO
NL1TE7WSALNrhQZ7PaErjFCAsmPNBkWEMmEnWqtD497Gf2TRejMqAP8EtmUpRDInlNK169MHcjWM
5gM/on877GV+zLpoiV5z5vdSV/JpYDPtbyCJ1FCmd2dwmUakNx1XyWjyrXLeAZFStvXrovcJUvxB
mDI7DiywNisUIyy6Ps92XhVZ6lCmYO6QR7Yj8uH8RiyAPX4/kL3X2ViDiYIiW5BrydHlh9IjeZj/
wm8Z+1gVsBLrfjDHFkL+mMRhP9I2OHiv+BAbtdpKdomqIoTN4b2Xk5znKwysru6qwBqqoc/PnT6G
rbKB/wL0WJ4V+bqrPI0oA03iYnPSpggEfYCWYvrNf4/4ckvOBH/ZVb9WsY8YDBCg+p4ksIA7E8Dx
82l9aMH5dYEqwYOaBlZzL8nBjJgnQCdoKg7QmoL+zO7fkZD1rer5B4YLrELUwLy1/3XnseIP2y+8
x6HVUix/ksLs9QqBBd83zcwxvgbp/ZotoWyyR7kuc+4vt8xrWLsl30fNLMWCxIZqoT/FnSEjCy2N
nAabgm4MGz2wD/LcNmC4OTWHOFcr3Z+FfA7/I/OjJu2MStlbY1OgVsogm+Z7BCJQPxPcHQEmUHjw
KkemF6hIJDklBVSizsDObQvsA4UFnw/5QSBSkzc9cA8XAyAMQWDRnbzNmb6GlMOcHbQZz+ytLMnx
gkpIi2O0WHgo5HerNMBIqIqKVk6ppcarif/C99GAJrKAKiTlQrFWKUE5s7D9HvU/NtsI48nFVgNh
4P3UdvBlDG6PTdTpCldrTX7MzUDTVi/duVUjTJ6p0M4tgK0+plYnX2jhVlvolLTm/mq+CT3zaRYm
1ylHII5vyoUDTLq0rl4EaGbtcpT1dXQTOFpEXqatX+qTKtFlHWHSakM5UYAATniUIimMj42Vd5Ml
jczMOCOOfRsA8uYpkg8Nh2VthA2ssbVyJDumbpm2hJgnXPzF3MSlP/83/ssi3WvGUGAqHyrQvKJ3
8izt/9BalOmjuO4daVuC9zIhB5KjjLIuESAJrdQKpONkrlRk8EBjIOzPF1xRnOoSchIvKf4PAdUE
zVR6V5L20f/kcsao9UOzV3FdFF00ZWQchMGz3bBUM4kh8KlaFmzvpDRHzf+iQO8sTd7+14/NIjEX
l72bIm2DoMd7wCy4AbpON3D7tQPV0AKuF0RF7tw8wo88gQh2j1PJKZwdzjdDaNxAsv7hOxIl1KuB
vxIprTfsPiK857LB6eoVpKW+O63K1h1kEUorOZRMAkwHXHSxuPw9VMd5dXu89BclNgmVI0WBralR
b+TT2E60f+suVpgA8+6/yxZvmN2okPLfhCePg8dGvj5esxjqUjSt8hMj5pGe+bMcM932dcUGEoXL
huIZMu0rtwYIQ3V75zn6AUYMwudXfQXzVTdWdGmIK0Buus2As77VO137jxDY92M2S1NeQkwmNpBH
jVNKSfVfSVd9U9klJetvcco6q0a+QtJdLfTiSt6i1BzniKQ66nsvi/xsqf7WY3vkze0IfeXqAUX0
NFjq0qed59YkRXPFfiEG5gI6d6SALGpvZTws2fbFulHeH4xA3duve/Pzn+KuPBJA7QJFnbUUeVVe
Ii0b5CMuKkUlGfn9izn8qcucNzVA71OMRJEbUlQhg1Rm0BoMMIFjlW1kHJlonvH8RoTSdzgnC3vD
AWkeZskOYQpNDtFUIlbyfwHBNloNPzJkcN+GTURbekrKKcxBLPl1WozWNzKtpM/6bf6+W96FTwih
XoBqc/Awg+kj1zD1Pt3TiGn+g7aW+M9X+7mbWvq8ZNXc7pfGOdyOpXZ5mRcZ2xw5W4uCZ3S46r7y
R+kzUU1ImvGK5R7LajQlXR9z2qxyymx0oMIX8y6Nswh/8NLHqhLImNjuWbQD4JFlUeBNQ0F+tPdd
pBms+vuxMsfuiyC5fDi2YTfknxf94sIxipL+19moqJFaXcHxQZfY6VkdjlPZi0bxlifyVN4VTPbg
OO2wX5KCrbmNjhhyQn7u0/2mKa7nHLXWnb2sSoTWb3cuvK5KzE78tq48tbEJcsB/owlA+7g7YHOD
86hJ+rZcmxQsZtpQCTJL6I4Ei2HlCH6Hn+drM2aNrRNX6DBDZGhLoohFtFNRPQs5M/Kk+FWZFcBg
xvXRsQNSCN1T269XV9zAegrlTMY87pO1Uw0cQ17WdYrQEmmisEIJVhKnNdv/EcyLwpLgbVyvYetZ
1YegxMsrmMg3ZTkoB5fTmLaOXTfFGij1z/MoZ8hHTSA5cOrMpRPDK60eZji6QZcQx3/IsmhaVyvY
P9InCLQIO12zln0vIT3ZaUBQeC1Hq8hjqkX1+fNyciaR19IJvQyEumC+QxHF83s6O94vUGE9EQXc
eiLg+Kl2fJQ/Yc3zcB3090zq+L/zaW2UcxToVZFJbkDeEfmAzIIy0x7Ay4LMLReyg3fHICDIagL6
MAjeJ2h8wHqyX1grijCImjwByoeDbZrp2OnIqwm+0uqn2CEcRS7EJwasyMoqgf2ix30EKcn8WGwI
LJf8rAMudmsK6ZqzKsPIDAVzOucpT3y2BrP+uZ4q9a2r8HQKImPLyTTb99WGZYczUjpyG7pnGFUs
m7fIZeE06ihdh4kABOHgCui4pYm4ewD40DAbAW+BpDEOGV/S+kMJx1fl9HYvcPzFtylz7z4GNYS/
ADFscs8wg+g7Hrz0MvroBqaUSXUss2MVzEUd0jvst/t2rmWaCg6/hRtY+gqEYIH4gLmiDbDuCMTM
+5anUxwGnoOcBmfBgIaGgt512p3NLExmuYk+qjr44zrODabG26W4O4swfJCINVAm+2fCSv4atJ89
EYoBjKAFg7wp35Ft+gL1z+/5uKnwJlQdRiPYrAlXUqTdWmZvlVy1WdOwznTVQBDA5Hxuys5tAAC5
tR6tjaY7KOIt8IGoPB6Dl/dDm/LxcaUrsLBCZThprgyt/a+GwWlxBWl8RbOu4zmZgiKj76oN9pZS
kpcLAnBmusZuRdYtr7XR4SWP1G93Exdt5sL5G+HJci4cjRXjzmHSLF/JGH5nSm+6AD2PVyYwmMJF
W5enbqUWz6a4xtTPbdXtream8VBSFjruRaWSNci+lVLT9EWzXAErdtLRX7U8m6pTvPlm7V2uoeST
5UWqkEWGYLR9VzId41mJJLOcrJY37ZXrb6cIGrqaxTB3Ym/0UiWNXdI4SnKL3siqmlYQ+CKBbT7R
QzPO9mAX6ZNqwOV4KDNrtzbFtmJ3MeQdFXfybNM70D0Sv9tPJ84Xdgcg2E5W+/b9aCK6CP/+lutq
LW22I8XtU9TO8/2kpsoNBNA8NuTCLdHPWpKssA+mBb5AoMMLYQCgog9404i2OVUDvkra+m0521Ur
YmUp+cRx8mShWu3XduAtMv389win5mttyRnzpRLEikzRhqLctCh9TwI2dZA8fX2grGnjf0yAXG4m
2q1AMrNODE6w6qNE7oBJbc7eGe5AkSyvZ4W0U1CUwBcsMN3kBbV8Y7Pk2vhIXupgaeZTfaOH/TU/
Kk9hFWfRw8nf6f4lSjytV7B6c1dfFVDQB9pdSi5aVb7nkrAXzC0PXpAzSpFAjtUVndY9aUkxEmEq
9YS2vRQISmTsVX4WCIh4O90yNq0814wHKlvkfsKH1eYcXdUb/SWmEpdG4rTJ7F+3H+bRGQLGFkw5
GEEn3LgjB1sTCTkl7JxXkSmAQKmVBEHzPcxvhyDaKXOYsM6DbpcJuhBGmvguGVmeMhP2D8N7/u0L
4OkCRoTEXMT5lt0rgDlHqz75ENdDbTnzJAbjEtSwGjMJYXAH+Pajz+YgN6Za1K1LjhwtP8X5NmDM
fjFBImrd6cltD5CwG2s6ttvYASN1PBIUtMle/047dl/jbdH3J7Nk842l4PWDNSUtabdGEclJLWC+
o2X0HS9ODbDzwIQ+RfPSm0Rt31L3+pXu2SAv0RA8kq1MYuE3m/WVtZPPKxhmLqWS8pmZuTdx/ht5
3EmFGuJo5BUuausz02Ps7uzktrnFDKdVCVtSo7rR1xexkWOnCmP1/MNz9qxYpLAhhW37w5HJ6krc
CCyODC3KvTdnAskPlB6CTiO4EaIWqBHwz8y08vfDJXUJuVIr2++AtsdschM2F58g0/Xk3uVNC/FY
9bIe/ArC9x3uH+x7GVD4CF1Rw0BazpkoP4WUyYboOSaXUzSzArJ6CxmcZjrYbFIE9N5NLgB2hpOX
e9bFO/egaZbSXN3BvBjNDpZnVZWSmCIziaDC7WeKsecNzxzHbcZr9BxYzUNDccfRMeik8OsHRkYC
uINfmhqDRjCYT7EObcSlriaRYOV+N4ED3rNTW26A6C9gnEEKs+XdvMImX1NtJ+bTH9s4hNzXmiTB
ldJqpla8hcEA8uG8QjwpfzZVMb+wdzMDV2R+qzO7sd5C3syRqwwV0+2n3xIGuQD/9Q333+BFNgGQ
8O9YyAyrVFkjtzNzHg6JiAf6FH+wtef7r9JutNOoDp6bMnJTc1iLrFcJGwrR6Ozs3Jo8O9FRQCbL
SxX4ohDC9ZHb3P3O0abP+cVNYewZ9Ig30Ntr0JbspzMpimK7Bx1sjm+gY+CIUiMvTE5BiGfMfXYT
eKkCZu9FA7zwicEO4+sH/yBDiI1xHSNSM/D5gdhh1JC+XkbtvEcY0i2Y8bkdPdBmXi867F5sysSU
75+dk7kBVV5FPv6ZV9XdlT5OdG5Dkcbku1o62/yobtqXsrRHzUpLtKDSeXXe5dkmy/uVH9Ys62d1
V1J7edrWJVyu963MV9LRh6+QfbOMJbZGVLM94dytOuOMKbUfCaCEoKfgCfcqrlcm0CgCEaLOwfnI
/W9/SMGNuKQtaZR63KsGyt3STtd/M3we3f8pQrbbXNpmGlXTE+Gx4lhl/kIBjoAyXebvhD6dlyXK
Ig/oTsKAdZjMr0lEI+YqGceKqTkzrQaOLWIZPsBMWFQHQ+VNBfaNygUpChJ8Xi60IghJH/tM3ja9
l/my6YwoT5VmgmqRzzEasg1D6MomTSBwebh9KmsVq6cXXkXqF9Fy2VrSYq0wtJ7OeMYUOtlEKZHG
p0xZbzaT1qWT5G/W5mRzlB2xQjQzutbwLNxtMwtMPPdYHuf07PVjlfEZgR8WrhgN1ZsFxew+OPKN
MNPHlxjaiKguV4Retz08fngzNA3tx3KPKkNyWAs/eyclsIbfwzS+BYYkQJ1vjeQbTjlRJdzoCkze
q6cPLspCqEH/mz+Z5jkEU79oF28DYcSIcKwQ2b0iD52dAD+wxtqKNPUYQEyiF4PTkUdRBfveX82C
dGfoUTHLgaMWhYT6UaEEddgdDCDqHf/92mdUV3Gj2rtXRK9qSsk+1AYJGzUAuzrBkYvlufmDKUrj
R4l9C8SVM8FC0Lt7tMea6VLdkRoSzmgDMjAoza3y5wI00qraTrVU+vYRgtdb9E6pgFPvXyTofr7k
YrwoRBzjRhA9gDfWKoXBC01sno8ITB+xvQd+Hs02Z3GmwbPklC4J8xXyCpS7iZ/o6pl0vgkCvXgY
xhAhaf4NWmiOgdg7tsymC0X8tuuXRWL1r/i3rBRpCz9QSDfrTaE1xcGJcLUQ1j/7BxfvKOZC0fx3
iXqOoZTVI4selPSLGsFvnmeHAnbzfVIaXnZalzImqSAEfX92VN2q5E2i0x+45ycomdhpcSWFhnWC
LL2J/ZV+pdnBeSHt2TzUHyl3xWTGwU6IkwaNkEMQOhqwuRVZMNfW5lP/GmCmzuNmVkzgi6me02jb
nGVF83gd5dfn2q+xsgjwEoYRT6k5LsynyrgzGxB1Cu3epI67/9AP/QEWpIjMHKwVXdjbzUFzAJ4d
JpavWtwHgeUCQxtbgRr9Cux6UwIMM/ubPaVecs5qbnMvl+LRs+Jo7hTmOHOYNGDBmX0crisqDxpy
PrNu7eglq8LhpOUCKZc1z1Y6SsxPn9ZaI1hGnujr263x19PKzyqbCiytxZJqsI17tYQE/+ZVpgsA
pzhgZEfNZw95SctosHkTWd5byf0CEfQeRK2H4u9dbMQ0t5Ho7DKdUdU7+bUUVzxILQgqbnEQYV+D
GZbpbWh/FV56icmg6xpw5N+wuOhCKz4ShrtaU1jvsSf8aH30H+wNBPZjB9mH7hTCg3R/uUQ+IKws
V1BTB9SEIFqfrpPF2UZF8PzeHOrQkrwVW6gCnNNPsheSDV+fPd90YDQ305SDmonDAshybqjb30Sw
hQogmuYmvrXJLeHt+hFB41arYQEvNGxHIaugRg5L3kBNzrG3FRX0OIxKbvue/3n59UNjltiYuYuR
n3T47UZ5mGwsR1gBI9vQhydvhsqjv5eAgwYcI5vywv6ytkbFkqRobCbfHRr4eQ3achgj8yI2sE1+
hQqbYBbtP2nx4rcZI65KAGOUnhPP2pJsL0NawPnk4+HaCjhiVNslW5dbBZAaWB4vfEmucN5bXDfX
XSxId2gbCrp7TalDYxuN2Ct/NL5R8keCQWIYjIsnHTyONNgx1HSZtuktHdTTwDYdHskP+1EqhI7b
OtJJs87tXkq8ZAaeQC9duID84WXWA8f4kRuSQeA56ECqPyf+TI4xZlih2WEoKnXzzLknojerZCFJ
T9J1QhEkbycFqlwBvsVXWBhfWfoS//gCVnIk0eFegY14MU2O/UAD+OxfmfWks1B6pjbKkQqnQEWR
LKWDg7tG+1RgEjxoG8mqZ2+6Zat4EgpYfkpgZYs9RBR3Bfj+4Gbu6qYARP6EFS4MD6lv2HnCFaFV
LBqnn+GlBKgrCyv+syS4TVogR8WAbIbPJ7vSE6S7b+OzRJn6eVCffI4gbEDg8ynu7f2KO/wkGF+5
NXArJkaxn7q+YNwkt7kd+B57tfT/O3RdDWNI3Fkzrc+0PkctjuiwcZN3+zN/N4IrsAfg9/pwa9ZQ
VXtMH+oMIo0vAWJ5wtHkFVCCpbMgU04WSKq+5O2/mGtqB4G/9tvnF3QAOTJoGF12CfAGiLYPC8Nx
UMyNOg5ADLEQIGtd4UObXKogSSQFeuG7U5RKL3OiRz81AFaYmJ/kwWi7KS01Va3rVWoqAz7SexeZ
N/QLuC0Nxnm8y5uFz+dT/VuEnwdHjfDK/IVGM4tBQdK57vVj/tmf0iqJCxxp3Qn4qyyRuPBATdk5
TOBu/69rpipRTZYgsaEHX1pIHY61oDifpnOT9Dipw/4uNxlEJyorZ9BSEoehL6cmNu8NfrbgdXPR
qe5FD4SH+nVV/XZqHoGSGHmC/tigFdNczQ27Kg3HlFC0pSfyUJjqOgr22I49eYQSC90LXPA6tWjX
+b3hf7WgC9hxP7OChrrknjQSL1WJBhH3PbyhwjwH9TyaXX6SvO1HVrO0mQc15bC0lXU40o+IDIha
fwJz+6SlC7ryHgg88JJmYcjgF56fwiVuHMrJdGstvjwSkJWqzhy7TIywsKg8l/ysn3OoB8Rz3d7u
DULp6NZOblbo2jkrcPt7x/OVZbTx468IkWeZRD+7SN2HuoG1DzZDeFFXd/k83uaPSEfdqS38qXS0
83QrUIqEGJItxx0e1vyGUmnWtvVcZSiH41op223wiUTB9dvxg8h7PGgfOv6uAGjI9EzRnj/9B1V5
LN7IGe/yTB26zEdNMUv7S0k8lMXcicUtrp83Vtp8XgfJUofKxoERuhkrsqW0V8y5eByMxyxDNytQ
X1i+UxWmSfeY8IodV36Y2JBnO1rLor0cgJoyLM2f01IHT3PWBDKk75dbzwgOynHKMkdYf8rpRstw
29MXwW+gz757pw//hY/CQNR85IW/reEHghGe2O1ftlebnkt+vR6yT07EbzYneIabO/BLi/UGvgUI
z90jsdsbhKpqnplXcQwfexdMy9LvsUJ287Xb5JObPeQ9y1P1D702EX+BtoPMWUqAgzUSAuPf1OJo
TgocPvlsh5GmqJdVjX++cIftGSZPLFcBlX4uZ1Rpbhi/Lj64p9LiblIr5LQYO2NZ9szT/tcJSUBS
j0PorIIAu5YNBUCyKTve7VL3tcgazKzxyKZBIdwgyPh0lBvA1RmDvt6NknF1IrouVvQGr1FKbwmX
BCIs61XIZKMr0XlLDSbSu9TCcK0/6AQ9DK0VoUQQ2D9u5KKNHkiUwyrRvpdLCeozjstNXN7EIr5b
ItPWe4o0jKlDmwKL12DzjrmoQuXV6QchtRGQdxLW0qEgoOIquz8TUMwphVhWAr8wu5vbMgXhQZj0
4tmZ4vUrINOiI+nKC1hFillTJciIHYF+Zy2H303A/uxT1utAsmbrCEB4y78vLpI17e859On3PfAi
PX4F18FClFhiwamJpY1mwr3m3FXMENv0scBYGIR8zEboCd/Rcf8FhmhlOQrjlHnUmO0eHwxTrMqZ
t5dxabUTTXAeHuI6U0QNS9oDaE0f1NLjy5Y2FoCAombX+GKMq+APsIcwzeJiTF1XM6foe8BLEgN3
dwmEQ3yevA38mLOE3z7zeZOzAeA48NSLz8GwIxRM4j1T2aWDuFM1G4PUmnBwWIemu3bB4uzABmAw
llaKd7rQrVIoUfNmaz/fDrODQno4IjbGT4OHlUvAdGlUtHO6OotYs8JJGVn5aogIqg+sjCUkf5Ob
eIKQhaAeygp1UXG2VUT0TUOJ5xcu6iwZu0QaHMNhsrez+a9+Dyq1jVJKRb/bfkEzWEGo8HlcQ77/
fv1BHF55ss8xs9/s8c/oK3uMEdxml6UH5KPD2/fu41uEWA94yOp+hzoIoHlKXFWuD0fg0at45Yr0
kbt9Pkzn59BNv3NwAb2cNtvEgnqCr71sVjoA/PeMoN3YC8gwDs9ocytMDV7O7+ex4f8RmNNj8aui
tP0OVKpdG7vQFPyZ8zCoFOm6Zi/jBHCiqfZsQ1b2/tPmJJHeeEJ5GVyvm9t0OTVR/PFEyHNl8CEE
X8iP+AcHDZxGENCiiNorZuwoe2ODU94xwMeR5RS4eCVxqvoCkLKd17BEQ53CccLbkfcw2RbdqlsP
8vAP0pykktxBAt8QzmYePr2ZUk4bKjTpFDcgTcmP1QHfIC1QugkPhA3SEXZvu+DStFgTQkDwWETz
1Y4u/MpbZLb3LROzPW7fFxoisQtG7uYf8cXxa6xLUCQOAxA/2HyL2DeumYwOCpHOy6ysDNtSYpmc
t4W14aPiy+EW+NdsNl3Q8ihxZMg3wPuD2yaIWUqS4es+45BmIXPQU+wZiWjvlNX9UiDe+zyGyWc6
tAO0UMthgXX/+mkFXximvku4BpcowNtHRCh8LfRcfYz4PSiQhFz/sho14lSDKOMcAGUN6u5Ljrb3
z5nLv7gunWgyHNt6Xx1hxgZ9NB+UXikeiUdVv+mwxTN5Upr1ZalJ8MAzjnOmON1fQLFteYfoAEnP
KjyPc+od8bF3CWFzFbwQO2cobyZZViXvnmzqeiFlecRZWxNF+6qjImjpY+DIyxNbBcQRz4rFZSzX
StfkbfCUEfP/jijNwEI7REgv9MWLbd8PKRiy+aAjwIrpku/nM4naiV/xbv0QHxTSd399rQ/draZN
VHv2UFciiMmjP0S9056zFyCZu6OldBtr04wzJ+p+CNrMH5XikyyKXd0JnxL7wGnfk/Ro+F5b3MWy
Typ6Tkm2qMXCd9qy80tHfmZ7wFqkYS80LlfEtatQwy1ViYIhXRLSo0Giq88HsQz36DcQ/7LnbVwq
KlmLHchT4cIaTmynetkzO2tl5MEQfv1JCGncE7GgNoCWtandw49kN97z7Xf9yVHy0azxjYpZOljn
Oce6MUpIY07mMBVMJhacRue1w3/gVNlq1PNyR1qgiIeFfvJHjmexl5Y4TPBO3XasaMORNuvXt/Sv
4k2yMVRxYD5wDzb/8vO3HfijMQUC27u7F2Ixwhll2vcviKaE5/E+4lYuLpW66pD1Tsn+rizRwhqH
e5KDw8d+adj0xSKyTqE2fdC7qsmE9vkHWaT07fo9mS7+15Ih+ioAj2Q45c1xEbMaAYf6cNWTJz0G
HCYDchbfz7NCg2GjDTDrESYdMe4eilVQTYDaUYJyIUqR076xn1kfiN777xnASzPqvezWDya7aE04
9XKZv4bEgq8DFcUHWbn5yxzH4tKOKtaTesXYVP7dNPbKpdXEsphQRzOv/4q9HZ4gJtVFX6CPb3fH
mjkhqyzDn/zsNIIvM841lyJ0oVRUNGaueJJAWPnbRnvLzItHeFwxUI8m9vyJtieVnVJvuwZxdvOE
Xk43wgUvwyUWzeKsHOu9w6UAwUI3CuZosb7Rhejbu1uDgVbDiwBctlzzt31M7jXx5ENdf4KeUuv3
uwfoefqPrtzLzeT6ZOz5fCB7HFKwDYj+Fa8eAt+wa4nxW9cADEvONW3amvR/BtBd3UgvHda1T8hb
eNaCKybFl7gsS9VlAUO1xmzFtcw8idC12MWqcBsJFL/tOC5Oum5m4h+nfN//WoeHhGl17gvYSAse
AOAZj3297nAzbj4ozABV7bKU9ipM6gGQ7dPvkiXcBuYpuAnZ2JDFUMwpAV5FprceN06gMknGolNH
rmp+mVD92beGQfHHD1Oyi4Icg+SlfjLsV2MlIOuTgMvJCJPxvCP8FG6+tUAwSNOyA8iOsqBqlLbO
l2MvCa7m5urwMPgfuEvHMqB4Lhlqalt3Si79YNJv0RvyeCXelr4DlTu5FQwuyODeRf2M4Bmxnaxf
4mrGWcMNxNPPus7lOciuXwsf9t0lcGcsnbyo0O0LvWg3kDN7FBtzaeJnjFQnJFjSt0XW5vt1mcIK
ageQIH00xpveObK1xHxkq0+tPTkXQwFIJgEY/XczwxV1NpEqctoYLq43+IZmVvrJ4yAf/fipJUFa
FqwrvaIxOCDnQnvR7t0aY3mA4Ujkp+eDh2DctHwPodk1qRZoN26mx8LiAFDYinmod2nV5OKaVC6N
ahCRvPeQi3AiniER5hHWQGNn693nZlAsASP79hX562YzRFquJWYA+8X1kF7dpF2E/KIvwu5CeSkK
cMwj8jFwztkYTaDiqKZnYenGaXJ89SikzW3fFaE3M5YcatkroMRfwCxTqsd8xeLo6joiAGSfy07Y
Nbop0GV4E0YHBDOTFYYPkqsSa86CVKIWbRdM4GTqfHO4rcbgPtRNM7QhqWOYW5vbIgHwXH2ad5BZ
lkZ1nuQz2qbekv0BX/X5F2LCCunum7mBlimjUhXViwaPLYHtHXm4Zs88v41RHrDiqMSMV+lbUF8H
BDnh+B1yk03Q+KxaZ2xzr/wJk3N0DMmFx5MB3zfqF4u9k/LrOSh4sSlX239pfWeeUKaJdjwYvciQ
7/pUXNBRsCg8aWYW0pdxRJ2Nd9O+gcEWywTo+Yqi8rteSlG3EqYdwh7aeerBjte8jnyCvmt1rmSK
EUJce9b6Hz60jbd2v4TsAtxWSC5QdyzGpyvzKyLKfmYspq23A94mxFsCupYudArkCNEed5kCBOuU
LI+kRNv1aNnqEF/+az31roLcStqeCASsdPU4zkIC+8PQM/n95InqJ7iDX3jYpJlDIU/eCJGhumnC
s1vzsOzc24XuDiW9iTty90JvLTUacRW7QXG2Od+vrtkrF6XR7Ozn3VEkyE7sxJWDvZOOKI7dCecP
qE1pdq9Kcib3HOc6bhQErGJYOvHzRyT37UxE+1GT5q2wPAC6BM1/93XekHtyjbkTzRA7I8/mUq6d
uYFE2bw2SX9PWkgmBqZUAHlWDu3o0Ibx8lYwGb472paoXG2cs5RsreRn1fb+5qxVZDZ9DsSy9doa
H8A5861nk7BnoHPOVmwAXYH5/hAZD9bqkCh/sUCDONYe8W845wP2tKLd1lN+ByfXwHOp93TSD2p8
59v1GCkrgD3w1o+Re00K6z4kfmBmCt5B+dgt9Aa/PyB+eJPl90g4nxxe5m6IpE/AEF4FbjJRrFEm
0vEcddJTwTgb+l7vjmVzeykGRr9WrkxDuSUXTHAoODFh1PD34GKi8787+bqlqi5+6yeTzRRbBAgI
1DNQ+acThNwmOEXDOpLiAqynpcm45vftPLyvZWkDaiGIe7kQB33PrNRM2CWqqUrqkhOtjXGPUOoR
hfTXvQ9+OWdsUoDqF3xLo1gbodhqc7tJsiwYklwFSsTSOntauHGdpnlvLIAkicoo3SR9YayYhudH
D9y3EczK/+J0e4NwQ9GayeH4UPTK2dfn40XyGm7KCXqqvPQTx7EZ0ZCbo+KNbciXkEbWZJRY0AE/
9ZM+wx6wXjWok9DhzrQoxz7AeN7NmLxaVYNc9m3bgPxZ+jOnsxJE3ywTteFD145izWLs+9li7rsU
rxvengrsmqOa6eZ6Z2hjOyhxMmOh2QqmFbYQ5OlKciAE2DPl6jV+nuB2rBPDHn2Cb4AoQhY78ZtI
TclqutPlgn2xDqFd8FZflT+iTTkm2hWYKLjEB63BgbfRSnYUBecHvD1teM7PP/YBBGKyUGYsBJRW
lCKywNRn4AxiK8Qy96Z4pDlHtH9M3SqvF6/U+wJm/oJ48AUJsCgug+2w1nrd/6MycoAlczL0tYFW
zgP0lB4CxnO0DshZ0DQ+jnAjhHspI9ptdu1ocpe6cPDr4BeMFP+lc/FCj9FX8X0MuQ9vXWfi+yPJ
Q5CN+4nzKd96l+AeXX2rkX4b0gE2QhVo9vLViF14VCnf5Q7NBoXG4lhB6agBuv1xsmTlq+jh4tdw
EfOqdRzkJSleliNyXw8N+RhNZVz8zwAvTOtjyXVu4/7f98cc+zq4ZV7PdfsXzeqD4jryn5yJXz3S
BTT+QmEQNgezOU2EwJEoDl7XQpaRNyKprxgGN6YyD1EKo6wQhIC9ZWPbi3z78Zv7DQFv658rl526
qKVnUguHXiJPIariEIyzaKcGnlBiI0HA1dCGjmYHa9URKx3eVU4fWXXAgydc29O0eV79kZGkN70F
8cKievnVe/VJSmF63RnTkjhDJj+rGXVwJSWhk+2LkpQ8HhOzc7dPf84Jj//Xh4Et/JrhIuL1YStK
tfkTRiSX0w9BuJqdX6HS4zOz/6yk8wZnoUjB/qybkJqUT9zZUqssv9vccyQALWB1f5ZdSyuXsI9p
SK6VryGm2T8VvTFFtLa7wWJmNfmDx25Gf+tlTISag4Qc3V5qmYwSlp3oQYMemohzZWra5nHcikBV
Wd50RgdBp0OCt+dJAgYdqRWtw5mWldKCpvsPAXePqKITROkUM5AbujxxOczznPafoBTOnXZFmxZx
ZNwyIkNBahJIDXsVAocgHwPyLm2XlKWpFo0qIL21JM70KHg2g26oht/JzLbdFEQ7ApvfB1o9rcB0
s7yat40wZWdgd5HbVHVI+ApnI2cLpYgG2Mx6szM4m7Hpnconc/2jnwdK7cbRcBxctvBCSXvXOOT1
ls8iA+Wr7ALgnY8pcDIwMc/RiQwl0bz+AA8wxCLeFIV0e2YZuPsm2vlfJz6HxYxwIVhYMHNUqOOj
Do9cFdWl8AVqDZI44hwCTGBr+vfVbwdLHCKnDwgQ2g5305KYI8dgx1ULXerY9piB6YEeyP36IDeh
vFPBSjV71e9S87ULkhfQlhFejpySTzw5KzxvSDHgfFQKwlEyTvHpG0Re5WfCxAEIDMn228YqLbeo
Wz64UzLltoMSmkDtv+GqUZvXWei/5spqV9RBNKewLV6hwWhaKlSuBMzepYQxEjkoIftjl65kTce0
2y+8VO13u4EhuKbo77y9lnw2lc61Hmimx85scO8YgxFFDzlZafjTHsSvSwL7NBrECFOEsHfNeKs1
ccuvNY9Oxjwc1jks/Tp5vOd/fEb9oSrmjLueIJk8YeIZQFsGvSdRC/JyX2pO7/YHhv2hna41Qy5U
I7+K4CzRnXTx1ojdho5YVyrEGcUFvVuejXq4KYmW8wMfQSCKEC+GP+DeeYvjDsts3T9fq/sqyM6r
QUCSGPTNHu2ldrpv2rKDVgUkJZxw+eaREUkEO0BdzlTKHqLcmK6IIr2Ts99yNOx+AoIUN8S66Bbi
/GpUlwZxc0ft8HPza8dc2DBN4HtBoEmca9FY8CkoIzDk8Q/FtzDOuDcEUgSNWm8qrPsHj1JkXLwX
eAn4mDmhIhgmBBVsqmwhqldugdUxe9wtabcBrGpbj0d+w3CCgFHQAc2Zpiai96/ozHhNIEE3gVUE
krLHXGVP3z/lniUBRE9AvL/256YEEWGNK/CFmrEqPVZgD1JkHGJiFVihUxKjKGvKUjTd/vxPVnop
TU9ijiIiMUOkqKJSW+0c9i48kxDFJjHQapv2yda0NX9FjuV+XiCm7bVunadQaEWqiD3k7WDhlKHr
UiKzZRG7oyQbJ/xnUXL6V6tin3achABoHhcKEcsjVvME1DfQTE3pLmiyjaV1Ln4RHMkiBqgp4XDf
q6gC2lpbrjt60Bl2hJotWYYuptUsTEbSkgIx9AwgmajjoG2flag+BrS/FyNRvpeFezLIjwtOeEtn
10ZB34vowMcfcyafpOhjDnApknmyvkNvCebupj1JN/JA3wOTGdIjzWK/YLkrehM9SykJCnm1rFtr
99oIHsFFH8gM+nLuZDjScvkUC5o2Crw0PUWyxVwms7RXYE04fkIAOZ/eg/SF+HFe4v1u3OVzsxRL
AMrHYyYSBi7NiQsPHILra+AzxN859YAXHir70Lus7hOAKU4pWQ0WNjfKPS0MnFMU8fLMHuK4ASbd
9zcv4SMbXegUVWJgQXxxzwcRAXoNmTdlOLKcuiwOeODrlZmI+j0j7/O+BjLgY0hJHbJvbCGPheDb
54DdheiQvm1XxBefbmKyZ2f/sFCt9jxgFNbGt40+SvmNCxN13Ih8LZMy1wnsc/RfbBk62K4ZsE37
4mFBRR9U2s5Tyr8DLcS5tRTdGH9abPS6+jPj/Cxl1DbeuE4NODNDYQ1IOZ5vpKC1emJnqGyDTDrk
AmlUpW1f6Nh0CaJrFVnnO9okBYO1VIWnJDCGVJgLbCQZV5VKDzP6Pm+/y4Q4seK6zJvquDSLWBCT
B0feMIap9MANlPPNQ4Kc8HNSO6Sgi9iyfUTfMXnRd4AXzObyqJYlbq86IX8XLC4MF5Zmq2cM4tWL
YDlR3Vgl2o/Cq/4QjNI1W+mFpBBPFMWOx3Reovffb0nRwSTFTVsq0skEuQRsox0MhAz5y1BrB2vD
aGIdR47gwWzl+HgdlxTFxj2Fh2JP90S8eF2TKHRKU2oapD2I89GmN1d3ul+xGio+FnTnXHXAdq+/
tYtPvDMpstrK3+zYzY15LOiBfUz03XxVk7UT/qy37P4qtxlnWceJN/us+6gUwO03FXARHtvmCVcl
KzC1j67MlIS0HakKHiCS1H2eOz4ZXyiz3MiB92qdUuyTSR7MlxHYSUM+jb/eL4ORR3GUjtmw1jOS
FUb1UyQpv4gEGf1HUFG6Xu5j3rIBi/wJHbEhkgenY7+DAzna6xzOWnWkYqp58VlBiPjytZpsAHoM
62vw+5c1xHz08DUbdby4LOH1mnL+PyXkNZvG5NHjk+isVonEXDXUWIuB5Ab/cWEx/D+xeRfkYmKT
J7kbGeXCKtnk7rRWoF9IDPUqpzaUIM/tzEIN9GTM1jI1VVouuyImPYuqKfzjz1hiyjlfcY4x5hCT
8c/52ZpGJZNzfi4fRDYkBwhjS3BhUo73tHg2ry8TZhXhlUWTCb9AoOE3EcPwdrLcCIYLxwWwwjHl
BCDNeZbiW9E8cbr2RfhZrzUOFSmOPpsiNodvhw6FGJnNmPJB+jLkiJOAPBGE8d+ZrFaEHWqSj28F
abvjKzo/4088L/MbC07z5Dt7a11yvvR/bxBY5aKYXurC1XrcZ9Fm5LjBOEIpnRlIka2IP2Qny9FF
SsvwCe/PUb31hTPcbB9pd7b4sWpFZOXaaZzcuRSkl7u2Vz6UjROv5kECGk5yL9LEvQyK5+M8miR0
WS/csNqDoBPNHvT28FcyQ8TfO0e6EDniiPcu4ohONUL/WgoNwquL3jKLqN7fVqCB7F0FOOiM4gKo
XYam3UVW30pAe9D1tEKueY5pdrPGpIYXKvHiCM5q6FjHdm7lcaSw6i4sgyV1n4usniG0K2eP4JYD
OhZ4hy5FUienf4AhETLc7JwiVhnKugaoGqOEb7NKR1NNfguASYMzbkL9zfUWVXk7E2O6frNAAnu2
OXE3u/84oi81+0bW2wEkcm3DQJVQedtsftCadzyBX4r2lRiu8bK75/67OS5oCXdjGG5cfRyVvXYU
7Aw7Bmz45fMo7Ot4pVjnYo4fu/4FFbcIGNV8P2qycFOaNoF0WNx9AzDMKu5OaQdB2kZ44TxrgUJp
VkgXj2UzH9iXaVEZRrDqy0iXUBFAmDLDhR7B84Fx3wdZi36zDW3zE74rtmjEt9wmsYH5pPJNFTPy
JMnJooUjvE7v/k7ZTRwS6DRiFvAU87EONoHzzAtramIh3Pxxz9cn+ucI2+JJogsUJO2GMp13TG14
dvPx0JTdrsvEvBze7tlf9O+M9b5PaLx64Dc7f8maOF3AFExWUxMyvMtnRQfAzmp+44Hxl0N6DRZ5
TDYHkgJe56/rpjOBgm8QE/iokulozSRLIYDg07WS4vz68ry5GMsHxB+S3VA0rFEBEI6E2ys4dKBQ
t72LaMN1MyUaAp93l6l1RpsYyhtrbM1Vfc3MbhV82plCTwcMAS6Kie3Ofk73GvnttqU6EsSqUkNj
fI9YLAYTexJ7NRXIoFWPvh8J/9zFW3hRBvtYZG4heOzIjE8E6tzbn5I+GYzDJtAVZJ3cXIotqrzy
uGZpxSBXc8v4txrd3oXpM1qGj0W6ApTkCJaCD55yqRp4Bf1xa4S0fv0lpxXDArfRVkwFlfxOhLr5
akWPv5TAB4cSXXyzKy87opADGkoApctgz3ZJzRGzZdm11PWa1zbQKw+6lslfZSlhk1BaI1HDO2DL
k9gXylTjBzkr5SjO2B2Q4Huo2qiXTSupWNfC8CPcI1iUBrNDSmrQiMCtmVx9+W+np3fwyqVzLP52
9ZeyJEvdRYJppQIjeNkzKIvMopTJV3lgvQQpgsoiZ9+y7KyeRe/NNvTomu6MIm6EcLgUcq/5ko7q
S8ROBPPxCY8O0VFju0v8wrGMXxEoxBgBCf+QorQP7MxZ/OWf3/zmjYZOKJ+ijSFBy030GS61BEQm
WNzZy8H+HWTanc51RZdA1RAnfSv+4WfykN8Z8Vr9am6T0TffC15c8soJ58+OeBCsJUhL3pcYs8dr
BhV9euK6XziE1wQidGpdD9kjxxE1pxGyzfQ5JPe2h+I5Vvz3KHsGW0DK2638ThSMPrjSewVOKCha
RGW883ZbVImyfkc1c6UMCujdDsXr9IJ5BHq0Wx0SHaUJoYT+JhRJYB3ioycSiGWiou9oIXeBw3uq
0HzhgNqy3hscsyObP6B0XyLrjst5xEI82/k+ERD2LUKiL5RyI2UZd96p8Djrk+5S7xh1CoqmbtoA
G2gd8n44mDCd2XCXCi/RQIHQIeDo1cEm2YuHDJwIxnKLNOogYcO8h0CJ0IxLxUoaMNGV6Aae11+3
9aD0cVf9WwAMi95zlnES7Efrmjxfo4YGfaB+Q5pGWqqqVbBKRkQcJldAe5vbgx9cUkJcNI4nxQ2R
T3/DQiPKVoQysAzfhPaWzFx+CyXCRgCP7K0F5iPVz3LqqdGEBr90Vg01RHNns+F55ZFTDknRjtK6
2g3YfaJnN6c8C9dwcIS3fJh0NCBHGggfsMCCz+Ft3X2nQJDwMPqK6sc7WSuCVuhAW1K2BHEr7lVQ
aAT97eZ32qFmMbJpfHxpbNtqbbPMavunOHkKJhJVQsw1jpycL0WZcOb1uYn4e1/FQFjEFofPPbAG
Tq6zO34RhnWEl+2oYENWo1VJkGxGO+PK7sR31qHfpKXrqj0X/ECwmJVuID9r66JNmfDQ952tOcrg
pjl5StASPwNpYShdhEoTQjizlkOxWnm1G5zQsmPyKZgFcFrjP0Xpq6sf1lrSmSpGCWDQjxwbIPZb
P+mt0ClbcimD4imFFVcp72jyy3zJPrsN08eAPMpyf9xHwHZTdCJy2XhMWWySeFkyDu3zcXA7wB0W
63+Tt0LCLDmcm5WSBOenIahL6wAwD4eDXXelrin9tVT/tD8rJ2jp5gz2m1tvvwCR4K0nZ2HqLFWO
vZEsm85xw8z1T08/TF2h2YK4V9d4vuU4K4I7veGNUc0ORaHE8TTjiBSI6KU8CoFSJgoc2X0Gc0t7
bgiQOl44eWP6IiwXyqbHlnz/DimcSMx5ZNJD0vdcpNE6/VyxYXiC+UpfJCHnE/7ojvqKLQbJY9+9
SC59SXg7JBZUOQ64pxAkbmWIfT9LbBc5aHpbJlF1bi8yC6iL1AfSgavsAzLrQ2ZcU/SX/MsUwUFg
eiv1Z6B1y/TFSL6Xm88wSPeQokpJY21BHKqgz6tGfxc2aOZ0l4jWW2Hb7w1sPA2BDh5j8XQqbbz4
ZUA8MR5ZOrdo+COACNiTuq5QAju9u2TAcpQcIqm6ozZWGNoR9eho7J+kOtpD5WEGUzD9U+6xQaff
jC46+BASBOmOA+n4db5cyZe52xUiIL8JkfnadFyC5liJmIt+sU65R9SbgvjNXAqM3V2h6YBJU6Hi
48uCFKK+Bf5o/zfJIlgudtg7CIwfIu8YvlxTVvjkQDi4dP5C53Bbk/19KJ4jGGS6osxFD3BkNurh
9M5D1WT7GD5CqCma+naBT1+7zNs2HEUEsmczi2cb99p/8hnQT1siU4qxBMNcfMYQ+XTHyK9uxAuj
THbd+Usml0sfbywdNTrI0YmSUC4qMZ6dMJgt/bX1xdN0IwcZGiRrQhgHYiSO7wewWoTYTVGad1cv
7/QtwofuOGx28uDAzB7lbdY9+E8wql86Jhqtb98JTDuteYMIfYcqpSLp5nypc6/aMm77iYAf5VXR
bx3D7bFejKIWD3xlyEBc7UY9RbXLo9mWjyB2HELq5IqRhM7ECRfwK3Qiz7RvkKRmSS5EZ/5bWN8c
RTbN/CbNJUGcm16WxpMt4cAlAoB0GyGEWRk2ys0M3cDX4BAckc1dhQdWybAN4DQxgo2zeC6NsPkE
jU6+2EDWlH3KqUqzIl3AYbqvgKMssrXuMaX835Y0rjbIrGHxm1OAwBUKYsBnLGJx2fyQIdHK4d6b
/o18bBbqpMfJCv1tyPhtnLjieGIR1+XMsOljKeQvQURVIZzcQwm8iZ2xNXmLxuX2jZQO6tDSuJq1
Lfk1VKpSfWItG1D9ta1aXaDXlvArNbX81/RkJ5dQl5/zpChD3W+7rMmWaWI+nQp4dgb5wQaEjQUM
dperVnBQ91jqzmnzeMt08t0kAvaqY+b5bpfatgy9TnwR8tbn9+4Wm0JtGp6phvepH33uMHq0nPqE
B7fwtrprzh7rq/H++xSB6+BybpMXUNGjtKoQ4MNaEvBM6LZlsa4kJh5aXANDZjeEh6P09yr22KKd
oBVGBtFsi6umD/hA/TnbZhmtWKsv3Q+/pcTO0UUgxTrJX9hJM2dUaGxx+niovizwyEYfwxQltIBh
amEGwmjMgFWvOdxa/xNWdD4nEp6Z6s0VMxkFQ9FQ3ll7Ls61q4kaH/66bl1XMUSlmdXzLH0VYphO
0+mDPbMGiYFYaFraPJKAYzwmu/UeXfXFECfKCzkXBLq3Cy8cFG8Fl4uTJN/EjKfMlIxx4WkIwzdm
91ZACloUjsEsFj2zHX48TkL8LWMV45fNI+tBElWL1y/U5WDyXsJysdxXealNH5U3syhMMzk415jT
RqXOEmWV6pQcZ5+Byve0ggSfSBO9aXfNz/h1tTlSZzCHCXrJIukh4xyJuqiPQfnWQ5VdFFClfyS9
37tcTiZRk2ud/9iNqUdRtOxsMjvSJa38QvlWRh2sa7QGvIPnc/A401JQBAnSXOXTAy7z17rEoxhM
enW+LorB/3RhXAWQjvg5ATZyt04lFj4SLof24fqZ5WtQjBQNY/x1e3DN9zUuDb27mabyGOb1PjKz
zw7x2G3DVyHw0QyVicEUiEb+d0NAcgd4zv/fXaizIYxyaKHoYDUunZAy+vxz/sWpN40egeDQdwiP
wM2aYhZPZ9Lv+wzrtNDjNNKEzHyBUnk9jaowgKYys2+wnVKyprTaan4pn++d4/nI1zF4thxr6+rI
lppZwK1UitjzLi2U02AKtHckCNwI8KXYAA0DNoPX7U68hwE6NWyr/r370EdHZMkkO9JsZZqIgA+r
p1DSjrlq7nN1hUxJeYpqIbjP/P/wIn4o/6sKyim2rzy1l261C1JuVGbsjI8GzPRzqY3++uxadXSa
HGTR8cIYZIetqZKoNgXZvYYfmmotdNGvpUBLbtDawoDT63slc7skkEEyONXJN/FQP2NWs4OLcChR
2DdB2ggAdIOd8jLnjNSwzrv2kVhrQPK3WxLKTUV91JBivXLvW9qNtuGBWmCFp6+q2EUgiv3CHbY3
vKsSqbZmn5yGTbgvZC2or3wL6ukAjl60AawEL5WN35w7I4yJwOg0uv4R4csDA+gA7rhGdh9vjtRh
LTFyTOTbuPBqd72QIC8mjhpYjvlXHg8KvSX8VmHO41mGOA3NAZUn18CbHXPH9eTZXqpRQ6OuPpET
j+mzVePpQysLmzl4l0fS2FAM6bgKCw4eewJbiJ6ZhRZlhVii34fZxJsC5B5O0M/TTRbSJaXmo5M3
H67dDZH9G1trarkJET6doi0sAq2mzWRNsU9z/w0BFkE4URwiO11VEzxBM2II7RcYgrMjM+I4WifK
UnJI8vcP47b9ApdVZgMMcdkT/LyjJEc5tdJaRLjvqEk0kqSSAOPVELTSH538xt9rOj9CByw0koVy
/bSYnSUQyv7IaenYm4cd1rLo1CWc4fuuUgmE2dSQ7IBF/L0NWn6Y0fViMT85Q8LqmRkpJJJtcuID
iWjBoxyUibT0btcgXXbCrLMtUCMru9n0s3Vz8VXsDbPS3+UCVSuSsoqwXAEtRpLjAwo5VN6mG5SV
Qnz598vcViKAjUosOmctfUYx/AlF/vqXr8wZ3rZV6lJW/MF4nfo2P8j0CfwyM4ZFsha3WRnVYraE
tJvaiWawidlJViv8Jl9j2BPZ9NyzeYIdp6bC7M/CqkpMJg+vt+/+spjU4Fj+0nwAv3UsECqWdldH
FomKMYTiCgENjRluP7DN2EdPwk/BEeA1f6ap13gxvYh5rj1VrHAipQXypBUqb8/XlEYLH7MCGhJl
MtYPadWcBtmK0fBDK7lRagZomUujFH/c1nkbukTtL1ol7d6wfilbf7iL0ndusFxfkC2s1fXXCcSB
0LaHZLTO+JVYvAXR2cbsa8qo6fqGATo4R48Y+gAEYmJqhsxg9t7lMxmfcAo3K6YxF+0zDeGxgP2g
ALhzxchIGa+gmPnXYnZWSuZZR0FR1UsITBHB+YlqPvHwc9+bSrDsO3ufgjJYzuOwhDjHDLYL1kB8
l4Ho2fQ9Zritab15Jf8y9FaruSEgFfSplcmYM5EJ6c2C483sTtnB/Ixg9abXnG34ht/b0pWi7TDQ
vYUMcQS89+mGAXWCTsto0676qUygVeqJOfaRuAqF/HkcyMPqyKwsK9Vu92JU3BP4nYvaGA9SUhiw
hmtZntlwoDwomtM3XqYuizLDwpNSsfATyooDavDsEVApo9HgqVDDXuZaH/5Exmq+wiy+7cPvVRut
a8S2DeeXxYgy9HxxTO9X+yGFZnmx6AiSOHZxEp42pBTe8RtupkAijaSu7HBBmi+weyfIFLo/bOz3
xOcOOP0Sysdkzxtquto6T+7GY8FveDAo8bekFE9d5rKJidCU2AXzYWKjNKGsZw6LEzdWO48xEhww
C+Mp7N2WwZ0Akq8hOL9jjJYxpeYIuqLPBDw1Lzlh8AhtLdyOP4YehH4qB2W6SipTGRcEDhFvBEhZ
fj3TQHH/bPwZtHrqnETa3OXET155GF2UVu0iKys9yW5dUPU8S89jTj43wu0g56jXqJ1lxoUB5FK7
CKr5opSy/MrUsJdd1xqO+jjH9OlzYLgizn5ilZ2U8DQwdftNWXBSkYzPGxjQoTaw4iZdtUxp0yEz
5qA3S1ja3L3YdXiKFsbQyNVsW8n27qJM3h/7RczYclTRAVdlqgMfjS1Q5cwVbTeVYi1fN1lqJniS
+3jokbkN5x6vYHeIZYSQcmAaTyHRFanox20yzaUF/OO3vah3nXJC7PK2GLfgh59z/D/tCR9PqXcB
uaye0svKo5McFAh/lQWZuTEEip8wH2y9I8q777bxlDE6ZsFo2IVLdXpym7sX2+VL+uzIqOkACmds
0TDrrYMaP6ONlm8qbLiubfSev7Jfo7xwb5PbETVwvrRnR7lmsN5YEl/6XIhH7+zpMwFpU9t7t2EK
7HhbQejoi5QgejvW9qPjGkiQl0azt8zry6rGcXHIj1JVifZtFUWYlJCqEKo1havbW3b/JGxj25Kh
K0CHwQ0vQovYwdmwk1znRHMkwqMboJB+2RnqVVcCl1vnXrLaEUqx1hAV4jXhwPWnAnbSVZvfsdhT
deTiIYD/mV238BFqQTnbx1ZoexY6ndb+8cLag55djvbf3yKp0Gjo1BtRgti7sb8xx+92i7eJUFHK
czBndf0bChyQhBuryUvLy/eFWsD8fsRNfFkQDFTdtA/rw4dxle0aQumc9KpGy0wThU10oSpOGK+/
+qgoIW2csFFu1xxz4G8fZ7wqS6WrGmK0nsvRUCY8ex+dlqACJBxlziFhEmvYpsLLUY91bWUN9q8T
1AvY9H/TtMl90zDNF57kNGQR5lNNSYDjsNS64YwqUCgrEotZZTiI6T6Ig4AaSJyHLhVR3PcoLAz3
KG1rP8/PeAzXD5fmtidu2cVvf8UdwsyWJN/yUOd/grTARMe9PTWK+QQpBBPw+iMz9HuNyeD12s9E
QqhYi7JtdSIjQTXdE6D9UOvvybrv4h4V1eyNTglO2rvUwue11OXZlMtPgBFfRfd71oNeoggizG8h
wvy0JL7a/S50t388OGeVscvspi6679YJG5lP826TIVVQyTvydCbXP0lmdFOUcMLLeJ1IJ3FrquFI
dogcEPedzqURKgc7Jz4q0IIfo+BqT0V59fKuLTCDVriVgYHIQvVI2zHcXVzxmAbBqdspc+B/cWxb
1ztJGJ8/JStitZ6r50nmRU3L1CHuay3EGIJ4PWvjQVfpxzJX2iIdVXjSm0McKr54JbjK6GjAZL/U
JX9sNhWksldowxT+er52doAi3o9pv0/eFCYg2UdFJ86rIycM3XNE/NEBRT0s8Sri79JXhOqlhdOf
aFss7CSkOKILvVJ7HZGwow6J+meMl5iBvEyR8+TE2FLQpU2DdLRyzpkD6mmIjknVrW91gdyj8hpX
KUn99W6jYMMG3YlbYW4FKHzjO9t58AQSSRrlB9LkrxNq05Qy5TI2eH/HZ5bG581/TPMMMwK3tHAl
n7lJmL67p01HTmgTRPtIfJAkEHzT4/n8pK/x7rJt1J5G2ZDs5VuosCfc/KW1iyEdBWfvJxgD3QCn
172X+H8ZARjRKfr7dfGK6hmFRokYGuaBuOlIKq5pB1ZasSJvr81U3Aa4i7GBGQwSmOS8MjNqDE5z
JSblPRDwrWvDPZs/gaDN5q0WgHHBNJYpTXLA+YlCOdoedIwAjMmo7VpgyHzqhzbB8QuIN02NG5xj
uYmCYWpnD+v1H3eVtx93TblbyedLkGa+oUKU9V7lCnr4HlmtJAEMrzjhiKMzfdPD7V+AjgUPQQut
bp0TGZqmKRRzsNZTY32ZdBMSzvydDTm1hWShKaX406URjm/2gV5OjkMMG/mcML6JYylV5Oy3ZpEZ
JRy3NfN/HU8vGiWJGUymNq1ws79c4grpxRcH7clmNhKxQH2NQx7SCu76nMGxf6nlB4aXa9olB+qr
7wmN+Mph6SNBGquYFmWZmiuMEleEiSRtZeYBswVD1m8DFsmiI6rfrt8DVFrlF31BvnSKY//Y9rp+
HauZdHsP0N5VZHASueRP68OQjjFPYUjqT8kAHRsHA98oRZpWduLGgAxb2NrmlcrrIWlqjalhLkR3
eUYzptduC/jjHAzVbu6tvsNUihtpPy2uaG6gcxVo1GGjZW75pUyWYP1NeEZ3uzQhp3mThuyWEonS
ZizpCdfMCQH8JzsiZAjBZhuruxFrSESV91SSijgVmAKLeFgiTrG/c9ZuJ//lb3CNRLYOQNnQQk7Z
+oAyael7L64VXnSpfsNH3vkPGWz3ANXefiS7AE0dnlidI90OPoWmB4aOQyJygKWeYVsLFBspL0La
HzNj7+Vp2qUUG16pLonyInk1aN4GyWpExNxiHQ+kD1YqxaQGIKPGEFPJatlUay5dTOkNN1KZI2U5
JVDS3JGQ9H2f1KZAwYrH3OnnnfNYnknRb31HqgXI62Y0s777YAHHpyOtA4f+Ycowgqdm1kkk9t7L
GbQZZks3vY+rTEoQokYRGuZVi4VwKVKsXH6AwnE10dXf3/Q146NUiMYXDPi3IGbm7gzcLMrCGqSX
RlAW22094kSE2kLfnbUePNKebKFU395Q5xdkvcLpp75Y9xZnW+UD1JkjYjQntdaYeqHqsAzOezGs
+LFiBR+xyCnlVwWPaFCF+S2wq5lSKKAWkbecMytNkp7LEgEi9JuuTW4uc8M+skq/4g/M88EeCRg8
YuP5394vVH3jpRPjLGO2gqhM80HPhkflNsmxqlbOhu4DldLHl86eW57sKlty3HNLEXxA40kyTkWZ
lJm/q28dyjxW/0uw1zG2wib70FU1DkV+TibT0BvIQ6Cy/p18B01WVkysnpWvRuSMbZzgCc625rYQ
kWs3b9TH5UFC28Ip+hxhBKbqDGNPes8nX2hFnxb6B38bX6jyuf55iAapio36Na5ah4y1mlN7sSZ3
bLHGWXOGX5Qqyn/iuwBOfSplxmX1kT0cEeXe60S0cwSD+nhbKS2SUhvWm67j9XU6Ee/g+Fry0mvO
AbP3SRajcLjBoddaO+wkCU1Wf7TQvSZ4D1uE3uegpCzwU88L95Pf+MnmRmxCFWEDASuEpSoUsM/n
+7IC2kli+ANk+1rbgejsGYUrvKOFhwxaVVk1wS4B5rZLm0vs+2X5UG4IkpI2laAIVoqbVQlzumV/
W/1Afm3k/EdqGkGLZVVt22Xqc4aGCV4W3l8Ngd0Bbv+/COJdLJQmdkMERTf/6eMlaTKzNQdU7Pru
QU8qpEkNWqHh6eOGUy3f5e12sa8lk4z9PWSAIqMFoENNxsy9fHwOadznUx+AWWpXmeLZXh5t2+v/
P5yRcbE9Xnk862+Mj9WQY5n4F0yNnymNhhlhXyefiOAZdqSvBkJawarKeEWf8iEBttF6b86/VNNo
OVJUV6LwV7Vh6p6gCJBppLI2ZQn1m5Si+qvZuJ+dLfX42mwkz0zMBeTe/o+WYiCv26YecLfoS2g+
+2MNWGkuUt/NZ2orawsJOGlOh6zcnwNNBiBd4rfiRAoyTUN/r+3b8ZTerlvTBy4IlIYCkBLObB9b
pw1ZUgt7ivRGnYn/Bkvv7U7LeRXvBQFXJxUhsAV+5IQBQeoMO+nhIjLnZj1DkF3hRPbiqNziu2eV
jtnZI94t7FdK/BmIIantr2hoTKq/3To8llfK0fMRvVJ4TgfdxzfXlcN3XfK0Dhercdzfzwc2mXG/
4hzxQtyTZp0etlrjSDzmo0Z5eSHAdexFysnh7/bu7UIFAmj170QO0rCaSB8jKiRqkDzlIzH00ryB
8mIRdqNE3OmVkZb+Y5nyUflD7A+RTA8AXSpTR8lWfOwg28a94aJ33eMuIF+0cm78BmdQImELdTtG
Ar+X547z59rCUgrwk6qDmXeO3QQua4lvYf5XuxNXycVhhqkZCqF1ObHWodaiyXVeqgNbeMwuLsjZ
IqfpgLTt2er0d/oHrHfKAaKiyk6vTCjMLIS4cnBOY1a/QKQEOmJYbD2fLilp8o1YRiVeYgt5VhI6
jC0VZwrNCV+3PLTJGslex3QsAIyRA5wFX33MiRVb7WtZqFBc5RFruG5Ym/dweqPbktbX1yeNruIo
LUMmr8f+UxmfT0mx6d7DK0vEoABs7cKTPPaidk2LaJsyjVhYsRyK9BOnfbbCBaMzooKI4PPGqaVO
qiz7/uukQCIc5fEhXYrHpuyM3tm8UUgHoxPza5Q7Aw/KONgzTcSRCEq4C+1RP2njwo0MxaI5pPdY
q+ennQIy0qxeK0YZoaz1DUkixkaWaFS4wsDebRsUX1Bq25BqGagjAjIPQwICM12qwMek4NWIenBf
R7msJeAl0OUhyBlzC/Rhmo+PVOhs8YrjSN6U8soCiLjHlsjeVRA4I/IApmAGaqku9/dmPkJclPHd
CDUUROfNju2n1XV9zu52zW38OYH845sS6s6oB5ZADsN5MNmeVWHnqAmgFReHWSPfqV9Ufjp+rwU/
EfRoACQD0zzFep0/TlrVAbWVlEv+6ccnV/AHdP+zfT+Mk70ZRUXujvb6RLiLch5FL6reuXKMAL8H
FqrD3gfmcrZF562IX2PZb+PJ4DY20XIsOxFRxY6+5RA1fmJORsYr5ua0/boPEZu8aeQx6Qxnlrw/
I/uBKanf84HzslEaUTo0i+fLmcLSvGRrU0NHgF4RygNaJxrQpkAi6eniahg7FoU73s5niYUCoTor
lfKLDLByg1fWT7YACd6FCZCldmv76NU5Ekdli5CAlhEethA/HqCxOSOp9JF5/jbhsBjCvNJCUDUB
LeQ+L7QMch65r4TlWzS/yJYqGhfy0bpivcyaiQl0xB1I6FT/cNEj3KRNuypYPGCdGHPwudmToywl
bz/tFoNi7eAt+426begkXvY6CDylQjh1S2aGNeSoxDsDrPwj6iabSlLL2kgVQvSN4CEQCP/eLPml
thgJwfItBN49ZrfADg3Xf5urgS9uhWQNmT37YSYE0o+ctYi657XSUoS/Ph67dVER/vF6Ujj22Q0+
slxzCTnbt8DLBasxqbY7V3Fkaib8Ebx1znQtk8EMOkVFJbUGZSjdIn4tkHszOCWkPfyXBNjWsDtN
Vu4lY/W7DqgvXIdIRaqzdSNW64RYiCkl7FZg7sZaE9tO+l9Zvh2EV1cmfoOupw2FyichZTs9jsZJ
gnqXUAljIALPvNXiyLpiSm1aFH0uCpXBLfyjg6UM4uNbGoogV5qJY12Pqx22a7K8Iro1JtEfGn3O
Aec3wtWW/e0vTWUh6O97pRGl4a3Laznyb0HxUEY0nGogaVIPu6kCiTM6WLehT5Hs3nHpemk4OasD
God+xL4YyZ7tl/6851uQ6l4/cywsVGpPvaiMVjGcf0X7uHxKH3w/wbL5W7NMo/vSXkemfSOLf/Hh
hFEy3ejFKJ/DSoDCQqkM6FWCQqfn4YyZ4Qdy7Tx/xhpsb0akvC/0xj1GftmiCG9f5vTomLPPgJgo
pfp7t3C+5oDqch/KxRstslbE6QIm3kENhv7KJxgfI8eHGOsvwSCw7x8VuicXA9en53FOm5lf1zsA
jzC1KNOWfhGq9tE0szfIrNTlOHojsnNdFwUvhnCLaC3A3tKTYF3zpQcLlqz+SuUDXNbrZhvdTHah
5jfvf7xLw/mDdIzV+RZ0izPhphX6LQUhQCnAwBTlGcKNf2ycNbHwc517LUr9Ae+A1wLEH8F3t6Wf
YIAW6YGLHTL0eMfWxg1tdxejlg4NWqirifp4zaDBWUTGpiWl6lUMDHJSRrZbAorZJ5z8o3tOHPQd
xkpeBJFeXt6jTfX7mnWtl7oqjSITEEwGVZbd2YX6Jec/cqkqh9iVr/h7rNduZf1xaetc6y1IJ4lu
hOQol22X9bqTugDk0snaSp8g53xCDfqBLyEQiQvUSkgFDpxEqmqyQG07FzQxKtOURYH4pRdoF+lO
zRU/FCtunjFPvHG09+3VE70gPbDsCYoqt8fWBhYUY8iLo1uZEyFFAURkh3tfgLy0odkxAW7u1iwe
of83wHEce/KV4NxSX+jBSloQiHu/PZHA8ZVxMfLQESmP887e6uezMs9onAwvo+MPi3XhGDz43ygq
OSVanA3k0ABwqrxxVI9v1IAZxNWMztJ+/npnqNz7m+FdCi+uPqoHzkGRYxK7W6/30gSQT0ABg0sY
MbStTfGEkb9GXOQ9GXVGGVbY+zYIoLAHVNrNwvLdryZWpwRk4mQqsJUV5sRFXOt3ygIzHl9Faqbz
RSYlzVKtCZBULVVTMgk+WpnLj9a8MUbTmKXIEInpZJWsAisN9KRWMNUL7k7IQ7UQXoea1GYbyeuL
BwxbDAcKUdVW/SDK0KrEuAbujz2mVHohoZiHAh/9Wm9bv4qFXfW369LgpP4AQazFQ4oymeJJFWKd
BWyh7xhPpO15EUyYyVQxoYfZxQuvxWtg2/3P+amMcHDVkci1HHpANVFUIw7LE4I0R98XEqMR5TQU
2JLLYTnoIeQ2XHbJSgalGmPWyZYOOhFZLVjOotS/gocFUqwjQeoEsO5rOsPQoFRuZwRpeAOqC4tb
BrMFImiR4qj0DsIEKeWR+yWo8mWE6EfC0M4vq0vW752sD3t4gMjgmpqqxdvJAWcAFfcgXQt5PHZ8
3iG2G+4Gak0e10qJvYFSvmL1KzNFwxjLBZfzBlV+FT2OiY3djevHb7uALeERh8yE3/mnh6a3m2EJ
CvsXKj2YQi8MajqeCIoXpoVx8/WjytBDg5qACSwCL4MNc+qtpT75j6eOh4TxINDFUAiA9+7VOD5p
HmaN2irx6n/AzD57gCRLpulMuLpgt7FUONkeN3JghsXtDSWdwqkPfH1Tv9I2Lr2K7Ncc+bWVpOyn
WdCqOlE3hhPz00dkgd5AYAgGKhIcKmCibrwyIHq+EfdtZZabBB/pod3otv4x3TDHa7ao3PpzfIr1
EzhK5QF8N8ZOAg3lHhH00n/uA/lKmU2G4Yj2xIgifDc8J0GfzyFrLdAECbYJFp2EUOeOP1B7Ro8F
cn6SFBzlfeLOuqM2f5iFvONqWDJh/a+kLpb4bAu3vo7VJ2+tZf1KhFZeeC9CvT5VINyOEzNEhxOU
gnpQA7u9gWAoa/P6p6iokdk4JZLBNFWl+m7SD+WnZNUzNjxkEUdIG7nhH8LhjlHHVJyPlCxt+kfR
IVuNr9PgTLD7G0Hf9jNGev49eF6ZjAcQM1nxIc2TGqnoPE0odeWrh+YXm0g/pMRvq+gV/EBc07hU
aXGRMxTd5ksLg23/Leo/jwR3wwcT91z4UATC7DaLFPRQZC+V/e9XkUVxD1x9kFiSPCKDw3frzO7D
jajrZJQKlsOdP/qxvw/E3hGW+RkjEpKdsFI42oD8rA8kIqAwz4lA0Qr0LD/Umnr8yyzaarRdlzpC
mkCFW79sBIfqjJ9mTiRb83gpMVYMevT09zjYTfIz8ysgf7XRkoHiQdgMWY9vQ9q3MlktMuJZtRDA
ykxUCZndTVREH6MiSFjp7iNfLIp75iS9D2ImWza2pGJ8wDyWUY2RCg4+KRBI6+uQuErnL6bcM8KT
JkJij7WTsHJEa+gqVCRFBUDRCHF0jPsi0Te7q2YtQnk2tOB4PizXxqx3DZl8966DPajpQq5utUCv
PobekFA86pNPCUyRZos4EBZ8beSY74RNgvw0r1m7ffRGqfWxLuA98jd2mtybCb6bXNpggJJ0bRUa
aZOmg9mVko1ppvPMw4uLKHypj4rq10cRd9h0l62ODqeM6SVkCp5SfLhniLgKmxOAwdPYoPV6rJL8
J2IJ9jgHY6eqAIOvgVdCjaS3Y00dpjDnR8NyLEyjZ3Z6ovQL9njVy2iUOv/OClRajy2bf++QSYcg
bZcg5VdgdAPKXx2DhqWPyNOaXTzHCFWQJNVtn0Ht+ChqoMS1ucESa211ORFC4NEOCGeFMN1f07bu
lDATcDj2F7cFpCkKdArzBhZH5u9kUE31u9lvHPa4m9SqjJcQGdcvoHAQJ2r8rWZ8whpcIgcApGFv
h80ei3f5a5HRxFD5gJSIMw+8pklXfnLE4k1R/+vMYGddpNGHJgZ9FAIsl9PTQSqtfwFQGnVFYw7h
RAWO7+uC6P0qs/I/6/pJpYPEzf38W7ShjAeHch6aJpSe9xwnqHpZ0rrC/dh7sMMvroL0ObrnCbiv
qt2TOwnB0P/8Ly8iAC2zo00QKRJw+d7CaVazx9OqAk7nRnEphlS8F7uaV/hH1n0wgLyjM/wfQQ/9
8Kr2AbEgke4ee59yrYWj2e1uOMi/QtKIeEkSXOjQBh9xsDjtfpwBjwZJ00Kxo40yZ0aubJ65r3i5
OIcAqdtcOF8KezIJ7I4navgXTumwC+b8G8bjdQQ7P2sGTzki/b1Wx0C2RxDT+AkMyGhiSEj969ww
7UTTdHrQ1Nx6t+NG9V4ADCFAin09zpdiuW4gjVOuUmwKxgRt9j3RHJ2sHnQTRPyKFVs7LJ+gqfJT
OMLwdguHMKDFVlRxgBLN06XuKQueAiRJWYoyg2ac/vNsgy2RsIpUNFjJssq0LToud1XU5YeWMozO
mx7YwcfP15L1cXVgigEEE5u0qnaKoPQoUYE+3AVzUcHq1mgngss9+UCvEYgZ9gg6kJWz8luBRbtH
DKcz6rG6OlFgTd+Udzk9XTSeKA2+MKNS3lZSDeqxp4MVgt4yel+FOZKhpwoSok8uezMpGCZqqMtj
bXFC1RhXvdLt7CjANQ2IGjw54IvlDaAoxEr1MHiXj5204PLQgV6GtRyPHEwqdbHtY4xdjirTtXue
h5v9jRryhTnDIDooIdwg80UepPaqpdWRwxxNIg4JDwCoQoHD9rl9+UnJtzNhDDhlMcfp1ojjJce1
YzC/XNaJT3GdFhlCUB6+zpADPMTKN4Vz4U1ppaVdTbsECvcYCVbJ+GcLfDc1+moEmhdVIXddROyz
I0adePzXKFklWzjZ+leU0fv+jsrxuhLELkg0Z6C2NoO1RTKyLh3/sZGpVO1J74daHQy++dDZARUB
yVJ8Pgo49yuO9bUzEPOAr1N87f3bxfaJ2FvrlDoCGF5FuCx/85RHM3IAti+fEhIe6UXnvkKNYhVg
fn4mjp01sHjyBvsHxmlm2F7+pLsT+bSFRmi8VJ7wnhj6dSY51a+HhtMood3Lj5jQf36VO6Sd9PaP
822UPUd6R5ftYGC9BEzyZeNxfhT85QYlbjb2514y8Ew0d5mOK3OWx6zlEmFBvm+JVh2AhheSvw+U
QlF46ueVL8Ztdwc3r/G5+JH5OQnEV4CzEg/JoCjOob3tiQjr/VGgzAxYT3dZm2xwkS/D70mEJDBp
/S/8gz6KWpmmy2bqMC82Ct9Mt52DL5+jUqaNLdyfpLS96gFtQ0OxWHQvyVoCsSkz4z18ZfgZRu5S
k9H9vKKu2D2VT60l2JKY/80ei9qF6iImK99AXkX5dlyFSMxU1QkSEJTs+k2EHajZNZvNYH5SLx4b
Zlnwk/5QtRaQavmzVSEirXtE9oh9GeueknNSiwfV269HYNLjEgk1NqJe95D7o//KKHvVOAtkM65S
e9IurTWJcBJmi9/2GQmQLmsJJD66obErHUd4sdnUcwas1JckAnh2Dda9h+G+ubrbok3QLO0+mACo
MhmSySmdRHwfrVHbYIzINfPPWsStLtUZCW31Pwl12YM/haQao9HmPdFq7tqlpFCsmdO51S2zsTu2
Q1ZstX6+BYy1nlg9hHih4QjTY4FlYxxy+pMBPWvxjGUTT/2O4eN+AgkOdKkkGbcSraEpRXCcVnwo
mdEIDYJ8lw5JnQGhuzG2tD0DgHcFIiWyU8PlxG4rPaD+hf74pBLe21Nxw6xkvNg+IEyy5DNWb8qU
bS3L2hD8Njqw4rLZXpoYECDL1HVwo6uk4npCr4RFjkk0cI8IEFiRAlyEv4gHjN3y4zS4NVSP2wZ1
oO4sjEH5QexQm5J+TLDFahm6NNuiJJnGHYtnEfF1vTYr0NNDOqYH/mRd5L51CsU7ky+RAORKVcu3
uXJ2FjwrO+9cQPINDx/lvJHzuIbLrxpkkBrT61hI3S5wR8FoGyBP/t1bu+IS4lNaJhQYEiWJkdzh
Up4xno7PBgYMJJCnWMUgIRoDB+h41CTxU3VIDT2ViWnADQHo5MyD144upgyfC+Emo5wlqPsmoFrg
nfuG6npT86ikIu2ELMjZIcaO4u3pwhe/Y+uCwM0NuOO10DBf32xbwV02CgYXUnRV4Um0dpNyXaSV
HZtwv4Wj0VBhoNqhMPRTYBs9zHH5iZ2i8nmvSGcpyIDDYZOhIGlXglCxh/GZHuPY/VqILA/+ZIT7
wVm7Nu/mIjq6uyUvRqYfFSapvIAULcMsBB9RpseXCTTH+40F8tYROpplUyUIRC53/oUye0o7yrft
SPqNtCtXfcgIP2EigNZJOd5VnhzIbdhr6salBUVqZXZonC5UPQhm450FRxImPpiOQQrlVqzs3mA+
N5xs/g/kC9gJIUQPyv68fw+GE4h/6HsdHfctfv14SNmcbFIPSVttTIBPSIsspHYSIbKf3lCS/zyS
E2ZXXgzqoJFmcOZSLeM7DNU8zpMjgXTBBBj4zA5br9GTSu6pvL6Al4uA033H78YqL5r2S2VwW9iJ
r6GrCP3btISIYDj/bBCiYggWEiD06hnh88dRXqnEAFQLXrSFtoXaD+O73oiMicrBvWJ+0CvAe3Ly
+etxpFdv4/AbYxZ4OiH64szpMMqWdbxrP2i+Dl5DrjaSK3Q6XWoL0lWmh48kyYMZWKq04X4OfTEy
62lZeNugvWMpAVA7lveVlqlXaUWMnCbwG0dVofU9p/D1i10vFWLe/9GiULUR09brOIjh+GodQF+p
U91k1JFEp+ZaAsmoOJII3wFARbbnaujcNSL6poOmBCVE2ZoQ7gav68csRUo7FQfXDb0ewgK3igL1
zV14nkVU46B6AENHFrWCEEuosMwPVtvC/z18udtSKpSK2salfzR/xobsfbDN0/ZPTVRYn3kh60qH
xQl4AUunNBZrzH0Qz5rLhoOwFay8K0PjYG9rxJfLP6ekn9tRWbyTB2oDTOapuuDn+inMyh2Og4H7
O5z0GelR0laaeKt5P7/sC0Zk+RL0M1hSoWEfJNJ8dktm7+0cInvSKuXCXLtO83QtABbz5EoPA7Sc
/VFHQDfuyBePkFuoQCb1ObZeYmLMTELUIg76xhbuxpmwcuFdoPWaFCFSwXpZwOykyUhWvehabWpY
De8WCQ6L/Zgpzq4Aa+pTAvEzpOTokUMt9TQlezefL63hBOBHsxTJAFx26svAj14H5Ll78HTJzU8J
fDTiXn21irCzCl+nQ8dsCvcXi5oB73fi7uKybwzwhLpAlJUo9dbtXrFJCgBXtnB5/qJWn47/BvEr
tR0wLT60YUCW3F591+PTzKFG2JO+8RMru4pMF0t1N7fx82JWkZhge1MU2FxvgUE+hYUQttf5gsea
Uvy71P8UkhKTZ1ZMHT+ljuxaztZeaNw1efqP7r8DnkEifO3O7Bgm177TI2Gl48/3xwqleEx9LBq/
IUlBAn942RK6fAHXnb2ZQe338ERxqncgLM6DIIInJvVDZigX3x7iiKNQI3y6jaMayrXmAGtgghsc
jioOVfO6/Jv9tpyxrStkhA+xe6euXDh8jHvGfVT27lBVVUjpfFT54bUMl2g3u+wnQlN+1VHoGbxm
WWLar7ANZ5BnBNVM5FMgFyubezjo0oa8ZNChSg7AALcZmf48QTFv2dekS+EdKSwxRpZSB6+50QKl
qdUEuESeJeHBd1H1jBN/WTTquHPwP9p7pIPTVzAsTPoi9yz4ric0Rjb7aOp5fhBWZH+kMEaKPrQQ
rkaiVxs1jJxVojcpoIzbpq5lSILJxE7XDGD++iTY8th0HvT2xGKjKtCMFkZf3x/Wuh91ZTCqwCKc
cophtCwE10JtIeLuEppFgkY9kGvFdXMrJF5+1bVVCFQCFeTbyiynawk9GCitrtbmlsg7VNbd7d0M
hLlLC0Gz1KMfseqnFWvBd8cORgZ91XEw24/97rp+Yw8McoTKZU7g6TWPXvPEWrc7CP401G266qQL
9zG2eJwe+7Xl05FYNHDtBney8YqhG2NOxZ/j140oIwHwESIiKdKo23RmXSHs+EIuO1UgYcwjLCzq
08oZ9Lid8ZDgjE9AMJbq19DN8Q3nPRu3M9Nn+7JV/YIGNksKk45T3S3nj3/n8uyenCobygdlihz4
p/EyxvoCBrO/SKrNWM2my9jgT4WdgMmYOE4ZEuyJop98cgLQ38Yklye7CwjqxQ11GsSHYcKw/Fqg
ZEfzSfo3expNs2iRa2rls2XxrTTGSBUIWrJV2YnJaNXIKOBDw4LPX3L7ufqz7UaqI1uM3rDZh6Nu
EuJF0PVjmTffLH2Go7Fz6y8s7OghL+zaDoXwN4mpF8xaLKbFg5cfD3tPl++9P8IdUNPNVu9wHR5v
ot00PvSgz/niLfnhgWxzgd+iUhSQ3Cl05zUoIsjcZpt2aIloriOaY0BW6L2gqXpgZ3kurK2KVj2/
UV0EuZMdPN1lvxqSEw/uBAP/fv6AH/AfZ2kfso3GXBZ3p905Sb/Pl4ZiRaF4tGTB09lwZHLwqc3Z
lBMSJLYrjCuhJ7MmUJtAiKlg4BkxPcxgT7H7a8suk/i9cgVkwiK2btnSUKC1BxMvS+qZgcWy8/K6
2K5bGy8k0ArgFcqS/3sMx02Vej+kcYe7jS4BPeTIdpb6b6sVm3duTTB1V8y2HibdxEmr25Q1dd/w
bxsvnsgSFUBNa5C3m+EuShvoa1VTImFHfpZmmHurh+h4jBVR6wySVbVzRhutIH29ejLj6sS2ydRG
FooyddVFhjHRMU70oBKLUX1lhX5SOdKYmcw7mfyt8f4ZMn/Rp8MTgi4LUIhjp71dm47dpoLZhDa4
tCb+jqqM2DpyzJ5ebGSp1Jx2kUgTQRd9maiarQW9zhjsr9CfZnonRxcm7iollti+fUG631yG0byy
n0ddC1roBXm3utuHWoLA77BbOtRPdGdFu4DfvMMLuCXFcDytc2VMHJQ2ggvxdXinRNGMOaeD10id
PuUJBagi6RfoGiALBuV8doUy7XnedrEyjitNdIFbjLbIrJFLm7mYVZnGzqZjOREtecWBGFQkrWpD
kgNCPqfV5zLSvkPaWqQ4jYDqFWgZXd0dKdbbbLqihzFmxwe7GxzEDpZ5VNm1keOdDhyQscJJsvne
+1uq9FszknWoUAU07P3UGbSiuWQz/QQrTFBWBIPIMT6FNKTeU2bLv9UZOtUW2YtdTQ0yO8H+45HO
mxaYqeoyONUzlbkjQU5h74OM+t7Pkz1iIhSO/T5OgEtTLpNyRIRFKsY1HwHabjFy+JEMuZINOWvw
DKZEZsF0gxJX1ABh1hQEHoOCasyupKtXxz3fntRBpmmw7ruMpyz2wpjQ3IBq3slYIKeZl7yqwZPL
iB+dEnyxJk/qIQnynCny9U4vn6SPFFfij43rShsI6gEa2rbcnEiIVWzJTgNzpS5R2jQ0RPi0tu+D
I2WmOaly7ZPAiDg+9dzFB+UV1IubdiIBDZRWgI9HxhKGESvroSZ+NscM5kp0PTedo/EqWjUrDEfF
CG59DCcYM7pYO7wBKdSWo2lRE8BUMO+AQha3BVkNbZwDH1LnYgiyfIo2MMv3xpskC+jmTtb8u5to
mat7e3ywXUp14P+tyN58xbsYBQd0n0vfD+GAfSGQulC62JAaZm4ZSAfKXMxaRlSB0gzMMZxa7lEk
9OFcZs3sWVjptk6350AJNhTXVonqNFmjM4yZSVM9+5oHCN8jgsv3TiqinYDRacnu/dmI9No7D/ID
EtvXPMBu7eoa3Zg8v9cms/W4SKTaJI5lbLPkcFrEWnVY9NaSrrwWKO8yakFscRrVE6QfuYyZPlNI
NhyTTxWyb+k1zakrvryy6wK9mW0LjLjZ7hZAD94P6UXHxohYz4YAEK6T6z3VFC1DvC1WEpStaTmM
BX5r7Yi8q5J+CfD65xRd1LYJRQn+QY8hZWLvVQQM1DMUWrNis9MEPt00G1uYSOUd1RSJFtXVnB6Z
nxrnnZbLPDbuuHJ4ZhmZZ5CFg58ZZ1as1hWCawa/nIA0WJwBz5lo0DWitSuczzBbBBfn1tFaYxQc
QFCc0SfqcNUkYLsio16QwSXrfZH9RMVeQ42AIYzmWySSOCtJNGxZNEehsdOOjG0slkl1H9P3P59B
JpUurOcfFaswY9CLOZ0GdGJqqFET42R8OpJtsBkEsucVkmbe13/LPuQRBMxMq4/GNUSlXF1yXX48
sZZ3PY+6Vtf0h8q0B9Id9nh0KdXQUi44eBV2ZZU0OMYTZ0Ar2Uc9gd/+ErUF38PTMgYG395j6SJn
mywgIiYU0JLXrlZzSLdm5B+TsZXcOljjnaRRPQYPzCLJ3E/+4Pk4sYS2b2mivc6TMwcd7u1mgNkQ
+npXYRndEB4T6OUeRFbm5ZEAQlQlNVsZM07ev0MnOJYmsJ9+ppqc49fwKNxwBghXlR9YxB006ysM
l0m7wRbjqR5P9r5OTN4E4D/FXeLSl/uT/YhrJbnqH4TjPG+nRTef+gKwaBsGllGszGwRwVJ2Rjpk
ktTRax+MDjWRpEZ0QNy6sfsdEYN/KoA3yaADlX86LtSXeHzTaBiR53ZR0zONNhSk7UM/oAf2zHlf
cSelmWJ+pJ6/IL6ydgFIZUTVuiyUK7/g1pYGpDhjc/ODvhiHjDnASQstlyfeVFGkf6kmUcfEEr6g
qsJBY3mCa/BEFr8elo4WFvbpeaCAr3rjqLuLBL/TXJ7T8v9MPKzho06RkhPOEjrzfYmRtoT6Ycne
NrgVQcYxOq0j65tofxeeNGSVfAmwYlyZAJYmQUThIWJfrRtgQwq4s7dJKc3Bt3Sql/7sNIPtp+8u
u6iTOb+2nJEKpglQ0EWRaHuwel+I8iICiDo7wXM+3u0UYppikU6iTB812NUKIo/+7c0ba8VjT7wU
nEiEod//akYuLKKBgz1SnUllIln5mky6SgBE7Odi6B06ARiPIc8SKCG36KvtLFdZySjMeb7MJUWb
H943AkxrJ5aC00oE7yL3Rk2qOhAxhCyLvmNOnOc5imZ0aQtJJsfhwwnaPXznOj92XVLH+C2KbU3C
XW5DqQvoJyJUXeeCSHB6VSpZsUEi4AtY7+HgkdaAQF6zn1ql8sczwnb+sTaph+EmwZOH23/YJQf/
DnFZKKloq1cyz0kEt3/nwGUwAqx47YUHJN1aUgQeioJFLud4TrEx+IZfkaWqAnkQtrAKirP3Nem4
IKBOXzE2vZP6Od5+EN4kCtLiWwKh7uBmPVrQbHHeUaBcasyK/F/pD4CJsi5zJn+gkx0i4eLPh+Ln
TKxHt1HK4uaxzw3fblNtzmd26Gasm527BRbMdPq/oS1Gx5xq9YdYJFDusbpKD2zHvMbL0T+j+j9T
wtHT+S4f0cP1x0+vn6oauwpPLLCm2L4p5/Vhz2G9uDxVYk594A9ur3pSmS0beNe5VLpYe/5BxfbI
M0UElgvXohv3TebcqxCqc3iAzx3zKvTGG+e3kKwoQKjO/M8ZgGpj6w3lgkBT+dJfzKCmV1iTc7nY
u/S8dcxk/kpGAgdwQoA7sQ/gXDy74DEnI7ZVnR7rEVXJlpJ2AvBuLk0NgyPAGv5BSLzgr3lzA/gs
Ca2PozUblrton3/nhzH1CEfI5T0joRJkoO88nHrGNdA/3Cmz2TEalYOkxFEfuT4EaCFZlO/N469p
XzF6N0HN0uaJJXPd4HgafOyaMPn8j5XnYBvfp5/oywM43fomKlVCpq4jzkXErNDZ/gHwWXWTffS3
UX/ZMWmp9w3It5YavrqXwXjalsgx4MfjPiCzy24c5D73scqB9O7Q+LSn6bwCVzv4qwLr+XNTnIdu
VmJ+7XEZNR1Jtf/F7ycuDmg1T5VTxMWOhJqROAYpEWYIwfo3VFy3ZEyh9wLsV25aUYFGmN7h/j+a
Q/kpYdJB4qVus79ToX9WwXgtxF+LwyRKKy4cgmqYnhCmLehhN3lSdZS54xG9Bdnj8eSR16NkBSly
euWuNbT0JuM5vmP4/n5vg8Hf+/kUFL4nbuiAmTmPcG9oux2vxarIcj2hpWn+wLvZld6O8nzvDEnR
pOkMdvS40HQN4MYZpb2rq3ShLxsjl9GK7EahG/+ueELQhSF2l1a40+AoKXfoAxuSn+xsPchG5zLc
YKatdq3S6TL2qLwAIBG3P7Lmg86ovRudZCpQw1UeQ4m56Z8mpTCr8Vez6Cr6HTQtbqC9OXe94qSd
Z1Lm19Wvdggz9vrQOSq2Ca36gYiyse21FIiY/517ftYjdmzSDEiqMe0QuuqJLmvzUHxTXwOqd74o
LLSyTje1RgXi33sAtOxAqo52e0AO9gKIdtBchSAH4wKDdeyAzZ3nQnIq4PUQVnQhxZgIDCJjpEW3
x1481e0qnkpW2lFyGmaAQYiWOXoqKHBDdWFQOLU60SiVTlTStY8W6SXtAQp5ZJi+h+/H7PSQ/Jhd
9a2SF74TsGWK5JE1Ncr+E0JcmoZvyLEBYg6Jlj6tOQ1FdgN2euPGR5Ahv3TVF129ZoCVHs8swzF5
T3N2ehSOkbIKDQFlIf/cmef1Mwq0u8i1BgfOoDy7vUtMOQfx/sU09+2PvA2gfivTy9yRu49gJ5Oy
GRHzMHnXCQK5n/2Bxm3q0z43SEPwnOnrsibGa4pCopJvn6bRWPM5dpyZ0bEdGGTVU+KQN6HH6NmY
c1kHpFdcSeQDrmu1DVAyBs2mbWY3BvwFHSGzb4y3vX3XKMvkmMzWpZZa0Pv1SXSs6p+CW+9eEJA5
hxgj6JnV3QqAQ1mABD+BkbP2PJzGTrIOhCu4+UJC4jMV3ty0t5ljlELHKe0xnlHmEPmwTvPu8LpA
gGtkpgFhALYFuw50qldET2J+tBh+DblNRenVBpzlSGtNU/r3oSP5kcDLkeAoYcaBMKm4aFhsFnKW
3o4xuR2BcFgjxV/kG2htSrOGSvBxLEy6ct5gK99reKJRpO1gxFVj+desd5sVY8jO1cHofJMNDAVF
3kcAl7WmAFWhmEgwA/Z9JABr6pl75dziBKQ9fxpNpOVj3VwoIeaHeoZc9mochXG5kSqaiq+N+s4q
hZPKYkbZsvuya4Ne4CTtWITZrKf8XqEqmFxslRh6wRBnyoCfqTG+XemMGANUhEFQRi01GiJRJXmL
DzKycAQaJCbuW0CSANQ21kH+sRFJ6nrNp7m/Rn6FgG2o4LhXzL7KY4UmlfEzi16GPojf/+yrNYsE
QvSswwg1eaKLk0ORDeop+DE1NRH8NkwNUH46RCBoa9gLJgcqhv4iIM9M+tUIgrt2gB5tIxg9y8Nb
vPt3EWPgQVvWt6IaLxpsThs30cnIZYMphGqJWqkKFroTRRqOQeIVNQJa4cdU1imMdZJb/tqsVutH
2UGQNZA+/g5e3lvF0G7U9D0wByuP+Dh0CzK9/GEUtKWNAWNUA6a6bikOup44KqjpcPCYxmXixE5c
4mE3rlPHp/DIQj+uiPRa/MPV73nJfn5k+UeZL37wd4c6bbtYSPWzyMSTX6eMdPU9bTQmEkeZiYS3
Rz+Vk+UA+1Defflm+7mGF++gIEWoiTIJWdB5c20W+SefARK/xZNx1qxcAexurjBmn0LJW/wPufhc
NkldInklEvsxdpai2vzUmpRxqUaZJmk2OuT+8YjiwdyQUa8/tcLHLxFnQ+rq/g11SGrKpZVcpLb1
xQKSsfpUX1cu8HXpSJ9ODCRm+gRN0K1G7w7p95VHKZGS75l4j753PYRMK1qnl9ox91g3LSx9s9sa
QA84KlpapwH+M9bnVCaxlD3y76/P55cLa6XYD2tmxgEBx7IUTDZXgAAfMrrkZdlFa3LJN0vrN2Jb
UAE5sAuC8bL62yMhfnaMc6sCMPJmONzXtAR0GT8YjBfsFfPFoRhnp61IJbL42Ibm6pnEdnDskLMA
VKj1Oi7Xhpi535r1MchKzrY8KK+1VvKQPz+gp7jpPR8M2CWp9OJ6k38EO8K+MZ6QHXsiSrg7edJ+
EIN9F3a1tgezU6fI4xlRhfVuVn97VCQAgcCqz4CxFxitTB2SFun2bNaR/5qoxnu5oIumpse8gXLa
vzkwqWXQ0M+mMcil2zhsE07YO1Pnw7Vd+6bU81X3MOomIYy6jyc4PA1RCcdu2riIP5ps22lxvQ50
gFFimvDb0zP340naasAT1haF8ILebI6F/6LgAXdmIMFDttdeyVXCn4wcdxCJxAjrZbUZPKT+1yOb
IjB3trx5QWJtzSIgecp1XmHdTPh+zr+ZjFc+FYbUiZ5ZXS+vaPAquj8F/JwCBOsp9aezRlH2YOBi
kSRUBP2+SWLUwUtIXzmzb+EPQbv4fkztWzB7rMTCWbrV9DcwTfE8uNvnmLwQTiefNFUnDbgX1LCU
gG4mEc1Y1bXv0iLAjFTKNMZPAgPJr3BSU9mFKCEc1YMFk/MjHbOB8fmF9PhIRFS4yWVwyL8WWBug
TIQgQjQm8LU6ZjxTDGyhCLsNzi5S76+eUtSWYlvpg6GMo6D1VBT/LDSAWw+1AxvYk/ZnPdUOtyPW
Fcd1pF/gsS15noI5LXpfsOZfMpf8HMScqESSm12nqSLP7D4QSXx1V/FxfiMIY+J5dEWur7yIiACz
noKZMLb/rzubuexgadL6YWQyUdlgq9Yhe2iDIjcukOSFK+8tdW75kp1vW4OPHc7o5HluyEeqG3gc
620ku3yuq7pIlxT5Np/tXBQ2shVA3N3Dt+VN1AyUnu9PcQhf9SzEyG22JWSIaOwvWM7mrYFJaU7l
3AEZ4yJSd2lYYR7vi4c8lyTC+hM/1sgiyiF/2Dwsogj+QFRj2Ib3nIQXfWGk6DBOhHJFN+O0scwY
PusdvYGQWKzxJId36XdE5bgmSHfDrzsEEhow4a2ywI+asbCunheUE0kiOjW8eGiAsGuN9oqFCLLa
crB4rj+PayP7/F8CoEfH5njYf54GSXU3MPXQSQQ0x5ZpnUc/NYH5gECS713IUmc4brIQong8Bd+T
TYQHxIg9Djvswi/KZqzLFGDXLaxDFkP919Ac9g23aJifm/ynfYDf6AoZ/GlSp72XMBTUfKrX0N5B
w4tlP5N6LnVATPH+6XvtzFJNZQFwEn1y/CbFnaR4sbYyb/NrRhUoAS95a36cbKSRD4LlaP8TEwc9
5l6gb5Oq4KvxB7QPTBBptWxcHk5b+W6SuYva7zuhwtDnSZkLi63Q5j8WqNXmZjoRo4XdfQKG0Ji2
7dbS7pN8AFFBTuaVvzhCCZZLD8xWI7Q81yXeRBnuTS8tcKH4JcwhGV5mp2ylXXFd07O+HXSLLJTM
Spk6VZWnVZXppd67RtpT3HM3ESeD2HQY6zEUFmdpl/8lrZlq0EYghvg8ysZ7lWEjQFHYtw2tVe8h
ASVd5h5FLDrN4le5nsU2dbb76Md6pusnArwnnsTscoxI9rX0FuSDEE5ybNtOnASMfLM54hqlE2g6
ZqiT4TIsi8gzWKDaN0DvpqFnFqkyb4q0GRKhxbAPZgr8VQ+fDakDQZ7X6wGZiMW4o+8XwHN485QQ
9fO3s5TpgWTFYm/h8u/As6wbvuHKqNMQjOCX+Z4QRjqmSgjG8FEoL7px1p9/k96y7C1njdxdqPk7
8nzqH11W/VXiGnrV0TtdYivW+hHIcRHCttqJy/JheKXOODmL1PHFj616Yj+OsidMltPtLKWJlNZi
HWgs3ha4fYPfVBfYS+CYHFSdcKtWx6lMDw8qtO3ukpjADW/wv9duSzeCAU0+Fxif1DK3ZaUcIHVY
XY8q1a4JSbm6Yzaq2sYO43G55Fdw7PpNl2hTOmAjD/3ifQUr7Efe+6jgBDbKU7uKKiNEjxbe53Jm
2KMAPTUllP/F9uAgFVqf4aZo53bdJL3pgFA7ZHd+h549RmtW5q1FH7jJ0Ft3H1cSMG/skGOBn9PX
lP1q0gvYpv7/+APJW3ELsS16zJqGK5hEvwEUE1UlxQpwRrzf3LJswj8mXfkxOo0N3JVkxpkYi3jE
Vj748ya2Og1teLRv+FOioWADNupdpDn1YBnxqMskZ5B/Kh6i+/9DBfBBEZ7nzyfX9DqEM6im3DCU
bM3LDOG9jiD9dnrjum5RUEPSA0SgMtmsMy5gg4kapTjqO0/mgsf433Nv5dUO+CZj0gBi+laKG2Jv
dXpioVaoyQ9Yd82qSaRTgo9fPYyboAje6o+yHBM2aKyNVtwTLHM+EB7T4+ybS1bHO0RPjcaJwyEc
n0zge4S4THjUwRRX3Fhvn54Q6cYmLXE2VrKKTeHp7jlmTUHHG3R7pm3Xd8Lsj7RrUA+iBkazmeT4
TuaJt5U4BPuutJuqbTeEmidjpQrtrxVKbZAHLScZHntG78dHfiU1OUMjfh5upE0FcTTjo6y5QsJC
QD1AoOwH4u/pOckcgN841viPLf6zcLR3LbUVviuALgIzkcE7ZEKh7GQ4SuwUJe7hE3VWUHQIjoWd
qUQIXpaYDbkdHD3YaxhKOaGWgSfHXcYh6owzc5VDD7VxvdAgtTwjNaL4j6YV4cpZdhOaVj+BBb8q
YXHvqqaI5S6ktNML45QtH5/cjmA0/8gXLg21aUpTvyTz05/shgCud1OyfuW9GI38g+HN2V90pjxo
C91TkaOA91FAwaVKMa3hEpnTSFOPK5WsXcYQuPuoxEUKkUg20e7+tYYiGzADFp9M19uuXdtCwo8P
6fzdSdFOcPuhWslMNN6PdhfF5zgdDchqPUrKciCM+hESXgjjMGpMPrO4fYVx6cTTEHUVtCvu5qeB
4Xn0xzvxVUXFgSRbEnqYepFeZJb2nc0Fnbl6eJujnAuUKM/HUR23FbCvKsQZBzMZ+LPlUm5NzsPg
YcHLwNr5+shfNkUl/mxMTqY1UWBvPEpgx5INJX/DSjVyCu58eru7qQC0M1ZawucxZLoa01AmiORG
kLivpqkaUQsafiWAWonNK3cXcgyngJ4L9h3TEscLg5cxZP8BMWGMI+p8V9pMprBGVxcfzuvkcW8p
9aBylQe1f+yReeXuLacwoh2AN1wve3WdaZGNdSs8uw7uvQMyiOn2DRFndFrocLBvJttKusMJDMbI
8JvIlbPirn6N7X3nFOT2Vm2UuxcM2vRMbDadCM/xpaXimniSJebr3CRr1sPU1GvANrAXPl7wJKhM
mjGHGekd5wKZHVQcmHYE2OmRHPXVUtdhSm6JDTE+brqZVOKSmuf6c2UrSUOf/n2IvK04K2FfXFA2
EA6KteWUAjsq1RL5h7hQ5IKeBr8WS0vkkc6bjDIrLNnS2Yh6FqqSyT0HxHjcR3ja1O9CT1KTR38L
g6YjW6/qjtPccb5F0el+v+HdAfVq0GWT4Ojtaiy7GEYwelRsv6/m87pWO42nT0uDhOeZtxKRFwoE
kt07rq5sbq9uDqXyQyWSkgIIW+TGChOIPKjbRLuzPnJt1prPShf+6KropaDHa8j6ulgx1qGBqwty
E468a5+88i1qseKPaRoUcHNk8WwnfA7bzYpKkOE1SiGDGhS3IUIyJlPYiTzAKsslGg8G33gxVuKO
w5wIIb9owXuFd6t1ejOl+P9IjMHTpfhHqSqMtxTM3hR3RshAm9WA8avviIEmCxFzQf79CG4T7KAa
7WNGuAZGtqRXBbnhTlWd3wCvFKloXsUEmTityOKJ3FPRkXERL1Drwyc+Q6mII/tmmjv5S1ZyBC96
deXVKLTHpbdv1dL2MY7KZeY2jg0qvH22uIryCPcXE9wb/qROkpMhC9m/Xt6UE95dImXQGSg8AAu7
ngn5FF2rRTTHOUM4fCewgS8+tiVCAG+upjUeb6O4ShSV0XfCqe7Ux1oeI8XH9KObuHJ5kF/ZTIHL
X+MjiXupzhqBGL/mLc4rVQPdm2vxgqZwahVtdhki9WgSnq9u+t6n0j6xS/be1ThwJO77kFMIMPk6
ouXSxw0hkZJLbznuo8H9VG2by3H26GlrbSLpKA2Sf4pE69Ovt8YPwKuCwjSJwuz8rTjmbRjBTCuI
wev5BWnw3mMhNKb4LmKNQ6V7cEyBfrEMDMhe1LTMINFqErjiP2EtE2xCVSi7wP4vfymdykKZ+ZZe
ePT//SvtNb2+I9HLJWDZx6AP1TR+HuapRhb1IYoAOzuRkbx62XJg5wbmewl3UzC3x5oE2XsK3mmR
SKExXQ3Mow5KpunOj4cAnGQW7zf08RjiAb9tHtp7CFN7WzgtuyZN0GWZpNkbZgiIJKwhvBCTwnX4
PBTqinNt2wKMecWMmAw3deUD9zyDjX5fkzznebDL/tn13hyaXiyqa+sFrVysdMgtm2h4IWghRZEQ
5c0z3/L+WnES0WuTaXV2pRXLHjQdI0PiWFxL5Fcwgc/skaKaZIdtvM7cneCeQX245NBGsSvmgNvP
IPpukuDQREMuM4CIOmQ2yI6dv2kFM0HohB4K1P7MuQgPPeVj1v4CoTuc9OPLJ55ImX6yEtHGrlp8
I0LvumEWkViZq2xkqNhA3WiCK073dlgS+pDzWLe9p0bQozPM9L97JH84KRq7zNgIA48yi6ee/FH1
YG+WEs8wI0yK4X+ef6bAY/eW0ZE3mSib2tGvCxUbo4amX4nh4IIgESdN3awnzH+bq2HZYHqWory/
3XJ0z5vhtpr72HD294KD9Azo+I57d4BaSVB4SX4ba6kZPnHXTRVzj5bYqiX6PDiu1yEbuBkOJ6EU
zirupWjpenbgNbCMEAEXPQZegjbEMc46CtaIZ090+ZQd1EuRBAKCL8gxoLOOMto9QzSGPvvHg52p
keOrsHMrJB7YV9wyet5fr++ES797/+u5jHofTWei07XnUjRyJodERz/CHwwQmwKPRAnWLlrD/hsD
ycNq+T2guwBI0EaSl5zy8ayyMJVVd4NjqSnDREuOAT1hiEXjXq7Y9qdcOQuBs7xuMegKC5IV3zM8
KNmtFiNzFBumohDdH65yyovISHtydAr46+5/y/OFc1t2No7Zqgb6eF5R5OmtOCANuWRxwzgCuXL/
HqO5gzPJlf1vG0kKlVKE31F1KUurztdAEcqVwSeODAIQUP6NnGigXAPiweUEM/NG4EUBcfAVzR74
/qC03Kg6WoWWPg3Tf1JKgnliXiI8HTMLs8o1zDWQlUGu+G8ncpRhOF02wP18Q9A92RRIpOjE2eLG
a9jWpgdSqrBUmxfnCib2o2Pc8s/eohZEySUqtixWlweI00vLNF/YJuAw2utKKRz832/S5NMpaa6h
jMeQmQmaYCjITTvx0CfalgQXPqPxNGhg0DT0fxoyoaNzBWb8JHp3a1BUGiS1TjfN3LlXsMHrTXCP
PvhF3L/RdHoPTxWefd/3TqLMqkeAeF+BzZfqg6j7ePpshQobxxGcCiduSNr9K2YOPszO/9LBSEFr
ksLCWWwLK/Pg5V7/B3mLYDTo2aHFbN5IIeWxxxUIuNyUXUw5m0JjpmnXa1I64orqWX8V0RBqP/KD
WoG4FEPtp7PjMZ320rciJ7EQB0y89lmBchuUYGJUSiwNX4x94U/mBApGFZWTWVTtjCRo2/jbUpuM
nHdkapLf0uJcMt5IkI3UtFNYbNbmnzurzKJNbMT7ocRtA4c6bGXVTJzUv8B1B4xax2l37fvCn1de
tnMcKaHt+QvdYzH5/gEfmqv+SlybK2+u5UirLegbh9IkfYGx5rMH9ADOoWsc5dsNWT6s+/6Zo1ez
hvR5iEbCocd9gq95GrgnW+6OYC8hVb/HD/WLpgW0QwrL90wSDNK8hdv0OOkaqDqHDWGiSoFy7YMT
7pjAj/PFyK/a+ZKcqmApGtZeaWtxivTlMhixGhMwFt5+V/oPCEZJQ7JADtJtig1ZfUxUIQlnJRHT
wJQEBm6r45atcqpQInGAiHKGrRadxrcNloYiIG1zLDbKRba8NhBBP+VO05O6zmrDlmbVlkGpEWxX
ICOs7wFhXvIw1wbjf/3W6hvDgjDMNfzXXtURXZ5EnEZbSkNeRcci98uXirj2hMlscUEKE3IMT0tn
pVnXfTFDCoC0uM65f94pbU+Dr1Zr7dwhGX7lQIc2Kn+CRlhLdFQnC3mEBmxiEw/QfDo8Rd60pj53
cPjR5psmFthaC0m8hdMABBEZj5jSL71s+t/2rxRceJqNPIsdlE7TgsuwSv62i2UW+vLhAw8m6RCa
UL5aTQuP+9yg5QbmnJJjckpvXoysYv8PR54kCQ5QnWIQghwMpmPB751ZLJ8/sJOEQJEYvU8/rRtx
rSKW1sxzBaxyI4BYAPrNOEOeNsThihNVtLDm2l0kxWImZFvORJIk08xMfehm3TQIKHFAOaNNTFP8
k5TtxmR4mN9Mu8e12D0jkJOoeEo8ErxB7IJ+JQ7TTxLQpHpmFvAcD2ueMOded5CdR9zUxuOIfviR
hMp0Nrd/yQTDAwKkc72ENriW/MM2EwMKOGsUkjFR87qfzDtvuUW2/Yryh+dfqd9GD9KcnkQ1oyUe
rsVoavIGsdPE6VLKxTgXEJhpDx2z42yTADtMEhIFGhXTGg1D9FRKPjOGZUxq8ITDnoElCFG+KAjZ
OSZj+GVA8Gc112f282Kc/YoP6Ws3drw1sZvocpFpsnj/A5BZXGfoB6ZxRwgzFQStqk1gWFxT2uvj
qMcNtnd7TVQBLLWxxqOkkUTdM/Vj+HmZRKLBQAbhx8XT4FLFFoKZq/KKU2MscKio/O+imlHWPSoY
knQyA0Yy5AelYGkCO3gV2iWk5hzL84vErTVZn3deXC64/f96m5dSWqZdQ6bW27jlsIees/E6RtqI
flF7QIRdryx5NSEHhYFTeuCmvaHav7VYALBa9o5UKDD8kAC20xQIJq4YmUeoKmfVefHmQ7Dlx/Cy
2II4HQ2o+kFhT6RSDwbB5FQB1/Q7f/sUC0qsDeYYudJv621PJ4VzTzw5ldpLlI6HOglD3kXDNDWF
eQ2b4jo9ex1oVYzWYsX3A2vEbxejSMDIunqWPbUuzBXL1Pmu2ZnfHaWtHOeqjefWaBmMqAXZT018
6bEUZ7wzk+MqBZNGOKEDrntZoJZsF0Eu2KGkmeZWB99o45MmOHfufkNQ9M2Sup23VDMk7cVYIVNy
KbiuImA0upEbe1oEgk14IUQENLaJxOl+JAhgLv2ZByp+aATqctatAhQTgCzGZRfAwtE5k+bcP0RD
nPLI3oD8ruU2V0PBHiNepHvoULsj8GswTJ9nnI2ZhKqDnlsXQo76yDPEx2A3rewA2OQq7bjmLGq/
15g6KTRK14b60H4H959LBnVxD+HC6IMAhzi5Wh6YhKxrBrFWVY11gVAYwJnkmjVGiQay4IOR87zT
rJZH14lztO4Za82Q64dBAzK3R+xjjbn/ewOAGzZNHwSG4tjmK1986nfbpvtBc0oEjMrfLa5HXgvJ
0jdxrv4+dzBgrIQPUUnp/kssmwOe9qUsRYX7ZzLB5frDildKEXBLptExMj46GPhA8LDTItUbFP2F
EpYYCH1YV2IugfPJ1EmKKyQDdEYh15PK5VMDmvNyO8vu1Z8RC+HiJ7o31nIE78thKOz+xsiioFeI
O1XIHPYc/kz8cMTFEt4Cc39rprFyUnWtWl2e7KGmgg7JaHn4GIVH0HEfmj8mh9bRhFuNZN3+Vl80
tZKkYQkQ5d7LjTXr42LhiER8btxZZqBsXD6a5mLDAvGGy+xV/nwA+XJK1zZrgesZPElrUWvAffM1
hc7xHMUqACNRiD04z8Kpg9sfVrE+YERxLObuzPzXZXGYZ8wOi2bDQAbM05d13myJTn9KI9oExIm+
1wYx8MgBPMjQlCt/UDs5RS+BOI5pkEscPb1+Vc3GAMlymFwqzqLpu5RD2qjd6OJjedZNCq/RIhFV
BelEsXeDRXZ9I9w0uxbJX3+iSkSs0txKmUXXod5suviuPz4dXHgVvKhUrt4uyrCQ6QLwwwP67erl
OHNLUXvV/wGEN4V0BtsFkStqZl5WzrdV2WZpQg5Twgr7oF0Jruu5LOyov4mrtah6N8IWASfn73dO
YRgdJ2ZdjlSMkeD5cPB+R8YSmN04F9tOH7waeidmgKV1w7q9XUR2qCnGf1UMe3y/28G3rCIjyPxA
YlA6RfBbF8Xbda0YlZ70JDg2qUvqfJ2lNo3fngB30OnRrse83GGEMJG9o9ovv2pbS9iz4LL/vHg2
ZpHRLSFh2M47assyjKu4BV9kpkL2nVt+3gbUcLrsx48lZTZmA9SpwB9QQ9D0QF6pDiogN5Cn4lLo
hfKmEgmCVlfWX4LZvQTFeaqxPvnMzjq/z0ILuTEbXapkGW882u1+4VNd2F2mu3aNOHWyq5bE62KL
uYMv/0F0NKHY2nhZ5ShlsOqxTNiURzIbxVQaELOTMqornFkLHCNPhMVSIfdEXdF/tqd/VA5Uyhhc
9AyTyR0ADLujiFhJ0Mqym0eWagfPLoFPReVf9Sut0L1bBEFv4hgzBIufUy2d8VXoJfGGX0q2q1re
YuNY0zyecUzr9JV7WCYZqIB0QsrA5WLnbxUatzPtwFVM49ZNLDJumn/7+TxHA4WclT17M12bZI4G
XAJSBz6ULJLgQl/FgKX516QrY7SR03OBZn+gb967TrD1Zh0QBEuDxlPdw9dnTDcEXPMt2EVcIejT
RBnLA74zS0YEUCJ9stuzoU5MowUC2Qh25NNO74yK5i0G/wVktOaE/xnnufOKU9/E9KNGwfk9mIGl
8TU6jG36oZwFy/OyZcRt9uYCthrY2ilYUB0uZTbsKx5MwkdNMIWlDLmGQGBgs+89hAJ7doNdjLbK
V/u6sNMYCvqTB99nL/gBFNSJ0uvGi5p12gRUkxgpLjzHiXJwm8AkbWmpHNzhTDo6bz8vcRPhoNsK
m2PvPI1JvtjLpeT6xfTFoI/IeI3J3kOAzh1r5m8Vk7neSy04Rpa8N0RLJB8g/VquzgIu2qOZvLwu
3rR+3Lq49Vo78pSJzEeeeXX5PPKooXjhi1qe1WGwTCs71W2q2jTd/TzPDkyKXRI8yRdRDGZ1XSYs
7KZEI+QPPuh/7zCWR52WFABlbSwqyUwUI49lj6IxX+Xhmucd/CkNfIyt50f0K7D1GbbNE9U+d5a3
1Q7A9sklekZStIhbpz+KuzYhVsBQg4A6VLBjmwz+qoWDO99A1BMk3LmjawXCqU6BsNx38kUbKe5b
ZS/nkDZCvEH/rjRTlv4IVZSa5yyW8LRvJGS3+4eZSL6nuhg92k8FYPnxRZB3fZ6VS5AvNMA3E5yy
z6sEEBd6Sv9//3hDD8E1urMPg3evUyuS5lj6IvCJZVQPFhnoZ8WNirZoAmjjXpyIrzoExbZbCJf+
ZStbAV+ol3JLk13x3DkXCbJ0xOusC6JkuRxG6sjqlOcTipziCiHn6EIPQVJWLsIwXRZLxAMJRUKK
El/0WrWJnpqY4ViL2qVQ+EJAVPhdaIbIwMsxQ4/dhpKvXu7uWlCYOKkiWcun8OwEmxrnMqg1dVqF
d97jFyKQv+lsVWDmAWfJlyOP5qGXUZRNXSisHrKU2wmfLGdF/kX1McMz6RISm+HVI/dr9C959i3X
V55omkcURHrORrewtUsWVhKSw0QjmHwKVqBMYjiEP4AjQmIa0SFWj6otQNMAbU2N9nPzKUDoaHRj
DLoQLyILFNif7DxSK70MXTKxoEQGAbt71YTPQ+CMSS4DR4Ubtg4h5MDsdtnvhTEi3isF9Tn1/lHy
A4Xp7Wbco9fFV4VelLkyZ08n/zibSorw9Y7T1rfecDXD/Kzb7Fdxh4npAP0oWxuLcOG7Q1WmuVIK
YT4oX8TqA+c3OfBZaddJ8wV4tMYNtAbDe4HnGvUBtU3plbU+d5/aBd1KmVPqzvAHza7VJHRDIoIm
w98q0CzXmea98keFVP2x40aHi8NRgPjJpK0Kki+JR4sZldJEzCr55nY/HWU5isVLG4N9d6YNYaF0
0k1V5rx2MtNrLzdGViS6ywv9u/I6NCo3KQ4tkH1pBt4vvT52UXWSLBTkfYjWOKbZFYg6AzgaxnEF
Hgq1de6T7IxfF2c9IXpuk6KfYN2Ks3W4WRxNOERUdd0qHybwR4Fml4GMf6e2zOH4qiivlPBPzO5p
08it7lz56LC+i3LJVHEiz+3rn48AWwWfJyhhYGZGo4aLptKxuONS5X/NgUjrTz3a32yCm/KAKnWm
USWOjAFpVhcsM7NHEg973MTNM/Z9QdIpK94pblJfunimOZGmQoybnEZpqHaZVv3f/8SoklV0hkRc
7JlFrd6dzdcMlYuIEmN/BWPkGeHjZE3sjrko3aOrxkXytfVlvJc+3+PMy30bKoOpjGKQIQitR2Jg
uyIfrEpW0/D2mSnxZQgI1BD08fHA4LioXr/Nhs8W8hkn1h8pkMisyprGpbEhQyymxUeM8lAlGdpW
D0G3PH5Eto+2aECid16msz6hyFc+zmB9bP4UVBym3+79/ifYScQSbdepyeyd3CxmJ6ghbqWItStM
UYRayLV8hld6P6YU8SGmWfmJ298ZaspSDxSGKWVNZlFc9gEqhX2p2+tm3SwD9ukgv6BxAC4bYR6A
d81BwSnfCc+x7G0u3Cx0B8GiEKR2NwWK+xANT5kp7MbwRd+3+5QgenFi7RvMaJbBHdwU8eu2oJ1p
Flo4m1pZZwXgjTJ8lilb36qyz/lTUY+OtkG/K/4GcWdKOXV+HBfqaqGorXy6fFYauDIrXNttJyPc
wk4IJi8hXI6iqxylA/KDWrZxDZaXRInILEhd8WuTAUPKYIrzc5EnNKalryfbBRAcNMgKs5EWOpn8
Atgc93YMQqIhtphw8sukIHtUVLCxiLMz0Apol0YKaSBWNAEderXmJlbevAMnHrzMWAn0gimhCJqQ
F28gewiBKA9KdA54OqIFfsrdHBP1loXV2p4e3KpjpJm1kZY/4o6S1IaNibFG2Ztns/SXnvYSktQJ
O8Ti+Sieg6aq8smCzAoE/j7IsnufUNGRNZ/6qSAJzGWrsiPnUq3GYTEP001iAg0xMHwJx9Z1V82S
Z40rIeoNX77i9QJ63uG8rivzH+h5LDy7jbOjvaDKYov+QZ6vknZFzl9OYgPq7LiMRfp7QNzBpG5I
bISci7sgScryomQTcu8yAl+AWD8ca7qSGIDilnVEVpiPDXCc+qcdtYstxusuCM+Oo/3Ur0g7W41s
8rChSIhQuhLGk6IdEQzFkJF4u53PuUoB/LSRE6Ldv69FfWAnrZkWq9T1c35M1ceagEmwfQBP5ioh
5AevU+mtrkzV/m1IC2hkA2sZ5XWhDl7FOxKf5wObqJuyLIxzN3zCnFEo+6evJwlK57aLhW6sVBOr
9vSDy5gDi9hHhUSlYKGas2L69esc8AaI3SsIjbZsE9iNNZm/c52Sd+OGajN2a/Z/ZVij0B8G4SDM
TOz9Vls8NNzrC79RiE85WBPVMvv/RgbSMl/myAF9VTJ9q353A6yXYQSRRbSZBkEIomWTf2zsTQRg
OIrJrBGxqzNcQQKkDx92zw6XY09jmGMH8QE8e7yoImIrWlvHno99Yaz58FhdUDUnZMIoeKKarT0j
2DrBxnOeqW1dvI9O7IdQQRQPnUEaaCKRxFcCqv/54k9jTAVA9iPA29nxXX8JQph8me0d7YC6moWw
znkMv80K6aj4mrMaLL4SlsLFL9zWvYS0temdyTvt13XupEnsCQvNbSykFShq2h6v5/0B8PmsM5FO
jdzDkSAC/DDq8v5om5Na7F/l7XcxXgxQZNaIPOuHAmF/xvw6A9pme/XqVwl6+pE1lhGW1sHQkubV
mmUuEV/eYOJ88JFakfXBkkDAzWZhm8bdDVBlIThUvKbPO2JwpxuDNFQs3hLl7z8mNtMOqP2zs89/
HPUSIhVyEb2pRpDDdekcKEhjRJjVRqLQGJLXw8QR5o9NUMtllCxMGWaw+OsQQSwYd25eWilXvmKC
JlYXs/vUnVDnmTte7nOde+anZC6avz6DuVQ0W4d5f7UQuvy5LKPWgIwXyjVcURMZZJuOVLV8anD9
Mjtmoa+0hZDUdXzsPal0WdulnAEZ3o2YFhkX+YS/IenE5+ZLD4QskBusgF/C6Ny0ml7iDOXLaLzj
M0wu3xV8IC7zAJOr1bxvTl3Gkd5pczcygqX+0XB1prU6BdeRPLWvua3kjVsCBqHrIsyH3xkRE2A+
UaWKZPg+rbIehMraIADwxjae/rOaAXhSorTa/HLx4Oh5MR7o8B3Szj9cOBYP8I5mw/YA7gYL8wSo
pHmDJ/eIICq2Ph0SA/F/2GV80Wrl2KICyZKsGFNix0GMKeRrSmZW+3MDanWlBGROTt34K83foXi1
NoBaZ3CpP3GJ9TLzEMm3syX/5cOyhjQouuyiGjY/tsDYcReigzS6S8fX2S46JUISS9DkHlqD/q6j
oU2P+55RDqOARZnuyW5FU4q9R5qWD4Y08SfPI121fHrQ2ZFjyDvqbjsiHwkakfziU8q6YETXne/w
xNI3Puq+sHb90C5NPPGEnaOZieYCVUZoYT2ZD7Iu8KFD8lk10bXhOXhBuFt19i2rKGMf8uxgnEV2
V8UJFwEt3nRwZU3gm1IKyxXx3TTGLxED4EAeT2fj3NbATwlo/ad/Lu4o/Jb7I92Jw/HasG6xjidq
TZ4NXn/VFzPzIQW5bQ7a07LDx3/E4ksdoklw0tTkpSSsKezm0UZvCCbtTBKQyWT6Z/eBTc/w9uMw
kIKi3WfUKaXKOYBdBYh/3AJqI7gxNszt77G9rU5pxm8Vhpf0vrs2J/6NY1vx4hgv8KjVpbmBFL2n
T8YluA1+nmB308y+TDdJ18Mue5kApGKuZKhCMmPl2LOyn5IgphrTz5izIe9MWjH0Ha5JvD0d2GaJ
qIE5eAc+3haV+Aisre9o7inP3JHUrAAwKXp+gEgUVbLsk0nq7XWEJEv1vowzoM9V5J5s4Iy2QhY1
TkPVMDPkZTgqrz7z4xUSsTwrS829BCeYPOF9iyvaV1CZc3fovgt6rVVGVDH6ldaJl7PjEcIRjgS2
+FVYDycWodczHsnFV6GJIzZg/PeBd9qfbgJ27iGRFm7RXNN6wDGfsdzT7IXK8sIVJBfEXqcHNxr6
z650w5D9RA4dI8BS8CEtwoskrn0ZWM3FlYuIQdI/94qlRhwc40AYwn3EGpmmLt0wEPAWMFrfze40
2xXjS+uG7Lb4ru/KrEZEW/9184LXFGrp0YPR5TQ94eJXDBvsOWqYfR12kkY6g4dGrVID5D8u0qhO
yoKKh/5KT/O9xZi8azARoPCzWwq3/8uy2phbv7vXf8BLSrAuhFN1dJuRBo4Ghh0OViFqtTAiQO2T
/tjbbXsUjC6Uy6RL6OVsppGXK9y78B1XEFaTS2IUZA+Ay9dJebH1BMemf0pUfqHLNZmKshkBCsS0
ft7uzGID0bljiTSimaiRrpH7Ref7qNWAXQFeN03BtfqMx87gKk0AEuSTScRQYPzpqC6y58jrtEzh
wY32t1l+sxuc+5V5xnwbfie4BKMqeQFigBdtdhhsDn5fwkBSb7Go3OPXSnnQICqNa9I3Xbcpy83V
QlKGF3nd003Ux8lI9YNFl60Z9LHoGySWN0wyYjwI6ehzWozvijFEEmupbiZYnfq3+jqEAjFP9t3E
TZePvrJY6/Ebd30Fnv09ou2BmnpSDntX6w3KcmRwv1jU9m0FeE5UxltrfVQA4/NGSFVZRz9P1BCi
sN3ds1WEzG5jxJ1EgfzjVNB6j2NWL/ZXkRjNdV4sikHO1hB//n1b1N0M70DATgyOxGXrV45eyjKK
otRLYu1SzEDFxxgnAWV6j0eR5k5zrqEKliH85vVSZjiyCtiXngFYVVmXckqSlraXpfJD+ySWKT3D
7bSpEuJCKkYrC0/pzuXqy5cWTl20XY5loo3Cove/6cc/na8WiE/6Fm/9Yo5IJp1M47Ao1bmjDm27
e1NR2mv2lvC92qjRnV7M2RleODRq+tLjQ27NlP74Dn4L1M5POiX3zBrUaEkKwTzs8GjZxJIkdm/0
Td9Ts5sXOja8093bSCdWdGmIzfOqH+woWv3Gh6Hgq0pHOwTWPatu3DyDvzBzIOQb4hp+ZogLvSVd
JAfebiAu65OsZ0spmPbu3kCREMFavmbjiww1H08R/vQiChMDNpbbNiviwTc0SRvOXeZksCkoXqni
tqMBtRZ8+XJWUDMaODy/YOaCHoa+WKt0796D/uCY8VImk+FTMuzojiAG6sEKTHQwb6XffdzyZr1D
Cckd/zuEngPqNcj8+aAmUEp9QYHoSSGLzcxsynNcy3C/UWZnFOdUUmQJjVb9IWwEiuIIp8mgUb51
BY+hphiKJxoPp/m3l1UF6BgtIB1Ylc55NzF+A+qjBawC+Nt17TPu5+/wme93QlEdLUFyoFmO3iiC
KZEYL1bC7+4i+wxoH2EKVmLERdKwOLrlkkoGJ7vaLw9jCCIR2IId3Y+kDBvwkqu+IeS2GHE9O0sb
WevDT1N/qGQs+UIn2mVa3hSlK31hsd9D0gozNu9uFSjfTvJ/UjsNE86wQSgizGrB/ePKopWn33DB
lA9ryTm+6nl2PyantgryiLppDHkWeZo1UZX9NUozwOz2hUp1pOIfD+ICBxpClj9ChXcEIxNBElUl
YTERP6MtB2GdmMpvec1M+HPIo1RlId6ehHCnU9uxMuzYo3gGiECmeEHuLaio/PZyLEva7Es3mOOk
pfmpsNqs/36IyhoQ3G8D5kWeqq7nbA8a0QMc7Y4RS6AfuUvyz7iqxwCU3+VgRRvb+R3qtqCpfTL9
ZLNQyUw0boauIpGGRVsE8NLKQCB5D9ntqIMF+Eq9EZOOjp0wVtkacxeg/f2J97lEvWfEwX+y5Uh6
dZJRz1N1rI7bPyCqCkgU56VZVWUfHrVfr0B+7AMb2XZ6kwL2MSpl5m4eTZNMyF568Zpas70+PTSU
lBv8w9KVtk77kcihrQUj3tq4sZGFaZ8y8NOY7pNc/DpZ02GdHvh9oRwvSqZhmJUgGCFerq2ERnZ5
I5YwAM+xtcgpF5nqLQngtM19ZZg2tLLmPH8j1eq0do5okR7vzxD4Y5rBUmbZkRR4tI6fI0jGWW+r
2Ed2ugdYYYSHo/GDwm5rgO9hSG/LTk81JFj4ISR3s04uxEt7e9yqR07JTtrplrlZ58b6gB1akGhK
ypVUd+p2SxS0G/GRtnAdkGTg1lDr9g005NtxBZfbenD5BXWwdwKAD3TZbMKhkXl0xBB+SEFD52ax
U5hhIxKR7lYfMy9A3qvNA98Yzx4SfZXdm4bD6lW2gJYzkbO+TYZdgX+EbEIT7J0JFVuEsA4ys7g+
gj02y9KBr2Sx6Hk4Am5Et769vwhhZyV3X0BnRX3oQMwAJk6y39zlOmY3MH1NjL+mSAz4tR/+KlSF
92kXOZu7G5GaCrKeeEc7RoXDA2+LGlBMi3Q/rjWdPwl0qydN0fCnqZZr/SEvUpVN7TPmZhWW9j1b
BJ4ziKvpTWv4jO9X/ejk4UQ711i9F2pHnaKrI4gKgLgCCMAhcUa2jKMmMjZ0916zbzcLhDfIpJfh
EBFIvgAvFU4TYAR2yUQzpEA6T5+AlWvfMaYnHVGxzhMfF/MGW31AZiHBRNd2CKFS6Yh6O7FWYGbf
APhHA8o4WwXLRouIchA6VtEWf7n4lIyGM2SGhNqisfhNjvGxeJhxO1Vo1Lo9ajHTnn8H9jJGtxhZ
nIbRQmuyylGY2J4MySi9kFkgDJpWCQb3G8mFHKgA3mgVnW2rJlBK7PrJtR+dCzkklt6V/shZstQU
g0n3mi7TXi7AewaOX/u8+aalItAHKTF6Au/l7Uhq4apM8dFuK+1lun65tl77JExDu4PlA2SnGo/+
OLivHJSTSN0u/bCmz0PCYbND1E44YbZhG8jCXpAPtTV+dtXfWVQZ1z/nqtmqLQo3YQ9pJC0DfnQe
i3KHXzpABoZU/9cDE4qYOeI0Qk6u2H3ulM7+GDmbDFwOMO9wdyVztMpSqb7nx/9Nv65dU6NFAzla
GDB1eN0c+05Q1VY8cVju1Zxbnsnr5GlMxZNuQDO+0BSezV7c0TdezAEHErdh4CgnWfpNUWJ+iCUF
8N8wWVnyFO+itm+pPwXeEBsI49mTjzvqRSK88ul9rYZYDRQag02XNxPfMcjazT2yPHDk0UgXMAqq
AzF0Va1fF0BFGAL1gcpLGDtG+BgXBE8PR7Micf8R36C5UJ7xw/ij/97Xx9RHpCSvmyArXMvDnRLv
Yf1PT/n4h3YT/Mcn2XubxcojFl0DUlqDVcvpRma0D1gGRzROHyhwRZ+QfYPRp3WqYDdos9TArSX5
UqpS7oXICNH5H850gaRsCGYmnqk3Ns23UNInYro7h8htVzburmOoTP9fv6NdY1PM07wGmUQ9OL35
DOPpEvs5qVkgsHW3DQYT2gQi046NkJs5PY3iUh6WxgKfTNmQg6odcgBSHMfobaz7vFDt9sR8w05F
l5RBh8zM7Q9rJjHKwmNzp5cWnzEy7RDmxnFgmOsbnKLEUhRMY5tMtsYRtpBj1LGHe1tRPaUkgMdQ
sKnFwMXSw6rdjgLGO6XXxdsICI+9WzS2jLTO8X2TrGFg8rZ59LTEkJU3+sHxZvzeHZaNJPRdoN0r
8P653t7DUWfzVLPG9aUFG85MKMCXb93bjJEWFBoN2NcmQ3+QsO4bCy0rmTUjOqFTX20zIP+R+D8k
Iw83579cheCu/o3EFa5uo513Pb+QgvN1iUjyn8vmXrZx20GgAvxE29weDkl7j38dqcuHvy8gJ2nm
K4lQwYXAsxcTblA/AOhZmIpjWDcQDtQ+UjAQBi6UMwjqZG28I3rh71Xt+KOHT6yHvHwHTOLnxzoJ
eRmNG6U32/NdGrgkN0bqYWM4TNbURu6/phCOP1TLUcixmBczJH6eONjw8gy64FOroi16m796KuU+
wUdpp9OJQHmuIuIn26NnrNRjdDE7wSUZ9vXo2eHIUVWiBCDjR3ya3/m2KTAy5ri46U9IZOcmK/Gb
PwVMMfElzV1pFTDkLdlOb6LbxOH9U4k3ydz3FwXlMJSGGQmNSQZcAJhTUm7eM0J1+It6uXShqLQk
XeVcNL1PCkp01IyBKC0CTNJiy2z25gSJDqCMpCGoSRkOIcMvnDrI166VQGuDARiw/Sepo9OvsEGW
dDv1Bp0PRJftq4ub+/VNn8ZjphvQVoCkRZ9JM89GvBKtdqT6JerJVHUxqu0bhR7GIqdUT10fEcKF
E++s9uEAGvQ1IAnjNt3kqD0hoQmf4a6yukex4VSIkIHuNLl5+R/y/8NT/JETKH8WP7LVspc0AxJE
CrbXs9vNL19PJQwaS156B9TKyo8D7cRKHFXgplTuJsCjgRMQEc7N8IpBM2aFugSPIAh8XH8lesNL
HCdq15q/XY69H+IxN/o7ewdet4fqdoNEGj4V1TV3k7c9OKQWq3F6OUqPVcnq8DT4XUJ2daxzPNi1
dxpstjEvt1IP4r18SEKaHECCs8NhhQduZ63hKkmLaTfqaHAFpCESgIzlw35K7FGSYPQDiUeBzyHu
UwbEb2CAO3ziNnuw19k/zk4p6Ws+zo67zHM81RfiUQjIgoqOXJSEkEoN4xbc/X+Ql6A3966Vxpx3
z4QSbK0qKMljxYpYRiHH3Ef07Y/RCa9nJfgg4m6Ubu9iNYkP8YRiUaaufyUFw5JlYLo6udfEsVnM
oFV+H/fl+pjtiF2/aqWTKBhDt1Zwbuyo6kR7+r0SLJjzCtDXcSZDAcXewMPJIttUWq9sY4kbPUxM
4YSe2QVNM9ajWaxwtPdOCgcuRIHy5LIes5J+/N86ty4Jj/Aq0MQ76TGSqyJeXmoL2dFOP+ibXI25
968eAdDDT7BxKMBKYtXI1PQZN9OaXZl+wUkQq1dDwsUG942+tC5vKiaeXhPP1qfIyi6JecH4yah3
OpUn2VQ7G8azxFWTBtQp+Bzie0rhRpNKhT9w6vJlw+DqMXuHYbRQHiR5f89O+wn2YzZCrf2IDD0G
tAKzHU+HqLHwv45TqdNMsAwsG2siznX+PmbXTGnT4/Hc39nPdJPLUYlXgJUULB2WrlQccfcUwRWp
A6XyFI8NIZZJCfNQuP8158cEG+BkpqznmZQHaFiz1pFS9+KCp6tdZZEtUfyqb4JHFMc4BjOrG+Gb
K8BwqRmey6U5ezzANMHXt7rezf2kxwHYFIzatrRP3vaDkbRf2Xjy2DphjA76lAD8t9q6pjHZNgMP
wPoZ2d5cJAwujw8v8PV0L94BTQBslO4iQGum4+huBQrZCIHgVWrVcV8sPqgsJ0Oz7XgiUsPJ2+zZ
B/6sb2Bb2Mm5SmN6qhBGxWSFmgbX5dDJoVsJWioeI1gonDGieju7/CrAmwkK2UAESdaPNDLGpZuq
XndTID+BfhSHDgp8fhuqt6h65Pe0p+jT45fltH4e7m5VBmdXR4pdh3IGRDG3jnrAEWJrgFpatj2J
r6pu0BRHbHTYt1D5AIXDIwaO3yrYZEYNHDgp7B0H9BElmvDzqIp4tuA5eal/P+EF1Rg2bcbfu6Ge
BUP3l0iZLSwrmlfhujgN+6VwVjp/HtWD6GbOLR4AEfRTAmenDwSA8kYFsEe7XuSKWL/vlesuVq95
YQRpUtL6nMSsP+R3iWz497L/zfs/do7w/k1D2GXFdlknk6JOv9CxvCEhcQXBKbSjO8DxbU9rv79X
EpGpYDkYOBBjxPlZ7Q8G0UxQlzz8vByq2JIquwi2Tjj+ocyd3RZ2pE1Bx987R9q2XurmJGplDmmn
rWbe8dhF2eDOkpDvglM7KAn7y4Wr0adq4jdiTj/Z20nlWSGE4rE0SFKjKc/9Y3oVl5XRdqy20Ya2
wO2Ajr29DqcBLs8IgoZdXJSy/kCcoFaYXByDQA4uv8V38mQ08EMHU0gVAVqhhtj4yB8vqLie/qnt
HqCKIvBeR1vXBAp1zISjF+geljlU6h4fGXuuVOixlaxhBatixf/9eBMSb1uuIYh/QeBnIXCneq5z
P/Y8b7o4oBemQOvpvzYn7y3PK/XaTcvYAuKNMQgE2WHZXfaIG9d4yXXl9lLDkVyDbBs/Dae6aeoq
PHfjCE0511XExAgrNMfNLTxoRBkDubbl6uPWK7JamptgKXiwNv+TbbZuoN991jO+El+aKC5XDzRL
82Z36wPGPv4q1+/rJ73IkG/eIn0zghrrygR/UNenRFdfT+FoU0avH3Kz1Stl6DK53oKsYSlB7PeF
wFbUFI/BPZrp+XEArvAlQOio7Ds4TnNiVddY2oZ3WHJYIG/cJUqEOgf9MI0YfFCIVs6frjHbXAKq
doh2uIkPmJf1xbb9DjO8dhhWM+13KqFFAINmw2yWE+BrQsaaKD5f8xay5bwQf7RfU/wwo96sjZPb
zzd0CQomR9+J0r0p/qxs56kGEczN9yOjHPNdOxQeh/htvp3XUzDJVWZ30xrPjSTFmJJKCBViFvK8
Ws4/v38WxJCYE55yz44EXW6xx1PyzE37SD739yWD4Ad+MF0iLHACP9eP5tnkySQgD28pRlGo8gkL
6hMIy7LZ0Q4Sae4p1RvWzPdDQAJhhX2JYJOYVKEM5qoS/JrxbxTQUuSytPmBjrsZgaUjLaqKY0Tg
x9yJbtEuvSKEQKP2COMfc4zp0yvXqRdDwH/BjKPnhkDHv3KemdZJvjWZx4ZDzNVwWqtKJ06gOJJp
BOstTkzKTGgfFcihPD1FPhsgfUxToQ6SBuEJKqvF8NKz8xSFfJDaBK6k5cdSUWsbEIXSBFdKJ5tH
ad5nk/m6ACrrW0kfsT0uTkdJ8fOhtEyR1QCBIiGh8MG58kIvJJesZ78hP14B4bjdDG5seRvfBMir
jwRkym8laX4ONrD7eo5mZw6HKmL4HeTXO/BVdzKn6kkuQMchsTvs7UepAzSo5Qb1gyPex2V2xhAU
iCOXZAb8va/Q+ahSYxU8e3tuCF4WGA3x4ZPvifes4Fsk58rsvigo0bZ3lcnFJIYJOiwiVBeRs6xi
GSwaSu2vwWz4E3lcZh7NGcog7kzm4SAwEhX1cS+EZ1MGTGtB91Bs3qwcUtT3SYcmc5q1VQbJJvB/
DMb/7pPN+fIkLO77WynPRRkYe0mEYTDDrsx/t0sH2aXaQ2L/VoT/vwMnM5fleRHrRXxGGmq8Jr04
LuSKU5mka8DhX88v7yGxYwGqR2aztjIumUPZbRjQQ6JxoTqhjWh0DHglCBBYulvkeSSSLhLo12Rf
5z59gj2CvRC2HqiuaRKi6Ok3ZcUPzNB06IHJjxqxG/XunWfPTjhAVTy7691NApIWgtuzPrJsdkqZ
s9XZIK9EA+fyPNuV9Dl2GfAYoqbDF0w+CjYf3HRF0kC697B+IMjScCziNzYONB9ZIZejiMtOsaRG
0lM6t/u+JA3t3KeoSkKIGXXV67B07QYnUPkxfM/YoUWg+UDXAE8CUgc+LUnYd4PcU3YFiXM/w8xD
3xHoPhihPZq93U31GEVpnKCTSuml2XBijiYIhJx90YWzu9+/fVsnJCuS//PcVwAT4yhi9TbYJbyK
jiG46Op6wOc40WOw/53dK4K22ZxSnBJMXWNiXT+XrUPsfo165CBHnwuUVIDIK8sV4bU1L6KRUPw9
GC2DNfSd/pL790azLJIOqoBA9F1Mj68ssRJtpW48Nwsex2/jmeJ8OkkbX0t+3VZzHBLfUuPh9eJG
OezhWHK9dxHWROU6MLupmA90139ztOwCwg/rsP2AENcgiN2JoDsE4ZnxBz5uNUfR0mIIQy+TN+nK
KwKU2BDAAlR2+uYaJoi70vyEMILyewCB0MWLiAetwD+A7bIK6uVNC9ylTslNqRbvKF39vbc73XmR
JTNIYm5RygUIMNkr1KnVCiDnpXGvZjOmLNvQpdVcvaczblIUjun8EyfwmIUWOZfS+CKqgWhotVJX
kulZ+MTzSLm1WHR914T5riN87/lCAksnLElby226Nbz95vO1DmJ5BwsLiGQ2RJ3kKUtsqCx9v+kP
BPLFCPI2fXuJGAnPvd+ExcEseSq8iZ4b4/ewiEGDahqML97E11Mfl0OlooXcPTMme2HZbZBl56NW
9FaKKG+HmINu7Dkcp/BSD0XzGBjMXQn2AAGn+U1o8npdWwBPsqrfjmmoVUdiAW3oHEuBs/2ADpUt
TQasVWKnXZkIbbYHNLMBXuRmsxgF90ftXHQuduhXSgbjGqsPlhAWzawjxjN6HUlyUXbIB39eavHA
LC4EYrUmQIgbjzkcrOuaSRM/MW67OWIcGPKobQ4oCpJLo43jhi4hjS6jIlYJ3ZY8bOE51PUQQnFV
4sHKlNlss557jfaDBCYwDDOVeSvuZQTJNLNafKXRUdQeLRdXTwTTrv2Q76I/X9S29FkBnBKSKcW5
kb0qrwJUu/r023g2fBtuS5JTDn3ZFjPRnClEoKlWef6ufczLPjpY8+fm6CCfU/Z7gSsKi1r7Jhzb
p1Lj6U5mepHvmOJ7bNdKAIRbOlEk+wB60mDcXQvLdQtR3EjQVmL36FeHDcwF0akmHvkSiksLRaSV
K7lJR2dmlyYN6ojhmC81BicZidWrUndtu+lCai8NEGQMQ9OEFADUHx23SGIBe8gAJz8WU2yWg4P3
EYAIvpkx4qDlw6f5XTQV6tC8B+fyzQ885JttZLxgljTtAFVRcJ1r5ivUJpsMFwe5UNTV5z1zFgQv
asBP2Z6Klk/hOnXL/70CRmFKdTOlD+JhA6snjBnW0FwOJHKasBYTZ0axzsRntchW4eeaDestHW7U
1jy9hB15XcfJcAbcv6aCxR16waF0Rtvrh347svNthxbC3dJVQV8kK3EiNXPGY4hGh7Db+aL2ZwBj
liwIzabmIryPxNY403UX348j/hx74OUe4PgEJZbX+fGtqfqeknd5g83b80N9IPGmj803FDw+dcHt
lzKPtPBJVfCqCWhRvswkGKmA4ny3Lb1mFJxbrJ1t9emdzuqsLK/MAXCVNWyK5Xeqv0llmk/qVNV5
Hp4ZgPGii9HMXR4E4CCl8u6CFl8VWr7jXbeJHK1Y3QV6iYVg61LdFI5iDprDUO+fEtKRmMWF0fIn
Y05cFhdoGtb7insLnRn8EQRxLNx2ggY6AKEKhPnSrCFMU7+898xerXHkogPWKpiaDREYGx4Lqe85
O0EdthWbDlJXu32OJkfUhV66THiXyENfhkFblbCukA3rfCv/6/JFKZpGy0LmabLo4V5jD/3qAePr
aFmg+1od1GlWMaPnWtRGxnMS+Z9M7GTR9oPVYtGzwIBFvgMQdp4fnHRpDZ220kNGY7MDQoM8VX8B
mCryiRRyFU+OVl2Fuu6+2+yszBzcJH+4vWntIJtd4j/7/aQeVkPk4+Dr6YHzMrjYUrVX+BeKeIQe
qoVUvKc0jahvXkdwa7tXUsZeqBYDRGfLPa5/zyNZZlNVWKhJRZjEs8d0BATVartw5ZgULIMRVXEt
Jh1dtmuh0X1vxogZ5eQX4H7cRDZSEcqJWJtI5SBxgeVnamWb98Pxw91mt63yq/LbwNs8jH95RQRt
jfvSspuiwH38aEEG/bG9K7CKmNrg2jK5sW8t7vZAxG7q9+oWD7orRMnJ67AUmdnLiNNzuzIDhzeW
bH08F88Y3rP5OYVk9phDMhG5VxrVA6GENOeOb9ZjWAWM7YXLKmnTdtPj9Zb1l24kFnh+f4dLYXkS
MG8vF2xxGNCY2ntX3GxV8fwKZVd214P0hmginsaRShfRijjI8Iwj+n1Wcn2hzB1SDedrFdsariz6
oC7UaJr1vXOG57MT6j/z7wNx8lrc4QKh18+5goQuJEd3FObeVB3r/lnEA0LrCiS3jLQP8LjyzkCb
QFJYSjszjkg0t8lBRLszXF+2bkoYG4MRSkWzmyrxo52P9W8t5M7SKMEtRITqEm4+5Rcxo9Ps7mvH
XtNV8RiB5jldByNLuYWJo9j+kEMDIQCK0aQAcLpRX/9dKgLhuNZxLYy03EBFnM7M+ue5HEsBJSSp
S29UQmAsIOs1pzrzPXz+UjT4IgtEkbWL7FmsJ/OeqFtuFvX2Ed2xF7qTIanTTf7AcZK59PJVkZ4n
N20kmRLAKkXHPiskkdeJmjPYa/KdN/27uVQ3JoJmmEY7PxvjX1Ce8C0QmuHni6GvOI5EMbjfVqUP
lLJHpR+nS5N3r7YcnoARMD7fzbpWSFFqQPsq++EA4Om5aiRDG2Jw5pheGeIJDB8PMjRDLkKw10yO
5LdCZOAAEEBUjK+7QGVrscxazuwQuokGIXsX8KpOSSixQd2p1RlFfGHRIhplQ4iYnH4v1w5SKBxv
YV/+NqM4cSljAvIhriWyXYYCMjXH4MdUUpOBHo/fRiGVwGqEoCmxVv3HESJjnnLLSpgzoY+n4Oov
kdKYNZ8grySNRyw2koRpRP+o6VuaVZm3VZ68WXfbJxya6SFXfqPrcDVWacS1Suk+YV5q5W3WeZOC
+vxBNlICDgY+V4jZvrtMKBl80SaVYFiP02KQOPbH+2/0nsRP1CpI29dbyrSco/kFOsus9p3SkYbU
mzPo/HSmC62B83oIKgwe3ueuXJEhQGPinSp3wCOuqz0OV32eLm+Tsi9OVRq9RZT9i9QR+mQgtDM1
KHrU1kmjaWnvhaoqBWKhe2a9DVbN/ALB7R3ogoXHfcz1QCa97QhiF8jAliwRLZCwB0/5VN5mb4rr
JD8pvdqeCawMzB8TTMCzNBwUNzLrD11zdXnrGGa2hWPzDso1oG1/ifv0Xbs0bBHhdIfarNzy46V0
nWlzgHDwGwT/4d5fU5KteinkT/iqOAesKpEEFSOa1ZMv2seiccIeglsRhjEmZe2Sk6bGdRfs6dNd
FS8KJ9bZ4G07THUrjWj4td5u33lR85KnubREFam06oW97xG80BgbGMt0iyhihFzUkUE2MEO0dnlA
V2CGDom341b3ql3X8qtcJ3YJQq8RbMqZ8qg8ExyRWSa7r2ZNiAVlWJsrtqStrqWul1rIAPlBt9D3
rb+4W649WTeFUOH7LUlWFY8DHyrci9oloVok8MwOBI8ailqWJ0eBFJKt5lHB/yycRJzU/0mEdvXN
FzjMcqVchLHkYlrb+7ELPPu0CV+NQVWMgdEHa3hmCDD3pqy9O8dlHtr/fRIpEAl0cDPmMqYzZndH
TAezpiqvfLcLOJcDCPHr97G6F/CAcvDwJNCeu624P8bRRncIB35K8ZNiRSEug9pWbKUvMvCVtjiu
Z1gIVgrxGEvKv4xY1OXIF6Jwnow2jRSYj3yhLEYocutSr5ynwFfDL74uruBAiP2EQrZOtfQcqh1G
c5/SXL34dVmL1IRKsou+oqzD5jWW0OXMS1TCsJ06swEl699HITX+ROkZjgu51YS+KdeSwK4aoqQs
SJjck5LaBsPVAlNPe4WlbUrUWPHfQI8ULY5I22rCkZYqj3DRija7zI1zWqbLtIJOjcmeinfq2CnX
Hcexspm1f2ZBIb9abzBjJHEctjcJy8sDdlkt/tZQrE2dmMixTF8CqMFxzgF3E544jS2SdfJzCj8n
Sq5ktGKb8iJ1Dx2GhPSiBTkve9LbDXfVMwYaaGKOQxXTQpb0B+2zffTDX9oa9JpWwPUeqkfqeM8o
YWrlembWa5367u8NRmceUqpxMbtzigR0wmrTJyxzRWONf3D/t7IFLyRyDT9s0r2hjsOqpyjSBT1O
O+5hpimf8mfXFYykQh57fOAdGUhBo9NmO6j1zkJblwTDp7AjfAbIBITO/HezPQG+v7+FbOechnqz
FG0Zcf0KvJdFClBLOMUZ8YLcDMKySIlI44nG+lNdD0WekJYk/utK6fG7miodR0pnnrDgAYTq96oO
jP5O55ngJ3m388kXKdrc/komnt263yMcraTBGCBuW7KPyrIOrZzClqit4oGmvlWkaYWiw8M9uH9o
zkpl/DaJVSqs1wvPalj4uzqREoVON7RM0dty/fdykZeGmADSWic/3WTOedNkwFEgvZJ4my+fn1ke
q0MWdpEmDI/0TYOdRRSPSER9PNR+XERnAFhK3J2RvYlL5QSeiJHhiHEvfIliZvSRlCzkwCTtLNNh
oQMjIPRq894lQVc8xA5vHsS6VBcO7oFiAfbAGMiITtRIOlbp3F6uZb99gA7yjt3iifnyIExkynev
C/wpFmu+CJ7JIBh9ZwX8HPTAq9JWLu08k2ZsTy+JI4thGM/lXTpgdvoZwSDGL+xnRKlmN2XTIuI2
kF95J23o0dmfalM/ojuvKG0lngu6sRrcYjw9iyQdEPUkbU9XwyVn+lue3KwOCqQ8kQezN0cLEJyU
JXOflyNrwJO/W7oS60LrDYuYjm4u4E2eIc5Tadgj/0TwusdilbOaxEdRXL97InWFOwbGDTs9Po4A
ltyTfkt19R1exnOLo/j6SMgundHjHg7mv3szJZC41IO6yy+eKVkPZTszs9GEBnoTh+e4bPltL+MK
gkzHMyqj1Znp76QQWF6/IrwEyfUUx3HSeNZ/1knHT4MWMtUqsdebl2COjk2U1lmCCt4SvL6txsy2
78lXVxSE0xCbYZWfWALVRNgjC0yXCJNBvnjM81f1i4VOM1K0PbndweiYB0D7qHvbxMQaWRkn6L4p
QowYFuPApoUgI1NQ1NSbZ9jgXYqh8/lih2+LKolUw2Y+bCmm906b2sG46h8KvCi8MVR8krkOI2GX
QJubjULXlJx1PZXyeayHHjrr+jnEZTWY3EyH5Ag2rgDbDinDLF8SH5nfp+mHdQVc2u34QahPUz2N
K3qQVewhLP432DqcKbXm79U7i3DEHZ4zdxpC4sFIkwextF2EiXNsrWXVQq7OKpyFcfosFmd6LWPO
mJp17pzLdQhpyt+626KdtglunvLeaUVtMyCuMsJ6V/QvQVG2pMvfkIKdo4VRXGWhWZjeTQcK4L8j
KRwS+GTW7RriswV57wlC47ityMqweYabz25Xp9RT1tuRpqmxTJHOG1IhzmJKycngFpbXqdTtWQgr
+94bwXUYJtUxyEVfBVHWf7VTZGI0k4OCos+smxWgYX7RxJMoVxLGnpgKfIwRTuqzZ3a0jZccR00/
/sjSOtKCegAquTIfVsyACrmJm+OvtizUrv3CabYMk6+6F4C8flJ2weqXLB0hiGRp7z5xyR23fIwj
huKnZZiaI8rVzw709in6MrWj8WveWRG6Wk4aSk+1JjM52i+vnaleZzOLDVRIBFST4OOFMmpcRSmJ
Dve5ukrr7n21idOoE7IPiZ8K9IHYAFCbVkgU/d+dUpwmuJgWkgn0rYkDKE9QgWhMb0YiQxm0wVeA
votETaRoXNg2b4ivIVAH5MUMh9vdsnnN3ttRE+0w50oRZveB4gYLffdMCXa2n7uRWSPeojDIfnP/
vKlPL8bm6BGgoa9kkAVlBJlTkpUxDQBjMlKwZ0B8qe+r7wDOo/KOo9UbKzOKGFVOT6cVHM1muvD0
08vneheQnzYU4ZsUTSrTLnBpTzDUWFcl8mf+EmkQkf9yAnknvlyaEmkArLyRUJemwVpDaq6g3dWs
WmT6gm1ysDBpKOUtY7KX1epeD4b4bwkJf1wIWN5uwBRRnonF3Tohqt5gBhexzNbowoVZTd7rGoh/
vJ1rmec164IcysVtKc6WBCYcSmGtDTz98qtzGqzurlGhzCtlkFHLh0w3rlaDCbCC6Y62Bi+GLj2V
vcTO5IQNL5WixxXlo1PwanoSNrJExh884Za6p0vXjpiIaq2oU8O89e4TMo7Fs/0oiT3yIx1Ku7Bd
6DUlq3epDYtwZFtXpBt1utlNS0fLvBQ0CwYtFAMNNC44VA+rrNQSInRp5BzpPyBkcY4InWkEkPzl
W43Gm0yGjR48oZTIACYYesBteY96AxDRMP221EbAtKcghascfy/iavlLQUt2Grw0VYGhHmkWwxVP
ToUWobMAgdk5vYqeS2nlHXNHhaNf8XGqvJutafGr/qEtsIKpVagwyOLDLUeNM99+5TY4DIJvcgdE
/gbLyd2Vb2UYqQH3ol2j6oV5wNjTqYgHDJFn6O63k4rNkpCfLmB6HU56egs6N8Sy8V9+KE9o9DiO
icSdQzFMQ4p/rzdSLkK4WKYkX1SqjuffgHCOPLRK9CPdychTWPq8HYvm9wehMfQq01y7rdf02NE2
0/wZaelaw2siZImBz4H1f8Tbdm+J4YdMtllD32WAib4GfBATrn+3iDgTRSHXx9WDNX06by3DoZHW
Zng6XIQFSCJDINJK+bUe844VJora0keEYgz/s4QgVnOELD4etKmF3xXV9mM0I/IaiXb9eyAXFBO8
PDZNC9E+1nPhnU205IiDq+3pYwrpvkPQQNDjNduZNpinq4yF9B5rd3ihf7ZGGameSM3K15gzkcYv
bugZdNujphxVB834O3EnF+a0U6M+QHFF7WkDd9CF/3bz3iqffJh8a12fUpLlPBhORkxzsT7I6R7/
eHrNAC/1e7XPeuVQ6xFJSjtu0VV3Zr9bp/G4Kp1Bc/QygNWOu9TChgZSdaeQTNjwm39ecVcnLu1T
1m5hcctT297E/ACn1avKIb4qB/H7CBRHZCiscbfh3P59jasNSeQH1mz9ZzwIW2zvyHEbW2C85NOC
9QaFFmfewMPY76qSC/EdDDJoSukCieUejDK1wHEg5Uq2VSG2bPVoh/UWc2JoRHuxVVhiuzOl1Zqz
KCAA7KwUbi/oHYC049VXAm+TqyuEDUG9GpwxnyrIOgvtE5rprLPXZ3m1Nl4ro2v/YQOdHl1NEA9u
SwBwYAIAbRN516UKXcU9IgRJZ9JUJ6Iy2BBMWTRQ/7BvvfSt87Hu1rjZR64CkgjtLGtm596OWyyq
zpFVqtZPij49JTXerP2kY0A+OT3BmsY4SEJSO3M31FWHIxaDd6AWPAo1HSNHedetF6TJQXJEEDkp
lvcTBa4vu/MKSaGhOM2UmI4P1srDtw/Bc+h4YeHfjZdAmumJErrZYEpaKi+pGzsz36Q/G8D50RJU
ba/kdQBq6H74RmnbGYmQYrQMmAXyGeB0abCBv24HsAWIf9HHH3qFABntjR3nHA6YGKh4wqyaaXBZ
aiXZYhvRxkAb3myU6luLaqcGvFM8KBPmDwe9761fYkQmZMD3VtG0BuA4n/B6lNrWAe+Gi+h0zztX
g7sxGPdLfbshuYQkVSCDvk3TJBvm2naA6eB0/cA0kWOQIFyWOGqoimll1Kp6JeH44a87dYkRl0c3
t4k4fZS603f52o9rLk8SptNrqEf2NszDGNA2agYvGyttcVgxKe5ybWDXrFpkpUgU0bXFyfEUD57H
N0L/nD8g2Tb7DzdB1bwxEKhqvPZ5OcvyU4UrUgpL1rz3Ww4b+43lY3EfCrn+jE/uIe3zoFgT1XkQ
8xmnIcWP5eR4pfUd3ubR9b25sllYYep5Zf0ydT6o28M1GjsajVXX3AvHhKgkhUchHUGJMaW5Y8ig
Fjih2oOWhGLz1KgcGR1T73XCnga4+5WamAcyPLUO3l4odgP8ESxcQ4hbkmBhepl8mWkacgpQE20t
lETzCclns+8O+0loLJydqGB2KxZT4jd9rXHLmHkI/hVpsAX8MP8yzgfvGVZ19TPcZ1OtKQxuD/7z
8b+xANnIEX4GEoCHd9AVCsnPHSm9HIKZaUPUnkmacCOcUc4ydmx0Bcjsjq91/chkYUvHrpaP5K+T
bY4Shl5jdr+obMrUCXgvby0tXNIeDbgPGLYYsG4B5g/YVVfePp9ubyrGuGkfAlwQyxgJrVIxDfb8
iIjmRMuMY1JhqAWpAG+rzXC2EBDhlXLoOBOCGxJT59EbenLzqB79R+nDUAjZqqAR6MxvaEx12ESi
2NlFUa2MWDjokssbSPKFXujQnSWJ27nSMKn4evqUc0Zy3VVKQ4MVYZqiZewk0y1NvwXFXPluDYfk
n4MF71EfItazoafwSva2I7gezh74hn0I27iqNbQ1jmNQr8XITZteze4HgZ4temYp/Ty1YhB3XAX2
kLe0D0q05QTGasSLd9MfM5V3cnOxuOJwVEQv5eR+T5Vn7Jk5A92++9qEdB9bV/2cIkXge7fu3AcN
8b4Rs2kN0TbtAWzm8WFEAxqTlRAY9DoHJNQ4ncPEgNegZ3xwrc4BB27cGKlfPoSPrHdQrsbzl5aC
T2JMK24IPc/qwE08LK30EyLK3LDpn8XmADc4rXi0qwBRXuf1D02zAHVY0mda2f2Am3UK0M2kAt3W
VE4Isx4wFlgPfbjfpLcyB5yWG1tqyo/pDlW9k8Khr2JRNnZyz4uQuQkslJEvlyPhgQka0wg6y2f2
4IhgzJmEA/3Jn+6FNXtwSc8KW7UeI+oW7TsMEgQjApdPVRzj0XLb8CBb+blEbiHBczaynfxRqPDl
88TV+VolQFNerf9HhkZ8VXLrUvLbONPfgdSrKFAIKAXVczUk5ztA882xBHQ0y6zVJuAGysOMN1uW
g0oJqgJuhtE+s9HRq4JBaC9EMkHyFNqJcpWIltxHi1ErzgNOOgsaeCzDEFC+d8H0pQaN27Iy2M3+
dSuzwRRFz1h0BePCqxdJZrCBUQxwITVyxKIj3Dgt+IqlYC8Yxvnn1psltCt4MKnnKYi8K3VoxW5E
O5Xoflg2bDlRAoFWcqi73xLjVU0owbBwtM9EftFHE8a8fIC0eiJ88rYxnM8L0ETXqZlwQzCdKMJ6
c6f3En8ytLQX64DrbVrxyPfoIdlhhKsNFyG+k2L2a7aTIdrKF0bfWe/zrfRd57u/bHLbzERFE8ju
bn7ltoniwx/qHjpKX04nXhNJg7jIkCVF0tEFxoAxiCkwuRw7b6sRbEeEcDj/uBsRauDu6C+8F7n4
3tqgF5vag7zjJ4XyXMuyX0KAMMgHiDy1rf+qIBfuTF4YZXFQDzD6bUrRR8aRbSKbLI5Qgem1CRQK
l/Mx/V/4poUkM92U0F0Rd3Lgp6O2/oYRsHAR9SZQceTyFcdwzs0roVOtqNZR5ldLQkYq2diK7cUH
6uw8KRmGvdn5yW8NHte3DBi1kQRU7nU2sx0mn5rHVd27n5GaNTmgr3ORml+4RCAcQrqTSCI9xPNo
LWATcKMadKMKLHsA/LNJ2rM1B2NnS/k22DfEMMGNWJnN70BqgfLmC1H5qO6xcSD4Lk3foW0Ja2ag
eGnhNh+AWAHHkt7oQjDaTYZiMFeU9cSCqj6BeAwt9nZGa0DLzQb7Ktmfe6zoCAC7BfXEVFJNDTdK
n9v5GvzX1KrlbwvRlCqY3rlCBYIZvAivxqtbOQ+oJd8gDo965v1Icc4U3qTOnxixdwUsr/WrNNNv
ZWPBnQJ/cA8uGkFfjEP/pOHtSQ7BVyggBupTkC/a/OyiPHY0NlNX6ZlWYqt5Bup27bFjVovao8Xj
ydH3wp7PRfdNgdD3nJwysohgqF/Id4cTQiDFdGhAf1Gln0CsME1jGbv6VV6VYyQkesfRM5ZTaVFt
+OJCPpEXVSTKbIpc1eGkEH7nJpQf/zCXTk1isHyu82LM8+9l0KmdRBt6fjOqCamjP24UCJbkPyEO
UoNv0WLFOsNSXgYz23crXXVCeRF1A924m20OlxRWdDXZ7+OmYz9sNUGnwqxwHuM6O37menCieiyw
CyTwvbfUn07K8O1JZWqFkwmWrKSMp7UtT4ckz+ZBipPwZ75YgBoNGwjqPt9pTbyGLvIhIxlSe4fU
6tu5JsPOBJlxIJRkPVzHsjciHpumsL5355nxb6llNk18Gk77UDPOHzPbLpCi5YQcwcqV85v2q2JY
Dv3WM7rmXshMNlrJsKnKGxD5BKLq7bPpSz7rYpWDeT7bgftTTpmpvt3dZ3eAqmij88m1DN5q5LeK
I1JhcIfvf8JEvNZIlcWQRGROpz50R8Zx6STxFNp5NB6IzfrnUSfz8Y+CaRw3wsRqDgAnwunH+0pq
Pq+YYa+CTgP0PzN0ggc7YuNNzjSU9Dys6UneIFkcvUg8qL0LgARU+Mnhg/Md817QIbGKk0zgUJOn
hkV/OgiIDOWGu9Of/q82Tf/Xe7XkIIvfO1RVX7MA9x7LK4fKkcQdKvewCNLlXfCKvgF6XZo2LqlD
KuUi8hNWVTAK6/Bo6/qwLpaUYzNy51hAvvUIlmy5aW0daGuMRwZM4X9eyMh/RCDWWvJZSK9CbV0S
t5FYD8OINBasFbsxmwzhL1/Ph+BSFQw6eYjRQDZek7jDehHZXZj4d7D3vNBm2KsDJn9WT/MzfX5p
smUbjbsQDjouTkPfxUstUByCuAdYHw9PnoTEh/zL09Q8lAfBpV2pTJ/GNmENHChNGRd41YDJBF3R
pttlnsQ3qz2AfCoD93G8w6GSYbiaN4bjOhaddJgmEF1LO3BsJ76ELETYgdRJv3j4gTmDp1F53czl
k9uRN+My6Rf4FUSa2IiEbodtWyZooyk22E47xe726zi2euXA5z89HB5+W4bLiGmqbB+o65aMozG8
yCyoFPjwCbeiRPqE5rzL3rEOg8gs56X9JCzss5jYKY9r9f6ljm+yurkAGXv6CCqcEQpPtdb95Emt
Ql9iqFn/0W4x5j9mSLlI4OZCd3whVtmNyMEls4YNuGPwTap9bX77Frv+DUzt/767g6iBzt3sv5bP
fqMWZE11f5Uov6mkO3rq97UD+RC6TnrmBK5Iag0mZ+Ou2YhCxD6LvtFsOJ6r2Io3YVUIyUZ9sFGk
4qgCk6hYhEyhHt0rZPl74rkvvP2FH6HwU2buyJwTQI0CvMZd/01rYHw3C7EcudDk2SRSWlcQDXdu
A9vxriWchWeSg87wvmr4BDvLdtPG4UqTMju02Sl3SMOCHvroCNvNf0jBivDEkRZE6LQeMqY008iU
DPd339jhQemPsRM6PEx6EXJfYlCEGtHe1nci7NiAFUADtXEOHUDt3ljtZ5384qPWdp1cGBjJsD1Q
IzgdGDMzo639XOBFpg11Z/SfTyV7xGACiUbCl8xCSNsRTVZHCXUDEJkSdpGZEFsyLf7s9UiQ1eP2
HHxjjdGII3GdUCCzMUo6L6Rw2qgOwj3ArffP5kijx71/D8q5nC+Z/bSfNmeQPFITJIn03pbmaL8h
qblFIr9g4ZFhNPiCRPTzJ9FOQmiNoFNTRVvnIa4eTpyGlb0JrhDQZfPtbB5jbgkaqWo96d5PvP2g
kHXzzZCyIxWtprcdQm6oGn0A6kDk1rMI4NN4TwNc67hhMkiJo5lSvi40g3ynbzOxLgAh3ZOFeWRX
nvK9jvSp1zdab4dr/wqI/IdzSr0pb/OgLF1dbfLYocENfr4KoPQhlk1hQ20qzs2cDO4VkinZ75c6
TEFnhOaR0sO08nyr8LJKj1tu2TyDQb90YhrJkqlM+BvMGpTWrsrTOh+mSSG9+4uf876PdWQLoBEZ
QoCP8v9ba08CFhPYNFuGoEm3g2sjytSoQH6LdIjDC42gjAgHRkHlmjCaVMqA3jDidWdL/AX+Ami3
u04fIQcG5uQPsuCawBbROf5IVC2/01OaA13fFVNzS8VGechuwwXYXj286X/HMswKlRq/8jaiiMvF
E27xhSKUtGEfug4szjWBBh0ZNpwdkLmaRhHkSgdTeaTZ068g0pbNb2dcF1rPxpFK3m9CzCdhnaK4
ONdAqLBZWzGE5BTUVFhaq9Uy2SN5S0UPwBb5kY4QtxSpn5hXzC53PuSLXpcXQjM5gdibwvqgmySR
GC6Cd/7wLyWHQkZosshXiH1Kd8HcUucPRpQyQ099o/JI4UZ7QoA0s2oA1KIO9aflv2+KqQWlyJRt
8tLEk1ndirH3Yy/6YJgCcWBBIUrpIfM9D76xkLX9BebUthqxXEPfLnVdJL8HmBoSv1QejrqQeZE6
T6+s75Obio894s0NpNd3rKPAgahaU4QHxL6x54v/WpDAwqEKsyu5wqIGbXrXeBRDDr7XqKXT4rzs
ynS0+c4YtV/kH1hPYipiM53KYnnGXbITWVTDQ5P3GQbVLiM2yi8sr2rsvBvmqmhDYn4qDRkzV3N8
bQDG+24cQyDZE44O2e1x4kjgjBRXThXdjkfGhWwYhotchOJ47LGNIOEj24UpqS6WIaDw6X9WbWXS
6zeBzSmm3J3AzAV4A+FhkeqXx7Ki/Ek3bU9neKUzmkZ2QI9vK/+SxSsTGNoSm1htI9WMI0affvCW
KJvVA8HsTOVm7dgDceNZflOlyUO58de1Cc9NNC3TckfRlbJYbV9KBF4fPkrjpAVukvrVmn4RJ7hj
EXgDpIPmmqc8KYsHNWvLtHiNn6NnrX6/BzLVswpsQ0xqkU0mOxrbdq/SBjWVhrNaln5au2z2qdxM
GeY2g59JpCPLe2pyaZ4QwmUTF8OQ3NtMFRShfhZ6RYBodyK3sdWrNfJg8blGzW608PxVgWCNwfc+
o1Hcr54W0MsYeWMiasUYnmoZvgLx3685GajManQVQU2EY4XrA6vN0pd/nT9LEt88hZLqVvLCRpW0
mXqOXpfHGIpULI5PIKJyZ1z4Ktf4hALm+Pws0pgZ6skN4mHWr5c5CNK0IW2iKgnpOtfeV4Zabl9A
0DWSM0h8JbEQofbcRsoHVz497ijCPQ+H34g7JFpO+SAVptzxiqDsymojX5SFqamtyhe648v4aDG4
qWVaCaGwG4DAj9m0DMrCOXs5sGjCrNavjuTQ+zCTED0SmfR33SJf+yOV+/BphzWm50WWkz9sn0R7
ucZ36O8wEPoHp3T3fo8k/HUvrp1FGxiAb9d+z76sQ8bfg5CuCSF2N5eloFzngccy9PNICKDYszaW
5eJuOhYtovWdeuved77w7/lTv6Efvk5jcGCJcMd0HC4V2DqWzU3alYa+6qGx6yPbfoCpiiJkU39S
WG17U5NRkrHtIFA5h+wxsVb0fB3X4ANlF7sa7Rlhx83PRnmJTeqgrgFlgstG+v9CTIBORgiT2Maa
QA/eR0V40nq5V/XoUZ57uU+3Lm6BQX8QCqMuzDy+l9QmjgYNiUAzbP8Xl6o+4mwpQma3/YbH6bwO
jhvj0y331+kJpRRBBBcip+KfsYRNbV6TM2F4BwrWBxvzaFZYSgDsmSZ/TaDaTutH1F2Ok7US53lZ
bTVpSQDZAtDxgExHaCUU0MRMZ4UdhCo08HqXJOM6m2uenE79w8JbxJ09AUFyyc8+taANHVExIgrO
jMxW7jfIjWsYsZFf8V2lBlxoMpbUvl0HhGz64r9fuQcwVq4T3Rn/XcHwSJJ/IQKn11r7UD0/4iCi
MKJcECFII6eLYqsjnJyDqgb0Jt3kq2zlRc5wIgfEk3NKSi6IgEyF7/z1kDQ7Z/TQvql0Cv/2sFOH
m0cpj0owdOd90jVPQZrDYIfj2IZXuGyeErolNzTng0CP9YFbRQfc0wUHJbdXLXHGwH1pl9lHVJVn
auu5sU+5hPkNc3odsN+jhJIuHV9zC+2qc245w4ao+BOR9P7kMl9gO6XMKQxFPwexIry9aCMRuHQg
uumyWID8xlbF2a2pN/dms6XfDo6ZcNcPhURc37GnMhZXN6XGZ/toy+2g0WeTJhaJQHhNdm+M6+4u
JC1nr9RKXk3AZI+2MMm+biuRjt27/l3dJNb3rNGdYcc4J2GTDcWI2fCWj+nMnlMICOGUWVElc+NG
HmGDk1W0xYDkiylSTLAAJUv7/ZVhTkL7Pe5EZUu5YsD2hy5gX/RzCwmqbh3//89+pLx+bgYlJYQe
nXOls5ZaR9JkXc7l9lAC7cmTW5bTkpgQdafXodxoUak4rNcSi3RwDaMmtDmu5/V3b4SxABhu9aWi
YiojcxpZ4HzMS9c0io2TIM+k6Mn8aRnZYBQzq6SqI50roPM39EKXKxOpMQjlPHvjg8CuAbucfgPR
0LK06EUImJZDFGDLJL4JioSbccefUUDrxnxuiPhg84MbUurhzpwXPQCQQt9pIRY47q4a/5hh9tKr
ygBJ45syg9gDS3y1jaLHpm7V1Qh/SAvST7CnkxA6NuQ9kzNeFDJ4yZFwgRy4Hsj6HMvletwO7ZcA
O2dMvQ1CLoXZNtsDI2/VGJI9XFVImJNwNiu1RLIJs6fTrKP6px6INHiuL6Wi45kk3SR6oKK2rd6C
j86xW0/9kuGe6SAlC0dr1AwkW28rspCcezwzfxkyzxe2i37B1XnCw04zOysVjavig6+Zab6XXTbQ
+gcaRmk9rGyiCvjoa/18YiokQnsrcIH/GwZWNzNOKzXO+E/w6jPKkBDJdTbjn4wAn17eOf6BY7bS
m6A1vTN13H1PotKBeNbN6jhwhDjXgUB3p6Vxj2J+cc24+R8Dxso5Ptcge6WOyJ05dWbffJEOSY6a
FBswtp0iJYt9K1/KkonNsiWhlslBUSA86QkWfU2VMS3SbrdlRVhEudzlLFjGSGUxmpJFk7nrUQeX
8VsDz+Lo3BRFPge2gm1IEJjQp0Pl5B7gRSwIH6wuwZ1bosECASobKm8TxVBI5F8ADt12Juk1Q0Uf
tcq1oSSF4n7eQDvSDAlyPckPnb6qHci02HX1f5zl2ssWV5D2BVzVaneItrNzHRu+hbilqzW0RqP5
HJfwmoyHfpXNKjgZwG/1wacqnY//WZi7RZb5TtgNAZWoNqItuF65QtVodaPUDAIJRzXMNAb6Pp1R
mPw5EW7zPnlTYPCC4mRiIveqX6L5jXSYzEouXNuvkIHFZoL/xy7pRWPYar4nYNQRXTQQwGDsiqOZ
dqUX3hfoXBkUwgsePHv/WjbC9gMEKq32lx4k3OACxFjHtdjMzpVw/4O6NV/oOUeFWofRkhUsy0ou
MlWT+QX0bbgbeyV+pqU4voLi0FdR8ZixAjr33d5xK7ZHU21RgY33N9LyBKoFZsqqasJytna6/WnI
Wp1mJEbMt0fFeQilOiexsb+jLX9yHtbeckWs68VANTLOA19nN6Y6J1UPat0CWgZoC/5PnKDGJK/N
faQvtib4mNlu3IRV9AZenH/Z1R2LFW+1OWOFao1XRfL1/+SJyYMl5cvFBk5gc3LE/IIxOq8Ac+7+
YQdWdhvEdmJXJLWRp8xUNI+K4OEyFI/jqHI/B0/XOtslwjDI6g3UCQYJQ6QIMkzD28MvRdZHvrrm
JeYI4Cyt0l4pZcFXF3yBPPOWC721Z43pYx4jJZBMkUwI+YLwXCxWF0Udq1OBTQr4RWpDIm96V3J5
uRxMXCxae6UBWs4YEFnoiy98hABmZ/mdw2qoOLpVMpEkFAKR0RN1UstW5geCA5y9CSLrzxCZ1ak2
oV6fLxIUd0ojyY3Q1Xul57NMHCiJUCsdTbca+plUuVySrh8vCgd5uWyzSRa648TCL3KlOAkDAm1Y
4wt6YzIK+7Nd+JfZPY+gO0kJ0cMbt5USOvz0BUinTLR6PKeJS35TLJYHKxqdjd3hHTNpGJ2QMXsM
LqXMUKdr5gszPX0FV+Wnt8E2n+dvmrudTZyRhU2BwlWJckz5M5Rhfp8kSnVAfLSWaqXnm0sI8n7F
dYCVkDGgwReSZkkqtS/Bu+NNJFqkvvjO6l6nA5IrYG4MvihZ2tBDVC5Wu28hA5kCZnotLauaf8WU
MBNd3b0AwY4rsASWgqBMGDm/LybB5iISlkt0WBcEwzLAg+89NGhApYu/X+u/un00b6b3nllRDaCI
AbcIjsCFoONadRO+xla25/y1Qh3il8LlduvYm9d3kBZUvaZP2bd2nMmVRZm4bi7XaQMJrDQ+nbuT
oDv5Mh4/hL00Smc00tMyvLNaURnL7ngxLWEH4B7prJVId6neUOfvI0c3k0DWjQJ3Frl9mFEV6Hpf
/9gaZCcqNfRQyaE1gX0fvqAdYsNojr8NHcjRZ6fKr7aGZVwQqKKEOIAgv5MMWVjNVn9Ah+7mxey8
bS5e2WWHXSUFOR1dmv57SpPZaZDxgyP81iOtrP+xy+msaHIQjhtLY26bS6KM0RX2ThSiezd9e0HW
xwdis3LopN5/MU1OZuzUkkP6F2oVQGEaAm2WzTz69wyvcS4WW663zgwZMijbCsdGlFltJY+/E9mJ
wDZYCctRBkcqKf4K2rqYWHEpzIWTpexQHaKFHXMTZOdtptx27/OgyikLVZeKgTBSOKiVQKRa7uIX
YtgcOcgb3LK/8d5RX4e+Q0oDu6e+6aUw6+tlZgm4EFOPqEp+lEGYDYkYktFnKkK3vHAy5yZQZ5Pw
T9eW5Qomv22CHG3uUmUV340J9NFlT/bI4X28+27t/3Q6TV2xawY0iiXfWWOSecRovB8hf9t2+Kcr
SuYDbGwnwP10Dbu/srGnBFjLPPdjS1Zvla6lt7AmjSeK5dEfPDC9YEoHnp521Kyuxu3WBBg/Kp1X
0jICtx1QOF5xM2B8ckE5o4NTvVjbH2vVlyMqg68KKhdbf/SrAdR1X99Sx4AyOeCXoIym/ELB+lU6
ScrHKMFmdwfupZ1KvTHq3Plyy+SgxgOKjq6R48cHGPL8+QB1AANT8m0AMFtVSvOX9vaAa2mgu94f
47UdShRf41wD0sTdngmREV5la9XALKpM0nC18GyQvkm0NIgry66jUalspon00n17G1LulVIdYvW+
1+oI7l5JY2E0Xhd9UdAovWtAb3U7xPPkkf4EiNm16JBwp84B87pgkapL9zyS+MAVx366lcQF1Fa7
hYhVRFxV5nLdHMmdz+xkjKXjVPNG8xojm+ea8QdxwKLT0NXFnjnVB9CA3DZQPTn4h/rIHsL4Ylka
mm9oX5MiNSJPiahvRhxsbQm25JtrLHeHaBpKwpw0NdYvyTo/nDuNm/PYuHrXl8lrVuF3o7ZyTb6t
xy4YAoie65XV5uoMq84P2l7fRavsj3Dx855MEtaoILZzDiEkQD2ZYbuovyhkfgONOBihnpD32a/d
lYa9qe5hzljwGbN23js/Dk8xJomFX/gwBV2vJRCFYngssXfO8k7hvjvoSHn9+cm2d4iAvfjmh0oT
e3d4WVjrMkdjLoPKoecdkdVOTrD9lD4SeoceqLX7SPmb85IUxjZLi3gH2OxxHnUrg777e5MkgTwh
p9LDqZsAsyAmWCJpE6b9f0CXVBjRfRjGtSkHHm3Jb4g2Dv6naZB4HcJ5M3DsMB2wqntApJUd4F7e
Kr34y4esw5QJ3+/YuK5mWVKQ2UNfMAejyo37jNYFl+H/ahWJqIyPp1jVPE49uCTx7/ux3mJGBqut
61yblm6mnTO5tyXJRXBb39z2VlWa0yMBlTNnyIWj3MBSpg2mz1tYXKA4ikxS+jktsJgOWKqctBF0
D3YApR8eIr0oQA1l8UBqxfCIz5O9LcG3RQuo9yS04+0ePoU6Q/rGGZS8zmEqGEyiHjh+w+Zt1Lje
IP5kGeL5/PnUqZSk1QuH1TxxURrKEOMhOnFPj1AxrfB+zJfbQKWe47oc1ZOtCa8+hcJjushAeKyW
QQwkQ0X3KEevYG7kT8hIaN2KCP6SpJVMq/Gp8SzY9743B/OYWBo7OEf9gsc8rt1QqUrpRn+bhref
I+3nXrS+3NFDhUWYUeFZ7uzyuKejAlP+NqCO8vHcdieI6xO8LTsDO/NEgcOkDwvx6FTyYGceWeDi
hTk/BLBQ3V2DiR6uY99QbgqMYc5dFx6Q8KAzSzMPUlGeH83lyNCKIT/0Wj/jgg9VH13t7aYquvfW
4zr77wx6uwyKszNbDIBZGFfNv13fdUd0J+eMgEYtRosIU8h7nKX8is0gDa7wcCdHi3EQEze+3ADB
k6XnyRui3eBtCyHmCd5AvajqvK7NVym47mOjuH2pL7w0gPXjQE5YI7F1D3muws1+olfel9ncRwZe
wY8q9C759a6JI6h4ZKl0zAOd+MsZENR1SFSHPHEUQydWWJg0mOWfoio6IcmCLmeqe02LZEYnuwig
1IuNqkEG2ZWsBHpEDsQuyl1a29g1i5zFnYVW3Q2T2bXFS/HClToiwY/F3gcUjzGbJavhdgsfTpDM
frOky7CPwgBsr/6r75jV0Wgnp678nl8u27YZVj+PnoUhUDayWVMRl6JYs6yzD4TJQJBV5uedMaZd
JwVfdnndoh8w692PhpN4asehmHe+VT41VBqKejnfM58D/3kP7WFS2sjiRuYmhXNZ3u8yZqKrLuFg
AuZc5zlFD9AwRDvijzutDXM2ENsHLHxty2Hd0YIvB30XmK1pS+vKCqoY4fr2Cu3u6V+QdMXlelf1
Fys6r9i6LvvssGbIREGvw+4pJKQf0xTPzuTrH7QBo2lwH428kMwiraB3BYXb+jH3Zpu3gH3u2kR3
S75XtCqzimwARBvSr6maWYifqVF49yTe5daej53Pv+pv0g1I+cWpNZIN3QPP656KZ/E8J1S5LicC
9nwN5JATb9bYUq3Oli/Hh8myNUZ/iDe2gczdohOuO3NCvySSOc1eLwZrquUAyIDYfO5bSbIf/W2/
arBv32SsbD2RZqw/9HAV5GpI0LZRnjnP8ZR3jUjYrtp/3/Dl0O3BdXUtHelVWob6nfj/8/+po7t1
8eKx2DFn3c2UzGu5PfbrcTkM1dEwgYTcD+Bj0G5SBa9GzHUVQeFqy50kPFROcfESg8HeZbrv/Wbw
4qOsCWshCo2cjD4k4HmFZREkMuWu5HjfOb/zoCXr1NUUgTXLapaV7slA7ndJ2rE0fq0xM+mi+d2i
8d1wv07oEQDIFpu+bsDrgzUJ3dQGPll785KLNc2941Gb4tLIVVVZ8n5zmz0W6oBTA+eerTeQ9g23
Jysq6efdo/CWBq2Tw2ZMFTwssoCrnXrKJvUe3WGdrCzie0lcjs3DfvsozG0PZmAlIjdMEUZXawmI
npFPYskIxNym/qfwug1JGW7a2GhRVLbiORi1iEQV9OJzLzrtyKwWPN7n+0tud0850p23VNzolGxY
NQKBpf2quO4IVJzIZLmPAZ9KiOJpTRf9ilGTYvi+hreKY772MVgnXBFYExbERTSB276mDarVxBSa
UCcFwFtlzHcWBra0BFN3u6+0IvC/oD3qOMeTraISlUcTlcDmXqiOWU8qYB1LetqvLpsi0z+ui9mU
vy3F9MLu5qcLoLxLzZSDgjq7fNrYUkwTUumUvANeZk63jy2yxjVXGhAr6p0dZeNxfGwwuQvFOlf0
2XdU0lhUy1YP/3FZmjX6DylX0tW0CbDOxqcyYaTE1hnqrvbpoHIFvIgrWn6yb4g0kA8mBfjdjdbF
ANdF3DrWq1f/rlDUCQhj+DnysNPiFFnsnCQH3eBQ9nWIP6wl8aj9Pyzfhjl/eIyrSeI7VPdUx1Ii
jlesWdR4pnPvZApQE3KwOULWkmK1mwLdndwiYA/JgyTNTx8CB5qBlY+4Wyjac9ugafV5c/mcz5XW
FX5IAEVQNDjE/5Cn5gBMHu511/BmE42TQOl3K/wgyJpA6tll7GlRtXJt/FBhgQpgbX0cwC9hcWf0
UY/E+6y3uO7uONkZmiqiDaZL+mqQu7lxdURDWU5nSp1CSkfIQwGTWFB5K+prP9EoxDxb3FODX3Wy
0pmhX9FJN9DRx4+PBOEPGJehjg0xGTqAf2LBo3MunSAWLYsE7YGoZc1mXh3ZBDqlXQYXqbBwZctW
AgMwiI9yHwJL8reEku4+j6Ge7bXlqT49Otn6Jrv60AjXFtOQp6AbfwXCGqiAiy6OItT5fEUQwODT
Rjy6rC8QsjTwB47OgGMr2kUb/Nf5/U9TtSWt/Ce5gjSXggQ/DNpCzc/H9lpIpy0IoUU0h73SoquD
2HgJuN5agp7FxopyaOMGKSCa8FMvDSTb/trAihEpo6F79ClCcdnlZVVGFuR1QtKRjxQBuCRngYoS
/OseRzIyEVb1gHctfxynY+pU0q8PY0NvvVtorvGpuBM6MtRrTmQKZTc7R4Oc2QfIkmolrmpqKMTw
vDWtIjkanBoECS1yolPtAvYDxJDNbM6XPmE6Zts32TDSRyLs3GM+0RAGmacW4tMRblaUfoBB7JwZ
9n+VTy2rdN5yP320kzH79nYbRO2ZWbgWsDuUBht0oXLDtGi3uCRd3PsnwC4W+Nb5aupStGB0cpTV
daO5OjSQ8xqB9JiphDCoGzsQPGeQIF96nSlH/cLvE5txQjPBPkVMMgGui2XWT4j2lFHJ+hJl+uNn
8RH/Om693dLmPydd05rkT1ftKGCMQ8Dc4EaYLKL1MlJX8x1127UzrilqK/e9AdeVcYmbZmPeO2Mr
HCGYAMo4DX130uzddu5k+CqoKHHqaAVv2ri69lKwQbFtsxNV+d1WXY0ZpEf7js5wgySdemaBF11m
Tit2C9FXT1JLsUKIoG6lm3YxjgIu2rHg7jEIOx1IYuNbisfQ/Wd6c2PomdCoFRavbu3UJg2LNgk2
RqmDJegd+YOvTZK6zUhwKfnpMESVCdD252ZkpwntRaVrkHYWxIyakP9It7QV9HK0RlkVaY45ugKv
1vfd4Z9z/1jL5tvXdCfmHR9GT6//VEGELFWuSd+IMvbNuCvyj+9FOoQNzaugs++CjOWlF0KJQ4Fx
1xu9Yg+ZbEGyjbfcMOdTZdT6OrV1sIRF0d13fEwWf7AfjylBHeFYiau3s3n/FfyjxsByMKPDCXMF
VgC++3zET7AD2mzPVHMDdSJSOner78TbYo1OotwuHoRh1awDQRxxXAGtfnfrKCgRTEiy8j5TDKvS
dmmk5MA8g8ddApd/eQp1+WnEbHA5hxlX+tJ5rXf5oOmlvDui7qqyM8CD5ZbetFrUG3d2YSt5itzc
qk2RWpFuXiirSTm2/yJ2lhcpTj+6dI2i1ys382dzhTIEcoibzbYEt/yaEIYZa0ZBGhvxTJBq+YGz
pvw4SobjNTJWD7sncX49gRWj7j69MQraXUiH/zgtcxcUQnykKa7EQnf9ayYUALJ3/iAcX+/JU6vW
HMTBJSgkuAPHOc5LkBhGjBZCra6BQUmzmm5M9q8e5Prh6zOdqoRgFSS/2V0pR7G2FuUH+nELkDqL
7C+2j5IrDRBpNwuG5/esObLLK8p2YwIitvpwi+1D7c/jYWKthNNemC2DvqiDdwEkmjMsOjxzZIsU
XzeIsNLW2eUwDb08Q6EGlzc/X6nxvEQ7AMvOdNV65XOMc4dkOgOVYYrhOI8JIsz/dWONiTcwvzir
+vBh1AyW0lH+jpZD0HnrnpfBh+kHp12aWFWs4SmmTBt4TztEn9Jl5vVeSaVIJ2DhffWw4PT7eK/v
bMbAitSUx+CccX5pKKjYvNixxwZSgyW7SqvaKpP56GrHXFrpF67eRxv1hiFN0rI74+Ibamt50FXp
kLaGiNg4UZo/DTMDUXIqxkaSW7ruTyQrN8ArC+filxev90vdLx93b0x+/TMPwaG5Y0EzxIP3Ey9M
4vJvbCwWAzRFUPxf7obkUaiSeNnLIp5hYy/MnrsrAohar2V/x62EAdlSbDyeox7W6yeywOckbvZm
rJCsnYuqrJdpOVrUreKEi0EzLYVH14sOjGtPp4ETvJrE0X0KCInOyWDFuZVcrGHL+E3E88en9xnJ
8ByX5NUmJHz5eqgjnieekxqxCdRuMPqSX2VF08V6QvIDvNwcuAGJeFPKXiLHPppYF2iVgh0J6PyI
1wcXMRjQp84len5ATnFGbv0S7x8JbHIauvvqPYYDpDwUHqpTnOBj+16PUexEJ/5i5k9ZxgXXNphv
TM6hWci7d4HUrtWC3rgmljlt19WG2cBS69+nnAfmxWrIXVEmRlDPsgLgDJzYR+KObXpkCzrWOmLD
93iahwykMfZu2PiNdR3iCpBD5qnn0mUFHPvQvFbR61mnCh8Ck74kuwjukdPE72JBZsSFZMmyvXjJ
jM7E196PJoy+m/3gLk4xFkZ7xi5zZU2vKPu9kY5Hw6mjciRHr4Yuk4RZaxtvHrD6EEF892G29ebw
lH/9e3oGx5fh3wj7pb2QHV5MVsulo4S623ICQMLwT96jge27/lkEjYD8DR3yiG0U50uZnJcHoLJh
AVNrhiSsMhZEdO3KOD6LiVGvV8kQty7j2Qgiw+S+DanUjVNKaZDKjetjT+N/dTQnj6WDwmu4UX4Z
bhRWoDbbYMDtP3PyCZeDy/iNtOd886xVlhWAuQfZTs8ssXoM/UbfpS+hvnLnj6rrIGaIoqxawlm6
qwT9FBt3RBehLr2hfkW5e32ayC1y6IXUp/6IwAJX8Wim0tH09B/5V/iSaC2DBo0JYhEU/AnCBz26
1uzKMalpZqi9moIu8xXGL1WqR3IVKfC7hn9IqADxNOSNLmv6u7NH6X9bSQAzkrhSyHY+U9kudhTa
uyUlh22meqvywGHaCb60oO1QDt2z4bHCmB/mcmLFNFSOKPuGRwwH8aP96q2YMwj8PezM6X0lGG/M
lXNNTAJqXCHNEW+tTBJWhgOcJU4ZxZmYT3yh51ueBVBKnur4Mwko4vDctMG0mZef0OVhQpBLsZ54
f7qKn2L7wXhVLGjF2dJP58lHwv7RcxgULuUWBEutT/8xkFJ3OF7ZkLIWG8s0uHl6+XPXOKwti1V6
MLzgH88NtBxgT6KCCNvc7Hapc0+CpVo3JPZI3nmziIcwkmZ58jkkOmqozcKOwEN/AN1giAX2M1xX
5O2P7ylOJMMogVuPG/wQ2pE+FSjzpqR4fiUaN2BNoqvW+xyrzLNUhbHlVMB3Sqmd0/vWLg7umkWi
iUKU5iMZX235E/xSRPWhQQhxmHPzABBNcbUe5CgfHAiDRnKvO/p6hWePXgh9LxPKZpps6wMvCtr+
kORY3IMLHdNtsJHlvkzXHKYPsrQTgcO3exxUuQr56Vm/jvt/0ZayOvv5ulCwQqtcB6stHYKBtzV8
Psc3Qc2eyhk20lC4JpeM9zpYR5IDx76JepNrEr8EkkVnWcwQ6gyiMh9/XL2EY4cBrStMQOJLxVjk
Wq8YFdJ+Uykxc+WZo3dTZcNKfA1ytPMlCTwVdj2YwNIlZUiKwImvC25/JfsbupjmXSgGkex9vJgK
gCmK4KHMoRVA533VoctAHCVl6Id2oPOCsz1aWb6BP+qJ/fqLuTqJcM6LuH6CckQCxWp35jls3INB
1Y6WkmLlPasM5L1qFvuw/Xo75jYHH9NZ6GgfFGBHQEpRRmtrwGduWKUkdEX4PhuMcUSgz8iV+P4z
tGIGGxlhuEbNDcmZJK7WGaIW6U4BhWwshRznBFvaMaWptf0gwgElMJuN9/SGq9bWOQlEzEb/iDvv
OICuKpfQBceuFd007fOggY20FC2XUgvir4Ax1yn6UStlpFPj+KF9e9QYHh9WOq8/QSz3/mRicqau
2eI1w8TvJ/ZAuNeMWmmKCKyNZmcQpFX0xjdFXq8EB/nFGbpfAshwI1EcgfpRkH46mqq8r3iCp/q8
zddl8qUEcA8l/vGkV3iqsAUkDbz1TwMAfTB4FWXG0tV5zE/GHdLh7iR+bvnSHTw+8oAHe64HzX/4
6tPOfMeXJcH+kKJGZn6XQZ5Fjq7NV4MKXSrKwulGOjAY20ijQbq+kUi+E7QCHJAuRdvz0sA62zOj
9hKJbHZEE6KhVfu5t/9nFHERiMY92ryt2dKtIh1PBfGvkK5Lr5VhU2e7Uj3t4f8o8rB2yo4wWRAC
IYHoE2BKC8qilSYNowyu+6+pLx7ovv14u2pXqvk+FnDRMuJMMAfKJYlLGP5mdZrxtJnZjXFR0C+W
bX//RKAdm80rBeXb7uo5U9U8w5KymR+5o0+qez6atz+zdZM8bEsyo7mSRRdWqNoaqyuLQWHlcbS4
MHigtoNEV6oqK5gTLs4kA+XSRpPVMVc4QKiXztcbz+XS9s8Q0bKU2Dd28gPFvXz9ZVHa1OvEYhcr
z0rnFJ58L4ol1PhImrDh4YxzC3bE9AG8dC6rcAs4CBTjV0uwWvsC9XWS8JeOVOORl+RM8k5Yq4Er
ZvNRZ1ig57BG5pZnIJnMI1wpd4NMvX4k8Hr1m5kHuKTC5D45UcS4NHl/bTF2FAyjFAB3vQvYZfJG
S5ItNSc+DOLq7dm5IQShjwBSBVjgEWQ2wS8UvG//f8Le7i0dlG1B43so8Zo872e7ok5AaQTS8U0f
DdkZPk3V+2UsAFygNkFN1ysxSecQrUIWySobn9m3hGXnT+Lpn+g00gfgBlI+wTIShEm0YZLvPwAL
cwEdyHxfh3BwCOup56OIrohWtGjnWyxgHtiZthVyT9Tegtl0881cQlA2Kx8q9Jp1ZRJlB+s2LSxe
I7PiCt6O9mDwIxQfIFzsuAjljA78UM2H/Jgr49qq4C4y3tfQGH77gkDDAIia8ukksjoyV4kQIgo2
Ie4fMbNZBf9rLupaLCXTLLjJtPfp4T/TEHR6mnG3MagItfs2g+6h7W2jjh1014lb/tgcIwjOcMGK
lXD2b0Dvja0Q9cSj3ifOe0H3N10yq3nhstNfX21OWtnOhLjaw1lP4Arvx32zkdwWWOF5Y6+dejfV
nkxtKdgywAnCbWaFtXbRZtZRpJ3TMLZnohAXdfBcjQTTW2nKnoBvZ1KhXBEkLB8tSb+5prNZE7j6
Qlw+Fx9QWZBARQAldpSHQksICkIiKPKF5QGXE5DVzY4B2jStY9gc3ZPijecvhv9xKGyBTqE8iEa3
wz9ReKxWFNZe5sewtpQmllMnBFQ+74UYAXe5ax2U7lfAMDH1DmqMVtR2t2Cey7GGUZnoSnqTzOSF
Zzdj/DYWYb43yOw2GmDjYGWUGO0gL663vHXStYgcPEF9MbU3CfjXVbE7Ny5yNH3qUZY2XmDHlfFJ
Fng0JvYx+x4+bCphPXwAq0w5fpKTAuQUtFb6k9EDM/gkIxP6jhba+gwqWbtxmL/gUUd4DRQWmsQK
mjBE81C0HNdY+yKy2wffOmgbXHx2svMcLg5ueAkiI74X9JMorxGua2MtGYlSXhto2ZR0wkeH0ku6
lq4f4pTbA8jPkszlaO74EazasMHHiJ/lcs5kWH0PVVHir7vwtztFpNhdcnxr2/pZFaq9KPW/dRGL
yCNO6t31r7mvA6WMX1AhHv7CmJWgYySXwAhEe11vxq9dxQZmfPrhBiT5hFRwS6RvQTa+RziTf0jQ
TqfUsokEwg6PQym4mn8oNDJfwLVUGtiAntchSPKotH49OAnAnx8lv3GHXmLHc9pf3CowE3JydmNK
zlLFWPvpClRiNOddLr8+02LqJBw9r2dGth5HHQfREEVb1TcdG8AH0ZIghsIy8gvxxA4VWtfTFLJG
ss80SnmV/G4jCwNdLVMA/DA5mGYJxgbZ/9aA1phy62hrVTLQzqXo3N2o84g3Py6rMtGHPIFdCD0S
iTDYwTxNn/I0qBjyVX5oajG3W2Zun05O+UGTGAFe63Fc0+h27ByYPfj4+gFqonjt//OwlkCPi/Eg
6imoJVxJTZQdel/TqDbGStfLdGlu2Lzce/HnGg3qiqxKd7OGn8pTzuMMfBmEM2ACk4rUQO+Z+VnV
RN1nPDCbqLf85+s8pF4R54I26MKNABwpI01DkSO9XVzEgtLfem65CIS68XvW0+SyKYr0Ml5fkkF9
N0vY0DfFhEX+Y6f6TR7aeIcfjI7xq4C/KxcwJfEwhPs06aOVPMQrfj0izIn4WefwjMokbNISd93y
SkGPdtccDE1h1gWnk6g1Z/LNHk4pMDLMZFF8tJl5EenK2174nU7WCp4YY6kcNDoMDQeJjSQxtj7Z
0WbNGYEIziTIwst7r+haoVcbpf0Fpz+2fnJye7HSacy+1ehzEZjeYruM2SMZ/V6uACxyvrpm6QIh
cb+eUJmDkejfwXP2VpccEtTjgbRodTL+DABEfom9qHhz7UmdOtCHGOajL4ltz3mSu1pIRMTCMbQY
ZU+gjmr4QajlRrF29Usa/LJcB/p1CMe6O4JP75V+JWJAIBASvdS9+mACZmjb5nXGl5WI46KYQy4R
Jubp4EkfKvAKaKfaLNgx0f8lmn/yqnZ+lLU53TKRnf9WJOl2KvLJgdOmvx7F7nh7m8R3YMay01qC
vOYw4+2UEtDHQwmOxxga4apH+qIr7YuGzwL5y8p0Yb0LpxGGnzgBGOUyC92XZ/GCtO1lUggLPQZC
4WpQ7yynTUGx4wkbtdGl3M6PsPA3bodP/+czUA+C1Z0+UDtXdoPP54LVqIguzu19RQ0+TAE+EmAk
y5gJkYBjucuD8HA0gRgK3lEWQ+nbf9LwjZY1FKyYCT2naJol3wosWb47AMHJxioT8/R/F+wkIItp
+nFMHfrHMa4vYrBDVHKFwgElZzWdVlBrmMhpTeOdrpgx29VadYYLsK5OLr12fZYYBWKcdTYx5cR0
0IxwwGmI3FEKBZM90B7TbUjdoq7Mzy8ODJcsUBOffa2zpmZBTCT4r2MCEw3wSZe01hVIXkCCdc6L
oPYWu1762v70nhoacyK9/Kn9tWXYOY8hyF7JYq0tcMOdpqv/1ucr9+GSw6ONiWJ2hD7YJEIP03XA
+y3XrFNiDGyV0NVwHighOneERvDlHTespqGnm7K+Car0Vkb/2UcThWzalfsC80HTh6DFO5qbvcJt
M3RFnZ1Gu1uuwfT/oa6sEJbaApHk3kT1/rpGqEPJJ2j+GLnuxR7OmzocGjgNgJsmgMgjFpQa4PL/
7RXNRYE6hJZlUItCrJd+DHzhqdNaf8pfxIpl1hDLBtrwenktLdwBOBWMq2sKhXPwOY1qIxNXLwfx
6rtlOURt1+rbwknfnj8zGcJX8LgwlQBf6TpXfj1fgCrMb0FI80CMf3kufFr3MivPe+rKYVl8i+o7
zxItD50VdukbuK5XpDBUMMjjogk3qpRko6fxC0RnaSWY72sC6yx7CVVslJn0y9XToX32WFejgeOk
qwefqw9CVxpZ9cDo+Ch8TOjwkt09kZzYu4IStcXPoCfayF6bTB0cS4gl2DXtuaFF6jQLewgj7Htr
1ggR4SU70khyauZPPhzBMwm5XQY/zBdKPpPYjXXE6DXGqP2Up8ZIVKDTIxfQs7eJucRh0MQarzwo
wH4ouifTnBy1x2cpwhYdt+EA1r+p6xepT5O1c6W7gT+S94rg31zjzCjT43xqewe0cZPkh79f9m/a
Rg8mGguh6KIMqrCPLw/N6WlhjZJbAADAlTpzvmyl4oWxkVr560kF5f742N7MoO8boFEQpH8s/eMi
KnnlgFY9GvbDCzQqzpubJ0lWjSk01dEBRo2stCYYmAnks3WjDjokm97mkG4+zR/XI8SNWOF1P47Y
a54Touw1Ir7/u1dkhP/ZazcBm/kR49kV1dpD+scT88vKmNomTk7emyfpnTbOMmGc/7uLWoxgVeCV
yAD+ks6paU+4g4MlbUyMPoYxWgwOpn1+wxRIjwnZ+0//JezhkDisPD9aXV6Llv5WI2tny8gjUf1d
1YT7vCOYW92YXM1qiV0UdIZGFCWDXTpsdQUDADjaQHprPFHscpB48tH725iFAu2pf2BOFDHK7cuz
sHkiwVwfWjkFgObxETRDANHpeGUsWw5ku9dhIYBnDl9LgwQrZyJzCun/Q3f/mW9uf+Tn4UJeEFPh
/x7L6CfmYZXMnOHUKu2FYPAFB3fjTM8U1vbayLNMWJjEqXeCLdft9ZFoVKLCJvboDM2jfkOzyfKi
hkDH2g+COED4c1+sEHzvUNTnYTA4z9Qm6stUTJpfKvFYnA8hR7oa6cIpT5zqEDefkJtCS0Oz++jp
zKKNcEL9yqAQ4xfdrvOXKcrjmcMXSLivNyy85TCKVdendriaZGlqA/EBzwLNWN3iM6uExom+KHEg
fxp7m7Oy7QkvGodAsaJ2KnoacxTJy7W524sdxeALvQF3RcqngShvaMoL8+0pDGjjayzyY3iy4MPw
4KHGWW/0IIXmMUkqZzi+X7+UeXgwTXZQgQQnVwbIeDdTvizYnMtYKplMA8t/yhaHlxm2nIKyEAfL
zIz5iUOMd5gHOng9WploPhv8vH0Kr7ZbMTN+NhdsFbFBimQ+5gDNRiiwvbDSoZtF0ssMdenTLJ0P
8Em4d7WZgvhCoU11OM83YR0nxS9XSp8KaVidIkVKUzhltv6dRArrpoHV6dj7JPgIqmDilpaEJ4rB
vGfH1hFO4drLuJD3soeySzR09Womm4z7eUTD8NtQbTnwBoyvfJLzWczJv/Kq3/EGQ7uW3nCUB37i
F1CzmJZISsFg3GZSejp7gqpj1+nTk39aFN0vTueEwMDYbUIBvmPMb4WQRbjvWKMqunwxD3cfifj1
kknhKN99kGc6LIrKCQCI5SYwE9queiu+CM546Vn94Nx7f3JNMoS0RL+92nFT9U9PDwZTL86KFHE6
Hw9FyfU8s6OA4tNWeFKOHs1mI62CmFA1ogZxrGXBmYKYcSaPJ9y4n5eWWTs/qC5OBL9/P/dNULK5
ivp+lZo+o41nDKYmCSIF+wp8BH8rw5V/uBOb2EM3QeVVGlD3Mfqaq/LhA5z49akZf6lE0oGqH+Ce
Q+rbgCC4X2uwiqSaqmWep7BatWoMXFwnbxoSm1sMeimAVzGfJy/QjBuTzOp3l8HJ0zSdKffcm0nZ
e/1hNwgMPA4vTumk7hEbwFofiTCNaivYzBsGHsMYR9u1ALhyj8JLT5kQtv9XFVsZ7K7gRT1Ys+k5
bLAhloMhP6I8X20Z/ZhK2aXPIGBgyI21NGaeo7mXaE4OUfv6dMJxOCTB7s6oMVzfsrAdN1+5mAjx
ij26H3vpINOi2Rdtmdcyd+dW0b+BgEg+ThvHTN5JCjoR48oapSYFwRalY4GUIyuo0O9IvEoQm7+G
VNfuzOgZLtPS/kwng0rQUk46/X8OZPd+SXvDkzf8hR2cTzXk16qzLcW3NiY2ib5s7n9DZa48HCyn
bHEg++ncDTBEXLV45txYlyoLxai6ciAhUUkllgEnbkUMQaMohRQFQvavacrPkhQrel5CLq0PR5oK
yV7d+q1xRFRmKNCo+0fhJ+paPuz/OhU4VWn/t2epPqO+C437nmJIusqXAdrS/zS4F0RB4qqb4s8w
nRaXaDVsSpWK0B7WxPZ6ccElihimZ7s0mmWSQ6OXMh2wE2wEptwMzwMMhpHoFcltX6KeA6vkaKI2
ZHkZuOM9WgpqdgCRonEFtS2qdOwh0BFU8PsNbsnciQGZSuF2qvX7IxzmbGfBwcyS0p9ZlCBo2Hww
z4zcsjNe9zyvu1lmN1aLNO5IGtiBGhf+5PzEotFOq9wXTFOQ1mOQtTAPOY8devaH/U96puhzQueL
ifEyQ7ZOj81OBs92/gMO0Rv7pEBZuGer6sK+zqOcC7PSf0fByLseAipz9omkGIrxOF6WofOgkwed
obmMltRlj5FVRoP2S0hKNpoJIXjFfJsfmPSVx6fDnObdVZJNVYhRwWWPZsXOLPjZRxlFb1KJr2vs
7YUD8UuqX6y5XOhAAMmWpjI6iI0avgDliVlY1njsL62TZ5hM4qPh3cmhm2AQoaIEkntOCR2qR7NI
aps5pbSQSMensnZE4VKGoJqawgZx9W/zyZzX4OofSgGeJD2dJEI8/UNO/FYYKdLwJLlq/ngcm/ND
hRtjYxIXVTe6lDsAsA2i56I4fkfADD3vKVIex15yxw6K6dF5uQh/QJiiXZie0gs1IqsS4WAlX5EO
TeXr0OAfMgJ3HFyeW3hculKbl78CF5JBJOnZoooLug9sabnvOhmI4UXGf0V2jE5crmqPt4tYz48t
XqFP7Lana29PmiU3mZ5/Fvmqq/HBPNslqE8hY52+HuY8ka7sa4sIcXHvXP0EID/GL8+b589C+FnM
iiILiPnzh38BucN0ftLnL2sQ+JG58B1qhucYqYyaBskyYxACUCvROagL7EQ+syzXP4MojWSA4ewa
iCRtYEkGqYC1eSoITCxQLwAwLThhEujciIWqppQ50wSLTdwr4OOKVBiKxR5EC51/w2Mq8WoL3hrC
paphbMO+3Fp6cjb6kmYZOFRVi/11XQRHhCc6AvgPJaPX+t62cfHc/OywWbfaBd8nBzMU6hZR38Ew
oJwENAVKKfU8EpKyi3AdDX4aJwJY6KFllx1nH9HnOvkDWHpw1dNK6NqIoUpyUX9YtFB6QiVmBZRi
OZ6QxATWs9iP/J10HJpwqiUid2BqYhuUHo18CPzwZ+yI0FpBb/rtUhmwmkZ8VIMfdX2XdAaa1vJT
71fihDsRZohpQnqVpCn0YXwvfbjlHNnM5DRJRzTnZKc+HmkldB3TmcaPAlMbB2zrLD2/1O1V32aj
pJId++waS5OIrX8Ka5tcV3t23U2KpcItX2L5IGajyiuLcAemDOyFt7AoLosdqeF0J7vw0bd1PZuH
IhN8UBq7za7O3IDTiBpSXcPxwqsReyRWZf393ann8A4oMo6j9RXlxOIcQK8ffQ1kfYy8t8HR9dFt
SFcL1+oz7pZBLWfjQBDIbSl9EZA0kw0HKwmaZhFxJEbMXmnN5IYzBEhpMdOXo6lbaP0tGN81szAs
0R8j5qxS2TIR5cQZ9UksSUZPEGA7Nb31jOxXy6EPmXA2QL4kzhfKK6qJEyR9djHjwFP1XEPUE/+p
28XuESt5zUcosupZC5QVb36FuwKDRIfThed8qEvSG3BgL3J2TrZXRLrOQCSlgu3Hfvll1b+0sK/5
6Mup/Os4/1PY3usfqy5t10zWEen6zcCNPAO9mOX2B2wK2aZf7wwSzhzHww7SObmqxv5mJ9a5k2C7
q9ylZANiDhxOquzWmy+Lr+Q4BCHkY/EiLrjoYutFgw265GEwx9V+H+tdR0g3SIxubSivN6VyyqRk
wgIVJSG5lxQ2EOfNoPnqlTafwU4+lznz676yXjiajjr70pkKOVmhtHU7ch872s2XPde1fwkDiQA6
QsS3Uf7aXBqYDgyAiEhjlmwNGHy8eBzMufvx1atXjSei8yXm7bKZfQe1z6biYmBCcJH29qSek/rE
Jl12KmM2uXGZcGOjiEq+i7hSr7aaw4kIorS5MFiAlg+sLzgDImm/MrlD0t/p8uCgv0VUo+PVtPwD
llyXsvMDziY7t5sF7dSZ/uulzHurdBhUhH86G5MVdEVN4EJcxEJNRAQLy/eSOrXT30DsYpqDPpea
3rd6S78/H7IvW2eehbSMmh/rWtBHM4xeY+U2J3tDUSPlvFBQJ9v01eJ0xYpWdduoNfbGV0wyQAuy
uKh1+MXisFjvIvD0gTiN+fnPy3Y74I9he+gtRRi3P9mMYuRMKWNS87v9pLboUle0APg2qDoxxsdE
lezAGhIaodbnyWsnlhe8HX91o5SEcbGWE21cv4I9pXLxcz6iw1V6fPoKUMecPn33avL/kA81RFTB
Rr/vo6mXI2UnDSFMM2Te2hUeug750ZfnSxMmbVf9DzxNqChpsHL6IYhSiIkmU7DYUcjkzKkMQaTC
5ypQ+FhIkPqgMF27p2TXnmpegEYNEgh60pUcBnbe+TkxM2FeZ6MWwlUtNAXSHZv9Mo8eZ8Etv0jD
YjumuOn4Vu/zwIfIGN5+G7YSxkd6vQ2byeO4P3yN53EJ7mPjYzVbwy/kmqdLDUWbeY5b3ZsxCbF8
zN5LBA+CUYfvt9mejfWhDIO+r2LTr4nFaiDjBAoFIHqZUgjJGUcSi+szR9ahBBNGJwQ0tCoc6Cmg
uxs6i0UXLARXaQKRzfYQFi6Gf1Xk4eBuz6Lws5iUppERgQYV/36evGHC+ROeXWd3wQQw0t+26I+S
PBeuPUu2KNZOwhcZZkqH0+16KBa4T9iGU7qTfRBdVlKUKn8XClp4MQLuQTsjY7SiZfvSclWTYifG
QeifOj5b4w52tUO6ELMVRFXZvl2LN5ncA9yS3vS/52k1otH0jQb3nkrRyL8cyFeIcjsUVmRb7g3x
FzcN+y6MpEYVMhvaUV0Az2/l+tgpd5GcWPB7NSVShl679fphGm8sD0peHG8QPOwXCoV/X3zGjk9+
DR68zZPgK0qx4BvNO9IvCCOQbAYVZjBXJLUs9O0J0h+WdDJC9SHQgODpXjOE4udzIids8pzX9hzU
ahp/qtae12koVnhpkeVM01ZqgxVATpUtuROMElxoHl5lb7fnXTxPqZIc9w//4BgS2Mqf9/TAIvTn
9WQA0S8x5SEEBjHD2aNkdvY7O7lHWyBcU3Akdc7dNr4VBM5adBn6PXzvpABEWE/PAHbVwILspsAQ
d2EjvaNtIfS4ADCOTF4uuAeDBhHUID62hln0ixBK1d2ImyXQRqwDNkgwPPvWedwnvNFZ9aBRGX9C
pTR+idpHiktUyFkMXx0Txgj0YDXomSqstCWBPnjH5iJQBkN62C7qgN+CAdTT0kDHcAdqus73c/Vl
ii+VYUtDDngsh94PX+k0YygfGlwTM4Dzk42oQmtA6fqI65lP4o+KrE7xMJpyPpLQusBNAQrL85WK
6Zis//Lnog4RVUZlMOWloILIh6UvQmV1SUfEybFpOOjHezlgRJVZSm+Tl4z7OE6YnoRN8CMDGb4P
yyE24j3UT20vleLqL7KF925B6iyk5iOanB8chpG8RBTEaBB3xLibwEK9CCwrAfqd+uuuHtd/C83L
5G/47ZY3vBAzUIviDCXr6czsaAAEHZQxBCcZpec9v7ucXrCAPFTwOpXGJYIp1Cy8rIkM7QUNFbtg
veRjoncCV5maWV2KqCM02MSeGTb35zFRRBczOZaWmzmtv/ElX4s62Mm3GAeYz5hLA/PfRDjRdP/y
4zXJmK6EGQmut5/cQ+SFrCjnZLS1sJWNbzSiMtLzdPUZ+nzvcwQ2NBQTzY0GpThXY65dQByI6Iqz
ymK1igAaoO/U55nyKZUyyKy79tWlziVj7+5IY1FgcoRJwaKsAUFEMEzDjTu/YWOziE8c2hApsz6r
dFMx9zaSR4MHvIiJ+eNm+G02wMf/mLu+onOQsYpuOeo3/n7tY731fTNoTWvajkD/Zopd2MWlbYy5
vz7UUOuU+PhDPAZQP11CPM74CcQ8IndXp691Nq9htfiOAWKS4T9ksMvu6xv/aIYc+u3c/UQlSBlN
0xq7O+Lna0G2HZQCEhlx2r3vf9FJxjohuiUOkUtE/paGaPc9f5hPjFKXpGLAGG7ZLWDhN1Dj07GD
htsbhLaI4cb0Bwt1lvGT/WGDVYiO+Scesi5HtarJ0dQ/hbzsUzTPxqqK1VQrplIVqkxl8+BRhQY7
8rtZyoiLEMv9KIAUuEs10FD5qRBOf6Aw6smpPOitjL1wMtk2rcwmwlV3yaiNP/daca0mmC82JXcu
j+V2u8Jf9LpU71mf1tt9anijZFOLpsJi6dN8qIuuydtt9MVEFven4pTVyp1GA+tfHYGeLRV4Noh9
kNxb0pbk2ReG4aNjXlX5j8gdxym72lU4kELrqV9y6Bu2XEzSsqtDA8hH88j0yI4fwSbhtmXicFyh
ZhUzYLqyWR2xuGWOsfE2Acraxq+rhDMhCSYnO4GnVoWsakyZRBEmuCiYBUEmOvCoBDNetNeJF9U9
VefutunPPOwf9lW7VBN7lc/y9sKteYRJsytpn3rkvCEe6575AP5DYdV77K3Zvh9BT9Y9pm0HbYP8
P2UxFzS8+0F8TBmcgKLKw1D21rudsfw0RJf3XVl1NscZrtBco1/q43X3k3Cn+tDCsDydf3ohMbBn
7vXT3l8oet13O+IQ04oUS81ENJXvoxRuf0DfBR/gQyKrDvsX90MEI71wWY3HC66CEjGWKA85X9W2
efuBuLTusl1NSO80shWDHWn9lx/rHaFHoqt9wwYvQFRVAzpiyvSWsl1q5ijmd3BrzinQSzN9mYWG
8REcsDLkw+2UnPJdZfknJk7Za9DSKsfbcWoESNxakvNvqJXvU5ioiOCo/89qs0/JcwvpOiFwRpKd
Y+e0Me7vSlnXlMTS5jDnGzMxgmf1BIGb4foBlJm5fHnLyLVWPjdWIM5CCql4PIY9S/WXP4oNFH87
ID4HDNBiaeMHbb1xOX+j+gJZo597vAlzpFtg0zBn3o1sJsQq0AJldQ8dfFk83jaAzuVaC6FDk3+o
5ZBA5jlVXM4WMqJUUX5exaj7ft6tVrYRbXNZmW3SH8TW+ZvzcOJd+TupxeVTZAjL28ujoUQgr6V+
XOUBTuEgljfXMjbagodEsi0KGmouvmMaoTBMnUSjMJgAfna9A5Mb1rzPTl7aVAnHYjf2zbFEPk79
myftvX0uX4JuuAn7rTRegiHYiWqhRdSKnfNdnmikzRYnFIypxmuRhjkdALW5rqPTNwzcc4g60aai
sARZ3k7l5A3T0SvUhlVrM87B18szhlYKXZuusbIanJu6Cn4wfFUQnE3sjLVYZDWl7FfaTeSIiP5G
o/UF8deT9ydk8wlNCD3zvhIvn7UV62OpynCyuVpBdBSHtmhw7acB8sx2ocshZqEZu+YhxAe2Ruvh
w8Yxmtbemy7oxbxt9GA5dNCIL/aizhgj96HNkTuuj7hg5TUuBMWUL2kl/NqQMUu48l48QaP63wfX
tD2I7p2NpwGh5Dgy7HnSCklgywiFaqyXfDHVNQOkjJ2QAvEtQ9Klc6JH/qwcNLWOIkgsS2RrCc8b
wfrF3QJExvkP6Kw6QW0xw1o23JDb++yRtLT5na+DRLF7+UEPiMneiShDXq+LoUdE7Rz8/M9zJ+f8
UjhnFQBGkohW/tYjddJMFW5TLgNqJePyKvkctlh4AulsBqk40aT6qOExxjHjrn2s3mmDcorJfVFf
TXINuwIHchIkLObdrCEiriiJkVv9MPq/8Wfr6s5eRt+th/OdKmG6HEaRt5wTJacK1zitjFGjUQr2
mnNqdo+8bXBv6oc+y3aoYnqF11kglaUTrRjKS/sSjT9z7PdNpEJXhPzpW+CwvWcdPm1hTBdLrps5
ZFwvK9i+4yot34MHQ8vAWhjFTEeSvQ4dvsPeM4Hw7kxwGzK2k9wdyXdemM0v+fGKTGY3ymZT473W
FUrAlHgugkL9fiNKL3xbIEhIjxjiCC1w8+0/zy7lLWVCIyznjzEpJPJXo1hNwAvNvnR56CSbRiPe
hZ8OEoIfUeO7LPjsKbLBofaSjSZ3xDvkPK1yAg/BIz5DlkFdCUnOca5Mlatn2JikTuoQY5olvI9X
oqdYEBuH2SXXzqssd6skOBN78TVhPhCaTNLq/XxJm3VvEHfWB6bql876K14XPLZLBpDpqnZYZuaj
FqFsYqh2DU5LK54v87gCqNCG8hJ+WE4IkTAcWStMmVMcrTgSrCEGGX+ShJsq4QDRp4OAzR63m39k
2r8LR1MIy5jpjSLKXf0tfnuSWNoyqtaIjeDlC0koQns/Vg2hOXKFOsVTIW50OG1gNPeWMwBz0Ng8
ZEoz2B1lxUYysq/SPqjmUXSZZXDQM2vLUSRqplOgC+jGUcjdLaILKv5B/REb6e00XOLAPzJade40
gsU6QFNlfHQbVfJEk043P9W8qI4Y8EUD66Mn00BSoz7dKWnRa8UV+YKTHkRouqAeQMBd1akJPpoz
+ZV0Qf6xzGAPltUHUNNPe6BkwgEWlQV2Knsrs7ajLLIS8T0ypIXn7VtELJgiKLnNr8q52vLKdioF
iyvquytPiJNrmgcAz7tksGKXlIxpx4ztWGEnl9us+cbjOQeZ0Zsac8OtXhHH+jRIR+s/E/B8uCgI
HNPjv6q6N1FBbF0E064Nz4kqg1PWDHGMMyaRKSZTbcERQj6isVD1Z2zdHx3azxRTJngXbrzdGqwP
fJd/lMhclR87Sr67/dGprmrCBLQOR0E03ZTl30mXP/kRztaoBF3mjMUiQhWoFaZjeN7P1Y+UOurA
JVhQGJDjRy9XN3Pb3geFSwUjF4+d420CgdnMak/pJinnd/JYWQ1ZFA3Nxs2jIZheXZv2cP/iqrUm
pitKhz054DBClnUYBeb80EeSAoOSLYrXB2QvgL7KbbYo4P3YQ2+anX42X7wfi+uZCj1xBPIYOesN
s15ERAV/BCStD+I34WIhybnQ4Ih2T0+K2XWvLxmNPSwiW8Y+dMfHdz89Fj2foDF/wXUOQyChmSAG
0TUyJH9cgvK6WO6AfsB5fZ3IOOD+Dxs8Zf9UkIBRBYODTV5u46YSY07056fr7HJO5SXNiDkMWgYy
RT/75BMYL/dmEdbyhdIZ1o+wj2MDA5PhAzwFy5yUQYS1zb62eeHMiISLt6818D3O6GGZiuUyalWU
RQTCijbTOjxiEiJYT1V6/0uW7QM4QOTJv0ofl3M+Y1F5FWbbZcXIhR8bOXJa6OwKeRl/f8jnU2ba
nogWJ7Q8/pVikz8Bt9yWzZhAFLhbKO4W8bm2+uoqnEUlvAv2V19UcbW5IYm7DTA475eXe9HzGucZ
j4JFX0euujr2ff1Mo4AAXFo5xhNEA7q6T7iUwGCRalouOe44P+wWBWYGHcdUtXNN2jYuKgGjQncL
KPwEP1rH9G+nT7EBvTAoVv0NnsMlnJHP6jTDiUs928MjT8ApAGlod9sx+TRhPczjRb8z9EAdfdLG
U5mV8OImCNR+Cdw57h0betw3YNm0QuVse++FF/EWe95bqhBGQOnsK1WFVKoDaQMmvHbiX7AUoFwg
vZ8hr64Lb3UkjZdmf2C5lqB4A3eFszI/KTWE/fE8dWdSG5wB09wbCs4q+3t/lsYZqiveRGxpRN9Q
oljT3azCKVXruFvD5zP8d4EepwSNKiJtHuibeTDHYTIOrIrb9prope4fo8lnXQ8SjvDHP3dSINsE
5p2HGL9nkxr5cQyhhfRi50dd7TLc26Kw7O0fk4/J+aSwlv5/enZDYA26ranVfeUNYCuNXgQZdNon
wTVV1mX7z2ctQlOpwldYtkK+p7Jo/+gofekUrDBgKAgEtrNH7D79Y8OqhmVqv1vyylGvcG1pe6XN
avwzVKgQV4K0yj+S31Gf4HeWJS6BTDcNB9UU+HHZh8FgAjUsk35RfyXcSYhGoVk62/omvJ6bQIqo
KqoobGjKVrcN36nLQ9eFOT4eL2y2kOMFAobVfZpmaC++a9h7GD4QpnmFHV+92nzZ9bwJwlU32a9l
14OsJq2vRx2kKc+OAgwBFDYhnXA5YherVMC7kcUmQaKkFlZCHn6tZQ0qwdecXzOTF2XU1Bn8tiuj
UoHO21PMHsYoD33tijJ9RrXk0izATXYkdAWWjtOYiL8EGQIpKjaKRuYmmUX2ZaNED9m/4Euap5DK
eTTPWVNCz6aNw716x33Rzwh0DYbaKWmms3EoV1QaRlnRRkU8yE3wTVGgCqasrcWFwRYD3YG225RN
z59+TNBrS4Bb4ijITbBKNuoaHV0EkZiatwBv9ZuGp0VO/QUi/zRaKu6+CyTzbSkLcbbf+8LvZ/pS
TWGkmeqswe0erP9oxHCMppVqwRtmXPA7tJ2Unm2X3h0V2SMta0CrzzvXhZDUQx1WdGq+KpwjjUiK
Sc0be2kaTlKHaLOfrHJ3g69gLAOrraY2CakItd60/9xTNmnDvYHedGDBtXKNJrZI7HXU2kW09vxJ
mcx8HiHJ6vClDcaAkU5jTQT2pJqOlW3Kig0gz+LAXz/r1itW+76SvxqwjDbw5gv6chZgVfdl//PR
kqAzCGzYmnTozGmStnAFnYkMe8d5dLqq/B10mEwB2oOY3lHNbcw/vDXmeuNIKj/3+k631C/gX4zo
70FKgNYAQ6EXFoH46f0eLdKTsjBVp6Bl2ls/WPaT8wCM+K/xXClOxa0sbqzHcXKqUzKZRP1v4d3f
GdoIcu6OlToRNtRAqTjn3WDwfVf1BVpu+69VW2zDXbK4V/CTdLZfhkTkCkct3OA7bOv/uYaQQ6HR
e7OxI7uTg4olUHWnJsD9Tjbx0cBO7sW4+auIYHPhpzjQ9/YCDvisDy/VWM0gchHjCgkzu+16bRUG
z+rJzzzn8IltZjTR82F/NGcSeKhvfe2I48YJex8fkHnIs+ayRjO7iHGi6MKRz+OTg+78G6HLpM0J
cMAL9rSUYl8pV+uKMDNnzz/T1jj4xARCXUBqOoU1VGWp3W+eApyu9K08jLXp74dzWV3U8NuH08Mt
mVv7m35tDaSIt1fuwp+el0wHslEZ7tffh8ilZxoNntH6mcGkUoenlfvaF+mndnAJEfdEQne03pJD
l26k7SW39kQwHyL9e16HB0w2SarkzyxTZhcU5U5fGTN4uI0SUZLHLvlHie8eNH5EHNjzdxLMvpXx
RxVP6TXqzuMd6qNlUSAMnkko79+FcuVT5h2CUXGt06ZjQvo48VaD58HZ+9VpaWox93AJD4Per8V3
1Yd+o1RUuNw/xs00wAVXb0qI2kZ4eS6wC/DVjO5aT9pGYe54ARr8zvVO6JWIp1375NSSyOqK57H3
DOf4jwK6CcyL+wHczQEFpuoTofxX2vtHSD5bOF1phpec126NOgxph9hpo8jOXDd1syrFUEDYjcy+
Q4PWp8siAoPAGOsuG2kX0/ALsouriRuJSfxiKFg5yKMA7m7YqdIcLKZc7X8IoDAOBXLOspFHNsO4
RcR9NDgtq+n1Ykv8GibuVFCDPMvVZ7nydfPL9XyCdnW3cR30NG9xQR4qUqWmI1c0gIdHl7CYyC+b
2KbnZ+bJfQHTrz/30tmbLusQtqIrzbgdnEV0/DiCs2Ue2yvvYGZyhdrd3cElLvCIgMrJCqCxRltn
br8uwZyx5865nRKacWGDohxwviLMVNC7au9SzVPtNp0hCEJP9d24XDRHJ0AcQupq6lpQC+HpFZ6K
gA5cL1Xh9Y2JUME/SigWWQjz0bd84wdjH5+KGSY+Uf7G81lLV8PAk6bt3ywR5/AXeZIlT6w0YLog
emuxrNUjB/eu+xLtbECpzT+M1/GlAx3vPD2t4uCAI+Zlgd1Py7vYBZUUrlUReZngLNS5UylcR0oP
6R+DMtd5hGeSeekV1H5w3u35VUxsRWE5lrltfL5DPRzThRdVN4f0+titjkTf0sCMfgW55UeSMRmq
gFfNh2XYBJE04NS1xeU8HTfUAYQAkVgJcrKdYO+eSxosRTRRiL2/HTm9F6WkEZHeWP/y+aUvQijB
Z/PMqNVRn+pS3oD9xPHC0dHj5jE8EAB2lE++998QTHGlxsSucVBWZ3ZulZHeJKKjM0Fibapusf/l
Il2KBF/dAzSDVp1mQR7AZVn1uRsAq2QmSA2oKVJvqg/Q8IUVLKoAe9i2G3gj5s1Q3ElVjYJE4/5r
1UfdUTXEbXoQ+vpfMzEGw1SCZ4pekjn6pxaGVcQVP0QvFJDVYO+LMN2SAb4irVxo7lobL2In+GyJ
FQ1WFuhpsonb38vmuBw0FIia5qqV+Y8LGB3AcTfKxf2XO4CUE7EB1n4xq+uW/r5MHgQ6QKL8akJk
gGEOAMhoEQrz5dt3nvHq1MJI/N2wyl34lo/rAom0QTsPheKpcWwmSowqtAJ42y2DAFeSL6GkpmEa
e0qsf8o7YzUvB6H3kI1XguPg8SiIylU/mVu8dpjaZMu1C2MpH9wEyZbw/uluSj3s6vvFU5dFeUqa
AcmIhr9NMQ0b0JI9aBW1vm0i5jPvlz1Q/mkvQ4voZA1xkPZBMW3NHCMdA0lIcJDQYD/LTgEAD3HE
oUsQhyvuM5TSq8BvzFdnn3W8/PThJ+KXSEzj1palvM15q4IW2PG2Ii/A0JPev6wb4VJfrAvMhiK5
hCDhjMNaZoJ2Kej+BAb4M58NJIoQcWvrLBSM2Xum4xN7gnYmHFunoP74EaD/k9L/VhQaUp4MrQcj
deCe3Uu5SpMyxyFJxB6NIkIB7AzKeOCZVqvPY5jL3T39X+R5bUyrnCgpVAfSFSSvb6x4fTS/sx6J
C1M2c6jNmrR1YCPs13oLnaGm5WD/9h+K+Ve5ej6Di9oprrxFzlPpCf2wWLd+RA+L2enmmFSsOPeU
vDn3LskJlNVE3TXlRtzmOOzG93Iw8NC1aWiHG/ppbVW7i0i0eTXC7UuBrnD+8+pvGRNX8WOijUD/
lN7Mh3ZlkMAUBhnCOCJGVolw+W7aIRN2rgqISqPPfjKOz80uku7B45Qmz2BJ2bJRfBr7JnEhF4D6
OQz86q/evOL3gDHVqwVde6T9nCr+LS3UofG0GlzApBZVVZmBIaV/WuTaUGT/R1wrbenWOS4rEWec
p4V7j23qo9ITsAZ7LsHhRJGgAr/zsn0fMYvL1itFrEQhMSyxUuu6okeEXHvL+whOmRYKqsiS+/9U
M9TAeexgy6CjVlEiJRdXnjCFHxYaYSIeer3IwZeGv45C8YWr6+W29cEdYtfecm7BavSQqN8YVljm
sASWlEyyk3dicZ4u7k+9qrR+HZDkt309t7DEEUJIQ5il+3++EbMq0V6b75OBK5unpXwdZ3kMHE4P
BIReJeGpjek4vOSCPxeNH+PKPsbcJ/pe84Wpfy72KdzFIY9B2vGVXrygqQ8GdByf1W+DN/9gNpy+
0pmQensan/m377XqtezgOsDZ0O2tFOGnYLDa127k1oeaQnRwxGVAz3foYf6H//bogxKqN8Amu9MX
hGBTTkd2mtKWWT9iNDa1Hy+gl9V4hw0ahus2QkGxQmQQgrKwB4kRADNjMtiTX4DKuIL317ByNXtj
fM13168901zOxHfkpBuxAZ1gHjLj06PDq6nWrYZ1o9sthoZDOTQJDi15G1/dMyeB+fKPOayQhlRA
+L2z4CR5PCyQhN2ZRdBF6m2R+3GBfrHKReEwdJelSkyS3uH/KHXyoPriAwy4p6YmunohVloMDvv3
Uq2tb15NF4U24rxqs3Zm9cH88oXIK6U83IjHLzJdQyi0Gw5UB5xrjFJF45w+YLO3Y1uwZ6HdTsiL
i7b3TOBBRWVaQOkI4wH7nfSXkwb0svTnzTslMqzNCyrezzfq9Vv/BzJEq2XSK24CodFj7XY+9kcW
h14XNtNvy6m8J901b5jlqQeFLMykrxvpfvEfeCQUfQGUR2q4IfWZZAg9U/28pvXAw/HAmr0tRGC0
flokvtNPUjd9g5KlCQEPF1HkULzMvYrYvEyhhpBnEEP3xVw5GxOR6XWfuzuecuBtkPc70ymIlwPw
ewCXCcaFkMbEyPsgCwDlfFCgCjh/H4km7QC5HYgwMq3wNY0uRu7gyw0l49yHBrNW6Ao4NFeMlIYQ
JVqfzKbZ6Zpl6csKFw6W0VyqW1VOO1MRSRqwhlFWeaILH2UOmQhNEgnKi3JZMP9QdSRbtI+cpy7Q
YkAZDSBZIDaix4T0TMzn1qRXxoAWkM+A0Tv8GIHTWiNZ3QSnTr/wMXP+u/R+T9UGs6Jqfuo2nwcJ
QqWOZAw8KC8cV/k0RNFHjv5LI0T0Xkv/q5luKK8frIfM+u4KYmucWjaS+cgRCVRXKpoL08dH+RNb
PjOotraPu7pUsdvrZ+PDosRPI6bN/vrsWW6/2s23Xf9XpOELogHT8FRy0uXAyErNOOBbXWfsUXtN
Gegle+MUvnEB2yfiM4oJMeD3/YOPkzNWfV3QzY0Uaj7TxwA3Q7nK1keChFymQH5K3yJEVDBUJqWZ
IDGI/lDYxo+vgl4ft1YfFdrkKRV7w+0xE6DMnv1XSPD0Ih6oICuvfFzwOsC4qbg2QdS6DLFo4UtQ
S1bfRz3d4qkqtMCrkyjENGV03LoQsDj2vhy74OpWVb1SgoDK6X+301181jQr2WykoUWF+SuK20yx
btL6AtwMk4mAMVB1KzS/xYtbG/0rNW9j8KCucF6EfhNxm3wd0XGXVP0YNn168FLdjo+c978BFWNd
20kxpGvd281lkICjcClDZ1YKnhka3/ytR76No/FO5sQWYOSHfZr0IdJ0vMq04wQ4JN4yccYU/BIk
4fGzbVQOoSqD5LAULu8BNzkUP+6me+GSvOVqbhVGHqPjG3hdyxyfbK36ecVOLVFLhJUVJmKXpCUi
Gl89YHx0HaY4/E9CJxqFnZuA3FJlr0OJbcTPantA8QgWtTocsvYPD5RBYriOw0z1nm3pbZ3brEJL
9mKCRaAV3K+Of7Ym7FKMtK8aZeOv9kM3gVadAFqLC0w3Eym48zJdPMZfHsYtH9SOwnik+C53iAwp
ngMfvG/ktU4s6VrhOpo+t3lR/GDedv/BQclRHbHze8tWWWYCyrpykxjmli+TiVYbXFSCQg/tT605
ItOmtPQp8/g5+mqXMFHIM7953wkcYt0We17UNfkx46n2idtJNJIENnua4ZTER7JGCTvNASUn0mSB
0hRCOoBJuCvd4GPVFBcBWjp9te0/yzJ7mFHEdovA0rlnMNoaXf16ep1tmVChiMFvEUYNSzaNIU2O
yJv2Ag8uaiH6Fy+tK7ozj1udOcmD4rbGJlD/bi20nPsY3CtQWbWy1zk+b3kSd6Vdp1lfrgP2dTCc
JPeIfurDkDwcJLtQNkRDwXzjjXJN103n1eIAyksxSIxHY/y+T/x7Sow8K1RK45LZgwkhym55aNam
st0HHLmkHnujSiy++/fcZ1izz9iGgrvYXQqJxtQWe3wYBfOpyz6lTCRCCrKJk/MuYh6m45z807Ma
MpxGkCFm9RwnG7iVtiLtYoWk2ipBoESt0rxvquEvJPmvUVcQW4VDuBIEDhoOMYQp0iDsI5M4GWHz
D1wBhJDfmKsshWXrRFnF7hgIQsFJWAPGcKHmP6byJOnaPDTYSbVNpihJq2OzKiI4MWRilpdGlW3H
xAIbCk7X4bEXGGmKyPrwZxYQKNBEWYcwWkjmKlNGiHTZQVEXPhEfF95vfwEy8DltR0+0TUpQdfRF
cnp3fDzMiyZU5lnei5cacqR7p7QerO+2eEbZZRKhKghIlgnsIxgDaibTHcB7ihi7VNofhQ/NFUmw
zPjKAU8fYcggkc6MFYeai7VvcTvxPDSmV9CWajKj6Y9Mb2Clp2um43DMsNFb/krFoKdG6j7YSfWy
Qdv591F1JJvJDrPkmsskSjkfEEzqxZikXJvTdU7xBfnOI/fb/2d/EtEV8VzLh5zU7vKBHPnhDUvo
CEgtxQnsdZi71v6fq4JsdzCfE54UF/H48s5NNFyEzQzr5nrpWvI6nx1qHO4P2wjA8v2jmPcwKU/k
u3ZiTia2mI2DP/AaPcld6DXn89Pm2kQb3yPSNZ5cDvMZalw+eWEUG6hTKRPvF51/MG3bnoGjDgKl
Ww+udeWeVo2AP7nY07wu79OpXdfnro8hhlWscpR7knGXGMG9IgpptTy4mfa4ItrR21yaczVdpQ8U
stIlHJ3uVXlPEeyuDAzf5TPzfUZpe9VcqO5Q86a+luF+2z8ggoZNOtH8MpqeqaQkYSQBlMmAft24
92oT/RzmCIMH7kuBRPjUOJB9mZaVIs/5UlrvEfuMnUd4NX69KZu6nVYo98njVFFzv+Ud1Xdw2AqY
vQdm6cVom+Tch8ELKNHC8n5vzCRTJhC+wNAI4toxEXQ+ovkh7Y55NDsn6fXpNvDFywDAYHaxN/30
Vzv9y0BgHo1rQqKa522Fhi6jQYfM3ypB3WDRuMZvmysrSy4kr7kggmWHKeycmW/RM/QaPs3ryW6c
7bJksiFaFZv4ewRr3Z02xFGNvtBVCsrUkh4FT7r9HGvM/bSJz0W3tM8DOga+IkqAk476at42Mf4p
1v0L+qc984XGnY0dAhW1RXe7ekpVoBgrgjIYuyNMY940rH09+0bx8ekmefOupjA984d6XAq1g/R/
d0WPb82CfGQ2qWxke0if88y8u4M6lMFPClG2wOvOgBNbZxOYfeOpSfNKndNGsU5E59gZdP0RrUPj
81SG+VetdxxPbS1iWnddk9dR8mz2d+AM9f1WPbxN9nK/Yye+UiGxHPyyFQVMey9c6jBXxn8Hb6ZF
sfpX+d0jrcG8ds4wQBP2v2C4tCnrw0pPsJZVnaga2N/evn/cieuaWKsg01zIihpsjwMWGafk+/YK
Z17YT+g8Hj5RM7nLNrK3tm9B0OTx/DbqC+D7TcYAQF1c68D6QAhCvR4wvC8ytrPgkGeNubivgODD
uWHoUPdqzNXzY9k5mKY2rQqW1Z0AghHdTY+W2ZuZuTbGnN04zqy+vFyRODuaRtDO1JHUyl3eshpE
KjufOzYcwU/etYWXfHRELVRxY8gejMmDbUQkIKsJ8wtpTsuzTg/B6LKlhR5GV6H86uAwIoZqL0rl
UFf1kHoBeqfvGSHQ+AQCv26vWffdED4nfhVdMWwa2qnucxJnnS93oUSFyfdDEOiFrICcS3zNxW52
ahKm4BSQArc1MhK4LNjhs6H3Vq3LEwxghpZ0Cc7BmpD+Der5ID5sNO5v0HBPEtjzi3zgtAdLIX5B
oj+tPb9FXIawdCkj4SVGkTrGYj81rX0x0hAUB6C+/4n0IYTkfR1yNUTT44GAeZceGzQENJ83WLwk
tuTWgXA7FmbFw+cl40o4Z49j66lusP5QlGMme7htvrpKE52eJI3iJRmBySH34PZSigZJAK1hEPPb
11E9NZOHBvO0BIxVc6kcnkVfDaq3n0iDyoRcUNO4cb5js83KIdcPoSfTjlk3eXI60s8E504qaDI/
RqK6u2gmqQxARMlZvzn41T7zAAAPK5206Ra546EMXC265JOfCvWrGSlMLC9nknsVdWC0VcPYNL7q
Uo9FC839C6hzivWvA7W04XR9jC5jocdDRugfZ81S+n21vM5SgUbHkGJtCZgX3f/N4l5zXLfwuJAj
eaGcQnmqVuvrwmRo7CoWX3D9Q7+ODrJM9gpVeglCiIFeopvMlTRUvD01psb6LURLe0BS+u2GjkI4
bqQ4Nv913rSCkqAwXk1n49MCYfKgA27KZpVb0kqmJa+BL03wMrrupIOiPQO/zGPKOQGQR8Tc30HT
e+Rg7qzyco5oxzTbnTnjObjk24aBw3Ko3v2Rpkhype5pmL9+BY2Hj097A1+1pzMop7kFmHFReCky
RPSyC+YLJT5AaGGht5odAi14Fk6mNOM/95HXCtkU3deXpzM3cl4jsW3Nj0WkFrIFE2bzEk+0pcFs
t2ecHAyD3AC1BuH0WkB6tyGPgoScnXQ9BMOr2DU9PPcXhESiG7RXIM0aHAy0ndGvug5O6SF8ttoJ
s51M4Haq3jTtE39CB7iVqfRAghq537+q0gU8sr6Ia4jIfempj8XD38KCDAfJqwN69hMq9pTO2i2e
cpM4qBEuR/o/qbXt/MBSajGLhJBsxItRhQ9VEGBZbhHlQ8AXlGxxwISuHf8vdvZn85SBDgnKtDQr
tQQefVmme7wi5RP0mg5N7s2ztuMIpxSwz7UgRpbBkJXpzyRNjsco9mPWtido4Ql8D2/dAwIlZHjh
Xr65gr1Mo9RrnTDw+0oAKaelVEPkNMmy20nkyhNgVuKSuYSCFVsROdPeI9tATXaSgrhxM18BY99a
JvvFHiCw0gKR3tXFSsCryiVd2yZKQgUel4ROMJXfHREZtu4xihGHvzpxGWYk2nP85xBOXrNGrC0l
X0O55+X7k3Oq1hivpztAMaAgN0MUnRUqBwXeBwH9Lt7rbpCAl+GUsVJmHbymD7HLnepJ5nBMNIao
krE9Y3aebvPS3kueciYgDgxNyhalSIO4D4+BVhN+CEp0WvHHOd/UgC46bSPqQuy8kt33XXkS5uiY
DoWSgAxS70sGOpvGSRsoiw32Tbep1xJjr2868+LE6B5XCh/WnUiUzYz18FlKA0JhdzkXBV31Whsu
yqu47LGDQezQejfWiOXZb3+CSoTfM7Cs25c5gPo9IT0PkCPy75P4QxsOSl9ND4boht+5rpVeT9ZV
n0pHXlCdXLju5Zf++gjoe3RrGjrq6GehoyO38g5Y3tqkFAwo1MVnnnG1t8Wn0A5gpoPuu7vZJ2pD
wugWJ5g7+pA6xpPHUuAUOYACZWk7xlyTq5hkNRde/y0ADncqwp3QWeFcXgY7edNbOMGdfS/O5uxr
b1pr6fr/Ot9tDMdfvPztVLKJU4ajTN5Aw2AnL0D6Bu5lXQmBbE6SqLmKwygRAYmtGutk6Eon4o4V
zT+QCkKbx0iURwZCthFoIm5CAMNe0Fmv8LJi3etQGIDNMXbsLx3v7PgStKUMI6c+UaOPR6cqaFxO
Ibu5nw81L3KFcKIHnYk7rHSpT2f3/69jNu7ai3soId+f+O30C5V1pf9WuXcdvaKHPFenMN67KoEJ
ovzwHjSp5kOPawAW8NlgWkzVQQwCdXyV/zmz+YYhJkHNvvkzd0+2kVobmzE+nfnDPgxdt7tWtIcP
3ptLNZv7qIlkCWby58jNnJ0L9xIpEcEMymJtdj9t7TbJzIN4HE8EDA1VFgIYxILaFHEv1LSIWxyh
r+xJsLW7/+RXhR3qcPRH8laVumd7pwluvXd4AwMiJI2bvHPWgKG+n8QHFwMBNAERsEOT4AdlX2vl
Pbs2nKkggmQ443av3fkQD/DXnaRP66OGgV0VfJ3LYYyL4jCTuDrUbJ545Ct3c2+3MRPz5HJq6C4t
qIy72kj52v9qtcxoe2hqQqaWCehuiRpIb6KXce4BVrBFIZdrYHjfpux59alx58hS/zXtWsRrkldi
TbIFGnUxjaghYrpa0aOo7DxPHkL4Qp7RZlyFEwXAis3b6XM5XLeD9hIMcJ1kPfDy5KC7DsipST0R
vxZmQbddIMqLtPOxeMv5q8oUWcjuCuHNVMjAbE2n4FwZuyGqb2tgaRPYML++JrAoTKR5cxISkYAt
fy8xGy2yOX0Jp6ZwH4dsS6vaJuIQnBG+3AAcrG+Xx66GuViX+Vlrx7zVXEAZQd8n7C3fZbW0AEvk
Z4K7v02UYiR7BixIBQ7r+E60hboXwYn2Yk3Gc0SCQgQcDizPjqs1HZUFZ4EZtGUVwWQJNL+RNoEo
KL9aRIRSH8P+4G3XWgT5xFRg677xPvdnN4QTDCD++3W9CfOoXligWQZL5rNB0J7oajEAU0ybHWpJ
+F3YIMcAY6eByw1Cu4UX+dsAbWz7WI7RU5vXwpawGM70dQZMa6nqST15ffVCyPC+xUj13Hre/IfJ
YecU8RBJaQjYO3MxSr6XpFTvcSq2KbCHTTDT0Zv+1HivYtGLKTznzagn8SC5sgR7p9YAO4E//g/r
hP35bIW3zxDjch7AsCQ3Ib1YQRBdpqokNrs+x4BWQg2CCJH8hLHpFCFXGZ1G4edJMhyaXYUY9QMR
84B1cJp/jMKVO2fVuwoZBeCGpb78HT+8NaOSAZF3sfIRPfz2QSnbW+0RfT4zVKePyXIhRpJQGTR0
wjiSZmJx7beVeVfaxsSUre189xyu33jBBTSi+cs/DZXl7nJUCmVJb2jirDWuAWKRCl4OyaRWhjRI
yKvZie49Z8anWdTed64ZPhWg96ztswc3k6NsWHWtokWXdNmKE+Ar9jevWvHblo/jKxKIZZrCyS7Q
2c72uK9QUhzB724hb0/XhBvsVMGbKDqaO+yl4lTdxSEBM2JlTfP+vZCGcI+/zlu/jXD4G+MEtlCK
sy2D6UX1nBlkxgGF1R/3VLtt9Cdl6E6Ohmnde+ZX4tZSlzrC/MkACWpcgzjgdmnGj+PIJCmgAhus
z8o+ATkxxPISP6VlYg1LS+VAzNOX4N7M0eL1w+fNUMthgYD054E7bd6jlHMiEAuHC9l+SnFwG7sv
ViuYYtQAhnKwxYU3ll/QJVorWZOnAWI6pq/zorVRGlB0vfihtEcCOSkZ3nz11epVfW14q1oZByHu
xAB8kW9RmmSozlTv/tMPHZgwhwpNpaPQNzuXKxRkdLxKn8M2qG43g/12wsif3YEYpGLFd1kHW0DN
db1zRbuT7Zba7uYotJQkq64rMjsntatQ+gYYcFIlwM+egL9I1o+KPSngnhJVz7zCoUHbCtWWgJo1
hg/N/fB5esBh14WQ55rKtv2wOFJWZY+oYaphdlMNzFPpxXlPI7c7Ctn6nlG1SrchuFdonT2UDHdc
vrHl8CP69PdmJ1wOc66W49JMIqnofxHwoVJV+Ou7W2nbxROHXkJAkGunzULMfArgaR63MU+VPXSY
jKTuiWCs8ZuE5VtqO8bEjT+X++7JBHFMmPVS7xBZYLl3Wk39ghAoYFXtppmYiUma9yQAK9d5CxbX
WplbpMgX/E32+sY0tgvSmeFFn3f2r8l8N+CdriVvvoCtXaFjWwCUOXSoKwSlOhOEjO3OSpvcFhpy
pTFJw6NJ1L8Y8TG/ca9tKUESMHhbFD3GYydBQTzFVru9mmJkK8dC9kOLIyc5UR4jhL7IhmarKJai
pkXeCAv09a4jId/VbJCHBJHaX+LT6rofOr3sI9BwigP+yO45ZuXgY4aRRbQZQLc8kRFNvyJRi9Dt
1nthYKaORKt4kcpJdvYdmqO67BkO19tOFaX+b2wqqdyjN4GHO6YVQfpw8RddkdoNR0P30uFYbMkp
vjAFZZV+Ef1vclhoS8Goe1jqT4iV75aOPowa8ARBXAr7RMAcmtpEPeXzws7RPPwRtfOzguUHmYGQ
HiaCaPdYA2BSO29ugdJZeyk9lkHXxx51G1FH/fMM8YGm5vVIOTGLBBgRksOHZtDEogfeTR2VaumR
LCebTz06G67yeA68QgEf5fqbRz7Nej4S8fJLcsHx93dq4oW1ym1sGLjPhwqFR+yZYsxYmUHEsmFX
Xh7bKZvl9pMFMUXcR5eIacSdcx4xs2XYQ78ar70PACKqP5vMd3xLQiX/6kl5QYX9DhtjsTD+WBwo
vz6f+GjW7PyvRF/qqr4Y1RZhmUeJ1F7TBV2ajtQvd5gXOFF0im6x0iPY/RbRhLK73IlJBeua9feL
fou92QIfJ7RL1W4pVrEtdWrgMyt2b5Dh3r5bXNEDt/iTJfNNLCsdGvZwySljk5j6B1OluVYZZDZe
N7d+n4TtNGFY+k/BK9cw9lY1xzCa+k+pR1ThLqN+aBWxxl8J6fGtJCy/bABYzo9dZwi0sNJrwo23
7duKTgm8n20x1YT+xnFQw42+MZn0Xj5sWZ4ok8DgBRQFL3qUpD+vaYxk/jgKzw3kbPXlG3L2qKPt
weuKvuOK4+ywbVXmsx3KgCY2yLqTrF1t5EuZRgZ8Sosy32LJojEXquWZpSRHsI7yT5FEcJV/0ng7
UXNJN6yD/2q8XBkVLRTYnbmkebMPtOisWqJsb8+e4Jra9wRWmTrhu5oGKSlJ9rHV7lhwoh0G0G2O
A98TGJ9hW0zImylBvt43RdiDlQQOx3Te51821xsKqYWWBQbFohwKgo+as47R6Lu3L1B4sqFFLo4D
JMqBv2oVAJIbFKLDcOMxB1XHQtvZvHl4qnMYXb67Os+2LGBqYI4up9iaSyK/Qo6vMyH7wKddEb3X
MhdvgVhQL9t4sZlxBnw00g+oMrs1IPersTfObcdJLIk1Wfose+ZLovYzrmF1XAdMxNaR5nYEnuLd
i4OO5nX6b6TPd/qveWCTDcMXZKNmYGpxLLMq/4mnirVOeyNco5PSI6HOsM6mSbjV34QPhVNY3Lvq
BOn7XmPrq92RVQkrew+B/ovZAe2mIX+YnZlZnhF7zKVLSnCHWQknfP6gj9twjVyYPCCfp5DRUcK5
iC4KwMbzPCsEOoa7PGM4X++5HEQ18gKF6CNlr5T3i9TE5zSH/xKsKM2DcNfAs1uG3BCHCUApTC49
jpEtCihs2SPJc3uER2+tQkXvnFHs9/wm+1V+iBoYz9AD/hSiyztLBVp8xMMQCvi3Ge6ZT/0XUc4E
yzima39yVEus4uiJGS8p1K093xpL9UvBklbW8UN86O3N2UIJZRCXIFRnuW8HZJnxFrp9YV3wUCN1
KHZyL77FS5rEbCrkefZNVXxHkzM22UjBEU7Wf9r5+ROs7biyZNHaj6IW5+3SvaRYT1qT/7sxARGT
LNjbgDGnOFrFgYjATwK52f8COQoIOKJ1clQPPV2O7jFWGhv6HW80bGttnjY+gh5g0sRApzSmmZWY
LWEfSwyN6Cyxnu+lw4Du1pnUk02YgXVVKzHtLKC+NEsaZtmYmkNtc+IG8lfvfbnqZyntLyN5aOzw
1qdaTOXez46u+p6jZdu4tSANTQL7FY/SNOURJw/NKQvWN9Y+AOn/IH2clC1sHZqEaOV4z5lMywBV
05bVXR4wGFJrR2cseq6AMcZ57zkkBxcMR8514fGlWQI8DqsVjA+aR/EKeuud2o4VBCHrl2rdSCHU
jN5jQ2SWTwTHkUu67XY+bfKW556h+grRy3SvFEcQDBP7YlL2T8kdSkcTYTUdz2Z48pNtMZs+1Y6s
/1zHG/PNNqOHWSrGmEw07AUiz3SG8nHREY/j/WJTHe8GvgYr15R0vBuvuKXs6+zcVyaRGlj2Oc1R
mn7SVoxfUaBumSFl3X+1C9vaMi8X+B86c5x6ysOFbHmdCDOqipDFTOb1WAoXwa2ZolQDMGSTpeBV
dtGRQRhysAYCqBFT8O7zGPYf9h4j5a2UYVVyEto/E6vDQfoCyjHIyleK2U3tZzxP1zSqXJmP6AJn
HxB7B9SZplf5cmhIDDKxN7VEX0M4wdr2RHW2Bw6znLRTIkUNp7ybekLJ0vrkDkF7ehfj3EXCQWkU
2poS5vhx9dcst9JqhZqLABpyqShaS2+AT9wxSWAcWNgucEbT+Toola5GX/UKAFbh9NA/sCUziEM6
Au4PYP2Ie9c1UtSFe+8rLt50ogTL1UVOi5m/C422c9gahGoCuONaBbf3t8LUgXab9xUfmiYbY0we
WYojmSXhL5h6KdNcUVKmc0VHLm8e+wssoFUpbYyILgC3Q6WPCqo+yhZ//9SwHpIspUEUsF6JzwUx
YbxAuVIvUrliG40DBpB8EgGrS2XpUbbJLvgzJL2lqPWm19qduZghxzcNW3MridpeuX+F7wuI662V
znsuOyx3SK/PxZujhVLzZlDwIc9uXqiuPip7fmRe6HTrNGc236Ulh5QBrmLTbNgxyVgyB6/SnEK9
2zW4a6Oang0VVICi00e39yM32qelnpOToP0rLisKUN3C8cb9AwxRSWiM0O9T58CqQ0b34nxJXdK8
DSkqlBSA/b9+v0KNcUXzx73hLh7G7AvkfCeHYskXG09m7pZTcXi3hg+PyDS8wxPxm3RD2OQg592+
mm68BN2vAhpg5qpm2yuDi2uzapmXv1oNZ0be6eDfAvoe51cA6zS/MxKaQ1B90q/4L7kf6MWBO7jt
1Cts5Q7/RX9QOCzYMp9zSPbKyYdBhPz8t3eyOQ1cBzu4zR8Z261WHAXbsZanx/ufJyJgyCtFClS9
PJprRLzB1Bq+scXuj7/YnlxLtZHO/XgQ0aosyQG3+XG+LS6NZoaOPDR8pnDnZKTPHIRTM1yxJIft
7E9WCB+ydso24qf1JMIREgjzjBJxtZ5MwSNWe+IZjdUl11dHZre6Nqb1LAjaHGaePw4Cg2LoPFK6
DRi+XRlITBfROQJE0WVYcHyqFBOo1cHlFkwC0i+6Uo0vcgCnLqMCjsilj27mrbh34BIzUQ0k5g+6
uUbQ9WgqJzxAH/AJjOTedJiQGq2sHYYuYpFoDzdRJFVpkN6DlwadOiYvSTKesy8OCfQQKWUl8RiT
ptlk1BiFQA0nXiKoag0NuNb9NnElOhsWbVzc5GE2XINH8kKOllh/cC227+dwOwiIaUa1cdyqLqmE
+s8XzFtt9oVAp7h2Pept1yugImhGCO++6EgzAMSnsJYFHgxr8viHXs95dDjWNohheN7/tEMHddqv
VKOsneJbU/3lrr7QvHHWrfobd07O2+TxYI2lBCCegQ/eb5q0l0zwh8KVoBoZPhZKwMsvFjzU1ldT
i2F6EwhvQxBxI8rp3quUf0QdNpoSBpMhefJqjsPgxC+hVwkQSVQ6ga5sqMT/LLMOKyLh5qGY0R8a
FgCW76g9ZNuHrRyFCQ3BlfPkXLC+Ve0GVauNjvmz5fdhTCfUr2uUDPN6KL0rNfhBHW+rQ3iYR0eG
bDx2YVteiIoGKItH30eX/QDnel4nCYlfLh6d2sguBEv3wDpjxK7zO//OklCS+ScWl4/g+x9/CoW0
LVZUQUb8yE9cf7RZRnzrMgOgyQoYEIu57Pm6UD1bAXFcBm+5fhVdPoo/aJWVUQYUKBBP+6teDGUA
nPgGAvON5l5oTwG9zmkztGdQ07+VmwtxkHgoxAACV3uJrhW3OeA2N393DOn0YL1XXK2N+gY9rXSD
3WJZXOiqXSviZZzVZUkPwg/ixufwHmBVBVvr+27Kj5PTQcbmDZZSmedCHQkoeSEOz2DreN+29JpX
JlZ1kgGm4o82Ok6ieloOTWCfQkeFmDPeXX3x71jLe0XWBpNnVgGeU6BWh3aRzJ31o7xxEehJRr5T
WDZiKY14fREyzhC4aeZyhIYCi97PIGAT9M9gLoRHLn48Wsd0k3JRJrf2UpugmtEsRiWChMLHmGpv
iimYsZZ9fTkSZeyUL+1cQm5y9MSp0/LrNnyFlYkdj0KRCq7IThlvkGmA1Y8OMgHYF/W/oJM+Y/bT
045uMlQJH4KIG+ZQt9MEWYv45NFPwQRMWY0shE7t6t5kgu6ni6rIADwok9o/+S9eJu14XR7MtoeE
DvqKFPns5ynJFMQALSqp3LN3ZhxjtB8sYOHM2JFS+5nfRQmVZy7gIIGd+t4lriy1UXfdrx86cQqL
5aR+2aLYEPQ3+puyZCgg+y6kr5QZrcRCIM198Y8KBSZDoZNnshRoR1OVddBPVRLBYjN2g6s9VWLb
yOJHt58rt3CNEMhqz+ir8mBRrbSiNzbYkMi1JRSK/XPKNMl+W5iHDsZXYo+5Y6ir6IV6NEP77oKd
vPgGs3NPDBKAfj2+FoxVTPEjw8dAewaWierT4KkSBezF7VdNWg1OD+kId2js1R+jTFnk+1zkz5G5
b6rzE20DmBpPSvxxWMvAVsGCtRG1NII1tShZ2mPLHrKaOe3cSSyXm/V6Ndj8wcSwdl/klAtaU7/i
L+6uotk6Ptrae3mN0KajCE/VsqKkPJJ8vJNINkr3toqYzlsUpE5ou5RpKIgrZ8EpTvD2XbqVfyZz
UI4UwIz/9hkxN8dbfRzeJgAsPbypPYa9Wpq6Y645ttb0g1Oalb04dEPg17kzcVHs8Zmp3etTJw6L
2ueWepMRMxlJw0kE5Au/+VJ4qtG/7lOAjfoTN8j8D/zGJIV52Ch17EyKdbWYFE03O9uxlTSVFEP9
qBJm6iN05cZPk7csETkjyL3FiYchQlomX6ji2ErBu2BMYVIqyiTkzgpkI7yX8Hd0tB2KKLNOxG6Y
PZq6L6Elh2VO0xAy02lbBdSHjmR3lYxxV9EzcNKReNNdz4p0y0wgvVPr0vPOb365ot7r1ajN6MxF
2V9rGMTpEAxR4d9pL8kFSlqxGyKs2P/2JoWO+Navuk8YBmnIo0B1iryQ/GdVHR+ME7NCLM5dDqwS
A2QCL/VcDsgfmnFt3wgcreE51oxWOsgcS573ZXTRVxsYidTcPv98/ep2OP49YbsvCWELsBea2edJ
qcA/Rmo+ZtInCwh8tzn8DmJK3YvgnnNBruGUvffOsGAU4LEyJ9duQoVJAqZ/SGSbmWoJwTBsQ6F5
Madhad4EIdMmlV3+odlLDFfnJS10M3YfOCNNIGwRhJ0qtxONF2VOv8eYM+2aEsOECvIUSEBHKe9C
e0EitOxeN1sDbbEBLOJPtu0PUd7iwveHk4aY9f7Zt0d7E1yju7+gK7JRB08BX1YUOaDP6BeTbm/o
eLt7PW/uhA4aQFk8cIBzKgSfpURtSsVCgD6JUl537B+2V2GM8dgzfbIkqhzUfL3qRi24bjqbfueQ
PkV6/cKDWCc4XaFmR+RRGV5T83Om0XpAFBTRX0Z+xEoWE/yN3bmXvOU1Noe+IvVvShmdJjrmn6iV
QKGS2w+Qu7RsGB4NMhN9zMJVxgWtzXD/28iVGkBzg1QkXMLqeLkiUq0T4VPGlrR5Ufmcc5slc9iu
ol1xhom1TaP8pXExrl5Bphh0GZVm52Dbgj/6G4uLHn5JH1PI8JXOxJRdVK47HIJZY6gzrgpgDiFx
NlVXmE6taNRawHzgtpISM6TI812drLcXGiSIp4IZL9z8TKooNh4/gKSS+I4VrFLS+rqBDdka2fDV
5+Xwak+LlI0aVi/PSTyDmC6SeSdlnmxYgpMoIalClmbaAQ8ZlZqtPUoT0Gu0CRdL+IpqN2GhY3MT
16hupPgwyqdZB1xSbiYg0BJPeNxoEBTt2pAEMqDS+W6NCEE6q7L13UnXfjleqokYx5TdvZiJiMfK
qMBWOyoHKV2brENDHidgpJ5isWA23pakJOfxalsffjD4PIAGYptonS1pZs0Or4S87pJEeYF7f7yw
eL9JfF2hT/KUd88bDr9yzUovjc0EdIm9BzLpg2nzjOBHypcKp6Cquzkbh3JThCHhehV5lRq0VaZD
1U3RwpIgA/NdSa1grtIoSgXTCkvDS7CO0Ch28IUFFT6ctNzVXrXpTv1/h0jrxRoM3FZnS038jGT/
2xUjBQc+hhl4E5bjD6VbavDZs2eOulQVvVT/em3dFaq2R5pbn+Wor3eNg/MhtLIeRoYNPJXgCrtd
Is6ds8mEHeSnHrNC6eAz37NSu/UFT2ac3/+SCaB0M5t1Q3DBW5SVLGTKhskeFmE2gidnZ5JZCs7B
xVE8NnrYT2r9OU17w1job6IyhxlN9eeADXtYgW7VgeUkuXb7naQHLK5pMEyWqNnHPI9PXYaxxX44
fqXI0mat6PIN240aV/cB1r06y4xtemVod07m98WlxqNUMa7U8pcnskTu5rAzQBNq0FBt9OYOfOpD
gfWyAu4InnlOQrtWMyQ447Q8kKuDgWfHnfsNf5VjNRfzkYe+2gscBlqbxzi6vPyWt9J+BL9uusuC
0gvBBUVO5r4FAbtrP5+a/t0GS3YcB/5f0Kmp1LEbCKgDwCjgPXOcfCvjGzWecX+f9WPdN03ubQAb
0oOprC45rHTeiAjoON8p6j8vBOrnJ9fUUZ8lm/77gjSWtud/MtYpG+xel+tkhLZktLJ5DvxKBq2x
KQHsUcbP7ns/NhDIjbuN1NGvJHwzrz6XTa2G8QcpVZesH/hHaInBUiB4eHa7/6WVrDJZ894ghOco
LUgYfn3rIYUOcIoNRnvaSGgDjiBkDfremQYBNSvfjth+zZtUg5ttuhYp2WeqxzdAeJmY+273nNfI
zKgVd/y9YRlHjADi30OZO2c+HC+nq/kGhXOiY1/WbTIboHjEv9LBMw8DgbmPGt2IeqsLloYqJ9O0
1nU49Du4IexKD389XTc4+AQOqktNVmT9AN2cEIJGj91n1TwLdwxrCtQzCoWOGPi2MKw5zy769RV0
FykrWLM4X4dUSS6KulxwoFjIVr9zdY7PiIqE0eYPyVcRIJi+zLELhDR9APE9nieZukPoDI6zP/ri
YhboldRN2sJIXzu6IoZdWa6KmUF/EBfHeLd9vtEM589gBAKlCCoLQM/yIf+kQ5VPMRTjuMBglunk
9KXPHKZprzoiw/UMM1P5EC3LpvXDPIx0bAhp1JviDH2B5ufrvJI7lbBL9nizD4YGLWx1QUkrWO9f
P5l/vlkB4L/mz18gBwOcVq7+6707OaW0dHtjpvbLoEL49rjMoehUm22yih99Vqn/0Do8ZKcnwu6Z
TYdGZbNWIn8FbZsbspNgkKMiIMHd9fRbwqy0nCjm5U+GBjp3F1EExdLIJefzoR0NuNGr9fR3YiUg
QXL2bymJpXaEse/NEo/QSJzfjLGkS/rVgtOxEQBhw6ZVVnGSk5t5WI8V/nQtlRUxieohGRXYPGcb
J6M1nZXMjARziGCQVlmJ0QCzz/JoNMv/lMoMBK2IBfdrEC3n7iTZjJUpehfiM40p4swqJnLshE5M
YrIIrhcmX+HAog2T3hk7yhzZDi+i32UJTF4+M9/VVnva/GMQnbfTl6qwnIHIYshJ2GrzDaHvh8Q/
Jz5lyu3YMeZmr6kaG30HAWSXO92vV917jADuJPxHGlbYkBgAi09dRRN3Y9wdEtFVDIuWIkBZBu9K
kyLKRRQ7QLKsQqrFDZ+CxB5e8N/hogIb3qNO0yKy9zksVbLDsMYaoXPTTV7gcTgZoLsQ0rFc4pG6
HOK64/PLJLO3klwpbErQWLTI4ItLO7RlraS94g+5RrXgt4AjDM/lHf1EcN5Ak24yKFi23J4/5iTa
N0H0tmv7FFSGCX6iGl/yKipjxKBK64D2CIpG6Aa5WOBIUpy3F9gIm5GQHyaipmRUyfQka7w+w3V0
4xXLhdgGfVKJF4GcmlzrHNpr8qm8MpGw/+HuwcC0Kss2ZSBTRB+iUheL05l4UYTLXrkMVkezDItc
dKrluvoporM3X8Mwfa/RebQWA+POaqVkPl75NfoEUG7QHl6LEZB2gcV/fyN+TKsv4AUBKJe7tTDZ
W9eaDAnk0k7lkoLyQgEmv4q4mbLas27WOyyFkmXgdNCsx4jQkVYBqVJ+X59Kf6y6XRigOCR81/L4
vmrAwvVqROXBIfI7nTTAtPuSL5mpUWGoOPB/e29xu/MAEj36v+XIGuH1K416QrmAdstQ3CFaC4mp
KlLcc8tQF4MFSwRFhk/ExbHtHteYvVXLfEMv17PfmMb0V2oWhYGCI0A4jQc/gXZBwh0OB5sd3Vaw
z3wMcSNQRMTfBbbssuNVqPgu6wG21VD3xHCs8qnfAchDthOpxempvURrjErpXiAEYkUtr7yQNX5t
5CDpE10xH3wDxWQMw/e3l2lUv3fwC/So19I8fdtZtnFPYkm0eptNJ82GFfbK2yOJaZopzvLsbxzX
fi7yhSMKpwm1gDHQSogKLdy/5CyLzLqYqE8v/BuWe5KOCZId83QoImig//DEr4qxvv8Chz6NrG8l
KJu1xGefhwkcVm+zVe37naoLxkmN8mtqxPXadHjn4Wi34qh/zZj9FzA/dNcNtBSCYPgy+T7ekPVL
HWTnxCBX5kyQKBwqNXucW1Cs7+vz9J2rLx2NB603W7XNY6pSwDiscgx9BjrKXt9jw6ct3nEQCCsn
xkd8zMsR8A202X1A3XLS0fVZdbdIWwwXSFETsOQs7tvQ1gMvIkQTsy19OfmiZ89ZeHG2AFypef3W
J8NyOYPFF40vtQaUJuQRCeA+LqfghL9GFUCSW01KWwMMrPVpNpCJxekNC/OrgdfTC2AvbDZN7VBm
WwH7qvn2lTWg2/xIHAXXz1xyFR2USjs1L0uNxbIfxlLUs70J1EsyCtgA00gDzMUbLssjprqGGSUW
R/CxzVZ2W/YlK2GjNwLeuYehrt6rHKKU5Cah5ya6w9XnQLU2ofdjvVrEgl+ObY7f9uURdinZKunj
MAdv7neV7mt9qGidesKIsjdD2hwjTqAs7D5Dl6ljdVRhfIhRaPV0/tqUjFXgsbqEl4Dkl3EcMoG8
96f0iq5fEwuyD7Acxt2ig27EHZxe3o5CPbsA/yexU/L47PeBTCfkyKVHKcLvCbOVQ/Oi3/NRFHzh
DXB5gDoLGZ2RgUDv3MJaLQharvbDnHkKt/ELBuID+BZgmeaPjbgAQKBOilIzSb5w7F1HLjn71cer
3AxLcb4dtyXd3QveWc21fGAZu0Ta3Au2I6AJDGGyqUbi/pp4txFdKNmBzOC8H2pO4KfyrUFPHu7S
dyBYFdCEc5re14V/dRDAkZtPCJfidB0XeC/lnMsOMd8XGed9dkRZFKrRbXfv3WXxQaE6C2kBTbPK
zsOPthodU+UtL19saeBkcxo8C+JbmKgheBWtMBrojL88OXuv0NO95CSUvclouhlk9vI98PzsHVPw
kr+PEWjHdxh1OE161Qc1LvNrdyZ7McqdmJblzyl2dvNZe2ojnesZzkuzJi0/egcbGgWC+rEPSnpq
Nub7uYKn15GNWUVxLSBU7bprvoFcz0eS8nn2uIk1OHMyZi+UJqloDgPpQ0ZoAJzRFG8MkKq/bt0C
jcwsMod8dvOEsTf3IgfAqKeYn+ROPZzQSTgy78FTpJuJ2QzUFCREbSK7BFp1aUyKESuTm4bVZ0AW
ueOTGERR/eapTk17BHbRbHjwnhLe+MsGbqIy4haywXZE5ZGI6JeQpaHLEvtsX60ao4dh+IRGZR7e
jMR+rZgiul1slltMrk0qbElNSCSruNOY1cNPLFt9A2sXFW568e57h7hYJkrak1PufbvIBs160Fzy
heQ8IF1ZJ0+i3rJHTzQK1CQRbHMGQo6hUDAlabHHzAQp9VNa+SlQjhRuXyRxe0T0PoBpXT328n1g
XWj1y/4KxOKjrYMtILFYEqkvJI1gtlSkiek3qYzMplnC4j+Zk2I0eFHuQldccq0H0PM89oqvvPdF
Pqi7REr3NGJN9+/qdPG1ieCewpTMhnf/EwRjEcx4lPMBZkPxPeYJgfIxEG4UFpQEnHjj5JDbxgD6
uCjLhkKqH/CM29n4gKsqSOaSvVs+BOQGrZuSwYmnsFhQlfyp3FKH4jFRh/9vhOGDvfGgskUVs0I/
UtQfPSznp6/IhK6JutP4OIbGdOYArOmF50IHNoDyPUEFL84JOrJn0+C1GpZ5/T56JAIrUClXF+8i
+lMClmLRHz1GK5LIQBV3LQD+mhCsLJKEInUh4FFi7rFQ0DQFWBfVZ74UBMh6CflwtcNGNq+tYrPX
mHLbtsSWJpxNzbajej2lPkyszTRtltIAkmDbXBjywk6pDK3/gmBGmE1VdlRk7LJeYMBC5Y02vlrZ
/xpfPoCf0twyLF9MY8CllXCDBnFvNSyCCnnEoTrz0iRRmTPJm49QK9Y79RZVmvAxPjmiZKm8bqN0
qWMYHjY7OuRIM+Rq6ilTKhmDzYdrGn8Dsk17aWc6uSHWxuLcLX5ASrxZ/NdOk5UmiV2vA+h7qtOY
DMvEt/QTdvBGIQGfWSOmg9sLsMyuY5LAnTTOmWxPBgnMgvNY7KVCCuMSltN9Po93PcPUurceUI4k
/2eLTv4OEzX6/2wH6NbAgy2KoRjfU91pU7KpsQGlDidkKARtNRGc3saxJElneU7myAYYcmerLnmL
LsmCN4WTTqYTB3NcZiVRhSR5g5j/4k/eakF2r4pI3TsylNBbgi/ET0hkATiQXx8r0NjwSV3JQAbP
VNGRcOuw7HxiBbDpIYWGs/f+W2aGRoX7990pkTwmywCYjtsv3QlunoCOop3eHAdop5S/lDIB7epv
7UWCfvgDtaWKTp+Of3uzHEqosMIs47V5oSp3hq2LxRl1LzI3o3xoOboFCVbw9HxcPQJIm9yE3t6O
Mj3qBdkBON3y67zqsdLp6/npKUtEJq9u7BaMe+yq2h8xdP+Dkm0sce4E/0NtyAjfVl9YH1wFCAyS
eKuYzlwapGOl1fPN/xJcBN9E9czwXSzkHuwd/VWz84gS/YEz7iFe+Oi2gg3o2zFG7T7YiCLcuTFS
F5OcoMlrGILgn1ciWhgzkDnBFCK9ZNDCFE3c25mBEMvSBO0/+9wFhhby5G1L1H8GJjYT6AUrCvBe
+F/kuCvsORFHgHmtAZIfg/As8Eap4plfEEZGuaVt+rGHAqHGQbiNMAtrf69NgY5sUxloNCjwrz15
/7MOAOSJu2DTqkav1rs1a9132A9+GkIkvxwP7WXRRxhF000ehl4wBlxgHfbZNvn1tY6Gk8X4yr8I
DM2ZlYHz8bAK5iJ62KohNgVPY0v8uUstr/CWUoBJZYeJtckX7mfr1X2ndXHXEIWHCmvfMsbummBA
FnCbQl3nFFCbVi3bvLE5AkBcbxr2uSDV2RLQfPCb8OgJnX4wsV8vMCvNGoc4Dqy0KHuL/jNG9wX/
qc5/5TTuPgBTWCY+Ys/IYsdpjPghkRlIZjeNw+OtsRimND7N7E0dsg8QkDNEMMt1gWeTBawfdP1+
GushCBjh2NWU8OCexzeO89hcuOQAFeVFEiOhsw5Lgb2g4WHcjlgdm2EXpVZ/+g2U0lGw+fj0YwKB
pSCQko5OUiI4NKN4nxlrUYFg+BLBzC6bd0OZ+cveWUHcuJU+KXF/hj8YSE8YLjSKYx1FRSrhl6d4
88ivrKXn9FWcvec2DZ89FflK8L02oSRvATmUB8DiSzOa/wLFJmogwJYHWXlkFP5mqMh6Yr38rsBZ
Vx41wuV7qHm0oFzVb5wJxDSk9hHk6HqIZ68xwR/jshDLCThAgKEYfCISc0ndVW4fQ8DEBhJKcyEQ
hmwHj2KsZf+DjhK57EYXVtos7ACSN+WHwhNmFFBFW0Cky1r1QZ2DxXcs1hNtJKGoWHu6/C/esEiC
DfFnCXKseYnACuCrAE8tkgVHkrhleS9/sElRWdZTts2DEbW3aXdZ6tjZ+EuwR2dI/6KNOE2/oZKN
YEGSHI61Bq4n8FCE0xJR7uAiLja6U28yr3w03M3gx3UftcZVCmqPGrQDrhXGfv3iexr/Yiqd8fWQ
Icp8WU8pdk0hVEEQu98RdXLbSq6Zg/J6WStRfW/UO1XmEs/ljpv9lV3552RyK6LN9VbBrExdDgKh
IKtCfTkW06Pev/fyE+HD9Gs9VMJJ1ikxhs3aVVAuPWRkXpgKWLpqePGVvn+oHuOxK+NPbOfm55LG
81opH4TUBvMINveEEvAK2BTqv3R6VcvsP/DdjE86YTQ3LAwswp3uEeGlQsYMi+6n8D9HvwvYFPuV
rA5IpeP+oiPn2SSYtYLoXTO3vOhR+NcktRO9JLKDGDCgW+x0fggsI2R2zEmum7PFO1h+XfiCDV2V
3nXr2nyxzW9thJDRnb/KQO/SU8kJmFZhzJtrLnGNyY+aKBhTsRobF0s84Iv1ciyoj3YEg1IlyBdT
zHZmjW2Mnk72iNoO4l0jHY6lWfeJmrHFe9r7XBbWZONyuh86X6EQUhgims5xZ0lXWFAdDvPfY8lC
Cs67F7iMitB5UacPcY5wbEtf5BOYVWkuRn96XQVDJi6Na2rNTJgl7vTlGUPHcCQR0efq6rje+tf3
5mXiCFHgRA+pm8TQvUyL22PBoRGVWZLh0v2dwpVXBijDM9yPKFlc+Cowddh8xKw5wYBLaguEGzL4
Ihzvvjg5sjABgdj+GlZSm8mOD7vCRHls0CXPPig7yeAAAgVqADWAzi0ky2hektNnNjHvERuMZ7jN
YFJewgWojNuBac5N2E/wxQxM6f5v+JjvZXi7QnDNtS/AMUVW0AQefo686mIhZruFDdOzKgTSLwIU
BgshG5W+4d3IQm9Zjtn1z5Nu8YNhhLbH0zionEv6/iaZCgcD/hQ2O7ZMqavujswINKr8TZnU2AHI
tJcSj413dJG21N2Yx9KJH2D8s75iatK1vaNAmWdF6Hv3VSp32iMX2Ke14gvPxis4+dlRJrRTfCjB
lW+YoF1YZlg7/ymPg/GSrn0nGfzFSowJvVfCf9kOkNlbVFW0ha6zmNwDQ0yIp1gXGK8fEs9Y8UOL
EzewIhPecBp6T6HnZzvAPN6I1AcT6s0Qv7JvqCIDn3OmLelDSL2E712C/BS5SnEayUIG7LmzvQxc
2Z39GPJSpcsnh9ioKuAGJGSo57gkRbFG6M9n/Q1+2gBktCG4EqroyRt5vo9auMhiPKLCA9511kH5
nQBJex3MTjS6Z+jdHYAf+UPtISifQJK7tPJXDaU+MTzWGA3lAsCZgGcKWqeQEOSX1NaP50yennTW
zJeo2JWFJpOA3Qt/dy/gKIiP96Omrt6vtt728qOaeCaExAMgfB04eb9v7NRWPJUV6C4BC6zsSbZk
+tq1YMCqjJf/W/Is2hYQjJlWrKM2P6lV+dtCLWCFtSOrVUsY7y1RwN3x7q/kGdDOOBLa1a9Uf3Tv
j7HV5fGW71ybgWDhL98i1hFyVlCQ/Oh3oF99RlDu9Ox7FqatuudluzubHBTj2xL0orgae3sapfro
/ifUjSzUjaVLeNQUvhOykIHVbPeYdMuAYh+GQn0TbpH3xsMUjnxiBNPsH+3Fn76g7KK8BGyKwGFK
z78sZjDQEZVr0rDyCacYu0UQk4eE0Zkwf5RAWJ6Htq2TYMG8U/TzSDouYOBO4Uac/3/zOp4fT4fg
Ea0WreFc8KNT+rhZja8Ikv5FV/Ou/rHrq2xNDsRYLY+GaPdVABxsocJCr6ObwiBLPqnFKa9Zt+oe
fnwlP191JagSoqdHSG3K0tfjHiWoR5GjNI4BiBFu+C1r3Qg1bzoc7krs9Gk4q2w9IX26BGqu0izu
JYOTefMuLhQtHAj9Ni3nXZx+F8JWwzJaaLOfIJxzUEc7pXLxDs7f8jJ2j8QkEKWElMOFOEyzm5yE
dOj1jvRAPkmhp8zZYHsNFwnjs37Z7+s28FwJnrZCw2ojk3MnjdEdFg+fQv4VykHp7DizrNbqmS7l
sZWf9p+zTtNKcZXQ4CicbPYjQzBbsDTJdvEGiYBMxdQoGdViuj66Jm6PG8teytCA/Wk3qW/6d0Fg
gl31UKL3w0R/QZTV1tHDhM+T724DHjlniEF63IJ7roOS6mkPnZdM4530R/Hl2qVCeblr7OCiDwpK
+MHHejvbJGjF0vwG20UgXuUL7I3Lju30Zp1BpVbzKXKLW9VQHAu7oqsqi1u1f1sw/l62dw/TTr8M
JpAv04CkeGcZY4vEXX6ldoXUKDjooPQ57cVMDVVB/ucuCcP+rS1I3XTIvIokICchmhArB0n6H8KQ
kiDpK7A02E6RhdxlVgfYSni1tiogOaeSO5Tj5Z6gNvc1VCh6S5gheyTOBc1ciQ292BfsrpWbjI8P
OlAT0uQbk7c0l4cLIwJrAGYtkj7SmnncdpMhv4aLRPj2JO3UeFjOvy8ShDWsr+KTwb0mHgSee8Wq
mLIOvtS68JND6aLKGRxEGQoj2H2dC1wa0asjEjE0mC5l2ZAZog2/PSC+8SAc2Oj5qVkRUBS05lW4
HFRaFqA9ITppKxBUz4Ct7bBlkTsMN9jxu8i/6wRLXNDffx7/jhYOQprNo1bwCA1MGUlzrOsPjPkL
ciJp9MLjb9XEMVTHnmYyEZWh+tUQSOvmPji7HOkvlt/nb4YbXBk+0bguc6whl2orknsM0zm/5Y5G
3t2x+rVNOl+FWudbVFPxVmeNMfu4fEkKddjPwZitw8re76EGkgPdzQKeoCglmPlLbir9G2D4Z/ih
OE1fqv98UyV7XZm0bNuU2Mi7drimoCjnbu7eNlJYe80vq4Uf5YjBpUdotG0Kp5obv5sJQt4a1Sxh
QkzNSFwIrv3M5Kt4iorFL2+DcMxH8ZhR6UiSx4EAWKn+qCf8Gqj0f1wyhiEqJj5Qbk+ayau5W7az
+dtfek21gVIgcmXKuptxyRT39T7oxZu9nyq1md8ZYgQ5KeC3MNlZpe3svU1tTqr8AN/CkwZtrbl7
P9VCB/eJ0ScrEptNIRoBBl0EWUXizziH2By/WzgxzJIh83N6M/k//U65tqegods2IcFuST4aTYof
DZSCFVCkuFGnJQ+qGHlmbOOyRoot01AUh/fPlLTf8ABsz8FtPwHH4DCpckREgiWMT/9J4K8coA/M
8gfoxUrR4WlT6QubCR4Kb/aPhJ7f5ConMN7ZCH77T9R1U6yoBjPaHGYgFpNyidyMnkCKHUKP90uj
QSIMjCg5EK/eXBcPIPKZECnon/qlK5HpQx8gLLdNL78gOJxnliGrt0b+hGOCoWRBLIIpxBc00CNR
/8b4PP4BCf1pO1D2fQfKD8GsqRiNMwtMmxjuqAjo/nok3XFHmxig/P5ONV/lwti1u77GV6onazWC
z5UJx1XKQfkw+vhdn9tLqcjoPWzha9VpGibgKw0QhHqNwm66WiiV8pqB+j5eK50NNJv5PTcbBJXo
YXzqTB2hCB9wwUFcEZa5lprUyKYeT+XKnqjS3TQf2axrhWrtJre7umVJoxmjKlJL/8RnrbxY58+S
/T5hvxFU/w7sIVeRUSbEWG1hsLRWujFEUtrorh+7Bcdy2+3y2d27JXe+YN3BpcBidhU4IzWRIwzt
6UUX1H6clpEoRr1qSAJKDvcQ59bV7KT9r110Yzt0V4aoNM4Y2i+ApN6baOxq9HMYm8ea6RIZaqpn
qLNEnNJt3kolzEqt4b/vOOWE2oxryXgZVyszW2TuQejK9iFyQ7cOf8FUu0IQPaumN7nr5nt8/v48
b7yX2MSIkHtoDDRbyP6MPh0AIXaXGjJiUSBhXjMxpA5+Vpy8dzoKnXPZlXUtycb7Ok/evoym1Zzk
VDYVxaLsEDItjiHx5wkG2WJRgSHggGZGBkiBcaPrk3uncw47VxAynCEj3N0jegBVRPKMISuV4R9Q
h1DNELjueTM9AQvicJxTFvcJV3Wltu/BoOnywm8axfzJIlyNXOh3nyroBUXU30zAlNR1eha2k3MB
7n2k3MPyqX2Lt8E31cw4CiJNHV7ougK4w+KjOs8Q3mseniBpUe9pTEvrwkB2olEUT2bpD9lgli1J
rWWM2PQ6Ghsk9gVQu9T11yhZNgXPUwmjRiinRSfct1queyDBIBWgmSwvgkGig8hYQf4Xl9EmVR4a
U4TqZI3V6mujo5586iBsFNJAXppXOocUqI3GN+Yj4IOjsD/6sZtshXlDYGl51bZ4bekLitbCdMzv
31/PeCi8IijGfKPvrFiX0f1eLQIyHHP2indw6MevxHoSKaE04DO4ZD8qm8pvDWpnQFOv1Wb0YPRX
8QFxmLJG8ivhGEhButcYZsjHeld+IExAtHo1qnbMOw1+xwBT3iyuWxNnaaWpwJej6wv3UperePux
VgA//5e+SnWZZPz50Q5BidBMopOQ6+ReemqSgUOrQP4MNMKA/NLQ2gto/YT4kQNltQc6DbiMXK2m
zInpvD6lSknV3iTqvFArh83jM2UbIuomxZ8n8dCsS4IBcIsnfbI0iuTd2lp5oXeTMBk5dTXz2ZBj
ly2jYUzfP3D8ooY2Wf4TJBgCCEGHA76a1ViOp8dlnUcNa+n0jdRPmpWBNRxC4++0UjohNkEsJjJh
tzKHhYKT0j+XmszKyiC5oC02gU5MgD6+wEPqtVJ5aNpNteUKfLZKkECAAGXKWCypJovICsheKv1P
uTizehlTopMdcK6NPeXCYC1Ki9+6WDyR3ZjDx95VPHTJ3wvEHVULY9GJLh0k3obncXVFnNiI9pfP
ktBp2dlBoINVKBzu9Zef0F+vV9Nc/iQE/WHNiVAf9B98naeb23Ak60NqOJekSJb0xQS2GEXfVGey
cUQgII9HznHdInJKZcL+ylPfRHAHWwzNge4pZuTzn1pLAIQL0HyDyMJ5JlHkbuUK3pVnKQ2GwXxv
S5WdB+NmMxtrqsZs96ub96yrMB2YEG8ooUs65Q2TlOG0osVUvTvW0zvrq6deOPz1sK6HVCWsqcVA
hIpD6XAyiH1dmttErqRTofPawESp8K4vmEiYNbOGUNYJJlSM1EujMcuW7DrM0SS9KgnSKYwzKEwf
KV4Vk0SM12g3ll0d/bngx8GIJd8KWD4IOTo2tgbD4S75kCq/aZJXoYtew0e6OVwg/YA9lmmOUcEJ
/7AB7aM1fDrhq11jcm+ZPfMg+Uc9T9OBsFQEOttA09r+h8Lmw1FnyUiJ9vxBiBpm5Qj1hJ8t04fQ
mBIQsAKew0DE+17z1sqg36sZTkux4yq9dRZL1S5tH5hgAdln4g9jb7Ui0a2zQZJxVQmDh6bFYU7c
x/y9ApCfzxqunVMWRj76SMnR8ELWtRF5+fGXmwLwq05RPbYh/eE8tBX6xu5L1d2R2FcIfJdihZQP
aDf2/wiQHAcJOuwNqX3t2cIdOn+BYuVRB2aNhmFmPOzXxr95GwO9Lc2f/F4psqC59ek21dN7/CjS
gCaSj7bPeG+eJSp7m23fyl2RW69xgWwFTS3CvDmePM62ieNGvSbFtrHcJ7HJhpq66ADkChgdp26D
HZRPLuBYPZye46Fpl+AM4oWuQC/Sv4J9bGjj61f9M4R+jQXaH7WzZUJgm1epO8qiQ+/UvhjSX56L
a+ok55XktxLda74pajVJK2Zi8gx2d/LTFebIdjhbm0ALVIKyfJpbz1eTsu24RV6oWcl/VoLOiso3
4FDT1AFxH/HE5Dsr+vv77zmS0gDk0kEFpTe0U5PkHSp6kpTHZ0jtXZ/MZAYUckW4z8DWpnEQvn8/
tYv06Mi0393+EZUr2J0DpTNWXsembz6bThfEYxh6JlVrCyLZamGfh0PLZfrDX5l9si46J+Yqv90L
VhRgeSisoKPlyN+w7mwvsCobbPKXT7q7znsiUzYCwVk+v/GPsb/oHRdZF4wU16FccvIyooYUajB5
4Il51aONkYX0o3NcAUwNdBKuFUEfcsThg4ciPll9U0q7+7f1N54NDZoBdndafEGlmBAV4IGRTrf+
rgVpf46fZErDcZGOx/LXpbAs10kOdSSG+fHOajqS/JX86ux2uxOJ74n9ycYFuT3vqMTD80dyYEfo
dfXOAqyM9itacI6apqz0D9eeIms9b39pIZy5sB/kyPihwqtNMt9a0/jS+w5MyOcOO5nj/aBnMBV1
gzrjRRjt+7LQKEdxdRhwrEGzwrKB0iqMlAIAllhSq5544pzywSpziiP6cL7mRS7TO49HYQuya4u5
mBb01uSW+2zMDtaQAHYFLQeL8m5/GkJ6LPq6DvUcO4tkZOl6qo66Qzm7xXLH+vrpK77cfcMeb0J4
+ogyy13XrZeIWrhxJ3CgKFrLh8KtoBd2PTqMpiTHslEf34y4DaoNCdp/nw7FUhbcp7dLvsW23bWT
HD40KVFP240awxmDW9IUQeMnYhPgCXmSRQDQtFOGN6bfwhRd9erKfMl5/EkyNjGinjULOUW7QWpv
VIFplH2eBPhqwbYjqPkEhcAGfAWSwyYRdCsTjL5kUhIDxI3COX91/d0NKQ9bvh6UCWtpswH3uYCL
iCrSj2Bg9JtQ2DA4dlsTKRik0EYS11M3botQBH1B9p0cWB3lDOeCbPezjoKanZjG6ZPs+j19dJLU
mkInoMV5W1VhsXQnCZ1FydlMs6ugRUxXY/PEt+cp+FQALWdA4YiFBdG9CT0g1HKa7yVGbE3lRY7Z
8jv+7jCvN4UjnNs6FusQI8jnu0XCKeQm7/We6neWAwB3UFlI2NRJZVSMCJirbA4Fu9FrAk7S7xVR
APJftFhC6Ks/xaPxA2mHjSgx2HFMR8rN5SzI8A83a3io3xFOkbI1MTNw0l+45292icKSwRN24dE1
w/mVKpfHQwnFIT9ba2h2qT0Tuqq91KRxX9JmCR6osqhNw8H+W/PnWAsgCneVgJfDV//y9GmKGbFl
jBla+v+91NLCcBgc7/dEPRL3UmfVQ90T+CrDy7yvmHvldM34WaKwIe2+WJwwbQuTeIgOdrG1mjLb
Jh+gwrK7F1p6dtxcFIi+R1CRIIANKgInh0hxg7hHvPChkW5qjv5X4VUuHq7fcPA1VuNPiTwjpVgI
WLtHtLGoJQPPT9PGyKCORuZp9MrfKk68qLRaiYEmP4/pmGVC4QLkdpYRg25fzGbRHKyaknvX9eeq
Mp7HblDbc2eLzayoFsx498KcSE60QecQHJyKdGiBRo+rUGQBcfCFFv5s3T7EZeEWx0msH+HYz5cv
/D4BiR3h6N7K6hJazk+vEmtopB/OmRagFXGk4keibd1DfukNObkwhL+xLDwgpeCd+st13ndD7kA2
gS3VvNvFGIhSCfGNswaTpcmQz1/8LBKVVH3J67FlyB0CfblkQNWfi8Aihl9PwbWyWOrcIfqOI17Z
aQfiYAw3V8vA5Skf176cGwHoi5dzCIY44UJ/RtUad55S1eacm8EC0zIAJvDgeoDefiO3W8jb6Lxd
TCswhlYh+lssefKBNn654tmXQKYPxg7/Qu44PJ4tqCiP7p+29A7aY74fV+2M2/PMVpkMKRCa1CIV
5qbibufkySVoRi5eXzU8g3Pb+UvjSqT9MvBtfWQ2L/5yJ9feLBH8PwHqWmzKco36nIAeqdnU/DYw
3K6lg6OXMkidmoe4ligr4mC6GtbylJG9m++JbLEuHP1ZygCuU60rRU1YgthJMuYoycdefiYu2lwf
HRG329d6wmWp1czZ2qaegJhKpynYPWlR7n/6Jko9jBbwRLCiiW5y5ZQCBKTzxs7tAhKFCnp9HXLS
zTjf6xupGOygPqLVVZk4LTcYWSM2c1W/W6a+he3pI83TAmiJ9QjL14uNTQPLnS9oqw95VjM2nGIi
1D0b4XewBiARWqpNJXEnDJwtfNXMSYjiu2Ci8bs8VxAIIiLAu5/Qdn5g2iMZchRygKeUvcLTyc5+
aJs6Xg+Y8/hGomNFEXCy5Kh+1VzWQd11Ra8EoSuqplUE8Ee62vfBJR3bjvrz64GFD0O3S9y9JVEg
0QjREY9b9zxKK36QuT7PYOriveir+uk3466p4y/wSdqoGqVENcKEWVv/oXWGua5W+cx0KjCDAJF3
Oea+SCH0GJDCxzzKsTiRDj5gJMRZVJIItF3n0i/2ZDoFj1VVgkC/Soxg8s3eSggjxmZorLaHE3cK
1sx2mphvhELWxgb+pW3ZYYZ0KMcDITit0+BWkbhQecjDoou3qN94vrYB+Bp2hJokxaSdpPACgfoE
UjX8u0LsLumU4Aq6v83vt2EO4zp9IU55/SO5r+wDqLZTvz14cZcAo4QnKQVL/mNg1Zwk/ebuevUM
lkCL8eTRyVFtTXheSpALuc+D3WtCp9Jf4Q+HDp/UAyozOMWh+W3JDy5NW7f8MIqqCDXiGjSr3ehl
RSqJzar2imAk1p0tkw33uiu0IMeLoxXjULbMvy2On8DfoxvvqPsFXTJ0D8YJqq3/a64fanjTnK9h
gGEWQVGyX2jL4RHmITz+yBlDnssL2O4IxdiE979l7I6iujFb61w6/saFjcYBgUxboLGGWs6j909e
vDlh2qKxIo/b2tbfVTym3EELzr5+NSOMVg4jyOu8XMOi4aTfakJ677cb5HlMr1MSvNcqWqKsS/cv
QO1tFCzvKIyM44eut5TNvE+MD3hYp3Rehn8UeYpyNHaPo0W8MWlEYM5NiLi6y30n1N3q/1u1QNHH
3BQPay7jPOM8q/Q34rkM1oNlsGkV0YIJQpDd5orxlvdw5Rp4/DS1oaNDa0m8EyeRqMWdMF/d2tu9
Q1dpsCZIU7AiCydtNbZaoLI9uU5PXir7iIh9HXIqUNbKgcenBIy3u0ewBd57m9MZCeXsUVIgXMI8
s7Ka5+Eb0oXAZcZV8c4eIW1Xj/+tAQDMWFFt6zlYrtIejeWcSOaY3BR+zBrgt1ee760sKGxWT0bt
O67YeJf7CfSdGB8REnT7fgLFPvJB5BCXRwx/Tied0wLXAZeaIcOr2fW7npLrqg543Ki9si6MuKpQ
cyk67uL+UrhlkGfhuWmCfgCjsqmfvKbiGGGOIGIgPo+BAwcnibe+B1RHVln8/xmDvxlKYW89IIBD
vEK94Exe7i9zcBuIVk1gElXkztSzolZrsG1d4ds2m8reSYNhzu+GkKRvMO79GCoA24ncGS4hx74r
u7GsI1Uk/Iy+F+Cwsby8lc58rj7kOwsV3W/4g9Xb+5+L50e98IECxO793rMZiS/OLSe3a8YAt5Gs
BfN3yS2r9wHQXn/BplkJwxY2baNQRc7zHovW0QGSyPDKb3I9j7jPHzw45l9uB+RapFffGX4CGDHq
6FbtcHIU1hwFuuhoE0FgKEco9VXdUrCqp8yQUKE7kncGkay2MhHxiJJxGxA+6+6RgBkTyzCUJ8lk
0QO3H5eKwdCBxQre1n9p8Rk/2EkGCJwNPKCTUOBWAXyDXk1ou0H92bfuyQ3rwRcrXPtX5Sy6NzrY
/FbvWW4NGTlmpuXzm6Es4xQtVKLwiSl8bumSq/OPtF/cawuVFYeitM6h8Hh+P1VzbGeVtOryM/Jf
H1f97kXNApg6ZVR0IcMHGfatf348JDNxchpIa2iG98402F5Fuv3bVjMSuyLRMBL93NBBv0yOeQo3
hpcu48DjitKiSy6uL/+oH82c6iv5EChU3gzUjZ7jCDuS7I3zGxPrk+fic1VBBAfa1ghScELALQ6x
fhfyTEGkiKYVZJmumMUdaPkpIquPoPNRJwDL2WsKIHmMf0oX9dslDVaxvI/fpT7YjQALW9LSttrO
bgvIlHyns06NtWWP4u0W+cbMWGzI12BsmNcrMNdU+0BBtAZUBvXQv0eRYQAIV1HRql9vCXfNppzf
FaSOCG0yF7CuO/hxDpFsUMsqlkHINsmWcwfsxJdlR4uMTjBh895/xheHwz5sJdYLPmXKhBDsMxah
J7tKvLTvrRlfvSmdo8RA/6K3KjSvKvCvNgqdeRvprPfstKex74qAGZDaHCnCpCYyIA7Of1Hw+xvV
dkZ5jCzvgwjvGu+zBf1cBZL81lQQ+zOPCYp6TMQ+wHqfKNmVEVvKuWcxhgEdcyjMiRvalWT5Spa/
J0wmpLAszqf9OGjm2hXEjcdb5OKIVLYdrBNslFtepO8mcAq61ks19AvTF36AiJEnGh5ys4pup7+7
BxAmdz4anX9Ciqvju0a4YbKJOSsofywN+P0zZ3GtgsTEDEd2u9R6IqOyBakUyEd/I080jwZ2RABw
1vGkNCesBepp1cGxtafwFAwep5+x+Bwc2OhnHXGhm6pu/tLHlxca/0KrkOZ6ydQN365YVb4vA7NN
x4oqeBQ9BO8Bmx7iQpEaVgeJRJCYcVLA7f26qNOMig+kuTAZ1nfsslCzMysPc6mNdlO2ARvAKoAG
OQRx6C5O9JqfFbGFM+VyhIe9TGj6ryu/GcTV9xzTfayDn5JRu459xKp55swDnb28f5g0cIixQDdq
lWFbyYzKrzLNu/19ggPGezV0FA6S9jjguMNJ+tvv30qGm0kqd6nCfzgIuvFXJXQRf8XV/55+u3ui
WHPX3ZBAvH8kZwZmv/tqOUKQR4e9e6xWerk4182h3R2nU3roibXC72J10PAA6ttr//yw+fSOlvHj
r/82qtNk60MoLedwMIz0RFnQGVp3SHK6QwzWy74HQeSRn9X9NJuOm9leI1kXvWiFQlmo38KUNZBh
ZqCQiEDDWcd8ldJZN32j2rWH7ujrqSAeAicr/IJ8q7jOvAIAHJ6F4VRQbMc9yG1EAfQqecrLUluX
UlDupEkXMiEsHPfFfMchqtM4xQss/P1ULAjeuRfoze/3qB6v2kdW/WXO2pTtkr5jbbXrROCzv8XI
pfu9QUgcq+ESLzlYa2NblNg+gbny2/RvU6sSm0CbyGM/ZvEwWIFyTIF2YjQotI+xAJYOyiaKiInV
s8ioYX6faf5X90gZRv1l4axC9h6B0VXrYVy234SZ1diDmDN/cfnFED6a5D66W6h2W7my78c+KzC8
dcCIjw6xkVF98xP82wnxJyXhmXli/wwudk3CVew1zy6ijbAFAcd+l3fO4vpOaCTX/PQQ0U2Y9hFJ
UtMz7E5BDWVP2JAfAL+sWGP7SFFL+nZIZD5eP8CdEmyELXVTuFyrZ8NUGjGPe9X36H3mJcAe4A7u
6Cnz98Z0kS0PZzCfJ/3KHh4q2+oIr79KaHh0znFjclO76W/H1XpbQKD//vBw7j+MXV4rK6xX2S6Q
b49liq/5P1dDerO6Uxec7cSnWQk+S8CavB4pFOE7Fgepw8b41hSoho5dXxvYuk5ONch5PufvwxNQ
PEwgr+WDPomrcUPD5uxgna1g4Yj5zNaA+zQt45GdT6AN5i41MF/UP3/FDuhkCDOHlmwbDS0Rlt9p
aPgKvxVoOOumcSVuuAcqfN84OJfaMZuHYNzs8yiI+SkOfRizFYbO4sgGekSNXWxUIbd6KDGumT3i
mYRVl6bUtYcIictXwMx74c1UbuP8xsZv/gNwMJ9V5q3VzIkDQD+UzuNbqDNo/LT9pmJA9xc4ocaj
eNtNWMz4g1CHpsv3NJGOVl8IQAxpBJbysSF7UCrLcMYsDKqJQldqGgz2wMm28ewD6Xh6TFkj+62G
eMHFVioghKPDvUoW7qv72GCOU+3Vk97v3TLnj/V/RBlgv5L4sXffS1RTXGjMjfH3AndLhTL+rUhY
HX8eSLgROfkw4jJWALDJT1krrr654hLKvhZgJKfTWmJm+VJlPZniyz4lQmx/8CgC9IYgSefOfLdO
DOoag7Bwuruh0giU73P83pJr6vtlSCLL4jl5YkpGpKNo61rMd6SDDeJkbV4bGvlQlV/gIQnMVJFt
imbiaI8G24qNHNlK9fz8RXaO/Z0lMWT3OFDOtPp1OE4PUhG9/7YEbD5vfLV9QhAdu972izpdsCDl
N1zDy3XW4axPVh2x6EuhRyUsAUZ5ALZEmL6ET5W8v4sTFg4Onx8o9t7TFvoB4CDxxz4VNH0DeXaT
1jN5QOOxnSGPK6QxN6Iz3PF10/QpV8ONSJ0magX7IYkhQKFMb9rp/+Cp1SrhqHIqA6cOOsrcDdos
qVbMKzc9EqsbgR3jyaAT2irUK0zZwF3iAjgoguBbJWVzyI7BDkBo1Zo14ho/BrelQQqednPkxUNL
u5HE/Idzhke4ZxgrJQaXSZbLtjPt6pb+pbiqkMRcz+Efu0WQGrBKOHyMTa+/TmyusL1PSjDbP9fV
nGPHb2HkMErEwUQl4hmitJ2P5IuT7EPlf66R0fR0PIOsruyDy56Y8y1rQ+HJ/dQ1XtaUsUzXtxZk
bp25FzKaZPyyB/v/SRrcKyd8KIel68af1pgN/fOYbt2Aa577zCCz0rWIfrKPI6hCQpYAhr9LVCLN
PhO3tPqyN8oKNECzcZBF1bmzKj4dHPnlQ1dT7nEr5qcL1eiCtVKrsKE1VSm6RS+6gtejNEV+NAqJ
Bk4/hb3/JzOH/7bHGSS5c7NE5Uv/KdtzsP38AHLFalFMbwO+nGyS35qAkz0qP2qwZu3+XYAwk5uF
15J9d13PcRGbNYn0QprNJOt+08o374sWPcs85JD6pfbVphJWnHmJBxPXN3ImsVBdrRKWwxWjZWMY
duzlrJPtxs2iip0dcfrHCESj7rfZ2Q5UXAEu7IDWABCFd6JQrSo8bvdIFvwDhO2JlU3NmWVs1Jb4
487BqjuwnkUVf5Og1ZPnrXZZrrcZCGyjijHUzS1s23i9k2WItzO7yqHgF9KHSBFxkn+tDYYCLezL
GFe6XvLRRvXdnzkWmnKkmSv0yocoMf6Svz91BfMZibyow6eHhzmiLXdOKDYlVeN4FLMbg3tvUKhu
17kGO8Uu1WZwR+YIgYDYQMUHNL2AzahLdL8KEpsZfr2avShXoJdhAPU8zmemeoZwhWZWpzS4Ejhu
b1ezgM+zVFOXYt3Gpfkcq5nGrFVXudDBoc5SygKlp8HSwIjvyJbfdaU33eZ+aVgPm+bIoIh4VyJW
N1XMPSKCIg1/3vKMijFuxo0K/P7ulNVn80Mxwfmsh6IQWx2RbA6ndK1tuF3SmGn4FVts2XlO5ngt
7M4i/ViATiqrmdgFY67BR4vylwJIHNnGAJa9fjLQ79XAfX1TSAyGyZ2EFfuSLR/lKXLjmfsyjtf1
FJsLU4Rtrz7jLtobOLmD6uJq5DNy3WDuJHizDSU5c+joQjP54dcpCM+CKjDBsdKuw50R5SfBnP8e
WHTEN25XV6G0tGOgo6SJ6s0OeyFdPXRKUlJJOnPCgY78eLVa6US8cfDqnEsP3Dsg9ANGoC/AtF8L
c2dgy171e3o/cu547utYhT2l8womrU4nrOHHe4/afvzT9VlEbI7nsJe6X9zrD0veXyCk9nKcyOP2
PyRfuPk1FumU8ZgB3rMsfWoC1NYaZRmuQ27hLPD/tk7jqEseJLDFcD9jgzshpEVRumjFDh+ZXtA4
LCaK803tN9V5PDRsojZ86fuIvD5CRMgEV/Bk3sgFQy6PIY7tGZdpWDILDNMJShdmbotxXwaPpncX
Y6Gn1LOWbqnDxmUVjqUF1IIlE2o94/qeBwPNr2VQrFYqs3lsWblfNkT4Y3xFO5nhE+g/L15fCLF5
otZo2J43HKOcEbKcc2HtF22fL5ZJPYO5/ywK83ZqWVQg42Nk0qEwVAAsGCLCkWQ/nrCoYfnBsBMQ
doAIgwUy5inbnYMOB7G1FLEQWzxZFEMoWvRmXdEWODoUC4U9VZMyfk4EXynOdCDY+QAVNiKaCOVP
0OG8rDrh3j/2Fso3Hj3HLXju72jI5KMqPx20JJ+yGLjwyVrRFWnHh493mME4w0hXatCGP02yQF+L
CXvAYw9PMXwZRVoi68sNpLWU6cXVU9ts8NtWci+oXntpJasO8/KOgdXX6NFheX6QZNeLlv50ytV4
xc8bNA7WPdQJTMPxpwrPkWN9D6hIclVDu0rzQ5BaTqTgJgci3/WTz4B8/qCqv+2dledsbsRCJqLf
K/cM9ou8ARckecvqEjTuHHyi3sE69DA6cYdQcO8Mvw81W8uGscCVbPg77Ywxctl77q9mADOO9tK2
aN2mn54FF+8vWh52MVZkKNnnLd7HCaQIQ13Ztd16VU2BTD37KNWokLllPnThQPsFnoVdYrZ47yAl
iQ8QVlgDvUhMphQ2iaZE1rQ9IKiwH1vO+3CXiR8qH+cKc/ajGeHRYgZth6HPAmJl2TFs2nr7R9mx
UTdy48i3mweNT5P8bCLzNl+rfGjifDQIDKrUslT7hW96Mfr47xgsgd92tLra2SLO1hPAekDcxJyh
LftKga/GwjNIGlzZVbUpq3KS05mXs1xjgnNx+xtEY7/Kgd/4J+uo2i3XSOgyWKQGUFzhxOmecWLH
fP27cSWLylraYN7bnq6Eljs/miSoIlx6SS9hWcr0x9OUfHKcKhBYDV9bokCD1uwLqEYnTR/QXr7L
Yat+pa0zGZOjUhO/3BBpYyzK4Ov4FCqPFfKg4pb/nP37S6jYOipAgiZgGSkVixBxq42krXEsqZPe
sCy9Mv/xz4Xz7emBJWs9S0WfJICG+ccipelIyq1vExJUDvNb6VEzpcQWI8I8KrVF8SiczQlGhRjp
i6yZGfX2bxb2UzR1yoSZmOAi8wwlLP1xAPhivGpYGRpAb5Q0aOrUebDMAEEPKhcGttQ2q39MRPwD
TPV0f3jUaPwFndZtwMJA9UzY7fTfqUaKKYQI0esdH/eajplgXv8QgcUMs744JP1Tun+eUt/V2BhN
cARbDfNcbQblQqyEStVxzE64UkiD2YkNRIDeAagt/RZfMEXDhrMbzCD33RvceW7YYGc4ZPdIJ4fI
c8WJdBOfedZ2R1mRmMxLhGl8LmJip13geSd0TC851LdIBX8q3A56f1zItZBeZEEbtVpp2EK7dhfh
LzV5G+Ji/GrxIblfLu8CRhniHFdNo0TWEVn8bxYKkjN5n3b2p5HwO86thecwlHHTM15emusVQVOS
KwA88U8bl2hlHybuQ/EdH7hfuGNAKN2VXDSmmzoxPd3eaTGK+B/Ro5NMJaHoaCAI+QbGyNrF75zm
ILxYr7ZK5Vk9fvS8VKUkrGhRy3yqMAxT9lNhkjxXxPIaauwoyookTIYfrA2WJGcOC+XJWa9blRRD
3XJ/hhGbY/pRPIkmYvx612vgiol4uJqXQReo8tIOxoXyti2h11MAwIYlc4PvQaZ6giKhsReVKF0v
mf5aWoh95QTjPBGt5OqPFMcPv99D1L3YEy/ChIhY8euTgy8K7he5JzHU51+olE2keCNLqyu7KVjk
VkmdaPKcYS62+a00XuVut8efe6nO5nDIl0ihDNsVMAVHrATsP9hUy3ZpQN+GnMvEX4N3+WpkWvKx
PBfXJoqRxNp9PRnuku2UpHsZUsODqQKLbJxjjAxllIk2qFTFQw4sho0bm7oabWdp0c/mbKjgj8Fe
uqJqMpr88NKW5627gJtGrrCy3LTALyLPI1SwV0vJQht96UWlYpgC5lBnHETCzi4z8JlvTQWER8FU
uPiJKDP+23YTvMu/1cYgfde4LiRQEbhvjqIXv/9qTqe+nRVtOGwB36NYxMMT0EYgmvDO3XyYFsvz
Z4+69TVp1bBhT52gjArAdp9h3KWdqv4gi2bXa49XhqlYRfHjL5sdRqhdQA+rOthrA+TfM2Y9xJKJ
iThXksiEeEVOUyjr8QsxPYyvIHIUje9U/gqy1o6Zq/wNdchUSa7oOoNsN06d9URYVsoVSaDez34r
RnYYLRuVSSdUuOswULZynRrTzJz+u4jmbWCZsxh6N1z+SX1a0/Pd+pMxGnvsvujZV9tQUr+WksZR
lX7PboTCniUvAH9SzPTDtuwWAQLhXernu7w/rPjS4e5OhVIXHuysUsjuo7OGHW13AbDQ3S8yHBeU
tuxnbULyIyYO6JOARFT6To0JWyBY5KjURvE5KdxooZOdxFneeCRx74HpfOx6DG5ibfs68y1YpI+Z
IrvAiJvnl0L2whIsTEL58k4fUBZgX8lNNKiZXRnw9NLPcUmUfTVX/XJqFk69d94RwN7qIAsd0UlX
genxhhdf7ekI0Bm4ayqHqPpx0H6aBI6VC+4MOoB7AAkETJhjxLmhrIjJYRKYsYm8Ss5xdxbo5WDg
Np6QuWOtJdutZnfj+klUrIFUsPXc69wYvCAmpsDlMlUYMulvh1nlpl+sqo3E/XNIgSc05VykhBG1
TBPwwMKKfUy6jjqeAO7MTFuFutMrVTTdHRKtlpEJqCODmLCI6OHGcKwViRu1qRPXQtdhQCq4447z
TIPa7ZVlZV6xuHqRxch3WGf6p3FWgkD9CcNrz+WbnhUZuxdaeOWqLpnB6MHqrXYEOSDyK8V1BS8H
3U3T3Po87R0H2GZyDNFg30UhAgw4NMUGskRnuoE97QlKr2B3agnc+gGHTWd0FsoSuI3SJ0f66c31
W/2DoS+h1g9uZ+qDuhIJ8RB0HQPUK+bZECSb/xMAKcbSOVN+m6RkU9D5UYii5z04wdcK+AMRzDi8
CATy6+kYjmrt3cAJxHpuvgHRcaJy+qNrXcjf4HNj04K4Vx887stJ4mXEkG9b/vgb3W2I9Sp3IlFA
AC0H2O7DMH1s+ds5tWeN2wmuq2uLo6KSkK5xzMhvTHmMOi2+qMY0Wg4DWjxxR1TgiMLUfBEAssM2
kZItVQHCPh7AU8SmhvnHd/JFMtrLiIAFrKq1w9Xi0o6glDgESZ2ChjviMBk72/zGB3Ok0w9/yXzF
RERpwCygdLbS4UmQKyBrECj4saC1Ugncw+NRzSPXqLThyFJ9yTZ+liGp97u8waBp5UjoUn3mNqMF
yCiqF6CAYkr2VGua8Pr92muSF369isuB8fmYIIPuYNQAff2niT0tV61MThSLQY018qJR+dreSKl5
I1TO/r0dqExc896ZS2kmSKfoeMbrGIIMhen97jDsB9cEptuye2umoLmhL8DxoRsoWeB0x9MDvtxJ
AnKCMVUdJLqUHG0dlqFKW5udxDqCRA2WsSg6vstzlGLiu/TVDCVafutXSZOrMv2mL7kkdx1vuGKW
uZzZ1wqlcIF32Sdm9BiT8MVS0NyVPQTNFzxSMN8ZySRaNN8Tn3e8Xa08D0YmHP5ePLyiTt8qqBu4
Av4W8XRjgoQGpyhcTDlOU7pOJ28ZPzz6oca1S24G2x/nYwdGN5gEaUQZsGMAW1UQpHRRDr/l+EKm
iRKJrSLEPQJo6OVEMqZm1ZZu9f+j2uOGICtPWOGctJ0vQfxOuTEGhxXhJ575q/yKv9ioP98w0+O+
UgV8jbKp4Dfm1UARxo8UWrFywJguFXa4oR0PD9uc9mg52S9VGGtjbnkR0R1GmcbKnFlT75nZvM+K
x16Xrot18X5V3+exIk6Ddx6U7Zufpb/+Vue6mJX925btaCgBSUYCWvNUt6hIJDOYkMpOCVdn3ZRo
gP9paEWrX/BMtDsY2GJojAnKI1Pd9XiS3oTx5yiUkdkSpxu/34mgMjhgmGPZmNwgfkIIjy+ucDbA
gCfoDe5k3eS0/wOcdZcgqO7LPj00J1hvE3iuHDfB3hEa7t8mf4FYelgnyLYHflZRMy5PBEOxwKoR
k3iPvUrzuDHnG01DlOMqEjIG5OFTQE1Z2rudw0N+VIigwjm1imFyux68H8piCHYc5w8nfIGyVGXT
mFXUIqB08xw8fSzQ/N+HWdpv2pyBOIduuoajcveNvSZytDa5WrlpQQrKKgyOosC0U9Nx4yZrEs8A
ExMUaFObFxgEN9z427flh24JIt8V32Izoj2xhzXP+/hwHs+CgQC6yTgn5vIz3dmxQjQcwN5DWO6+
n4vjPpp7kA/iEnAlgU79UkgAFBSi9tME4xucdTvT2HtTp3mbsAgZvYHtzpyRMoBKBzGQrJsc4juk
SsPcar4OofBQbFa0LzVp+7GuNzXNxTxwCZxZNK1zlIxRMpKDwoZWS3SJmnDR/tLBLtv748cHWioN
pyrYiIjLAVt53GVqmN+c1D3PIlepUkMJiqA+NHtgzsUHrbDQJC1q1lzhgrNyNl/JG7/4BLXpbg7w
30CazP2LaSBIIySPwITwUyYmIK69TSLnOcoZdyZJIXSqJkSjINM+7P4XO3SUney6+s5qjpZyYqPE
q3E0r6+etw/Nxf7TSW1deHgBc5cwp/Vl2C/tNKkG+1Z/+MsrKrlyGLwkd2VkKOB/OJPSqWrpsstQ
UTJq9CcPemiEPw5yoHG5lTuG1XWP0KSGMqtcSDzzzKpPPG2SNunJsDUembAf+pYj6yjW4kvtMOgY
/YbGInFRsBVTD7mNCy+UNxtgy/HmMpfXmCYKJUfV+F+WULz8Bz9/hB4cujubDMcLKgHB9nPFmpkG
K6dDUhEFUDNbaF6/KhGaOGKJqsUj/104/VcTo6ASXoahRCRLdgcogNGz4D7iqDF7B8vBePdDuNuN
EuOGp/wpZ54LxEYSomltD30Fcny8vbnCxJqioLIZzZfNDJK9iFQeOfm4Z3fzU4KkHgU+4AY8U1G7
H+cDBDvxOzgiO3uBFaOd6pRlzXK1DTj4KjIBzdQV5lqOH/FCR9db5CVtpRnWuTxWNYj5Yxpv1U4G
j6rDsRURayNYcWpPcScUx+eHLZQthIHFoDTRp5YhVMCe6J8kGh+3OTPP8pTmukJqideCeKI7kd6I
RtkPqklXfCd/NO58HLJ5Kg5BIqqEZhc4ghk9ccj4okbjykVKFTeaLGTnDivHDGfkgMy9Oml2nNuv
pHXhb+c9fzre71gk2Z8CION9Yxv83iQkkEuQ+hWPeXpnXLpL4+OsN0oFvPxJ4QG4EMOFb868KJHE
MTgD7C7A2jF1fWoH3hXz/asbpJHoWbFVTPf1bQv/2C44MVFPoKCfAAkcnE/22ZUd43CnGPrTD346
zuYnv8RNks2zIe9xNjH0mH4WINvSyRrnB+ME0gvFd9vvMiG8sJHWKxrdkrX+iM4w4Kpsgilh5iE1
APNP1SpJNRaRXqxqDIepHj+INl8LxpEnkUBLTWgivyIJNBkD/qm7dXoCBd9uRun9IMMLzMcZZsEo
1HV7aYwm75vboMa6pNKNNBTsgUSVtSFip04t75zVNoLwrp7pnlHvahG/2cu+yuI26oVflJ7yYdyV
b/OehWuyeAJEwYHGfQwntK8UNcgFPgyU/UdLi6TW5NDhLMYVRTFr8qbxbwaqhOiPIij1elE2tNEa
Sspu/iOiyZKwqnsSUYf2IyH44gtORfVwUI+FbznsuP/r/vuQcJf45KNeHpDGM77DzYDJeb9j5uTE
wZQ2GFIBuU2djdKZhB14OaBk/fAUjNi0YDg2mN4vAikD6igKs+SnMW2MvTEDQ/udAFI1T8c9ABsf
rAnsSIRq///1GxD5SuvzKdbW+ghE/kA2xh3DAaQy6YNMOM//eExZK9YZwCOFIrzrG4vOBH088Oab
C/AzJC6mOYAY0s3HXgSyIx6J68w0WUxxTCIvkvYoNEBcWj1IKXczSo68jBYCzV7ev1akpnApqSxd
OxPSWJuALImzDbDANEnTEaLXUWuOdrARhjV2U2YGcTcpRN2FHWqMWBydU5KDe6HF/p2Secs/lRDh
vfSlBdefgLpjm+mML2ZPUG2dYzhU1TcqbDGyLHMMmPD/uoMcAWDXWJmmqNeev2sz2pPteE1grPVg
GKyuIT8XBgsO1F6lBYyOPyJsjxibNHkrXqoXuY1i3OaogswpdQn3PIGNp4Nv9TOLfumGJyFiuYEZ
YQI9amefX5JaYPpSSa5qjGo8oV5k8Gem8lR/CBpdBW70YWjyu7fxvK9zxmFNB4qkpZf6AyQWSfAM
cCh2D535W3Nod6CGSjF8wHXeZ+1uqkql7oL6ogxOwsOu30KEi/Z0gzXTuWSehCPTj4mIEJbDuoN3
8VR7cKg8yzOOUyUzEiUaw8qlKKjkCi6Yzn1mZE4fTYlv6/00R7kbGnBUJIfcr2YY/upqXpHdVST3
ByGDdn8qRrheD6PLA6NRjMFVm8v3k2vPg1nv35S54ZwwkjCxkg7FSkXu3g2gf16meMoJKIOVlkLk
7LlvDqNVPxsoy18d7FEI0kMqay+n1glIM65ju1ctjQHmKZBL3a/Z4jUqgeU6WtSn6beJ1WLOycgf
+p1Fhn8jib6ZXat4sjrkktLp94L/u78tCkPJ18k5xWJsfKaZfMOlhTW0ZP6JS2lpyaBcZTiWyTin
ct7MRMS2HXIBsO00lodIzGxF2XstSsFG+yqT2Aa9m2zATuGd2+mvRqYIuVOXoXcQIpKQp8/+Q/Es
lW5SvW5jfzwrd4EG/g1rJicinIbfGTv0qTL7HkUHZ/MPQTa9YI+lLuSkKctEtZpM5BKzN/BrrIQB
qJ+8eN4NmUtvhie6vbh/mx3O7dguAKAh/3Crsgyd84WDJBZoNLYc3tiQEpp+NvIL0tjF8NXNmXIQ
q3UE8qlRDELC2SJUtwk2mqz6cyxHFUWbCelgSlcf/KbmDGhy5V7dEjl4eOMNXfk91i4cTWZMVwN4
mQdjaA5rejtaw30WLhfprXwyl+s6Ao3HUIGN/3dnUzgZfbLbcZaJB/x53dvh2FAtLE5a6qRaUUEy
gB8FWFYAutT6Er51jNrJyVxuzic4MyJiP7dGja9Y0lPuo7/UF+FNxGPUB836KKMVPmaxntNM6GWS
CGXcA0ZyeRCl0fSJWsbldqN6a+qvXf0OZI2NoImPCU0xDOj4Ip56AkdF3tokGJWPbxv3m4+TqTit
lKJ2lGjWIEVMzFgKGRhsx0//JqkPSe/t3EBJzeYht6XrzvtBmsFaXMoeGLBLRY4rhAaRztOKwxbd
AfwKRTuT9tNgVS5Nsly2Yv4VNZ+AoQhMKWl7bvch7bO/y92H/hNPSM1WEZjDIi3SX3ZvAme6RYpu
TvCUM3xmROyaSFpM9b9/1PYuisiDffO7lT9ZwqEl7XRbRdyzL9SXdEhr2F+uKvk8fA5UxOelhkJN
tYfezjHSlCBhQfrsuHsIO5gItFP5f6EagetdK/Ul61WTUyLd4Ij80AcEUG76lRuG406o/7szQL0P
wvcMaM8YZPKjerBV/ihJ5+T7O2WMe4u/d/B1lIxzYVEj/SM5vkg8sB4s8tC7XWTiowybIU7s5Cts
laxu5aBqwAPJOzB2r1m9D/taBaQ7lzfhQGN1m5svDKP2vtk7l2vu77gaSz7lXUi4LQ0yQdD/de3c
VfwbArHXwM+5SDjO7taisO5ma7kWV920da27DpWGIko7XvUdU0oMkAwG1gUp+jziXKELEiwCnMW7
xXa4tadDe40X3CP9CUjwJU4cpDo/FsYi7J1ypmbiCM803zqJhJLK1jlZ7mI5przpX/4umXJq6Apx
B8C/s58HvvTC36BUtuE3gnVdi9h2c5HYskvtRtybYXgEjlbHiEm6qOwRQhq/uP9+rPhXPocxCiRI
kkTFjg0HT3odR3osz2vvQru2uV2eP3vLnr/c4zTL+ATlv3Rh19dM4rMG/ZdBNZOXxzxXAeR8rr9x
u4ElxPkTa3JVMqvkv/c9XSuhzmb2IDrvlJ7lnQef9k+W95kKeCvRJwEleTSDwvrdOY6PcsfYcrIL
MONi2s+eiDnsKXtMtbXJgyl3wlSjgbUck+4c4iwaOZq7C2E7eUXeQfwHoy8tgxs2ZKmVf6oT5Jgg
dxSNwEeCedY9yGognZ05S/gRPpQndoLtpFdp8rhOUvWvK8sKN5iW6a1YQQdxIsBwS2ZR0e3HpS8t
zuYgSIKhPJAeGJH8QtA9rTvI1jAGVW+EIs20NoSEi7E4CWj9tOLg9rXVrD3y5uUTHjtFaGx3Gr9r
oXFiuF63uG9ZB4B4DSBWrhm0woINa3/sCA4/Sh1AR7GnL/Si4M0di0sEClhp5BqT3LzwV4zut0bR
1iSm22OjLRD/jgaHDo4s8W4pZlUcvzsPZseAafTM+l9tjA7on3uxoNeJxE9+SN4xKEd/MDx1cO3y
SBL/iQAlriQITQ99f9mMHaow/Tc7hHjXDgmBuzoBWoweuqixipzUaCs0X7pl3/SjQGOGRNnK9qxG
4wQkR3nhqj9Sv2YNjOxdTDlmn1+g2bEBtd52qYpPiKBoNONUMY8pofa0ghxZedaTU1f5mOH45R59
SKvzmZa7fo6tzMH22L70+g1tgew/B5tEVjTANL4I/+JE/MZHdt0HLfBygwi2C4nW9dnArg5XasSC
tMgwmOFmKu4RcTdu8pjbcnqHSYipNqmi6kI0IiGzUrz/B2LQwrpfJ1tkkAskYeOrGvOYHmpUIEEs
cakc4rV3kzyprHtiHivN8UUgpqHgEvj1z20G7pQD+8lxLDD85Hbte0RUuCHly9qemoPYds8RA/Sc
Ll4ftIxurVNm/gXlhsY5eXOLaTdeiBFimz4QFxDaEqzh7mz3/ogUcxkWJ7L/GrE5BwxtFL/3dtmZ
eMGDqBkNS5STHF/E+pPeNvKP2WcEKlci6gLMykTgisEs113LNmvCBm2Zo69nUFtIoKYWO0GkWLPc
ABtVC8dSzWcKhTWnQ2ZX2+SSiiuP+yJpAhYt7BiXRNsDkMN425qtPCh7+2Ezi/O4638N6qTn7YvO
I4OmpwlS/evx157QRN9YcZmQtHOHL5yCNesy+s7veAoPWCC+sM9LnJm3sn7Q5Ai2Uof/gvO3pANP
JBXKuCBAOa03M0YMNjycXPc1kQpkKCWPxW6F9HSb1/UiE/gIYuygrK4FkgMln6p5MFRlr6MvP6+/
FaLZqYeNC5dBK0Ve4B88ZHod4iOwjX7Z/i66cml8r51D0wEhpIzHqNqTh4dG4LOu5oKV545dXpwJ
QHg3z01U9ChFeAzcNFXigzm0kusO1aZlL+RdoPy0K/6zXD+28oUVwrS4U6umWdl7MR2SwXmafshJ
XJ/KSgFQxM4lGHWoohbnraX5xLpebGZbD6PNGq/6tQ192bUEQWGpVpYK5i09iMorXhjoVg826vM6
IKpEtANO8v4sIV6ElQLBqJBXSu7mpxJW+0kRf6jcYfzPhi/4Qf1RWUW0EUC6dZcu0OkmUs/NhDjB
4VpWiSRXdB6IhcGUDIPPB3Rr7M/2zA5W5KNMZqp0AriAAHcGSSmVmWV6DSnj6w5paFDOURICS/kx
n1fu/ZkOSG72r7FwThpv5TVM/t9A6bymw22dLfItNAadU4nnm1qEfEmRyRkvBrW77Gq1QOB9gugj
iF4W02IsCsyEBHDzbMpUthS7TM7g5+uFpznwIJzoPy2MrgOlGp5nTx6AQ6e7YBozO7SP95eQbKZr
jAw77uBbN/P05u1axu4qFxsTuW9ssOKtGYSUGBwJ0BPPJpcM4GYJj5ok+5UfxyPHv/OmydXgDaKe
Sa9tlX2uWznSXVn3+qQ8ZPBEnjZyZ2aZtqGWTp3KEmUDZei9O1RJeeemgrzMp4QYrRe00Bh7pJ8m
Bxq/kimmZaUIzTARy0rNzX5GwDzCs9+j0iamIrQjleEIi4oJcO0Cp/2fOht6qthWQasm8rB3slGX
XzMJ/0GxIa4Ev5jNAuQtwLlRkpnpph4bygNLPVtUb6FAv76IV9fFcb8teZGeDgtmSFnLxsDhigaZ
C29P6SDWtxG6cUoBsNQvB72dex2dU4HiimP/qhVkEohJqymlfXcIk8Mg/gfZ3NbDtzmHk4nwAnH7
MZiCLSbUD2qz8KLVknh9Zn++rtIhesmSk0D0Wdh05mEfx7v6saFD8etRmcLSMaDQVesoqIiSUDAj
jJENKHPNT73ReMBYynvxVr9VNc6KaXGM5I+Ivk9DykgFkscCQAwcRNBU3MsbAZJi4AofzIJWLPzN
pkj6wcNzQUoRV6nN97vew92FJtizwOqpqCnwDL2V4PIc+PdEeoawHPEjGWRobcf6i43MwRyFoT2W
xuJlBZ01kHF9w8izLEVWtHmqJCyF1D2g1gFX75IQhaA3NsUHgerBheTuanDN9i4QzYx01dDns+08
NrIDiQsy4ob9spgiGOFbOrUUBnPFC1W/Fjphis6xCUPzLziXsAgGipsSzqJQ4HAN+Ewtvfxo1yqq
wVrXbL3hzguoJOkXIkYqoPLuHk98rSAmzSZqChYQ2djqF2lsyZO/ONJFfWWv99MjJ0v4v/ZSXz/C
yaw6Uly4lpYnUIZ7mpl4PkRU/LGb8/AKaigulwjMQS1iZ6XY2rWq2pAgc01opnDXYDMperkh4T0V
w+rycC7UnTfqwdFuJeUmWwiFJENc+0s/mOFpnGrXEwMj8W6ZIZBofJwJUOEOFv8EcgC2F33GVu2F
chqSE3/fVuM227mEXyjpMwVPmvb9ofYeTVBt7kGJWm54ysizSPBTc70hSqer+U3Sb5UqOsU90nWh
oWQrOZPwMGqpdHeu+kLbwLYfAWsfmwNnYxPXc529ld8/mMXa8ndXsIHG+wDiNfnhbc34Yp23ycmd
99S0c4+LVRkI9e1vEpuUrkg0Hl3S1WT8sNJsLUh2RzQYylpekCsFWY639Uyy9FLZC+MdbhFm/dWd
rg8GcbpZY+6Ykxonz1g8iG9jGksgIMI1PqpQ4jDw0NInjAO0/gkt7+PAi5uQj2gax2BoGwpFP4op
GG1V9oJlthNwtcO03gcHyWCdDaZO3irFTjsKeJAzM4bk1UkM3e8wXSij3hi598nX9lxnrZTRubET
MxWT56szQbnH9QLFoBvLwBnldw++SxU13oKIu3cvdl8Trnk16tZFmJm/PsJeTrDWrql7FUweIhCj
5WEKLsDNa5PlIMfXPy0TvcR3y2l4YQU5qm/qsgp9yns4CoKjgadoBtf8vsQkFGjOP2Lm1LujFe++
USUVoyPxhlFZwgVQV2r0LkgoYAzHhSlEIkL6NJ7ID5p3+iK712VsZ1G3tV9tJfDrDa8dtomdOERV
TknEoHLJ2FlIQf22YWDapDETdIZs9siddug6eXGveCwL2QGM719VqdpUebt6KV6lyg4sKScIcW3H
ghoTZevKaj5C45bSxgtbUOZJ6WEridY5sCyUXnQvIbmaeODueKusthAp9g88Pn4ioaO/dNUUy2T1
6yakPg4lgRQuQTsTJdFakJQkn6TGYOKLY91/K2twuQw9T+MV+2HG+W+kj62QnwxlL0T0TiysEgHc
LsH1T4attI2aoUK0tKd4aEWgJiBZIjtMYrxC3WeREhemBTdmRAOU3pO7Q/b4tBGUNJIBOkOEm4dZ
o2xquYNZIODBfzQ3vesFeIoik86SToEHRaBPt3NSqf33wgjmirEc++Xrp339Iab9Ni5zqMn3UgtT
X/3VuxxQb6pCc5sO9AbtpuBoJQwf2GVRXbDkfaokjqxXibCI8pGj6SPpI+FvLmwbXXKACdC4/3/7
haqy2x9//kjXwxhmfn35SgMbB6XtthsbiMg7Zfk+2ewPgvthd3yrhWGyZicucgq/huKdIBhVEA0O
euE4F4wRrS1Y0aCf/mQ5Sn1/RPxRdrirpeiPUdeLEkZSGG8hFiRBNMpfE18ZatJBWVJjtyhd6p3K
lAClFrR7FzdDSum8kAUDMjuvrCrbZwJfSWjv1VqHZor/XAkWD4MZcxvqtGD+i7oaFHGbPsSVXZ7P
ykRDo+hARRBAr8ydWt3g6UFVDcWy1ZvnWWa+JYzxm8QGkUQE8t/x3+1LfVg80D9ljthSK6ouz1xf
jA0t7jrODl92HVsEK9kVR4r3WFkNTn4drph1UN/K75BSAzCtdR+1UOt7BzWl6ycpBys+1P3KGST7
y0MIqDK+uEoUr2PUIuqhTvl6+atAjd0Fpjs01nUkLtCXp8D2ueDT+M8mfjm0gt+9x+OO1C/uCvI7
sOtwswrV0bBUiTqXj3ZN286BOWV9Glnf06qHjzAJHauTjYEjnfjzow1VTXmQl5CTpzP0M44YyUxl
F9ND60L30oQNvlfb5iyoduZrwaEkzr0bVt3r+LNgVyJItWqgPoFYnPp95HzqnnIiksh3+oC+oPfn
php0KylVM+KcZfC2oOj1dGw41W/4tCK3r7mzO2/j1qq19y2y4kGAVhzbAozYmhk/Q184k5YyRQ4m
WMUlm267z9iY72hnENQ3xTf9YBB7wDTeWud/mHN2dswSUx/Fiu6VXnzhevdIIbcjBVi2K3y660q1
r6KFo4T5gNJIIDy6MvJfUhoN6w8YNRbOkJXFZuA7kDHAcmFgkJp7g9Ze7U+KbmpPh9un44qbex91
7eZwjT6ClXMYLWKRa2Qyqj6HI6UcV/6uG6TVRAEJq28Z9qYtosNiOVj1utkaX9MAVfhw7sHKvDb4
mdIMt6PyyJ+hhjTs5Vl4jXQZv5BeqHRb0BtmK8HWI2QRWuFXBF8x8HwBD5oYLhG2w6XojC2LWVCs
HYaALA4kDa48Q+hppAZfXesgSmfXcv3R2zXlyt119NMyBLlVsw+karU9ucuwzCBYUobO5u9mq1bk
C7mGzw+9wVp1E7K/DESTWW3jEzdrF+DJE2qme7N4XMxGDAKzFZz2qSFnf6OTJGc7rvuTYRXJ3428
PMjJ8ut1SvFz4Irw4BcVkIxgz/iuxoMootP/m68Yy6Rj4MUxHk+UkQdLNgzkH+RkWlV8LXaEVRW8
liHU8SwzlPxpapknr/6xii8qvSsc12VgvmntGVly0l9Bu7JCxebvF/67z9c9dGhvBsTprIKnovl8
NWgoVYuc7btDpMA3lYEFHT7T4OmxnXef1H9cQ1FceHkS7naLSOwjrZrSgNY5NHyLghivZ87FJrob
TknUdBZr2Chj71aPRozvcQrrLAp+/tg9Nvw0iNRTBMR6ewPg7x6xaxgmF07g25ObqyWUBBD5ZZqZ
OGsXDJXogR/qH4QEYqYjfST920hlC1VK7boNg97EB8/luDWzahdKgnvCIcb9dhXoFhB73iNkvkCM
niAs/PtbJIhvU77o8Tvn2Uz+F1isSRklt2ERzAsQhgwyTyb/Qc/8um5aDvmY8Izzrz2Z2XABeiEe
cg1iMD5JXP3HKVyu8oEIT19W/aB3oJcUoZcFFG2TbS4VOStOY9NjE3v2DQUAewAwpcPlRPWgLtXM
HQIv3HxL1A6JVLOtcbUVdz4cKSKFVw/lOXH8c7jhgUs64TSAR0pjxt+lL0QI9x9P7rsfM9GejZVW
6JMkni1Dh8L/mnjNowaRgsEc9BLaxmkK6kUZFo2MPBaoBkal8NugqfFRRMEBaNTK/AoHhXq55qi3
j4nIWwsV2v7GosyeV184cIbynyT0BeTLWIzH9ZEOf6PDpneWvg8SlptUZs0DG1tF+H4+hqs9CZs4
Oo1Ju3/AKQiDzu+xF12CAB8cTTKf6aAQ3ZlY2dTtCjoQrq4Kz/BbsJUwzfiQ1h9nihXiJE1sF6b2
sdaF9jAbhG/Y+267mcnA3twybRa4iSu29fu+s8ZE2L6w8hoZWPR+cGamLiV39SvkZE+Y5vVarLQ/
qCjlWAGyAYt5+IpEuschdzWj6iBOZxES8l4l8QNRfC3mTnijjj8NSXQeE00W862QXRJR+bMYnpC4
cmPHaV7lJ6rUzwpv7eLHQ2PIjdMyHaHpkcOKJfmhVgKGLQArAXF//MFOaXM9BOHYms6+VBTkGAkU
bC071fXNk9LdxdkE+WTefDAUwoUDLTakHIZ2PRkoseJHRuZ2vn6mZMANDR37G9N85gMC1vmXNjpc
TNoIFOxv92NTqnmTJQ/l9ANc52rEsKP1vBr7RcRPA1hifCEvOHqs37PfACUeZexlLsgBnIEXW/4E
BhEfFdFF+w5V7lCBP4W1YJpy7e40ofOPEBQ/H7Qbm0wX8IqBSnw2+M8EE3BnyzL5S2+xbNXqvwtR
pIRRYOZGvy0/T/eSXr9Ihh9aDpOt2nMuqAXY1Ylgth59mwH5dh/3kmrtY1ZKzmzOEnu51uZLWuVk
MBfjzgHFgsoGXvUfo9dwQKYtMxOG25In8GHwzQN2g/sn06lGehWQ7zMnWNpekvhIjNdCkOFMBW3u
oKmxOC+5w8PoGJe//3wY8G5xFP5bdbJwM3tKNCNW+fLFFo06Mev3eV3eUwRszS8+kIHxebz3ZRpp
btODeoKCZ4hbjulp+jk2PmX9faF5GkGDAIyml1Lmjfsgz0x46PUXBj0cpVcKmdumX7wLefh++whx
CBvM60f0kb4RIj3qHkJZekbLClGFMNQFM002jV0D1mCZPGz+ujcrQxvbaNLN4CfgKsaTEl8t5sDg
cM16pNTkFHtqZKqq+O62AsFq/zSQuSQ4DT07WNk+qwuC/5D1v/GT4rOc9VMPLjJtgMRegxwi0ir4
t6UZQTepwvwLmJ2wIRVtnJ6r6K0mEPY8LzPUcUZW7lCZECAy5LW1dKf75bALWMSYkC/NBap8wKqf
72lRU1l46JVvFT2jeUtuHlFp2XpbaxRmPA78VJXTx1FDZxxdurEmKy7xkkDZYtuZ0gIDUKkVdc80
FrP2G3/ExmMhSoxzxdfytT/8Nk2/MKB4Op+GGqzoxW7z3iZ/ipIO3dJb/G1uwAFoc/qTaHLo9Srg
2flMJtx7eXT/IgYfs4hRkk2/HEDG0RkInPbp4mGTEK/ImouDFG0ztV63E7GnmHNBc5Gj6vXraXoZ
ue5x2oaEhw2I8Ac5TXVgGg0TXVS4dgsEOd/2RPEXmOBC9J5/4yw4A4vJEY1CZormU5c0Y30Ed3MT
MBGmVV/m/wnFihLe++DF0SN3OSLlDLZT6svWj1ihYY/B6Vu7VrgVLsHQQ0GbTSYvH7bWYDnLd//6
0sJ0SLKVhwE9Lfnho7P/jeieP6juU8NSoW1u3d4L77/VVxv2ZU+oCye9PN4GBW9K/v9YYgbh+HGY
Dl4dvqGX7KwpJA77byWVFDgHSOaZ2AbvcclinrCoL/+7JV6izygRn4R/4AtAkFjV3PUqpnDzurjP
qrt0z3NSGpwi+1H+UxUN03Sduaj09cwQaVfmsVcOa6Q5pCR2ffUsd8Cv1vd9dRpjE4HSXkmIqEgO
ZOFnJkt84hBNzG2OdSU2AvKIWfip0X1nsEC94cBsUTNBBW0u1IJ7B2lM4936bQA53KSLqKl3wprT
l9cn3BFbbByX7fib4Ye3VLfN20359ukPzamO41HczbgNgLGJP3cpfakUNiV42MGfsFKYTZfL/XP8
JWKiMuRAQhiW8rf7VONn5mq20nV4TWnCugdN2ff2GIwS+8W5fvl1gSHVJXqMYWfNpNs2AkBBn4HB
3B3W1ohO7wHXvd0BEwyMubMpIMIrUg9LvESpVFQ80Q38PuCq6Xmah4Xb4/QMJUi9GjA82DDhAv1q
PFK/hB6xVxV4sINY/kPJ3Ka55EOs/W1yUuiffeIVv+CLtVmAQyCzw0G1+FEMCMEZoNyDQkSKZZE4
GevPr1HEYINmKcOFc0sV1cBf699bl+I43upShLP6RrpO4gzyt/wMxJUEXTXE4R8F/7TOWwrJvUfl
6Kn65UJ0te+ssWje9RIuWioIWi6w99rbBfM55E8PAOTtZxYln+UT1BnSi684yCHCzkWW1UIu3t9l
PZ8fzkYVLFniBHL7mULagGonZmWzTukgu9tP/eGvOMUj7bKvQtWF9J1zcDcT5O3d6aZm7/nmGEzJ
IwmqvbAxmnuWoVIZrvaDMnpfbDGg8zE1A4GeL9ciW7mDKJY6WNGuqq3IezR7sS5m7KB0uI/txJNc
ONLkVOudsF6DMwqmAsS5HTqh80SEW+xxb9vchbSocoUa3it6Mr52M6IFVJp+CTHbBbalKcmJLiPz
gMImZ9XTCV24GoLMtelbN50Uo87auDORsWmz0L7X7dkOxEBYD2GWQqQ+xiLcfDg0g/WewVIk+tGV
YCxWi49/+m4NG+krC2hNLJnq6mVVIeQjTy2JGMH1resthpMDIeq/H0CdYdY9JtZl8gPx+21THcPR
C886R0tUy65io5PSR9VaTTfrBH9tJRi1zbxWGrwaR7ghRdcUWWmrhn6//dtw+KHLVrv7w4mLyO07
nP0qJUkHIvyZEacNqkGTcKq4lr2OBvBXaXEUefdD9GoKwKh0EYpX+ho2lBfcs90a0eonaZHKWdMt
GrdRbeujV7oyeWGsbj2IB84O2n6UXhtWorUSP9fe443rAvR85yFyVs+31BBXcQbfFa2BGi94I7cK
XTwSEnCYKncEA6hQslRXJDIuPkXMjrvqwkLmE4XnTfOoQJJn/iTWT7InnMCj1pAP3p1gcIOgg/sw
o7TgzcL/IcMZD0UqaqXxB2iSJg0ScxHdahd1IoNXthHCaNVpLfzt0MKmp8X2U8qKmQBxRK/YSYEg
LZxZ2Y5gc6JAnqH0g7Qj+i9bAzovVGcwjOt0lgcejXunBQI1tfcZM3yEQtzFJvRamFXbFDCoTfz2
2W9Sd2ln9b50gyJFerlXltt0HKP0y0GSgiaENrMp8C8UaX/YHretxIOacjwps244U7gVJWrpbdgF
0zzZlwawa43WVdfkt6EQmv0C0BlLFX7oFcdW9OajBEvKEvhAosngptU2ui1nB9E8juSigZ7f+HQC
P8lGnOSQkkcdcVZDvEQXS/3PMURHhpBXNbyVvYA48wN/Bq53qUJ/aR4Oxi0DlNoEFWwhOY0aFLC0
4wFvsl/5Xe16GcO94CE01J+wIdsNC7gXGvJzcxD/oH0CZ/mjS+P+wHcPOKmWMR3Y1QOu9vK8eUF7
3cLW/jMDZhYs//Dk1z/TDytwDutP4drRKdqkg832I020KKx6BziY647JeeSOhXp4c7nvLJ/Y9FvX
hZkEuCHsBLlSKuaencsifa/7V7dPwG6HfJiT2ABebIsS+6de9xtUepU4rZyceCeMSLmLh3HlH/4r
vomkWlNhCn9lfYypYWmL5TnBX+evnhRalmyHxIqc/3pnULAg1ilzxTxynICDpNVJM/JwHI3qTCvT
86+GqlS3oJBPagvPEGRVzDr5iQShULJfaWslQv3mAXqoB3pINTg37+rzu6MmkSjYvhFF37lqwcam
HQEgsuTzURWWFe37fz56JYTmEh1bcLRWroBEPAejHXGhvR9nwMhJCoO+BZg3NTxkf1FyZloiYlhe
d9Nr4dfw8QPQhTSomzCJ0JlwXAt5QoATSiCPj/oM7Bkbycaipv8PCOc9w4xf8RdFWmDLuy5qNjcZ
q1Y/u7CYaDgOsbynBj8O+vtgOb3ZWyzcecuQf54/tf1Jbdz++QRsRjhhE/7NxUrLElEP4LR+EBcp
he/3xO3dLtd6Zg5Q8SC9C2JDkR/SezxxlZeosNNT7f4WxdbYdYJ5qOtTPa8cHSNGgNwrhaAFMsTl
NOi91BIb72cw73nZ3pJx+zU4fK4Wk7+uesmir5MmDdD5SHFp/zttpIXHmKKLLwpbG+C9HM+Asiwg
rZeFcF+Ci0vqP4kpMe0cn/Ods9XZvGEPyQyTGMhjNXuBUgBzoleJoMWCxEdyVYmZlWuBoGWmR890
EME4CiT/FVVHtLhqwDKNrjUntxjXZPvtNHLduYj2P8iD78sSWMm1jWc7JJkcWPVakIxhDQZcVvoH
QjCp452k3FgyLlW3MZXLX6LwqNT07B/eSskjc9tYiXlGdge0k+mbRFhzo/lF+eHgtRMGN+/nzuew
y5MHmIv0Jascgv9Ho3C8aqvom6Oso6mxqYThK3ggBAWu+KsY1hffXRptQ4z2m2CidLSw2OL5cW/4
JGIEf5KtUjjcpXvtT1/KsvuyWU41shJgtQdKwvkP6EOA9tjWYHC9gzb+QYoIxUQif49NftS3hfqm
FkT9Xj1O4LKlHEKtK1IBb9saVXRF4f8U0VWaay2eRmUzZ+KJGvDkA9wvRNAyUI6F1yFH62EDUc7V
hIaMtaDUIXFnOVY/4PCSkRaNLjyXngaRpO7sCTGrYTH5tjBE9k9XCOkO5z2K838tFs8QyLpWgEh9
klm9blqNfr7bj8hUaZLFxtnNEBIH8YydKWhFYUgJ8eRBFGMlUyEo+I6A8lDqfM5FjmOYws92aCHh
gjog1NkxSUuuCYzzsmFPO7upqA5YMwUV4Nj84wm/aO6mVM635vQPMiP5d7OhC/IeLctsrWsc8TF5
Icz8TKemvSAlTm25CZcyt0yPv6xWfL+043uKEUcxYv2s5NzAm8C5IIs990CnD2bltp7tPa4tkGEH
p6Kn7oZQhsubWlotF/S6bxBqD60ChhHS9+YfrBo79chVxj5JQoGA9YY7jDmMNmP79uCziVhNmA0P
fTig49o+Q4iW02KTQXiUlSI8QT47QgMmOaVeEP3eSixBoN6cpo2XrWOaIseR6M3KaR6xz2MSjFQy
00HhUu1rze+upNNKS1C6xrXayMSow+eBhBxJxv6F4sB+0nYq53r0GPFKJCiW+JytdffQrfwTkc+p
C8szXua7/cPJEE4ldIRZ9PUaTolabdnBDWU0woYViRaKLlqgKgZ5gTKhb6gfQGGDYzBtlPDmz34D
Un9PdyXpM+uEqiUJwmIfoi/l+tY5cwdXUQzzrHJktSIShP9nyuoh+GW08fndFrExfsKtStTzLwTO
VR/tLwaQbzeAIMhjNMOUeVnX0zj3BQFpZLq3hbjht9f6wO3FF7G0YbIKpqERvW1pVwgmoeV++TtO
tNeqRSWVCr1tBAtL2SBKN7SQlgCUMN4cjNFGtxrrA5k0J/IRvwm0cZayJJtRrAfiCks970AyZwk9
Os4s46/YyJxamaE4h9yYYF9F6g+Ll7BIYOckSZNrPFrONpkrgMJvVfmT4nIj4OUjV29IGNDvnlvV
SMJm4VlT4wvNpBuTx0TZJXLBJvvvFqLTDJgk+LHYfl2wYdkgYq1gVAZJAuazss/4o9h67/jN1rrp
Y2GMgLhQUpwGm/FKB9gclilQwLexTmA7/nQXX4vMdRHJBgAHvlF4fuk0sGIEBBUuauV76YzCxGjy
heWMcv33gNnfXye2PjZ0n1CZTjrP96HEFhTHbc5n0YACygQKtw2Xbm/uN6o1+9qB841XPFjGcHCq
XvcYQwr1KJpuHASAl1t5QwxfeGSvSI/JQxP+bbD+OqH0TRnH0gpm5eWo5ONu1MzzfTq969PnYUjm
ZjoMg2cxMOz/vvdkyaTzrbYuzKvghmYnMcqElZjkKbnztcZL89qRTXCXCotXj7vo4Gmwg7Bjp1jY
jnObTtrvr1KeRQQIezmFZV9tofhbkx9I/dIY7pjuqBQjfdPeM8RAfbNsuzkGM7F7Ymdnii91w4vJ
vSS6WCg+x4UgvbMmBn4ta1+rLHWBSxPGGK3iYd8m7NwEQMMwO5zH45KsEOoBhS06QuUfaZ7IKdsN
aBoxORE/qIHepa2t564xJqZl3BB8ThJNb6TG7tuCg7oSw+xSoNYlAMLaRlVKOqauZkdqwa/2k8jU
TR+RkTi+JxZGLs5l52a5RiQyBedGJ32DdA3ytTBvpmUzCUMu7JMcgweTQe/JVLqNMQLTXu32AjQR
FuKjQ0tKHQoLNWJHZrc+YVitXKPvks2u5rdeMn4/U51EvN5mfpguSrTNLXVLUddGJuO2/6YHAktY
buNW8eZ0b0jVX40i/9OHPq6gNNRGSWfTY9epc1aY5zAGsvjp4BgB8X8GF6WwJLC6ca/Cvf8fFIK+
aUOGUYtivP7qubVM/yUk8amalsqLWIomgyHWSrPQymWBwsfHdQdLo9Yaka5AjB4tjWbdjFUxqg4/
mS7oUCEI7y4zDr5LZAuVp3uzi4STKKERdQtiCj0MRevqn1Pv0A/b9Vo2sLM5zrT0fVs0UdEcAEvs
/QTVrC/kfxRBRtayYdQyl8fG2v+empLMySqePSg87xsw1jKGvaeNrDioqQUa3ftjoYnuuSkd3FwL
PkOUKLJy9q2Xw2/rDw2MQWS+BoEsZmeODl8NOSqlBm/QDglQDlRZkspfh+kLTGNG9pivCwrrtzJX
WT37yPnVn3t/SneT0H4fY6BcqFHvs7O5d83uST+oEJ8JTRTIj2/w2oOYtTMWmbPSlzAC6uWyCq1m
eG9x4JSmPJqj9Hl/mPIKJ30DEU7Zyd3U6SVUWCnTh6ndcN1K0OXpsQX4HbLy3rwu3Dj9pnQDKkip
1PHvh1At7WsyfllS3BOmlM+967sx2OQBvtmOLEgQ0qSTTBo3JMsiC9eypbFmYwv3kAQ7EHRmKD36
LCMmkCcriRx7hEXgU9Mj15JrhMpdaqt/Jdgi6Ilxo0VDzb3mNDa3+8ckh0Kp6TJ8cdtATu6YHjsH
zi3Pu7SCcRVnWcGwIXploBPdsV3SMZtTEhmHaytIn/hkXYJvp0zsSpD1xWWf/1pHQwBlQnnse7G6
xd2V5eVQcl+mjzSrbfjHndY0jvhAiVl/VTO5d+hjomsHzW3ogOSuUw4MjDdI0mI4+sw1FKTj8wxD
8Xb3shUGV4GBvCfcG2ycUffr6gErfx2t00sH/GzfXQLfmadsQr7+Kzu8ZwQLhA7hLkcQWbnLSgpy
YzpEtfdLHYakcVhrbpCLKj+EvIYVTaKrQKw1oxTbI93K4AzmiTCzSFdGGKP0kxnXTkQe6KteOaRu
I11F07z+/iJ/WuybEPMGxUi6zGVM1x5rIPQcZiS4dVyMyLVDAd1N4PQjiDg/8VBj66ht94uk7Mea
XSbODGPLB8tE4fPzOl7/v0yEYnR8KnHGxff3BmSkTS4DjMStH+8rIZgHnmCW8q0l1hCCzKXpn6tk
Y5dFMMH6i43QfqwPGpMFu3uvzhxRIGQ4sdF1lVCPax8ZIaKH2KsEQpKdeObKP+XiqqLh3f6nE/JQ
g13lkb7gk14KBGNayzvVoeyPRzmhI81Jt55n6F/r1K/4OVVsWpnelVCk+iUJ9EpUTzY0cp8J9TqY
5qlgz4+TsqFS9qpaTgKGd7OvZilzENDrxpR98VvBpStaWBvwGDqCq//sf8MvEiRhuADX7wVyZqGn
Dw4VU5dNjjuQx/9J7AULeQLcOZmUduqHXEl6pzvX8Z3E/rux//tNxMyjLuyMvBltkl4yly7cQnQz
Q+JoeMQtDCMKAAIS7ZdxZmIDpgHlq3upviZUXtF0y5DbHynS+8rOugTkond+TgOSXZR4xwW07MOS
+QMjPVHxw2IcBeEwalfnmbm55fhz6zrWtMFvA+kVm1ZEgW3HFfHwP3C6pAby8LHA6R6e2GX8xUIz
jMkryEZhbbFU3SyCJydRk/E8cFwnFO0WjQ1wqLstPcaOTgDd8QwB2yjKENQQwJn6qTdc+roGMT5k
6pxzYmOLnfBb/zJOqXEPgRt8JC9dsqfh60+aorauErkMJ5DCknpi6aYQoY+rXpzQxnIdmjTBYeWK
9PxWBUQSeBcWndEE7ZmskuteGGqgruIgdQG82HcEkln5Nttx3lkQW6Y84QzBdM6ugBayGCtNSb4Q
cfH69VPIbzrlCa86kVbzB6KsjeJUCEa+seG/cC6rdRziGCq8+uAhtS4Rfm/r2GYKQ25a++coXuTz
IymTaimmFEbFMHRHVpuPa+SiRGczsfQNEkYedHXT1HXqv6QYU0Te4aaO3zuaiUTSwJOQVnjjUdC5
6latj1rZQ0qbTKyBkWYfZeu2PXMrtpp3d/8NxN0HLi4nOmP9NCpqj+7NYqYS5hZLxZoFZFCc1/k3
tHu4tetameOXNHyqGes+Juihri7UuIQRauVJYaY3nC8Omhc6CwLVfPyMlYNVkL9D8fjJ6zc/855k
ikaEw6wzeyQv/3bNGQb7juKwLvcXCJkwtO1bN+t74pZnlB7Is70GDc2nVZdN9Q+S5l+mGF/OQulR
VvKkMwQ5uvK5MPszTfu5pVznzknjIRrN6jV0hrYhwhxKvFW+3VGZpTizp92uyecMLpNiNBCRsEDU
gIaegD47/eMIiYIucudmYWjidAkTib6K4OLV2RevhGTHzInKA9hvWK1ySDOU/D0JkP3FRiPzB6nM
AOdYOXkU5ULZA+c3ok8lOpIKuqaKEfXnWLIDA3InvYYBucZI4415UAMlfkT7X/1m4Ny/jB3dWMqB
cv80+WHfYdQrgHKFFqFIXobp9cAzzPftUhs5P5Wvcd9fq54MIH9Hb4fMwD58T4VSkU5V0i1kIZ11
oHa4WIy/r1s1GkOLOnJ9NJPMUwZ283Wa+UT4S81vN91VWOLIQDRN39OLKlwVsbaCGjXZJVhFM5Ag
k2tLIxtH21QfrNiZMplhmDJQISDTFJKekVW2Vdee3r9uXf6hpy9sHYDIJKn69r9bbr1X2RMYs55t
kCcRdY9BrdAfuJIz7MwPRjsG1m+KYFyAAGJIlrJPrUP2sCDC7jWTgLB/pZ4EJFkG1B/dDdmhXIab
HV7NfMwjBqLYU/5hsNirFPcI8BZTuEj0daUj/kK1mwiYoHnsOU7C+SvUyrAhbQQ9rUJor4PTPnX1
UbJu3Zs/76ba2VGYlvHnzbVMz6foNJoWuEzRobEs1ZSRv+2XIe7JYBgye6Uyyx4zcBWa2R6nC6Tr
MqztTuzhMacfz71k0o61l1fArgjE0i0OahEH9FNNTxoOhIZaahJuaslM9Hbfwzj0vGbG/H1XxlPJ
eQDYIPJbwuL8hOeASQCgg55VkT5RsCBFsyhJuko61oii/MkRU8FXnwdlyKq7Vsjof21BsCkS+PQZ
XdLA5aQiCo7k8ovji9nq4UmfT3VLmlldqExTEm8nP+AW0GBeIxL1kUCXXWw9fNFqR2YSRubC7HWy
QaUqUElU6cs5sVur4xO4c6xYJwg/gh0K3oStxc6sMgVSsPogpDsSWHLWF++9wRDJeBGkrhA9tDbt
RY6fdOmi5e75sxDO7EocUDNqztfPdhQrZt9vmhh8aUPQsG771fTNEDfMp5qvA1lrbHdA198rm3ak
TuFwKgebMgfY6sOeHCWLUdQYV5QN8Du8uSuhRNFx/LiF1Ii8+xr6gJAhLOe4pbxbKtkSW+mA9gar
mJqaOGIkFODHKCQdX/O9ayjVSarVfR+odEosee5PyYTP2IpHokT21KOPGf2+AJajAjskpi8nALv4
BXFHovCtWAANr3G3jvZLAnalwlI9EebXIkDebbhKh/r7GIKRx5rCP44B/I9m3vphFFX2T31CXSNf
ptQfuPnKd46X1YOGSVAiHtHq1H6VxGREaaPKbLNXMYkReupsvOabM+MBVxf9se35du0ZYYoFPiWl
YPvW2tLj+cySeeExp3cjeAh6yzScWx9bjoUiacRTxSHcZhnt3mh5PNCdTpmKjyIojeItnhq9eCLG
jMbTfS6D7PWpqopVmN108e7k8rUiqSq/MnSD32aVAi42EFUI3cjwhsj5X1zCHQfTe9ix6YQtW4R1
kH+KxDrtbSY3HQ9dohJkUZHaRxs8jplEZLCeVflhGuJ5sLlN7dXtswy9YFq08syM1ZGhqPaVM3Gh
Uw3VYQWamj7nNnuW89vjkTptVy44gXKQILoFdHfbIdoozh5R+6EZzFriZ55N4vLhtEaPnK6EYFdN
A8Dyy29UGAk+cIoVVqclODGguV/UZyRmpA2hr2RWHTxRpqNX1BypQYwR1DZzSf+UP/JTeJuFEoXN
lxOBp3JSulu8Wo4lb0Fgz92/E3BXtocUZgAA+KbTd8vS7TGIUlP0DkAOEhphmAtTCdkTZfurc6AH
VgfXNjxr0JIRs4Z/KIYtUZ2CEHE+irBnSyYdpQviKUx9Ddl3awEnh4MiJ5iBcMZFJd1uJhARgw/3
cMPlozFBBKF+KIsONaap6OYNuZ3KiUR52ZxneJREhzjl2wSjVbxU6KZm2ZcLh3eGEkJi65JHmpOZ
GZqgi3Dcf/cGLWnkzf9ydw8STwAEMi6d4uyWNG8mG1yG2/vd1nO4mAX1rUEErxYpFsmuEgfbtnUk
PrmXJ6D2KpMlJsG1usxghApvs5elLSPR8ks4fFStc1t6JBQ4btY3zs5IaqQHoIHMmpDFlipr47Vx
7IdjB+GddBr86175HLak9idrC8Xhlgh+jiBmgrlY3G2HeYzPR355TS90t8Puk8QKqZkzLGwN3UTa
PpFyAtn3YQhDfezCTXJHUdbN30TyvQnuqcEoS7Z05Fkc6o1c0TrgXCv7lmwhD1fvaHLjqMEwMjiL
IINjYGOkkSNNlzrAXUuNC0DoehYMQdn62FHYFouhfOsmkX1apNvff+GLFxmtuhmojo3ONXh5mp/H
ZP7md3MOspWwZaAF6NnacVbnKfWjpImI9s3n015K82dsFAOv385mSvJMSknYbbybfvXUtqkU8Xm6
knUIijH0YRCSUvUr0m47gI+BV/YXa9lWLowUy2jIBLgf7j0Zk58esjGFGlvAyPtByBq5LH7BRKAZ
unf6bCdOji8GaDwX6gUQyftRGG1FLVXFx/gpbP5gYgs9cocmNm55YKoxzfjkeGkrmGP0AReUD526
LAcnPL52GkXUlaoSGriO/OXI5XcmOCB/AEWEY9HY0Um6symrEZlMT3V0dXMOzYNCAYLMxTNRwvvH
xN/0kdRWf1VAEnKj1jtMzLiyW5GYRt0jrAvt7Xr4Gn0dvUYJTpv1yUPl5fzn3JqhPQdTOaGHjb07
jHsAve2NAivDCu+tqmTPkOgfj4XxJhCRSep5Nt+KBOsFVxfSob+2xdmkfss381npIj3szdWS5Fmq
wrDR5JtneAg66TOUPHguZJbtCVAOfJWD0Tjp9+vZcQ5rfq3P/7xyvdDwZnwqmw02WD0zGT0+ZYIL
Ip4c1lPMF1c7iVjS6gyAUa/UbbmcQp6UfBBz2B/i5JTuwdOqx02NkbEsCyG+NOG0b3/rizEAMK3U
ubeUvuuqdCraHmmFJ58UP/RPUNdhol0xQK/H97gNXiLRiC6fWTI+0fLsn7/g/85XNDti/1CmJstQ
N4IHYXFJrvn+uqPkuGRAsKhOl0LbisiLPdHmlD0iFvGCAXwtjTA5BM8TcvB0aIxkqjHuUouzQMkK
mEalRwLmLIuziud5EgcHYQh+aaZbSYFcJTGR5PgloI2v6FvwNSmjgJbx4r5rP6b8IQzKcwlnLUZo
h8gtOyDFzE76MiGUCU+j2byIaFpEukB7QpE1if+/6H/T/mY7zkFhHNzp54Pi/YVqNNLS+WaDnKV4
PB3I2T5+rEX5zYx9ao/suzKiTqTrVlAgxOo+XIpH6JRrb73yOR8sJbSzSzoOD0n5aw1jz1UFc7we
Tn7jzRelJ08+vI/KgE0uLZUIftUzLYu5F9Mw8qZL9WXracnjBhp6osScRB0GWyrt2kaZEEjAQh9o
3TdSXsid3X0Pt2wi2knOTz4gTLiocJxl+OhUNsCC9+WJGkZzZogC8r1DeCBYWApzVdnZjcjMUYlX
fHjmuTSZX4lJUNRhl8EhRZUnMrDN06r3v9ONZJ3SbFKanBkWObXUEbEaNuwbWiHsl8A7aGR2LcJU
lxfwMEBpkdVUS8Dcb/tCI2ZOvl8aLJUvttQUjW9ZgcSJNBQTj507CI6D/oV/5cWPKBQl95b7kQWl
eZVe3xh2BS0u0YnGYv1uw3WzzpawkFwMvAlWICvXl2QJjOZAnEXyS3BN3FEO2Xxj2xLPec0ZB9lU
Fbzxy5+231ZJnukKQgVkTjdEhM5KktVp8sGlvlZSqNGArYcXpbwFduPTglU2473RUQcERkw8nnPc
L0kUAr+FZE/M8GC5wQSw6/Ah2SLDXlVPGKP9AQSIAJIjze0vFavW8kkYpEIZBoh2ub61kWXXXrQ3
AYRbfHvEnSGtrs1dz3XYDlqFgROkqhYZwIwRmZYXbiSHWhNf/QTCeyjLMYEx6BF5EyRoS5i/oLrs
Wbk7uIP8ZzHxkuMgmLntMWBSRFdz/yu7OcBVQGXfFnv6w855GhBXJYPmNBjSATwmoJmBk39ulZHM
sDcanSyjK9eLRTrp70O49SJJZU+Bqt8wLbwUNX3/iH+UOW8AnlZLEU9AGeUllQ3KWYLhdHKpGxP8
aIEE4sETaNJEO3Wbe4SMBYGhyBSDSDUlmdtR363UUqzT3eUKb6o0nfjmMEs11qcPYER5B9Dih4Vq
uJuXDZ6j8IK4jukaFKa2AIIXi+2jvfwSFD0YRoC12/Q+uyRlKrDLCGnUthNC4SpsgcdQ3jMYL+Ry
33xXWL4m7CdViQDAWkxyxoIQGkzOQ7agTQeavGLTPOBgzhhG0x+4mtvTL5Qi1bV9I0mHmo0hls56
NPoyoKW2B++xvNBKdQE2hsnBYsUx3b0uXnQC11mMTDUeA3pp1JHF3i3u05m7eExrfxkavyuA+eqI
FWRn6fML/4YjL2Tci9HQBEMQluFZRvvE73JgnCxuOgD79wSTJ4U503k2gQth/iJLmAW+KCWW6TkP
VURho0hQIxtHZ3fvywntFxbZknlJE5Iv9pyyDuQxwIL5FcmovosBEA/Z+ke3ciUPnPbWRxGNRJAW
fb375oDdalAMUJK9pgrqBTr0C6SvNHVwPi1tlD74sR6QIhntVvL8V7YLC88IPFNeCr8zNh+3Cx3E
S3N3Fve6yO6hixA8KMqQ+bjD8HRv7xyKm9o9VKABECBFIH6vsXfJnL5vMdNTKaovjD/7pXHlZ7hf
OjOsDOEFxhzKwTfCPb6s42lmQLl2+2yYevtq8anbn9bFFzMBBuRWTQJ8CToWdE8BiL08jkpG6cDd
YFC9dSR4V2fNcP4MWx4FZpZpYuMJpeeUt6S6j+ijItH5dKI3E84ffhEDMaznLv+Qgjl3X3a6p3To
Sao2LMHXtXl4kCkVwdY6BkdSeRrLRinRGS+QASm2acpcUUipRVjA/IIQk7V+fvR0FdH8cWbxr511
ib2FJRmV61IeVMTHWT2XRxHAdy+Kt00TXSZo1iN1Pb0vAZshqHSeoHe69SCC7tZFNDS+NZxmCBEX
aAsCvnWrB6ViCnAkM6r6Ls3gu1SeCBdSimU7bi/mgh9iTEG6ur/5G9F4g1vcL1xHboVcAsLjE3On
0R9QSMkfgxH78hjav+iOK1AH0d/SadG0PsPgseiVMMTPhMIUArMWiqWq5rkZIFLGeqJibkZjjioF
hre4+WGmFF0TDqQ7exDLowWu1IrXl0j3iEz99oqmqkF0LI6Ep2edrx+mJEG2/rkeVkUvn+yPvGX7
AtcrO5jzbw0PpgqskOxlhl1lEHSRo4Dw6wxXlkz3fZYCXYZqK6b+C7EoQuI+cOIh0FYoRYz4/XBn
yVsvdf4OCeQrdgOb+XRfHlGXnkBKMhXTnKXMY+g78kczFY/ENVPoYvUZF1BoBJgazVutTjpc/DT3
Jtbf1IxSZ15c3pzQtAQ73w8ARIW6+B4mFPvNujOg0c/WtuRO3LRozGrg6cAzv93rMmsG3+l/6dEO
w4fq5V+vUr6k9ow4VRLe/u4KHbxfE033i915GGoYA5DlQhvaxHEAOa5eGy/h+eXVDF8iZqAdObBV
7hl9uH4yDoSdNNulPpMclLgmYW+WmM/61TiXsGySgAyXlzb+1qdU3GoXdWQ3ms6wfjSlNjC4zGrs
SVzGNbW9kbM8aPZSnJCW3gLFIDJOqypWDYgZlyGW+pnankLQm2RAucrW22GVx5eFF/oE7yMSPZCM
DySmhfXjU0lqj3MrEG/IAYUc0p73k8PvVcB+Me2hI7cbPdW+q2nrjqTQ//wzjXTRXv4eCc3Z8njB
oZeaiWr15w+dAjlp7ADdI/1c7Vw4PZSKnuse4TMgQReBK8Lo2QEyRbDNm5kUb3Iwmose3JnkojfU
f2NbyW1X3w7ywVZ3Lpr4MaBrH4q7A74qW+aeaelPM/3goJNh+Kw8U/cSAyqIqY4jgdmqvSWJ2cBd
Jh7hTrVIPTjqRpKfZKnNOrle5Q1oma/YD1Nn+V5P6Ekp8yWat/yrSSpRw8iVzRYLlWpA6TyDi+2y
Rcqjp1OPtZI6aarxnVJ5h0apKLo2KqHKAJDuOGy4ej1h6B+io9q1GACP64gbHKkHYcCUf1ElQZK/
y6DGzT+nlkuwkTCjy8XbU7R98d85O4fuHFcohdI1l80jQcbf4dml7y29kuqDWRxIcRK9KTc9ZZAJ
g3ap2sqrJFbG+4Hm4RTKyGh7Dv1luJe1BZfQIoEavB7UkPYq+Xu0AyDDhunkiJajB2OhCxrX18m/
5M0ANjbTlL98QP6eyuvrEf1Q1dJxhOKMbAxGubzL/6oISbcQoMypZrDFoyeTWWIclYpoXiubUVJ/
ImSw1/gIkhn3jsJaXYW8/Se9d+2cQMrras7RRpuOdF6l4uX8MmYrY7UHADzjsXeDjULglAPZ9dsP
F3gOHPfk23iVeOUxspj5s40oQEpnurKGmg5ccVu7aBTk2poeDxW7zVD17rPZfgrQey3/KX83tXmm
F6AaRa1Is9vgcFubw/PASyFMYUX7GU4/3QJtHUGvJ64xu9WFJGw3rgEXMiF4sBvXl5OaQSkB7z/l
ElbJA0y0fwm0Vnewbu7oXKBvqpqFeDxLQ2QX1FheWui3SePlzvmoKrmgMBzZfGBxer4UD2qhjzfj
U2SZj3BYpyas/pU7QC/2FTU0ef/CgxvVGGyJyILPZzd0Db7RaizuCWVvdJ1SwL9ClfdigHsMxhly
1nFRc/0ihpkexZrqSq8BsbpaWSQDN5oObTYZFeRidiEl8C6tYwcB4eyvgt/0M6KS61ezp3YKyHLq
D6aXy5SPigZh7yHHOrPhvYc+IoRXJbgeSC7hhMegg2gaPu+R+NjfuLj2nHJuPij8tnYRO8Iucylg
pxrcC4JYCYspJ0EOf4XxQNrO/IDDu7eHYCp2LkK/T7VsUbeBx+afudsm0Cp4pBpLlLW/79UZpUnu
iLjQrC7asCxbXw7OPRPjeHL0mmNgYXIjHIrIVJ6MS2FUHqspgybDgakEsfCY2jHcTVX/pGiyHw4b
qyQZ3czHcYwIaPGyYvFJ6DiOu7JhSPmP1Iyy0abapWyRZJ/EB4+intKUcExIQUtx9OskPtewcy2O
M7BdfH88HwjwpmPfHq/7iJPOS7vExPnOhyryxkYSW+59kN9TzzrWfE3UI8DgCXcJrbJq1WH/tOEG
ewYJE7TyOCelIkHXknMuP55Z68IswptsKyWMJDwDGHZTZPdOeMwPeENDzwZyeSBXZsieVVSWEas8
Xab5v5r//TFNQDIPjOwyPvRxcYQMiH5p+laaKtaH/PvoMtCcwKGS5RDWd7vBdz0ngviZzgqowDXb
fbxcJuWjpizjQgofgsaM9Njaon/Z5b+8n/kZXvsUHyHaS0zaUAhnr9Jki58SmXNgGBFt81ocN1ek
oY7YPz5ooi66p+EQQNcM9KI9XfZWn/pYvvXPYysQ+xez1/t66kfW8cObjvpQBvD3/Nw2wpJLuv2A
nRPRUZHxP5kdSlydu2Vw9L7a86OrsIM1e6T3LGN3RmLDMAKGqmqvFmaoPpHwdfgeLUYV+6etLkck
LEYZZV5gv30o7dwW6bNFeBWtQv0TgjKCM7m/nHrN/jwhhd3jPLHAMWX3WhdrLjpHGjH+TBMj1ZwT
jXPLKXEiav/Sw+9oN5AzD7vrdScOXDY9VvgxhqeCaW8pJDzYX1kZbY7/e1Hx1vC1zIEAPD9q4dJn
gswG015Y1q/meZXUVbExb+jP/08SEYACOEu4ukV4nZSmlIiCL2tZ64+NF6ojGKsLAvSB6BZTFpgY
jKcB/AvcvLonqJPs9rVfZd+DO/TWW3/yt/8eaUSX0xIfBxlhL10uPwPfnz2m0bauu+CpwW0QbasQ
i0dk2fSBt3MX/jcUaYeV1mNjE0NIOvSgwlcj9P8Uq7M9h5r/AiWHQTT/8dgmEODnxEoaXQ8+UUmH
g3WGDcl49RiX6kfaqfBCPYQzhetz80Ju1UiwlYg/1x76in+8d50mom4XYfOY1CssjdfRkjxMf/+5
i33iqJORSigFGHyO+vko98s1OCzWuNTThzo5UVkFqSfNDyHouUYldkcZ2/CbNG3i+/e6pepmmBbQ
nPofiUumxuPwOUsZZRlzjt2tjdTJXtcMwl4dR+cRLaTEQmk1G43GOdEs+X0bpI28MOyfRnERPkQG
gs3E7ZdQWjUDpDEKjoBOkA5GpF9fRzyAfSGIvenhgC0VkLrQaFMvFUAGVWs6U6f/vddrl/SmfEBP
ot+2SWCbWVKQtY4VpPgUcCGBBGzcw6cad6dRTwPMeo1jel5QK6aKwqwIZnC0U9CeVz1/35qTL0kn
Fj8Zi9d01GHfJXMV6y79S9gv+Mii7GonXjBShoFehKL9xM1RiXBh81AHNV7b98ZpsbMM2rpjV5i9
v2TrW8QOtBijzh/fyEtISujslU1qoasCRwmwgkif0p1l0v0nRbIVbW/J9xSVGYagQlprbspLnB3Y
7I8DrBntbx8gXugIw9rCkV0bHlmGYfcW72bTkBZRvtOMFf3z136Mq4inFkeMqaulSgWo1c2uhq1Q
hNBHgq3kerv5F+jd5xOscyuww6OLRmPi7S0+b3VSlW7GKZGUr6Qvs1Lx2WB+hfU5OhxEgxKflUCy
yQrZ6m8G3cy4as54Nc0r9AIlJV9U98nIpasDB7UlLtVqhpPlFbY0Byt0PhZjGKgKSkxnbPv0UmI2
obpgQisEgV2+EmGVX8Ma4gxo9SVp7OKyqf95O8xY7ztJ71tFkzbDOABbE1xWDPKoLU8jXhTNBn7q
cDQPrwAVbfTAgC72Fi2ZESMzrNBSef0nWyQW9VdqLDqf29YIKjxYEn6AIU0ENiWd72JXnzldbJYS
sv68xi381VlGaht7Q+XHjaBQRCVeqNmlWUTRWz49mhwCkUasO2ck3CdpnW4EJzgo8uDeM4rWuogj
ZO3Zrkvv2V7mZQMmNzJAlDnZJnRpMYFIc6fdR8oRi6ogZ9DpbfCwB/ypHUaoicGzNKB7B4ESIHD+
EgqGPh+ZP9Qsr7z9KsfVxdmirKevgkyWKzEz4a6cQDf2AwdivplQmpLs+OfdPuc3S54np4TewqjJ
0KJ3w8JUPIjsp1MJRAPHyRGOm4TtgMT6Rkvx2fB1OgZasBLGN+1T0vBdueYVBK9AmyH5Ip0ORCkC
9wTXxn9+xpRa3bug1bS3cqlbNHWIL7V4F1H1rYQEW8EaEQ29n44m6Rpwjp2DubjlDB5apA+8O4bk
6/7Qo6J7hre+ZlGkprpskYIhWu88/woAOA/SkARFxW3kOPYfHm/XGx9KXvtiQVzDscZU7NVClRYR
ipxxubkMDVQHhkPZ4ZLqJsj0FYY4Cxmk8bIcvZl7/HjxxkAucvsya7cbmLIMzEI2kAD2chfznU6D
KdC63VgmppJ7VHqEb13xUNzUrRT8sByiA8Ku+5PC3jiydjtnZ0h/3zaP6xBpvxNFraz3i+nI2JAX
8d90tSTKENrozpu3mgNj7srBfEqZb85K0XG470YLM8XXEJ+g8ZLbpqqo1dMbNtBt4qXZqH3dYdLy
ZpUxqRSyJPFB0910uum4p/AnzQCJpx/whJaF2/HTGa2FdnS6ICXC31Ot9cqALX8yMO8DxIGnPtv4
zqjhdzkQM7YCI7o/PZnbykNJvbzk9jmqm0lcM+SPo8GLasGMLu1b7FhD91eX9CluQi94EA/HHjjf
zQhcsh4EBPRcbtNvS78qQvn/79P+9x0X0liTfa7K+bjOnISwJ8ro79CFOMPMF5AsMY3LxDTN0cls
EcJiB+TsbmXzuWUBy9VVRMXW16WxqsqQjbf2yUl7u28zfO8zl2yrNpkM9s6rWc/hBLQ8HCdOqSkW
YM58fbm9QNYPC3JmlMQbaML71m8Y4U3jcLiO8ihKZn29ww/WMd/pwoD2VK7o7L3rDDQD+F+KsQWQ
wNzo+ne07lg8UPULcQsw7MSBn2RT63cXGvGu10/vU2UM1vULtwubST+UgOW8JZhFKxl5TgHcbdVV
V7QOp34pHOk1IGDJexSHt+ZnPV6nhJBNAyNSU/jTWRgSj/6xcVK1jKHDiwCo3HH5DqsYT63HA9Dl
gr5PGgUQflbHQnltqxySjc9M04725lZ5H6CdClgajEflAzkuLy220k0e3IuS9QFFjfm4yR7K6eBQ
kfXUt1ztSEjg+VRfSQOf3NSnayelliOqKU03FVlRFNy5FMqNdw7RJPyb/n7lpl+HDOUULJOLUTt+
eDxQNU7Qyuykz0wpicuscx+QOb7F67uqx/3mA2CYWzKuDDOzUiXMs2zoBBpVRHwI/QR1nCoPC9o7
po64KN5w+lBt2Ueu+rY+DtGP7WvF/ogqMl3vC8rCoL+lDdp0OmfMHlSQycNzCGK+lXlmHwmnGdYb
1UHikRjjf1wjX8wjr526xhr/5PJEayqLmr7+pSwHgn+6nLgYCUD2v7dnjs5iaeHTUVSo++FmrCol
eA7ijSGa98KwhD/XM5gMpGDanRNjKA6uaoBm3snjBkYPLKfV16XoU3toIRCFDphqxfWmE7+Wzvxv
Zdg5xEsal6wz47QP27upK1BgpnkhXRglIyhA7056CNzuvkfAnPEbdYdRPASNL+pBVdz/hKqt2G5X
fZ7wmqEipERh6wbbhnrXYwa7lFuXMe80NdDXmRxkkIK9Q9pg6RvCy0soHEBFPxZUDt9OY3CrkV9S
QyTvh1ifzR1BTKUBspKfwsksZ53gf8vrSxsyQhZ7yBvgE3VgPoGcPjqlnvqo9Zxw2dV1N77Anc3P
5Cx2t5HfRzgAy7ttUNftdfUBKILxbpiRWVEFkAvawV9Im1CWitGW7B53B7o90d9erg5TIDc6y0fU
TsncGNocIfoa1l7Yvhj/3c/xyVg8HHf7rdFzqtY4DwpLp2r43FckDGzO2qq48LeeN8+5Ozn7YDZV
ICAJNB/b49XpgeL+crrsIxPkuTIyKdtxxzeLke1a3oo7KwPC0tmk1n8tVhxhAIW3oR320ddSP9TY
6FdcHbqMjaJPMhg9DAUvx7nL5Mae/I+a1c4iQonKlSct3j7ZTtX2HrwowN3yBr/Lq6hT5BTqU26s
HqKlRwnBPnTWNjPqCDay4uRD4L9hAEOQhS1t4bHi/bTkBSxRgkDrXvzKlM22/hdZb9OClPrLqBZJ
00sbS/3hAlA92df08rvL4+O0MxtYh+7+Eh2q627jSo2s7yNjnznLEZrzGEh8x5J/kRWYnr38diAZ
617lort39G0+m7cJNznaCrVIVIBgVfl+lkK3YVSrXH1ruIxQf8QviRXWx375Lth9nC3d0XDbCIMB
4juHwvdNpdp4Vl2nh3XbFQYC+yRNsU6eCw13awYrptxNoMqybTj8YzV6whbZY57+E+C23ksTPmah
dhnI7v6EqNGU9DPdAyIFHAKHGOFCwlN/VGTQdxSEozLH/6ImVQ5lft82I9e/qZc6kSPRYhlIXnm4
I5YdE/9Ipp+ZCEn18iTtsp5AvSJgXKMNH0i4CeaQjbfraCjd3YgNrZOGhNnaeOiwUvS+XWOWhSst
lpKH3LC+wcqF1F6vNVH0BGK6yhNbYlVB9q0d7RrisLcQPTbVvsWWbzxuuAAJ1YJqdwSDNmRhZtdH
y2iZqycsANMA0No9rRdAqT1r4l9KXMipRbI/oisSa91cGfM/eeF2DY+XGlKwlNUJl+YZmDqxWI9U
Q89aPJm2BMWETIVu5rxRuVnhkmP6rSGu5KkpI9XcsuZzJ4xOFZvG9nbp2W1BzuLVVgUkNrYFjPk3
cWyoJm0G+mQXnn6AzFBP+89YF4LIYu+Bm7TcA5F2z3kALm6aPy274dSu5n70n5kkA20CPI56TdKc
69OplZob+rE8NBNPh0o3gE36BXgd4Cziq92ROFpjlp0I9Xkj0ELltQw9fFYmkl8zzzaMtNlOc6VM
TtwKk6z2FgFFLLlJ0p2nIy1v8fk0VzWPDqF7oyHR53iM4R87M0JDxgsZddwieypxDvNHdTkYd77w
gGgjwq56oYhaDDHJZe4GuxdtAEuNvTOgjHGdE2Ecc/NxQgmakY4Jx8SdUYqJ4vMBaHYhbDvdRwoI
0YlOtRvLAmGtRGfVBUTyR3tubLwcGhONeREoEw16cfsjwU+car/7Vwe7a4w+m93h5nljkQtVtV8W
GEr4GTj949hDZP12IUlA3xb2HxON7echkUJoFwW0J1gNafxEodfW0f7vkea+1sf+CxnjlVqVtbJl
11IT5tnv3Ep6ewHemU8UjgzZGK9PxfN/eKpWO9cgRpArYF6sYetLKME/HUdf9DLORf8InnSo4xnp
bvukwFP4oQ6iYt/Au9Ry7Y+OTFjT1OQU9QVzLBCPaM/5/1E2EAF+/hLi3pZITD8MobPbxsRbGWkK
S8d7yV7kmKVBEztk/evFbt+cntExfIRNlVLMZ7EPe5qvxPNcOpF8EYRROddxYl8ld5Gd8xKjxR9v
UoHPn1joE2VC+XjgquCkGM9aHdGjo+DP91g84K97lpKKf90E9HP+AetF01L4D5R9t4nXTmeNNSpG
s3F8qW58uXxAAQLUkjAQNvq7rfzMhwbJmiPwhT6uqURQ9vNozaKJljF5Zg0Jx2ZJ9BdFVqpjs2z5
N7Dz4bBYQqImrdbhFm8ClORcpV6ggaAXTJgMfEYgURcqYSKOpyKTbG2nQ1ppDDQ+Nb2gJ8uM6bxn
RbleHJqWDvDiFdfYqMFnjEDbEwv/BbhUWiI1rsnilF2fTqqxY5qoaA0nd5jupZrX05GIcJ2RzyGf
Zv/L6DA+trwXffylhxP1bR/AjeSAfYFRd7gxD3PkPfnWxvHchrS1nsJ2GnZo5TQvIRx5GOfHJord
V0jeFYq0PmGlt/YajEZ7o8/rmYmjI60HE5GYEWPQgsb1l20AaJAn7rMdxnoG2wJl4QStQQXaLylV
Yt50QD2am0WTp+k2yU3xpsPEysxTXgu8n9JUYWwhUfzrvx+mDdiQ9ORRfGXcfHQCWXPlCYeIFZj3
N5ywBWGoJj5Aq5YekV+q8K+r3v+etWmMj953P1q9pq6PpoyE+HsiZ+4q/juHsARWOlDUjBo/esxN
c2WbqVfQbyEZHpLPOMBETtb96FcO4dWCR9tVd8bV7YZMeDqZM6rmVTsXH6qYKKCttYe7RwAH7kvD
CB6HYcxNNebl34XdwLAPCXobKA27Te1HI9lARFpsNKm3A/WJsszBUrv7UyVkc3OqTOULNvK7QbMY
oR8pVt0V0WrN7vYeIllnQlG3NGLe4JDqqB8I064lPTrDno3lz909KIaTgStRACl8opWCrvUXj2az
KNrjc5JdKrFhKGCHFAQsfsmsbxqQK+GHAobPqSOIVKAz3Ca6C6jR89TdjVaQvHzxaYNFIuzz4Q9d
1vc5psOH5CtzL+qzfySisJfDq97VDYNqi2TaKv0NrG+aq9007v2ibFXaPJfPo+S2MqtH+DrMi2ls
gKu/jcVPyJm1D3l46UtZWhhv4P9t5hY5XF8JkL+5NwnHdCVBSs2CW1t6mzc+D1dIz2R2FKpx+0Kt
rqUcSceeoCLkSNx2v8pUHCOG/IZWpwgROqk4DT8LjLyKnqK6E3qxqbrqpKi0oTlydQJy367yqZMS
jLwR1VpUFnxIu8cfopzpmqgp03DOtrGm5r1PrmX09M4vSfEuu+ElBsBOvVEwBk39KKm8AB8/L7iY
v83EUqw8B1GEf9fU5BWTLugtHnS9dZHCCJZ/N8KFFiYhRJ+Mp8pGern0uoKWDR05keU0ij0irhnk
A3Ku1trDLMvY3MTE8AYn4uvavrhK0sI+Yrsx7bN570opdj9uICjxUM8ioyrMQGdWxv0BDCtw5FTg
rFhpB01dTevOJyXX83GI6oQHuitGvgrN9AXtnZ2Ad4N6HzXeeIFx75f0ElF8ntCCQOCex5duh+Lr
/RYnqkWzq+TD4I1aIG1z1OuO+SO5LNuib2dz3eztmOcFu1Sxj1iAvcpvjzhWxfb0ITNaOyIcrDUP
PfJMjK5ezibpNaI6pgIhOML1ldkUgN8qIcseax6Eix79uxMHkbzFeiMG54vZP4HSQwTDbyOy3J3d
WyWdaiuAQLpuRutdcEbwse79Icosh6fxpLTNK+rxo8kHqiLt5yxP8mcRFyUXGAt+781ZOkefWBNq
qjKlu/1TTG/j0xpHuImmlgCPDAPcRrGf2uXPTyam4mippcYVKGO3n0XJmis5ajAjOKO7ie2Unkpg
QbPd7F+9qxSCpjjCglxjeMt2NK8AV8LuK6+I6/LoQr4J8gy/tk/+GyNOOtT5HypqxSdMtkGD9uD9
RI9XQSgiXJ3XQYD9H/30X8L2BF1QLZwGLEuJ3tnT360HOlTrARvqVGGlUN17sj9DPI+ALrvVXpC0
TDrAi0DjPTb+Yaw8zaM8GcMl81cHt+N2YdM/Lftdi3IQmr1x7bVFhKkhCVeok+qBU3FR4UQndeg0
zJbCan0HIcihT4srL2u5/sx34A7bPBM2JAhARkqU9RLtqpnykn/dlM48QElAI5kkCHcjgiAYwMlO
lkUXnDzJtfDwSyLFn1wAl+mSWhQ4plh5j4FF/e103X9SDoOx7MUZCCODX2mC1nSPRHGkP32cDydZ
E2kPmG2wpOdNOz1sWy5Hmd2SvbpqMZ9ITBvYTgt9KqoaZkfo2fcFdlfcaAVmaPogFGSZW1PYFTPO
DrHapOsgY83UhykK4lfxYQVdjmxKPZF3wQeSPwISqfKPb8YdyS3Bs6swjVl+PoqPvIfjl6+DX2SG
/M5D9ayurs/NdajnBn60YYrzP0e0mUtV3NNO9HE+ao6NQnwHrIozeq9JH+vTdBztIPdvUDwOSI84
4DWM9J5SLXcTC3CZclim1c/btpFnZz1P2//gYwW+IhYSOaeTYq+NJFNeiWZaVKyTgeoXKm7oocTd
tzjmmDp754zSlcLFAmDhNBXDpXmGud8aK8osBziacjOgMSGk74wl5N628FbkG6ZT24xwdRr6jnjM
8BPp/5lwKyY0SeNPAZcwPPSEFrPkc12WGfLo3FfHqYwDd2Pzes2siB3tEU10Tl/E+SNWGyCY/vSN
Cnvza8mwPt4RHVy1VZizVyZDbqExxqQHQA638VkeivYLWyDPXkUMv/rm9ZIpgoT92h4oeyhv7uaf
PGLMcziQ8RM63Nrdl0jVbfPeCmRXRe5Cvd339EUvKRBgVYYhXFYa2gOe7614r9oC+8bmNMM3ml8P
296beR/nMthejHe5mDG/2hSSOb/wTolX51jOIV3uXlZJenGVXNSLjuFlv2NloRPCGkfkMjsuulDo
Hed3HGY/mAwrFao03nm4sqFrSHjZaK/KGM/6CkD1EArU2naAPjjQR+++I4oUetDo9M2eDV66R1k9
6xxSCY1IV7oBIjGgOQnnDZIR9J55f/BBLkDJWV9Lp//Y0ERnUZ4pQIAAVr/EgpLFHuUnWDYhT3SG
7ffABqf5o17lyRdNVHW9/VW5mGH1TsHYXaJOagEJmZSedPeiV3VNaskFyKN6Fz24LxDYrMC6COA7
dcmwgtya3tFVjKAeDHnoqdyGtA5OuyRmLNQTQbur3hMXnzT8BN4GLz6gX2qcDVNZ9PKthdlsMOHz
dV1OHerfbmLSf7JH6UABNmYlZXQ8p1pxprUxTiJToD0ZB1HZN2ZULjwG19tHNpkYpTQ6fAakqXvg
ovZgdAqn74FhKwoTcD8PAFsjrvPlsmgNOX7uvFJ//g2/8sO7uPY8bDEjsWoNQT3X2d4+O+6JJPxX
A2PDdsI9lbrDzEwBmvC23UurGrvqi3QPFS2jKYKD1qkyznoCbwfvzcuO1TWpPVak25g67xIy1Czz
opuSkqopAD+NpATFtKGwKFHcvFHNd5ok578i7oPXkNJY0cNQNbwcIuvjqZW7z6ryf8adFpixOTeD
jocC2u1+gOck24/rDSexcJOUqW0MR9vdpHyyZL0HVNTQ8XMeC2ajpD/AUzp4MoKks7ZVT/s7D98j
pjptL51lpomnx2IVTCTMboRsZpPw0n2dcuHONxKiRtXftPyYT6gZNpqTzqXu2nUOWieupxNdpF9s
FvUWGBvm3ExpCcw/GR6gbNAfWUxUmQXk/WD4oOHLo0in8v5+VmqlFPa7BnSVhvAS9q02kKRWk+l7
7ktAgzXYWQxo38I4Ww9YVaBEHUBGzrah7ukaQgQYJE7+X/ziNLu7FVsXmx9vxXf9JjoHq3RL4FN+
7NlQlXG8JPRwOV9iKEtD57M1TS7+Pf5lEk+Coe3Te+X4s2ilnj1VaHVa6n6u8Y5mB44uFM9W75oF
D+ZrW0i819AqZF1pkT1x5SpA9heTt2GSrPRGxeZc3HxVgXJvlnBEssMlliF0VwRC0/ixRqtkyz/P
8konQ/syzT4WzwhNS3Z6PlN2RJYb4a39EBVTTFiGuFJKTHb1/NRXkIJdH8pSvOFNCv1vMgyUx5Es
hUvEiNliqCpQi7KkjyrwfAgprtArj1qw1pa4k3CBqISq7CilYFdInmbiZVFnFOr4iUR9eU/v7NGN
/aOg8uU4t9j24CiByPsRRvhIg+kqeslV7yKPRmdKII4jZWM0neahKIMIKjjylXMFvH7D0wMA5D1e
lmNgPXPX1Fkk3puz1Ev6bvhghCO5A/02Yk15k5I13PAgL8/schTXjGLgo0y5PuFwJoDIiIfzU1+4
4Ab0CQLgxjgOYPxzRp96YumHx8++M67kxg01VYaMKzZfljDOtKdyk9325gIS5g8hKwnNyLlxmmuN
vWCYbXVW2jiypJ3rL8h8LclXCZEFS4rriVR0nAhuY0vuEvvA8Bl/7UOvUa5i12f5vKZGSwxG6uR9
QfE4ueQewtFDtePs0BEz9RwP7+N/71B7nkr8Bjj2kRsyCtM+iPooSFcC874q4BrcsMhCIz/JRJcP
6oQzfPgqbE1TKtNZfJ+TdYnvqDF1OJbeQtKBI42eTKY2sXKz/oczcfQ7mis3/v7mwFMIProG7nHc
rzfQPUAxmS+kgRr4UFdTsVmrPoailIKreXYA4mXEnBW5kwyzdIWJAOaMzZ0C8M3cebNHj+htIwn1
v6sM32tl7LtnE5+ejkbZmVlKsY4BlDet7o0rdvBCAPdXvoPSvUbB9Ausytv+11eNU+9LVSZqikeb
kY3EbLcsMQIVPwvuQMI35PqqBU+eCzb5cqY2M19K6XEsBpfuD6OQwtOybCDpLDkYCmGb4EBD9sHY
ZJRRwJsgsBvufV+9k0/OL2bqsEeNm1Ebtl6EZkrkf9z1b5BWvCIzr4HVLUMCviF30M0hKvU0JZUq
BcoQBvkAbAjSSot2AkzO1PCnk+v+UTza1iEFpMtusL3JnbSDZ4YkpleJ1EPincMNdLeixeTstoAA
JClb0fDwJCMNcCQpDSy0vXO9KEDX/4Zio6cTvpMGYDf+wbM43rZ8fFCPV2VjW3CDQkUxdPB64QEI
QYdJmNDKtGJg30FpgQSLjcr1Oey/AXew2oL1cG3g2g/Zz8ql0tcTuEqyv6BpN5I9DrHrEyNeGryP
O47SQBhV+6sJL5FIk5cF/Da5p82tuo8D7MBlb8OWNkutxhrhQTbi1PrlK+bUWpUBli8KmSlwlP+b
wF7qwTkIFlj2lYBA394UIVKKZX6OKQd2BgFicJhewCzied74D8qteMw5toJpfiWp2ECGXJsqYP0t
ElWjKyzLDTS/lAUE3/JzIOXlbUv96d7vldxiB9t3GgjpbQVlchtIOblbRl36CqoI1GqdsvdcqmwD
1szmOxafenJOkILsN6ND3XR9S5En0Fn9FORF3+oryZruO67zzUENy7hWbTCERAZsDsuwZgfMHmbQ
uUenFvisy2ULp793BsXORL4W4dqoBsnTroUeevTepZDnyr2jJ0lLtlWTlNUO7c05A6hHeur41cqH
rgjr25UoTqsmwRmEVZX6nDH2Q1P4WxJImEgpPB4ZfbDpLWEYDzHnwMkYrmISRl/WRKD9LVK4OFcB
s3G0KT3Fd1XUuY5d+MBVZrwakAg88woPiblKKoa2WtRaYkzvvf0mqNVSN96YxhpJI3l1bu1Vztjt
YlON+/o7mX1dvM4L4bsWSEAB9iC/y3krRX91x1dDSNB7uHEgYdK+PfQLTX0N7q7qOgz3mL3KxhBQ
WsKaa2DbleTte2QZTyHb0UNnqSClx/tpjwJs7oZgL4XiVCwOsEGU3GFeSa6Q0jwRDzxzzizpgDrX
sZkt9Np4w7XYQBhMSwaqbxYdakXEYgvknM0P12rh168L+NRTcnGqVjSrMdyojihW43YqD5Np4/xY
Rcm+dLGBzxmXQk/2nr/nDCnxfOvd9081wP1HgGZSP22x9Qms0gHO05zs0qHwR6pOkqIN8mGSH1ei
KsBMyjU3PNofVkKIFD1glHWjTYkEybUm9bpE+0oPczePTojc/a78YU7+Epz0TYdF85sYKt8MTBlr
ElkoFVt7LznBKVrAlAuCwjuNb1T6AbxgRIPH7/M6O9NQVPHY5Fy2za4RK06aL+7PVJXTC0VUWKOr
K/chgC9LxjALfWyvvNF4JRHpLLFth0MJZ9/90oia2Qsa8QHwgx+dVgMnDSs53zgMK9TY3gyqRMo2
82FQAO98pTMFSgArzCMs3VNHfMp+El7l/EM6zL8Zc/knDpqxrRpbmi6sfClylOPGdqqnXbbEgAc8
mrocfOdaCJpiB5IM1VuLmLRjzQZ4U8qwI5uBiJuHFJAwVokCLkUlU1D8u4rdJDnzHIkETr3Kxeow
bOpu3NYAlwnhNGnnicEl1PhRrq1ohKHrfX7kR+do9OINWr2Oi02qFvbBr/K+LAABGrQmwH/LlStq
eiKxrQ9jop3ge03/rr4Wc085Xx7wF11Ol5JXYmMOW3p3mN9M2uHDiqrr0233JVcSHi6WR5QujF2v
uOdM/SlvNJKYOyw5kfnIKJpE5x8W9Q2UPlIbfLiVzt8Ii/kw+HhZT5ms7pXL2OEtUqti8nXZLUqX
MhYMZPCiDxYMF+BB6U2ltm+u11/3i7WhvL8j0QY5A3N5gV/bYYb5yU3g3Yj597YgrXTAmna9I8gE
XMwNE6Sn/P8cDG+HSW+Zm4beV85lQh1/VyZjb/czKpBV76qip7vWt1niYRu6Un/Rt6h9f6T9AMuM
HvRB1PtdRQ+GvkYOWCqw1N4mR3M3NzGw3WYAmmovNxsDjQYimjV1s1H7ZfRja8GW0H1w1igrwMiJ
UpGahOyXK+53mr9+ii+eKD9v/R33P5hMSA7nymHbYxd0IjbX7WgPa3xUvkBa2Z/clXywsvcEIsAx
Bs8fNOCqtF1i72R4ua+WrFlYOt09HCg5QdFRnBb5CElbMbRG5at0Hr0tKYzJYAeOY2KiS3zq2Br3
UPXjC5YR6ifDvbPnX4QvFZa6HrVEHAsbChzbuHCCUCUuS+QHaDc/EG2g7AZ8cIve6XAa/jH+q+zb
/DHSxhfpsuFs2XbsXGEydEZl4QuAWrqhweOiFx2HBya+TaV8uQwnrjK/p2Jz3vNScMLUGZlvoZax
PuEKSkfVkthdzvwTNimiK9QigT3IIQdDLyZ093bAgQFRK/dMwlmG6b4rrMkiRczINS/oBGBIvoH6
HJjQ8q4AkNFbIO7xX9+fnr9DyvpNHBgepcbfi13sqBq0PRD46hy88NaZtBdNaMVMYeVXWbZNyEA3
4+9sWfsERu/Xn38mwwAv2KoBbU/06dHUuBuKUKaIOd19PIpSXKgepuns7X9QPaAsMCsElH1nnJB4
VGLmCEq+8GcP7P59QEmmyiBQ4V7WI09SjKsUvv02YfzLe/z7dABZnH70nk65euJCNde0P/nI9frV
qNR1kojunPWuMsmfURSGV2SZq6wbJ1xgc4h1EOH7Wv+7HnFDO7o0oD1+ZLTsf/3JFjqXMHLsgGqI
dlje78Z8RSYzRNYzAN0cSZhLnb6W2YcYlw+ZjPOx/RoQ6K6Wb13OC5dTcZQSCFRNG6iIPQn/hrBf
Won5CjuYMQ8hNZrY3Xe9OjtRlywkkpaIweq3A9ZUMHkofWB/Z0Aciuy4Gy9Ac8YHr4RvOyK6eFbb
Wf0TPtOzHsQ35z96KHY8j6Odok8tI8JhQtHNLtLXDS8H65AQuxS2F66Yj11GJeR+30x3dfcooRDS
k4oKXGarThuMIrkuYLppLO5sSVfPnBfWdGjlOE4cjFYwuPaJnOLj6ffVwWU9KwAb07vGaGjvxNMy
N9nheR4qgUqMot0XZ/V1PVDicJzWyTfmwmHW0ZjmaT97tOnPO7bAwe6SqRdiyaGtohEJzC8ZtCDu
3D0mBlZHL+iHz/4r8U7gld1piNjjdIEaTzIGOfyZD/6bzGR+Dsk4JVFA0iJBrYK0DrKPHX1t0r2r
mj1dJKCiDtxzlaComAchkE5uQ3aszXegw4DdRVRro7exBAQZ8mTYhIsDdHi+PuCzZNT/2BI5kDTF
mcK+8DC+JLUSBaTOut86uuawvF61zBF6FQo50kb/hj4GszJWUo7kOtyTQPDOcCf9gXK829bqB3EO
S4UkwFidgFmP/ZENaEbHjw6G28FfPmOqIOz2IU9YaDVnaN7/KuY99tZb/6CnJ3YrCXv1gnZN/6Dx
z2i+FRm4XIbDc0X/ZrU/uXvVopANmRJPZKJjNkt1Bgq1d1buD8AQOmR4iQRICwqTK10UMVDXykN5
KIb4P5ZscVu9NOfg7/rDxQIWG6jZg8uiZH9a+TZS9A9y/tFWapr28psmTq2RFhL7ZVaew/owLoMh
Ti4+HY6xQd4EWERC+ddAsVisVXcVNHsqPIYQD5QZP8A4UtfFyIfTbSTbNXA+Bicq8YlDr9bhJyvE
gzu9vxkdrGOKOKK5uV4aowEySl05P1+aejHkdXCjZk3MUqyVriXqcijQJISC3SV+0c0uAunl+O1D
GI7cXx04CEsQ0Ssagxf6nYbOIdbMskh8qzvKrk3U5nfmQe8WXD1tKpaGcI3ZauLvCOuDiCVVArGa
PlescLBACkMv+WYWPTDj0lphOLORwvCUHiYUgTBbYthMo1cB126MHBdy9yJf2FOb8n/dEfqDDpXc
MHyUMnv6N+4cpids4ryyRiYQrImxzNiPZtwRzq5iZO5RAsq+lkyk4hzL8ygWeXrEVOpheQvp1hCL
gIGK6Y3dy40wFSSohIMRltJnxTmR/9Xo2WI3ewYfN1E0kCn6Yh8r33SbaO+lc2CwU4tUCSdX57ym
10Rjmd5RNtu8GocIqBQzakDF2bGKqDx/r6SFvWyXwYK0VrC8Mbkopdz8gk88oQVq6nCXVlMhbz0a
K8b734WS10CzRWBcOx12m7ZEmsq2nxClKWEs/LxvHzTAorzScn/l9XmVov7ZI94qqtUM2HGXNEgq
0/VAzZBQKLJGYjN9zCfhx4REWu2Abqxcrd73qVK3kv3TvBu9/HldB/mw6SE//d1q3JqCJ6WVNCd1
dhBTI5sttDTEEN7oaK4aKxHm995AABMr5GFuzXnAefQ7G5WHCHK1O6D3iJrR6o3ug7VBcqM0hZFy
XqqwnOmKSYDS5qmVszQc0dltzYWUScZNisB3sNceWse5jJZ/wfRsI2nNfuN1Wwds2pDauz6CFtQr
fcg6zdCpDwWJxDeOzku5XSLjA+mZxJWRjvjerxr59rXLZ9SZcbfFcc7zxY1HBBZvtpr/nIXPLzO/
v93B6tfYbcI14/SOVOx9K8EEuOAb3RCu0gDSxoClxXNU9G0k+3LpCsPqLWv6Xlb5mHTxO/BukPjL
PyNqCqJN0XZZn/Hzqkz4AdA5N2e/brU+wzVYvBQ8Zm2jelQEsyZ+2lS3N4RrNS52Sw2rRZz2J3b8
BULY+GMsNRly/dzjG5vGOdxfaidZcdf9Mg6iFdipRUk8IydCYum74zKAsIA1yitYgYHI+KRznJut
l/2gVs3hpEk6kHdDz7a3IDqYyf6gAeOORttww0EdU5718O49RBiMywxVuostQwuTOAyW5rzaveWt
6W/PFOGFjJlQ7W1d++Qt+crlUee6DSxAgQCiu+K6E3wHtz7UumDJKW7BI0MpgHpWlhMGnGTQDN5g
vpKOtuEAoklN7rNbz6IrW7CAFj8TCYM1C4d9wpv5DuKmqDwTSJwns5PqBfv3uzD6lhe6weNvB4In
OBvUnn4GX4ZaqJG+KtuBEN9uBb2fIZ9AZOwhvBX3yDjwpp219976YepxnNgfqFXCC4JTy2e6S3ps
vj1c9+9GdHAPbR+sXbiaETIszrO8KHTDoFhEN0zjQ4KRMqmwrwkhntQMNT8apdXFv/rKaNxRRnul
vTFxLBoxeWoDtbrV5PQok+0a8OV/AF0LZtWvC4QcDJ3UxXVUGy9uZHThg8qAavIoCd/8OwSn1alY
NDKl65lj9Az06j2+Sw4YjFLt03gT+SFx9MRr0T9PkRVXg/zUBFfdnfAd7cG//s7hvi5g7z+GfG8m
rlqhY0maJ93oJJbRMZ5Dy/UOH2OCMl1yXWZwZDm3HQvQ+f9srhOFwHC0ppXy4UAm/036Enftc2zX
LamtMoge4sn2G1Ew1/qktjmE5x56SgGA1ZYJ82WUwYhHu4koClN/zi8ERtPi30qyqEpIOCM0w91j
h+e39w5ivM+ffmoLOaM//z/lXxMaLGcJx8a3TXg3yoeodWbPik4c8jAAAchlHydAj8Ab/EPaj9zO
a0lqqTE+w/odqKSB3NO4cTPwrg/pTk2oc8XoaVvwNw7kdhJoxSma5ODiEeZiRH9LSmhRHdK1ZcOE
7G1wVfViSQO2g8KcvIUdzfuULuvmW1V/Cfh7ynJ4xVs5ZYRtiixNoAATBhe+QKoIXUpUgHH9nPXU
3G3x/+RMdLb8YdloBbg7SmGsN+hiSDo9aNHkuiCrAZkIDp5ybiP8C5gGUflAbHq5X2h/p71husX/
gPyilddfwajstcNmxmM7ZA7CoopD3sB4ZjgrJ1thNzXSUPn7LJYAbprNCGJ0FOjEZbFuAaxZu0+b
Fx3P1FiAbjmwWwLLsjJFxgc+A4KRt2oaCKT9lnJLj/3DiZ1qDK7/wSo8t062GnOZQnLtYnTpf7DW
3do0nYuz7FoASKlTeAx5nFKCiBOPM5k+m0xe7C8rVD299uCQayThZU5EzI+2lIqE6VLBAofnXGxt
FT8imXnA5RXRH686C/o3ZfqLVUyQaybsjtM7UFInPjDJH2WBj/FCigdSd5+ctTlokFCw3fLGmy26
H11fdkowIKYoyHJ3Av7Hvlle5iRkgTbT7g9MzNYg7VGVWZez0ZykMRhUjow2sbVUN6WHBmXbD6u4
AmIYsXjI1C7ttg2ktAB/OFbTpyaFYK1X/j9g+/jZ7/16bQSqBykZC+qSybde+bH3g+vlpNj2BSfu
rIdTk0BQsBsPKl8/BW5VeseWKZ5WA7ADmZeLuD6de3G2ss7CiY/Y4Llb+9vVs39arVbpcSAROeEO
X7N7Kv820RZhC+gwy9GtUCfYvviHbORr31mWXGYVmeI6qSawCbzhviexY7GH9gfNL6H+cUTmM1X/
Oub5Ggz115jNJ3aA5suVLsenIUj9rBwnGkCXqmee878VngNgtxV3tGunIg7TQvu8moic4l5VtfUk
pQdsiNFW72LuHkfjplE7HXI2O9BH9gIbvf7FJznb3o6XecHIOFbWb7fxG/mVUEoaJ2ddmRCpU69o
MK6fIa6hjDhvyGhFss9ixWWcjrOFDel2TyRkCkFtGdV+5EJN2bmzHtDza7+sTH/PPdVjwSTTdpIP
R9hSPw9rbJoCRhNZ8bncOYeoyx+e2innk6EMDgR6htEzSRL1qdVJZmfYEYWvCfjtcOb2sWCeVBT7
1sAUmcgo4H++FbGJGAuW4UI2JEyAvLteHxRlJJmyxD3EVyu5dYGvWyGOo0lcwtbKdtl3kEioCi0a
yxz/6As0ag7HAFOiOtzKdBJMRVfSoxsH/RwGgskEPgo8pJKLvQ/VvgGnghZiZXsRU8bM8IouDktr
fUo0oOXV0FNASU+jyX4A9OJBqzwraCoG19irH85uYJQfFmMRfRQ/OyAhl5yl9fHZyzmzTGNWstX/
UOCmZKKb6QOQwtqGh8/dvAJ5CUi9xt9bAD/v+FMOvQc/NyaZA8c4tfl/MZfOz0RUfoA95mZDmc0s
e3aMChikkR6EnKyIqSjXoFYVgo8qUO7pauCif2gXidJXP2IRjBrExo1MPoW9VvEWhdivEi1pVyGi
3/UjWgkyvydnqywwk+jM9B/jES8ZTImB15o64e4aH0fT4kOI5gkMmDRxH5W+/vzfG4hLjezWfwtD
J81oaVI0GZvIr7K5kCDISFZMUTkmEi5Z7p60VZ6epzXcty5qyFfnO8ijHH/wpi6rHAwMeSNsDiDs
Txp/BZM6jLS5jnZ33HXEEzidKZRoPBIO4wfbIR+pa+2r41hD8fCYApBL2p4/JsIsuJzO19DPOAQb
2+uzhhVJQCkdyXlgSTwXzmrcbIoH21OInTVxEL3BPXmY/m28F7RD0ZDoJqaKua+yHFWBGOTrol/N
G/FuwtDgx5WxPM8Aaprld7qFDFDezczN+1n03r8RPgtK2ZcK4LK/xCrOV2PC4qBHyszHk43YakIC
u6k4pZrMsaK/ISNTrjjLEWljLh+FPcrlcUsxdJL48JImbHQga1wvbEGzehchd4+w7U/8ld7qbgXL
+4mDu2uQTXn7LZIA4HRmjT0AoWUNmcskDN+PDQ7qFL6cnIiAe7OAyUDjDKCGuZFqr63DYgJDWSRi
rmSpiZWCx9shFKdzSXohhyRAuuOvx0kiGFtyN+AG7RP172+V/iUes8GzyloQNt7m/OFF8YYt52F6
tuVYPpkcf8wJFsgihlkmX2pQ4H49J4z+s9ETzbOPTzHFI5zC2mMB29lohSGIsWjoxBgVpGUspSS3
s8ypiuc7vDxL71SjwRFXDsqfwn3CSYDd980nDd0b28mazNP23OGTF31/e6+QU2prhhTzGwettc2b
sIfiWVoRgCQDsI9qw/XHEGY9Ir6hIEU8Yia8epL1TH7S/O9xfDRmt6M8Oc2hwZDMn2t4HVY2IhOE
2AfoQ3FBXT6i55vP4HkUt9xfYUptkpWYuzKNhE5Hn4xJ1OxQ7Dh26PKo8IEhtQlLHT8l8MQ9M2ST
lQM6kQ25HRQZlyfYT6nGgIdM/sZEzd56RntQ3n2oaZLCU7ZiVe3iFwUrbPFNjHmLcjpIJNrXis/5
+Sbyz5jO3dCXxStdCxd0NWBMrUdFCoh5Yicyq+Av7l0pe58pHD58HfkLFVfcLZrSF0NoEqb7ILdM
1Iz2YlmvCOE2au0pCIieC4ir14RWmptxfJUQcm3moX6uwuOJnVjNZDGy07ZKFpAxXU2f8V82d1ih
s6aXeQt0BKmG9Nu9wBEl9YNoGpRKZ/JuwOGRerEt2EciUGvk/G5xgkhKkc0cstDBHjp2An0FV9tB
g4qh5pGJwD+WuDtZbOx8n58QhxSkeafkbh6WdR2qAdd2UEVO0iBk9fEvZMoajKfXUZO0fFb7U3in
jHDtZhRY4F8q7JPl8X3DmbtGCmjeP2hX1Kou6aZCTP0xGL8qfFeJ71WMORHzfBLW69b5xQ01iWqI
vi7pEAaaaqv9swISt2eP2vBH8Ev9C46vnC5nowT+S7YlHKE6R7REx6VE4LDyBF7N1HYNkOR8BauZ
SKsGV2YcPKjIZT9H7AaPC6AsAtYpb3UHdubVDwiyJeieQhJPtnEl4IuGcKsovL7bT9v/LrBCnbLY
PWRkHS/waaQ4UbdNHgNf4unwBwC/QXQXwQYK3OkpNCB8zoe7SM5lp1nGNDfLQoAmSc4C0UWLrgvF
QAn4Z1hdcORi4ugMnHs+WdOTKZtETzsW8ZwSXxdi+w/hlShDVli4a2yHeViVvZ/eSNCeDc9Z+HIe
q3FBVTVOeNWSmKr1fO68Oe58T7e5UGLDShVnneVlBRO3GHKTOkiqELzp2SZl/QQ+Cglw9tssMLDv
mRtl4xeOBTTLXE5k/QAL8jyKBR9b3osYknslSylYHZA19Q0HCkhUwuiwSgD3zQMVqtGeSa/hS7AV
Lx46zfVS5U3HXwYOcoJexNW9IIMjNlGSijONGqOKnjqTwPXnd2BGgaQwMdluOnra77Cvxil9PQZt
484SckfO5RVyt/T/aw36fUOD56vsZBdDzPyprVhWoMPG8D5DMJSXoJMp0Wt4arkepPteZOpfm513
ho3AA2+jwuhs4itmWBBS+QAlWhMQ+hZKz3mDqoZlOq2/9cCWQfzKNVnY0SMkNHN6f5ajYQ9LsXEr
xd/OYe7hSd9oU1eUz2083LrWQtBTtzAOgEge4Cpj9lUj/luOTvYtNJZcb+NyKav7miSBxHncVZUr
o5TuZ+v8w7p+0nLVAQRciRy1nQchfEXr+R3MDzXqrUHD+9EKsbCaqtU8Vmamd6hasGkKJKyuTseh
skLQy52N61WqlpDm8J+AHXfylaEBiH95ZvxNEftvX8vs9107W/sRYDLv1eviNUfbzsmZZgG2bBj6
WmxGmV/9R7fBjGxZpuh/D3QJNV6mkhn+ryiWlz5b1+4s+dpCNjwArxMIKwOJoDCJhYAV09eigWvy
t4PAkzJ0QhYHIVoH/0ajmwvUQeY78iIy4Yqqi6N0+a6SD7SVe3JAHjjrg34xqBSOSuYPyTG4XF1g
q1htTXeg3LVYRqqQyHYU1AItVZ54F+poL5oCU0JNGn017Xp8Ad7TcQMhQoiELSmeA3913y9gRi4X
xQ0X333pi4sLgv4Lxobpmst98fKvLtoq6a/omSgdxE8lWOCQ7FZShtiODAYebvyFwGv25Kd1Kwhq
KWm9zJzBCfVI1Vu4YTmck1okCNp8Ti0dTz9X4ZBSGNS+Y+9ZFDPz6AaDzZxnsy1vUqdVC3kV2AZA
sNPCnSzNEsNyApHhgfNt4L15BYqwVDnmM7ICveBq9spDDycpJ2mmJBRx8gCcsRbpoey1PJodE1Ys
BO7Yu897NqGJsMOzoUHBJArJv7bjTfs0Aewt/rs/N//h4CkDWA+Z+S9x0r7QZg8bkmD0tqW55hIe
XdenBnYDpMNf5vRDpRU19cW/W+ix+zpq9aQMgCnpBiQv5pOAs+kZhFlzHq7lcAAWXlVHo0x4jXCo
vobNa3F53bImSelLLtXzyh3kJmpVtqlGuQNQ21ObsflhC5cJJ3Wq9Fj4Or2SfTCF3Y6Q1441YwrA
91U87PDSr+vHHjwfvesekv7DmsNKHNjjAPpHVl+zvhn6oUYsL/L8J4LgtjXRwpIP0oag1Y8rSriU
38xZUPEHvi0qTDIatf8vE0/r9YqrFHatc3X2jBMif/SEBPO+mcAAhKrOjPn1kO4zAIAWt/FkxYWS
+LDWWkWgyDm2wTcFDogWqgUitA/qj6oiu6+AWCMR2v9H0vNM8VxX/m/50zEz03IYe9FehvlShp2F
5uuuICpOxYf01U8Z6tYEuzTGCVPvk7com3GDPNrfnc6Cr7s8j+87rc92HM4f9Czmu0zI2GQ7ZVn5
e2w/umf9pF5LNfX7xxYKyepvabMYk5eFyZXp5Vn9AE5eZhbO6L1xF/w07kZgnH8oD33PBvi5Ptm5
FN60Ip03awtr7Av9sLmcqZSYI3jHjbxRN2qQtas+gGdtNgzIyHLVSd50z/Uf9x74Bl7lMS5S4wq+
6TU/eFZXTZo6deyqhGDOtoCsDlF/wLpKUQIw8LjYL+zmZj4BvrQjZQ7bb2cfvNfDAM7NwCuutTYK
EWTbnu38Kseqywp0CkD0fq2FNemToVJbU6pGWG0piqQq/cQDUq7MwPVfW5v+bmrW0lpbgHnchEei
kEZ3n+XuA0H56TDwLCLO8EouJX2LAMgNQR68PakM9gEFinVMSlD20PwIn8M5iZ62DZMeB+1HsK8s
ZkXpv+LubNFCYyUEL3EVeGLmh2wDn0T4URwk/59YkNQokuMTdNoMoDcfkun+uSWgDx8zJa4XroR4
gIxURp2tVdul3/kERAqOlzE96ALH8xVkeOOUvgfUSzN0ka3yFK/RxK8dEQc0zDOhTPzC99Svh9nM
0xmezRtIFlxw0J4jJuuXGCiD9E3IsPf0GwwTAA+z1ZOuAm1M0/xBLetnLRGNmNooWi8LxtTLC2kO
NtkvfAvy+3MhzsrOdNq3B53gWgZZhgxjRjlQk2Z1eGzNPXriEJDc5FoxSjSBbZIs4Zc4bv2pB2LI
Qr08hnLK+/woNac92hDL1izCzqzC+crTbr5I0UeBmhDN2v1NyA3CmVZOj5xeW0ft7R6W4McQoRsx
WA4w22qlIcZikTJWt3VwCNy6GRzXtfxSBHEQl0uSNGXlgViwOBqyKCSiWM4mR65g8P8ao4geffSR
2TPkd5Ui1113+25OQ0ZJep2UmrRHZ/lYraRquO5W+IHIkV0C1KCjsuhJf+u/njGF0vOSy7CkEkqx
nup1KxoNOZTHYRBmjOfc3LCnA2KnJ2Bi8HDoUjkuz5VlMVl9CbgTDT5AXfx98Bhw25LpT3UFqEdz
q+HqeV7J1vDZIic84RVULeBjy2C0xpB/U5YGZvFJi3oLo6DZRGFik5JNO5ViU9lA4Sp8mxt561SI
KigPpyIEXsJ3BSLS3U2XoseBjFxBFQOL7IN7QFiLGLJWnJDLvCHXS91jIpt6odZwqnpZOl1ZTDU7
WBRnUMP1FFYUTM8xHA2EPBVAuumRvggqFRo3lr2PSGoLdL3LaTAjfL0w+petqisb/1wG0YDwv+xi
DlVVGiEhRkepwWYzWB9to4sDa7cXYxb4nNFVTsO7KnDnKw82HoesL7wgLCbbXGl1GK4prehIz19Q
6imtmw4sk7C0iNZJE5vOVFukBZvY+l6zXkqKQxLtyCi5VIFwIpPPhuSiUrtWkGL7XvfZ7uX4xJO9
H4Q23DfConyCOz6YJ8dEVJ7eS0e5eptCTEZPDnz5BU5PxHWjLz3lppGFopqxbB3K8FHrj15siUVJ
qEZU1i9/7YCgTQp0mdhTv31SqmC6FTapNKGsfc2X3LH+t6PuUgaB6M0/vo/4kHeRo72BX8WNI6ME
G4YY3lGJOYt6Ca9tkcIUE48rlh7WdheG/V3KB7B+/WmN2y9fEHkURBLevnSUrYI2P42qpCaa+VF+
DmmmfD+AtIfmcb+l8/eBvAn7otlDc8wp8kCoAtmJJUjpJ6rvbc9q6/HGy44fzYx8eESOmfmLcUYV
TgflkJJHNl/8ddLP1lfAr0T7JE56AxUwWRl+EmEh4miEokIWJq4Xvu6DQ8zOIe7AdAkSUOUJuxVq
ArBgY7EJAIAErBkAkXvpRGN+o8aZ0lpg4oYp4RIDQvPBA3tzieoerW2EqBALbWotGEs4D9/R29xd
UniHl2oSYkK2HwlfRA34qCQOtepd5vGmtulbhsYTl+aukaz4m16BZQIqZdTL2IUZPLncjfla/Quw
jW8mLRbvBNAbzZsO3T9P0liKREdLj9pF3Fhx73qjfIaVpB9A+scYGpbUYPDnoENcuo8O8u8j95t5
14ZUo7IpJ05XdX81hqZpqI6xJ+8U6aw6ilNPhtCbKhjD9Q0ug/W4pNHW7EBvu969XixWtLZYu/gp
CGjaDqX1TVSBaLpWiS/PPV4l64sQw1CauOyvpr2R6Y69GI+FPg36F8cMIdL7VK3v5Adr7SCVdHYP
a22sdwCct+P+E12fRjfT1UeIR1MuRKKgDVTClZNAMFSjX8lyqPC4K8C2r6RaArtEqbYnApw7jWtq
zBTXNe/s7eDBoRx/PE3KzXkz6tmfFe+PHTGtiJLEADnDCWBg8td0a4/+Q/7LuT1rU5kT3puSRkwr
8N9vZ5CvmOhoxVNmM5qjemH9G7Ms0ve2iVIrDE+VHLVRyZfDrp1wHnJ1NKPaixaWcagcoXEFMdh0
RDWMpLJ6OazwTbTbr3B5xoHO2f3loUp8Jp737WqPINmBMzMxO831xWKbDhl+uLn1yxpyo2fVMMOC
HwctG7FgUixVNraqvTdwjqeOSIIZmZ6XNZG0EVByCBc8zw+oRthhBPlOfkbtDwUGrY13hizz+wRw
4tx3X07sZ76UGLezDN/hXQqsW1hyPU9aifza4OcljVCjS0Mffvwfm5OPUOeVPZIV2UqxqBaYem3l
CPnOBwhASC0qv7grNaban0B+VqyCzJ72lkXF+aswsszz9SNZzBB59IUMUEZupbu0nn9TOUXIWQoV
uJdAyRAAY62FYbDTLF33n94jKL76X4/gJquxTIPgDQYRH9m2ZYXVFozCSHYpFgMUvT1xSQmfiCtG
AYtu5DG/MqtjvnBsiWOTXmK/eRNxvKYdEY4gDivngQzwFUhN1505doyXYiEESfotkwTkA1znOPzG
4XhYW5X150GEp33VTb9z6TZJXldRlevYyNLi+Z5cYFIwWgQV7DmAFxrz/dzR3iOOV3YuEbd6lSSp
M7X55nszV24f02vI21Jt8tn42G1TrJYPayluWnn/u8Jkd1KcpN9id15YvzgwRXEF38+qCQXmdNzq
0YTb9jg3QQ58RKhMTWNee+hp2EWfiklejria91TurK8vC89tLlNpYwVd4LXkgdl7JfgTpb0JXWxz
nQe4RbRdtaF8cFNvlPVfEZMcjcYhbpRQWYbdsan5olroYfyje5PjjRuKk1pZj8q0ZyhoedV3kuzI
riHLWyroaDgSX2qtebeVEhWWlat9AXD36EOXtPH95Um3Mbkc6i8JggwjBwhmClsKDns8pfx04oJE
YRJHuxKV1aOUC5dCF9w87xf5K/g6Hg+IzTGTkKhErprTEkUsSnHqRawAYn4rzVZSu78bD3vNpbyf
PWvButkXhgp95iZXMfZK7YbZYISN3X1H3HYTH9GSMXGWBCm+ctrhv6PCfnsgk6yIRInitJ1lKs4R
7Xenk3E4J6cIzKS916gU4cbk7ROJcmYul2heLEwsGvaY3TTA+duWquGxgPq8CBN1JtFDluk6eb2+
QiUYJAB3Zv1yZtRhhU9mLjCFcl+xzOx5Sg9AbCu2vxmfc7h2EQLF2FPayTLCQXfOUJeWifnKqkA2
pYHWMvhSD7YAlxN7DeHboQz7POj63enKQUa8fvcVqjea8X5YHooLuJyz8E6cCp08JCjJd/Gqlpkg
ZrpivPn7uMDEmQTWqsNV4+8xLbGdAu7fDLIZKLIe/URybbJmYzOcRk79afkanapBqYWoR3u0ERvq
NOU0urR/X5QZ8wwUr+wIOKTNu+90Sg8HNEtpLWb/nvIw6ZJ3b1t/qcotzq/3pWJqjqeycYBh0ZOy
vezMAJ4e9TihqcYZUTH98B2l56SXe7WJ737Vjl0mfjii2vuYdTCtkVw91ywJpKqh1+Maqy8GTEw5
5XiQg33aI4KQzqIwAqhOoO4cjFa8l5irmmxy39oYGSlryC8IvPQLQPNgqA3XZQiquPAlpcUBkGQs
X9IIKsfl1d+rrFR/UfAIwQxXV++x3oNccBu7XBnOd878YSGczCku9UQIKOnnuVwwx9jADogL4oeb
jzezuaKa+BouDa6WUQoYequXez/ThUzSkSa7wAzdC8hIMamoO74UkDdrn6hUZzAuIzJKFAO+M8MK
nI6AMNCkOCOWAguq3t1coTQIfGzUVClT9fxGhuUfbUHXAcQCgZiB4Zw3II5MPyLx7Ro3u0LE9TF2
5iPu9fq0eSWw2cxnnaQkvTfd7zfomQxJn/gkr3G08NHVgy4QNvSk3dBpIIEv+tk9U8sMStkZiP8Z
LMYqM5KrMwHC54crbIr1KwUqTyhn9atSRoQxj6xeSR+GDQcknr9Lm3CMcouKS+1kg23N6FE1hDj5
50WgAgxPZtRfQ+EXW29YLkBeil2tX7/6agZURw+r4tWRNHowimICNkLHeA8tmu2OSR/fDo5tT1+k
QQNJY0WmLPTwaqeXOuNDWyMHqzeRAlwUreqtjOvfToVW++IiyZNd4GSpLtp+TX4AY70B0+iYho4/
LJznWvNf1O4QNyd8xBUDJe99u5tRU6/v3hTEKwAcZmnt4hD9gkE2do/kkW42U5LGWXaCAk69hPEl
9lbr+tfbqhKC8i2cT7bUd/Wxlw4z+OcnPrK/tnxEHF0LUx7v5GOz2/wRZRgYdOPO2wKxZbgSh2YL
P/xgyEym0AUQpX4Wom3ZX9bhk+ErkbGlWmFcHv6zuOsUt4xXCoViLZPEdbGpMbrJlXoW01RCp3Ko
7YiyTx0MGVZZFvAqQiJEJ6q+vuUXOvQdT4JOTupZRX+cyiEfUhjzsMOuzDaF/7PKU7GS8c9jUHJG
+H1PIcK3ZGn0BzSqrX16tZk8lCXza+QcuU6b0NjRdTZjB2zqyS/rRDQG401yS2kcWqIA/dda9h2Y
hjmH7M5VkoAWaSgBMJsmdJ/royMc4qrF/Ygft4EuCCMwRJIm4HL+MDB/C90RIq2oYmIGR2+EJdCb
0XvXJjDYDlX94wyMhLgcyWHlDINDbwVHzvhAiCfY056OFiYLEV8ezDHxKujL0kiayPaotNr1nerY
GthXNhHPUssjkzaL1Zj+yyPqXqCW1CNFpfoOvasSqvHeQ1UxoNDGKJqJCrJO2bpPd8vO6mt4kUgu
cLJAb1sJcnytkpGv1GYIW++7iImGN0OYuqe1f6xmVcttfCZDBFK0V1QR9BRbQMl6j34xQIwvDatN
Q+fdDCdPw06/Wbq9rqw2tNqRebJVVsbUmaon5KJESRog3X/ZrgocKo3vgHC6ZnVbx0Xch/rq8xMP
0g8DQJy/8flv5QrQY2kzKbJIqQOk4eazQw2Y7bEbA9YdL2lXFeah1Z+LXQ60ZrD4SuIeJ3x/OZXI
kOlOcI4vodKYGUlJrT1NPuvg6B4amYwFHCHPbHBE9ddacB5YWW+5f1IbKpOAohzb0QRx1VpJiNcm
CqZcSC/SMqrPVns8OUzPhs7miJPmbZ7olvpJKmOk6/AWcS+QRhmRu4rvZ4s7BuMtzAkTHnhFgnoG
6tp8r3o2Qgl6LYIFh9s7STnlxSgDeG/J2vmOUxJuM6B+O+dTSDSvO6d2IXgJxqFsyeD45RwJkynZ
9SnJOykHIHy6HQrrVWic05fVRso91F3Ur+pgYxkX/lnvcmlVZtfBCzdYkaQky6LFosDKVDqsNAuM
ifYgHjAVYcaOqETdrGfwq7dRt7iKZQCRbSz3dZ7zp9RmyG1w+5C2414hYm4NSWNTQrqJr5gcOtWI
vIMxwZva9aT1uSKs1rCcwKt1hGCiEo18KDrJBv8QmEbWAuCfP1aUkUrSvES5XMAMwkD8Sws5dAfj
tb+6IVj6iSnT6oeb1dD5Xoc7+5kw0C56G7etcZSG5SQApNAd8DLjkvXgDIHI07/ztC31dGP+Zo1P
58khSYhkVN+9y4Q7i/PTa6twtmduDBoiuQQq9s/Sc6/iZr7xRgR2JjpciXwU0W07n5pVtgNS0Pa+
nXkFkvvRsL1JtE4hDu3dK3X+BY8iWm+y7cSiogfSimPKppo+Hrv5T4T6EkeUZGef6/n/lFuqeLRy
/neGIClRwLvxmIMhyl6eNHzdGOWortQv+fiB5gmiSZ1iu/L1ld+Sl3llr9kieSEHtn6NE+5CPNrk
2YxxUPTiSlnTzLMgTxcDMY7j9Bsc77wqpPL7hLaX+3ZSAzr+uQHsYjSe+B4pStOWwiVFsghenMsw
nduOp/Mu9tT0XKssBhtoCZosIXvSnorMqMKOSrAu9+vkB/s6NE4fCzVV9kr+eNmXo1YjA2RglyeI
rPgZrabxAOuopeDtkHMkcBqwObhK7b5G2I+mC1bvR3X+ANddNfDyMfVUb39VruSFnQ5Hy/Y/want
o8YUkN4E8p3lW5pkMvG1MPlA1IfoCxYE8oWCR3uj6eOp4IWLXE9xU5mCE9SZbDUrxtYbPkdxrvNG
bp85zX4DoEoQ6W1at+/tVbsvmIExcu2QcEBzfBnFfmE01iE7AtS8zDWfKxON+QmYj1stcQnqLnGX
NoJVrpgXbAy6jLHdHYINTIO7FoW22sVtz39/Yw7F3g/J2MDb7cJaWGbelgKZ5tDcSPMDc2rke9JS
JqzHfE303phVi+6mQmZJEV3p+Bn962Tt/Nm1gWaFE+TwEatYUSSn5rh0g4Vrx8MwK8O+zC4LMS3T
isw4kjZBuO/Ou88YnhiDU3FrPdxYlFpFTRwSqMzxzn5lBpJx9JLr+E5RvKKWbS6WWmn4/OM0MfLL
laTI1wzEDbx5eBf3O9x597+GGgURzKcPqQIy6ch5t63RsyJdWA/l7JB2pjpWwR7gpkKKJCSHaGWE
FAtiCL0SPMqs48iCo30PDBW1n64lztyDoJ7jAf5CGafQJXzNctKGO/1iG9e/l+eNutkWJ1q1uIF4
UFJkMK77nqkjZHMm9qBMdHYQlmnGNqqMwNtJafkfMVDIVqWMp1YKX7zcxr8OprTfXuqW4g9MiMR4
VWNZLhV1W4aK44QL8q3B6q+w+UXP6acn5AUHNfGa9W4X2oMC+AfaqrU6fqIGBxhp7ui512o9/Lua
5D0nuw0QaZ0ujOh8ozzDpQ1H6lxDMGQv2rOq1q/CE7QKW35PFzU83TukkqHZ+8l7oGUOUTbt1qpv
3QzSomyo8HqVNeneqId4EJilQgDiUoSH7E6hiQQi3Pc4pSZc9ST7fIseVJ6JxaOSdO3JpBGglJhU
m6dXP+6INt8BGBZ7bb52sutPjFU1pHC5ZC/eQ/134/4r/neFLtYV+Ra5DP0UrfEJAEI/7D9mtd0g
qvaiUJgLbk/vKU6EcwEWUSwdFB9x+u+Vb9KXCEJU1t9vSSmgxz2yZfsT4itJ0gCXKdxT0IYTZDNL
2a+aV3C7rNM+mJtkcmlgR2F8tojPpuedCTw+1a+5WLgzsjG8m0GEI6Uh4b2zhyNoknxOPVREhYxS
r0eNPaI0NVyVx6oX0zaheNVoydWe+5szF+iBpCohhLWjyq4ibNJPFxRHjWa5/p7qiQGUFcFrJXR+
gtilPf1Uh2iVfmf8Ig0QYhJaVTsUZDRwPI14/46QwM/nevm5zi3kYRJtXUIgc5+MlQfeWiMXJOsy
RmyvRjxqw+wcn+OJuWD1tCNyqCvKbykIHLkz2efu/QGxVXuULWyAu5WkvaOByhAif3OD5sRLdOOd
Jf3B4nBhLrB3cc4812pP+q9TG/QJJCLgAPcs67ztscno6gObz2e7Z83zqO42k/3mGzquu01x2NJk
jLCZyTYv6yWq0aeDV1WMnDdm+w86d1juYhra4gkwUkwu3952C4afl0BERWhdEPBVwQo3yB1zLMDB
fw0X2szzAY4O28xLY1ChsO8SBXNLWOtHWa2Jvi0sWmcTd2xs4lBjrmRKuPMveZNc5rgz9pC0et55
XdjjZrjINDhz7orj1mDL9LZ0AcIqlRIKm5Y5S0lUHZK0tAfvRMd+tUvuke4JTeV4t4B2RciItqTw
eppJsLkgD2YtMpPpll0aY10bMOJcESZcNX0uJREqOKkjDzP0wK2E7cZjBD4qEjjoGhs+/itSRiFr
DqtAcdYQtcunD0p5dF0qLVCyQqEpJHMNB/hiH0i5BuwOaiJnggxIbTn501Ctublp5O2kQbCqb7Gv
qdV/imXhrEWGBHtaIR6lfXSBBRAymYccjpUEmjVkubpIvW9McyEoiFhHIw4QfQsxWU7C2P76VDK/
c2Ip9xrXlmVLoxQIORNW21pHLYm9rPGnswPEuBnVXigi4cHiJo3RwuEtVudHzo8bD82AQx2ai7wA
dMFht8k10dHM8ZaIXTexTOfMYLrYskGD3UNHcbBkzvpiWXOvOvE4z0f1QoyTaQ5cqfMsje5GrUH2
IncIQVezAu75QUsTm7rvc0gAgJn7d+XuHzMciuagNZyxrPiQWSBhP60mTeH+HUCeEcqxa8KEqpLo
utiiXRt4sD7VxM9WadkvykSVCrP2HdP+WbXPFxFvR0E3B/pB9u7JRbWlS6suB3HfoNesLfr3tTr9
14bg1XxTtcRLE4ROmgfxuXidJirR/ejDKa5u077ruO8o3b3gZWK9qR4BXYN5k2eaq75DDLbqNalM
MTd2fYj2xCQjqf2H+OQgABxeJLhWgwrh+KOdG1r00WkivTvQucxl9eNvxlWqrjRwIcclH8hblwCX
9KSRTtFRNdYtBXX1npnvOjjOEYFbjWcDjafKarwKb+rvHMw1g0fMA8zsU2mN5JZWhGUDuStOiY/4
O9HXZEDuoJVZgnI9Wu2JDSXyYK6ugCaAmDJIVZA/66sq4qQWeXIzNUCFiiBAx4KBuse+3Pm/vqwv
rjrNmNmnmxoRjkWQB5X97LtTnYWnqgf/OqUrqxlubBbZaU+XLDnp5Q/weHeffXR8RTGAWZTU+PZl
VEq776zk3NyU0sZcc4e+rUJacwCt8qpkIuOgTgj8kHOIHT9+VScetY8UpL04oZI3xTnlDZjnGayZ
fM2MWsbCoJIoXBF7c5q+S/Ym/H1nVZ1v7sPj7brezQL/ETj8K1VfUBvZxGyAjaXdJ7fqg4mrrf0Z
qMIhZ8tv4Ba7FA5Zvz216HAaUDnxOmDM+HT/XjnxdmMYX+cB5/VngXEPjSl+f3OZwh7FOkWeEcTx
bBqchJ9h0q3Qdw3lU1MYWYMv2rGUrUcgT47aQ96QBZ1IgUqqrOAO54/8bK44F7/69Co29+z4S1Be
Wc+8kONRQ4hZ6PeRgCEJvMbuBT5N9NJ0n9aMA+R9mnQg8tg8vkXZZ3Bwebdg2Nw+4va59NLDzoNd
hFMGTgnQRX70M1KkMkvkImUtzVZZ5elQUaTMWowUHI0OSG8jjG85mu75AnjdxsonrIeZi6QSY2CL
+HnNWx/I5qgVKkQqDE6hh/87GMUmYZxwXyYzqe/uwJahAPNuhyZNHu78Xokdb2S8gyd6aBpes5fU
+FHIBf0KNIwjAW7BvdWr+l+rG956eriNJXrHGEUIigwD3pLkrV9hNfPq25L7F6mbfYNPr1hVVf3Y
ug3LlfHrzatIC5Q0ibhw6otXa2dgQIscaB7PJlOmx5OuH0MfW0Ixv/huLJsLG3ZOnN7sO/19WL68
VkKLo1yORgqUFSrfS8taCQn89BFP0AZEcdSQD0Dnc9BusPSLeW+qZHOmRP5JNc1NecRS/jrRVG9h
03v+jgbY1dXhhnVv/u2jrQ15lEACjiio0pY+QxHtVSC3KEoHZw7e/fgPC7AmlcHb6hX9bb3ws3QI
ElpXofjwSBU+qI54krjBjQ2emmodfRWRyj7IoNWD9jmAhdhLDtx4eQdxuQf4jrMciEc3AIKsRSjE
nkBgM4qVLOepAKR+HX+ygvGu/7jvCDNLkVDm9Rj1PgVtCHg5rkkRacnjzKilHd+nK1yvQRXBEpYy
ny4D9Ap2S9BE/tVkHXIufCfCzyuPwaJubDwNNsHO+cEt6dfGYR7QgV3/bVABrqQzNghUGFG76S60
0yf6IQQVIJSiHUgbP9I94lCH/Y56e6JolchUvpLjQvjOJzYtVBNTaZeWyeLTDLTrML4wRzNZBsf8
7738HQbZH3sE+wqvptZud7SBAXFWwtRSovV8sMj+0wLG0xetzRpWXmXVpy/JVKG4PR2mgPQN8FME
fffhlvIB84yIz/wn193+p3RaatTdec5E1nRQ60kCtoh46f3sucp9xeTovLupsdXvCRIw8VmZF+Zp
O4BHMwtwmxK9eJaw0wP3cHbwyYI6KvFacqolW/U1gSsskaa6ArON+qPq+dXbzf1VsviYo0XphhpK
fQvyJ/HX7SntXKUWkKwCTvIoXWvOSA19bTSvi5iDRkLbRLywJVwwBopLAcY5pcBItYncA1benkKu
uQ2I1rw+F5eGHPUs8m4WD+hkO77QD05lspdrvRlajyqm693ZkSY+Sx92cBFYXWzCFLtXT07y/0PI
0h/lPYp7bg+lw1swFWXRcOTTT6QujEZPWvbWphfXAD5BEpKGMp0wKwB7Wq3cRJaVHgBy4nlbe7d5
u0Q/dG8WrAbKjkhJlkIYBZVbFjthxGs5zSWWZ1e/6fCMuTAVFOresQTWdrKOTK6+SrljHvGBa4v5
1CUaRYJWjnDk1Mz1JNwXyeUipchSaJCYvRioHQsWHT/zG02P7MHxZjCboL1f5iCoUdLcHAXpQyJn
MQRSx5g67c4WM26sZHNwOxqkX8zot4ds65oFPlaM2XIKFswTAgfF1PYwvCr1l5dQsZi6x6YntL1R
RiydAgDJ3gXsTPt2vfhplTwcKqzCNOKPFg9yh3ZjsEH6q67K2nWJQ5yugRsv6jcMQaM0yFqwYH/5
CTwmSxpmbHIDI5n1+L+6p3tMrKwhFlBIax0klCcy7lf1KmmhJOKJ5g85Jw7eEFZvQB4y7+eJ5mJr
jisKFz6pEKK8RbOj2+NnSie3TnaC4+y9enCJCVLXFufpCNCFkNJWacXdxBFZzhFoP4giPp+2a5Jt
K2HdJ7GgN/BxEGbQ3T4pUutWJbTgDsQlwp+V8xXzUQKtxBd9+VTbdQNrA7Q+tMtTna4LQqTxn1IH
7WaycEQBmotE03yht2ry1SLwbzDOicPVZJX/7d/fm43xNdOo4+NCFcGEkgpY8u1mNaF+e8G110sG
wM9dLv+DjcujCBkfOvTiy7mBrqCDQ1tLMt5dqOYkWEhTu1lSfvgu/uP2CLXw2xcDhjG8e9SbvAO/
FlgCEfypBmgxaI+yxfvRWIRzDmWk5pcCFr7zKT9Li0sowLOPVbsBYkcqDvAKzPtL8qJYN+PN5LhS
MwYsqS2Zgu14DBAtbshQcYpdN2dzQuPkOlQfXe1fOMcj7liyuESE8g/ZilZDm379b/grsUfp8cBV
3flhgoxIhrNW+XhVLY/8zkIiTu0hhiidGyMFAkNJAwezJ1zx56E5qaqvg716Q44Pc+y2/LHv83bQ
9ZvnQzp8XSxtzMXECIpRzcE8IRQPFeJkfsXyHycl+yTWGUpLi2rSCAs/fHbiWlmRWBYlpPNw+VCJ
AH4cKX0bo2Uncuy/vPn2f5u27n+XFqBxr6tl6TJjxRKmS671kAhVVM/SAXYnnIkUvO+7TjEFNFXf
zOyOqvDZ1HGUAr7nfpiw5ccvxMY7Fp4pDgAZk3grorpESsv6tKPF8/7gYES9tcnV9CFeilrbKYOc
GV5dWSfQmNHFhP9t+PVezx9Zw3tkaJQt/kFAaDS0oNTkVkNWLCusupCPLMXAJA6ZRxo4d3mrjmWd
C3thmPZLPrY+baR8so+7GTIcrabxZsB9tt1JMHyRi9zbxdK/dTyJukLEO3r5Q8pJV+tcEH+1macX
q69OVGttJzjxsulH7KZd6cAE3u0VXUfPFHMt3Pu4w2V+ouCgRFWx6mi8G/g1CwaYM6/1pVn8Pbqp
iotCTD0Isfy6w/5QEK2yxgZAtkoBErgtlMMCFzKx/YQsdge3bTnUwbRg1c05AAUgGkXFlFbJo6A4
+PBRyg7ij9dh08Ih9GP11VRBFrd8DK+bJE3EY5tbkG94dqE5yiBN07I6T9zB7HRg8X0/ru94MPTy
MlvQhAeWd1spCfGRQrIkwE0XTQx+i71cJDPPQOZ3UxLuVWHRxuy1tlE9fVL+3DmIH8TwoH0lSx3a
LAmarlJaKYmWs7ESIk7sqKhE0dArZbf6X8UK9G4HZ1E7XODAHaHeCtKmV3OfMFrYYJn/s7UEDTz9
qsybL9qJywMQmRIabZ0UPHgBCQEOHtVhm/Kas6VZNH2hObRL3MMPTd0Y4i5JpihCddri1O3EiHnc
s0PHjE5jD7V0glen3O/JqcyLCWtpo3Eq5Z42TqM7ynBT4jKK9wxDxNju336rkuesm3cHukJ5dwz9
Gf2sRSZf9DnXAaBsUGKUAc9krAAi2BWtnl3/Ksw+5a4j4aG9xasOvOEaOpymFVH3eZ/w3Qgu8vBU
XDcuxXEyhcV4TnexpAA35coBFyivNdmUiry9PRkcZKOhT+82heuDp+f79wk7rxm4ESXF0dPXk3fb
PReNlw6TTP5sVUnR5RGhvo2LTCcqYKpFTFJGElVJ/oB/9fRQ+SIDg16mqTwVc07+gKsMSxgWAxHm
SUzyBlJs/jA1bFn3nPc8VE9W87hSy4DEsE5YVr4RBv8qOMny4LHKzldQaghHD06xcpZ+kquAg1gj
cclROWmWq7yo4+8hCUyiuTQiaxEp0rZPfrgnjgRW7f+tFGf3yNdeM9MieiHkqfLdfGg5UEAyqOLJ
0/As5DKydwlQxVf4z0Xuc2TXw/QCDsaYw+TxzFRL/GlmI0VclNLRUMQqU2GThuGRcizZLRJI4WR0
KWxgj5JsNflQ6z6v7dGzZHXKHHa4VCXswx6X4ILhJu99o+eHeFnt8C2YfomV4zY3rdW01wcUWBCt
VdgPmSf7mO83fqPGZgIv+cPmyVawU0SgOlgRTHb4I/Ou9rqIRJ0VrVUsUlYxgPDZxoZ6AeDhpZJ4
Xv5+KCZMlkd/iVMpBIk8jtgexm6jAoHcF0z84F0WO1ttYxdAKwmWIpHWYvcwIKwMj7GCckZl+lRs
DW8HAgRMY0RfsQQWIu++YAgaqQ7co8N2rzda8C0W8PAa/dVEbHCy82a70l3iQ8GX+goX9Bcj/Tc3
dvtowsSVYJzAnPrOI8zzgX3JAIejsifnJWLKjtiL3mMQJpvBz7wIU0HfEyVPofgLwVrUIfFYqTlo
lM4B7GqWhqFNRrEIh/zThtJ6XVn+RmlfF9T2DpKxbXu+lMhlXN2g1fnOAum5hbeQELJ4dTaJtESr
HhBLAu0rC6quTCOF/X1wC35a9y6xfTsP4RPai7UqFDtsMSlxj7HXxMajhdqYuhqwN4xYr6Veil8P
8m1RY6PzR//99ANIzAqcwqjm0z1FAoxGzB3TXxNyr+2BUuRsRfNSm68zNIhm08pm1NxXp0oL0UMv
GS1BkKJMC9LDRVfpV+Fb0zKAQFYtUG+oV9Cr7i27YS0QqGvtvosGHUiTVZNANdzhlLuf+qFWN+x5
7gH1v7Vw/9/H2aJlb9jCKQApfoydWbZcO/MTM1LU55NiQ+HGeTeqyU6yATPAQB8vD2ZLvOhlQUuA
3QLGVsXvWKFvzQ+D5AprYU6kUUyVY5czBkNG6UBN7oRYksctgFDqeX2a4reZBVouJ0dLHbHg9LB2
md+eebki3+6fQYgAHif4XmdG+qf4abvtslGfzWSv1SweDvBz5mwCStrymXwOvEjPqS4EOiSRM/IY
vnfGouWHWxn3yliQ5taX71FTXKuLdO8bbgI5xOpxs1bgU8nxEcjYfRy55lBQnx4DGeYjWaNQVzh7
ElWOQxtQU91lv4IKJe3JJ3KJ2baXcELOZvcVh4r27Ed3OZ+m+71CHzphdZgpvSTmqZsDBdi2AY1N
GCucduL/Ky3QOkhgmoPktgsAlmMO52hcuUwMy71zX0l2a7PcK0bH/z6TcSARySyQs0kYDgEMqQHi
12+cBnkOTzAYt+uhBMQZM8PhECk1sfT5p5KgIXGjY4EV8b7RvOSMZMhz7JNk5Dbm2ovzT3mfaNxB
YDi+da5sM90QP/GT0PV0YHTLh98m6h0PRghLBKZvzSYnjPjrlJ8mSkwDgzKiKeKRODmHotBs82xh
WMCMCOh8o1DQHDNKqEFRL2SbJPN0S9YH//+MxzjlSdJhIdkQ8AZsoRxrD3iERMJ63I00188z5JWO
sUZ8R9NQo/oFnHctMm1I4RYhqDDrY0U/4//k37by2zPhsD0mnSFTrRICJJTZt1iHkEK3fJlcLJh/
TrBsyc2Vh/wwcttn5mONTpVpABK/HQCqrL2rDX2tMfv5RQ0j/GV25cDMynQyq85BYLJWswBxoiVi
lVjsIv6GUnWcxxszHOGma1kRVrKJUIpxd+E6OKKORsMev5eBnaALs+U10kpJCsqScm/qEH6oIvp5
FMiGhUfvZxgQ9JNbz6zE9IqWREMtNS4ZZ/iOvEvRN5dQHSPxAJrIhSNJki6Z6DlKfsCVCC2gtObC
M7wb5RArwAzu1jC6ZW972l/CVeNoMZ1k5KvJsb8BHpd0o4/wFyN+M9YrWWpf6h5LBlh2mAnYMKrg
tEOZcln1xO5JZx5eOnnwHEYLp6L0XbyC5vWrq2p7TO20VKyNSAeXZadbj5vpWn7ZIiSTujSHA9BK
d3CidHeAE843fxcYaVlwkfoWOvnqv6bC1Dflttp4HUAyW9nYn1A74/nA045uKHe/9C4UQi04rhYq
NGHAHnPKVu1ha/KdtJT1NtBAp6dUcxOyrbKsrZLCxXsCYIP7UI4nS1cNj88N2e33bXiuc44iOXyJ
gQIpSbDNaGeHOfN6YM2wOvP06at60+WTfllWCv56rq3fmuIGOQKOZGZtKpnun9H53d28P23INtNk
wU/PskCrPHp9RjEm0UYvJ9YNvkA84UJq7lnvf1xSB99qOrbstEayoISuBHPBlG1B3LB8M4y3FhsZ
yzaIDV5AJ71boDei1Yy/D1y0RLr0RTlEMEGLzNxSeuDaHWuBs3OX5AXwVXYSYxjymXPSeII0jRTY
/SaMmun+TZcN/cAQO549zDHTIm+uLNMj5tUC4OcOyNVS4ZadvV6ePOFItoGcJPCDjJN6glJIczqw
zoF4d+zntdpZfnwyzg6PxeSha/MpuqIt1XFBNzCpvKdFy2FAzF56KzhIp+Y3Pf3PflriBIDLnyJT
1CRD4r+zPjzI4r51edmD3rIKpVL8KZ81YW0yW17L3gw/6bVBvboOGccwKU7192q1lN1VoC1LLlOJ
2AUt3ToWfC/uXwnobEpYmLciyy1ODOcGqvIII0X6bru7uHXthZF9KGH1mxUbAlXsI6T/2UBl1gXC
ZXqwfT5nbiB1ZpjiJo3jXMbyE5vH+/6/yA8oV4FY7dmZrXAjdG3I/Cerv8QNf7Jul2pLFbsV1YX8
p91PaTeB7bwlCXICqbPhD5LxSapiAvUrkW4sXeXa3ywuK1dSLV19YsN6RpkLd1dS91AEKh03niyc
l0/h6rqlfD8FyyQaDd6/Y1srl54bb/lpK5UaXehTH0HwIHVs38poVBkOIhQmc+R3oeBh6jLIASpx
kdcXRC4Hkf6NfA64fht49/6qzZzBG/lnepTCaCyEeSnINl5CM+umVayxInVpYb6jQTtTPwGQbuUD
7SEyT5QCdWxQiAhK8YXxESnLzE45z4NyxmPpXciR2edKsO3q2yoX2WQ4NxtvxamYyFkUXU8Mjkhu
rPlHl3zZMkf6t36VeRlr8woXw/G/jgecsODFIZrKXs+txFO8ZHddtTG1UehuOSqad9NijK311R1u
nVi4qd3UDL7o0JYl93e1JMyzHs0Yyn10JkWIRX3hO+Z3j+U9G8pmYfTSgTaoBGJwsOtOrcNrMrUZ
WmGWbzUcJlHGAgHZomQRRb5Q4gI/c4RstOtYzbJ4UQyHg5JByIWGkB1FW0jDu/VU2J1qhOtj7CmG
xGPJjYSPy1nOCM19nC/+4jxgckzxrF82aS263GsLh9k8yWCCm70PtrAmN4+dU+5XhjN0tDQlfnMt
P2veZc2cX8q3fFjpGd+Fp1X4uHRH0y/1J7sL88LHOwr8BEyMMoEW2LnyeF6jOB0A9IVjlx0oVC8W
C+77EVGHMS6I/VDbelDij1kz85Cm9+JnIeax4vwbzf/O+W4b7liq0cLUkrCOz94KevbYrpJSJ0Qy
rOgNLTGGaDrOClHYy0KwvES70c/Lh56Ug0erGuVsDMSgTgVse2HVYF4J2IKDUQA/MJ7Y5pv1NLvW
wleken/Bjr5B8xm5RRtapkScQqDx3wFb+LAtDG0Q0Of9Adkh6ShFgyYhEJmXSmj0fgpinB3J3h76
cC10WzxaI8tvDYsWSj2QnGnVhwgPHss7wmxbtzUKQ6wDC04Dn4HLqXW9wPhQjf3ro0TZqr8XW0n+
9cf2M2cdHXsxOSPytLZWHMXCLDChgM05tAJJLgolIHxE5D8Agq+f4i64TXbYbdPOLuUhfBc2I44R
1Zcq/FyHrJMA1wF8s1RZrgTpYYE9hJix0W4kBjROlj6cZsyzXy9CWZBasjo/rLH3a0XDOy0k/BS1
baozx0TbP/bA+bUQ/WtXpOh42C/jnNKouIbhlo+0/ifqK9ewqhVeTJ9GuXk8iTngXgRv+z7zKRp3
VKbV1YDgg0get38Y8QTrmcn898/d1o2Nlr52mW/n3WLJQJV7UIQZAQjhohe3Y0qPzgtBfGvvZDWG
3n6lfRQlsO+CdsUN+7ui4aAYL0V4QtaMsTzACMXWaesh6NF5IlkFwRNcNldq3xl/uZFT/vGn9p44
SyL/8NP1ieiZijXaK2izJwqPIj/7I19XXQMsTt0OcT6m6U1ulSSzhTrZ9r0zgpKjHqF4CZ1lhu/y
LbYBIJzKZiVaY8B+0wGkfsBC3S2c3DHYR1sor8bcOgBO5QSrURUWUGA5EdLqdQs3kiOVu5w5lB1J
VxPAfu9lm4vCyaONkt1y8GJ8tOCCTPu/5ZcTUNvKHobgsi8JNVlMUVN/tjpEF0Cs3jVmcDkPGoPx
b9u41oG32bjv5luwP5fTdjh2SLGge4nFgET8XEoX8VSiTQKZM4tKd3RqViZT4NrqNu8ouqvHM/hB
rDG7cHr9TBVZiGgD6P5cvD+dDs0lPC0finjxauIPDJlWKqqKilhq3JSd/30FaHxxaKBV6HC7FW4n
7mAtPlCh+s/tJQALfBv1wI66lTXYEhK8BBpn5Yc29g8Xc5IddlNCFHF4maiW7xHFy0HlMNq/BBj8
s4PBKPZXqSnH6uvWv/lDcmRt68v1l308/LQ5HMmQDXU8ikESiMQvsRH+UyV197qsXhSpCmCF36ub
1h5ihWWmsrcUspT5BHcsX8HLYoVpgasI9Gnhhb+xP0RMJ8yTDVvyUS7YsI0bYFL3VV6P2nR2GF66
w67HyUDAwMiPo9H1bvDiypJFGmojsbvt+9g6+OLKoBZUzAZG8MXYNS1E2m5bIYzaTkmtOhZ6/JmB
RjINJeKtD/57LBnshfib0c3r+p0N110d6DG9A+bZ1+or7HT0kGUZm3wDd0vsr7ahO0P4TkvEnOXB
6xvWMi8jou9kPwTBq3EIXE4rRm7nF3N8hFLaqKTG2O5qwPsXWtqnMWaWwQE6VQxT9s1d5/gSf1bn
82aCRdK1oK97HNIqfCkWze6cETYvLMvmvfzuTdWNMBMNBFD6jsMfh+DseoulaZcMDao6eEb1pvtP
9GZtofjea/yt9ONYte1LxWL7NRqtwG7tnHxRuAwwNPdgExssQlYN7HtrFAuP68wPjUayrmhQCMTu
vPyTmHkP5v1mPYhvGJLoY812j0PnDvjgRI2m1Dw9tbDZMy4P29acuDg+3b/THO9GnFXIpO100Ut3
2vcEiOxd6LnW0WxmMc+L/bRroICJZsXqzX+C2iPTxIoPIHFw06k1cLzKjXs4maC9D7hXWEm3VROk
08rvW39NHgcHqchi9HNhLQxJN5L7w+dum2xS9hyMZWUFhkTHp3d7oFro7TMlzs36Rrplpqf19Wc0
z1wCf69Pk6UJyNouBHKH1fDtqz8QAUrx8gAYJKVK8NmXWcPmDSnB4U2Rh7bGBufbhsAZqJzubyUw
/i0cM638ZVPk0VJLbF1lq48RjnFaFbabmoPOj+77WIMvS+A7Z7kig0vo+IiKAc10+U4DZFgoqZAO
73nlsL5LZAoz3aKod6L1Fh0hAN7x7JqEqG33nQfaM6kjhVdbX/GmAwb/kgGtW35gCRAfF1w+I5FD
fGDHnv4Ls9HIZwHMWZmj1wscZtraqUsxWvVlny0M+iBRph9VHstzNKvMXcT7Q36pjEam3OLlRxwn
4TjX1BiOLMvNdVRsMxkTWYuaebvDuhsyj0P9btGsIngxfyNsIEXeu0Hh3RDEBImUaPaAqQWFkByN
7ul+iiQixBSYNPCkcIEAVu/lLh9a6kLtT4RD4+yuzIx7Li/Bs3HR2rcTrjal1/mPlKRTKZe/6S8+
2VCuXbyybsry8WktLZ0he1+J38XAfSaYcfwpwftiAv6ctzFWT3g4PUmN5JfbMLWMufTReT5Ui39F
4hnm51PDHGvSCNl7o/221XFDNa5KDGLI7AFGDRwQ8DmkCYcgtCRqzgXsFKnVYTCJwzBXXO642oGo
5B9nX46gegx7YVYMEKikVotdsEKfuYE+e0qkJpy5OzdYM/ltnRylkIIrnthov6q/OjkVtlVUITiE
WY+vYB4tIp0qpiq/+9dQVvJOu4lDjUaOSrKKE1tqiOZ7A+lB4Z+br7OiyEtf0U41G6orBvU17egg
1ozbh8IQXlDEBUOscH/+9E3rWCIiLevCVa1oqWsxumcWmCGL1Nh1A/bL7r0tKWNVNXtHSYOcMKVF
40hRu/yne53EOSqOsWolT9c+65KHFAvQWnvBQ6+VJfltfQ82YIgh5JTXif4jmBrzKqqOsxifCC9P
0RpPuid3jbsXos1BfOf0lA5qXgJxJyDa3KYY4PYFbfMWMd0301ZJo7h3wHAn6EqJXdH+3rCK2l3g
NP9ItZzrB4InnOURLLurAi984m2lv5gNDpqPHyb5oaUwWEOp5HqR2Pkk2xV4GzYp7NXhJaXS0Edd
kolQGVMjglXCpln1KkOqctfBBtQBLiyFxUMIAWdS6oI6bhpiMD2OS1QG7RD3N/liFlApG4QW4tYw
l1Pk3TSyI7SkNZPqIXBlI+k8fhTk4AvDDl23nfj+Jh7+FfspYKvofZz/sQ5NyxlB00tGzDnTJ9HO
7dJol9/CuYF7nlUTuadns7g/woOCl6MHVQxF8G7TzvlETT+GTqVpqhTo7g/850MAw/LMlqgrhDHs
mVcwL88QdykRIZ4xqn9KyTbjAYKBeW3rwXYd/Zr1Bt1djI2YnSf+VloHFf81SaykDKSXfdJ4/Niw
/Glj7Emo3pxL70tvuVIKHV0otXKOyg45/jwQPcm66YVoT0L7tcz9UpDRHh0bpzLDorEBgeK4Eadm
xS9/994++KpQSRkogO5y6kOEjYITOeQG7N50JXM8lF9U42qmyoROJfH6O3q0aFDmIonp9zUfCc2N
3TUrvBmtzrAE+8UB8a7RG4liwEsFS/EmOdiel1kVNzslM6uzHK33fN6bK9sl84vhyKX/E+5FjIQD
whlIv1QCadfZnrck6+0LiRlBpabtQeIeh0plHPCKpdta+IMxYE9fpkMxlkvwhX22E68y2QSADc4B
8+Yd4dzgh3LY8bvBclwNOu9t6iKJlM7No8lxMhyig62o3keA/foL8HUNgAuM53rord3KayySjLzY
QouyfzS6XI65DhPPpKBhVr/vDoZD1489fFoyerVWzcZy7CMxXibdlB1M0xjE3q1pxtsQ8zGOxyfG
5wECbBr7bDWp/3T1bwlEd5jPcnKUZbvJkcwTut/gCxsZ14CmVHXBYvF0qNMnY6SEdqVoFe/HASNE
KRtoj1JqgAVs/+ziSVGHkf9GEyprsqOpAFcG429ZfYFipSicNBzfC0T6ejNtKA5+krnwBIrpbBRW
cox9GDP5Lv1izDh1kky4CJY/L4tAZquhjqk1HF+djNFjTiJXkK15No//lm9+nB2Mvnw55LwdzbjU
EWau830np8aBV9OKSlv4w7K6nMk/koHqWJd5mCuSQM7/Kou9bGMkxV/clZ51YZjdSY7omTVWdkHo
va8uENFOn4bWhxe41WEJyVw7Y8OkWAKXv56IwJPIn9XBbEuKU1H/poBOrxyy+SCdMubJlae9uN5N
l7/9grDp7oIlMN2DCDxl6Gi35gsa+Z6cq7QWERgrKBoxyVhTW80GNwE5Dlz4P6oF0+navRBUQrBg
RX0i+S+rDY7dEoWp045khDZMXSxD5a5iMtohJNq2ygkvR3BJd5r8rq+9o1vujrTbHYlXVhzyeej3
/EHTtrJ/iyfI3Sriv9yxl8ZK5T369p8OUMMFZ3YHTogqd4XAAkJRYLdhF0o1niacrQnQlGssseyS
pRcsXSQMRNBBNsaSBKOAt6YAs9zdc4+wAwltL+cE68GstmKbFzNlCPJ8W24znpa55EIIQOSUF6xZ
nSVNRWfvO78TJcnJCgl1za31Vh2jlJmR0fln2+lBkWjW4ZVo180aCEaLpXzaE65UE3Jeycb/Ja//
ffxbi555gEzkrhtIJ0+TSxYDuACL3guHoWhpDUb6kbZ5LIWfUO7tUFHg+77lSN6ZtWHJ/ueyXpEj
mq3o/WpguJ7kR3F38ml/LqCsF/KSKSaPLhNtFnJP+XzhpQLnRsS8ykz6RCg6DzlZllE4Ea+JY/wQ
ODTDJHSlq0eBMHi+TZWz8rESh5u9zqf5LJ2eKjdEeqKJwLlocQ8uAe7lSUeEZNUnVZsUgrk/4vYi
DQ0f9FZbXVKVJXXGbauGZVdZCUmOZuMlTacOphXrS6sfnj+Bz8NU6PZm/m/+TFYs3JsuSr7AgaG1
KEWuO0yNU1ugJl7owPXcGTNtmbk7v9xVjqNea6nI89sskH+3haFi5NOHWFXkq4yOryGa9j4ZgnC/
qt1XD6yNbC2TljwEPpkBDxvNHlr2BPZlSzIGg3eNzeHpkWqldTn+vNhDNarIx4mc+qfJGlGsdG3e
2I/N5xnFZHsMbu4HZObctnhDU68MVad67vYdWIn13RW3mbHfT2XSqe9Nn/s8eZoYldfNxsQ+zTkG
lGbCc2vkuWTg997P4heD5o9nRLzlQ+l0NmE0gI4+JEt1p59xr7O4/gTs8n4G2Wqn3yfsC5/1pXis
EDwGdYbOVTdk9m9i85TQRRTIPbTE4cGBz1NoOhnXVFQrmp9Ph3IYAkCquU7AvNgyk6zsAMCVCcvf
AHIidUfN9NXFVqev0Upf24IHJd7e23EWtCSFAZOtW+qBaB9XJXcI5Yj4X/r/9esljvKBqnYTqpgA
4vs/87QU6ZwwezGHyaUkGoRQu8POBMMY7saBTLCN9LTappxxITCPpeGEYuAyP6eEoE/bCL4E0Blv
V4u7+N3ny2zyyBnpev1dNfCujHYxd+jJr/cZmkbgpfHFq263psSyGwaMWrtvj15YtIOHHvinCyNQ
Th+sbvgEbVsJZiVrpGNgZpF7gugeBBahY6jRXUI9XQ/7ox/QED5xLnT6hiCMqVKYL444NcUUmexD
icfrIflPMglfHdlAnEJZYl/1pRPiaPo4ZEPA3w3qOhdkkHEQBsbs5ZJvJ2wOjt5kdPxHK5xHce20
4j4C6W7fdHmysADF90rg8TuKvTvdaqQnnpFI7FO2z0m3bTeh+0p+ISSmiwdJ8zioc4P3JS6L3WyH
Vh1fhX2ETTtOnpqwbGEgj+stewgZ+AIKqoYJ3avw3xfjF6J6zWTlziucZej5VsUfI9IDCbn1377o
4hDh9ba2hxlTraxjGgAG3abw6bexRawxDatkehCgjNpBPneX8g1GnAY40uOSQITX8NjfJaYuD/tJ
xKC7lgkVl+qFV1q1+HyHjbA/Q4biiE1rt5uU478o27tVB8H9kNOhI1CMaoIfIPAuDDN+uPP/4pUs
B/Pu+1EhQL2P3wWvrAZzvOPCO6mPjgne7IEl+0UcrVpPDrSBSu5kzrApF/knOR95Yz9y/iKnlXZe
Q+HP8ppHfxNw0rIn0zvhmBxpTP5huIrLqR+hbGt+5hNdGi/S0x7Z6WrwnntQQMbqxDADMQ4aQSu+
arlWixx28LNLtVWwsU4p20c/SO1ALbGKCjCzG0emCs1hf6DWDjN9HQsg3clYPHXCc9uccNqhT3Kk
jZdwCfCydf8QeX8giM1M+v4b57hlvnZ11dmp2Nf5hqK3v/r95muTKsCr1j+VNvc7SiqJySi9i6R/
KHbXVRfPHacT8mdqmakoytMwSZ2DMYwXbfjgsaF+1FBF2MACrOzFvg18OIKZxICR/VNkytdIljeO
zMQkZCtkDNNfrQikYqczNYxf0iksZI7TJR0TNtcv7n/5BqbIiq2v+xMjgrjU7JhZq1WaC/pBXRdE
XrrobTBE4SYSOTxfRhuVnHlus+EUPYdLSNj76WRGAWmS6l7RCRyHWFWIfVIPJbouLAZDVDpMxO1v
ISWLUdDLJoqEcKV0TTWgnSVAJSDcw5F4ZLolzMndPKwlk4pulPe9LBgsATmP1jTCTgEyu1n2lZPV
1OK4CW56Gc6jZC83vhQTLb4i3LKyvEyiV02nj/MJTfpg9FxCfIGDlkcBfHQFLVF+Ixbabh7h1uP/
w56p8uVLFmVuanzEKXIZJfI7OR7j3WJKaI/ub5gZs9AI6xeDFRTz9AGSOYlo0+S9g8WsfQ/kQuOv
OF4+BrwUcwu8vVCJd/yw2ScclRsbI01NXYw7XBYtyAJvdq0w8R9T4PLX+g6pz0M6Hi974vQgOmZ1
tAaVu51pNUhPZmNXFu78WfkOPy/kShlYkOJjrUfykfBTGnEcGLkJa3P68z7kgl8tm8APVGE+DvlN
1CYrP57bz8Dv+8cs9peeZeRvZHdcOF8mwCDUnT0VBxWNBeWX5O6l4VF06dq/dM3H7daUkS6ZZW/M
AjggclhdZphPZbJBzxAxSjTbQeHFJ9uv3twUZ08GBXz7ZPMRvAdwn42BC26lq9k2d2g1mZd6adYW
ZZMw0M5hwLreuzyfNmLJ7xzEara0GgkMyKehm09U/REk1YUgpVFVJ0yCrNro89PZJN11WVA9jDzH
DMq0r0M1xRwFJFXN4t1UhOidkaSuj/aQ187SFvqBuUds7xvugMORrwDi0DudwN3sTqFMwez8XT6/
IDLa45e7arXiMOYyaUkdt2bpvQfqXLe+nzQEsnGxowBgY3g8bZImIqsvWeYiQJCEU4CgmRacQCHi
+AEJfBNjf3TR1OB72xDOXuvi2RWnurb3BZx0bKMkvAmFVwvh/JFOF51R25ZqXXBxG4/qOo0PUwJv
cj4F7r1JQ6f+QR+T2RAyhh5yS4rw6deJ8Ertj25Zsrh7WD7HtflJ1VFt+oJ1GgSKytUi4Q8PCLZg
lAHWqayvuvqiCNZEQwsaq/34cc5EvdNiTL95lr1MWOp8kpwKjCSlQSZSSlFANyu7bIYUAkbff2V4
K473lFU02h5tNX8C5d5eUkA7qyMSToRrHtc5Cp/RAxj3s+ALpfAVqDWq1YNTlq1fENrR2bmFkEOY
RqzDFGGH0QBPw2vGJ5UwQnAUFmf5EapZaGajS73nnee8iHUif1kYU9rJcFTNovC+ZR4DHOIQhgrg
nk1ii50BO4+QPimZrhk1CZiMHwff9g0h7C3DMTbQW+GiVM86tGCh6KJgOysudo7dpLyOjzaFfzDL
KC9AoxdiMPvVxsfGk2/NuQsEfMOg94oy7u+9EIVQSoG2ZM+fK9v3duyRa7KQL5JMHxE9MSgrawcy
N9GGtvk+W9xQkQOxn0mhp+gDXLqNtX3MqLeV2zko4ErRnVdgU4jquwHVXqEQ9aYrVehoPHSMikHD
ihIP5GEKyX12yXiD/oa9MppaPfsVWQ7oXNSSLAlz8DuaTk8wX6c5U+EubLdWx55e6WJVBfLsAHAN
iPc9IrSKY7d/dZEFBKNal8JxeLaSceNLMShOpiW/whbocNiQIZmLYCgBsRLkVKsYN8gQwNmeqGR+
sFb2mclAKOUgSrJT4Q9btvgIrCyz9VT8nx+mVl0UfrY0KrZFdpXlTEtun2hO8l1ZelTr5UfVYroT
Tjzs8EwlmvlGZov6POWpVzJHov1Xv/d805sXSa2rsWQa2yU5UB6JPUVYd2JWHuSA7ocjWdIEVgUX
LNtK4ZvGimTDXKr2tpm2EvbRHVOXF4Q0uzFgyrLOM2LYhl7Ja8y67eRFZ0l3MoftcDcXI7k3BQ9R
zK9dnjQk5SVt28jlNXVsBVp+KOVOnj3Zd5Zb+CEwirFp63eMQhckF6P8gabyET+caC3VWjm4Glan
8g2MlNq3IH/HfK0SC7wONsJFRlDsm8eSk8ymLdHXV1hrtpjgYA8WPDf/mLDwNJkPyFNbLdPpEOBs
ExuYytz4catDFD4w+cdnEhlqSoqzOyLLhCvPZalKMTIh3UG5or0C/c2GtEgq6FTfToOTTIqO22IO
dirBFAfGiNEXRhLIU+moHg4bnf7R0HgjCCgG/NY7Au9KGRHJPx9dKhq0eVT7BfYSQz636QCguzJt
sX6vR/ZVc0S3W7YOnsq1ftqLBtJeXDCGnKCLV9K5X+/ZRKgskV83JZ6uH9r41dQ2+LeqkDHmdnQi
HkcfH42Bp2VzZlGbKxikKy9q4pKmrJjK6dDCkqW7giiatFGiekSDKFXYXTzwFC9HrcvRLQWPcx1p
P99owh/p8huRFfSUvzEmXjtugL5PGokwWHe/3sBoyr6VH2sV39hVZV/8LsCXZRaSORoAJ6OalOhP
7u6kjcfKFXWb4D+wc15EZLy0TpbfZvQJ2sEKdCaipXbAndVKjwA4bkG8rWQsL5NnjkflVtOHCq6H
vvuFg47oJV6wpCcYrpGyDilu5ir+n//3d/apgMH1b2VYbztY0Fw2dg6pAFNDOwveiu0wgwkqcCpg
/JTXquUfickHNRkmj5Jey8+5iqorxzhKmakuDurhIPRRV/Aj1AE6lbSru5anBB1qCD8odcLRX16p
K3YLk91d3L2ljjHIT3zh3CTZE6Abzh2Hu0ExQ6hM+iX8f0kMiCFATx1uq064K2BvCudSRin+1pgv
6PKCcqBuJmdhpVmUgvkizShpZlYAxDcW6GQzAzNPvRTrNvpZDg/6gee/8QfjuS6luVvpnYeLGMdK
HPusn8PDXGzZPW3XmODusVwfDFReW6G3doiX4w7HnRAocCJFVqfK49bixTXVrscrH1H7ZSu+IX4J
CkS0EfKVsxWXb1mwLQqZ7Q6D6f7x+16UPHDWn677jHwyofdnU7Qj2Pr4pITKbKUN3Dl5suQ3glUk
bevAvJZNTqQSkzFZkpEsqfgfdhc9oE6+sYuzGYGz4U6kYejhsrJjgDQVxGf9MpeHSPTiyu1w/hfx
KUAUHESmpQbIRpGkCpNvfC1Rju6ryLe68iIkzLirGme98cygHaUaheBUA32mIr+tB9HP5lew6nSO
HiO1RUwVaeQRYpd1PckDfwRtnk0/ZZ0yAwTt0DOsAZC6U18nc90YXb91E4UFRjmBETasU4z8Ge9H
868anLRzuSKQZ++tWLhw8K4rX1RvEpzcoRN+Fsac46mQzGhQB0oT3FlTqYfLSKtfydhXLlWdQvZK
t2Z3cCjlghpvAiErjSPfov2TjZIrEhtFdzB7vcuHjz6P4l2DZuPHdm/JyFUiEnF3GjV+/wDr5vLW
penP3DKsatRvosKVnkMtI86a+w5y1+lgVc1hJO1SMyBms3HrDzI8Nte88nxPCIAA2JLY0z3DZPmn
WaH1tpvVJwrGfwqvcoHjd0Dn+Af6j6ladpqvuJmbooNU47YJ6O6FFo6gBtTECWJNy3OpgBujcVy5
On6Xtx1V1BhNrnQ0VMHK5P1Y9UntQSAnaWFfH0Pm/yJfmOpKupfgb/bsYhnSYSyRqFli/y0TocpN
AE7ceiE0w5/nWfm3DmYBnLiR+qfSVsUQsFKPFemyYmbYshWLNdZ8GIkV0efpTHaCBOtElnzYAntb
djfLY67Tdl/eNR0tsa6qALs0qFpMCWGPfS4s+6gUxtsYf2v07LdXf5iphrpPFMsba6a7vRZx4Nl/
Kr1L2ae1kShDkK4/obITv7NPYp+1b1DzxZq7acd+GlDCZsp3jG9uTneBDuh0/QHWMrcUZuqZ6mOv
uzrL8y3xTJKbtYH+cKlVRD6EOolhnQ5ES87g7ehw4b/uCqTLdyLV3rf2OJTbPmU7zLSfgaNMMuBQ
kX50xnS8O5c65dYGCHfBDUKf2rFlnqH23OZ2HXKzUZUHubE/uEjemBphp3PEnkER5Cu8smasxAKb
cptASsFVVXePJVHMje7tcinyCqBPs5uAF8AWRMBgCaWFZ1cwlL/OTpvpw+UyftnuYWrIyNawMVDZ
lzot9afy6kTEa2bmE0XUq3L4mYA2H4bXIqGo/uKWBooP4a5VespxvJ5xMy9GOO0mL2pHQRsTJlx+
v1IqAlFNTWaYS7vmcinAZDgU0EtrzUvnQMdIl6GOEj+XGHmIPuHsn99b2y+TU7o6c+08aBPOnjtB
kcNbSKhaZIM/pZ6QQwKgyP5C7B3/SpVCdx7yii4QvCSO5GcCyfyJHRPL/qdCocpsJ+PJpSMRKXg+
SOLaQHAC1/w+JXojWDDib4eYnEJSYv+/MKTwlWaUdiALHZFubclg70sIgFFoxHG+6O6qvxPL6p05
fzeeGFCovdtAPyFEr9we1K8R1OY5IjZDZtyep25iBQQcmkmThqvWrYOWLVgDRKWad8G2bQJvn9TY
oJDsxgnDAKdqANhVsq/7T0WtNy4H90GwBFeaPPub3NE7in9Mgo4DjyHAaE5dHBOaiPLJFyXFsuk7
lCNDmpLrXqdZcvEFdc+jKxJTbjITTa+zHBUg1btadwsjoMKVI8xy9PrzTPU+3mhU0eFDCzl6Pe2J
WLvY2yIkQb6nIK8u377VTM+1ahrvmlYkrn2gBEg7IFwVnWWzu53ji2+/DKMHK593hnDUjiKTfYjP
P4/4sTXsBdzchvzIYfyJLpWrj/VXaNPtj7I29E2Y3b/FpheFWJ7UldIFlwwjfGi8ZLDSMw6cj94q
Eho1ZTR5LKT+yicJSONVSXxIg97ZrZUlMtsgTGAeR/Riv/dpUDvsvxY5Ea9+g3h3xL2Jux0EVZuF
6hjdO0BZeHj8uhzOahfQwvFUwxYx2SFLtPYEB6mmExoWf3hYLrtOAbvuiPDWxeqpsknjaO3ix/wB
gobuvs/7sRiCAw/LJdWHv6OYGP8nHDjiFkvwgami1i54cQwPLW7TZG7R05LRPlHfVExZlDm1u5IU
VLfKxhLrvFQOYnQffzi6K2LQlfB2T/UTRecMk4Bj9BYViQ+F30dV0x6wy+BXIYJWqZmt0GStdwNV
ZBYX00do6zQGN0GcJbWDcYqFw6souLucZLUMjiFRx2KjVgD2W3PS0AqKkELHkZAyuQRp6K2iZ3yn
EpL54n8lvons0asBx8s6+4vfgTnQbyd4LVRPIBR9wgmzpUXikhDKZS0EghYo5EiaK7IQDpfHZNvX
0pF3thwjYutyx8zUjoaF8uIJ7oaesML+4ldQJY9ZMbGmr1t9PFryHt6s7ry8bstnXrgn4Jcct092
lU7RrWlMUXOpVZGoDQiayHIxWltuLaJ+tXkYlYNUJ4+s4YUJFZlFwqiFIK2+B1EiUOBkV3f2zIqn
fW6DUhgZcSyA2MG3pieULCUDOHDXJMhRnAA+6PY1T0dD4wfBzLR9WyqiNySN9IvcNU2R3F7nbog4
1doWaRwrdAglWtc2H9g+Z24r/jWCMVXYNGb2zN87/FVtgC4lzchiyNZ8F5v683itAEIaw0uaVUt5
cYGXIEP2y6xTTlC7so1otg63Cet+oca7pwlYdnl5shBpiuhLUiehJCsadpyJMZMFqsG91YbR67Ri
EVQ28IQkbSaEC8720x5aqiXpD5arWFNttGayWg+Imaz3q1ScPLLI51TcsZGW9IdT8FVCFcorLjMQ
USsNmDA2bwOHhATe7HaKrlhiCJbgHS+uvAfNVLIpKatucPwb3BpZGrMWItgOQ4e2TmKWuO3USguW
ghg+VhfDKxe1cVpv2i2aatd2g+fjfIs2XY/8wRyPx17M0tqI1ljPfusYKHjP3ikVtRSBNpgtlYuG
SYU4zV0kI/NsFO/87/2SlUe5I3ELWiWnPW/dp2IBpDipnKE/Z9BfGaFvqsSAjDr7ZLCS9q2wpZeb
Ga24ojbwSePG+i6LjCeBXj1z7tvJtPhNZAe22/SY9bAy89BNcj/WZNjVw5JmfASSR+zCTccSNxfN
5Bsyf519LphvKde0H/s0HXG9fBrBVxJ1+bkXdTy8LGEnZX8q41G35cPTXfpnWGu1wsYwhjrHAYQw
1lE5D/MKNTKpMldS6EwlCHx1NrOcHVrNygFSI0/zMbsqIqAXQK8OjA1JSBy7YvTmKvUiGhC4QNDv
vtegeC6vTx8YK44T5aD8b+6s7ZCEkpbP18mhp2m6dYzn8D/ls22w2F3n+Xn2KpvqNlJxfYd9Ykab
AacMER7o/VOcVKjJDk/e2wnJMmrHyta7CAt2lJVIQhlaPXj2Nck+WFi+HYZwiW3cffia3mwRpR+f
cTuNSr1EanyzBuxM44e7J2zuV+1amZ2fF62RHBrWFmWqWIvdHd18pZpcv3zOCm8Gy57je8qfnNFj
XmT7MSGAk1KJKOQ+D7JDG2RF7ccHLbRi69aWR0RsZKbhQp/v7YkDl7IfkWoKpfKxBOSzWgTDDmX5
F8G7vzJ7BCJ5U9bJbI8ne2jz0faI8l/y0VQcgSNd61r0Rzgx/2/zorFMs0zcqtJHFtSWL2tDx4SP
JJI/HymzfMrVVG4PbgkUL/N6OCyHGiivpcBctrEXWjNpPaD1LamBFFRFtN3Gz7tMUSJ2YvQeetPZ
0pWGkhVqXAj1zHkM45DQGyPWgQ2/2FR8V4znPieRkfJBqbcoGLZveACVNTXLlFyIWchGi845m/ak
grDL4to9II4wOT/XBO6LGWMeqy5qMY2re4pB2wu9s43dtpCVbTr3uRXOtAiWCfFkZLaTg/g0u9Mo
FFPK60Vq7YzGQEVtDWXHMTcOXkk2ScpK+PhrJlLTQTh6ou34HTygP35w4NEWnvxMbWSFVLx//9jY
At0VjHBoLEZG6q4StBP2DuVOauLI7TTK7+Xrnmw1Gso6hD/naqAF1EbLSbxBTDQ5dBCLA9byUDHe
2+poQEWoeDSjn334Ip2RVY6Bm/ybCJ/oeLwvY1M3UwBEJs4RHlOthxzkwi3WIq9AKSaRIm/Z8BJq
LbhRThDJOnmb8+PJWvcYa4Fx7gvbBN5bKN+YQZhcmGTqBYJaoOr4KqilEiIL/DAl6ucbia+s7Ppv
wvWt0uSb1kyOf7PUFehAZuaoXNY/n6peVzVDiZMYr52qkQl2A+O6lG8dCPaWo3ZrM2+ep2ZmHPTj
YmvG2QHuuOkhEV/ftnhjDel1NS7wD0B+SfhnJ+WT8nKBdU5rw16BBiopmmcMAg9tkLyZ+sL+2HH2
kXXTZbuVHVutXfswP8nuC4174iZArbOsRDBAvOz0n8bBujILCkdtb/ZLmmn4Re03tgnW8fQUlfT2
duYhfC8Pji/xe687sUXTwkO9aguFdUh6Ryj2f4a3WrHJ13prfaJ5X/l8nFsEDmHc47GQ5WAte4Zz
PXe4Uf6R4HOLA+rIPQSzidfEtUJ42JULVTRaI7lBFy4oWX4/Bp8k/0dNTk4VcMiTYehkPrUXIV/L
RPSFpiSrttwU/HFysBmMZML4KbPZ3lGZMsy8vI0N9HEnlw0i6LMOVqQp+bxwxihVj4/rzhHB4s2V
1XslU3iEniNxmgb0jLaO/YKb+RH1PZWBOmmle1YfVMB6Jox08LA3na/xU8AfEW5YvZj93euAFtjW
iobnzj/SwBJM0oDZKCSPIBN54N9bJQ9mY3mLkFMdHB67SubGFzaG4h0ShwHEsDl5n8rik9hX8t7O
8nECNLiWvk1JXNugtZ7svaNpsOLJXB+NOrIffV8fmKS/gacKTCUckVBDjc+uI4voXoMaWgI2SH59
N1PMTwTAkSNpBwIuRUxvumdMRijiYWZVm6Hw7BFTAgQ7vt5zPhgvnBcMd6Ftj7kzT4SFmRXOJexS
DdhO08NXVYMTW9GKyNZjtq1bdi/WPjcfnqKpM+nHaoOLylHGHVf4/36Rwaxvxe4w0k8/6OcPC2hj
YH943cMWzbuEfqz+vFTVzhK6QPd95Zk1gDcZnSCLw3qe8+QaBt3I1Rfw921yKZUbRjMzRnfWijz6
KpOySXBUKeRC6q/hAL7h74VdMTGClYc1VAFwcGlThwX8r9bdtfcmlI2B1VE536t/AQ8zWBmztEc7
dtwPOF3qXX/T7UJkAAauJZorg0Y7OeK/AbFSgaWFj1O3v6Fk4d6bCKPr07Ivc/Bu4XM6Em+9oxbk
mWVx5GKBa1uzwOVriYpJls6VTckL79Ld02twURroN/ZMAVYzq4O5nxd/d+5NLLOrCkpydXRGxix/
XAEgkz2nwwJbEwn3ehHYW7yFEOnMYlNgwwlClCTWKkVXyAUazpKecl1LK6SLZ6DqZmHxyv1ExYOF
4Htsz/TY53DeYrh9M2NvBdr79R+3H3Ii1IK8jBlu2YOJliL9LV1+QznlbH2anv3MpPS+g4azoAz+
nYJQTJ/mX+n1YGFL/qaTdf2RxaYCOcYoNoi1zFW/QUVLq5KV77YfHNn5F3GmoXZdbVWKUev6OCS8
dcyaDQb9v3okCygy/14EHP4TTc3xuLhsLdosDPyl3p525BirNXpg4Mrla2+kwKIq458fm5Nn5zYS
/NzeVDFUCIwWaofg8U1P0HfdZhbxMuzU4t3KIkDP2PkS0v5o0Kd5k8cQQVABhsPf6k967E5xbV/g
xLIY/5cWE1yyR9lbhP72ZrkE/yXeYH2w4mky0Z4I81cCS9Cmiexy/pQgwqKuiBNmd56N9S0kug5q
Gkeky2DSG838EZ6/25bDDGcnSOqmHpuB1y29RdPk7p1i+H8kA+fmL2MVIX0EIxU7R1G69a5qzSmF
ved3Ucz498wg/aFlflXLx6ilmK1rOArkK9WUxp/IpnKpTP0w5NhUxijksux/VHlQZ4SgyMZKKOmz
qzXbj0chrkZjpy704iFzpswWVwddRpSs6A+rbqyKwTnTdw2Jbz4GMIuKafIUp4Zvg0MnP/VNGVhg
tRgiIDVo0g5EJdbETZ9XS97GYl/ge75ow8GNX8esMiClVgZwpN3VzNDdG75DRJWyNWjlM3Lqvreh
vMZsB+0s90rwwwbOVOVuuBXMc12IlnvV2V7p20ZTKYk9yQk7tiEE/Pnrn2hTc1R8j4tvMsGzdBQp
6C9cD5Q6NsGU4bTL7GXE0cAtC3gv8abz/wN87vxqAWSE3vi2wVrNxuM4HFJ/F6r7VZf0+U567Z3w
f3BJ+XUtaZaTw86c44a6j6NEO+S8bkfEwaKYHKmhCP7lgy3wFF/yCgIfrk8ZSJPkrmb+6vO0/G3W
0dx+kXEzIQo2xE46G+ZgNs0wDASALx3k+VSHaXWNx0n9+WWtTAnlIlPBS5mGshk+7tQiI/GsvNSp
ILlS/Pu7QbltlpXcYwNK1GDGUn7VeHt753whhuEUTNyDkSuiXiMSf5hHN22XCm8rKPAsylTfGiOu
0341owbWZ03tdzKZNKAXwkp7YA5o/8UGhmnIEmfbi1xsiAe/U5AUUmX3zbX8YfzohRkzAGw2jBqJ
/VxoeI8qiZjbiwvgMo/GihjWRH3zLCidxqRS92lVsCMQ1fvXTaoMqZgv7UFLz7wa1BfdLyeST0UF
pg+PzC54p6VVrmFLE3r1zZkVWsulSko4I8F8vREvDF+JGHeYL85LRW53EFSPBtFZLaFDJSOowpVo
WMUww9qqqyPLSAs0SPUHejEsnfPflDa2P67VdbersUz5jzcLEyXtrZQIXPC/dmqvypA6ur82S53b
j7GHUbzU2emK0c+jUXIvwh3VNlqCrDUBN/yb59D23ysikClsFiz6COTAdkzOOu5TWRvYWYntXy47
i23zvGOA7LkTMNsRqP3SKOc06DKFnowPtRQgL3MufElu9avrBqgnJTxgMrwwRke0BW+6ljWbNHge
wHuVNhkTnQxZxUucPzlf9paaqOISROXcVnMLV8xW7yIR3p2NAykENgr4upSMY7EhZWL290n/XGfZ
FL0GXempcUrp/6qQvW8w1yeWiFYN6S9yIvIpYRGGs3QRsGduOD0SEtfB1oQDsZBaLCCTEmDF/yFV
sTH76F+m2mw4XkMNG3SO3CYMG8AeJgg1xMPXtUwV9yKvIykr+AkIrKpQ9y8WMzdYEdK/CgWeW7GJ
909UQPy9qvIB3rbkupRibRXyzL+duLlhqnHlvDNqhtHZlW0tC3z5sPNj7iDuBp73Zcqy2bVQmV3Q
rDrjBfHb8a4ofJEjtL0NV7e4aZ97Q430kElPJQtkivejYjFvEJP3ZkGkpZf1/rZEOqiayeXqFTJF
b+K0IxVz9NymXm5DbCK4tlrbir8juwO2Fvv9mOFxMg8a7I08T21/TKvEP1EK3Ub5l3dz+/uAMkIi
UCYqrYZVh1ZkGNmVzH0193mX+ZFIZwUnuMJCefiIkFLQt3XHcKht4gX0r2dj5hwygfS7eaUlpTqK
ufZ5C6DV4axElrHJRYQfRyXGMvsQ1TbPWSsgSl4UsHGc9IS3FrOHKr9BsbdbmP41BflI28qecrfl
kSCQNPNI4WE0Sz4PHOBZIWUp7ugV4bZIEWB1BB5qLci2+A4wl3PDm+o26+jB+2Vk9eHzYoDmT3HR
0IIR9KNcEuK3/HHc7QHkNjn1eIUwYOZnT5m9E6tjT40yJQHjWHSH0o/893SlGVcdPTR9UaZd9GwU
7MOFSZ/QACDpc7xIu7pk1Z8GEGvYmLImswNpqythgxA63iV0vQAIQq8J2pfxtlZzwNjTjv4sg9s2
HCD96Tgasvgmy1jq0Px82Yc+ck61lZ3qOOpyNEK/51a3dFmGAXJJ69i5NL799uUcIML710oQ0IBs
nG/BPP20VUv15Jws4CwsgPwZm8DLQ9xV7hbVymdn7txy4MMBpgab9yjNxGZxyYVAgbEpIMbnI9dh
vfT8sI8mi53UsLqWKka4VCiMmkdZPJOtPWO3cYDTKvV/N3JLskz5ircBR/Gh5KtuDf40GTX3Hf/x
Y9uQFDQcLSlAwSXFGYcFapD8SljvyrzjyP5SfnpKZhADKcZMAB/i+z9aVB2W+UQ5Sgg1KSy6Qun+
SET2q0ZibFB+33LcmUtgkimjR90Lc+jwsa1EpsCF0/Ru4Eu4KzukTUhSuJKUSNaJsgI6SigYvfO7
d/00e45MW0xdjF1bv/FAxnfbr/VHCI9R7wIeSXzrbJvyoB+LKtliNMhqPr6ls9cjeDQoxebo3JOr
CmHwV7vZG8MNXyAROgTc0hGysNaSC9HPb+qiHQ8Flvxkwj99cA3YgDhMoCTzF403MgtEfvDpBhHT
X1VNwPFo9FjVaxrKraAG063ExsYYXxbLC62d956H7oh4SZGB8i412VVSTkLF/VjqTDUaGEZaeTV+
BnrMxyFMIgDM6SzR7ijIDa0gQNaHWsBzTG5Mgc4UY1+Qsh5hrCBmMDYrAZ1EYwntZVEbJzthwOW4
nPXGWI5BN6SsteJ6P5A6HT2QSwGODre0vygZ0a29djG72Ihae53OXFZgeVECTBjlebNZ/ZECLxg2
nelBSiYflq4UjVHoM8Wp3mrxHfxMapZMVW5jN/h1rsSaIj6G3fe3/bKseAoqy7zoBvlwroNWZOCm
4e3zGZ6r07VWi/cn29xfnmI9W/yiDkiUvPixTcxDY6ZHBrrs04BAPsJwZ+CglXwNh/zQCl/S2mue
VgtQdThk9aLJlp3R9iPuZ+CkAo1fs1sMf/amROwHNvma7SSeeysvGByXg6+2/mVsgRYUPeQWJNsA
yj1OLh0HTeWuyzz9Xxq1YJ1G4fqj5VqYL9nXD6OMm3wc1HhQM3EAYnHHAA9Ji6vhbX/mHT43Qkg9
QPB0IVqR31hyQvQ/eADGl4EMgayW1kBc7KOjVgRfOocGB5nhzNikCxHPSZ8bpCXMyZnKiG9FmDbn
61MGZY6ZaAtdHR5XRw2SJnTC7XWikktrujRk+uiF5tP5DavUM9dku04SvtFZoO5yeu+6VCSzslyS
jv4Eg2/CfIPuCmWVgw3b4y87RC3OCFOgOSdA10zkPRICnm/rMOKwTl6lHQJgo0DnSafhvR5wpscg
blzXlNKfBSgOb/Z3RezOgbPlO2zb9bNWW08j7a1a5fEnEN+D/7Ihy5VE6IGSXM73V9HcuWLMxiOk
ck2dBkrqDDUN0v2mGoqxL8mnPxrflnNtze/4C3ED2tBxw9v+/pZ9g6rTa80SJGUTmGAM8GBgVOgE
YdwBhPdMCX5SPTYAY+2IqIevjRp8MI0Ck1AWPhdW24eHDwXdpqTnmNlLfHzftIC8Rh5CsFlfrFs0
1RWyistcEAUS4Sjz0PVXZs/OiFSekNwVnLjU0BJ+SlB9Fb5Hzz7n7vIZylAtr7T6hIhMuOfOEcEZ
UWm+kwIhw4RffszJpD6GTvfWto9EKZ910P5mSxivsqBnPJo6YjhoAUkiwvuebPlgsgJEjPAYcYF0
ynkRyBQTE8vb8k/9+686GF/DRW2C1tgtzGgZC6ZsT7EYgTZQAsLH/wZiiwJcmgpGmbgnRHQsmSL5
IXdE8Ad7wtEN8eARbffQL4crIsBWqrF29NHta3RRhLS62kphIOiMuNt6rNNnk+CYaJY6lFxTx/3+
G3uHhHDZlYPHGOH7oiQudlagPf9Ci2TtNP+L1Duek4HuFZjfVEY+PmNaxcy4+QW+hxY5CxVhcebX
uCzPann2OzZxejCO7w65rPgbKgfb6K6XHNJqLst8RdjwtxeRDVa4M0DAi8uJC0VSPI5KE9lgrRHD
o3DXIe+gSHQmvoaMNvHlWHoB4a3qYNaG1DjWeULkCCiYLSk9kWmXyb+qeeISf4nfdvfHbBOlvqtn
y+wO2XmFiLrNUrUTNoZs8JbY9zlEPGgKbkLtWd/czkL83Os7VkZA8Jq4/Ne857P+O1pNZb02tRBx
7brGjWbImZ0o5qfTrVaeoCeuM5QP/KPOIDV1LDNDtU/64azVIg6C4IUGwVasT9LoImoiW3yUJh6n
2SVMFgXl/kme8W3GcmAfX+X3EawKuh1Ix6ggldXyuYWUpxreL5yonfht/jzH9lkyaeh1erPA2can
tN3EQ5w6TEaExi5jaCf8oqtmqFX6B4zRsX7nrAjNRMURrNPnufsGjOKUwbkHVvXlnltbrDNj9V3D
/d9ufm8dMutnBVydtEsLMgqhHKWr/eqTdGle7/nknW9xH/mCNxYvOlOm8Dlx8wDou2uFC5M1/Alh
LWuxh8XGlTD1H+LjsQN/TpGjBNwpSF+1Ir9YN3EIBumFl+BG4Z/t2fUV9W4D43Nwhv8bCA+oVy6M
oQTkFXgOrSY9fskKLppXEcDmacIRHcjrIwzGQkhZzpirDT5G9g6igDOb2KSV0R//rtFEsAliGTA7
db5nRNXUVztkNRW7EWwMXwjvRm9D1eZEg8fF/LdF5qo8Ds9cwxQqx6sPGU0DmvC5rFs9pZUFawRm
5VRJQnUCPZkNjFrqkl5Q3EnyNXO3ctqndRCX2kjIQ6aEsjvNrW/5Q2CASeQ4tLFSms9OvddC1ci9
Yz5FRdM9VXPRzs/GJZFWl0iAqo2SyAH3WI5TtH8gJNNwWd5QuiWJIML+fmOJR8GxLxld7Jexidj1
p/in9/lRv2QcLXjjz46jHAsPEVNh3lXHVeQ049gIirSBhxbwtWnpkYm80a9nV9t1mNKTq/r7/b45
QxAD6M1vXxT43fBdtfb+zcjUYEm+pW+Be7q4e3kw/mD2qBuihPal4u8QHH47fnY19cfbRQAPi9vA
wCqucnKGv/XFeJPzEQGWFr3mwVRvxkJOWnxMEvBWo5CY04NOps0PLmuFYIQFxT9cee+XMLojOjZ/
6UpjRvrZF+YIEuW5unCNRcWHG8p5oml6ArCkK7d/RZBiN0BH+CbitkFnKy7/z8AxsmS9OQHmNX8z
P5RcLUVHf++gz4PcnXx4lSAlAiSs27w3kizHl8NOAG1XklH8utbROSLcWFOY00OiJGZp4hbSzS4W
lwAynSx3xklK9MOUyXICorxnWo+nq/MW/DOH0yEe557puT0bxcldodNqsiHSImbp4DNZD3ADTo3Y
HZ9Apaxatbo118k4DYSyrjSbOXsJqLs0LbbXSnk+0dDRkBLiuep1Y3k+B3QCfLQ4ImAvw8aMBLuq
Qhe3eVRROxWuG9XeiD4EEFbU6yLz/5HBuDf7hVd1QzUt+gk1kzM44SOab7fL+FmmqBc6aBOmptdX
W8pPS4T5jkekoUbPZZhj4eSFXLikOMOSGdfYTniK9AXV7SiltMvXOBLkstwMSB9C86cZmTMU/XIX
OtvyEewvPjoJ803PTAPjuEk+AGe+7rGaauoH283l04zsu5pzUT4gsjyRpOl1UvIjSXb8qCrk+5ga
kQ2ZLS5UKSbryCWpmKe1vBHATTZpFDPbrq8nCKDL3N3PC/3SR6boBFEtVA7IU49ZkNPGaqCJBJ0f
IJ+rUBNzpL25ogoPzbX+v7Yd5XIZ6YHbOKeE3naeAyH1ELe+Mtw7A6eIbx2aaIeH2WWSwyFcDKzz
/rn4gaTJHY1obz2J/Bb5gaTQjSA+zl3o0gsPfgSAbrjLhmZKLLBBHrFNTHmL9bE4cSMRej/isq61
MpwmIdnRjAwMW2xom/H7TBRj9fu7UmpyjgRpXwfx92zkuNMGuTdB2R9QOY/LEdw2UgfE5v6GvPXI
XPfxrn51d91rpDbxuV6UgJ+N3B2K0C1vT1TIiu8LquWyOFNOP719ABsHyDsa4HdQ8RcKoNQKmM4V
lPCdMrmiZJFOgN1CIxERUUaOMsFUY+2u4X1qH3v4ApwS9Mye4gQ2xNNncrgUiIlpoTGjgPNTmY5E
69OazxZsHn2Lckp0O4woV6zLpNhPdbEMsLT1dAA5Mh6Bo99b2UAT98cv5p0o6kMiuzVxU6YiSmkj
+n6IWj0Y7S4+7A2hVIqi5nQNqNC3GZccWxtDdLy2asqbtkfTj+RpSuWn1i5QqKbEdqoyp+40MRqZ
/wKkT02kp+YxI38Lw5mizE+jiGxii6BeBsz96HJ0bv6MiHoRWoHkQ9qCZRcgmzH4rFypllXInfBi
qyuk07VbVg7PGCgajIKppiB26PLd3X+yqrqzrEr2NpF8fS/UuUp5I+B9xHAkDEn8D/rLLj1qZdMs
6RcYbyhJt/hKJgzfrRhPE2ZajHxFXoFYL1caFSJqjTI3naDeNmxNTi6tDjjuPeYdOJTJOE0IBoNc
Q6iHo/RkiwdAVPeSfRAYDd88YTRaOrSbNms/h8n8rvkWmI36TKkXi5GMm9BM8q+ZkMvj4fyB2TwS
9/uT1fFkQHB7US+sd0AtkqoeJ1urEXTdlFYr+cwxoOqe5oF8GWzPIfKJk9snBI/tZB/awNnW2l+v
5YgwfH09agNk32XARl321B6g0xt+UanQJYo/fTzraivS7OTKUyo2YYFmJtot+jelKo8P7K7v2DGr
VdTtd4FXuyPgW74E5gbqixw9T0VW4K4HqkXBzFHMuS7lt3qt5q+ainR5wehWIcNb9mw6Oc6GkR6y
yG2e1GPpKMf3yCU9S/GInLlkQQVOuIWhBr7cSkEK6AbsNMQSWL3vrMtIepFZgz1RT8LcMGIIVsEi
BnkPIlK9sLTWWwWKsKbE69BetVWm0TohJcKvQm9ND0dMXtqw8em30IKVyCp4JeBBiWFxJU89HNVL
ayXHp4drTeXsPDv9jRRlzQYrYcopsFByAuSuf8aO3cNkz26t3X1XWcRu0/lgh6cg35RgXpR7w7g5
5VMx5biHzqs4eBUVDUbkC6vWfe234Zj+0wGFdDfWNdlrBhnmneWiQBpgWDlIVkQH5CXgB1qirWLr
x/Bk5Hum94GIzU1wuOHje5DcO4Ye/mq2MNNV0+0KSIC2apmCh9yTIFaoydEkAoLWf6dp97cSFLJK
JHupJLpK9xWmA2pFdpbNmIrxgg6cwyfdZyQTO+hhbhxYfuHyhnLD+LCvgqoCcjcLmRCI1PndXK6T
pE3lMlz2CFcUk7jzgQtpZI6W7fnJvrhcNrElkH1rYgbOAiP1w+PMBNGa3QEzX1rX4LAHjPwgdEsG
RVrM9paSiPltHjK0nNptk+RNuXQDExZeam4j71Sb19okF201vHOwLvKrovpmIK4GSjfqsBTMJUmH
k9Cd5YYLlHW+LisBy/tN0aaPH2thzJZFBlPNp8Ny+VV/lDgvO2E/4zfIzJRNRNQyiltFZy+oVK5E
QPeMoKuypBuIXoWE5bL5YdShJIRP9KNMrU/KKcby1MogeFcepcO0UyLeVSxGiPZHlWxciUIICwNa
mu4bWOgW1s+FUzUN7V9MNhuB5ur5es8EuUjwbutLUaFWG30jxmc9vaFq/KOrnSc/sv+550TuoSHj
Sjb8n2M9BmBeiW39t64ZzrktYyADUBwYFqH7T51T215R48raTGWr7JpIO8UKucrugGfJ/W/dIP4V
uWlr0m+B51yYsXeIy4mbqT7GbE02UT+TqYN0+sCUbUyEuf4FbhqCGs/lplm8/U2mUVQ+YBUlXu0U
V5z7+lC3VgXvDP0U+8vzlf2kcuWGDGJ5CvYFC0SR5TrTQdFmcaqafGGgw738vHdMpD2ys5O0Jphk
qYYY5kg5Db2aLlnuCFppQDKm4vf/+PcpfbvHKJoXiJVuODs7yBMk11OdfskMr6TRt4RV31DR1tV0
pNl3ooDE7zjFlstFjA1gLlezj/AQs52modChr88m5jwvkYkIWWYg7kv73sWLNvnfFaNMzJCVsSzy
I0cdKOsSWX5XBvAMqk/kIeZagp6G6p5ts5acnx3uv5CoN5FiiHRQ2zLgiJwhwQrzeJFQWwjsA/lP
x+P0iI4K/xVRRJsZ1kMutouYR26amtOlWxsIN58kOvtWhoqS6RNDxt9HCUfezc1PNloVYF6uqqd+
w56UflNZh6MXg5+Ui0h/qjXsRU4rPR9mLTyYaCoR1iPg0e9e/5bf8UNO8sgy6SlTGDfwKu4OFtBk
ovleFyAaRVzmq6a7ffBvI78DG8Z8nOf2kBe4LSLdmIRmMhQ3PmvusBGks9n3Q4GK+bec6n3zRLWM
KKPGz+R4gjOFmbBgkCB9AxXqxI2Jb7E/LDupc+t9K7CNt6hVPw4wzyc8uebiL/e1OPIHkDd4c1oO
1LrFtugc59W11BNFmc/vq0Du0VT6XXy4Nzt4FJjJ46YULhVhqvyRcKrIUbujdNaSkllseW0Gqchc
CMPxZD45e5NJOJZNDsLKybsxz08ppg13GlIxzqIqjVSuI4tdX15OMavziLZ6xXnIbmD/2dKpk3id
vhf78Z31oWRNnFLnsH6ZylGOiU3wywCBVz42SaOmCYZsa0DPH77pyv0M8lubiP3iUkEBnEebCF8N
3LwSo84SxvBcAe0xRextQN4WdWLjSZCt+/UKElGe8+5JN5glLEBBQjhsHoihXwR+RxvE4bgwqxvD
ssQB1acWfDoiagzbJIL8W1GZeghOTvRLh1PS5dgiQmSvjEvhaUMajTXaK4SQUY1WhVOYKjKF6B2d
Tro3JcO57QnuCM1sKPEVCkauRSMCprhuw5gwFAyyjm1Gxnbh45W/iRBS6D4yyOIqAYYoSwKnxT8m
jse0+IoAiSATJ2nlUM2EKQsY1NsMxVQqf0PaDlKtR6OmpQ3mqKTjaPNRSNca9n01jeyjS9BOsn3T
aa0W6Ps13J/hd2dlmf2uf0N1Rv1BWlEFR9OycQ+/InUK94wHcFZAA6lPqin3RzjxqkEbdOJQoMce
uWumQT4P3uaH/7g/A99Q26vgAS2ILJ9vdmJzsDyFhz8CcXpozQ1Hk/q1wXcVkx9dIzM0v+k389h5
sZCZxN9mWV/3MsmE7NqTi5iM0MOGRIdw1yL84VIj77q6UXKNDWcaRRb0Xkljh4O0bf4hNIRH/5q5
gNMMlkGijSjjI1STdgORbgQPM+o2FAU1qv54asUsms10YbOP/XCwSaayF6g91SD39InX5eYvOVYD
J++bqOW2QEU6GvS3UqSKdc5HT5hWRyYyvIwIzJIt/Ou3VsBzsoCQInUF0dshdij9474ftXtRQJTx
aTP1OtHHjLZxbsxWAAO/f/p9F759b2y6MlMlXRDXYG03fFob/zEukfrO33BSY3eFH2efujjGkCR3
tYp4q5IGJ87Bfj1m5sB5y93ZxW6GTRfV9etsfiXlhNd4JrzXFvpSHbn0CY60HuotbdwMCEGCmBLX
DpiFxSZYz5ut7BfZhW+86W3KErdv9U/naZFDjoKIWNic7oHw4wVHU2kGWcFbvyPibYWYgxy0VDd3
nFqQz4fb1aedJNK+tW1tSjlfLat5W7n87Cwhr5V29DPEpP51BFRIDRMPfhrxGw0FtiaAu9Difct8
o8PlIpQcdTqqe4qGIUnpNtnxaEoJaLVKH9w6hT6gojjSxXygpGCivri9iuvRmO4zzxo6ehFzl6Mm
1LfaKEFGQBUFsZ6+BBXxw8TJVdhVUbTFZ5LV/yRmVm/ZK2J+REu7/F56zGd4dQkZ4RzgQqQIQJ0C
ph4tNWT05F25sE0n392uEBv95AsjECXLecUQ6Weag5pyvsdPXhbe52pgS7Pi4FBvN4I/+YMx9Svv
FPAWlpuIww+YxsfNUJ1v6bJFZivTN+lQ07tupkS8uiUCcg1qJyG5sRYBMrNeHXluS/nPr5/EbB8Z
W1FnTZJBb7WcDI2sxIvM8HKgn4cr6jT/Ns3+OiJaOhUo/E5r0j3ApLbe/4UAFawdmAaVSOn+vT53
W6kBARID6BZ9fdud99+FKlevuXoCDPz5G+UwKibBzy7Xp3zqlegudiXTlvDqXTdoBg95DXjD2qkP
G/Knr9mJbsfSN2DQhRnQcvCwe2hQiCrW763QF4WNeULAwR/tgSGK/JoqIQ7QQUaHb0bHRL0NaA9e
yoK2KToLXbw494VeldVltkBNwPSZDjgAvq8dayBBg5kAsOl4zYnwkDkFBDZhTfifa+mxZrS6of6f
vJVAMrvbHDTyejFu86aRd44cX6tzkuKQ8y8Z3AgQKXfAT8xsoxYiQrTInoYfHkpp7uedl2bu9GnA
Tm7M+JhSqspiNGHEpYMHOUwxUwx4Omt81zmwpXuuEmyYhcdY0saA9ixekmyy6Ctf8f3al0LdolyS
ZWEMPulVHWFedFCAUkBDR7gsk94YxUCs8aWHWNlGOifzRlcotUJmYkE5fEmJmrjn6t4uOTrxij2F
K/acThrhcM5jKNmX/aK/lA8s3Lp5qg+NzxCd+m9YxIgLp9XSQY/qaXtVvDePiZ+mXWKsloLcFnNm
BiyxEVxJuVEkZUhJZ60jvpP5pz3MMhbHqXQCu6LHO1pMf6ORr/bnXC+LFRCb0BgwV1IbRjxAwTkm
c5bP3pamh4CbAtgjQYh14vtT1jFUzTy3fule6AqMNQfe7YKYQVrgDMDI9G1XIGTTLPfappNPKEky
QeNm7Dzo2knDkMADiGuzgDh3WHENprocQbPHW/rERZRRlzmnk27XI2IFbN9M3bBX6k3S+cojNQop
RRKp/TxXM6l9rzrqxmjsToRi/3Pv48IuZgxP0zpUmZpPqLVzF6foF/RSWlgkhJwaKJXwxSKObX3m
VSrL9OM0gykNN8tBj3d64ORzAnxmznseHPLxty5Ty8LH0sQiMGYJirtKyMJJfTUAksEHu0EUHkZo
pFOx49vhx/0xBEtstD+ApPv6fNIff3FLEKOMgzRhRcrcDkoQwl7eKq0QEtNm30v6zkm3YnjrWv/X
uYEen2UMrsy0Z1CNVCJ5M0aDbAiv5x9eGz9QAb4Hic02pj0/sIbXwmVtI3rV67cjwMKhV0LCaRVg
Qdg0oLsLUDrvkWDHZtGu4tcbhKrtaia4uYUlAjRVaRMRVtRRkyvvYSdvq2iPe6PmaJ3ecF/s43Mt
zK2kDaGtsHbFsRy8Eifq684Zdp+cccCQtzkjwfgM92GijbVrw13jU1stZ8Z5Q4nI+8GALF08TRlq
/tRQNJKH/0paPR/QXLmJSb6XnBHKYCRdSXoNaZ7tjP7wQc2xfjPZUe8Ez/YaRE8W4aArBwr8PSmW
T6ReOa4Oc+Sadz5RPaoiPc3qkIRDAQbbgt1eucrm2Uq7nCjqwanXxoKyxeACM80eAGpssRq8BwRy
SpOBD+ynCCwvHV/fCxqYXTJGqPU9r1Kwl9N1/Y1K9Uvnb9qjWzFY2SstiokUafszH2OXBzVwYNBu
+8TiulPA+xGhHvGdmQbuYqHLD/P5zCnniMzeXDfccw7Z74GPfPkpNETNXQPTe4c8uaxCDMBRLpNc
UE9Y+tM1j+so4mT4XRrzkltoQmcLMRYYrwQUTy5BhGole5vvd/RzRY4hlnrWqLSWoV93K2qJBx83
5gUttHQ1msCEt4fIo2vIvxjr86SEoE0ZF/5zQcjppDuCj8gkTem0ViSovEQrkHrcjFx9gSsneK+n
U4HCMp4q3raXQcasMjYOB8D4l3T53a8+4+ez2+G6CIlKF3Zd8xOBvYOXEr0y8mV6+FmsPWQ4ctuv
3KJuIuImzeOxpOI5lfHNWBYOpvhoIcd7KsXUGO6onpH8XPrjFydaPvB6Et0cg6ixA+RiqsPCB9m5
6fj35OIw4skWgHFiCAJZuNzsM9SCuvC6pKMVxd15MfX8nmOFuSS5tuZHSUlNfS186z3ACplCrMZc
MEA9jgEWi1EZMQIt6J33wbjW+Z+SzKRupNgxYJmEH5noyGODZ7uYGVLbmuIChoE2wiJxe9cv7C2r
X95Eqr0rEWjOWnUf4ng549FDd8hwtKHmv5A1moeJcX86EmmppXY5onKsvPsNYXFmvlw5S/01JoEB
ViW2v6ANtjLuFoXrVQsUQ9KuUgmkstj1VCuWYHRAuMMGSEfgMSiUVfdQK5H8HLqE5JcclJBG8Vyl
qMkRQFp077PC8Cd7+6G/TjKsVQT4012oVGKzId04NXBP0Z1o7oqq/EmM7lwEeRcYyzXHFIB52qmF
WndD1cEtj+vrBtzE2C0yGipQDL4aae8gy8e4GZy37o3FJVq4/iIF73n/lNcCZFj3hDs2FNPElvaM
nRjLYkwbBq0FVyDgYYlfxkbxyDMkC82a2leo8q3yCz7Ec+Xa0Io9+eSev/YMSRZJKKMJKSogYFwh
EVPNwGwG2m4XzjYx7dsurnmWNtwZOV8NS0yYA64df+AeGcGoRmMj4Fc8L9gzDH1t/x1vV/ZnkXp+
XbI+IdCO2KsceOAVA5q6NHPgAZrHFKzdch+BfK78mV9nUzQGhq/LYLdwoDPqWGd6idtjMxE/f0q9
+mjvPUzqs78BFFqyiCPicr5qMZlvAGypGyvxHUthEM4jbNt02TlvYcnyPaI3N3uLiQF1hsJjjmFN
VZgZytY0fFCr4TtW7Zj+WZ7hnrS+qsXgacsRimz0q5eO9tFuAvLW4qpDi2E95V5TcUYUZFr0fPvr
fJos4X7eVm/jYTMXUkul1//ebI4mSa78nCo4SHt0UpktVSNn+9DQSwFpzvLOlJkQCNYkfooMkaxy
KAuQyvUu0uPrG8T5TVC/4awzWEP2shKy3KxoGWSNmygrImM2WvOZAhn/5VBlpA6pzrjLWKjMSzRR
msmAgU8hJTzpbz29WbRJRwCo7v5X9T+UeK2fOZ0nWhlzbA9XMd0DzhhEUaVNnVb5S1TuF1K2Lph8
iRTX4t9ncYNiy8/yqcOeB1fAcAV/Mb1dr55SA9X5dNW267U1jsRU3QXNjg01rG1d8f/hTPSx9Aop
H1tAWkpsgmhQiiC++ay9auyRRb1j0rGG6nkUUdpgf8iQJRYJ2BCz3jWKLnXR1yH1E9EF2uIt6gjn
8UlBmZ3JJuPQBKpVZOe6gNfSC+h1AGUoMDTGuNVTNW151B2ZJLcogWhnoLFuZWS+oOlMx+EuYn4Y
pOGWnI4FaRGA2WS9ccXFu3Z9gAlqkvtS+hZ+ewKwv9WfanU67ixuMLK5zarhtzPqCXunCIXYnlTI
cF11t+5DfZwu/hgUGpaWW35buGFWEcopxSyn8RHdir53iZREUuWMQxOUeVrisQxCoffyOuvsO+Ze
s25wboLAe0efw9dLexy3pVD1gAVccAKpKZf6LGaMEFIJD8ndhdXH1+rtcLEp6nHPA1SO1cE0eoyZ
Pa/rDxQVDbvhv5XecjoxOr44Ez/hcPnR/AOX/diJqpV8hERirDp9NfsBuRFFvf2XswL2wHFLK0pO
HJXFBJ5mplJrWSMH2SwmGGYY0ohL78u0Ecn/4zlhhMwgsuf8rKG1aSHJd79mFgw6/u3zqEI1UXVr
gQJJHh1hadG3qKgx2tcuGSuCITcvOLTJ6/AFRM+UmNcBuuheij2aDYwCNhZe2PdTAPG45uIVL4Nf
+Namg98ZNrLlexaSfnpPa1Hi0q7mcX811oNTrkPJcHosB1DxYYE7hBnLmNnvVvjBWObSFbwUDrYk
a9hv8asHVxQEA+9ZGGrkkd7COiV0+A8Aul1i19j0xGJ5VFdyqL6LUz3LEAC8ysrucm2wjh4iqwm3
qlo7uL7ATso6KyS44IX2omxSu5LsuC9wOD0edqVw1YN8oNbxxn/epIX3AYE2mxy5xjd8MGplRtuq
EUJgPtANPl+eZeB4oN3EuR5JZptevqRfK5eitUK6nd5XrpK7I0+E6UtrsPa6riLmrwnHk5Nh1fws
HlT0dSBk4IEJ0ibq9xXtwK4f/KKcvpSabSwXCMbLuZf9m+DoMEG8rmSRiuieKdzmSJd53McZvBNw
kQpwrewoCGS5377Ex+XtBrnxrn6xAEbqANzJnS78zBlQQmeszE9t5pOjwKRUKEjlIN1immP520s6
O/WJuNau/Fq/smBddbbvrjTrIFHvvaythgQDgRW8n0COS3J85au6ClT8mu4A/dIg8lJzEq8V6lSb
lYC8+r08PjIAeZjBBCpWdRvT169a2R8rGqqoN652DdZ/4Ql/DhJLpJWw3LnH+gfSEFixYXsxtrVX
40QVIcnSuvOHGE4lO0Wjin6P53/kgWp1wA/eM4rNVzblyW7xODqGxrjYKIyDo/N4o2LRTAj6rYxh
z4a25DIDaJuv8U6EaLQFxgoNOBLZU8rX9RoHU8CZ2LKaDZdnOyTzbNVXt4u6ongWivEiim4YxLwz
wJ2jjUuqyy3VDU5QjJnoJxz0dr8ziqI/I1kyrR+KQ5cUOtefkqbyesJR+6uWlnQ3D8fHxFWjVnlr
3WvSX/8W5Op2b11kq0RWug0Dx6D1cpdBq+1S9QCKJ+H4XZNQVp/98IF0s0c6oB7RnIlRyZ2jbIjZ
2Iq/HVPHVIKuCfBuS4jghbXZxHvXlYJOWm9ROSSc9jYkiolBrZec030mjFq8cfiz8hFdKJwg95/j
erzSWgWM/72R8bMaB8IatfMDKqT5jgrNBuFl5RnjWI8do+Uw+iHKVQoMRCPn+5UrGQqsZvPQAds+
Lk5F4ukLGR+Od/1b0EJwK51bHuTdMeXrxnSWb7Jpl9r3QtwFrixUsSXss7dOuI3awUkaHmW8q1Jt
sNw3I/AaH27SNygNFXOlPQY42xPKC0BTjpiG2mCoZUjA202/XHEio9QNq2IE6OF6VIz0Z8pj8rYg
loLZul4hMXatgjMZZ3Npl0peX0bQru54eKXwBWk3LvtrgZqW1//gz3V5XKX5ipbMjIeVFhCeWjJi
C9SN7pCOnJSeGawOS1vn/8PHVIacjANYohxkqLbv3W6EIfCgS2zXlnPG69hIvN1FQembssSmlGns
FFuEsO56uTDM/rj6KCY5E9VfUr5TFpO4RN2vlqxCv0yAzSlfamApjAuTEYnnl5svfbyxTeJan29y
A7Tc3kgtk/TWSTFVwLPzelGWVmQe3j+QTpoBpj1G6dVgUsdJ+nOdDDxB/5+V3Zf7NHVtYNshxvmW
iIcET6Nf1PYc8j5khBEEEu8bOWr9k5bv/swjliza/3DjlETQcgHWNJbaVhaZvhXVOF8ZpffyGZaT
Ap1HBjxckuN3oVbP+Y6VoqgLoUNflNRC1Fj/yiV3QQAdefxbgszST6ukSfmNYV0cTs8ssepr9zvY
Jpu+0Xk/74fqDz1KPG9XOx3bdRE2jci4mNw2e4Db18diZtVl3MGwc+5WSGiNf4emyI71dOPzXHoI
MbBVXHiUVvReDpCH2QhNW3HRvY8MwItzAtpVbv7hVnDv4rhICs9BUH0RFAcWA1pOroaZIqzmHwIq
vtoLaMKbvY4vCnCYdBn5BogTZOJq3B3bDsF7et5jC3TQ76o67mV+eOg1pLxc9fCyJME4OsbMzCxP
d0f2+QgwpMKbfyKWA27rPSEgIJQwuXt+OQDrvhwXPnbaUsqfi9KIJ1WKye1IchOMj8vXnUjauQCe
uqVUZ4pDzdZE+tFhafQUN6rlV0WwXFmrv37m3wL0ZSPH0fl0UML+ptXn6xttlzOOIY/P7uPqQyUo
rRXPPfUVq5cIs9eXFvRMdpHSySHNx4R2tri739BOg0ioNm4PL/FbzKK03eSqlV6phqFO8mfH72pv
cBx6hxppO8rqldnNlzgZnv8m6/ibJzptXVfdGCnRHSK5LOzOHQvqFH3oJwz0XZ3O3Uiq7ObNj01n
l8avFH5ASA1i9HbruD76sdiM3Ytl5gz3ucbTZQ3yeUZWVW9eBbNh6mP3LCjSfFqMBLWu/EkomWXm
NQ6aN9yDdH2dtHUtmtDmVDXKjEXxq9WM2KH42yMNMqm9zPxYfmYc5Rd/kmmKNeZSSWDGohoTb9l9
vR+VpbCbkYIAb+fzW/3CsxpBzemhWGXaTeY0ppgmsu/Hv4E0LSceckEmZeymR/AT/CKQKERXY9LX
pdjyFfYScl930yH+zrmaoFl7vTHUoXTByzRh5XwOBFP78KcyMyz4wkaVdFmQstEemEUxQU+TLtW8
WTGRg204CoF4N4Me25ewr37Td7V5XmmggZGe9M2KLTw4FtYvOf8HHrWGxZXAi4xQJVhurNU0avuM
65Kpxj1Fucf+OhHb2R48Q9XRN6Z9BpTNml0kjBgrMIIcKXp3atW8Bi7kft8IHz4AVAU26qPWTGl/
CHndzRo7uVXoBqsjmPqq+Gsg2ulE4tHSMTToPT+QGsb1NU70/pxUytqFEGesomEG4LxIVs0EKLxV
9tPwQlfQQv6hU2Ct7SaXa/N5n/UrYW2otMhTdexM7/l3jXQZryZ68LTzHHqZsQ+VJ1B9ECtK/LTI
cHLjCY9sFtlLpnkfEEBHsA1lhhpSzgWZ++ejYf6/HarMuuW5/VlKuQ0zuMUJJ1F0Q3pa23tq0oyI
PQBI6F0FYD1psaaP3zjqglwOrj4pDu5YF/cjrHU/dOW5dO05HZIdeM81jz2Qm83CHiDSSlpqP//B
ajjtH9XQXDXTAd4yPDvQUMKHRHO3PaR0XSk95018yhovnyK03DflQwKTum28JcRoBVrX7o2daMek
7OiDMcV0a3zm0PV+kC2tf3p5wUtqQsCNQRcs/d3t7Z6WPk5HMJJTyGnLIxqi+bznU8v7QZz4YiP5
LxvrLFe9DnTWbMjBRP8R405+C9a8Nkylgw1fVoPhAq+su+aOhk8E7AJTkx2jVU4lMB2ZcvhJ7zZj
gpOg4EJeyrfMAtaGS2W31MwfK/zqhe8DQ31jkEIzI/QzUHPZAnONBVqiVtIDn9y6b97gnH2KbdbC
55mG2GP1OL+CIH71tyqXM9REfUJkGrZxsvB8nPeFJKPtr8sO/mueDIewcorq01atoTljhwAaNG6n
Kd3v5cfqR3IBT5vYO9e21da1FK3SxlXUmJFFHQd+ixRTs3XXVfaWlTDby/3KRRHdi+nhwWbSBy/K
yyVTSHX+zRnfTMnI9fx9JVlwIr4nsVbNI6/8ZDL+v7FpD+Vqvz8e/pn+GuFrNzsdeb2ej189clYP
E5RxT/ULLbUWh8kI35HI08Pgv3fWbuoQIYETXnHpxKWPTP1VLalK1i6naY+WGStb5Cx32wBPdZ96
RlP3/O0K5eNpZMI0j6LI65jGNfd/l+S9rhS8pvFms+8aqNq90BwOFLctPKN+wmUJRTTYZTZbQo3M
XPuEMvhM+/Vq3s6JWFRJSsH2plLR54enICPG/vRpbn5QiWC7mnZvAV+fM1aRPaEZZ64hddp3Ou2U
pPqLm2VdwFZfBA5FMl3wd64n9iay6dDkcx/i0QxXjD7pB42Gj4ryacAis4eBz6KW8GCjxRDTjgXt
erMPzgL71+D6N/F6YX6xlBblBQLOCxjXLqMOEtXRsBHGoWfdFX/+YuWyVj/GBA6ciPjxnSmbz23W
wH8zfPBZ1AvsVjh/uvp0wKkoHWUPU6SLPueuJ6ooH469zrOLgKiyuIvuTAec0Y5wCo3VI18vc6Tp
vKXuXl5NR4GjkoQQYJw02c7AZxUUvL/oy2N6whLB59HhJmVYQ+6T1tgzWgHHDwkPpoVd6Jwb6eSk
YILLIOMZ66V1q6T2A19dbcYOVt9c/nAbONG1nlZV7h0F6mxj0GZ+vM3MFhsZ4TXmfOvjTDziTa+N
6X0Lb2xg3DI3/nwUtNAvGYleuuB9srX3+M83icnzFCODAhCkccHtFxwcg1xomjZKghnGcm7XayjZ
sCreCy/3x/JtyxYof+lvz9Yfsyfj9ND69wTsErpcE/erX1824x3oj7ePan5iMUwcurvThvy3l7Gp
94I6BZPxDFER6PffXl0eqDEy/Cw7k6nae12N1QY8iz2pjbjJjX8rqJVAjkJrv0AwkoTgrexFae4F
J876tC0rnPabAVAeGalhTbPfbQyFoeW05khlrHrPQDr2tzR4NVoHwKiuito0SIRtCUH1xc96Yg5N
Xx1G1Dsj7UWlXLDM+Q/wm5KAnItRldYhwvSGd6BCgPfbupAzuaOSx1MMNIWAVc82b2r2utYccHa6
4ZbcZTY2bwblFXgGo231KYdVmvxsiy7MZTImXtr9Z/YwyKKGQRPTnu5zahlcdfvHBVywTwht/2wt
PCGw6/o0sHD0lVSyVNYe3GnSv7CexnvE5U6PcgB1Xp1mN3XZdPoCe+lT1mzeA8AyhGYYzu9/Lbdp
/zC+808xsxtwPwkJGxE8HA5XaPFsPW7yjZ2Vc+Rkr9wGlnIRknQv4hqhLLpwESXGCwYthX6mf3aj
AmBsZ/0csm4OnlfbFRH5iVVw32YptHolE9JmQLfM9rSmrqKmt3IOz4mmhIuI99I22ALxYRsuy9E8
uKp/dkVs9oPj941MQHXzYtB4mBs5i2P3ZPY5/HlnByiBvwm/bwFqnI8LccUprMzIoEmOdmHfYCCt
z6X6FcjBLrzMqMUODMokLBih0sgkyqqIm6JMrMc6DL7LCRLYlBIHQgHqpBKCiah6tXrqfSKfGDqG
oJwvcFLA08NvVWcP29815uOmM5pwLgS/j84/Gw5z64um2siycHqfk5Wi9tArJNsR98KGJPbm/fYx
EcjZOCeZyrQ//kZwlIleAHYSG6zZwY12D/DFKfwfkCUgpvIFwMp9jNp20PNH8ljMCtvpsl5lJMoo
4iBIPz++Bv9HtZ34vNpplaL1L5szd3s/MvZiPQdEajAXhrLoSp+GWcr3uxieit2Voxgnyn9HV+yV
kOolIBweHZnJVMecJ917IVnWzzdo9Hb5DHX0JQKoGCwHfZGWmLCcefizX6SISwo+WdFYM0d5Jm2A
eLnZenufH8h16kpNbTZ4XdW8sH1JnupJhOADjC3NhDwPF3RKGEw4po6vTIr8UXXITci5r5DAZowP
UAwSHMdkycvj/e5InAqr7tjViyDEu/XIRpuW/vBCSLoIsTjOpp/HBWMy0S4gazrDKprBrSXWOE/N
xHRCxjRb/9sBDFXYrcjPNp0hiHtrWJpFg+Z9uoMJYOblAksuUjoanMI+6cNjDdhxwXbdQxsyuE5S
CX5Iz7vBqh4STfTOh7FdsJrZCbThUGu7+WT3QXLUxtPGDCphloj/QPWkpgN0ZqptA3di5SAykO7Q
3jqBGWIFB72BlE8drbnoVdUJHJ3OVwb/jmtXm0/Ovt73SphaZaxgcxOmwvj4SRWrI4BLw6YMs7JS
f3Kogfku27K3KuTU+ZWFyqBCcNnhEAUCBy8VzhirDUnJ1p9WGdPfbECrg1x4p+gMyCYZbxjjNf5e
haczOVeVEw5+jg76lfBPRoI6sVO3m36ZCH6ctjc4dJEKbjl8nytqHKvF+FmAGxtOl1pwQKpKPmvM
w8aEiomr0zp8JcaX2EdD4rajtFUy3VGkbLCfC3h7TIYUsxgWCPw5cmxOGpmSJn9pzbYmCPu7Y1NQ
XGGbT/YwcZW5b9RnyOGk4rrrhZf3bq1DFcmnVXf2Y/pNShHb4nxzY3KhJx2+r41P7aMs7lfEl0zA
spVvR+jZEWFLcVhefrxgq/Rv95chk8XbMUynCdmszmst3ooWFKPXYSYXx6sRaRVbqiiHVYC95uWv
bvEABf0LPM9VK0y2W6BvhTuYt73pr5yN3Mpk1E381DooId9GbIMraHSRgDsmF8j1FS8wFkze6UiY
n2s0Yft67O/jOCblDhqoqGyDuPZAvtYZADE8dfakE9vsQ0V2RC48WMMHkutco6p5pnvugPl0Fakg
zs8U5zFLbvDLEPNTaCBoZafLMdmCO36d0WayhaYYGJJRscqLUvvbPsrZLNIoKdnmLHOnbkefXFrx
4wWUHhKaLWrMCChV0OAIkX4cvQqnj92DCsfcpiSq4KeavB7wvCza9qeR8S9Ifp7HTU5pGB6QffMy
6NKiJ2+FP30UIpnRcF9qi0AxNzLiNHT4DeBjHJxdHmniEun0dJAKB9wjmXgN+me3u7CoJ7o3Nt6X
E9PSYb3eQOKSrlp7Ai5zD0VCIA/anqhqjjmyVggnW2OM+K6TkY2eFStHbDdZYwI20Z7mM7zALKmT
WUVZBDjIJGBDR5+9ttuQbnlLLsKzi/CY7FcmN4zXiwXFGew+4J1lGo8X68B2mu1VCc1uFfpXgMZw
b6oZv45DEn8Nc6vItKYYEy3lYMtN9KQw8XSA+n6qpq7LKSyp4TLAfwvSJmqs/S41nRTGePdaIqD7
geVTUkWkS7FIf07rsb4Lj3lX+h4KmayyceyUW5SdB5ecMcHvMjxljuLgwmfXeXF47YeK5Vlc+3vV
BcoVKQGbBFijTF5pM8atDRYLIewosunTmurWdAh/EXVEfArBnUCiB9quTiAEJCgQCnEa8hbFcFWz
/+Q5nJP6aE4ocSM4+EHYDb8Tn19q3wyva/d7DJ8saZ2HgxaXSe0LDjarv6WSwOE+8XJBtpHno0qk
Bi5USxWJpmwaZa76VinWBC11s/dQ++MsOhDa4/zOoxdv4pDIkd1SqX22NyWIJdRJnef0RfOOFXSa
7NJxcM7J1T/RTRaSm9EbfAzwTI0Jesezeondrfrf5uXEFr2jrBlxUl+h1Wy5IET4mBSLkc/TWkOT
dxnUwlVTq+QP0JtKZWxx3/IOltiIf9kliJlCmKafp5C1wB2ldMkQtPTtM50lBS8+lOVlPLxfHEPD
Dgv0IRh79HtS6j4CB47qpvp/AYJHXf/lwXNd/ZaIzubXDeU5wBz+qQn2rOef5BTYQAs4hjA9OUKO
jAPZMQBVgKTaqzrf4MXu3ixrq8Z6PVLTPhDdX7RJm7gXB9voZg5yDNdr+Msw8+nLeqnugetUyQm3
KXMNt+c9s+BeIjvNtOA36Psl4/KeCgmQc0N7QZdx9vZiOvb3E3opONPZ1RLqJpqSoTe6bZq5l3+k
Kipw5N/sHG/N2F1wdxCtEq1nsD0jO6fbZ5DKaPIh2j8+4DemetkafXk/95Qzadz6i5x+tqBrDLhw
BjTnFu4DTutov5LU4mRKpZ8EOn03IX7ly6nxG4U/kDZ91Kf5DU56k1v4mmRcnaSaNKCP5dlX0vIb
l2f9MOtk/uaQbiMzPQma+91oW6/ioI6bFKlauHRiGThaF83iWBEmuOtvYeDYAcyf/GeYuptrEDus
Epk2i/MZmsUZm0co2+8rjaxQ3SI7o+9wsfn7Xq4n8eknifTsDBcGb+UnNF3Vn2BJ8unYFr7eT29p
0Uaw/5xOgGJmCY6H+yWuxECVEysVmvSr4CBoarxu8TBZ0D03bqRKazoXEgv7zdwgG30q9tBKEfyJ
hxzaAHMaH/KMvnc2RpNQWXLkzA1SLELH3kTG7iC5VVfmSPsBHPMKx2MU4Jvvm8bwMKEY7e9UOCJi
gmn2aJjjoPYVpve1tBpUQ+crmhwQPx/EMLKTvmP5RTRxyMdsFtDG6c56hkFp+lHpInLLvxJo+klm
dGer15TxWMiOWkMfkV5O+GLTv1wQEOOX+LnOXdQXphLRvzRJJ7rbCLSZ31Kis+HmogdnRZA98Gzd
L5BeeKGLpBAh2DttUcgycCBF7ILL89HTa4bBOTzdvHRBQxnSZ6n8YKKfMJocFl7TwTYPR2W/BhkH
+SRgiyVjvYepd/gAiUhCEln7fXWkgKLkmvCeyDNYSwQ0VItMZZrHMqGW0xA4sRfHuG9di8iDrC08
MgdijvtHvU9Lz5lCbYwmkDz7C45Guq7Jn21lmBKPp9cQRP9lQ1R0q6oHLWOMRQOAsoLqtq0HeF7h
jwCgJn4vwJ+CFSh3sgHcx7UT1ldhjZmmTDXadlFFZWW/gQx5Iy9yqXtoc79PQd1Z63i2jFsapIfw
SH3UARKb2WibQUROsMwwlKULTquCUAb3oQGRDQwSOeEnCxDApaqfadFpO9PiXGSqrDWd6KwlkRvJ
OfiyTBxg9mZhdIJNVZzSahmKQzpBLO6W9w8TWpez6eWZf349zk1wBRrQGsUwehh2xeBwP+H7ovwS
Hxp5ylpTSFELkbckWpymLZJA2uMV6QwFbFcY8p9X7qdxz3ixep6iyCTKkKo2FZqnkmVDmXp/TxEK
J1uz4Ah9i2SIPjoTFoLAkNiFnJ6s5vEMdFUOHA33f+71vtHP6UwTL4cqvT49dPGWt/MI4k/MWLer
9J/IBeOhy5iUUYmXblxZDrmmWXLqGROWfFHDAJav0okLeKJuDrb6385XgDLNO335VHCHg7zBeQtw
RL2QZomFrxkzltqOd53vs0oV73rlxK9FFVCaz/RG9X9Hu58dSxFhe/WPrIFzd9/XLesZMqGxRew9
IcIi78v3XhDVZLRIa4mrOcd4jQD1nCX2eLQfQx0YOgZNqRc5I4OtuMvYlf99iiISXeGuhL81azVf
EzFzopV5DdI7ydHibrAfU+bbEkLkbFF2JDr1mxetg0dAqmqysREW+OWPRmaQVlmyPdUltTLkyAmo
o+bNdhIwo2gu6X0WMkCgKcJx8uJoV6ZIv705yDl2Qtsx+VtHfX/8sDQJVkmbyV9AGrMRY9yRfczk
+QWlFw+8NgGdcdIzxT5mjci8VVG9HeKNEvv633yELG/P3Cg0ycs/gwV8nATJSFCfwsz9CioSWc1J
wW2EzehV697ZFDBpdybRVftivz63hejH6Ky0py3oc5z0LpTXPLsK2emXbJYpiTl7s8wfbKJoRo5r
cvQtkmzhWgL8yab6oNkQAXQmg0EJif501VbM6SvMlEG5UI4N1JBJkM/nsLUAzyVy01KN6+DIme1B
F5mhc3f8YDTdOV7ieNHndpcn7pIycW2RkPyaXMskfgX8cicaBAB5QK4egenUOIz8Sifdtcjk0UYP
TKRWrSsL1y8Eh+8dhwPbfJkysWsM+wr2XZXTPIPCw2dZhSHKlraRQfu4INBhY7Cd3LRkKlqaqjRr
rIsLyI+z1GTlf/lbAqa6CicyrAmxFWp3CUMmKeVOrm+R0aiFYAUHuJAm6zQJlK079toWoymmHxwz
RMGPWbnTyS0eTgGcZooebxva61GJta0h+mYHRSGmT85/lHikl/IbmNgRB83XE9N0sAmKv3B0HetR
f3JBS8Ao/0UC52B/G2Icz4pJMS6Y1h0PZU1DVwBteaED29da2UGvnHP8fb7vrgn+KeNHIymVVTwX
gGDl4JVNp8+6oSnXG5J9j+Zbxo+k+VHejPUVrQhqkXA1t7nRUuzpYBnfjfCm7ajggOz4lT7lYGQT
88ZDOqxQ0APYoATJsfUz4lAa8obF7ohKvPHdOkqydkPh9vdGEXAuJNdtXf92Kgsb/Pxv9MEu+IBf
lhkrdseizA61YvVRnnuHGB0J7fH/8btd/Nox3ydgiYCyPmRdCeNomOVu02GRNGEAzev76sfedq1/
+RPdQ53xkYw7m7YelHBcskVvWfqkHu4UlVIwLBrSuZScSaBJaRYhoODgL6Y4O/zU4zW1a9tQWmWP
hC9WxMtTPEzdCHxvVmEM1PskeNAZ1InExmlwmqxFKfFrysuJY62dkenklOzT5SI/IdVSaU1+k3wZ
A/NifUE6825Tz80J9YJVJTmAGnSSb6Sxqk7sg7hYoLuAXU6y2oS5AEq+EWVltWEuVkidmp8ScTfW
GOlybmWxFi8kHkZ13/P/We27M3n/wWQt1+1pBF07Wlb6q9ImnOg36GsUA7U8fc+mLNQcW6Fybmdh
gLExmSzBwwSGDt0TVdpXEFAEWiCc4GoeQ9SPp8JO4XYrpiVDv4zgtq93i1GNoiJM1qxk+syEgew9
ckKnpj4jOHHjHX57pEnMle2ALPQ8KhblsLD1/20ZK6GWlXxg8qNzNG6opF7XAU5bAs1yEvO8ELBG
YajCBwYRcqM6fAZsng5dXP5bkLu7+YFmu36XxegzslpdleNWscm4UiX1Yw1N7f61CpBt51eqhD5t
Yeo0bdWkz8ahsKvV815I2X1T3AZSni0/BD946IlOkRhhht5+Y6p0DgeQfZxH4ZpEmGqlqu5gAubh
y+3LofSbQR5fuPbZy6ZwXfy8k0RQcN2sH7g2Dgw1NSJdCIuNGns9lj+ONZvUIdSlRHF4JnWb9Hws
gZmArEkSncvsHV7Yb7SlwBdtmJDZK1lip8mambTqvYMuV9W7hDstJhOF9GWmVREyxNAPKA082uv2
CzLM4xuZsZ+0iTBG8JkXIScHRLWop/2kgfxCsJD90WTbwsnBFlKxzYXaKgUJfGkKaz7Ow4bo1Xir
qVl8o5BdYLdy776Q20KYMWd7PG0WLSCaIB3g51Z92pE8XYQorCJAO3+btKJtmA4a3IC4r4TUVX2a
0MDT1wimjcwpQOLRx3tDcbVjR58j2PTn87v4Rs2dkV2Qi/5yserTtZDpii9KZEip4nnO1kkDZbC0
0E+5DQIIJPGYgkaZoZNWhqdpBVPp6XpDUdvn7fo0G9a1v5VjPOs3Z4LFxgEvobi3K9eBcfVUNOti
29ilQ28T588Z2sVRXzWzmfCUpkM08Ndtq9ces8lm5cJTkxhoGr/aXq5Xy6ypaa6HRlXOa99/7tie
rrEg6Csj519snTDqdBCH9V/7zuJKF4nmcrCTAaDJ5RbSh/g/M5GLfzMjwlwwV2WKj4CytYZji4cr
hqVGp+QCnfFUlLJn5XG1mIdzhPlWfaBonSQ/WOxGTbSJdi5ifdNVTTn7TChMCNwaiEBGNfVL43up
6loYNAALwHQSObRtuUDz3OATJYefI5Dhv3gp+iM4DciPo2TnkVK+wofedrU2DOjHcJKcVhMKNFCQ
dZU/YgxD1dj7xJfvA8Vr73aCw+A3VtfFw73XNLlzzq2zAAKbyh8yd7kz9TTRbm9XbSFilY/frGO7
uvWWjPb7wzLGh8pyhjFFB+SCrrO6rfRnnDRF8Wswhkpsfbj0w9k6wnxjbsA47eNAqcQVGZhSLMu+
cOaw+rFLArh02L1IvF2qoDm4ynEzYTxVMVvP3quahHhJqBs5SatgDZAVHVOdLqmPQ02IdTxHE7g8
0gY/D6rba3pdJLZ6fgqLLjU0HO8imwLduEBXeoVyBemScIwTrz051n07FMn1oAU0liWM9NC+GC9c
r5Y5ynbo5+4iYZ/0cawpcQZApvKJkAcIPzyCeGWVZldX+6jw/nhEoHtnExghxSKQ8sdWvEvY3dCZ
mqltB8zwjaHdESktsnyRud88AfFZa0Aw00XEtR2epDFNv97F9Nm3jhJ10Vjqpjb5CofJCwfZQH6Z
yrxxLhgxAIWyIlCPBtgoTrJf5Yr7vJdK/qfg03xxJfPX2W9d+Z3K70mjr88eElwkt004x54eaDX4
5c2LKfOvLh6N2t29vx+2OFE3p91+GdEfIrxzEM2VfeD0detQcMaB6K4qEMqNfoyHoIbM0IBNVSEp
QSySSiu3MvvEwiaF/R5JBuqVbSQvIWUjv1D6OpeRKk3JwKGtG9UyQEqBNfhFetIVFRWUgQOvzrDr
7STwtTDPEbVYZ4mzpsKycwb9bf9LKmrjQuLV3Chh1nW1AniO3cdSLQKB0TmpHpwxUYEECdFa3PhQ
xQnc1eWfxjlLCrB0ca6cSMTy0P++yBwiGYDgmEZfv04tReoZHHLgDonQiGKZg7ThA1XobmaJ10mE
q0CDH3CgOmWg4Z/k82b5H0c6Nz53/dMsYDfaaOsuFWQp5LHnY0nI9qWp5YQbi6W9uDBD1FS3FRAn
v3UojzfVj7qjF8e5CC6mqLWJ1or/6j9o+OKZXD5crwgnCs4sYknd6+geWmCJkQPMIUSOmIy6HP3s
GZBLPftw6SgSFUlbF7sCIwhsM3brTtQgwS283inK2A4k/NwOSzlVqNPVgoy2iMs4f/z2E4of97HM
ubiH3MSQmPNFI6UDGEYmFzCcGcS5ds/LtorffBsQOhmD+xZcS/QsV3PFnY89bn2bEVYE6WL1hN7h
BIBB26ODripOxbi2spAwbCjG98gyzALuro3bSBYuoJFx7h9g2BMxWrIxo/R7ubiCFXQ7zhEXg+6S
p4pEmO7d1eIN/SeHtTUs7qvz6JrcU6b3ayACStj75XfEC3/THVgMdAztkxlIO4Z86dpQfM5McqGp
S8XBLT7K54ThUDyKHO4+dV6OZC5UhIw0F2IVGk+CgBC1jtKbcbRC4355vDprlkGri2fVV6iiUnNT
P50fKoJZYzaM6hNv2N+UaDBpPcydCZz6b71IGtSNBMQYRmHQs7cy1Wa6fkCfhmp8jHQIXnClMM8h
l15RlKTWIkb4L0d6anY8bEYP6bpKsxEdQl/tOkKzEgVmRAdIO3WHyRlb/7UnmtuSqxQJskuZdLPk
nbauZTIu+qAIufDaIqmUo5x1QRwf3/LXMtv8qoexcSYUklc3jrxmBJ3MyNy3eyrLv9zKkv25ws2V
KUZxm2A8AUMb0DMTf1MIa0PDBjrmxdL2eKelMEvqfYw4iX6wPX8oal4DQx9nKFDEqtQ4a1cAoyOd
0fldMANse3/3+DwINstK+cvIbC10iSzorOqAfQMQyz+ni+8g3vm4IDx6diux7kRlGrQYkzqHOoxD
96EEocC0eQLVeWz9zlY7D9qC4/vRIpWrzFii2hYsK8GgKkEwLvmEIC1D8P8KlL8pBwLtMBVMOI3C
Iu4p+k+Md4Kti4XTHyl+ClXCP3ldf8b3wQglf4Fq8ORBoG5QAZ8wCWtbnFry4yAQWZkO2VfipIXz
aejj40NoZPpeL1ojOvd+j1m8MPzrxJf86IvYAFL2l3ugWNH+BMU80kzSp9Gov4/JMqtwqZkcS2TS
i2mBW6xILaPXENruXhFlZgH44JH/FiTVLjKIdf4lQtP3XfDSfSGP37JRLZ6slLFp1++O2QuoEoVu
6tnSeLO6yTeH3Cp6GMGNFWN7TF8ALyxS1q5KWpgRvT8+35iP3fIPYj+JV0z4YlFNF0DV2PN0LM3B
VuUb36OS7FBGHPUBPFVBQNflNZrRHwx3REzqLBq+uR77v6jJN7Q3s39VWIPflbA6ZLVEQliq5wE8
aeY5EmCS74gPnlfrfoBuNeYuJkSGo31A2wcqztM6+d/HiGPU9mP0Y2p+zRgMCTQlfKP58eE58vT/
9wNmIMbj8nqa79aq2Nh0NVPWP+SaVm2JF40T5tKYbx4UTJbg/pWkt7gHe8Nx2hOly2WqG3P8ZLlw
8Q2lznzyFro9mC54QcOWcU9C7xJuPZNasG50xrK3jOwLptNA6cNkZaZ9GpMPGTMFWy2TEM/vq0yt
uk+DOolqUv1z9MoOL9QVJc5q4rUY0EP21wXIkPKzr/8xmwim7lF9lRROvYPFelXeoSwPSmfxmO+h
NdE8FKuOj4zi1b867bRvkiWOjVb8BlPfeybSzzZWzFIHivvY6B5nlDQ2MSaHPm8b8VwZApG12qWC
wjX/ccJ4Am/t7JGPCH0MxtLm4JCKm/9mrG/0EY0KlO/OHbBKi3RbTYhKPoKEFOnGLj6fx7ek/7hi
uX4ntbrnDbPISWNJ9pbhpQvNwkPDeYHrI1PBa7oBa9562Y/sw3S+H9bniPmnHeVZz6lwuYmfZ5K/
29oR2CAYfFDwjM+kKT/Ge4zaz8RMA+qBWF5DfDUVrQd1dUcNl3GeIynd1qM4YykwBfkKp8XKPR5S
ZpnPMLCUFgCW1ZtgkspT1cfnDnKKd8gpEyBzWnzXdMjuL5brXzWbnJRaTz2VXWKkPsvWFolXfbP1
gc0FGJ98fznYXQw0JNUIzU5CYZqoI9wcPUF3M2DYgQYB5UOEWzrsV/FcWNLFXpUGg8q9E0WnHIsE
8f4K6Gp1XTCyT/V7ehlHxr5jWevZ9cew7d/9b44GeLxYa5PO68xJYdXTtMMIV/uAAYSp+a6hI8gb
q1Wcpfv0nV6tZy1UxVgdfqFAaH5mGAR7/vDLX7WY+scAlJEStoYMPgbT1fUcT3tte862QaEVqLky
uyjficYYo7P8mADuuWtAMVLloVKa1mWqeGfzRz6t2FNtAJZCzK9XK0mUNxHgVG20Mhq9eEL8PtYR
26j+GycPlWVhwtlkH7M4t0E4NQif3i/pB0sSfC2HD2bqo6dfm6mclLdszWvBIlQ0B+tGfVqoeA7K
pxD99vKSpXEOZMAVzZIz++oWXhtKA/+z33/z+MWHihsL66vY9tcEMVl2RnUhtlvjCyo9Bmm1U4ck
Cub9+kqdkDuHigGjIGgE326bflOOfFSZahjn+/AcL+kr6ziFX58dFpvpAKJeG0+yAVsRo4COrGoG
yUekaMCmleZFDCN4b3X67KjGOOjwYf0KiBJ+/D7tVctN93TXaBng5LVBNi0tUYBtnhO1HrIXGFjh
lDiuuIZ5t7OJMvCjcfuHyqLzLlYX9rV+duf57e4wvNwhHXiTY/09Pbv5b5t7HtClpmDzVRvNNn3P
OliSa7XfsRtNvFklOhSsg+0fn1hOAnoNNDGhygvNpMyHfjCzhqqbqkX3ugF68kY2lbtoa3HhL+nK
NKu8+bjlScTvA1HrRctkg01mYMblLVYgOYLlFoP7MqbNSTX4lbTZjpi3OFKnutZg26Rt3zVvNVPW
FlyftPPHQI7djlH/6yJbnVX0vnwroEkTm4fcdmBkpukW+hn1W5pd/uycTWEOIqj8P76xUFi9MT9a
W2MiRBYBpx2iacCJPVWCqD75PIBcmBW+j2jkkdDnbP9KmAIZVSxpG3z5sMqe5sUCKbhwMv8E0dhZ
N0+RIdfxA07gGXYSM5E2oy8pnOY0STLZqRzFRQWXpyWGn2vPQOWgfoh2LrLLsfHsjUWJgQEG7EgG
CpDALbm7ExhfSEsEJM0NcPlEe0qwKm9rA6W7SZXsqRb+3nQqcOMbbbo/a9Ug8Hj4HHrKiQpErn6O
HGijLjAlzeHbt7KEC5741KNBwj1rmGH6ZpWc5U7RdgR4tacQ9BpeK+00cvC/hR0Zccm/DviPsDMc
RYQuqElEd1Men4ljk7nJyDNDTTar11XejCX2GQ19+6N5heUKdqk50AbVXh8Fjh/60gUeCgbCBvmq
OeIXCI9jjT0OPIe+eCuzKj7M/djZshyk5N62+FfcRZGpLHtoC/lOt0YR4d1e/oA2PbKkufD+9FeD
6ee1YYNGlo6zspbLUW15EH0IkKA9Pxyvrj6uzYz/wedpThhsauPiFSMf7qOkI2LUkNVhGsozyCjR
0SSjOYQ975O2Byyoq34zrFDiGoETlwRfR2erKbxHTUmALdL8HQ/H+EAi01I8QkFo9qkh2iNelP90
BIGxMFX6WgoNFjiGr33mO3Rj2s0FlWBCgxKwxEp7m1eE1qOJ5ZsH2ub4PdDIO0Mn2PgstoE2xBDn
czP1xMN5AvQ4LMp4bc2ZYJNenPSyciotjwxgOcwB1/Mj2FZPERu32AUZAV2AGs3Ur2ELEJ07WqA6
omyX/L+i1+tiz6itigldq++P9VixR2o59NtT7UVZCLoqvS73oOJSZwUwwt7FzKtTejO6zumto+sF
rCYzFgt4kl7VByH66YPjSC5J01RpqgF5P+2FruichIq8WigQ9fUYo1rmOWJ+difxaTSDb8likSBe
S8uPv2eVgL8oUMya5FcoTzTV+WSeAIzf4ruMuAQDGMFRXa/RGQSscg94MOSmZHcvWeYjidwgvQgk
S/wlihEsGWb+kPOkGNL3frdvLxPuK9DQ6sxKv4qIekAaCIY9kY7o+qQgusE/Kv59/ql5czQMha1/
Cps85Yq7nofri67S6xSRkeGI92mKdrDjh95rQLk70zzK6P9E8au5Jjg2Lagn7ZMNoVIPhE2/3tOp
q1Eh7Lh4S5WDxv7xPAT0jtVHxDZfSLK414GYHHJlZgvFRMGXPQaSctzOmGMh7okh770c9lNf4pS2
49PZXeVrEZUcranFKVL9BuZbeWmefbq18aYKlsZbWRpmsm/BkzSQad5KaeDbldjW1ofFlL/ogTvm
dRnw8viE7/1aiMjlGQM4FZ/IpC34ng26fA/v3NtM8w5MuqW3HhJQDJhXC+pDekghZZwXf5cfxTei
Id4Xqr1OYcCwZc/u6btdfAAnFvujjaabx4tZf5WRUsVszYSry3JEhaIn0fsl0cZKX+6l6q8pq4EQ
3fUAsHh776sUt3fb40vOgXeflqqcwCiGjOx4elSPM1oq+H6ARtkFmG9h+gR9aNCoKBJAJXj8AwKV
cNAM/YGH0wJavZMyTF33EnBiDoz5y6U+R/KsKtcPk3UCYQnHm2kt3AErxB/55RHJdltr6h51RScK
oBI1Z1MytEtu8mc1oMSLT119vWEOYjDgD8YT8CVAOFh8XPTCXCOWNLwWh+cnQVERxwQz3xBXICQv
muaYoNXpRUf5eF2BdOUT7PX8+k/7mvkbdI4vj4nLsZbNIoshesU6uVZuQlo+rc5j1NhdtceFxPTU
l7qxyThBEZstnfvR31zQQ8vDMlb6+AWYxOHnPGuVJl/MltBjtQiQSsp1V7/FcgXU8gpFUbcaG4cc
cAkfoX3PAVR3FoIPNy+X06RfhKHRHkE07zoKXo2ny2uVWgRbU2ZwVW3415laGl3bRi7j06+FWbqJ
/LZa+OhKrBjclD93RcSpkBaX1VUHZP4NlHaTeHtn6hAYpEktKt8VuMeEHviyTYynVoJHo5FVmzmt
gZ4rpbcX+slYNAttBMiyxy6tOfZWB5SN6x37Gn3zdopNSAGc3KNqeWoncWf9llQSOEzikEl6h3Hb
wP7KGYfnZEVznd/myStdGKufDZ6N3coFycOSQ3RWzW1ykKv8JgpPKt8+11sYsO2LiYc0c5ie2PVg
1AT6LU1Le8H0yRKWFo2GaXgehZo3ZWp2jWkeNg/L4fLqYPsW82/koibFoTjUDcXAerXHLXaYBQpY
AgXy/47o4YxrRcDxkKR1SJ3gz12xjNTZ+mMnZyM3ZTk8FBXwsrWS5RJvTOZApfWDxbBl38IP3kWP
42mWWYCahwJsfYuP3oYE9Be9spQyK6XSnoNLNL5J9SjVQUQOjkJtO1EID3xa+vIX+kcQDHzCRbb+
QZ6B/Yl0u7tAa3wHPPtQyI7n2cJ2WTXELQdb7d3W86OaG/l7lHMQxX3XHeiRadEUfRleV64Xyyel
qBDzjT9Zfqw9SCziSgt8yjjEzDG4lUdNKM/rTsClPL6IIb12q87c8xBL9ZDvQSNFDFyE7iAKQ1y/
crWba8FCFIvFzgP8kS9UcqrxQ5Nyrj/2eluKJpauXXsYVjNqH4cWs9wx5uUHJ1/qnQpfEheDg90Q
D4oSPwvyce6RV39ANiKbDEkPaeUXWIYQPOZMRq5g2Kd1y4lXV9Wx5SuhZRfryFMZZLWGn7hwRbo/
W6xXOaUJL7DquWSCCnD7SdPVAj3+En0xzcElA9hN2KJQLaOCkiZx3B8jOS6APuTYEKSs0QC63wjX
hZWcqOxzxzfg7pZdVgA3pn53qVHRgkiLuPRzwAjbUr3mvVByWNkwnF/KqDbI2P00LRZWhXDLt519
A8Jh9xZGFwCr9ixqGUn8bhsVeLGaJxW6mL6q73HFlgMTJbyJ4TReo3pHJQ6n1u8vKRF6kSDYNAVn
5+bGG48m7QEKtZ14PKIhuVdRYpcqIFpQgQ5ufhfNNLq7k+IcQ+udO1EMx+Zi+ZUoN2u/L/sVG2Oe
BldGLMq5UfLSG5d3roPlwJhxVw6iYB0C8wHqARye4JuS/CIuTrNTVLG2wKBTz72OjebPJc2BowMw
ybxsa1mPJqwKN48OBF5US0HZ349obF3rCnc6Z/ExIQPUJp0dAW4L7ypPBBTfbQKOaXp4xGcRuqmq
qPOXqBqPwLnViMD1FVCieXvWMLn8GKmvFMdoiFI+lwCxLmwYj/S8JoUDt/cMz7/9wJTfrHvCXa9K
BAKaAdK5eGOwhvo6jE0B+jctPKzeLROaYaRvkYwLncQxSpNKRruBuc5qCSwreT7OkCXpbxm4ulUL
8XD92X0H9/2NjiLCTtrPjcCYPEnLPXHd1vR9HUrc/PNk3DtkHjScvPiPLGXUkOJRmiNyxJryFufu
HEvP9rvwm32X3cwxaBklhj1iW+DFMHpvzz2Xm7pLL9EUAFM1Vb141feYHLsiWw1c1XVhR3WW5rX/
QEzjtizNh37LLjSclk5vWtrJP9n4qUitZyyvvbdUyhxQEkfJQqaDhLo2eVjHOH3nCnXxkD5SDT/Z
ZYNwIv67SXGcdbrp1UK7b1VlucqrzzZdVEPQ3tZJcWIrRM1JqDk3SyWqtqFLxPC8NBlYlUZoGltP
Cq/VkJgkgz/xVx8xvOeQUrtl0astgm4jIgBP2K078InKjvpZtKlZFD0fc4AiAE8L9qETITrJOFgu
y9sw3Q9fmS9f1SOnyovozO51i4jX2CUwcYUilR6OeveeUVTBOlIsxvLR9XRXxMeEpaWsg8ougEbd
AdWtlhMqMsR2LvkPzPKWtLBwcMNTD5s6nmw8L2Pe/5mRYH0Egfp5Em9XK+NL6lPUvOg9I5rU3tgB
REjwGlQoqoDbz8wSJlr/7zHR7/XuAnvLEnsDtPa7fWSnSOgbKYceAI7q+w1VfkXBp+EM9YApmMkM
FhsEHcpvQEoz6t4xV9TIeVnqP5V9eijeJIQbvAt2MY4SqHgJZjzGChf4MrELfioS959ISVaaOVsz
AVRYjdrHzjTEeHGAmhiSHja3gNPBYsh0Em9lFgWjKk1Xind0MB7y2YjzRa9NslmFSYSgG5iVmdIB
M3etebkc0J+6jxIGO5RmwuL0t5T3mPjqKQOxr97F+bKms3lXxGcITBCbj2o01sdLlMBgZZNss/PT
jOei+fUqWAeALXtqK7ohSTLayML5k9pjvJxUBe915d93HrvGC/wYgCt2OlVIr1cJMOlXF47OsOPq
hiXm1GwnLDs+b5y2M0xJgq/Gnq5wDtzXnzyK8zs3ZPn2/H0i/7LWAtt7nUQOK+447nYhjm/4uK42
AFzOhD70pIQF4fpUOI2DKo1Gq09IhoByuIKRt/YNgXc4mgr61iUta2JWwK/YRmg6Ibbdbv5IB7SY
PQ9vxwTcazoOW5ib/g4tgOTTqTzgdg+vpwW106eY9JxTK0nx5GuTU1v/Aw6HiBXVl6oJa4nPpTi9
GEOijfPhI2Q/ByYHj9KKPLBCUdiXS9rSOllCQpkRzxu5Qh4kcMjlu9TFP+ymsanmDDS3xYTedEZ5
6TK/8072SG4qcYGDeAnOD1mKSAiSqbZW3Vohsy42JEy8/bd+BMoqR1VnXhk8SmzWRZ2aU7cP26cT
AGGg/xr+9vNUNiU5hilcooAVPZLr+fyzmWo7R38g958NP7I+NcBWvm74DqZLEo26UiKK4j5GfDPY
2zjt/2BFP3DmalCVpdWTtB3w6gVmXll5AAtMljXKQ5x3EuvZmNEfMr4m68OWyg/Hu9X2FtciojDS
GQRF/7XQ1+1EpgORet/aMGsSh1rNcHW1qqyFAviupPMcPdDuISHOVuEj6wvrehWr1knWDouffiau
5Tmy7ClHpG7ch3FxcteZvw4c6oDIY2Gx3e1skvrubeE7Bb5Kl+PgmPS1NijM4SFhLfUR2m80FWYk
cMkP/a//bX0e90eXpdCclpxHn521CrltGrDiuJ0vw+sO1mJF1JkWrmBFh9IzW7oPJovdXNagXRbI
t8rqWvlFMfq77QQRrB1n8/ahYmHU3Dagi+nzyIwsAntmDOIIrUNgCHfiEmCKHt0Jp0IEc1u7kO76
rXKomrmZ54k+myt5WDcqvQPrycGq6R1b7hvdK6l8plZ0PYzcfgroIiByukYH1ct6PRsdaYpYBcP4
lzLadgMoE7VNEINZFD350UyoSNDWtgDDMFFRxNC3qiuQORsHbzqKCEMwvz8K2jr07FMhGRuOvCM2
gMXWjLS+tGnsp/Kiw/FI8gMntCGkTlVAyqzdTaplwTZiRrpIJqYiQnhEdk734IG/N2YsBfshttX/
eIFZIhamh0IJMmpLSYLUi8NlZwFGrVH3n00FiWMgp6h/0ikxSmTduu+nw3OVzAAgYjD3OOlgR9LI
yGumm37DZ5k2uQ5KfGvRyZS+Vxun8JbOqtBkPhyT14VCL1UiHPqnwv31C9ZQb3GFePMJpCAtq1oI
GiiylPHM4VBlDYpnPa193a6aMytaEKOKSvdnlSyFz3GG6GxGd6RNowGTsMyG48MxWYl/ce0FMc9i
x/sQnUh6wiwM8Zdsb4+R8q3cw2MABFxzr+NX23OsBB2v+0Vw/9r9n1ECXo6U8l4i/m+lt4jvm2k6
wjUndWRkdcX5+dcJ66lin8RjHa9ZjaOaK0LERRn5j070Qj81raOLhBtVA7qdZXet2akPxJFiz51j
ySyfJCqdkxvTXGc54jQwhtfK/G5LYFmmt1pQ3OOWQs2dv/dAvvX3Nh3MNRPbxfND5lN9RBmaO070
MBKQzKhEO/8unGsRFYtC8cFgL9TerJtuHh7yMgW3MZUMYHHsGTZ1jxXQIswObdR48s9rSV8QNYWj
OojpeGnCDQ7FNNaWFOj6ZvOU3eBYXabzbV6w1ve9LH+vP4f/pMBaGQ6R6ugwh9QK3TAr9ADKvEDm
esHG67o2DxMf/qSHL04Xnp2Iui7KfuZklvliMjqCiubSyKyLMxOFDq9kLPsjrhpo7SgXTFK5k57N
O8UYMrBRU7ILaZXmk7tF33mj/o9ZWHbvGxnWk7xGxwHkXiIP2YxHRqqK5MWMA6Agb3tmo4oLWDBM
OmmvleKarxExrAxQsuCwFCI+K7x9NFePsRwgav/tI8tDmbRKjqUajCM3ovceBW37qmMOoV+TA0Iu
qzeILRIdb1SU4yqqQDykN77Zaokh+Krrmr4l4ifwAdcfUiqqEuEXnu6m2ZL2FhIbpnPqVLRnCsI5
RPLBDQtzl/GJsVUU9dihwlSAZ/GChOwWTZp6Ysw7AJvtdLFXTpfFAItD4OVprMmcf8V/vhBfq7Of
7PlpuYhHcCGJiLDCM+RQ02GN3kr09dNhb2CqR7w+Uh5zCPUraEMTxpOQh2yHdyxd5bDGtrhZYs07
86F2RaPbQATl1Nh4QAwiQEQojJ9OCm+F6BxLViGOv1rl5jSWw0zsrP3E8nBRBIJRqYxbtFCFoi07
C3sxTeTMzorrQtTDi36UoE7OQEjWhTd+mCxC9Yz1W2FIMU3Ah0w6UaZxiwcIGobFeJe3i1344GxX
Ga5nWNpKRRO4YLj3G4cw2gCk7W84A8HBxaC2FrAV3CS0B8EA5yiS4NKU+kCgypLST+mu825Eb7IY
e3f7CTnj4qxo5mbVJb+lk0mSnrUmMEJfPv1UQU/iQ9snyEejbr9tjuQqv6mEOdViVgcbOzGax3Ht
G9RmvU54uiZasduETg1yOoh/9u2voRSLE9qdrhY2mfIq2dR8gsKKtC0uxN3PnVfSYSpv56rmxkHm
u3u7i9/Lt7bWK8IYaRlOqoZUFFxAUcLG5Wvi4zmTQg7Qgn9m+ef63/l63P7CrFoyOBvMszO1oP2v
5iKz/13eTABaXMYfx0/jzlqVXcSN7DOAWPGebaxScqCjC+5VLd7Mxuv7xNZNLrrZ6TpJTNWnsg1L
DCJcIykhqK4B4jh0sJIJHP/Ew57oJvEa1h5sNnHxM1Rv1c0UdzyXQhyyrpRnKtK6BgF49izlqBsV
ySzvhg1LmKqxm7fovTbm56FJ7jRxztu5h22QObDvfSgzFSeWnJFf39FToPUq1U/5u/pTHwXJgUB4
Mrr7D0o5JuA4AhHr4IEB0+lQkRiZTuPTHxamW3SqwFCjJzx0ICC2SpHNpYt69WiqP6c/5MwDDhni
FuYGpV4sKT2O9YkVWPWRYUJUAcuCTdGRgesGNIvZEbi/cqCOwicwTQiNj6LStHIRkbWnuYRUr4qP
WDorbGKTJjX5o1I2IJgU042jjHlsg6eSJSkdzOWw3mRm46BEp2hX7NcmS9dflBYFIGj+70K4Wp4w
K2zUR+bA7fkBafqvcyEV74t/FcUnv8X3Liw7uZXgQ4bAhaZNf5FyTnZYoH1dzdxRn+gi8m2EtxeF
JrBzCpw7vlMoG87hNBmt1Hex+wyDHO6THDn9/BWnLpaSQnigmW7wDQoAtI0oP3SeuFt3K/XDJqgr
kC9rrpYPiUkm79ytSDQRxx0uZxDvsbXtkR1ksiWNjTM1YFlijxswVh+w8vT7aJXin5Q2FYPqjCDP
6ybhkptARtDPkrNC9KMc5ls73ujOpuHBrsTWqh74mrD2pRsaVbH+P9RF1wPTb+ksiykFe24sjeD8
3yS28VPhPCULUfHfgiPF3ivf0eHcqIzRL39pENx8Nu0bEXRP2dQgAQq+1zAHjSl3M55IBEoulEaJ
70wCgTlgcXY5iJNk6I/slP2m/PghlHPRLwXJr7AYR9SYR8aoOdvAC2BIuc3MUOvmU/12OLNiuZHH
wxSkOu1gsuVFSrXIhbMDmYx/feqSbEfGE93+WtAGLtmrPMrnbYg2nGwJ2o1RVdihENUXh/slTVVg
TtM4cH00dQYcf0lEUPt0JZdJ7VgwkSyRZhtklxZ6fizZHJFIkaT9I4U6dE7XMsqU8EEAgbSuNAgY
q3gjaNR2XkgcqVx8frx8TDoHSQTroqB1R8f87pYsvV3yIU/s7mXkXybpf/J/q9MUudkaaha/7Zit
fU6NSeK/uO4kOHO3Z/20f9airZkYL/zCryFKNy1dVvjHuUn1DOM3dOwgivqrxIqCCgZKyxQK8h4c
6krBqGGQnscsfwRfDNnwSwOd8DHhGbUIQO1PGb/FzaD2cUMXKOkMUiTeVPRqdI7+RQmi3cG61K8G
Hz/zUQjeg0VE/KDAqH/5LJRMvUBhxT4/q4iiGhmJrp9ivRvT9SBNq3KEdQyi9xRuuc74bSJDTY52
KeMXw+wPnhtE9NipfrLKmN7c2dGx+/RrUEq9YTfiiGpkdk0gpqC1bSbxnY8F8uGm5Iz6Ck0QA97l
0uZsLZRpVIvVISmfhY0n2GeM2JyqG2ICsY+oWtRi6ToZJNWYicM5XXcHMS3gM9eXmfuyUqdcSWq0
LnCKnlcu+4qD6nKFotjpYdta0lGFy+vEq8wOpFHa5/sw7ZJ1HFCqHVs/3WzPYFl8GYbQRtFFj7d4
xov0nN4VChgHsKlAid1CAaBxoQjWaeiOLvHLw96ix7ojeHPOJKr3gXm86xCNLeKKdgidAPdTXJ/W
3FUzue677IBjCdXM8a/g3NijzPF+YBGZPke7ZRfAYtBM9nFPaLxHCmEzFPsLSWN7s8pSLgkoSlBz
uEgHj0JbTiGsWpmmeE79e4tdCVqM3WMnpr+jQkeUGQEWJcWlJsA6DxaNNhzh7RFYFkS151zCeR9q
b4kEMXUli8nHRjpVfyy+nSUboac6hZmTnWYEq4Y/YpjaovY1IRY8HGPW04hJwdvpehzXERllVeaK
xQkgVpo/XiAqXAI36fUe4IcIE3dq8qxw81u4opRCSB1vRsqQWRjUbNBIJ6ZikLgT5R4HKAZaQ7wG
pHv2Q6Z53P0AQ65zza3tO1VFcIFEpeHZT18TJ/gwQah4mR/wDGSSEH1DBQHNuRpGz8FootFamF4I
IO9JWsHTFJr5QZBBDUZDDtdX9GvCqbXC5+rlw91+gP8Qey4YoIL6oX9zmZcV6JLyoXpnZZoCc6Pp
ZSTDtWcGkGhL7IEEyy1RJud32w8YLpCV6YQMjVpaj83l/9icMHPtJLbg2B6kQh90h98yNI+5cuSv
HcgSuNBuHwpWfQFuQmYm4fKJ6X5z09FNEED9TDHrkZ5SdDU9cJcpd94kV+W3mNAjKaSH2CiN8eRC
tzeX52M5C/FNNRq6ruTDNy6RVVK9mJP4Iotb1uJkKf3cHilw55/GJVjaMnFo9nfUlwzk23VB+p5L
L0JfePc612L6qzoVgVHoi1xKTA1cQFyuk9Bcs/EfAtbc/ejj0IFG/6QtUObyk/IcTL5holIFbP/C
tKfVwrk2hfOeejfTBxu+6TKcS58IJ+lb/pPzxuzjQKhp5jQM8mf4XWhw6jJKq1pHix1vo/L9ifrl
yqFUsR51ogzCeqegDEZ3YfnvIEa2GFy7IYvVOcDcbQY1IOpUQTEgeV4+r+XK5xCJUV4BrDYnsAZn
0WKgE4kILxVPYF6EiVHL69UUgdKV0V+WCpCuSRP47uVPu4hwivqaj0FPfjltefG5hKr8QDS/ZlPQ
0Bbv3iAJ4Li4TmCmMj8+6L/xyEdc+6vqLlOdTfU4KMWwD+CAIHRk8DRa1Hp9Puapc1rSqFDlNgp2
4sf4dYdArBZSPTWJ7yLJTOL9Zrxr8m0wBO+eRIYPQFxnuc9KeKwI2Pd/98oOfzhPfREhDkgZGgeG
q0ehTpYYiJSspjnJP4sTVh5CHeLZ42KPKos2864T173U2ExMyGVGW/Svb7dyNeOy10jhKLLWFv/o
Lr0QuxPCSqPXTZXRibMRMp9spi53xYhXu5EOlYRq0FwKCM2z62y1jJEmHxUqggXHbL50gJPnVgdz
TkDaHax+QyklMw5UKW7wu32fmcUr1Ann0nEIVubh7ZqngRKekLKLhSNntAynm6mrwNzBOsx8/BKP
qTuHA/tS3S76Rin4kzee8U94IiMlf6LUk2P/jQwrVMxjgNEekuBkWVitwCvLX5M/GS0gVdPDuMSd
rOPytxB4PI07bZqJWGImFk4mfBXka3iQuEbFl0lTvBKHBYLxxq02B1ALTxXFrTRONY6yf+RrUpXl
CgKaqY3hcmRsI0mc32Gxaxpsg6vZarSkuUiwQvDoA08IJ/MfTlfjTTRST4HfegRLsphqeQ9lEhSA
R2OFeOJ8UyYyQe9z/1fGVZv6QrqV1i/6EmWAd6EW40uD1oBdhgt+SdZEGHapFBC9CYQ2F7g6hFtW
RStHMwf9OkhnCKNBdmojSuNJ39K3JvN4UhSq84PrrvBlSyXDk+ikfbA35sb1+d/vjJ96KsV27zuV
2zTVBuQEwzN9p6MtfSSrQSMmcldmVZ3PsY2NyKN9FisSNl/zksutWEGIAhAgfAXwYZE/+cNVP1hY
Oz1iwgr5pm7PJupPiurvLsqXN2IGp+giCwWEGxkqjbmUtFNncnuAnCh0aKRjkfMdtoe/xfgpOFQn
RvzrvVkPafvTpXx9U2u3YjcJKabbcNdhyz+yOHL08u065L5HRQ6EBBuw5s1XcdAaIY7QTfMPpwoT
NTFyIoosm0EnWbamMpDHoV5Ssl5wbQKoAjDUdASUuWTiXlHD9J1yuZd81spisbjg34Lachc7pgS+
+ME7guv72XJbo5DxXUa0c91T3j0Ud3Fe5Vfou/phJ608PDlx6B3Qq1OuKyrBl1gHBlj1e5NLTHDu
a5THLPc/7ziaayavCrhhG63CU7DnRGNAKrs0bR+Sv1C5mECGxSgr4YUQvd0BaATCm+VK9w3AhyHL
VN5FrBNO5rFWNn7wl6Nji1PEnTGgB+9c/3AqrvIZUp3K46xp28FAjkCLZ3JIXGs9g7B4G3iZxTos
EyzGQwKQ71VSRNhK3gsOhPCH8S1eu89qdHXreTAOhDm5bvVsznr7ed2bc1MIHgswiE/7yJAFVrNG
S8Qa5mNDsYoz6pTOb8a5dbdrXSPCH2Kq6ngqlMw/fY1K/N10E9Qf1ciut/DQczQeHRi00jjMsHl4
EkSa1hiEZVa4FqkDFCAKhJmcgcp2NphnuTczVFgTKmwS99aGW/K6DDz2zEYQXxpcs5vBqHnhzKnU
NBCSoePcNlxc6QORBFJAztS09sVJgJGAUG5z7XCQtm4y3pZ7Y0aK8yTOh5EGspZMRbetcSNJazgq
T5WHb28tDH4KoLaDBnrF94yXt5jl66Pv1kjzXQ1kG5pEI2Mycd7HohrY72J8nQDZoL/6IlCpiF/o
3rOHEn4w4J/4aIaZxpZlTkSMnN9VsfpVMWtH7s9hNjJIpYcOVDut6G4a/3yMb9JDHzFGONufab7N
RGnVGFqg8aeKwb4mOdlj7yzpWVz6gpGfvYuZ1EHLw7YZrtqcQ+thHqqF8kNWcmcan0l5to8958fi
FIOtHlzU2CwoUWHGNWJGpsq4sRoVYLDh+Paw0zYBT5nxp3v+y0JYrBtBM5IvtbE39qNvOYZM0iM2
4vGzXSG+Hh+8hMLBi6MptKIineZOAIGPTYWr8GSRsGUNiJK//jbsco1LYpBzFudIZkGg5JINi/R/
0QnkBIydG7oPDqAL7R1BNUfYmwbxToS3m3CbYQn89cv9SP3fBmFMGShWlBb1im+usvROgxb1+wUb
17yP/De+MBMxN53zo5CXxs/WlNt2S0yQ63uw7mIF5ZqY0bHmJRwGyEP9/Nfyjto3XBRvB25xqXwu
5ny8QgwMU+l8Uw0SY2W2Rq+2meNt9C0nFWiswLNbyaW3XXjYuxxLxkVhvwOWlJDOsj8E3po8CRnt
SJTpHBQcuOeFvzXp3vQMCIffr8yZxAD5396EF/6e/cx0bSmqL28DFmmI3GHG+8y61lcw7JmEosRd
by/ORiLAOvh7Sa/7V5T+llfHppvt/PHqlhsF4BXOUpxp5m55v7+Lwh4Se+yJ4/e26uKat5AEmY6N
kGFFOuc/uZdsagnvVW8jTFJpe38Fz9ZwsCkpEMSHy+CF28lkm8SO0Q+q+QdofBF+N0y8+bny9+96
EjEo/bFUbkCg0OcFTeAfjpYceFeva8LiVQK6VQRTbsWvEzP8LvevlFuVbmYpqYc/b5Vb9n/csknf
zDTD6FRNhxAJLwxOfm5WCE+/IlPJNy1xYXe6UedtRLg+47LYG/377nJ61mDSZN/vUu1rhFtXWORR
0K9MOaIT1X+nghR8x89oLQ0X1dU4pBUA0Ssl7NQRQTQrQL8qdguZvpeZHMKA5HndaCO+lO5TvpP8
2Z4zCAX3EJ45kL0Bml9sNIX4NjTuIeH9ZrefPAqSUuUG1Tk8y1q43wGsLBOmA5RcMVDQejCMv0be
q+XEk34887DDq0Ku4shzIlnZgLPcscoZErUYGeRZLZYslmIp1myZUWKuaCWilSS8tZhYQ0e7LaIL
aNfeB2iknVwZHIbWeJ1MfYctvE3jlc7vg5ymXtRQcJKscQCRGmxk18WN5Mw3b2zdeUUpQhFUpmJI
CFHyADFi/ZF8nwknWH4HcKh7dK21MNnE+d6eW2nyqbMnVx2RKc3zFNmcUTUxjVtwFuR6gFR/5aSj
v6KNfdwDDuClbkffRBBP9v7waZbaVWjUPVYZE1yHjfaopJkjU0JrCsmtUirhoG0EFZZygb38yYbV
wpS8dklco2c/qJM7JwFrtgAOe/cZSvnalmzITfxIBTrcWQjx51hE1u/byCGqxpIJx1IdIQmio5SZ
uxSer1VZkzNaKiMzgoMy0gHoCo8/4EBkOSeMOiSvxxPrGHwJYXNMrDuKZ/lc1PkwSouH3U24D+jU
KjvqJJwy7xRoXlE/cpfqCMZPCIFsvSzGr6YImt0J3aVlcNV2BNccorbkvciFTVb8BjxU2HON2N9I
/hC9R7IvGBVqXd6ISA77ZPDwtPu2WQskEJJ85dYisLmJnvSfQQ4G7l5YX53Rd3dDVwuArFvcIm9S
KDVxgJ8oZtwVsPewEDFcjznO2xPnms4ivMFLxuX2GEdA0aIoKOK0vwKOv5gXRqv52VNSNOJKG29x
NQUibM8ESirIk/7E/T67lt82/MjvZsaVVI2q32NPqmMRuNWeG4g3p6PpEKuaypmDjotBn4SN/u9Z
UoMz/wiGUb+Ax+0UJrQElyf/XzhZdOHgJFUTT9VDhqZtsyAQ8t14rnDn3dFv5N1mDHCEiF/dy501
Gf2k5MxGMhW7CEewhh5pVh5Ob+fpyTtFIW3MhjabscRy5to6D0nwWZL5SkkPgl8+qpD9xwQqqPU0
q8C+N124cWpH1hA2dXhXWFZ3ODAbk9gLITnkZs6mL1Oxj/Q9SyFUIOxDRIJ4jeIAsVapGagW+fPX
MNyPAQdNaVx+lVSGYZ0zp19MevME1Ixn6daoJnigAYWwhsqD9t8JpJpb2I9jGxexOATZngqDPE/i
RjMDuTvUkGlqqTXOwzQy+wKKvDGdEiwqM2ofGqFdZNrzbOgIIvtVUS7rqH71qSX3kUekIZ3u9eqP
7Tjvex3nqX9m73DsDwOEQfea7wpVc3lR1nkqrXfeHk0XA6j9gnMVFqdtqbiUs9LYJ7vVw78RUXzG
bPcOY1D2xMFPXLyynLimlvFGaSLInMHXbIXkN44lsLsolV2oFiZLEbWF75j3TxQjJGebNa3VTpXy
hqa5u9iq8mWHqGDxJRttAHnR29lXG6cYeEDkkISfmyEDruLhrCr/gOp/LjcrW1nYQHJMKgXD7SGx
0lOq2EYtOzi4RYc5U/fAEy25KMYOhBTcIcW11z2pZd2LOXGghuZcMoR8CBiexNLZxGmgQlIGIjzU
7ALhHPUgll2bhzE0BYLe6LxB73ffpxsEFS9yU+6xx7rZf8o9kpgdJo1dOkPNuMkUsFsgInaC6q/L
yI6ZUhPGHSshx9gcWZTE53iAV+ATzcdJz1aaxU0x+yvTSSu0E2RGsRff0Do3D9i7jlWJZPtcWbGI
22c/en+pq7ctKjAEWqDd71n78JbPdx2Ej1HxGgSmKiNR3Gsh7SE0CPeAPiIXr2rwq2zxKxINeMAV
DD/B6yVuCoBSlaIuO39fUsqE03GTEY+nzxNVK9TGH0/KmH7ip1zLTX4bypBNIwNP5Kf0c2afi2xH
4Xi6B35mT3/IT1GwH4uPE0UUcD+6AlUPDcn0NIZTJinh3GS+7LFCOSnireZhjRVooRIqpbWOM5Vz
hD2wS5GdwRV3Wk+3L6Rs6a1N2STkRPvKvNOcxaXH9ao1S+jQ1jRGmTj3WRRjhOsExwOZbJ551Grj
dry8Zddiep6/eAWtC4J6pqaLS7is1TLHcp4wknZqDLtIe3bOw4zs6ArCTMAzrfx4TzNGK+MsADjf
/GhfVv3dMnh1HK2Jx/HEmpP03Em0wQtnUxB0xeGWH8gXuRSzE/PovF86BVpaOAaxpG87wcwkHC+V
CXRxDH/W5W48m3S/Pv3mi9dTW3DE+jbK5lslCSV+VqyTA4svmKRvJ58yh0vd04fvKHrMzhS+aodM
u3yJ/13z9ZNdv3wA8S5qYGv79E0u63F7HtKtNj/BIkmMl7JShnrhXfDtuVFH7bxwFg9bhR4Inv6L
hCdj98vOxlm8G+0nJLmo6m2Sy+GL5YZFaj6VjibaqxFriGjIbM/Xxwno1jVDQZx8M7BRwL4QWWoW
GIJtCV2yL8KhXSSGvG7c9P7F+5xtvwvXJXBVUrzHDjyMixa074Ub+4va5FijqIp/IG5LVxfFtziN
JB8hhRYQb6cFK4mZCwjF31lNK1oqK6zxN0jZ3NaytC1ea2nTHNPVj8ASS20SsFXaiuySZ0t2WoaH
OkN700IT9bHzA7pUctO9wF1set6Fv0sCZXqgorEK82HurBFh7bZfO9RSEay1G8DpS3GoN/45VcT0
40qPTLPAaLaWwquzFgxtU6rMD+jWRqpJNccxDuKdVtJ+fnfNVZ9GiwAf0Nc4DJZVy6PAs1sunikD
louTP18FQ6r1fA3qXIqArN3sdR+6BpK7QpJBDDRcedLYHAFoyipoCk3t8+BmPuUYe/0MD21K8kNH
8jU3msFHLGV4vP26U1Fs+gDJUrMkGynkLO+PrqWVhw7GTAGFSZbYfz6St9hhwV6ODt7sFqlLz7hM
VAiZCyn5JIHp1HL6Q1HOt5NrjPTdXxYtyZ3sPuFxpcQzL7olhNO0xmhUJ/ZGs/mTu7e15jf6kUra
crpCHQpZPgRqb9JGFJ6xlYbhpwE/Ujsk+eH+kxIQAFhEwX9+L3GyxU9ArpILgV7pjtDw7OUW5qE9
SPPZksSnzaEP72X3oYWaMaLzeda7OloOUy3WwY4gjaLmTTWAMmevswDN0Ftas1Ik3J5XeEBn04pH
tezk0y26fXuvnXOaz6VFZElJ7KgYtykn3bHDR3wVMP8wOLqfbjEJ6o8N64sDywTd0Q4nzgcroSeZ
XHn4Jlx78MKTazuW8B52Zln+iqXfkyCMItdx2mufIOMHjc5CotcTeTMZbiDPIFW9rDeIP5CR4oZO
O7UlTWBeia6DGB2MVmJjpg3xTaQuzEaeNXQaSTJRQ1R7MIXMHpNleUmdQmkI+mD03rSIrjJ7lixv
VBWRCtR3BlhvgftwLLEiSkFvxaKbccNXh4tVircNT+qd+mZ8alF6XZFLcGOOCxX0MRVN0W79ws7I
UfE/9NTp5fPUal2+lzimHjFVI4oSUpMb05+2P/oR8ph0vppbotwi3dV3DjFFgQXvAtKah3gHARZP
Zj4+DqK0CUKUmS0I3sOW5Y/md2E5znrNYRhk0Lx7E2sORH1k3e83gmJZVytEq9WypzCvN6FWqpAN
T5o1RKoNoyeyIxx1l/++X0x8+50tJS4Sasc5nUVxCwZvfMc64G9YuucrFxWen+XA39tYRF8qr0cw
FEVpQXFhKMldmO1BlvFISgUWD3VkzJ1bQUR+QIV5OydHoVoMI7Yfx9u6tLZl2AieDlv6oaqf7z7N
bgXT2BvFpQ6EzbnOPWZ8xYEyhsz8UyNByreWTuFsprlw8cyPoXs4wywoYT7BJNBU1OH7tmNEJO2r
re7e4mv/fLGnI6Gk9vZhZWdyVw6dIXC7FRIFDa/lK50kDGP0iaX2nSl1m4CGxNvA3QCLg8Aiz+6x
33/94DldWx84TmD+QjWlvo7cunJTbvrcQycpseCeG0wn+jiPm2+4poEKkvZ+TU6FrbXQE6gx599K
wuavmZJAdM9mZ6a5cc9MLZOgTXQe11LwstpWPWxhNuG4GCxGzSnfTA7VbJCWzE+Tg1MP+TI2NMzh
4OXZQBb47t0M3n7GBEcXmgH46StbDHce839mVAIDbzYw3zBExLpsf2JNj2u5nsKabL2VVlVyB5ns
Wh1E7oJxeU7088ovgHVny3/nOYltoyImq40uDveFGqS0T0TOYifkU2gKpo55tbC5uFvHIfsG8SrH
cnfoRorui/UaN/+49Vy7noHb7sK19lzKVHBsn1EX/q8jkiv/4X4F8Da1+418/FItR80+1R3NKxJY
IS+Op1c2I0u8ddUaS0wPQQOmuMedvfnyLGpGcc1KcpOjYlkvwzBp91O7y24jZCcIxuY/eNsHVlFc
9Zqw4H/XvRQ6zVc16i7hddXDMaARudASsuDwuLdKkUR+3dWmY0piqj5QEfx9yO+EG2zIYchcxEfl
/btY33ifUCXKrp8ws9utuEV2C8OM7EGaZNiAhK6cApsSBRbRPicn4ho3wXMIrHzYETC005jbNz0Q
mZBSFPw6LZUIEXQWW2fNiEcVFpQsuoRZE95639H5wV2fKK8Zl6WHY+uWiO+jT30zQA4jwNV4h6pl
xFWPus4w9r5M3VCwJRZV3D7wnDMSRz2xODJIs2uf/uDBeab7f6ELEfdT7tsPPeguJpIa+MHeeeL1
9bmTleG624frDqJAL436pI06XtrgXB2ZxyvIgKQYcDKg5xpLgGBTvZAGDR0SZBKiKLcDruggZSdi
X/cdXinSAoHLIpLBspya+7Du5ZqQg0i0vPlTdExJsRx5VDi0vbBgeeHFrIUznw4R0r1laYqTa0hT
P39QqT6QWBV490TvFlBbPidJZENanm5sgpmjajouMaIHWYlGyD3AtzJX2xvn0wQo1dYBnuhfl72C
wVJQKQgOzefih2ctA3SJ06bc4vTlCbAlERBscnufEQ7L7mewEvJApieE7lITE34OZmxEUekqkGtT
HvHpEyhnn/ExcDM9zi8FPeshUq2iLCUMrVzc7JHpcAOUsd8ODQ5V+wJC7lZbRv4cLIwRBsqh7PDr
78yt8wtDCkEQHchdHIztAUrr4u7sZjewBI/hPwVLhHdY1rEEv8h0D8HnpqjDvn8LpUNC7fSxmsw0
/tfREFnbKvfGCaE2VlpOB+Oyw3v5MRl8Q66qZGTHnnkopMSZlqrwrMyjc6ZiigCULBbWC4wojb6Z
wousM4ARB/M5ci+WtL5dR2WE/FI7Z2s5zEJtlI0tDU+1qm82wtESfet2mGj7i1FyTZuoRJIOnt/X
w6Hd2j1YkIhPpBx9FSytmGDWn0c6dHaG9achOhPgUvgRGell7VR7wYTLxO8Uquq1Zv3jq1JZmvu9
KWzhc28nJFvqoxgYaRgos8MCc+gwMnGfD/UojN20wvV5xB8J4x+1r+X1zdcbTL8VmBZP6hEF5Aqm
sxiyEEGUNwtdxDA1iLaOyATf76n28O1773j4YdJJSoFotGL2KWT8dzbcMRW+dHYti8e7RZ7Qisy+
6jfTwucrPwGmh0Z/GWSDPX5Ix/t3XnKV/e8BUyeOnh2CU7enGUnfLhyPYCacDS3yLeZWTOCbqCKZ
eXztzpzsRXSmYaK6TFIgJuBkb8SctrIGPfPqdicEZR0joehnPBiGWuPBMyS6EhkbWLIHXUyL0txl
xC7sziwX4mO0k3n5nTjv9VFM3OgyeQ73xb23rFJuuoKmqsaqsoe5IWY/GNcKTUWXOFmBsoDvRj7f
tP7EYzWM0nWLkC1kOIJqOHU9qSorsxu/g7DvZOkRIuIrk8bh1oSgIY1SkUVHbH5x/W+GD7IA/IGa
UVuqor9N2NocR3NUQp7kY0pV4EPC+mZPgQxJq9d/YwvP3qMU1tqwBJkcPGV9PZoVaDW2PgovFix/
rZ3vARP66xFH+mOTT23GO4vhqLnuOv3imbkd0hVi8u2TVbgF/kIB++3lW33/jgyrPHBND4Fji5Sg
CIrFhF3DmekCKP8pKk3ScFYd0HASIsMf3z/gWqhhX3t/8RrxjJ0wArsN3JaMgkKlxP/n2GpNR4EB
71dmEKXWq7VML2Sio6q5YxQwb3lRNN4VftpTL0deJVNhDPEp2TFm+lJn4DMAH6usLLNhyChFlRbK
kwGuDzuK0PHyOXSHE2GqmHrFShiPxpTHnsq14ZYN9fxIcM6KedVLwOHcEKsvZQVNP2M3VUQeMsie
0GoErWUIkLtynOiPtYnoozf1jYAao9GzcDBdI/HMLw5fQtzB7BzgHkTiNUiz2ZlCN6NS7oKv2I3Z
mLIkfwgHDpKPO+7Ss4D8c/MDuC34kY2ucdQbJ2diCFBJKEc4gP38vDaGPev4P43zKVmmhBTVbubK
kEkO2IPLt0SHH+F62XLeM5K7UrBke7ayxzm8K7C3Y6DCPQ+oc6DJ/acINkIB3KYq4liX3jFZhWX9
fHhNCec3tz1dCwgDeGVZDYktF0qBimfDtpOQp1k7YenFCcESSoNAx9YTY4zdAaz/dX4wXa9pPRb0
rlIJve1krDRu5ErrzpqVlmOE0CY1JQoFkQjWckvBTucLLfFiDEGHnMxWung/We4GD5BkBIAh8z3G
16ktMG/uj8ZabyQmgOV8GXYLE2rrU0JAZnt/4Hn4dzWreJGUC907rbgMnfIKt9bdSflQ0vwsDBsL
TlDnZ8dvKfRptLYAj24Os5I8NrdTac5Eq68JM2CFyINlMDlHwSYzYz34i08P6RsEuMCvdxCpsrKI
6f0mM6jIQyV7a3DjXNiecE4qxVw4Kudi6sw9MTq8dgxxoZDoCnQH58G//x3nzqRbBqpQgER1dnDk
gI2EB3Kve717K9VXNd46wSPcre9U5BEmehsJdH98Bb8ECR4Fon0Kr0LvpFyLslRjy1Fu4RZzGN3e
Q7AakvLOT1mB6XJrSVbCVTDVl4dW3G2s5EEOr+wrs+4Gs3Tr44FOEdC44hOgMi1KPJ6hNvNUmy0P
cJtWRP0pBpg7HkKKfD4GzcjDgi2xtv2W3SfmtP5bVSN3Ujt5qHQ3ht5jwsS5lXNinL5bXjtfpx5W
xjK5xUAKlU+eVRCIF/lIP2p3AsHQysht9712iJiB0txYFuhW+iRPcIc8KivVIYXVGUnhb6tDkLQd
3XzIgo4oPkhzAs2U/yVs/1e719u9dFsvYXI6j2L2r5N9hUGnFR/jQ4zrHl/qO2zq/IMygjdMnu2c
4gDQ/3gClt37jIMM79JuWySILe0wE59lw4erZGbWVvWPyNHmErbQgGhcvG4AVIj3nBCeQkEBd43U
Tyr3IL+gTdSxfFyzZNsZWimfuMcIn28vXlu4h4MdxsOFGwIT3IlKQ9LsPY/Y4DZhTGpIyds4COzN
OP96kxG3QM8V/iHrNpa61ZAhMlnEoU2NYWkO9K9xrcux7aAMgRAj2KIvtiWcKj8PyhooGvECSDC0
pvC02a2zh3E8gmV1QH7tgzty8SUlF4cG7LU9p1pE+0LiYgpDhAZva8QMoQ0WbKrwUYr97NbBixnD
WowJRzmnO/GNSfpUnXviDxvmLinIW5jsWI+RoGigK5fUasV49Y3Tsu3aIEGGIkWd8FSGDk2VYW/U
pH27ApV+Jirotn5hdO36qGOYSYYKWwo3/f8ndfRnM37XDxxvbNEg1YEhGoEiJdOlsgqmURG2+KrW
Pr0y7gW6A4BS4B1tX7qdecYFne2HZH7CjEkdysqo1kJrCSDYNXgl/UdddEiBnQP56btI/s2onOBJ
+bf4DzB2EwBMDBLoscCNkGnvAgIJbRMQ9f+YB+pUOVq8QXzw4yMD0wSbOfF5V8z6he+K7gb6oSog
g5sKcOSjQsszyDVyv5HPXXzIzbvIsJfgLo5Eky7mEWBWNUCN4nVsPxtRaZT4/qpE79pNsz+TGUug
lhwjzlIFYXb44Gn5PFuWOzROT2PkMeTECLaAQPeES6qLQ6DWZgCfc+e2KW2F4aq+UC9Snc1N4tLh
MhvW4hrnTSbsNSQ7NaXPsyWsJck+ejvUpAZPILac5SOhweUh/laROYpB2sP77VEVX3moITx7F9wM
3Khjl4DkOupepXhR8X6Y8X1rVFC54/nBWyfK3RIb7/viI2i1L+AmQN4EqREud5FN9Y34uB9n+1X5
xO6dVzlhKY85xwYvajGKCBtzqPMBX8PMZKT1b3yG8DEJ2Ijl0DESp38jw/wgnz2f6DaCfqOgUWut
nIYUW09YuGu3qSK4r0bDmuW2MbTEWk9YrDmJQSBXV468SQ9g9vCsWKNETTLBiyXe6h/SkJ8JVP/X
LuAEVqrv7ioI166TW6KwH7PmvNqnUQfM11l2dcg4TIoE2aquj4E99pFrNlWi2lQXmy1s8OE8IW7k
Ix1xMya1Tu72gI75zJHDctFWPZtepG0Uo44gSkxoLMO89he6Vsj2CrFCC3u53KhlNH5N7xo3w1xG
fqDd5uwJL14yZj8b/bF1r2D7Twx4saSb0s3qXsbNpR83l4n9gYhl/KIay+0U4tDhNyg84jtIrhki
bAOeadKrfKM/6CFcCtRBlJnLjWZzpzxIr1m5tO74e0/DjNGTSoeet/Ra4tCsVeeN29chUpTr6tNl
I5aLU+JoOU2ICQgpJUrDkWO8jSQfDjalDzT5ljGYn0bnAucdSK5+RQIZMmHdyeYueTq8P2MaJy8Q
cN+BUD1BkjbFdK9zcpefHlapNqQF5ZcMlwENqq/Mu4CDTAl0CcXyjqIdlRbwEhsfExVOrKWMgNsT
JC9hoD9s+/ZHTMMKTErqW6QcMYw0cYN62lI3TgSoVc6WBsbTgP1rzo/7uX9QW4uRBUzPo4qO2FfN
3pbeahoPPw4KGer6INzS7FggEY2lUMUFjFPDL329bBRE2tmVQuav3PYIIh562q+c8ki52i5Dpb4k
30iJDk4in80wTEMBpZOs7hmnPZJcL2rBLc7eMUlCYMWdF3oS8sTUuCaOPjS/J9wi3D2f3xlNNi1g
YXn1sG7Pc71z1Zz218mKo5pkVITPRjdQjr9/WOHgqqmRlL897zL1Q/MZEBk0fXskbwt0+DuHs8Ic
KTFvtzUtTbF7SQpYn4Q63t8tL875DbLEv4urJUHOkSpMfhiG35LOnCNBJ2wyFacMexEHD7ezF1bV
iumnJnfLWjVqt9sXDXORuQsDOd2o2gklHCSRgdvuG1t/+/NIpRvUf6pHyAOvtcAIhoQyQE4MBQDM
o+IdtRNxR2WWKMN46SHwZeTFReRsxyqnMkwyk6JCvFMNKqTmIHSk5KQrquJMY2VDAz2JWbmW3nyG
232OOOSwn/BdF8JShspvdtXkon5cHJs/rtlXynN/7KptMT0uQJVgqP0Wd7UhgnnyTySJZMlJTQop
dFMe2uX3LE7JvsyiZYxFjHZ9I1y+o+3tbklYDjViBfxXYFI2ogtwA2RBeH9P3HHgiWBZU64Oe3aU
NhfE5BVaZ0VKjsk5NwAhULz6vCH579CGBShZUC6r8eQBnqbMBTyLN2/bOoVhfmSrc8kLojHJuHsx
w2nYJjAUdsHe8uiofnz06V0UdMH+GHhd7Bcl0amKApe6tFyCD/b2uv1K0GH74FnGKq9TP2+/srmC
ck3dX5WXcZNBa7c1TKV34D+IPR4FVxZkF67ixlQ0StEfVfUXRij+x7KxEmyMydAvPaeow+VZagKY
wJM+yf8g4qaRoC4wuv9sHt2VhsNK+RazPwC7u7Im2DF1ThvM0SfkwwTOZEeCuf/uCJqfBIhZjkcm
WtlSgK4TGefUSMRLhtl8PNFjL1Oah05RAzZM3HAu8A8mpukBWJ4fFhhTwFS6OGyKMsk3VEuFEk+r
dCmpV34iCtmDFblfuki3Whix9ALhjmpmAIPzhs7wQG3+sQtcsH8lSl8BMDrB7NCJT7J+M33jArTf
/icg3wDY/mRXxUN3fqYlNvBxLy/yVIpTZxmF4ppRI5oHaNOUr2XakQH2lGHqwcwv6vAciH/hnU52
ZhPrFKzNQPQGtVvjl6ZyV2txdrVydv4SVLqivF4Fuc5cqY5hnRUJ8xgVRVaVHruJuO/snpMsKZzi
DiQNRc7dGdfGRjEypugPvOu90Fpyl/Q7vzqtszo9EwL1MaTTT/Ff2vYZratO+jfmWopaEha+cm10
0XrW3dIqj5aivxKRRE7tXEpaSJLv8fWZ+B/e8Gpp4a6Q0SfMENVuBwgLzUIY1Zm/1iZQqq8oi0e3
wDUIp8MsAKWZ0PMu34+11HpSR0/0gIjaevxurCB1VPsmQQSUXKwVqH2CgInh07BJ71Y7zo4qEIld
u27vOr9DyOb1YIlVQ6HdQONNgfo0jttAopT165uLCCcpXHaJ7s9Jappmg5f9ecvC5JfIjnKX6KyI
FgS0jcXTQndhZPIFhLqKREm5G5tgXnUj3HE4uw3L/DlvDB2ShtZFKqNiNykdd3nCtWwZsb43JjA1
/mdiAG7PTn1Z9IG+XYTHjzjk0ulV1IxQugFjvob64SgOjysqp8aFS+nNqALyUC1Y8ojmZCZmZoTZ
UA0XsqOFeF72hh4Y9xM/OdrodLzAoFQV9awZlRsU5FuAc+EHqquMwSfICxjddz+J6YKsrgN7i16P
FPjSfFApUsoZ0R+Hvjvp0usUUQpUU1ZILqr3mjo19bNVri1jmyghiDd0Oid+OylM8lmuOPJ2DOuF
QAbWsHFXfIkwrHodzKKAsbeQabj9dyKzXSoFMUvkbhx8mvDID42GgGr138a97nFMd10TYCvy1Zad
8P7URFy7goRFXYbhKhlRnKUkLnjXRUymhmkf3US1K0LOX0lThmV+cK6a77Tp/5tFGwxKoXMQCOnC
Y4jtVcuZYLQ2uZY4SuSSwVoYEc2X4Y9s2piMh/BlvS+/zKPOQs+1UNxyEVVgs6Y4zBdgzWnNRNnl
ybqlOodxb5EXXj276VXJg1sM9vtD9eazDx1ovSzYTgADuFjWagMWvgDjy/UfI/DFpKojchvXy7uQ
GC/DFUH/D4h05rgBJGWsUhlMxA1hs9hUkfsWUL2wCfpJXmQRSNm0WW7MGghnoe6gj8KfMBpzjX1Y
bxF23o2fLFZOYfOtYZrf8mMSCwIbMFWy+2r/p+KT0wc2yrcSudBWaaDC8zPg249qI4RejE8ckffF
AZl3zSBp175tRhmDa9jvs0qq5W33dCwyDRV0ERar1ooNmWIxmYcExZQIrrk1kEXto6AgU/cjJU9w
rHrqs2B3SkM7y4FQynV7SjGuufKGY1t65ZVN6Rb01enBiRQzqyAKFNlPq6bCduirRS6e9aqsILpm
9hKPWWVmi1YNfVJmiki61PSrrtZntvlsTtqVmTUoWfCmilUxqntbZoQpzgFvScD9pMb85Cge8p5t
khBKxcJ6wRli0AuwVpHpiHEewH7H75IWL2xpfbHsU8Wiq6+AAWGy+RGWX1ATAGBCsX/rhL2/mX1M
ghoL7HV7QcQ5UUGzzVPPrIcmHeU5dvG9Qq+RmPTtrcp01bf8vLl4Kqvra2IgMRZ1WqI8/6vMNNID
n3GxZUFzyqLPhkGWY8BSY5HQ+UuoZxsOBBCmuptBPzexvGDTs/9V5B93Om8uupOaj9VizBdIk9qs
OhT3TRyl54Tc0h3usueWngpIhfU+gkvMPBmPL8yCdJX6Xv4D1JbjgZYz/eKu52MNmNfg/2j5+P+n
n7BTL6nfKcn69jkQRm6hnk7Kn+n6PtY0xtfLxJBW5BrEkHlMGfJeF/613gNxmgY4g9rTcohVTZls
qRqE7oym8Y3+Tckn7Ez/JF4wJ/3VaSsuTPwhZHdJQgPLJpgKjw2JBIwD2xSk5vbmRjSVA/zab8Eg
2JEhrf5OjFDoquSAHbj0LZrgTi13L0tL7RXAmiMIfkc7P8MdScWGUtDoyp+mnxGyxRXkZfD41yXC
taxpFjCdveotgae1z0S2FXwEqhFsxwbpw3F7F2Hq3Aa4zVtJyCK0oN2cZWavYshvFqaY2du5rk+G
UWgydeXeYMbMS9uqCCUWCmWz2SH9XhYOyj9Vp0kmiYrh85QW1xJyG3pzmp0Cs+slIDHSmj3hZXGA
0NXVK2t4fyOa4DARqMZM6cnVyedY/9Pi+hzLegAs5NkfC3hrCjokNMEjMdS4BUjk2BmaSlFIWOq5
t9lFhI7AR3OUIuBLHfl5RgaHuCGx2YdNpYOCPxlyDvY7KqKb5t442yMP7mU3W9CmHganrKEK9TBA
5ZZfUs2G5T6QpW+SXHvuB29KOH9WTn5sWfevO8xfjOV/kuqlRPE6VyIUZPEujLckBZyzNNzopYH2
PT0xxKrcaYjrGE0rCdh1taw3D92mglajaTcMUawaXQDnHA5mMcfpj2bu+DGKxutETOVxE2N//f5T
lLJYnfkuwj6M6FcXQVeqj6oqZDl6jJyhhPJZ9bfW0tLJJchQWpv5elrbp2ygvK3FcdOox1nIcrdQ
ga3suCQVOPPksE0BGOmTTSabry6ljcFdD0YIMzmno3jltr8C4laD2SIZTpqcVd+KsHJ+3QXzP7xJ
2ABCvgp+qAZYd4krwLtrFHkEraWBJMVur3RvycqY8SSmXFXjaPmZWBWwgoJ8ScDBw6k0QE58e8JN
k3uO6LTalzSlC7Q+pNEXVb1de19k59mfVL8ZAsq4D78Qu6+iGc/8cDv6eGcwVvzjOnJCEWaU8TQ6
a5ZMmHgNjI4cBqw47ENu0abMjCuZNxZICMWpZBoI8qx9o+cZR0vGOh4PXuA7ZpKFR/7JnhowlBVr
R4sUc7rZxL8t/JoeGhPyKQT5RUia1SsaQMBX0xOj/Jp4m/N6ICbbsABdo7T5j+Z2NNSmezW+T9gj
zapixpT8dfdxQE9tC3np0zxEtFWk8HPyBnVB6qSC81dpIl3I5jZ7nHNL37iP1pXQtXiRf8vYTUD1
+I+2TWldPa2oO4UCh2yRAyFS+eMILyhnDnWBtEN5efcRdihmX7kdPX6dXOoP06y39oxsloZUvI9j
Lw0t46wAWuPIik59y4Au8r7bbvsn02T9RmYKCNOWd4aBrG7plzOcisoo1UBBKmvxFtIBcUwJBJ7p
3g48BM8lNykSz/9GpeYer0zA0D3OtHY1K5XUnmUWsMyyM/DIEEOZPhSjVj/S+CxKJMp8qFKssf85
juhfBYiL7nVRjujFpMAn0eghAsCIu2asoToeJUmKwF6kQ5xPzof6c/6nH+NTeyXZ8Qzz5Re8kcGF
vqNR7twmP/Wu032JOGQTFDXbJPiIEgEuyVyI5u19j8593GbZPi4bVXR0vrG4HWOwUFIaB7ApZQ1c
j8UzJ6YSDA7g+BIkvXJUghdGUZokSBWlwth++sbSFEDFLIvR5LPkPjXxFRGlpKFKDIutaluKrfYz
mZnQMizCMuTCu/mWcRRoBIsbjBwAAU4kHH7GCif6WxF/E+xKIVceCDNfDhXD7SCPrQVLlEkWhZQE
qKLBbbi0tnUCohiVmn2dEMV1W7JJJr3pXkUY+yjoiXBJWX8cugfpxfllRvVyxqLwcOPh/2yMbqts
vLY/O6tg7eubYUKkL42lSwRedLhUdzPsi6cwVhv9KqBmUNpdxwvr4neVRk8eN/MyLyzbO7llCSVA
cd9KbFIABgpzOQIdvau6Mc2ptNB0GwgwgsqEusbIIUUi3T81Csh8QqRkpP/fBG6KIw0OHcqkl/fl
4HmyOOutaTMdknRiE3+bA+QeOZwALulOfAffeYZJA6tSMScJdM7uspP58pP5z5vZwoVMwHiMAg8g
PZy8TqJuSkuyPnHLdIVzU/bU22OGsP9QP557eawQNm0pXmyYM7G2v0Ux6gk0au9sQ0HMoPRfQccH
DobqPmcU6tiV2q1z3zpwIApuUS4YitPvHou7uNL3V6i5QNV9mkt8sO1GqfMOcyRHf9VCKwI3iBgH
sfVG94oqbHor2rUPzGL974NtzekPS45KQ6bSODJQAKkD1c2J+0XbOCCtL062mBZS4KWUXE/a4oN7
eLIcaZ6+p6VhPLbjDLFaGAI4/O8t1nezWYXaFguLXfRJlYjH+OgEyDq/6Y86oOLZiKDXClaCO9QW
hIAJzIL+Uup3FBSXg/m73hPt9eSrkZ8S62Rs2ipY5uXGK18IyXLS5jkBZHlYJdt+7xizxvVcb8NP
LW2z4HQJwMyjJcc71AqvZXvuPiQvRmqY8aJeJGAr8xMFftSg3EQDW3eoemBhfR6oyc82dnVaFtsG
BmFVxv6HZS2btDh4PU/yKihKl/cXse6rsgRNmLxvM7b8zEOZLGacH10dJkx8vkr7fmn6wwxLbq/d
RTUCFEg9s0JNo8NPd3pHOMcADz57Adt8QCFoDD0YjEuPrI+YaDZZ2gefgVSOu4MwoS48VeFgt3WM
3+JVbFYkSkNJLzeKZObDGm5ZiXpuvP/4tHykykOwKB/QVCYSSdsKR2P975lKoFeFFNDw0mWSBNVN
hJzYP/9zVaPd4gSKvHWB1jqewE2wnF28WmEHm88qimf0l88HQ7gZAa418E2+fR+8YYXSR8ngazej
g4jiT879OBtprCUxfyPZ85EdP8kJQRSDEeFqdleCvCKWiCT0VEPusNN7f0+NnEBPa33D1InzGJ2L
ArPsGrQkJj06la09hiTb8OGnRcOUFqJZWtPkfNsWvHzBYwKtuqJYwtt4d2yYiAAYMmlSlsAyyq+J
Kc/NsBp1kgNKS05xmT2Kd9rwaoc2Ejx6tC1LpObv0bK2BizYXyuKzETzKQNGPWwv25HkUYHQV46x
loIv31zGwfQP5VnDVSS8EH8m2RBAiWxONmE+D4q5E2tzK+W0GoyNlUQ+s5nlP6l6Q9YnPVD4LBHb
kEiQmckeeoqc6jg5FBxYSZDVDsdaxsUsLUv1PddgwRdVw1rjlGTbIpEZlU27hQ9q26BsqfCN5OOS
riKtGYrGCMxfSD1HhyjI4nvuaFu4cniy+hOvk0hrHzv+i580n3etoZpwKn9L9wecEN/Phd35543v
wjc+UtAVXanWsxOkL7IWwpD/DU0D2va17Q2IspBGjyEGeTv0WvylTK1YaSTBcAI70lFiI0NWLM6g
q1CEN1+Wo3mYLcBudg9QQcHebqBhwiZeSP3vUQw7JLyQ8cXq/9WBIq5bnHukV7f7nbJ5bYLxtxB9
gGdk39PRDjcpTSSjES7l4UW7+nV+FX0fGZCfIJt/tegqWXS3e6K2F0xIeY3RcKTNh9NEFsijjH7Q
H8IzkWz2HrfeebebghN6HZncCE/sNDYIIzrPa5Fefe6UuiXrLAMM+K1aAx4QkvVOvl6647bY5btN
x/k+yMEz5DdyBXncyvgaG9wUnjhxr0NriezgPKd0x3DGQF23PDxK3aW7429qtwf2L7UdJALxk7S5
UFbxvBoyPBTWUC/8cGqhKkkLZ1txwCEoQK+xLRXj+uMERlqV+aGdxD8sRiJgWV9idYQn2VkseAX3
L6jscbuzETaxTCIkDBwTGnDgytfAqVx+f4oklhWnSU1YnelVmejSDG7RldU0f1g6ESDWOJ3MEx5E
J9e7C8MojD8gEE+i7Igqv+ZR6QPO/Y5U4rvAF0gdUJY/45ZLI1NsYzMF6/UW7n9P45hTjc3ReEJH
GFjqYrzTtXmtTTUe3GVlQetvbeTIi+d1nXfFKWVrE9ABoZmzIx6u6lKjWNNJlP8P9+A06EF10Bpp
avKPR3w2xnYUJpKR0bPLL7jlQQ9xuZyYNW2dy6uxV86lvfucr6G+bzWAxYBmnSjvAlyhW0F67HkA
nR/tdkx4+8J4oY2ArapPJLQgQis58+onM0FowFzybqA3deT6nlQ8VbdBvG2u/oVOlqEbw5vM/OcD
woq509gB2EGMqsN9S8c1dE9FOnEu/nlVvj01CpDvOpcBdgmFJZbdEqIbPpvCmKPsVuLhGl6ufNuh
4qZ12Z1nUCSaa0aIAGkA9wiDl/opThekr+jTG89vIyXFlNyrj7GO5YTyIWFzfYvu+VLAwcq5B7J+
xyDESbXF7vHchyP7ngQ8se+TH3gepMFa9EEDCG/ChdI+EzbfWwYIs0L6kM1YTt1kYxeoeJ/Dg8wa
SNjWceHE7ExRxyygbSuIsr98Sqhb4biwTyDy9vfQuXHLQQWf29U5qFbc/JH11G0M73qUX8ixA7oh
dxtO9spM+sE26G6x8cAhq9yGbJ3eJJTAr05sMcwO0OTgqXf9KWLN1agDqzpCKn8dxk8jCWOAt4Hx
V/oMifvVo1twbCodm9WvEasMAwwizN1epjNM8PKKyFjQsEEZgGS6Dd0pe4g5kgJK3PFnxQwQ4k3Q
uWyWy/iy/E0MOwHoZu4RWixhaZcb0KCg7lUdOYH7x5aZlCnVpkvb4dTJ8+lc4hW/LGpp+A/4T41k
a5gEsImvICcYAzHDZ/IidN4TO1gMsPDIZKqHuHqSONkrWNR1FGF9T+KDf7u86vFxwG3/2YtgO8Yg
SEBK0hIOT38rU9RN6ouzx4ZM1Hs5RGkRcBYRDx4RmwQBEZySFAomJYoq6SlCMTAOKYajIunavJxL
2DlTfw+nzPzDmxzbxGOhiljoCAryu9+Awyxxn7OMelcl9Eotuu3BuyT8R42ypWHxuYpKlxhgozNF
UlTt64mDEbYbX1YmcsW/Jef7D2ORA/+GiuH4BZre9yyxT8pSdelqxuoUgBrWnoNNzFnUo4+WHIfT
qP6mxNUzfczBTkH3YhW41eyRycJIk0zHbDhDfHNoZQylMfd9ItrWzmPjGPYvwxeYrMCA2Mxmoirx
hoXRy2Kfid5GfmUaRBGaXMtUMGF+gLoK9j2d48iahVq+8CXAgRW3Ch00LZaoh3O0njel+fnWuzbm
FDCUvteTgIlj2Qpyb2dCoiOohqOImHd/jTZPSjm9xd1KKDNz+uK2zUIgdBDuUzPkI+zS79HGmVNr
SaANPYNn+NbAaDUCC4xrwl8Gu8PSjrQXQjKUqMFNgy/knx4NfKxcmGf1ml3+OIg9xvwgaaD91gs5
SuzEXarxQQXAy+5ANUZ3g1tttUbZReszfjnSyJ0CUeogWYNBkDznthXDIBzPsOEMH1CSdfwvHOZI
r0vSrMTt55qktZfErTFUUl6YDUY2e2qC41Vy8xmpIZIhdX0K/W6D9UjAkMbV+F53mSMnNAukVV+j
5Q+p7AA9mIwH8ISuWtJs0Lrorez/lGuXOUiMcVGA1C9R/EKeY/3EkwAVRILsz217hKzn8+j2tONA
54Rvg5WJMKkb5OogcsWx7PCzVyn+fGMc9+vjxU3umGUhb1oPQaQZVRkDgiM4fTAjOaA2r/WlWEJ0
A2myCtKi2oQUne+lijHd5e1N1X5BXxPPsFmiDTZHbi9fpb1+2xDO8MGbqLk4+W6eACszgPNphXGf
ssx/9pyL5dMGTgpiISIWuv85Q3jYJJ1KkM6jk7tm58AU6bBMT7XBjl0RG0ihNmCYuEfTMePgVPWI
xPG4ghF5d9cwfRgCHRcat2lLavCzkFRxSyWcL1AEYS2hxmrK1RzkSz99vZaIpUM0QVdpoeLA/VhN
WrQulTYyB+XP7pFUlbgOt0+kKIsXGIcrU9Fhb91SKpV/jkcmzyWxYgIivyxIcfwfQI7ReKaFwPOQ
1VUwHA7DTs39pis0A24wtsliW7M39SqgVl/DbFauWwoISddgnydQU3wtHPyIrZJ2TC1wNvQjU6V1
4XQQ5FSd+zrcSqLM2Ks9MLLqvdp9lyf3kl4KMbDnPcyk4FBkq/wMwos76vJ5rbTtukI9XpkUo2Wf
K0SBZ8RokEyv03t14MvYo66+pZpaEV2DhLTISYhH+oHIDL86F2UNyHZ8sNFegdsZUhccDUc9XBX1
okBhBCHdo3GJGkX4GS2WXRv5xwo3ujLEGLG6xuJXGDNvGPDRovE+pMD3aoHpHlAGRFRDTV7l5Lmt
5GwgsTt5EIyYdPH/PF7JZ3RPbJIHNH+teKB5H4ufqTzLMjvqQMH3g5OoNUOLyOngV6eDcwST3ADM
sfETa1X94uSE1DsY1OZ2iTuWAFfMzwL6gETUGAhK/p92DKX6XOpf8+DwjXOw0YuY6ga7wp3Mnlo0
FA2FjZ/vN/QC6y4BL7s/oPbK4ahTd7TT1bEPamH/PojhqZn7aDdz2aZCJg6w0J8EnTA1OMu3cSbn
t7Xd59d8og/TWcVBHHDWpI9X7qg7fSLg0X8wmT9zTv7Hbsbc6h4CsSy9VFZW6MwuWNBCPf7znQbS
z6NJPy+4x0GWE0u/DZy5IwNXrKwaww6e1pusIs13Sb8NhmDhMG61sr1Fd3qzsa4B330JwIYMw9tm
ehYHHB1c+dKJJ9bZujOSDaNTSFK7/Rv/2jSTf40/erEh1OCeaM2Kdfvow2XBV/irFPp89y41PK8/
fjBVQGmzVVv80JTwSR9fTFCJqFhk/TITD/8YLnpMyLTk7VhBLXAiUOix8pNGoqa6gGz5t8TF9tei
HQqFHrvJjh8gwQyH2ttPy7VGhBr32ZTWg9GO1pz+ylBJ9g1qxrYrOLqsG5KXIi/sbqiCuJFffA/J
1B1NFctQR2kc3Qoi9O5EDDqZ4iuU8LaYFx/N6rghCjl/Kj7QCdb+5BbEiWxpuJyAOyfZlFO2MFqC
xgTmyTOPyoFkaIhixBlhaxglntiz9/r8T4aSxffN59rIvszvq9dsdbanR7ntLE0RmO4Jzy1u3jU7
1sv8uG6F4YUBUPmps4Urw4qMtf57mWyScYJrRxvPUuzUvr7CrMS9e5wrrDtX074n+BSvz8ps5M3G
shmNizpxzq+/+4BKM4H4dMkZPT85X9X9s60/f34vYaDi+QqQ3rp/RY19xFlrAT3cSmSpMj7QJmsA
zZsyjSr34cI+wYu+IA8GnLMhyQpjq4d/txH8P2cAoz/ezPPPY5DGJW2oTUXBluKNjoPsEUC/hNWx
O1GNIaPZEoQR5R1SDsZymLSMp8ryc2+n5QW8DYP+CeMRdPDE4CsN8QbDfKtOi7/b0JH5Z1NtGn5p
gXuje36iRtZ7fnFWRJSbOqcKwiwy4HZyYe1V5NOSGpzXC2hM9Pgk8OUO4giS9Tl96q1rswSKKRTB
SY/pv5oT4otzstgIzg+rj3FcOKPRifFvFMK9+M2dCPJ3gGzukWalfK1zXhG/4sFy3YR8uqcK3OEf
U5cYIEyKd1xKVc64ncaQZyQ5+mFBqUQUtIPRil2XtQ5RyfDWFi3pP85rNX+TkUnXIeGNeGuKAkqB
UrD/yOvoFl1n3hfAzyaM2PhzaqIDV0Ki+aBtNQFnc2A24LIDiyVsPVahqBXkGSKIfNy9NdVrcKFH
V8+w8t93eGrpm0qlazbwnT3xhAO7UGbXCzBP1B2foL8XTiG9BtHXtJWtk7yldn7Y6MYVjUgDa4fN
QRAdJl4ZwLaQG2Ivx5OvF9x7sc8U0gRPdiAN9gXtW6qeSu0ml/NWSf7fSHvGqO+sOlgbLCvT7CeE
QnUXnkL8r8tj4nzpie3tD4nQ0m0NYi4Uf1fWscOwJtphtEZap+AtaMyqhHz+0r0jQhRoBEBpPNzY
mW03yamHRANxjpjCHYu8q3qpq7zshe+NITcFEEsXG58oXL4840V0jeYEV0DOaaxB34dHP1GYkqns
uPKfmh0OJiOreEObsHo55CyfLInQzKI55n5f2mzZwhnKkQry8TycwOVw9lFIiDXTHSTV2oUOqroe
T+R4jlLFcJHtPB7AvpW8o+YID5+iFKoUaExYRB4MUbg8h8uWOBWgHsyMIh8DDGCN50w9/kdRALgl
b/A26MPsbDI+M2O7KtKld/GI00QbQ1BSmZXpMZ/qlcDJYXgsJQyNkkh3oZunENCRpMgahdTdrOw7
kHFgBpAR6MNgKj0bfuD1ZbbAaSHqdSYx+E4BKzM7dBBhdzxWmSGc2KP9Hhp+ha0+txTpq8k5WABh
uF9p3GzzQHu0EsL4HXgEa2T4MXeQ/s1VID0xpaU7PrC3VTNtkJ7Mcp3B9eC+3erFGeoa5RXNUiYQ
yFHItIglpWY04a832XTkSDzhJAvR/N1P2b+D8diUnwqIOokUvvJRWVLiYtZv5C8iR227w3kSn00V
2UORJq+59wHz5b5OqYOaf6steIntHqgjmx179R1BaNBDpcLGyWWquVJW+x982cHpR0bjF3p7e9x5
7/ijPo6tlyUWvTsj9GPsBBSZRuAkNX/s/2LXOxAuQ7Ye6ymXfcPiWD98gNN6Fyzq9xLj6BmaPH4W
k5C4EnXYuWgmgikV1zfBdM5d24bw08/i9bExBzP3L++jqHZseZWcphGV9zELo/+SoCLME5BGZfcC
vAQBulMAkzi+LKmV3Q29NsawHWWBtMzaBP4OP+ezxx50mGUyL5e+5wj6+xBVp6EPKtb1Y0gQOWRY
cpK3r4u0/lOVRumQWFz4uwTE0tJZBLozGUS5rchAF1TobtB3B+SyDRPZ26blLIOLWm+KPj7Y3JSr
tIoHjKfLRMZJhpLDWZti8ykzjMQgwaCxdH/K26hRHx3HUmP6cmrNBZZNox4a+/IMyIYpUuh8by2z
BHO8DR4LpzvoeizyqsgzkY2JPsQOXtIOO3Ax1h3XEBOQDn7+aWVClu7pVKyb4G6+YDj0oa9nnCLX
CwY5wj3hKN2ARPNqi1LxG64MBYUMMrNBQcK1FC4fSaybyMJtxZnfNLUO2uINkWzmDaGf2dqrLJta
yDLfpCGLkrTcMCl6QgH3ZAbdxYXtmji5f7IKEhKwCmNXgwMM4vcVyGwky9gmQbVRR5ZdZneoPWyt
6jrHeZJ/uV7V50SGFwPrrpCaiRR82E5FEtLr65XlXKb34o/R3VyKJ6misS1S+Iss0gP81jnh71sW
0dgaZrxFI4uVhoqjcVThBEF3rMWEaYYQjFTRoeRvcVmrZkXQrtJhhVF2oM6s+Xa874SrUqEkzJq+
Gs5vfVihWS9qJcAkLJ1ckr0+cR8715Y635hc0XdGwNaLr5k+XRONf818ZFFJ9k5a5XYiI6Oy1ZxS
iNeO6aYNC8pYQGH4lt7Ldd8Q8NU41nckpIozZ18tKRp4U+VUVPe2nPP8xBbTb+KG1SL0ThfU8p4C
cvZpAREW0BS9It3EJDbRK5QIXtrTRBG7Q2N+uNKRyI4opi5FdQJZa1n3QIjO+4ktaOkowVfYi9MH
mcjmB/i40/Ji4bDe+nZt2t91e8+PLnroEw5MByHy3WNTxWKiOiAdt4BiOJ0YEnTJKCKh2Un+eSY1
9b7bkC4Chq/pPwuC7t4YThmMEUlh7qfi6/Nr9nnxnb7eRu1IniLzxfktaMgdY49kR9cghA1SIExg
OOIHtnbSLz9vhDvDW5MPcrJIhdvm+cCu5sUINTRQ5y+bE0+ynxrZA/I9+pEEJuQoroCxasPPvEDF
Ro6SKgP5EAZ+jwWVmU/7IZgb0rnZDtvCSpPybCIjl0y4l/iyPDnicFFtW1+4KGaEptwIBrWJ3SuM
9ZGEjQiiActyQHyqaiKItGP66+LGv7znDB3auNuCdps4EFm2EUwOI5brtbMeVf4vE4AFtDrMFINb
XMeIxAN6kXiER8zGNeG57kzAckkC+4mbXbXeykh6iC85u46VEv5UT4U+wRIndITOUTGKx5t+riT+
ZU4O4+3N0Dh2P2fpcJF5soKb7OnMUxWbnwYd6LI45gsK2EAAeigRDdJA0neZ+VWqvSJy8I1eshT8
HuVGzRoRO1wqyN2OV5LRzCADgryriEz+NfSrS/CXtMWzh6YfHjYrHdyJWxjFQcpBrSJgj9ldJ42n
KvF2M1Wd7jgUMbrgfwJS+9DWQo+zoRravo5GEPabjyF99pStQ+gL3XSxDNHhRVkJT4YmTMg1THhQ
kUxUPLprYyKAasfunncg8FdT5tIXrN/Iq9usNX2eaqmp1WPoI5SuV9Kg9UkwVgEuOQ32mzIERrP4
Kou5dTnDys3GiJZRvy8KAJWyy/ZbIz4zKZ21JuZ+BGNae+KVEgjPGYfaMF/eJpag+uTB8vfWwrcc
yGJefxS2cR7sZSVSxm20TtRU8UU+Duh8f0IM8fFgCKhR1ctBYb5mDfFwWvWnItk9clE2wysG1wYg
spNUe/N9SJc4EPsRd9Nu+bYX+UQU3ywGP9I/liC5C6e01rM5mAX1rLr+tRBm0JAN8Zu+ZpeLzbCW
0+h2gwh3VbuGr2/bjZdgxzEldtPS4U/utru2RycLU+mPu9yP4B1bpcH+cM6s/IksNL75tPw4EsvH
sV6yVIKPzgjgrFBQQ1IQnlCRPqxL+7WKAZJ1gn6XQQkpWv5E6hzl7hZppwv5d68oKa60zcOL3hBg
NjCWbx5PQclYSiduAd0tabQKM9PFv0EKOJuIuDecl1yl28yNYPymR+ethpdoqWXry52QGoAqLME4
lIzXTMQvNqJTQ3FvvpqpfU4C0balTzd1g/3PBjTh2LsZc/fx3fMRFH9bQOE6IvlfqIs94jeleIIN
T12Lm3WCtG8OheKaP3szmTRkNJ/HDYivLHfrMATE+6dEimJZCu/v2/+RS/EIhK7F4e+yt8mozEM2
wzPJhmFoQIjjnkCmAkIQx3NhLTRGFxjrvUoXr17Ius/BgWurtw0Aa6Z3DdKkRRUllRpvr8Aak9xQ
cygf5GspFuVc4GPREPT3QiYV8o/1pCCePxZA03JI2HrwbD5RrOaa/yJyYiVyMCGQ+RBN3QGoCdwX
fyHKtoG2R6oGcM+QBbv49Yhj7N2cJ59klJd9n76CH9B1dQKhAEAABjSojl2ZD/MfQupyOPRQXrz+
vj/UH+sJ2JKY+ef9WktSLbPxGzgeeLnP3Jg4qEE+L6PAtUyAda0GYybKzkmOj4aEwswdQqzNTjIp
j3g+7ELjIqYDYCg4G/dewh5SoRa5DIStd9GoiAsN97fL2JqPbMPKGuXwMw14vCOrk8j9iIjW5bXu
X9JzpbQBev7hgNuQdC2pzeYcBcSdN/rbEOP9qHGBNhNpC/kAu4M7F8bDU67UJMjEDTr2DzGsgB82
UqFmjT6wfMwO215fYLWkOM3J54mSc/Lwcg9F0fCeNSAz3TjNy+dlb2znbOVyVmLJIhSRYVuy1nIX
phiTSwYFknkUocK21VEQDw5IFMBRrfPaKKJT4kDZW77mahrlBlD0XdqCLxYKrm5CY7ufw4cAnk94
yuG2OUDkgBhHK6KF6jiNRv3UANcqAADcctxT+TNQH9A9LyRuzl0ieaw1pf6PAR3988pzOFGuwk0+
voMgygqChcPi7gm8OskafgWI1rJyAk/dEb9WfsH1bn9Yy1w4Gm1Ik1MZrbTA1DFg1EJAEbGNfrD4
mJItsBOEpQs7w9qWue4Q6fNQABqfE9F90Tyfrhw9MWBGMFMF+AUubOoAlmhM22syUs8U76LS45DR
0H35iZ2t7nSs5MbGQ64zLE9xQcla7+3V3ncEKxj470+4EJ4jXxHxg1WktG96vogYyytnDDCMsZq3
ZtHtOPknnMeiwPv2l6nhqS3WWTsPIStGKI6F0ay0QJ5F8DFnIMgpMbWADAjG4PIawpIfjHEcRelW
DYxaynE4rzpHY24+O/2815dCFro0dQiVGGzQwcnB5hE0jsL+9iP0fTLh9b1hksA6GTqq7j4XPri7
dIgcNnTx15YDr44If3WQ8yIcMDJuJds0TYf6kqeeEZ5ALs7EA8eNaxIz6PzXcFP4siIBe56/tXNO
99voNTbtyWtOlP3/4hRDDbvx5fUZGGvr529LouqlZSLN5jENBANB1WMIg8DyOpMi+YVPdhW0OhGO
bOkqWJ6YXSSIAdSMsG5Ep2WqFO8sw+eu5mYMuUtJt6D/4VAUJqf9Gnni578cbbJUNk0Ysj8L4ffu
pPqX4CGx/cXNhklpvCf1HuW9+Ca9yAQ2zvV+B2pE5QVYvupqET7MOefwspxpJFY8zEmtSRL4nMFx
QmJI49BzYSCUHJ7JH58CkhQsHphe9HJ3nXA2yqqym/U+bN3ZupDWAUJFuVJD9YfLimoPATFEkzsW
KIUBD2vY/Rx6A7D5nMEqyrWEY7Kbtt0pJVI+J9G7PHrbgQrh83mLZ/amsaDh8Y0xaGZmgLKOk4DX
qSaq/AU6ih0jEfQYAcBx9YTFPTwtf8rM9GMBX1D7n8mZ5REJRzgBkMR1NZqFl+mVg2bSKJF9KpN8
Ci2Nj0aMPI5g8Zq6D0v7uJmAdBwXVztQVMTi7WeNpTCsXWTtbn/6xES6uCcYpzcYgBbF1LoimylG
YFi+mpjcoES83W4lOo49DlwisolJ0E+VmTRg4sVN+q8e8FN7uYCAFHU3igqrq5sG6e4dVeHFss9D
4xEWRSwoy0dPoMmlYSDn7p4oQVBfg/2HH6zn4/alRvqJv2um14CCh3HLqsJ84LnOfzEKoxP1oUYg
QBvgFMRzGGoO56oPx4wgjRzplVRuRNEI9dcu07yKsEuxW8Xxt4Kf6Dn1B/vJ8mPOiDwQN+aaF2Ek
u/TstakGxmTXcesLP9O75lD3lx+1NTU6ypp/VjeB0VpUEgscmyxdEwsbBpxd5Gd3N2FQ5wOocuG1
c3feSowLIeZPamhuluLpvM2RkZkEg8sxvFg9axUTS+rQDiOu4v9sORZLgzL2d5MyTtG7PxWZFA5V
dfkhWBEgVay5qtPIzAWStGOVob+pjqLp3xKMmU8H9il23wTw5QQpqX4trZvop/gar8zslo1D+5tm
giakXohyuIfTAjWeBFfYUbBMmaSdustX7Y6wp7HtWitha2RwQh5SW7iPuZlsaOOWKpA4rcgn4DuB
Ii4TM1wLCopUqes4ObohUKy9qZ36ivtZk5lcaKNxFv7PcqZKYC2Wgsg6+0jXk8u6l22/3AGZJNKN
10OChd0DEXV2HC+DUDCF3+WePcRreV5EwukFcPyhUfV5zy1ZDnsBJtwqMaqU+79othOScCC5Qb7m
RntCAEQl+8bIwEvO6riXSE6fNdreBH9IJObOE24B+UyFbWlMgxjby82CspVRAX7etzCGmWOuJneN
A+yLBr/ezHYD09804+/INhHdklo1lojmRaiieAepYIYMMcuEBRaAGBQWF8Xt9FgckXKUaP9pR0dI
AoOWTeCuVHO7BdAjaOxRyDsiAHXG+CHefEe9IKn43JbA0kF4ZTnuoNEsAw3upQNQWX0CdPAsJxTy
Cj8wH2K8fYNiplSRoiTeoUoSIhpxczI4kg6HVA76PLsXirEwE3AdotZ3ORJpFxEx52byuipeY7Gc
cVslgyw4qFJpODIjqCGBOPJzQhOySqbdTtZdTaUshgY5VGUfmcJaiRJkUztrZQYCFqAlpkwlRTiG
WV4GZIhfb4D29IYJ5rYUZ3ToqO3wOKHWqgrknx4+IOqosISToLMyEbtAkWpH1duQHYtEio60IkaU
b6UiTT/1jiwmGr6HyOXleVNqRzd0z9BpnSn0K5jkEzx1MWEfxdg7qEwZoEEViPhyphuq2nT1+fJN
ZsZ5Bs8R7vzTtzA4Xj983vH6nTVpr77NFp+TvpE70FV4n30k65O076siUM0koqrMhvxAv3Yc5imS
vfoky5vnxs5R1wyYbJxuTpEh8YjwlOniJOVBXuWpKffIpX0IR4JNzi/+Ile6fSlB9zY4ojLLisl6
G06OI2V40pru+IkXC5lOaXgFq4HBHxO0WaoGS2lGP+Obe0EkCqpeWSO2k81MsRXx6Vpfe7s5BJYJ
GSCiVhlqJS1cwEQlrT8/umHBJcfiLuyXvEpoAe59JYAysThdWIN17BabBXWD7KpfRb7W3XFrqgQ4
KqIYrH7a1C1Vc8peVIhuqhDkhFNmNSm0hXEOVDcwUce7962CkL+wygmuKlRzptsjVPGUtM52Oaa6
cxd5Ww6LewwXs8nBEZgrlSrqCSjI/Q9NsmPhDde2j91rqNHUBEn1J/xb5vVhMINFkcEq5ejpqpvo
/1f6mh1ySDvn5xI3iWCclneKcIF3jqfUCz93EqcnkwaNxMkqrK6sGPQIcd63wdoZJfwhYaVsY+2g
8hCsblVBuhJ8AFwELF4scPkBXMIdOB/bMWAXpOyfLmTYXc0rzdsITyPMkQ/40vEzvHOFH0GPR5vq
jGZo4tUhonwqAuPJC7NYaR08b5NMMHKIewQFCvPHTpl3UR/+h4N7JevOCKvuUNDdWhSs/MvXYGVQ
SkEkyx+37eNInST2aGoTEy/bs6O2FSCyFlzK7Irji28gYEITxR2wH2+nb9uMQNXImMg8MbU1ro1c
ofzvIEk75sRN6SHhcJz+MkHfDgIl2Cnpm9I5cGsHLteCBI3pocvdhYIRJ0FzDuwfQVPIz8Xm+iwu
3H9qRfMb2J0o2F6EwxZkgF2rTvXWbx0m9+7/g0OJiHykVziePs+CT0ZuexFdX5d2MzH5k4GzT5+u
UzbQXEBnQ4yJnXLbb25BKEQnIK6GpCviJUmPH+OGATuax1dRq7bVnMVju573cGY9XCOzkn+gvfnk
ygmQV7jg6BcWWjbtKbxhyTsJDVul6SaQquTaWsAZLTHvKwrE2evg3RLgQ+4oRKOLVFOLpC31qr7v
863uAtxCHw1dOeTM5jgnJQzBpaJY2js6LFd77xskNY9h4HjLuaWtus6l+A+FVR6g8v9SK78fcCEM
0Eo3c6vmofLky9dtQ/A22wKeVVho42ibds8eVie5L5jF7HBCMDKDqI3rvbbkmKOkH6AQzf+jyd4B
90D8X2sgleJziBiZfou55NBwReI9aZZDds6+254KnNnBrlBZ2iVgxRCf0ukCmXNYvQwA7ba1aYCs
2v3vYR16BRtsh7WAIQeNI/Tu2qh3ycUpniduFD70u5YhFg/o5U0R18lIMCapVD4HxifG3w+iSIxy
r6qw259REiKCeYpmsKlVuBhC08xSyDPMAT8juW0rXIYWj5WsphcThn3GBUbqLsTVowtt9Fv9hKcm
MvtX7bhcfgS4LyuXv7ZQuhhRiKrsjCZS0RAMZZBCamPisgh1lf2VwO+FrCzMridOO5pvSaQBxkkV
70SqZTYk1Yd2DkW878hhkvaHUtQsHTXI5aMZYzGdDsPqOMEtovPm70bD0oEOW3tsVUdxiBSnFCjn
ACTVwIXeEDd+dkpx4Ypui5wDb9myWnsmiGn/VFmIxRNUpUdW9tK0ILnTLqkoQD2GlL/QBe9cjjVO
79XUyDaPY+o6eEaOPmwPN3UzA+dCfIE74ESbKluckZlZogXE0pVONm5oP0YHTtjGJQ8fkzhK63iW
rWLvCP4x41WEEjW8HIwId4GwxbsIkErobiSdGoNjTy4L1S55MAoMS+VSM3nsMMGglXSD6qUWC8F6
rK70FVD/6aeTO3f7IFipPJHfJ8SxywdTTf588t+/dcsKBrbhL1FyTyQ99d+tIr8ghpTIn0k5oVxS
SSfmcxEfGWVHxIwEbakHD0ka68fXPkG5rBiUGK/Z36oFl30mDaHg8WOV+qpy4g5b/LCyOlBhxYSj
VOXQvBxiqqHCvjuOYHqGcD+RypPPnpZTNyF3G+pcWNaCcL6Vot7pJD/xkifIqNwIzTGm/brARMX4
Um39lPvGRcDF40IJnzqTaOQmGr7l5ATxxyDAi8oBdupeja1XwOGwfVnO0sUzM5EgbxAjZF715Wch
ZibKiNJv1cjfCZ3foVFCKQo6T0zJM3s0Lzy6uPwMfmXqcc7vQhFqxG46eV5x5ar/IbtfpeWhI4oc
0ZnSCTk5FG0iZaN1FQXrHqchPafkEEUn4QaO6ikY+JfZ+xgMfULO/m6imQg+GIunoWrA6QngYM+S
9yjxhihmE3v3z87yPpLyvRhHzcV//DAul6YsdjBooQOR6tgmtAlPKzR5HcFRvDYH4vePPMn2hISj
g/HyktA0q4+LyWbaWlC7rSQ2Z5+gP+NhpC5ETjBTb7G4uF0i8u2Ok4+/FttxASe01K6Gx6CSKOZI
hFdc/4OxZCXKn/QxTFPIMS7l1LeBkCqJYKGP4Z/3vzXZAOC4gAKPQZ8tnQifXf3HjGRGLqZV9JVk
TdgPav2tT5Ew42jzWX7JO6m9SkgMEcJ0rC7WXnseK878mVMEOnb4w6Ho82iDfYI3DxUiEp9hYO9b
ZHPym7Lto1+dHefgyz30mxEqVmor1WSY398iUe6jGuDaLOSmvRJeowRGZiP85ZUGuu/uPJh8YPKY
5lDEe/QmmoXINdADp51ezEmyLqfb1lryxNZ2LSI3mi61Q73QTsNrU1dRrLz6POsI3d78SW7puup5
oTHkl3WZ6nv1Za2+1kCyLEj/18xhydWLk8VZcD0we/HMscrwQjOkl8T4FCXnsx66uaKim0dDPbxM
lGeBSUYbYOWI5PRNhbk6rQOcAtQxA6McuSvxqEPcI4HAKRpmg/RhF5dEl4eInERNJlvDNN0Jqqmx
xO7jJp+QKAJ8oWjo6XUkM1+kMWqWh7OjG/AgJ+T2ldZVQC/j2Ezr24mcQfbM+VcKQ8YET39SxQzn
je0nov4TKWtPD0I3I2OS/BGfoExsv15/eCYfnbLBoK/eSh8atux9sJfaY40Qv4+2/jLfId5WaErS
0ynv4qxnO/D6mutMZX5f4c47sQFXGnPs7rgBE4K6Ww0Yp27okQzamWsk01dAUUuS/tvSq8PTM4vM
CAay1gSb1juWwwzlE+ZyhYSFDS4twjDF7m2DllyKsRgrX04f0m/sn+VbVPJ4O3tKBTYz7anfFbK9
0xM7IrPtPF7vVVgnYpv4klpLrdTlnifJYJnBr+o/PO4OabZa9BEOhtImZDYCZ9+9d6QctSycz8qI
BI6MnBx5ebqbiE2/WGRkz3cjjUz3E2+zuI8bsPOHQ6Pkxj9bGgzHUuJuVO+UvUeYQwNgpdmPcY1z
sPkeikukngsiwLFABpRVZ6u6l4VNqfDyThomHyuUsjqsYm7VnAWUOweE5JNhC6zLlOBKs9fqCOTC
wqVnmoxIM9e49PVztDTxDtdyPi4aDjWw+sRmvYxNodxOnvlr4cK49Gtw3Kd/NyaRciz0m6lp5Yij
dZdaQxu0Tea3NzEiOkebjuRRuQzH35uW0ofOiuXcJdyOdmkYeXiUtJt97v847uvyV5H65MjzLD+M
mLRmKenfUYgB/pnhe5GkvnVLUXnZBBsBOkI0JQ7e/W/5AlK6EQbNreXGDwzK5OnnIQKJHYkoGHF5
2is7oH+z0aBS3BpS9pxSgfDt5Wtu6v0wfqLvfk2VGAwNSvT3r4a/SsPTaY2pBw85aunHcCGOl+11
v1qXXJm8tO7BrGBF0AAKoE6/rQ+s4gH/LlSi+7+RCm/DleG69mF8w52Z6H79PFWlbv8wcPVAawT4
6kTP6vGGsPU/hcxXAkwxYtgyBgGXYF+XW+rJ59Dppv3GqZf41DjvADkOCp1VoBMWgUQ6X+Fn91Rq
7BuuYJRhBSUS2wp/Xed+FgU3nrj0DfPm39X4iV631oQu4zJHKkeJ5/5zOdmA1BEqQ5AGnSLnvY92
W6snKohCRDI2N8UxScc7Hag9yiOR76m9ZlITjPXpol8Gb4XcdmuJjPaJvFvDAMV+0HZIHzMgECjs
VXn6dgre5iGjqn4x9tx7NJ33kbuuwR+b1lTbCgp31g8E1RUU8mKUTkRNJsJRG3a3qTYm5cezjoDd
o1E+75m3+dgALwJQT5hXEhFIMdtUYn4X5dgOM+4GjFnOB9/BO/f7px8Ve/kceMNDjVGYia8qbjqC
dqFHIQGnX/DG05ivnQkkMhNtyIn5/wzaHJ8kwXJ6XohJZrLGylbik8YWhgULMWzvC7V1tWIvJC/c
NUGbO3tzH09mKQX+xedYHPJNnqFZQYD7FGaiqFdv9ADZyOGyNARhWqwRs4gG1p/408D67SvDraX6
aph2cXPso5eQWGKObaoPR6HIQz2JavcQF3bgLsRRzRXRCxK/HJksIGh6JH+Gs0GeJqrHtXVAUwEK
DICiiNPUJOGbomN7p8bZ4GxpZtbpQjkxDdqVjaKwmhRDLSnYYmV8xvb5Go4QPrD10Jge8FmRRkwq
8IhVXPz89pkFaXgs1YlN8ztjoeObD8gnDK11egjEfyTSl/2K68yJ2UnZFsekHsFT9I02rgStl38K
bwOUune1v9ME6edHJqKKav8kiqkwAS0tFJKeCYdE6Vez3DwDSFsrYoHIsoiIWQ2QFB+IQCCIVrSs
HhP3I6JU6ZKmbkpezOwMsHfmF0IaZnr7vZAmmLi1Jnse5J8a7+ErPAmUVXHYdi7y9zCU51wJCBwP
4hEN65QCeo5VQAgcw7JoXKjFM2Cg1rTFUIyCYnBSJ9SVfrVegkTt/FpUwEydl7yTEvl5KrL1CTfk
E7MwJ/L0A9+7iUUn7WF5C9VMiuEBC5Jb4mqbobF+cNPhHoF5M6XM3AmrZ7/9RzUOFmZUcxcOnqWM
KjzyJTGfF/EKG8gkuFRpOGVNrMa2wuwmGNsUrTWvUfpAbqfa0od9fbL2GSo7z01b3jGWF9MaYGuA
sIgdxe2ok+z5LcH3CsvH/vH4wDs6788aqVPTNTY6+ijVs7B0b8H5kUfxO9/uZFpT0e0yXT/2MJxY
JTNc/hi0UZFzfXFtht3igY9VWjWtr8dwnLyOYLAlDvpuUsCbFz6OROGzBwdE150d8vEihwzxrPka
1ohyRtqOi3Rf71iKnXnV8SIZtVGPMOUUWg6JcMCTp/SXqZye8StBZV1vPm7bJsPhR4wN2M9YGUhG
n6pqUA0HLpxygmNmznvAUUmjgc99gtP/r6pG0f7qtBqocMnz7gVOzQWYWQoGKgIzYclaKcIpCOWY
knri8eG+pxi+u5RUlJyK8Hq+X1uNlB1aj78UUQ83v4QQ0URR7t6ZIphdHjq83J8L6SAXuzahEYkT
dXq8zujCeNDKDL83w0wHhK0plXoBQ+pDOzH36bQom92wMNOAjpKiJaVUUFqav3+zNeMgnVXbmdiG
YJ2xrKwX+hc4CotKWQggcZI6ZVvj1q54xQum3m4s03dpFwvCdRMllkT6a0nFiKQfuxq2OMNmq+Zm
J7dmidhQSNrY49HlswIC/VZv9GXs8pndN9UVZ4Q/A7UZmRV3mdrTT6cfteAZJdis2n3b7Sk20D9l
LvFkL1GGMFsERiYuJamIjE+RYIBMCfz2nr9517tmbC1uAoEl7Xr058sYuSXAlSUtB2wGsSGtG764
Wu6Iwj62YoEGpUtpFlXhkSB8geKIgkSxRKy1uTdOZM7PWVO+u06hTXv2MA9qecTQACGYRb4K7R5H
eSOPKxytLbvmXGAzYK9uV6yQK52lumcoWnENuwQ7xXjVaFv4TltqeEQHAyArqF8AzGXSx10sXSRh
d9K2ElqR7m5MfNadyWti8MxZ2xps7ylC2TVzlUVRsMxxLeBwq04nP9q24dR7Pg43e1qlFjr6Qu8m
8lAdAsTjJIgZm4lrBytsfksIyzYaBymUzZuAq26HX8Y9iuuzyx8jH7rEH6Qn1Zrp7SRHMEG7Vpos
mBuV7SOvYSuLzXIEqY5WiChtiZJB3JHq8B8Jp4qIHjz5dnG7lsNBED0gb1qIvTzsvlRfDfFOvOV/
9z+x55bCZYC4TuDKLr+cVLsqGjf8epaYzGMFPtjncocKW+N07b/vlDyo2/NWKZQgf6QUq6kA905j
26yDe8x133TH730hfGpB+VAtq2vxKqj6n6GJPAXSqr0BPDfKRSAAQihUl6N5dblloawX+owDkXw3
PUE8bJeJpABOw5b8EA0NKOE2yHYyj4S30Ol4b+RaquyXdkjuNhRE7iRbPts1uLsJ7iYgskt2UM+H
IzBJjjnsCRuABnMgyzJJ5hKFiJ9WI9Kse58XZKL6qTDQUPLhxkpQzKnuZtAw3AWb/hAPOt3v0AEr
6IjU8APiijPTvpjyw3DpaBFW/ycUah908k1OibDzW8FOGJ9RGnXTx9mzpKPc6hn/eCNcpj7VVaF3
OAj1ZYMDKJYIR/KrVI0XKYvqjqPrUWa41gPH7hoTqOPwapdTBi9S8yOdnGrntZZXlQq2eJWRaHfl
zv4GASkdKDOqVZXOBeNdx2Jcqndq5vrOUpY9nYAs2WZ5TcdmaqqHiDNY2/pg84u5CX0PT3SwXk/Y
MVqNjAGb6aG68KVhI865ExTOLmrqfo8VLqPIM722FJiSbMW06clArtV6ZSk3Cya7n266j12XlbKp
h4u9IbuCCXWone9BN2r/9TFY+YCxQqLFEKnAExd7JMSvUKvj/L5eYiRGDG6KvUOD7pzrMXODGMkG
Ymsa00W17KguoykLqoX7JHUUA9OS9qizS1hoeeXsrIG9aWgaNrEnfkSaX7Wh5Kwl//gAddstYbFh
o1EnU5Asgz2T1XNIRjNfAMBzEO7UBAjkB/dExdd72q69C6qYA0M+9bW8DBLZy+Ie/Eon+emNoX7C
cklUS6dETfYnQBNV7PCw57tNvuyZL9RJaEdBIzKFpCa7Qs8dM3sdQ88w+60C8EhnHEvqYhEdrQDp
F4pn+IRcoZOO3mGw4pFcJ746M1W5LZSUuaL8tuwTS2uq7mdNraAisZIDkQZvRSFmXb/GKR7iPLiN
IFBYZw2SRaB8R/MVLVuInUJD3kimpfRvmfjzcaCQ9RwG4eA7T3S7M4OzX0JNW9KRbHKtP5yZO0U6
VejK05uMWmHeWqgUPBrjErwW4aD+e/7uDlpliW+5IIE+2GCqVtRMd3r6fY99ypX7b9AhNzmvfZm4
1coQBzC0gPbXZF7Lc8zR7E28htVKcGnPNNoTy6eNHDHwoJX7Lfp1XRi2ZELuHvoMOWxylCNi90//
5DplUXaLjlvLueHsKIOziIcLbnzICHy9wlL9LY55yJLbcWObW/uQhE0KfLgDMliGIEOdiMI62Q5q
800rdA4rHmus5+7ZJsQk513xlsWK3S1k33KRLI2trsP0I/ZgDGxDCD2EoPXmWGopPOy2j7zJdZ6j
ogTS4sNXjWMaClVW/RYDBWHhzriaDOqHJ2Db+/7NOG+DaoPmDXNJ1SrRlVPAfWOGDxkfHumZGt4D
4OYSMr/99OyKJz2VEKLxiLe2B4I2yRlqVV6XfKV41BuFkpYmzrLecVrBIeK/l4h+nSnjyaSQ4t7C
gwoF4l4ygmxgoQ/tAfzA8iVhBlR1x2RPoVqA9y5t5pI3CatGxn8CEOeVaesUH9wvdy4DSb9LQc76
n2xCSpFK3niTvMsX/YHTzDUrLipZru09dY43Nur+pbRBtXXBwFxj665UtCwuxpCyGuRxRO1ugwHO
wMBn2Ae5twhvJhKKOV1KAR8721bWmNXd3VeoKZrdac4emj7x1it1F4EJcPTDu59NDSaUxdQdBxFg
Mg+pPdoqCtw3lH40XPXT4+x7oetoofxXiuqOfzN1ZblYDWj7xcK3Y3rkZJ7v9yQWAjt8Lu97hxBp
ZUPkrL2KuXhJ3DXrfVXHdQr2GgtlUJFOpz6sBo2AYBURCKLXp14I7a0ytUjc+BJKAlMszaU/OtiJ
bgwQYnPVPfvaMOZr/K7qXtETa0cpA19416vJgWbS7cmgdInYLYDhdg+T15zURTvEbUKk+7NMwJkr
LnrIvkEvh+5U1sBBtwjs94eMZ3kqN8TH+yVi1xl8j5JS/+Uy0ZA+FpYV+8alr8qMaxHLzcFrof3v
yYIUryR1Bh0Blk2uKD1nS47JAjzLe2o59Y17SjXq/4i0lyNW5gqqm5tVjlKXjHbPlYPo9Pzwtuty
4XpGZyzKcjkctgYq40Zm2nSTzJk9Fuk4HD/HQrrVn3Y7sxH5XxxowyKStUHtrAt40QHp9/+iIfBE
cwvvN5XGwlzOExS+xq1gPI6v10o3OOiKOh9gUN1re4WhHBdT2Wg2jx1zTZINh6ozqkplswLdsUaS
9AschixLza9K2fDs9Z43D1WzPZ870JEmhNAbTRTj0AYyxex9DT6lgD9GDxwUbSGVHErkSm4FwK35
PKnD4vnMq2qDJySxXULVpd7+iRr1S8UYrdM/oHAATnwCozimvgpfIevPdo9sXTKwY1irR7xx+4rQ
HxRjelfNe+E/OzlUtILOyZVdZuf9oKMhj2PhRUzozBwYs2C4MzTJIdan3DbjMqzqNVr8Si33viYy
jc4hOWhFRm/Zz6Bat7m8hI93/cDyGLGce1PpOWEM+ZJHCQQND3kJkD9lzUhMrJh+Zz0YeWIMSsWU
H/nv4ZZm0G/XXl2XxZrCEf4cVPPgHtfnWyjg1w4C94/WrqiSN/WJ8J6HtumMfLeeu0BZn5+GzI1B
BMV88Oevp7hvztOwTQ/z06mSDKcpn83FZSTqeQcTB6id1CxF5JFtoFjPDwlOq/85mEq7N6fKJwRK
+BCcTqAgyDC1fFoKKZKQJ0yzpVNzZuDM8D5i/Hb4Sn4D+DZRDaRkGIQvDJGi/e+r/1Ny24t55K/q
KlsF2KVL31UQyrr/7BUFGcpxnlMo8mkszJlfGrIyzmx04TO4XEP8BZZve1CjEVRrhRcgBmTD56Hc
9IThv90p9xalfsvgqQpwOAGMBcfeBrR6Pzap2mCluDAvkZXH++hWN0jWPBgFcrHjesXs3nH4fedN
5TdToKwaigQK1sxZPSsolU122FpolSb/25zy6ZfaGfvg0lb79O88Das3781Wv5VZUKJPZoy2zhw5
yL+/S+ayWAzGvlskD1fPXJQOXXq01hGKFsZgm9q1siMJAUUrfyrBdfvQzhpzE+p/9FeM8yvgCVZs
oW5+v54fPqozJgEU2H5iWrWVqEXzGtokRy3WElaLIdc7Mp7LuA57uFt3CV0OWEs4Q87mwJhmqP06
ibz98ELBXr7TglWlVkLa6Z46mBN++9Bbku5x3ciUsf3A9XgZ8RdvAXQ8kAELyTceyvICqt0+Dnm9
Pa5ShRoSOrn2ILv+PiYuK820u2wF+ix9osrN1vs0ulCHfjWObOUmlPPF9E+11YbLc/6hc35Q9MV5
wkY1osGc3B7Exszr1r4aVPRIR2/11ivpviDKiiEoYR4iDUtfpblJZkRzV952N4T7amEqSYcz2i6D
VaJgLG9NMiYtJ8nd/jdo1YRKPoMfKenSo8sQNLhyARTJOs3WXF162IsCVovO4Jsn24TsPqTmMMgO
Lglht8c4fgxqnMvei/JdPd1wNqc34HtFyJDp/AAbAsctQ/3GBlEF5pmd3X7Jh5QJHTX4ABbomHJH
nGQGHIAr3HsN2h1d3DCTIvttzGKVK+ehOGldko8/nfKPQOyFF4MDl4Z+2nFbbpmXLhmLO49PrSJU
PpBTahXn7C/WAhRiC5w4+XPm8HTb54k0eDPRqrthgf+jQAyJ9rYIOB5d4yzosEBk7P8zCJ+Rm/HM
28DBGvj5gPiDc7oYimkCTFIv1NHmuVyLL2LwtQOT3o6RhvgPHqpqN72otf/TSCuE1AoXIPLWVTVU
hjtUqxcIxuyTqZyuqIi1WHCMvm8O6ndCXnjsfv/bFeMUeKRqcTLEJ5BdVb+4I1qLG+7c9l9GZrLT
UOrKZt2VHADQkNlyQbaIJObly8vK/LiB80rkrBLEf6CiJLJ1UkI3tUBbavINKqmPHfLZ8ySpP6rC
aLPUTG+OEqGE2J/TmeHXhIp6FwgMfm6cGosWQW+CHU9sWm6D4RuqECa0Hf9wq8qTlJgUdzlLCXb2
UjuY7dlYh8TIKXYMy6gw+Pk4PHD8QueyikS45pG9tQ/ZU4v3rnQ8wSXXQYSC+EYie/Jw5Dw8jKGf
ULxdFPHubZKapCZmhtl5NeKLvtLPA8j6F1H/HoOZGwVhFNaIJIDXZbFLp/QaJGV0oxg/kLPqKuXd
HCv06biaZX3LADg3pq3QTdfyWPngZY7ivwOqYQuiMVY+m0WvMJ6AIehNLyMdo4JJQTBs0ouIN7gT
nEecqillaGmIY5QsI8KMDtA93lPKv3FG0hqoZ3YrCq9bwJQlgZvFFnfs/tAP5UnazG8Q7ckQkeOU
ICKuAGTMVAzvJRZHrBhlhgXQNgF65IY+tO1zkX9Q8eP6BzVrGNzKFmAdYHltlm76CXZ0UmUPuGVJ
riXCrqGXF99hpudC1u12Ehniz4TtXEqCwcB7aFR045l6zClRW6O9cRYohvlGimnBg8IxWkThaOPp
PTUgm67tO4Zs9ugO+Jl9kzdVCCNeteb+ae7BaoR5bV8fZN88pNRTBlZzx14wz/54B3noE5PGaeDs
+GWjzehFcJYtwSWIxWsi8MTxUwgzTIIJOu1VDG+JSS6zVaoAfDxXFXwRxqBd4Rb1xi9zqe4VqEHE
Oov0X8Iql+jUAZVX782A71P20F8wuejB6OKA4yxUlP5HEUAYuSWs15QJVkd9JpZDvs7twc56wo5Y
t4+/TbkA/5Q+5b5LGgiQ6WZ/IwYIBB34GUWv/S2vZXt/2WhcAjGiCmChtFbP8EuxWwFfVEeB3gK1
bvHeKGYyqkwRNSdSmlQGHvW8uJ183AFOgiX334Lw959a0z96NxidQC0tpqoCP9YAQh3dG++Zx+l8
F/P/BCFZLNpCQfjHOdBAduAe9k+jPOo2g9IOjWI0JQciwAxwLBTOtkYybaokZ2cqbDRbvg580+Ee
04jhmNSeFs7Avz/LVOimwA75XO3hyqekffi+57qzabb4r3s0s5udOBa0rYiWxbsP1OBqe1WzDqU1
FIvnkaKUFmWmo2TTmAyjaos2NcKYblvIPnPbjBIW1pWy5Yqo/WVNpwDe98hYXIDDU0L8E4xlB6Xy
Bz1sXKWEfRlSJE2P1ljy/UfcXmyX2d9qI7wWpO+9vZj6yjiBhtMdeL7jKxxD3DqKZ9hHJtDG55/R
bJo4hkV1gnuElTQoZOV9Uyg3rquZ3rSp9JBIktMkh2Wb2HUuq/35O4gWETt6oRLguq/Q6dCZLUTH
bpUH55Yt8/Rh6I673fmACvijtIHZzWu/juzcee/+LN5PCyIN7M458bi+C/TMVnh5z5IqhVGqR3fU
vvpgJGggVI3WeFmMjjytfEhPCpfO2oqgVyupYkmv3sl/YLHNWsUTniUjIYOir7wTQSY25xSrJDm/
JwOHPgeQKErJVMifb1/Y7aWcJtZwdSHUjY9nN8rE59MWFVWZNDnE4og18m7s1WMbkL04PNJAkVQA
q3RSEXTJ3LXflJXBapPKyVltk2Yc1sjtcmFhoeFtSANEcLThGXFbgYXWyY2KsKVlm2aq1JeMrhnJ
5qMA7d3lfBW14VtFS/DG9rxB+cBwwJJ1/4qCgrVcl+RfHFqFloOVBbgPbR275pGhBpJlA6z2zwKZ
ybcQkYTDfpaAa3J9jg3c3/oeOwurGyDd64W0Eq7kT4Rmir5Npqyep5m7oHGnaA2o6ejUM/rEraY8
8m5M9k/KFjasec7FG83BgvLvKSHVaUqhDBy++JJxL3QvQouKXw0B5/ewCC/l/R1G0GDXS9aB4WEx
VtOgsAe9jdBNTLXX8+Fr5z0Spsw3Nj9xlQ+xFZpaQ4CW1QhD8h8u+6HKWO0YRjoqYRKQYcz3QR4P
4m8PujTEsdsYwjsWUhqwbsoOVjA7J38C35nKg6mYr3MucjxbqbBE3LISyahMfBtzhwAOfOi+W48I
Lch1asPRLnWEtzlmXqPm85URl9IMjfDI7DTCIP+lLE21j1qsM+Spi+pFRGOjifLvKqX0QKfcLvMq
AyURjpAHyMhcH+n6aDSOCQprQR39SwDMmowahGO73Net+DEZxEpKvtF5rgGPIv53cNEiC5qb2kkh
r8ISN7oIGLJngY9SWKz2LQ8tb1x3R1cs7luVm/woU4xTtPBpzyWToLHSXbt5yblNvpEpVw36TAqK
aJsH/PeTJdjzzHCrwr9eALofF+5xdHLKF+cJaHFkNZWR19mx0bEvDZy135fpfrEXc/B5XUSnu1CF
8L74rjZofX/k6YEO2dJKGblu+m5EwOJqJ+l2ezpUC6uYV9lj8+iCa7h31oNirVYRCWcyfOp2rohz
TIJ1DL+oUREnQUa7B41JtlKWY7c+GCmm50k6gVA/2LO5cyld9qA5zOMy9qROGpvnHLMz3YrMk1jj
CjNU7ECUeFu2xQQSbzxCL3fUB2cEbu0NLQjNczlPS8CxGWt9rwNO/TpYv7imx0weLOBnFfQigZNi
aOky+D+CIFYIrxFciXg+9Bl1akBacXfMyBN6aRV5mzt+Np6tar3PhljY2O/KCWQ+kdmUx0ydgiLu
lS9NfK3XocFFW2yGc37m2oJAh4dSIuzYGCVZc7lMxtEbl+vqEc7ZO2RqBYVRuSQpMjDhxX/Nzri4
wWbhN2dKxq1qq+oo4Y27pN0nsWcAu6Sr6DHx+gia1lrBbXLVHpzgoAqGP8CXRpblJTYHpUif4Tx2
Jf1r9AAp2Q+sUEVwNuJF36T5gsdzpSlxLZYayUSll4mxlNTf1UgoZsiIPeiAEnxi2NXd7DBzOhpN
MAspHFiQbsvsp+VTmN5D1sZg8kpgJEO8np6mtHUaQYEcty04CVsDo/mjSRmfKmMJrl1Ldso6R2uI
G0AL/OdJZhTyUIZemacBGe9RZkc2bzOUYlPROpt1xJ9FKmERTppvkG0n1hslIJkJsLaHX/DxaVTg
Mh0LBM6cVyJcjMNFHxKurZK8eUH59vLKz5jrsevl2ccg5Wy7ZhmM1/hdFxMU3WqO1Fyfq6gYFw4z
evv4M3OQfLMKdehKZ8YhLZIzPBl3Wey73c+BkFlRzyM8sAhe9aQn7nbb9IUTr559/ivZHIVMpm3q
yakWngCE24ir485+7rw5AoqLDqGxELBPvut9Pto5pbhn0CbvDqyBW9HW88a9de3cab+EQauGcHsj
eRTqwJ/0RKoNneItXUgskGFYqi+lz167DeGGvvvVC2eooeg6yuVl9rGKtgT3vqZxwEd/frPRhs7v
H8PqkKsffbkIKRCF8HvJm35ld1FTAeSCp/LYEf89WMSucWlkF59Q0ZGCSqh88rLOF9p6vzYLWOSi
QAaN9ggrqU6Ca5LSgfyi8YkuuJ3Q4cr61H0hzsLLj7dxhiV1UHdhqvC9ICMi9ysylsMdpqVLjuQx
2WpBjDBaBbsMBtgNIpe4CluQ87KsyLpzBCTjMRU0qDzvYP6WklqLq7++STUcqTiisUADITs6MoUL
n8VpHyjCy/cUXIZe+GrOGe8qKfOJYJjiFmjyrF//HqcHmJcAOZIJu++xpAK9iLyRyTdz+VIJKYOE
uQcVvXBIxTYU+kjywGFnEPbBskPkavXsTxR2KyX5t167sWkICgULVQq/vma01j5biEO2e23VSUWj
Dmgh8sH6W3F8W4cUxSqTUZ1w8OgHdOyJlmIodC+gvdgef8CikAkLVNZH6Wx/HabziBKVFAKFj+yR
2fNwbnPxmTe5dcT79n70H7NFOQkzN8g16QNaMkAY6uxizZlgGrhTktD6sTFRAlpSotAxa7sM25c5
nQ58nnD0dbg7MrJ7fSNCugfJ9pDpublL5IsG/hBwHBc4mTqByaL6hJZiwhd1em14IvRq1sIyfww8
vnvoQCv5/+/9AOghFqyR8zcFinCgrMGYVwe26oBDoBxIQArtnMCYuOlAIHvwlA+0OYo0Nlal48QH
k2u7ZmIGIYEdhwYKLADfVYIkwlghcID3hVNjUOybeS4zxD5O4M/am0FPBskZF7uBXuXqPsajdTgR
u4RBQJ/az1AtN58SnO9K9d2BObFtbXOQ6WFa/EiYNkPMV0hFx2lyEryfiLSGmJdgv4WOS0f4iimW
ZV8sTzt3dtYCg1xotUqSvy/nGZ6elLeiDyRS/7g5lRkxebTRg2iCzJRlqv7myb2mKzUp+DYqDlot
5AcB5imdE+s6+Lky3mhaWcNRCSeSlQLoP6bY3sXQT46NXUDqbHZi20PsPznOOjmpxmrEIVQHZrf4
1JcYWXQFSUo+MHSW8U9K3u7Z2TgSns2qmojiObQEeRB1v/ig413QVSFZnynR90PxjMjyQolONsjZ
WGFoUDQEXTqxyvPgsFa3iccXDYj+gBa7eImfsJISh/LNRFymE3vRrDgEQcD9UgR4yxewULhPBo/k
zMRR7B0PE2OfBBig3jgqsX4ySLSi+yx2W/onqtJx1XcG7SSafWyeGWSa7iwrX09gRgOjl2FJm0CY
m+p7FSj9I1pxZcJcZqkSOC2R2DbrDf456ON/VIQnVB5+6i8sigEi7EPEt9l1Dnpkl4IZauRIAnnN
hAB98Bs/YW+pIOWDcr4+MTMcF4kJ6pT13BWr9lxszvZSD/bQh7bn4U6vi+KNNTqOrHfp/DjBGS2y
/FW7zet5ZvPPi2QHRhDz0vSllnIqgnmYmKhfxH6pIdAEa6g+GFTlAdM5Y1C3XNOKr+Rb5WDvkBIc
Hq3QqyA9T9XrW+PnuWfzBSRsErw6BBTf9adMEao0tUjdR205Oxj2RpS0AIbWpLYdc5m4D2/4L3cE
A86O936pko9lxrVjF3qk7LqcOI08/iIhh5TN/eN2yVcdIPntzuUcjoGTRLsDPn9m5686SgVsAH2t
WP6Z8eV3vv3aET2Br3YJ4egh4CcsOBCZKBrJKEQLzxs7LgvJ56PzD9EnQ5fUFceNKHLa3k4j9pf1
gAI4RHRWgszdFA66wwSQWCgdDPIXlnaNh4NK+ls33MlsM6SF1K5GB33YNlOD2KEMe5nPDFvnH+Z7
29dOZTiYkc6DNF8ODHiULkH7XZiBK0Jqyf3EOrC/mtyLtI7tkVSSFwEOgYptZmFIsn2KUaXYpLco
uv/2kemJGn2mGCnfQrgYP47NCn/fTtoXB+xpx8BxvAnq/dmnap0l+AFJDdtCQlsABV10qsLkpjz8
Dpbjm+vBBZiEMfNlx4SeoRK0ZjQ8n7HHPn3jAq/7FN9PixiH6toe1CqX89QylyrgDAUb3TYJMvuJ
KmtsXZg+WVHMer5/Gx5JtQKDhx3m0Yw/46otD1OrGaFXpkux+J782550KuD2NxbpgfSbGICOe0+o
FcLMZL7K7c0HD3GCWgIC6EGdxofAV3sZsZm+Ti4jGxRNPQCU4eIGLLWmjCkCT12tB7om/YneqSu8
7YgKMsWslTSduVo4sRHguEX27QiiftXdf5Jbg02tslf6t/w49MHgRadDTttwWMSAExt4GuH0lPhY
lC5MZgkkGwFDUe3yNz3W2ZReswO+KxtrFu9eLRENXuSfhx4WrxgbKlAt14KWoTPI4WG9DPJnc9TP
Nj+YVdjzjNNNsPWpiK2+JmFFH5hCs9wL6zVlwiPneorexLp9XFnvKIYvVpz84+VdJ9XwpgbB+CPP
McSKWYnue3MIWJUFITgmxW6mtVZMAS+gecwQPP2Cgari/FN+EVEEcG18BcVDReYrHZQf2mmA/01L
/cOHVcHtJoDam13sV5ovS2zWdg0mYqPzG6djSsgtMaNCvBgm4db7P8opRwgojVQHge4ap45y+OS3
rV5W6OrRP99hdDVHQNuu/IRFUli1EgxfN6jyE5DUsbL3A2r57XaKUZTZBXtJDhrZM6LQUaG5QkXs
yh4olsq51tgEB/eufbJEgkA24timEGpk7k3Kvu7v2RLoQsvg4/oNBalH7MJTsiwerFHQBtSlA8Q2
zAggMOmWnF0DF6OgeVJx0+1VMRTH6e3tOyicDKdRcQXuI6uqoOnmEgoNDdnwijSszBlBU0p/ce1F
uv2avXz+GMVAlfQrxstu0pDmNenX6arfy9Qfw/bD74l1biMG9msbpGRI9wP9QMA63RNmxWi2gGx9
NNYs9h4naLt/gbgGumbf/oIBR6tqDXW1L3SuQEHNduJE2aQA6SK5lig43t3NOsjoinIeGUbt9jy4
UwAyuCmYhmOwMhqHqD5VsD6rrKdM1eKmOcX/lFYNngnk3PUuK3ddxmPuRSstH1vAymsfutNdPv1e
tRtTHMy0ZJc2HA7WtpFJutHCc9t39g0DEiQ2UUnJbHRAWnTh75KNZ8ndlivXwoQS9q9tE+InEXMa
ZEC4tP6HGjnIEOkPXu7JG2mtyMhQvNBAbO2KUvUlnN7ToDokOH8O3EqD1WTGOREdhKvasxW+Vtc7
qg4Z/BsiixRzf4tO+NJQJOZlwzSPq3r0YDnGW78nlBfc7Hel2Cs//v98ne4v+aWXslPgmJEKIAnT
dimOMdLpNbfS0XwiPF36JuhBjp0UzNXUCleWRED7FakFOeGPZmMnZpis/jWHNzkjz+giL5JmeXG8
wL1zT/gmf2RxK6y+iJ2qxkydFz2tAjCCcxnNeA9fDvziVMKaTeYKn1hW9FH9hcXgxtlSr04fev1d
IgbJTb45/uZTpNXaaGguzC6d5gUEzvka/0N4qxdXgPfu4Z9jVnPwyGlhx4aE54w/5/5aa8DlQmUe
GdvGjCj+vExT+rF+pYl6jCswcWtv02gzTor/KI7IGU8t/mDFI2AFErMDsLzvwKdEx589iqsO2Vtn
vwV7TB3qCy8P3Abikwc1CuneUUCOrK+5kGtcoZdKlMx+bulfdgD8bNAclgCJ1sq382NIF9P+krAt
9l1jaPyygAcPtPXW6F3lLzXfScUDEggX29+AYHqnwIkGXnh/1xaNF7JgeHudaJrMXocPatbfRa9J
eZ4z8YoxHN7cPm/gKzMZVMuvHd8ULFq5KiR3V8hjimtcbrxyPGgr/xtng9/zvJQ2JTd6/ghE/MMr
iqekse9tb3S0gKaJXQd6YO7cRtGGsnsD3KBARNjNCuMl2+tsWE/WNkTKfAgYR/qWn5oSw2VI8033
9HoSVMnf5K3K1bXixzj38soFUvL+IHJknulVDdrtt28Z00+DJNElNl1VQccWEUjPGYq4wpebNVR+
3C+gdQ3iRnFScY3TRVjfZOZu/rJDvmvtllyMylIy9GKE3FovAxS4BfsBUeg0C5ZzdvC8pUpwVSVv
uP9ksVQEI1yJXGILbzq0aBV8sAZTwvoaiFYr2K3m/JtZLgzRTURZaxcwykRtbQSc+8gsKDWDTQrF
LRDGL7mxgJQJZn+RK5BktEXg1qxgMzMinKvJnvGrQy5M7pUdsoi7PAHUECXMD72H6IgPkr2R4hXU
kY1SbYZlFX5+SW26rUuuNsqcItVErin3P3USeAFPuBr8jRqi14ixY1JRraSDDpdoKtJa+uiJWm9P
UBxYUf76mgp1hcC83QtFjfj8V7xAZiigtJQijAztNUlU1thHORtUnl3WALigWpzDlwxnEOYhmrYL
mokQaBF22YvHjyBs/17xbUnWoBoHtljJrlbIyiuqpX6n3zuGXNfGj+7V7EnnotN+qV2e7nXSeNJG
ZJV5EPC3vl2w1yFa52LimAEE9hKlB/t/6d3/VjwfDMiD2nf6nJJLPgr+w1hac74wwqXoLtT0FYtZ
1kZNHM7yLHAH479fCZE02UWvGKOzjd6Eqt9fcyU5I4Y6hj4NV5GScXASr6z75jcnVSjRzhgzLHkP
eZ9cX8ca/lJSwpUORTjIycCp9l6zFCtD+A0EQAnxAP8QjsX28lGse/re43mh8UQfDfyTRse3QSQO
SZip4yRXnP40F4K1AK0oc93wEM1sOJ6DvUc0LuFjJHknlTNK728A7dcJZN3RXu/tLs3KzGyvDfvb
9+rJPPuoIzGNbarntAjdVen5Hj1B8LRIZA7aV0ssW9a/QoCyqsRzZM0SSWh+GiT/76JOo9bEkL4i
r/QaoRvqBKx+374hqlnQaIxHYQyRU/KegmzPmj7LQt6cK8SB+rilYGNpDtIF5dBXHeIQMikzA4kA
IgnXZC6nGL67Gl+jRVNBy/hUAkURWdQBVAJ630PtN9D6LUeXGYsBHpNQcn68Q4x6GsYHel7pgVFK
ryKBPSrCiwwN2tVBDw40KZAp4L+WHKCnnT0sS4e6HHq2YzLDhShohA/+PKc4pyZrYnnAotx9Fhfh
EiuAACYtKWzSlVupov4+uihY235d6DPtpofFvrP7gzS1OHQeB6V3NfxWMm+F47jQPZ9Oew1SJ3ue
kbVuPqDRVkr65FuRnlWUVGFTVYfVYntFIg0c8QTxdHZMfqI4v4nWaSKQ7MfTRcBrt/e2pwzXJN8c
a2LUn1Py+qa+bTQ2Djg2TbG1VjpBDXy3Vcd99/++W73ULpgpbJv1iTRm+QKqC9C9hLL9MQFfGbxg
/dQas2gZ+24zPH9ME9CVmhpv2FoKRqZTIbrkDLz6YYH5tlTIbwxOfytrCRECKtMNhfiAmBhNadn7
kXaQiS7yaok0DzH4EAiVoRt1bbun43D4LLBUULM7dTO1SS5wSkE74/WU0yuuEzwfF8yC5l8eYoXI
WblBQGGkb5I/8yzzJTUftvUeys8l5poELbotf6h8lpxtk+f7uiteHTQzZJ6Fr/zgY0DIrs4ZComB
yGDVIyrinL7BrHvhHbaoOuWi60BgTW6D+7LJ3926axvGNV56VfwXpBsEj5rlgevyn9w5Ca8BVz3t
DkVSLPtSnhe7lkct/KIG2BewwIAzdBmNeO0vaO8AH3qTAsKRKOOWT5z7rlfpabtu0oEyXDwY0PHp
dHmVWO2Uf+n0lVpdN/3ImYP/FY4AmNNs4SHPQXewpg4UnpXQGf3fQm4eXOTX7ykufrclpDcacdhw
YzVDxY5w4mfL5UhvkO6ZkLf+WRRd7Kh+rZTYkcNZ9PK50NHqP1ZO5ibvOzKkzVmVXJYBlO/08UuH
ezZ2eFDThbNn7BBPNPpGzto8kBr1bMLWvqoWOZpTqV3gKIcnTSPYY/AHkmQ2v+gCEZ1T+AuzObyq
O5fx0lhUgVs79w/TwvGvySgRaIU2Peq/fvPrwVfyTzEWwlUMyn+fC2+XBqL968/HPUDUClaX51V0
8M5742XDASsJUb0Ic1NtJSNf6gyVbxKnf95ESenidJWJNA4y7ktferlRzpNN8qDEcw1E6nfPXyqa
XKeoXEWjqa5ztPvzmgHmReo876j3Hf7S4l4k8EryO1UNkNTgPbthLzT4DH0hy2Li4fRYxk8tTFuh
yZKP1fy6SQeeI6Mcg+fWNsJrINLgE+wDbrA9udJKEhZtEZ9zGiZhXiXvHEp6NGchr7gyCs4xKXl+
8nytaFzmfuwgI+srnZnJqjJx0VUc59rsoWAdPkDprwHISHCfvwvggvaCu6oeSE1/dortEQ+oS7eK
3iOFcseXXDgrx/uC3jt7O86bIiVzAIR0MnC3RDm+Z+dOhbUUNjdDyIyAHFtqeoyiALf5i44ZPGht
QmTMczzQ2aWq9tR4L8y7gTxsB7eKM94IX9UPz0kB/JK1lUvj7yrXpUC9iqGxSsgI7OXWR6ehMAjo
mc5sTlVElC22is2pq5LMf76nZqI/xSiDu4najBoH+5R8u23XwF/35hImj4EcT6zJH6DNeK2lOMkR
hDOsGDdbzxCB0jRyEnf2aOTDpVn2eBZSfxHPdb1lywF5GTT2GzMrA/Uyo2GJBr3fsO2ZGqcoSVAi
leZcqxBwbT46+2kD6RIFWbztOevmU1WlTNVanIKqY6QwnmIdz8P9QJmf3ZnBO7STopkaQgiZFzC7
NoEOcdvmnNfdCjcB+lpvgyroAhXeHGsCjnBZs6STfQhUi743SDy91tDmI7q5w570+6M4TF2cHtWi
xcb57NaUmqyakZNehbSa07XgPvsq2bte2mDwS2eO6OJYmmC6RJgD+W/tOSrOch79CeY3++cF06zG
lrGcEgaMU3nKdmLP2ug+RdHqyZU4fstB84u+lEAC2ISmTgL+qY2PYLBZNQpwCFWxZhCgo3KJibnp
kkoHz3TlZIiF6iBf7K1Ydc+tbsMy0t9TfEuMPYHpHKuWTrkCNNbhFoICAQHnLqR2vCh0MTJUzX1k
WUKgiWfAUat9s1q8cw+uTmJ62aHbmErqINj2gOgbza41R27+y9yRGnfppRAU1RmfBrCiwDoz9PBT
zCkZht7+2ES0JfxBBUBi8S5DdUf6qbNsSw2LrqvqGPWu78auPUrbfRXaHrnpLDfqOGsxgOXtwsVj
F9NQ4nOhL5vkMzns5oJaxk2NscZIKi9GLXoMlzMtpz4Lv6QMzfbVhtgLJuCkJC87NVPIecjXr3V0
i1fxXaSIBJh1YNvOUMb8Vo5GhW/KCW0KNd3Xs+MTCCtjKfhsAoJ/j8gHjxBdHKpVrnsfLmZmbD+E
af3pyd5gfC7eyan/6Q4OjS7c8cxdPwopc/F38lHY6pCa+rm8Iyn46TmA33Z44KeIdYRYTlYNcU/z
CfsM+kw1lM7x0DF0sXaUTz2HoFgUbLHnf1UyrcBqgAe+x02Ap3okXcuOo0dH3jtieBcquKBfLvgp
1s1kJxSBSicoCEXINl7qUDaU0ZHjoX4je2KRDUEVtZ02iFKcf4BmTqQLokT0NLhXfLEK+xb9P3Ez
rbE4EQBQb2IfbZfokFrfaWSutVNiuF/trsHz5bYUlUk/p54BcfbLQCZ6vFC3dR7QHlbQB2xIgVsn
XRySfjrberlHLyphdn1h0VT1BNLxBf+N294cbbO4bNpLwewF1cipiavnHfAozkbWQKiL+PG/0E3b
q0Ov7wzFT0HEx8K6mNWUYxG/xerX196RAR5wu4+WOtj/MUsJ26ubzlyNILbW8GhqEU8NnEr7zNzx
hy1785HHMd/yZxxLB2Qoex5pF6KEGNJvPRGj8LRH/ZWsRDNcSNakinpM04Ln/GMX5RnjyJbVvhE4
jXjnn8cesXmQOzhMg2OImOBv4tiE+Tvqcv1/4q8Qv9ByIKm0TCBVJ6YOYuRxjMdrT4hiT0c5zXA7
NRGGSTzBAJ7mXscpmcJ6UYlxcpKrs7U9P9muifDa1bjZ1TwC6IsNp/hEIBfikqqegHWomNXz+bLg
vCBtstLjIzbZ1tsCWfViAgB0+uPE7h+SjuqY7LNwYv/KxbzKGJA4zMrb1wz44mfZQ+flFHZqyn7z
fyuXzLrvINXp7rBgfqhUObbCj6zFVNPkphCVD5lyihTVHqOZSSbJtAtePkkMGL5pkf+d5r0MaAF2
IfgnEc7yPpSoSG9NXUMAxuvOIi8oDbUSD0qNDxDidZbwGOG5YLt98/veXpupedM/M2bsrd6TKXjo
qLfW9gq/81J1DRkD8oa/pOS5LH+58eSk33jqm4GgyNTG+ODlaQiWnTxz1wp+EcRGKUxnRvnSNohL
s5KF1d3i98Nj6PH0Q5+D6TTFoNo7gh7tqT0opFRaiZt8DMqv5vIaE449kcfbTXwTbzWZE1LAGCpU
o4KfNscFXqZo4LIwGqmK5X1CLfRdsLDcBm3OjLz7LJG43xzahWpr57yP7qpg0RirgNX+FJgyrvfw
YayzZ/M0DBbgSSQIx2STUIBUAUzYuRsayjHzyzSP6E4pc7PKvRvtN/YLb+BfsP7Z4FvdDp5tnd6Q
lE2PRYYjcwdCR3ySNw+KvyLVHK8t0KLw5/Z/0B3iygCkUYMXrerfSC1mvGScTHe26kgf3Zumj01S
mT9WF/Q5SulTddW2qPjnHHKHehPIErdJjg4U25AYhwLfsz2yeTLQlo7KYAxU6uS5c+UyFUt9g/j8
6DTNtBYUD/4ywHU8fl0fCxtzDbzJl0d4wymEi8+jhRDqFoyN8dA9IlUQCK81z/TD5TpW1V2C6B4r
7uBxTgSCVw5J60sF0GBZjNpgI1WsnVLOCm3VYHEpRoCubSUEdxujuzRoLxr4N0NwYy+sYkf3HjPH
h6zjRaCEQFffZrIfRRtDU7wOmVFBNJcMVkDeoru7p2FfZ0yr0Nr5c1jT/8wf1seMxyBWjt0x8mZS
j/o0vemaBpVqxLPz/SzkYlPZ07zGw3zfepXwVyAMmlllVxa8viOlHFjK1Sk1dRorYoamj/GbnL3H
C33h8BXREj2TB/Uc49qVBdBQJMXJCw4RfrI0/ubXoYESgl5paV1puModBo2eqIoUOVkJ+kw+d5qh
JzH60MbBZHjZZPu0eQqUeLv96e3cTYQ2mL0Pf6wdaV0rXLwtzG0Q0ye50FVvynIIIRc5qPD9J+G/
djodBuYYb/lHJWUeOkEWv2/ypBXmMMe7MJrypUQwziRolCaxyv3xoJXkfqukjcpSnRDzNt+MfQoX
+u9laRVpyhg78JVxGUYyjAFXyWkzPN4+XGdcxNz+2Fxvh3HI1FCcGIq6Rui3d0ru2FPmsV5q7G0K
mgF4M6h+SGPleDDmWvDXqUfeUemA+1zZtxRzs0+8wOiMD3/01wb17Fzncg5v949fEtFChVMGR7sV
dip4BjjQiVhImv3P8v0EqCGhRLPHetNZ0JTzekef5/wzlYTVs/yCBZSTeFt0r8eFJJBMNrmyB6U0
pwUD7Vz2fEZWv0URofg6Vgng7NmkWD3saTHTTD3cwJDPw32wmRst3MUotdGbRu4OGnvVtrYOpPmz
kkc0ieSgH/uzk6Zvo5aw6X6yNwNmTUyFAT4qGmpFGcPz7/H0/mgMGQDXEfCoFOeJTFo5ShQxUzWb
fSiE6eVs9sPMuKuddW1n9XWkwl0W0Lsl7JpuXImVUdxBlB6+2Paq9FnTOqQ5eBycIQgsExTD+EuR
PcdQ6rcYdsonTolkhS80hUdfaVMud3Rvh2zf1tpDThtl2avoUFCMAHbmCNzRQ3tDH3R9mKmX0kNb
0yigfVVTe5JRMmySEcTGEyRTqHc6kJqSXzgjzg9rMaFRY9XT7B0kvJFYWJuoKw+bIZtDNe3Yz1J2
o1kMijs9Qo0yCkGLyATJBC6xji1FbV72FYbMzqF3bqf9ekLR94w0j+tv4XN9OsiWAAogNkgdxOv2
I1CoYDLrgXdhPCuke+dfq+tusPxKrZRc1tQZqaNkBt+k+3RhGyJtKtm+MrwDNapB5i3twp0kROsq
t7CZQPH7AgLxGEvxFJbxCWfHNi45B0JBWZ43n0T37gaOaABATcRsTUxzc5A8vUnFJXGcTVaX808D
z0xJr1/H/m8jwfymj1Wa4YX+4/lUMYxZy8C7JBMIRZ2PioCXvTMiKkbCNRoSyjMdIsnYX0KeM1D3
H+foAH0Fpsp46IQ5+WG1119zews3N/a0plTHNJzOq4Ilwmofd82H7+PzvBJVDQUSWdiAqPFUYRdW
qQXJI+hfsUSPLBI1mMaJfzWy0iadvYyN487mZbFxyHSgqIB3wJ8H0ZaeqRN/9bAyu45Al3I8KhZN
muSg5YMhKMeHknNIwUO2GwQf14f0Wcd+V6IWz+tsZ+ElNZVAZcRcaxDhJIfgT1oJQqEHtu+mVCKZ
xUOlkOpgYI1uvcgIsD9pHC20t5w1OihKY0VyD5YPoeEjvHXPkeiDXkpawGKOtIFGGCIzr9bFr/4S
ydRKiwl7Fs8p3MyrOSX/nzHTKYlwz+ndXZqmsluH5G7pshP84L7NNFM1ao+dA9XsJxbPRXcZfTRH
EPb5mX13IZkIHz4s/cMaPUbpORWDcxCA5jKeszkhfqHFqmfbvm3C1GUt+7/wfms2sqHLQAj7wBfb
idL3TQ73P+GFn17+aHwJ0YO3Sz4F5fbLLDjRFrxUdknRKOEJgHB8W6w32Ch2kMH5t13ZG8lpF9H8
VjaaiEUr9pBqF2nWEcHYn0Sh4oK7ks4ezz6jtPq6w6Zanc82Glsokorl7h1ws5O5ZrXSOk8DkFEw
Ym1wMEE6zChXntjHlTfQhc7ybtpKk7tTOrTyckOpzlIhrTpz6/LZokSdu2DmXeuVRhoCOtKyhR1P
5aiRnZNLionJAiMeGOlZDdoMOgZplZt4GM25sEIK6mf5QxgCxjmtfuIToCH9g4eFJdnthiuBBpLG
ZDJJueqHddxxHwYONvtUee1PFZGAZs1ZMHrPn//3o9JogMSUyOXUhZgnGKOaRB6PI7xx/JhDbrwz
PFG8twViMv/nMlvv62urGzkcO8cCA3pfUk7ZQE2w6hitWQU8UE2sfHMMbYRf8xYJNjBAsOZQ3QV5
Uwo8b609PwFJXpqZBw0T1zVcqtd+BpEesWGWDcfsYu130JgxLzk3EbHaHXPs9+/t5uxg5UB3r+AC
++vZFHjdBisjz/VxQx9pIDSeTCp/fS2r0WmLIu2Z5xuAZTrx5TqEp0xUcSCgXZjW2OJUmnjGyS1G
AtQnXE7uoo+asL7rqKnHjYJx85wzBInBIqmqGauMhRrEfy/KnDpq4BTzGImtb1vyrznfdNo6/U7Z
kKFTWV7zSJfyUCf7nnZoiQ3p2YNaEFF3RocdEziRu2XQqkHHbhUPpS75QSzHNdURCVMuAJrRsO1c
FVgxlRsko90fF7BsmrnC7uP/KlqEXUDgZsw7Zl4MaJSqDsieOPN5grcDG2AYOtJ+kga3fFgy22+g
hwMx1LebenbGWm7oYes2ujJoHJPeN5AaoZrqxRVL6ORNVwqQc8+aPat3t2hGKxSAkVsA4N+gLMDG
g+EW27lRp5V32O3MVsAYILv02O81aM44U9MWqIjdSPSPqT3LkUAcLLNv1yrm5Hwg7kAioIEtdhDN
t3ShDzFsVPeLqnHbM/Ea+DGyyusCVU1HPbh3+T5q9ar2sBBJu/pvSYfQijLLO2ozRL1hbRT8OUcY
4YOf7Qt1iYY9I6RB8+ZO9/AmTvEXLHBiS7oyKkucOarjiBA94if19a2qpWrOJdDq3ISaA/tmtJvi
xqKoCGAi+jusU5i45nbBN2436QH8Rxnyl+wPeLw48HSw49LWRHDM/rxk4Ydf5nrjMilqPE5BidCF
KvK8qBYk9ggaWbfYJu5oeqgZ0DGV39Wq8Q9hOP9f/TFCy5Dy2vZrH3LkxqE7eKLyGVV09YYCOrFz
rUVS760Viq7Uub0ehG3TTpcUIvjdGL80QapOSDGB9wHw3hul9nioQRUzgKFT/KdJmoj09VHv1Ecg
1xaKEWuxIcvyZq3xhckqosBYH7+b6QzgeHaShvaxzoe2jehi0Yhmr3gpL8gJgZoqSZBeRQyIkiXM
BnbzS4IGln5M6mMOKTlXWfosJE6jDg+b6XnE8WjAvjvEKQWxTJxXD4M1ExmByC7waDNUpDI6lDVz
Uz05DuDjO+mbbLrrM86AAqwbLkyV7lXvJ4Aqoo+2rlLy6XtH3nlyQ6iMGvIihQykMzxslb6/OIal
bkW/vFsZs/LlclT0F6S0WT4Iy6SXAKf4mWOrAva8fAxxHSdebT9j+otCoiuaG705Uko2lolojq6s
k8wwkSRjpADYZUgEgp19YMNiD7glLgmA2b8A2A2ZeAw/RS/evDo+jn4o0B6OxF9nCUWvon0duuNw
yLdmFZ8qn4pz1YXuiitjsoc+UYN5ruuOMLFRAOgrlF1BBFiE5Rb0OzycHuTxmFP3rnfd0yBTlNDk
YbKXyVQiwZZgnzGtltpts5d+VJpwSdl5vgJu+V3swSAWMVBrBTyJGRM89zJikCp7yc+ZIHX/elJv
9GyeyWtCgI5uklsrKwPiI0KH1LdVfFRZl+6mUO5YctGRZj19VIwEqCUtiD6EkPAvZ/OesiRUhzIP
BbeLfseZVVtVPY50EPcC6sa6PYLt5Vr4lc42E5RKECFiWGU1tJSe2uCKH3WoCrBxL20LpQMEPVeg
tGmtcEkFPdWaAF0BRTpJTKmyDMCeupIQn1Ug8EmP1ekbrSTggHu31O0Rq9OibRqcONfAfT7fDUUc
YxYMLgeF78DHrRCgE8h011S30YWtrpvyIYH/RNZor2oYtEKVJE2ZO3y7dGuc74flOJ82FgLXJ0xb
eQ00S1XExMlu9PM63OZcZJLEonZgNKMtpapmkgAd88AMRh0VrgaoD84mWFKpZLtUU3T9AviD5ZhB
VitlFfbYF9/lR063+0pRiDrEHj+oggOuunO449m1BJaGBHw/aY6oH/WxHeum6NYRP3vAuAt/ETCO
Cc6Amv1qDsTVjSthWnGm061y2SyQW7cSy3wAX1i1wB6ri8iwver0G+Aa+Rgrjy1Y4V3w/wpcgdwQ
QMvg9cE8GGpury+ZOoy5RQ+AnekSaBzz769ET2t6I6WcTJ6g9MZrSaRYe0PFEna4tUjUkw0S6rVJ
hIlWM4d7HjMzThqPIuMuVwwh5sIWrpEuOcjtVb/B6Ka6wUz0ybG1Km9PsQ6GsCxkU1x6Ef4iH+eN
hGBlFnkPFBEflzsos9Ot1aa2kg1aJ3PPvuSw2FqDyD5/awuJ0ICiVUh8mVSTbU5mXMXziOZvfn9E
jPcorYy3uQh4pWFdYLSklYSdRI5UKFKB5TAPzsch+TvGM8vUOYVeR6rd4NQJsVcRplDOOv9w7Anc
IovWzaVO6vSFHQfEvhLjlRxK1Ec2p/noa+C7EpW2nxBqzrku345L/MNogRhZ/PmZXwNgY4Dj4rJc
O9PUfQgFMejfcVh12vFgt/I47KN0Xa91UBntQc6vUhuPqB06i12W3n5kYuwpk7CEcS6WeieQf47o
ztZgIg+/CTbugUQz4Tq3vxPX4sVVsXF0COm/AgakdiI7vvSXME/m+Sf2HJz3wRBHI4Gc3IJDmHnO
5HZDlWXfRFRNf6d18TSZLF3qnFyjhv3i2i5zn/5v+DPah2jypcH7d6qRQlNPqrcUc4rABBplZ5to
8IrFFIM0Uwir56a+1/dAH3XT/HNGTmZHLUXabveiVVjA/ntAk4Q4BR4Y8KYFwwNVY1BSfyZckiOO
ZbGQYwNQLGqpMxHE67BFhf9p5EeZ/qhb0Dp/s9TZLLEB6phyI+nbepi9IZunnxR0mr4uCK+2p39p
UlRKbk/8ZB+6T2EZWoL/dzbHCBX4FXttq425pESOAN3G8jq7CEuYJEWPpOvHz5JlYqj4dzxX7k5p
MpOTawXB3ZlYg4evttSQENbehFbbosAOefKZKu9tGxE/EHrY7Qf7jYCnwn2x9bQTBhlYCVRF+PcH
9xIxae+EEMMmnifaUCTmuZTGNtAgLces/pAU+WVNIuXUsgiHUIwycoX5LnKshpkECNQ2sxqzfR52
rrlmG/loACkrSaBDnHs0w3cTYnmFL/0KsyEicXI+obq7vH+klMlSf4Clzp43X2yXCncz732tvz03
R4Y8HtZXeCDT80CqQrAcLjo8f3+a7HxwuyZqyPC88vvei+luRG12FX3GUs9VsY3u9NAs6P8vDckg
JOPEk3fDwmqFOQL9rUbrjL6twj/w3uVs0vQDqvV6x639nAk+u8XPnMnDybFPWbTpZhQxipaLZGAi
8gwLLKi48JJPEe+yndVDcmESv8yVw0na90rXTuXHjyGw3x4BWnD+iUZ00QVPcLwXZrbBh47vbKFL
dDH+oxjirSPsZQ/RW9+AcdhLdzpqU+e2Mp0XVqh28r8+TabjZBqdQeze940OwTN0m69h8vmKKpSZ
nMjtuFRG1S1A+Br5hG+6YD3Rw2xSHOo5EbNISZpVx2YlrZfGph0dMv0pJ79f4a1bL/vXgHO3WUBx
8Qy3jPPkFQfrG2fzCiFn5YcaB4RSBpUqIK55AvlcniZ/qLuQGsUORfYuD3edyC5/znkdhssZFoz7
BlCLSuUsHMH1nvFft+dmptMCDzmfMvvqETsq1RJnZuKfv1SvZOp8VPTKS4e/1QQE5p5nYXpVQbHf
vrh//5LS++Y0HDOcLjDY6dB9Rcs0OVDgC8lfhNr3Fqk+orEJmioxTmGWC1M3npK8OF19elXOEZb+
IbIDUCCLVDBcfRGiOSCc1lacdJkTZSKVaXEcrTZRyay59F9PIepPRoNkoX2VlTnCcuHbnd37OBOl
bVMqiR+C7g6J+b5sFhd6tkncRvhoNrXXgP9/WcyJbPV3ytUq8ShxYK4jL6mqnUnPJYoWwe+SG4oK
wcT5ePrJcGtz6eRtInqKoXvYWzjpqKdxh4vjzW0efy108rbP00EQXRvxMqHMA3KAKEs1G9GHsgPU
mH8rZmDN/yu6Y8w0vKR2ivWY2mnk7BIKYS6TMWcNOYjSRCGZK8lVkGRNq4LcPljqx9+yiswiEPRj
VDhSk7yHVJsKcQ5yoSHyshboXPbr+FeW31Je0DtTncehSSiGb0NSJJjC+0NwhpUYt/spN/Z9h0of
gAX+qNGin+JnZfvAULoa5dfYTrSeDKjM+g/9hAwQplC5fmF4IVGIvhxzPKyFLYSAsXE45CZI3MLU
S02gDVi00KL0s/ORUuXrMYSP45GO13hlaaSFdYhwTxcqFBNDnCGxjQ6v0qxIFvD4uZM9wgER/ibk
ThMUSfX9+kgG85Kc649kJToKCjsZ6T8J9jxghM4fMCF1ueWe7WDu6lHMkKbj0LoVuFQlEEYCMLmI
3tOxm8lRvaEMKIfzUuFqOLDCckQyW2+q2iH4R10vE7sw60+ikATo7iVyWZIvy7T3ve01SDRPvocE
k7EyFWwYFHMpjK/5WRcjXDIUbIvlJMRZny/hb9W76ZGf2k/JA4vm778sOzE3544YVKvKoS+oR/EE
SGCNFiEURYLJUyge22gQLcZKgPJv43J6isDJxg0HwC56/dvqolhJzOUGI4MMnkvNsbtFmPOMyNus
JrrP3/WRnFKDtMawuSTCFCdkCHO4NQkW2HPVdlZfkWybDQcFNet4jFCJhxbFzeprTc/51Jn4i0HI
DpLdk4abUREHc9HL/g6dFk8gFjGtSmLZo3oOYDTe067AJk7Xw9aZXocEXwD3pGTk1yk166rfx+gN
0V851kuL8TZMIYNexFaN9ZmhtRI6jkksg1+I86mixHoPSiiyuViee00J/8IKRUqc4ZQElowVh6Rk
FddY1zA+X1Y7Z8CwwRL9CHb9W3ws6z2AuBMlpg6xpHQxt8lqFG5sHTQXUDtZDDxfHgYS5TZkHY5L
MwF7YZ1eEliwyyoC0H9ExHjnlyIeLQOvAduvTfOoUIf0HFiyEnpDjdLsWwPt84EEIZpgkiUGKeX5
XugJK70/HkqfsfPOXi0TD1wp0k9iZyHPdRtmo0rirJ5XpOwkvr7j8x6+LxkvH7ejxEjE9pxonlIp
HSZdpxtYodeTGP06c5K94kY9VB2zuFej64Bf4jRjI+vXRx9avyAohvcBdTos4dOj63nZXPHoiM4t
U2xpXZcto5h7+064gAc7UzrSUU/zqj3uOJQBmyqACGppInyMH8X6o04gX66w9Oos9eiL3GHyTUVj
gYlm1uBYuUOv7+bbrjGYZ5L3VShXq/zvPl9QPOT2ISjjG2827EhQpyDgB2P00dXLWdUa9gVznSiy
TxgLmeh5Yu9/KuW4r9F3KADfMETT4bpFU51D2iatYGXCNKq3H/pgJqARq1dCw+GHMnRnNU8ZzR4I
EVyE/MzRMHCc9Ikiy8PvEQuIm+Ic80gsaC8rxiI0QtbUZt9S7O6/qdm+WYF/xLZ4Rjq2oHwZGsdV
F4glOzX0RacwS/z1Om5GxNooq+CpH7zuj1M24uAvD6VixDa+ZDed8fRRDgcaWaooCFt3rSDRckEh
Yi8JGPKtIMKIBATAOVbtyE+Ew+TTgZv12Lu8JuMDlNQpnKe7i4kSLDYlQDinGtKDcV9qdmf/Ksdx
/mGdehu1nFeIfOSCuUhEhg2NaW+1dwHggp1yA4+9fAqskueDPtTIWxevxfhfDl8hsLnhHdLNHFa8
RausXRU2PNOL4Jv/eJJch7Ot9YWE1KLEzJb9Qa2o8YU5ECyZGzlDkibHcz+5Oo+AIpVQIHZDbvqg
1mk/7FfTbcV+l8ImSr9T8/CrbpZmMX59oOszgQRynLlLLIaW7UxpAblES0ILlaS/Ag3BFR8LysCK
TVlXt3jdhW3EP/bGOScBp0gUlbtsgDbC0L8LPMhprDoLOjw/U7QfRnNKbeL4l61vBBqg745X//PN
BHTZREYu4UBH3hrj9CKHml8un0yQ2JEwVOYtErSbkEytrNx5XjBFVQRUhn/xLUkHCeTlbp651Iea
RM5sd0MPKRzrk9efytAq3FPQC237vF3wbuKNT/Yl7baE//uaftrPTzDjL/c7wxUIF3H+F9KFurBH
FktiiNyg4VRX9K7jLULDp2HWSHzj8/R03BwsvskwN9R62Tp28z7oNbXt6PTmUYE5EATWZOAEQhFV
YeAyZReCJ7LVvuCMIiRwEJVJ80jvi4vLhX+3uFbzq/Y85IeqcurmtrZnlbO+U/G+zmbG7iC/Zhvc
WVimmJaYGw32ytra1QhiJ4oJvPyKKIcPffDrIcOAoVo9JzgFuEiF0tdICFDe7Byo6zxIZmV93ZAt
/c5K36/+c5IfCjVEeRc0PgXZiydfD1dKDsxQb9WDz5bi1ZlvEiiy0K6qAeBNnoU3v6xO6FmHoGCD
rekxvz6rZLbEB5DhEcGI0OzU36YYN/HEH66ZBpiYSDw8vgZ15hq7NfNr9u15TjEtCSpf1U9qyqdK
NTQIttZakxjBeNU1aJgzwDiolpzIWHPM6cuay29f15iOyaY3RY4whQMkueVGqwtCOcIlQQ9EnPH8
uqblMhDMabSZbCQTFXXlykKuoT+gW4mz/ieQ1GBEepxug+MQy92SjAIhl1Tli4iHFpmbWipGWR15
lum9S59CC/N0xdD2iv4wPtmNKAxpiTDw2UftD/4mYKzqRxBLrllCUBHigle6j6aPbcK2cRKUU6H/
7fRrEYW3UlgQ/vJJ095C9tkgQdaTCrpxEyvIiixGV8R5ZDaFOv8TEy4o95bSSirRA51c8cwEckXp
VjtTK5PFSC+d5VX80QXQt2WVE7TVH12FpEckdzOyZhq95DELtymkaPC8i3QKZk/gDDjBWT5pxyKo
o98QstYcYOEwRhq5B9coxpyJJenXU/nTeZm/bz2APsV+kFJARoHxpUQBrraaDvrIifw9DgYu6rMR
jZhykI9oK4OzpQQN9ioFvNpyIk7fcNYU+nETuqujC+B++H24SZdQZ5eLX1bDSp5X8ZWJxAU6f/s6
X7Yf0XmMjV7NrLKvcNPazNDhH10zSdCOB7S0tOm0+xcg9icy2QnwXIE7o+KR4LFLcM+pdP0Y9b37
iuF4Lsy2z1dQiSeEWfxXTf0N3bxJ2F+anjY6aI6D1caLp/vSEntWgOhv0ogef4d+M2puuKF+35SZ
lG4x2WZhqM02fo1evuEu6sqNorx02J6aDDNR2bwIi7/sQEoZ4aY+Kv0L8rfOBx4Al9XgAEcqUV5y
/nRyp5Y2xH83/Ab37n+5//gRMECDGT24UJOl7J6CrAyRZzbpDD/JOuoWw2iChKsIFHWkZpetrRtC
rThYEh+st975fZXGi+Mc78N18nshA5TvDxbdav+V3wTu7+1JX1/3+jXkfmucHNe0tnT0P8aeu8yS
/V92Ig+nZZekOV+nBRtfYC15pVRAPn3nO9L4l9UX2LDpMG4mVKNKEdpb6BEccj8m9M+gI7GMTrMP
Ddf0gTpDxk8maJ0vNZApHSvCXTzrsDEeyuM0x8zgqPP8YBeGKT5n475t6q0dz0DwC1HPWKgbxefS
mFXnq+01YtPPEpsEYBxEyy+k1pq89mxARRaoseJMSCvL0z4Y6c8vq3DtMhWWIGXEy8/Oc3RBaIdl
1HJgVCo6PsKeAwegHnI/3tWAKo2766LX+B0rzOvcCmj4nCe26LzPNAl5Sj9timYDpPPI0rt2ogq0
IhsaLp1FjOv57vXYK6lCZ1vqByjTKHD4GjQHOL+nPic2d28758DYoIc/Q2IDMSMqlE448NU4ZDbJ
+7HNEnlQBj9vKG7GF2YYm8sP8Sl9Blxb/oqoyxviWCtui9BOCWp0onlaRFldv+rUyfQ87V2RfH1z
pIXX9E9JIQodclr+JXtd1PF5THambXfiOdRp6rX45ALBSzefj6wgfvoEjzlxwZlfh2+n9Crsc8ZX
w4nqJH5Z31RLtZOYtcXsw3lHWDV12X8+EUzOb3JNHaPtKZYRrJQ/CAy2CKWxqsS6+wwrYix+lwcd
/TmJovMD4aZ3UGYYvQsIX7WpuC9atqhtP41DB3bDObSEsrf5VTLQuJMJvHL20F1e4koM8Q5p6bA/
pE+XVIeyieGR9kgm0eCNUtjI/oddwABVUTzhw+Xw7rSDOOoAC0Vf5Laq+bfcwL/gy2S+fhptI/5O
duo6DniMQi22PWyw0qRE63I6zjruarYeZvPDOG9Y0CIRRaH5PdTsPXiJi2C8NLljXt37Fj2jEyo1
VM6c2dWeF6APKgeC13R+nZcUkkvuoPeI53VLNJk0Lew76287813MJVCkxLqsMJTsJMVsA9bMqCnE
WJVeoEw+JGIr5KJS9iv0Sw+zkgsWzkFu+NNsmEf5QXU3vQM+lfdsZt1JDLQqfgKSQniMcwcu6hh9
kVK6YIAgPAZK/Z4Cstl8jgzjlrVLaxKGioGhscV7pEQ9EVqPVM5cRAogTW9cNXKoVANigJQlFhXq
Jrx6Hizeefd0Rv0c4IkZzNgplNvAAlZef4H//sjkMsO/NjvAuuxolE57pGAgnVSUbykfPFsr/8Kv
byYdxFzlYpIdfbfK13lONuidOy7LM3znDpvQ/kEHkgcOLB6HlAhRtZ8dccJuqB0vgU4nxF52G+Kc
MhFAw6YFGnlJVGbsUsBPJ0LiuYa+DrLqcFTRcJQHgaAeiJi25Ubx92Bys3/5nAQuHhXtz/50DWxB
HGK8nGs0Xaw0z2MC6go9BLLs75nvS6xnE/9jiO0DtV1pR0dPL0qRNzPzQjbjqx93G2vvZnLRZNQk
HjvnJnc0iRtIZ0XWn6MFj1ah68K6jMHDwdW/6lkJ65/LlwDzSv3PlvYoiadTCKbniePX2XDi9FO/
Km15hMXpjWX6nqOe2DUJXr8mrqkz0hQeAt79ciHrzZAsJ24Zy4H6nT39HJiz0kt50TCKgTycMcCo
ViOtzC/Xof3gjY/OuU+Og3QK1HobU10rkegm+jy3THVa3QnGdrldRCyu1zcE+Ywkm6zX8TDD6Dw1
hFlqwxiZz+ANZfOCbFxxnmT/86fR7hlHEhedbfG4LsfCLKMUrFJ12xzsxfUKyLkF5enTFT2mGbBa
39pIG3g8cDTAIDPAECfXabuRc2JuDBgvcYlQnXJCPAe8T9XZHwci4EpXJTCgToyqH0f6Ex7EdKPl
uQPo62H1S/sCBLdTHlmUJxxcYYMpE1U9b8uPUodongfKWOcRD7xJ8G7lg5ravcgoPR19Mvjin3uM
4FzNWzUIg4TZ3t2UlsaMN/y1CEE9hLO6YsmRxSxgaWqIxoQ6JW6OSSoDFLTFmGnpqrnhMKPWt260
BhR3HM4py4zuMu7kypz9awHxBiFCWMnVIPMEbX7wPCaWtVerISG3fE/jlGuLZIarthnTf2kXfEi0
miOYMRXD++fcNM0Uh6QkTtXBgURgOx9KsQijujknuiw0x+f+myHm7uhuwzTdbK6f1VrqcubjRh4J
yrpEiEkq/bajFkOqAcia1ekQaA873U4Jw8J89gHmnqs6lkghcT1WiSt04rPOkFb1psLq6FHAQHpd
+hjvomXvaQOjP1uPF1U/mA1B/oO3Y82YYpkFmv+4HI7YW/7C4kCEezqVWx6szNLBBBd1OHFpfB8x
DaR1vptHpLg4tovTpVCZyYRhjUExdD/OlfQFlF38eezA42d+ITBJ86RxajkeC9Kh5U+heoDADBwJ
lhhA2R7dsRERffGvt8tAKX0dEnFgfi26Gx7JoZu8+UOS1BNuTyBhKZXv+FkUMRNMN0XnHWJ0hsjt
YBe8ifDM6DDXG9ZEFCqP5MTt0O6dcRNyiRNMsZtuviANSeIy9q/EjYGXA0KVgGN6g/5BhFjs+SzB
UCvjmIKsgvpOeOQVvylX7fEB4KhEuktg9b03vcd3hfw1RKek00iB0OvNeQDAQ8Og0gHtJVO/CWC9
Q8OBFpaJzsEyHN5wiZ0ckvPA6U1xft+U2wACn3jKbsOwKnDF0zj1UzFZJyGPwCEOAeLA6moTVEy8
pCaYTcvDU6gN3jmZissidg9trlm1DFdkuPPu8Uz8athj5n1L+dTZl7Kk/goyfHPLm/0poqdg57q+
KAaMbhFnaHRJTl2JRYsjctzuaq32MWZ92ruid/W96pDzpBKrwmvWYBRM1xRTL0TkSDOLw7olT6k6
EdnNVpV/7xcJWsQw3a69ET8FQNU7wYVJgdetjry7HxsG174k/YqSXA9pDWuzQmmr4wadAPzaHiQr
KZzaMlg3yTEg/pwVwRSAjs+8t3wRuIsHlJD3QM92B1ur61WXueUCPhmPxNILp7TutaVwDll5nUoj
XOJZsA/64ZlsgXNOvrx0sVlX8cSTYNAPEOV0UpZW0Tj98s2c48m3SN+M9PziDD2+fpmyBc1REZ5B
bL9VixTkrOdY8EQlxhoGnzQBRRA58BY9xwRYISR858E6iQ65ohFdRK1/T8+KeQZXRNgklf5baiLi
6lKUUEFDSNy8JksT/TCRDe2ezjW6kuXEtltQLJWPjG95sfySjLxdKoeptQ1J1wJgwz5U56UkOA3j
h3T+r/TA0zPctALrybL3YC0osUF6JCPKAjRBlIEGB1WS858xE+ucqfad85cbM/dBiqtfH1sDWpp9
59tXikyeM72rWnNVnJgxFjw249QLvtxNGwxqiqN3hQ2AIOIVPS8J2Pk/vqrk7Q1SVs5reCyBQAFj
pZxQxdleHSZIcgF5lBXjPxt9b5cnKC+k6ZJTcwEwOL2sES9ePYFHpx5yEmwLbjqpOMIlDAvAH96D
iFunpS6GeDoV/+TlIpgSazolbeDihvvUCQpE6mI1Z6XonGA5JZGs28RaLzq+0pY16Qnu9x/UljkD
2bLC/uYXo7aDyT9SoXkujZT1IbKWkKEh+H6QZYLOXrlKIznImt81RYW8cWho1SiWRxKow2kdYrqS
ZUWQEGtuP77IkEwBLBxxYDaLlnIQ9w8JWvyOQYQNYKGvrpNIf8zf34g/EuQxEUo3j9sYXHT8fZgi
nr4BuqTstw3N5AIXphxR1pBq2yGsbNMSvDOmHdDEGrAw5kFx676F+MT7NFBUIF+YBLCaqZMEc/71
zc+FsgcuC6JHK7cQ4FGw2u++T5oers9Uq11EU0uRdF7ijCmdaCyyWvW38fAqVJ/p23fmfhPsDFjW
87faeuDZQrmOmsNW3ZIs2dtBD2Pb6ZurdjbFFzDho8SQMJXFCUxK11lkyzS4SjsMIdcSbq7lS3dC
2hiZ9n8MduvX7WgWn9MvRuOB+U02MVpJASFDYcHpDcbfGuUmH3e+LU8jbwCixiuDPJVbM6/vzzp0
cCgaiCJz7ZHUy8GKxxI5raWaNcCzcU/C3GLHGL3hpW2jYfx6pxkUw3M/QTjg9YmdJKpZ/5MBTAL6
DKgh2CRh6AJMKP7NN8AuDnyBf0MEyADneNOSeBH6oElKF0aHkwd4RzkGHhP/bJU+e7rgdNqiz02M
t0tpBdwAqqHsHf54iuQpBXGcizsXwgC2yHGUzGOyqN755GJGOVv8W8ouj3Mq1ddcvpIDNCEoS8lE
PlblxSiAiyqLllBJinrz4EQG9KW6OWzN+2EJchIJamWGMjOPSHQF5FO2mltDA7y/2PFYu/lXLlEK
VUeYZC64O2D1Sgimh8sjdtjd0mEJ+NDhy7xlLDB+PFiRqIzW366k4ghb80gWJBw5HVEMzofAnNbt
OlnezZ3QlWGfV0dch1XP6Jsd7Mjr5Cpe0Fqi1tIrUb63PLpZa1kVVWrTTTsm4Geh2qAX3Ex9zkKr
IEDKezzfvR9DMCCAefWRGCO4LhmWPYE0oT/6h+t2IyTAD5ox5AXFnoh3+RKnlbn6hT5gw6xUpFZT
ZWC7m66r7f6eSofx/KknZ/PwnzVtS86Nz7EnHL29pzoGEK6spVVhmLmm3dzog7jXKpYieLcWky9d
l1zW0mCEu328Po9d9WINwG8hnZYavDIz7ro9varUK14SCk9V10WKTco9OlavOXaUbMRP2RrIv+Gu
2Y4jZGUvWcJS7Ho4EgNBCtRBZHBGb52jtjdVPGWdfspZDrzcBCTFLSdnQ/ioYVeQvjPAXu09MHAT
9tfO7ns17w31RgXNMexFGZitXTk53QcGmk6auchmUC/2SOdFiV5DUmNYyzrf/O8rhi4uMi2dJ2uM
PYsaa+huA+0BzQsihhzFQ49/t9/lMuqU0eluFSwFpYriLHLQ3rllcpAYv9GdX/0uTRwvQ13z/SNh
27ZxdOLsOPHFpfI6yi4Zkga1Bf2+CgGNIS9T1NSCsq8b/OAARPhg+N1jdO56DX632XmEi5xZjpP6
JVDdKIbfc93tM/lOuHOxup/z/EW9aBNx8EPUYiuhEEQpKAw3OzXaYMKpMdpIN15UakxNdrypklpw
O2fq3uSj7tSAvXLFCCSFOwSfHzdmg0d3ECKsylJso1WKZwu+iob3DiO5MmKgJoIKultwqoW4WjZR
Hr7YhKJEYVZD64/K7qzv7lLigQhu2zvCNk0oRwIcdsEz209yGvRxNqEw3DI7jY6jn9wk3G9f0Ad+
68JBfVwfB/ZErBFV2sdSCH+RH80XM0gdOY9YUSkTPB0P/oKMXp7OMrKJEq7RSbVJ4vdjB60b+qwl
UtM+EGJp6j9Vr55Ir/v+mVzXO/C6QvfiAcOUhIuvP/5TmlJZARe0COA+blEoAEco9nex0Tag7Rdz
Ohysdsf9PaxwATB52uYHI9Q2SPSDmBLm+msdP5wHywx5TEy6d8gXIStRLZMpyosO8bivj+Cfdz0R
ZGtZmt8PU4enevBcYdElTWAFKa8sGJ2BtKcJFFgMUo2f9qv/k+aL6TDEkKGcnytU0Fv78TT2f0B7
dH148hFgZmakqENBA2J+ShzxMhiUS5o1M34HjACW6pxJmpuDaBemvsXrJ0aGQETwlFhm9nVhi5NU
7brALntJAwY4THfFyFsvpy8YlV81/yy4iVIXPWZ+bOCerLStJ9MyJCgZF5Tp/hdpa1sa712/zCZO
dZEUhsw5Q/cjLj2HDjTyiqW57CR6YgBa9MWutD9YCp3Xem3P4W+ltLqaT4i3hOQ8xhWx8Dwv6OxN
HucbQLQvJsQFT5qxvR2Rzgkjt5ExkcbYVUYou5JU83c59GV0ojP777KkHEdz8Fseeq/ikzDc9EzG
oghGs/qGrMPYQqgEsk9RRcITv6EMVEXJnLiv0LnCnTHMbRhi0UUtlbAEz4zoGT09rR/qjAf+AwNv
y1iRsB1FVMJaqWaPt0EHXGj0Tak+yVaf1FjA0Fiw+8oO8XHUB4NH5bMbzp6ht/V7+MJVDAjKsxZM
A8e/2BmZy6J1Ra8BaKKKxgKr9bxz5Nh6RhF/z9RUXHxMNSfuF+cPYQqrHQiM4W3a9vt8qEYtTkM+
5beCBNmtai7u0tKc7/Fr0rRv1fOfgRGVrQmQ02O+eT89W7DRVWdYkT5iXapUZLdhr2x+F9TO1BPw
qfCyFKQP8EZTKRSnbX0AM6TOvue9Z1MNHHkV0NTeLIRiARVsudkk9ERXQTOJJqmV8oF7+DrNIJjZ
cGUppkEbRKjwZl2PwB4o1BI3kdUuUFDOtEuRxZOUM9LsrZpGXwTiPlaPdWF1fzfMRGe5q/hHuvHs
b5KSxhGJUBBYwYc9A3pBkrnpJBwu1C81q6Fo9v+sA7yKGKFwOLpzFl1Eo2xTw1J8DhPp5coYtz9a
aA/00sKIoxDp7zve/KOhSbyg5JdFm+eD/oA6hrK6EUTOtvtuq8v7Dd3E6AbIADzIVlX4Fsb2EiZN
1BKVEL3mhZkd4b8WsPWC0sKl27JNDP0pfD/EtMyJrbGGCZEDUutLHlf2trHvzaL0MGKRcFZDAhBB
jlmIlWEfzdZxVkCGZHjr6wI99zSpyzqRL3dfHp8HOL8Q7mzkz/j7XFNfDZ5GN3t/7/dGNml4qcov
qzIvRIVb20Wq4Hc5Vrq76oWJ3vLVcHM1xSVx/JfGPrD5nuVodsshEIA5QVgBbXx03dqbB/n1cNkx
/VrYYT3kl/dwF8vSET7eqJv35LifpLEFxtlAggHgYAe3EvsBk4b+yAtPfOssOwrvkyX10xX8S4/D
yYP0CVHSc9jpikVt2f0FnfpaJ07JjEOnXS45qgkFOym3QxqGaDgIlx6qzt/16NqxRMyxPDfA875u
tL9eUYY3kjdaGSlT+I5JmUs7OMrHmTAIh79LfsfuHjawL9gTO7rfrfYdr1Om53dZwqJblh4t765i
lMdvQJ1tNlB/Mkt1Kd7f50wW/bfFjvYkKqDA3NIJGhz6gAuvwnVPdJzgxICnTyYH2byl35cZYnso
fOuPiUXReQ1U88FwgcZQpG5aCU7u8KnnGPIcUAlg3kuyYXVI3T/dMbrIgNRl4ANr4gDnInivJD4g
nRB/nYLdsGoecV2z9ZBCw5nis0kPMEGXZFnHvQnZihvaGk9DPI+O5alRDt7peIj/yvS22ptkLlS0
UfDeoK8YYkAdppi8aIgLCqxXUoYoT6opEcgZolNpZsdZ/TqDZv+uG+DMKuWzU5uMoytZxWXrJAdp
7QX6zh630GSTK9CSkx+p+hq/IAGb9hyjiKKO7FtTrhFhUqhXJPEd8DicqFAGY8nV+HO6vScWJXXb
M3qdybTmsz5VTH1dNKWbmtgppkwQ/9AU7PIt8frKck05wseQHbRqSjqVxhBg4jp3VGO6JkK2ZXyL
2791yFQE1iSLXar91CSWlfyDVb0NZBYKSKr+Jk93CTJTTjqcKYGXS/7tnyPF/ewWwH1OT2mO41Ht
HKsC2oIsjI9ocoqaEoj+gxN2yIlLRYtIZnX4JJyIL4+j5FgV5hX+xwPcedspxCaP8jV/4mmkCz6x
sp5XXPcfsBl2zHxG8EcyyR/cq463gDJNq8Lqk6nHJuVBMXhzW5rFfgTj+9BmjShK1NR0KRQ+/6Gk
daD5P2ndFoRZ4WFDHF3DS4oT3oVGtas8n8fAEChQOjsim/pPC1A9aw8EcWQHF0AuYxOE7Y+PUOkQ
1kGbGrOR4IPRvjq0aBxABIGmbCY02E6MhInz6/9aUdhaFp52y9mBqOAsbEgZRsEejM+efGL80Pgr
BRV19crE8fcB6997Epg+NagNg98zcZk/7WfTAvZ4fGJq+ni4sqaUorA+7UxR0tUj872COayh51dT
JGZmzrd2DRz/Yjnd2Ocx0j7eydUGfCVqkMWMgkWX1C33MaNVI4cuFxKULyfCL7FwHKKsaxxM/HRi
5rxwq8TlNsMLOA1VFqlKhZc0sJyoDp2D/4H7k/sATKJEZns40XsUaat20JZ+WnrY4HlyiCg7mk5g
SUmGw/yVd2aH3FPbY88cuXs0Hwe2vSMFWEpAis8KnALa6mVwJVLo0rMB8fxh4AwpUlLpJz9EZ0x7
FZEvLHV6ouH6gBiOBEwQCIFFMbMHEQZp3DZN+qy1zAfMPSqvtEdU4wjN13O9Pbcsa707t0h4/vea
/5u72/yMtORHDRdBFiuNd9biRP+aDtX0JdhtG4LsiTQwMwaydbzjZ3qPzeaB3R9GX6yZHhL7xxyk
ZlWeTmpiZmd6En3qW5op1VRfEAHyakRIImGJGZ0isFP5E8nx3YE2cFqXv7Qo7eH//6bY0EYNyh+Y
8LgcGzqM3YA9jsUMfbvYYW+MoV5awiRECDWziUgxPyjfUOgq9PsmiXXarKBdssvCXR/hmBcW5r50
Xa8tklmd/KmT5jBNmn/8WEUU1uf5xSBgDPG9XN1mA0PGmXOBbbjMlEy3cHf30U4aKjEH+9HNpWvI
kxfcvvUhF5glnwtGfleFF8hGXbbbAeNT3qXmmNhRGV3URYNUBk0g7M5MjZOZ8UWf1cs0WKS8S2Gb
cvrSMv3urAWg0TnDPjC7ea5govA+jr3JESDtMI9zB+uJ7cu8pk6I6s40g+AVntqRqG7O3r7EQFgy
cDT4PiUQpCnLkUkb802nlsPMTn1TneAYBAxwoFoZjeY9Dk6qSjfu94LgQ9qy7WKzYxPPQ2LPKE1U
dUFFvy2Z4JL3U4MJiPNTZFwEqG3rfGWFXGyEIHBjq0E8Bih0cqNjCtIN21waXtmGpTwh/+nT50XE
Xc0UT/BeGQ1rOz4m/sy6DD5XVGbcukiwiIUrQxE6tKbl9Sh5888L5msFCKS9nH8lWHwzXql5kBkB
lKG8TXATgaApucRhqU/vtO/sQMtgYUcFZ7AU5v4c9M9BaaojJ9acKIP738IvG8sHMYMgvlWqNDOT
o+1U60kuIdjP9hvw2UyslRaPOgDoE6LYgWt4Ap73RfMcjOfC81piT9DYsruMmDDCMj/ouanXaADN
Q111V8Jt1hi2q+/KrbkRo2irYUmBuJMRMvUQ6pwxEFeokEBhs2glhbbBk8rMu/yOg3pwJZ7M+Xwd
0yczioI9CKBEWtZRgueok4/Q0Kn1qsZXx/Yw44m5Oe+BHna0vnkYKOx+PNvER77gyVcPsqG8G52B
cZO96ad/c6JeVlZJeez+voNXXBqDHiwkJjW8Enfx5Drwq/yeDp/FPQHnSAsHEUihP2BGfxFUoXQo
PtqHvYME8FcrJhL/IUXxEh6KaZHeqF+2yf8LCIUeiotgpSIYLLWYzXh+WeIttdm6SxNr9wJIWTPn
Pgqn/OXw46dpzAodC7/jXg6WMrKxPJKbliehbpgO2N5+Q6oWKOEGRDtZzndIYfJzolYN0/NNsJ/x
3bCTJien44AD8fwfdUxNv0RnM86m3p99eTy15LZoPccn9f9bw3z/06974nRp1/MAmIHoaiJW1s3v
Dw/BBfXOzqKJVLVy9OaWo2XuAn3zTISUEKv2jo+uuWyOyTv7FtaPLpdEMXb/3VmS7FaYVk+Dv/11
iyozxPpX54+2qHEB6u7zfYN1j1dRyZkDCZvgxY9dO0CSTFWP81RP00BvvIsdUD7DH8qWuBjg0RaX
gh/PE0Y1/JwSiC11HVLgSEcgY2P106cizJREmONwQbYNOkACoraeASbwW6q5Oo7PmN6/gn/Z//qC
4ti7Rj9k7s+DcXHn2L+BMQ9SSduxVTyISB3PFHvsKbfofj0sSbfdUDf2/X46dc/ArkQf1w3ZsTz9
ixYwy6HIxpC5W1j5qtfi7KYUOEw+bDSjW87X9G/Wsw15IJ0DRLk5DHHhHam78C+HLS4Yyv8+WvI+
3eIwP8pEAoYX7RyPreuLyw9U04+cFP2r76eidLoC4LudMVevdlQgMlNrWa2t3wM/l0m55Sm0hw7c
/19DagvJX8uophTfEyAgMSPhd7F0KX/cZa7IguCUoeJYMMw+t6MeliiwjqOaHWK4jtyPWFQDl4IX
DJytLLxePnZaMhVyhODLduIge8TxCGRmAi6gKlmtzNQsdK+H1nRpo1otgojl1jkpPK985wtKI95t
4duZbYDGOnmy2qxT/S4S+FEa4q7XcZAdn+iaO6jvSuqVHtEuXsXUlG5gVF0+DQBvIlTiIT7lg0hz
az5aWl4q+kny9k5PV/ETSoXiK2pNriCt4CeXk6JMHH7nQg53pQO03YBSYVHz/8Rgot3GDdVXY7pJ
g61VyAFE/MJY+vsXx941MyiJbdYv+esOo1aVEk8lbKJAuhafrBX4GvGhvIHnsi/QplIpXk/IJsjD
CufLcdPl7t5JhdJd+tnV2OtiE0dAcD9S+cL+2UJ0jUhmav61KAp11YytgrpzeMoMFLZGVIohJiB+
ul1JIflhL0m00n/2WA8XnzTVx/3+Sbw7klBtpHa3Jg9vxcfoG54VLYB8iT47wspNqqkCZ/iGFMA6
JiDjRYxYdfHEX0/2vHQ8G4l8/B5H+bKiXyS8lLYLXdNJ1B9jHrgjLxhotGSCxGlsewX1g5ryuvfR
artrze/RVh76hOA5I5klEmzoloj/xrPw352LYnFm8r6jWuySKCKa2neIfape77wnBhu1hE+6qOVE
WpRIobIj4EkVW4cjIrNjrUgBQgQ5Z3FgHkJkGb0ernqbOTSSsOT61mTfqxV6pZzxd2T2lcpQrI8v
r0SFp1mRndVaRkvbtikkCnGMOHQ2RJPPN2mTUJwzmYzgkNvASRrQ5eoinMmoAOWMI1Iqin3TlRle
PTMFUhrDAeMX4quHEGMrioe8dgNedrV921ZzJyPGSknLWvlPBCrcNwOi5oBJL1z1qv0uZkukSYNF
Bk/EZm73VozC5+LZeo/wNLncATEfe/vNuYBWSkKYa12KhFYn27TsmdYNb/0cR0OqIvBeo4+Vz6xk
ddofJgvO87zqq9gcp+6U4HCDvvx5Re/cTffsCF0cREmhDVN6e6uEYgti7xMtd2uQMLqsIPlzJmlV
8Su26dsFce9FraZ3Ua+1rXTYK7NcyxVSWd83OKE+Qz7jiqySnn7cq9yF41fhc90HzCP0EzQX8jC9
XZ3+50sXAEC1/+pS5M2Jy58y9I/q1dQQ5HnhvGDhykuHTYuVa4fjh0B4uDoSrrvF08NL/qdeMFLc
jews9eIZ8Tr9jnu8ZXlBGWuRVFa79avNnpNicFfVPVsBGu/Cln6KPuO0D9IxVF4OcpNlWuKp0JAV
zZzThyx0GE07LREWUsE0X/JEjPIKNmC/Bmu7j7mA0JkQdq4A1ymlyznPAq1uYHvBFTGdK3Ew9yAS
wkpR7aWvA6qf8TDXhD9OdS5JEtsmX9DERy2F/Z1KuHbFQaZKnddoMBxaCZvZSZ5StANpX0jJo8/W
tYZOqgXn3dg+MVoZAeIQ1qH3bNxshVnAQBWLy5RQC3gyTUwPIQEimjSqHqO+sWx3PTqAJ4bhpNUf
yeRwnE/myX/oTWnlglx6aIfbU+fezTUtToXKiqvo+/4lhWdGm83igjYO2PeFTO+DUkjppZvjpDK+
8s+TUR1Pc+CbNbgLuRH70EjE4at1Lu/joPDrt2XLZ99TgVuUz8Ru/NDfeUf+SrZxnL811JdW9ZM5
MRtbtsNeWMoFtEBTJi5cfBkQ9TMyrKI5kRv+fw3zUSDWFgGJxl16baoSvN3HbT/HOWsbvhqj2slU
l5nNW+Xxnk6myUERH4zcy1RylOz8WpexwvPTSbCvvnPXoKpMSo6SNi79/v6bu9xp3dvV3ZSb2DGW
vOHjlMtu/1wPbjC13zryLxSPz21o9TRU65cKHf2J7S9ELlzizoHwt5gpsVKciNS/EEt6cxHJPtLh
sJOFF5f35KMDSFislK2CWBZZMmTNZtYkWekA1VrYavCgcoVk23ywIw6Gsw9Ur4GxOPEaIjp6JhLt
vj6aVUiEju+B5Y5gZUc27lr4qJaVRMVcpeVs7iro/95YGGo2D3wig+N27ZwR8CEw1N90/Hi9lPUn
W5Q8mLck5D49+DQTeC0EHAJxByWoKP5BWhO3cKpcuLUHJwFJ6Mm4vyx5MJH52vHqBHKMh01tcl9R
AbBKYZcZ5Wh9wpV22nl6yFZO7lv00buzKAyx4x4HPJP+NvHINd7zMM8kRxsrr7VMKNOPAjfXqez5
tYDnYo9lKRpEpNG26oGmqwMCAq9rJOvgVpfDpkJqstHRrYHRt5DMS4P1gUUdURpWOkih5MGkzMR7
ejfe2MkR+lJ2Os8jXvSnhFcOFQ+coTZVprN8kWOu6u9PUzrBcnpyWzbv+f7q0QuWcUUTREsqbRNZ
IyW08aIkFghldvAvY4RvMIYv+qQp80Mjzyfn2y+fvXvRdKmijgpha19ZbitfO0o/FHx38dO8enI7
fcTnmWLLR3Fp4ffrKLjWORQc9Vm1QLoINFie6vQiJMu2NQ5gpaKy/KPP0ftariZLurj/KVgftM1C
sPaW+iVCBpqJgVF0Xs7EIYEnATY2C5hVH4Dhm/AQlC4TJXIcjkB9jGWbgzMf/cthZrHqT03S7Na3
XusCbOdxmHGkzsFOB21ZMWD1Ra9877/UCmlHhfoeG1GW9iG7+upFyW0cbxWhqcyJn+oDGQzPU2AC
2YG1lHaRpRcerITiu9glmZ2B9koi3hjU6MUusO74Kl2YpLHmpreNZ6NVV1oGzxN1u0JonaBuj0pW
4pd6QU0Qo4uQhVOk89Ibc2VwefGkVQQ57kj5GRnx+7JbhDZNVZzuvnMgziQDrNpkWhU+e1/xGNPX
DParVf5cgO4JCTMF6N06zeLTL397jlGySd7ZCirpSo4elTdNsOefOvLZVj4VmKj1uuUmHeBQ77Ni
XiAYMFhpGPogff0NZg2F6hsLyPCQ0wuHszlYHpdCGUXCi/ps5s0stXyy9nEA2tC7jsxhovYlNF7A
krNGcIGCIff5Sut8v7Mq0pVBWh2suXzOtzXpJ/mgT8vuwHulZ9dkh744M3sfF25/t8L6sVsw1a+0
Enm7PVc8cQt49glAUw6njXzSMXkynUFqThA+Gftw64iWddLVc5zoJPYOGmguFaACZhzs/sZAlxtt
7qGx+PvaWBSo8aDC6ursiZBgDjM2xXhBqXkFSCrATHF91kNbvR2keGffPDKgHF7qr9kbWFXQLJGZ
lP1Cg6hGQA79IF4r1TcbSEXEBsg6bOpYbA8d/bfETaqReaocOzIQb4pf+VFC7EbDZO+TCNoGLGE0
RFmOqI6yA63uusOey88DAwabmMJ+L4TPIRhr9joiRcVTQGucg1iiOh4r9WKcpvFPRILlpY21caHt
5fJx+8PMgoppxuau28UIdqKpu/C07VgvxcT+i9QkNoO309ADaWezQNGYwtGZNUn3dR4T2TqN5/9i
fBXdW6yYxYswVNWcB9FLSgAWfPjYW8DtXwCXwmpjKxfFZVkWvcie1O+q8dhARHfdeHLbSa7fRpil
EZ3Z+ME26y/gGNfjBNsDW9zUZ8HhPc2g0+RqJGgRKLHLKLSUV5auyat6euU0XZz7CS5LiXsXF5+L
05xfuNWzjITXdDcX9uxrt31C9u6r8RssvXHOwib8kB40iHxt7y15cwhsDuBk08qX0HRfAYu+0S5o
BudbjbVdvBu5MskYhVBszXQcT4LW1cxLia45yJCmhgwgu+i3JnYIFCkKnflc9SHcEUUrX9hQVwy+
O1DTgyAiFzj2Bfp6NL7c8O8IRmqJP+n35k8I4wknA3/GTrDR2KyYckEf60u9UID64IFR7crN3YT8
1iOiR4HzRXEAqp2CPPhe3ILeAxVam1nJvMTdKHaKfwlUhME5pt39fOTdSYzq/TrWCgN3qXcqlyhk
QISAGlNepC+celEUZpRfSEDEWd2mR9Ex6b14X1pqWxbC4HU6/hwfJhtn8tC/eVdscymYdM6KEfrk
TY7wYvyOjJqzmyGG+ex8g8Hlaki2SaIaJS+QHBUeNd0xRpAg4wkVj94l5OadqF5cIFTWFMULFd/Y
V6ZIiDEjWncK176+Cp/2MM1ZxIklRmwYTIYG0bCuRBXWCwKPFrFHc+JU2DaWDAvGapwFB65gM8J2
ZbDU1AJIgWDYUiN3i22pEKVz6B2jlsJGSNnljAeIVDv0lfui3yDrpXf0pyvA8Xg41TlKCjmvstZQ
MMtJh15vp28MQT3eb62gXJr1rGr56QkgH2QYv2KRQg3/z7aHxBwh7qEwjWuBbWFZV2tNcCtxxp1x
yawKi9iNdHZ2mR2lChb6Eb/dMf0fMUKrAOzr5YRUoPCIDyD7O3I+sS1Okf0IskPGnajxt/gvFMdN
QcD+NmDfz2RzcJr9NI9Kb9eFIO+z4/Ic3/uEt7VN+ZRQXxPdB/fxhN0RUu6hDILZBR1PYptMEhyq
YqGH0Pq9mmcVL67Z5i5W3/7jfuF3W5NN7PFPMVyKFXUbAp4S4Bd8BHh8JSjyPALfFYTw2+Tqf9OP
I/onIiNnVtEliktZdVmvYytrSieX8+GnEqUSCkw4rrE0z+oej+7cgu1mwzypqgm6jl/MHdjFSNoC
myZk1w68oX/Z92lhSGqKFJP5LZ9UTLFX7s2DjZkJ3l2FJSWDJibwcy1FnTKmRUmfX57zre0wUunj
jkdN94Mh7Z9QA+bENMZOAYm7PiEHrbVhavyDy//lTQsjvjqBqXQyyX3XqFey5UZ2GR/eGP01W85t
LbkMpcr3rVyn5kmkvX2RWOdj9qnR4AHzUtF3sVfZ8M+pTx/377S2PkAwWv+8XepJ5BdKBi6kkvuK
KOuwQ8kOxLRYer9YC/TM6QyaVRjGQ9mBJvOrC0lRnOkUE5w7JAJZQ7ldHLDBCIZadgF/ztS+eehV
pH7A0nWMVYMXG25kXuzOZZrX6ltKCa+Mj7jnkqItKMToaP6JMOkruitg/rzLiFMhwFmapQX5Jxdu
ANl81nvYTajNZKqgsmNM03lfr27onR0DCKS3zSFvU4BmNbUEfAnL/fFPbZcFWwtaxVR5adaKS7Qg
iMJ0BfOsGcS9hYLaFuMZbzSlevBfpT91n1qzORvsGlmYYZPoRu90+Ts8Ucetcwqok9tZk/JZ4La5
n3m8eC/53DDrHPEPqfvWHWEifDwXDjnOf4z0s1TqTI1Fveh1walXZ991yvXiMAQuQye6ZZMJLkXm
eCyphLLoBDcKgyEd537kaqY4nbrgojUCSujgjhW9Pcej+dFGkJoGx9OEvmppvoFdxcMVA+o0J9+v
ULSaWioJTbzge3mEWWM56W7oJgyaOHHUg8I4ti22gHznl+h5lRZsxHWdPy38a5ILyEIYB1I0boNl
s8HO/4s78dbxUtj1ZszdPsTxv3R2PTTbKwKhS2NffZgu0YHRM0FLeM/oHNn7YqAxP2UOg6KrcL8U
umpL2VaVoIGjZeGU31HsCMlmni8ocx5gNExZnlqPpKhG8jINrQ8qEw9aKk0y5HH8JHLCb7DEyCCx
jwFB1Ybiv6d6ntsWEJ4vRBNmRZ5QJfbyfektHprrpb5OHl52Dw3EOfPBxf/2vCn3IhDQJZXsAP+U
izKVzh3LrA1oFY2xh0rFYM1/hgM9V0cSimVBOeE0UNDEr/pZJsRRKYQdkAj7x8lbUA+JIdmtbTde
ZeajId1pnjdLgYmy3Ke1aDMCggSzNiJ8mEMI+saXfb2Gm0H41EiOT5hsXUIwLzjvVYHaDYlgWUb6
d1AC7G8FOPtb0IyQ3jkQ5P6xPBa0/0bpfj6flPeeOHuDKOU0jQjiuqUlzIOJGcBI++cPztCpBiZv
dVcNNoAgLfZHZHsxxva/4xkuAy5PwW5XjjtGy9WGCQ0i/GgfbIkSm1x10gr82iOmkQTnhhOlqCqM
UzWV8J2HodBCGjX+40Q4fB2FJ7z6JE8zmQHgeMQTgfOAWv8z9rjtyMp71XTzQ71iqy3uTxCShOvj
NNK9Xe/+jxuipI4JIs5z9pW2t7lVkE3hcfYDL1BYpb/iVMEYIiEq5HHzr5j74aFKDj6FbxZL6tGq
J3M6yyIrY/jTmCXRV1htwwSufmlUMbrG2cM4oCfy3d7xUmx5guYEWMkqkG5ovWOs7+ZUeO4+bgi8
EV82wLGG7aU53i1J4g+MyV1Dhq4gfeLgxZLtNEkMI5n7XKJl6S/oej8ZIUaaubR7aYv1aixodT7w
h7ytzVTgM5+AfHcBwNu3X1bSysfYrtidqTcI1jhVz0f4ioC74Ug6bylPfh1oINILKpk52eOVYfWY
lE9n8pNbPSvesGsQ2UnAjpZ0vSX7TMv5u4o3ONqukaFoEHVDd8M+jEfT5UgvYYgfnJpmy/cetWFI
iSOoyzpL8T/Rn4QYKsMdXzjNEzQsmy2fk4BltgEy0aMFXFWc1BPZCCZwWZF+Y7jvQn34qK7ave+W
Efa8v0Py+/C+t5n3OqFnL2kB8CkKc8QXLpO76PSShV632xr3fIElWzPov8Rv776BSfoetbOIVJy2
fCJI+0wfPPazU0B80/hWHGMmzycHf8ngSn8asP/OMpVZTuJRBk6pK6RU+j6oR9lQtOu94gUyOz+6
/4/sOLUDq/TCSkpPMlg3h2Id9Fj+aMwFYmfa/ACBUO3yLGIZx5X+U7cDM0uLPEcVIykvKko5Y7xA
wU3tppK4oUjVgcCLXbQnVaV8P/XKMvQhY0533IPzpCYNGN87sT1Mhi2zOsSmfhUtrQwjYXCI5DIu
w8XOMMYkMN5KbSq0QjjrwsKz1ggvxgsI5LZ0bGIAQkcD0ms/oK+sOmrf0lnxrCbiVzUPUt+/nGSq
S2c47yeTT0Fw/2Qwxl0V3Bp50jpYNyhdYF4ww8vDWQDXQ+6xpT8gsKCfg3skd3B4eSzFQW39nIZc
ThM60YijbbowwFo/+CTVmsb4YfLb1GucW2eYgfYF/389cK8XwV8Y3wOr7wQL4So2kFzwuebveq/1
+OaJMFUPat+zdPmw5sqe8Ku5kqyXizAVHLmSTrEP+GwYeSK/7K0TSTY3G8YMLcGg5gvrG0fn2KcG
xfAzl1VJtU9VsDY8QeY+1WNG1tvKDq6OLQJNEqH5z5GfnBu5XWjQabH7HrYCYZznjT0gzU+ZDKJ9
0HzTMU6L/Xy7NF0f2JU8bx3cWtSFL2vg1ctDXx7Nqnba49YObyoUWSarAwfZC+3FKs68mDYTi3aL
DIBTWh3F3EPTxRycCLXEX648hWuufobwJ0PqOR6Mwyirlyqkuikr2wcxIZ0ky3C2cRTvWgYiiHzR
hIzLJMesv8ZgX5T2DdwSAr7mQfY1mSjmo5GnkdktBk6O8IOVqGNB34CaQs3ZNv25XDEzukgUV75K
776T+U3ptpm++TThphMadDp6jRrgUZQnQ0llA5t8TzAxxckafRcZzbWkg293hR4KFh7HWFiHx/m8
IYbINep4GGU5JB8zjY6HpUNkNbWzkBgK/BSRG9wr/Nx4458sBMGhvGWbCsQODtABrh5lgyC3pwWq
xYe7Fs2oAxzM+Ruch04L/6ybtzJyUgsI4mWka/yymDcL5Id85wkNJpGXo32D9a2q9x4Tv0CqA1II
QJdgiqsI1RMpZP7CRrCvpMH1ED6c8orDm0l+agWQi36SpUMx32ksnHr1i445BjMS8vlJ4MsXWO5k
u0yN+0NaM07BFLzXEv2r+0QobwJEezCQyWwgttR7kCJrFxBucV2swjkfTmzDZrJpZJwtSWSVIOJL
5lfeOEY21SkqyZua/iw/KB54/4p5l7EKnY2Cc58f+mt5nLyM+It8qaDhJn5ICMc98Brvm/aOjvt8
c1Bhx+Y2b/ABcdvzmgzb2LBoLSKXwA9O6hL4l+H6fJO2td+4hnKZq9lJxgBwPZHcjsoFJYva8vi9
+kURZbp5GAf/NrpF8kpcb8PVEGCsYnoqiw6ywdx2NprBjjgJB0zfl+/HndMkbAncXkFN+mFaWNPd
jevgkF1e+BWsyb2nWfyRsNivVvU54b4PnUMkB4VXyy/TJw5bmYOR9/k51tip3ixWRNwDV40PxKeB
9glQpkdyGq6LcTIp7aGJxMXg5154U83B9fwvmi1J4yjxmTrFej6BOYLaAvIsIU3wQWp4OQyb7EAX
1JYaxzvEh47w3MPS6JqK6I7NxFbjb9IVkYrYkwr/9NBBv7Sl7pZplAAuORY3rJEMf4WWJWjz/pb2
Q9oYI95RKHNdMen1xVRbsx85mkxavUdQKfSSoNIZ7Gte2Op9jrjVJx60rqjt9AhNR9AjSJTOzIrC
snXaGjAn5ZE+of3C7hQE70xqUZeLhOW5qrQedsJsOOHcOEqRYIUsoigaeSgdx8tB75Nx59YPiHW6
3QHMaeSvXmKgImRnjDVUizqEWWzBCiTR+MGaCav/cvVbugP7H2Vwv5bnLiLlGYd2IiYIMbGAl+z7
4i1RMQFyZUHYdOv8uouOa4f07y8jZyzqtv1IyZCsGZB3fA6T1Y9rdXRThUgCE44SYxyGJoYxB9at
6ymsG9pbIfxDUmA56xzgIQF5v6gsDHSkV+dkObcO3a25nd0vqPOC+DcsLi+Om0DEFpbR7IoWHdqJ
fS1QaHXrm1RM0mzg7w3TRrApCuRTyjQxek0X0vVa4upBDN0k233D0M3aLk1cTZweFDrv1z7ebXsJ
5p9kuMavA1mPMpwEfjMtzBK3VIKBKmgnZAnG3JynyZnu16jXDqz8nOXIx0cN7O3WmvDi06YH0b6j
ul04ZiwCNZx9jSceFhPM65RA3qwDIRq9kL9ijOWsb6bqYgpkjbq5VHNBbdo/GWG8Dw/Y2L7iK7Uq
DugzE7IHd86kGNCpOueu8FZKVoHm6g9Dq97/lYIgTggFn7byyqNAC48JXr1F/StlwBauMFV1p1Dy
Wh+DifWmWBkJ6QBcwrsp6TwXrDNjS5G9XW5eZzMFsH+5RmBi7kUqqpN5d6M2MSYBkvos8yYRJ9+a
h2kQHJkROvDM6KCRNGF7+OQoq1NL+SayR2JVYAx+ApC18K4HxCJPTZef4xtVUp+QYnXFLcsRNsJX
HrXohdHBVOPAnQjZcNlBiAQlrEnBasGdSmr6HCwAPau6AXOVo3U9Nmy5MkQ18l7fZHG13glraeFE
8NO61txnzLm+vQ/6hhmmCS0Ak+KgaE0pSV13mQV9jzYzEyz602O0IHJq4Z35IQ+0BZRVIcwuXCNp
eLGIuBPbpEDuMQTMN56SIbL+2foJBPY4gH86oKIKeCdx6tuqY7rm1CrfIvc9DoAMipfkjRAhcJzs
DsP11ypqRqgoJ5dda1x86G0/X7q9c4ousT/tcFUiAYisNGFTjzFfn6fCt8QLp1iHdWWWU1aVZ8cd
wp4/PlvmgEyrSI6fRcoX2jS007kWTa3flWmOA6ZPLIR+7IPnfhRwemaGsuGnx/NV07PVCe+7cd87
KfBk9v3YmHD2dTGu45P5uv5/6l9SMIfMjrUT/m7dAQi0bmsTQd7Vhq/3mNc6med/ScUn6SzFr1o5
ZADg/rzSclZ83IMKFDCkwDDdY6rpKNVbNtFeocCiTB9wZuFmkt+Q1dl07lmmQXjygkEnt4D8m/o9
QrEb7v/5yrr9VHcsnboGMtBKy4VRO3Xyh0Qdbt/p65MlurDAG9JnJF6u9PYajXQEr4KTnQSTRBUA
iGF8T8+N3qCek0vDBLbNQHaXMrTaWFrltPIY5knO7gMEWvtjHBdlg1L96QAck0CwuxzERYB5C5Hz
DVjwbP7iCwzwzywtviRCqx4CWrBh6DuKiicPqy3ElTXUndIwCsiNwehjWh0G+MZ9Mtq02cQd51c5
0Qybwj5jCwT7cxBanmQbDbJGoMbC/cPDAFaAvBnlHtEKv/GPeY8+DchFUBcOHiZY/8T++p65rLqJ
J2BUTqdT/k/RbufkAPnYkwXOtPJBSJA7FzYkJX36m4imt8ag6vRWu4SlGG7xMaYarryp9vnJAZ5G
E5/T9SFuOJGSASKLnBtHytj4RmNdwGE/+2BsllYF0XaDkWsC7pYG50cFF1jNxo/tjhIZ1V0kjUUR
+UmYilcteUW2WMJOmFX8Ln1tyJts+7zEdhX6iDZr0+jNWvJlL7YYRWSyOGzI2t1xZNNvdWp/AgpE
902lVgKD7UamG09F0x4/0pqaHbCQsldRDRZzcq0jZMJGzO1VA3TOcIksMapW7l08JDzCjR1cXdFA
dKXO/UdI79q0TthKUsD5817iPyL1xCpgtURX1O/CYiAvcoym5LlCg9OT+1LdLc+Vn7QXWOlEjM0I
f7ckd4PYg4jlghN6OH3iDGrBuS53SC8cD5FsRfQFzyReY3eqeCig2N7BvCahCiIcWxbkCe7S3+b+
IfWJqt4Tzvv6FnACE/ENBSGbdkpttIiDrPoWjVeUwRDmdb3IjjIlVtyma3Rn33qWPTUSysuzq6zd
xBoUMY+TrToEIf4I3MCcmH9SdDLj92SjJXuQ+kpZyTBsdUDsWerXcsbuFdZJI4UvtKF+DSri+ay8
Ir0fvBmibQuotc3xNxs5MJw4r+wBFY8bn+poZCdpdxwtwJPaC5mc5/AP+I2VjSr/re1VzubaPGig
fkER9L+acwYGxfYwjLW+FIsOVsjU6ccFO+wRqT1JWqJw1vo1fZlm9LNTkwc0fYPDriDY3ebjVQQe
osHulRJerxDgEjK9zVUMHb3UVehX6RHAPU6lwaGHlyg6sM/0qRAWVo9BXdfvjE7rYIjcAR+C0Y1g
1oZkJWJnAp/Gg1AFn9+gyH3Bx9LtCRq9gBzsGYIil6scVC9wO0rMDhFCyXpXxS4aETDHPZU5EwZd
3R8/YKIFS1p8qVHcawEu2ZxcWwvTvGAp2lYQmRQkU9bvVCmJVWt/aPaWbxx15+86nqt3eLnQbACw
wkxnAqdY17+rmKa8zTA8HQROx0owPrTPG5g9846ct14jwnD6WaBOcyJ0BVNK6Td4i+ExJGxT0or6
a7YSPqa0lbrnBSoavSXJzNIFXkEWT/rRe3KLRB7L4l+r/xGwumIJdw4NPFzWZ3xQh3+OJzshqngX
bWcZda2HU8HBTCjJfc6g2WjVB4lQ3m1dMJLi8qXmpKwi8AB1043iwH63ONdrddG8QGYLizcuEJBJ
ZkCRAxo3CpN7/WYuqqdmNgCyi6Nu35l0zKT9bnwpJG5H6vUKtO6CDluPTF1Nz74zPrX3XIsv51A/
HAkRh+CVZKgDKndUgCrhZCy/R0IbXB1nS86S957G0PIYzcRv9uLjt57UZi3Q6SBQtQ5vuLalcl+r
dxjwwwiK3rwc409Qj6VgGWLB31usPWqbv4gzDZXdQTh3+t82aNCXcDxaoHdancSXTAtD40Bzrgwd
9L4qlo+M48nQ0gM2b3jLu8XGxJlBkk282KQ31z4ayfdD0fPVF8MMF+uFyttICXaas3C94Q6/Thm3
VaNl1wDNK1WfDDculwZp5rHD2pbPCUshWCWnCVnX28MTEqWqipI0WGqxF+lxhD70WJblYovBls0R
FE7pTT3obpuoVPqd6+Gl24FJNJ6a8ujg9IGACELWqULEo85nbwRYCvyBy+n/rGYbSGc+NdgwuhKF
NCozarGxco6IGudEzXHEZOmNt8+3gJCM5QhhaLEeCK6KE0tx/HX15hteSuwdJPpUm0TCgAFR9Ano
8iQwj1Ate7mocW6uhnd+tYIYrXO97LQInChOpVz4mUlqkOTLvVyiP2hAmBwOQQz+/wz3NQAcY63H
I2+h5fo0LgncuaxwRlq9k5L4hRhMnOjEgRc2lKUgtttdd0WHj7GTqM8zP2Oq0ybuUJbPXRdhpuok
aKRsHqBQoY8rU4V/Ie0+wJBHIXCiPNuQVXs9OMj2pgKSG5gKxnMwbT1uyJjy1xmNhHwZdSiFeNaX
C80jmKe8Rm9JMhgUjibbpV9yawuG7u5nRTatlf/UT0trYfborM0UJuOswFLmT7ryBc2Wr6mH6KGo
UCcxGwI4aN/HuzcqJLDGOo3yg1+1PyGq2UAeTwWF8uuiDPUXSGHxSkjMhchjFGJnemZ+Hcj/k+AH
Trnb6PsHPwSjgrxT3CL0yejCoYxRgPoEseHq0z/qyl8hJerhhBr4IegbIEEXoz55vEOzOa/w4uYm
qXzjcSzbs10+nyyK0HdsIWJ5lp/g6/yMEv+krkcvNhz8il7eDaoFHQWtTDEo9EJWlcv2ygQ52HZk
fG7Xih9IoVR3F5cTp4RRYomwj3nsJqJxe5J25GRzBIYpNnqQvQHu3b7lnjwj4zA8p6a948iW3ems
8ewPztTIIBWIR9aVhjo+Chnu/2S8S69O5cyV59ORM3pBikQB+VzNJ/TIBSBNYyBf40/oAGV70P9F
dibjAYbISXs/vhfdjcfKYOQAf0wHIAl5ASZkmoE1/6Y2b34eaF+odkoLro1m4acszBMm8gn7gpuO
m6sHNlAMtzSPV5cOy5k+fX3x0NDwK8yy64RlvThx1YNNe8k19chcVZA/LRC+bKCbCKpPeiutwL0B
gpT56adXJib25s+8gYjfPUfNDT+j5J85d8kSlmU4zvYhNRRAC41RVQvsakF80wU5ajbGEx4gq77s
etR7G87mUAzxlt8d6WPSqX0JrGSpwYJRxLZwHlgxB8L3aveUtqvwa7OtzsTrzO1xa91V4LoL7VJh
ePs8xgFjN8EijuRPMxyNBNWZy6TrO8al3u4vJ+B+vgcXoiPWOM407oYxCZ+KTI9XT+PEGsRQyeaN
oYrFtbcDPQT4q38YQYSltJ0tjjPNTtTJg8mj1AIPc8DsmQFdcBL9CczjLqwXEkKnrcvQzhTCYRew
ECsOvS0wJMre/K7tFDRskrilhV28xlZhHLRsZ6nULWo9/hj6W/X5cgWrpbYDyF6JK8WUPHlzFQwr
44AYfporkoFYmqJjy5nIvjbYXMYO5xTV0LQU1VPuj3nY7cxcGmfG++UvYwjA7KLg7JMzNDeKG4Dm
I2JWWNZNxNvLosK0WO+Pbmf8yGuP6NUOk2ujCnePbjp/IEj9ODQALlt0cu8ggYxodnkDCAKAUvEV
6HNmi1Q7GMPOAewc5DuPZJb1TJNl0U1wkR0R+IiEo0/CTIJ/AMQb6s7RUpM7KzGkSuZA8pqqDx/d
5ebOuycurdooMw5t1HboSxNEXPD07b5DAwdGPSNI1wLGxvPBqKVuOc4clZexeXfZsgfTNYZK2hsG
YBUWgzJv9jdbadlFpdcKjakMo5BIMtY816bClxTp1OyhT7nh5ClN9p4/EZoCZnkC5m9FD1TPrBL7
atqht9MRmWGa8c9tsKLB6vZQBajX/BuTlI3V6Ofbj4+6gogGtl22Zw2+mfkTKBCdKXyNPjBKCLj8
SXf+FbJul5gHvVWdbaxsoCljdJ1OmEwG9aAzsydYvqKxvoGzD236TelkVfTfTAgSFgPrc+/518qM
2ZvFSZl1GsejPl4EAQfpsOBDF+2XIPHyxDifXNv4jzf6hea3oeU6QHNRPygzwAs/Xro9fBtf/YH+
HT4k80u8GyCDM9YCZvDXsHgp85uDhfyKwQIcy01dwRI0hkITO7WHtMX/hbaCNZdO9+3uRa+Z5J1j
F0Q++NhcwO82eGfNrcKf27nIL9Fwd4xbY0NzUNvNz6KbYdWc7tg+iDS38Bj96vw8ELzJIvfFN1GP
O4k4JoJ6stzQHlO8CLaQZ62cZrnTfQRw8nGet+kXV+QOkw7jq8Mu4haAqIuujQ8yWnN9CvL1BTIT
Ex2ef91+UgCMTvQRWWkJvCI0IoMxO2QZkDUS8DQ94r52bw7YNuOu8DA7GMjG/BYsPYCbteiHK/nL
gDLEcLGeyGgm34udiZIfT+ZYU5cirtSNQGriReQRFUpE3mlehcZJevpVrZZocN6R+d5BwwukahLK
l9M7N285Qn4Mbr/5ZM3CzgvPP+rBMZjxhncING3NoVpy15Ar2q5lv36D//zvqFf4+OGQ3zEgfsza
lq2MtEj43QVLUtq8Cbo1CWZXmZkyOKJQapmNkjuC2L6jAzURYC8LXJ250paf1sCeFkKEJxTpXqcs
QB3Edg7j5NO1MLYsezgMUlGNfiK6e5ISBx8nCOD8gtwC9a/6tORFE8vDenlXAVyhvDVKrMjaaE4X
txUEFVPFzr9mobS+OGKGxgVJ0wOHUvFugD7wB3M7cG1un9Xy5LOcTbyzfdUjzJJE5jG0JCS1EaIo
EkhIvYUdhxj0/AQwLH0vcVuTYkgCQ1CRkhqBPUmx70itW2Bm7qwGxeaYpfULFBkQFJUIlOZj/0KL
0t9T1qAMKBrpqR8XFUvOHGYwpbZQ0Xr+QDJZPDA4UYBU5h/KNjwhhlLJLy2nPV6MBkcJlxMwdWYv
RE3Pz+z123H5SqGMWHmylaHWJABD68/6wSyh5f+iGCnzdo2e7H/xUa3eWa41dOcPHhNYih1qQPIW
7hzESnslFkZ9ekpFO2P2YwsJqLYCP9UcliCgZ4fuJSadj0W6GCbL1oJ5i65VYCl6mLj3SKbcMlMy
fEwu1qjFunRZSfYm8x34tBADhniwQuEWDI9fhdOcQa5wtSyUfCDBIVHBAnzGuqB9JdasM8CJdnwg
vSgzMCjARvQPtKUA20ZkVhxJy73DOpP404FjNeMgduFL5M7pCfLVj7Zhpm+p8janRl4H4WozT4gO
zFusA3Zz/4gGL4CdNiW7wkEsyJBixHc4SJmMdUuoZaSOPX6zXy2DPfru4D2YN1wn3ymc1aYCC+jm
lc61bHXs/KhRFRV71sP6QHLR7mU7SQK0+YYvKKHWN3Rb10SQTqkg82827hc3GrQXaX92oA1Lwpuc
3Knqs96hbHt1DQ4UaJDOpVcrGG5fgdqu/pekreRMcAC15QJj+k3g32/Z4cY2+k8h1aC9kp3KNQsQ
Kj+qSyWpQ5A+3S6AJiP1cfFlRPo5JSLq+yrwcRiS/SkrY7wR6LFvqoW0uhfueVg2U6AwSd6EEZoJ
vpTMXhNbWaslMFaPoF+t8JfMZ57h8A0fb+dxH72xdr5aJBbJvt7mlwcAH11mSSGyfFwTQBgJiUOr
g77Uq8gCB0lSu/doDyjnxSVBo1HSKiNoo08Q6OOA0XlSdNkpZhboN1c++1VDMhuZfoiF8MBYQ4FN
41z0PM0aj+RNm3zwGjdUyCQDJkF5oFJf+eJtOudL9A/95VbKQibggG+X4h3hYJWoq+5PHSqjtMT2
ICqYjaNlVlVvn5kmoTN3RcUcN76WoOZaUCdkBGm0VXKtjBPxYwtcCbPpDK2OGo5BYj306OPrjr0N
h6LtTi+UxQbDrAFp1e6d0ykogqXlhkYXUoQrTGVER8JuOz/Grr9TjdLJ6FKDmIFD0cz0n+XejdMx
9IRCPix+wRocVyH0YxG1aa6Q0M7vvbYHSJc9g8gBk9QeXJiyz9OY3mPGUbH44lCzqIfqBtJaGb/0
8V4jbD6joyUotj1KVDmLkY+6Neh2dlp8mYMQFLu4VmVT5H2JltmCfRoLrgRtw+rq9nX1IRPvfNYI
0xW8AEbEr8dwxkHHvMQi/magxIfb0t7q6+eq6XnhIUjxcCf4iq6dMBu2xNelhmNcUs25ybiSlx1q
+j2RU5a04evG63SdYoTw3m2RCuikDKFGHGWYpr/e9Q+9p99YssVPIHoSkuHLw06PVPlmN6MyXbvl
oicIW/b/ISPtBkirjyzECdKN19TPxMHggN/7czItOn1SBbN8JuNs39vL0dv5v2P/nyaV+RmqMR9Q
6Ze+5B/D36DjmWUS6PwE+7jumQeFTqfSox8Ey1Q8e5vN1z4StK0A2S65VIUloZYkL5+DrxJcuDR4
skKzdD/JTYYsFb4UhqFppkOLB7KjyLi1hhvqi1WS1wtSv6ETDJ3eXiHq/9oJXDKLKmoZdBtU7NMk
Ge8g8IyHN92y31hjEYzDI3WbA6jMSuZRD21w/tU3y0SkFezGwvSUWKaHUcBfc82LKqh5yK7WVR89
DsbGd48z8QLnmP2iNlIuVJI1y7Njmua12nyfXpFvt3Wdu5Vt3nQ6U+7wOGslLPDYnEaWoRgK+Zvl
MH69xITba9B1DHPirQCOmVVGp0l2J8p0cmJz49tNp8dmbtKkQ+ZPe8FalrkcQFz9re6GTh9wUQKM
ndm1ekjR5NIlUvfXLSS1iNbfMku9e4ibyaqzM+PO26OL1JZ5zGdiP0FWFGDsR3Rl61m450r11YfY
ybLfrDSvbBSNRCH8Zm2dnoEw13RmG5vTHVtLM1+eni1cJN2mwJqqQFkXkytewaUOSpSo/gWXyvbs
tXzZf6gYomWZbQ/ali2rFe8j7hb+zpnssYtuZfZg/KkTgaMo61Ti74oWvc4MMmWodGONr9pP2+Go
bJUopL8kZu+v04Yc0Eugkb2/xQO9ZhzbZYe3/QU+ne6lPNxqBvhg6NC/Yif73WEBQJwD0Q3lGIwL
+x99LMasaz/cc4XixjD1b8YN+0oc4w8xRYO/8/YlTIuX+y4FvZZ1oMR9uAgKh0xlVJTALEh7kFxc
Et8Veo3Twef8Mml4KJNvr1EyChv+jQfNa2P91oSISfmGsTyMfyGwl0T9TTQkb2XNqaRZZP3t1NqW
NJbNmOY4NQtrDr0SmO4qiunvY0n/EBbBwn3M7rS6pMFnD46uPmKm0ASAyO22FEsH5axJYpqijavw
Nk6ZgpQjGRTwTEAN38lmDgQOphujKnsXoGEpGSXRP5a5MkMBl887M9ZCSdbdI1ol4WI/j0GzbYir
j85eMLQY0EdqjQ3qEZ6ujZODzbzjhemXM+0hcHXDhaiGoF/193k50zhT5h1UfqtkHEVXVNp5bvNi
OlGdMcvjAU7DmNJSLsUmcPA09C7bXYgq2sbdv8nllaKII8HriSz3a0AaoARWRdsxLGTHWqw5swe0
1Ns3CC0tsja5gfUfsZHxwshbSIeFgpM2MoOQZY5xPZpy9HoqgxMiAEyze2d58yLg88oPyUciTm5u
X51ODtef8y2V6kOrSODAuTtJIDdIma/qyOPbnr4CjEXCXgh4ogJLd1hH34Hu9fdeEsZx0dVKHB+x
HrR+7tHcJR1I5U3ZOA7gKm2rzJvvMX9envZa81eNPF2qcMfpxWXWsnJuO3Wqh2FYPuTQTBAzd9b0
NZpKZwourz0HeQpGMXCfOsLIr3mFBqM0+H28hKaFjmUvwEa3hK9EdzfnSHXvVCoSKhvVc4b/ThG4
ritAgjvgDFCLFS9csOcXF12bHdVPfuE5FwDC2VBu6HtIIvRXBNbTKOQfFkYTDnyS6CDo/2gWP90u
gFZ50G9jXJ+1lgylY+obIxF7SCgi4AdzSxUHGnplD3y7C6jy9U0Mqm7qKpW5Obzs2IF/CByk+ee4
Q846vJJIM6UrcoiB/LBOAzQTPBSNN6nwsmn1OqdiKbaD1Ovoyf9XqWDmXBwoJ+dtnmNDxBtej7t7
JUD1ibjQIYPbcZltuxg4Bsy5Bd/A3AaCBrRBKNBZVUt6RsrElipfXFJ5PoTfdaaNXykm2vPLIdPy
9xCGC8boDuV83gKy81BteCj4KTRiXgMme00lxsVy+l9pOZXE7eu+j0gx2ut3lR0VWdOSFIF74GhS
AZWubZ/N5MwfOVL+RacSfA8MfX4cReR1wRkROKLSP/m53eZJzsdX4wT0d9wHBXSxfoLJoXAPYrfp
AL2h69GaaM9V7L/KKwXgX31mCPCoWB5XsTFwtMYMLI8XY6J3y8h1Np0Qa66mfOVwYOkVCRuetNtm
Sm2VIOn9TFw6eQ0rJ4IBCNwNnD6J8aF+Bn+MSErAqsBFuG56sHO0ivI+k9PtV1vYZPDZcziftCYu
OAJcfzZSkO6KKj9CkCKDNPQg7Ctx8E7Js99kB/Nk7w+jwUVw8Djym9/dtM4MrsjD+N+43PshlEMd
9Acar0WzGqWxS/dAhYP+Da1j1T1NH0JJEwadtbeojaS+AUU/ut/SGDdu8CtO3y7K9HIlS2krPcNa
mJo94Y4sjWbD3nzptoTUdAddv3PPqrZtNgnHA/PObqTKfwbVmGoRL42KLANtGBTEJHDBD2KmVRKI
FT4YCNlw3tu5/2mE9/ePoQ31PTG9ykzGFavzRDrLzhVty3hulC5enQUhfHdbxrtUW+dMXSzzIY6r
KdNhdno5eE1jmwfLdVV8Ox37j4jJ8eY90ju/ZH+b3kSi/ge85B7FEeI3CW6I2oj2V0uqI5tMa3B/
tAaC1J3h879W59dAE6/5qdnUpGqj7V0qyGa2n4ePpdGzlXyU1hfoPlAFlpKBQqtNQDXL5N+Q6oYC
aK6btZ6WFC08vYD37TpD/FMLjdSbdEhUZ75gHJcfs+W/j9dPIlqLhAVXVlYicJ55OfbI+psDBv1O
LvUhUcaxc/i9o/Ld9S4k9uXHvPGRnzvbdaw6Ic/UAaXqjVBASrWkALWAZEmlU+E+pUjel0UgAETD
TUd+UVW9W+1FNL5i6Ec58qmHr1tUI3PEQBzECTqNoW833k56eIxEnvsPYHIn8q47l2FZ05tRwz28
w9nHcVBf3vGcQTmE0h0/ASP9BOS++8kg5qOBSVKFOgD42A/HzibOuH7cBYd9C8hzh+1xvkr+qY9b
0TnAaXglUIcXVTIhjxBXJ2Z7Ki9QqSBqrjXlONXrkTlbL7Splc27rGAXkBh/c7n8iB7iLbP8rUmQ
CsUu7tAngU8C5UyxgWJnHmko53qCP/Ei2AIzIneqSssv/2Vmxi0HBcdQaY1Vdx1rdqRBMVhXX1hE
BC6L95iNfAeLg/VuUQxoBkae3bmE/3V1gsmbqXJ3tz2JXm1GxlWoACvhv80l3pNoct4q0ZnXWcoK
Dxik6qJAnadj+3DMqmm21SYu4RaNUVLubZDUPpY5+B40Dthow34z5Y/giHO4EMQw90UlO6LtZ1Rd
RTICmytYHIQzaAt2Dcia8bjToeezv+vL6hMUr2Typo3F2hPTOOkJrJOguK3nXbQMJXiyMLbMwdzD
pTZPFvSKrdQTvw7qKbRpotUByusVI+Na4WtKba6rvyuO1GHSJaVI3tdeoy2YYsca0MsTQpLLEUo+
Np1spXX82s5sCF/a+32MVykY4z56SZYB0/sybfUM7k93bO9FAotgKck9zDeT66CHAz8l8qdcq13n
MvfEhxgu3ERD43mplKE8XgoAd1HXaV78ropR1QXIQfQCPZUSlJMVso71bkqUHxUthlh0ycRYVq0a
21qY4JScDb844u8Si54J6lF9DiAXgizYW4Jbo9ru4bDBiSt5i31L2xO1aQwyYt4H1lT69TgPuI3y
rSHBN4hE8G+mce8euyV3697DQo2buLvp6FdYB7rFb6Vy2yCEqO0B/X4oCfQRcgpOKl3cj6LEWTc5
af9Wwim248HujYD0hUIsfGP+3NWRHOH2a1UKXwG9hZW52aUnkn6J+q4Bz11oA0TsAcDFACtFcEC/
Mk0uzAN0VvpBviARB4hidfKQeEYGVETMc85FbXLSYlWywPoevKByDEAXPL29SbV+F4KsufNie9t2
Fx0cUIWIv44iSKy8bqnDDXZOewEKCUnhjDga2aAbeiW3vRhbjMscrvLTlrz6KQ+CORVa/FpMWrae
HeiAiA09O3g4Te8UvrRlhuuJYra0Q51YA6dxqmR2guXmqrqnHLww2LWMI8Uqf6VWMQfWibYUZn9Z
wDAsk5fKkHzwseVZI0opcjOh5xy0h9SpljOsNsfarSXZdm1ff8jBqDo8JWuiOe61ppAKKMaMNEbQ
MkxwMFlZq5nRWfzVLZBAvRXRGiAtcvaXS9+91/WCf6Zs/oQmXqFUYFz27rslmJ2zRXd9sMkkF8KZ
J8FR7w3Y9pVAAr11VxROSJAmXSq++s0zE2OnyJME2Zgt0svImnbKOaSZR2JDBP7bvxPLjTylgDAO
hKCv0QUemBFbG4a8fck6gBVFFfolP56JreP7+Hhld01z0Y17gon2SZ91xTIONoJq6wBsZZMyPDFZ
jHIvJHb70GKVi7oFnMtaFtR/aXC0swwy/0uBKyw8uwalKiNnWeZdaVcIKkEupWZspYqdNQtXQX1f
JJgXLWrOZj4v18hPcbDQ2NGS+FOusTmoeZoj72tMPcbHsg21vGFoAOU0TJBilGQSgKd6iyX6xlBT
EgLJFA98wJCYMwSak6AlDG2Q59GthRtUgGvkbWXtoMg4QuTawmmtUdbTcd88Zw6b0i5JTPE/DWmU
MI1bTx/Q4Ix2AmUoH9bnw34+5vgaiVgoGcvy7wEYFiHBriAMEpjSFuhADW9aNqtlX1oKPNHi+Ncq
xzvU3moIzZk76kO3e8bOco1ZBgTCLD0tKDOulXzH0Hi0V7o+/fSb2y4AKSW9D3ViL1W4zi/o+Gf1
A79GbhypfnursajVNL+NNOwZUM68dSJxkzCP64q8uWbhPsZ3iAYXEKs14ziMCd4r2zu+/J5Cp+9J
OdbG4e8Ehq5TrTjUMk/2g4XFmtYq9j8dL71VWV/dZDoaBknhyCVQeEbyUM1NFmlFE9iZxJLfTOR/
10DUsPVPGamkZpoe8HIWZ8IHno1ADsJdpzl1+sqBjrkMv0Tub8e47dGpQ59Ur5yuU5gR8fMKBYQG
uzaW/bZdEhvT8e46Y2oo6wRRcJ4qLot+L64ecTShqc9izG6Hrke31iDMijOrJ93lXHE3Z+hWymdM
l0XGFkhM+ZF/pawYliJqklLRlORAE4whjf271RCitAhhztCQ3ER0gfC5yiPb4dDWsvvW/438b1oB
A/vtb/eoqRoP/UsOu7LqwESqQo6/Ow3xgcco7mw+QNbevC3Y8bxS3WX3Q9yQssKmgFXf23CM+alR
2KYblHujj13gUUnAE8uO0M+GUz0RSMegkqBYoUnbSpMywBMEtSbDuBl2Y+T8qYl36hoEXfErW2I2
hilYeL9DVMTEyRZwQxphbtFAmIOypHL/qc3pp2nFo6JdtcfV8c6pnQTqdneXRwzlS13ueZofPtkT
PC3tAa9EdXTz+0XWIrmbw8PWrwjugOVHxeMzXScJJtIDONX83hyq3M2nW/cwW82pXWaClVKX0Ipn
C0k3243s1SkB+Um5Yg0/huxEo6BKFBB43wNLMq+GpH3SaGEYHtuEzwpX1vGMQYd5jkHhkB7J9kpF
UKAv7WFDi4zqHtQuJNCjWFp1SWP8wLUgHBg4eFXgDmp4R8UD0rlDM90qaNy2viZCvfwGo2mPmbu/
z1Loz76z3U5n+OahAN4oPitcYiv4Kw8Y7X7pbV9FpdBLFnq5mqFfLsnZFtabasdpqObWWIdbreum
YdDBYxKa6YNpKGwqPh7ik8AIcyym2051El3l3G57DtquOxJPc8UTwQiPhfENxqBpIJ8xwTWv7GwJ
6JORXzKYm9qgksIRRQ6sFXA1D/eZzNxBsPYd3p4lYlCXKLRT8MMKDOsSFCIhEibUEmC7bxrbz2b7
cARQhuObRelxrX6+sQLaG9K/Id12w4n9YLFDvW2bnbU+zBTr8Hzmx5JlRHy7ajP1fkGoJsCsHkz5
MPnMLyLcIG+RjfVJA0glVyC69aGZIHgt0WBdpiqs1irfbxpZx/CHTaplLKKWuQPiq9B5GasYmjsd
e+ilTpjP3faHRp9PRjHh1trgvVKXFdmCOzyYiHcgBulLcd+c3IQUQDcPD/kzqKaz2VTq7kLyPcM1
MxWUTND0mYAXn8r2sq9KBCm4+fDvW5dGTRTj4kspw75zyPgHQJ7e5MC1XeDLNdElRtb+XuJu5DGO
3b7/S6SMcKBig/zm5I7ksE98Seazb/z8F0GqXasJlOHwtxmN9v+Xha7YdRgMS2fMbklV9lU8BKhr
do16HaOAm6pE+Puhm0VANw9dvZiZSFcDKRM7ejQW9jXJq8pUnjz5cGtMXJ0tWbT76Dop1qs0ULe6
0u9OSHJ+/odaDtsmNAx7pAQMEGDz3h6Ta3U3rWNWYoGLytJzOc4fw4329szFHaNkF1gpIkpeCSTT
ygEJNNhTm2QbvoxDcMmkPB8TDb3KMHzexxNmMEZmX2rIiUhSOruZktAYvzwhDEiYQoOGR6JetD/a
aniN3u79caCBDo3p1R5OPM1knbc++83WC6rk7blsT87qFA8wR/2zU3nWpGSKiAlYNpnIFB8CjyxE
4fzzFIkKU3oGf32y2U7dJzIC+Hse+0DNYScGa1Gj+Km/xMFqbSXI3oJz7CbSIeW6y9EclLd5s6BE
sS9XufOs41WRmUgkDB1akf04u5mHMmvHkZi9tXyrxE9+zgUD+d00P96eC9Np0+8Yhg2TQT/NUmLc
3sOWccEgRdXIGxuD8wZSpQQwDE57puEVCjhtGwwRj1y8wM2YRv2fbmGHcV1nSSPQzttoV6r6dEAA
p1oUptLy+QP/c5toXEZ9RDxq0jymleTBQgcalRieT7Crb9rXXFgXzvxR/Lcb4iRXggg95ZqKiQH3
ehUv1JB+Up7835PEZiwvCe6ytAG5Er0FUtrcMSEqSrGB6wucpypwwyiwPADeZ3xw3OGJcldmizYx
oMdPmMzu3l3C+Lhe6GjQ2ZsjHo4MAQjvR097JgJivtq8MV7HGAxNtxlCwepRi8uiB9CM1Jb3rbhl
/FI+3KgvZb4LcTI92AV/2yXnaOcaIU+dZtBwQxQOqUkyMHh5Oqn3TiPKi5ZDp3xXwu10rOI6IDEz
olwFuOHojeuHUlnio/ZBWpIhvRFj/0l+yyJG63O34KEiTMNw6v670RXNq1gfeWR/gu3Fh9ERaJyY
3XTH5VEtqTQp6mqTXbiZCvM0GenF/Szw0tYwvPUJ1vBvEGDKDr0Z0b/pr/p4B71Zj3oqUdFrj3gl
tsuVB3i9a7Gk2hOelBQbuxFQQWUZJS3QCvDww1UR0lDXkNjis3mX6emL/Z8KqaM1yJ/PUbnnulDp
z7lNEzVgWqzpfAAqeqZTrQN3Kf6TRPVtCZY7Ikc0WjYcmyr50athu5cXv2SD8phLGsBl2bXar1np
XYA5b/lgamxLq1QxYSgj7oRlx2hXzIJuT2PpWS/LpgbWf3aH79KdeR2X4JSD0vSjnrdwc4tvSK8c
cgGZ1Fsp8sqsoAlhffc3vgFs5iNNbjyRBOif1FCmlZevYvOwXfxmNda+MFka51GIjw05wIu0tazJ
kKjXkAPzc7jc4pTuqMJt9wrFyuBE4JVfQ88RpYSR05CtEUZlCQgw3e+SsZw8K/vqt255Nx9Z+cyv
7UYRPCvBchcwGfHJ9H2U010aNXUc89dm6VKnzIbAlljWeF2QWUuoLJ8kkuR1mbngJ8p4ECR4YJPx
dtIT7eazWH1diBX3WmZBYpZeSzp9LglOBcC0gNTOazMKYlIHEsVMWeeSaAzZvt5Fc85eGx5hAJjc
/FWAr+lIGJ+pyqyz8thDx/ZBzwHXhNcDNztqNt6GKvbtjH97udJ7YeTYY8SDO0phfi33WONMoyR/
BysjGSXy51o8a89wk2PPlORi79V4sbZJhj18XcaJA4X4IuERCRa24oP+5iM5PMqCulSc5DXp6te0
EKTJN9nLih4lQBDVUKl33rpzoi/5NOvTvJdh0c8gJcJMX41oxFX5ThqGEx/45ODZmLWAR/akh3gS
bN9eejJ7RGm90f4s/M3pt6g+51936EUJnBzBp4wEwUC5v3xwDnzObfaG52lPi9Tq4g6fq4SzX7un
saCicom+Rc1L1/Cun6J+8hPRPCsyWOfk5J1tK6zlr1jRo1REG7o0NuIJBEoPEOlj1EgM5a+ukWID
hLISAyNDYCfnEH5KlrktVpcMVRNq9Vi/7fNK4m45gy3su77tX01IHeW9c548u1atDmGIVwKv6UZf
s9h+V5ug9uHKy1zR03U02FgCaksjygX+4kc7o3tpiADcVBr5wSHBcwUiH8eehEO6ZTcyvWKWaLm+
QpjKnzHLuwM3Mopl9KJS5DP2IgtoI6pP7oxp88PjcdhfE7dUyCqD24Gpl4g0RhS01kybGO2AzolE
7129yf5Djxq3NsEWy2tFNPE8EPCDOaOhpcQhfaMw5Mbe2q+o0LKWmHVLNDkgKWCPknXUdDEvJamL
hNOUSkAKQnUt9vF0kFUxi2yh6Cry/IC+jXaZS8MYdpJTD01iCd1FxREKK7ul/5qtIWekDwO9nFV9
LT7cmC0hPyxx/m58nhwi00VADecaXaiMe8axXSk81rxYVhVDyI3uIiblMe1fd1ThLegt8MVxdVNV
3w+3f2fYwWu/ZAlyUd3dT3TtU1v7vsZVHW9v63A/38RQKqutK4+r7t33D+E1ZCVkPqnmA6o/d/Bc
ndITZE5W3FD0JgHZUUeJqHLVPdJynnE/Hg9MhUoPFfjiq7jsYN9qC5r1MTFs1nag2d6UctNn22j1
RcvFwM+IQX6V6YFJG6NtIEd0ibop2/QvQQQHym02BT4B8XhjIisYMkeVWYYr/yca5te1wDGlR+vq
CTuqCa0hHe1paTKFoeKWsZCliT/b/JzuKW4VaIR49yGGFbyK3YmYLGDkUpJPzomfkenis/0ZZjyB
9Aa7MSKrQ3InilJ8IMfcsVOmFOpDSGUpNzoyUWJd2ZyXJ3vJ1L5ApipX47NSPUOam45cGjct82cx
YADBoT+lMSNlTwVJ6OEWPiGslzb0+sUO07nJDfVBuCS1LcDhSWiD5fD7+V+bB+7hkdgPjVm+CtIK
SfS0PGQ0WbiUy+WIhipNISBaCXZHdyKQP7hRkggUHz5g+E8QUKJOdSkAtwzTB+zcpmis8vAZz/19
CosZh8JchluhFzByuL1YCWG9pcvZtdtFNfFY1U8Tw+5+yUH/7ygDRQAqn1wJeYDyPDzW1q0I3fcO
FoMzRUpBWPKpVz/QXNixZGqKpXja38TckJtjHko99+FmFZ18jpBsnuZTopuTfJXJAgnxplMxzZlA
JsjFFnD98LXjjaZK2DPxyVPsJ9enkhA0jGZ8c0hUFjgXdor+OXPuXTQLbZpkNuNU7y+k/0Rv1BYD
/j6ZcMUEOsFXM2/BvivWnNx7J/Y0XlxgCqxRIbC05zCy7w61GLXI0hq2m5sGlW5mX9nBfZVPr/jB
AZxRiiT6PO62853DNvxXWJapmpgb+a7Bfr3mbY+bh6WAKmMBsbipx/jxfK5gXZtFAv39DvLySsoG
gqIDZLKRkQJwBRMW+tHoPcsKBv2awLpB1ULRL57S6+ZpupHq+k/hMTBe1sGVo7/GoC++bn7qjvhZ
VfNU9RlJsz4NH5g8p7qs6y3UqstcgdBldICndCa7X22hwK26V/b40kRuP7BbBa17Cb7LL7XJB4rW
sm1Dk/C0uPZbTkib4C7JNxyh5/UU8OKRzaeEtCC0jK8l7aCuZpCpSZpUSmhrgz6DSxdT6lxJ0dHU
v0REJDKMITE/bGOKHJ/WpF+6Dvcffebq8VysxPRk/NZahy5TqnZsIcQm8Ynp09uGeoYbwuat2ucn
8xbbAWjXJ2jLmYc/2LvlGUxrVwlFHNCB7K98F9W1mnnBTb+efoeJQ/WaUN8knhgIbplMa96SQGRt
b4x0UiCKQy2pnBTM/psI/H1Of6tN8S+r32S58PHjmFI7wW5WsA0f2oiYlxnhVM3KWnJvSNEbO6tg
8Zi2oCJV8+pL9LrwtwdSD40VaiV9EtmNap+E0HYVsqI3+vXRwfQuJ50gGZuAetLh6KWuHghZdZHa
/3nNgXhNMFV7uCZyHsD7FCDT1msv6QCjozwNFaSynqY33DICucV0ztLYf/FecZ8tmmx5Q/Ity9fS
OTbG4o+qbVdQKG/uptuhLrlnx3ymBWxLJ92JR5Dhh1l5gC0CoQuz5nFQuDidT73F/pUkYtyBp0O9
oaHkgO9oc22yPh/dfCapeh2nniWByCbPIa58IImnD5gtLTq9x25Obc7Y2Kop37vE/FLhIkkZzWN8
1gaOclzxRP6UHmpaXLYIeYdVwZM+fvERW999YFmuSN3eIrvrRqyeNnxZm1+zDRPM0Z3MoLohtSQz
DM+Tp/fYdnEjAHjsJjVmxspuT6G/OU9V5BOiSC8e42/sxIqEyfr8dMlZe8ogHkPpRP7/GYfotdI7
FvHV6jLinkc373QEAygAmCEWAESwunAdNFx4cpNKqA8YIl9umyBy/ti9zxX8vtCTVwkM4WpUQBcG
Rk1j1k548aaX6mWFCD5BnAtCchOgSZuy6055uSD+x70uXG5CD6C05oej4x4JA5nIcnpu5OQK2R3d
4XxNwDrhG2hSqBbS7PFfYBukfVxoZuYAti5uS1470nwr3Q5GMf0KRlJl637g0mDMPjQWq20tMhsm
IqxvMymsj/8KsoZu3ZMsFgt6gdZ2qdFVQfhePJAzYJ53TxF86II+TGaLV4ju8iZs7DhMQsnS5r+L
AQdQQcCMWwBPZPjL+JTbNAF2PDDGGhi80wmRopbBJWkIdWL1rYvTfwhFh9dQnPtG2xKBwJeHwWSl
AwsdRT1nGaerkJpcdYMYE16M6NldKOBEeRQPmlM+dP2h0NpdKavyIeFCLu8uzumUXGhu8wNqS3ib
e8j+LSNGrWimOCN6EqH0oKUHKPbtgmgazrDBDW6wIzisFsv6b72d30Ii3JEQTcMUWeMXu2x5L3SI
IFlsHVnQitYthe3mcRUvoT534PNOiSKhtfLq9FTpTv7DnkcsZJXybIMEuf4fnA7KtwoEDYdZ5f+n
nPuGp1BDVwF/JiriCdzSjOZq+3FJLeO0OepdSHtmY2VtUT3Gh7TBWChlGnV5U3s9Gfn2xkZSYjLi
iukE7I0rUB7UnxwCimEc23A99VaypSamgjN09B47JH1QzGm9Uu5ymPUrbzIGpYIwp/Aa/34nJ1X6
ITEQUB1jMZ0MhmjTviB8E3jXSgbJX28fSjN/c0QKGdni0tQ1oFKINBQkFA6mC37nPiL/YaBtnIxv
e6XlycQa+U/b1UxSsLEQUdjBUalILaAVK4R16B46OIg8z2zqGxEVgZKBFQ4qsTlQ4f+ZcSXYHdSA
Sd+5iJc8/x3iSrZg0XAzpcwopPoVPvJjEgpKJHNKrOqru4RiK2qvt3ixU5+MA+EGAlgHyjo8E8rm
FpJ7wvn8lkp0N3brgNF9crlisQG81DNTuwAS/EtTYYUfNSUYAy75iD6uh9SBr5P1pB5ppoDTNdto
lVXVo5hRIWZ5Yh/Wnv3SSzWIXMWJSn9iclINYZljMAab32OKwgzDpY1KiH+gNkrll1xumTwKDTwP
Ye9GsuGJlH5/aPJfq5bIpqtvjnu+MMqbGuCXYfTA6Hk6N8lMfAx5Nk+hIX40Cqzu+gcZtD25vLyb
0O2KeI7BNn9g7P8wi7OG+Oxfyq5B78+MRwS+9csyH8SwzCVtjtIGq/QVhfZ25jBHAacuXDvGWp9c
+TdC7iDJSJinCyNNXkIfNsXNbWXKuyVLWaylD4KkU/vRXox1xqmdTpTfgujTvzXceq/SI79kJYtv
GHE5OhH3CEYXtX9BMiajodDmwGoNukbW7cNP4LsQYUBGEtM4isqKAOpS011DN/+YD4KKnz2lWeL7
+kfr0nnLvsSY8b+vfkjEZ5wKKewWJx23Y7NaacQjoSezBI2BteZoJiGi14eSyQNE8PK7FKSQeusi
5pZiPKEsAIdxBXrCW7afrLD2MyDotF2panfM1Rhz/ugc/M8kmUtkOntJPcKCe4paLIJ1FIkE4zEW
0zyQNBSQlV3vvm6s5MPlIalzx+pqJc6OzsxNNNW2hasiahj8EWNYkO2mgx9QtcJnQ1rVyi7jHltM
icAN05LkyYj3YggmREeCWTYtqUwRtG3Dl2hyFSMNmXcQU11LPhvb1MJcxT0uxkOrzQFky0tJG6mb
cMtRF8DtG0lCozhnnVnqZ/c9wOBfA2FDVRL+OSN+5ShqiHGRVmXClS1rZ5VEWsFssWIJqYKlwFl8
9SrtPu7dx/3pQo6F9WUTYkmxiwvwDFD1LQyhvsNfSPp4KY0ZLBeQoAhWtFakjmUJ3gDFMyxX3aJJ
2v0T0Rs/T0p9A3oiYPjJjB872iKyrXYfmvdAdDYmzQXO7z1nT6db2plajCOgP2zMmTpUOk/t/k/G
qCt2OH7bPLRTpWJzBywZhzsv5r0KSFpisue3Eep1P2uIZfpl8HEmH4ypqYcTgAgPZ3QRw8kt/pbh
nPWv6i/84EkdlNMaZZBjAIxWR+qo5TK17XDCZTTcpZuRvbQEiudhbaWz4n6GRDELumq0z4DmLpwe
khWPGB1E8gXMLxnWC/wqnEp4HRGcZ41XyiSeFd0KLUh/UJbV4HojkWBkihP0UmfDQJ+enqr+gXDP
mPsA5IifH1R043qQN+V6ceLNehB0ueyhwME7hRm6q+byCOY0Egt0Vo39g6yAq4F5nYysZZthwaha
Y11pbdAbz4AKyKWEvZMTc1kZFCdk5soHUHdaqDrJZyrRQe09bjfB7Cbl2YguBtaYBWlRZVCxATdd
pgKBnZhpahvXjJ4v0Hc3I5gkaP9K1kQc8/cDq1YPdIWxm1RubTVuF73Lh96GHjSQYXIQ3Mx8Hktv
9qdZmV/60OgG85qJzCDI7Eu7mmu7nwTFk1ZXXBc0zbrLCOqAYogWRfdEY3XR+ixw6ZUtrp4EIfD1
QFOPHfbPY0FaH7+FvanrpUpsBXrVtDpAr/NHxL/WSMfJIK0mx7xKJIggyozy4+KTm2RiA6zAgkQ6
8a916W5MLZoCknFaGaHhm9rKY0nshyApic/vufdurb5dqaWW5UCd4BQ6Yg1AMVq22r4ta+0Drejs
2E41d2wBWXSGJ5qI0dpf8hcBDSu8cLvHvwcg7FTfbo9+qHZPNJmtTZrvd3nWP8Ch41bvf6pHpIxB
eb0JVu65frpR5OFMi+jMJ5W3S3U1DtetX0VcTziSafQaOwQdFaJ9koDTg+iKXCHrgG4KricdzYSE
vdFMJ6Dx2OTYy5F5M3AwT5v8GG4bhkZUKz5nz1oQaIe+fC+V5NUoFRJ5iQ6tmxIcuSwa4bXDYA9z
JNC3EgcWYCR/qZlPbImlnc6WZ3i4rJauPuyDND8S0Q8k+ALvRHU3K2oXjrx0sKk0utvTwfURVmyL
aFtkVkkDf3d3f8BYcVPe5DZKRBfFUXCWG3+jYRx+GygsVPxAf4ySZ+XwSVuDdrvycZtO2ShRxb1H
PyVNwpsU8ENgYseESZpvjKpycbzzi82koMMQDE6lKb2ZVDzg5tKtKb/G+iYdv7eQ4UVQpRngjguw
Qdjrmqx85l/GbTd0KIzxKBjr+LuHGtu8sPl1IYiRt13T/o0aRLrKbqhPtg3quzBQccEH7H5Z5fbr
OuE8g2VgphSh5ay0ZSq5KVS0L7g4bQAfFeX/DuxujWtylDcIIQlmGMsQ5/aa4s201mR2Mc26O7jX
HrylK0dHsBNYJQMgdFl5Uq0db6Tw1CTwUP9E3SX2EsCd0G2YDa+u+0xo44ji5ICz5wnC6Trx65gI
CNJ4rKxtPnmvhFU64stOpBVaPTtTM4ZzSgO3oi35JArZQ8Tnf1FbM/jEl2RxzPHAGPR/ilhOugEk
sQA+c4EyMvJhf81Y47tHq1qo9y0l4/iNJ4/k/eQTO4sWk08ENVJeW4NQLo+K+sIlX3rBzgf0N07Y
FC4RglG+1AW1+UySC3lRSsP1nKbTEO/HxLfxgoQLrgK94tdB2HHRNPONu6v4jm+79OcC25O0vuud
oP8j9N0o/aq8FIir96xxb/pwub/193HNPe60AI6/TA2OCO6/BMHJCbEeY5vhLbTA7sLb+M/I4yUe
HHInzQFWPdCruIIBbrmjFxojcqQL9ItkdzvufWtHkFC+6jLsZel/01xmLt2DYBAMSaWdJic8oXa7
ienF9sMn/B1t3+vZ+JKtt6QpO0+O7hiN4EEuxaRj3Hm2XwFMcKW9dAQHELP9r72AqaWf1apwqs6j
7zbtT93MSLTyFUwwcqlHCBRAQxbZOn0Kki9lkictEmjUNcoJFjniMwxsJ1ewznGFm3GtuEf/xpPc
xQBYvs8pbo9MVNVpgVCs01vhif74/48CuqeRQe9oAVrbs/uONjMdyopYAyU7rpFHHECLIRzkDu7s
tzZyFsbBgzomBi54jmPgCFvSnLqm6s+Qia8Ot/++/qT4+jkmpJXe3R7oV7q8LWM7RVb/ZoaFXkyI
4RPs58uhkkT76sfqC2SJz2H4MuonZrkO+D14zB1dB3bEe6MnfDtVf4F/BOfifvTlDRPm3aNxaNtd
k6zkgKO/Ri01e3gPTkav4rfEQHlrbedvtXTp9ncOeAzTtX3NwfnN5OzhDGCjpPvLX0q/kZLbSSSk
BlGdx70WzqONjJiosRtreV7epVvEUU7Zn+gUVbKuRFgDOf6EXFpw6Z+2WUPFyVL47X16HMegcRzW
WW8WXAV4Iv7KCuByTf7Q71g2KaLkkEm6mysmNQpbfz0kaqk7YmJr5EoJPPrnEDYHQZ6JtbtKZXnH
KoMSOA4rIQXjpk5xtISiV8OSbymgC1vzXaFjq4mpPk/gBcEglcMhYSy2EcMVbPY6+GlD5hhpRfig
+Co1XHj9Ig1yCtDl0iOamjX4Hu4QUQs1Kq/tdlAXMIjQquL5r2czDe+1zM/2zGR589AqZwV40UwN
0+3OE95vIMSIuH6EMjpQ44ExUMYJZ9RBA21GY5Clo1SQeLZ3WtTc5bCwV3s83amVaRzFVxD+rLKx
Ys66lyJTZ4/aTXiQORiKZDntpavAf86Q5YfAAskg8PIUOp+izKYYwd4AtXzpB8ZP2NbW9pu4EzXR
9tgFXfWxJTHpZHg3UIrFJbq6VP1I8WeRtjKkNODImqIBYjqqdXoOrmh/DE2AwE13LLAcEDzNS9kN
qPMDCEEgqIzLGaiFveLoxoE+poZpWfgYjE9CYb5ozX9cDWPMj/63sdTkIhdeQy+FCW4WKSxc1s9A
VfKovnYPnCyFJyCUXoA/u8lOUOillZ6mtUN+cxKoWnMiawgLEHx0bh//oHLsvORH51211MWv+5I3
U41dEfkwq9E1vlgPt3R/7+EoNna6Km793N0CLl7uQsrBdmtDnjfz3A9UyNZKbUPdudBUE7RPE3GG
gvJ0Dc3p5l4EOjMIeL/coBVSJK6kg6g3Onm2jRhxhOU2BZDoCge1nUOd1/QnIS4aH7ti6eL9TmNN
950V3JhsxUUO9sPzT/W2sQIsmKuiKvfYB/wap3wdZe8bFH3ZcqRGwCOH1qa2ugXZAWeFWyIfyoA6
nKZSly3O3w8RAN6WpDe8dmxSZzofBkirnl/phN2/lbCrYRAohp6oypzqDYYCO0hwxmx+yQ9N2hak
4gD/TAyU9JIGIc3S89I5I3CfXD30nl31jfeQNVBrSRiYHqJXwWvstuaIiC+u9pFVJobTRan4xlnb
sq7Kd164i4dVONJiIiicaqdQIKHMbflMCBm0PV61o++HWOO/tFcmSurk5NDTNMCe0ryHLZVKWrJS
etyWhMBAhSsVkXtFGB0J0lpLQuPiMfSFtXB0MoCMHLRj4/sbwe0gkRaHlopt/wluEzIq2WFmRuhm
qbZFy5Bc/Yf8VGyynIv9mhxmvyPdU95heUCZKPDqXJ2aC0JI0Yw28FWUDdB6Pfp7+0oiEEurviYF
p4VBASlRud4YLr9afdnomn5KYn2szMnE4PUgwdkxRBrYnai/49YK58n6bSajyd+sCDySlYrMN9Pk
VtcPE712YHDJXgireQjtQOVMbOlmvUXWD1mHN63YO88jeaH7PAa5cKHX9aDd3aYeYlIc431LHlQQ
7tCBQTLj8fYIKOX/PoWLdNT1KpRsNZC5XR/2nBIWi0qEPG1XK9xPU9R1jyBsWi4Y+FcTGiWlQ8vh
WoSs8Ykt5NDm+rZv7MYT6I8hLl8/f7DxvmTEc5rzjCOIWcL7FA+bT9TiMzwAOkDbC7Jdf6Fd/bvI
Et/blvxa7t88zE7/dJRRTGejAmUDGSysRiHMZC+jomfCeJ0m7NuiHY8m5N9uU+TB24lVYAaHyDrf
GsnQzwg7nb+yLE2ontKV+NTsecpFhG/rYOjRRnLseNvKyQEFkfSUT2GLeBouVG2mll+HPMC/wflg
AAowQRQWcG0pjlnN4eiVMLU/8roJKUIOgBrmbQdNplrHzUEGtLjaLLJ3dpMLdblBuHqjYmdVMfn8
/JeMfb2+w2dojhPRAMV3vCzLVmbD4EDYLbUn+7jn1zP4JNT6v6vf/pjJzVDgWFTprLW0aQZ54fKb
cp0znPbIzsyQIpPf7LJ7ue5V6fCz8Ri2txxWF7unH1eB2Z1QfwDwP2LChxP3mTH/92HqwhXoQqfM
M1v/if7GFkTouytd5jFmYAYetZE0RofyJKQeIrlrCWoEPTYWe6dxYthgd39KmQysdeyjAjwF/u+4
+eR0gQRjjSGnJeXQDVX8bM/Azpggt2snKH4XE5WpoUg8oiJWyNS5EFfHsBk0L0j2+Dkt+Po5zPTN
nHf0DY3xSj7iBFlVlfZWiA9cNlJFoZVES/EYgUNP2o5kEhe9SCM/VC/n830Gk+vAUKmUVq5AEC8C
tjPG71pvgb+UJe4QqSN5/exgzXbjkVwBsWeBI1KESuTJxPDqggABZlOs3pD+0Yd5OBWHH0qiEjPt
WmPAiZe3qWDmCyBGBBI742QLh+kl2TFJDajRVU0oNlUhJCPYdLpDl7Y0fGVVYaBks2lsYT2tlZA3
uKErP/a10Y8L+x7yynOOSKoKGrhlzCtjelC2u0Sz3KuaHJ7oUYiPf5mEZA8Vpe9+t/ETXhg2ca4V
LIGVzpjZFeOxX94aqZSEezWov+HgXP2lSUW8a48Aq+kvAkhkYVCcy5PV57fNTNeSUUQ0LAAkoD9k
dHn3Vm+Louk7hbgMYzosDXlkfbtqn1fWK0nZ7KMQjCHn2HJ/3cb1h7PVK1x5KLh5nx9YopRM38Ob
hgrvqsj8eULo6g9REdgzTJ9JiFIYEbgthHXRDXPpVjnwab1scHI8Ya4PZINEdWkXBFfjmHfA0U4k
Na2NnsfDuK6OUriUsXbTqd00zqY9L1vKxs9GgtqO/R53uD5juYgMQN6kXbvTJcY34ZW11wvxWFrC
VaF3bo833PwQSm+mhajdX5FkdERmwlyuleGaAAeAN13Zu490ADpVtGXBVUz08PIY/8HLt3bO2nng
OJycuENKovZlO8x7Vp4JGUinotDeTnrXq/ebgnBt/lsOfFLZsw4xEfEpcq6H0q836GyHGVDIU/U1
u5XXQ3pv6bQu9Dptlvtp/ByH5UPWPCoJf8EpxLVGMQJPBAWaJMEMN0uilB1a3gzu9VGgFO5MxIS9
/mkGa/GqXlxjl4kTNixnbi8r0DEuOh/MaxendKEdKDqDSAN0CVKOeFTn4W+HrB4YoyFRuKP7DV5Z
5qfJ+OxUDPi9vSVU/qkzcPgbuLaCFNcW6q8nSfg5ZcB3i/GUXcrpeBFxm7XZcofechcTDO9yN5bs
BXItAlJCOKRe4XMkegUh9QnX90uDZog7Zhvi8iKAPJCE/Q/ihEiwpTWfjgrITWrXJ81zuGTc4LsI
c5x0+aWw+H5Pb6lg0oAPCNNol0Wm8SxYzlgC9jMgDovWCxHDWRnevHOkf+2Z+lkn1+U/hN446dvO
jYPbHTX/xGRXlCarZ6ZQxIIVxkMqx/kR5H3Afyx6h+p4+XUskU+X4Q2pog+suHVLBIEAnGpkcb6y
6odcHrIUCKg4AB/TP65IouG+s71wR8OMOm9CuWUwetDIDbHyQfPCpW8QFT8dzJhDcn5VlAxmEnHe
4z+E3jWoGdj9rNmjPweS1kcBSSSpKyNxPJObjoicBDLz3SL2kSbbRVM1ThzVO0McVlwaFGlUVzNQ
a5XVOTh1CPpcO+eku47hzkTTbXduV06qVP3AAfC2AfmVspZQ233s2xipggP5Fkz9UpZQugAKSlYr
0i/mecZGWFQlyT4clO56McnaeE9FHWOHKKqio8gsylrdu+ky/IQf5iSk78MQeenbyf7QoIGCo1hh
5Sod1fakapmxUrihSSwLp9BUgBkhmorUNm6uk4ACq9/qMiDIMyPtftf1DlFm4fsVLvCzx6vMNifm
ZKUeY1I3I6RUTp0k5lTAs3KjBi7tAw7haC1ZdZLiSnS0hrl5OECsP609nxvVZgIMG+CYssQ/JZ0T
/8/BuGGE064EydSuxRtRZdAKIauqjCCeXWvK/m60Y2pLL6SOkxGn64mNOwuASuGvEASINNm4VIxD
c8Xhf9yKkEXSbKsWWSmhYTjqPJy9ZWWqWFZ3Ls3QsRRnqfwYj7ZYR4sg3bBET5TQcTnhOjJdI3Ax
lBUmn5eVrNrGUbizq7tVgtqrO9BiobI+yet0ZyrJWH9f9QIJQE3hCGPzNVBk0owaxoER6RnOFXO3
MuscgSzffp2UrhZr/XJzkwpz3gTfyVMUyYUgc5LpzUnDn01ue6ikJDjkr8N33afS0cLX0/Rlwe4b
5SPKpCM/e9ht8e3LlYuD1QIU/u22Ta/hSn3iH2y5nHttIIhLaN+B969dhO5w8aIHNjdYW6+6i0sL
tjL3JWnMQfCbHZCiktK3KmxSwC6A5Qyhu5ZPZWky7qQI6ozlvrfE7aq02G3co/NlPlQor8QxXSSB
kr3sb/vxAaU7sLGxDT4MiaBiGS87+X4zDnPpsfWGZJZKvuaatOnHB/M2VFUxDF/sS/Bm+jABDLq6
pwbiJJ35AAHzeutxX42RAsJJ6vM2KD8bJyJqolyIdd4abubFMoGTI/wgUKX4PqBmNAa2MoxYae8X
e5d01voRVN0MC07+aCwNEL26Ob0xQCa9Vd5Hw9unpigiZTS5MZIv5r4l75pXHF5bHXpz40KiVis8
QQ9B4DaeJl+R03kTf72UiVfg5iJQpN+fOCGU3wW3C1xny7oihvD6yMVKu1/pjkaOrCexdpZBim6z
qfNwEhuvFftcsjinYqJrmggUzfYTJi/g+bOjriMgxeiCVk/qsdYy9yuzB9EWz+KPr6UzdtZ8zvJU
H9nf3YhlJPv4oZ71WckGoaDkeJfffL7dPqUsZ085xGjYyfEq2cQbHUFIfX0eeuI+Oiilk2x7h7+i
Dtq4SwJobG20qllLisevdj5FGjnI5PxeuWXSPdmi5fDBFUTUOLgVN2GXlER9gaGoEr696fcx9hVB
RZEX0nYsohCqPjmqT7O0Qj0eqVSThT1Ps17wNtZ7bMAY2emJx4HwVesaWUB6ilmIBVVQQCT3d3vv
ii3O9uMnAsjHNx7aGMZq7AHsEoZHGhVnYuWmBO80wyMgqthRrex/rtOFqLBsiomlWRaZjLISFyYv
S5IaeMkxcOmWV/fV/erXPXhBw0nERhByifulVcc+pdoGaJdm2HDw14pj1bCNmBuFgZuCg3w5VIck
cygPJ+b2YRmIi2by1ea/NwDAQhsK/AWbHnOIOaIkrPFm0vvGXaH6/VOzOuCUxIhSlhtpB10LybbW
Pmq78ffOlQhQjNVG9i1/ap8S3nCaZcvDILJxEkde3HPWEXV8Ctxz6EzNf6DN1g4Ei8poZ3eEDGnG
h8VxR5882XoGxxPGRc9EE47805zkTFJclxH1aBZzaU/A8c/pBkBw8edJnil5lyyPF74PwNPkcIVK
hi0I5I5TYiqFCizZFJt0bVY/zpz5TqF+utRASPf2rCnZdneR2W9JjZSXgQHskFvjsCqSHI+tWXKy
a7EhSYT53ozVdWWNHKVWoA1YgJpmPKtO9KpAjahxRKTX1ZqCaslsr30UCZqLLwkECfYH6Q8G8i8S
IbSW+CxOgq8AEk7KBboNbRH/lIus+KN5YFDj8QhqjLEypGS3t4TNdHvu52m4nE6/iPfevqq1eZEq
nH4CDxeLBHUT1xdG4DBGJjubMGMpg2pcqKpwrl/LpjNebV+AuxYOVRt0SdRCQ82YviGWOlCaa+PV
nWdspvQs47KrDb9H/ieYGwc78ovlv8MN0gIozSZDDlXhX+8cimIJDB3vSELA8+q8EZrYStmk99E+
G96JLObn8iVEyBsskfbhXAIjOk72RHgSrW2bxM+eJYlLewrXl+nuUeEwulNG2E3lHuVwk8jVtrbr
cGN9BFY0fFWqqiBVU/nI2Ct7eMHiS0td2p0+JCmWuMKzz9XEHd7GpdmmqoI1uT7+P9wFae6oz97l
OCXYWD9QJD7u9iNVwi01j+pMBGpmwKLmPK6Aic9ohWZlMs6oYb5DQRUjaSjsv/CaQf8WmA71g7+2
sqOIK6MQf5BjxtiJm7IJYX6XmM22vqfl4A9quW/7VyWZh+uCV9E2pKtA6BBp//07ROuKgTGX8RAT
3y7acqKFt8epVCmtgld3LFllM9fE4C3yugiw4LfX2wdcHWQtZ33sKgZDQWmrnsqcLYSJ/ozqrXTl
AX60tmxQP+77yHZWYEFlitfSLeQkZqSEw8N4Fuh+56elyk062SOy2CFMiOlJ+xwnKJUuQ8QY4O8V
bHJasX1bV6q5l15W7Rqr78KsVXTnZ1ZduYTqWbnr+gPN/Mfocl5orIb++SIB2SW1gldkzeYEoOtj
WeiZ0ao1WbJkPapi8+EZZIJL7Y0/VfhDOeYqup7gsziiPu3nB1fJM9fmTsdhmlwDEZ+fjlaKXGqp
HLm+/3ASBtIWr5Jpp5a2OkMqRHlLCii3MEWkeqTza+RErREqgSH05OXjQJVu/+3qvARDYLbgM3WG
GOxn2oC7QjlVMxjkse2vNYd0Vx5DD35lmYChDIt0gduHFHZKmsUdmQkqqMiIZyQZ2pjHPGiGZET1
AAkaVwHvpBmsBaZNUzqAmgsoOsVnhrFMGJc8070A4a3DXV4DCGZztWJasazLLqsQJH8gxI9iXg64
k4Ge/Q3pqD+geC/D8cJxRFwfjjEeF/dFNZgh80jBbZS/0gZYy7isC6QJ44xd8Dj8JwsAcAjog+FY
dCdb+Myo8wR87Q0VK5jAC4zY2xJ7fOFncQAGVXu4jXGjRin2606n0rEfgVv0YZQEX7fCO0sun+Hm
JmfA4AbF2+fURg0pMr47bsAvT1Zw0yihgbRfIEhdjl3srdZcYS4PXDN1IVeBTIC8BgnojlgmiBa1
jmEhdfWNe+fFanwibxQhA4miZc/DKWFnBVnAB5lpulQJXdZ8+6zgL6WgvqA3wmGRCEH09QZ6kVAy
lXl+gvdq59FeUh8gVcSP/5DD2l1jMVTuqiNxxmjk2colBLU+fHYDzKzvo0XuaZDw1+FhHnMf5Zfl
7EQyXxnf9dHQ2+veMtm6hgPCeUyrPoXxlSnZWGaejj/iCtDZaxr0f2e/JtUVGEV0M4a0URfyeXle
eQmrGydHY/zZXFBqZbeAgZ6OrdiJZaLwGXSMOnM1H91Ve6ypt0VwFOo3LmuY7uPJhVtuHIC1yRZu
+RSrPDyLQc7EsTPMrfs/4J54wbNymyvAUpX96m9vrWWRSkT7WTB4KWQM/icNwM89rvCeib6FpE0Q
YDnNPTOhO3/7+sNql/6bLAYVmTaubhlxvmdsmEVHbsqpLwmBldPL4QM2MEOPSqDLxXcRkmZRQ/Qj
VwuKDLVl44kgltM/vp4a2EgXpwbG1RJql5/J0cqtdUIgmeL/PQG9mWwjVCZmizHruEx6t9tG6jVG
4RDqyMpuT/ls6qj0V1wwAixPgdTnSRxYPQUiAPmJ5mmgD8ec8UgFaAA6ZL80YIBnYJassvbDLAMC
GFfdYr6/5LC4rb+NcZip+k7efXA5G0zknXTer59SFyU9rATrJ/7sMoMiR80uZO4Zr2ml0kQVS/de
FySNAm++IGA+cPZ3QdrDUEoL9jzsUTwQ5nA/vkGbGBB7SFLkHDdiZUSbOkHBN8mn0DOThV7BXT/b
Kly+Ypsht2/1wuJXoXE/INqsLfN06YSfnVBd6Yzy96RS1MVGEKPN+RC3t5xX6pLg4wRzKJgRvc/C
zs7Ik9T/qIl3/9X7GSsM2+gRj4r5tkQju0p6j1gx9R1x67vZs0glK37NQQDBGSyR4IezyipPjjH1
S+dnMmjEZ/KaeKXLZqe08vRf3pmIDEed9auly8fmHEI/oNCYBmnoGLtGTvIsfQPisKctY9Bh2aSx
KE+intRWw7TJA24oF1rrNE7KAEndfkPAitZxPfnEWFYei9sTmRnIogZfIAkPiVws837MF1c+idUX
28HCrl4khxCy566e8IegkOrjhxlKAAcUntH7DIh8N59kIbk7iMiZGjJfQeCyUbVMb/tftKMJV9n3
1nSkwsdxw5k0bUrioNKudfsmLH6rCzXhZ8CjQgoc9WryRnBVcKbNTlytSIYZoFUIRHBH+UwvbisK
E9bgywTrNPPylPspV/f+8UIp3DFCXi6Bjbusw9w3vSu0nNkJEb9Tq4f5pK/ivOBRfekcAtOCeOnL
kJgVh831fwovDZgGwnQ1eVPL8P7Q6vtE8l1TEFVhdCTo5Qhd/KRe/7THQ1Z5YB3i0HlaHVzZvD8f
C8fh4qGeeOmX6qg9X/aeX9sdoPpIQfSiDnOUrDDb2keCpeU+F9m8bvVE1mtcxem1VBU8ltu6GdL0
t86RL0u4Hn9oGCtr2pTECazSfiXwIe+7l/pbRS9SsoCQVfn9frhW0haNHIqrPUzc1pwPezYG/F3e
jGHCIYmMYwWXG9jEwYveQNsNwSbgjuyFq5Z+m0CjtfCqVPkCWZyyAx6gs4Mj8URCthsr2V/eX8Lj
34L0b7F6FRzrTNYdaVW8a+RxJ8J9JePi1XOnKC9mzwQDpXxDceUuEwyz5GQVZDFfUA/BRtkwftdC
OxnVcEH/twPKTDAJZDCvLqIniWrko94GlCNmTHoEId/USh1hpkQflsDSvoaIB5G8Mz9j/pMHUiue
dcAhW1krapRbz1LupsCoJMEZOVf7z0wBCobOtv2GTkWOZaqbpceFyEjEKCigH/PK4gSxZLd2wfoN
rBtUU2+IE8nG2JBxoaWKKJBWq6ec5LIuHgcBB1yUCaTanFwPxVQiL/hq4SsM2wfFy3ISnuN+hled
o+sVvsQuLzU6GKoK5U3jSuP+V5vii+JtogEksr5iQN0fP1g9avq5mFHWLjvUWzfYdlQVmY7otDbG
5bGmePNtQ/lxut3dgBfnSfSB0VFCRpwuMWJZvEOR1170SEuxvmjrsX0qJmBuspWhXEUHVphPQRXC
fadrJiw9GLPzrfEx3+Q6jaDCbA1I8N310A3HpSq8GswPvys7D5z2htkiTcbDJSdcduHxE79Uycqr
HlHneIeCeaDFsfD2ekb+xG1pgIp/nZsurWkZ1Oq7ecD9kLLya0QjKX4SjXdVuu0W9fTLBJrAL5FZ
ymrEi4WXpvaVjKLCH8MFFryzky1fhT7gMChJ+EkO+woeTwd12cx73R7CkznyeWKxk/mim39+bIh5
YIzlzcJkZvb1VmaF0rT1LnLfl90yf2bJyP/N6cWFSe1FS76p9S6JJzWD9tGvcrCD4RSdYxhpaEJ6
sSl5g7ov5YG0hc7jF8/hpDXgjrKJSN2j1ibJ0e24hDc/qfXa6X/RfnRQd/nL9y4g/pV6hkjolpXu
zL8fEQHub8hoPG3jJtn97gZ8dpnwwJmS5cr546tT1KIy5OZnWPpfQQLpoiWiqxCmU34b9GTzIMWK
uMcEIi0a5YDSdDPlv6R7PLDbLe6nbumisU2ia6v2v34waLyTyyFP4cvVVCXq9AEXp72bnoGy85zp
XtbnHhvwjRfhkPiYMb8VPQJHUT0s0lZdIuYmObpD4P031GiTEgnk83AoDnz5YFyfsIUB9PtwvOyT
j4T2pBx9bfnI2p2ucwLtdw53rcsutx+XzH5sJ8VeR6Anhm2/gzBZ2uFpDsqPdRWI2KvV0OGnjPy5
LRpw3jJh8P6z31OXB3XnYTvtZ5FfCEAMt1UwXE4LQKMTh6Ziqq8bCAf2WQfRNKeYU/EUuHv54fQG
qcioZmVhc4IrAW6Yb220+fJyJABWZTPxA9wwBeRYppWVmyl+zkpmyDqKYQ1iq+WyOcdQNd4vgHX9
71tNjoTmay41RHAaTKTHoI19lvalvQ7RU6bSA9DelNmhJRkt73yJdzcB+qyNiKN8aIo3uSwyG0An
RqbQdhCDGS6pmZGDl2SKw/1atk2MKMDOrYRpxwFFC78YtdhjAdJYHBmgbXciRNeTkUvGjIuLCed7
e4Lo9shm3a83J+dF42Lp8EbQvsAK5xahkMpCgL66WLB46dHeym8wtKS9nhm0rcscbzpm5nzRjcci
JxRv1rQPSqpyYUTzT/OSxkmm5BoJe7GcIjutcQM69MCyKl9U/eY364rcn1ndF0wi9p37VTQxtwa2
/D1vtrarKphfedxsRw6XxhqvnaqkFVbRLXdVlKLUa2CZHLlkaQCjdKEC6btVbZ+ZxiRsIxWYCCA1
7OSqDZpeIw3YG+97F2BpalVc9JS9Z+pJHMpFbAmznymZKyISKUA/NceOjofVIzkVLYy4FJoyFQ7s
gzBf7UaSQU801IacXlJufO5x6nThmrYJduUz7IEzZJ6SI1Ezm3SgXBjzaTq5oUCUVQMiqTh8pQam
HDIRWKFepXWJsbeumC3+yaLY6QFXt9Md0c/VFtCkG4PZ0Ixqpx52K0h9uGD5R3pWBoM3HmIaNhyT
QAaCfFH3TeVLiEC94LKiGcy+GkwOmMQsmN/bIJgrNYWx8+MMzfYrACFeDARXA8TsMhFCm0IvNpmB
BxyRu0h3nyrdUHPHj49MtkXt5D9mELZ9d7tBq14PcR11y32u+G3DVnbfTWDBC6/Ar1L5XtR43CmE
sH/AZ5XybZHUCdF300Al8dziOMlBdxJcfd7g3S4+hyl/eJQ4N2xMpjV+3LZYNmJj/77+iePA4pF5
sHMeamM4hUnz0Wk/o2cS4Z1NPv+VUdF7hJwKC7V63+ztd/GrCoirOy09vqDkdhPm0Wz1qKbh/RGo
SME/UnHku6hP9d83bn7x1MZQ2zdkPEWcFT+W+Ot53IcTYw+xmBk/gpq5f+iaTY06uh2lE40cvCXc
VGUo5tkSdv4v/Fx8SXRJCqudJzNATb/q9PxNSP/2VYuFNPI9UPrRnvHRP222xnSXiaQOxTUDLoLB
gucaZqzIprcVNDLVvCbTm4/5W8aIsoTWC9/I8eVU93t56oeuXaKtGexRpSeMILeOSM2lqEklyzaW
A1zbvboN1cEANROxqXhbj5davi87cyiTqSNj2AAUZ1VJxHgyPN+b6EzKtsGuuhjTc6J0PltS+rvV
hNizzPpDKngbkZAvevGWmAkeFeph/hTkJ+2upA6OkCnK9z1GSJtSMrXp9A+8O28jjKH2Cuf5fVog
K+ZSA7fysZRnrLrBWUgHHbfe2pHTqE3QWM+OCadNFuDfRfzBeysJgjQGzUsVt2gJz7RR8k8mUMIA
vMLMLFkmfRFETzRAu6dCHlYAIvNcKQgri1KeI2evbCp7pXxFmXAsqarS1Om+IRaBHiEkqQmrqwRz
h16cnzNxmTJQ8F/2qcC1tUeEfCfrZP4W9v+0aVpQe6SUrZErWIbXXDt4HLM4NAkZPyJAnjgv1nvv
LnlK36mSLqcWbHEB9JTcwUHv56eUOMpwdiGMO+IDprIgcdzmAIZYl/FufbaIm18F7Vfm8MAiwDEP
sDXqbxz2U6VsQuNoBpUIfD892140QkN95lhCga8+QwVkGq9NtY6/a5hiNNak61GiLjor4UWyzJAO
mXAjxWgSBPczJKoOr/MMZcniXmHI4bfeRgM5alvIcJcSdJg3S/pn+yTP3WBB31GxKa6k6CxkCSOl
TPaNggRARTz+4h43ofLL/2NvFcLzGBC6v4t84b6iiq2/QN8weInp3R0ERlDBFjMYVImBYpyJi7re
pHjX9fcAhDL5wWuCnGu8ayRjIJMSvPFkpAgDLebXnJ4uMFBY8/8HAbQDXVfNpAewihVXIH9PWwXO
Y3+qCeMTAA2oOVdIjANOtJA8mjGySFwxwDzzanXhkE9uo1SUJUjA6gnmSpne1nlZBEV3/HIzsMoV
cncAKZHDJ+VZVxDc6RRXuZIizBPYES97rShm3Hq0EFn+5ZZ1ylrVhzbubszL/ucjFEzadqvZxo31
a8mtjurkMiZZQh19djwrex4DOtXYayH8+SLPmsZ2FmoVchX7QntCrUlhT1XQjHREXeTUDZ5zv7D9
hlT5lQAlHCkQU/fS0qu3hApoX40QgHMFucX6dXtAZiDvpyzepI+lVOHFyTXdEcoOUGkfGvTmUv5u
3eAE/kr9uRdLfOSJ9nLaYQp+9Z/ffjt+3d2JLK7Ucp8T31QMllR4kNYenUG06iiLb2j7S4XVlH1Q
1GdFHwhgNakLy62w14C8VhBY6N29CxwHFji7Cx/iK4MwIoyyDWoDh7V0VYxTgtpyzc0dfNziTrpd
eQb1BkOUt9MWUVcmLwUmfpytiDAhKsl8E2ubP4LYUq3eI5RrRE4spwunmWRpN2oyB68GFzKOPcOt
phg7EHpaDERb71rAY28FHIQjRsotwz+29tQtcOOuEb2y2b6h3gevOQRLpHJp4Qs/Qx0yXTITAcu5
fBcY7QJihDrpsvNZO/Duwb6SWGo5GSt2HL9EWdRb0Lwauer4FNMmvqOeaPeUYf5gAo0YOtQss3oz
a7n5kMHrINWn3hI01GROcrU5QIgROPMrhqKKbILKPBy2N4I6YvmS4+MRPmsuAdpkuSWHS4tvYj7c
z2Gx6qW64FWsazi9cirT4KbwAGpPCYarIBjWTqsosEb9Gg92czmafSLVdPKmUR81r5h1QAyHSflb
1MCAPNA2+UzfAI/f3RBhWe1hXd0h18ZYCIjr8+5QKooN0beFGv5XJHfJ72Fx+G2tauQB0TDOI67e
U4D2vCNYdjy1ivx6pUGBes0AbJQTjMUBs8qDxU0GrOA3KrFpyKOQCQgr2muFWdhhdHT5CusKH9l3
Y1Kbz+0IiSEP8EudkiZLmfl5iEt+3/m6T5ezgSO5fPzlXVbiZlvS/a93uhAOnSHwFWxNmTxxD30l
bVh+zsYvhkv/WFAV0HFpGraOHrnIEc1ArWs1RU2K72f2WmW2ynZKJS0KKgnhEV1rZ/AzQxSV0D7l
MsSrpQXiay2B3uGwtNbHUb+uda6T43iilgmxYIJNqkngNB53L/vJiQG5t+Q//VUYAAoKhQst9Bqx
Zoy5tLldMH7IFrXbxw+Cs3WlDtt4/mBARjpGOAPRYK0SDHiwWAay3ChwgUNRHRiDzGnh3nHs0R4S
xeYHyZsRaT0+ISiu+Bv6f4hpB1iMw0yfP27vcNI2jOudI65SqnbsqtQoW2bY6aPE1gBWRVBTSuoj
8N1kuoUd2W341fiC+r5w9FrC0ucJ6An+yXpH9ddebx/penh7ggrUr3W+rn8ofVHzwHCe1IoMMAPU
qAX7jRiZG2QXUW7NG5yoFzfxNkmHB8lm6mHUayLu41ft1uJudEIBIbxjy2v3HMXQ9otasmONIEDe
IErNHPGiPJSTs1m3NoNgIjXdfWU9c4uVlyR2acRYNUbWiD1id8QDPOvU3yifg1uPVbTgNtULkoAr
ShlIb0C5Dck+29rRyXxqT6N9ipodFtoq1R88egmOLXoebAj1HurVQzpYzsogHDoeCCFxfrqOge9m
wcWaE1G2JQQnlQBIVcOtBaysi4AJz8PEW7toLq63FB49V55SNUwDLYQBnxuiNsGugCZGMEhEEa8h
1+WMp5Hit/R1q5cfcNGFmM9r5Y+6t8THMEyC4o9N+m1GweX2NkDfPBJ71x1SPtj21VHGc8om0vSH
t73+U0hboZWPVSAT+IkbrITs2mYgRMX+Nyzv/+ZwQcsvRZfKf7n9v0b8AHlQ6R8XgoTg4kxNZb+1
B5LpOx0+A5Tkk+Xn6EH0HFuLg/IHAeGHv4et2XSrsXPSjDLNmPWTK2Dy398QN/ucGxGPWdFnccOk
3ZnXdMktBac3RxYyXqqsUBtA5sJXYWxRqZdUHch0iH8/PoBXDeiM91UZEoXr9+ESnD3gNlrkQ2BY
P3jlr6Pcib/5AQguuyvApAqdyU0AjhXjmbGYC0x8TydurPBqZek12x4BnuX9BmB4uImWIpOHg16k
w8inN6eTuwwLm5c/M57wbcSBDP1IlCYcRAQAO6Yrh4Bot9x3WhR84JSgzszA0+Eeio96rVgd3BBq
XkIXVUPN3KY0n4DHShcxF4DUgAGWzNtddV+pCD9VWdYCsQVt8fhsAelvej0vSWKFO1BgMGsuFBh+
hs676i9RN0EUxQhN6d4pqGptGrIljyxKpFYF8ejwKrDqhNAomYIdcjdrLWYVXKv4Vuu+U824JspV
Mu5n9ZqSpBmwKJSc8Pb6IG6Pyu99ClZHBoeYDK2SbCi2mYNB20/om/acf5XEOU9Rdfk2clZs1nM8
KuJPGBRY5zdCjXiisLEKwpV1halqmzb812ewmsUW1X+cmhtgWuBvsbXV1cLNr05QK7d6cQ+yxNk7
TjZYW1VOHMaKZgN42M5PYsnAmtfR4oFRjJO1dGgXBBPhEQ0RSoKSehHBhoRegU5CsF9E8Z2jHCqs
YWPlE3e3vZGVN92p9K8Les+obbMZ4d4aLyFdR8SEkTduWamGhEmCqqlXNpaNurG/q2c6FFvsxYDt
q+GzDevf2JChPTaEJ0pyC8QbjGgeOOnCZnPeelrIduXtOfI3LweFJGfBcFiLm78UYw9h2b6pWptA
YNMh5BU39tbgBZTBygfkg76etQkeHMNAXZ9yPMoWmorqKODb4kTt1upwMFtDKIY0UzVr8fSHilT8
hu3tj/UGYJpCgCSXwCTz3W74+u+jLWoectqhZTPM1Bde6jD9labD9EOKsMWTGbFjuDeJYbTe0+sB
1ufd0j/mk1tikQugjvhb3H5sGwePt667/EjRSakvFFihdVIIRKa2rDUw+05uPh1pN+4G2At5a/mo
n1nmMvR9igYYxlEy4s8uejBEplMUIG0KmpSgzMUNlDz+q1dZSmfAjbQ1DduEc+HHMcGIitMapj5w
mg0xw8r14Q5m64KFILoWELXRpewsc869qO9kSeGJ8lgLBn4eJa3GKML8avsWtTxZuMdm8QC/Swrd
Lz8l2XXAx/BbcDswO/Kou3HM9aDBolFT3Cb9PJ9thiDpGPOmYViYrEJlvr0SwVIHr/+eHNgos7Ju
qyySl3xEfOwiEVZ/8Tii2u1Svrvl9BBHCKT713nuxb7ENdKr2mc+fVL2ht3qLH4mjY+/ehi3XxHA
ntuDIaz5kDYg+xWh4SQkJwLFLQChAXIGeMoSd91Z9UgC/n9CvFA6fb3747/v6c2sV/jechu7llMq
wb+PsAEOl4eFVp2yKolayFVEvZA1P3YSPhuH/CsKxFymsklvxvZPZQlJPQdzEXVsGk5sYxgTZjwt
Nf9TFco/EjCU1Le/RlmUhRoes0HrKTig7u3VB+TWz9tTqBbATgDDnalNkOv1TJCmDSal4Aibbmr9
s9VyqJiT6W6oYEy66ktvJFi9uF8x3JZYuy4Xh54PkFJPmruDEZJoCLudBs1QofzOL+xb5tfg5yrT
I9t7qUjwJnqUM8H6BP7HRtRIFhbs5Gvwdv4eknrj5qMwUpuEbAxlkNeJpinXCALaocJVxMXhhhYB
DNNAeuFwyYaJAtZTvJ4cpE67CQb/AM4I7yfm9YzDvzhhVmBGh8/lfWUSvasQoQI86lq1BxkuOX2W
SnYtAAZyAOCKG6l+seR8GFLxSZFUKG0hPMce1VefV8F/4aPrviI1CdMwavp7t3zBa2i07GVOinTa
HRwx3O6PA4gb2hFgfUmMaLnEcVpO6Zoo1TmWx0umS9i9Ny0jccxmyyenNXSAbn2rk3VAv4xlhXjH
myAHkfauoCkGS//SwN0rBM6djgLPFTC2JDUQ9FvMPtywOt4ZXB2up83Bwo1GnFfHfaA6bj6dxhYU
BwdkVPLOJfs8ciDd4ACSQ7Mjd8bIkf3rL7KNmbQvfgKofpO4ka15nrtX5OF3/gAbHQEmf3dn6u45
AXN3tHImdixtRDRNlGOoPZjNAUFQwQgNj14KHnoZblUdPhH9PQv72l8I8SRa4dnwQT4UmsYbkBof
DJGesB3VQ7wicYrkgIP0qi747RwheQEbzzvQ8REVv+J3GxjgYgSJsxsZ4PRAdKInIVdyqkJ/Vj5U
JZAdZ5Bs/uxMoYpEufYbS4APrguHylSrLR/quL6XPMJ2MK6G3h95hnmYBImThTKJsmJ9k4ClZyaB
hp8fEndGGDVDc4QlRvhg7sSHspJ8uPV/mkuz5jcnf0/o/XG7Jy03ruMso+U23xfJ0oacFkCQKCom
+VYVhb/Y2pydxnaLIx3yVuoTM9ZHR9P/fwTqkERW6OtwPKRCRB8GrmwI6Sre4X7LDBvcoUkRPQNb
aAXHpPSr/zqTomcNYNIu8s/4MeRReBhtUGjjntflzfb/vBMCNXB/RDfvyY2HJVlIJUckV3KGf2lN
YEZbD1KT4W6QDS+pShwJdyqy3+i80pCWMroizBaIEpltdzE5IpTqiGod1WTe1RUPl0Yc2s8PJzrn
hoIwdqfW5ZjzP927ryjl7eUKb54U3k1XoGB78sznSOVxZRquoTi0UjOJNuOlQF15n4rJjlevKik+
QV9pzvo/A7+R8mG3uUaFN2cZIUuEeQE3Ic8HGoo29geiwUSDIyN0wOqrOzlEPjcvuWQsAaWFOrYt
JRZPvJTgnDvklDMaKppS4T+CAVxXqA8Pf01SGkDo29hcS1ceB9Pr0xamtPUjG/VqZtda7fkaxVl7
gMvmJlfbwGcRZ4oLstJH/8+u+4twZd8Cj9rCnAvyn1QObS6j/bWhYBcLq5gw4tSdIGBGHArQ7Wmc
63yo3SIfOUQNbZdhCWOxsH9M5AYCsBAuoWpAmpxUABkIb9Un7WShehuJyBfJRgjiwevrSK0voBx0
b3F3UwvFuAhcYZnJozTxePSivk2jdPPAbT6qZjRdsjjillzEGVmRzB3Owiw+itdu+aGYBiTBY1OI
GorQLhZ3UcovmtKTnapPG4mGGTWVcNbeXCZ1ggQlGTbAGAwLhqifM4lCvaM9BY2iXLp81/ZbZeqf
DzYkvgyXzEDrPgRUnqM77NnWWzIYMqkA4IJ/tIa4sHWc0pqSSWpmrczwjorbbAPfaLBLxwXnAHes
0MvT6rgDct0FyjKotl2dSOuCtP0kxc4vCJqYEFCYfGbzfV7MdUokFeYfSkwccbUr6uHt1uGKpiNI
RUmmEauRoi7kJOe++mVbD6DvhEkxvJNW5bsW+p+q7Z5T8KnBeJLDkaZzDBDr1uV4VsK+vlH2y+ow
bBzS4v4yqLt3vZNJ8ZfoE7Xb9jGU6X7T2xhci44gZ2FkOI/lR6jYFRR+1RGGxTGwgpCamBzlvIXM
qYoUhs6f3wfL+7WySZvmEE/fbtO5CEI7VKT4CTXojFRzZwUiyKRHe3RomWmMagwiYzmYQ2BD7zQ/
pOoK9GaBPvF/ArMU3+IeMk7LFl7fJWGUXMyXP1Vol6fyqQlHeNATwEsC1M4nJRA9zlA4nTPi54//
dj7ndI0LJkkwVS3ZyQZ9wGSYOCgzX9sMOy+NJot18YxkweU0Fc4EX1rt+ulvSQx/uBLhbOb+xzPe
ZXqxKYBsv058XyHftW5WefSvGI7v7qFGOx4LPr0Ykgohax9UoWKlCNZAFz9Jvxab6272JC3jAneG
6E/nRYNKKakDh+l6DXBiV8tZ3LBOmTaCBB/uA61XgNQFDxXEzZqEwn5htS7TUe2T/aQi8dNlPYAg
A33wjdwK1blSQUN7ne4JdYE/PDtqgHcMWWBOPXdSnDmMpHAR9Z3SJH5U5OOS/6uS2Imc1K0+QfGb
gu2B/6O68dX1nmDb6PbnyByy9tZOvJ3zCCbDKRGjeLuZ+vcgF6yaz/fbK6pwqpCLdT2h60fWdVbM
DzJwmiF9Evn4r/+0QVZRG0uxnvhELg7NR0kSo0Ol9Gl03QefizbOxJ1D1Rsuhmo4ProfcSwvkGzP
mN6MqunOxEQUe+5kZwrAWFlLD4gAIbE5DG1GyCFQCUAyXZKDMfm7SAWtJBAY4Zc6JApv7Bj2f0Q2
uoiunPzT8Ltw6DhbpSxqRpddbq2uHaOMB3GcEOq5fuymYjC65xTQ4axRONLKfl28Vp5Kpxnz5IeB
nMeKEFwQowpVe1YU+jpnFBSrLEo76Lyw0JUgU/tWSKR0nbab2UGbPyddKRCbmS9j4fSnqnAvvL45
tqDJ+vCUHDOv+OD2bnqjdsjp/QKB+vCnY+grnSd8DO0GrFhY3pwtYaUQsNMo813pVT7/pfisOmXn
pepc7g5r2p6UPo5o3jyx3UdtXimm2BdYsf6qCBxwvgEQanOpq8Hba0CZTrLK+bNOPlf8mFvKCiTU
IutiGGsPgYiCeHCcRvU7bW64pD5TNOwmezYfoYhCDqOm6efEjQA92/hCICsV+U+1CVyllApYDy6C
S3XatRb/rXpEe5VcxLaVJ8by/vSSsuEJ8CV8RAZQxcyTTY5FIo6jwm+8wTsPf9gv0YzwRX9QvXMP
ubBqKqGwYWL5Egt54NMzzJSTaE1E5hiXq22ErV8X5Wwwm6HEC9RHU4zyp5YFfI0FdmcaJHc+uX68
y+1GUmgogU1JAxM1CInpWXXCMyirEwTnoDbIC0gHwDYryQBdkRW9koWbkxIjz7SloaP5QyIsoySa
SZha0XyjeayFPDgMC+OlZ0giDQxzAzn58fgPD8bT2ZO8ycxkq8VLr+QSzf6N4dAWsRbUMmHXDk16
i0AblIQ24zh1dW24KjqCmrSMr/IoBbjnpt0YZaJNEZ93IWyf/2AzcY6sly5CagNIF3LEHEJgbhSW
jCxV/6TQQjTbkCpkSF10jCqSEpIrkwlrGgsM5u2B3FtewY+pfCht2qKWrS6o6A950LckOmJXv5wE
MS9GnuOQW7XA7fMtI1/MnxZnTfgki59LBGXlaouoB9XNJXmePIeMJUuUWbUbR4JMpifsEMF0EMtF
fpgx41WWku2EW7b520lMiMfAg9UVHSnWHtK4pHI1S0SRDk++UgGk10n4ytfZqZN27uwJMNdiVfsg
mrDRV4kh4L592x/Q+j1PoX6EhDPhzdUMCp6dk7pMa1HdrA7jZ8BW78eWaUaQrfa11HWLAR6nAKQX
TdPLJT/NpzlF0YMgYh4ilvDFApvCN/hlI4cngD8T61K8couIQmpnXPtkxS6uXiQRqr0RvEaKG84y
9UWoynU4RvmAxMfXhU86aLpt7mxx0yyEXmQT2o1fjggoXWACuJrhoZdKuV4cDtH9ZLeodOJLUK/e
m3egp09a/0JniziP95Wu/rR8L+BwZ6kl+8lDEW6PY46L3V4EFstHnVZLErai/SdepH1i6NpioRTD
+EennzwidJM9HbTE2FnRJQw+Z22sOgXHWEoMpGq3GB+qb5mbC3pqmFLXIK2mzZu6fGaQaR7Egk3p
UwJMbhUuMASRZVSRa0Ptyv/btw7VTVH0YHyHuJRrt450uqO72aTej5WAyDh1cce6ZXWobztdIyB0
Crx4AmYzofSy4pPPUPO2y57eqXEFXqBWFN23+Mffaz2gkplrG03sg+kBn6gZ6Hh2U6DVp3YJbLDI
HZXmQb8FvC4S/cvVrIfbcwfi93KMCH2anS8rZfi3hKoLMHj5i2t8RVESWVFZ51eF0yi3gglUetDB
SsV/st8OPM3ki5NcPG6DTLA8Knb2TIjPLxhbIkMxNLkJLFXe7g5jpay4yaHX3zMCpIEWp6dMnyjO
H9CikPf93whQQJbM+5YwNCjkHLPLtMMl/xGh2M8fmEzWLMg6tEVBL0sJxwXu+CECG5I1X8XqQBXo
kui2uA90vy0wFrwmZC7g0wT8kX9IpC1e75GiWZX3MJ6Su/Efsl/GXBMao2aU/c1ZIu4uYGmpkVNk
v1qAVMaGFnLf7v7nOw8zMFQaZ7SXSk7aoFUcMxxQaUFy7kJVemrRzEGVbScVt0P+6WDPOwoa34aB
Ww7ZSzW1y5eNGrVETxXB0QHXskg8tZnEu0pGZvb/fb+Xvb4lpQrj6D7l3DnYmD7nbbF6BBi4C6UB
xYRVXXc9gGSe6aGqNno2v8Vj29buGPVkVnoOPPtztKNbYonPkcsoblmJCxFzvble/xgmhfl4XQVs
HpcEQagT5bSqwyfrz+obhrVUnkqGTimCFFhRbMalrHl/z2mxHU7FvVduzRH/RxdODl6Yye05hIiS
IaIbBPOcxSU6l0lHQYmlGADyJrrLCzRdeqwFsyRtuBBcLV2OrQiWrzQ/gFKB/y46jWPGMTByNISg
AS560GCNjZVGcsbk02vYypqU022Gm+8AQmfx+DiXRguWL/stHDeDB/YxVb4iG02kvHynyPX7fAdf
zL1b12PfzqML9YOnDHebKD6o2ZE1PZsvpn+Y3Our+2X8SR1fPAkmg5SiHOm47nI+QVBR3hy6uByG
S0Em6T39Ds3Py6otYXxvxQUtXZBgb9rRWZidK1OGpIE3TipE+nQaQoqBKBY8zvz81+t+PbkgimFD
zu6VF8foy5FL+/jAydnETNT2Ro20bN76IF/ImgSH5NkJhUYqW55Zxog2qcy1eoerdo8JWfTd/lne
S31jtELaupmaHAVvUVxU8eBchXXguB5GG5ofDUtzps5fcSigzi3Y452lR60zPloKe11PitCeB244
OC6UNezirseuyT8KmbGOT4Bk6h851B3QRZYBYmLBR63kv0xNr1hMKy50usjOqVVhgklMQ7//pgyt
lvOy31b21j9Ois6NJroSslnXf5GAwwL6Jkvyqx8noBZROwUIdpCv6YNkTgamoO/5rRszUeESRiJs
ekQfvY8EP6RAN48IDdy/L/yxXEqIE3DmJDdMrVyVDLMKioa5465erBsCcI8HBzCHSOwDfNj2NQxi
TF2DBhOMLu+Ix2AblhD9kQrsfG/aMqPdch8V5tLYnirdM3fMoC6Sil2tG4nqLOk/ZL206neEK29V
E5i9ie4LkxZ7Zz5rbssk98cNkHWetiHqy81QlbYfm/cbxf9LTByZYegkA2EwWo4LDYVK1myiFSYW
GPK8/up3YuiLbSSezLv02eBcHMXNuwdSBvVn1Dp4HgKck2lbJkW2e41MGaXpv37Q5KaeF4l6+Zzf
7RnUv0cgmaVKWOIbOApcLoKBDSBtA0mPuJwTHuJiDivAgLcJHAz2qPVgY3v/lnZrY11sehS3+ITj
L6xu04IYIvktd6zzE2e65+IuY3BUdET4NaVrPqsDrIahiOkebHuWVTV0kmk5HgW76xVHhadKe5L6
FtBimf88MTt5hIutuWgzM59Mco5yUYfk29eZda9WHihaa32moQilH1Q/5biqJArzlkYxhRZBj6iR
eberqpmUJta5AQruW0cEP64ZKHzRjNyUyUpje5YVRz0LmVdWZn0Q3xJSHnBZ0fAHwIJmwu0Pj2b2
7qrPMy4u7LoSMX7nvNKuXiPrHta7GZd9/K+hNW9wJWCEyd5fVZKGqxmvuAoRaTwR6UarVVVt8rR7
2OcLouhZwMlBjtLlBGd1EsRhk9JmP/8PlitmIf+/vEDwubCRGxNvj+1YVfseBhs9XupESjPTcRsQ
WPNOfPWcxq+XsUJF6qkHEfhvtUs5H6XK3w2k+UreNsW43nFlo+JlHpJGdrOpPzs76yHOR9g7rFEf
FL5mS94WtKzYtngytQVkF0479b2oe8nAeu63AIJorEdNpAE9ntMn809u13dwK/m8MnFPTe+SOTGJ
ua9oFfnBeVId082Cp8NW0z9JJZxPLTS1xKL2UVc8pkknUnVC72nLtEgb6b7+7hPNRpVVr2NPdEMY
O3l6Lc82A88Wce1u5c57vXq5HkukKyqKgHicTEhyty50cjKI2oam1Z9rxRYXEBG1zSMxGZp0IbuV
ipYZAp80wmv7CC2YMgEFvdnRK6IsrcInyEcu2Y8mr0fdlXuehw0vlo75tLU8Umxf2lRxChB+XNJk
4Ru2/fpINqj+fPBdk+I9dj1tqom2SWMSUIgvGp7X8Un3c5EBUE9zjDIx+eBE7LBmcxm2MgIX97JH
kKEeHsRhmku4QK3l+OgbcbyLzpeaT/tL84TT0apf7MU3lF+uGxTN1x1izN6tTYdmm5cCIhiG+lqf
fbpiRaXiz69gmEVh3nbfpfl/mC1HvHx9BYtsT6iKKgNOGPLJBfD6+IpL6Pfb9RjTiGPeM1L6ZOTn
qbcOyWMYgQyED/bTVOAlWEWg4ZWeCRekw3+zPFhiXEr+k3z/rEQwtgaYCM/vHF1+1ugm2EdSqe0m
PG7epjJu4v76eK5XGXYcOk6M/wTwgy2ynU6RUyge361v7ok2vH0Fs6VWVL6TDBAK3w3gLF+QPH1z
xdQ7wvBT0Y+11SOtWNrWccOjnbBp3jMWGXftPQJSHYWfsx0y12RAdDP846tmZSuqsb8x236+AY9t
oLsriojqRtIya00xGP1c+lfwW4w063e6fzpaifsVLEUdwYeok9UWXi1L31GSh0aiESKwhjtqnnSE
S1EawANj3KgIMsQA7g0sdC7z8Q8zaguIU7bZ2f7wz6/3W/LBYTSTygTWld2IlprWVK/6y5LITr9p
AfHyDst3F2sO20cbEnaZvrDFoxpF1gfcEcHioX0/zMpCLvNeKbO7OisYsJcJA15s44ALnqlEQXLa
MXmO153i5vyre6KuHNgUj5c1dc7OwQmUCq0e8FuvikprNBr65o9lltPw4OVpcUNxRfDrRvt8a/bi
j9fzemLFSZzqE+u3hZ4MkI4b8MHUMsAhuuKP1VAJa7KrhOyTP0Qa3so+v38n7mlxACPpcx1jjURm
BaqgnVyVcnIxaV7ego3LjZ1GlBOhihlBE9QAYPfyohBcJrr151XZp8/FXxIfrC5l2B49YIZIYb3D
P86txO2LorL7/pNNQe+JFjXR2tluQ4HF+4/Zyd6l4s/xFFPYHYNQqaB2EG9X/lfLfMch0+9hXxkJ
lE1Aps6OVXVM8TD8UUAlB8x8CHFnX6B928S4SfMnu/OdvGmV/bEB6d7+JahEuJUaZs+jJecxPoqA
eeFqfzg7ZXEFh3ANsh6onBId0OjWaWDtqeQAnjrNuSEqL8bXpvNcZiAE/1iOlVDrSJZAtf0FyrMk
vImCmqzHVEOmkGH6WoPxXz3TgsROSbG26Npc3pGjBUnW0x8k17kjAl0n/y/rKuVCfViAhU/liHie
36uzxUf7B8DEAMKKlQoKCVDJfNk3tJT5olsOOdu/nKDZBERyyuYgGqw88q40fz4cT0XhK2wLMLUa
ty1UJPAIsVlR+bxFYPlPsnCgadQLuYvGODT6lXH4LMqXVOrXZIamxyJE3ESXHWFd9OpNQM/0PJ0G
sOxs28bkJ/KuWe0dAL1ExEE4oHmNjL508iUfC+tWYKF0ht1ESfJRyEi4RDd436bVFXxIQy7CrMs3
z/U7NyO2vH4c/nZdqRczYtwBoHGxKV4J9S804Vdg7UnVL2P4sAjgWmioc9dhY9UCdzu8+gfoCJd4
CRyXYTKhssmIBTsLHUglGwZqFAl8aUfQXBwLpAWkrQbwArt4j7AeT1EJI10/l3L0geSXlmwmZsM/
ZKLiMaHmaeRYQq9mgn/PmBEiIKJvAbOH1qHR/ObF3uJ7LcmImRW95EWPJEOjOwaqLpT2GEXZAxoF
jqFfXHC45L/HiITIn3+5XG7/mp0mtfT3vlo2AloMkVJ8hJY4FFBYTfojYTrqaAxUqB7nbqRzMJbk
6vCdTm7UyGl6TV+MYxdBV0DOjyyyrW7/lrjD0trgLWFOzzQw7fSrUdZihZRqFOnKHtvzSxMrFQBP
Q6N+aOmictUgvwM2dkizeDaJPA0jQFO9HF+MFxSJbg96G/EkeVIV08HLxv9yXxb+L2iob9/XFd17
eDQwPtS64Q6zA3yyVzcWAjXBw8hq9LrHc/To4gdrGoOmup/QHxXkVvfB9C+zhJ34sa7CBuGwUOey
crVHYykCUT4UNE5JKSw+0rpEc25ni+K3iWuRBm23zQbmVCaA6N2iC135Au5pmgdtfRu8IEz7A8uA
y7Vy3gJFwDACOSB20ObxLknqlY2SJHtQs1hzZ8gQ8cr0We1MjjxGwcT4R7851rlBUe6YKrv6AQjh
mKDkZiiIY0i4gF0o/lnO5+fV35VArdXTaJ7enVKkNphhdCjHIXcgkEgfC/zZqwNIX9Fy7Zx8rGCj
N192kcRaveWX6C/R1vwAc1pj+OeKkeUoC8x8u0hbyBpjo50apBnCxtviIG0ExafBIP8SMElxQnSR
2HhzCg2DpPjgwTrQt6Aep4US21dKQhysB8CBQShx03w4TvOz1Vm9tIHT8sB50L6VRBsgr2Xq/KQ0
Aa1Hj+/pOPA8lSELO+T4bAodNE4OLvaRVmxqQ6n0jYbPGRcBPbbKPGgjjjCTydIhdtRBkwh1TmG2
9iLfXJTL99nI6Tfy93knUlM3yKe0mwDwo3wq+DsNy6/LlD/Z5aKj+YAiK4Yb6qVXqkSnPMXI/Fuu
FMc0GRjxuqKTYtsmZjSOIPJm5Y5CrExIbfCtHLPh+HLktsdHVKo8NN89OJm822oRu7dLDKRckm0/
FUYxCxSuYc7iD92UMwRA7zIUTgvJm6uT+MXV2bt9Sa4DADcaUnSdHjmJlNCZtgIrqjd85Oz5u5tP
wThipKbVXuupCY9mwEwqzEgzgaeJ2xuERGUb1HFqE4GDdew1LzTAszZbcwpU/Ld1W+VtmITUrIzh
n/tvm0OoV7nFYq7SMOe6dMnSckYP83vdgUHc9AG4V8naV7FtYNsrFMqK0TZ86Vfv64IJ1TDERAC/
eznbo/KDs6gypLBTnA+gRz/z7n0TS0PyE7P0Vv+FnKAJAQHxayAxNaM74gWxKzYlr+pgd1shR5g3
yjV5fVJdOCIlVK60DitiBbtdaIFKR6/mthKp/28wzEyBHe+wNcctAle1B/aVSLyPqb1gTfiAIQtG
S6qQbz07a5x8p4f0ndLY/EpAEcXTTlUki2W0yjRUT5VLf/wCGAYTyBHVlLZmieom67U9HgqaFIwp
yHIg+Rmh1FCUvw4xLUaAUgmdYbOwss30fs7NdqeBMxzywW2pz3p37S6qBG65xhyduryGfdw0wqlp
U0UVjoeO+GesbebbCo75zn0W2VHtijYJISaPBeip9cIPyL4bIGlOdL/JWBDcFt4RQBq6NKYTCVvn
abQX7UwWBKCr7z0GnzL6EdiDhnx7MWHH6CYBZzqdlIg3WPiWxcqnCp340LMnIq3bKk9lYI7SOm+V
yZPBftad7s5RpAmFrHH+BS3s2kGYwZlaarIWreuA1L0nLozimxjbJGlD7q+EzMdAkdqwaUXWQFK+
83nwV0ZKYpkYU2EXMzntOUxnQF/rJRLAl8XEcLAgG59+9U3qmDDLdhCdvdpYTg/QDobmkhI3Stow
qOmuGPggNtV4e3id6iqC7O8umaeddyx7AF+NbTZw61ibC/zhF6dtuWBUdhXUpIwGmwFB4NiJZZxQ
QpTLv2ltaeFhOglXkzUgho7pYOYm8qXxH7+A3+kWesm9QRXpvckRcWUlKZqLjnJBKrLkurr3FuJD
klsNQq5p5Sb5UJYSUbmkijUb5AH8psuVXjn7zH5gCbapvotsIUyV2Uj93OuDJDPYjIwCeBJj5YCB
aIsHXjGkbd5AAH+/iUoHKfBdnL56uku3j0ukMbJyoJ+0IxiFE7Se7Y3EH60J3nSa/ME0yexZ9vNW
9WEAyIRoZsFr7A1hQb0T5yJfBqZ52EUdgYqra0eDiG7XT83jSChTRBJXw/QHpmbMrYgNsYNSsd1t
FMomnYRCroX+78CHaT1+5JQ3TVzZ+SmH24ITnLuff2x6OOa2PQE3W1HpJ0kC9Uznd5vOCgcS1iFY
TcGszL9b8QmaZFZckmpM/ZdX7wJjw/juUIA19o7mvcxRPHzxXJx3yJ/tKBuM2rq5h8yW63H2mk9x
zNSNeRF1lnqG67lfCNa7HIIrQ/qIFVPo9Kv6JiZQTf172fEcTRFjjcf3Pi4aL+Pdmgqy9SPZusq5
bo9B3ClwqgV6mNSoe4BmJUr9YROs7j1bhg7nUYh6AuBML7cPufOeHz2RHWSLxxjfYm+N/ST8SNQA
gEDCKRt2b0ntpQX2Q05nTaH8kr/KZ7j/1TVzmeh30widRWa9ZFgXjB6EAIEChNDCPOF0NCHvo//j
5bPZr2Ce4r/XjXNhveo4PASFZFdJ8Gu3RnlZUvrskWTCvfSYBASniFLeBYsWpaQVTnnwQShi8/+m
lnYas9IJtl90nY84JileZJ11HWN5PvH4eLdOMxJdrZe9Rpgs+qYYaxj26DJ+FCHBdbW9P1eOebJC
3PCyp/R81x3yKEd/m7m6jdKPBQIJ4LDiw64vc1vsSze3aujfzJIi63v+9Z/a4PYNqv1avB8ikSKb
rsyn0vkjq+hLoGYqS4Xs1ONmwik52yKyVp2XIUdnhv3ACWzMEx0KU2NzUsqcdmqSmsbab5Un5LRd
A8/SNsJ4Z75cBQJyJ0A20ydzw+AVJK7+x2XwlQ08wBq1Nhafr1vNrBAMVE8N2tVbAW3AK7yghege
lEBrlOhBG5O1XXLGfdXYySQCpmLOTSF5InpkqTNqRyTeRFJw+FSSs3xIo+8mzixoWkHlxLJKx1J+
Cj5hmNG4WEsM7Bz5ASfbijlyHDIDTNi3HId/9hz4bic3KfH6G6d7tPrEfcOQmCZT2/wViHXd7UyG
vLjS+CYm7VSL2ulY76iOgv5SYu7mypT+p7TTEy6rUZ+wD2c1vmcJMokaJSubMd0PGluKjfHlcq6I
VED06R/oLI8Jlfo4gIEuc3GAQZmhVi+G+DBh//Fo6ZrTSytNWtRh/UIuHFw2M956yEVtiqEgqiGI
OVJq5oxRNw87R6PAT4UngQkGn8xZ4YxSTo3zh4pHd8gd3QMRo/svz1RBsQS6pycQf88zfWgQb4wk
4CLXONF6xhOMK/KINdJLdb0Wzajbfb41nFKcf4P8mTJXnkmC3IvZH4QTnlZMzfhyNxKHThAgKjdz
c8cUH2OiLldwAHYPAwXj8120STOT9iX6qehM+3usRBwF0bnnrylsZI9q0d5cjKZE0LtOH5MFrJMH
7bHjT2xsgk8uSKq2a+AZoSLvyfVzPxHh0vkCkxRO8kBXnqk4GzFKKNNbcCHt4trUxeCR8teezTma
uLvjjLGm9FYqaqEBYJ59ENnf7MFnLWmzulnpN3lKcKx6Nkv/6a/V/4JoI9Iubca9QvGu5bJzS24h
nl3wh4CqnBq8qj+hJj9hbvQ90/3zVCr+W0OuoAYae962PCeamoFbL6fR+wAgJfWPBrif7Q7SiEEI
O+fBLH60C5QXcdt5jPbJS8Qd0ouD/yLT5VJ6oJ+wYEeSKk7lfZLWXjjbcQXxRHKEi8SAUnCD0UrG
bbzoFec6x2EHY0FB4cZq2Si3Kv6F1vs8pq5D+f4KsKZQSghnnQ1Eahi+aNSd9z3q6QNuwEKD/vtr
iJUCGAL9rBmQAg7sbg2t5tjE3Pxu4HTssVg2mj1L6Ym67wTMJ1SauqWC6Ul3k1aZiWGZYN9jvyUn
NGv2VRe97z1Tx+bA0zsU2PCVZr/DEFJ5o8ulaUaQEJK7+Eh4kXiqOiDqx4R5Uw79I0kjouPtiwsJ
P43+zZynp6vyW3fZtw5/d8YV5NVMgNOsZNGMCIgOrE7y2aZWh2ozd+CM5QGhcYwyQYNX2/L6TnPX
tlpq7MGkCzCFmRj4EmKtRGfLvf2y5UzDVU22DLG9ypvkxjTcr0X8Ozgow+GQzB/AgbwcF5DATpL7
w1lRAYu3IhfVVQDLrpiwwWKdXuYZICWrEvdA9O2BVyboQ5DSrdGJSzXwYmy90eNUVMA44Zx06zqM
Idwsjk9vCSojcgU+zZDXSLe2xJ4m97DAHesZlFq6800QWdV1Vlgg6ZliKmgvkT5gYM/Xb6Fq+kDk
eylUd/Xq0KwDXHr+LMilHW035KiB7Xo+zOGHcddYazR07syM/wMHGSwqjGgogpzzJxFW1SE/cMHS
xOSz8wA+q2KpCZQHtsK/lqGbm0g+K6SO8/oawlnZRG8DcMUoBAVBOTBPvoXtq0s2a5ZyNn0FAZ0x
JJvc9MkcMqYMtqDrmOaJdG83moSGftgtuHr5pNDWqU9J39RhqWbvZpXvq/Ebcbwrai0BjFO7SJhG
7Wg3AgdM81FKP3v7ftUTGj3EicPcZfgnD/ylK8nltk2vPosCpjdNKjBIs8qidiRrutdZyKOV3inu
wuRPp7MMHBQGJMfZRaM2AyGnaT++rMJA2TDD9xyGUlmS+hQccbHps14Ug9mRx375SpUOlWCpV1sd
UrAUMm1b8A+fP4Vyj0cR0khgKanK0rJyAqmtrpim6JYEkE7Zcdnd0i3d5i17aYdyn8BgrREQtJR3
31v6TuXcVw2RfvzqkXPHftmE36Gc/lQJl5aAPB7kbw6lCzGhoqqrk21YpKd0oFJtNE6Pj5Ngsljq
ySXycCzRqBEXrpt0ysr2LonhFvUJuBCAToUpRfSon5Dk2Dves+BgRwF0LTVJ8ywXtkTfg1ZHvFJS
e3UQpg0KlaAzWq8+fa9pPFUjBp3rYulGhGwNDceVbs3+4yKlRM+1aVgUAHDNWME/TxIV6CsRR030
YvQSy+Kzm8wIxrDTyWwgGz/1pPCiMAnVFlHMqr7rRijWsRYnquA9qbx/LNrRFk1pK2q6qiL4BxAE
vUFunYCNyliWkBWb19g7r5GhP9F2yKW93p8j5G1Dhj13TWfgCEFV/Vcgu8J2WnVxydKxp01VRWG4
Pgk+p0uHhr92v/qbIBIRzVgGjSYmyIguSbM4x1XHIPOw7Rgr4YjTL+NykoyimmVAUAN7EA4icCYr
SnDCFlVG1as7yCiqD3c9qTcgdlg4zq76izU1a6+JXxorTt6jv+9Nvb/XpFbcVVP3l87avVY0KOm0
mOzV5S88mte35njqg9TPd9hXqO4qfCpAgrsjJy7lcgJCKnDCOdzkAnOQqgrPUiv6U2C5HhlVaYhm
eN3ySid7lrmNR7UY6gnNT3ookaO59dG21FkdwuVeOGQ8d/QqRDrtqViatj4FkCMZ8cv7EdbP+oYW
QLYSeJyKaMr3Ylu0QpliC4ZbT/tSxJ1888KtS2Nvk4C+tLf7ImxT4iFt7O93FL7dVC/R+NsN7d1L
c3mxuDF/zQkKoxPsP+Nsw3FoKrgPiDRCZBBkvaw1SY2RKwgOz2pDSEnTGPJe4QNVdTWap6bscnaV
nr3IkuyfUJLRVnal437qP8o5th2VoG4o6ieCUrewfXswxvpijYyTghwHP9fLOS4BlBd0J6D4qY2t
s1mBIeUVfSQUYPPsPtBLLa1dJrWwx7NYoSy8QyFoMUfE67Mo0zwNkSiNyu6YNXh8pYJFHOEuKv+b
fAplYnQY12miMv/j9rYss7lLzqDXVhlDlb/c6dcHNDeyH5ParHTVgXXvxE6V3LJV+tdm520awUJJ
UQEWs95/lW8KJDZAE0ug3X17RKhbet0KMyLVeO8l4S+SEOJkVLs/g1C7LYTFkEO3vN80WWJURe9b
q/v5U5jTykl5l0/q2UplwLuJleKcHVjNh77SBAFHEBHd8Opo6V54ab/Fy2yh2Gdl36esAMp1XDy3
h2ys+gsh1Xekl8M8vvA003z8v0HJ+eutJSH7Ms3qOg1fdhgSkdJ7zURD4wmJLwYuKhGGsCv2CRQQ
/o87UdJ9dO3QDlX4t3C5E68T8KKt3CmvIXT0XtYs63fZuB0njH0DPJyDbFh5dqn8EEgW6pDCC70h
AJ+nG2XDkFBh4QFit1FuWATdd9MmbSF7REPfHZEKlHtfmb/Seq6WbvfAcijnRxOS89Yu6R+F6R/c
3BkSgYyt49eT0UP04VcJu3DCwk6lYdMkkydh4zevpk4R98Xz9Q0ZJ4wRHeGTBdsR0iUN+Ry0q+3l
8lE1rZoCf4Ph3c37zBV02Dfj6NU9m0mzVrrV6OORXWgdjFoR/nGnBvSOag6m9Rm6e3pF8WmU2+ds
NdSq2hRRWVnYT8g2gZGxQUM4fczSHc2rKRy1brCMu53c0d7Gkl/EkjDumjvPGM0jMEfEGEsl5Ro5
U7yTTBr49WxWmC5P1GTgyiFH2sQxrn7p07kNxxKCi2Q4kyw5l73SKDVc1DgrN+aP/kPyRBZLjnEj
xNFUpOVKSwpQhBlqFhmtgxiwJxOGK0/A7LE+QT3JZGjXNlgXX+NG2Ch8lyx5q3Ep79c4OEKYFDWS
BLUQXGaOtMK6qzjl2q2h9KsJn3FhnKPJCRoHKgmgrctxkIJVhCbBRxFcip+RZRsxAHdowpATJXJp
w5+XeQaTlXmHQ6+Ark0xidAyclmTg9qD78iHnZNpz01Ozut6L0zW0A1rkXNvsoRJ4RwlT3yeSihp
gQsuQIGEuB4LboBWrEdYz6HsSMwMgDBDKtimOOpp4kznOCT7mpUhkA/ZdV/2roEPy6RTzhl04cWL
MZIx1PzzpkuC9e/XmWZg9VOuhULwTSdJEraYN8Mtfy22+c3cKwx78Rn9Qn3GLBEDhcPjEs+D/X5y
n21mLcP8AHMT1g2LmV6GxI5Hj4AePcXed+NHdXNVEH/RcUra6vCcmJM+RF5Mo7lRk21SQuI2NdTT
qDHZhsegKjG7KIMKEyZacZUCDk36Wgykcwct6/In56n8zEBO1AKNPPo+vQRUalsDWLNLpSSJSJKR
kUnHcU1X+owKBLsYu+egegGXXH5v8oGp10By418+4/lWfnmm0u42/sv3V6KmmFNIm5dWZZyt5JHT
yte8gb/kKcj9FCux3BZRkCGStKtjQXvv1WsbKmlbr3KMIbcKu0TS6rrwhTWQkIpdTKNLXkKhpFQx
UJSqqryQWbXKGeveuXo+7GmC85ODgay+dpTkqiVWozlSRcs58s7H++8ApEDdWoEk7u4t0PUhk7MB
EgXV5vai6dV5YhoO17iN6qRUOS+3mDFHaMPiNRGCgZuOyGeUUbWE0GVf6wdZoF34r7KKihaF29kK
/fTUPAvG+n6D23NDMPpq9TTFviRDtynw033FYUfIKw1tnbSLXWLNg6j+7v2TrrWA4LowTP1f+IlL
Qti9pBW5Gg/V4Ql7Ve8FBD0KbdGZ9LdOOpFA4T2CcngpXeveNjFBs9puBZtHe/sjAfH/iG0I6IhT
e83tO9jnTLC7d1067YSjCaMbR8Soaz1lLVwe0C5VjBQZnu30zJ1+8594N3Ei4FzU7rEI8UDbK6LB
+YUVmE9iOVszcd5d20ZO3WSF14lxym3DhUEMql1PrLFe6A/yVeOuE8lT7p0vc2osZGTpazSM+/3k
tu5KyJqeodcW62jfOhpcJy8Z88LzfFYTksrudoXTYp10PBX6Eh8T4UtgNyCHeACZBRJPF62QwNHx
OfRCz5UPAc31WZmawMregA4RTsmdEG0qStTO3ECriRh+5DaXFmUsBl1vZz6THa+Ye41chVXLTWP3
jOA8IGhSmeKxICGLwqv2p1YJi9RJWgs/4qWVGvXqLOTqvcWHJ9tnVLExJI78Dzwbo3WkTaGPZiNh
MTyasDZiFoPMhXuFjUnpb0VQDWMRzmkjhfGDk5Yv+W2iMptuWvN/75Fwp+ogwj/hHHvTNHV6rYXm
DUID53+tcyxRGOfU7f9Or4hG675P2dzOzuhr369aNVAyhLPo+ZsR3FlOT2Ol0olhuE/sChoKBddk
CFrySmZM0UQLb6+bw/koimul+rxi1UAUQdUl6FFgmUuZIwuFfxo/Zqlkl+F17tZl+E9sbwje7zZ6
KXsL8ZYK/keUJL0VKcF38KGCVYRVGj8uukKISFYLxKQm7oyLyf6n4IgYSPjjX7rd2jKMit616lfR
1/ZEfmg5CSfyzevMaHL4iNFUcmMIBHYK/rT/xYD9hDXsfP6alfeuUVbZ8QZ5jbMZtfgrmRxl4JYM
Qe55hq05g42Ou+PiB0e4wsZCk+tUZVtW7D3DKEOL9YqNQ20gocWNYzXdp6VdTq/srZR/faRhD//A
hvepu0TUGkcbE8ux1b1F5IkZdpkrUPgogEGoOBnB8X37LmTDY3kUexdN05+dpLBa9vQ5I6U4mw7m
lCG0U41/EqQJQQ2PSNJv0Q9mX4gFJCEWDyuVTEXJR/Fgh7CxMKqc89kHpLLc6PE245AgfuSs7a9M
Ct/42v1sRp6iqg1WQGTFalAtj0fVqliHZC4dydq1/1BWC3Ai3ExNE0f5thnbMs1E/dh2hKCr+PTI
bWwSZnzvPpYW+18jLRBbxo+oxW5e/3/BW7rKLg1UfpaUeazRtK+P/04s5+nAhrCjxJrmGvHod8k/
ueR3DBmu2eJoyA/dwKxssQA7aSuFcSssoI1WkyKutQcYXsh/O6aqDOtbylgMRSZInaVmgs5UaOB7
nDoyp6OmyejXI+TAyma60I3l3fd0qGlGFbEiyXNLdWWNRxsLUYML6z2T94+S5k/aYlZauyz4yrks
xiWBBO68b5elgKACgo5/vk0iIBqXL6HIzgFqvpzx0ubgUCjJ5+X0c56iQIEcbce1JPHBglXK20ot
Qx70XpqiD5blbOuD3xB9XEh6IJtkSGxpYRiPQxvRSXn1dnX6MojNdVfMdtmyx6iQmNybqBVd6VCV
svRV9PpN23grKajNLDqC4nmNM3CIXd7hKg6t2Sb2LziBJXTiGugHrJ+EQ1H2laVsleea72VOrZEL
VhDc/WJhTNZgxUSeEa8FI94RnIy7FvHpn3Si8BKTDhfnQ5Pts/TwX4cyfUUzUNn1trjYk5DSUwYK
ZLng1UXgAKy9jZBF+mN7MRE/IT77AurMSWjzqqAEiFA9UdiseQmH0buqoAZgMU/ubfINzH2l1YCz
BIzQzmcrkw0xHKKh9m5+oOozmkzvCfAroGASDWILKEgk951EqyOqztUuypQdWUTCfuinv/2oyECb
7PAyxEyNaWdwAEKN9zpURYgeedyE7ZFhjtKuDLOt+MG/rv5rre66TbsXcHFyR34nRHyDBDTVeyLI
iAJlXYVfoqA3vVH9HwN+KYU86Nsu6mkfW5qkfl4Tqa6gyfAq5f9Egp40S9/du9mBIXnwmP61nvrW
gD9KlSi/Z3THk8eX7WgWpVcUx3dQkI6xuCsk64Zu97JZ+npwCmAJ2YsehuMudvUZboqWmkfUeuiQ
VU9nwSxIm532ZPB6KibrJJgC8kev38qH2QlewTDFUFRQchNHxpFJArxHvR6R6y4u+69EDYYxXvDS
fJDcZBvZiYsVcWUsVscmrfyx+U3rcwB/1lnhhCR+SQ07gCPkuheZ3xSoISQmL+bfP+BacuSz3XtU
Z7K1GT9g7giR5PG8EA4/PtN0rn/x4/RnbLD1khSKa43W3gjgNC/3mpMtT+0i7t/LJBW+No79/ms7
/MSCabQfhHD5Sk3KoAXPWIOSMjYv6oqZnONnHNUx0GKveZ+iDNzvoF4rv8EToygeq/M7QB0nhwHi
tHNFvQajp+fGmTj6lHd5CIrsoS/O6y/lvXicz6Sdif0aorttN1+/p0yDtdHGqcfMh9pSmLrWd+5e
KccKDxgD4Mij/1V0pCJFi4XJGmjozdLvyXpqHG1/cLl6qqn9rQoAZFKIF+6b7MxdJr1tGqNjUHXQ
kE7hZB+P3gsDreYltnB9FP73C/vFHL11F5EJ33i+eIxa8XLRHnTvGnMn9PYuMhfcnBZBAtM9KyLj
lxOH4QPVsYr8LFDx1+1PKwJY87XHZcLb+eAq8KRwRfuNqWyHDSln4XWlsmNj3GuwWdukRhlqlnll
J+N6WX8iFRp/xr56go4wgbCNg/ynvU7c/cqTfSKDnyNl0RR2PDd1slb092Ge2ud4AzWuclLcKr+A
ydwsl3LBqWR/+0tCSzbDcazlvQvpSGB8NSDeLcnOePqvwJBrUJKH7KjnaLw+Ln0IZvz0JoHBgBhN
LOekCrGb7/gEoFL2t8g0P8HNGH4GgZgE0d4/4hNM26GK5IrSdqrJ0goqEG05UMmCGup0o1NNhtIW
EVFs6O71AL5emxCfH3/WJ6kXeNmfJpMoI1c8pScGk2FL5lT9guhO1qHl7/wpUberWGqHfOJowJYD
yodqfyKcRmtKlrSusD9Q7D/Qn0G5ZwS5fS0zO59qaIDcWd/ZOLNbOJteCTRrjeuQ+vvmhjQ8raGQ
Q6XF95Yv7Yq9ZPWyVC+/a5sbAPZO2jTkRdFX8VkuwIFFmTS+ZOLxPHN4G3oMvKOWn53nQMXOOJqY
LoUnpEg5PyipyTq+gzoObhJO4PVDLO/odS5iGKA73Z29MzA4mADRA/Z4F+Zxld/AHM/x+Hdo9ifD
uQC2CryoLa3urPNOyBYFZpCTampBWILzvcTFYTFzeJXzKwYsfHBZouZXL9xFcTnExNhtfS7/K3xO
i1UkwqWEXHZeBj2GHADbOaHWJk0lslkcJaG2GpdUeeYhzijry2J5wJexoD+GrCa+PU2qUZeUW5Wb
dSHpQUvZ8wHjNDyExnKCtd5s3NqGWKveeR7YPmu6A+vZO6Q+SMIW9mTB8XMFH3x5GFdEVC6c1FVh
GhQe6qxUHfAZUg5ZpTQBG3r8ysNCZ7V21iqoep+DCOHu43EPgJrexEE7jS6hhMc+SZoMavHyy72O
1IMrT8NdK40N/2R/P838hVwHxmWPGF2lHJ91Wf6gGXkSTzgKh2g9Vf3W9QOYsUVNzze6Q5umacOk
s4Gm/HJDKiBBHOck0vlXLHcWETyPWng8+GJ/gWWYCUXr2IXOw7l/Q8ioojKh9CnieePWlsY5FfSJ
ZoUVr7KYkfCyuF7pENIErolhRFxduwLUlH3SAmAz/JqnJ8Q/zO6M9Vcb1TcKO1r1GxZHSBaYitaI
pkA+i0s1pwReoQbOwp4u8eDrzWyS4Oc9Q+rE//feDKLcuKIXBE5TGpoZg2HZejmknxMIM9+CuORF
dXbYV4obgjcBjdxVc6cphBcWDJi+E4wYujxlKQafAyyAkSCM+cq67D6jolKVreP2oRNt6ipt/h1F
i2HaRGSmiIc32+ZfSfrNzF6N22HQ44GRgPMuEv9m0vpvvXkyPPlq9Ed702FXZAH2nc4z+2kRE8aV
Z8WIx76lwFdt24gFX5i19rUc3MVNbLtWX3WRdhsvDXL8ghI8BAw0O4hmiWlX2JZ2Fyx/kZE52Aam
EFhrhzahoSsh1GeU9D3pwzxu8tLJsjYm58ddgZhDp7blK7VQgmyg70DwxxiOsFtKCCBQ4dFTKESy
Os3z5WWovyar/Wd8w44ecps9LJ5iso+5h0lAlmA6OxABM7dJ6abBaMGuK9iQ8ZzMUFqjncJpIKCs
qhxsR+NpJ21JbRawE2GHJcJpKUMuVDl34A3p3UI/OfRLLW197d9j5NM27EhT92aB04c0jV9Ki6nK
wT4P9NH56LE6dZKd/thMj3Tb/I+SJU2z+5WeixKl2OwwsU4ezQlyOt3HL+kamkesNK1IK4+MTTiZ
Xo+W+0nwnEoH3HkIEqkYi37EHTJgHMiMN6l4XJk5UjSpLTLT8R6eWtYQ9vJT9d2CmnkNvHawLWnW
3ia2oPIaWpRxCzq95/lNLpLzuXMwJ4HcO4q6zuXHa3u6xNdw5ThR92xlloxEyZJncJSuLUa7G5AT
joblR5vH9QQmQoCZQ55ww+xcx9Q6lDNpUfkWHud1yW2dYt7tE63TMRsBvlR6uRAhWtVGlOhZ6K7R
9tNmQEo/JJS9NkOAC9FcoVJrY7gWZF9dQ0OiPtAmNAM8eT8eeL2z2fQxmrC8n6pD4+cLd5x6SUcM
pbnV0VGplQq7BWpEHAiO6k5KmGJaOONKQaqbf45F3Df6r3ed0YNFhh9cgqV4/6ncPPNxHSm5wWgx
BzslnfAYv16BK/1KgLQW1WJmUCPfptjtoVk/BBRTIMUfqThUpVO1oa7lcser3QQXLepfxEwDL8vo
Q6wcXmtKcGpIzpyj+GPabIRjH13jsV+AsAUDBJ25002kJSEJOkBTjKnwIMmCJDJyOGMUSvUZ/TSe
vRQWeWDSrxp7aV0dOo7O9s4yS7cWE+c+gevaVzRjEoZmEIXc8Z5Pv4ADT5HSTPGo2JrzRwgzs3hk
LEWlHPfS108n8Xp/5pC6YEGfGrptKzz9BTES2fAsyIzY6KWxUB27xBZP45qgRepzGcCfwNegOy98
W6mF5Iy8eBsVFoU42PrAGL2ipWK8AQsE1Bv7M34kUVf7Zn8mkudtYS9GIkMLjmzproZhMmf+cPXS
jrZz94B9Y8U+dnuASWFuM605H0w5rLSw85ZTis4VsDyT3sdMj+XMXaEemC9/Jif4ogszDFPTWAG6
v3nLr68tAf5ZmFWMkrYRC3L0Y0i2XVcLCB1FRHBko7WAbLITFqxj1bh5cS86+1E/S2F59FxJ8SA4
PAzLUAmlpOumfxmxT1i13KVsgieL+tXfmKLSNR4761MsTQBOn8MiEjY4wZ8nrUA5WTxASn+SCu7T
12DvIEN1g/r0RwmeDOzaL/lo7Fu122S3Qb8zUlzMHRAOByqDxqc0Bp/UtnGD+1hkK9QotBVC8nzy
AGhEaD/1J+OZwY2qqsVF9VcxXHKMrdcg0L3pYCa9eWuVxf3+RkfrYPR7AMvTSWwUo1b6HS5EEuHN
Xrxkph7Zzn2G81t4bz7ecniKmSvPbQaU9T7AcSdSF/OZradkKhkSNI64QNyI+js5sYzAk7kR1Zsy
ldrQJvsESAr4sObB/FzJraz4RWM5aF5+c2pj6qtF6NU/R9C96OALg9BkukEPaDbY+9FLF4qbXeT/
W3mN/bZB3kjvn8yaOeVoHRkOHvLqJ/Tsa5cfD8ZOJrAh4S0tSb29+9dhbyyMB9gquhc58LMgFj5D
Bwf/WPPt7Oa8GmqsiPJuFVBLYBA0HsDz+v1ND2jsU0shaoI5Dbw1qmaRRNdXvS0F9ltuVOKfR9vb
CZD0fwC6Eyju/iwVP9YBwcOxT0k5JT3gz+7LOiMTTPqeVK5KAscZhhqgs2id9pvX+AAcSWCFIZqd
7//ZuBFfy7vUPb783FvK8OX6QQVf1abfQEyu/clSKorAZVkZiFY4AW5+fyaw288l6G42K+1b1zfb
LX8Ap0CZiTIFujlN6TF10UTuHI5ILLEl2mNhph06ADZ8sc4ArXA+RLrdXbmEhDpKVGkp+9TbuNjk
BV53cRGeNDmvUNgWWRtDdv8tGVdqA/VPTJqyH0OM1kvCK3Sw3eNAQ5RgxJ6Nfm1dHgBysA8g3UA2
VeBwR+1UXexnPtiJzs49DzxB85ewLfAMsyrgoOcgo2CV2jOrIzZjsJR7o1ddUW9Xx91SXZN2tDtz
1g31CAt3Z9FgBG1/p6LPXK52LLuRUBX3WI0V3H4GugP12eIU3zn2VXz31beAxO77sNXEHm3EmEb7
qb1i+vmcrlqzKpOzelCoMKwDcmhw3BZqmkI7+m+pa+OhmQNChmKYbL6gA2MJgglsI4eiuP0Ffj/1
uA3Xo9IwXD58AImFZeuEIezhFhZoiOTVMRAKxiMTReiaOF5ftPFXUvSv+kZk3NQij00O8/4FoUwA
EvMnIExZdanEGlc50HFngWr+2FNLab8vIl5Fw8CbdizYqZRD9jpRV7MPTB1SGKXOIlf4cnkAyQ6L
K7xY30R18yYsPAZt8buC1DiMUJ65zY70Xd0L4ehs+zmfQT1XWlqfn3ZNGIRP927L1b4AtfRDCrpJ
Rs/izG4aWWsimj8R+awzCeuG0NFlWhQg9Qgjoy0yW9VeeAoUbSYFR4oaLqxwSnnYybosGTQJBiDy
H5rs5gdXfc/R7jZz5B2MCoD6L0i6rkxgjqKkCwFAV8ZSlDWoy+QKrfrgTBVDRVGRxSeTVjaM1Uyn
BF8NTVpxJDVdw6o3ScuEDqvNqrtUrOcXCSw6V0hXdbk5eKblhFd7hGxSS24ElbGGIKhi9J3ae1gp
uJ131TZXuqfuRmfRO2kIySzOvsnLu4QUKmWFHHYV+rCN7v6mP9MU+rQAzjTBycIlv6zjG9wVML/T
4oMp9Qd5X6/bb8s22TTmA+Ciljx4fEEqndIMF0EqjDWufVcNY15An/cTuL8Hd5IViz/sgBA1J9+N
Qe8T/X9rBVilSgmfpDy/gsTBNFeYVdEMG/KDG/VyxLbXfxcg/bxRJLgmstBcU8zVw2sZx7IdIhdy
gXFxWBstEWW4hivJPpPdSjPdfudB8R0QMl383WgNSrzt4+312fE97jeOgJAXz8XQPcEd/HYy/iEj
ogzA61A1MgAI/uStLcwW8QyxYOhL5FFfZNR8A+QCrDdDjT56bTZgpN1ys6lELhuDvQu2ys5uCjqT
A7kB9itwb9yJ66LwrnWc7VIRd4H0IGl3UbDQEFZKBiOeVfzJVDxgGnIAL2KPzNcK+LvLA/527Zt5
xzvVYonGXE3klJGJkfK5d/+WN/fRULh4Ugsq8XMYlshi0ZDfzFuFlNDzdYEYUsozPtHthSoc80DX
nfPiA8V7BjrxIw6PWq/bnOD06KWMQy67bQj2uLFEppNqQvHoEL6Q2v8aYe7Dm0jkQe7ie1Y4uUP3
iZwhau9yvYKH+RWqaetJDrqcB/CMUpiHVvRoECBnEICHXTeZrdxGiOSWCd7/xVFunVAzyLPs0Cx5
YdoE6NCuUA5DGZFPuNzRvfGRL+uYFhVFsi4JnYWObaq5DZaw72Kr2P3cp/0vw9yKC0CmiM5q5cSW
Ua1fblbhjToFAesNmPZ3HD3HplbzNKrdhe1GUYonQsn7cMl5RWI+ZE1whx41SLGK8s6Xio4YnT/8
LL7w61iE3A/I0Cyfehsehb4DHIvQsbye2n3p3vAXX2+z4DCkenErQpSMgM0UytdP0Kon41JyCp5R
unfaJ7DJec+OuOiO9YWMiAbLOnwC9/4a1+0qcc34Zs3ZQD+WInH7Yh05RoTWpU0C7QycJMl1Ja8A
cWq4vaLnVL9/i7ZlRhBwYPiu9dxBRUJrrYRMFoiokzbgDfMp7FzlRnotEY+ol+KtlpS69blY3udq
H7TH5dMSBFZQwn51sFGgXb7hEmMlm52kucu+nhV+SPPld4tskdjwmTCOzjhNwq1Cgsyi8ougLmWD
cPXTM7oxSxA7mUyvQ56Wd1FN0pOPS0oIHC+CX0ZMbU8Bp6rRsB+M1HBRTY4mMYJz5fGLo9AxmHyP
ssip8Me3c5QrJGBFJdgNUbeL7maijXpAD6XXJmJKSE2d2XKc7zxnxAz/XmqYsJx6IElW7Y1Ox/jn
ErI+IfTu+Fn/39oQ1ZsrqB/qjGOT0sGsLLgrYt17aMiDyPCquU1G7NThCztCG75xfGbgGuP5prVr
1tu2Q+Ab5Z9RfDU8zRIwN7ykL9OfFS1E8KDXVkHF6mnJAYOdknlOH6tpM03hGWg3KTobdFGJMO3a
CgtDq0EpI/icWXoThRrPCfFsDnwKqV8DqHyf7tD79cZi3H4lpX7UzGBRGlzz9fSU0WYlrF+ivmOq
2CPQBe5ZFkeLOIzSmJerppFlm5lG12BYa0DS6bQKR84yj+bUHSGtfZCw+t4HO2uHXNSdQDIh5CiZ
KThGW2IMpTeCDjwFqyW2vG63WqwqbjZvfu9UHVeZkviOUbuYTioVOLOo/GSjhx6GVA3KoD3I91Ul
+9uQOqVxD0ciZ3a1KqbRNDTUIQ6MYksqBzzQ4K8phaTEoyKV1QhiydfQP2JYBw8I/McxGs0o91rS
kQ0cj+9RWgT1UakKLbtgeteI7/oyitHFssP5UjL/+9HvnBeFTobB0OQGvypox7ng4khLhF//zSjp
dOih69n6Ize5OPTD/qeptGCvJ54SGUGOoDS4Zm6RUKVBIQC50orG1d7GfGzo04LbSXSFk2k8gsTc
tkr7OKPXJTvcoCN0g49acMOfzylFujims2BXUmLqIemXp5lsCyCIVF0xKVUcCW0NVh5Kyg9haQgG
tA5TIm3Ug5hvJQLB72poneowSLKgckC0I3Kt4wbZpb737p91ZCAy3idOg5niPZoX96PlKU8kNU2A
HAtQap3FRSxOuS9NdzK0NAbjLD8e6wUPw+rr2fR/ifS1cpVxb31/V+9N8tZpYwFLq5aqK9Re6zXp
wa/u4os1jMKvNIlpWgJgrjegjAahNXfBCSxiEtEhS9MtFbgIP8BLIHB0sbBCAyaKBpbdkIBLsmC5
fh4vAljEhr4ufT612BsQQI0CVltA2/KXMzhCpN1fAfHPvYBzDcrLXFKCizuVCN78p57fHX5IAAft
1fIUKwOoIsgz8yTXTaDZsDSQGqnFdJy9lvK8qdTGc+JMCKB7+rMODrsrbrMhCrldkDNUt075MqoX
lQCNBbtBFho9cX9YrfYRyrvhjURDoz/qKsYIhMzMfPe4+9qdzLMKQiZUinRk9bAxabiY8OaCb0nj
uSQYHpuVhxrCAkghdOdsi9+qOFGpjee6J6Qya1NX/OGH5hv9/FQRb374eVn1jNin0u+zBoRFTgNE
Y1FJppWycMqfj36pgEEEKJuXLG5nFhohNlNEA7BlYn0BxvupkCdBrLffDS6ItgVFZguVsKa7xvK+
O+1FLcSJFKioZJeW9R3bqmzPgXCJZrNt6wU5RIYYROziDYtz7OC2WOvFU4jcgx9gWMBg7DenbY91
ji1DA0kusDejdOY5ZbJravFiR/QWhhJR4cV1MjSlYWHpR9nmnC+KgMAZK4vLxRh9waQYknhyWw9k
z0KtvOyMIbbC0IX5oiqhkvJtGzAN6+CGQDrNKM6sqRxLqd+XExZpCCuePl/VcwQyedlwUZRT4/OJ
jHigdrt+6W+qt3PtC3eN8LhEqDzZ/i/zfkUCXdGDMNTNu2Fh7YxkMX1HrjD4Mt5nQvgJKX4BVmMe
wHzuCkk/wEEY7NnNGjgDdxAUdsILs3jRLyGhO8sQp1BjZkfcc/QyXWV2phgJSk9GJc+XDvusxIcq
tcBK9p4cD7oA1Kh51burYMMI76IJR1LCcWpxl3gYxVuL1xSJTTrqMKqTccqEPnyGbtOlsZHwH7/P
i/VWFzqmaumtgSKFQ6Fo8H7RbNuW0TATsgA6H/QhJuuGXHqi0ZpXALDKHQbdyH9ZAL1gRMykWyrm
ciXswg1P4w8EOfxxbgqBcYjnphWo9EEM12F7v4MN162G8OiLcThfPBGmPlaAMgozcv90BBXW9TMk
g8c00BX9f4q8aAoirWFH3N4jt8OCbf3ppG/+rGO/UXiinlfpFMh9PjfXO+zK3Q4jwp2lobacfF+9
6EW33Pr/5ljlKgkdLYWfL8TpsAJsI33qSObgRpmWyYG3cuSwNGlPXRfLYASI00ffOOrg53lzzwlm
8h8ZZhoqohCP5J31u9OeM9Woq9/CmOtm2dS0gcId8Gbe8DdPlNBpa+nCqOh6zaciRVE6kwmSjFay
SNPdWDKSMhBkVQT18XWgb1VDoW3WAz1ncPNM6RvRJdWs2RtLkbJyBtFMjn6ITuXhXtVu8pKyE5C1
/UJVQxPfQguRV6DuFXf7VRZSL5YBPwmaikHoVZoiseiowEg5DZxk+WUrx3CoauQgSHnYRZoj1/N1
PfCbzhvvqG8Z5qxSaz9xC8Dut7AYnsDdOPa7NZU4CGKgQM7fNAsVBHrtthdEF+HZMmU6f+ipsqkg
mNkaQ/qAfRxW9vp6J6Bo3D442/gamvYRLv+psQv6qkUdzhIPeG/wpmHDt6kPSC6WDmGGR8UBHOSl
M81m9oe5QR6mqgy2j/yWGlZ1unORPSkMyUY5vQmATCSF9NvzGKfFXb34h8scJvXnhiJNwFtO9IHO
84kRN5DzwG+w91Xwx0tb/IgluW4UimRYsGc3A8ZwnE/OT4OZaR4iEHkRL6ubq8lcr7+L1fFXi9pY
a7rMjZneM64Qd58Mnu27BeG/zab5wFO199DbDs5gi1YPeT8S9dyoXS2t1sLkQqFvBJW6+20+R6AN
HbmVZVZ/LVFj2svUaJA/DLGOgj87NY5+HHb8YixN/kSSIpRaveo/JBLl5jq/9Lbe1Y9e9dlYGr1o
R7OkYBELIZGXRk1X50AkIqT8qMCsRznLmZXQjQJdnsuzDFeovoSjtuvtJhNNZCPHcIakohWSAbbo
5LJiw9YbsPMWsacwCM3q36goR/7ZfL0k+AKW+6kR1HjEQzeTKHGH1HXiAlzK/+RP5gV3LhdNilBV
9ZMNzicy3npBLaUO+HCBAelwMQ6x5JA8rIJWlPAv0dBo0thVgdK7f0VFNq37bMcjxMR70lfrJ+Aj
zcsCp9dySiiepqzLnqF+5Wq2f/MRaa6dJ8zDfW2tWlIQyW+AkOEhbX1R/GwMiZGAjxPXlS4d8uwK
Y/y/MThfvE6q5BuoGya5oFmbIJv4pi0WW8emmC3L7nOVVTPzn6vYiUcjJNMb/WLGkBTnMDowKsyS
/RvgOaTG0sxsyum+r0OqXwRmPFw4e8f0cOD/nPxMUElAUxmeT4sDWgTRwQpH2fY5oRrvzC1PC0Qy
mzXs/u9JgmxqZN1kJh6lyiFSZwRTtsb9UuVpiVvJq3V5ATmSOyJacsabHGDQOzwONhhk2F43kfkA
QW6/jfSIdvsxOkoOb7e/k5P3yLIPj88v/ly+66tyZxB0QVUpKEx+UPO/xQ1vdk2G2JACc9Ig8Qfz
Qnm3BHSKv4+o5DaoGZYCrfsxlEKjZAJFo9umh23E2pgKQKiQF0btwgPNy2CBtg01+PvgyUjuu8PB
pkKbsFi6jaMIEe6PpAXDfSauEuS+MVeLtg3nghy+OHTfk3/juv+thSM0RiGM5ZiRoAg5FbIT4GZl
w2elfNXJbRK6mUTQravp8hTab2KBsBtbfommTBrMSq7Kf0p4tL3kVl9aq50rITTtxpLeNSppkntw
wyfv2DmhXIFYaEd6o6NezqKoK7fZ3U48pGQzB3Z5xZiDr8mCZmnqKNnSZr5jI474ag7B3IWiKmVt
RJ2juaec7nJr4VG9En5D4k30H2eiRXCSNy3Ij10S54R2IwUB8WAcntP5iV9eaWwrzb8vfS2uCmPz
a0YHwsnG7wJEq3C604TrwSoxrTF7JvYrDFvMUXJmeG1pOltXCMwdc0TS/tb8LtwsGGd05+x2cw4x
7o2sDm/z3zjul/DLFnhXmQErZL7aeRPBYdUZn0HWE7FsKOg4Ps1HNnd3n/+Ufu0leNDyi7iyBwo3
OYG24f7+qiZmbsiOHMvuRfv3xtnWg7fsoqTmkOEtM3FcoIDdD2lULl0nE98xfF59lb89j4LoqLPW
gRId+TI7rlz0Lbh3lQsS4KLiA2PCzxmv97WALBXIM6LwsutlwyEX+0UYYx+Bi1qE5NLZBWwgeGoa
t3Cg6Q0asbuWkKSmA2WN+AweH3behg/UdzhpfrckGshwFA9Q8gbcdvCxmO03jFxnG3fGXQFjU+1/
BcZMixDNStzrsDzgxPNRnIGBEtUfH4J0DGpcl1m3y9E+zibOZmQl3XjFPGLKpxhnXixe+UoWlXqF
lU4mHzTAFgSphrkqc/ZBbzijVe6w31LMa1bCKKZD1rBlQK/+3q2nZkY5Zt+NCkOb/r0hsr1YS8LI
5M90AT76sWs0GXr4nkp/nWS51wMW5dW9sqT63VeahZBTj8C4RBsZr8UCX3GYpIYJd5a1m3/OE95g
8qOnYRkimslPybmBQgOxbmCEedg/c7tJX7KP2kkuma+b8YsIIqIalfGlusMqrdhuHWN4H7mfoi84
sX0y63SC1iMlfZW8UTFQfmHT7JaqmERqNjTP4WQQ2IUkI9w4P9gRdvlzZgyoqrfVr8nmOFiZPfZu
yudAaCFJHYZIQqeWGm4MHzpBYsMBQYwsc3RP+xDAyOgg8/Op2gNeh9GGV7v0fqvtMjeA9/R5cysu
BqESmM4GzWQCBJljCtBzlh2s2amFjm3+nP37D6eBFBvsPFKKt/8cX3xuo78G7ESP9YBVz4lapnFO
Ae/4/9eGxtjTUZ7wP2XtzWbqDUx4S/5iPN7EfURI89ieiwy1F0rFV0J2W6TZiLCZ+fAhBJQRnvGo
FTrqaip5InWeIoERcli56gZ2T4CI48LsaiV352gvWw5wbjGVwe2dju+4izt8r2JS+3s75S5y2dqk
RvD0daW/U7UGx5ZKnzOG74CRJIyi06FLnONiWXxtbDf30XLBdGhV92H98E/Ost88Hwn5ZD3ADT0f
D4IWzC+eEp4d8zaZWuU1pG4DI3QTOrqLK6i8470I608KiFSuG9bvu7OSATie3aAEwq4rk5UHVdFE
MBG3FZG/ciiVrWe986T3a+itXXN1N0RrOAXeaekuvB5NZfySS4dVdVfhGYePxYKJUO14ZALKRPY3
eA2AKYEI1LvpkhUHHUGQQJ0sUl+XVtYH+6WV/3T/+b7qUJbWgEmfAjmSYqOfFQygmMWGYjILU/oL
kGR/5wcmEvEinbjjMflov9+PNFsGbWpe+rt1vwbEBbJK1JR0WsaA3mwf/7VVVMGr8lRjWZ69DYsX
9GAyZpP+xrMx1W88+IdVBCGYkjitk1WWDDvdWBcL4M2S1Ye0aj6PBmAqDnLG1OPQgq2bH5rFY7Jk
gglMiTGD6aUw+dJsP3MtcSC+cew2jJup1KUEdZQIg2jyPLDRmPASJePUE8ySkhrYiMwBpdXhY9mv
OikYW0hl/OwCwD39EqnydHEDXGtM1H+p8WJgQ76UVNmj9G+K3lY0ld3rcZ61us5i18f8mcCu7CBg
jWDTWGvlYksIV3y7dO9ccvkwH1sjx/q0dYwo9IOfRHyMw4soseo+Uluprf5Kk7Wy6FBvjV2H3wZC
FnafyLm/8RGbLEpmgNVBemg3SCGC7/Gn9BoQw/tKzDALQZVFrjunKcFBotRQw5f1Lwh35W8bxT8R
bzoZRohJlGHtr8dzO7DAsQNVD4Fx7DzMv4tLpjY5OqHNJOXE2cPNoe+Dnc7ZhhVJBeL9hszFE78Q
Dh1pRPYrSRBOQ0mYn4GCNF4okLIR9yN9NNd24nA55kxQ6brw3eFVqDo0ezIFnPIc13e5J3HdE0qu
PphEiLP4zJLKsiqZLxdZa2p1xYRjj5dP83xPud6kW6pehj8pYeLGImMxfm6w+eB0P2qGaHtgmpNZ
xeYxUebnX3X3eLJwt++gN/zm7ZmEiMAtk0U6eQcJvD1TVGLpXmiOxZnyp1qGz/qpJc702gN9DjRh
KBwCTErRehl+2m6xUQuwNJ2X+bhJRc5S/H9H6EjAd0k2QoJVCviUps62jpq0aX438J8z90D7mYFP
Jdh9hbhf1BXyqoUt0P7+VAJZQAgt0OXT3UtyVUrpuS7ifBmbhXM0wtvBmQnPcuWH+3KmgR7D7Rjd
K8HWVEa0CbvrqOPMzwbFM1Flvx94c96oDSHUn5uQbDEhuBxjqowA9ebtIewOg8d77WOgUhyz2118
qNODfP2W8Y6k2BUnSgVaqtsrWStsOnSOqOHJeT1F4fuU4sNrjb48UPmK5Qk6w+/HbHlvvugkfM/h
GpSt82st1cP6vane4r0G9rnuMLD3sgmQ3l4l35PyJmtTb38PA+Z2t2xhidU98J495kEfKX9mXq7E
ha5OTF3PxBaXwTypRqY89pO44hTK7+hYE43G4Ylzlz55UWB1hwlkeS+p6Yu2zwuOr5G/jW6JDkK9
rEyiZ/Ex3BX4coK3wzXY+TlCz7R4E+n5KVlZrlVAB4ur89FBE7oJqVIEnSwIMWQpZyx3iersvYeB
1Gxw/8DRgEan2wY9Vx6/NMhFv0Yk9HSupj9bfnhVUqWv6GXvjLFH+2HXS2Vhi9YSjXShW+cgCJkO
eegTm7VBIOjlMzW/QHhgtFnaoBOutbIoeyQ/9aZdCKhm3jslUbN363PPzxScM8vi1wHNsZjwzcBK
rfnVCpZr+WiNziCPlwKdgnX2iYkAYm7zoDlDoUujhTxOTEKmus8Jb/C96SR7fM599PrAP4pPrsVA
cxYaMb7EVdZaRLtWoaQAiR8YH7kdj6oFyHZwgNa24kXiHPDVqbP/pmI+dBIWMJZnmzbV8IFBZJLE
+sEubLxYSQ67C9KJmcx4tPijmjeXuhBYVT/5Y4UporY4GRC51858w5VMOl2oPUB7MW/3aQr+6P7B
hb4Hz+TLfUEiDiUx2Mm7vpkWGfYexdV5ZmVXRAfJupd3Ar5owzULSl9+BSBluPct5Hww2h5OBC6V
1bIkG4rcmh+U2WDvtLKQwDPv6ojGOv6vAlLCCq4Oy01RignvG5mAUnFcfIOj3/j8hVOM9p1j9i8a
t5nrkG++jrZ9SZoJ+rwNlG8Ysr2oNAXnkMW1Cf0jQ1fLAcd6ke80v1jUKRa8CneX82PDVpgOEqMC
bvLAkKeByj7D6u5wyxddShnXvX9mWDhTbmJs95kbGDKxBUBjGhy7Vmo8RHXBjFEAjxuXReSiz3gA
NGTOAObzUJREDLbqs1dTsmDGRH8AoRNxPZJ7XR6m8BsJC3mMi6ciADjJk8jHkBJYYWunLNiaVaMO
q2z0Gz1rRTs9Y0Q7Cn2JezpHRMqRdURGhDbZdWPjTt/Y0At4JUelf7u3vKyk4o0nzi5UAqpTE8Xx
eAD5/OlobiHoyUxB5OIr43dO1EOhf0hcsDXlvCWgTSUruGH65FrJSy258kGjtfqRfJ09aEPjmIyL
9D9xjtfuDOnBQmcKvgoabqenwp+Tx9qlTOzd56FeM2thYoQ7rFKQ44ViByhVUUowTncWNTNpUofl
NqcxAX1c6ePMrmrHuQZOv7gosYba3myPFWZCYVQ/wPoQdZitqUndTLwIECFkugFZmvZtL7jCtFSo
Egu4g/U0AckLPLyOvCIyLuVBuynaQ6yVNbEdeg1ZPxTG8Lkxp+FyfkSlo/X9mbvudmJTyQIl8WC9
bvkqjWoKg1bib3guesCcgeaNYrkvvnXHaaj/h/QiZaH5Tig7dC9IyOBLAhmPg/APv834FM/bQXtY
yb7FgfrgKtLXjQ+scRoC1qL4O9grUsIc1Fy0Gn0xV/UlBTq8/eYMzD0jG8YPbSmTM2+grU6hVcZk
tN2XYpgM/ir/Ovr1IgcDJtdWGn9yLg9eaO/FMwHUjpB2/u0qpkjDpO44isA0rYcvhFfUBmf7L4w+
r7cvXN+vik9hPZiCpJItbFlqfnWSfTcEAdfGAcJHEHWE/HrPYWPi/G7fRe8UJCPQSNPJw4nJ6j6Q
BoasSwbl4Ou2gEI3oldF1Xj27kDxhPGT8BpXJ4hJE1qmX5hW+W+FNtnCyH9rgn1+xeFA0DA/RMdl
PW7hXC4GyuLdyBbnELU+47c0qleE3K27NblaZImfzHXy9LPXE38CbfZaHzB8e0xLKm84J3tmbIiO
FgcjvlS6Zr/DvyJ6pOdHxkTxsgGPY4svOKNnlc0OjLKqMXgQNJudfEH+yvB8Hy3k6/S8TCiT7q8i
kXGBUs1s8ABCkMmkYRj/zyPbcyodsf+UJ+cE50Bt4tehewUosvOXsOBuwqycxdGAIiuh/kj9lHsg
BvhV7V9rbElSif7W+RlgUcf6sg3YdeLF59WbcictxamPRr+dEympkSXT0TyTwPHbEv5iwtBpdOLZ
NkknBA7tRYDTbMG8USWIyD0uvS4tmdJtA8jSgdwSh5dajlk6yTuv7cRvIeqcjS+MFaY59xtJzq8i
iXOh4D0dpqdGpNbTp7BFC4FYivy45kJlpWCPbEPBUECcftmwHwnjNCwjBytZKeXWQeReIIQr7A0L
p6yKVRDxSyIQS0Jfkno8gcVwBHmEUh7zyHt7F8GBnbw8AkaDlWRpfFWKy4xLt9CnqIfv9bQb8SOl
3w9T9p94GvBvwSvljPSEOk6rfxNufYJHdz3VKuHX0C8zLU7bi0RUNjG19l6Zapp6Q75V+BhdBwGJ
VJpi6s9eZ5+8DfaY0CTpvVnS/89gDP+mW6q15bl+LQDwURcs0a6RDlFUiXVqCOhm0PwCeD31s9zT
L+FVM7rYgcaExG+sGQfeSSMzWURr+cYdwNRBy9S8wF+caYNu0KYM9yg5vFksL4DEl/q9QaenlS8m
9xbHh3TqYI87h/ec3je8MD9fmx5phIKkIPef2qeLfM0AUJdDRG9HrZf2u5WZRWHE6ik1y33BTg2l
FUwWEN8Jg/QcWC4oQgksG1x51mPkuhaX710ljE1KiCbWT6oldyrQ3TnlNMV9xBSECdxZJ7ybW9FC
W5UR8BoBbOEEe6rqrK4pbHI+jk+ClXeGiLu/syc1XNzyt6+tNMr0FiJ6viZS6JjaeJ/zWGWAqgr8
yIErUEapFKcuP/ms66NuwBsnlCvyBpWT/7yglfDB3PCQWj7CbVfclviARguiqC4txUNQFaJijmR+
EHtn+f62iDZT4iQn73BSW2aGvgtzZJx3LKexppt/T53VtZ3X26hvCDkqv1PEDJzrq9c3Dkc9eO8l
xSoiw+8gbeiyAE228CGeq68/isab/FXVA+S+7UDEBtx1paE0ycRglCmCDzbfXjMFp6ijOQEfUFT0
pVP1D8rEurQ9SSIwSjTsT7t6akGuNHFzCaajLYQn+BlChVJPmvPQN69dmNgR+bkWbdD7+Oi3+JLZ
dLksptVMiO3DPIgfj/uO3oMFPInlsccODPHHNVQIs8ciEjLKkYCw7fS3pEOHpIIzdwWXwGJYqMfJ
vH88eZe72RRGuFYtMxzxrraunB3tuL+cUU1OcgM+T8sDcZDTT39dt1Kd0/+1vADc3X0qQTwLLEYS
YDeM1/QN1LsTugqcYZ1h/Vw7GvCcmyjaFYVLek6aqHcSyAuSHBgMgy9OgNnCkHH+ckfSwEwMNJnH
ISYlwxQA9HsVATjrPI6Sbc8/q8XzIXW02X2BwerDfmJAOY1WNqgJizLsitc8jqR3MukwJqLtVSXj
jHqL9wnbx303xzTSQmJVCVduxaCYEismF/3DgzqlUIiu2tUNpVnYmH5D0DALX1hphZiM0bk9ai2l
2aTrvf+1X0oN3YVPIfNqKaEPrnJvUGdRYJ5qJL79upEMciucYHasH9xTMlR2NaJcqFPTmwjjMDAC
1YIgWJwz/i/D3ws4zc8Sm2VT6iTnL8jyFoFNSftCjLL7hL6c1HnOds0OR9oW0tjiGM+x43QxiCKs
IgEhTndHSm1Qdtm9tExhQfswjlCpMVd+OKKE97p82VAFay5oNv5IYlrdamVLd9HZeSEYX9C7rmZW
zsNG4r6Jrzttpqw6SyRUILSY3YvwPTj68xyP2lTQEdKjMsH9UAfUI5h7lgnpGgv/6NszCyRX8keZ
FnjvJfY8KwM9MTa0g4c1n8EEf98R1GYA0tqv+d65Gw6J65jb5hD0VhTRNpeCe8eI360CvmiKioie
rwdrTPuH0HX7R2FB4bwkbKzbNDN8DAFXdWXDwOYGPF2wn5xYWDGA8eT35G0OkOfX9dRCPOSF+n0v
w3kdlf35C0yAhdaHkVMBXibbmv6EDXX+KCGMXnYVSRqc4AGNZw8ultXhqvlw3QKZrqSDJAPJeq3H
tMwugTG+HFkZubi9/AwS8GanTj4tkEWOG2ilcwlUUMh1X8qED4sUvdjNa4knWcU/0SQIJlMVBBu8
NIVvziP76x2V7SOWWV4lsEy5Kg6+/kHQcUohQ47GdPADbJB1uHew5bXV7RpMqRyl+JW5IwOkOkZS
M0PWLHrhmaDqtdppZKRulMwTXOq75T7GT5K0ZIXD6FkADkXhf07nAwGxVANEmh5qM1sH5yXabrHv
UaOu9vI1yRQNej0j3e8C4bPqLgZ5jyR2fWVF06jJXPLq2yOC4xY87qrJ8Vs5H5wkrqnm1EtUwtmS
9Q6E/qN4niyCq1ACRuj8YfcDZX1BTqio3QKezptify4DYIQFN8G7xzHxlTMBAkmRxropr1rYIivf
/FcGBJyDs5LpOp4Pc9u/T+noHwkc0lQqyew+5u2cTc30hb0jSVyiaP50qh+lS00SeoIjF6CeD0TZ
0ch/lxPyZhOqw3bBdAyB5qT2nAjUH8rPC7jwSjP6jkLf6yayTJbNm1f11OlFGU28Rxzhnlw+KM1j
QfDWLp7vEn5fyEAaTDI4gc51Z0BwyWkUAAcw/3ak0/ZONtRW73I7lTZ/cwpEfCJujRhvz5unGRlR
3upiqxC5sws5IOHxH6ID65mexhvZ41jwtGVvD7svkRvADvS82klRHdQ9UfVe7V8y2b7lBc62zvYU
5lyqGb/hUbBxcJgzNytICtzZIaxEx+eZOGE4zZCVXVuLzklIyvgOSFLB2Ig5lovnTlArESjd99X0
pHm3u0v65Gt4+MJIXW2cRx1AvgxA30J3rdSm+rnVPRcNaMgdWqHR49opyTtjI2uPdNBVo5tKXxZ/
v8ATSkuXSQm9ORw5nNCH3ACZebdgQuP+KK+C3ZnNrUijtIB2bnxwpcZ0VMbwn8nsOjiJ8GREuVlY
BP2tbaH0f5QGEaRB2A0rcSGHh1A6mvhAAkItHbOaJAf8gYhXev99G+9W3UI0n2auTuzzZJpauimn
aWfDL3fOYvEHFmtBGyx7egYwoBytdKnBHUW4bMNBlqVzlzrMaO6uBukSHpPTfWrtghrGheh4Iu6q
eYL2/oSCugMOcuIqA561pu/5dmJGZnx59kzvrNcBifXgebBIsOfg3cunzH2KARa61IWt2hSVx3xL
RhGovDSf964izRr2A3+uyszCnyne4Pao53QgnYODpPrDsSelT65R1QAztbmDAqwxn2Zv724kX+Px
3s2q186ViYqLiJqVC77rMVpKcTKjrH142gqwEwn1PSpsDAZd1ISukz52N2hfYAT7/Cx1a0TNm440
Nvidao5km1RInm/aWWL0t46RFTtoyWpoKt6fgkr2VdCkCCls/RacLLggk4CcBcYIJkbKJqwycqKe
k+O3z5ptI+6BPp6g2s1O+csX5zSZBd/TwTyDEVEBUmYG2OH/kKmDSIBRBzMYgxpUXTxL4/05cZc+
jVqdLC/7FsQJYFTu2IJXdL+jfKUtXBFRR0gDopr/JcgZm8Y+D7tvPofaFZf42a4i3iAyzwex+IWY
fkeYy5ejCbP6+ypyFpSU+QB5pW02hWJemEiboybxMNbQ/rNgNAYk71F6Ozzl8cmEbbqBSEUNri01
Q9Ehk/vc8zzzy60Xr8S7z4WTVZx3MZNthB5H3i7ukyNCAIOKlwpGEXLTo4x6sENV22cDKKsyIvOG
JAYSkZtcfxrvvrnJO1bxQc7fG35D/KY0QAMnbWyARUnSLDjKluHSBMsMWUXijKtMhystV2qTMEPK
IsN2mbpYkZccEvHR1nMQhQ03PJtbE72QFkgsAzTyhuJk0wgqEw4qGeaZVPC+CMv4mga3ZYWXUnZI
pixyMxTDVS6ms1VdES/t7Z4uU/TiVjZCH8nKc2HXN8B4LehHXNpaJWJameuZZI0QHbNR5a+wJw7i
q5wLZs9GTT1bjmFe0PJTubgpwlIAyYTrWHIgx+IKR8MujZbAX189+q3R9jadKynvY1lm0ct6C3zg
vGqwNJQHi8smBB+kceYEIWgRCKqLghdk1si8g1zPA1MRpE69l9duEI5Lnn66Gd/Hy50DANFJFJKN
5dKi592Rp0eUAeHx32BBKapq+Co15CietkA+t6kpzClNbc9sCKpvXyBZghYQunQpVisaL232SN8c
/e7Kn31ioJqiCqK7MG+U6737S+du88k3KC4HU679KcVGQlydBimmJ93LjLNjnDpiEEtfY3o2g6cM
b29GMZgwNRtUYdrxHM+hO595eWHYRWFpW4USdKcRyVOzcYWo7WUnpggC0aj+XV8XlfOlIhjS6cZn
uvptBpsF/WXDnR3yOmej7XYHXHBFBzzQ80n3s3BhwXXVO+JX2jKTShK2YHLm03N4WfWgS4VeN+Pt
W7laJWfDKEI31yEzhQZRAIuGJi7icJfPNTW86uHF5iRhjoe/vsmmR+mzOR6tNU6AOueSfY8Ib9A9
j2FKlWsfA9ijVm2xuqlBo7mbXcNsuFVR6y+t/DDrZC3T4AuCw3ICI1TpPtDxVMlg1yXEe8n8LJw4
l8/Jt3xqJXoFyaJC89FHgVpIsXCCa+9yq5qb9fHQ2xgpLwsMsNU5U8eudTDQ/vtwEFOEoC+UK03H
fWAIIE7n9q3MexIfPsNsu5Q52GGypXtsLigMOy3WcnRPuHAUUo4yWzTo/+SO5dTJ3/uVzaCt7VgE
u25ZZ8wKAEh3ockI/kCfbXOyNOJEX5NJOuUlHoFp93Tjn1yd1WYFlwO2DITJ8ImUdj0ssrtzKx19
G+5HQ3/oQBlh2Oidg/e4NDjEFioQqmO+Z/YPwvUWw0C8z4Z8YgZ4FNDHoSlFUSwlqg81SrmXqU99
X58b105mUmISoWjNxPhD8sdGZXN6MbTFORhR6J/E6fex20SL5HU4KZAWmbV+IdHcQ/w5SlS6/DGt
TYZyXrua92VZQaiYnLTYRVbrUae7nvitejaAMBdKwlUITmGQjC6nI4y+3KGE1kMaMPfMvlRZdYME
Avj7CI1FX3shuGg9r1oMuuC2jve9i+EZrWtejM8DN94n0CykpHYG1nsCqNkcW5sAJ66KIUcN0aZT
mN7O0k4R0+oDrhfxjtfiJedEpcpjhLbypcXV5RkO2c/ugrOEGDjUuXwRG/2RNh0axeAdlCHMGJSD
PiK6UR/j4laHcAF49EYghv32+cTQJUY5+nk0LDFARgFp7Tq2SvvENeajWUFL4z83TxRTkcMU4ujr
zPwzyPoMMGonme4LSl2qIlyTF7hl42kwPUSRz/sF2V3nwHELkEgvs10G+asuXbbW/vZIsG7wI7lz
1YBM/LMdb7bLwlV5isxdgMPXoRrKzF0yegnq6T11QZpusSmnw2f/ZMksyk00IIrQcsgGAnwsbyB4
W796BXwqJLz0pi0FwMDkmaXd1oj4YpMdsVJNW7gxJK5vzx5bwPIIW5M/G16ROcSEZ0E6U9AAQOyL
h67GcqAgbfu8ClVl1k58y5A8qxGypXxRCLoq+2eNu6yiCvpv4ztkUfE8OKS1OmrvP1POpzL1ps9P
nI5xhuzx1kHZQWVt9TtzWPG24ixYvlscYy1JExIwNFMeVM0+BDeWZ5A9OWJgqIL5GUCIAMXMcZbV
uDyrMk0RBhpeh4iFLEXVmsr6zY2FbOL3lF1iUSI3Bs2K7bJndWwB5seMXqFnt/E7r/gukGgwnXk3
a8GxcUsvyoiLydoPBMeo80D7kakgMiNUOTbQEoATPjF5CvJ0VIbFUizc9SUrycnyS7z5rFFfaOG1
XefEKlt/p0Mo5a91JyJSwkwLCJkh+yj/rKUHdjm3+4kS3AX/i96G1Vpfi9m+RrhTPkXI8EwmIr4V
MyM9OT+4mnwAnUHFCqLFkN9wdkadeRnsfEZJLT9BJ9xETuWd6mz0Err4Wof7NapnKCkJKWjBsVI6
bDwIwsBSKGHJufxP2yV9e/hHHsAkNE8ACeSNVUv3rCSLhhzRaG6RXEfeXOUBFK0hp1LdaL//St9O
VlpvmTpzRKiPe/brTXq0IIvovxpHu9e1igZn+fYMo6417Lp7z28ja0kNm0GWHG0iRkHQKUshZJi7
OC5ejSvgOtsp/tcwY4Es0l6amDkz410O5YoDm1w68r9tBkmvckrPj7sVe1RjkkHgxSJnmEw460wb
JvZn4bk7ZSWqnjORk/WeI/InyImwSmr2VuMwSehP785rWIJEyp989TwnYOJDy6aiYmdC9G8iCHmK
kva8WjMZTbuLdZ6JaU3ugSZDDBujZYKtN59UtYY38cszbfMo9okzREZn8BPdmERaj+toD/Iy0VNW
c+fBiLTxHG/ov80DySQEX1Yp1++C4DSA1OqTt3fO1Wgjo/bN5Htrux9LktwzPTuT2CJsu7a5ihPU
nhRPOuMVq+Zw5DHuybRRa+0vtnWye2NeYCwLDaqWv4OVbsTqW284DnPXLGzdrrPxH1niZ3jw/JxT
7mswO8rSJi2Udf2cJMSD5dQtsanZ559YVQE0klhk5zncTD7bDmg3u3gaJlPX1BYEd1kyEw98yeUG
OQtvHD4gm/eU+PcoTKRb7b/DtrGIikldG/yZFAGqcPttU2uztdlh1yZVELvqe2cR0Mu0eUIgvuWK
ZKCCHGn2x4zIAB2py9SqE2EE96ogl1w4opOff0Ymb8cMe4aNyePKkqBcT52YMsCG18Dj/qXxSIZp
8/SteTToBwBDv1LorrjvJ1eeQp5NyQkUw6y2RQ+qCGPpsGKv/Lq365ZqGKYBZtlsiJTDh5Z6d9SL
+qu1J+65jx2mcKnSX61j0eVikfH3479CK3D9EGwvhCu3xN1hv505dH2lX1zzGEUcmPAQkwO3AQx7
eBLSMBpUSnmBoHJqOHGLO5Z2YmCDdUUkDWJUu/tTH408Dx3ShCPnBx4BCLsyyIKIWT0+vB8y2zu4
ai8egnp4usS+MM7GCzKUhTva7jX8C4ZcnkYJGcj4vmBLLnbiqLkvh0W3nJdvLQ0RWT0vVpMSaSNo
xpmraNrLzGclrVp0p3UvPSTB3tLMys3P7mCm9GOXLbCMLvyPYW6xXq3A6LfqpiihdO/SnvdFqzaj
kDVQutXIiqN1PF9hbu3tsxVN+t89BGYCd1nr0MbTryDZ9vj6fAARyrYZOo8RW1yBnWaZ1W/pJo9C
EI/dhCNnWEFHBPyeuioRxtkC5hIN8huZoLICIb9oIn4ROXFbyVDKDX79StAoIz3iIrNxTuUScwLu
yXOx+FPjOgmjlz1oTFFj/xzGunD2d/jxqAObEx77Oe04gJ1UKuMC4kGDXF0zPpfBVJlEVZQoO9MI
SIOPCspBGxeXUz139kGJayS8zEB7SlvbDWf43nmwY82xw+QItogp/n88EwYA6//IJtJvqqjt9Atz
d38Ocg760Zd+RxtERfeYu/boTHXyz041Yx1KYGEiJUgHIRG1ByzjtJ4wQKWnIICsflRxxjZAuPzW
EWjew87xu+gzDw+8akuJL/CAB+uILdRSfRr3soR7WhgnccrX/ph+GV5p8u/XWU8q+5LNfzXIj2iC
bTg2W/r53gtpcbVGAz4ckmLidA8o0RqlgyoX4s9bijtKHeH+ccBGHFyfKkhn3U4yDoM/6sqGlxny
+LZt32V8MI0OFcCtvF0wAtSSF1fU6pJZeCr7qyBXsJjcvAjw0BAvGHHMl3urhhOAXNgPDB6ZHMif
fVscBlKVTl2aXkJ77lTlLjxwbwfjSaNXnFfw+oI/lXbR9g9iOS/ycWKVD07NlBqQKGYwdSUiaMoF
b1a2rmtNWUCfdLmf3cwYMIByAV+zflYFlN9tKwse9rJYZiN/dXFCjwuGm2vL6BsL2S5TUoNlDJI5
ZJyCurgilgYFuNktkUxYR/DIULRVGTn5i9u0FpoOZy9LyS52lKIxsmY7/JAwObwBtvpnwCFgwJcl
6BFamhwcx0G8ezqwejG696oeoQ17XDb8VzIjS/Lc7HXe3f+8sBNmUX4yzEvO8B6QKTmRFObTIW33
CcJy1PnwvI6JbO/QJDQRiQWP6n6/2Vr5LGsTQl1fZuOHixakgx4r+m7v/xJ27oQIgTXbOkldCCqc
FFNsX/ojYOtO7k32wCzaY1CV5vfT8fA5r996T8QYkW+2I0mErW39T3AV87d0fzKatkV3bxIvwV3c
whxQxI3yV4ooe6nqyyy1MWdRw7dcge3GYsQZU7UnMX5gDrdMoNbHdCshTj2zAXegOuh/0bu/MhnO
6wyitIFSNYW1daNkSd3pJCnkFR1+lR09Z22ppCG7LiR6tTpxuPYmLJe+s+7VtiCXwZTB1U88DlDE
fAjjZSgCtGt2KiuIKy+OIDr6g8nI8ktktPmtVsj0y/Yz0iKubJ3gANrAt2EpCNfxzRh+eFgudm6M
QlCgBbEbKUfIuIDEY8w3F6UkOJ9D6QwqZDQ/p3+OBzjuY5uJf8NBqJur9cjlw8qcvjJZw3uFXMlR
Dea4NgE3FmXQXr8sUOyjOb/5OCKvDAyAzb/S3X0NTgSRcoBA/O1ZyrtWTKFEBBBW2IGL1UvpuVwO
AxvJYlDZLsc87KRVvJ606U79CuiBoDR2NGK+oOX+fKVio8bmq7Z50JYG0jI3uLcH8JyJSR6Ai3Bo
rMCtKv3H/A5W6/3enMT9GuPRcWlvra2SEvJeN7z1nmcS9DEkcxcbBhat48AhMhacQGsfQeULVDSZ
MrXwnzGcg7YgaOiutF66qD1ApAc9Bmbg5ftu7UsCRmye2SYXYcr6XqrEAO1VaCDtY3bHoenIl2g6
ZaWYGUmZlXgKZ2pE3CnqTv2338DHP36hO+AJx/01wSZtHIMS9V5GaO26BIB1/bTZzPsI1MS0lYBA
nZnP9Lh6kMh732cBvo8C+NE3fmp8azNInSjXkn0YYK+rXHQcttgQ2CVBU1pF+yv6rltvcczVO3mp
v56+ihMhw8CcAhpJMzOBbiKgLtK+bwj3OZZvVy/eAk8bxoKXXxndfo4aQkw3X3ZuOBv2l5oKKHkp
ImvR8akp/oQ4RSsG3MsYAf7H27GMYpVQxRUJlFvIeDRz/913Kc2N/SXTwnkGkG1dYXejV4hTPbS4
OO8R1osX4BYZxPE7hPMR0VkaN1YTNvsxKORyhpdnTYcxfszKTM3qC5wqDSI7Ecv2dMOoNNsexaBv
jfOATdmTFx934VPuKQSImGYJKueZoxBmnmxXiR4ZUrmUjGtVGo0/rkh9r1rlwQ7u8MAXf8C9QFo4
otno6GR1IUXtaWET+IjTBmq69MbKs+gLrN8D0058tWAkhXIYF/PQftVRTevULvNogyyV4xzRjC5J
nQY+lnLFjUnu+16yFrchO5DBxNol/obwcYmGZw1D51g/oX36h7plaMaKJODke2hGCy9hwkvFtlWV
pN1xxK4D9EGqzlnSdctwaqfka26uGIv+5Cd/nwlnezNCb+CxpKyRrqRPYeelAlKf7xfAwP+Wv8ZQ
bsjN09Id9ILGb+T+o8eN2nnGvvyvZw5D8vBcwvxFrIb/i2t028IrZWnUe4B4x8Vj6etsvD6V/5hz
28rJhRvthrVYCZmDmFwiADej3zvEVgXYYqj6qX7biLlemDygjwvXpSEJ4Ax8fLfznS/5K7Tu4Gxh
+eAi73jYBm8IXutWCHwVruCzkYUaHDv4Cj0L57OT+bvOS5REhEm2l99uhumR3L28AXmDsf9s5Kay
2Jg794cGbt5XBuT0YzOInsIxbS4lRQezOfguQtn56GaJImA1/Sm6ONm4b7dbkTDvYhDB+St5CYkN
Cd2X6v25kjcM3oSHUq6mRM6kDJqnp93gVwa/dpd0+lkiEd692fZ1hDsi1DOAPib5KcB+kLmWnAx7
COyQUDSHT8Zo0E7gX/9rGgM2RmHUcEr4b0Iwn4MhQKSAVEBsGz696/lw27h/uD4Ryd6ct9v+yIT3
pwIZqQhuKSQtPtMZFQAhqKEjcnrTuc6L/jFZmbUeGmo9XCfoPt/lHFuNwf40XO+7cHBFjfewr7O1
6brfdMT7WXGaEKR6AMWYRgxWeJ0WYepbDVOm5R2dhcaWGMsdqGGhQzV1VhnjVFxfQ5Bkr9A7eOOZ
j4mmEH3zJsVLchjjhVkuOgU5puLAhMlKwUaP0hB8QUYJMMDgcFylRjsjVQ9Hf1CZSe8jlwqt7Qac
d9yjL2iDo9mkXQCCNTJH8u8XPsEUvjBbdzEMuem1Fx5Sh7W2tnGf3/o9YOX+YLOYHjjzNZ+p3IA0
qe4rITIz76XtZhoe7LVj0+aMVDBGNRgUm4nobbmwSy4NV5+EgByVAhxQQUQg2f5W4xVmE8dFtWKh
cSg/dVi7jkw33g2LaizM+KPYLxtjb3IBpYVqVQFPOQaF3qyVDbYVY2CzGbMgO/Yg8IKUHPW4+TEP
juRN01+rqeoV9MUbbnuaezgAapoAvgdwRsrgrEE3gGWmuLrm7nvXa9BNKwKXLpkYoNAFpqOKzLZi
O6GzLmrjpxAwJqHEfq6GZ8YIOG7OMc+ciFDw+Rfykvq3kFKCx7Ry/W9PFi2yMe+KUjutr+vH60Wg
xdwX+130xkefdwgn1H6aBYBypkJAPtdlFInuEOW6UWs87dT2kQ1xuC/HFm70N92t9fKjQaheLVzQ
kSqiwuFUr6VSxN5E+MANBVlJL4DJyEingMiU90I+pfbrLdqJbHW7JoJ2f85ze9FEZsUuNU1ateU4
MVVudqjv6+5X6vZ/9erk7iQdKh4/huLDPwCXToCWy1VthSDw38nzNTt2m8P2kkLg7ckE9lF2pZrt
OK4jxuCUGtBxfIq7MzdUL3eeO3zUDtpIe5oQVHklGv1AFP/U7XsB9CSo23f6xWkydzWdkCeta+Ax
bDOyMw71hWgkamqkqiM8NngB6x32cNikpOwgxUq2qxALrNLhJXDg6heqD5gUkkxe+VFRcl1LYRy+
+59v7Y87tlLQMT95tUFolVHjILxqAlpcwhGuGDPFTwIVZXhCjodBD5S+8arzm7CyndFZ6kAG+JRc
+lGkYTcf4ySgJ48QStdnesf/lswSw3To+OpUH0+6FrqihU+x9UbTb+vHD59y4q+kKYkCGd+/H5YV
YhS4UU0Q/pFbxrmeFk7cg0TIGstzRjQjVu+PF7b0r4lV0/V/Zjv+lGggoGjo4aWpYJRHf8r3fLAq
0Lrska6EWmVB3CPG2P+OygD5SQYlWXaNScXtDPDcs6r4vDaHsGqvi1WM0Tg+c9oeTSlegL7WTCek
LYWIrDp7iXRwrwtD11f+3lRo/zxKYvMyyj+GacnTyA33/bjG0SuEkgvEdCsiGI3xTLpoZ1YUJy/M
EBqbJi9xOOh8aIXZXimR4DqSIdjxWrrc77EXRL4sOIUXYq73+nRqHnB3rELoV03tN/9isHNS7o8R
tbGlLCGGjiwagQ6MyDdeUbLWvE0s2Rb2nOMOWaX9VEfTT2YRBN9hNLrgCGRaCNZdQLc/iS2f+m6O
QXNC1q/2zRHekClkkJpaMQPHvRCSHCQjL9IqYqcfk2mREgFr02s9fc26BYYhb4QlbH3O68ImfmMI
hRKQMniXur3uPJL31S0NP4FvdQepFbyh5fQmeecDuOXFBTOd/ZR+mDQzA6F37x8SshtsLPRTy2D8
HgWoB9tBcuaw8marLO1jwoFvZdLLsac3OwmdcVQPgAhh910G7pbwSmevydgmIegt0qaTgZNwB6QW
4blCbwsVi0LF5N6plTKhkL7CO3NgkediP5xXcbpyAXMjgjdTo6EkIV2wukZdz/ybNy4MvS29GEWJ
sU7xG/75JTBTsur/fkwpYZQJHvCuqnN3oyW7RdWdS1Ot4Vbwd3DdjYMCnEol32GmUFlXrx2/S2Q0
U6tTrjKFaLCMCXfn75IQfk/aLFDWmB0fXx34gxK7Gake9k9Sh6OvSBKD1yaaNG2Rb5zu0QtrzRjC
8yezimqTVSUrEmKiXcjvdpx0rBUlu43k39k1nEnKEUMtjq0w39PDpUBbx2QllFg6UVeoSzi/1/rZ
GwFvZLH7pD77nn0+SgJDEaZaGol5K9LO1GDxzU9bfHpf/e1Ea/MDHzOcupu0DjkeTSHcA1PBLS6S
S1Y3DjnJoDzL+8T11PT1ibwffhk4dGgiGZuDM7To99iSYU0itTKhZiVFsvIbTInd4L+K6Z5SBYQG
rQQNVRZIbQJcOZ4/ttsZVJfbNVyGfa9oLHDgHL5AohN3CSJ82IBzlyxf7a/xCS8xCKfjfsmHIC1x
es3LEqxCOmMKmJ56owKBcfjdcRyVwVrjtCrpBNWDAFdocsBGs+miP4rHtCPFIFCzthg4Nb998dGB
pkWobmHo5zPF579LWlo4vpzMXXNpc2fWzvBqn22t3yr+Jc6E/m8wUTzknWMWg0/n5IuynC44lQEA
MFn8toudSTgWlhah/8EG+xvR4XyKDACoxGA2eC3L6zfibsHfhaDGfm9CJBp2P053TzoIypLs+Oms
7+Mytvhn/C3dcuUwQUp3gXtMNT8fZRcVCi106qDFp1JTiRqnHuzftNesmgG0egNq4Wd8qq1cgB7+
9sLUw3Q6kN7771Z4ZCfeSBdzpdXBoUdq9a5Eg28DTWp5YuhtsSa65qQkvqLWTfIFmjyvS2wmm+nw
WYo6Ick/IejLI9sja2Jis1BRoIdFqPOs/BI3RKsM3SvSn43iI79Yb7FdHsMYZhcpWUPJEuRXqEJl
WhAQT15X2HjrwlPsWU/L9UO/slAATHHb6URn5I5jbByTMGoc1tYwWihqknRgflaZ2ZxxIBu7OYDT
UNsuVHK1l6cZS4SBOLF/dp2oiI4XLI4KeRRAGU127I/IiHu8Tsu04CU0QTlBV2+ZC4hLhQb7JTOu
Ke1xT3WzqeTpwTP+r9thj3uK13MajkLq7QdGKGMIhdpHqtSUExS0vD7+7zH+AuMgN4yJ7J6ro7r6
+iCf/VfwpJM3S7NjbLxBJ3DUwRcVsvoaAgtmMtzxVI1UdnEGYASLr+SVjJN0wWM8GQcPptYsNnA0
iNS4TERXjFBpFkPuZ0hdBN/5Pm1m597+qr39IBFyibU91ksKKY54N8q/mCyFDBJ7Xl4Kb0qm8EJJ
FzHydv4cecWsy4OQNrXPTDWY321pud4kDKx9MHxx4zFA3uf9LbSylt4yULV8izTqUsnbsJg71jM1
CJyKFBVTmkqDYfssQbfHWXwpjWpEoI3yOGm6QGMWsKpbAo17ojeJjoICNoEEDzdmBq2DyrDemcNY
WxhiJYWxBNVZ96d+O3TBTw8MfAXhwz6Fc9EYiO1xpNjFuV6RQaHjUYEJ0zafzSALyKTUv9ckEm4u
ST/NPQKog8z/HJjCxiUveNC+LVM0is55pG+nDCJCDaFUke85g3zgIDyKKZFwNEUjxOwYfGuoQ1s7
iTZqeS/5viig8Ym1KBgFX2SFnBRbm8bVXQdB+UdZ+tpfvNQBsXSRbAuu+fCSTUhs4b6C90OKy7/0
xJeCUjsl4OcoQJ1Dz6IKh7e0E7Azs1leAQFyJHZrqLA0SzUPkut2Fev+8NKYAWxBEVoI/Zih0ber
W6xVwcT6t2LZIhLHCwV2ZLjwhC04q1RKQuejLvFOmtTqrd9GllPUKLf9B3US0uRlWVQ4slrIYhqq
KqKirTsbS/ylXfFBbyvBAQRMSmiQclIcsfCjAZByQ4hs/U5AawgxrhgRPKlfxvav7byRxExckyvY
ahbbJRJOA6rTgNgLg+WE0mmww9zPJcQ76qmfpqU4He+h0JmcmkaVaexylIV9xoUk7WTXTraONdo5
GXufFl3Xhn/qo6FVQZ1/G7m6+j/tvC6eBybPsV4IEmnC44JWFkRHqcLiVA9l/W1X4yD4sRVD4hVm
m1c8YIxe6HsWTKuefMHN3sUjT2TRz+FgMpRRWXaTQvVk+iTBoMuA+DwRxN5TnzZajJhRYQN/Gtlm
uERKKfNO91feFz1xee9gM8wcjRuDjlDJ0pFEY45nZJ7el0U+p04uZoFJibAISjglR5ZKtz5UhIvD
JFN5mYYnIU6vcCh++hk9zB5gJsodoK4R1J8LmJX8sb+7O+f5YE/XmDcxckRaO5AqG06cWlFtlmbY
IB24fR8Z3XuL0Mr7XgbJLxlAZ61s3pRKS3Oo1lNocbwhG5pzmsxul5a4LtJaCmqa7n6sHh14fNDH
Ato9a71+bjqtVsJ4ZvneNHxa1NOkHRVYVPxgd5Bcgea+shNeZLR1ZHZpGobDfEI2cHfTLtS+EK1X
iF3DvjFA2yDD2yBWYI6Z8PFt45EgAPkFA+4m20iY1IVqCqc+WS9tkJtqMARolgYXz1VWD84Y7SMs
gtnRwV+Jesa+gGuIHTQp0kYlFdFMz0RQXj4gWKqtiTzuRe9PpQ20ubIcRSB3TLXmwpL4jDSoNz31
grG88GIb2NtoZM7fIQsJT9AvQgwl1QTMeuneTgD0Dc6BnsgsD+Dy8guDOTgnmbTKTZCP8t9UwZAM
h+jxU6n2urr0V7xj/qd8A4BWUmB7eMuPAlyDHyiLH60GSzoj7ilYLNq7F+lQwTZSzqPHke3voYqL
Cpky9WRBtam/eDvFdx8cwDqXX3b8IZh21Sxq2JZg2WsccFNXpiJ6LrXpgMJ3rj4nKEenayRmfW2L
QW5j/tte10Q9AWegDWyXiwEZlxqoI6ZcC4kl8qn4YABlWBKkQhj1j3bcpr++xSbhlI2kUD1Pusig
/RbACJ5jF2jYebhPgOX10v9eRXMsmji2ly9Ki+LwC13k7ShWvfXaqwudCejalCShZJhr04ISKhM+
+OiwcXt9PIs9GYoXUw7KHRbEghgoh7XQK8PNU/s+qaOE4JmZUM0muP8TT1/tBfrwaxNrQoNVo5xK
hYX+l52wedadC/IaurTL49z9aXmD8hGJdoNmASNtyd/ZxuaEvCY27oCKQx3BT/o7qa+4h6yLhCig
I5Nht2H7O3fsfo02/0Uytvjr+3OWjH0pXMzdwaKZU29wk7PkIVzF0KeSYthPqDE7okfNyuVkH/7i
FP99QfcAMX/NbXOmfJSABSFkMqysTZ3wWiNcxL4bdpSWLBmKpybHwoNeS9OYUvfBgfhG7aOBI/7l
HklxV6SkYGJfrbXLcL00s1kuz8QvHGLqZicW4KmBQ0czM/6pZT9vWHWIstFQRS4CCin/0x/59u90
ecljeVZ+XLPkOF7T+1Uxox8tTqeuYP9B2Ne8v/eGTUhrEOm+/jFdwpCNhQnNQItzpDtGEWjHcDjO
ietPB7Wcc2VAjrS23qQdQMSZaVDI8Kj41ejirpey1+WfTCmy12C5WIxMBsDiqs8sgvpO717yXXqQ
BGiBgZOljGdjyXh8AdT8m2VzDacXWe6p5Fd5b1kO2qHL6gNGfOL9SBlKULH0vJrCzGPaOtk16K4o
x4o/0QfTwcQ5KNdluVLSIrDB6bM5QP59XxW4VrhbccIOkflTI9oDCYPUp3WZsQb9gl5vsb8g+zKt
roaYbHickiJ9VnmdG8r4PJGXNZgvGmuDzxDLhf//sG66pbMaB/RFxQTa2FSvt8AHtYwnkb9xPG82
n/A0TJxom1ZvNjsMGSjoWouOeCnviu+tK3hmtvKf2znSZcxy98ZOh5cXG/GEyXtsQmObLqgSIG7v
cz08nUcBnz/uc/0VA30vQByNm/fLqcfvHjQ2eVNs5t0aB5okZmncPTXzG0ceLD+dlatK5fATPxVh
KqUq41IKu7uu7ArKCkJCcPAbvBxwknfAvxihOaCS/2aZuh7Oxh7P/hC+09cvNxxxjPCottShIpEH
RBTkKA7PV7hcc6uTAzsgwO60rnbWeTO6LqMn6STLDDnEtgJjj8BJ+OsfJJZ/nEaMK+aO/IQFSbyx
mTxOTtMm9WGiLf2Odk2jp37LM/TbW4a0oQC12Ditt7PD0WNjoJEP4jLIN8+hn9LlnZnNmJJqmheg
StenBacTHOV1gY4sDf0UehkjCeFL7TLAKe+WW6l3oQuQNqEAizGCOHLqfnDl5GRLro7ETCfmlcX5
xzo7UUWoreQZnFZMoI8OeQ3ShZCBgks3cx465mA2ZBQbukphWHMXhZZl7hRNXjBW5LVFsH45+MJA
Rb3H2uNPAUPRkXtHUsf9lTIFWe6/urJQu356BBMDoDesvIrhIsC3cNrz3dQxNMqDjAjXXCG2m7iD
M78WGC62Gr9tAUZHFey1pkKpEPx1/ijv6KbPI87donygzI0kzw+Otq3mEArMbU7VR4E7gp+YyGi6
lMj5T8sYViVDDpI0CDUMYR8ObfNP0x1uSkNV4ODs3VxN1kdOl33/5HX+1xoQAH+0fwsfhRWEAhwZ
GL+41zuapx7iHgexAPTBsHi2V/SbdD5bR80MH2rnf9w6GAZeL8s3KbHMWVdOfXn6miEBwRxJVDaK
Dsy5w6P48Fk1H7IARtYlmxft8gdswkDsSr6OZf56iCYWrq5S3o2WUsfdUB/CM/6PGBsCKe8RFFRR
r1hXvzFUp/APrj1Lik2wabiU4cKj3midzCgeVoOUPo6nnm0uidImPDEbjy9x250b5ZNBjCg+3Da2
ovRZ4eTsudLifIC8B3niILWI3543gIzXMv+tupDtCfd7wNUuCtyzU2rbhzMh8yfsow/INarw8hVx
AWS0qrztqr/hdxePojcY9gffZPXOcBnjy4o8u6NhqgUET4tbIYiZvB3PKAk3W9srh1XhIvEfhPFC
g8fdu5wHurFubGRpNxqwKPY9ue9pYIWTQomlAU4sVZU0sVZ5+U/mz4PwjP6Y12m/1C7lchjdsQPx
tdUoJjGZQql0f840eUsU1mBpeQ0RyIxFGPBLmIR1pBCZ6WHPULP0HFAaq99m1waAglAt7s7NgbzC
+zBuXtvK7aOI85gNElyKKv40tECnI6ETO+7AI4tvMxR8ZRdz66kha12F4TMycjgpv7wW505Wq0Fp
MF2UlaqE4xb7rpq/v+qmL+Mi6goFK47iCgO6BCddvERAU+15exo/v0OiWkEwRMBxXGBxkhZoLdnr
z1aQP0l9SF4BvX0Yu4a2EajprF4t2mt0vEqgNE1pL7m+4g6BcM/C86M9wh3xPZytSP6NJJ61OvaO
qPxVCQ9Y+x+gpBCh7WgGsEF+b/gmBrjViVBvYFy3vLfUgdkjb/6HhoHVwEhaTbKrv2R3cKHzZEM6
2SmhcMYmP0utqjguOqJDc8O0ThFW/ymWMd5t8a1KRasoasTenLRbTvz53nNVdddWYQ0yi66bOZQD
dc6ixpysoNZK03nfu2b5mAVrWP7TaXuNmXWiP2J3pVl9Au5KQCdsNq+nZcIKKjn45/u61+hZ9vda
oGTCb45YZLTTf0zSJrQ55YXhkD39aTQvFFjL9myQCso72raOpf1FlH9G8u70IHX9CsIlyeINMSoE
TBJzfta1o04HHU1M5Cj4u2/OynFqzh89KihqPJd6R+CjajKGSd8potp4+wuiXKF9OMxJL5jz5Zoq
ILzdSh3ZlrXimmASbnW+AowzY4VvnE2f6SyJoI8z++Cyew5y66Ru89pqOPHaWGZRr+ghmjNBBqbE
Veu9vYb7Hofd68Jy8L2M7h9aygh773LP9wDhMALUNvMyWg1GxiD7v351URvmT7JmMdhdq+Xsb+3Q
A1WZhnAD7yfY08q/UEdGR4SRXIV3S+HOeCwQtlwiFtqjY31fD+ue0qv+wGRNiUdXiuuj0UV4dTI7
/2TKhdIkGgOWkRXRtQNextt5rZ2ms6DCTrpUcDmdAF2tHF1EhFc1o2j13aH3PdjsUkizXdpgEWHr
Hz4ryDSC6U9KqWrhfCuge0Eylg54HFNHNwzythF+ib/FSDBuz8Mkqd7oMMB5s7e+jy/UC98/MulY
HRGCyytQLIVE4x39t2ApAQSQpjzlBp8kZxuaJuFJISX4vrDWWpysYaKncFp+HDjzgRLPce6meo/p
1F1uVnzrR6hQko6usdhb54EiAEJ6Zz4Y+NiOp4l1HoKK96d0gmsQcgGAKen4CQ4hIWR6b6KneNvq
cwbOfCEwR3HTJCAk4EEX4xBsTKlRqNQRu/xSd/VorQ5iQc+L00O8NvpnGk8z60CwH+KneCkqrb09
21ak5Jo2vhx79bCw3s0Ozh6/kcvYOSvlXX7u2dM5NK5l17OjtJNXz5pUI6iLG0R9LidHAUjZIQGA
TG35jYMBaA1f+hpFGZ/QdYiJbVeMmCWxSgb7kL8bK4syjrAxUAr8QtPJ+W0rMWhmHnbWe1VPqXIy
qlCVrCNJEpNMtdf4cnHJa8sV6/qQnir3yGysf44GpKoClEuNtTrvtG0Vo6Xkd49OuSRQP668QNU8
7kHeW6KyWPr6eO6gaWrt1xxeXN9R/bbOxSc84+OMzWZWVXm22zCQg/HeoD5qe1QxSQeRNKlwSm+Z
zYx5mlKno4IhHVpyMANXSuBt9TMrDK8OWqElzeO7ivdxqG8zc5bsMPqEuv7aMF0GFn12xT19Wc9E
tK88TrrdkrPfwZ9HUNytLYjSRR+yFoCPAhABaOZXZPVFG2X6+yMNV5Wn1zkd4EJxOJeavhJdxZJj
0e1MKx+WGHtWvPQx6VonAVCrCHnLGBGY4ZbKijSR/PigO42ya4zCKibG1pcRx4V6GAikyTWjoCsH
wsz0h21hKJmNQPFVSqdP2lxkEdhpJ3Z+8R3A/3j6SwXeTLWWF24KBTneKXIuWk3a8bCuYENcwyfu
ngtLxMzkPC+fpZbf6d3Pu4FdJtjVrVzQLCHOVvzxdUhJJrNi/V2NjQXvt/A5m1FSfcUQJTm0WPed
pv0s08FuDdCWfiS9xprzpDc1uBv1H3P47SjcUHsnBLNkGcsmG2AnoHVT6Mnj86SriZvw60igu9Ch
BuUPpRrWWWlqWPdZ1ZzoXJICQpSL2FjXnSD7ZBZfutbKVMjkO561Syoey2Wk4k7/n1ARQCu9pjVs
/X9ojRSvMHmnuE+zTfg2V7mwI12+fefbiNOnT6Wi/b8pNs+/v5CE5ZOMB5gGgraud6xfduBavxP5
6XJbj/mWvpYm5kAl0j3ZsFZAgz5XZobC8fHbc4Gj+aVA6UyoDipjrC++2B8B6o8lElvytFxlKZWf
NteoWP9iXcK1yWfNNvGxHSirJvImYHWVRwEoCqwE6ldOE8c2Xjv/Q+JlVqWIzZF+WfrdEE6WWT9S
PlXLXinaR+nIajNKRTx7GcmkyZ1BLFvL3bOj/YUrRhVEraOHRazQklIJPOTqwIjvmmNvoBFhewGl
2jo7RI42P9gmJwRGM3unGN0oQxDuRbT86DwgPcL2ir17B14fbAUKI1p7Dy3QWFoZ6kilPJRUoAWT
VKVWYAgdNpb+Jb9ntxr6tG8hgIHueVhRSL/fEbsC+NRBlh1WUnvUMhh/OstGCZqTqIVBNm7r04Gh
POJNBxoPLsnGBix8u0W/F2mPRLp4qaYFkrz2QTQ7W1DPv5YoYXYd/6ebhHp/ETky+LkSpPm8HRUp
EBeVgmICN8qrxdcZzddgmqQakUVgT1n8kya14germcrFbcw9Ye4CEjEfeCKBDaXOnmVJQXR5Xtl7
5kI0oPnIe1eg4CYDEzgBFxLGcLLj3zcVsKpK1viO3iC5iBRhPT64jVcrU0x75arS4tpxX8iwDT4N
m4EGC9MsOKXpWwp6CFGx9S6EV2F7PAxtGSRJ4tOuTwnY/U+p0nn7RguRuYkBe+9ZgvRRroUM4RQJ
DCNVhCC3jcJjvWIOO9OPUDTioHk+g81Dh+8dCWl7GWLyUmh4vSyC9ZiRFbr7JI341xAQYvVdmcf6
2ocuM8WufVwUwxhA19j/D5/WuF5mRPFAqmdFpU/uPsziqV5XuAZK0aQx3a7H3tS8ajKMhK6LT7V5
/dJkYSM9R0udXFv3Y03GKVyy/Rb5B1K9rxQ7JreiLncvBPCuTWbMCwYTOhCPlRMXwxdveCXEIEHh
Igm6rYRSIXg1s0oboy+k1c1IvOr28Dwq8aBLmq3FiA3Q28EBOr2ewIWbTmS/cmiWiI3C/ha9bVED
2aUsVS3NGFpwANvOxUYTpymaSQ4zcTn19YciEZwiv3u/FxFT14SiMyLsv2Qe1IB+iSm4ciIi57/0
hMDRnboiluoVtS6jwjyTX2GBlZr795xUfj8xtGDNjkgFzy4IKpn34IhQ50GnlBTEFk43hcZWiWQ7
gAJKBm+ulJedKrPc58FfTUV+Ga9EOK+HxSGgWVkczhyc011P5Xup0oIAJo+C1zL46JMfeTd7DVjJ
z9MvHV+oDeLEFIsdT1Gbm9ZJPn4iDNT+aqD/aHMwICsK9kt8u/VWEK4RgYdkPAl5t8epW9htcKKO
Yk8PfB6m3AEjJ6YQV2cbxmfCHHi1WCZlI75YU+/czmg8ea3juLbgtrmQf1lUf0Wua49n0W8vECcB
bpCeXOcfrqrm+pemlQ1HnfbjA1L+xfJFfT1rEbGYet4z7uv6qs+DVM43HHfwI3kwBw1dI6yPTZj2
Nr/+LGk95u6Ormc+NCKt49rEOFyShroP5HSwiSYF/qS+oiSLPyDVv2XRqOJ/uPj6v/qq1Ayd4xX+
OhZ0ccK3MRhNabRn/f9ucdMw/YxGrmnlXixRJHzR6n505FJvxcZUddIlx7ttL0sJTKt1dtTC6M7q
lgXlKB8QFAu1Ri70A+YeLVydyrc8FQTnp/9ztYTOQauiV6+aaUQ+bGtG25YizkbkWTZ1ZGlGFoPO
HGbzQNOOd13nroAP8k5ihpFvC2ytzAO26ictnkYh6kpoMBZczu7PDpxXV40trNPRYtHACZmjS8e3
ZybInLqk4pDPbnzWQShKrdeUrwGt9q8ICidWvhMZI9akv3HyH9+IOTGCB5MfvfOjwusLfjdSXk8+
AmMnX6YVt4GmwjgxsUvws9xF7uKzZSIcFI165WIk5ZTsRz84mgBdqL827ACXqH5lJwl0VPIEsrsR
ZwIJGByuP5rADJ9YI6dG28rpyE4ak8te/lG9jLTXUE5bu/0X9PAgHf3oHdl7lmOcElj0ClPhQYZh
kNV2UyJiCsuohYT5AwnQutbfiu72GPCUQGB8T6lN0DjvZGXGQ9+hYUA6OWFyVEqzWtFmn8fRGYC+
kqQJxqLZfDp9X5k0FikEE4ZpfxVXxsnqQUxlpIKpbcfa9t0vpJ0Ecp29zuo+BB166sIiseCkonUJ
du/1ABxmr0bmKkS1e5vCW7sOAshzD3a96G246SOa4zxYKw1nnu9aX4Js27RRw+YDHI64H+htZ30h
dwPxsQxFC91V+3HM6cXtSZb20awZgboM/9bjRyi8jJx+PGpkswtV8FVB3xRCHYXL+IOKU7Vih9Ea
BStBTl/z3LkjRL7zfIAvUzTu846EW30vZpU8rECvEA4VURFVsu3eAQ958UKjwTyaVsNAD9eFKrgy
M2KWPm6GAlV67QuPftcK9TeV1h5oHgra0k7fqysoPemw2i6MA4Lod8EpAT14QdKiRagEAGfHdzvX
pcbEFkQXsq4U/OgtRE4WvWVU0T5VrZNrr6/kSnb7SFxP9QOig4Yxbyx1e35TrXZAu4fbqerQ2T5m
Y+L0ItCObX2XkS6cVk4b0jZ9nSl2J3pQpKjEDhW3WFqIeEcISZf4t5/a7LC2iHYQa6ukOiBZYtU4
5dVXjxOlcIFXN6jntNLMDzaVRKrplD8mzz4XYJ7b3FJLyJGK+4kEgDJS1i7tB3It0M8/JKViulUM
zN45nujZZVciUbuh8jfX+N+Kbbfd2eX5zJ5uhn6hgxbRCwvGrRcKoC7jCQPs8GNWnNivRuHCfeOK
00kzzgUlUVTI3r/Xq1uiqIzFykSCL5xyxttH+qrgUl4dsjzYfNKrkRMohctECkO420Jrtq0w0VS2
qYxIiFiHljeapBdJjnHnpjSXf67hNz5oSgvsAvr4+hTG3AzYiR7be+jjKwzZsZkgkWGUd4ulA1n1
rbMwCPaC1OsDyGMv6hIn8d6tdnqL4VfmngR1q2IUgvvJXlvsbvFairYAqmn0bE9USMAQKDIVnLMQ
FDJ2CSlxQJC/wNJeziAHpoTkLbjiVJqTu2SKdfo2lV4oZlh/E0WSjZCKXGI2bLXK2KYRA2GndyLB
ZKKRz8TpHNhcsqu7m/F0aBmpE+6uoWqDLizhQw2+0HYCEdawg3oi5r00qFyDVAWJc7LEtgaKpssY
u7SliwzC+0Brm3q7HkmNtaZTCzq4YpA/sKq4K3V8pERfc/ePVTPLj002pKugWziVhMF2q5udi286
8cbARZRjMfo+bV3Po7npGpqlo4WAT5cWoR1CU8rMsKvgGv4xP6QPGVwQnoFLcl3C6BPwp3sXgCYo
7zxu9nTw6TeEmyYHh/XlBcyOZV9t4V/vTVgfM4nkO7NSceTeHWx2aJJCsNN6/cmW7oP3xlLtObSv
Fis/ZxAhXhxPk8PGjri/ggo0eGvQ6zonbHejNmjJ0iS7cguF91jvqNga7MWAwof5Sr2vokFpb7gb
Wmuu5pjgBAHzzKM6MoHJcgwn3Bw0cYSFScfhLoajlHasliD/3fwchL4eREYjjsw2//Q2lOPmgcW3
BRlxLpKl36W1dnfuoE8/XEYy89635hC7Bhz3iqJyM8/9267GAcIKfXXNlrb/DUO7yZmBylipDSLd
o9GfmcFYDzeY8A+PHqRPDVu7rXrzl1rU/JJ5AzWL0kLn9cywn9yHG2tdN5R/4Z1ZwAMkwr/2KmEN
WH7cnotZbtpEzzj/PvrK0e0rej3pEhFpAv5lCFS4lNYjIDw/SWOk4f5ni/Rsixtc09Q2maDUNbne
WHxtEfxE3S6+bhhiQXmRLm8qucJDP7F4penmqWRETqljhGFkLpbP2VtoN1Wto5wXtNpU+7wtsTAQ
UmJWBSqfUGhlRqFgD7a86S1fBNqqcbSC/J+d2JtyArqKcErZwVDn8A3a61ON/SJ7b+K5cmKoi8oc
jxinHqBMEn9dzsOx2aaM7IDF/RvKqZDWWG4HbcLWC9p7rMOlkp8e51hievX/sFt60k8nlvej9yhc
rqAFJU0G8+FAAIXcorPTKTEjSWGyGPrryKunptu9Saga/DDDGIpA15eo0DhfvCdCRVKbBkw0UXat
xkMJWKu1S0JaomxSRXGn0wZGWXoYgkGXTm8yH5JeVEJaN/3+3zszwzq5OsP4TJ+kOGFIAP3Bkqa/
cj+wWUd02eXh4OwlepxlLokpszr9j8ug8DmvLXMKaIvGcUAzfMn8x4yTt+62yCd/rgRg2e03nyR7
U3VT0SpHkmSvkDbGaZm/02o+4d8EP9u43bYBgd1LX6fwIU2u4t8s8FJxg4CtPLwiRvpFy1tuZB0K
AE2j9zMV7Jzs4HlxQ6FkmQByIhPgnSGd7kKovyVKzyrvk4uBL1ecy+s6hYKbzCFKeDuCce5WjRpL
7lVlJa6/SbTWxUlAaqdP/9b5VeX9YwCLJbVrVTDr/aFaTyaLqMl5LclhlD2aejwbK2PDgPLFvZ76
bFrHzMnjw1XUNnbcZ2Q7Md84lWjgDBuuAlMk2uZrOzYHx2c4uPm9f5WLYqPKX30+6adzyVIovEok
BLU8OSVn+ZFB7wFvQZCA566M4I4ETk/YV3zZaIPdwcT0Eyimaf5YzKzra5YtShkRCReVdUgWOunG
H0KQs/smds+9XFPnZyJMLIWDCjhVUcNRBbYbIem+Hdo+ufmOg9r6+WDZv+6o/GTzofksQCKCtoBd
IJauTyGYxggzoGp6fp1cUFjbrjptgzhkjBev32Nj97S/h62iNakuBxl5VCWYMj2A/JXkNcbpn7de
JIGUfsnW9nzOukJxMiii9TU5RgQh3bfgw/TUTyLVKT3pb3owuzjDIH7mp7pRx+ZkjxsN0rgvENy0
XscjZ6RSKqxFbv0MgPx7ceGULlEpLD/1I1n/XvIOJjnGIKNXEcuyEwV+d7GNge5UvmK987vGLm3x
K1DOvbWJfPBmEVjO4cEpvj7f8teB4sSGGtL3jepm0huWnGWiI/CqVWmGSwKVAIjg5XgHatIfrT1r
O/D2h8NRnumKaHbyxicTGLEMYC30di/Pa4isd/7axVDHegBdrTKJYXuAj0hMvdpyWvFaTqNfkjBL
zF3SgiWjPfrAQZIBq94YPXZ81tqyYl3C50x2h3NgZZc/7m+lE2wtK+dBQrhhXApCA5mcL5d11uFf
lfXobOgsfjjZIz6UhG/uVpnFtoOnsZG751rjgtmpjZYR4p+Dqb1ZGhiw88vO+PJnSlAPQKVeHI7E
BfrHQimt2UM5RB9cwmAASbGdi0u9yauDTCxwymv6ASMj49rP8wcYyGbJPtHQCfSeUdhEGd9iEPqZ
UbTgu4d/emVgMKPRifHJhjnmIovGdjhVnCh42RjqWlpCu/OT4SuCwbBHDcSbLFpMha5q4Cyobi0L
9Ant8WM+Bf9dVwmagfXzdrf/dx9a1JQ77wNuwg3ysWiNUvGnddr3V6YHyovEOpWhl2qJtoQ1uBZI
s0v/5DAhxDiVcxqlRTpol5aCHD3AqfszzGK3xQhirAimAZmzQaudxRaitdjdXrBdFSZVsrIa/GFf
N1Gr6Ywz2crMOKd7zbo7VPfysHpwRcaQSKjPgq/ctvBV2pgl+nYDkVgnJ6+Pwyot49mbPqjcizz0
V+msZiR14ZyS8o1Bohv7WnxFalpNch4VvmO2WgLswOmD53X3SMWeDW1zIYdKSUcH2il1/zYc8Lh8
+f98p5AFzHpfLuFskZHMs/JyVf1VteeCvggrgTbRblibEaEsaBxnBLB5G2xEBrX1Hw70wYPO7ZLT
5WjpXU91yr5cfDmqgp+WIEMCJITcQ/NG9p60x26rXcaaAiN0laa6effJenLLvQnhyYhDgg+RAaHC
Gs61wx0OO/v4pswm5bbSyhtvuZgFxpBLGfuja3bUDS51lI08IBhcjYUVXo3UDNK0Xyp0ZmfhQFib
X8BtjtcE0un5a64fkMMiXAl9IzDu2CylEoXQ3X8mUd2aufuoOp7kqNKQW35wWiXugKLoW9uhGbp6
R/4lGBY0H9FjCOluKA8XP+48ZMQGAw+BiZ13wBXtEFKSy8n+t1XRxdZoyTsTXBWV5bUMwX+S7Hg6
TESwNEZ9nTVNrS07mg+TLjc+wPV38LX+fDdUjWpa97lhaadZnFNPHbemNBAgsD2jcODC2XgfZr0n
JcQK9aYR+Buy288zYJkU+qeV3Yene2l0I8UYbUKw+qs761zedkj0zI3k+DdsHWUL1/8OEPlFPNgF
20glN1kGvSohCIS/wcmwYwXcelnTkgGWS+nQmhsH7d9XYmWf89sxe/l+5X1mtkK8u/iPksKQ347r
vBqUI3EE6MWN7Z1mFW3vedaaeVGqf1QLvNtSVSuEgVO+n5uslH8CSRo6UPwCiw18WzOl66lRybub
wfiwdCpj4t1ff84kV7Cmtk01n9eRjRS3iQTxJRG5BXbuk8WZaaUQBi760jOtt7V6HNRwJTENOB+r
QPZfa86YU9SH3gnBjB0J2tqnz8OA6xVAHcdOT8xRt1MXjjGSbtG186Yo48XRIkstAxHwwq9XnW/L
OIS+T9dfG7cxoj1TUztPoxp1lgHZqKHkJ0SDWyy/4WsofAICoozMjxuiHYzoOoKdKMKOU7rLnRrt
6kAQP7e4onilQhPkfnmE2YA9BnPXBteAuMumjEUcePANvXeKimuE+/oEhNJAuciE1oBINA1bOPUr
S2ZsZ2lMUVMWC4H3BUs5S1vmkT6mO2+PM9mLN7I2Vu0Ocw4KZ8uXg2Tgt45N5amVB6vpcFYd+hfL
LVk6KCRSqMmgujJZClL+fT4To+vCJZpMcWxRRAbJHN7PpzWSgm39UNrOiud4eyz9p1j52tIE7GS5
n/fFvVuUE+bKywtUcfQJDbzKSWftYuaXrTD+ZCKPdBZuzKkr3+qMhkCqLfDoVR9BZgipkLTvJF/F
2biISIGozc3tbuGX6wlfGsq8CsA8U2V5OKI44LJAZTPMhhqky0K8HPtuOgZttRh9vJMF9QWszmUV
8aNlPCWGqeuEEn68E3cT9QbWkKkvkAvdJHS1gPuaeFLXRK8EDmgaPxw96dinXV7ShGhnn958rtQs
ceCxUyH48zLvbiy0Ear2yqF+e15srEL8xhjwSmyTVVptWRV1XaVqjqgEvs5jJXKkzrBouBG69mtP
54nAsX7waPElNjM+2eiXD/P5bWWfF3itp4LV5pvuv8uX/evbvhwd3tQGJOZ+GRaTThgRNZXDt/Cf
RkT4ShB5QtjSvNl6FI/ovd8gyNpAt1xm2J6MgWgqkSmyowNemNxnZfFpINRjHxe7mjMYpL5381Yv
NYdNb1mi/OiMpm1e9ZdV4isma4Zhadz2YxivKuSHS5WEOvzddLj55d4+hLXUJwNnr1DAReb9wHJR
w300/Rga1Z6v0eg5X30z8YocFRXn1dv+AUa9YNZTnOIBd8KyWryeTHc74INb1g8RTiWtcignmEyo
JFtEy3vI0PmGY98iBjvjtb6gZb67qcyoyap1gqh2dJovi4CepC7rjBwXUobYpz8gsVgYpWC8CT/e
SVOVVhx7K9E88dISshCZNxE1uGsER2syB8/+dqTnw7ie4wVbAQczvwMT3LSN16lyCBUHzUU9VtSy
g10RY7SWdflknd68k0orw7uFlsNPGrKYP6BhNbSyy2tKIQNIXRSoDERFrTBxjouVRgThLSiuu60X
Ck72NT7YzaNCK5IHGOugoXCHH8Wb8aRl5TCwajovk6N80Gf1YKFPQciQmt6XZP739zf4uqLNwsm1
ON4P/vkAZ6vNXES11lPmII07w42bHVOhBWjKKFbl0LiqIU4xLx+NT+AALHiCSsCn0R5QlCIV97PG
NFZeg4+gZ5NZH2vWHGm0Wxx4EWkemarilQOY2bRm1UVoZ1HVkp5osecEBOopaHnc4DnfKkJHw3ow
+JjsK7/+17heF/Jb0uzEfAIWaTGqnLz9utrZztvANzmccP/1bHoc7QP4HGI7617RsCT9r2yB+34W
RgAPEidfrQ6e+DaYuccrftAfaF7HoK+o42sqLen53dtEJ70XCjnHp29p1ge7THd/18Ocsh/yHawk
2GJcuCWbozWc87rDvpIBfcTWU43ZpLyztUlj84v7HmLD73AelawNRBOHynMvthm+T2Fd16gI2/s1
JYx98BLqC/hPZf9KRPqMQE0Z+EAykjtu/qHMaZU2EJlluRvudYWACIY6RzWahS12pJouvjkZHlYO
o2G5i2VBHcE/F+avrYjUHH1QqIJHGlNkQgj9l5BLHedG9yReOr52voSuI2LnOwUDbaTY+pZ9pbfh
MhDnp2ePzhCnKf4sI4yhMCtLehi8vqvZpZjeO2H3DFE3M9o9lTWMg5xN3354eCtfUjB3VuJc9Udh
1ogk1ox49zV5tLAgjT+0EAwcr4g4uBGiPaHpQqCMG5TVoQAiIgfUqokryfL7IXbq+BpWBUDelhCl
Z2xk0YEjb+f9/DLkyjaYPuPngZRL1NoCLjeshT0sFd+eJbEafSVzeC3MHVKwfy7dnSN8csyg37mG
511Z6cw9XVtlS3Gb06CtesQRX4kSnyTNfGVO8Z3UcLdW+wDiFTPgsGIJw7/L4QwXP8LFYjAOkGDY
A0eHz0bjJIDYvH1DBjN/ShqRgNmbLA7LR5lOHP9ps7LifYxqIP1oNp5jkiCtkX/qLzS0aIXR4vnX
WuhOkdYj2Vfy6Rkt+aZiJ+Di6svmDM+pbmtU7JYkSiC+1k8d+A5s8lEyAmL2GBesqgha9zFmiF5b
0wa5V7KyTHSNTnnq9MntIb2wxVmCQsgrGlxtRoHd7+f9JugUQVGYNL/RE4K4eka/D5gqU8SA+MiC
Eyd1MeMs2PPYmj5KOpn0HlQSNnTxFyW2I8zJcF3La5ZhbVKrePXdRBVapLyve9/44czXVyh9Vy1H
wArKjoYIbzfi/lhlyRo67cNAFgkRFCfBzF45sasAD2jgG7y31JTftY7ImJhSrIYyDfUoX9mzLuUm
nxH6KiqqvryxCxwVPhhbyhnWxxR+2MoIC4OUk1hO9+7LoUuMWQEs7yJYk5Ua0ebUwM/PP5SbCx0a
tSWCd32Rgu+8HeFRT77EYC8hbXyr+ZzPvem6IYDoBLqAFPtJRULcEb3Eap76knbRwz7csKioHHXu
cQSgDhEF8BJK5/Y5duJK582rF+EhqjbBUmN4R7yw+4lFGVXn5uEU8Ryhjrng/2/lkW8NVMjpfXFB
RceAX9LvIoqXY2Rch+6eIVwOZM90g/3FalqsTJLKZhUXeg5sZ3WfhKbaWq1PZLC5q974FRcxtjHZ
QKfPkWBfyPNK4P4Y9xjx9ptKlKV8iRTWz1irgKxzRwwQqd4IrYAFFqO4dzLqUKGRByhgD8eCethO
OWVee7Set1g0AJwhwKeQXl2Z4ie9HBsoZx1oBGicYZOQLEYtCwaK7fo9UQjueTn9FaGe6b4laz54
ElFGByZ4rS2NjPCkKznj+RQMfiNmCPWXBzBfeCcZgsokTvxbgwWrXS0TuvHnG2VvJcbG/oj1RgCT
aVUWGkiPcMAyp8aolykDLJImppYR6JWeJAY5tqtHamMNzHQH4Aw/dEyOzTSDHtTSXLWiUQSkn8Hr
sgWLmDE1+2sPOoUWy9kZQxlhzUL6O8MMUAr44tL9bFD5Sgru668XtbhitDe2t1Inn3JQ/kyl/Dy+
gxySSIVFkF2DOiK3NnqiRx4+LOb3goX/+8PdWollw8IoRNFBqCotUATic7cCRW6Q3I3UEkjOsKiD
ewKx7P+JqQ8B+gtKAesl20MCX0PXC7csDKxJd7iI97bccZOQOXuoob2k3WgXlQkcvHSCb1f02OQP
2bx/6TQ61R62TAyiqUp/uRFOYeVyBEaYR7/dqDXS6qYSIO7IwuLctua1QH4FPkLohq+x70tyFLhJ
Gg8c6ot1W/Ys7O6BkLz/kOXyZAvqpo/2MlVvjmWF6f5TTKvQEKN+gjFrSv0flsDB/4Ar5DLTvL+D
/WtsKapLJfc7tYrAyiuwNsQK7TuY6/fQ2hnqW5FwquIfU64KhCJFjpC0jShqD2kBmEBiJja/DDUG
rzfMN87ZBej2HoAUuybrlt4X8wkHN+L3hA+ns+LPyP7odY/WSAlo7uA9KRqeSKuAch0oKhKU2HYv
6MueL27nQIopweORRSGG3+cM1KGxmGk49JDgPIDGIxT1YO+fTBiDXJWmDl0pvgPW5AooakIxwtGW
+On9Wc2UFVHRnM7ws12sfHgk7eDCFGgUWkKhgo2oaivur3IGctl5WgL/0zIUTFbxAuqXQV9uNAsg
ovZh5IszXsE9ZjEfqRnk9Jvm+b6I0dUIo/AS+dKdfj/oq4EZ0DFXilbe49xDTPJR9iVAHCUag0RM
zwqimD6FCMIWAowseMpwqpvcgA8+pQDukaxk+1YclqHTc1+PGjdeP1QR09JBxoRxPesgRVcGo4LA
/0raowwXtrr1Jm6Rt+E3iyyppYnL1WMr0dSPZY8chTyFqovrQSKdxanNrAABqNCiZESeMyNs5yct
1+D8vVOigp4OQ9dWAl6xSDOmlpODRDRpFQpeSnHW2elqzXdKzV0ghYpyMde5d83Yyz4YqwO14M4B
MFuqRgziJPmHueN0Ki9u5n5ntgheW7qSr5Zuzq2L+zRKzej9bXxNU0jT9ksJUpr1FmtJkE0J875u
lpMEVZIQttKid5JI/3IoCouHlaJdD/vMY+THiO/GZROEWdxai/RS1y86ClLAASvdZBNijGniFzVN
0gdiGagV+lV+U23/s8IQGvYnJ39NqI5C34hDDxyE0F777QawOrxHk2jA9xlGx1un2ULwgjvLfe7P
jXyn3blVzG2fwRtf6s+vtoqG/Ht/K1JCEYIXXXcdf+Oj2rQ9FIoiMAiitr090ypvWN4FVL4loSWT
fduSb/dZLrlYZYRXJdsw3ZKwYUWTkr9ZGo+MO02EWXnCJ+V1Zg3k8vL34DtgVHHiEtBuhfiABm4q
sjBXExobYV/MemJC0fRHyhU1szgDkgPF0nEaCln0hSCzMxa5OsbiCdTV9zFh8nZkv/129HgOvFeD
7jJU1G1Z5D2xFfr/bi0YKflqyk0ts196ZnbVsX5ArtVmdH35x41G6dzbYP2EIQ2qb3m8qsWe6GDG
nF2SS/lT8lzlO2caqmUB6SNLKQVbIqotyLFr8oRCRRcJdfvOfQIhlL/frei2ChxOaB6xJ6bXpTvO
P+fSFmrM9Wzb4hPK+kU01yQlEZcuvRtQ3sPrztZ1vmvOIogTJn+7cw5d7uajiDQgQIo+XBD37d1l
hNvlMHIkcEsEXlVpK9lz3X/mCJkgiiYDlPGnWtKOw2ksrbh3tz1gmmxGURkPgstN1yU8gHT7bmz/
qO5OJh5c3wtOhDv83cYgl4zpARQeVWzrvosy1rttb34rdr+2vR8o/ohlDr4Au3kx3K5PTuzQsrXr
46rsbAvzd9F1O+d130T9RFofgarItZtJbAZVIS0gc410xXhsdGo07r8C42nE6ZJlVIn6rq69soFT
8iazstBkLdNZuKwMfC1f0ocBhuQyLUqzEFkFvR+O68/Ly7OeS3XmMT6NNhkng/I9etEa78lfAbKB
rZCihSqw2rHqlWJukcsR43mv7vig6Urb65yMdnQAuBpnphCc2dsIA1jctduAI4zJbdB23YL25Cip
0H8b//HjmmKkywo66YTooPufyw9P/sk1VQ4ULMMzdjzA+BvKj75l4ZFm0OWEcwBZdrQcD1Xw1ZBT
Cr0NK0BvURgA2CeTPLvfRN9t0x/cBwmcRCfnmgcbJuamoU/GCiqwlTlD4Z4vjkEW3PQ2yqe7wg3s
LJfnz8JaJ+0z78KNTueoITxMDnppySYW2teOe4WjEWR8VFokeYMSk6+ltnZeXHneZFjxN2bAzwO3
oE3tPAPMSiS6i9lH37cFPz+f1JEDQtN95zfeJUCO8Q7jftChw4VRggda3inyc218DLAkKg1ong6i
RMzIPI6zqqiwZjaLq40M12dX1/yJM9rM3XoRH4Z4/px/C+2mbO3W95HB8Uqq2+sgZfl8D6a8aHzS
TYFXzKIkbwL2mrDqJWZF7vdCE9rEKdJBqthnV75bvgvjP3ERQExbcmt3ZaW6kPzn0PCTAdE4CkDV
besarBUodICvN+FKVvjySn4B4YkV9+7ejArZty4lggAQ7KcvCIfbp/zGrDsC20bMi0PN/nqfRQeW
69EzbNpyD3nE0pH8WM/NGD3nkfg7couelNQahD57NfZBY6CI2mCAsbCj9ENRcp6i3C0yKpS3KdgD
noVbB6rYKXqc+RrVJ5MN6DSo1jH5kL+2dJBy4AVBETZREOF3QPedZciP21erznc7xnPP6Z4gTowu
6aamuZNbHZaMbIaMdrGKxErYnF8I1PuI/Q560bC1gY2gD+KD2qNMbmqu7uWO/aMgkWH2BQ49w7r5
/K4MwNUl73+wK5Ejf9joGGMU/A2Hue0pWrXPLqW0KeauFhmD3HHiqSWYBCqHUWG6CFRXH+b/DPzR
B//jcItahAdQaaCEUM0T0w4jvEt2gqZozCZUvyG/mQkdeswXclEaCRavO2A3K+UpM2KkcQfA162j
ggkrAEdVZsx/2RjL4Yymg6JhDzS6mkMjN3CnYdCHypISmB518nV4ENOTSToNP7L0uCnOQlDgXVtT
N7fqbAc1IyVeEzzxV6Qxg586AhQJLQvCetjcwBm4RVYp2xEhxrBrzl37q9nt9tAxaGxj+EeDEJKo
rflcwCRieAzgiUQixgxIJE75aDY2HWohacG1f7r7G6DgSB6nL+Dlw6u/tZI+trqrMNdNJ24Qt1wH
g5u8hIj81nYAVcI//U+UFsQITz/Ajb4jgwUcUfT9NzpVbkpq9BrR0YXjST77zURZ8nbfHW5ygrG3
uZQ2Tp5+rm7yqq1YJGdo4djN6sKBftBfv7l3YwZdRSVh/l4XQPUWr0hp20lAYs26sYw8e1Uip3Vz
jvxE2mL4PkxTzzGdLJl7DE0rTbEHoVfwJ2Sq0tuuI1pGL3h4X/t66mpbR8SWoTdc8dJJMczgE3ML
Ir8UeWwMnXqfS+4EQsX3b+63pE1FhGlKBgUuAb0co1gQttq/sv+oDaHLLdBavLKbJcZkmY2MbnP4
IAigv6NU0VBL4lAiuLklE2KC3RdltqBARoajRYteMl1MYv/4sGFIfNtcMI6exSvTH2rgn9HSVfvN
jLAZg/n00HDxLvEUGhKdjOiN+fK5+gOu/hrHNFTKbTYIBvGoOlJCwQox/zucuFqyKf8ZutdiTZXH
mbSH7NcMZtV+2fh518wBcKgjQhM3Cn8wi16358w1VnY/JatPhpZsa9bJPXEmUJSyyx7MNf1KB8Uz
1Pc1YvsP7JVvub8kzFHP0v9VRBY15J0JQAuVk5a9pUWFFNFchdOAoqJ3uE90vWc3iJnpYS2kBxJp
Zm+LgCkXRt+XzG/5DJOuTnNJERY5OIKJYT+y/AqKfZXDw1RWx4izYLHBaB0760gLawjV6lIhmKs+
S55UmKv+uhOAdwbBcJh1Qk3TOpX7TNhhtiJJ2GYT2DpTg7ey8JQTtVf7eE4t+DF6Yu0IYlRIVJ7A
QkoCANUkqiDKOIn1CSwT11/DtKEr+PcphxQPeJxLrdrS5TzsnBxFQWPX+8af4/XN2wJRMltmT0h3
oawKdhV/ICmCyX4cjOTjdiYhm8wK7kRYu1GSGgMTlGcN942fcVBJ/wgEsrEfiWL4ym7k6tX40m9D
dBgqlmO1Fco1iimoiPsf1ZdFkkqnWYJJlrF5tmKxGyEYLikZBIZMmYAERDjc3ItIHgyOLBl3fQEt
xFCm7SEzbOTRrjbCrxekEVqa/aAJK/aZGiLzTPuOhO1GLpFZjsBU5i8SDte+J9o1A4oxLnBS8diD
OhiMZhkvxJAnub90f++PUxLRRkU5KOibT7igEr2wm3zPadAa9POLMLEhuV33uVJS1PxjaxoAb5+I
kcMHpcjP7oHNhdSXi6cACc+vTbir13jVxLAySmfxKPs9cjpuntlZlj3fWqHkd0SVyCk2CY1JoNQy
VHvlLzEGv04dfZDogiBu5/C6ZAkpY7njcIsdqQ79UjM15l2u/pVwiExrHKxfnYFyZPJFXqw4/Ab+
SOKd2W3RTLJMsZLle9cjfhNu/BCGBz4p1Kg47kHaLKvhzsZNNlr6EZizHkpxzOFGM+9CvTIluCMS
ispqfkRnuYLRUrNP71rRG6wRLK4NY8TyvEoX84ONw/9idjNu1jscsYFPdStGqLj3C1SikLzN8Lpi
oYnR7MI9wNs9hNH2v1TLKfeOuPcec8a59HwFh0QylnMEqaNfy1mwrNxBWun/C0h3vaMIfRkvEkZ2
WQTOCfUk6/72OXcdisYNDyEpJEyQROJGvTe8ht3OXn7R4zqdjEigd7J6KZ8r3Zba+WqyJ+iIsfNo
6rlOM+4/phDYMkMzHsmpMbviUlr16rkT/L39n+mtUS+hjtEl0PrfR+BKn4b2LhQKfjBXqz2ULHgi
4JBCJoFIYHM+ixBg6FUPhGBD8j99Roir2XPJ2qSF89wnLk1z6pFzpprrr2rB3FE7g1zt9ff0MIIE
+SsnXqsF2sWkKUvyOcmy3kPr5ia3sSl1KYlMTi0E5N7FRF1Obpz/y4/H9n0TgkT1R3zEsWb4wUXZ
vkl0CIp9auGwF0UPvSLeBSiuan92eAXayxcC1kuQh7yEZy8WZwZHjdVvGY5cM8rD9eEuOsfyEWAg
+w8353AvKC4UEMgWf249kkTHgHjcTiIMsfDJxhuZ9EIWofOQmxNZpLF8Kr2s8HQQKs9aQmX+337p
aeUu8OOzBm0IMzv++k8R7kCaVF18gmSvsJXdKfji/nH0E0/YCPUUZQdOPtRWA/Y7LvM2UQZlH4m/
n87D9FINwG9oiko7Z1yTht4wLayqYpZNB7s6D1PSCh3UmLjLjL2wP8ex0pleURwjEai2rqsoeGaA
wDssFmdH3Yj5ENOrfT8+U2rhli7nX5KZySzLK7vHHPOVpEOIPYR+FQSiZR5LKcz+Ju8IyDSDoabJ
Wmr2G2gi01mEQzqEnR4Ixh8PSNWcpST228/8RrmcXmiU8VE5Czia6rMtGaptjWciuvK/kh6YHSMQ
rnYyhm6NLj6SI56XclwfnWkYFRmU9VH9LKh0P3rLntxL77W5tbMOs45jiDwCNE6hS5XwrwssMpyT
usd9TbIPFNoBelL3o8ExgZEMdeDYpIEXi1k7O1vWi5eOgGg4Ju0EDiiYXEvCZN3SLy12dVYHBxWt
gj5Qh67obrQV/leBbiq/dG5EWSJGF5nEFRDkj1q+BTEHGaCbgySWOXVCjWmvO+Tx8tlo4nIIfHsP
GNM9Hm7jVJgc1tQhuwGb6bKwAyFMTIXDA50LDwyWrl6c8jbMaUyVWaNIdahfHMZSBPRWRjlntkn2
mvuHOkZi9TebA2hOchiDwlR0+0s6iqv2a83imJNavZdGwuVn8pCsTS+dtWZE4BRcY2FhPzc/hEer
E524kzeV237n8zXN+G2VVpd/x7HGmoj6d1b6HSQKxVR0uL7CrhngkuLZmDc5YHmJm8QfDV5ggs2m
5BW6XUgYpFF4EBcGTJofDKPA8XoZ3JTjj/i8csmLq9kTSMm4Mbo3HlBUSs/Al8wqN7iG3GU76Sc2
PlbmKrCIMsOXcRV9E5Gx6AodJLWVyKsqLjiUkJZXqsoOIy/r+eIKUw9BASDRZ2I744lrohfqg78j
xOr8yBqcKAcKwylVgmjd2paQj1+Nrb5nuoWslSmt/PhuRskTWo1LTTIfngJtoYWa+jSp7YhgcmrH
SDoEms4Taa1JFCtsCL0lh32WUCQ5ZTnh1r7oZHIuZQpX2ZPoa9rJjXuh7keCYp3aXJeueQXOiFWp
IGr+U9gj8/sOKxzcP6WkHaxgeo5BYc4kWmVYYmf1eK/4GnnpqR00mxdAFOmBM+uWyQe2Wye6wCpS
iJ4FRPvpKOJIpersFH4GDFYaVECDNmvegTgs3rUCOpHjWg15y+DBxZeLnrhGk54E2BVQ6xEHQg7w
nntVkL0jKLMfIjwUx9HG57QUC04WG2N2d6ljprQSNFNi7FW1r1afVVm1Laq2kj/tFvFo2Y5wOZ9I
+xLUxyxr9+5EM19SzeTFgcTvXOOzlnea1xZ4ZmCZyHLkhO22RJuEmWTqRb4Nti+/8xiRC5LQNNJ+
5Cjp6zIB+v6IiB80Mec7eycAfnpAXtSRhrg1QUKrqkMwFcq/nInZt7HjIew4jAlyG1bR9Krzz6Xx
oV6NOT1s/JCZte/c/xhY4VJ9GPoE//ihAo7SIhKHDzmaPnC6NBsQXOa28Fr2HzePb7BUHFwQXk5N
e9ZBlbo49mZgTeRXeSeqCMGvrO7/kzwj1oNVozMRtPOjD82sFY/zkjaVEJOljV2/qB3fhoHf1xUr
V/RYMxHiudJStLyz97grh/GwUGVKEmatLfRK3oC3YMJD3Mr1GU9EG/+3UZN7eRhjqv0aJmNGPxym
u+e+aTb1xwZKbXg5raT2MZjSEWn42D1uEDdu1+Um/r9BCy1Da4KhuGxJlQ2e/q1Ok94Yx3D3GY2S
cBV/JOlfnvQqxZr3p7aNE8k4EGIjp8EVrjpu5yik+4YfWq++ARYPmiCEQoTOWX3FhXWEeqT2A5/i
GARG62Fn49ZP7/kyJUwH3hCvZYBcHqjEo7dvttHM23hm+kLvitMB87rF27AkPIaqlTa5qxc+6Hoy
n5yeJ3YkxaeDMyrmm/S1XVM5gNfSH1OtHUc67zbDAQ/ObFlaPH2PA3kQNyX65cXnB88VWReE3JLv
nBGtttw6D6rmVbUu8vDqVFd1y7PbY7Qno6sIUX4zdaggc0qP6agWqMTlSFKuVcDTHZPL4I72xnez
pLxzjnNuDaUANZMF8k51Sw7Qt8ldp4MIcXggklDSrnB2LwO/CgYrMLh8WL1GtrF7CUMyObATVVcp
D32UVCYeH6ycRrwDxytZJWV8Kaa3hvDwMM/E0lYiB/DTv2kWwst1JKkBkIveBM4i6uBrpfLFRo0P
sT0QeAt6atJkvo/AIcCFeopV/DQrC0jqrJuIy8sIqavIvti9VgLsTc93TLkvbFwKMQkuQa9K3nlo
g1igR3BOuc1Lz51m5lcwuw06SrQWadJ0VKPiXV2RU9b+SdBqsLLYrB5sTRY3GdEQhcsNmFvO39qo
JPLrePNCJZObGnRwZ8FE7x4vrPpMPb034UrN/IkSrb6AKaisd8G7lWIBD7qQDnOebTm6pbJmJd8j
nRKOwUAstSwCG6cHTrBWcghXoFUDAkkMwca24bWN+J9/PaO59/ZZo4obkurdg4Aushw8aXox0v5q
6b5KBT88lsxktCbZjkcfJHmCBhnF5ZEERDmu/pm0z6dNWo/9wa0waV/bxrPeQy30MVt8ucYRz/EU
DGrlmvGx3m/uauRTvU1HSJN4rOtdIUAeJ/4iOxoEsA8lG2V3v1a0Ci2xMvgnh4VqbU4L5wUdI92l
tGT03tDMVzCkcIZp4ZW/3xvfnp/k1ALvWPqgoGvSk/A4EwtU5RNxN/g21ucVaLJzdNBHvzNtR39Y
PLXfEaY/r1YfKKAjaBBcZH02iEZlt/gfxUv+X+ifWqYW5nNV8k2AzmFcVzy3PcNJRbRBlUEf7ogG
gEsqtDj0vzFz3eT0QgWewMn+2Br5ETBchYQ9gRfxgU/YfEx5k0xJcft62ooNYlbU0QIuXJvOPZXa
MEiTVDX2vFBfkictdJZtX0Oggw9HHU1ht2WUXj7uyQLXsvcO5UzPz9Up2Mk9e5mVLlJegSAgfNWJ
ILdvWnYeIYh9eEsVt7E0TU5ZNQLYqLApq32CshWY2o/cV0ulWDmJRSP5v0MkY/eAWMjn7dirfIo3
+FrwJ75qzkocf862xLhWMYTcJuDWx4YlQFYKAg1El96C6W4HSyaq0aT8gNl1Ksty6CTllLdkL0+K
XWHH9rEuAePFZHWsWrh18sCD66rpeg9ARA+R2ezcosPA/TwtdAtye8VmKzFW/v1H1MjcwTpXxHe5
kiiyXDijSubGxa9yrNVTf2Hix/t/G0u1E3TrPcihh5sjL4cu/UdqKfIHpoQ6An6kwz+e5wM0Kuch
BeymWsJ1FIOqlsOhoZ48h9Zqsk19eaS+7uMPSAtGZQVjy6xHbTQNpvYXBOqosPHMw/7E4iRZas0x
wsaF5xbaRWNSdGbvIJdAM8UaEXtsr0Rmpokp9+Lelw/mBAm9onmakzcsm1HWr3SEvkKBQcUrqWX+
6m0aT4UcuPcxhDsrIk+1PjqS0IvC2ra3IXg//HEVOa2dtYE6AnVsixPkVMo5YqZ07rQfNzhOHA8j
e4CuJiDvtn8SO85jsHgjEUgr2n1u7/pL2xUCWT7atugJUQGo26SdaZ/L/BFqQi62Bt5nsQV/jmso
qJBKgxcnKxAa8sS7THNebnfIVmL8vyc6deg4s90l0QE8BOlJLOmxO6Oe9dwGit4/s3zmsN19w3O2
kySYmVZo8EexPmunKPhr8hCxJLFKhiyfu5ckB5ZrGcnef+fKL8Z5n2PLZhr3q7blQxROE0yEovsW
neb4QPDK7wu4QtweuyS7NhExv9ywG2h0rvENA/YsRXYDDuyx86zZZLSLFbiN/7wLZiJjem6EhjDt
T47Bsqlk1HZsGV6kG6gNTH1Th5TFq65Nx30tVRIgSC5GDXk5hXumbx4fS61qD3snGc9qS70jdugE
Tff5QYycpFo+KOgg6aKDY1oWasJqPZphk14rus0kF1/8ZH8os0hHGEcOL3kiMw/PkuCrn07zE8oM
smvVSxsiMMs71NKBgcSHdLfz/hSFOVzBCxEZoHdpmuZVkq4RqmgHb3d+8ion+t/h+Wp1+3QrsXOr
usC+K07AsUmYM4Xs2syvHjMRpgUjijEcbyJxHVxiunmkvDpcIlOuqx+BfprMto/2/kyPIHZI2FWk
xwdRHystbOIl1Qgk5Q4nyxiNbjfvnxv3r/YVvSm5K76DRjwZHzOV02Prq4D8FoUrZ7gcCQrf8PMU
qlhqs9oct/eUUvUlZYxXQDmOGpLkdMbYOLJ7AdDNJYNIuHOZzW529X02iqxR6irLnVNtxIFRVhAu
Yt1whZfQ0dQTbLbWOz6WYhyK+bsPcV5BieCtNfEJZfxhtHkIA8471hAKhe8VXqzxsGBvc7SwHQNF
M7fqBG5nfvVG0P75AdReOeAF6ii3aMKr/0jSE2lRYtzvk3fKGJbRNUqEBykhoqIWWXNUbtjM6CmL
9sHQqiCiFgFuOpdHFx9WUkRPUL76xTx5e7FwPa8kCFdo14rZ/mhDsg3h/jYD+qfTjMdVGBk9K+Ad
1YXszP8df1rygINaKtNcI9/oen9vZfWG3EhF2j9IdCjMXiry4i0X7Pav+aL60qZAPQ4ASB+h7HY7
YBawi4fO/1D2wedQzPqRUImnIgvKmvQdntZIjeEX4wFqmi/YPDPk1Il5qLwscu9rrf2OSmvHiqMD
XIp3IixlNKOX35I/FR+3UtSHkOYJ8pPkcItpYmifooJiRBdWwE6aT7RCe83brZEgPVh7pILJcyn3
DMB9umqvyW6tf5keWdh6LEIvIG7dANATL46M1jlY3Vt0fElc+vPnt37xa36xb6DZNd9g7yZ5vsHz
7XRMqZyCJcNDfmW4ogu1jvULI1AaYsy28/gHC0SRTr4aYeyxrfGe0cFHmtCd9QXxBctmhlRjpgRb
au37T1tYicvolCi1YvylSp38ZRiqh3wi1RnQqgHFS4VJtJTVsqzE47xhZmo/JIEkNQlGNzMyQgSP
/E7EMxVsVHh0sPGTmhzcxBz6bCeEy+Yu+Z9pMKWXk3sCZKGZTDVmOuGQ7OeRmPcMP3Ur5Lp73WdD
s28Kun4qDokKU79pVfAVt2whQ3cRCcmnWvRCcwtGET+aHA8uTrXJYO+hLnVSXk2GmiivFkkIkZp2
82NFEdUSORu2q+S/pI9cHMs/sH+iFzv4ENP4pQVBOSslkXI1iSoHrWEg30K7DxoqqdhgdR3SqBOx
YHgnwAAaViCALZ+nJoBUb+9vjnjGPH+f74Y6rithdvd2U8fxdYkfjjmiECbtPX907cQSHKOx38yb
YKbzOrOTVgv8gxnYq0tyrgoCs52LS0IRYQ68AWhvK7v5N+zlTp8Ca05b21vMaA4Y4TYWPxEuThYu
rID4txagLiUyCYcsp6AG/e6tamH4ofDiiU6w6GYMsOOABX/wKROmXPxpcV66q1ebDrHaJuKYfQax
tV7Ztuy2PSlhMF0FSZR5dWUmx2TfZKCfndiCrdmaXVuTygSLRDiuk4Ek3tpC54PfqroAagjBJ5Zh
CqnoEuaB3Z1/vOhKpg6pkhV4nkXre8athDC52lZKFJE6zOemN/YvQItN3szLIxD4WfdXo5WWAYtG
cUWfsKVTiDud868giJmL5Try2cDBsaPu7pf7xEWEIk9HB1aLz72glodu5LwZLWsqC/QkTU1wycZ0
q6uBdKMOiqcowmt6ta7oBwlU26jyLbG1IuuNvZGs+pqN4/P5ozuzpyPPll79mVcSlaxbaJ0ueB6b
S8CRBXGJPSoss1MH+lN12niMjrkeE62J5qxukAT4iOsqyMIr1Pi+z5RPQf8R0a8MqtLg9vvdIEfE
KjasiBEX6zVeypE/Jm1ZgMzkg6MumYB4EhZS2nTTdBtZzh5kIgn7U0C+U3sNHCp3UB1G3FiHz1lq
LTtSG9aAavYbwUpX2vXOlcaeZpQIADE/WYcX9o3ub0IpdHYZFEXtzVL5xjQUvqmkZfJALWwZGozk
AG8ihuxk6tzyoaDVQ71cP1qK5gBPsJqPSRbkipThCxP/ZszVUNzHwv0176QkMtwNKa7ZXGWbLiKM
LtKjVOMZ9OaUmXY514NbVJbCu68tHzLi8sFPBGYtXzZ4GaeBWSAmgk3bMSZTfry+0sEIfoQaWujN
Zl/nezZwAvaO9NX48QdU/6TAm6Mt1pBvH0ufFj0U0RGp+vfssAlOSAbvE7Bl3UZ+ujLgve5W38TU
6jCZ03Db91GyJk9MG/jW+NLkhMwUO6L3QtXOnojWEvCfJ63KqKW6IktUYQTUn8Rv9kyOmED2xVQU
RSO5dvTCszk8dyvOt8okFI/eOi6luBPCj4UKB0RaYU7D0T+GYhULESBwnLvuM6h9rtnKq9TpU4kG
5NEn5dPkc7pDC2mkItyj/IPXdfgIhWkfhirjrqjoLWGntf2sT9dVhhyGVmONk9qWvJNqNBH7TSnx
/r7zQ8fieYxMpWEmWXBCFwmefi3mu5xbRY683Y6OLpNAh5er7oRn8moE4Llh3i8LAMQws6vxtdwb
cRCu3RdXDMZsvTF2EZhvhJkeE+9I0Be2uulUFqNBFNKAa8SywzsNyHgqXBH+4YtlqvbzCWE3go0o
apPJHNFJpCwbZDeDV2m+vXquIQgP53gGS9CH2+08ccplOrNgUdatDa/OqtsEKiv9oa/Ys56EtdqT
RQZfqEJPUmkFHyxS4AIEtAmJia/2Cq5G9aBiE/NzTqOs5I5+f/pr3423uvSLVe2LP7D8m4urjV7T
LbYMsoT8YbNawgxDSAjlsCl62VNapy7rAlBolZKvLK1JmDBvWG3oqrkj9/FVU3HB8H5v+xh5HHAf
syzHDr5ku4XRHZrieDe4lCCr2iNPqxqk+T0kjlXRxWaxJU6OdRJB0/wquXij5om9+iCVn5AleDgH
AFiBuW1JAp9Y9Ph+zXXw5pFAVbTIa3zPAr4fiydeZ3ijLsc1fJ9QaO1XlBDuvTKW3//+1J8+0b9x
y9JqwO4aaLRYQHE8XtYfSBhsJ8WKCwt1vIuK02f07RfFlytSGkCvBNuLLJlWze6RUcbEHfqsQEsz
aAC5q1kRjE4N6Xc7Qef8iVXPBFdPjBAGsb40DEOjfLOo1HhpCMMvEmE5uS6q4Pn3xSP+v6h33zDy
q2XFHhnyDHEf1P20fzfA8Wc2ZgejA+lrZTdBHrp70k/xkC8qZhvLTLm9u1UBuSZETK2EiTCGkI9K
ljJFd1iPQRnukxKxmJbUr0IODWVKFUCrwY564yr+6Z7rLp0TQNTQW8788I4sRui0QnfrgnBQ7An2
R3xDFlkuYiCzMu50rbwjxOFrYraL+hYdc7OSh0BT+auFMcMXnQOjz9PVALKl5n7G4nIMzUPyrlHO
M5PngomXp74LUh0WJO/cW4NmzcvTDwdCVDcAwkaNJcgDPBTcbiWDWLnvZnqOXE4AJz/vGEPOboIR
G12ihIBAs+eTbr2kf+VyalU8cFjYavVwjACUmj/p1Ap6QRJsH5OLpBPMB8zJf6J18ZIGdbcVcSfj
zRxXaE+dN89ezRejPi7wy+8g+D4utORNBD/XRNn7JnptJ/txbR44WpzzC9RzF6dtg5qW9dTuM4TT
VwEtwfUzAaHJuKxglkWSvO2XdGGq2loGSJeyxASN7t4ujucAONe/km2xbapI51bmEhI97LICeY3d
cqalbiTMDonuYcYdYLGsUAFVe4nsa9VKcN0KiU2JP5zsD4SCENvSYyYGrSVWZZi1AuMj8QQ0Q+TO
2jsMN8pDCYdjzNWlfmmLcS1enx0j0wbTt2aRf/fBXhHrvAc+ezocxZ+7J4UMvtuZZ7jlGAo+MwAz
OO0Cx2KJ3ftXfpuZIScfiCi8c4+cTrlIWyyepdiKh9ZPGfD/H82Fnjuj8ne3a8BMIwLHjuVwx/u+
c7pOlc7dK/01198Izh62zKUvfrlzZf1Xrf0omeLNadJ9HtfwTDew+UR1ToREyUjMleYXcHfksEFl
HbyG+6b1vNJkK+TV18wQQyP+p5Ma6+tXqM2WfPOFod8Q5QrlhI0+LCxa4AU8kww2c/+HqEamxFLf
95Zp6/soNPUolLmRTJzSRU+KL5sII4bHJd3SaBUQ5nmjvGLYbkbGDxUoUaKP3aXzOH/+ACiBMgfD
fOFOppTWtGykqDlI3cyUHtx7ki0Cx8ba4gXN2BfkNBK5/GvXRR19M7LMjsJ/se2oPA0W6Go6qEIS
1XR/6zp62i6Xe93ahasV6IncLraITIYf4ox/4KUxJ0l5s9c1uii91e3sTXTtZcEY/RxK7B35w+x9
RFbeNQNR80d0Vm3JZLizBDcWAdISSNwjZsxQ9Zpr8sxC2KKXWt4hwJ67IcOrCaneFKjQ7BZ7B43R
69tpqKFF5TMNF4lcBPX/FgxxolANFLKwXTPlnTjftfa2e2QXplPA4zimktfMEmHBnpo29nezXPJw
a2ib0A+R19ChRfEpapDhAlf6wD8JA+8Dc6Q2SJTJ5Qc5aoIzjRWpp2kd3DJCL9WgdC/CORM9akhY
uaU3v5eVK0hNMv+w/Q1ramTpxO7fqQ/3cgY69FkUOm3PDONxQ9ah5l3omJ4DIiTJpKkAyoZhY0yg
Ohay6yXMDfRt62sLPHyRh+JTn22/stdH/MrU2Wb0LJNCjrcmjtMkYJG6DOnJefGOZrUp3iCI/QNx
TvqrtJxSeB1qH0FJLPS8PHCheTvoM+ov3AFSpOaBr7NrF8YlGU4sDojkGPu6gTnzT7Eriy1Ij3Ic
+4nh0mQC2RzXZrZTHJzBoIX3rYkKDZMv740aH4xG+ckl/THgBf4rMsqYvW2m0kIVY5bTNGEl0gZG
5lWO8zVurriA6DTK62yWUEP7w1TwGeWxUy98RgSPgw9a3QGslv6SgZZT5V9R58ZGuf7bQ8BsNS62
fROe0Ru2V3KiDV9COAQqOsrCsxUV0sMjO3MnRqRcgcZEylYYqUq8Kl1DXR29kkY/9NEbOJj1DyAm
u/kaQaHoNRwW/41tSgp6kWnumSSwvQ7P/3B+CTvCXMDthwbHpoJv8Uu8PtHKtNMbX/BRsXYYO1vJ
l91Lz1r7ofSZ3i5z3prTMoG/uO187R1A58vCJ3WGD6LwxLVYDRKHWm/fhI/4G2G1a3oqfwFe5c4s
kPN9cIZlPD8weSMQ9+NJHX52QvncHNlGo5bB4v3YHn+p278QvJ7b4XLgl5qzbsn4DAw0OQG/ocvN
DQSV1WMaGI0A11IgibRrfcAxD5ix8mnu8VD/XpED+eRQ7UfdhjZ/mM5S0wT3VlXfj56TsIgzia/q
XAPkksHeWs3/AvnJlo+4mmcKTtMpMb/zYS9sEkfl8M9zwuHVwaBqYu2OgWT36Yed0XQ2FQ5gzZFt
Zbd4cpNMwLEFq6nZggx2kkshIwSu8XQkx7rXf8cNizz10r9wPl7r1c3vhry3SmtBTE54ZoLU9+FU
QsKTgm27Yxk4wIFgd0/KhJ8tc78bdGIlL7tuH2jTCZkNtPF1tzwi94e1oVaa4/9dUCrLvwZ7wZEt
WWn0f343zy7LD7HWxD5LCTm8lcGr7/sHIM8YcyfnkGTS5ahxMsArVf/NOK7K3iAJJm2gt1aUiov7
zD+UfLE61A/Bd7yqxxOZN02DHj2h2pjAivBau/04sObO7Ce79dVctoBXUrOnB0SYTnUPIhMhCglh
kgd0xmmRU59/DHMN2uPO+qYMljDQEdZDWVONiD0N3SBGrlaCl8KyFZZG4SblE2TjZu0AE0UZM0Rq
jGseLqrDqB/vJT7nK8ToGwAVTXqQ2JvIuYmkhAD2YTKeFk/+PVUNXjBgh71RYi2ZODKVYpdQU8BT
pGZ/H4VSO775EAtDL4lv5HpIK+QSvbeFD4wHRhkhLYA/dpIcowyqQtAMXPQUKiJ8JmSURa1ologp
ah8MOo0EWoCIp6ipUZZjiyTTYQPtkI59PWtMW5I34/mp26SgVN17r6hYX394RVvabhRX7vQytVk4
7spvjzkP4S4PPRZDuVyzX88mGSj9CoK+TWqw0G1C1ILDPpCHCsER76nvsEAmzKNxHt0V5+/VGo1X
ENpcsNH+Zb2g5fjIeQmzfc87KkbYBo9OdEO3mwPXkLcjrnel3xxaIiE/21gQ8eBcKev7kGTrUs0F
uIW/PYj/bIYNe6Jtlroa4EeWfCFt8durWdLj0ZdPSsNp5EYARlwrEb/3KE+Dbu3oRMqXvbpoBQYI
9zr6QMbkBl0IHbxzRxvZgv/dJ8zGxUkIvvTgXY0CQOc93uUjrvtsgeCcuxz+QnuG7Gs2ppTTUMb0
Kyy/BrXfqkBXEVJ9DdhG3wIZg4ourIXJgcGwkryNnWC0Yrbo6jk0NFspCl4V5DqpRd/UZH+HcJvo
Rh9lFOjV7mQzWqNm2qpko9goYaWlVoM8ZZC5/lDhF8zMeaP+sDkRDWq5tAuiBLcJuNucLaiBZ9HR
ZVYHy+6KWUsOTPq1E7p+/p6l9sm/irPPBW4d8RJP2cR23OZ6pPaGvU8jRImxg6cON+KMQrLvC4cl
HKXymfjbVTtx0mxPB+k3KUhEVPWZhfrAY1V4w5o4i0eBUTV+hY6uI8EEU6oWGfHt8IjSdPsqUhBY
oLXPoqqPubeUC0tlwnu11EI0mszAN+OGY1Z6o4fLGBbSWStVC/KT1/LwGdYRx/iIxqw9fIH4RBX5
jH056cwKJ8Va294MUb6wZcJkvRlet5XCgyvnr5D14rRNyG/+z2T/T4V0fzQrfL8tG4713aTqcVXD
hMhxkiTFajl+4I+HxL1NyBd6GhKnWhb62lWCTILzqm98TyeL3HYK8VfrWbILiIk/4CoVlU+yJ5Hf
TrG8F2yepn+5HJ37yO6T4F1HWXD75XITn9G4AXDlKj418hJ7MT3d+IBlHARDKA6CmppUWdJcJplB
8CU+19SfGSKVmY2b+izn8b3MXORGR2qTIhS6lbLpunex3egLAeOHeDh1bEA6Zhb6fIAgcmmjATvW
NKVPVIKFoTXJlBpUr2hxdMq4jHMxpam5FA7yiz5uKmxKgLTU/RTklZ2Ftc4XiZCZVOjmB39Ys9F8
Z3oBHO+B1ZnnXeL66FC4JwEwyOnlJWSFCaW1Zunmo8gJ5gVplfoZYSJJ9k+KUQ8Mb1OL7Zqw6/2q
GjS7tm4cgwv3MZh4jb7MESIdaFU98PcMPsWiGiYsUxMrqtxE0+9+wX7HZe6/PH2+9CSfYk7m8NJB
ayCGgJV+QxbS33qihb1f3IZcjUEwpyQgNgj/ObGM6JM921Tn8L1YDvo9KUlr8a6exvhwAYEf+q5V
deS46+4d6m5EOTgKDRkVjtsd2xcsUokQ3jPuZLRk/cHDw+IxsU2UYRYb0YLpfI81C7kPDZB+ph2G
rqQ3qJ8nxZ6c6PFhpfpUSqjsZ+l51izsQMLclVbxoswXy7b8lCIj1oDAn1xNVZDY3a4h6nBPfok+
iI6fDMg6TKljOh+PLrK5jx2UkbQDEg1uLKGbK6RZOUCxsDMa1bA7/v4dk4Uo/lo7HJvJX2gzNgZ/
xpBdH1xKx1PstDSLa74DSUvt7a14/D8NUx4Zi9WRVj544+s+68X4+UtDhOusZdYY2J3sQRO70hzw
v8a4X7ie8GkVBxrmmqnQkHAHaShhfob8q77qlPdTUPQ8CGw3aJokQT3hFhtrKph33CXoP+fvGdET
xlbTiuMQD0dKbLXQ6rs2whDpv7AxTz8VJMjEcSJ0bq49/el5UsGQkDxtBgFG3L06KchPJmPVwxks
9xc29pKM/c46irlhBX97af5QFK5qiW8dwQK9CwiVNhe2plSvJmEMnGutBrSDMp8ZzJjTXdDeIjR9
cHhOsoWkB7eOwAYHBGXCIWVfAi74+a9rR4zs9PTxFytisOj9m8+d0C5QzdEr7lkU5wACp88lw+K+
4Zmm0Luoe4HaRBOXAmqqVV5UCgnd5jZYEdZyFQBJIGVUnVQWEYUF4gji0KBfWxVcDZNC2xvKMlOF
4UuEeFL9R3XDgicT9g4IJDETYZNj2XKf2lObZCk1ImvUlPFg+Qq8LvHx+oBUnRP1HyM3xeyQKOmi
f1HakiKfpbXRW3/ZalqTFxsP9+eUun1hyd3O8QFwSwKwrqqGHBSYVULiuYF7AoMt4S7CcuJzdU5r
sp7K4XyrujVL0q73/PUquWpBzMhOr0ODehabym6hxtElB0jF0VirgP8aylaVpf3wLQeuqfD0cVj5
Dqjt8WoYPM9kEPq7ISlKh/In1pQnNOdx0L4BOW1ET/co6AHyCMEaCqk/wNBQlROGvwMWQDMRL0Hv
V77KfdjClNetrkNhG6XU5B3RVXJ0iiloU3C/DXgJtwtCdKLohvDNQ/Xymjqwv/yNGLK3hfA6v/5u
juuPcIf/lD1mi7WFohDvEjuRj51YeooWwavloqfSzjMr0qq7XsPS5h2MfS48idlsKcDfty5JxUcC
9xMTiR9IynWvwRhkuU7OGe/CBi1bCJKxDJOhZkCgmprS7XBU97PSS1rnJLyhSuLpTISNe5G85C95
DxmwXrEV59k3UkLqd7rdvSfBmgZ+2spFrbVzPq4BJYbTj4joFyg6Qi1mbWCgXQEfiP9UuxMDNTI9
Vy545KtRquv8N2Dvuq2gbyNTPy/6onNqIQ1ftVm0AUiKEyTRvj4cq9gPjOnCWDt7vUcvxbM7Tquo
HqOyJZiVR86sX5EVjly08sB1X1B1h6XkSYk7z6K9VnWqsYmsMac59bWhYK4Vf1vAfTQTo3jpIp+b
jjSXQqa13A+Ca29mOBWlUCm5uigHlVe5SabntDQoKmrbP3TG+w+HpD930O+7Ui7+5xAHlk2mvO7f
7ANAJ9loXbGkg6mE6zM64iteFR4qzRXP4nW+i4YR6XrXpPURvKuVX4j7eZjL54T2AHb+c+uXxhZq
AThCtIZxGZYoLjW6dfMHA1iK+cO9R3OC9n/tDLOCCxarsQXOgAZpVcvtJVjAmgGSxXCWR3DzZJXH
U7ZQ9WaRLPtjlJzxPpJdSF7gK/eLT6c3r3x/ZMH26n737QNXpAvk/mZUWDmYLlrRrqtCBw7PaDGT
p9w/pT91FPeMuu7Rpd9f098fP7/Qql2ls1vQNkAGm56kKm5eQnsyVdjjL4hFMZTpbOECUmVsSQx0
5Ngd/oNEhfAygXhTx1xXzMgeU6oYPxG1rA0Ehi4bn/FAl7DAp2cjwsZuzcWOMm7qEuFcPkMBJF8N
7WdX5GP4elvCWGC6GajJNVzks9QNvc0NHu9Avj2M2bJztFy0dW2n0co3Gks1GG2HxJqm/o08pXev
S83zPJS3BD4cDELSaJRJPdh4IfqYwg4vIzfwdzhL7O7tHOp3RyGoWSlmcfjugMC88iSjLj5r27m3
9fsBNSuVfu+XY2u8zFs74rZdWyRE5DPVGEDlHZVS1GV7Fjak8VknDXkKW6GpqxgwNeamb5Wz0GM5
9vcepziXEORees4Gb9xs2RraFAGtp6RIZo9fWhsXFrN405mbOhUcoMDYbAZdQQvvEAAwVeUc5TYS
lKwpmiw/qY2ccpxMIxIt21lOmh1cAFjsN26Ue4UTVt7dR/F/SKg1sw6iH91xCrXtaF9sEsouKAw5
WTHpfML8mSCKZDi9mFOumI6f19XdDFatP2lrpoxY/vwZEx2dSqU4JHz5sqzUzv2iUYL1fPCXxmV8
qPvvWiTnF55LtGnLspUL2ch7y+xKJiCE3nQ5EK7Xwf0hUeVueFJV28H37HYhC1+XsJXHEavMD907
aQa8yjXdQyzl9lYDeHMHcc3XIDFHzBDKVqvKQh0oH9HNlmMbxnVifTovC9URS+0ExyMu7GVew9PE
TWHXLNPWrpb4i/Kg6sJDIOLDaI62ePfFkatWyS2nG3KUkhHWQ//eq/BKzY7z1Fgb/P1b2HLR2tHk
FdD3MuqcY2vDnUC45tABs4LZFZ4PTXDyj0dKXz2ejEhGdTEx5+/CBkUHzfvm5Zv7sh4is7AY7Sp+
v6j1i+zFeXcthyjaBIR8ldQcuRYsAfAULew+EzYHJJducHS/qB3VC5efBNj+SfREE1uxz6AMRUU0
rectgi6BzklUHg5l5pCJr2qJcMQ6SODUrD1RUlnOaZqIMYPnyriabI/P0Gz2YK08vnmyqWgvZ4Ty
KluHClYE/PfHRj/FzLDVPk0g+wVUM1GoYxWRs+5UDCPlh8ABOUubCDnAc26F0KKbJQKyOZMvfvfr
jaar3BdURaJhXyNmNkrVRY4Uuw4AgJp6+YFTcPWeNgqyoRLuNfFLGPrJyVLQaXTnY+oXLUum+E65
qpiBnH6ntBYu624kqrn+9hMAb8SXQmb8PcgpoMNUJfV0VcivOAowwXn3i3CeYsKyN0EwVcdUurR6
dOucpJzWFv9zjI/Z9wIa5BE/yiVF4cDKFlf2nekv6xKxOZP7W6SgoUb7IbVuAlh9i5oI4vjapfbH
Ee4bF+OtOn8VSuv95CBM91QSOZefX6jSSt4g5mfq6CjT47crhThoj+IOdPRDVmRt0CLG8ce5Dw6X
FlF3Hzs0xxBcubR770HLXE8nTopZfXIWAaaVfO8e5ne0KPGG37wwtS4DODx2GTe3Qx3ZIGX/tjtH
D1Z62r5YLVOP/rSBYhDav/y4iNrHBhTfHEa4kWK0R+yoLJmydn/yWwFnzMBj9PWXAtzPsDq2jtB2
Wu4ePaD3/QzQkFWP9G/+3RGsYrNrCkXu7FeclplZcVTqI3rGjAwurcLraU02aDkt9AgfscY4zikK
CpfhXDFOBW/i0l3n3RUzmfFS0WIV1lbvH0XjkYTzD9alvNL9k97wnW+PuSeDUX13PZDENPZHnntQ
c9xCM0/qfKiet5ZLKm/R2SHWshUThK2i+a9bmcbpBdjZdssu2B7IHAbk6QAKhSJ2n2IPoA0IIE6g
5ZMKlixfmnqzwAEcSRaERRo3s+W7FrasOIEU6jD4oC3RTTHABYVsHlFYQUC4xHSZ9z9TBDRoQPv+
4RTjD/9qrq/0Tl4KcfCvPYYw+eCHqhfh3u3Zau8WkZD2PzUzXWMeDy0xurSONvwtiQW9LwrQfXic
ZFyvIHgFycDrWHuFzDSHQBW66aU2blAuB7gKYbBVz6PKjgCXojLJaY4tDaxKf+gldIBezi6tiV4h
o2f02+222MJVmhF+Fu4zm314gXuS+LMMFt3AmDFQ5nBxTw4LPLyKwF1aebIBvF5fn7VZp0X2Iomz
eunTBAx4hkt7Z9OSSiiAiZNrtYczqmEI/Hi2UgUaT05CecngobpMDsEmLjLmOuVFrUYS7evzVOGd
yK0CBGOjqi6Bny44ww5oA5EiK2CNJVSZeCG/cORI4HDDOh+E+a0pJOaUeVGI6a1rVjcZMfFGenTn
Qb8Ep/szT4msbrqKTmvALvZU0qqa/fpWR3U8WIbndXXeauz/MBJhof6Ze/5JBc7WadwPhSkmANm3
pAYlP7a8LHT+GJGu0D8ssAjaehOkHZ7jZYR9kU5zdAZwW2qzrcTZPtAAszXGSBv6XUZH7NsqnwDt
UoYrIzoZ6MpGy8OAZcdOh12tXcFsp2tVYFUIncYaxNt4P4BZZAxRTjuMvgVlZCJRtwrFVpRMbm3c
CyaGfc36o1cW92Ef343EkHFk6r24V2aqvvK9RmEPllvJDNR9np7GKplgdi6pBCE5m58tVk/rao9p
dy1/UnYhjhrOYLMIVimUoPS0Vsf67iw5b5R729REURP/H5c5kKm3FQWTEkerWYGDfmoWqlTnxjs7
EeN9LR7azZmYlYJiaKTJ1LutMcsXgu3mEPlf/kJqJD2csDInJyQJN8k3oA97RToKVumAk49FHmY6
uasbwkxdSh15+MiuoFjVYdNibxG1N8vLHF/XJ0dKWDiRPV43fld2n7PinUDrNIlow5ESQmFDMczS
ZrGszsBo5fveHZKrjMGwC9sKRc20+O8Ql3GYYoJ5soHfB8GNg4Obva/y2G43quXHjZgr5CG7kpsc
Avj4m+Iy51RQEAf0Oj95iGuvqgOR8MF6RNpP3LxDqqs4FpZThOJ+Gl2U1x6d3yJhKOEzXeTdcsJW
6WbTwn44g6hEXmmTSK6DjLy0uctkLex5TDzRW5hSbQHmOXMvVC2dP6Dyaxk/B4bR4Yasr7nU2fVu
6D4JsTxAlsRX7vm+5gUjBDUE46haSDMnm5g58fC+tTBlJSE6wjlLaFOi4YjakNBclvu8sX5UPASf
N2b4VK8K8YysjXtX1r8ycjtph3vJmYDZTTRAdynqGmqKN1GJwEKb2J9QLkashs+K2qRb7H7dtdeQ
M21om9oDrf2tSfOPkbBGCvQvn6JZSDyNEtva1002B0VqySoQcSFDfmktYCdujULPho+I2u3Kl3en
joyczqMfUK+3U6iHZNc1zX924pe+KvpGkfr5TMe3bK+jttmDyYq13gUk7LMs3grjPS/DIOlM4gK4
oFOCp65vP3MHjAZE367pkFFEcCTXqXuznWWipslagb8MmTrvRmveILG1aM3xuVJrm8gXtxZQ5tig
Hv3iRxmydDOpxovEhd8z45Ulw7ckcMy69ZKPYDJ6meki04KExH+6OsgSaL0VfZPn3P6hhylluMqi
mpdpyvDcsgoZKA8lN3Lcwuwm+arqB7L97AbZ20yeD1r/hC/JVmag7fHnK8I7xHgScc/UzLzqpbYQ
DIKWHZxGNRJYVhletTBYMDyUnI38GsS2jYXmCKFtBc90pi78lAPYKWJv7zgrEiVX8L+5ZXydqhcf
j0OiinoVpEE2K/Z9864penNeGQaJ0i2jxfxacTy8tt3XMMj3UFwgWq3S36x6fSFSaxck8Y/fL6dx
FJ1fG/fDeZ46mkjaHjtCUOE7VIrjfcs+5Y43+Sieq9luBuR5hFo1z/Gp495Ph4rz7cQn92/Sc5r0
+IWnsRQ+9M5quPa2pfN0HEz4vvnDt/rxPJOAawDec/bMatFUBFpmcD1pV6gKT7xgDxxomKt2BqyO
B6XFUTVAuH1jT9qqeCu/sjo2H5dTybCcaKn1CM6kO445IMlcO+chmuYHe3iKVGd+onsGk2BGMKs5
NQ39M1/QrGhSy2m7OtYj/9LRXZHR0PgQqyHj1kT+ie29kTEnL4S6IroHDwssbEyONu9/UXVcctXh
b88ZMG5kr/P+uvcCfGjK+NWcU1UPNDQNH21KWSpE48bueemqGKEkVNvQx/3dR6OGL8Vgc/ujjMLK
DMiJptNmYbiqgmxsLNea0Vi28QVbYM8hLYip9dRaVuI6Giqv/ucjw7p/4XJIh/XGM+7/fYN7zSkF
Ggr3uqeX22G0gK022e3KD9nj00Qb+GuLFsJD62EqFkcayylHux6iozOsWdOtzTSduDxALBn1zwTt
CExikq4gaBWAPRbskrIBjY/xkHAjGOuk6UrDvv8JeFDM0jNmre11dV6Z5vxyE2XqnC/u0D5vy9tN
X7V1uo4iMO9pqKZuqG5V/0OQH2SBJ4kAd7U8CON4WhP5zqH54OeMweyQmF+xn8UpRnMlEuQLT5cq
6wZpTAHv+dWViRlo0cauOdh+HB1W9wgLvz0A3W6uHtEKgfIvwrTRxfAQRf/AYtCODC2oSCmFTcrO
wUCpRWmC4Amv7FnuGehgNPHmrvNu9W8s8dBCdUR+13tkt6S9PpJXSA71u1VM1OmNVgVGw33e4GDw
oSMldWa5bs9m/KMhNd3vJ4S+nFZvLuoBv8Ejsfp63C74/5q43cppTMHU+tBdzTv+70loQ428SAcl
TUQBHuD2i8xpb9AOPURTy+xhqNygXtc1rLvzy5JoJyM0qIfzLHmEnKuvTLiSry67vWI88X0rXSzn
OO6G+AjCgsh0vtYuQUPUOQNzMAfRgtjMJn/B9ZWDV6jIGZ3octFcNRVQVLqU0hdbzdgzTbnP7RQF
SgJDykgiPUIBlamB3E11/0zFwosgw1w9KhKPGE2LZG9OYYZmMaRmqYzoVhdtdvOOkStvrC2gbHcg
BeCWNBFtXMUggomMRMKg4cEptweOSTpCz2MwCwjl4TEHyUaX5CTc9GYwRgplmXODsfBIg49g5dCb
eCRSGHM07Nd5I5IH75phH8p0uuya1MXH+yYy0qy08CQWqdM9DlFYs+ujgAAUEgOo9N3qqjrJASuJ
3QToeYtXX4rQ3d8nYpQ9MtyFu7fXceOPSdAYZL2Ci8w5efY3/asjXbVOU19ZtHSbZ8OfyaxL1kli
6Aq4dHmbtJev9HIx7hT4147dwXSR1LthZh0fgZvVsNSok9j022i5+Bh6JPxXpwdKkuIl3SwRfCBs
PJttVmI7x6AzXXZ9rX95KEXlDruZraM/vhefW0kzz+YhRDXNyFjjC/d0tNYfIJLQWqnlG5rRzky0
gddTd1vbhb9iO264GZ8zfU6E3BOiD2ZXIUsBKALNIPIGVhTdnDaUsJbF44HLnKPunbesvLFk4kgH
BisF1a501KTQQXVfKhbzrhv4BFq5Dk+IXp+i+xa9Rn/Yv//MWUIIfl9ERJXKGqJEt1szMTJu+4k1
Nxc7YcOjjLaDFKuPxYUDmNpSAg/z2Z683edb8cIXJRugHr28vhJZFkReE08t6jSwPMAJ/tXd2AXC
S4ET6OZ/Ew92VI/Zk8rmqpwbqgIm3IBUiSVufJZHXldvod5emhcg/MuFgGqt3yNOap68+awafdCN
FIu//g8ZzTJdOtpHxOTBz9pC+ijYgqcRZO7QcBFQNRaQMTdC/DEcSrZb9J6yog8zld4r1axB606m
dfZPsWsR3auXE2jK8BPZfHW8sTfnvURzRVTPd4sVffc94YwtN702e7e0GP3/vUCvolHx7rHe5IP8
hR5u/AWBiiEkhIhH6NXOqdi0f1dXm5N2T21t0lU96YpobEXdDqW374va/YXd4amvY7TuhMCoYo7l
CB+unj4RQzpqES/OdxSSU6da8Z+bmRhFjZruwVA+Awce8EDCGO5IlyBZu43/CH2rVLLSxKqRmrN6
lV9XBWtqm7ScUXqP17LoXi8krEAtU0X/qWry6Gf3VRGzrFAq05sPke9bdX+fvgG3TYoFGemA2MBh
k1ULe8rHaFY2RwHRsdSYzcYv+A/oFhuozTj4hEAtTxGp6RVc9opNFEoVQYwo7/po5VRNOrrWs91B
3iPxj3W/Fq/7Z+GYn+aSwGhgljsq/ghPZ1yCUPXJ+JuM8oXle6lkxGWhfh/Lhpxf8Vkyu5U9R1//
usrOuLFwGy1WDgWUSTCW0N7Zywo0SOPPG5kle8rJBehcK4kSp48lnLAKJxvRxzwDLJ1h4uLzlPSp
K4YEI3FrT/EOvsKw9dh1dofXDt767lwI/AUM7HI4LagejWiwbG5nYDPo4oUEeQBkskEVy16bPWrJ
2VXx9IzzXkfhbLYNLBt5yJ4nJKCxEJE5aR0o9w2r+cNFxmhHDtTMtBiou3MUM33PgTGLF71NlRoj
vv7MELAVr4rXICrF2dsAIxVaN1MmFYhitWFhxT3bUAvh1GWJUX+5S4kUq1PINlUCdbNl/b5ZmiRe
f5sH5jc74cTVV+8wJoC2y/vGmOwtPO/fh8n9PhR8Ke2fwShh9PGVc4s8uLGyTciagnKvs6gwtzAG
b6102egTpyMdz2pSnaKG9EtvFjPyMbtAallfknFzMUo3h8Dw/z32bQhr9rRhpeBOn8bJS+vFGFZX
He+AroWvA+WmckViBS3R87Dg7m5rKHPvq0yaqYoFRA6SxqCxx4ZZ6kNvDenm+YkxuzzbdlsDfWZD
mDFQF/Krqi4PDpfh8N1gWP1LLm5sZhIvRNIUGfdL/ICF+v2hbs2oGD1E8jU3KvlLjCioAMubKLiY
xHMG8RZAyKz7d7gTR4Eqp3vsMl67hDiNMiN6Kvwat56ewRty0EXGmMly3uI4/M+zJ9tbty6bwNfJ
CCMuoHP/YDmIHouDCWId2lua4gsq++LDqRRXYDCzpr2mqStGq9NueNT831HMDpkzyqrfuXGoM8E2
Mf39D4gcrwUIdxrZJzIkNm4gLIV8dXaztwX2RdVJ5hiJi7WxmoNtkH912xD+nyZjWJAJFIU/HSI8
TZtRR/+zhr4EfsdEUk7EFtFI9nI1ue3OchpN/Crn8xzZmifsYJuuaLouKZ/eaXcUkXQYlgi7KG9q
GWTxxzm0WIwNwXdnJqbaT04pFRvDUjy0o55VyUrc1T0UDn25hbJjViqVKhboZsvzWQd2Y9BKwUql
+Y4Qp4RsQiExsXRfn8G3W4fvEP/wr2hGCprRk64xudR4f7ohRV6zv+TxyLMyg0FtTj5hylhtHyi7
xXZWR3S00/bise3Lt2bnMPpHZ/fb8/C5USyOc+hSpPWOj6BwrASEtQbvft9uWNVdYmSphl6G3aqW
Cof+fpp9v+zC3YMh1E8pozh3dgWF42b/TWdDdWq0yw1Sta3J625Lrf1/QlG637VF2+TqI/LR8HbC
eazWrDC3nTIp50Iz0n6kgT02p0iv3uxlEK3D/kYQQv8vHqvVpAaze96wHA1ICNg3fJbWQCtZQkmh
zOjf6tqfBPdfvolGE7G6x8RIP/WIKlUy7Z6OOFqxha2J8VH7ZKkIEKazi36rhduvLMi6DOaWZDxv
4RbukveZxnLXeMzSn5jbs9DTZGZVhxNfjNUwVVFyKmJ4PDvXPn2EIkGsjIVlM1F8B8NrxTevn0wT
JFBz2gcHibgUGB99rnL/Tuzqzg01tYplp6OtXEq4pUiZzKOHmJk+jTj6XnE25sMbd+tAl4UaNJUD
4sQQaaR8L/uf3cILMu26JvCu0J1Pat1UVJsXHTQLhwNzgHqhoeS2viA9wcM0ykVCx3kQym8d1216
/xHx8/ZdicY/5bEXhyghAOBPAdlsgiEGKojZgCIK35v5XsWyVhOAAdje08gvGP+fpIGIF/4HaIqe
OmzI2i1bOmGkRj28+Wcj5sE0Xczjfs3fkTVydh6bYADhUjKmRoGzeFTsULjmoa1V3yV13xBUxnid
m7rmXd8qSZpPvwg4Ufuf7vl38GK5JlcwUZcADH6RDrGx2OyHS9GM5tUnZa7oZ99Qm0eqN8mAs17F
tYzFeUp9fhMA3owJEfeUp5qifg7D+fZY1JNn1GUCgUxItzT2p73f9T4+BuXBLgqIpo4AEXuT68YB
5ODxu5LrixUaIzwMMLKp7dHhPl4aiwZLDe/FXyiOii0QVUaeD99uDY/UWKFya+F4SaLsPABeLUnS
xZC7JbwWPCX0AXMFokzLvEFb5NObVGrQ6DU233HUFu2noqPUokpGPuMyFK53rQEzQ6i51UJ+CbnI
fxvYIvtoovfeqXzVrDak0VeFCfBIXP1p5GLoaNjrgsW5hF/48q5uNIXga9/gjPFyBbbkL57QWxPo
9xKtoz+xr9tW2kwGOOTKK5y4uJ2DUrPswQbHCb8H3n1X5VkSkBJ0WHy1VJRZE5pIjNeAMNH18C+7
UsqaeyzRLy81iRZ9zuFyz5zAv6pgYBmG9PYRl4xeHVZ4OxZDOvbUcYXE2dgo9fPqrgqYV2HWhkaN
KmXmvejehwPv6nbDX7rq6eYb1zY+AqpPHll/fn7h5q+n1SEP/8ya8MvhPsD/cmUnWDFxNluFvUZ4
Bvl+1dRl3HXPTD3zpxIL0dgRPnMawvaBYoMjBTnEzSUpSBw0tU9ZoErvYq8X/0lnu+Ptcv3KDKX1
OZMqo6BloYvUHeZdjqzjEHG+1oldOLdTEIDBkBvVQt/s4Z4TUb2DWOWxwUYKPmTRADKY2QyuP3v3
eVYpkXfivYX2GxOwQ+F3wSlhAQcEjKqCCFo3BIn7qXffkYR9X9KBE8sAmdc4sqAtH3bFRxCoUeTc
QA4lR0oeQcZBY3xRk0ew8AUv3c776sBaWL1aGFgblF+T4kdqWv2ITseDtO387mvA2YZVRu7QDgEU
iTPX2O4ZD1k+3BlvexyZTCK3QhcwbgFIg7v551s7kWN4dPl1MV0nR0q4/GkBtP+z0qbQzfHQqkzy
xilWt4gYnzLD+u5hDvXJDeO+zUcIn2XEtXxwYbE/YHI0Om4FkQRPmWhfg5wm+IGFhIeqs+TszuAI
znSlcr3XtfG9r/PcMu3/t80slqeMHpHsL8TuC1tHDXleZLF9hQqX3AK7CxpGKFzRLx3pLmbJPeSQ
xccR7VhjeVXr9Id5ItjFi5gOpfCyYd2WI/fFlLk/pFFmDPz69Ypdo878Q3GK9wc3PcQhpIw5U2ep
ujQqeAQ0aAott/ZMPFnHbTrCY7knfLz09ePMZN880bvIqoSbX8wNQmAk530FOZ+9m4aJFAtX2WZi
D+N2ssoegfUHsxysA3cc41sP2ziayDKoZyWtE2+VTesXZkVuwhW2HARGI7vbHs2L3UD+8EBR8DE+
Wl8r9H0Vp/gwhTGJkbgmR8IyrISAfxJ+kH23LoK1vVzP3RBG+kR6TUCvH8vq/oL833ESgQd0jltI
meojZ5AD5CL00WpHRARwVhC+/+vZ8scZwTQhjdFW3rtvPyeO9hV5JbEjCt6naKBaZnsYARuUtYWD
EsX94MPUK6yIQjIbjItpNvJfdhLL03VuRsj6thD81FmZ7qkSTZCWFMIpLUa1X9iIsdjpEVSNErBS
tAgocq/ulmCVhWIXZ09uadBOsjZiDf//tDLpRLvuHwmo/g/+b5tXtELaXOF6IQxyaW1m/jci+gSp
iXVbMXbHhW3ZBduonpBo0uvBS3XwQXHGgj5q7NaLrrWJdUPPm/ijsi9q+snlxw4jDj1r0XkK+cIm
WDKZvEPZ6LiiLCv/Q1iuBmW7JaMGqwrt2sDA2qMlYZkB8UJIhFKxraP3+FWy2PWsanhYSW7rcOtv
8/2u+SArdwKPGxJu5zJl0Hl45fawC3PILwgZdR/biSlykfYoRuEaVov/o3CdUzA6OGc+AQhPasQz
Y/iQoQg2TTWIWxTcWVnenjBeSlWolJj8v7uh7V6omJfsFxooXBdOb1zK4jtb0mTCWVbpGW9QYmuT
avUCc2ug5c1SVU3iBBN0zufl+ZB851OhcLJZQvoEdBcSfGyNYhP0CpGXOSvinL/69O0i1IeSTDnx
ZpOQgFPDNVdu1Rb7jRZR3Kl36PjHA2+0JYBJEz/vsYE5QcRVwz4cCOYHrDrdFCgsp1DA3aldFSYj
5XfW/9eDIHilxg02MlAryXcl5YYknTwii772GmwJboDSKVq3iuSuWusRieAyUZS63VBAJXB1QeDx
3InJM8m3pmStbqvBlb9Puw4ISR6iUhsjfCF9RHuA4WsqJemCkj0MGwi2BYMG8PsfNsRCFhrQIlif
3sOcK/3YxS8KQUw80N90SVFCcf+sSKytkr24vD7Lbk+whkKymRO1/qgJMud+rmALmVoiz5iINoXm
MtT9lRGg5PEcW/hQ3YMXyGzpC+NW+qwcmadpMWhkpkd8eurzONYqzfgr0OYmC48vOWeFHrIJ2qfm
6bmWfkzNGOe67+R4Mo4PbSCEXST++D+KTZPKc4DT9nG8kZtP2NL8iU7dyoh2eR5xNxKBLR7veW6n
HvJrY+RPaZkquJwHd01qFIc4Oic3ehKVOAzEtRRYIXadIKe1t38xhaKkZIcScHjrc5jHeP62CJvf
UWVcmKIhc6cyn05r2hqbv7li6esR27rHED6hTuiE+S2fSewnhCWPgef4ezBz81hM2iDVd4ZMGhc3
AxuFnX/ZtAwj0nn4qg53Bvo8KwscK0kxqJWpDcQMnoE50krdTjnIgmEsqoHTixaZlK97Re4/0Fbx
DtHyavN0o64yhQLN2CGhocj8UGkmyXbUqh2alWsbxpXrvZvWgjYhc7071QxpK589Blo90/9JKKka
L9KcOjNbfiRlwnYDSI4CFUO/teG3XR45EUuyIZZv/l/MZXV06Md2GYH+X96kQTTOHEbIvSCowwRb
VgORUNNnjevFYo70fgr9xSAtYYbVl5UNX/oNyJ6s7da4A93j/CunXkIex9QEM6l5g4Z3QTWRAops
kqA2+wrzfXhmGc8EgkIaf/5ox4ajr4hQkUSu26QMMQWlbm9wVjOI4JcYgniP6kM9PUORD2tgaYw9
pu62uet+a1aR1BiMnhYQXy1EOREvtg2AHKvqKD2+dAuhdQ5qQbjdxA5J6O7HKsPn8rg7rK3CKbY1
6mRxqgSqLbd3z1e3t6xNhMS/gQ5BeUAs1UiG0vvRBNCbObZv2LI4vaMh3mxXDKiWcdmeZD4a2Hfy
KaRy0oruH+HN8TZdcR9emK9om7dJUmeqo+ctsgnA6vK2DSEGBmci/M7lhbY+Up56rNYCvvL/+lZs
wnBu76bDEAEL/rwZfgcvuRkWVOX+v44oiv8s2r2B5lQaALvr2iLSU/2/MdbzGL9pTbc0wDR9GQUX
moNPRrxMl9tDS9k0kDBbyFcLPAZF51U783CRsvazdRXSI1dFhaJDaT/d0bYzkrk50tphfiFctooA
/5Ha27/RfV9r10jR0MVz6Nm5MLQYSBx0f2rOh460R04CKEq6MvMj4o0cC0zQdlPD8EnUpW0J42Nb
Fg5i5q0IOOYefbtOKHuO+g6hYauCUQPQGSAfeEl5XxVyz1RVO0efrtoXYyfQUZrGK6cVWxepd6EO
CnHLyw4eyb+O3faUCWI2SnkeI3VB0ziLBi2LmZ9rM2uyjX8aFx6U9TmtKulVPx75CnfNxlox9/3+
OSnLtj1O219LN5/Iq9umLY25PEP3CmBrUV0yIlz9nrun+tlDJ6014HiRbHJS1hGB3N2m5i5PnZVr
alCNHw3kgKhWjcNTZdbxE0sAmsOCbJGRYPhktBCr9wMaACHRU4AukAIBBddWPYssIU2YTYUaCce9
YeMKf11tDPXYWHVBHm6ZaDSJMC7GfVAFsNBFzHWd0M/hzqvipBo4+hLw4p+v2uFj/Su/oHktHGhI
fcfgWIj1EC3UFI4+BsCf4hvbogiocioMtpss3O7yYPdhriWvBuTaVtqr4Md3SQqIannRrN6fvZei
WFNA2i4I/VzCrYvRUS7lUO2u7LP1ArBpiWtpW3nU352TMjABH5SWuO6VQGeW/LIaiLFybuFeuPde
Em7qiTuzjX3wLXj8fBwDBEZQ6jG5S+bOaVNDKNIFCnPVonyHbyacroYj0veJBayfalhPpDfvejHR
w0vCx1LYeYHz5JMCTeMOQHM7trrE9KGVvpTiNDUpHeKBoR23T4rSDq8nl1tyTLVakBWU4gYmdHo1
8kuVK00mLYjO+LTfxJugubm0VRfgCQOgmx5Ol929jG9NhwZWyDuY8bF9PXsPIdgx7HyS9xPs2qql
pdWOInFd67Rnnge9gEoCWungrqmWjlN6TazJjdm3jlZlVXmZm0vke4FJ/RfElMjZ3igVbsVU5mI8
sydZVTdfIu54XZeqmW4AggTGXRU23a6Vi+pzLBAlQTaauOkVCzETzOyKAE+idwErVYgLF2ZKphE3
8i9TxOBhfGveKFnCxW6i9ZuzrtOZ6EUSLgBi1UjboNBjI0dHzgbfiNw3ygatWxXkVAyLa8FwhC1z
9Qv/i0FNBB9MSOR3d9iOAzRoqj3YxDTDYax8klcg6AFOEcdvRdxbEdDBl8HvpJLkRqyM/jYWhDDe
4zqsuSft4Oeoeqb9G9N562Cs1Rt5oL2TDucswMwkicilnC/MW+UevM+wgB4AM0pkhPunzDwBDzFw
h9JfbRSAWR+lImjKzsuWU0uhWh/jxLysrx3C+jIOa4iVQ8sjAO2kL83EBZvu3n6YDJhuQgp0X8qw
2rfE4Z5GnPXiuxXb/P9PVtfa0nKY4C3+POSOy1oRtxvKTl4H/wDEAkA6Bs48GHsJE1BKx7ju9QHD
/HwClSB/hvzIeJbwYthE/YOk8nn2aN+z4ZcV019ogV4DabbxPFo9DNVMfieOqJB029NWrN3fRUFN
B4x1ntltcp49lRjM8pZq8j4FXl39BxhX6B/711/AoTE2lMBrhJTCdRH8XOlVIFGJ8EdA9ZX+25ye
zu5xjz80SDgNNrj5irFyySwucNcmL35K4UFr0rzAebGjbdzbBYTAbX3cm2a1ylSoWB+Uo4KOB288
BSdc0UZawrAOct7LgmAyJg5BvkaCP+sxgb7rP13lsAut9/PvGqr5y3mPAQf2NHKTR1sMwithrsA1
RtHyIrf4bUcZ6j7eJZcQK+GiQJF8y/JwqilOB2UlMl7QKZ0drU1H/QJ8rrpYjaxHFm5NboPEZSzH
/+kDgME4tF0p3IUHx+e9Vs8+CRFzy1orm6eI1Cr6YHnRJS0GQwH3DdH8nMkNHErtmvUJMip6fXyS
fY8pymle6e62NsZzFnD/ettE7rNt2nK0HB0LOe5fMv7M1vNMG4e4RdLgnL4IeZKZOIgr0pR310g3
Shq+0ZT0FcZ1FqT3Pby7qLdBp36fd7+mxiwPgqURu33/crHIh7JnAZuIh8A7TvPaSErRhqONlQWn
HJnmK4W4I/ycPqOyTOhdtxmm0LPW4mkU99Y63a2SfluNpDsf5TQYhVw+wcmIz4JYHADbbX3zxnO9
mV/IJLiBVFL16e24z1O1JIq3gv1F7RDjdrbKNL4jzt5pwZofx6JXD+iHW3m8J9TeHARnae5Vu0az
yc/rfhNAPIjEkOCKwbF1NJRoIwIdaky5fWCWNye8sozltCV7nmK18aSB2qcYJo4qjQnBfpf+NFJx
JxZ6Xe58PZv3KR9ZT4ptsXaeCAA29MDu/nT5e7DbNLd/Yuv2gHiM5TcW7qHNjpaML/b3bEJmY9KN
JveyhI1MtvJIKyJCJrYTsJvW2HB7RFqC0NMgz3l4vkG2HD1LZoVRGw71v96WjKL+99QoHOCKZ3G8
3nJz/BvAb6w1tmXpV5OptioMk79xohNkgFzg2Gus1P15ly7dBmGkPXvXKdgaeR53VXyflDA/qiYs
1/QfE95ryj43yq4/imSFYliYti/FkcfcIkn9JR/D5bfigg7a2trV7oO5NofGg9f2BVJKp+0TD6Vh
JotjATLtP+MdpjoGzkmqMyXaCa5vvTI/7Vncx7H3bRrfSF9vYkaji87Dh6qdKGt3MmJb8mn4R5+X
ARO8I9b5I4m5zDfDox9i2Idc3bxWthkmRkl/uqPUdr7K7P1VhpiX86WP0FmW73asJQKwauJKD3AL
sk9B7H7uWpX8bt1msddC+OVKUd+rh1ghugbBRipaKDiv424KvgW/XSOfsJ/QWYox5m8T46v4nvfn
jdamTfKv2MWCXOCwloGCe8EGqtdh1yVJcqMbw81u65+PVs1bHagIYA7MrltphwO0bKSIIg1drJrt
YzFe/fhsMuV798qNLesRWnOdbavsP2NGxtfb7t33+swcIihRmxuOMZtv31lFBsjlzt9eXVwes4Q3
7YVLx0au1kSO5OKhOAuoxPooRfR+fJNALJWJ+M3bQK1RuI48gX2mKjUEhsFp9F2wzH5LXTae7qQK
/3EQSG5HidocsPZHCymvUYHPK0asc4TxC5FeXnFNJeZgrAQTlJPOcwM433oeNGbi39aS4g4vPlqd
jfIS8O5frA8V4SlVFfTcu3GtgE2z04Nkh5nX7k2Mh/+axFqhVXrZTrJLcZhITMoivBpUI9cXCgt0
zvKf0yJ3dU19L+rvz5vTJxWvVqCND3J75nZG08UVcVA/FAuxMmhR9f2qYUvTynEwja0kF/NmYKtJ
mB0JQ8sRyhIefMiEdHP0c+xcWtnz3e+KgJeYvHeu4EUcQPkxZ65vHXY/YOmr42dj+oxAOtp4CQaU
ruR4J+Kdg7G9psjyMrio6OYquZrgWhzlmiGE7kUYdyUuzMZPHd4W4Oyk54lIUkzLIrPXSk5/3EFe
ivbUcaBKdGphtEt2EfB3hGAvzOYUUXkxFIqJ3ziJkqXRD05C0cfCeu7RkpbmA0vkEUqhlkyXWjR4
6+H/vAZh2mXtr53ljva3/9vsnuDZgPHVt8ZfpBDo8QnW41w6BF55F2PlnbmgNOIGSeGqXJu94xi8
FkVtMLQLE51DcBd0hQjI2NdEldBEq+BdQUoGMMyFlIQu0z7d7hbPOgxGGTG8uwFmvxMljfu5K4du
xAVeigluqydIXVP64z/O/vg/C9cKjnEsR6x7kNoI3KYab9mi5rHw+HjnzCBY0Vdd969TtnLVo+Nx
DmA1qI6D+eSc7eZ08cjHwoCUhmtgSL5mSxuIVIyeSMULPjJoMQ335yyhf2HFbLOuiZ3ublaHduQg
4Xkk+f29zSKfqQbykKSrdw1tUORXvAggYjY55RBc9kJE1mH51m99DzZkhc0EeAzONfbaPi04yzVf
byfft8JVpwTYwOXXmoFrKxXzsO1KTPa1+fhVSAu7vsFfx6ISufaig6zNDczIi6lP6F8KXjwmGyEx
uPP2u6ylJx6Ru3IoIJDlGC6XEDq3gCpAZ8Qo4DpR+qtPQs3fReNcJMcMtW8g35THILjn4KnI+fKt
7DALMZDl9/QyB6JXc/zEIZkfFZhkVRM1h6yMAdntxKlFymYrSvZ2ptN1GCptR3IiGeV3bO215yWV
7Ik4S07OAKN3SMO/c9uxu+Xd1KaVqUPuqqjTz/nt/GDcrcbthfn3r0KAuGPsnIUp4yeQxL8oQQgu
ezOTtDjuGmfVW6HrfKNpW18AU8+3BQR0/c00w72ok9RRm4zhad54yGkI59cRBpe2Qeaz4yAAhZNw
XcBWf831mqQHFw/CxPv8Jy/6kxgHElLO+sgA1hCXEp3r6vMrePmhhVawXL8xSYqDBPl4qveqvEps
x1jxC/j1swASJDmLg4SGYX52mJoEweyPqKxGMy2/v0I2HLBN3NYWo0sQYwMEDPw851jgI3Y1cxb/
bHTguFEWdu4tOYozjCyNBJ5l5HXqw4/0BEq4WFcKnHjP3I3dvnmFAA87mbyn28FDfe7PTksRTm0k
RcOBRpIniHoeDIALosewXqE/BqtDCJHVLasj6Z5r6CWak0hBH0oVOu/3/k121dcCO8L86Xvbcb9y
UIXPzAtfmcEbPLOyCoJCl4QJ5vQ1WAzeAxreSSeMVqksB3TCoTwZTo625md5tIAodiD+y0YEXL2d
eJQCTFa8dmuFKGfLpbLzjB4isC/unCc92+gEZwoFTUrAJeTsXz/5Q4smxzZYccYml2/pQPsuW0/B
et2PiRNqbPZ+vcySiFB267ZCPEHf3+OM5yAtaHAcW1b5Ktr6TqP65I21penAixcVVgoQ9R22zO5G
SI8CutahRd9hbQOyiVR63q9N/jmC7chZiyre/6tgXRClfRboQx149iBZgUDot5gDlhTTwDlnkjTP
UzBkJ139uN6LRyRwsY/7Ce+tROx3adjweLVbi/7auWtsIOvPyWD7KEmPs1uBOo4270WuZKMg0yhZ
8s/oott38gPtqhVk7JdPVxaHkiJIXw9wKeW4lo1JbfkTc82/QqteHt/ODj+np0DardmxJEkL07fY
z8w7dVVCwSuBvmNL9c6dhBd/FxK9PqVXso6R6NXKkSKTZQVETOJeY0P8WBLI5kc3/UvjQwFGM/u2
uW8Y3ppk2KskXcryYAiiJ8XqzmzbirNco6T7F5OcLNmyBq4M8zJ4lyum9wu/Mh/93SnPItWilL64
5wz3psZFRhNT0aw3KJJpuKD0gufYY8gY9p0jM6hIX7p274ge6h8R5ZPfjRytG5UbTKv6Isrotn2r
HvmNaUanvL+DedpEh5OYYq6CyUcCsY2NyKAlAnQWBswD2KgoXSEmDtL7Zhd/rIQgx2XehrgPNszl
ZVNW+t4UoVlLx9xkxcdb8BEAOv5ndf51vBbu67rbxY0w81LaUHdHlCGsHTCo2AotDXIWrB24tcVE
PwliLeMFWD99a7nArB9s+5JlV/2jXWZSC/yt+0grRqTGkDFoVYw7c+woSYexm65+xAJscnp7dSIM
DLs2X9jekaeDYWh8MjWJybXqRpJKOdH6IN4Ytv952tlXB9wyi9GKqLxR6z7stBavSXmzTErNecTK
MvlOasE8rs18qfhH0JPgKmhUu5yyiselu3EhxtvRRirBdIrhcoqPQjdJMt2MSXi0r+ytNrnVDx7R
F+topUgLagg0Qs7n10RmGIVFLJCQ5r6J2gy5lckp5q6mL0wJsYStTpefdQsEDW7CqUCzTJU2Lw7h
TbDoZCLhTXgErOagYVD9l6vC9jzfZ4TT7Hk6HE3PCvdQ1YHvIhU9f/8Je2l5848YLwf1kwaw7Fhq
gRbBrUDD5qY7GpQSvd02RgZ1ae8o6KEdvpzzDx2h0COrWT2VKgNxhnmJkkH6qjzz7yclIIW7AsPz
5B5KXO4dMicS7Iqxy+2q5iTb95WXEPQ0evmU2v4NxvZ1eFNU1Qebor1JV1kqZ5wts+Vtaf+MvPmO
gTUskfT7I6uEe4yJuIjgWzammKV4lY/3oJU33K2W3SdINVJbN2aW7ErUnOmfZPENVk1odULdM+Mw
WBUhG0PmI58b+JuuffEVMeHZqESel6NSw7kgWjLws5a1fzuOVlExykgiBdZdizsfj+/x7g6n7F6y
MQY3LYEYcO4EDlVFwUOD5lcqt72EiKTLtIDUNh+FjyrLybzdNYuV1dwVal5rnzlDMmcqitQA4u5G
aGgCm4dHLHe/mEdXXkmhfKc1MQr1EBAxU+caB3NRxcHPtMveFcOXGsvvQMXMeIA4n8xnsWAH0A8U
VqgwnK1GMYGh0rUdYC9brs1pFzYXjs4RuHy6qt01YUEOvSg1zD7ozdD6KFHTzHsbI8v6FypnYOIA
RNm/DFuIZ28aRRBVU0Ocxz2wavdrr7MEKUnTmeUUgupT5tt6VtW81QBB45pbXaL+RDDSnq18u7lj
LdahunF40ns3t26z/uZ3+Wlf0W2tAXfhPJhX6SC4pjVwZd0pKnvGLvTQxdNom0ESeEbS91lCKaMU
kFrtkUGItmjLZZ0LzhnLR2cRKIV0T+/I2tN24donbxyotH40yxB+y3iuUu4PV7qFtDKx6fTnmJ4Q
5OHNoALoc/3uQ0/CWfs63CaHGmG5OMLL5ZajRLP2Ve4ttYKDSy6ZUpJQdwYnZnYFTtLWv90mIDW0
BKCvQ+/ZS+BerNp6vbZxJ0pI8h+120ejqjp8lVbaMh910Jzhwi+f5y0Mh8WPsiv/oj9T+YQy62O3
aJCaxwz3JnJSBA42GvK7bjJ2dEBeWuAJYDblUhOrPFIXX3ANGoKJBT5siEcvYu7cauhS+X8N5g7d
YrL2y7pmtzOtJvbQLQmM+sMxxY6yIicAPI3gNetFnxpJeXi31gwHj1ImuuEvDhc19/HpOv37dQ42
hUAkkncb7MFtSbXFCEcqyxOjSMqdW2SutayeBqhOi3fh2rmwNZnuu3h3Qya60swmzo47PkM7rWm0
V9j3Md4jChzIgpsjmrUy/3bvUU4HVx7klYmv+xQHD07vdBD3PhUTuLo8EmwJnMM3dWoNT3Y+jgVW
uEeFhandJ0IscwHQlL8tFL5QeFM8Bux8Azfqksp33nbAGtM4sQGcOiQrJ+ClUaJAr7R63130kQ7/
eqzimAlJlrJ+wShwXSbYpTpus0QTzHw+zU+fToYMLCHdfGbwzBVFofOggUiRTnxyvaIrWaO5oBoa
k2UDAFlXU+IfLckrhjMWe8hB51JVo8qQZdf1vZsB68PyMgmXo2TQgIQdQSLLuncPXOvPz57Amyax
tvf0X423ifdnDo8rTxGnYXdNraULa7PCTyiBSbU31re8iAtPSUcZzjfsa5jB6z1Lc8Pb1c2ENUe6
YfMhOTz/8rNH+DzTeg2la5QxBZKPbpC8CSX/fsuaEM8EaI081Rbb29mDHgaJZMFHiov7c+TigO7M
GGJCBDghiHJl0jl4+lJXma/wt49uO85D1Frt5NYneRvIXnNF+t9ACPNMVMVVp1Cj08IpySrRfYn8
AzEvdmZKeVoBi4C/Dw0LaTMHDyw0mXIadBIEUobpb658JKjxlb/QWEkZGaSSJrE2uZAsLo+srdCL
XovxbzULzciHnmyLb5nFMlO6DgvAxc5c++D2qogxQ/zJ9SOYUkG/6afaR774Oty6VU6MGWmmJU1C
utamvHfhPvVzGiyd+LyRxhLZNiO/r3g12BVZfEHblZzL+fZaPQIsQiFZpy18xJy9oBWRkS/fFVBP
cxhKxfmeTRrSmv8pLEoNU63ZikBC7AmFo8sg7zl61vPNqpM8n4RGxp1pEjm7Rzqprl7OH2ohrvvS
zDj/bOvRp/Rb37yYztlavpTWdD8MnJnQP31A2PVDQfmFwdXPzcewoYbw35MCF8ThK/j1e+4YpffS
CAGsz0PL3l6fm0ZaJltdsNql3jjMJEgz2yD4L3+9EkclYjbQuWSPl4iKzZjsW2FijTWlXdC0jxIy
UoK9GbVxm0oWnwIxE9RbxDkdg3hJBiplALowsr4zH5278BLQCVWa55W0BWdTi/tR5p8DUeMlVLCA
sewiZt4rGSo+NdL/ujMj8JEGKzskv2GuXZ890OnbAEEzZ4enksm3wCLPXDc+OLYMKyVTRvmqoZ9b
119nxkox/JQ/rhhtmdkzxHb3u9pyeysgK9No9cGek3xWeywV6PSKajxbtDyquT+EFBE+N+qf2ny/
1FIRT9vmDThMLllPDoCumwXGNGhVV2BiTG4NjLl/1YPkosGFkKn/EazMoL1DiG1AUlHj5AuL6Qc7
cDuJM1YRYL9ZLdwJmx2L2JywiejnRVveaCoPh0ltDXcPcnJzNeUI0HRxsSF+Wb9oAlsmlWBM/wvA
/r75lcwTiAqrqb0Fesh2yLSzvKCFO/N4Uft+ZtfKmvbX2cQBTI6S1ruM5RFZJOWR6EaGqT35czmv
b/xCQF0UxXY6tAOVRlix9I6u+hSXtoaQrM+qfh5M7wtJ34Bsxjy7l1acD9nngFiNMIHl7ZQTTSfR
RQpFBqXmwFSn9I2knG4ee96wrdKhH6a+TdGcei/qWJKdJW+c2PuC9jX0vaDjc08m4u3AnNqLqSaX
CA3P9tI6pItIQsWdvi6uijfRYO1TsmLvAbgfHy1uE4eeVBqKqIBOG7VRIpiz4hmO4J/ZI5wsmRYM
kiEjN/tEgZAJNKityB9imWmVDB+KJMo3NHWgOb8joFgcJ0/V2HDxg9uEZXmD8z3PONe4xl29tG8+
w0c+FMhBmUbCzmv5cKUcfHNTuN2J8n0ciNW/JFDuReogSvr36IrFSzG3Al8jm3uSA3wo3AD3nfDl
PrI9fMKh3L1sMOFefjrf5S8JKWDI6mTdzna9aQa3+nNVCjE85tcEWrCv/08JpvlezyrGAeQxzt+p
314YTsepXU27jPbj7u8LHuZdMpXz3KM/I4iiUJllWsKtaluUtoeqAxrvquGxF2wSsezG+cBvBIeR
hSh74BU3lzhS4mtMptd0w/j+UEZ7jytxYz+sqjsHoTUka5g6e/h+M2C0utyiko9mzxE4vFT6EeKo
fLDLYds3TJm0cye4X+O11YtYjwCsL1q8y0AKZ31q6ytprM92t2IJ79PFqG0EvoZuWKlE00dKB5vL
xvboT11x6ofofFOmH3VXhYBhYxw+aLzNwqlAMUzTNbzMgrxUMGjQmW85yV/9qC0RTIHcUo98eGK+
U56gIRec0uGu+grtzTPm0n7lT/xchVjsNnHk+fk95Sr/BwQEv2BdqN9E8VDcKYvI0CahD4da1PMz
oMUxcKwedEQuDLSaqze3PPg4rqN0NYGiDF+vQ9IBOvO5BX550US4h4/GDkruRMXmNzAaO5RhJcyj
rMHkL4KitI42fjum4lT4wm37W2yHOzmjlHWENhABTdibptbA12k9AEcN1NSoTyso/YxcnGJFhvdP
QwHCC9Xl1+Ywmyu3ccPZlZ7BAQl72PwQVsK8FMCQQubIh35/2Y8JowE0GN6W4sIH9NyqFiDzXSj+
00qGKqwnq7m8r43D8G5BMxDyP0eBAYhhvPWR0LF/BA7dZnIky2qNFyBbOT/W3t19lV0RSwyzriRy
1WZN+ZYhFcxhan7RYoxYamZSBjlvMUJ/CWEFIY1GHUFvHkvwR8rQOXF8SW+XQ1GNPvlfNejVzUAS
9+0eaSFWACQfzQ8hROym9z2gTbnbpUq4KjGwqMb/ULYfDuGZOlf5/WbC54LaXSJJfBBxj0aGNKXI
tE2bCD1kPIUEYS8ooEqQJe+Wzelb/EHXHXhgq8iOx9eiZxh2dwJxiZOuEKL5rvvOAmAojUG2ZxtV
gOOvpILOY/8F6UzYtqrU10/+aWHnvPcwPZeLVa7lteoEXGtFdCR0QeHI7t8kbW56iRtUHgY+eW+n
TsZCJ9pDvWyoxdDBQAT/ktf/S7WrqLD9F64HFyCZPTGEvjeME2QEJ1Lt7UnBCilM3dXEB/Mk9itV
tnu4ubZog1kdRn6RHwyTbf+7f1AD/xZwuGr+RMIo5yJK/sJtkMwrsIPssFohfG+FXG/NE1IBuJdB
9hZWhhc/W48+5X8v0tQOP5SZCZKur8jI4sIxoj7F1acOwpGAy+wNNeoBs2bXwVSzngLvlDYPF1O6
kApJqciPkzIJdsZi2LShA4KXgeRQmjqPly+DBDdubuLMVkq1kUvcrwvzOpzdpePz5Va0bUq6N2hy
X7i1jlsbOzRCw3OhRT74ZKdPkG4yu0N2InybI2W1wkNPYPt37C1JeP6fzWvQuIH2IugA6DsyBMRe
ZRqNUeawXP42g0wUYiBcvL66gWl9n/OVvvvGJLbmneMor7M+m03oJQVtHlhoTzidc/QdEJ0JD4td
miNnFl/s9kU4jCDZBNTavOCasv5Y408DaPKiHJfKHcunwr95qong6t4PSJ2igBL+Y3I5xwK09xuM
B82MChLRLrSb8tZWu8fZXo3m8Vyj8QETcaPbW3JkFRhd7/6zIf+lbTah6jmdgBBUcJDDHjKOLqm5
h4oEsA3mow8WHXxEH5akSwu4M2Bd7SPU8tThOz4WfTrLqT6EoYbW2nAKXzVGypQUAE7i905dtckQ
gvT8r2eUv4T43s3iYkL228/R4W6vQcKzkYF5u6fqIk+5OlsP2tEjcQMfK+P8qyDrMrXawClFiMB5
QZdd7GolKEXVWwARsqCG4uIJIKgBg931rcZfCCMpUgeElSB5kUkjQe3JR36k58JUX3xfYZH8unXe
d13cV/bFCtpiOZ0XYkyHgBHSfCP+l0seylJthbZ9U3JE/qqrVq/7x86lxHS19VGmBcWoEKROu0ri
ArMMYRoWiQyqu+OznvCbS3e5ypEOX5LxNTpVCl1i+wKKyhRVJ4Hri9ortqqZLleZ5mNiGyfP+xg0
NssD9eWVCcZHC0VyFJR+b5iszgn+LyEcV5tNrlIb/cvbQIGnNgrJPa45xB30zHgZ+qder1HYeCXf
1dzJmWMaFBaJhTjWaVM1znpiaCoREg6DCKb1QLY7hrGhz1Q5e4Toe0TElVLIncTw6KTBbLnwkn9o
pJfU6KMiT6w/X6SECwo8mQng80YX8UXGZQfRXcu/uRlDzZ+tMjuBDiBFJJ+qraTkMTNBeN1ohWpZ
ek6W1sRmCWIt+OD/O4tJtvjDMpzaMZ1aJA8/Y9OxV6nZ7jrBdSQEDm9vLhq7iZGwK4Q5cArxT82o
7lg4XciJJNzHmivJqNbxrP/C7O65CPD6HxJOJiJ04aLeS+sArihXHx0LvdscfJoQFndhFFp3Pd/C
fXsxQJXLTSMRPdsUiuA3wGOl7j5pN66vR6aawEuF9R2c9ysXkUHOsdH7Hz6d2x2sOPJHaqcFbeK+
8rp4yPPxN1n7fTZww+If93ukj5QMrlbG02eQlejxs42FmNKoz1Hxa916mKQ/xJl7xi8llmATNHlP
dHyt1eMRXFq8Z89jFbr1yY5zHKqJA5YXhGxmqfXmAcn32W11WI4Ttxd+BjClz+CFI7FzLK+Ug5a9
HkdFIeBlCRss6rVyNzc9L9CisjSHzNNvA/lYH8BflpDtI16I9Rf5I/kZRsK4gXh4R0tmvfaQExCD
Arzv1WWLRwlAWWD3bD84TF8UXi/jOyno8DDHnbj8Fckqx5m8oQsR1uFQiwBpqkbyi3m5TEYD5Gne
8J6+eq6L/ZUKSPcH4f42gdKDGdNEdPTHtd0joB5MzHnuZdnsW1iS4nxGq+cdlLvrZ1X6z0JTBUwr
MMDRnLVyLogLdwq0OIHd+WmPVg5rtuTy6BNYf/c843rFRkleXLW3ky9a1nNBGowMOXRlzF4TkYvu
6cPhPVtZ3shnxQk0cvhWkHR3omw/T6BuL8/fRLsN4p6Ae5T+80vRP8gE2Q1Ke28bEgZa7mAmiLcd
w5InwNh1gq5qoTcVohXGN/tTlh4ARyVZLZ/aS2Zwsc80JgVgxhbTo5VKv4OHzg15B7jbXwX+ajqK
eBdaG2X10E9gKoIRRvV3kIYdlSa1moMkWZ4+pghk/ZhyFKyQdm4XRZQUNJ+osrB38RkV8HkYvVbO
n6Wtw8b8S7PY73Tz0r/4q7g2bX0sm6dC9zrl2Z4Zx+B+lDxucrsvqgjhkN5xTQjr9PTytGW3tBL+
/bJnvtaFjSPvhseQxnaCkWHVqCSfrAcXK8R64Yoc9GKrR6Ap5mwrrMZh4vaUPfo3pc0CRhjQE9Xo
Nm+AB8A9xiLvxo75Ot6ZlFd/VOjH5ThWXeJ+woMD+IZFYaRgoIVX3QgPD9LH8CqlmaIeN1MbXUee
GZlhA/XcZ9841XXJcV3P6AVj3EQ+dGcdxgI2P+RBQtnYGIr2UZWB94af0ymvtg+t+14OBfd8vOzV
nidAmv1vo5zBM8NiKCZ8012xryzRhgIxMkxXGbROduvdL2Qcov5eR9xZl/SU/tmHSy6cnuwJhnYS
LycrRpdJuOKR9NjnttC96/uquMbuq1aAPI0eXqoeqovOKVK8unPmFFUOHirPwaE8H5898aOW8xMS
nVXnINpeF8kZyXCGWMo3s1F/+rs1O87ujVIqgIrxryWNSm/NcFRMaS2asZJdR9UpsAFfRyiih3Hu
t/o80UZXdI22KxQmBvZkz1yd4f3xcaDBqpZbkqQ4boXJdX61kyrZ/pGa+N9fJfPbcLS/1Kw+e/Jt
Dcgj4gtc6OsLgPnBT6XvJOn7wC+cHDTdT1XPuStUzadvkGjalACJ//thbvgIcR6Y470DglwWRQ7S
h8WmBW/2f2h+oDyFSjEN3jEr5BVFJ7iGL8Xk+6YLFDplogkUodxCJi0ZmHnkPy7SC+YZ1GPAHCK3
6htgBT5xW+rjLyWuJkIVmM0Be8NonaKSK+jJNQrvgGL8a0j7vBFi0sUkYSc9Fo9aMvqTErtVU8/6
6W7NEI+k1oNDmZAG0lIxyC7og4ZYMhpbhNqFQY3lW+mmal9noDClSST+TUXJsumXugnDUzV7oJLf
zOwiwJuOUItV8OfYys+0yZdJtDdRuo5zbnf7VdYZi5UW/obfPUrBP2uS/mWhaHN06RSUBC0iAMca
ACosje8iRwy6sGgpka1rQEbZTkGoGnOhp3G1u3WXszIw3zZhuCD2zOKZ25w8yNzYlCiH2/P1VoU+
e2tcOZcj/ArjzElqxGKJPc473i+J64M3Kd9kD0Mji3yEpCtKP68RlT3yhB5X68lb3iRMy5Pokeo8
vfS3sU2ZaCCQawCY2ugUDMUQWqCqcKLTccMZRqhYUGfYyswsN6aO6IhSf5kOfSwo+N7hJxdeueiK
REPkmwK41skXF4FYQ3lAT6zzI5yv/b7D/CbpezXytQ/Y8A2o5pd5/Hg4cO0Ue72X+sQ+Bdca+3KI
cFcsHqoZwC8Pt2tBCEqYeCSy0x519BzvULRaQGH3BcKNd/5jc5Kg4WbMs2DDK+hBGqMy4HjQhV+L
bAVKDRuTnnuw4s3rY7KfC5DfGbNklIcMxZgsQh6nUL//wnvfix3ORZy0Hv1yzNBM6S5NGi8rfLt1
T37KaqsCEN0RAtMzSn/F7Bn921BuD/8Vh26/ZwcVi0+7trAQNoAWEtCKU/RszZcGx9UnrOuoCooh
PC2VjdH+LhPaZzg/CODJDtEXEaJY/ffLBpoTQNsoky0loW++QTmvjY30CbE0be/qF0BEpoCIu6i/
HEP+ZjZ2IffaWGSVpL2NuQ9XGQfowncPG17VmfF0btY+GRNlG2RdFA5PRpgt2gumcjN5HP4cD8+Z
oAl7H1FZ4Dc6xFEAhWw6HQAaF9N/0NPafNddp5OAgOhUO7zVxamySpquYS8QxrNa6ZD/9U5PnBe8
pPaWgqoTtU0Bimn+YHYJDl8qzJLv6/zzVpgDRlD6RP03yUElT2qkeD9PEXwq5XUjkh+HXSsCnY3j
YhGIqPFBJTulMAPS2eiVoXFHcjWpabbwsxumcmxkBTssvL8R+rrRWnMdrQ0yNLhkhNaObPQ97GwT
b/L861d3IN+SBNZ817Pkn4mtQLs/6/hpWm1lHo8Xp9igREJS30/c2rvA5Psw91GGcNuBT/3x2Trv
CXI5TPzI6czWa9wspuaaP30KLWv0OmRAgRNEC33n2F9Xz7O7h3tyMRJiEjP0oIMy1zGubv/v7EQr
hWkb9NUEyfleuJc3OyQe/hkyfNVURQ1pd9MVY9SKGspaf6djb6MzBwTZ9twS+Q1QZLEYfSV/tcSg
UiGo+dzfJsOO4vkmJ2Zj19JlEufru7+TlVDclicNbQvwWqX7xa5wtfzALtKojgGWkjqYX8Ho0oKz
oQJE0cOTxvhqajc3fFQl+lo8KQjptGOGPHFNTmaKrqr+X7Eainr8lOCHOV0Eo2W9y9P8I5YzPGwe
eiLyycg07Gpwy10MRKJ26HtgeofeNgPdt+bTZ07/mdNzwJKMjmfaUlJOvwsxXzURkIkSxBC9pn9k
SjJchANT0bZe0OZSXxqZzR3y7U3ZZtotSV+KxiqBVkxG8mXoBF6rbrCbtYp8L7lASDkGznabh65E
ubS7svaKuI7G3LMbIqD5OrPjXyaFUCchMg23SlPqd/q7RkkrqMEcBhXHNkFbSITsVTRN2XCuNTfJ
RbWzjPq99rlqJSSM6OZQDZntV3/7nPjwFonIQLHr50nYmrf4x7I4C2v9VxvKDjJF8JY+Oxcy45J5
NLgQRlTSY4IE5Uxj/UAd814PjZRaqWY/jKfFT8YY7+m3+mYJhiSF6IFS8g/WMFXfxD7qMhCjci79
OdZ0C4f5jJh5qsmcwX3fOlByijIdwcZPHbICHL9PvaECzrLL2ijVmujfeXsyid1RHca6qXzT+TzL
WaeQQZoOapliHYD/nuh6pDjBwVi8Wo/GrU3uj4fnHt6R5lb5gz8rpxN+sM1eLBaBeo7OmBIJzbv4
u5BLVufSNFxcv7Fj5IOUtjcP9zFt2rDVKrM0OBRujID5FxydhyVMYrz3r7xyVL3JtkaMbMNStmr9
RJN2oc5ZSf8VnovTTzlosB1HxaDWapo0mzPyrJrvorPyjISspqEf0/v92h9OH2rPsKReKECd4kK2
MfVcp/pwdJpNgdgov3wxYfBoA51o5QtD2Uw0sWM4O2CIhdnmQnX+CHwdssFpPnDbBqbwFcklC7h2
VvNPRUUbCSji3Ko3Xvn3fba/wlpA/YKPwLCqGqtlcetV7WTBGeXFj0kmiJLXO9H57vCimvLOASlx
pxtJpgImhbN8qDi7CdL2koQCQnGVmZLEOyfIe6of4Uwvkh+tk/V+Fetjskbt17EsF1W9DDsHqdcN
wr827Ld/jEQdrAXJJ9uMMf7xDC45ZRxeHr3txvfR2wfpT4xMbDU4Yaa0RiTimAorvMd8Ry1MUS27
rh+iuf0IUjsdzpH+CiP+LOHys/gOZV5Rq0i8BxUxmPO/pQDoIX4LwrDNafIYrBTWAzPUzvm8tNaZ
fauQsujyKqQhDjZgQriRmefYxF8hU4NLw+xhPnlr822tHpfDEimyWfb/mj5EByg7+TKMU6Y88i8M
Ys52bQDQIMcQpUWn4gbUm85XD8EINyEvSaxf4BkqzmpkIsZC46ekOkROe6NgU3sHHGmmJrBbBlRl
KJFgESgz3mnTcF2d4uc09xP7FwEW4uFSTGtRrEdJGC3q0fOr+XK+/ZCw8O0/6YzjTcerCNlDZD7H
wKfpobByW875yOmLcdTPCEyIwk9XDHW8M/WHqGwgitp3vTrWSJtG8fVoo0Nwg8n2UnOE/x0L63su
M3IP6oo7dLXBS969d4tsO7FSEbzEt0Vl/gyMRxu3LrIzt4IdiNuMHTDj1lIjpcz8cr2dGg/LCc4c
M99vk/w6+TPWjc+s54nwqNzncKVm1bzoQRFIQPQcxiB0KJB6VfO7cEM8/h7rqUdDgme1E/pOLhMW
gTA3SxyD3fLs4s/b70kA3mngN+pCkuz5zvvTTlT1V/uGgG3xxqwvVOJxT0WX5dx2e0PR1Ui26QEh
toYEq6zJhjEhSc78HeB/yrTbQsIfSyYh1EwUSXOeq3BcA2kzELkNGlNuulfD5F8cIJhubXHcw7cy
zHtuGdkkjjtX4BmXthZNrtqh+3ZsiFfjmaG3rRkD2M0uQr0ofmSHbTkiWWsX+Hq00XgDizFFDxqu
zG/DmAxI22zMdGnr+hoaCsErfa93gYRnkdpVHyZqDQLq6v87PLZljTnFk/kEWdWyKb8Uo1JtT7/B
gKUIZgRwnTHM6ATPPIhPkZi7mk+AFawfZSpNvnE3PZlOtR+AuBH57YuiHsLSQqEdHc1IxsXzN/zG
koznlV6+FIhTf4vZXj/DlVG14hMTUzq4eUirLxzL4juTOlYrYRf3RJGlP0GexFusw5sT5lwTM8Gx
XBNimgBiRS8DEE3twTAW+cUb/SD7AogU684RG2p+UOoTFmwcaCwdfYa0+zNyUHyfSwwTWyETwpGV
wD4w9ZyJfucE69tQTXWKjjDfjz9HBfplj/INTVMRR/vfoUDcr9MT2ziMA+pd+2n/K9ky8dHYtd42
fx78FSg8AU9kPEOb/tRtB5gPWEUmdG+aPj6JC89a4H4XW3iaTMImQcy6gZerjYZhPEGb3XkVjTvy
DVjvhvCYfiJ8sEAjaPGdz+Cr00XK00wxLxrZA+cx0aIKYFOjYNQL/q5AcnGPJre5zJIHk0PjiNol
aR/xRcPXxNeorVAtFtZqac6EZte/8Ml81DLjjAhlL3s1Ez0ybA238NL7gYq6mW80TByCA6G4HAjZ
7j4xBSj6YTT2qO5YzMiYjblsKhXx3edxtgf9SImeW4k2yejSd48wA/sZdaEVaKBJ5rFWIxcjXGMR
M8XEGNSpW+coZPS+63l0vZKv8dl3LqYNCu5LESq1Ch/5ltcGGa4x2N1JNsqLJinkSDfyLUde/6Tx
N6HPT3DU0QSywpKGkIk0KuZuTHrFq73Uorgax22QE+ReYgMrOoKtSkeNRlDJysR3dXCu3iQo/OLC
IKTkR/X67DPo9hMBllS/9F2CQaltULiKsVjF1r70yNQmiqILjuJI4g3wyUAoHECRBaZ29qh74Xcf
y0y8OzIGYSlCfA27u67o8WvUAjO+7w+pqca0AzuT8flXVb1laNoTDs+0paN0dUV7Z/nT/ZHVUSxr
ZpZfDO2oS4OEZmpnlpKvvKtHbjLvrUEN6L2RFYZVOnWt2FRse7DzwydEBDbNURnUBSJCZ1JfpX7H
ZH2rQINinnObuH94jOOEl1GYPBXqz/hymJ0JosHVAVPAaIQE3TEMAxMoKUr5MQBsLUzuVv2F1CFQ
rkFbHTa2W+u4sEHNov7JwgWaOBE0Zd8vRod7gYRsXW4hJ5sHLtGWlcYdWUimBgqSCA8aFqL/GgIC
7EQ1Ac/hWcSaZh3n8XYgVDvWnltXFBaGczrKw5uUEYQHKnWXt3q5iGH51nFXsv1QerhtCwPef8nU
t80Eow0WkgDJT/07q/TDFy4x6wbS9maTGEC0JY/qglbwBDiY3la4SK8tZZCNYlP+ckmnzVvjcZA5
7mD453cP2Gz/DwPp2yPeej9sQudKKNklh2ltwBSJ70uor6vzHX+WecN3FJsB14cEJJwMhKUeqAal
IRI20r+Q/CaX3fNOwJPuxqY6KITdcyTdt0prZfXTYZ5mDln149ZqLj2YWX7TannmTzApHKjE1iY3
V7iSsuS/isM4mGBy2djfVxhFOD9vEplgg0rGnboBctHimLnQ/JKq0x8l/tN5HTMN5kgKOTJOqR9U
0T2cT/VLNwR6RGu24AJ+isCPSMJBKqrtspQZ4uInFcOYFXT3q+rhT57/xih8dLmlAFWWEUSMJB2N
C0xKWOmtugexbp6bXXp6sA+0iB4TWmd3i4/vDK8bGZCTp9+dcutITc9k73iMOkhs1auBRpv3M/MF
JbP8NXbbGpuHQjlzj1J8o69CFBbTzMU3GpA/cyGIFdq6b3NOwUnfCYSdwUN199WsK3csyn5dysbV
BjW5GzlJzQpn4Z/r12G/FmUhcZisE87xp8nKaTWh6XNgNZSUCUzuZqs6Q5NbrBZj+nyzYJ+SYR94
V3llrnZKHc/mrydR7fRuKKCU2NPBlLOSmcClS65pl0ivVrlpAK1gPOLd9or3osvIbOpxGSI72yhB
IoInezgQvrDDmpK+dBcuVxPVywkBXH/Q8n7/q/A7k0wCDjD0LiOmlwrZ8PwHDlIqu0JgFNeYUU3L
ZyoLS59VvBR7eSTlsBq7u4KtltBA0yxMdcFFCE/EMWcv3g5IKEzznO9rGyTO5c7sVfGLQ5CFgYPR
1DecaxGBqYz3WnKmbJD7cf9UIsyibWQcCKFej89GsBlfNB2Lz94dTf7GQEZIrE9C4Sk/dwBLM3Fw
y39mYqiBevDruPzCSlIoloznVWkveYjck5LKEGIl/tTCcq5kCglCywVfOqHBLOkLtk3BI56n5aQB
8PnQdAQ1XQVCGliYmvLDvAyRj9xTTKr6oLXK8nLr0ByjGHxKm+KUt6jisG7l0FCtZceL7+Eol3Pl
kmKbGt8Ecyew9iPtjjilF8y+GourDSj9+eTOVWqmOA5aCzIRw4wixiBFmPe64UxQd57yTZMWb3gD
yAaGVUXHJilAytxAybTm98il2o5blmEIsGrBmHtqzUZFM4OqE0MFdEgp9rymKYCTJwKB8tWcg+g+
Ye5COJvr+kPvHDbPC5GTFKRnMdYvusJwaZcoDLodNXfe0UQNWmwaQ6UOhz3L2WR/KySCzqAe+VK/
lIR5mDPkDid8swcV/NPWWrQAeUvI9gfKXqK8o0SAgQTidDaBtcnEFbQ3o/IR+AhLefSjlIShFNco
SLaDs0zODAOCNwT0zwWUizZSXDW/6FBPX2ri+9eyLYC6bSeAadYGWklhK2TJrHpgF3EVo1Fu7FsL
uo5A/vIxmBxC6aA8qku95f0tnZMs7Qy4OjW7U+lCOiakaNY9ORSQL8sjQRMnnqp8zPYS1XjEVfjZ
3n7msbMjJ6wc+ciFEjHvYeXoBOwXMu/8YGFtMblfQunpJRHd19U/tWo6YVn57JxQHRtA2jxObaLe
1mvtTPqKjaib6TVXqaDhRuchMYkqoyROMOo2CEXO+MvF8InCBaPH2CS16uhIVsIpdv8pJmvVntCG
6diLnheiXke2uqEecBH8CHm3fw7lkZcPkBti/ggGLZBWFk8KZ0KL88d6jDS2O8XbXhttS30gokpv
u/9awHAoY9ubrMJ88maYl8Lg0apBUEpeLrwHVXXnwyLWxHz+7Qe6NIFz7czY9rNTOrfFudsuDfyE
Ym1Ov7+EE0hAwqxQ6Ci+hshrHHiUOKvYGIohGf+ct5EmXzdlDY0+0S09pTnMQuklWNCWS4L0waxA
APTugYIiBxWOY6lYh+w5iMGDMMnI/BplbHPIgGOK40JWMEyxyeqgTxMbbeEnKL8jHgHzs5x2g0eS
CPYy5nBADJiIikMGBVCpvhYlz8P62kMJyg0Crg5V8kHa5CY2nSGSg6l2vdroNGVOHMBRgqQj8oyB
p4Hs4kyEvuk48sHK8mr+ZymBWSvWY8x4nb1iZA0oM3xDMiDUNHHf/0NnTQAjz1aAwkLsaI3ptuvw
L94gTqqmTvOYy+LOiVjbgwkGeyBo3TfO0gWGXWmEcjeHVwIT5lEmWN58M45F2WVNKAwMssZMfenp
sA3YyXqQHr74KpDiQXe390OdX8f83z6/8uMgZxCTvLpJTD9jm8Xr650UiRRI8GRbVYjIhVn0awG/
Lk5/zkNFdbBKv/x7AM/tE0RplKVf0gPzZWv5ZnVeXsrPTGYiL/JuxYR4fX9umvSoQ18mejLPeoFB
Eo2Cl0Q0LXmgLKN1H1IkHoTpGJ24vVo7zPiTNSw1n9WINjnwJl34DJtUiki0PB0EsYfJJidhxwBL
2b1RCGAgJpCITreq9pHYIVrYTbkIPFfhV7UXrHhcwcTcQLyIgbWO0vapGzjhC6ijg5CdkCBAwsbk
lmXqS6DEXD4k7azVskvOeNQOTjwFe9FHWNh5UyU6ZTXOdasBYALN9NwbVFt4crjS0J9PoV5SGfsR
gF+n4YkE0EVgB9FIntfh9PeTFk1DvQbV6ovVIK1f9QAQKWnhRDNzzPmZq0gFAih6Fh4cmaVbKgLt
L5fOp3iW7E9SkiovFL6ah9knXDvpD5Zi2kSD2aVpr7vYs0k3D9EKV3gjwyhTdaieaxMNZD1Pz7T2
7VVWvcs7IvUz84a+KcTeIj4m3Q0jkeEecNWqAlCtjbaf81Xo2wMzfHNvRPIHiqo+/agoX9Hj8YBX
GeJ3p03cRIyOoSrdgfiOrqqGq8dJJJqmwUJThwEsnpBagq7GCDAUZD1fN23vf7KrEEMXqYn4Hmrp
FKPqgak2t8yD8970d6al02glWt/sTqmfrjmDTc/LLNEa5SvKNB+Illkra3F3q/7r3yDiwjADRy9o
yUBPcycsfTme72F/zbzR39mI5MZFR3V6ejYg8+l4FrUexY/x8bmwdYJj+bJ8MmfUBGN7Nqr3jq5U
FL9Z4jwU5bJ3sPNMN3QUznFTRIl/ZsWf2vpZ3Qxw9obo5JhLh4kCtGL+XzH2cywev7+AbQyn09Lz
BPWj7zgoHeQHdOE5tpdDsVgpIzTNBBLsPnUq1SoN4vpvu04r0IaXLnY8RkkOK/UUs8cMpdjQcSNk
ot9TC+5xnryt+YbKiBguKCGae94X3y9kvp9APiPopkkfPUwJ2cEHQjC8Zf1TBEGNl6U0gIOR7Sse
bSHhoyCMK2W0m1CAj0ByrHmVFLtK8ycstE4S0HbE81KP4xt8MJYswErL+8j+UvHOXKzWxP29CJlQ
IXOlA2XKaYZS4Emv6DiJgTNBcbK+/dNfLfh/rZUD9mXAPnnaTzZrrEZjiDfe/yo1fKu/f6qOggo+
nY+nPCEr8n76nLWH0k3FW6QQrZah/JRUMzFfTQxYhdmdIqU+8P9jlhVhCwVF4DjdH/kfreLt4Y1F
Oul5U+wH293AImNcyFymDFrB++bMoWKUfzAcd0D5TRXj3qrEgEUQa3IdYlbs+Xi5vRZiCa/qfLgw
vWsKJ/esY9qdo+QqA5waX5YRHTXtkmfOmZM2aIZVScqd2hq3dliZSBkTHfBOOi15rO0Te44xIRm4
BwjAesEb3lmwhwJ8dSp46vwpbjAyTP1E/ys2y6ULwcTp8yXf1Z6gDF/cmG+a6xZWanpn+sWbTbKI
wzbzet395eTJkGNWBtFjnfOU2Pr4Qxz5RxqY+eWI4OlfdapMclmCNqTCxg3wpvSUFqlBlv1ji+qf
RBo+VLergOcf5f01szQUijqBAht9t4YALWbR2PQOtfQiosyyuhR/LgzbzaNf4aOBSRjc8Vm05TTv
+WnRGWiKZOsTKCEOP1Gyp1CBpfbOQ4242pQ/u89twESlRFV9Txmbjp2x8F+a3VfyfWqETEL1dHR5
pcK/RK4XpTKh9lx9+TgHtvV/gPL0+bUIkEYwt/y6pNblywsP+YhSx6Jsy4EVv/63USMyJ2fKcFyV
CFX+C2rJs6uMhEMHYLa9DKPTlJA/dCBfi3zhmYtXU0/6ox6B5W7Eh8NX23smiel6UNsavmT3BvP8
9ByJv+ceTG63frrsRp1fZfkfoPZngo/G14pslrHjG+OIheqeoymhY5HIUb7OChr9i7Kk+YCp+uNM
95U2pdJ3WIAGucLfiDovDSwE3B3td/ouO9LynsO9TDIoRG0V1UOGOF5aQaQ53T/+bxeW2O3uQsUG
PCifDTifIuIdh7NePJYANEBTUTDttGbpfWhZsao2tCnC2X1VUJUF8YB+kWLg4rSWtBpPKKXAsRni
sOaVl241iLHZ7clvY8j40tZepBxM6+1gb4F5MbI3LmnG3E7GIEeImS3oUo3b5AuR/ZQXxfausgAU
oSl1zX+631RiMXlE7+g2d6T7vMPIzM7UXgYyolq4kGWRrlUnrdyfFVXzh0vdhnZ179Qw/bBtqXLw
mzg813SBq2VXeD8wN0NwtHBUqE8haaPDbHmfL5hi5SPonMtTS+moryjczqoPKzoqZbYHKYkVCTEn
edUUd3ZxxpLqKn3LW5dp903n+vlhhHYE+zCoHJXe+aI6p7VRLCp1anrTBB3ZsRdbcxSKvtEdOKOb
xVxQockiZwsLFrXmzspF0q8aWIFu8zCNAmJYHR7AUuRMigQ6k+62zukljV1DrXw1/ujv2MOylb5D
XOpVfdJD0IePEb6/xg2dbB860h1gRxM7RclEqDEGljodlZum2H7OzC9KXtzNpvo7laJp4CuTIO8E
7edSjYJuihh4/sGBlzYnAas5Mg8tuf/UMyxtUweja4Y3GZXjaqi1LDQyGICbqdh7OySp/uH3RCDp
HhSzTcqOzV6ggIBWLatswJxXYfV6A0m2Fh0WWNeQKkQhsrOLwtZmZPiXuhtz5fMHTnU6SXG8O8XU
+eWvcdBK07ADLHstKiXctbphrPZf+zkQCjiXF6kV6ICp8qfV2gyk7TKgNMkha1vJRjMV03ZZTehu
NbVZy6vLf6HT71ez+q5XCF5aL5uljDkMpb3lBMzfZNYqymSD5qYU/8WrW7zLL0UpRpygqxfXus5K
p8uC8+gzVX4TVFdO/lWXH5i4bEb2jCZVt2uiCScPTmy/i8n6W2wZOvrFJ7kaO0ye9ZywfJU3JBLa
UvLGsgK6Lw21bgxjZVMpwaHj8RpxGivFenku2rgHAcJZzCdDmg0adc1nDRDrR4M/dvsO29Xkj36D
HVQL/b5ykqen3ee1p/EeyGyV2fLUH4WJVYJgIjj2ZXW3a27kHkjTZVajTWOtRDwzhJyTAwDuGLFp
kUNDRI88iNEVK0o8X0szqytjXWqNnS2AYPvhzIoaZlqTEZtdymIk0ZWZLft2DSf/8mGkjEGa58F/
4VU9CwqKv9NLXyF0CxnpDXl5pxc6mrEMCwBbnGdBnSDiVvwbLFNXsSzemtuEYRG/Zmc4QOouYAmm
t0sZZlA+zY+Omnkzhj0Q/9EJKX/vWxPR0DDvww+wurjYVWd1tHjoB7uhVpT68EFw6N+wSR7monOF
U+4h0J1WWvzoOkql6SvgZgQZkLAM1J1FoDELjs3zbs/z2tHHHm6basuOFOkGICCeTFqPSNoJD1yR
X0IgnkJXnt2mIraP9LLkY46Jp5nq0A3pboipGWdiS7+Neh3qREIJfcHF2uxFyUlSsESMfNW2BURp
N2d/WNlgIxYQXpNAfsaQ8UugSytZWMIXieFaqMemmHuxBL5a8q5ieeXYIInw9KMe7ORSaxv78IL/
tjv61H2zGcK51NHgX7d+9zPb292/KE39F7zADTSYb5q0uZaVovFPtB2IxhwOy8Ocz9aKmhKM+xpU
hJsNnFS1F7L1s0Cx8w6YZ/pRa1ANc2Ld8/bhFtLVsDTpJEeNCFRDiUZHr+Os8ypWDKxl+O0BlaDQ
vrJmZC/vH7nUgEFHghwJy/5SBaKf3Y1rwu4bPbctaiDLYryNgRH9E3zq5QP8KfUOyHfAXDdsM5ZY
e95i7T0KGNxWFAZ90B5WaP6tH2xclMVt+UWUItD3LBcOOU901WGcn6Jhs8z1/HxSyLBftmmhaTPR
nD+4pTWFqgInAsmE45hhOLiZLi6iSYoaDSm6HLzrLsve3xZJ0AOux95kXSUpUVdoYwzJbtQ5Z2yZ
FF2aVo/MPtcLqGNwr1HBxCX2+jzk0QBBwl2DYbPy7yWuHk3skkgqsEbyUINe0wQJGzShbfn0RXpb
YBe2VQx9enClp4vANLMzt227TrUgiVm7ptLHcGA7HQOUSdeh5EC7+XEO6WIBQ6QPLMCOoU0Rr9yv
nO3z58PhxcAFn5sQmqf09Q6dBVQWV6aosg6q9FJXDy9Ci3Tuttk7qoA8vA8mOKm9XfC7J/mJmEYS
jA4g6aZREStBAkntI+b4+GcjjKSPBCt4T9BLhtMO1vCj1GDsT7vvPzVHTemd7O9UYh1JZbQXVuDj
0bu5GrXQbppJsHAdXDcGOvuhd6+ZIXAHaxlWWvlga+bZ0E9KmXb16bBCfWSyD5rJuE4ZOS0raJDe
n9ZzuuIrYgP1lzQj1ggtUTsSAUiuCsLGOMBKSB5VsEHIwO+25vXD2vN7gAdriMKCbN2G7yyOPVka
nc8l3XltfnDryTDlV8dOJ+O7M6IE0qCQ+d8Il1qrBEQIS7fSPB7p1i8tD3EehOaZ6ZmxnyAYp9UM
Dyora9J2NOkBDv2C+J2YrM0EicGWIyHVl9QNRVSczkNgcNDX82OPZVMm90mX6sj+flAtl05i+NnP
bKXDZy+LdveHlGZPWO0fYRC+Fgq9NuVJfDGLM03G6cAVWUF3AChK65L6KhFhu2Mmt8PzQc/ykNSp
tkZmGvpxUPcah8UOsRbyFBZzQJ4cj2Ec6eyozi+Bo2nTVPe9kUc57fUiZgx2LtFwblOuHP58216f
GcaBWXHzzIMDIFM1pQH24tlWiBeeRlogDq58tHChEUEMDy089JqgzT25c7hrzxw56Wd4dzUemaEH
KnAvz46v1Tx30I+81s3xkSEaazTcVOwiomNBOoljgTj49TH0JzTYs/EsdeEqyZUCvO+KVN5KX6xE
7KigqIEC239ybJUsUIkmY1h6QKE7cezp3VB9ZqpBmYoeSf0Dq4Emw67F5wTg4AB1IhLeRfq5RtDd
9rStA/CaADnQasGLY1uJG7A1O1nd9JZiq3Z7H7mqd4WFZkabwn+Ysn8KxB9UGDUArY/Phv7INdmH
cHGdn+4I3RaOCcLu31kBI0D30kSxs7QzCoYOxpzHXzImI0UCaOZWehDgWy483NEVsdQr+OoWqAmO
tCBGJCn/p51lKll/h3FrY7XHpEt+9wCXhsTgIaXvUCR+N11VhsT5m8ICMdMNj+KHwG0HP7dlLyus
AZZcnv818yBh81GJDOn+6pImnpB/q9gEF3UGNVApl0N138REkLNG7sws/ybbb72eEg90z7MmYbY4
OPoaFYsWgRQ71LNiSVym4sx+OUb5h1XsEmKOMBEcffP1aOyWkDhtGqUzZPB7dD4Kkq1ANtGPKmAH
jf62u2Fp5fv6cPQ+eYZ53eEJHlWWLSO9CkpzUEcJ8+xnKvfbizYPF7K3F/jQKcBuQE/JR+IwmXJd
yNQf+Zaruscur+1WjnmidYbpQZgN6YAYJfI3RVhhz6dnvXlyRnWSqCU2EQhK1X4yqHqlpPXcTJ79
9twpDht5TJtQwQIQhfw21ERQIVW+ASL3FKkun5HHZgNLJuWgQTeD9Fa3smx5ObMeuPgOxiuC6Fbi
9m16VWpXCPuQe1T8WwMpTKMVwS21lQs3Supv74sjQnyfgPdpK9R7Gz7PXeyLp7UZ4wFuEEfJmMUG
lbzZDbdrEDGyowxV+PSJe9k5v465pjCRJJ99XfCyTLoG3w126K8vWmE+a5tM8oCPMs4NWkqV9+W2
CiRU2d29pwWiMWKRBdKSyoal8iTTw1/cJbQOALJLNG2jdPhQZlXA9tUGUNiiJYVhdim9TgwOckgf
J1OcHE7kXE4haERz+jRT+2LYSzNriK0PA+VTIaThwT9B8S9xkumX16m3/BOd3jKAoIpz4RW4sSqf
zY59vxc1m8saNPLHtxgf4hC4IatmXK9M6ZI/rnDb0w6EiQSzsrwq9Z1Zu6SaTXzm3Gq80wFC8Lz5
Yj9f+I7KWQ8UYpsXwZznN0N5dnExTQ6yWGmS8S9+02psqjznaqWrZMG5/d74orJgP5VZZaPWDvxC
ZJdRKcLiU/OaAEUnmZvhNXCxtISBIa5DKgMfjeFFYfx4WDjr0RbT1Mw2RcsyMe36+PHAugkb0v8U
iCH4pjQScdnVfSjAmh2nH4IIUGBxQOuSqds81W/Hk+BF7NqwjcdiBc9yFCeuNshwJL0DP5z2xulf
ORdO8IUiKPTyMX7PaJ8+3hPh+1+SQNFwkaLqGYLxVL5g6p0Z5d3+f4m+kfVCQDVaRA7H1/LU0luM
1HkrWCfFEQbXCjYfoHjnCPaB1aVFLHNYR90v26lCsiBLbhxutkGsy5T8jTfu+zFwJ4Vvwp6gestP
4dY+4Z2OmzJUpfMuoG1rDcxZbObYS8Np5KJIZvrj1oD/X+7/50SIFohnGNdj2564qx13wRQkDrqX
EubK+8jlXSfQdpNq4b/ziqwxmkwXCmXMDbQYrEO0Wsl7uCg5Mb81+gy5Z0lcRW+MXwZYyqxwaTYx
aMI7uXT1Q+02++BZ++muUlqt4Zj+18QOaTlJxm94xG95scjOR/pmUgbosfNM3gau2JbzVe/rs6ZK
8IIfr31qDqWvm8f+iyCLa8wnccnNLCeyhJhwat6x5GjHo7FcLkrJzdQfbzNVRXkW61hRP2PlzFDu
AXz2sCQtP6ldvwIeOdHthj0VO+XIWpSXkS/VtXoGXMvKmFdRDb/UeSjJhlgZ/jf0oBszRvGveB9K
M9GuhNmx6NE71LQ41onHh+hRTZpTQ4yw3tMS6BoPn9i12IG60IDBmrw8+yFgRre504JOZA/IbFBO
qkVcUITYfskdty1iz+WfBACG/hQ1c0FzIoC3OTBPxZnKluereSFlPY7RLnEggwOIlP0JzDZ4hS4e
y5Xd9Ox8liSay0USPx2ef7m1Nj1/XLi1sLpwR1mCOPRQd10sp1P/kb1VGtB6hFPCiV06nNk0ciBj
zkY8NPyxutXpZ5rQedV3Ro578VzpkxKUu+VZYn67QLdvRV2uFjHwgl+IOM4Hdl3T6bxiLREDXX7e
VZExng1zAZfnNrrdwFxZ8Z2M/jv8D9gxUtqFCQu8Q0Ze3UzYRWhvgSCyArVwpYfWsAoSo1O5ni/z
WqJrwDHLxOE6vTe14b7oMZE9vJk2Td3pzzzYWdYSBTtND26v/Nqr3ug1+jUK11txkGc6+I0AQRSc
NagWKe6eWQfrECKzrpjBhRK/3OuE+fCX6XsmPSvWgEqJVTddVifraBLEvFt/ayBJXCQZ3XQJNRGc
lKju0Rz7oaJpvhgpj+m9T0A+auH505+ilOv6LczK+Sk3qFKd9QS48QyiMjd0G64ZFYPCwJbfn7R4
uZYM4pNgy4ZgbzWYe6qzt2MHIcfsAsIuOOlik7mAORpb0d3NjHy8pvN0zo7XJBcdV2VQGQIAFDLy
miI5yedZYiBO/SnHGVFjOAWv4V7ot/4kWO6XnMR4t/xPhUvRPQnueRz119ol6WvJ81YWSjV+RevP
wzmBOsQMokaRger2vfivoJfumANXRV6m0Q2+KygNR5Cu/lfvsyb9fYin987qiVpyedLCOroyRLSK
yrO4GsWInSjh+7G0yBVMU3flvm2mUXzQ3M1WaVIoUsTMQ33tC0rbbUFK+w7juadShOWkgJZB2g+P
GjVu13zNGzC/HmfVlR6Iq5tcD/2W45M+plLSHGQClmch9bQeqLwQNnz91DmEsXF7T2SFN1/QzukL
7CGoNvUpY7Nc0TuUVcZiRMfAcT8A82iO+VT8bvyKfv/+aHL3V8PTYdXHN5NG/CaWB+vbvgh9LCET
YxGdv+eUhOMyHiP6cvu1vWzvS5uTXa1I+llfyq0g6SH9qbEBFkP2w1zGgRPqIy6lLjMmmFgrhdXl
tZ6i74c7n7WhI6+Mi32j4Gwh16fdsYrtfwZn01FLWh0hwOSn7on8/lxqoeNE4vgKcEKc439dUUCL
4mZRvoXXfVc7z/TS+Fe5ztU9Fbq/RGm0ezjYLesGSsHOD0aXhhsyvm1D8MueP3g9q4WXIFS3XOUj
o6+KME6y4cRqvQ7okPSp86YnL7LW7sdSHUyeYZyNRvPeMAqKzyE0L/DYvzCjyITxgYALI37OJVEb
FGNQnEoiya8jDL0a0a78M4gKICzwbjKVgJZBjunIe5LFRFKePg6KdMPJVOpfSVjy5y8lqod83W7N
KCzRAOKTXub/RzsBTHKWQiGtTYk+5aRgtVZ1k5zcEDoaYOWaFsym504GczCT1HWSOxftJo1AGHfb
brr3HSS0sr7ZtHXQCJzInyaZ7/VNlzimMQuPm4FmWj/zZwE9Bl0DVZ6w2Xy+YQCQ8U8wG8f789s4
6hsD66zKlNynlkhWMdS50WFOP92fL3syMX19RYdiMRM3NQZBlsBvQLpEKhWcorxLzibDJkJRBLmc
3YYRvZM1UXZTuPTlaJNV/0385qq36mNrUgva9feyHBEoqjsErm9pfCw26hDX8+GE3/G5lDbwwt2e
j4H6Fg2V0bH5ri+OczqyHBd6B+c7maSOltvS7c1jJTaCZu19lr+EPDsb5PPU6xgPS05B60eYKIF7
I8DltG6zXnBLfe//0KhRTSV3XhVsg1Z6+2VWlRti+NTmniPCchRkzCsTbrcH1D+rN4nIvJ2OzuDG
9fPpPityornJLezGjw4TRQ6dBMt1K9v7/S7iVfL0Tkoi4vZvDp52YubjNR38W8m6Z/CPNvRwh/hm
6K/ZVzzTG8wRXs1tcvWCzvfEcDpXI3kQtsIYzFqzNNidoaYTXEw9D+MOOWtUtxLenDeclUUFfgDP
4nOT87oF/yznFJWBm+eQ33DyBS68ZxZJPCVYw1Jnw5RISeUNvrkTaZQHuQ6kJ/Jn726f50BlryDc
5AUGVtakV5QyNZYh/387b3bSmSBhvrXhrLR6oiDfkjDfZuEMIAwsyd81swBdjUSNmq0/Vv8XhdkU
U9i9WMG9Y61qlqixHR0mgvtMnDcN0I2DPRDnr1VwCUiOCnxaOl01+J65xutJ3cuEabYX/lLUBY3P
o7E+Dp9+iTiqLgsFqiRttfHaMnDdDC+TcLBXIQJwVo0jGAxgs5OrjCKyqbtU+ZVA2913OTqAbh9m
5cHKA78s9TH+B7A6WhN6RrM1V+fZcRslqGNzsjjT/13ozIg2tQVoNI8q6r7iygJi237VIHrOuagi
axbLWzdwKRSvH2tsIQ3asQQTfA7pPp7pLcGFHsJUgXrvPQ53CuxawQn3t+4xp/evVAeQMTqnA3Xf
RTsFHtYBAIfetZ4hKBrWllRfMF7o+mwc9qTF+lfcP1jES1iRIuQf1/mek5PWYoDUm5JrEQoJwpoq
lpd1aZ57cHXXgJa35hTyb/W/A4MU3pn/vwOFLwNAu9vcmq8Mg5Roh7Ha/0x/99Q2fWqReoZ65+7A
CIIg+PMmWE35tdwFTplBLKW50GxBmhoNEkSP1s7k/HCaryAc3y7yk67/4WExG4jMzGfnOas+Xhnb
8HaI11wNsIAEu6ZrdRl4MY1nhLJIFG+ikBYjdppwYmwXAn7R/zmmHTMwNDcT7x8h69aUxxYe+BxO
n/jaak6i8P15UWBLLfUTY2d7vKdiudswJkUqzJ7aHCcnKWRji4ORHLXlEMLkF5ADdpiBKE02wcCc
HJ013enAWc8ZVnBiPhr/aBgES/Qu/e+6XrCMF2Bpl7Vp0UpkCiYXbi8dwDNkOy1K3trOJN1a0oHm
X+13bRw0flFqwTPWBfqyXJ9Tk5a+U9sSC293EedkA8FGhSzwWLbiEbzxayAkam46ZO3ouhfbiHv1
OlB2Sv0GQU3o0SlisI776Trl9bAAWu+DqC+59d4g2ovCMc4lKBgAgvIe0KA/4axzhlc1KA2XGtm/
JdL4YJuUwq5BF2j/u+Ovn9oG28+MFf5QAED9J4FEFXTrcVZuD5ttyUYiVKATwfmnRwHUmA2oRJOb
T37unQNvLpy9IjZz6Yz53UrghIzmpGW9YhJu1Ef3wVBTfr9571zncIFgsgvp7ZS1LKnwORKZcWnI
uVm0hp75gipcdKBw5TBu1vPZnezMe6qTKmZCeCrtCyTuo6CKep5mw6UQ3W7DCFVUc1IKBNAQJmQP
IFKXB6gPsU7JsooyjPQdc0BKGY1kUIOqqy6kFljb1LUMJEbdLcbHgsU95DARDd6wfym9FS/UOctF
/8Dv2kmSNGyqz3Xu91mLYWzfwP64c1a8geccHNd+GNeyWZwOUod5c0EdaXQe29GFWIAs9lr9CPZa
qWYZqv/Ay1oGO6BAIAzL+C1TWGTgq3euJJtPNTB8buBifSxT7hLLIHUz3jpX2pwSrCVNtG6iracU
gjuOiGBre8IQERMpJoRaTu48eXVYuynmDY4W+Oj1QqPQQKE2GeM3CGLE085JmFnP/4FCFKRPQ2JX
ze6crrrmosYTeiteM/ds4HYxd3w6H5XTW2jRRznvHMJqKN2dI2gT4e+3bI3kq1c7yIzjg/jnEME0
qMxU4bwb4u9h9u3wODn2rKTbdv/h+zpZghwh3TVKToz1VNSk9/NfxX6Mz6G23ckSdm8HqItXlJU6
Zqj58kdHlQhlIVV94RhSFOxDqY3OLm8lMKCmRIsDK71E4HOeIW6RPgyfQmUhQ48Ji9m6uqD033vX
bHoj+bdMsDey4y3UDjrBOYcIkITzrGS9Bm2vvlua0zRlEyN8d6oiUwsO1ShlObV9NCWNFJ7ODnFt
NhYGBFzNF/ZE5LRPawQadgZSy4kIayLcwhT0zsitVcEo+wX+/hrs0sHTNGZTTl1iTluG6gO7JEml
yfs2UZWPTN0pC9rgZL+OG7CL5lyoLTFWpRPuFFEl+OeUMRhSw4e3dkXiIyNrVZE1TEbvrEocTr/d
1/QX1nXI3WO7RYb3DHZOoB6nmdFU9ZSjEG8SZMkCUEO57gdpyEsEP3tsTXXAWAZ9hwe4vtSXZTGi
qRbGbM+REi5MkDf2Rqasy2Y6wU8wD5QOTXKzMi3u0RgglamIe6AoZJy/G59KNqD3QlQeBwUDTiH5
SEbZEfFMgyvOdAJOS8zCB5n2fdXL5xKNWmUpAiYrk3wmDzl76V3h4ALIYnmM5W/XanYGFjH5OUCv
np9iw28OF4cl0wrYTeXBAaFyvaleAzI421O/JpqxPFTNSEV/YF5pt9/jDCus2P94Bg0teATUszD0
oZ6aJG39QrPisBF6kwGsC5UK3r8xxHo/QDfIahD0eSNsbTFJbf67e6V/5+a8j+AA0Htpqw26jhH7
qN6u5/+65gkNjqtcjbzXePbo2LUmxBuWsw4nRzgvhqQkKvoI5NgJkAKRbOIl5vHE2F8zl88RfcfD
hHQK/7xo+zgGHkCzfHw8wVRU5xrtisoWRtVX0LZ7CeVUCYFqesey3Y0221W0DZ39Tg8k/haFjFdT
s2FLBk4P5YsJe2hH4ElkBOMdKMvqbyxdQ9QyJN4bPltoWraGLstP3fx0MVifstxXx5R7HXDe1/iM
oV5SqQWo9kEkdDRduWVsv3gQFVdv9Ta3RshMKsEE9BeGkHbirYC8AswmKYYCruOHXBRRSA0FtL+H
tX1SR3IS/UNhdF3QI+PgJHMXEbRKMiiQBkFpv4z1Dvdy/fJf1lxRLmm/bfCWqzkAsJgRLKhaAH6d
GYDQZanBKJ75E4sIeZBxBoIx57fSDwGJPQ6sZgatalPT9AVvSgVVW1Zuqzdn5eGHKOTnFIV62HzN
XYuPZxVYYYuiOVF1/nmwu1DqEengb2GieoQdh+GOrDh1K5YLF65gx1sEd7L0G77DsmzmhUADsvU6
ONjNuy3JcvUCFtuHwtXNzoYRX05iCQkwRTHo/1fZXaquZIKDiUDRak2QGwEEt8wg5j2qh6KSnSOF
gkBJnf80mw8iG9WCWXjC5t/csHSBcNOgTHuKWD0UuUhRUpI7AHwG6M1hkAbI3TY8kgB8Q1UeeJbI
3IvhZz9rVSghWMGoWXGZIE07vaNVfd+YN0XTY2y4hGi9Y2lNIH57VbE2ehkS2p7rxYdUVKQOB6XE
76ye41nejVM6FFbGywCAPFQYRMrgvs8PnNcHNelltWq/h5H4va6rsDnt+tkHGHw/HPVIqnoL4P3s
flg73d59KwZwW7DPpotYCgPetF0YNcBPGwnWNSVQLUWxby6rZwDMdLzGBwYwV//B2PiLcFQ11Ak6
0sGgLlgq5T6ARHhM/lv0SDEYCM+9+FXKlOrNQN0XZ+lkolunXWDjuQZx4olRl5hbL9AtOQFSSBeR
74ks7kyTSrtXyE+pdA57ys6Ha9cy3hPMSF5BefCwS012JVkVvJSD/coQ9B6Lcs504q5cFMp4RP3/
ySJs8TCxl6iACdxupQEY/m2QVachBGgpyzbUFhGYkInF3Ne0YytrHzUn6/pvZu1MqNsaZhXQqRkW
65613CBrUgpqsccdz0YqoF9G3J6D+OiJa+LpDd/xNMkOMBb0IxgDOL4JJ+2GeM/O57+pN2AhwSH8
W8YldVddULFrERh2RQ77ACNDzdzixg80fx5X8tghCYTziD7//8pfecM5fdhMuQxCajBKkkuuYMak
PPfnv4dX9+InI0vYQiLECb+7+n9gHLy5jrOFXmSu97MmJZueziIHbPy0ehwAlr/cdKCzjtVbHNiI
hK/BjnQEDVyPLXeN26GZLTOD5A8sbm2e3JMxBLETorQpJ4uHjU7JJSdsEa6wHMIeBT3Fcv0rwbk/
/zEWZx0hXDY+HvDJl7iJxfzdX0FGq+8f/BnXe2xWoYRT13ObuTWYFXb4GuGicKYGs2541RAlzMfI
4PlGX63QcMjJKuLprQ5C4whP0rRxKFQyLvEoOwCXxlVQDldvITCeS+t5eNFPf4pUPWJnJS6WPw4i
RSowE/9hKfA0zi3qzEsGNkYKXnhVxRiJujN1uXfEUl80mghY1fNBr0tyNBvnKh0Kur1yIh3btpO5
4yArephYvrbDPOySyFXGmSH/MUW7XI+xfTw3TY+OGGqh0jUELAC0sEHkSfd5yTEt55Plz1iY5Dpo
pBD2UzTcYgUogxpSmkhIKwQWZJ04q/3bIzsKoS/16aU/RbFUI3u9vuekylffLPCDrq7XvhH9Azz7
LE25fUWij5h3m1rRxI55w3DPDQnP01paxIWzUmnW1KQOLOKrddFcD+uOE8bEq7B23YL5cD37txtZ
F9ztUY98v0T9xccnpxvwMAUDGmp1CraU4IU7NkI3Fv3+QmOBmKl7d55AojMYDNukfWsPPnx41A+C
JoNFQjzIxpjBvn4G5++lqXEydAPgsATReQKqXKQi2n+sZt+JL5OE7SAzzVxWkv0eNrvoRJaprm+j
CB7OzFWEGtK1auDzWwXIeBTcf/M9T2+35QicSupu8RRr4I3DQ9Zu4hE/t8ugkA+DlREgUNmPtviY
IeX3MFJxOWBjRgNf7s7GYf1YTmjQqlFiH9V0/gqtzM5Q4ihJa3agOhrpyT/JaTvujcWyCcPAFzCN
4THxH1c9/knoOUnW4ZcWfbyMJJBJVyWTCarM91tMxnd+6wHClKO16RPrpZIaNddEpPQYDbd5ib5p
qkVipvjHHvMP0euQxk5VXvna8ohsRxnXd9gHmHu5aklbkfgphlqsAXKjqdSFy5e3hHAXQpAO0sQm
lEoIB9pbgI1RmdcQxPs3L0dWvdVGpVuJ1ImMXgq9ZvKjsubl01i3qmEx50od1O6VX/yZwQ1eufsw
3Ys/QW2clEVVgIvr+goUJKIz9ntP3XJGyBJ9sc3nvvrtaSC8GU0t1PrggM7kXnKwnjIY8qeYohN5
VZBDg5XI5IHiuQfLi488ECsTmZXflJvEFhO0ijRfs3Uq+pB7W5sM9Xlkniy5scjOYWbqJch9pNq4
5o2nzRbjMP1e6BoPbR0rKTMqcQ0wxAy3FtU/TLHz/oDkFxma03mDjeO04Bp5h3UbAf/XPZ6eW3Zq
jCLW8PkneDKnTI+2aOCfD3Mm/RfMdBfYo1Sxz0jyRJ5a7nZuEvsXX+aWfHtJwq2YlV5I6jC6dTYR
7FJOQ0V5nViXYDtmv7vgAxSVL7tS6mN+wyRJ6bebHoAmA3bo4ZfTc2mm3LTFFcY/RnWWnrNQqGj/
m3TXeoVmMNb6xuZPXM1kBbnwH/sLiXFFgD6VmFhA/1TFWOL0qSSXNZlSZuBZfkbLcJJlv9k+Stj6
SDgJBETQgoe6Aju/x4M+N+5wI8MlOoemcr6SsoVY0cjFI9pe9PcR4qKmYC03YfNuUWL+Xt26MnpD
z6FnMokbTIagSNDP3/QFqCX9aE+xRuXo5jcPigksghrpApBxmdVBpa0dmadG2Cq7D3/YpfJ2dqA/
A2VaLsnNPfzozbhoXiqJzDj64oCtC+pIjqnFZDxg7kOzXcLy1MTK0dOdPvoTUP6VruLSi/d81Zw3
1Gq6tgRF946DZJ8nR3NRumrHlOMdrVwIQVdJhCBIW4RNBe7TjHAUlbwWG6zmv5QoVNgSB+YTPIXt
RYHn1p+q0ieVovJ30LWmf7a5c6yBtyNzSx/dNNpCo0ypffzbLxzrrnTLO7f6jiPWgD63MrWR//rO
U9hooaGbGY5XGhyaL4/rYOqGS5v7rBwRSeSwKLePkj76jJgV/5NKEXtf1ud+lEAHf7BsFtqPnQSl
xf7VdBRfHY1ryum/1awhxm/LKWzNjgkAe1kjpPLWegCS0XO6IJ7ZzsDV2lbiK/hvhwRkeAK5EBo5
UGiLyd9VuNQh2Cowt3+9gk/ZAqH/LPKjVhkkvZYTiG3XEtJYHM7T3n+/fxF8AO+ryhcSckNKVMMg
cri9ZfDjTYaeVqYatLE7tTc3JuU+fmTs7VjsFAJnBbZqQIoyd12HpLwp8ImPtl5/zrx2gxTB6sZW
RqYMAXRpMdn2TL2G3P1dhFstqNEmOSV2wbMxTvbPosIJ2r7mEsfa507FlOy7N+8VdcwZzsu7fbX+
RqS0BQT/JVYRkImRuCqs2BvO5hQuhZeDiPpg0VVLcBDUsiqBuekFlwqoYu3V1Rc6MOaMze29GAWV
3WhoIlbTK5SZ6lpL5/IjOVmjlgeJYZQmfVNfeZGVG3K04WvyAtBaNblVYMyKk/OyV18JzMNADwmg
JdvfAb+GuF2M6awX/PsOlaohHfQZZNOKDry/lYOwYI4ojmNQwdBLpSwoYthAzHtJPQFfV5v9xDe6
F1D9b3g24uwcrOJzbND9kXVws4MeGxpMa6xYsExUAQBqRYXG3PrqIIptSqSyn6/zQxMhrs4ZBzFd
eomHudywT/0ftfszrfylcmD9w+FPfRyWEWvJ0y6EpDYxfZGXS9FmalTbyopMUzpydUz6E7vjqOAm
DGT4xX8tR0YLRvI/s9C6KGWFPtMRWvWJRC7NJGv8ub61GLf9HuxCK5Aog/CNs2iN/wb+ee4bSM8Y
rk/OU/M72IpN/0GzWfw+CYEIBQHvZ17kUCdlLDPlvDUdnb+SLy5oy/YmRoqobgIshO02XwR3p5Vi
2S5+fpTglyaDHLzXJ4rgwayhgEUqMVixSV+ZbKjijHmEQcRbdY99NoBgBlZDshKk4mP7KkNcI86v
9finFVzkshSO6ZVLeXupojEwevUsGip5hewM9Sw+MB0pWfHE13u0PAqkdKQjV3W6cD/H8guDVnHr
ncRKEKX0j2UuL2WhlvkY5yp9zcLlDoACOnCdLHXFvQNZwLGpws26O0guAKgoB3RrMVL5maeB0mFU
Gzz0Ulw9bmcysSIJVrfCSp5u7FeFsGiarleVqZXdxJYt5Dsgw6ts7OuFdF+QQKONJ5cH7MmpkYGr
Fq+ZOF7aneEHFrCcn7YfaKRnPuua18DBCAWtcF2xJXyhaseLq9Z+P8qN6kdPAKHGZQvAVACD+eak
Pz69Cf14B02XOVaokndMCrBo9ttUPcIWYHC6nkYk39HB+CT8US8uD/X4tC7aKrVaXEg6qUdJGB+d
dJ0gZRVyqmtfxZJPKzXVNxtUu0laKEV911n2UCaolfp6wDZLZLL7X3I7+ft24SQ3RJRg1Bc3prhM
luOxa58STXYBaSB80wY6mPuW1Q5m8homK7tK7pwvE8QiavD7eYbinB+d1yKrYxpK5JT38p3yWPfv
H8U4SaCzPSUI+zUl2LWCZNr2pccQkhS8l3PBG009jmZMFI2V562GD4KsXUfkgTxRj/DQoQaIEIdZ
97re6Gp9EI6nFJmWhiGJouXXTYno9dX1KlYTI8XJFwfBdEaxTJwXXoYUIaKxr02lwV3UgmdyH2SL
OffdvQvyFNC3Xyy7VWNGVx/gr7mj+YakDirQV/yNvtzE4a8NJ1MObL4NTGhVuNksJ3Ri7TE/6Zob
oUV4vH+rZZnttHK8RdJEAdOagUdLv3xObkK2zCnBXcLoj4pk9BFJvql6QqYZ5Glg9tgAg58SevnT
svzdBsvfioHwpc+8bbnAdVB/Pc5La2BAizhfaWXVdAJk16anhWKF9HNbJeVTNtnkW4FhdUfn4ViQ
ch2h2vIb/oZUNuGAZs2GG2Gx1RDf/h/ESi1h5e61xaDjAFbck1a5o/gSFYXPGuOlVQ2vQ0aal3Eo
542QlTUOy5C8GcvHrYNWVe5ukqmOsAEgkr5k3gyPm/0eiDwfDlK7d4qRrMggrk/lPDzQCzxcdWIY
bbEyz2lTmA7aG7NIUpvwpAXTG50Y1qKrO0af49mNI+IqSTjdy70mxyYk9penlxpYckFOkUdY8UcP
aD+o9TVSrw0Ab25QxunT+kxGErgPeV7+kBu5+rRsySOM6t5piwvQAIwkSqRyYLpYrV3Ya4qX7iYr
LCZhjDyzAPhniz5bNQXgMcZ+XBb7Slf0txjrZec82MBoyIURwLrYEXBd1UxdgApH8nQooIeME8C4
KHtJMp75HgLBaMHhC5TyqQjg7mEnXOLYeziTepC5+W1DfYqK4BzzGMZiwqQ22yLAVnOh3bsoocNg
HWyw+oKJHSO+XbIL2Kxi1QSkYLKX1PVxDr/ENgYQ2xjkn+hU0EAFqtJ6jriv63GS4si61XhR6DS9
szN+n5jg7sW//KBPwic+xujPChIqixQZ/qGCdXQDo/br2Dgea2bz8nZ3JQ0hcqds8iFjt2zoRFmN
fd9E3esEMOGwxJ+r/aX43rb1vmyfotc9pZ5vCytctRYm5REshDDBmlRC+66a0o5uGsZR471V7CXn
Ht0Atw0EQ0HELxiB8s9yGyIr1ZJARTLkaa+fe23BHp/MMOxiC75nZzwjy8+PiDjQxZlNacukP3fG
YLgGvwUGVDzzbvC8wytordzDbzmgq1dfemAUYZANKQsnpBJaTn3jkEzlE55CXXYjEXiW8SPiX2aE
ur/Oe+XU9z4J1UzbCS99pQ6tugtYnJNZHV2PA/pSD2cFtO/4TGYaF5oKx1kgmvCf7YHXaCWe71pe
EjPE8XFXNmuM5wKK8Xok277GRF2fpUdvVYlYRPOW9Kfigf5301jDvDjm2vmcsVxzi0fbNuZFHMOl
+h8YrXVDrV44TTKE5KM7wqd/ZSSH9OYjVdTeL1AdS36UUlxjZUg56FGU4H91e/t2TmACGr8uHAlI
osixFp1SV0zyVfZfTKsI/0So+1fWWrnjGVdttvi7kuw7lPV1JA9CeUPPIAGFotqshU61zpwWcZA1
k+PEfo+6qpCad9hVwGqE7k5LUZRgOBFm3X7S+tAgqxWh0197CC8fN0pFmWnLy4mHk4Fee+x/dp32
W6rLwRIYLjnfuOOpCCFZY0CEvf/nrsn8sdRR1O70eLPlrldO4J+f3Qg8RKPYSEArKpinzm5HWO5+
/uEQhlq2BXR2fnMdlR9c1jgyi+B/U5zdtoH24FYS/4ePQjKFf4aldr/gulwfWVn1y9gCeQFkbV5J
zXdP1p4edcQalLpCQm8vdR9OX5d/ZK4P45L4qiorhyA4Azqc+jEdlQBi0Ag23IwLNNj5dFHEEeno
52F44IQ/djS04xvFX9Ba6VL5aVnijqQX2j3RpTPWYYISSRH06UuHGHfSUWiJKNbKct71zvHSWG4j
03qE+EOutXE0fFnF9Fe776mE0A7T1kdCRisx6OZMccYZVVNk3aobAGTNBO92Jfl0LEQuH7G7iCLW
ZHmbtLu0cjk4yL2G3Zxl5Ym4paD8ebaY16qUZInN9UeTQwCKTsa0Z/+OeisFUObE+trvRCZP8KzT
Kn3No74kZhHNVKTwzl1QC43u2OjYAxGX1HtnjITadiB08OXkR7ys4R1DVylmt7aNJmorvFELyB9y
8jSJ4LWGywY87YOM0+/1TOFpbxpsgr5QNBj23FlFCXIP58maOytgqo2e/mtuEuwiSBAk/AS4AyG3
+twWJwhS9b3ZWPiIDZ/ETWStQmttKXZQf7wIFpwhaeIw9JoG+Sebf1PYJL2Vks8Y/b5iVONzAyxI
HBHA37kBikJpgJG2Rz2wP9CbmAnizJQGCimPM1uDkpn65+cqTOAdzUf/q2WxHsb/PC0OtCVOI6rn
q53QGBvNYUgpyvhKVx6mvlGq2NWKFZBINW8iSH1tP81qOpzFr77eCLBW3IG4b/ylzVJujpq/pVeZ
CAuVaA8z1jiyJaSngTU00gLtjKE4/Ebbv3QM/UCXwPT0+Yo7HzSK+ZWd78VwljfnHcc11W6w2OFW
Wc0JdcE+OvZ5xbBsquCqKpLPlaQ+JWHO5fLI6eLMN7KzPKxKXwG3Iy0rqec0/1lgZrKly7moP7CH
GyI6Ydv33Ia4jw4RN6S7pyjEXELR+3j7tKZxpv4mOpFUCvjYVkhIT8vNAmg4fk4JBNVxD8Sxb29N
ZgFvTPXPYmj+OnmGTKdX1qgy+WuYcjXYp3BD+wC6XYI3LGrSe19447LYn/+gfIaKt/gvsqo1mccX
Gkl3yNOdToCdt+GaD2m75jQzyc4QuX3SgsG9Dpfk+gS4bma+kyk3xMB2oFZYGpFsNvdF37Bsi6EW
56JHg3DsDhZpNjFZxWpIXdGOhtJwXj5M5wxrZvJiWrtw1dOEhvzkVzH18Z4sVUrmEqbcnZ1ECYqr
A5U6CldlIG1MRt2golm++Grw08GG4SqFsSgt0hzpz1Jmm3i4Zv0XrXvmuTeDgHR1WfjBVCVtdm0O
XEaNni1wLlE0Ki4W5ACRjLcggzsUyeCvlexQydoKoFM1bo9hALD90TGsdfHbYVgpw0SzkJYc6cJy
g8RW+5gbUGh65jDiao/Jd6supLY9vN+SEXPSdZsQeAuDiuEXf3g5qxG9fixNTAqmmukwZ7Q3pgnS
wQJ5pRkhDOyP7VEdEfQWXbQNvs/NPquT033Ko/xV/saVnb8hABE0hyoyl8yi9sXhQI8pBza3RonB
lLXZxSgsC8gtcqb4EMyj+4gEgY/wzqirSktXoJDXfQjdEp2wUKEO5g9r78L2UN1MXeKZT+hTtCKf
pWOt/t5CNvH45KKn6V8HEODr3OdDBOB4bUvA+y1Rm7DuxbJNQ+qMishqbbB4Lx36+zeV2Of4oPH+
np63ePWt6yjC5Zb3ygQ2rzH7DyFZVh38xLlbYfbE12/w3r6Gw509KIJq6WW6VlOQAOSXj/U429WP
p3c2IBYgcIrfUkusUSbCbNCSaOvAKwOML1NXkafiUz2/V6d7V0njVFUQ6V9FoRAkpt4qugFxnnds
/N5KpF8HBgN80MO2kQOQ8n7QvdTTxdg7IbvjqQQ19aFlLb0RdFEtfvopcIYEkYIF+1pMi7sfLrgn
EO/j6XPzJLFbG9apzpb15sPcaHCNdxXrqWp6C9gvpqw8NlIoZH+7GZZ25t0NLDCsvmfR5IfajPkX
b5b2VPH6J9N4UF0cQZz5GAtjN7slDhu10wyOLj7K3rP32+ZsNPY4VFjKslRZhcyPrKLX8fLX5ifd
N+OkNhIYxX/hzLtqY9N8GxBVVrMWABNW0JsANc2jo3q2o05rJ6ZZNyl8L+2StCgAr5/gxn4+TGPO
2mvYXXSLLc31Rc8rldiYaeNXnx1WjbNxopi/v9ZxLEdK1X4JNDZJ8sv0XTr0XoIwHWM/zaJSuQPo
9UmHmXpkh/lw0xFhJZAtv3AyHLk32pj4JOdubRvukwN0VmzNqCJVWQhgziK9uet8yxCHLAeHmc6y
eNAeHXWvrrphiq/b3fGuiMcc1IDssanCdNJ8jYMN/tv2J9dKSrWGLB2pmaqn7KPOi24ZvPS8d/rX
Rh+tPSYQaIraf5oJYgTEw7E77bD9VCI4FwVYYu+3uUV30VlgFi5ihUQU7jJweQ7U6rJjeI+pGLmg
K1ChjsYIuXwXW7aFXJ++nVQDgSZZFiPZGELRfdnanXm4JDbps+E/Ilh93+kk7PyFkbcu3NwXiN/0
BMNJp9TMjfhJK12a79wXaBO2rNfmlHaKkQW9jwsi5CmlLxfFghokUCJVyR/QPPKPkl4bqVerapiF
llTo+sG1Lq/eT2HwHaBwitRXMkZ/HCpYiPsQm3L14vQOa2zXPae3mwsuLxfArByxc4QG3Z3wKtXu
aIxcme14yLzE6rWjmk5OmCPIc/HPTUnu1OnmOCVBtAY/zNVYmxzFSsDlRo83WrEoEWFvGJExUtD1
TTBwYlCxzTN3PTD0VS8L9+50LLLYG5EiydwAlh/AqFd2mSUKIGuxqJ+ILNu+RASH+XpLbzF3jtul
saSKiD0MxZ7sYO7LEGGdy8C4n4Yk7yy+1QLtZeLKWrhQILAFz1pSHxvtEQ9UPS2bAcZ4kaoy2V1N
OBP3q27LtjAbyKUF4Tx6/179FPzjJrgcZJlD419F4ziAGdV06qshoZRT7iWej2uMTrW5GaCrhPp2
dSJ+lqVYTj7PUb173RsaCDbD82sakBCvNT3fIuqfPnJ31lgRJzE9Bss8wSh1Ewe8xt7FbzLgAEkj
GnfCZZdTLiULtnbk+IYr1pNCnVhr79HUeqGQzVCA0uFjnMj6rao8stOhspa5DDlzf6sCeJMFoHGG
L2FXhLl7o053EyHrXhJYYl7yw8WAMvxuVfVECm1xDWRVNYsU02w5Lh6wjuk4ZtbjNIxQkX0Bj96E
+r2x/ih70Qn+J2foMgMmfH5yk9u0wGik42F4b9c6H1vmYPLhISaA/7cR5Hy0uRwUO1oZQUBSs5zL
cXwrIwkAXAaBUOaG2pWDqnIpaGF1H+8DPUGAYRPS0uezmHWkJgRp06bte+fKZesVT1HaGLxQEzw3
PLPvhcvx5GAayefVOXgTnRVE/l8P1Ud6lwrw9+Kjo/6i7yvADLIsdsCp2mz7uFfMwQL5pAvHev8s
OLMvXMqLv6JSyi1o85YnjajR2bco2Mo1SKlXzHpME2t+q/yioKybSE4EeCaHB8uwqZ2cl1nyCwct
dzJn9PcdJE68ISYRrloRz+XcF4T/6EHVBoh2OxEqUmLli3zqm6OgqXCVPFSHkJOiBQ9n7IzWyGDG
DQf/QlkJs3gR9516qtwQbJx6ITnR+INgBWzzS+bAKeN7pSYE6eF+olj1jmLkH0spH70FWeED5XFS
lNe5EDIxNozsuCEuJkJkGF49qkT66N+i+IgSK3NKnpLouRbJ5PkxhODdlQgHqysNwZ804jc+oWlc
Ob0ZwLJNjjbjOXREQL+ZmPTtJiPHFxMo+xLKbLMYVLF6xl/6R69HAOmwau18yYFiU7z8d/gxeFyQ
1cr8gwqwkDGhMh1Ew/fsUnUHsAlkokhrqY9gfBmElBAkRFp9sIg+SrT9brOi0Du6aHW2OH6hJRka
rsESkJ2uCTk8oZoD7CXE71fGeUfuFUUaBcKb+HD/HOYxT2N9thDolZHRXqA8bxnE/AbWNM+FTPVU
1jk+pVY70M3+jBCruP+rkihGOBnArm7PyhAwg6gr0j5r1CnqN49w2mLx/tw/b3SMlUFHKlhlPlZm
YjMV8mLRRqZklen3EiIKDpYRawli9CfNk/vQVTngmD0qnvALFqQWl8GM0sLMdLEOjEocDKPEGg3p
3Bkx7susGVyqJuFlsjn8Mrw9lskaqOLAOwEMZycOpvFqBnfoK+46yNpoRCWP3hlrnSUWogRyDLac
1iVkUR2FDGdU2xfGZRaUxnMTGVOOiwrvRLaYtx1dajeYEH8XP4DzRtq8/mr1NOA4+QOmYwKL94f7
YZX9UU1YbW5Z7xb1n9/HW/DDsvjdQekGz4lYtzMiVknZH2qy8jho4HbX3U/7dYS4fjdorSfnnvEP
rFvCXPW1dmWEn825nHOEGhb4SZc4krXauZOLdLjrKiA2Ew+WMEdelu/8iNCk7artYVgX84t0S0HZ
WqvYBJfFMcj2CqVxfbFz87pP/bpwL7qUNzQAROKhWXrY8plxW3lw6HBAZMmw5bBsaXXiCk03z0wS
cjzj5pwp0gJz9hiX66ZlRUBowBnFRZDx7ySxkrFI4bItQa5X72BcaYdmYnD7Nx7jxhWAXIPYsdII
4aL0ng/kP5JTgwDcjgCRUfhMSyheuPDmq8222Ezj9htG6Bj8BUgBBeh0BvqA1iZlx3n8fGcZYbrC
MsL2U+P4eKwqDSxXZBJI4xM2zIWN4Y7nmms25xJITx+WBJCwX0M1kiP3JeU5Zbaxm6wz3326+9R0
8Jjy9o28FVjn+8N8+9KsYSx1CFeRfB7GPmZQbNh5fN4jl8o2ex/EM8uzot7pBDo1ObJjfnKIyoXA
hC4+muxre0Yrnbe145AlBgduBjSNts2Sy+T2ZBsCa0EaNQCVrqwkMRzz3NPB+J+NIZX+8NZB0UDJ
pB4KKgUgLAvxTQo4xR8ppeKTa2La7qs13jhtqeP2Rul5VhYa5ZkM/qDTEOyAlIR2mGt3NcPNt79q
1Ao02w87Gh9S4b3KNDjsDI+aIRs5ybX9GIti6csH/UQFYfr2DqI9rNeB9eihqQ2TSvrh7Okg5kG9
+ctR/Ot0ZHuS0qy8lJcT315Of9yUP+PsnasEOP1Kjwj4Ic6X18D0mUrjkS+RTGuPo0Zt9Vp0A+jz
J6kTiULdhPWzBp1SXlue+S+Di1fPk+dR/Q/jC/z8B2cn+PFpmL2uQPqTt6PTultEleqskgArQJyR
BmcgEJMcF2QanY/6nOd6r5c7ae3Eda1FYgdZsrZ5yslFvb/gh7bI690bUd7L1kWRdxPAAODlwPuW
X5j8qqPKjXPYtxWF88ipCqU0d8POAbduX1WXljmJY+lXiT0F1zlIXp9pO+5t/HrlAb/BfxXpn4B/
We+/ZebkCpPwU47DadrLNPUhPi1Sp69SN8tWr1QcJz7TBbMjEQut8UQGjNTfZ24Q7JdEd0QM803g
Bf4SqgQlXFQAQTJ0mrxDmHtygFpidyQQeGA3Xq9qe1sr90Spp763xMLVu/ykNVWxmUp9s5xz1R+H
BtdkE3z1ldgNocWkm3PXq8lctAoljgYj7Hn83Ah7Dh4MhDQRohkc2YVwQOBa23rv8IvwupMuYRha
2qq30UbjbiTi2tpjvxpoUXC4ZK9GnoXs+1+GLQehGfZhxe2aLUiy0eMEvJH9JmEpnxeDBYf7r+Sv
4ey4XULI0BMkxsPbASUcEvL4rpJgWDM3IEmo4lu+bJlyEbeBYb4bFuvJWJHcYDUQ9Q5pSWAh35OL
nwX5AvFZblS6Vs9hb8CdTm2s0JFwdhOlMe+x5pjiQTlaeXJ+u/gEiFokAAycD91ZLHrJEglDAHNb
QYnOqz4DSBWDkdeJA0ccFelU7FUf39xzgybnvlAE8u0Sl+2qALgjRu4KAJXPtAHo9x7M1NMNi6yF
hrKU3HO0OtkQ++Z3/e/vLn8HzOOoREfvzJfNe/Tk39t72kE+0PjKk8lORA1Rq+BAuQDpwfIpl1p4
//qCzpTxiEjw6DnmsJnjyx6UO0XaO+lklIB8+HrbiKCdYS8dKgzRjx95EprHrjTm4CN1BLbAH134
uEVcpSmRYDDXYiSijIBZwD/NQfAIDsawqso8pS8Rby2ofbIiNM4zj8/qoOW2WhN3HOqCfVyZCdCt
LWrVwdY0az0W5V2hp9yy6XQrDc+cDgXEgp9ZrQTPs8vEZhYDOCKrscFHTYlKKro8RiK1thEP8GQA
QTXie2fYWikAGJyhhMHhGdLFvBnw1+SmUIfjaBBvxpgSGIgG0WbtAn6oLZ584V6zddTiW1l3oJRM
xVfjWCoqCsJO0WPqNCchZL1tMFalq9202J2iNffx64F1Jy2InTgxRyDgINHBf+9wnFEtTrDrWIw1
qEOFPuRojyZ0IT+N1GrY/xqHi6GEZpyTRTM71xfEztWxfDZQlecyr7z5tE+MWpIrhCBTHcNa3GWz
1Chp+1RH5oSiJ9BtrYpM0nT7ybGGt1e5WMHPbAKI3TFOBB4hOtufX4M1DSDf676UHmZ76TJVLPYB
tptdY4FnhItfPqeZ/bhYrwB6voV5u4p6TNpnb5vj3F9L/wyCP56HLMsCFSGrAlj7oPQ3WjOr6UIA
f4MP8c8G6qmRVBrZeztllXy/TERHxmC2jQ26E3jjxQMRz9EYTM5DKsMe0abSsAP4Re4fhy74o8AW
/zsd1QFiHLYT7QOBoBCw9We+YhJFq/2Ug5Hp4mlhQKpM8Qn6dUyK3JVXj0aFUzRsP8PxEBdqzjRJ
YMpIaulgTBq6SJPQ6+2rxp16xAQaKmOlWHDmr2U/3LWExxWo7eU+XzZIOeK10PCz1vpAUDTuvurO
A6CCS0wWbn7Cd09j9Cae0/Iy9LVILDyaGXq3IBs+/q1Js1T2duFqeA1UZ6Y9h/yQxcmqbV0A0Q7z
X4SIPKj5zhLcn8iEKXDooRKnOoZxrJ00abFiUikgab0reCLolf6HL/AY/bB32yTwj/cQ0NLE6Xs6
siYsA0xSaAPkY8WvDvESQTfL+b1cCWbeayma+JX2QMvhJpLi2nzt4S7kiJ9M1kngTfDo1gEGvY1i
RZ3VGrZ5vSaQsKq8NXnz2pl+xl0XLB0jUCcDBYpMNudmyKa7MIzC4sRQIrmvLVMmkUTdvPrfZplO
yXu0X7ZdUdHwD9lGqpT3hyJmWqLnfETYeHm3XdcIPhnenQbCWzjM6lM1F+TkhBB1tvxOWubH/veY
kS6o12eiC1I0iN2z+S5E9vdijhLz4I82EFuJt30kojmNeDiCjqbXlJ7Jfof+VR7Lwa39gWmcaFoX
QaiS3OPZu0YVKLYSwiOV54/KZCJgRWPNwPb6JPkCY951ChnvY7kVYfdkneP1UZ4EvPFZ027sHYLK
nDqQw3xFb+sWNADFKs2IPPR16KiTlVXW52ShKbKTeYLyL7YOoZimOrj5PSa/sb7+eoe8lzRecZ0s
8YI3mQv7xfb6B71sIuWBaHb2734kJ4cYWoo0OISSv/jXIMZUVhW/wZ9+4qM41fffmeL9M0DX9vn2
+KH3lrLfTFmXDWaf9ZYL2OjWY2cH10xjiQeQIgZdAzkYpEeSQ+Dbp/V1pGvWyByWPHRB4xdSzw0v
qMeUafZWgxYHLj8iiWcWIHWCBRfumRFiEdDE5skyK487RNRMHXKqTyAUWaS3oTMu7B66JKiRbYkv
G4LwckEB4mUCDdsvW/EYT0us2TVj11mvmQ1RqaF2qP1lHQKDwC+6tmORK4kNVvSApvUr91KMns6h
z2SsbnVh5h6j1RyvaqJ/y/zX+31RUMS4maqizkH9WWQ0aGnLZoEml+GXJCF0/k0supUVZ3jNf6Uy
CWJmoEquXiFRU/MQ309vXLgRbFkCzs46RugFIDRJQzA1w4uSg/HbHpUZKND7LZGotVE3WwTYIN2q
HN5EgNb+UIwup54L0JPkkNlgwcJRYpUGmYnT0uPn2k2tgjiu/Utg1/8BqBdANNY89B6JSkiY6OXp
vEqC1JE4lusvJl3ISbtg/SSsg6fricpQ2T/mgWorkd7wV7TeZTR0EDX4FNgzA17cKf9W83NZSSvf
On1R5ksH7UmC79qpUQGbq6HXU+2zjA3fW9hhiguH4BKq3rMr/zLHLMN98AStsndB3EwXZUXNbqOk
0jvC9KE0q3r96qI8uqI5zWnWbFLOOOmjTxqclGN/FwtnMYj29zs5JbqGZRHqiMvlSQrGU11IbH7M
/xwJHLD+yCWlBO4bfo6CYdozgsvqsuDzNPy+mQ81Tf5Q1w4DoLdWyFRJwvN5NpBeg9bU0tSB73QX
yZGhxTjIyQzvCNDuE+/Rm3ljlX11n++e3n/FM7K5OAPOfeiMHRBsLCU0ZODBHJhtMm5wgXPvZq/8
fvEWUpSjKJOaF5kodhHsrkc5lCOhPwbBPRVJCfldaC7MU25kHa8z7JxKrk5AaB6HWf1gOaLwCYQv
B/zPZoesuUQm4ONCgfqO2tN7jp+7BA6Hj6/S/JWmonOJJjvsMOBQnvcx3RobxaFCOQJmZHxcA3s+
YqugThANqhIhSx0GXOgZfeoX8fUHYl1Gq8ezp08mrIILkU0ULfCMkMb6x/TVS58Bt+CDGyH4De0p
AceqBjY2tSsR3L+j1ImrCu/XYnnJV6Da/ktJGnTo7Ydp/gVOL+1CRq88c/QPOacg5pXxvbiYHTbB
4PJe8QeWN0N1DyL54rzH6exKG0tTiCFCd/sQdL7ustEK3cilr+9wRP+NtyszKsEXianex2FTnUUA
CXDHQD9wz50gDI/FIoFQEGO2cyjZzYBeQSlthIdDQ21toLnVO793oFNOGmIIBfVx0jFfAU9Eocop
ndq7xLDL+C4qyJw1+47wGEuFlPdSWPEdPXadoX6lh5IYqY+Z3Im5Argfzcnkeo+uJdDiiOuexxa6
/PT0i/ztOjYhLDi2AOilFUNIeGpqJHY9G3vqJs143sdReVCASiB6Eq0lJDyaks37wNN2ZaRAkgwv
l9pdxMzb8wsffYsLB8bMK9oiOfSo2WbuAFWNbJbqNRVdg0lj6QQWxUwnlMduVjJZ0doek6HEsFSX
eAuy5J/v/KN7na9Rjv20ZnmIiHaaUC3HV/wvCNtU4q6a0xdhjUQm/jfEsDBpgpvtYYpTClkNRETa
cQQ0U8gVvlhJOmMA0Ap84HEzuMxs6pNJR5mDlQNwwWsuqvynIX3nrMCBRajW7F8zMQTcJ6BrI8lV
QU1dUDTC5tQkLIskU5zw6WmiEUNMrfWvG9PpHJxg1iUyVYoktrKQwt/a+BvSqHPTCCivpMFSEBfS
bWsSTaSBDMdNQA/YFG3DQsQk6x97cR+v/EUR6HCxFFVLx3nHhVJOnMBa0hJMWL8sGB1icto+yZge
AHJw5MHRksaQ8mVLy2rI0/jwp5T0KwciGcUzclF6BSx3IbewtBnp1Rg7+TCgN6sZMgZnAuJRKW63
klQR4UOWt4M9y9io4YTavNsXDTq0jT0S1FMha7QSxtk/YKZIaDs3+CJUROb7r2iMIXP92TcxgpKi
WqN4RoSO05YV3NZXj1sFkF0Kd4hSoihO3vYmp/FzTg8o9aYkcwgygy3c/rba+iOqTXteNK9zn75t
JNOUdIRAJ5N7prfQs/QVVgz6o+K5jRc26Ebtf0/0tBsOi+DIpg/2oEgCCyYNasYUAHxiKAHBZhBA
hmDPwJKUDuktLNF6TKPFVvBTcnjbnNHqv2fQi5L9iWCjTit9Ef0NqeuTtMK7M7YaKX3H+L3+bUvR
MRz68lXe8M7GxvKzey8Elevye74cZqkk48LYGL9jgWP2EKuq/T+SBlZ+JFOspgLQK8RV5XdJ1VSD
nHHXkTGjn/TuXuZesFYQDMp9lCVEhc8xl+U3mtI1ebzNOaN3uqmkddfv6Ubig/iSeCnxzmzm3vUf
VH4M2kOXVDLwNzXJjnzpUiW28WoQfrNMJGdyepcJ86QDx6mFnd9lYoL3hhLBcIM0vX13HqJXOyTl
0bLjib7seBwzZpybZtVFvgajF6IpPMgWHROh0RM/+WMbHNHZLhZwG9zGiYoPtdjieQCBN4w8WCzy
AvifytlzRAwdk1ligacFAlSCeIQsbUsbpU+Px51LNrnWS6kNEOU4hZfJnM7oMd7igZDJ/z1+BWQh
DTKBL99iZRV2iDiG+zs3SMQotMXzvEGwE5KdFb/IVuh1kreH/z1lHsNAu0PICoQN4+QbfV5kOI9m
3jpkSgmUoYQRhZ1Ivb//ujc3gv+gRMXDXy+waihR/5NLVikAlLuY+t/iUPJLCU9HHURn6bn9QQGj
dsID8jGdPl+PE/IybFeeHXwG86ythC4gDowQNHTrXP9rL5midLppBs5/cQTo06CtY4jC0lDrbdeP
j8V6LE2PVEiKLdr7jUFo8R4AgkGrMdF0me6tXFdbFKd10ycYeyd+0vt2kKwMcFTtwRZYJ+1Z9Of4
HIyrmjlYSeU2BiXOMUKfGqn0Wyfycljp4ft2vffr7ilIyAZcyXik+oQb3TmR1maUTggbC3GE77Mc
Va5OGu6hiHOUdMAxnzm7/K1ck+LGGQUWa0ouRY6nDZ1G8DyrOXg5YaOwPJT5nawjlNLP/mXjDHKG
mfkmES5Hik6vHB0T1wv7bGVx5XFMLh/+gI82toMbIX9mhdFFGmoC7Chm4z03PytBhU7/J1lskybo
wrnJqmvoLXt8/tWUQ4CXthT7clDsiEz9z0uy1PcfVNtXsPEm1ltlW9/ncF2FToYV8q2MQ1II/fD7
DnoWNLiTIAtn6It709VHolJRvtZp6iP++cHkuS29RjIuQo6QlGbnWSZcV2lbbVE5UAMcLZin9pGZ
lj9pA8nXeAEggsni1TOaUbDKe36NUTSxIs9UttnucVCEyBL5DvtIteQmPBwMd+xbwUwVatpTTOfV
aOPnJi7Nz4AiKwtfAwtxQ1yxbg+vsHzAMzRsCzEjcYXGYJw8QehlcdiEobczwegctROjO5ojgAzU
NEeRr6yGNgbbMNMWMSWVDrVwHtBQiqwSwoqachp8zCQ4PfA8Nu5Ku3r1pH2JX6olIQ8pCHYURQar
77fNKHk+ABA154Zbc36hAWX4FZfi75kgkmqhw9uZ4AdxsWsBw/p9B0UyVascEP4RXuK5anLyrmtJ
yog4xUsAwcwsdHI8I9FCCNPKt1i0IZV7YiV0f/Gw/HKeTsnJ7oyJNvMfqTIccPAcd/7HA2hsc3CJ
Wob6iYEJ5LAHiEAWdOixC4xFVKq8RXAMgbeiq1XQEYF6DGYuAdTOhlpa9sIAFi29y2hz5OghZHL4
kCgWoaqEJQsDAqRXcXNzYvMzlZj77UYsUFDuVpGUnAnV+Sexm8yZquOPID9anxtXSwY0i36F/qK+
NIhmqY1w8MRioSsPijAcd52+ouomd/HVbxts5sqsgWwiCaFAcvjE5gnFRbr0sYHPnW6V7w49PhLm
y0qoirCA8oflPEIh7NQYYEmKWmS5iPW0sj+7WWpCqxdoD6x6K/Jb5nraygbehEPm/Wf/twSsW2Ey
qk1GvK9wFgjf/DV4ZvE9KkzywbZ94zUWZu3x/BNjM4Ib8bsPbhnywibL0IEEKRqWuWvfTD+Nq0uM
Yr7lJXRYCS4LinnwFr2/dl5BsyfSpEO8gvnHhx0Z8UmUkAO3P4vIumb3oEgUlEDajMRDv17V43qQ
Hclbnrh5pJma7vkZkv7082aecOlP3fAyQD00Xci3uPwP9fs47BlV6iaIZHVGZ+X+1TgcHQ9lV+DN
EM5VgP/fDXkBQSe9FHBWziXPBrAfuLoYEEWPUzxLj1OKMP301AFibN2R7fOAusxFcO+yA5LKute9
tIvJwyFEfUcwDea2Fm8CdNhBad1ESAyZ/9RTjnHJFyrySSJgBgYxcFzNpvqaV27K24A6sfydneDk
UzluYXVq9blrjnEMKwFk5undJd8nA3E7wcymrYl7YVz9s4BjHAxdrRcAwFrWd7VQlSVzbphXymWG
F6/ygVIDgIGRY3AqaZRKmuqRX6Zo0S7+7xX2R/oZno2R6h3IhUzMrjnYjVL/Tuy8A3FYeI5VG/Gu
p+/2LF7OCR2MD4Uz+dGTtmzzPvDpr3k4KeWHkEtPJSNQ34zOJXIHOxZT40t4545O6ro6lC+PSqh8
6dKSRjp6rUrY4yFQm9B20T7OaP7WJP2opJM+MQMpgQJ5qwQQaocHD+rwuQcauNJRvfgLDI/KjJEe
NJ+UaumpYnNRMuzAqw3DpZh/g35wH/J0fIOSI2lk/ByamEXykuy13Oyq5vMU9yEhvUTYEwjuZdoC
653Cafkdhsch7OIq9AixU8OAp83mgWMxdSh9ZYm+sumTKBh2OEHE+R8xr851tXhfT4B695Rz7863
1XYCu56fIssDlo4f+2hoUi1EydV4+Ze3rErwkJZ/wOF6R3pu8moTN4hm9/4CkprOSCT/JfX7cv4t
YIYj3+DmaxB/pq8uc+/ytyAMF85zjZqKBjuJO+pTzWc8207OZYh9AOcx6Hji7SHLGx6o6E9k2BKp
RWRR98Zb78Ne+Aj7ZHWbV9pyRbBTRpG3nNEVRa/whdIk1m0EGe4dwMPxYYX9c9dAuoppOSghVt9C
I7XWNojsaP4iU9GP6IyzqaYV3D0pZ3J41dQGCwhJihiWVh2LTTVLf7BSEbyN+c7bqtbUiu0hQI+8
/FJLf0IIC0jeFSvMKwMJPiY8uXF6zpKR9kJWbhmnPsJb9QwFBCxIjBclzfLoZb12UK/FNAV6QJYj
VyI/fARxSzicbywkkHlA8Ff7sL/eqlJ33O+hB/JpUUdsuKRnQbphD9twOzmz6ZTmHU2q6wZvJWYt
rtTKMau3kXq9lPijr85wUyEA0/mSWtN19LlX2+gZFKcUdxcPFry6YwmOaZLyaVboh/gzeoQS0eXW
npTVm8MkK1RmAgkseGoRz8jPF9lKeEMjtUqR85aH858CyV4cZ3QAlcwFrAHusFoNkiPbC15znQUZ
6rLH64Gl7aBVfRnktFWwbzdXgy0eM1AiLsJpx9Y2ggxRxpUF2BXMLO1L9u77ViuZU+crYoYAg6Dt
AclqoIsp/+LmU4X71UZLIxZPieYZW+EK6P9KeKoqqyZbKJVhWhH/W5b6yKxo/cXBCdmnFUD5w45a
SOmP9LFWn9BL61rsCD2PVxtoUR0jFbcm82EC8WbZBUZ18Qa2vL7YCKQsXKvVRp1hLyv64HoDydTz
/laqN5/Fq02YMFdL79Wl/SPGY5dX+j3Otd8sKEMbqhu6SvRBeMOm8E+iMZ1IDXR7caczJOUbEdTw
PIESqZYpEJm4tX+yEoC7aIp1DIRC54PtNk8QFIsqQZXTjrHiiGk3+m1+w8UXGG+jFhjsNeiC0vGO
4cgC/RAcwPGAMfED1NznmoFZ2wzKf7TjBdrSXtGj88nwvwG/9WW5N9ZOk+5lMNzUfdrKoCT6lDZo
dmD+DK47jpf5+ZZWieRQNr4uCwPj0X+Erjmq4wYdxZZtnTDmly9E19FNlroj69+kzpRMajO6WEHC
J6ZetnmGE5LoBMB2vWf40r0xaxvSIRjVMaG8rsBI9k1K72kLXfd2nD6KE4iJVyQR5Pjn5qrzH87o
ThgmAsdTXrjv3puOfFa/Ees4Y7mB2wGfaR/5jL7je55SE/lRE9LAh95Tq0pDif/ajGSMB64TLO/c
seqesQytIJjNvYTJS2gsUD81H1WzaXOzT1yAEjLG0BCLg800fmm/VR0HMyx7o94904SISpGgImTQ
QGQdjOQ5eRfowFkyc3KDxDtP6hNNcU+vt/3utTGoZ1XxTfXgfz4Z5BvjXQGlWe7BmoTdaQL0ydgu
CHCJt3JQrMKo8bETlv0NiOslOuEQv1/j0EUnEa6dmDuNcFzvvVmm/rCm3ihi/VqF0NYEIhm6Iyo+
zm+QAEP4zUaILHOxOVsU5re0bWmapMLtyi5sj+K0QBoNO1rYtp38cPNEkg5xPo1tqTCn/dzscDaH
KvQBRLv+hmh6blEM6MQ7fsQRSfSoZ6bHWtbqTWU9cI0a/Nm3IP97vVjxH09I2fxXTI8cmclUUc7f
k/t8bZRobJL/RFxg4swU4yxADNSPmFyn9yfNMWJhCEQrjXNYZ2XZuusmp8Kex4v83dvZmA0jGjpA
d5c+yK5Vw8w34uneRZIAAkmEANa8HWQLsbEcX7FosGz5yPxyUiDpxobK74frUJ7G0W7m//K1agqh
LTAkyyaHkemL2qL+6OF4n1Nv+pB/lpj7a0uccVVIkFfwh3usyeUfKU2ilu25FacVK+hDsKuhpWnD
srnakPdsRNcF1nJHRsgfb0EfIC5Mxp+036hUWDLd/GoEzSkOvhZ/CeqJW3v76+TAwm8rN4pFPHH+
4j2wIBXfKsUYab43WrvPqSNCUhX/U7SmtdJdG42BzCWgLaz6DQ1I15cmkk3LxqTBK0lKwrhYVUtq
NaNFe7wYDb8mnAuEzswpem9zS/nbdRktNQQ6uhcuIJImU5IhTYG0Hn/n9745w+3dylAGz6mbL06n
IEH4c+Cwz5MEjA0+vExyC28BfPOKLZSQXU/iIJ2O9jNzyJYVebA/LIadESdLEyayH1k0pKGD4ODx
f4zIVkvqPk8THSrBIKk+0DssB4wyte2RhzxreAaZDEDGF7i5us+09c0N0ZDI1JP0zrb8L5shIelb
aW7uMgdsV97NxurwR9Gh4iCZ2AIUE87BykvOHl4+vOZSoxD68ZnffjXmk0HEdkC1fKdO83HclfQZ
DkHI4XPky8vKWWG3o3W3X7q2+ADliO+Ywl0K5zQzUjQnPM3GrD6SZK+UXZQ88iopHtODzch8HR+W
GJ9XRwsI01D/gKGsPkoWR+2hTT0g+LGhwR550r18PrOjFppb5GKnci8sze3czauO4llvaGsTgwbB
o4BIMdSoTaWU55+y8jU38LTdYo35k9raLlfVl1bfj0/vQAiCkoJR21zBhpwFQvX9K89gs9ShTt7W
3OhIYRto3yugc9d7K6oNqwunYfW8dAJWND4tmYFmC5lxpcvox1Hkk0Kox8+vKsTqgic2sgAwX2vG
uIJL20Omm+t0/zNWXdwQzTbIfp7AcJTKjo1+ZcTMSUfeLwa+LQqm3P/Pu4CUORiPcYH/Xyo22l4m
1QvuBO4NlZ9EtLeGc6V5tMSey3BqEO8pJ0kimtUicdj06IoY4FSVfReqnL46I2C3g8HYX71O65FS
mxob6Uo/2w1hRaox+vPvUgq3KlXMubkpv6J5vvzxnGmPTmp9VeA6/gCQTQKb4nL6II+Q9cIkpbs3
5pqYTCKy3MRmuwFRg4fencHLv3ZEVEE4HFFVZkOnl91RFpUIBpSxbFgPUMNlLCR08o8fN3lmVmjm
9aIQq0M+B1LzMuIISTm5IUJL3Hxggmh7xcGCH5lGQlt85aINLQynad3iR8JFjlcyRfoqZ/1ENzpc
cMyhxgficDE7wanN3yUZTh/bxaoZmUe9aI8tqwaJ0zETlPo39AwNZmunWG1fLzPhHah3//h5KCe6
kD74b1pJnDJzrXJI4yUolsRJ7XIzIQKrCZT89GmbZD8xjjvdvUTFRH/XywIjXyrfufizVj+58vvj
2AleMJfIIwxIxR4q8D9x8l4AktT9ygInzagwr+Kj9KjpqQRXOviAVPXekDFEP/rpuITtCCn49+SL
NoAOC8r3pZM39vfpxtyhnMeqDoaLSR1RnxQanmo/PAyCKuyYsVMcVE3LEGStA78qv6ygI2CVRg6S
ao/USOgNLA7eYwRm3Le1gxtwBKSOIu4wGtvW+fp7AmI1IA8kIH18/EcjlxPNqD8i8DftStZPCxJW
rLMmjTWw6X3Qw3HaKTRhWSZw01eSlYPY4ouFrDOfQrWpNVQCpf94Txz+991UIEywlmteCHakuLF7
W+rbcaUEQbE+04PCGg5nw4zN3+GnYWxiO3KRvcd1dUb5STIy6vHBDmmpabaYWghzCVlum9XWMgEq
9N3X8/TMRYS6JYarda+gWaU8id17dtQe7t/rJOFqgHlgumG2ryEK5yZn7P3pu8OP3XtXFf2cSzJ/
6Uo6mNL1KNNXR055JNtjBW4PasEdtw8E1E2Kh543vdMkAGe/pNyIVtdZFsk1WRgWbxafkWaFBx4/
RSweSiSfA6jEYabsl5nvSEzJOxZNIQZk2cwQnlaIjx6FJ5GOGDEJL4Xu3HnxtbVk8ZGUy2g8rk46
et8oT5ljFwaR/B2QffXCH3JnKkYl8/9oHoyCw1h7V0avw2rbFAso86AWZLXPpne6vaimeBIpVCkI
+fr6p+xWg748eTnFXncqoD8kN9zUXkox2NoTr/RlS/STrdJMQZbKWC0OS65Uou7aBkfgwKYR+O0J
kovbjEQJBPi5GNUV9YiXseBbv4fUO18e9/yRWcMDDGUHdwe/gPhpoI9/0gFh3EnJ57Y5rtl+aC8N
hatCIWlehgSHee6zgIVMB0hryq43s6XG+3yLkCjpn7s6IiVVpYFBOslvkH9SiwS6TuYt5ko3vG+T
mZwWxiesL+Q2lMhTycMGVAHiJmD8bo6NoaFT/L3HOdkZIiF6gescCp2pWJpMxfSKoM1aWYIXQzs1
zLe/Zv+ggSI9+p5jfeH6wjWvLY9gmjKWTqSWHFv3c7axGVbVOJKR+FWbC3Gr9S7me978BU4XMiCa
1RJf+AoWgPENIcHDHLhOWBYaLguiOMB61COMxGz/bRUOUyNnW9NrSyuygE4odY4UAqxSrmo/YFr/
kGsEYMX8Ugy2NrMAnXTaXj/W3QzKuifjEQ3Bch8bvPdbn+vzQs524Ijigw2aeO2r658a03FTgGjf
n4N3LRegXn/LK6S0YBNVvsCdfsym7YoWmiFbT29fIgTG5a7ONXV1TrTZQZdn6ByDLhPaqPDTEiqA
xNn5cIHL+zYc3MnV1HhFzauOAeTZFlCMK9b081AzTS0KQ/h+uymc1QqmNPoCBr4YRWPTGsSliHmH
zTwwv1fTmAn1YhLYp7Dr6SOxjJde+4WZCJF71boUz0TPYbOTY7qt9dKodX3UY9XbRGQh6f/N/Umh
kZaSWNWfK4NbWkBsr4gk1jrA61oSeq0Ml4Ye58tOEI+gNEwVD1XNHBvI6s12zObDWEgiz3p+Wa4R
1Tu78U2YE27J3hsfvWKSKHOhQNFslNXI/dfTnIX5Nao8H9aISt0MAt24IOz1Kx6GWJrCAq72wDoy
XUIqkwZKnbpN+KU1/2Qu6X3QsR3Foj1qqmG7mQPPv2KZhI4ditFTd9S0p1eVbo33rleWNdPzPwlZ
EmY2F8I1wlZS6Sqh//fD5HXvSoyGEhIKidZeLALX+Aci1OPTIu/vhRX/LVhkMS0KZ5F7mf8jfdRA
BmrmNhjrWaU2rRsIG/jKn1xVZe6+CXBZ6v0hsi6WYku2/HbrzttVfFzK7ef1eyJqPu37iFmrwSBt
CHV0T03nWbAxbouLSQo7Knt3tjeCccgs3LunnZtW9TV6JOnTjTl3D6qMg9rgUr/VqNx52XnX+kdC
KtXiW9Qfexv6r/hy2fBXD/eHwjN9slHQbpTCHG48v//mJDA7/GpEwHyBMH27w4kg5gtED+alhjWV
aSU16Ud3eTpZMSZ+5pVBQ6QMIFZr/U9BQGmrwunce/lMmVHNuUk/dERzgmPlEHLjYXiC1ltHceUy
2ToFwF3P68Ev2EF1VdZvFViJEpr7cQgHVgLP0Uw2dRT4ax/fSNp2kBUE8BiIyguzAFHP23MQwESz
fX82KouuXJwSF6xWxFHn+oHaiSsAlS+H7E14p5CwZGDyBLLJI/MZQA824AHAb9x8PTQkc9frFSlr
AeCF3orh2yh9i7enlg6FC2cSTTSNE+hP4xHCWZeHucuDhlsTAf8jdt6WWeJqPK6lMCvfVvUzgYVg
CHPLCM3rdLgiWd8kbCf+aRXZD83/IgF+q9QFPQwwHbcqFn6VOoBG3+7Q99+sKQw4Iz8xnYoz2EXq
bUlLMeZ3XpA99sQwN+TADhnHXxq+Jp5ICYLKiO8osiO2ZLea3tFHk6v7yUS1y5PMAcvjNG6l7OGR
BUQPhLFc09yJJ3NOvL9Rzzo1/ID2PwmQ/Qw0dexr1ayGdINJn9cHe1WxjYkYzAUPWasbtqiIkcdO
cQDbzBUsxKdwSyExWL8NGoCwOIlNyGORZ/4uiBxjoG4uJLP4J9H/lW2cwwM1Am2JR0PGbeBbSccF
FAL1zCacxFH16o2Wv7e+AXW3eLVkV1poBrv6z32I9aU00dzOlyXFQrMlcE52Ih1F50G0Fi/WSKuL
UwAkWFM+aGlXDsTvBZiTTA8HA9NOlqkkSR8+vyjQxmE+qAklruaw3MoAP/1Xjo9lm+UzSPlaWYGK
ahSlQt50Gk4eZ6gsa2J9Ewca3/tITH4sID/4y58zZQTMlSut57423JhR0pJ5R2rEk3x0cwgnWWWK
+cMFiIEhlQ0rymQQ13oxOdtwxDt/iYqfWyISNhvU4u4f5zB2w6STRc0dus0gnaDWGf1yp3J5nZ75
DvWPtyl5gx1xQOgPvyEAEvSuodcIFtH09UsZI0ONejLZ/8jPypzsfiQ8GKOYM23az9lJjxCw6q6s
7JsSiwH+SQTyQnOvIAVqibi5HEUDzkyw2q9cmhpb7zrnFqmRfiGIPgWbqfdCoLN5NXj9spohlA8G
U11+5NwwduGMyhxcDBRru2wFQMURz2bZjsMxCq73NP/lFrSvTYDD6LnfiwnHEA3ZGASG5rK2Vvwt
NOW8RlaejP1aDusSTZcvyjKlohx8DvUpO73If5QUdZ2pskpGyjBP1bAIvPONd553KHd6EHCop9b2
dG8AOTF0ltIbAdWG5t6VxyhYCDsqYPOYJ5l3vG1M+og1jlmo1oN713Qh8to/Fb4gtv8hPd8v8Ssu
3ksh3CbINOoBf44Fu7LWrCPI008uCejNxGerCmgfJhGguGMhPG13M8xrwohD0vGKbJfKieROEQ8u
tQmGyptrHq0kG/7HdyBF8JQt1e1VSCp3V1YgWs9OlQYVWovuh8u9VQRYB8kTKNx7KtlPFw8U4vBV
gUD1s5yxa9AxRHgQ2xF6CPRPwY39FQQNe/nv9RdLb+1wgH/pRv6ThGa3os9G997MUBJ0sHb52q9W
dYA//CY98LTyykMsmHaIiDmB6BZHcU0jilb0JuR8v2pqSinl1RDFkozCdbZg+OEbY7Nb3lNXEuBM
zyPzXyaGJx01Iqn/XgVcl+9SQaSYvD++AoRrMKsT325u9mR2haOuOR9xET4aaLKaulp+Qh61z9cx
gbdVytDs0zvKm2PVAnN70C1Nl/23zs+3T5RsOG3HPKS33K8Y0nRsJhcoRyeh/hHYUtA12olIhhm1
catmHWpuCrnYddqaQI7n1YKk03QHVqDYa/gUiWZcvQxL8gWz/u3eEEv5NFC5UNxHbwC1SYejozWn
58IbRRIiqTfQbao8n3bruQvM72So7oj9YL6uqDRk3se4gPCzyUl/z/fqYSsihRyYh171UWOfzFjU
XNiuhJ5m3onbF9D3lqgXzHu6em4vhu3Bly1XE8SMJ8b5/AOBCojell079Z+7WONWe5D7cSftWFAa
Zae180nf8dJVDsdFUufxs4AiZCjxf3RG5hjuTodHK3uaKokH/SkySSjAeRuwHV8+JQ+KbFnAYKWj
aqSgrT5zAwjbbzfGAyR1PRlqZrc+jpcjKKduj0JMZpqVXYXHV9AmR2LtO2mdSDRomFlYCHyd2hed
Mx51bhSn2B3wxzuhBJ8WLfy5+xHLFqO1shDNXCOBIdBLC7zAo1CgYQTZEXZr1fXGGXsXCbvbjGpm
NuWzhg9YC7G+WIwiTcl1v1prtWX7wSqSKoRTBnJtpz47G2t2GXJ+r+9Q99ektNuV+QprkoxaFQHL
ELWm3ySi5GO1fBcmBQ+fRjRW7jpSzD7m7y95vcPOUqmBPoZ9zSd2dHocf7CcffqDdx38es71RZlQ
jD2JrTdCED4y512BSmjIkikqG/5M05ptpshqmqa0xWtTZKwXkEP3syM0qGipKWcdLmb8kNZ/t+ym
AL0TfsWLnzLQii2cwA7wWX/STr2nOL6hKVUe+rKtiYlJYe4qBJGgCxIfGvrRbbap6+GK/B52DOqy
jjcfKhvms/veKFoNnflQg0hgTWbMqjyCXLR3BQjBHyT9VZQX2saO2uiN7drm7lT6606zTKFwBA0G
6mlXYL83C5Su7YXHpGiQq+ZM9UE3JmD0lPOIwblxB5mS/q3wm5d2Ec1FdPKtrFqZWzRTsKIGqaUO
qYJ9HkTD9MXjpMJ/NLniu2s0WaXhF2oA5nZTnPA59Aa/ZshfH13uvJD1mETlM0tjt4WiPtOBERE9
hTWhjiqz4ISwRYk/278rOOT99mfI1n3KiA5idnZNHHTDGu85YlP11SS2+DSL5qN9aFSk7EqImnQt
acgDtwu2u2w74mNwuD0nLQzdhe1bWP5wPw5ZjwWi6hXtDUhe2Xey9rsnFJEays4xqR9DPk2HsAZv
wjx2LsoRc/9b52SHcfyjZZ5DlodnxreSbH6SkHgen7+alceI3bQb8maAiffwTbTinCtNYX1kf3T0
JbjJwBEYnh3cwXaFgi8bPlgHwlz8lVDu9qRbY/MVNBQO1D4lMqk42FwFY42GK6PoVLRaRkez7+zV
o7EzwL4Pmg2Cm0olKoplxuoANJtpm/n4LB5mmddCi/1nsSENxi1PYWM5Uz5B5RBQtvDTDoo2OnMa
tTuR6SKHK3ximDawL7va0uzsuO/Al4QQUFhgX+DCgtZfA8sgWneJJDq5E9EWsDjuS3TpMkEu/p3v
h8tOUki+huh/DBSF90Co/lI/Kro+3uviHu9rcj/T/cMQ4s7razHdyZ0pzTLBv5E/JWXMWqECgAaE
koDTZXjArE8wK/TCXdg/l97gJegrC3F0DEmLon9rR0lfnqfCJzezCkEYbU9AZztnRtzzIIfJSSqD
2OoVWLwgRi0AFd76ydCZrvnCIID9gbKGdazkArYHcDEuYYv3owi4ZoeR7vAIF/iVCGixDPPfiBTI
yp6H1cKJkeOSrHxjx30JCsUh51qqne/Ok+qcAGvDRQqlzKCxYZ5zpgrT9tLRrSrdnrDf1cCXwgPy
yPVAoDChaQbvixItCq6yQbYR2Nkq1Zvdbkwrgf1hW+bBg7oth+Ag1bHjLOK0E0tEWYHqA87MM43R
Gk94/UIkEE/oldWQaYfBs26wGwwDQh7fJEzDqC8AqJDXnFMUUYv463PfXD0ow/m9sCEzZKf+EoNg
RNRyZidortZxjMpvgvVVq5vIn6pD3QEevLOngMziHbXhKEOU7JdNlDVI8BNM0v7MBp8GKS/pb3QY
sjzbzhRegY8mAdKQ+CQPruqYeJ0uopKLhPa+GdD2vo9Vi8aV42HXnBoPT6AXOHCm+YGoJUJhzg7b
vIeMWX9oHE01dCtN02CRfNL69U8myJbVMs0T86BA0ADkSR/qrICjOGHoN5IHoml6Ix2H5D6FW4F9
7KkOFriP4A25J31iDzUEUIc34TITmdjpKNpgsm9iaXvIQooPoY2bjJ2bWKMcQpbQAegwgiUrLcUl
rPf737TejoyXMWD6hGnAt6LZe845uhONvnu2DNR9MD0mEoGoNw6vW0AhY+SFbkewrIV1Yg1moyM5
x3AuzqU1/wbP52AWZdLB1d1OjkZSxgPewF7cgLQXMu2I7icXXcnbq/s6fSJyIsi3FoMi/Q3R0MDL
AhBruVVO/0LsF2gk9YszAIVoc0Wb0EHyiaOqpPqpHMrNf4a6lB6R5GSgGZ/jZXoq/OcclOiGOKOe
73t4RT+VkVoTfHSDvOHv4xi75wxFsTRC3uFS1HdNQ3b0r6e4rbK9dcWjmdIy8EF3rWU1KP1363L0
CtZJxzs6iQyv0KsWbJRk0psnU/7fyqzmwSU0XvqpDO549Brhq9QiaymdnC72eyRnvW16UOmtydAk
vM90RZXb84KXFL3JVPur550TQqOiZUKWFnI0yzXWvy2QA7hK6CCyz4um+0e6FVjUFB5bOlUabUzT
IKDkb6UmvhbiJPBH/prGpPju7fRKdCTKGgE2D9y8yCNsS78X/gLYttx50iAvG8KNa2COdl7FS1Fv
/aggSQ4ARfpC6betiJxhn2sl+mH664lpm3cuLpKO+V6yV/Ol9PrP/7Uq18BWdVIhj4slLIPAWLjX
xM+yUv8eZyE+7ZO56Of6ZwTjym5aiNayEjPtk5PptekIzikiEFTwEWrdhSEHQUqwuwICwaiUljMl
xOxquG407UCUwnAhgsIizec0keuXj8Qb9hc7F4ZT6bFjBxQoe/l0lca2PSbzUkHyXRTRnMqCKFZy
ZPDs9EREnn+l6LgZLQ829Npk+lqPoLPh7fIACAYQureDurcJca1ax3AZEsyRLKRhaWtxLHYg82g2
k+sF8Y+gY+ckexvOqpdSrqI09goD3FQhmpiCJP/+EQfaNq3IAYPhcrUz+cUvoLeQ4bKccgHF/Tel
XZiRU0qY12Uj1dnLn5G5cyoQrZA8PZfmGoLLloEDEUx+vut5Ij3ywLOXzG96lX4UyzSSQdeXuR/E
fCPdklNkhiSjcPqbfH4BTB5+g57pSnJO/EDmBVRwjiNTOkOKSyxXhgF1nU3k5OoZhoq99Ofly17h
9JFgVqOufrLr92tGNaIHBnpBdd7p1MiCO9xFRgntAnR2UwhfKrrmBGvPv8SFkRXM9qHlqYjbHyRV
tvlj6ZWD5x1J9F+UDGAByZcd3Fq12/eNk07GeBbkmx6ggu/bkQncZjh8+NKRzEGW92V/FkOub+6c
lZgXL+ST2KvCwqig98Z3B2YvUoDBxv+wK7f/400HAhyfZZBDOl1g+SMa9vr3CZ8MX2r90rKiKVIP
6pOnqD/CO99Qw2uxJI+8WMlpveQKK6QDzCdH0xG1V79kvf+cEDSW2ThwPWcUtdtUbKoH7RGeb8SG
keDatMCLy8znlAsZuoojsOGqP3VZhdvWePoW3xaCVMtKK6fS+SSG/jai27Y5meeuhI5UMKG076ME
NLhg6tS+BzEmJAyDiQ6HmMYnkftCU0sex3zMWszaeR86P+swiH9/edD7KbAMvTyUzIm8o2xYSFun
piv3EIFHPUyZTgd6K0bSK3hw0Imb1kJykI6bSjxHZ0B3IDEX2AWcJpXCp0uuNOFlc3HqntnT4RSC
2f/adelsx9r40mDM25WyZZT9phF21cCTPpzzwY2xUBRi0pDwG0AgABQpuF6+qFE/DE/7j6+4mIPE
fXk/s3YroVuawc4XmxF8XjyA68m+zfMqtCRyPaBSeO02tGwXnfsqmuMyUw0NEVVZ0zIYqhiqPpzN
i9QAfDhnN0+n7/1IIDUs3lYjrSVdVQoi/PHaXS7KGWvAF6aB5DB1o8iXpGnZoVGCA8twuuu2K0Te
an7mqdNaWJsoN8BrQS3QSzB+y/onbAosBzEodrODkulxjBmyBEmcZlW4KmiRHAmR/UaRmwLlR9Iu
H05PaEq8ad1SBxRCYe458r/uT8x8G7eYbV/GiiBw6rvHxa5LT0w1GWztctJM5vZLdPx34DwKBxWz
lHsE0qM1sysQNMEESulC8JyuHAqRByAwsAyLuuXpQZ0VdeqndWgnETLtsO0ZOEXt/YsmgN4cxNZw
iui2SmJ4ug/k6diEtKMnAjFm9DT1OCVBuG6jl5BzUCJilMCHCiJCMFbBOgmqir+g/8p+mMMoH8B1
wKPxoj2RYz2sBzw0eAoYTnKOT5LSUtqAwgUrHwJEhn0UODCgDpV27v9AXLjpC+MF4EfSres1CVb4
CWiqYbeoE50JuIsWRYapjj6yFWFrJBrTYnzdmZaCQ1Z/2mej1f00Z0y0U08NzWDt43cqUY+O2wdI
verCHnK4vounogCEhvaWvStMrRAsHKN6W6D7nMFnsjOANydMTRuHCsiooJ2qXhoAXRHoqa8BtMg+
glVwbecMRBxUmjZ8rjHLeins77QlD2lNtxO1hzr3wEw0M8cRcm9czAFwid/J1btiFWn/Lm3+l6CD
cCRm0f4mv/B2i3bmHhOgCE0lyBu9UOSc2CN2sssrCv2eXUqOpX+eQQ06wfbpvRgRelUrroeM30m6
loj3j2kzQkcCpgiPyqYS6F+Jt6zABC23jfD1nWKLjWkn9e8BQZljEDjtXp9P8iJ/p/1eMinqiyUo
p27Pi5gxC/Gz8+EYu46DPRgBqC15EkDb/HC71kAIVkHH4EMtGOnjdlqCUxxNnp9vg19kNxxviPLR
vTVK5K+xN8B3K8vek1Xp4k/owV9aIAmps+ml1ucTIK3nlPFgETBO0btLBHvErd/Uyj7w45UpIOzb
G/rIHV0lpz7pvAZo/WxBIigcnhJw8NopjOT7fNt7onoagPuF5WpeKMzw9MvOwYGqVGmLPrLzavlY
v1XYh5hECYUSVYCyoIMZa96md0ODbWlXRUU98q4mMMiM8OkYB0jtwLxrhhbVXfwj52GlAsFT7g+6
X8XKBI1P8nOptKr5ORB25KtHiN6pIRKe6GZ6XkdfHSlKbqi0HoONuCPCFSj/lrlUVJqRb3cG3DPh
aBwq7ybbcQY8V6m6z84wCVCNopHlnGQXIxcmDdv7/XL+rP8ovU/ltdXwBdduIj13hxKcTgysBd0o
2SVx4Zk+7pPNxpb5ztAnsP39FZvhQHG+X6GVLjQmTx2bcCvKvdwhzOX2J2o9Jsw36Slgxjw92Lt9
Duw5XH11/jL6Iaxj+4nCjnu84xRf/VK/VPoHbz6viNCMn9fyKb3jCXe9GAKbP+nY7Zi12WAe+0Qd
VOQGb5YRdCVT1qK+SpDPFXcXt8hl0deX1+kQBcYCReN8bAH0/Zj7Jl6zFy2RMlnMi7Nj6jM9WFH/
AEM82uHIIf66owGvrGfjVQlK7/G90NcPbjZDw1JXF+8CX35gLN0w3uNUjgWsinPyqWizqudMvUzD
MllHpkF2/QceNF4Rk++CqSUuo/JwfZLSWL4KasUbjPKIq29J0f9DnudzkRnxiEw96IwIaKOnH/Qh
mwAxfwHe9fwgNw49PXSeeDbi1Rmwx3I6fCKqWfd2us9CE2vF+4WBxSljYSDGNYhgQ6ZnsFdkqCXE
ebiuG2uMOiIrip73UJvauubAZTJodSn/wEZsZgthrYC+7Z3thjNOFNENZveoryn3A8fVAJOXVJ1s
UJSWZl0nlGByAD/RsSq/SaDfLaCTereAeKuKZ6JYdH6fyNwkSgDbwnm/uj4P8hll8y672DtJH5di
YJmLk77CFMpbUkddfpKI5ivRLU6feZsuS3EHSeo1oXizWJHaNAiRJUno6PKLcexzJWay2invfTb4
3ABfddfWu5lalUQg7KAsxgabNaic8pCWVnnI4ZvnzzZ894K6BP/ROYbRqmtQYGMeMs4EdUytXK/f
aLhhP/ehJwtwWeBpOCmOuGm4B5POCEKYDp8cJ2qQgERupEmIccta3l1ExRomT+8As/gq5KrEPO+U
KIaeGaioMO8Hfl9wNQGyNw6u+ZZyYWFL2CfDoJ+7eNm3TCuw9uP6xBSOHyqvmNNNKxUa7NWRJZI7
c37cfM8iBOIjA7hPHze72oQ9zGzATynfPdpo3RuYTOBhzVnvQSNVZLiOrIahoHu64c0HYBDnpYvG
25PADA1sv3lRx+EPSgbqOVn7pS5/4e9xtUaWcnN75dq1wDAq+peB9xmS4yS3EJIJ/fYoE8VH1CGM
KFTQo3z6vTjFkxZx/o3vLs3KYRHR5Sohao87T0Ri2fw2yOpv23rsoBAOjbCuD1lSSpvM6TJ2aFzX
C17mYgm25y/UHF3rvNrf9PMN5qy4FXOyBMR/UQCiS+VCieLxvj6ekv/UuCNdvP6pbHGWsilfxlB7
dBALTlT6r0y/s4+nHZlt382UBGVBoh2ttkfv6YGOGtOqo7s6l41PRDPb5jc5ubVxlOOZ7iGb8RGm
jwhZdUwz/u/ohp9I2oBFRH2dTePJBpMFqH+wEm9+xI20Nc3a2/eMtXAkCLpV9e1w++xTdURaziMZ
PVdRPf8oeIwXCs22SJ8gc//N3Lu7R3UHzU/5QJ3pH3XgFltMOC9jJj8cxI2ju5y1OYP4fnbxdd2p
GgwFmtvj4nqdw8mrtSSexkLWsjI/J3FuK4new83Cdmz3JqGtFJkEmYPBfXFBSZ3TEik+ydexSK0O
aCCQq7Mi6jVdOapZaej6vJxH8xVSe9BVMONPP/2ZpSK52QjGQcthkEPV+Cnl4Lc6cyyDe9kVBJl7
Zg7N9LUDZ6uurhbdCDp9BAd9cGsoZ/WiYAmncF2xSbPsUKTGmpJ5/eDut+5ezJrEnOyJsV8kYQTc
SJRPJLdHfI0c0EJy4+80XZNwRk5o0e3cTqyMvAb2z4f65WjVPjIonA4tneUpHK04UVXZFP6SpliO
pK/X6E+QxQz+Ses5Nig5cbd1q5Ij0/fjMsEk9v5qfACkGMDEYydU11S1kBzrNJs2E02f0sSajRzx
TRJBn5Xg9qlFi11+sXB7PfDvw2asPJq0mL/EHc5nbdhybgdtZIALcra/d0HDoCdNDBFVKj8Taxzy
Z29mWvsa0oeiG8eJPZf6fa5ho9u0YCsmIa3BSRzw2NcoVD6nLsd19/2jendYXDZVNc/LxeEpp6Mt
CxtMNFNEq+xRkdq1Uhasrigqae2VLyiToUlR5VIKwSaWcsdXKK10MNc2SkAFuK8Sg3PV/94k8Hsi
cMO17ixQ+VsB+ZluJo2uaB6HfqnYqDeGmDtPPgnoC/gCfKYW59cAPfCO6M2CMPe53evifGtZCxUA
cjqpuPKSqj/45TAA27SONjqRVN3sH2SosHRtYNlcyiXC59zwc3DXaBP6m88rwQyd+JWs727lzm5r
oITGkY55sdaeELUyR3rTnttr/KsuJRm00iT2egktYpq/F16xoOpv+zFA5KzufG5FpEuLtUTEK2lv
at3sWxzf4omi1iSG5IUC6CoRMjIGw4P0OxEUwHxrSNjfNWq31uBF+bjQvbN0IZIqYr+lj9v90Rtw
J0s57VethKap7cQ7L/d2+30AQHagUTXnSKVVKOAbU+pTh+LxU9hQHSIjKvKLj997xSIO3zeFbtup
NA8ixvSMkGbUOyWqQJrTAB4ncLR9LoQutA7meFiSNGlLnsxzLt4JIG3FLdl9xEh68k+9ykMrRw0y
ytOJPWsqL3sZOLw6DCQgaFenlpYo6Bmxik28/Y/RHSKuaTl08IAILWr6ebT6AuCqqeOd/hbrPDpj
A61j3mXpDAH5DxnK6R5JgC7sUbV9BIc306lGE1TZ/M7rLXjWedJg+gALQdsagwKx5l67gKw6gvlw
05DvxP0ZQxtL4pzK3mRBz97kEfQH7l4hTBqCugqEtIiMJBScAPn7QaVTFj1ZT2h0oF5Mw3sMAys4
5FaWVAQBzdM4FwYxA+Uv3P9qcpj3KkoFu7PXHa6CrpNBv3w7IdOaXRsxcIChaONNlUHNkfEDNevo
oHFNIIsyn2NswvVwFI0BM1e+f5094bDs4xVx0GK3wmmv7eYTCaokUOJTqjCi0BL5X00U6KT66Fra
2I5EOi3WIdeHibmLDg1XB/He2u5lR6kXpLJZK1bMYK+Za+umuiNgNWqMozxYAEKx3JDfXWpDyfv9
CCUhjs2vGb0/avznEHzAKtoNY9PoYyVTy/4mRFaamds+T7v/vg+K34UPvnK+cJarRuA778VifLik
eWz8+asLK02Z/VGFqhKhyF9KyDCF5DF8/+YStRN90kU483jDrCglilHxqt2tHw162KJ/NK4MEguh
AjOU0JN4JRaunqF1TNEgHNBNF5p5yR3nEy3beCQUzI0o2WS0vPGhmr5YTU3jM/EK0Y9hMtt6c+9Q
HD2teWQJbv/hxEvcuv9bDdXQIyIQJyndjeg1bVpJQgtAbR5k6d2fQ6neTEp1z8th+7364cDfKati
YViJsTKZQs1YgG2js5eeCbPOWSAoMG6VeZzKxZUYj3P/xmk2WhUJxX4AJtLGSYdWQYQiCGRMx/jo
K8tnrhJ/1hpVoQpelI+4wbXJwFvgPJrA2TqGnsJbLNTrNa7MSKMIBsYSaAKRuKkdf6Ury8ASR9/U
NbPXg3ZZZd7GE+r+sGIYh93VBvthjOJCurv3t0NBNRDxnjfXaX6vJp5/jrmQa4xWtQhc8G2YJY8O
9Ib280HAD7JewLi6oGGcWGpdl9KYQswjFlWpP+Ps7E4ZwKO8ypmZ64qn5Fn+RRcg2iZt88jzkbuG
iAieN0lo3YL1xa42jxRd87EqseH5fc0W3dZMwkGSZZAHm81iCbn7DRgeb2VnJ6Rm6rQsGrE4DBXT
EYS855rpVsHaVqpTuEcwZJ8CwRQcAwM1R6keEuhmVxl7fy4/KXEZEGhOrninElHS1NGwJfaGAF4m
nVkuiqoAzBFuL2JvveFD5XLHxGqmiem+7/t77ySDQWpIYT3LloEf6YCXhbe7dzLl1lDCjiDMb+rs
OLCDbh/ntfJjqXS/6UWQpYuQgf4QJ0zxFWSWsUXsJHWFv4CkBt3bxQyyKZZt7ypb1AMyzT+xFWvD
oYj6TCsxDP+dBK7+epOprQbVLzav+B8lvJR9wCmAD0IhuyE9NXKjWflHl++cOoPILCtD+hozIUeg
VfdlLaCp3GYWmvwkxlhZCN5862dX/YkXwFjPkBRO1adMAIrD1QfmaX36JUmSssO8E0I0l1WFFAMH
yxXzQ/IKqZH9RdjzXXqb0aLBSpfzdz2au+guRhQ7nICDAMTUvlYvx3eo98sVc5uh1faM6Lfnfs76
TbkwKjJ2snDvzsyUJ++Uowrv6XVVfn26YpYemDNkpt8eh78d86h8IECtqPDQVDL3LsLSHCOMPS2h
TH4Ifre3y4/0f4zgBKuU6GzXj/fgqMcxFQlj5GVObwvPCk3RdVHvJlrLn9LU8uXM8janhUN4DZ8b
Xxv7Z1Q4ZX56WbAZGDacOD8YufoNlixEnmLHa+9kYS3L1coYI02NR5Z7lJEhbhL1KW8fswxpIDg4
DgMm4MGYGEtPaC23+rGMJnNc/eWv07rIuBccDOYHeogEZgG9t74fUGLl+4FM765zxvGJi9WKZ2jw
9rK+FN6/E8w5+2ioL2ieg0XhdNavj8Vwj4Zd8THRluvItkHZbg7sfLe5Z6Xt6ad+9bkZxIBRTZgz
Sc0b8QJ++n6xUkFeSZG4sG4Q6ne3174CDza3VOyyNOfffrwMkZ1TZxt3pv3g5hX9JN8KyTjHJt2M
WPfXyTd1pWnBAg77Es8LItsSn+GhsGgDjfAJLYUH4S6JRlwpSFIyAcE6Uz9DCaAl0MPrgz0thCTB
J66zkf16VYFpTbY1L356LLhuDctZYCjKJw52Nx7Y6KUZIoYWT6MVhAYGg8T1icGOMm9Tpl5lxhL7
WpJ+DiruMLXbRCNf/v36pw84CLU3+vAI/kxEZaH1zZQA+bZBSqIRhlU/5t0GJyjzaS7dlaHQjJti
Qr1tRNlRKUZaMy8ERWK+9ZjDRjLN08sTVOG2TRsCc/a2fWX5X4f/MXxmtdTjUu+Xe2EBwqIf4oMN
5egittMrAvfRtveO7f+aZeXu4Tb8VGiaV7cDGKO+9j8OgCeaQrLMsu78jbCnSGHUEePIsmXquCg8
mSTC8Af+QBLR/cz/3woui2xthQYz29LSOMbSb41vsAeodF4aE16Y6vvcmy4aORbw2Uo4dhtnY390
Z4mo2+uzeVaOovuHPSbtWf/WsS4b5s5dpqRN7+b9dEvh3bYWjBKFGXNbhR/GzYIJqEkYURx/YPDi
87Hlx4Ii6Zru+D9Qbv+aOPw3BLCjM8GrP6JV19jTK4+3pPN+j0vvUsE/9IxietlpmSwmeb+NdWwe
Xka+QZt93Ba/11wkF+vxXD1uJSkiiNkkYpV26mUsJAAbd0foZVPDtzAAwDlZ7T2XUNnCB1qxUzZc
W8WYce0njWHYZezNZ5ft9WOawar+SB8/M2m2KsUmRyMwEVbEdE4ov/gJPzPaGuOLa5bUZdHc1mEQ
vrq6bW8vYS7uoJ/gDFBbgjVTXypb1Z50dyxrV6KcaT6FdA1hxVzMuCBgR0g/BA+pvDHNVoYt1KaS
EGrX/scYOWK2vDsCio8rLz7Bbsw8cHE4E3eJtWZbsfbsYrOqfR0dLOpMdqI1MeoZrA7mZZ8L/UiN
RYuYzRxpScKwWIbWQePtWUXRNJlVN+TgZUf0A9fshQISWZClMJNS8YAojHUTbeexIs1pAgNLOSzF
mr+1dJcHgSguFNNVXH3H5CbKZpC79WL1SOpxlUzKqmZ0m/kIsdL1sojcujm0pJWW7EJn3tVDs4wW
w+vGXPPABBDTnExm+hIN+4xz4ke2QEkS8g0eca1x6Z2rLTi8qhiGCbkyvSxs3C9HAbcU1djfVyoY
QtGNqyHxlA55L968L7q6pfupACyTHiY58sHvZKjLtW5692keumub0RL2ukbkhNqTCcIjo+8eWDzA
INUfuA6i5yhuq5hoXjqiWgK5IGCSXjbOpvkQzi96PI5UtksRrm2K01xMXwSj6VX1QrNzcN6zZFBp
J+g89tk0jpUVYauGrxyJOps9xyYTcscqPPVAAudRKTje0y8KW84H1kInUsOj5oxNE/XKCYYayeln
l9gIf6acVBTDLgM/AMrVk/x9tc/Ln9RO1rmiAvo4b52mOtHrjppAoIIcBzdW8hY0PwcJwpu7d/FT
AHeQZoa/+z7/EGokBr2WySfTMl7xYAo7sYpLLpR+jrcZZHkgYr7Aw5gyBZgzNQYSUSHfQqexMMF8
/owqx3pMiVZ+saOF7mcnwEyZ0Sx4OpPoA05nJ5j2Rh7/8cHr0C3OR2kZxqZgZlZ5XbFCKRLV8kpO
78u3ft/ub/V8b1VnAf2xXpoxPVxCiiy6GRRFTGV6roIXLTwO86IXXymZqJQCucto+HMwWSQi5GE5
HK1y7qcN4LtNoBIIGyYl0e4mNDHjh5D0u202NZh9pFmPwoSGo6DDa+eIcy0JORcv+/6bwqGRr0up
cwTQYqhviZA5wScxmTIR62j/hht6ws5kG8uG3buXN+3B1nNB4pkPB2JfXidAcy7t54mP+aASeOwy
JRj+UN9Pf3bKp0ZtsbvzGF/NZ+1UKkYbDu2f44JTpJTicaAcReIlYorxLgUH1zMcZodkuc1Zv9p3
bh2MwZIwSAS608GP0FSNGyjFsjRHukOBMF09qlLxsKd3o8S3IHCY4Up6RGQ7FwRlefYTYGqfL7xQ
crKs9j/ZeYgsMt1z378Hhn+MWkDL48sSr90crTNh7mAow5VlT8ggI7dJEIdfaUaMhFQE3jC+XtiY
fibxfAyvZLkO1umtH7BUm7ZlD/l145Z1yqPADZ1oMeoiTjnC4KsFU9x79VouLQAcjabdmdYzvJkR
3j18HruYVFJpxh/IZRH3RBXVoHjI4YAowRGq+TLwf+jAyqNUdEFgN9q+nNX6KnTUNf89zTfhB69J
2jG6Tt6sU1BmDpDsBVa9wVTXP8WIceyLcu2FI1Q4X8l3cw9mI1rv9H1Es5XnL8cAlGAlkzRFQjwV
zAT9KwOe/vjEHbOEGJiGZNmLgz1E6vSoWJ5o6eBURqiePrRU+AxeG+NJ7lj/oTV4Vw6SAIdYlRA8
zxSqfJg3+6vYQfei5xteR+/Ka+YtjGRwBUwGqiwkGTC6QbKil/IEguAFzNDLNxwVtogiByYhmk7f
Nx2bAL29m3AGTRNTsMknNv1e4I/FQNS2pI6PN00RoZuM/t8OO4ZL1QF+H2G/9x+FS59njCJ1lG+s
lpXjg4fQXWyLR6CxS2MyGp3sSDBz/bbvd9zgUpHE3zJ+4CZmOLF/7pAfj71197c7kTEpzv9O5J1R
jls3EYPSD2Me7iiNZQTs/PXQ8hfz8n8OJJ7aX/dDaHbcZtPiLoeAdpqG9IPMxdT7lgOSBpgSLK5B
Oe4A88rRNmu4oWO3fEQkHYwhjdxsiHyOaxzdm2sJEpQZx5rNYBVIE71xnTpIxD2Lo6eDev/vwwUk
U03GKxDFUUZmDxEp4AwvtQKu67ytI2Tm4MDe5YMUGNh6U1OuaqZUeN0QsGgWsStxRzxc3L7Abtga
WVDplbe22QKwsbTNRR9xCHS/UbIdanBBqbWxGi3NRMKTMe0pqN6rP2Pn1XBdY1RdJOfWb2ibjG0w
pAKWB2/9qdabCWO/2rkSyuocTpKxmweyoo3fpo4lkoaguSdSmafj0Rs3X2A9lJOK61KnEm3e/jCv
Cn2NrtzRkkJ/6imIQ1/6q+U0TSs4RvatV6/nVMa5oWMwreZOLUDAJZ33Fdaf9HqbWOoPX0WbuwXa
M8Y8UInZICQ7gNQa2kM1Ux4Bqnm1aKChSAjKnK/GM4blNCO6CT7ntbYY4emDmqZaAAugR7MO5uvH
XzDIT8SFchtp9JNQD8t6LIWPU9vS4/pWHeHCLq7VYjWIhX34Ri4rqtgl3aogOK/HDruly5Vumomh
H0FQ8Zt2aVMWNRUCcBMyx7GzSMDc7wnvccHwb3bg7pI4d2JP40+xn3n4MQQ/fqU+3P3fUucsurzP
8lsxzxUGdWn3Gc+tFQu99LjmaR8AzkBQkajc00dlqzK8lrPyhGYyQbvGZh3qFk11MWnIZub6RufP
U/QQMCVXWoNRnrQDulkCWqediOOM9IyJYPJ9/cLapmzryTSBgN1dLvqyq8H0e2p3aptsg/Yw7fte
xgvdaEV9qDRGMqYoQlcrB5fpCDp82z2ilhVtwQ64ZSRQi5PcEF9hlDsM1JOCrCtT3CwFboZX1EkD
ZNSuY+dNwXRpoCM+bbLFYXyCCOmVts7MDYn/luLoIRzqntZZRhwg3yOqXI409CVtbBdaqCV8jOwv
ss192t0UCi5eTB9s14joHiJoNIXunsb5yGxxuLRjbRH2dJLM7qn7AfiZkor3DqGHi4t4zznmpRor
rSemUjceATzAPAUDIJpzfoH/5Hf1ccQ/Cp8tEcMxluoCtHzxFu2KRzAAXn814mmfcSRXwwjcFMi6
7WdAEhKSqbp80g3d+cFvH0rIqJT87dTM344EJUv2zge2fgVtFMHx3tInHA3VUU2wumF+qLNXHDPg
TXcHiguRRt69nACL6ENgtzKiQ80xajMEq+t76YmAquscqaoWWcNsu5mYLbCh0/eX8sjVDmfvg9Yh
S6zW1uUHQByb7I4/AD84mnQhBy2PmOU98bIxPLIQhnPodb9HTeBRfyMkToAF+00zWzj2gJCyy2KU
5LzxCHfyqfomPUP8whhuZtaGzZ6C96AHjc/Bag88QosT3q1t1r36tChreAWhupQ3LBdqAtSuVkQp
ap7WYjjsNSL/lpfDz9bDq+Vkca1X+LT7fsFp9BUKaWqG5zFTFqcQnPhx0diawNpOsYOCU3lOQnTX
zt76J58BTOkKTaMwpMHtp1K0qHcKwx6dFJimbWtQ+hpYLdH/T8yCPkZVdBnyb5KCpTIFf9Jh9z6N
gY6MwQldZoB41sLwd3rp306eGdVtO0nwp1osTUbjw70zWaB0Ulol8rThtj52wtpV6LzXCGcbXkCu
wmp2JkaILytSmxAwaqOpoQPJPs1u1E/dsWcOo8nA6Iafi+Ru64EyMplO4qmxHMCvzbkeYTnZ/w8V
x2do1TLrouUJB4FJauiFVmwlTRY8N9auH/n9stA/7Mop+MPbl2IZHOYa7ebMAJYH+YcWTUywu3qc
H9FYQHxeatHkYPHkVfFB0PBtp06abNWCvXYxrjyzdJyZ2bOkYwUOdVjz0PGR8Prvip//x7gtrU+y
62ZjuuP3Md/n6+KROZalUwfsp8exoR7D4IrVEPaIJiyB1X8xMgyoYRkvAzggiKYbzvJsei1s1qst
SDCpQZLlUAf192CsYR1OcPtfv8n0iK6mV8HsTXvRc7wi7RID6x7C8TGJWAZmjcMZyKHGh3fE3iva
cTA1cNcxxd09AEkxqa5w89V8+owufySdY/1dNP1kTjGh9XpWbr9jk5QZlcA3h5kQ/2wUskF4iswg
zSLmzwYTyY5D2mTiNqu+/cj43p/FizBNibaX93wkxjDggREMMP2e4TA4bM2EID9uzhjUo1t5DETb
Vq8xcoYCDEi4F3iC44j10nMhtLR7EzakMnpzxfRY2qudaDVO8NZsGxC0Dx5x2lMv15H8fwGOwS8t
fkkHLL6diWcjLEJE2a7lEL9sxFy2HJcntNXqiBFz/8CIogZOxD6+BL25q0NVknDYnfwM1uHnrOBv
+8p2d3RodV2l3Y/ev9iE2zVEqyDFy1lZRfsedoYrqgDF1GMoKo7E+ER/RHPL0+4TqlzSbVeJrbfx
IEL1faUxW/4E33VS2kSvwMeILmwJ+gUC3OShUJnzW3LGncf+WFLIeF9IWmeODQTnhI2SGTky9b4f
Z9SK7dF3v2TY2GOtTxbriWpgt3gXwtqFLW1alDZXKYb+RGODasNegT/eMjt5pFAVmq0vDjFy7zVv
gHijU/Jp6IoAlCD0ftS0mvbUQgxN48se9A7yziNk2EuZaqrVYUARZ2rcA/tVJ3CpAVNpaAEabAu3
7BveKp6ZIUELL4pEgzgphV4ugTVCG+GWa95ZgGrM+P9yBSjof/8ESQYZPS8JVfIUhe2nxYEb+T56
IpcFv5od+2S4TFg2dmNCPMMr08Lg3oczCxrrtwE0RY9tdZwxGi62Y+w8dYo9/o5ysrl/Ovd+ktN3
uyNZYmX2U2jkW8s2FQ8fRABDZhrzloGYpFDVEMLvdkFRXEZLZicWagaF1ajwzvXc3TPWXM7/FwEU
GsB0n2O9L2tFaDRfq0lHQwlE/DGgA/OU6fn5q7oMHUoAzemnz66zRq8NNItZWQCmv30b0reuVqoh
VBW9iD64zybPd28qpM6ITFW9rhjR1v6RFGLX7kSjEyCKOjJmDlij+1eB0IsGClvMKq0wVgTt+pV+
IVuuNUfu1WPEhgnQFW/g2wglocaRracXNH4hTlvmhAbj8FS+elusI27hivgxq4zEACYT6DmSU38t
EKRr9iWJT/Y1Hy5RQLzaNHq2lvAPKIOMocLIA5XWnnMIi0PV2zvcWdz3mudmoxM6hLaacG5aiWXD
N1hZ4Vv/Wbv/F07Gsk0Hulep6wIIGX3riGwdXP0mAt9mCiGdlOiWy/cs4QoYfT2Np9LlQ0oXgFwJ
bGYyON7jM2ueiJNKCN1cHeLq0z/TMmGbOkksor9pzDGzDkzdYdnUYw+EbbCvMvI1hb5wXE8l7dyv
+z5Ic3twgsLMEyAzzzOFNqf+E69jFQy2CFnaQZLq8jZk3eV9rBAEf+qpHI3kIciZ8tKQ5yrR5zDi
pTjZgIHnqZn+KD9mdLgmlHS3V4ByewlcEvFUtfxdPY02gPjHZL4B7LlMUSuD/xzHhbOh1Izrujj/
RFe9hl+Q0waUyu7Qs693fijsRN+6nokxR0faWItaFZ1PFAjUOzp74nEUUTtGt+Jm0mzBsR2X6AYY
9YuDJcKVmg2YmxP6vvlg1AU9Oj7KdxdFHrehKMfaxoFCOnEV1tomIuXLvA+GoZsARiV1yZWA0pkg
1MK4zYJ/K6TPDeIcfQSQkRk/pLHukWkBBPeDHcXjXjkZXvxKXSMOsYWxi0IdTrZk0TMfPk02xjH/
rezcrQZtZ3D1I8ffGNXoU1jW4TXF+OBbVolyGcfX8Ka+Tifnuud/JSSE/NICwZsojWhYNh5Y7VNe
pNx4HWTbTDae+JvOiaC10T+K79hwW7USxQD/n/bDdo04cm1Iu7V/+CgwuoJDZWaMihvLqkTzvGkT
6XWitvcAzzyF/MuYlH3bqNTRkauGqjjI4UEGFjKeVM/9PSVPTBMbDUdg9rrkR+w6p0VVy7XCQak8
AfszcN+h5jZ86PiXncKZ/4t7Su+rrQ/+HesdbcInPmfG6kbbYlq6eqCaae4WNk1o3EmB1050HQpl
1hTTOWYTsO3q45GY99ujDBQMgVfv2CBL5EeGUuYpO7ZKBTpPrVhi+QfdFdM1u6pM4jNf/m7fKaJU
oOXjR47T8u5DRTmMa22YlvbIxdeyis1OqN2B5jzdiLKEaOjHCxiCWlnp66x7OY3lCUuPysIjyj41
e4PMbLLJ0Vwjfx4IvTcLXyhc2fHLeQ9zFXmZqyidrBvP51KJz4ntJdrQZ23zS7I6o2oA5hjkR5dq
ofovlN4edZ7+SgVtVXNBid7N4GYBfch0E/e/idNs8Y0qXeogtmz914tkTMauD/u0enZVNTE57zZZ
2p2mU3s3ns4XWIJ4iqSsVU2lrxRsmkfJNwIn4GDKBVI9WMfIUJa6toBsIpTQOJmyW6LszWuUtGj0
xieLiQOpJAY7Nk3U2+lEIjBk708MRf45+H5wnsZJgOVu+dBfPTmsrWItgRORh/is8q2J2qkOcKjl
9m8ss0VrVohhZqQZ0Cuje+7B9PQGjJqiJuzWBjliks8dhBTnIfs19J6ESH5oqdg1nA7VstKUrUgV
AJ+/OWSde4Zoyhu1LoBU0ujvHAncJjqHCSuT532V7i3JfFXG0ohsy/LyEmMBUDe+aN+1GjhMiwnF
KD6nfoSnQXH0khA7sP5Zb1F/BnbYVeID4JbiePGWRp9j4vRuyknqi9ZOvvQAgd1UlmVLqilNqutg
KRcxP/B8vAtcVO6zHTzYY/92aFYIiMW1JX43bVQTMi8AAl9Kj8GEYzGelMyI1O+xeycxxvc3NC4r
9PwSW+PmDiQqypdp4uNowp1FtfJ5gFSqC0liIQRkAwprNAjld+nq3xkiXDNEQYrSJq68QHb4V+wz
GoG4scyYdPSt7NBhNND54FRfa0njEx9psKPqc5UxG0Ccm6MUaRehpg57fADOgF0aXFlDNMgZxRgG
Aq2AQFhKOcp+ZCcLCjUdRbUE9d5Yy5/oCZqceolZT1h3mKTSijx6F9lnAszu+zsz3cH1Htt0TZYA
0rniI7m8lzbkarPpUi8gcLcPcjk5mVI9OSd8lqYztWjPF70SXxWzpMDNcsYB+CvPe+rLfWS8CjAA
5ugO0aKZbKelVObILcCLaqEcb5FJ2yL18XVpuNapGR4djFYiI5ExxG3hsmXsOweHMhbPi/jUlvgW
JPWBtZ5wfckRzzhHcNzGdz5nl4sWeKue1jKw21miCBYaYLU0bdS2PtNfVPgNl9N1uMDMkdso2T0P
vh3ptGX9wK1DOPVdwm1J9Bi5D4y2KJAReXH87lshnVq6RQ5NAYOB/zzVT5brquwtne60AbE4rEEp
1IQgvXYWK7R6gM75RQdXPrjjlkSkkOyTBZx4cXAdxhlORY0BAmyFcS830uRcIvVplrAf/QnO9UCD
seKrVOMyveR0DhpbvEgecVcJ5pLUfJCh+lOK6oHq1WMLKkbGFoEdW0wm64teyN3A6HP6oNNNQErs
UqvsGDX9ULvKx7K423olp2hSd/gYpHJSpQ5pjLeSrDRa+xWEN0ywKigUcVN2DQ7V/RR6tZj3pKrG
MqJ7mSwDlp6K9aICLikZWua69EPTYaPEUoslig+bBjp2UzGZGXv2yqldYVtpDxDG+C9h/Tlp/wV0
NW780dfHpVOiAn6m1fstvEnPruvlrFVklO+p38weiXuwejgEddDeQB83O0aO2mnM92Hp+hXtBj7E
6OeHmkrlRCsdVIlezQNk1p4fmixf+nzvMporudMrDzLqvYGFpLaBlAXz7lArbuuIEiizgA+BTfUR
q0MRxukI3RYjVfM4PCibExLmPZusfJ3jvgkH9riAG6T5BIape3DRLrdrbFeLVcXVMeBpPpCbrzou
8seVf3ZVDvfHUUlHmJ6VYZAKEF2j716cSN5SLqQ5Gfycma9SM1VWb4cJgZy0ofmNvrPhqwA/zNi2
lsg8htkzzCdEvB1BYpnEjka7wASTvjgGYDRmY3FuTR33DE7IJti7yPEBZL1tAQSnEGEP2mluPopQ
Z8/sdMNl08VssuPeGpScwPVlOHvfn7eOOUbpK0aIWJ6s0cwhnpVfATjslB1FNwgCBdrH6DvQJYH5
oLsVVZNGEo/HElMHh73fkXcf6XCGQyYQU9Wn3b/Q++G1OmuBMUCUN+p8KCHBT3bHC8L7jfskK2Si
RIfxrLDDMA7ZBYYEjG3VSp4NYR+nr8NGrf19PlD+YlG73ciaanV93dO1CTgPE1G200uKM77NnOuU
YgYb8y5NziBeBPL8Eh+Fro8BHvd70e3RxbvUuH6+5Hhw/4rHVLVfyVADM+OUb92CC6pHiJfdAoqD
ByZDw/ucl9L+iNMaYD1Rllt9GzE4Er3jJjN71GCbNQK5QK5eAqJQ6Ao4vpYRIzYDSGpEhUQmTh6A
v5ibh6rwD+B94dfEJFNbtRIkXkHHtUssb2sEX97oj6oWdG1/T5jy3qKXhRPW8z1oGDgOy2BGg5Ey
JScbXopMziiOA/F/xOSwMfrM0Ooq46v/mFFuQII53uqiEG1xrDgudFBrBF45t0xda+w8yOCqKpeT
YldWDgl9i4NXRDK242JsyY8W4GeaJYx/feNaoj7JxbJSNeEmbxtJF5BDI/PYzAB4Gx7npReEWVx0
lpdpcD05+MGn0sucMJJ2hAIHwn/3k4rBDVmKteU9t0X+Qvb/YzB6o/cuuTal5W/3ZAwc2oF9qfeu
xIc2kgGA1Z/RENrUYlmvZqYbW7ry+rW2tITa0OaCe3SsxOt9UYqpuXw7maaJ9/7E1zGsJZuuw8P1
9Nvujnd58+Q/iRC2ahbfd9BtALH7TknFuQuOiCBArtVJOIWJx2ie60sXN2eb52WXzsBErueniuXM
ZxZ/At1tFMWJ6X3eQIWfPYOmDYO/zaYPD0FGQG+7cwg/v/fSuSFqJYrWTtAZw26g0WT/CJSclm1j
7SkkQ0Xy3fnj9yosfzxRG9s0vVEPo9bEFxmAuIFAFab2hCF0+CXjLLVjWwGGYJjSA8Pt3p0KIAtY
WOUpWkOwpFMm7F5kKn1rIQi45VYR66CKmsRo2yskUJGYXXXNIISySGAqD6qPwqkbdau0Yjm3R/wB
nSrkkBKNrYfCJDlNHSPrPiaZncLxeq7WjZKxnoC2JkP+phlU15YWd9Huk7v4cnFaIVfcsRsxIe/A
tUBUfRDGvFldoa843G4XnbEwZDjuGre5j93qEtEUqDLAsdRlgP0dm8LyA3yDcOubJL4td8b8rQv9
rQbrZPA/MIc/X+YSqm+JcK9xIPont9sH7EndeqkoRAU2ObLGrVd1vl4PNj7HCmcirr/D/VnsnnIo
5aRcLp2uOP54DvnwgAPNT5FsliY76X8KLRZEVFN+AC5mpqGvcGU0VXolK8d0jcJn5GxBN4quTtYf
SnctFE+q8hfszWKgUln1RLjVtofoSsulrSy3cZsxj3g0tPg9ijAkKkH+1QkCerHkZTlvrdgtt9ho
2dD57Raub61vCQiRrN79k7a5hhry/m61NG2DZYxv5+Tk5zffAOJQUbBMquY4LlmL2FVnMfzDfHPF
BGs900p7RC+OBjs9SJ1D9LhiMcu8FY0uI21IMJj/Ztlsb9ucdzunndg7KUzlDbRAJAShCEk1/rN9
c8F6cN5GbL9x67MCTjXrP5RJI/SHi9earvPQbo4ZhdvRwwQvyF5D6I2oiwrpUAykoL8HLMEnmjAe
NX7wIQb7PnY+CeYIKEtQnoeihBXaXHYV74FsTzE9ssr/4fqjru+79gIAMG3hvrjKNS1zc4l8XbjP
ppkV0mhdW+W+8Xaf/fVsz6HLLALlb8ZDpgZ1XDCd3ltb+7tmln2gB2jZIjKR26zz4An+mjO0LR5W
QL1XNjPrSmWpomKYa/dlMB7nVeQXdiFFUobEi0CA+wJkJ20Kv/INyQvTDJ63iVA8u/j1ml8mt5Vi
sqv5xhbf0xPzVZVXzfldXeeH8zlkU9K/UYdmJd9hxl3PQHWhmfb8taPFjqKYpVU/ARTt0OHxlR3N
Ury12rkr9SNNmAgt4aL0oIT/gbE25Fu/BXKTYGFVjhA8ecvsCCsxsAnZv16eQwnc0uv8Ikr2x4/A
zyUuYa70hiPyaKvtWLIqq31nsMyXmbbjLBXXO8MG2kvF+EpZcCgJB4H0tJtXJDxD5ODNoj+Vu5i+
Il/aA90D3Fht0WXedY2f7Wx46AL/yKAHy5DntxZJSwohzI8IwzDVp2gmYafiGJI9CDC1PeCb3tVB
A+H4kJry8anuglpb2Gz9Rt435vsdsj2L4g+pU2+sF7De4q2ejvjLF1Z5qqvKOUPqaULoyf6hZ77G
/qcxlaYzmfTYLD9ZIMttJnoDkMqf8qj7dT/v5xu6kdsqmNV2tMMNgUacRBWtOZFmSsqgyNRBLX9A
Dq5FT7adxvy7LWnJE5+BfbMIS2zBzkqbfuoM1wJK321d3/xQyIG0gi2SB6Z5F1gfLovdKc20q1dX
i3IybNikPxGfRrXUH+TmXz8+y259G3cSbE0ajkpKrHArE3Kjo82GBYDL7MB0kbd1U0OdsJPtZ4D3
OJmB8GwEncRZhErzIN/S80VAUFfrnSgN2YZ7W9dGCtMy7M9Pvi2NxzZVYI7re39V5UGWWdFbXDhf
Z+L1iiGQ+uqsiTzqJL5chFcJ1WM2uJNXMLS/HiD0sIthyHM9nDiee8bMgPuFFXISY705Aqls3ctE
v0JZbGmWg2+DDGv4/pRnyp0P3wyKmgVk52/4rDWoK6lMt+fOWhfKd6PW1ZvAg1v6iOH2xRKQwdPL
+gbxcHlDlR49w2NvEHYLonNtQh7ngoXBfT/tpvySIUqA1WmtgfDUCkisMYs0X1P+jK9f7wqvkOcW
n4OKuGEtq68OoYWgiiVj6GjhovPPPLrCCx+43QY8x1/f/e4NoUYAa2rQF92GVyO7oR8rzImqhUMy
7Yaxb16sbWuYCnsbpkrRuW/2+VOCI91ZXufsiGvLqFLW08JVhBWT/rbghU6MQHGzJOf9htGoMJkz
B8BeAW2R4UencAoKTeppVRgpe7DYNpXmocSpJ59zpiwsHOxlzvZdLFnVlbQTsCzbQVTvCuZoJnFL
aJLE23ql5Ti5FQ+OgwQATwBjyw1TvfU6fAXKfFrIYg4tGv3stvhTRGiEPkI1L9micrzG5EOqNxkn
BlhHtWkOpkSyl2DD7tTDxrGvnh6HNPQfQcPEFF7Ux42+EtPI4ree3y8TlRrT+AyUzLuGm1+FhDV5
uqZHW5aOcB4fCEJC482nDDRIcmeZUhF47MiExIWc8+tFOvZuMh1ZodO9NqzpY4LUQZ+c3CCD4eWV
TbCGER/2koEwXmY8XV2GNOrJi7QuqWTrcqNtfqerlGu5szUnw1P15CtSw9WiurlMwHTxb1iWuWJj
kzEE5BVz3o5QUdnuPfXQCmiZF/Txt4CZPb0nWBVMOK3+shwjjOhSZcqe59pB1XXHhR9efgjT/hiV
ME+36EhRrFXJ8ssbdPJGQraLAiDgomfO/aBXwc1voAh01rAAvm8LZZsPyKaRE0hjqxd/oSHLI6f+
rjYgCqvsFRRPbuotRiQXHgTuoVASCSRqIrMxSkiEXYeS+2BJaOpuZ3XqkWHuuA+sXkk98Tg02L+l
SLfrQsIRB6FDEKg1DnKLe9pyEjShfXZKmjnFdAOD6+0BuFFBWRoczxoYeXwYJaRsKBfdyyBlu4wi
OO1AktvPidAerDnfrfRb1ZOqyXC7Q9+HjjKZLaBKkFtWXZMX0WSWocSudXCPG8spYidK9cs801WJ
tv5zbVC7eGMSQ8f1QBf/9TwvpYVwl+PN8qJhtrxBfMaH5ZjpTV2zeRWLemPzVXx2I/0vptjVBh1j
5PzJGx0mTTtoy6Hq3zbyp31sctHPXiAibvwrKPoGeTpjdif7A9+xIu9OeRJcWB5Zp5ZE1S93SLT7
u8uQgJtpz7mxErAzCwcbouqTPrO/IMTh39OKlhE4Zj8VEzWLBg2+CAa/jWzwltzI58Ovsg+vUsuO
x6yeMeovmdWuEiRykWwAl7eirFwXXpA0/eo9eGlj8d7tFUn0JnbmRUxuasZ3gVzHRiAf7sTU0EDn
i0ZjSADdXfne5wdgm+Y5c/1CDSGkyAoE7RKP8Ih2Omk5epRcdmLVnArfiypIaaMm2ihUgocLH4oY
XQSb7IK8EhkBlat2u450tHuikJ4Q8yWTGGmuJE81qQiQhvDShk+/Z4jqpCBO1TT8I9pQSZsNokQ0
j2C6r+n42+KnrgicMSoS8EMU48I+iuCbVzI+CSelFtUgXbSPWnU9vSGIzme/lD+oXca5t8Y/3dqs
FEM/BEQRZOE5gVYQ31hVWP2cIwPX8SjSA4Ziic687gbgnPy1hSNnWQghJmkEm85Ng3dzNmzoIbQ8
NbBzbUDZbuhrwajU8hPztIwBMMNLi2Lr3PylWlv+0iwYkNDwoUf+dWEblZm7SPgBfJ7oFWam5QDW
ZIhcMU/eaSU6s7nFIy/uuJEJoyI0tO/TEkO+v/YP3j2erCGKLOJ14RKRqso9Q0ewNmQ0GDXbYBqZ
Zu/oi3BhJSFZ3z8fySDhmPu1VxEaLzM6LEgtqQEo25UyJWRKVBZYV0wLGjseZMSLEn/+V9J7gcuO
7AiAPBDhiZYudW0E9guMxo1Iw/E/bNWVBBtR+3LGLGA2i/5BiDsAXAdJRjXIRyj6UuRhhxM2xocX
YvNGwauMYG7+v715g+fgllt1ZbMcof5qBDyNR+Rk4Ecns8v3TBkR+CcYzYXJMAuqxcRpwHdtnlnB
57kwn64yg7/iITnejaaR9huo6sxZILjnqILsoIzX2mQEEobnlmgY5GUmVuSz+A2rDJujtG1iF0IN
icKPR0/JA+HVj125h/NtnUcQ7cgllPXZhCp+fpCTeUNCU6HBXGuUZ9wo0iBCHStBWRWkk4oP7UPE
vmwFQkGDOBClnCIqevnbFdXnzcHdUT0cXTK5SyqXFMBztT5/urTt0ceEcSq8EDlLGXZh3ylBODZq
jl5jrypPE+yGZO8La6C60WoOY6R28F14/im0SyhYm67euUMIq4C6WtSGREQy0HlIjmkwHpZ0p8Sq
9x+xhKoCBGNtXFZ2mqPHxPov21mAfldri440r9ngBQRTcFPzGAZXYT7cpYuL/EhjD93jifb49w/P
d7F/RqMEEU0INaB1mmjqKUby1XsKGF+mPwNeJVTI2B5sYJgSJIbbVRqgfLrilt6hJkqlsqa4N8YN
/JgEsNz9uVMJho3yrlvOHi23dG2Uky+gtT3wGN/eOjOaWlSC+gl/pLK9gRTOimr+crT92X0jlWY6
fdl1pogAh2CuWEpHvLDlYLOe8KIhZRwUVy71JwHx6gsxQqGbkP5IjKuW+MkuZjj6qNqGOPMOGN7R
jE7OVfwWgc/no3+A18BbG/hq3Ff/h/uBFFErPta0S8DaZuBDwlv6DPUnQRQ/DsnId+Dpw8PzJVRX
9WmC7yygm+Z7tF7BMTXLUeJbSDUOykzUdGpx6ZLOw4qOn3Vbrp7tc2JeHFMKK95mzhT9yM3rQ3hp
239pD8jYnJVX5mM+p0jaxQpMIyWtKSHKs4WZEj1HaweXFGItg21rQsfBBEmruux+gU0MOjKBfXX0
nIhHWOaJbo4TZ+VfWc0zASGqHb0RmvaeUPKtOWMInhT/0gAAEypP2xmaXwhrLspR7d3b+Qx1HKkX
Ec2JzRqYtEsY+BBAjYO3VEfayatyzcWxldSozYktk8LHC2RvmgK6DJT8JTnCqNDJL+jhZL/g+tlH
qZrajA+C/vwa+toHP3s5OHDnyugEdMiK98we70xjNCcmpMztAouRr4LzQ8gpBv/tkMm5ZNqAlDew
pPsc1TxO5rl1VaSawpMCEghug3HViYsPg1YSAyMEyrxxvtAAW4MFNSIn8tNAtq4lB8XkZzTKJt5H
+uXIcuy4B+rFL38ccS+sALdvxFmuoBtlUXLPd8eCDWjECQUif69ASbwJYOlAqLTrXIQF1K2Mm0NZ
KJE9E567v68IWoPW2ZZEH+4ROxgT/y9+NUyKfBLKN8GZqVlYnSztfn7yJP7ceZLkgNXZgVitc5t4
lE/95KheeEWPmGKlq/ZYOOmKqUXlCwwwR64u8EyTZrWNCpFmb9uMKiqtUGmk1+qwcS5uVvd/cisd
oLDpsWVmsWlNZ6hnmzhxfaAkNTiNW/xbIPwKgiyAhgYVdvGQkYpV2sq0MzQkLdTutIAZ4z5zz+NS
/larjkNS9ys7VyADhc1TWcTTh2d7z+yxEh8UFIW9PV6pOuembRwWxL1m3lrzNoj93r0aEGKuBB3P
kzRkcibtbJ39Pr5Fv5BDuzPw3YCsvJAuZnFHz3rJgj1ZSIWF1ijHEUh9/lh2xg4M0jxQzOMFvh1y
+dbyrKKReTTgQ/skA37Cors5rWaa+kGdn6Ll7l4rt3csBO/Sg2fOgqxoRZlvH8gnJXZJvplOE72a
aZ7hCclH8mZANxq4tRfU8fcfWghqsa6NNV9aFdcGe0D1rtmJl3PyJK8RS3b949Zc17ydy9Y3yztT
2Mbf4L5Pysnq0V+3RW/XfjmK5qwhMpW8ZlcdMfoUUeH+h7gnqLqs029pQ70Slr4Rs3iEERSuJHQe
2xEr1/yyJmL8pB2fh1/6wDBg+wHbrQUJXjYMYGbjlBQ/IpDIOlvfCK3SFLGLUYWnfA05XyPxAIAc
pk03e1T3jX5bRxf+fZ/iH0a5wy3Yw+NcDJP3bIdIFkYIw0NYXcCEo0pwzdfaF19PuJVaNuPGDYh5
hZeXvQu+EP6PZpMtGKy7svdCyGB/5pjLbQ6TJUCE4NHVsXmhY34ad3nychZndIAaF0K4Zy0N/w6z
4W/cPD8ZdQqvfiBqjRrmATfyZPaZNH8rov8hOOQ6NE7VozhCz4LXL4SzR9vqPZWxkpU7EECjYtvB
1hB5GK6UmPKrQVVkmT/yE8XIJwgDnVg2YlvTHXeoIuimVTNf+937trawT6lVDgReZQt6vOCiC+Cc
XgSy49F9wQtBPa+yUUzV1RiSs+Jpm3xnIfwCnYU1cplxDR9azV+t9I6P+XipW0mXx4fvIaNQsXdO
0uu2efevLjPVwiXR5VUYNFXABkQhbr15T4mFeWZnDWOrJXmlOh0pJ3cJWaeaYGojoEx76rIbCgqR
ggqOL76cfapyhLtfI5hvc1SoDYWm43f485sVNVRHJCW9Y5CvPGPirsw60ULx5BqXgieO1+T7E91e
ZgGSJwH/mJxUq3wIYAXCk95KDAWpuFyQaJBAACtUL768fKbOIf+p3kvGfHx9lX3fB/p2CpvzaT0G
Hy26u37rL3JYYCjavCx+GljDTVsInliE0n2ENUWntN3Q7mUFHEaCxPEGVbvTXnozRLhJ4ChCHrPS
MgQVJRa/AVHWRdZv6eswg6ya/Yp4zQ18l9mmQ6YCENPFQDyQTYv0dcrJ+zK9Zm0Z3yS8cwchVskk
Q43iYc4p7QKAwu9MUleHi1lhZNO3WQ6LWw82vWqJPpUyyAObmn+cqjLCkv/LZ/jvjIq2KkceZdd8
4v2svE1Ow8iewIWuMoCF3FS5zryEM1NkjtQjHT0kBshCX2J0Mw7u/6y1MgAIAXisZX+4UUvFFbaI
GCL4JXPWaT6rTlDYusCfoYPm09XzGUmSvkMaPZ3RMMD31NJ650tNTQdq3WVYlX2+ipNzgGEzHf3g
wWvo1pTmgrLAoKWydhqS44U8JaICo0L3ZX6N0+B/wOZ+Kl22jRw4hr8rMxd1T6EgapGqPCG4uabi
GP5Jt/Y9KYrQq4oc58jtDBiuvJxfx8MBvwG7exumue3X15EB2+UCu8atFlduLcNZmdk55t5jrMVu
uoJ5Btm0hE7zX2wd4LaKucw8WuFqVpRxVT7cekOFLAY0REyKCSwB1rRyFyRyAGz8sF2lw8zeQ/uK
zitxwnXiFB3mDUAijgyoazRpFKOM3qWJ1L+ooAna9VacccFZQU+AfcblVe9byLZutr8RiYGDpSL7
UKFFyXHHaRqDHDs0Wcnh/o0D65Qc5E89hylro8hpK6uQk9mZIXvxOmJLgTs5cKKxlw607wLx4b2a
L8oNL4DB8g76KXvfinr5B+IyzokKV0Ar7FsLV/430seiEQRrByDTc011KP1Zxto2rN8FVQaAhZxq
djleiU7BmR5aeOlpEWtSA7YLEJGtQHb92VeUDHICS1l+kI74r44hofE4jKDMEEeXjDuDv5AypdpU
Dz8rIb2Q7DIcWzhvMkNRXf+EEN15mKyLd4bmvHOthg0lqX4tn8dLiVyT3wMbLjIiCudP2q3k9HRR
fkrI8fNci9fgCsX6VjFs+8ZtjBTEk5mVWia/9S/jPTv9Jdh1bWSN2uzCbDfpigjqJdCkP3eKBdoH
HZL99HTpHHaTL7jGdBizQZ5/avn4NMgvRk7XTrPZB1ceFqkWr4SWlYCpB/kAVR8vFOdg3nQakHCB
qOWqN4EDjHUpdUD9AVlR/Q/bJf1B9n+1ZtGf1JEOsQi4+9Fd1H4/v8UiMoQRRqn+EItrvGCIYSKt
R3edAZjG7XfifdzDEoEPHAx9OuTER0yLPdrIh2m8lxA8WfnoNgvtao+0b7NsIvm2axGktos+G+gx
wnmt0NJyzDkb7ewe6P16bP3ma93Yd0NDYiKNYk6fX69fpwWzptB3/u+fSqyCoNoDWDK8T3hU9D6b
8mWGtjRC/0VJoAQuhG3bJr15IAUR7RhEQ9XD4Io5BvUSvCyfpFfytjzPHYa4RWsbGPuqvUHSu+ZN
EfngP/rFFCGsRP0Tee9WoL5ap1LyFXu4tNq24uBUhpHF50p8kYGlzelr6g/ZT7SjvFZBCqSPtKWa
e0yf50IRq3Du9NDLJyES1IyM99x0bGN+vI+JKE/eswNO8CWc32oQwdf+GS1L7W7m1znvcgPn9bke
3bwjKupOmAYqMR9Y5qafx5fUgHpV5xgq/OXrgQheoZBLK4f/atYqK2DjmEnFAePIk+H/7bx1dIpK
1y6sE8EBlq8nG3Xh6eouvVTe1Z+CGbbBuGIyT+lZHTvMtOeTEou0e4ezDBiUFFgc+THIuanTQ2cH
hHFtWDye2YMWsEP6W62JHIiQj/SkcF6FcfEuCTlNIWuIw0iPgYBH8RVh2N6wkwJv85U5aeqXHcGM
JF9/GfPBFn9U2lKYpeyZID7Y97bqOfNtZYLFrgLS4ihyyQW0xBvTadC4T4BDCAh5EBVdEpKrDv+L
Ntxw1H547nCpXT1O5l1OT2itD+cRGFm0uxnzJvx6DcV/nqTdlYddGKgjJf8RF7wfMlwY2Ake+hjM
hCdxoGi3TZBk2qOVdD7x8Y7OT0nrjNLR8D4lGPssEMN5SeyeT2nj7AL27wMPLuHlY1vbbcWZsCie
7ZYieKSL0miOxsM7bvJ5YAIEX4uLgGqok1lNwk9WVPyCFLqgQwhhAEkenTdmQ2qiEVtW615D8ITD
8isK3pTl17KNqsTkEcI1/PPV5ULjI4zHyNAzNSPCcU/RN48x3lCXHESYbuVyGDvUbXp3OAYJDoCD
MEy6vaIvy7aV0ljNa4zUtj8mp13pXxhRhARsDwU02hZtGIpQziIH1KcdYzp8KD+OuMIJj2SJD1z3
P0U9vdz8qTUMop9nkKl3HaAP6LMVxv/ja9jExc3CZLZfbuLoF7XNjBdPJK/JuhLSLL142ktEFHue
OQCQ6hVhCMMAWzwphvDasCb03xE+EaZlfC4yO2bCrPFmazGxVOkkq05mEAzVIXKwVIR/SkFyt0K+
ofYT0dnEOiwgIQ8IjQPO/op8srnIw28stwLCs1/tyLAbTBThMe0FjAE4ddw5+ShUSGGRqUXCG/Gu
bReop83V3FOjoGWHoZ8IUyQUxuoGk9PgqM4oXehA6VHlGRTfpvfpK8uWpYZBelC5jFl6/RHhw2gO
g6T9DDdhqnbxy4nHFKBFNmpFxmWFxx0wF61qBnetCV3KtVhm1BQMf1DqTWxa6+CsU6jaHVRWqRO4
4P2jDfCumrGkLy8aTD1nMLwyNeVmunA9CVBZVLRZsvpKarxRbTn4o/IAQs1tfjrPaeL4a0Cp0THY
KfrPG+OwYSHadZARuoJ0gTbSOCHZ8Eb5nZqfEjcPTn7o5e4SrbF3L7cdzhZXkBvqosr5i4EGufkY
TBr1BD2Vg4IzHCb3alvRQpsYQYm9Jnt4G+pa72bithJa+rVp78WzaZc3yuSJEXv7T9FmCXTTEESA
UcfXPs/+L/8wOY6b0P2VtuZUTbNA0nxTF5e2W1R5A2abU/ClL9sN9JbqKGHhUw5B42W7i7upe2to
eR3G2l5y90VGL4iH8gqyJ56JlBDyl5j0jsrZgInlT1guvm2m71dn3jJ2UlKrUNwZCKwLGSPuc1gu
5Vy2myhqer3ZIlATSULaZ1arEgxzYwgpvpSFdG7kfvZ+/vBYmRXZpuhKYr8lMoNiq0awS44/rn23
0uoGJXM2AoHht6vkPyOX3NgDYLJiN/Uu9HOWust+YVQTXgLz5aYsLwPB1HBKsQhOa4Wiu5Q/uJB9
mKZSN713nXIzaAjj6Kz1EoYDSYTMjSnXtjXzntP/m7UbU7erHo+egv08wKDo7M0/VGsIYKxJUvLq
1Zz3EZjIuetv5YKI0G0xpjhCSs4CSfzutI4mEW7gwrPRzFryfetocYOa/YnnHuexIXX1eMW0nSj8
9MgblHldVyvtRsJYBqdBRTQCPydUXR5E+iHHVEhAXaQXhDxWb10DUhkg2KSI/3Hp64qTOlzwVVBL
1+GvIvEOcx/TbaaYTVvV852piz2ILtEa5e2u0yJr4klnRv1IV0nLnUn07nQ66FiHvdi66C1mQAeF
F0GJXmFS28NGPgLcnUnJAF2laZjsv3fJyXg9S4S5+oNXmr1AU2n0RzQ2f2afaVqRDPMklFF05tqQ
dJDRq6EP94wBdjrjviB1LRS2e0ZNlIxauz7WBVxGK7cYcG4euNzJLaY5rxq7IjdXZxyAuT0l7dZn
F5Z40ZUXMrLt92cdk4SyYazKGPZL5qHHtUMRJUR8/FKS+OZYSXhLrJxV25vjuQyS2/6u5GpWfrGH
G5jQpeKwo5xeOH/LUU+gB7h1V++y71XYofrP0mECCTw2FFfCrh+HMuHP4T8+9JakAFTQ/BocKq5q
XZfRGllrpLR0tbnloc1fBCA7H+Tl2+xWFduHZ4WdzODljbA9jbgsRJQ8dbwRLxVZL0bqP5Ck9/zW
hE1aHAUkrhnuwCrtCsjwHF3ebYTTxl1x67yxY3aUkjy61hIGp3uBSHGEjl5JDqctBsHNyx2zZSOt
1X651NduqZ1CbPaMDfaB68yaw8QbnGOv+/MQKlLgRTrKGNfKK1nb1RJ9IKIaQ0uOWMEN8DmOfqZr
XDsmfyRkmAnqVYQx+SMvRqLx2rDa9GoI2kz/yub/1/U6hwID7KkH02iwmztLjc1SxcpcZyt7gLAN
KcYyIZ2jdJrvghv3wSs0OtBnxLpXRbyG/lVV9O9IuuF58itoA+Pg0DIKKLdtVlx4sqXfCMDR0MLO
2T+gV33MXWMrvWCnIOCiMtShzWUTPg9CuTe/XO84i5i7egc+Hf63ONDVZLd/HT4tRoVjiP7Wu3ym
oNNYlaknKgAyy+0J4eTMWkoKzjqAYCd484/n+toUVk5pCsGraXuKmXq/FHda2gYoQ7G5TIKY0GSS
hQ0KzfhDAtn+6wUH2ih26uYkMZp2tQXtCLqp8kdq2WDYamoeWY0F3ga33qqLJSCeqlqI0iTvjIA5
ESI6vwIb1xtlTywC4oD5hxvWiQYfzW7Hazm1MIqVOJ2HGaBJ4K6a9b74V1YcCFnS5or+07Xb6sJk
JQFo1EpYXVNk7hf3wnl3aJRnR24FaFxh+xzyfJ+eEmoMEJhSVrxjx4PP9NIrBAIjvfHztAmYCpeH
8H6XFqSM1bkCB4qPIRCumavw/+NE0j4Gwu4dgUjlWe47g/mc4pkIGHHmHhtuTomxE8wmEjwJtUmO
KRyVCrGwDPFpdMSUhLid5tZktydnKMAbKmqPHSdz3+7i78vA8N387AJWTPZhIYTFwrSW14CfWPmF
f7jXJUS6qrAk/CTKrzMMgkIjsdprTvaAMBXLFA58F/Id5OwsQSPFs043Q4BvfaE3/1zGoydi+Jkb
6KudLw4J/J8WzXYJreH7I7KXN5NQ5j3TPf8VgAYOoMffs0nphZfSR6zdUAvxfYMk9XtGcg3aDICF
HZb77jr0Nj4VDhsF3m+fDcCZrN6IGvrxIDhSLV+kUZL0USiFerynj7m8f8dqZfg2ZcWNTLQ/CrNS
+OKx8FJUcEcQ7TWdfLejkii3LNuU8RJzqneHv5Cp0WkEQ8s8Sw65g5PaxS2R4cUhpQAbiuX6zS38
oaPURtD5mHaKvv9H6caTpGcXRnPXhE5yOz14c0wS7xKvGCMBp53cIMi2Ff1Z7DqT3n0Xg5nAas4D
LUZlY90Tx7CAZhpZlkOkevhg7nP+Tie+ZMQ5SCd+48V1WcH5Ym9jiFos56hR5VkjJoRHpElfyP11
FLD/PSZj/yzl9DLlvjGH3cdxARXUs3T1cQWcunQ9QiJRJLCbFH0J8Kc+0PH7qaY3OkhlQMJ6sSMm
L5BShcZGYu3Zf+2dRZD+WJCP/EHBIUnawf0DyM79+L/Hz5jnViUqYpLhgms5GY80l+FMO8qJdkiq
4iHumneZxHw0Bq2KmPODEwzcsfgX6nKpDRjb8QAtZDEuBB1JDeHcl6rTxKLXcoG3DfzpWuw2JKCK
D4RYrlieODe8f4hxA9EqNuobByOuV++18hDGA3kRjlGdoLXvm1whlo89tZ8FCS6EeyD08Rm5YMzm
3fygnQJTfGNJzKEAF4wQzEj/lP+9Ue1YTnXpd4AqV8othstCm6oiTRa3LRxZYYY05PwydDSQoIUu
rSqX2106b9WMwnkNEMNRJ84bL3+2n3umLN0S9VW9oDHJyAE7Z8LB17SAuBFtVkVIh+iEn+M7r+Go
BshMgB8nqotPB2mFOO00ShToP+bcuiphOXi9mBq59vLpf7rj/VQIzFWCf0iDe1IWyZE0JpLkHpaX
Da+v+BMSgVbxh6k5U/y3iY52CkiWsaVBkUEAdac4LpqBgEOnqfmcdOeh6Yc8t+6D7Soq0LWkXFlL
r+WYPoL4tf1H+l980LhiVMc5tMJYr3o4hsW+HmZyASl9MDhaiT6T+qSIQO0qUJ46Iiaq5913Owdf
ERhxnBNTKyzgIizQWdUnkZ6gG2l1EgJhNTt2vTUHk2mxn1zbgMS630fbdzjikeXqNCzsCzzF8dIi
9ZJY+596UcDKltBvpFJ/chih6RQtMmRpBWOT1TR4HOWKxcn72SY7wKeTWT7zLj5tMsuabavsmB6i
hxiWA3RvxvZ0XvmHdbM/BrZjSpDYmpHDDmXKGmEyMt1b6p9jgpx4nRNNlDWuU9qjdAc8I1Z0rc8u
9WldfZmm67y5hW3eM/W7tOqQglKQHHdMEkG3barR5GVW8xL5UlghlzEYoahD9sgUaqxObey4tPF4
ERpfElSlFS47GKJhdWxBM3elQgDn9qPe2kh86eo3e3knWi1vhpxNGkfWS9HbMblmZq9vanVViifT
Da7qgVAKjsfgEwCBCRhg9JK9KuUv6FjrUzvU0LvrVQrw0QeIuve603ajMUrL40PijQPRcWGTwOmv
TZpy42Iwnc13Zsub4NmhYCAF+L3NhDXHzjYWS1xFFNfHVpq785e6H1flQ4+LvwP1Bo0q+R336Oox
1PfyNbujmofQ6AiJTp+TbE8P+L8zqfyn4fV+DCXbz5lp++GVOJrX3jwB35TCCK4qUgfifjAWdfcZ
9NpLNVg1ZDCbL/SKHAPg4w3SwXfD0e10tnY8qELmakYrKV4UQ1tTfzgl8STQjOijMB8ljHKqZVRN
b1h+sZIiB9F7GhaP7dLSlFs7Lz+tp3CA9efSmxJcKRGJGeVfE1TG20gx4FefrPTe5aYZV7UBIfxP
4KRVjj4B0iQ8B3MBq05gTX/OWYZu8//d/b50CDNrmBMkioEm9npsLBn4fAbNFHxatIYgmzSROlYK
6FphQV4nEl5JMFJtdhBlsLyLyRMl7XTnRS1JidRG5TLp6Pehucu+CM0yL0qRP/xcqSiKQ8qQfZND
Z+lfAF/q4yT3dFopHXNxv1qDE5zeWk9YHcKqyLLVvqu6AakMp7fCoTn6XbkqIMBUfKwetYZRJoZv
jzhs8/G1asWVooEoBw9UkThJT9ceGNnauJkWiM19U76u6BdHqKT6n7YFtALtRLFUwoNDOwefdNKz
iZm+/Od7rYAaOtMwBjwzIcGcFBjmr3M4Cp5/Lc8wVd1LaT8cgOaJiO4wAuL/YbLsSFGolMOcFc1d
9xitoAqgQYpClZ2ygxrXVrxfWHAJ7QmAmZqBxCNCCWite66got6/K+p6ic/35N3zGgsz7YlDWFKX
ptgakAb/Bhn//xK5TjjYpgiWcYjaW0y+qEufeHE4fe5GvUAKdgljTknIi86D2ulrzdZ1ylkfpVUM
zyK88Uu6Cqn0Eud0dwJ9hFSSgxaKqyuiGFfQOld6X5M9vYjvrkVpTVTMznirj3BR1vQxbabCJ0zw
l5+7borGs7RQwIVKglSVRjKGGsIIg3akIwmHyQhPV4nL6T9vNLflzhNQD8Z6WDU4fTXleZC5BjFH
w5GeFTVYvXcwN6rpexoOsGTR1TRLXfDHxre4tuJUkjwPC0mXx7g+uoSH0r3QCZ5IwBGGPhptTZFN
6Qykk6/rrtDBNOUuoyQirFLmn6YRptWBT0KTvaPKFtvNo5a3LLHA/P5aIZJeTpfEOGwlXI/WqP38
Wxbwcl9+L9mQzdMZ1s5q7VvQsAZ32KOR0Kgem1wOtDkobk2UsHvM8bg1MfDuAdYQf3WmqX+0nYQ5
EfLLHDARgRckJewtpwB5f1dQkVWwXvIL/6FDE/TSqieW9mSuYSqKFniBhanQ+hgnf+nnf7GMC8+C
Vm52hvoy7Lkmt9gBsqWEs6FkdDbwvgeeIaq2YYvjqEde9/tS656ehw1Mul4ct7Y8/ex7z/gcvkxQ
KW0d/JtDIDtuv3raGklcZkmY4h+rDOncpQfMBphuE+ZgnDx0sI89IRyjDpht+sBo2OQUHhXCREj7
akft5yA7ACutZGJJtkgx9rR7VfX09ZQ/QTNun4Ya/8bgKnIgCjT5zjiFaJQRXMg4vSPSFukbhicR
E6cZTWmI/CZFr0UCg5kXBTrqJaupunXXXWU6AJmY6SjH67OlfrIX1dLk+XgeDz/+9ZPqnJI8pKQy
V+PzCjnAixHggak46PqQcHx54lVTOQbqeL6/a6dwdcRla8hn1GgX1xbkKBdJxP7RgJe7wzplvHkh
ngqaOvagAsJ+1ki8gP7ku1+tPpOvGaDV69fmAXoKlQIYMARXuGVEgobBrssBNO6uMCC2HJuiPB19
a6jAiftJ2x+KZKdEN9DLKujDUDXjPnlENcxim5BT08vYL9VPzTOC40/wN3oDx9xORAQzbDd+aky5
VxpC32K2I0TDXD+zNN2VMkfDRYijR1/kbtclcHJjqEMSFgT2ZP2X9198z56R5ZGVRnZAeLiyx1r9
RZVI1/rdA+F4g36TsjHAAEfGZ/zbrbr22Yj8u55vSsPFFX4lTSBpvEv4RSAWQp/aZMpG+4h8+2aM
jag5I/48vSbESsfsuuVchevMdcBEQLgPtSvU9nBgA3Yb9gR7Ug7XFz1DN1JWK2kPonsKw5DKfGeK
F0vvpZ7P36HWPriPfXpEZhusFzcLxf/duyMu2DCCpivficbUgPkDOtHwoDiVd+Gi+vUPVK9nJ4UV
1vOzAsBUCSHCsU4D0Kr8U5alj7GsrGl+e8mgFKho7Nx5hLMBuuoGE48OsgtJj04T7b4fna/t2mJ/
0sBv88d9YfzmVAgFllkDv3p8sqswyPnRfgaqWCJp6OX/06+U+5fQauP2ozYMhSShMZTtB4wiYDYa
nV5O0a3FKKeFTPt1NqVWbXxf1M3TPWmPt4+i0n4DuLMQ+qjRmUqX5ZKZuLRof7nGaxAJ2L4jrOn7
Cs7RNCyrWszKumIQNrFXkpVja7X8GAd7aEK5cTuvlVDDApyVczmkPUftA0YJUhem6uernhyKXwdc
ITNkDipuVUZs8Rg2YcUvYpDQ2yX+LtxujRDyZUQGwHUaELyqkECFDLk4meWBeRUsBRdQPAU9V6gM
QxYR3vYY4J46usVZ2l+uZXyrgWpxZd9os9N7ps5gMfedsMv8qAjnJN4J9qbEDKl6zrm9HBn9WybF
kipyRwY112k26VAuWk36eckqlMXYpCckU+1YBDIyz9ExY2dk5Nj9XWlsG7DUUrpqn6uQtUTOnm/C
bQ+ZOLUjXuM8f9pZOoSexZrWvGLMrRiX44ml+4TaOAoGgIyu+1hmsjjtSHkFdGDVF3kUzqHH8TRb
DWmT+i6N+s2JJcH8fjyq7p7oe+ithabHH/GmxqB9ZSv4QuA7t5g6oLGJXi4O1bhan+MUaGHiVjzU
aFoSroDkf4hTMX/gLIZ49jAQXHbSbcxGQ9bYE0FXYqhGpoodMKmAbSvMDWvGkDRq+c7SJ9Bwzasw
5JsQgHuJI136leWzuubDENgajj+3aCWfyafLdGR2DEiAITwjlzlE+U8F0K5LLigAn6ULVBf5nbnZ
2c6oax+5UlCQFMWAacfMQujpK3EAU73RP+Lt7EI+KIED83Uj9nNevtDL66Zl5JPCPGu/Otz+L0+D
0sI9+qrZbFe2wafzlRGXPrDnb1i5oRDLv2XKyhD4ugXa3ISfSoeSB9I2WfVXSFQXdrqsFnAjTpPc
PkpRmpjbpcW7NkkCrzhukM7OYUqvxdyYnG8ufsHake/rjps04kzJ5DM7Sj/bfCupbAg/oe10MrVM
++V5+Vfy4T0GGnK6n1kbpV7DV6uOW0BgUv4qDNjT6TdICEXFObdQdt3iK6E37hzBHS/PXR66TNBI
UYQtkTyelzog7FrkXUDUCaG5o53VR6X1VibLsHfhwObc9JajkhNb210i+mbEQ2JQVWfY4hdEg1Rw
hhT86Fdp6hbLNtp6vBtOaQhMlx64OJ3fNZvcrq3vSMuBfrDA0wfXeKyZojvBhADxe5lOpWYGB3CZ
YdxO0/3MA9UNByvBibYDyEEk0aYpBSziy2UCv6nXob4qexNvBmym9dckjIbiMEBD6QN2t0/KHgxi
8YqGQ5ry0GNgBi3hzorNVbdHjtd2cLNgXSZBNSjHg094h+LpHsVAx5WZ+GmeE8IweNiJG5EyC5rU
Y9KZAz71/1xL6qf8V3DRWRSN19Ub0eUTNjG7milSVjJNAJxy9gnF1nIxWaXFGTCiLSR/x8fYi4Qq
MmIQUZeZ16+CeWvFvqE3LUdWYceQTSB8QDcSTFYiCKyBZiewyOpVXdc8eDaotrLffAFkaZa0AN4+
N/9SunxBkz8mGscOewgpwg5oQgUoS4gKEAWfFuy08gr+o7rbxopS/tjYAxlzrEow93Rk9J6IVp4u
86QSJ1hINnd7PFef2fuozIUIhhD+sOq0/7VfSCQxB6XcXr574yLoJBllnAlGiAkOyz7TsxxfROJV
7BxQ4FU9rjcTcsRZ7ja9QzLZrimLoL9P+E4pbXRfwYORJrmWlFP/uKGi+zNwMTzpRfhLa2yVtzCS
h8yCT3pwtNYc+vzaTCCjpKLH7ZKWz0VHL+SKNWCPZ/eZ4jbkGVv/t8+23LuPZgVjOIc7aUpvhko6
o8KyiTcjFJxtm9cFj4ThP1A0BU/gSNKA9x+RqLjIH2pQ/LffT5d772HDzZL666rek/D0Ohj/u9bc
vV23cfqnEVfkWngQAUqlVZh15QAjNgZ9CU3ojXXQ4rg4mE/nRSaUpQAbTaguns0w4q0HYFRydc8G
8y7MeAXyctcShWb3XL6g+8pTHiV4jftmq71/pS3jITyf+tzlAMlOUNm85a7WJnOGZPfARaRr9g4y
idfYZD3Mc9KZ4Nmhp3eqCsYnMAdpSKepEZ7+MRQhndrQLZ8XdvUeC4w1/JhDLKDhZ/n1G1f2W8/c
R8XOK1cV3GwXq2Lntn0quaX3QoJ8tuvGirRWHRsSeGpR1b0I2xhYHOjGBCHATof20H6TBplS+uuS
hiBqP65d4NQQ65YNRGlZcQWSrlONdYUx4ttx65TeQ60IUAiRAhRy75WAD6m1Yjbz0mjRrVSzfqPf
7RltU5EJeVAw9L0r7MInCZ35wLX6PHYS0Be/871EQoCjHoYo7Pp0x0QBPJfZn3JUb5qrfJI21tXI
m3dlxP3c+0EdeExF+BnLFsxiP3/ajOzJsK+dvlqw5VF3k7QZo0tgXuUP4BNAz/PnitvBV42zH71x
IxgK66UR6T/B/Q/uJpD9mPOwPDrXcL3nVWR+Y4jepU5Pcw+NelN5xgdMDroa9aQD2BahzvdNNoXn
lWFboHlbANX4wq7grEuzPLobk8gQUbTGkf/IH39Nxtom278VIMci6bc6xKNPcJ4rHz+4OhXIzFQb
8FnPu1cv77uw/WLs1H3fmXbsERwG7Lft/OKVxgukzdf/84cKMsvX52ze09a6AMWQVDmkp4IzzrXB
vJdTnmJ1T3Kk7DMhUnAdt1yetIKQgEx+M+tanXNHc9hwVelAEw/bHUjMq6Sx+0pCJzYmimW3ScMc
8SQ4KbpuCArnmqt+IdOG3w6Vc1IMVQh5FMrIpySPX79evOfVaCbei/EKuwcq/IOgZ4OsV852Wgym
IwTgynmFZRjpsQMSkVk24yTs8aOrZ5Q4hh4Xao/KAgePgJ2TgULFwDBL8rBtVjBQuD0lYggYqwD6
SsJBhX1QZLc8tGHpFoJGHE5p8ooWqYutgCzkgfZfvrFc4rlzLq6tWDSvcRAZJAx4KNbve3FDbMfy
yPJx1ruECzvJKkctLwp46Wt0eMwId/nb+APtWQcWsn4EDxSDa3xKvW2ip6Dq0UUw9KTJPK66ZGhy
fnLlsZ6X3W12yCRkMh9zcUT0FoiptBl7VUpdYNl7C+ejhS5y5OIYsyRQk0ZkvzCojktwoNLSiW0q
IA0u39fr9raHGIXBoP9C58ufqka44hLH9p/ZjRdSiDqjtc4t0NU0yEKAVqKHzdec7iOffVE75Fug
8Z8+1C6DbyjPVmDaDSvXdmfE1y9QDBhmjXYuTUxh3oBz+BNRELLotbyiqlSUS0bCSHMnXW9Nakiq
6IzNkA40iKZdt3hhr8sheKC/7y8OPa076W2Zggbjv6GWABntqyx6o/VoUeEA6r6eIAp3D3h2fPbN
KSs+SGLdGLxd/3KIoItSIb39LYRjiuVIw+lR9Z1zo1aRF6MC7+e6SisQsm/qaTnCUIl+JSygrTLA
BbY4eUjtOkLskfnMdQJghYDHw+oZ0MPvd9UxfhuQQm3fNCI/7R9KOwCrkEKquUZuNrhJ0pcMEzpP
/BfTm3XxXxa1Yc3bQ0QiMRlUsHGqdQuR3Gbhoww3/lbLAvHAbn4D1GStnVk8Z5DgQSe2jfRTSk0b
MHOAglHWqHwnTzf6uGY7yBh6VpjKVCVT5HgZrJVR/XRhudnVfHKVd5Wn3F1Zk2RNre6liv3Lc5F9
gNl6G7KTVztvEhJa6l4Z8bYkJVyGMBfQq0ecXqg2h4MA5FfQaE3tZDTpAx68axuAJ0CXbGssikD+
ip5D9PJK8l28ncQXKUeEE7tRullfL2hYJWGlbadkpTdIUZhvJtjFYhJmmTilxZlrvUs6L7szrQOb
UwGiGCOMA7flJL0Y5FPVn08E01OvE4HwRqe7y3PghmdIoYgePHk0KT5o04wMrhhOrht00n86bZg9
XqqPqgmFArrpNl524uR4NLG2DGX+3g1nJx3P5A1+TAUVEVo+3jblTqKaX5tQVVy700Wxkw1VjJKl
sfDt5ns0MS9kbBGLIG8kqywXz0Hw5F9stT1tLzYaL7BGlTBlxaHN+ce+PQoMFp9RhBqevOPwVltK
5xP8+2+/QiJhu8UUIy/MzRMnmNZaGXmmEf1M7jhR9mGCJVXHSmYd30Y4qnwK4B3fljGyTb/9KPbv
Xt9b8LPH7u+ix1GmOv3OyxpzqDOcw7ZobPulaDv8J+KFjY5txTRZ58/G7OlMx4yQLEFnie/13VRz
bvu3hwTWRUNMGrdAalq6NAeEUgMpgojKtNsGa8AYddoqKcUQzNh7wTSF1Bybd6DF+Es1QtbCnhzp
LC5o3WAtImKarDlieoyWzet8E9JsOkq2Dj5pveH8fp1qdnIzjM5eSSFhLc+vB3cY8MJRv21WL/n7
94YU1CPAWPnYvuyIZ1zWkdtCDj3VZ7r7XfrullXDaS0gM3K1Opksg6eeodp9pmOTRAZPG42VC/XR
tbh9K0QgVUSwMdSES1V5y3eqb0EcqcRME7rEpQhov3iBel8nae7qRs/0jNCIeAYYftzTTuv3mNC6
KMgIZZG880t8vi0FSTOgVahFMvtY20m41uUexThey1XdDuFdBH2rrNk0VgBc7wtsO1I3IqFYFH5S
KcwGu3yo4juNQiZXuPX+mps9u+8SA2/rs1f1ZgR+5xNiVIcRh/AD8MAmGSeRkefEJ6Y9qQotkUc/
CSUxRT3OQ+N6MOcl+h2f2SrR5iHUDLfT5SPz+RPYsNmB+twM4IgoNjPMnEPSHrUEBw0wMBSpyucA
9Rg7cjzBAKslhvjnTZyWDH4riD2nqO+OF9xZeNzuhH86avJjWBZgb8+7XHdcdtpLoIZAxZvEwXYD
B+Mv5tGDiEZJfY72rzKoZCFv8/jLkLk1MV7y/LETUXLvODS8ZVCWE5vYgkOedVwHIxfaiPT96Ver
ADQaAKVadrimPT4rxR63GwRNgwGOB72sF/CjdLnUIMv1tat7Nce1aIWLas9ec+YHDU1jPMwiLSEA
j+7mx0lzKFrY1kINv9uTnA+C5qE3zg/WiB2qMKi2TQvMyrXa+BTPJMbz1a3cMbvVnSB9ErJD7ROL
gcp769bCtdnsqAcHV1ujX6u0PehpfiGe9JfljvCRlWE8QeqTTQrV6Ev/rBObjBda4gQZZ9rXNiI3
Utr5IjZJZ1dwQvILdJmkDGDSNkvNq3XKENvmnZqDIEXhhXVv1WQTGX4sXltKnmU27I0P8M+F/yHF
6QDy1Z6r3n+WdenfUs0EpshshMSbl8CmOPPIBJm9/G476XxUPfKpw0aerrF3bW+tV5/pXYBuOxa6
aRveaqkK/LnQDEen40mnyU8B2Ge2JRbZR1JZYLI9b3jiKYV2ugQPNbDovbJUAw528GRRLkzCoWiG
qykajg27GkGDKg1s5N6CdkBUhi/ZT1hBssyulKG37F3ScDYIY5SzC2QEMAz+TVRrLDov6FmlxfBy
B2nqNWIFoiiWWKROEnppcThdCHmjRgDCUw2rD0u7a8u+T21ridHK1QeFD37BvDrB4W63POuh2Nd5
NVJlTfzm3KW7cKI0aY9aWrwf9hVROsQCgxqkhDZ3IpN7c9dvpp/L3HVLjcfOcNpzattjwv653pUJ
lhkr+KRuVpSrGCuqQhI1CR6IT8Qv2dj+sFMNQLCNW8KK1x9752StqoDiKNQKBhCyXxVdzWzKE9wW
O5cR0ikzB0I4+Z/X1oOCyjX5wIB/12F+WDqiSpCsbIZqpt/YoYDfvK38qwgB5lHjhhJolia21C5Q
s1UI/Zu/xcGtJnAOZavdqyM3yXnoexkFHB6gmNv2CEX8IKSyAHQeXJcVUsXRAqXziMoqG/0h++ZQ
W5gjgRvQgYgrKymsRNwwIqDd4gczCHTEb70vQI5y3SwJXqf+tRcKO7zJq8R9kwKfqCd2GsM1kNsw
4uDa3EB80PQtLExoS40EYWbVJG5x2IimlAHOdqsmkDzc8w3sVxZQpHr8DMLGY3IDo8M3FCmdNGFu
bGFY51iLYmsTDZqim/Sg2uHtuqAIpIEFv2362r1oq1AHZHvLAOLom2r+57Qe2Aqro01iA6TQlho3
SVHrZ35QChAYv+jL9bSmpZVXMZg6ikT3xxx6jAcuc0JNqrljsVntThZie3+vKggbmHl19Z8sGWXG
nGmwoyPYAtBDAI8S9m5gHlfN5mekOMoSjaZ8eGX5jckDhHsC4WFjXfI+UFS0RiffcmKYV2kv/PvX
h3Mz8oewjhHCUlwjmcCakfbZD5WC3Y+KxzKb+oRj1wTwiPPLYUiVI/Ha39GXivMKdgb/yH7onqxM
8PXP9MhYcKrj3LqlHtSi/P8C6zfwclZMroXQlP7h9r7MimPmP/18y78QJvtVZu5+5MySwGfZnd8F
7wSXlGB+RawHn8o5cT9dHYFVqSEH6yp6Hb117cN9Z58kgFOHjlHPJnO4mJOsu45Zq7Q84b70NlVn
eb6Dk/JlVk7HEhyiXgceJ6P4GIw1I1Sdt8rynE1NIk8AejHIact8tbbMDwykentnIhPOULM6nUeE
nF76VsUTFDcU9/v7eJ1mXmw4eNsHK6lVjhIWtj3THdVie56BvBIam+/tPkMdnM4J3Dul/yemzDT6
FF+0U92kh5lE1aPVN5byuuBHZ21Rw/IIEAqiQ6wXo1ZKXa9fQEltmRsgenH613MjLU5Hcn1qJSJt
g0SqeTUPMP5lJFAZMc29bNjsP19Vjfskxbev+elg70EjkuvwiAvqBi41NHEyDlNw4L0aN20Jchd0
783boh+XPVyPtuRP4xC04Dc5LCfqCPUAnyfMISQ3hX6Mflt62Nicg43i2ujwWguE+do2pzzyyqjG
CHqP06sLdgcQRZCgndJOk3Kuj3LUFh4ufgHVkhCw3+0VMviLXBQuzPw21OHOb5+vGh7nGjnHuLub
9K3HJ/AatlzJdUrcuxAFB/wK8WB5i8P8aMlsxjEgWpx8i0sbPbcL30yC3qdpo7S2efhHLhaX46UN
x3rUm71MxGRnkaaTXBRSoofv7ZKc7D2iaLzLMACWdqwKT27E7eWuL6a2FSnuvUrP36lvy4ZABPsR
MMpUxzCXBQHn8V5WKmJQkjRMaYSlsizgDAEC30Zy+iSCNlbADZdSoog62wtk5hxhE3hlSCi0u24D
gT5Xo2SgeVJ9kUEZumefaUAgIGEfylH23DzF78yzDvW9+fQPSSrGgFBr1nV8ME1+Eiv/7InP8Oqz
WbtjUlpD0A2hh718OPLaAmCvr569bvu20ypJRTyIUgIo7yAmivwjUnAvxUxWsdALF/st0BLsQQVz
mY8FJgwr97z0xzILkCfaHEX9k+u2waeuqvzO6efd+1YpnGtUMkE9N5DEDWDwG1APAvlMFapdSi1o
pzDT7fRgbW98/qz+AxBZDtj1FokgHFFRuFZ5iojHBsnggT7Eq5v8uh53JIa1dIxuOvrR0AsLO/d9
7+oJPjQv+fjn+aLl+90Mg9Easut0UFBlkbBTTUIwwKMYn7H95hiB2NDpsPMHTc9RVtkrOdUif1Tc
ZdAQX1/3DL5XUpCJc9njJVV4YvsbNZ1CbqQnsciQlVNwyHpYddQeUBgXsu91hOo94GH640BnZf+Z
nbFiWgJUXmsjHRZolo6XRc9jeusWiSsWmHxb0IjvpSmc6Cp5kSx7JJ7hdWEsSl8fSqfGg1UPpCtq
gqh0hXmg1dHV99RX4ufWqV31GwDZ30Tgz+fP6saGuGLySMmJNUu8At95jX43CrbXHLdY1E/NsP74
MkVhBls8RR+n1nS8c+DwX03Gwemox3dAC34796uUkyAUqUU0QTTnBCWQ6QBO5a8XMzzdm8byCCA2
BJAUzSjwYhdxo3O1/qdAOL2IiOeFDv5un18e3R/uKbptzH6LQH7EJRPzuDsSUKPhFGFTbonyPVJv
Hm70Q76yyXwjCZHiWJZ9fvOz78hDDXpDiVdefS94BwYu2P37E04WXUzIDkvqW7GALBCleVI7vQky
UYsFd+VIXAPtVUc+fkAuwFHXL5NmHgMTkYGVuFdUdsKBUd3A3k2+wCIniT8+2R1HyydoVM1bLGhc
cwoDj0ZHBk5psLVo2ZUrwKDX5f5A3fCQDBx9Kd6vBpc7TWi9/D+63syyQVm8Y1n/oXGmMjwywKI8
iTKRM3/hbQU7Ub3dmYZOUqzlNN9G3is/op1Q8aKQZ5QjP+F8Rs/hDC3ZdW7xPwsg14rqPD9o/IuE
fUnn3/i5nFdWyhfxxPob16vXx6VCHUvhubOPM//NkYvYpojSp8heq/RNQn6MFrlCRkYFzZxqiSck
z1uN6YMgg4ULA9p+DYeG45KCTBs0dpHntC2Zygmh7QxUcQL9KKKPDCFiUAJVEbRtIsCuc+p//eeQ
tzQsTT7Znp8a42E4F2JxyDeBSeukmGMrj3RCikAjL3vrknoFSHVpaAhpvpE/NGiqP/cdyxDWnERS
MyVpMYsfTmtSmf+5zumMQg7IezbR2vuFnbKtFlF205jWf/VtcqwSx5bgKbzzpkhgsmOfH3JsWQ4x
yKcOGLZ29IZse6oMfxOv8uJ3O6M98LZKtZD6ySQmphcrhdKuZDM+AC+nm/jRXZow3hKA+VRexOoD
YLux5bxRXTT7r6Nqw8hy/qjQbrKnhB/nrm7qjwXJz/sWXYe9fMTjOXA146Hwtlxbqv86Ec7LVdFj
RZJcaPmYCRB6ZhyA2l01XDe5J1ynbbXF9XxZJMHiOsTINS7IylofWnBn8vdylDXTNBL9E4V+IIGQ
n548Rb0Vxzwka/exZRtiStHdM/ozR3tRGNYaCg284bss0Utxs78yT3mIidVc36ugzgQs7CVFyeNA
JrBUUcF+fRC/2dTwIPcqrm72wKG375aP0oDczdtEsFmjBI9rIuJxeM88Hle0mPOZyDZkFhhOt1+V
LUTCLhSGm4ni/neM+EI6qrVUJqjFFXf41j2YEsNU1e74pZq+CjX022I9Uts2xCfboyG6LdgK2eGJ
6DSwQmZsMROBmRno+5zF4eQkvTL0o4WC4gPLeW85orWJh1VnE7qQgEzfUCvxt1ShfOkPC2GIlb/m
gEbZJfIuTbPkmrBF4qgv6rOis7Fct/s2aYn/ZtI8sWv7swrQHGHyhNNVVt+iKYI901DgdsVXzc6a
PzqCDPXD8u5XtWPwdwRbxWlig2fQqvRUk8eNgW09zUIAj/9zfIOR337M4poxBNJOWjmjLcnxvWye
1MYmVhNtx9yi4hHgdbweX8O+4g95ko01cfpTuse9cQAQwpufrIndyEW6m46+L6aIqPgQErCAxtDi
H4qtJw0WrBlCbT/FsCaxI56RIfIh0BhUE35+dLt616ipSLjlNSVzkEz4uIkWGD6tA6APh37epFsV
hXKGkKWZzxoAqp+O5HSmfsspnAjeGHtF/50T1yuEYkH7X+Uoz2wSvv0dY25EXBUduu2qj6t/NWOz
ftbttsLaOXpuj2c2htCA7PvZ2b8dcd4i6bfP3KKZMQ2jKBaqJNj3VdLPvXroSCGk3MwyytCQzozX
T+0eiFlyjaG5fCRTk9ycl7ThYcD3a6aTbn3Dx6MsjVU6neczJ079L0OYDjgeCqggo2ZTBZcrx0+q
24T7MIFWBa1O7IgCPc0QvLPqcRAQwIUwx9B5JNPYZ61B2R7BnwxuOfpeM7yKOx5Z0XBKSLmhZixp
X5zK5Rwc9BbHBbZUgoE/yZrMpNI/uPHBH1Z0LqnP4+fXUoW53HeifD6cOe1mtHDCUL7Qhv7mpfiJ
/6oNsNckwRQs5SRO4F6oGuSJkU3JFxVyEs+GPjsdpJ2mgthmYwVr8enVnmBaYs9E9zukHLAQdI6B
FVTPHrOQ9vhMOwV4jSLKaiFQoJ0upGdw/BIbmGTisLZNqwkvMkeUBRZ2a6b7q1NABLrWRWSQtWPF
QaCsbx/Z1fiiPBDjFCHH7+bNgUJOJgMzPo5NEShKJbU3AUPo8Vj2MFMNfymBpw20+egOVoctp3m4
tGg5taIg/VS5OgBucbSdlNZyvEXUmzMew8jUkMmq/H1xz4lH2v8R/Jfkd7Jg9NC5+xI6ufyveIup
l4ZMwttGxs/7QJwr8jUh6eoRRkBGmN6aZnsI5tYvPM6/oExQwhueFqG/yFm2etcocLx9tA9cWjXd
Gl/kLd7HM8cqgwqk9mJUhMjMxp7QrhJGDP5fz+d9wHIhk5UPvFx+R0y4bkn2RXMWKWc0Ytms6jJJ
QK+n6eEiRiCyNwDunKKRj2ZnXv4Ej4GDnT22dOXuJgr/EToaxhh/h/KhIGQfg/lJemHdi7zGEDfE
Fx727l7EIM2SuW306AptaypF3SZIT51sDEYTesAO6ZUO6ZwPnB/SSqrXz6A0GKHyO3vE0HC6H7n1
cNfk9W2SjyTYozQ9U7bt5L8O14g96+7erQ5P0ZZgB7NTceAFo1+05QPa71V9BYUA7SNZow43oKX/
Nlg/fzV8T48/bEHhwZuvmm6D3W39gVi1rdWZvNRSshDtvqzAlV4cYZjjeSmK+xnF8FyWdTzzvRjs
0vz9ZzM7bf+vTg0AomGQhavT+MtEgaUHvSebjq5Fj+CYo+HvN5n1KPUYgV+NlY46hPXlXXDN4/bt
7U6HxuE205kSxeKpFsHwjdNMC0Sm1yUTV56VIgZyFeJqGFbCbBZ7qJLhoBq4CaIJgkBZEHxYsjO6
zXcX4JShkvz/y1msQWattaV1C9NyASGCVdvTnx5kuBsxVXCvAtTyPMiC5JQlZ1zsNAxG6a6SvPgq
6tcwdYmZqDWhT4kwID+QXlFQnLAS0PSroldr/rQ/NM2JTuVKdcjC20mWaQw+LG/i6WcigHf80jej
3Nxy1PcNOOyrsuu0EzPCmIK6tkhjKPUjZD7H6jlwK4hR+hyF9dprmGPPgChzS7pTWP4aqNjblOaV
7sstcUb2AcqHKBwVSIrXamOz4SETSf6z791YjU7o9xiuAblgxWollCXeXXVOwAybgESEWmCDZiRx
1k5bRDtIIwIu/7kMBHKlFBs4qMm2JVi5F64pH2PVajDyMEHGTA8RFKMpPXqwCpYEr6+JAOF25Vms
2Pdda9PRQIDh5MDv70bPJ5ZxOc9XPElu7+GfiNabjZmH2wHvaGsU3tjKHTLgoEY41LpTOhH5/f9X
IDZksMwdaq0of/qJh/fs7p1zl7oxSPPT4lfr3v4cUnO1LT99g47XRlontQkh1elRbDKvfHMmU6q2
L8hmzt7zVy14OjbtQl599LHoP1QnZktBRxzGhx5fmo5OAm+DQJdyKN8UM39P0avUkm6JTh+q5BIN
AS5VSYvfPeMAqWTwgIcMfbBQyt9Rs4iJIIjfpvKUSae7eREYaAi/VuTAtTD4BypJ6Ldquw8/y5a0
FStZojDVT+Gz4lPC30GYK5gylUA8Koc1oxCgFho/amNMwK71mbumUSZUToR75rPbqUDLr/YlJUPc
29fynna0+BrzP6hKmO5N78ydcIJIGPgO3GP0xebqcrGqAxormp4OJVlwKXdGDk5pnzUNf0hGxHX9
p4SAo8Kes6ic1FoBjZlMMWxmJpCDMgjoI7jn8Q9vrWTLb+pDN3jJFlTQ6/xIyEVDt9DKmIVmU3sT
PR29wf68VBv8I6BvH/MFDsUMhB0iDesOE5XX2BgeKyM7jzpq8iSkQx06rdPz6vzTWrdiSN2d/f2i
AvZc1gcgOA4FEAdAz9OJEuCuTByYJ3JqKMI2FnneP69w+rBZlNtn5HEr6m2J/T9VRR9ImdA+LKDH
3IhPqQm4/PhSLX6Gc4ANFudfU4/+FVP3CNIuJRchXZMPciDxGlnHbvzdENsBLFgWBlpvenYfNbPf
9wIcKdmINEG1NOXUIXuvlmGJiiITVrn/hWkUQE2jOxfKA04Bjf+PcJyliFMrC6kshZ0fD31ikKF6
Rh7HbJzD0OtmrLnFBFT8inkARJQOSCtptnvNR0/I4SOmA2+PhqDb+LtGOZG6KuDJkmKWMrzioum0
ivsrJBkzUELlcc8FEwAYW3zAZ9lc/Ci+KzuDE+E6TgeJwPz+wtuecwhoEAE2qPOFIgu7dRNZLaEX
vzVa3mENRsrwjS7ESRdEN3B6HV8x7mjzypj7U0shOqzQ8baqiKWIQOhUV5+wTGKHed6RkzwBP3wQ
tiqdXTlelz7gyRgjiiUk0b27UI34Fz7gYPiSixKaxGXjGmz6T3FFGpJDcKQ3DvMTJxMu2Hlu0Zli
vUJm6a4jozZbAn+WOpP//WEAaKSyzLScAjrhwMWsFqg11c5bUYHrQ07cGR7RWmLVwugDGX0aP/jo
JnI1Lq79KJ7v2f4X5UWDs5jn8eMsaZQJaUwnck84kRltMXAfbRe50FJARgBJX1RvpCwdCod3zegK
U6xaAgpFjRalcGfQ19WQ4wNLUwpfKgcepPKniERH2lOIQ0V/Hp9Dj/VK/hmnBePuGt62y3+npYGF
j3ez8qV3pbSMOQ+W4Fi4HRwZRIw6GI4MO6eX1vu7/2SFVvTnmbcVy4Y/essktvFqcRksMqkxZBkz
WRzBuktBgrj4Ed4ufRZCPh/v0Tx18oxWgaG9Ry/3VFp9le4VSyTShGU6m/+pN7OxDangkdujnFB6
QHBigEwKIL0wuGwzZITqJ5ux+BpM8DK/3GMhl3Q15ovP6ZrzQeSQVwmmiQ3m+8qsfnd30fNuUdST
GV8OdTnwieTHXOd+kmMKPrgjsAwNWf1H916C1pyI+ym/2TsPHMqxcXZix16LJpl/nLD+62toQB2m
0hNo0JexaPdxlFzx1AmnEqY7VD4pKnnOPw1mY5gIFoPytcTWlu9tef3+ud1ElTOxQAhnYA9hHvWn
PUe/PeG76RKKrA+RxDGfxo05j1pp3Agh87HySmxHyoxQ2KRsEaqZzmkFiUJOUce8fF4YvFvgOsh9
zDuSHm2wXkmkiTmt8ban52oykxAoDW1ryJZKa3Ct89s/9e1FCpmqNxf8fbCYh5JFFcasAIXERcPe
ej/F3kLYUg/t7HTGuFZiHDoEbZgveJQFwxbd4dQ3RQbdKL8hI6mVSHBz1nwHQ3DIj2BnsdOBNZX4
iCrTw3SDZlIlSdsgao4L6IT97MEiOPZ1Yk1R+eBq5OXei28i3DqKC0cinJFFJPHHhX2+S47o99ch
u7Gm2K9MmaViv+/RoMTRZTHWnH6A4FdV8Pkhgqav0I79ApLEO+WJAC6E7veBg1umD0y2A1TpqQfW
5/p9yr8Hg+exMeuwTiI/Fdy1Uxy9oofVH0SVH40QF7YGnVzktFK0P5DYtG1WXfkiz90oF+TM3Qkr
cpoV2CUKFEPqefbzpejdIHW+sYXwuPjVo6Sg5xdBVqfVetFXsLvQM4WY/qBB4woHGKHxujUXclBC
Q6dwG/bt4Nc4Dk6CAkFfAIJBCfLk1M7fh1mQqp2cbpE562ahY6223EhWLoFTPT3I3PcoXQkPr4qv
QLBpy4DEIIcInIFoR0g9kWTNDOcospAyFx28656WjfpiFCu00L3JzMRwqnbSwGb50yHL8Ha6aCFA
gzzf121v34yFpNiHnF6u1C2mAAkqXFESeRkNsc+XJksNXlF1yfWZf+DOuGxGnJeFJVmMlAZd76mx
U2m32+fo5W4yqLaTw6rWIkMZXxdq5L0iiODS9pySPg2ulDgRMTF743A2tEHVWKZA6crwGSdOP8fq
ixaSQZMcpx0ltFj6Mt0xqjqXsdatc3aJQB9h8DUKCRyvIQF/z4NhpgRedhR/fNje5w3Lk704tupm
gf/X37xuaeIu+EFyA9ReKY68gW4+ZVNpRozQwAIaaVDgJ1i+mBxva7K8+c9f3TdyXJsPibtCUDBa
E5DrYrRj6/V4bYjDGwzyg2HLj8D3tyJ+M4gpCBETnQlhaGAGFuInVMdPwZJB9xBvkGWxzd2j+pPR
AzY4Ggzaers/72cJXx72oty4UqWXyuAxkX8ituVkwYgmKHZ193RpFIub/icj1ULHqMtzIK53qpd4
Tv/LyDEvV/rPUBQ6jUlgK2AFn3t4VJiUH15U/44GsLu4fqhcGg5sz5LZVs8fruvqPAUUPKy9lkn/
Lvu4hbBCuOIcFqE33mrdO6OKaQQGdBGilogTaEGBkN03BxO4sRyVM0uOdkzT05JLUs4lh3RrCDN2
bzTJG0F9c+QaLUI7Ty/taTLjGArh4LWl6ivJG3KzNXKER7jtKsgC797oA+7F7INR7g+ZSO/QuHzu
nKKFSQ2JaEiPWJ9vFbn1jf5NgErgmAkc/rIgHTrbB7yM/J8gExugyIlxjmXsG59xdEYKhgy+esl6
x2uKbiTiQsNZsR3MlOkIp9kXrWrG5MzAUDvGupmI7hcs4s/GbYclV/UpiXwpr3J5iEaOle+e8kWc
I91Bq7qYC2K4Wdmw6HnFoDFFiSYyD1eT+8SWtQOIMKB7nvI3D8cRYUfETRebtunDLaf6OmqiqarC
VDZZcRE3wAxmrpW3WEo+3eUhxasdOK2RodMrLQrXLXC5Fud/i3TaYVrrw1VXQ3NW/Wat+RXRQHxD
nwhsh4nlvsujExEjl374iciAJOJSdi3qyOd4wA38E+GELOdkUlHQg/xjChX5x6i8wrgNsBNGyA81
me18Hz2yMx8/MllFp7BV84TRTXoioJRKf0gabmQgulUgykHJbQ1jwp0OW3Bf+9P3oBCI7t4lRWbs
4yeN7BtKb8aOjUorkcThgvltvxQ2VVsQtGkhGq89WUNOKsxtvc8TXrYWXdK+r4QfOijhnyofYKG3
GMleXRp9rdzT9/aM/wLqAxU45OPs9eVrQ5hKzLAi0q8PbVSs+Zf4NNxwftygOAJfouxTRYFEtqTR
5/MLC/iuFvwjL4EWNzp2fKHjYU5jJ78nxtQpVNRvhDvXOAn6PXjFaNcnF6UgJcg/Qbadx6oyFpRd
W4veJyJNjKu4ZUNKs+J1YFoHZ+Vm6iLx20EcnmFj2f9ZDAFDC4iehQubVx1Z5KWCvJcOKe4jYT8u
aY7nphBik1wrtPq4xXvY3lNfUSU2bKlUhV2AfqCXCwhPc/8rGwAyxJE/tzZ6rxCrkUDgvCA5Olv1
41YfMaiSeYq9AOKCu2F1p7UZE9Y/H+obYhEDg1YuCWNAMf/YI+5MIuU/TNSn0NLj7zVw4TMGH+0p
UzDoBwNxYgMTeM65AYmCjOO16YcXlofRMa8DCM/yMou+Fubc1QywzXIDuzWKFCdRGTS7TxCcQPtm
TbWr6sPDFqEkTiEsv/LXaBIgxQPAFTs1OneRQhnQieGj59Ww9rwxvDLEB+UQcIZzp1/CM+9ROU60
RQR/UEgLaSJEWRUmiyN8jk9qVZFkdxFJbdxPpBMdCyXpiQYDOYF/v+v3G6NQhJr6HOqREQ+77ybH
sJcoThmG7HNyghI8E22V1VKOYT8ZRutbhi+BqXEO4UYMfF58uUz3DNNlukhvBCRZTqw0ElV+1jRR
KfyJrDAqwWtmsbdr9zbEcTiGb1P3hqdYXKtfZ1sXAfyMW0cLqL8ib8YEukIOjMzOZD91kzK9X9Bw
J88rHr3w9Xayt23JuOo3dlYTAhm4kT2mTWGq4Zp67nRk7Wkm1pg0XDULKMcrud+62fnK+AsNkrWz
t9HfPU3ybt0mDsmUZbzp2y3wPhTdTYsH//nmZMUlnRGZeIUXqRq96/B2cPxfaNLCTjp40FScy2V9
xH2sDLa7R0+8DCkFQ3p3N1Zgrj27iYeuEMZqWEKRFHQ8bBS9lnWKjA1O2/b3VZqH7Fg4S6/zVkue
yz+ir+vqauoHOniY24lyNHKAm3hDf/KmIMptln6ilCBOgrzof54nRHhrBe13lSFVTHamJAjC3Fwk
u9+FJs61xjvmrbxYmt9OQgd16LsoNqYLGjYcQjwHsHmaXI7jj6+dKFFABk0MhgpcHbv2L8qPZe0M
a7ec0CJyxV+2PQa9LxA114L30WBN1jPbG4MdOaAmn6sJaOKzTL+TXKWQNJF77isnWpFxdn/OJ4LL
9Hx+MZh5ryNGCyw6Jlffj7vW8aoaCG3EDyKlZRe08+t1+oBIIvE65MYwgEEzMHqXvPLEnx3wWG4C
ozjfoAj4KE2YR5TyhyrRz0dWY/JGJQFuY6d4WRZpZaM6BfWBVp5K5nXM4OAsfF2+uvAvxiUsr8aF
CMsZ+pVjtY9efJmrUIOgQTeeO2XneXCwCRPceGoukwOa5JQzwMrqgF8sNMtElZADMYdvGNzvftV4
6NExkqTvRGrSzZwkEqUVNopmg86eEaZvwrWi6PM3FHonqYYKywkbjEFDFVQyah5Cpjyi1PfuYost
eEeLDp+sC+aZJ2YUSE27YM7rKvtaSODnzmntqQwPY6+GJ3jv2cMu+9qT2h60heClRI6dCmEc1ez4
kTLIUsUl4j+3FpRCLAJWWIkXvYGrZ0pMH1a4SHYdO4qmlKbiQiLrJhgxfY5VA/TemnsF2miJsVNs
DFG+h20Uuulxl9sqRsq+R2LqyH6+r1IHqZdPoOZvZqP3tHXZ+cWM0CAw0sKMcHPq3Td3jY5HTCHa
z6uHKmc1Hwc2tzNQusFK9hyYZFFMi6oOo9W00Dq3vbHmfBO729FTYxicdyT4lEQUQa13MSwbkE1o
204Wii4SvNJsRRhE9xGrmBbgML5porKyhJXxE7mUQ3lit5yD00nMRYAdtRmYHfDmoYcVHm0FJs6H
DO39m12hwiJ0GTS6rUsdCTM9itqKRm7gx9iB+bpCZVOYBhjZ5IxQ08PZAV9pVMwDqUDRI5fJK+e8
zpFgKW5bTzxMVVxcYyatGyQL27qDA5EShZQ+lOkBWLn/TNTa3nvrdkqf3MZ5nUR/of07gwFQHTUt
UNazA0OjPKv+DZvUk+G4BqwfQ9WzX6zwFa7kvXMhMS2dqS3SXRJUpk8DgO1zq0sSPuaH/6tHwt97
YymfR01nfEJ5OfXYrj/LNKGgidP1yf+bJGWFUyiGup/vhhtcxWFR3DxVrcVraqlo4c+V8p19ixv3
lSaaer6hPU52uePPuhDgFTzoXBcp99f9evay8VG/Tv+LAWGMSDYxopmTK+JmzDlAZ7aVYHrnfVU6
WC8nf0+fjfB53emHvlcxIGYe+S+ea3j3PS1XikKSwlhNHUbOAeNgQNJ53m1mC9NzufICB1vOm9Y1
78gvr4S7/e+RJUssb2eza0DTO2xeCy32emEec1mXAZMNNv5Z1DsRdXCCzMuJ9Bo5N0PDM1CTFIu3
qz1qE4K7GNhSocxOLo5wnjG3wUEVvQuJPFT2d4N195UlcVsxO/Ss3X64YjPiOLTqLE/eReQIK/s0
79ANesuuhXg+jdLPY5IxhK2Ww4ZhVg60jc4TTali8DffIy3EY/M4dtR0tiV9GN3sgy5hoMLUlEn1
biIzm4HROsz8WKFwgErYK7hWleuwBebl62Klz8hJjtolRfD6wNtG+MOWn2wPrpp4Wi/cTj0DgP7L
GjLmG7kX3a6SLxZ08plyB4x4Z0hFo0A/bUeyqbooeRgiordzxfCQybIp9pzOnFiy0lY4k7MMpSBo
jwCM+hSKb48oYHqqRKN0KIqRd6pwxIk6atX0MdTSBcSOqO1ufJaboX5JACfBm/m6aEWgCem0AAEC
08VhoyZKQmH+oonszDME4bh+yg4RU801m79lhpuN5E20ikVd2cxDMlk3MLxMUuZhHRSwftBuZhJ8
Q1TZ3M39fOekskIXGT3qwI7eAgVY7d1HiBYtM36gwvKr2kug6r1WlCXbjw+Gu8a33ubdLkie1Mya
TaZwchWbHWlghbDJ7fA7npsykfWG3shnZNvNLpgPCSK5EzfZlgw1PFJYVLsvm54FNO72r8XMMkXQ
pv1549IlUhpKN4EKHd8VpAkMwnTgYrGJqpw8/WzccPD/X8x0jeRbVp3plXBUd1H0k827Yzj553Bv
QhQkEHigbIHwgIbQSCaDQmDZYE+jEQZu663DWIdVOqDkH2PGDmMEa48H8VomZcKySZlxjMA9pK4V
zpCizhp4Z7kwQiLZ7eppkFIIroXsoIbVAYBoDyiGjkZbmJwLz0h/2lhahguAYrSeNnpnz1YmOd4D
QoK6jDDVskk6MSJM4a7DYVFzRzuWm5FscnZyRn9NBpS+ck8qwBeFrBxoScTrbr1SoeJ89gCBeAV9
6VMU6eqWefe4ghUAxP/Zfhlt20lmDD3l31ax1ftJfFcnCMj17Cb6UDBDCO24DAnF9sIYJNcbBrCk
LZlca2I4rcn+1aU1+/kelibjjVpWDcl6+BUmFAuVUMOnCTWz7UXxQYlcPUTbVasel57UBzCqB0h5
/1KT8qJzpRc5sBhifxWJ61HZBsWGunyEY1WPcO5MioeoNU515Z3tzb3VmxUr2BPIriSmFgSkDo6I
7/THjjIH1yQtkcCgm+XsT841LMxjrnOA2+L4F/NWNHUOOL4+qY8vS1dt5kka+iDQ0xU8o3+jA1E6
n96Foe/5v8+BsMrl1h69CuG+JXkPxh0OUpIIlQ+xPXeDRkcl4ikU97fztioebuzvvS4Cr19hGgbJ
/o0C0giNoFfEvMDcUmzsaFcUXuc+r/9VEy03WzlM1lyVb9X0L6QCGS+7bb+GSMeKBS+jLOmG7srj
ywOa15SHGFRSBH0wbN5AhAiukMNG+2FccytSFFlk5OKr6zA9SvOYGQsEa+n7O7o/+2Lhzu48Y2cK
vPjmdISNeYW7V71gPuVLQ45hSgzUK+/LfJTAOUFfhP6J4pXItwc1qY3mqbWAxNJzQR5ZaQV1aOWS
2ZtKZ/t6gzyg+laFyFNCPFbYJysqWTptyCY3QwW+SQU5q1ym11rYF9NGFmGWqGb2YJco15jPimra
1TBLIpd0T05iS7XgHvpI5hm4DT77IOs5pxjjO6K2HOjsb3fIURcABJ6dT9zb+a+dvrndsWruFqYx
KvK8DT0bmE+P5TXpVn4pKROlPgMn4x1yLVrZnDFuGD1Apfke6ls/wf0+3nIxIij7DnmRwksSrzMl
56qyO4urG6NWb6QEX6JBacnZtUw3A6mxSrMRSg+GD2zOKhd95rriDxDokmr+pue7JHwcTKVkz6AC
YMT/6I4Esbi9Eq8KZXvY+05VW2ypWRF6MYAn6o7v4Ahq7DvyU6tn9t8zc0/pKv+PZBX4XgFyPpLq
XlHXl71CF1/tkrvULuGmbm109mahj6Mf4YTN1IBOCmpjxIrr41SvGMHZkcqn9W9j+/EDuNhVpokF
hnczMaqiviWKw3s1tU6Z5CWRGbT8ruKSsRy43u1JzEGcRQBIGBDTyoj21jN8pAumVAKfvPn4mKd2
rwmp3Q5GGiCUIwJ7scHqKGcrv6BNMpEqihqKuP4CGc87ec4JeAV3VQVv/YAykBhOHcFjhWe2F/YD
ZWK1pXTIV0Ioa+T/oOG4uBO40nM8LSbk/klcUnBUPclL0ImaUHzrR3JVnMteHUXZyucwfk3P4BIJ
XJD6Rg5ZozVGdJ+RUceZeNDIP7sIM5D9OTcQSFk6une39zMfJdozi9h65sBxkhqtfIkMe+fRcRtA
sVbLbOq0KkvDWNElBcX1oOTt2E5cJwr5QvzfhBJaCddxETfSfHqNlvRzAWT4synFnxM1hB2u4rdt
bK2DTug0w91BX3RmsSQLs8l75oZsTebyG2l1dQD6pxDQXsPdAU9f32PcoWKmqiNbEaxZySNbpUgE
/rynfaF0WTxCSh7V3ZsEnAYH7IgtloJlAKtxbVyWz9hF8j8a6ZvQlaD8w2LxrajXKNxKdWM89MB6
KZ4Ga+Z4pn7r7TPp0ulQcL0Q5rD9Lcgpc8xiHZKcS7I5xnx+2bkurkhp7ePLCGHQEzRQmjCDyEZZ
q2wb2uOTop5LIchOMrRvmI1CJ/S6w3GYhl69fuxRKlBzlPVAamc9xW5v8S8USs01CXKN3afg04lH
9S+NPuMyc9dN3rS7uzk91YkmZsu2UqNywiAoy+8eQ99s/6AplVA8HcEN5L3KjNC0jHpAgfzB6VHj
zTvUMxlZxXVuhp7DDuXn/uYSAg+Bg5PYo7Asqih8DXSi8/r9afgvXbLbM0Dda8czNIa5bcY354dm
7kXDQTbA6SRwJ95vBmJggK5zfwMhKPLZ4KUHzj7o8IkSL29Y9pou1fh5S6Tcwh0wk0EnPTm7vNnP
emjUz2bU1lqw4RUCkbtyysS2LhflUUSnxTs3QGV9y8Pvun+c/SDeZhBY59ccWI4Z77g62L/ewp90
vt3n1eXrkbfZYYAAkhMPiwGvJxS/HHlqZpJ3N3orVhlMYvQl3H7LxD51fiamBTnV8AbjbVmI0ewB
EPdqPt0fdKNjzUL3u22jVAy+xMmGk5cpO4n0KIcKZ2/HGPYMDDVhsCryH9sRT7NVZHR5/5sz31W2
fPgwTT4A04rMqPnzimHq7zEgfu3UpgGltPWqNtkqOhhSYPyKiT7OG6m4xhdY4iQsJyDCz0IcVgTa
/bj4PhKuXAV4wfBPIJGDl2eovEr6mIBXocGVgF+3zx2n06NhmekTidG/vSEhjCNDf6ogmAh8lyJR
sTSKuj3E3CSE52I8LH9ZhE64FKPUnWseB8VnfFOMDsLI9em4UucRMvPKptyMpNBFYYR8zkCbqL83
J3OBhcYL8V2XZrOkGblVLHcrtX/rLortt7qyHedn0JQYMovK4KNlAVd9F5NlV4LPsYDS4//dAdMP
ZqD9/7KXbMcgwg3CmWnNoGOOFIi5V31UhuZWRiAJJlS82HSRK/wF83QiJOamFNRez6MLIj4w69n3
rt4qUUMZvkKpQuU8Io5JQ3M7B/wSd+YtxmwI5cZbdU9di5H2sDY5xjh0rRgN5vfmVk+PI8sUr/94
DDD+N2+jQ7MhxzssqC7cGbpaTN07puG5aSjAwa0VcZscwEd9iPS2NoH5juCC+zSZ86nXEKcfx2pN
twgkmSL1dpHBHTyEXG1MEyeoFp+7FSr+4N+6BF6kHHD+NmQWzyTt2ePG89Adgfc2prfvMH1yZinL
o2xSqf0IuqnP61qtWTY11JIHNORkUubWIo8VN8/IS/Wgld9LfXnMMOdb+sRyzMQSrY1nTLVHk6JM
nBgXKti/sDMFzXK/pwHkubw8SVmmY8PNZZN4padRGdl/cYbC4e9GUEX675QVa6FlD5ZXZpSLAoIB
1eZ55CsbrXmCIWMVg1uZ0VSltKoPFPCHAAPDFXxUnIb6teaePrHt1i9uBZSC0JScHnbqno6Wb60D
WlgJAFB7ToRslpzHeCeRvsFj/RmSH4rIVtIfgzyO5UXux+xBxb4P5nDKrTDSD4u4G5nBzf7AE/yr
+EGRxvv7skUA1x0QAIxpPRnGN6vaZuy1WugE25LWlL8p7jKqCUb9dgqnoaJrcwolf6rtQiPFxzOk
A0m8f1AdovRjGCr0ENICWEyHP1tlkaT44sWoh97682a5dR01Y884qY+9LEuFF8cGS2w1Q7U7U1GF
Nsg/GkKHkik/2dg+f5QxTlEj4ws9wCgjtRFhNXz2JbbvblFeh1shphtlji//jVOakUjw3kYZqiuu
RSdnpfwIDm7sphl7bgr+WjXJkzNf3/Mg93G4IUm58oQyuQeR9i0TWHGDoc/eO92qnnPKU7rqiws6
btTdQgNaLFNNDA3O5mFHUVz9pRU18nBp4v6gozFEL+zEIs3Y6h3VFGJ5jlBnDwZQXace0tJG42mv
fVL0Mg2Pm5afxVbdwSGZiQOnLS27mLUpsAgGkj+Tl/Imqh5FtiedoEIE351CVVpbMgVM9JEsO+Ai
/OVcen+v/sMBMaVCY9p0V4NMNpTY9hRiBmMqv27J8RuLH+lB5toSyDQSmk8WgmzAq00ppv5CQQCX
jcNPmyfS8mHIIMcD1L9C6hQrYMTus9dr0ogkCCHN8D5CJq7HkC67pfvlb31+QXhpLty4S1hP/6f/
KnbaQ1XmzWfJl/S+wm/ZcLTyRtWeprXRLLiQpfnTiJ86CEK8X4gZiMkD/11g1Zw7T7ga3kGCdiRe
MEBvkh6eBZBBuKtnoIroRtVyIqytbGKfZmhz/2Q3t/Yla1U7QnPikIUne4F+LkSSJl6/dqn3qR7W
B7OYq0aobK3Bg8bZjat9Ir5wIu1lRdGiuH0ePXHRZ3R05+yHmTfspcda0lMjMhN1WxU9SjP+BI+z
EtN/pnJn1TRiC47ZvijTYetYdujbmrim9frhNceboZ7ug+7t1mSWUANSlsGCBuMGsfk0mr0faTXM
xT5DuckVR18QIlZ6vW8q93NwDXCw0LD8lrqHoRYBs/z56PgDYsYeENlaNSABdch5Mytr1GRln3FL
syRD+UEFQMA3sH09y9OrS0BhHaBhKc0TMiz5GS0m2ldAIAj+r7zIL3BKCi95O1oWhVgrrl/P1NAG
ftucvR8FX52yUDVK00QR6dedxLwE/xptND4cBe2DBKua68bQW/F4hAYBc52WrrDTe0PxXvfTx5ct
y+1PcC+gdCEE0Wp0W6gpKDA2WteH2xFCDeovE+/lji6EFzTKy0bweC0bYuHfTbeHeco/i4WE/9YC
GsDVv4nFxxKBIiyASGGRj8bOBopH12zvW5yvD1OdaYVQAL0732AuCuJfym4s11W0wFVvbK5enqQ2
6y6wcfZWNNNHLrQAYnSxUCghV3UFm5qgTaV6ZN7PsHz3gfTajJFdrrdeDYfN5XYhI+12khoUdyRd
QF9sCAkaCuwaYT5sUB/eexqGO0M2PYx5ZVs4f1ixxoq3xbyFq/KMcoB13YEf9+jQju0sEd3QPHl1
TOBwLMiOnyHLiMchBOcVXwXF2hcdeOBMuoQ7kcjDewswmZeh5IhphYLIzF2IJIj32h+gJpIMuJtb
JCgoFYcvbrICVo78jWRCwbnhgw2Pyi8oMSGPcZyxwJC2zMc0X6quYbe63PYqiuHOLqmkW7j3VPH5
6ppiaLqp3p4p3kxFwcfby67Guj/9mj7WnhOLZ1tuhAruQzF9ZTAj6ovGr/L7AB931Xv/RB0UYow4
7Dp+6t+pzB8dxhDiRkNIMbLbgK4Vk4gYOAKHPDS6zDXbzUPzbFuFi5qnpMI/qBFaOVIlUABzMo1d
KtMpDT2e9vUsetbgvac86ooA8LvgX5ZpPpvcUrns04ZjRWZ+Fgvrz9I2dquiSYEll6a9gyXAngea
qoDwDhXaShOXOSYSXOafJxucJ5J3w66LyeaUWdO+OIP8OScecSE0onHTUxrBj53IPohRcD8+HKcl
T4QoebdXMx7XZXnUM3jTGitpROdB5WIlIEkB2dxIEQoaHAFZbD5T8fpe9aaQvvDFEekgEEcWezrd
j9R4Jp7YwqN6GZbT5+T3wXV2XdkBXkm+692B6tMeQ6ZIOsgATbSBn2Hf0xOSE9zZRr75G1iy/oWd
5Y2gu8UgxJHPlQjAdmfyP4l1LcuOqLAI9QK8b4sBtA2aW176OemYYGm9DhjVwMUQeMhp2LxHrkMP
F/H0b5AFu0dxxIEiBgpb59WWxaKOLU34uxNya96GkFckb+uHT/xQ57XjpnMsEjBzjzPzjzd9Nnc4
4XDF03K4SDjanTh8h77EwHY8AX26u+pK7lpx04lxbmV/iVlciBC92Bol9R+XbhwbJ0K0dByaWrDO
M0kfom8ESz2sujAPldfacdCfuvkBlUlJnnca2nZwSBlHROSKTVQLTlWBN4wW3hEFo+o4XY2J/c+j
tuOB5UrtRXRUhU/a8ITbDBizqc+YOolnZ8MCGLaoKHpxbi4Uv4D2D1toC9cPsUgORSKjpKCUeYWd
YzEJFjNZHbNlNzU3ynBtAUyhZTBOwd+GpoOkhurt2KHRImGUvbrksFZI+Q8rLQgVJQSWyLllKo2Y
P1pkhMehNrDJlW5R8KskHD2Kaj/DENcG0PelZ4Pyh+7DgUJ42xgpGGeW0f1CWC0hazTZ7HpUbRFl
DAtnko0Ha5CgQf7ELLbAVHvW4gVgAOIzs5Y/Yj7qL7tZkP80p+3iBFOEXO8FlStHUXltmTNfvLg/
/zN8BmwH9pGkkRcoyT+BhS3Kx+v48tRxwZIAAeYK8tzKt13rt2KO3rkvTYS/38S2SkNW6gjB8oXW
tVfQzCLvs1suYESSPUaiYwjPJgMjbZsnVAFSj+3/yQD9jImLnzJYFqMtabFsevYvinHL6HktlOcQ
n4J8m74KBrwq1Dh58ZFyVuKBtEB/co6NruVgftuOpAZdgZbtiNeAMRCrjv/f//4d5SncK6rBZgvd
9CjPXHFyYV/2GkX2aq5PmDJVSH9QqojeAqLRjoCB7squisdCbG6apvQyPyTlGjQa4R5E6Bl816BV
GFCh5yMHDFJ7LVyChx9cSDliCrnK4hTRKjR2NPq6eXjDgP2EYGa63M5q6KhDnkPlb0LtZcFPQke4
IIIvFhcSaLy90VrdsfFB/RfVIMtl9cVY0LaG86itkGTwb2OvbQPDD5DHo1GePlgEFpucCn29Ntp6
uAJWVfJVKe1TiNzFl3O5AecQDw2UnK9vVms2AFMc+dPv/K+sfbIzCYgtI0TQpkYdY7tzaiH5f4ru
LYqyP6UlMriBq4KYYgS1douAkdg2fIGlwm7YO+6BqXvHBBHA2pGzQGaNXRnBzBEYrUTfD8IX6nR8
y3uVGWTQOvWtHYmd0hH32PvADtDdzvQ5hEqx8TYX/GdAYtlrjVeI+9rIukmk8ka9+b8pZ+wsv3Gk
GeQ6PIGVJ2pnF8Emh0GXt6D1W2qsMpVo9pwNYuC0s74kpAOfCumy+vTLjJl0XQfqoO4aGWzdQZ+R
WJNY03Eb8LK32NWVL3BEKhk2/eNKq1JZgC3tG49j5Xk/fw5AOZs1zwflcrczyfEywdwQz2uzF1no
3s8U8Eeqh45sUmoPhh0E3T4UgJslTXfnGvA1QkqAKixNt87JmNwdwTvdgSQt+pkQ4NOq6XstZhyH
LJ52BbOoPCZqnUjVzlqZfi7CQTnIaWw67GysUbAN2Wr/6ozSlAPPnwtuWh3wCIswMy0TT35F9ui1
P3QhRuEAxOIqzVCCWeQsczRm3BfRTNDCImOz2wXdPHEsHMwHQwA6mO1rqBNbkXQPkUZUn9aKNbiD
BHR3rSunfp0zseaLnIpRGZkFNK+kfXOqsratNvXjSGnAQUhWvkp4yvI6V48sjNgbjGrYMx9HgDTA
SlECDQzlv63gRykCaqwXVa6qifg1hWP3M/icQscjfU1OI56gn4lvqik2fBnBNarKTWYyjs0sl2aZ
Mpq6EWWN0N4Q+eakgWJAzqidkYRtvzBnWkbRX1KAHKtysJIZjowIdCxPNgUdCmHZxn8UcGgbXgxH
gSbefNrXH7eyqs+S9p5MlF3zO6CnpG4ev7hHK6QNGjjY2AGeisr2aL6+SlVTQ0mkjfHIXW5qJmc5
hXEzEhCZFXqnGaAK5lMfj2NYBaMw9T2T1WBdje8ODxxsPXTdGn7GGkC2mfwv9v7OWqVhFwltVH6b
NIGBWTYuaNKkOx3FKig1WkAxkLgqNxocVv/Kt1BL/sFINAHhnLVPfVbJNtbXwSTIJR++UGLEDXfQ
iYekerpB3Xu5JQR/8oL1ZJxC5FmYJ5v9qH+qsHRXYXcNqY7FG16QQYDJoLTjYUA7yhScjz53N1Fi
fwtukNeUbx5WjHoNQqAmaMWchagGU/cMRSzX5DCHg03dbHJXJbiUatwPM3TUHxGLOxH86jhG3ZpZ
lcCpOxaBf0SJQf3dbsmVWkrMuT2WdN3Y/iWvcP95S6z2r6RZmdWw2A9t00babgsRNw11tK2y3bKY
FaIzwqMpNrMxDjed0FynRQtvm9KQp6VePoCrO67IZwfrCSKzZhBCNkrWSDIQUX76FQb9lnDTHAa7
c/64433Tos7mWeiQo36MNL9anO2vSod3p+SlqDMmqDeIQe+uGpE0L7Md/hOZ8O2hkLjqBdssGPq2
EurEpKUrDRa9qW2EzVKk7mTz/ku2JDGTkqv0YVt7j++fPmnjiXwDnul8u7gt4ux4Soc8gkQr1zSd
b9USvX7BXEUSELTc2yzBsIrunyviTaZ7eB3Ug+rP7XqBEEi15l8cdgfhGrcdFhTJSmcAP/vxr/aP
xXOvaq4GEKUgNmEP5bsQ56EqmosirkMV/+mIp/9Bx6tPjrM3/VCCnZdAzwXevPzfSlTehixAF0SS
fCL175m78g3CsoSMJi7PpHqsOCGrQ8WHSLXi1G5Sz9EWtUa1cFqcOw3BQpwYErJ9WpDDBHFgpjdY
z2I7nWJ4HG/0xCLnqTP8FNTzB49rsqWTk/n8hZgZao2KedHqtLnluD27ZJBgmbX7AsRqFzetPaoP
IUeYok4aIWtry42M6vsJOHQkzc/Ic27xFD/EI0Fo/trVyvKcRn/TSthYqa+Kqj0oWvMA2vS4fAd1
YPJhViC0z4ocZ4/cevW6nqEgzjUl5pR5lEs4uNodr/SgGG/Y9Kbob5YXYJ480I4BiyP2ZrIEJahv
l9lUjFysHAV27x+AiLgwFmfr8ceuyW/klo3zvfMnQRoFMiK1m77RL8ycwJPNOE6OxP8FrFf7vAHo
yD2p9HGHtnMBZk4NRqoZW4rWJbsU3tv1MGUa5RNUPPOFCD6RtJ/3TcThxX5qj9PNgv5yjDkfLhlU
D2SXaNTSg82A4cRiiaNdz2pJOgHIDPyAj162oat72wH/8ZFCtLpaMCymj3dTMkgPVj0Kghu+nGNL
Dl5p8RmPbjRVzf5z1DZreNXUXw+LH8DUOiV8PeNRwBx2TPxeq38lAke3NLgLPb6mCuNr89RQDoBe
HX3z1M4JF7BZoNUjANi3WrMdG1ayXcKN/6z2VeI5VdLW8ZDFVnMRvZDtVfeLJLOGH1MTvGqjE6qi
Kx5eE09IpYBYVAZb4MVpYXvZBgC1vCLxDp/gTtaXa2dZOH1Z4AXSOk1CD6qLGbA4ey/lCmXvnIrT
Mtmmd6PkRjnL4Rd92DNVP9xdDLhNgvc5H0NGoQr9+ClzDh990l7md3RTa++TOO48bADBE1wk3ASo
sp4gqW8cDY+G4eHMy9hyAaxMxUs5RJGTPUsIE653FHVV6T3Tgt/lC3N2XGkIKW2kVAww1t5FMiF/
HPna87D2Vw0Y8xzTpIfdQOIRVTf7x+f6pgnhoXdJ8KPIi8/1zBnBR924+xGYHe5a0QTL3Z1Dh1j1
ohJrW+kr6CTwBDnwZt0pfxD75VoRHnItF0j3sDKp7cZvJ4scasgbpmv6rIqM9IHuT99k5aIzkQ97
+4u9B4d4zwHtMBqqBeMfm+eMPzLCqqIGSnEMFf9CU3RvZcXjQ18e9fg3o9anUjRSFEY82ezw3+/M
tRKZTM1L8DN3VQ0a0oP9HF+HbpLvb6jE7hukyO/wotFGzUmjuR4YoYnXCPcHVaM+ectkt7Xb03f9
y+IKu//WRN516K6QT5K+/TmDn5tfMhGnKSfqH61kw2Pu7hSrJlORNwuBViIIHIQK9kYuiAuiJDKa
b4k9YPRBaAReO2684DKScx+iK7ntWOACeyXE/+T9sp/H1dZvcLbEeepE4mXKzKfVkE4cvK4Im5Tm
LXLkbtN9js0Kbor9aZXr8KRO/kZj+z4E/90V0eQjPAqGjTC2bRBXRtX4gwDJfU1n6tYim5r/WrvL
kx/llq9MFaKlMqVHXmDHZrUb7rG8k/+t6jAwkk79xCaNuELEAQoJyE293OqIBzZIDDTmJlQYDeOc
oTAlUE36MgtreKrvXVKG1WFEKUgY/SLSWZ68KDl1jjsh7t2W7LBkuCVjZJcDlM+Ynwv02aCnZED2
LASH5JIuUUKWU6+ek7+NaOiRKzWWLBdV/SoIc/KnRqkcRIaysYpSUqvTBmUBIuV2EJgyoLNGfrtl
GSXJCwLTOpADR02eaWIO3KWo+yVCCHXqh/L+e2nCWI7Enp04vVuPAhddPP0YaNMLxHf1iea9+IAY
E8GgrDXHPQBraBRRvT8vpATsx4YFfoI2qQIHTus9Jv7DPV6MXdD+n7XWTyfQmxKIFLsU/XFeq9br
ZUJ+riwyPtG5yohmpfqdEVcZxB7y2rmxk11kJyTlllCc3hf6kXt7qgMIp3CmNwBZBx9JmENGXLr1
ykRNLf9dbiGHeJzGfXgNOBaiL9xM5iMabM3v2IouC0WiORyYGemx4YO+6RmslNOzrO/b9oPfsivs
6jllnE/onnvSfBRPd1b8VRwuqPrGt998EIIhopVGdBxNjzvzKiQJUlValNrAgQH+AIDn4+RAY2CR
HUfyn4+oXmwIeZzuE2ZiXytr7uidwJxmj3R4y5ulV8aAAAAC8EwMUEEvokopuSUcq1EEtq8zHHSx
WkkDpP99P3/8g+ru5b1xxFAi7boDw4+bt7Iy05lA7C/jGRmOUAv7EGbSkzKGrvnsauzH0mYO2HlP
3sKvsKoCQA8D6SDulFRUQfx/83+h6rdUgfPDV7YQo+/rrTfKV1wqG3KzYim63lCc821anSm5Ywxx
chwl1l7TXs5VwOvnh/PWeNWYH2MPqDYPoAs1o6sAHAbBtkavOhxCF/37njp7H8xfRPBpbw0kkZcK
bnEDCyh9JzK9aCmzDmQQNFBuDWfG+NruOVnNah4OIcYdnqU2RVOv+Q6yRLaq76VaB5AeLniJOTzm
XBo7PQ/co7WBIaz48YyuymD9Jgbv/EEna7F4Il1C3Qc188gjFxkpDyVSkvUKlCrOf2k1apiIhZUe
KF4okAwbbN5LIrwbTcuj+grK1BM+9VIlwLpH05vq3CopuRyv228cRLhdJ+6XLd9tsrSUByFBs+35
RMCxNeehtjhyfltzXK5k6ZAEC1y0RvO2qX33Wfc/RwwjJ89w2osdPgWs200zraXLCmUSa96on29Q
q9lIA5b3DgMm+nR+RmCFrpCu+IruAgOoJzfRkYLwxFMwkvJzwyZOJLfB/LVRBdStx3AVrm4+lXMW
m9U4HSWwOdz9OQJG8I1UIxCgUhluLxIE3REeicifZWfPZ3YqIo27/IZUOZcGUWHhZ/8g0yHCbqzR
1pdAt0sZ1rcIYVevS8dephP7h7rEXmolpjYhQXK/bj4EOmPovZQeScsP5OmRRQDv8+nLV1Ubbf0S
kROiA4eRE9gdI20JRZbkSZNaWfEDzRIUoHRAmNVC7538geQHjLVGtYt5MHTKxnmMlSw8dvfGmuyY
x11e/lPAVT/uY5AyhEewRoCND/oNLnszDJDnQ7Eu2NkEN0XBqKo4tW8X1OECrRaVbKz5IxTE3PLa
kE/sChQQN1JgQsYUpWg/adxhtxMcB7tdyyt74l3AVVs0zdbFCZyvtQJ/MbyyyGE7GYhdrE9piD40
0JkQmpWz1qoJ04yTZD1Io1ASE7+Mzx5LuSuyuQ7gLRa1ZhJ6LC0C+rpsC7hzygWf4iSx8IBi0b49
n7hLF+pzaoO4gubj+1mdKB64BF7x05+Zrh7ecCJKpQ3x6tELgeREGUM6fOl+MoWuSQ/J9mn3TPHj
v0muWnG6O6izzNupkJM5NyhMQHCcOan2Orh13xPoPoGUTkoehYxfQorGCE4w8Q96v0hDja4vBLnb
GAZnQQr+Gz57koaHE4gyia4oxwh8g9vzvEygNVyvfWhP9KTjMWEvgsuOJz7nbNjEpWFrb+BrC5Hw
SZUe5IL3sr0Rjxjx7NKRTkz0biZvLjg2a3I3TCtKZf+h9orzxlUud4uMWefzVZrbj2W/DRyUy06p
xxD19xkEziZgeTCra6oVp3Ulnm5BG3AVdg0OE0VF0Teep7x2IHD8BVb0khBqEDRK40eadwMNV24l
76Xv0P6WMNM48Jh4rEO/9bFjPT52Bfnm7hW/wBtheYOqgo8viksuXxEF0m8PWLw1iD7YaLnf7bQO
ewdqNsKka/QuivrrSvXUR3mS5aT0elG/dHTI/BAr4iXCaI6kWpxoeKVNFplP/vWcLVN9Zp+645v4
twKlEsCM+mJWalHmh2qKEofkvhV6MmS0dYovlsw57IpOYKDip+Bbe73oSQ/sKq7pCO536nJy/+8d
uiFG9quP/kmKkdfqvsoWkEGOHl1gwAGBydvvExODEWoD30Iz+sV+lPWgv/A2fGN8kDXj7hbj71vE
NJqUeOfbry/yLbG/vJxvX6onb95TG4IfM882O8ED30IM75a8f5xdmqNkHU3KQelD3JHDIdbq+o2x
6+wSG7Zfv6dW7NoODHg7fNU9oXpyeTEdYP5vvEWDYqm8htkhq+S197xlP+FlhuSwz6+qqRNuuEe7
AOz7wJPH7IX0JYH6xSHZTWJqBrta/Qkrm43kVjiGRbybrXzij/m/nzyhB6j0iYVKitO6mWAvn5jX
lJ38jQgtB4Ie82ns1UHvjwJMIztltG0o6k6CD+SHtTqM966qCcUBHNWTYUl8xIvE3lDpa1AYGYDf
RH0C86ppzYoQjChSt5rzRiOlnNMMHatr+x+Gk5QpJVLdmDaK5uIaWkFDJP1Tr8dRj9L343cFY6fg
/ugs/lLCBxXRrHafePkpF6Pv7kjEPNjW3TM6D4zOjUk2rUD4y/9CGojFTVScMJXV7M1+5AXGtPtP
eenqcsng9gqNkbbCcrV4HtUwdvljGLqYMpS9IAKgUK8GmBnGj4fagiKPadpzfhBM+TUMlBPrzs1F
FKckUL/5HdJZB+JAP2FauQO0UznLC7/nICt62SqncvKovcrXCIWB47N6k8PGbn7zuGOxrZoObByd
aB+uaH3QuvJ8I8radKOpmFxc2A853Ff1MLnQ4e0Sxo+0kC/sf+DuDLbivjq1iZkTHuvmWj66el4F
PVVmSi4EC9522IkcHqv1ZU+QhBJEIJZCcmma9/0iizyEt45tZqT/kMB63ftqIH8jJ1+Ew/z87VLA
UfhAcSM+EvT54an0roP+IJAxx5h8g1jqMW9/AhlBZhSOmwxhhgm7LNi5C8r23V78NHg3O1bf3N/A
QKyaci0UwXu1l5N4OZpy5sO+Cnok6J/k6yRq57Q4f3C6TM2XcnnT1AiZtf4rTFYwfpp6xm9HQ8yt
rkZVUGXhnUq9Jq5TdLIyD4j8+5ZualbGbEMlmcNSZ9N913OE20s3l9nE0p/oikmzJifiYzftZc2h
ORmEGAXV0U8No33mRiqoJlMIMM58eChRnX9ONk+aVoCD94alAY4Jk2J2IfoPQbpGv43vnspqeqeq
zAgdoFirBIXn66eCBy/ml5EG6SLB4b5v4eSnyiqqFnBvyVFq9VF6XMm99rFfIS7D577JnB5iZwwA
WdDZKXrGG1PTfdVkCS8lNN1Kd/oYpWftqCVjA7ABgLOFNooXBDYM/L7m6zTSMokAkRmORS6uwv7u
uZ6vxfza8vrQ+sLBROqD0zIhv6recbTmMOTJDsJzuO1iv6J8Wb5kMysjj4a5YwJswxyLFhZE4woJ
bvrORprNlnHBSTIf7yLwl3at/dI+C8MQ7QkAizlNBEEU+leFMB/fhCy+SOKvLtMY0R00XF8PsMvx
bISzVR/92gLYfuf2vubUbfCUa7zW2x/p1z9Pd/PKaHcR+Yl0jhq47PYYvKaqaYEP4KUGKEap+22E
Mm2LU4oCxYNYAXBBWTLt3J9QPnOPTWfbt7POVWG0XI6i9WPXwnfjkmiZdZa1tumNgdJZaBZe8eDf
bv4IdwiCLr7ooA6KqFz6Cca898ezTzBZ5e6oIllABe257404D4NLlNvQAbpJ11+9AvZru9rh0IYL
ivPMGg1XxSFAe2E3n8TmkMxoXQkBaU3DK9evLl0NYoKeXADY13GY6Qq58EqOUg6HAFNAGVOU0CLz
bHXKNZ0YcDeZi3twxChd1auKJwnQ9mfkr5dfhYCaTdmP7fWdVUC/0FA1VsubzL/IfB6cFvVNhxuA
ZPMVoD28x/gEpHRc0oz3vbFp9FPrLfwH6gcXI9dNqqWp9UNCmt0wJOg/vq/9DOCAPMFn1XKdmwFp
nc7Si4ywlURdteXUgLZG7maHN034yP0uWhzTZ3P6lazHG1G3kERcz6NF1OuyBM1mbWy2tygzf159
k5zQFViTCczPjTq1iXfDnDnjZ6+S+4zMFsN4zXgZuGPR7LtA4UJzk+20TtpFbCQToF5dBZH2KETH
anpMC/8VEanlnWiTD7dqISEa8dxYtPL6CgPsT8CTxSYlRRlpRyqMdcAj0eLRwVB93dnH7y512Bf5
ckrIjDdjAkBflnV0kAp+EODTKF8mg8yQ/1q59Zi+AZ7xgvGC73gveYW3/ca1+Nk9XHszdv2/0VI4
ArLJPSDhnFHgaME811Xt6a3YtTU9zC/nwYOeAz8/AaDBMfiIDYXnErzc6Gd1pnVCzXNmPyVOb+2u
o5xmLlOP/b1TWLwvqDeGmS996szVgexVggkYH4i5Kg2/XqICRfWx7R+sHNO1ZlfegNT5RA0N5LRS
EIWHsWiL9NEKeA4FuB9V9l+q4c5b8WcFtWoggw9L0EgFFaDkURl+xm2joZL8bi89nyvZaDv5fAp1
uT6A0WtcWMmEIGGdX7HO7MRFNrC3EDrs0KSsEmrhduQUjTXi0ZUrXIHYArOKSfSq3Eyuo2K80e0Z
Jnti8cCqkPdWaqYg1KHitRlMvBcp3+XvrK88kaojIFod3qFP8+VqtNsIYgif4Mb5QFPf9J6ssmXz
vxvLJoONUmb6dkdRGHvTLP5vnnZrf7etjWjC62WTv7iMc1EKjBY9d93oHvCp/6YmblihuyOaobR2
BrV/JCiCct2RHNLCH0AvIgzo/zb5M89VtijTRcNmgzkhe5uYnL+IptoG1pSIKdRXizp8I/drF24P
WhAqtQ0C6Rqe6W/FTynrRvCtVohTx2XyjrP8IqQo/PWSIAyhSh/Nkc9e90aHpEPJBCXMVKy/lWkc
F/yubV4rqp/xoPdyqCb5PmNYF22ZD4x4YbFbsMfHwnRWdHuMFSR6d1hrDXSomYdLrn0osD+GrloL
ItUro6UkWPrGD6iEXJ/oh2ooHHAxAzd8tTa6zX2iY+SDqzjpr5t6lDgaXg/WeLYHo2KT6lz8iHWC
kOsGP4vjhjHnF3wsRU8wDoSE5N5aXORrMtxtJEdVS4bSvDa+IQlNwbzn0s3pJxnbClG3nAHqGvsz
qSZ7qkHMBe1KAoSILmCsM5f8GRyfG66UytHjSWq1Lh6k9YTa4PXaxAedCh5L61tH+e8nlghscMD1
F8UM4VXWHwFgy66L+76NIAUeP9bGgO1Ph2KibVjHlhAyJyDytlJ+hyCSgtVq0n33ehEfkW4GMQoX
xq1cvhCF5T+sh4AdJUP9hVwzYyL38273Sb2ddL3Oks7GsKJsuQ9RtIJCNAbOgSZucIstAYeJI2vg
x1KELo6wzwMVU2xbCkPQ6UB+kHiTXr7l6mUOOxUdWXf24nJ4cb3RdePRZRBRDUY4oFYKMPv9XD1e
4a4/Smb/nGagyVc97mHrlNDDJtEYHC57Zj7/Ame/Ab5I8YXDOPfJTQnLF5EvafhztHYvvSFuFXAe
TZ/2rku0pO6j7vqtUootikDsvIZFKXkdLu64PbT/yeuZa3NmZyKa7RGeYahniwIqBUMWvO9GOuOY
GuBxgKDzKbJrTNwhPZEBP3W6MmvuXQzXVF70EU3i7zfhJ+kE2E8zy1chCLBYhX+yI4z7did83kmc
n+olnoPA2+vBe9UVNLjUnG5iX8zpI0dXnKPnRrDsPFfO/Kp2bbebDudE/bj08THtjeJhZHil8QyD
aVDKpS4mKkrc5SUXmOHmWjkd67ILOxxd5VLVAgtSIjNEeaYhILJcRgNwN4BVvLm4XFSic5JCQUmW
s5LfAmaedoHUo7qFkILZTXWaZDkDINcr/gog3xFI0i1Nf2pPBjC5xdz1FMaod2eWQWeD3gATIQbH
vUcSgykjQiLfl+cy1eUGI7Ccin+rHwY+gq75b/fseXd75WrwIl122bX57iwVQ+Y5wgceF4ZtymC2
Llq8dbkIJfWgQYQZNM9OnmeKXsXo8bd8F4q81GqFzKL71AW3j00XRmVBy+rQW/Db0Uicwgd22vjb
RW9vAclJiri2b3BGJyVk4E5kotUPdPXYubcMbroBsQgwKoCteZQuvQl2/XKPegv7SGnnasNVdBA1
Cx9Rkf7n8tFt11GeABjDgHNjNfzegkUOtzy/kK89L0vLJbAad7mhsFtesCvLMj10JeNQhe4838to
iT1dz9vwEN3vuHe+laacEjjMJ/0Qlw/G+pMsKRLyz5qlE1ZaGcOdhZzvcEbue7aLtdurjLrh8tdM
/s7sudWKT08BzAQwfogJhNI6eR0ERhU8AXsQ2J6KBpvFCDFeZtbAj3ZC7oKPJ/5+SgWasefs7bE1
ppBGi4d3SEHguZ7GU3YCqSTZ9guuhNf4Qo1oaj10nQ5xZkaRGSGMrMwwQkNgJXlVHPer7+Mujq1y
heVvhVKaUjK+FuaNXdQ2HK4QnQIejWKwQZVcUuvX7QMPbCaD4/pD3rNNU7wTFSU0VX5wc6CHez8L
dXFRqZ+dQpSUnMtUxCOBL4aHF4AszHh+U4xs+BQro+NkKWCa+zQJkY8kJb8uHpPn6/Rm9FMSdgQl
l588xMgOoz8AY/4NHFQLEPOnwhJzY6XBX2hq6VPippvnfU1hmvSdT5qD3dt5X5e1gr7FUjIh9FwK
LQI7o43kIadBbICwY9KEvsLkLtvGMBmi89rfdNq0sT5Oq5oOe70rf704/a3wZT6rimXvAQg1wUtX
14ghnYNYpc4a33LXVsPFGftpKjeU1DjwsXc5ALBmUHlgP+5C6YM+1qJzwsuIup4scOQe4bQTVQ+L
xeYHlHi+9yGaNA7HzhYXrS+F3Dcj/XmcLNpmCXNIyG3SUex6fyKlAgPzDcYmA64m6GZkZhbHg212
ln5P1iXMyk6Q05oYu4bvDR0Dm8SitUy2Z7FmCLF6hVOu5fGOHeT/jjCWhHLtnqbOxqhGma6FiLaw
VvpwJtAO0BFm9okyICDupWKhWr5hfDXPMNXAuzLsp7r0q/tXS080UO6uqoy/7rQYbS4Ik5qpXpkq
mvnMdTE7GpOXnnrkMqG6U6gLyf8c+6Yndph1v1Ez2WScWDQjQljgmRBe6jueBKhQs1qOqA+lOZL3
A+UrV/lqf4PVtgItSOu6nUOwTEJmASMbxTMolb6p8oos1U1xisvrKqKUzLjGSaFArv5X2lBKtQJ+
W7n980KGc9+P0N4UBfaRDbfAnfkIhczxQMXaBcr+hdTpzEVFqPMEb5XZmAv5Wb1fuMpxlMlWVAGp
V0D5mZAnb2IEIcIDU7+b5MtrE97WJa7xHZm6mhVk8WYOkQKr/2BM/0BN2C5Qqx/m521wZkSoGFfC
iU5mAMuEj6C6Rpb+VI9O6xSDIqBrvOeWZryouzi3Eb+XITGMBXwSNSSGFM2rew1UHnzK3Q6oIgrC
oiui8ZjDhBt+qwA80YcB6aXmeMkFe7FnNkJaP8e9WZqn00x5gU9sELgrgaN9Ridz2C22k/iuzYXm
qlUtNqqb5wJPXz9i04hL4jKM3qPvcwivxXnYWKx2Zx41MSqxTZFEfKOWPVjvLLhq/pvkc9q03StA
pryYGylfTSfSsXhrUhd8oSjwUdmfRQ1jeoHP2eVGM0gPL6bgjtmzZxunR7g1ui7zq/xeBcF+KITW
LGCfUujOSMSnHY7s7Ivl3VVq7V9CJuwoI4+HNCofZpU2HF50swUzQK3x6w/9gY1LTrW4gPjyX5p/
q17VGT3zDttMEH0hukycwLzRKBwq++DRSU1UmeHvOlM8OPU1l4wjB+eddaWXLS1x5VALFiDojciY
kot7pwOsjaJSsNU/t4V8Y47FHwHM+5e3/rXBz0raUNL2PHXorxJbqtwTmXYhEMlyFZi1qEALfgCg
wCaIUyodgZnWFcSuQ75cMm0dH9FLE8UiCczq+rEnuoDpMOdIXFTDCTAsWjbdO3otzDSV5h9pARka
tsgeHOY+eb57JuRoV0EsibD0RqPNQJXF6s0nvcIuwKU9C9qOJQXVzlBjtiVQDfujV4buCnQbNSKi
Q9p8ddwh6n0rUwTU5/9ZzLYaAIXEUOue1b819pdJqgslUFgEKSuM2zIFwRpjtx3isSLwSIrLK0tr
m+FOtVShBrxigV/94n0Nuko8kpEgUvjf/reQxIo0GSKTHWr7qQ14BRXO9j8r+7DEPKMlB8egGa4H
CfDDY8tm8kAb2HT/0ZkMkCM+WsKvId9sQ3UiuK7LJUQ7/dexs5guEMwYZeXgLhAq2uqp7eCmx+Rr
96zsOPbF5foKaJjKc2t2+Q2v5+rHb56uOZ4ea6CeMa8CtR11vCc8o9wYQT7Mla3Qi3BRq8CIHOf6
Gh5Mi5EYHIjWd2XGBCpguxdd9uN7hDxUNHBR/v0zBRR8rTh7E4VF4lwt8S4M1Td/5wSe+vh8pql4
h0jWgRko6uWNn3BrannlhYwAXGj7NtWqsgwbb6hIVRoTL9a8Fv4Tol39UKP+ZbI7SBlDwOPBzCgG
V7EetTaNm+mARCX0bnpDV6n9EphlFrnycm2VFP63erXKP6nMUAfi0Ss8n4zj7Psjq6lD2P5kjcLD
ncauk/UMH+TH+LL9j75rMcdxlY7P3MgFuidMWzEqgaRGHHoqt8m16qKcM+BZ0PKPFm4yB3rLxHjD
tdeHFZzKFTSPdYXkR+cUJNY2LodpeJ88CC+sLj5GuWmcxGuaXqHix18hIqFjr1kWuErHvP1anLYo
PcSOGQFH3UVSKWUbNZUHAYN24RQoxNW9tU4kD+Kiqj57BvMOhNoRNChETtE11kxnmT51TL8H4Tjx
z4a8iIfeM2xwmh9YsE6ZH0iYmGAhrgDRFGnKBSDByLH6MJ9YMM4tTyEf2ouYyxW5rsfGy3klgF+S
iJq2AUeNhBc+AsFxKJsLwAhImfj2cj+xFJZFO7shrPHgotHoqQ1gX6Vpd7cTcyyBQBs6kDAdfsV7
AL6mPg5CRFFcZgadtYDpesyRCrIGdPcHWKkSBZ81cTc5mN+f5Mgzck8Pz5lrqL9q8y8mBixW/mXv
V91iMOt/5lBSbEP94PPryB2/TId5d0Q9dw7W5TuilzyNO7mZpxWJ9Hgmobjp95anGq8JLS/uchKi
soODtVqL4H+VreKtVHRslfDWygeSASQ3trPKhxYKGI06+pNPzK7EDw4LhEkN7q/UyI3Bkxe1jUwt
9SSSzAWXjTKvY3QPS5KU6+1HKgjIlCWUeBLvlXK3EghTSDhcGi3y7baH6VoZGLv4P9q3a3/b0Cw5
YzUbRhjwJpt10Q1c0HysQ/xVWEwoasAMgAdKz4dPEDpiL++syd9p0AB6cVIZllLI9vjOt4dbA6rU
aAUKRTf8vJlLJ4VQ3RTQG8yDAb86z0nszpjxJ+b8PlmC3WjNVuK2VTAPtx8IJmahTAgsmReCshj9
rMZGWOGxCqlSMo2Byi9IraTjlKVO1rMcXuDjESO9V4SLPY+E+J2Mrt0tsvkWR3TYRbQwFJiiAVAH
FvQlwG5Dx7JxGX5o6qceFOod5XlzLJb5J1F+JwFzn88258uAlPU9ImgNko0AG/bhmF9GkcXTDxT7
zMXYG4BAsPpEDLtcVN7MpmxSwbHXYP5pMBZu6WJyxntet0E3rZnbSj79540bIjVVBmetdBj/0n9g
gRE+qXJj/9XWTLne0PeRzP6NM2a6Yemlpmn9Vyeg1MZnJETg2d9WG/QqONCfbusz23yIp/FEjoT2
K5UQNupu328xl6a185L2IJ2fyepONd/1CgYDIylkwLIMvzUcecdPT9rLKmVE6xjs/CFFBM8v3j6L
aQvvm/Ad2XaocJjRCLZVTmYrEdC2kZoRGR7QSiikgryxrbcSSdOKWPQj0yq1i4fzh+rvd2vS0ur4
2jNK9nliQ01LqMhU6CEQR4MX98rX7fDmttC+P6YeIlVCH3AfsvTNlId1CG9z2kAKcF4mIfDnKa4I
ABzKIO+jyDxMhULoDrePoN2v2EScC62YE+lTx3HbKTxdK3uG8103+50QMdiEQTDS6L2S3EOjcQ4U
b1JJF1+WDVh5FgFIeIsTbrb38Psee5CUaX4o8zZaFC9WVGDwc5/IYYU0SLfezggGGidzKFx/Z6h1
yvMN6YfZtyTwOKoFPA72C16cuF1SyyWW3l65PXKyLajznp0rwE0v872Jt91SoroQ7g2Vc/x9Np43
hlhp6S2EUrXox0B33tgmBXiaFO3Z5SR9yxzepEXS0S+n0hpuobRv5+K0Nf+k4ApsixuPuGIEGMff
qB9VxNxHKSKP/AMsZEV2eqOdtSvBzPSTFRwF9PjYEf55UO0kRI5sG5w80YVAuWQdBmMLNSZWAfOP
9Eca+8IeLnMRQ+dInaU6jkBhTz2yjg99kAa+U5jvL5w76QH2sWbVqEN134r4/rMIcDRybcRBXPbf
L95LRjpnLvMUXKu0sMT4UM0zls4NB0HL5fSSyaDxtDXddipjzc2te01Ac/nvAeA9fU6T8fg8bMJz
8+NNSogLORrHAgk0eBghI748HPFIJw90Vtn51O0gA1c2ODFGUFufuKzXw1G+/BIOyRKVtDTtXS+J
JgqGoGT1CPBB0hPupxRRRbFPusa+CqeRyj5O8TqPV+YT9zmiQzxNCXrPS8oGKlzurB5kixWI2p4P
2x0YTER3wZiPwnPvmR9PGZshjCyDGmKwzctipWlGLr5M8vqsHcpEhYxeVA1bLh3AJEZKZUZj7Zxj
DphK4VNF51GcRH+0ONKyOSLm2c6Qy3x+dHFP4SMg4HGQRB8es5PWqTCCE+VQc4D0GfrsNZGGc5Z3
sdizLRs++DakBkqt+r33k26CrBmbAkMnyC08WBkoHZJRurZEbz26AvpxRZqs2J5ku4Qp0AFPNHFO
y7kmeWLSLKGq0fPjhzWOCyTDGkH/D1zE2WftGprB5ayEq87OKZFS7Av4pAD8SNDR0ONk8hXzj/G2
PhTa6fm01trwqWnxZxx45VBv2OnwXra8h9N00GM9VevzjPAUrC1Z7VjtU7zBXlvWh7GUb6DmV4qf
MMtglXBG5KvPSCsNba6JZYFq5hj+rAKNzqZz+5LALlXRr1VhSSL3wS51Faui/ESYK9LVHXRAUHcm
nZ29jpfcs15ipm5rF7I4YKr1IP+cU95VSXsBLtO4bx4mG5YJ8JBHivTzi20N0StE2OMU0oobevY2
HcmhNcrXsQkNLVIOC6HotMuaAnRjZ7Yl4F2pXhfZq91Rp4zau6hsdrCKuin5QF4rSXkBBufc8yLx
R0tCCZeIjlQ+sz6/8RwW9zvuQnKJUcDAo8NUIGpqK/VtqnBRQs6M94ktoYdSsWjdXcK3EcHGOixp
+ZvoONdOvAVSjERf+nFxtmpw9Cjt8+RAjKwPhgPZqzS1FVLjnRQJCCwLUqlgaE3Rdg/WPN9/kOpq
trKyCstEd9k7fJACrXdKEJMZXEfRaIU0LrDIcBLE8+Wzr6LP2bqvouVMFGPAK9nhbgS3wwciolhj
0dP6V5VjFB0L5WZkk8wdoT9YXwo5w4TBvtPLFURLPsnhhDHOE75LaC2yTMTBRBeXDwcoTk0iAh7a
qfUvgqMH+i+KYZmFPuDMWj1SWwVGm1f+06wcmJ20mSSpzJvJZeLBON6QCE8XnjGCPY7XqUlShlEa
u2E0NjrAG59Mkz/IZ8g/miieZSCbojF9YT9DmEVGRBTB6OgEsYMyd0bZ+WxeYOy/5jV79q/nLIz2
dbQ3THRUb69a1dhYx2t15DqveKmqbI4atShhS/CruhEK759LSnN5MusElEWaOFHwxl8MTb0OybCg
1lv4vaOhjchvOWn+bl7tq4iUoUHGZLJpZfOazl+HKEHuzzWvuOfDpMjYn+CP2a2eIH0/WG5rjPRJ
DGGsd4ervWvj4/7lsaKazHmI3DMBi8VsFRQyIKrbteZmq5BhGxqZDQ+ViCKxbUFcPiGNrjVHdGnS
rHay2A1Oeg1+GQ0nS9fOHeOEw0N1R1GzT5zkVvRJLwJSoRsMYhVKNSIZXI9Osg6MhJ6liXpF8xXJ
Y0Jo6QeMuzkT0pcLYZ12ge3yL3UFQWzTG6oYaDpn0coaVTqE5hP6BR2gULyKEtOcnW4NTr/M2o/Q
tEg2pwkabfABKSKxgjcB03xm0nsuddRgbV9MSwZMaElabO0gpKl970VZAGaCMeoH4INKk+ZldQHR
7sje/+T5/UH9aMHcUt3aIRze2r3kwzBI06SvYQg1jFntxRgfWBFaaZRjPumHfImzDwky0Lam2wlI
1Y/Q+YpAG3GysiaxUcUteOI36MEylGr6+3HkYWk3IbHNNqrznS9tW3OvxmcfHffpP4fZR/7MSAED
h3bPQMdDldJsRN6fJ3gR9TYkD9Wtt0ZMBbQkSk6rUN4tgn+zJFm9dP9qN7DPf9Aki6lvIlCjKMdy
csWOWrKy7i2e2HVPrZeQkJeYnWuqbRcwjhMF8ymvKFHKYxvSjh4WVuPPl49ukTDwooUnpRseKcf7
gChVJre024EXXmiqlUuqh6gNsFWqTJhsHNl5PxgtUg34Jd7WNf9khBBmgjYW9wHVDJsHIX/sQm9Z
dr7YsKerF5hsLMrHoNyc06Q1RV/3DknVMBhpt273xtpRG30vaCzpn2p/pU+US9ysBc68ssIYJP9c
deV59Dd6hj68wKJbm+P2HGgTR5ySRkkVUfnwaH153bZxNDYtl2IqCv+IbS52+JvVe4YFyg1AKM+R
ZguVZPcqJWHqyKIQNdfJcGe6jacAOUz635TQQ8y1JNZihPo9If9FH+b1C8ABnBj0bquWvYVLDmSS
JmClZsSY+jnpIhU8b+EpzNImJFCm6tJgAkzP+c4yh8ytDM2KLcF39CL9JhdTap3q8HJggTiio35r
VTz740g3hbedtAWWwP0HGGJq2yj//f1VClOf+up5lLCbiUig/xkIzhQncdCKF2Wfm+Le/4kmyz1N
AdUzPPC6YC/DFSoa302Rx3yihh7y1gPTMAGBYDDYTOVqAFTv7c8VSh/RkZI0SM5+C2NBcgNUksDs
aR0KqVvXZ5kNtu6VAYvtsa/Wz0pj/dIj0JrmCak5Z6T2OJ3PV8MXtRvGhzc3WWxpjD3GvsRSA0z4
YSua7jmWyvEM2xMa0ipc1i+wnLQugI7zyU+vEc3ok78HwyD6caQEt3rq8YIZkD7DhJDy8AJHCRMf
mxYx7tmSsuvno4pNvRUF1Y1WvoNfD7WFLhPVPPZdyhbhKVKc6gB+Up8E16MGFvJW8yodADUcLYO3
Cs9v+q18HfnUTvl7uKh7ZJcDwxxaZZ9Fhf+ciD6yH+Q05EVqZZuP7jkB+DNdc9es3/ux7NX1ntHd
oIggDRl2BKkQZVLtPA+3GDnmt90MxMt1k4lAoCdb/0P+O+bDYYtaiY8rJ1AW8Ln1oDWqbe/cK02k
ER6IOBLixFU72z8H87Rs8/PqhA8nyoSGyW6oU84QaEhldaz22v2DNynSyL7W7XLJTpZur5VDL928
6Q6I4KiMxJsMjHCZ9Y/O6ZgurqAKdnVX2qZWHOXe3MjvRqJrpRTAQhSGZVzt5URbmnJQBBKZw7VK
j+AuR7Nui4hkN7QXSKqhTsOvKQ1FBCdflm+JCqyu59o6ekFArn6gtB+DhhYnqW6bo2sKwuTz8g/R
RhNsdy5bf2cNOW5Tu08Wjw/UMQgHYSLKFiYWySYKYeD5yfWaO1Valt+v49Yr1B/CZuo+xN71FUOS
ytdDXFybGW70m7QTjqJE5kN8FR2a27yot6vArv75is4Kvf005+/WbaVAH/hB2ELn3nk6THWVm3hi
MLhVi/bx2y3ft8BO8P8zRJjgvqfMdqVBPuDEwo+jdVbP+ovFuY5PR2th/JtIrjRUZYWtLf0voSB6
kwo6laA85oMxH3aXdd8HGKX3WBoFH4x0Sxc0mOd6hcKwDSRsCTgTYn5WBYvjmBEKFGbvQjv5D6Nj
TlJyAVUaMVIbD2hxJUsM3FC3mGeDbhhtbBhvlZzM0+7gYdTsjcpbDm7bv6nVHfUDTejNPjBeqBGJ
2vUrRlyGVa2/WYvRKMm8S6ozeEoXR46Gc9cXDpgZ/sILeYVGTA/yqIrOx186J44KbO/tJsbwMHIS
JvafCfUzNaTZJ0t1DxoreQY/lXM2ZNX+5f2ulSYbovRJ8xkcZGGNtQz/Q36Bu+0hMMZmbb7yLy/A
8ZhDbmRLPgD0qrxqu6S2XWMNyvhV6Z9Miy7pwNZYhraeGr7yQu0YZGKXZbBR0OVQ88lLG79laUaG
cmSkW0VfnH7AI8ykV9Qu2l9TYsVqsbsDu4fHnYIW6JG6MQ5mTqxTSsDXRoSqanzC9A55PnLTihzE
8RExmHeYaK3gajntknmTmngmtcJfWekgq9s9CQNnb+ih0C9x1ty2MuyuFE7m+B053HYklHDbm7tX
BdXSJ/inRwj7WfVuubVw614rYt883eu70jB5Gui3M+DaO/FzsuFU9sWOgiJw6OHrhde/hAzppia9
ga6HDfMH0ej2tIZWfEsGsKTCBwzfUK6ow5rahDyJY3N0VGx7JUvwnLGnsCgVhGikNIYWGUfYSy6X
Fr0csn4isfS9NA8A10ggqPI2c1KQn+fevSP8K8ej/m9FDc6S9p7grmhTr7Dus2IM4jG2PIvWiZVa
wfThJnO+WDbiTR6tQsDsx80F0gInsa8y3UWKgxNOotYTxqiTvNrgtMPScfLz9w6FdgnyRKrey5nw
xpv5Ut8gWS6iEGeWeOy0FTocKyHhTLuGVSWYeDZeqB28lhUpVZA2o7Vvbvh/YzvllU+MgABe7tUE
VTASOiZIpKuz+z9We+5bOc0KKq5zNlW8aordkr0TvXyPVC5DcIIHptaG6fsSRG6o0wQyDNvalmjQ
if6aG6YsPnmIz8CbRoNeAGGfswPpqk+92t6VxFYs6bwfPrXh87YmmHHlZ8RF82/18luKPRhBHQVu
sDhOUCJrCZVx/NHXwucOgD/awB3krJuMFHajwU8g5AwVPJDQPPpScKFJzFrP8SyMCfFV0gsoZ+Wx
upAJIWVcMs+z0FYPaJEQ5e6Ofgzea9lJYLnNm+EKMO3NARXfGjAkNv5Q9IexYJs1qa43KS2XuzMI
5hPQZJV77J94Aoh1AhpzQiiAvYjTwKrn4aLdbObLaEGSzsb9DzzOapXllFps6zgbAOQjbhsC5LN5
dxC2kypPz3BQvnEOrzJuPnNIDWqzViycu6ErX97DvBj65PGVRhQFOCUi2uE3nzofkwF/idmGEIsK
/fWHJHbAfIoUZbt5Xqo9rq/T6LlcAkWdmX1rMMFKVh5Vjw8cB5mKLzgQzZ0Y9wTxdeUZORlbtffC
UI49hA2gdKDKj3g5yB9advJR7RAznJZXFXFUrT19JHT8Nw5qFbidwtlKmO7oKilEKeJ2hhymH75C
Cijzvu4IWSqJ0Nutpwgnqw1reMChbVamTKOVcWk+UouulwnKs2CyVVSKEGGQ608E7mMxOkwMLPWb
NKVIymaeQaykpxbskb1YXCLauu9we92LBsm+TzqzwMKeeAx3+HXGk84L1qGIfLlR9Z+EMGLmdWTB
nkENJa3PpxF6m8dCUYQTcEq4uJIlYpIBvxD8QWppFBnL0WKKGvyBDmFMxcwM5yEnekB0gc+Kg7U9
T43ZILR3haAfn0ck3Kmr0yzN1eM2e2PurPgRNzRXe/hasQgCBMpUYeSvwvwYkaPnw+gNiXbEAlJy
GYn5c0kKwEQMc3DUiDpt/qGOWBJzPx911cFRBrdPr4gXynE1x3uvLjhwWwNaw6dK/SgS3WOqnRnO
j9JxHRGK+0xOaKMcBr00VIXN9GLdNnYURz1PQ9Qlu16oy+4pcfu76ediiSnNoR+MdqDG/6jUeHZ3
PJG0ukSW69trV0CCiX5VdhvadDi49pUWut9jVf5cS8/99g/FZiJ+3EuDb/cpo+J169aK5uMDiXqW
MdFuFpMNJLCccnRZgkzgqTDL28JIUZ2/g6R8Uo0k4IrrT84deQP7z7Ro1RLIrUFcIreCB48+OYk5
gcYu7VjJ4lEDEu93/PlEtWEQ2ZiLk+hR3QmqQySTwgQiWQlx18x50zk5FaqpycidpxhRQXS2y/cu
MWYlmF8EmQaFIpijS8TET6JMmpMewIo02AHTaqDBTHKPjb80dFBOcA+b+wdcDrF5JyaMWjSxl6/j
4woRYTxpQ/RIhhEosqPX1MsjXeuUbiegoMclTCeC107iFXxn60n1mL4Y92W3J51SFBvar15th/Ob
+E78fmx3DycNFiATcFUtUIxS46kvGie1iQmdErrbBnT0F9U1PjwIO4bNuYgeYI3r8EKpM8pgN3x/
/BZCyYL8AVVMVjFO5kkT/rAaD5BunvLx6hD3JwUXscX3wlgz4G6i0Bwhkx1mferS6egqeb2b/OSe
qxe2aRoI9un5FlK8172SSilZkn1FYXp9vx7hOOLBYMMkhUgwxCgz+BgXKPV6rxJOQUEUdSYxKrvI
Tl9iPtRBbCDMPYVe5gj+wIQKlfnsSENujjbApn89bUdIYhHm8NOE5zcMSOIgXsBtbeBpBeY15GxO
1HpYCmM7cdR6SFQIZeWVDyIqxQrfDN3cLVvKNKV1FNnz1TM+YUgE1EX3E0HHIwRcpQCxdc03mtfw
lxz/zCg0eo1TrJh7/bWahSlpgwa6OUPiutqUL4cJ/Lz9wrfptTSBftTkVN+aSxOJr6dPpoy49/FS
3ElyZYR1/zcLyq2Vec0lyC1Uoo1+ry78I23gUq4r4UglBnCgFZ72jJCZGyffyWmuRdnWbgMG49FI
/0VpJpo8sxdthJQ//Y99757HmUJeTWoVM8avzMN6IVmtBtIq23az8DIzGOcTMLtRHFq+9D5WxIGW
AFGVqsW4Q/IX+/+yI2N9ouXvI0Ai8P15Ln6PrfnZHWoSj4vyvShmOv2U3XPkrkG4Kvw7sDKDYjcf
UJb7EuCkpSMljZVaU0f2iR+9AzhxP6hrp6j7BZ+MCB1FRnkvG2eA/b85rlsDQ1/yA1MI8K2MDZpz
XHL5xr4/cdeqGKMCGuZTkMn+QnA0mFbKaiqbPQk+bQ0Pf70RY5+NlfK/aeKvJWoyDi3SUFc+JjV7
AOWBrvsqoYb+RPe+0ACgUBy7WyFbxMROinfO8jDWym58Yb29EM0iY++hJ6Imudf+kHuvlbooKxzM
ItHH1O+plHLsr29VjhkW6Wjpzbx9zm0A+FzmOa6FHyVsHWKiXPoa55Xy6vAiuvf//xJtItafloKq
3tu6EhwJOEBaUxznnAopAY9CrQ2mAmwZbzxaHWMNV2cR+xsbOAKkA0i1v8/4ZNSMtPIFrzfYqQ7a
oK0JIkYaiU8cQsj+jSmw/8T3htaqNbIk93Ky47n3XmQLf6zuypr+2prfAmI32WrlCPIVoqi8JLOe
IiRS2VM6qlZ8nHiogxJirVnWuNKjd/e2zaFsOgeD7NgxH5GBEVDRnxd7EIBLFeV0mspDkqJReoRY
7SHJ3KJ6R7Yff3rOJDxe+tJRy3nOhV2V7uBBQ57B/afrVvskVTBqdvB7dgJZ/UdC+/Yg1lzACUCZ
RjWamkvWl4UWX21f0dnX2EwdCCvki07kz8JfyQZVvIRwirB4ffW6aadN1CN6CPj5z3gKQ5ueyT8C
pBLeBsljEZD+2mFJI8oYLbGrba1bkCxtcBdsWvv/VNPD1X4MT+6TPXWiex+TbeUiP7qAT1qkXSGO
fFBOPebPxuySunmdNKbduowc6ubaor92R7mGgwNjyo0O5fc/OAy1T9f4SpvT4RyL1NPoo8sTwWC5
j3WMLvGqZkMnMp2w0E36Se+b06eu/ntdDraEC1BTL2Y/zAdHK35ERkEaJYmUqvcLtwo4m+WnXUGj
vvq/MwMJOjrU0I1mZaCCAuuxg42MXD6spVAuf8GelA6l1WzE/OLvObUTKwZr7d0Zgtcek0RqQ04o
HZF4pTua/+9P2a5uzapAmC9ew6AqzrxO03qXqFnVuFxHv6LZyZkTvxWcpoJPLGwCxSILMLlvVtuE
3E0ADfYBQ3QmVFPRKJGywcoejvXcUtMezZd0+2jrY4WyqBrpZKgUMKN4I+29whIf/OZTGJlJQ7nA
KTqJ16RZorZVYkmECETRq348DheQCyX/nQtP1ryKhFFbdDGwOuC3csi4v+b7YiUBGTxKeltLj8m7
05+ELS8TxweN83Mdia/esFVfpLZKPUuNM1SMoGgcTCGQWrEja7ksqzjcjDjTNe/kaWA3W87g/0KS
W5t18qE/a+eIsvWbcaFMtOYsBN88y4EqrKTCSl3R4MJyuhQrBTLqBmdr9bBZho7yE9Fht2b9aplJ
/wbHZ1Is9SWXlCBPLCkI47M6ay9+j9eUH2vPkL2mlj9Phz2liSBbNxTxHAhhhWtftm3qAthN/+37
BJDKMPY44wfWGqcew7IPGwRXaAtZgyaA1tuJZkIsDszirkKEhaeHWLy9zTBZKT7RTcRrgRHmPVqg
7S695qfqbrIwZdE8Lqd4Cu+EqAtXCcrFroAh9zbl/e6a/u2x7J2WYiaqdJheCL49OIc3bgkptvgh
Cu5BtjFEyfQhSvcn0jeIVPEPeKMaz8VuLOy++oJ8Np73ViKTsO0zSH2Wv6T6MP+inQveg7Xdy0qY
eSLPkjQFsOOdHAcZomtNGPBKnTNRMoCtyEFl9nGzrY39IZMwpaiLeHz0ZgKUiEbmra2pxB9d6pPY
d52jjlh5NUMtBHz4Jn6MaheQaTVx1v3/yZC8vS5B0nAVwvnhca8zgziryXeZSHTdWkd2liIRUOiS
es+DHbCVyk1oN2qvi2b9gpIN4NBx/oAPZOOS+fhK4fopKMpVU9iZFhAtUW+ksVyS6ud5vlgeKctK
c9zx3dtYmZsktASNEJN+vP09ZY/kdjFHrhG9kLl02sZNeFXl9lSHuYRc71naOKy1qfyVTUQxWC2F
hbsWriC5kdobqIhGfFBokB67ta1hHyA85b0jPnc5m8GchsEcENwKeDKZiaDGDJJ414vIcjgCNJl5
ONw3LPCIa4pXWkAYVb92BY8W5mJNosSWnQWriv1Avo7ltbNbA0tSi1MVr7qtBYnjaiD5GUslh+SY
C1sfWZVOVKNC+QLhGIkL7vu/LKkV0kWIeTg2oNVPNJB6AX0MhHVQcOKZl1F0PlYJHcX6j0pcBiRF
xXj3EHb2blbvgqSJ8ZeooeUZ/7U459s4CLMVsMGeoP03oWBKJSE2thxHHT23cAhcyJXloKIHxjrY
0HRPAtWiCDc+BFlQZkFsVqnoknm5IjWNMIjcWIUQmaTW3nC4unayEhLx7mCo8Q96qtCtuqNMc/hM
CXrlAmNSEzyswnoo3tcafpBdsI0KPRCFiZHTmLpUf20ZViGgKnNwLGYZhf4jNZqHfhyBpAcJGWxa
HuHDOglGgyiA5NeHlKSqk1eoXWiL8MugLRoS9mzO05zDMccXkh0y5/VuXTlcg7fwcxTucXG7GltI
uvLriDv7EsVOUQ2DXkrjCA2UHlrzZNeVI53zMJbZjho1rGRNk9/3+dy2DCAcDNcnigXcMLRI0hMD
dLpAHEhxCrJBsjyycMhpvNibwZHT+g6KhPBT8JRVc9JQlvdaybHswVreZNiw79csI2cMbIncvPZm
z54ro7dQm5n/LmPOW4D2lDud37Djr6FolsOhzV6rgf8lS6f9ER2/3+Sg2+oI8G+dcm8NWr3Wh/WZ
HI0yoRjBtkh1ygPDgqQGUdPKLkLqY71YA5/YxFV/LA5eWJ892a/AaDTGkBJrZDXRA0/+Zzr7yQBN
EQpndnNUnyHs3Fj5yC2ZzPTFsya4Q8n/r2QVc0CuV8LPeWkaUgRaOGCZIO/jec2tOew1+z1cdLsi
UGg0zsdoQ7ws138iQl7Cb42sKpFLm3DoiicSSuFpfKmbgZsbMfTReDtAnT9O7dTNMFNXdFgUIKF3
sJn+LFltMmgVHzZEn8Q1ML09VDhuZVMmq6jxFI6h1UVDOf6hPE2O+Lw/GZlXyNd1UVCdNNhFMO8L
8eyu9bYXsHKlQ66fnLiTXxVwg87GxmIQnPeRftwiZ+maYyM9g0gWMGs+UlSyclZAErmxjSo3aDiU
nGOtyPlQ6FHqoFo/PahMWLFaP6A4RBUOogfIQtnK0AGrG7SlWmFfRHAFcQOvbeZIHm2tdjxFJRgK
PWrA3RcM0nrWkh3a2NOjcjWOc0jvP0MB43eFm4ED5O41h/iajplxr6GwjdUZjBjb77bagGWZNTnx
ORnuqvDiPwCgkAb7QqMGwtxoKJJOjJmsyI9CpmruzoLtGy5k8wPWwRM2JA5Mhwbq0FWTxUC/FBqr
ocWCV2I847CHwc1U7dN6Q/Djzes+sSpfQF0m+1vh5RQ/dv+GXuBbHqO4o0JrX2ybhEqsFvPvzQKC
5Tmo4zjIEDBOkO0aZcZmXnyhp2avhComQoSZfZodJcxaxT6Nk6Kl01Q//KyH3JWxBkzfjokvyfny
rXyugZCdNMQF98WTu2K1U0+q/CIyv7JAtdJMar/KYqQlMUwcRrKE0HnQyp2wcP0MBFjA/f2K0gMC
UCqIIfN0UsDN6Ii6A4z4fM43AfAK6qHJVfh1J/RqXui6vdo00YGLVR6S10C3i8nttnTwAujouAhh
XXx4COouPuWnixSXBpA7T/CQ7j1EnZsGqidof0Ges4nTRWygfYXjNlTp8g5gppq0zFLQfN6Ex6T/
yD6dlRtxuGrdfnSWM/2ci9ocidc5QC8YjzAmZl2lOKE8aFEQBcdITHEhDO/cjTY6nPIw2Cucg68O
NtlldIIwX7d4NbvguTqRUrL+GCxDjPGh1eFxWG+DLQTyvksuRoSpvalJPIac8mjzp1HYYURwvd5q
PAjpZMOTccxYxSbr4sDh8IyPmj1WE4QAs9M4Jd5IBpGrd7K4cP1hopkNizCqmDTXxbgii6d1gLCe
NwBn2YXgKHooJw+Z7iB2dhElM8EKxSktQVqsuYqsQ1Uq+GMwe9KFAkdsUpL63Tya+twazlDdZ+2S
eiBsgHi5qiQvr7k+KlYmdtFGfvkia298DkuH1R8otTMOh3dwM74J47TTWQKNY5wvPxiv+FDysC2Z
Lo6gMTYWVJGOToVEeBE8RLRXSCfSl1x0fx2oGjeAJbR556+lEcelMMB6wlTpN5jFmGrOrzhYf4Gb
b8L6TQhQtGyo4zksY7l2ewrjbIkhpmLTkcu7o1QqEvVMUARk6RFny9ZT420fEpAJzRf5F7mE3KmX
/SowBomHEH8PtlReqnEN97YmM3GycmGHAHjyr+yO/y2oPdCjvv0Qodf6oBT0DVeeFNg9vmPsZdhZ
OEFUwb6mEz5w1xVAPtmhi8oLo67nHCoGS26xZcA8b5z+bayS27sMydr9O753Wz29nnxSF9RbUP15
53DyfyApYe9SHf1qUrcamFJAXGuG2TJX4z1AUjdOEUtG4vgm9IqN922zhxwy7d13LL5qpcu7pCAX
8Bd1zS78eml4SX9eYXppD9vlt7y4PmGFr4oExcvITr073otLTbrGxUdDuK5pEzYtydAt/WaUQ4Cb
4dw/ANFXupQVjBjw6J+fVLhbsBE5t8ThcEePud84nmE2wEGBFcDOU00IHM77kjbHntDQ7AgXo1Vk
XISXW7XbVTJfAJ00vg6DytlMdLNRjP3Dg6XR9KGAQ6xSDDMil0/7apX0tTeV3DayQS5wV/2MOYOn
uATsxxlIIg7j4MBjz4SN1+3MY7rmgKqoG4sijH/VeLGEW6nZXf1jUJk9syXr0YMJrTHPJKNcpyv1
WDoyxGfprKTtn/xEMmeE5XruaQLOa/Fv0hVsKFq7bg2WeuT2Bnamp0VmJWKbkpa06XCLOHkPYE/b
jsVE8sRu3iXohnZLKs5AbwXMLMJWM27y763L+pN8ibptZEpf0rSndCF3pLPk43MBXYH10kQnQroB
uKoF7+ccDZh7clMyAKSHxvOtmwpIEgXpkAG+gqeTH3XVfuQSzjxwYDajFB81J7fBVM4m0A9wOOJv
yz1xtrC5hYCCYmZ1aoDto1ldBIM9leKAf9JjS4PvVMdpQlM1U3MkusE6Fgj4ntUOzIf3Vh+wAF+G
sNo7EHqhYnEP5SM++GMocch7jd2iPwDorv5lOfYFHp3zTaotRKhTkBsPRXvhEAnKwDzPwxdGBq+Z
f0E5+CYUr/bkEbV3DJa/TGO9TBP3MBWA0AWlXe0N3Bz8B947nAqljqOgod3jdaCE2kUiIMzQnv9k
A+qCvfmIC56YMg5O58sUSZNHr3T/oXm/wSzBoheoFH9eOyHgt3mXQLAGI2j9vsVlYwcwYQzRsVpX
jjDbxyqmpA3/bYOvyjl0vhjjMCLIx8cjAsXOx/9opmS4KegPZ8w3z5zik1FrYVLK48N3GOnuIWYW
vfB8dYxZ23SE0CVp89oVHmTkpF3i2uUPmSb9kVw4kDZ/K6Dwt6ezCQRF+3J6sS6TZo0MWpfw4Yo7
K4ZCSEKGMmwM9xqLP0HaOg9x8AAn0Hn4snKYqJiH2pYtmxm2ZxK0VIKDRG//VjSbWP5ZfTGTrycG
zwMZuTlFhATqH8XE+R82J7iAyfMmf4kyFhLfXMnkCXLa7jQHb+CBiv6U44ryEpIkxTrjQ3n/AUmi
lQIpCqIV7JDR3CD9DBC+oqvyIVIxc6IkCfj4gBkCQWV+ce16k4JP04POKk/0U3F3sRaZZYl3MtV1
j8ZqXjE2MyZRRpjG4zkTvFQyhXx21lUSmxxZZtsZuz0sYtoa8b/ndoeq7jpsGLpyBQLugKwTk/SE
GCNN+R29vEFXrGOddkTeMTiiBuPlgZ5/iwrW9VzslEzPHT/I596z4rEsguFaE6scuJOxlZtnb2Ea
4l1El2dblyTLzlYfuzsrBngRoc/fFI7EMoRAfs6WwrTuukkkeUMILWC/uHg2nImAWG+QprmLR2yP
6fkwCFPaFle1spAYtBnyv18fRnXp5O1H4TaS/3nPuKCDo9igcrjlpfnM8tY8+ZRvYB9pimzBMo4q
0fNA8uxVm4PFa3cn3a5hWBMdLjwLpSffXgoEjfdOv4rUczeFbfTnQ+f1TOCUSza9VMIyvANLyd7k
6w7Dr1p/v6DBzZFSD1vJPSOiAeZWnUIGnlOCuTpPSecWksOcWIY8nBpTylqsJX723LCkZWCFHQk3
Ejx1QQIMJ+Kemk2cBj44iIMZNGqi4BLC4HiuuM1LKDAsC7mEMtionq9pPJSzpgNBHxdhKAHMQLKe
+JCwSSbRsTsUDHPf0lcKxpYTkxFb+w/Mhz4CLcJ7ewQGSNfDmkq8vQvstYvP6kVPqTPzo0xyckk7
YDFXJz7xc2rLeX6SMygrhPwB2XRB/iQZtsiwS0AjnK//71dDddt1hD4vjGx36rL+6wR/QOwfiHj7
r56ZTuYIbylJl+fFiYxazEYfSxLmyt8+Ezanye3c6djAQRyqJpqd9i5Z60h+VNbZJxCEifLj4qrW
sI9XbfvD5cWn1Zk0e1U0jmx14KhqC1nT+X3prCsioHA/trTWPRKf9AmxDXoO8uKOyqlzKDDSwOvv
9hmEaAiKxR6IF3Bg1EpFDLOLJlmvr1UEUp9271p3UJI9VYGzhtTJwa7KW0neSZj97ReDF3gwfFRb
VTXG/XlZXt7y9hkqxNlnNYWWHgpotTAdyjjrGV7ffPcQ+GilJd1Jzwag+r/DY/MNsfIHqNWGM9kE
ZEXbypGU+2wC553GXqn1Kql8Qd/9GjHcMfIKta0+xWUUYWGIxskNaOrDvqKWFqAWSdy6i7GbjgqV
5tk9siH8zvy7WJSPaJjAKKrZU5KRX4H70IWER9e0arERsbuMvy4/rNy319UcYf1Q8j386Dm/hlWe
dzD7bjKsOdhiOHOfrkJ/p+/9OjnzZ3uFkUyMZUKnH93eTBUkYLaZYE1m6uu4oar/jS/NAPkD3N56
gPuLirsukiecVmO/gihPFM7Chr4fEGwfCkNNPsYoIKYHSn1MVaLZJSeFjhysoou/uhgO/ojJU7eO
JFTHlgbPdZkp7BEcBChXPN7NBAT09YyPOxIoPnj2PJAZ6uCsH77UotA5A6Lb2SEzMdQXBkxNKo/z
z5sWvccn6hmnYQlrRej6gdJmrhoZEgC57cqTSPPbR3PvNLKv7o49SSy6rWgdfeAxSqI5LqBH+Eaz
UYH0mK98jXgfBmT8rqRSwcYSh2C7MhZVvoBWewzp+7ePUZx4bhjN+A4vVHNYhP2TzTNHoHxtlebQ
qyTmXCNXDVvM0uwORwjI5MaGJGWYjvxPvph7Oxeuu30APaIp/TZBhnnmyvruXX7WfOAocInmfW5p
cUEAFwJN5OuBelb9BbBx/ol+Sxz90ggUZ63HEpd9+VFb+M4xJxCIOWOzKmGLzgX9ttmDtpU/WyZT
fkEOkU6M0uJZo8f5mic70/HV9fUdVEwqJ1UcsdwXZvG1E58EJmqK9Lw7sa2hXuCc4lwsyjw6tvN6
H+56VSdqmhRGEZpf+W6QGrU9Z+ehAIvSJM8GNsJlO0ylJ9wvOjsYv3kSTlBNT40Eofldc6fz0pEE
3o2X3iX8ramP+5RmB9yNw11AWRqf3e91N+Ty5mYlzq+yCUpNwyWOCDIn94szC49P/8tNoov8N8WV
stMX3eQ1wBR4qIuvimUGyevccUZcGzd4wnVybLkWKztCM9IF23rYRMNhVb3LhDMxfoaqTCDcgdD+
UjRC4pyhBLI/UoIrXLhUZhXZs8JkX9/O1ODn9n0nI5gd1Rrm7emuf8rTuSZf1VUPznerYYQdd25D
mFMh7uMfzOPKhhyYUguSUNtPh6/M6xScCs4yv0MCJKBeyHkWKllxS2TOmJ38jhtIMj1LLEZCvqbP
uNE0clQyGAs5hZGQLmycMECtwJGZsaSwZP6xS8IecvdXer0jcR1HNc6hSQuM7Hjd0lEiM1ucZpYY
Brb1W1VKNQ33KGB+rYbDjvQlnxNrchqdrrM/7eSEb1Hy4zu7obfVdtT4jROEKdr+8L8Mkd8TNXwe
JKj4QE5vqw9UJPyge+DZNSI58RAS9GPWSM+aEeBRHgkChCYxtL+V5K8LoxvN5fALfig6pXfH0tGY
hGLV9cslAN42rKo7k2wf1HcHSW/zvejP8q84nKlRn7wE8W/hRKMESSZQ9ir8uJQaZz5ZkWotZltJ
LCCaa9PEbINoDit9fVOoonnXF0KUXUHZ4Wfto73hJ0jSRiFmjMIyWBFXqrgWuat6ZPxPD1b1dkRy
cNTvmFvQySD4Od67xQWQ2hepzyDRdO1oAfASz/qKTCQQWIRB5+7334ipVedxGN3ea5y6aEkfBCeq
Gp+pYjISAjAHih2/AiaX9TBlaZfGKuB3Esl0Ktnj8aTsK2pVIsildXY8p4g3nR4JoK3j3czQzas3
+YJLrgyBgCpWCm2/0tPm2DmtgljQ7n9l1CtCtVGhsg9drL0D1hzhczeSfD/SSFzivcju1IsKCG6Z
uveqXVW6P2FsBZLENa2UIjN9gU1g9C8sJHsZq9PVmE+WuXZ97N0GEKl4bv5QImOF5P6SJB7GAoB7
mroGRONGIDMtEZmp2Pop9t6OdbMgGQf8qSJ/HaQGUx5nOxNjE5/00adhTP7pkO8stfMndR8LGqPi
4fXfqcV+U1Ep8JLMcC4UKnwACS5IJPa0hp8yXbGlmRabfsDmi0sp2HjZHwerFZCIFcjnyWnwAW0z
nbfbuuAc1Rw0DvlSfgy5JLmOh2V4n/Cl13oSEBr/hunSpM/BNAmJxc3ftciMTPTsaGToVl6Lfp92
YO0OPRLRqFGxkVGE2LvK9ZgvTfRIwZlqdluAEShXfND/GtYxA3Soy3nBF6uWXSr1ExwKEOqtwYXi
RpORl+JQM9Fz59V3OLeN45g2m5P0PTFdirST1QV/3CmJbCA1pxt8tT14RH50MvrVnzmQ7KRaRNjX
WctEMfIKeWykoyDdu3liEjLqxkayYx9OVOTBPVP7RY6+u6y3Q1OhVM4+BHBvZyhqPxyFHjTd4Q0M
BOuFyRohWojFVEbPDY/mZgbcWqaEotwvOOW5XvtFY3nX44UPA/azw8r2t37Tr0Du57Qy9YTmbxcO
6gy6Xa/P890SEXgRXRiOQ2R3x9B3WlWbhr/HIosfq+QZHJIWoHGWJ1EVG2ngFcLIl/yu/6tJu/Uf
bFOz50wVYyM2h5PG7BZCLjIFvqp/3WzTLIEYsP6UVN3tEOEDaJIpduuu5ELan2wfx1D+5FZkveAW
osfTc3DOl/HgLJPZAR0M+KneIuuHVTuFlHOTWB6ATYB1J/BwJODQ4x2FqP02iCjCv0sempihOfdI
Wh1W0/j9cRgU92AF6IzgBMj+OLS9KTlgsQrIpvRnoDM1Jd61T5q/FmlkBkYsczQVE279o6BGKcdH
oDdA80AlOs9Jlw67H6gVoN/MxEyUbbGR92f64yvyGs5JcvKqb3UefILcFyTE4wYVeVE3MQLY5ZU9
U2gZJLRkYIvTK1vSqQgrswy9Y+MBP/Y6r2jni9GgGCFwgIrhR28hAED1LkSZ0U2SL/7iJBdVz2Fn
zzVQ+0KKjpVXPZf3kk7Ncj9jQUHV3+XZYcXVJ2CRJn+lc9+00kk7ekEsmeMhizgnWuE0GqhHlvTF
U9YBvWUiggVhyB2bVoqT75g9rC2hCyeWKr4sR4V4Rr1CZigJt/QP9GylN/Ggwyfm1SQHTlvUJhs2
8nYcJ+oq0s/EYiRcAaPLg5NiVq+6cRDzTF2AWuURXhq9nSWJyIIrIc0F4/vnDXLgM0Hetklb9cfz
uO+549eTY2XzTOgQVA82GOxnyjL82GmxUf7XR3UjD2hudaCgIwAYOsllZ0ZGWaE+XviQyAE0AVqp
NghTO+KBU/PibO8hwcEyVjMpCi3tXRjiJvNxOipWpGiQHE2zhqocq1eoolkHAVztxtBxEiuQPa3+
HMJ2shTGWQ0+noEjCzWv3K78Xsx61H+fSn0/vIxaV3gd1aIuuIbVUYxZ7E+fx0JPaWQF0tdwE8Rk
LGZr+Kd398fl+gUff4pgnI7szpmlNBgR7pmlvS7dR263A7cBmszTBAZbmJFRWcTHT9H5OqBMfRXV
K+cbqxxrgN8zMETao0NVXnIKB/JXLSab30emEyUh+1InZndDOH51/7LNp8EAr6PBhs6BqvDPFFg3
eilkR3xrWKmtb1TRPVLOL1ixV7o32W2HA76dOyuuIRlP/bD0LxLeKSx7TnwvmbzkRkncdC7OYm7M
CORveQAt250awjNNZV2qiv2pgoCKH29l3alatfMR/pFBUIXzAO6tAtGwNGWuvgsed83vk4Ay3ftk
u5PsUbnrglGP8bD3WsxAh5k8hYbHkbMW80lCjjf9F4UHfFJp2n5U9sJnD+jwu1b0zGmYmIjydfJl
M2rbkeOaHDZOhM2wL9woRUndTFCQ6gL0655dsGIn7Tdg6B6cDFdPVkwRKMx7okbU3ms+MU0QJKWZ
sfA5SklJ79dcJoxO/wwQ0vZdGsX1Q2ixrZq/T665voLPeNTWARrlbhcTb9HabiHKnvcWFger3l0Z
uBNm+Ri38PJ526cpOuw8NZ8vmtlRR1lBNJr/aJXnhqL0YxFC9AYJzEmBrhLAAzSHUCqrAAdrCONr
x16wg/fS3+k0FxHbw3/TxShcqIIap8KLDqlJ5oq3UnIdiIWStzlahxXw5W5AJZ0tWSuBZdfuH1x3
HjwvLOjZMdPQPi5t0tO6wwF6lN0nxHuNCFYDv5UPmXtAXRGWf2GibSf8HYb1mYiSrzWN8Gpbl+yP
X8DdVDZK7xMEc2CzgkCZX1TKP+yao/7nyxXfVMQ75f4a5rZ2ZTMlrYr5hkid13LZVO5upe/qUdYs
0q/96h55EozXXji9/IP6srM42aBVzcx9pFCcNgRC3n7waW4WzNqbKxtjsbXfRf+9xItRK8nybDWE
rfcEPcI/SmXzZq9yqHLsFcSYopvTpM8fPjZD5aNuESHNL1tNDp8KF2yUqbtjIlduzTWiv6HwXxez
A1ch2F2KlWHIMFj5v3Ad1eekJRXY+WUlwZsJP9wfS/iL8uswdcHcQv4YPib072NuKvUIGlYsEbdA
f8hrHMqyIJwWifsbXncoZBYoAN9Sn5ilhaAN910t7rq2nAvgnk6Oq8q44SVKpWD3imqiOZvbx/Rh
TnZ/Spo4M5x4jk6VWMHEvUThda7mG/IwBaEa8DGzcxXhd6MSNZ2pNLe/hlr4iCpFdgtS9a498gfp
PIOMBCcU+aZE1eQTGwexAJhoy0PmI6e0oxsw/rB4D9yODHYpb/thdet63tF+DBDe8Nok2sdadV/k
W2YcpyrdCOBxSLsxS4amxZ10Zrqh51mOnQRl0Uz3AnJotL8wSw6Ya1iwePrak4v4DlyKs0+FH8x2
izLWNVIClO7Vo7qf9jzu2yvKbFsK/ZvmjJMJufT21LrSFnHpa6qLama5rePJpy6bIRIbI+p9Oe4G
rToDfBIcNBc4NlG/mpR24bm4WuDCuoIA1/3ZZiXI/7yfdO9Ji7mpKHmXV+3jJ6uwpMMx4L4RArJJ
GC2tAm+Cj1bfvfD5nzQLIh3lCvHidZUP4dIC0FojmwLlGThyBC5wrt4cKYzrCllz6/yPnvLoGjli
i3VT2wsLKDxigg6az8lmJK4EgoLP95ne2vNWFvq9MfDygZbYHoelXUe8ln3jgeP0kCDssiwCwflV
aLluWhDUplm+I3Ee7yrGWkMq/BenJlTC6khc6guaYpgxtcJoJsj3yeC8yX5MyxjVGFiBlqScqf9x
IXrJr/MT/MHGjwAjx8aXebwUbB4nycuoLVv2cWk7BUWrZ9R0AKOlI329XLLQrOVqreJkAxMXO8Fl
p1JkPLurQauZap5cZmjvfy7wntS/vYzrSaHwi5lpfrJVFOEGViInjDSRElPzi40BcF7FlkTkhFlj
ktbV9xoIsYiOfs2nUH2HINSTU9qGNuOhZ2hPIXGLiXanJXVr4qIpAzoKj24qvChJPFLWj8HwZ/fY
O1GPJTyTNwQzEPUQrylyR/Ch6Oj3sfpCECTeeCAfQluebpizb4vQMUjfkEHDEje6+RAAgKrKx2bY
iuLSj9pf35u7PoXIy7R26oLDtrlw4eiwatTbbV9UYFjPEoU26JadRpYst5Eoomd9Db1Wv6GoeHTK
yryQ3IZuE25Xm7Ap9wVAcIsHi7bwGjvbQ2gTtu3NgG5aNtjpdtscLKya+JSXuafAIR+QotzGS5MP
MgQFOYI8XpSMWEExu3/5WisytCh9Ypanp1m1QupEaSRXS5ErdLOcEhiF0Pb58yB+EDGr6X2YESyq
K0dCNdUyqPA8Na0uVS3jA0cRE1Ks6k35xNUBKgDvYJydKSiznO6xci1afIYHm4U//cl1TYjSBPhF
PATd58sYlmOUknGTnvLfrxX5SofUwXmTE6ujXRLClaCvTkPTg2oaznyPDXlUKQ5jteY8y7NlrnTY
56ZDpDeGEDdoQ+rKadLGrICW63yRaB7qgwf3Wp66rszPeKkcjf+VdJtjn/32SohF3SrhWMG6bvUE
LokCBzCG6v/LsSzqpWi5LdGBs68qGP+vZRqLO29zG6QkyrY1WN1t+G4BGAL6rKTjwJpDnFTMH3kX
PqRWZKtgfZqokDHZWJXSMi36tEOqoNwagrX3vpIkeqp+hlKID9lF5V62QZQ3VLvlJkRSLZcii3k5
arvsBmLbzaGgvfkcEKDBzr6Wn8vIemE/vF9YOQwTrRXev65PbUqrYoH7PzbCUMemtdpx8/byRqH+
qDtLbyJ6OyZQI/aK+HG6GCmHYWU8QmvuPo77kI04iVWF0MMSWA1k8NVfqLTKpxb2MMFyz8AE4drw
IO0WBdQ2YXF3oa+IfjYda+0pZECTMsrZ5I3Dw6WlToT/YRA8IeAtrE878v/qE8ijIS8hv3jBdPqD
/WcAsvo4Bg3G2qCDdvdyg5KTUmPl856pmS6dpiBb6HbCefB859K6aUYZ8dzO9XqioC4XMmqCH3Ya
tncdlCR6FQ260DEopHnP5Vvx6F8B61xCCMcjXgHmUJFscysZfF5bof6N75dWI3X94m0xOfM6lEBb
qZ9Hyll7lC+fPRl9YB3GfpU/lepqjKGCK/mq9wOJgBR4fBxE1xQ5J+LNPg6djPht639YwkXjj4NU
wi7W5htQsLeQHZlIWhXtPh9tJ9jviMbaElfHbDgsKZfm2wrtCgHJlwnasQP5ysbgI/jEosouszwF
+SFVFTnlE3cm1AcAY9aLY3Ggn5ZjN3Jns/6nuE6+z8yPLLBmTLWgJGDRDox9tmGs8MJWSlbzpy32
feVnH16DYPYj2z9vOc2I4jYDFszp5bwGWdMi9Srfn/8Q5TSDGO4fkOiYGsydyPbQVsU71S9Udz6X
a/NRPjvEmlUZSbhhwWz0E9m1YeYtE6xa2gFphd2SjMY7Pv2tO+eEToZruGbq89g/ivArylRZmthc
kIa8l+qHW4+zr8ysTdVSPxAvcRjIiG74+T4aPshfkudxL/PXt3Sakxa+H/UcrBogINpStChDPrRI
HVP/xaaJ480yxzazDosDTVi40AO6rSw1rQTAa9op+Os3dixc2tDDmwhq564abRs8EahEQG+VSwe0
2T1ioPzHZpg0Lko/sXr7W0AduPPr2EKnTtijsxmJ6y5t/IH6KSQ1X/DvA2dSsDwUGJcawcI8ABhV
kuGmJIiB3oO/xkjuK/LQJlFkolIX4fOvm6kZvI6ESXiB0uM96k059iPxim560KGWhLhABrFxGtY0
xM24lP3b/rBdRs2HeHxELINbF9Odh+Ap4GSAhI19cgKOoH/sisegrumz05iQHnijJeRWZqBhs2Ml
V4nuBN6ItD6t7xMC2t2FK8kJkMDULuthshGnKvE6qyR/dV16UFFNYPsTQ84z0hcMDx2IglfcMPrA
IHbNa270MC8zwvPAMEsBC0Bo8nWO8Bx1HdjmiBYA9u0nf9dTDEWbjCWwwsd/l6bGWrnmgYXJg4v5
/pbdL2hPLSe/OE+LFPAg1LqNvhzkCiVRbUjcq0tFZNujSn94+IMIS2i/3IhhO8bekw108PGFbs83
EbtY3t7W1hChXv/nK4FSugi4GGpuLCNvBDa7AeayxMaaAzLFrT9CSkR2Zpa6RMvm6xu/0cCLncBm
8NDkhbPSqHyC9WzPXl/TiXpjunJ/bxL+q2KLV8t17r4oUq3tBc2Cm3EKo02aJol8e1Xopi8G0/c+
cqhWIQ7m/55mgarCi+7RxJ3+lSSyuia3qi9i5FwDbUeiB0LR0UO9KpKBvB1YyvjpYhW8jf15C9jo
qP82I+wf9DdFPeS5aUMcRb5Wr6MTQMBVe0VhNRyfMz5MOrKRvBMzBKEu+UotyDwhqGZWwszhN1xe
TDEn59/NvNwKxdrBPJruJHKUjXKTVPCAiDxIEQ6ZDXxp2rF7dkkuxc+IyuBbMgMo9LGCBzGKk8a4
SVe+AZM5XyJVEckzvehd2U55L57HSUzrpZ2wg/qOMJCPf+FmAdyvV1UC+Jm0BdlzZ+Xk7mZ6X7eR
WRAd/RzJItrFQv1EhcytB4ravtGhc74xRUgEEsy1xvuaZJa3iZSSIGKBUMNOtNU3c5xQqefww6rj
tUnTeyT2RSeXy/W+/TP1Cwpg3ypQEJL25uM6qxwQMheIKybHQ2MhHZFzsZslhcFUoHROW6H2tf5H
N6LMV2iTF9ndjr6qXDs5E43VE0ETsSsku2DO3/T4fpdixc4oO5CORWWG3b86jdNEgYKz0A+UXboq
M+ov/DjjAcDkPOiAWfe0Bq1I23I3pzwXUSS7o8K27qeJ0oEcsTDxd4uRixDNc6khsAYxV5sd4ReA
r90BJF+N7HT8sG3s6WNLY4jQTpxsXNmnH+6pUAorG1p6EpmYSfiYpVnKk7rs/7GaHf0L22aVO2SK
FCydKLPJs0OfUzzRg/mLd4qu+MvAh2xkme8QPWDAnyxEWNw2rDfmWdAt2ZdizQcrYI/kelEgqHiD
Dp/YscbzDwcit4o0x8xEpLRTs3Ey7QaY4xyv59Iu6KkBmrBiUzKR682nszyvIPz8i8Ytjgi6ySTI
PcMMojSar7PwQi/NK/g/qnAofFuByEgtPFvC0/6HtFS/5i16mWujRvtJJI44IGR2o7h9+MrNSiK5
OWBlDhthvznUV46eZ2+b8WTmKGK1FSE7kJHFnQNEto3UgkxDTE862FB7N+pB4aTLK+Wwt7viJljC
8zTms0m0wMrRUiIre/mx1pKS7E3SB5UHnIhpjC4ZiQkcEI8Zdy08dzQFhvhbgiJxwREduGIVCWGW
0ZrLY1kULLbmvmOm/5AWLY45oXu/0SfG8hKwNzfR5bD7U+qAhpOvttANTzvwRFHar8eSI9yQWvrI
O9G7I98/ebwc67dglcMm2ef70W9Ik7D4gNwcwaxD1d06VuHO14qEWCn+KaEOQQdOx5LD6ZUnAxw7
Y/aXICyFblzUQSA0H8otfcNSXt9fEUl1+WxiIyviklDIS3R+V/8NVUEq8yUWpQr7vUGLbUmLESx+
HwdYCWK234MbGEAltrEV2isNLEehmCoN7NSrFNSDPmc8H3oMEa7tTpcxMA0URrQ7uvEeJQ2Skgp3
MkdNKAJU14dWL7bBKSWoveWwIZXrCSCLXNH13UqX2jQlLK2jRfitB6hB1hnCAR5/dB+WFcixBNCq
SdP6X1myy9BcupQzkENwrC5H6Oy1Y3kAOG7feYOqEMQn9nG6tHwPid61B0ld9wa0sOF5Ue/t4iSg
aG60Jg8bAd/nRrVVpKeyVuir/3sQwe1Il9ojCCyNsTS5eqS4fzCyt4QApSHhpNF3DrNUbUhcvxWo
3u7YU+K0A48XlyBfL+1xkRHdlsU65BC1BjQc9HekH4KOc03MW8mA+DpEn/y21XLdkm3ocxovQfmV
JlVpT0WzCn9MTm836TTQL00NHPgLQvTYNerbG5NpGD41PqlrYdPXlwrKLx/6CU+9wn2hIbs5afIP
NfBjs7HBYx4caKvbAMtSvnD9b//PDwkn7NTxka5IiHCNb2LYuO84zhbM55+KZgb7TZim+iE1DWSB
i96/972rIwPmwH4PozRU4kqHTKqI4LBumZUwdFElYQHzV69a0WSQWJZdE7R0HgsFaAP5kFtzxauK
Si005ZFnIiPZMOxdMc0zLFmgkfdyKs5QAeS5gpUIM4d0bY9Kh231jdU71cz8GUYacOBV+iDrVRjc
eKj8lyiXq62aFpHOrgNdnGXE2A5bZS2Vx2cwdqIv9dZYYDaRzLFA13aC1FqE+kmHpmzw2cW0xrnV
nTVnp5EOj9Qsjajl734/lqNJgzppHZbdozFAAFdsLzSBMX/qTSuY3tFpKo3AoNp3kkQACjYaVzbf
kari1XS3ovVWRuV0o9EjXO/Nisp8KXJrGQdSjuDuMctydU6HxZywhBHgpojiNFNDN7FrF5taKXcn
wEukJMbF2aYtKlYfKD1d0g7+G3uwzSlS5h3wRhuhbqJhB2DwrOuiYmUqxg/RZpcCzT+KzA7Rl9Nv
83L1eqaYnFEGGueHKTQfszrPEQMfHVjxK3torhNraCuibzi3DF5cbQrLBbpflDMSDaO/g0FA3vtL
CWTSEXDeRXXXR3rMQwlTZjzm073HvTG9BoPlKgpfix4O3uGW6Ss7PgMqKnoklztc2f6MdFE/cbf6
OXSIWKd7Z8z4L0ubQBEorGBB7e40t87B5uE/jw3tSdf7ZNswUXKYzXbLRtQOaZABFy3J0DIDk8fa
8RwsW6iktdp4CMxfBUv35tZcXcvM/qGy30di4a5q6oqOX88X6h9lJ9+HZ8gAfvUv5HeoEMb2rXGe
/9S/+1VPfqXbOztNSqG9O+AjCD/d6+ER+fIlWtopLMgKrongKaetzhH4CJYuJt86+9VWcsAMgvQ5
0UpyWF3hinzJmMu4dXJ8dEHIqP1hs22BTySL4/l9JFujEPB0PkqSEoyLFr+tT/sWEJAyhKp7SYfS
xWdstBnkJWloguJxfTmil3S9WY7xmpYcaN1w0bXnwRm7d+6zIu1zh2grJLZiuN/pvz6gAeptsXx1
N1L/tyv56gyH0blMmBSwCMuv9If6YbnvNO+rgCszJN4XnDNBjuAnUScc95NITKhMVNvmJg5G0LOQ
xGZXR+hI+7noGEMc2ZGZvhZtOOaFqkBdxOTc4jfuOIpiA9jYr/vpVMxUcRjpYn5XQUDMdLeg51YN
O8gAkvDzhbK5EnFU2jldINmWNIuIOSq360T6QmTzRDU0dC8hCUZSICKhnzjDuQw9UIRIBNv8PbKd
VlYtha6VN1njv2BqOafhleUbB+/f8mGZMCMu0CW0HNtgSII1khKfYA2PaYMPxc188ekw8nXnCSql
pgF05tz/dn+Xm+dG2hA7XKa3e8rVkmVylSY8TyXJdvH3KcZJx79lXireZb5AbBCYpvEJVFjRnvkw
sEFgqrv7v3rQth8ExH4TwlFAb4CE/JMxN1IPSk9eJgFUnx2q9+4Du8Xukf8R05DINkGWIcIiBIrM
vcjgcUmMzR1oTQe5yy8NK/sfIBDoAdoDCTJMuyzeibsggY3+NuO5ruJEoxkIYWRxdfr/S6k6Btqr
D7+U4G1GrAbApg+u0k0zRbXkeaQvJiACgTEC8wUeonMPDEwBQPr9fnj8NvBrxfTSH5ZuQBy1mttJ
FIB+wCgfdJOYUgcSQdAT1V3YO7y3/1Nlf2//UamPy942dEFB0ey3wD8nTQyCj1Ozep2wwcyVTNkv
P3z6m1yWLem6Zfo0vwGRxZlRm6Jw/Oz8l4JVwm80pOTBS0W6v4p5FhIugyi+ndzQNOGwKgISQ5MC
LdNWCBIeXSSUZ7mLY5q80D7B4C9M3ylOHeLTkGZ3XVWYtAxPGHkzNC/Z1iRhT1mc4kCagZm3wLQP
w+4MCIp1CYAsqyAemxo25KpmAXYg+nzwUa2O7bfZUnO4OpEf2R0kv+jty96zs2Pzq/v/YU39q8jG
ecvVausB0tVX/+WwrdGkQlV2G4GdBolzCFZR55pVW9+qb/JdaDjyt+Ad1I31ce/yYFb0NcZ1lTat
FVxzINZH9xLWHf7RokXmCxkDoUOmG/dFzdm/aNyH5zpSPiSERtQa8ng+TDtXSJtIbzoczrCp5etX
jv4VR4UDNLm/+GS5F3qvlo9nk2h/+cRgwbFIntavYjqzoqdo+c2nEpBwRvzNuBZlTrRUQtdGMKg6
ji1nX+jWK+J0zeByGG/toQmSWBqq4J+6M/IRAz/RPCgO7cuJHJQ9yVAt84D9wcGU5gusNSCQECSw
+yBYm1zW6QFBROtJ5kBH8V54o0keXsgCU4VPIJKMtuFVvTKLYrQwxNeA+YwvKSlPfJPIlqg3wP1O
BZEbgDQpIGDi/+QmqZTtx5FAAG7dmvYFOHzZVTR5ImOYhhwZIxEnmJ4BHjTtmfB4gnAf9M59fl91
QmzE20tXxRE5kgRuB9/DZvfy0Ir3Q7hf99DAFqV8qUiLWdA2QKQ2Gp5k4UOpozydct3Zqmlic7MH
7xU1uaJmppUZF2yuvx6h8mWzUcQy/ue63D1JD49No2hYsERcxhbTIMGH9r926ypohxvNI49gojmu
vTYp2bkhus49YD4PFnHgGBMVdSQu6E63ij4pmZICHCiovpzM8MT+LJeu79OG1lzfbQx0SbXix5TT
6EDsQWcObEBSmbmR99zJ+VThV5IE7RuY/VDXYNnqbmIIe/OmIjEvIQEDZXXcRJHHnE8oWgLvzQZj
m8cGP2POhvxQ76n0mH6VMimW0ljwztWSoYdVY3218GqB0xXajor2rRX4fBQn9HYQaGtPBC8Fy92f
1skB/pzOb9oABZFR88rtD+XLh6DPtGr54Zn6yAZCvO5iLNEMVa/PctmjGhquoOTl+PpBWdlcdpNQ
W7/f77SQNyZzKAHGcYHTl3e/oSYvvtowb0Xnqg1HSr1h+ROsTfftmBoTFuU2lTe2cJOKwa2PXE36
AXD+4AtYeIlMXkp5tFcdfEnazZItyScD0ft4w2I9pi8YDmHxi+0mu1ifUeDNnqDyits0Yh/vUPJA
fQUF72lRIEBiNzlYXO7nz1kqTysUeTXNmCKoF0/aAbXWMv6VwqpVWmxzIHgLGY6Xtx66Binlojn4
98Os/VGmDzzD7FbQRgFBFm+u2mIz4LYwPbfkK1h3aCWTwSflZ4G4/XtA3fZS7aQd59qOtv0eluWv
4Y7OGpYRcRrmFU0zPwbUOCX25uJhL6ot3NedyRyZEnKV2byb/MzoDPEqfHoBXsviBvoSTikjmZ10
25CGeVS5ZzoLWmPsd12X6iysl6clQfdlUlEaDe+OdA77UU/mQ5RaewQc3fFs9sTNg+tby0b1kNnE
X+ZOBEx9Eq15jUokOZ+XEuDDRT5MvRbeNUXGVOG2yGBZk1bkCgXUL8iGK5xntHB5TJMgr7LIXjhN
/OgejVipp316jRLklCdZV5hJ6FlDODroZ/xZjvwi+7RPz0WWhBilRNWX8SLELxyb810gh17t86aM
ARBHBhnM2sD511btDlOLaJGplL3q4OwDoQQAIB05sRuwvyBLgjRzmpGsLbqaf0y2yYp4y4ZHDd3m
5ka9wQ04iPvV7Fy6FquP1+fBbOt6sEcj0cMBJSkqPhplRTzFxjnQLytFBUvmscc0tNrYIh9WDRGj
IE6isiNdujrP2ieYJkTuutbGaF5gD+Sxeb/SbGUFq2nlhvh2uJRBc62H1s5HnlXxXS7oOz/nbkkj
E0m5TAf7lWk+k9crebYJD3flFYNV3AeUPBpk26IM1yEOuyFFfWqYkaWtXpqJLEYSUeAPT2rVZl1s
wiZ32OLqJ+7YyzagAwGzbWQI7JUxVRYps3tqrbwObeKplUfdETNiPYDqcMt5msDs3OktC01RmtBB
jLY/e/ehkFGNRrCQ57aEAxS2d6CELf7W3A/tq5/RD2YwxW5qHolgELkA+D6eumflJtwVD6HegPRG
45iEsF0iqkOjGiHUn99k3og3dEIAj+fSdECsIH/sgr/13j+/nVcFaWRs+7oMK6b/K6MJrOMYWpZA
pBqvXWi3n7UORE8zGPfu4igPZkS6CNLzpmT09wFp9yGQbXpdaqRd1iyGbqp5vVaz0ujuDdQdg4kp
kG9bWhd8AreneLXdyDtKVmcbozWIcB12b9spzoCCdPVHjPSZ0G91PpgV38JOsSlnbypsZQIZCW66
AbDbSHmc563wkKiXOGlG992hhi9crJLbVY/Hf2r3sISk36LjUCHX8uKS/vD3f8mJIv758dFdeboZ
b34mvBgrfgXP57kHv+q4VzDTp6JvdmX75s9hgVtT0WRqms7SujDnRdoW0IW7iAPLF0WhWvNEIyr1
mP54ebNpIxKuAqTyYa5tSL3uUOtuaRI+YksmA0WeKpIj3EfCFvE4jYXFT/nRLtAFHE6+7MlcRWK4
8eGCD/jUdEyWtggIxGqW4iJJAArLAxJUjLmOK/nT+qQD2WMKB7clDOjTX6lt7X4ZLBCxEQrOwzr/
nmsd0tlY8IVeHZUFq8ii/lsNVeE+ECtGWCoXGRjW4q0u50CJdTjpWNwpR6qL40BG1O2k7WNhLMl7
qdrMXBjuo/STTn4GI/l9R2gI+xOiPR8ZtZ9HJlLt6vUqfVNq0/NREkAyhpTu9QK2aJqDifxqzJVY
czHDWztaRex4GO7nOOt+Cb8S5N+qu46ZtiJURqfBsa+O9UNBZNZE/veo2WQ7sCVff+5G/YSjyc/7
685m+KsE8L2+yFc+bcOB4fzPmZwJ0VcbxNNyraiO9QMa045azr9t6F1Ky5XrB1nQyTv+EvR638H/
KpdX6KuNFXoyI5xh3IpGEv1PvbVsLeKZYNhfakZu3C5L1FdhZJsBkCDSUm/bGi/9pdqXnbAapIfe
GI4cp5pKDGyyF8/OHmdPClxet2C8Ze0YhvA+/Pdt48xTpeAYWDrTcqVZJvFB5T4SHl86yh/gxbNA
dyofUO8+H7sT5obnNSKzGNLUGqzJ0C3GCosdhoSOMZle7GQYe4aquRA4QJdO1qv1EDr3T6qkpkJc
xxh9Ei9jUsB/4R4frRVzw4Nmi9Yi4Lx82+BKfRrtk7Sm0YSigT7RXaAwqpsZC1/t1v117dlilC4c
U6R//wIfcCv7M/VrGwmoYaqm4nW8kiubVlU38rAqA2YWxGqUxox30FBHgg9i0hwn08+sCP3Fv+ul
XIGnoU22L7TEZHuGvWWyI8ubqMSB1pjMlTaFxvZCNYPxVvunwvoqQMdo6ha8DWSdc/8ZXf2WMEAq
vObP3ifuLCnwNFUSjiuKCTfh5NEsDPhEGzf2Zxq50cpqRmzs8s4OTKlK0xDkCTO5bX5oQpEWJJ2b
vs/XHNBC89I3fzB9vXBW/E2RMu14k3YzMINVCTqJfezn/n7SRjPSMdzDRJF6H9/FyYE3L9XVOYT9
+rDfOlFiEl2rDBbw6pNC6Y1KIktRHpQXYnkw2a6G+i2xslhbbQWbm0zql3zOnu0m6W0Ki+yg1jP2
A22DUUbzqhNzz5SXsOMkgL/xH4EJVCbIgH1W7ED0fG61px1zpQ9lgTWhpAjp3WucbWnwp7TWnnkm
D85pNutxC8cYYHdqXKregX/AA5QAMLx0nBMXTH7rME+z/NfbW/U2CrVHyant6tR5k+h3neAstL7H
sCNy/mqlcKPkf/KdhScBtXOtYyPjB/M5+SejMGaI3IaMi1HG9hqRqHd9t4cHbPHPxbj3JezG/PZw
08icJ7jvSUweDVn6lw9OVtKPdcBQlv1wkFSaykBnDiGmP/rMVrj+KvQpNxjTw0bjzFVxYOLgR1PQ
Ff2UJIOtxFBQtAWxYB9CUCHEBJFkqiyJ8pNnEVG+5qSzz0e9us3zt1xubrN9XHVmS/8ZS9hQqScF
bp/4HSKAvYDZsdIoeGOHuZF3uSifIMBr0/YEgs1ULDPoHkVETk9YQwLLlpY1gYwsIAF6vxYzRYF8
6i96w3FDCBJycn30CBXyebtjuac/4nPrKJ3fBd7y6HL4+UjF7YkJRLVuNcbLz8QJXzrSozI+m7mA
xwbxxoc4ufsw1OJCF/afbOzPYrgw1QiOa+MZ/ZNKHbJqzv8aH1gZxfX5/vAjtKY//gbf40mOpJFs
DErNppiLRm7nXxBqWhknP+Ql1Fq2gmqXz+aONtt3aaFZM4+1McB3pAWLYlz6gnsZR5xQ0A2LiMW0
hhTzXmuTt0XoT2MZlYkwNAkrE5LNM9htpxaWilrS9gmiHOBGtkIoJFF0m94Hawbb9buKJf/lS9Rg
dfCYn5Swz0UK7O+KIn7DcT/kN33dJpqyWxBBzQkkxU/z0i2824Q+jgVilQz4fkyh6hRtWujT1LWm
5q9ciBpTTMWNcgvFdpgs1y1M7Dh312uoesFo8HW/30GMCQCTiWH0gk5taqEz20QRK12D2S1qczuA
5CtyI8lEBsPUC7h7ngCaRiCdaHl4iNKLC6jKJm2jNNb+vTOheZo6mPc27deNcUvivXdAuc2w+Jgp
J/KHQBj52J+Z+Ba9KD7SKBIDS+am6cRJTZ/WOFr15IGyb5PXDdrpPrAcJSgeWtwHQJ1KD1sQhueU
RvtM7zoAoXSC5XDq2mx587uNrKGHEVRravJYZhqdNFRDLywPs1FVakRvVBzUhD/lVQBTJFuc3NSo
ypOT51n5UmxcVDyatWWY9YV+sPxldYLK+WjyXRVdk/yJIWkzfmx7YeIrDx32Xx5Fie1/0kYlPnrD
qPHS+T2C6hKvuunizsBuoSIOiCcU49OMQJJJR4NuXaFOSlB5Nkfp6SBFSqcCuYRSdV1ToSxWWvqI
8U6SViHq4+y5+EcnrHaOYH24KZeQXCEc2V1/+2QnK6eEaWUQlUtWGX5otBqFpGRNRNTFG2NrQ9bp
mO6m1GxzNpERvaQ/vcsmkFvSMls4u6Iy07SEFseawrVU9LIQZ++aZGF0xhLmLJay+Z0sBE3caJbp
vhxQ8KzFlYflepQxc0uppL9qXl2sEiDufyttixhgKIm0r65cKTQV2bBTcoiq+pXTN9YMLlQnCzww
7pNcAk7piQyMnEn8CXUEA2eyVgToImftt3x/mEMzF/Wr9hx/maIKukYs9UrawOIsG+uTf6SQPY6w
lW5vBkd1kTYs4ZbhX/aXetTl1yd3fJB1wjRCz7p2QC4HNaqmaFJ2O1qGm/NNFQQoGdWph8lHuYXO
9Gi4+qxZNgFFLttx5Y0omjn4xda0uwkOg9vWUvNuIn8pW0sMXtDU7mbZT/A1Ve5LDRRgdBWEdlwL
KCWTb4iP40wcoxhRYH9br7ijcIXhgC8kvIr6vY5K349LZnszOPnEjTIctL47c/S6/iEzZWOd+S+d
Xi7fFy79Fxg/8kTTr2CQoHVkS384/n7+yjsgnn5jRcpWXqaI03qLed6jOQNbPvyXY+n+E44xwNjS
Zi3wZ5UQHdEVGOIK/0Cw6KstTArMpBTiay5Y3D8t7lAarUnSqHFruOXg2c6HnQvjWP3EwDCL6vyH
A+lRNliRERGZ1dC9uzEy+7lfmkO84OxViYV8AQbJG4VcX+sSHQtttask1futp2TB1PVlkGao5RQK
6mZlWQjJ5oTDcaRA5wJE4On/uy9Cc/Y0pxota9Uh1QkLDXou8qdpd3JByLS1hKBQI7Ux+m5O602J
A/gxdBFkgI6BaacYHkZkRSpoBStNp48n233DrB6H+j+o4ksNwDai9pc7zFhTvXIxY7IlPWhyiQw2
PgKNglPgsW4x0aZ2n+xgqxz3c47VHcSXK9l3ytXFc27xAazjQmgDARUxkD4hj7gJNHVQiEOIhuru
dbTIwuE6iLWf5mn5N6C3219qemXYAu0rhESiA9rHPoGsqdbDZEoLR0jKYkFF7EUkgdu1eSrGdeZw
lowrQoNJhxa8shCwffJ3VS/K12/7S9rkVQuCtNZWMCT4EnwefQPQ7QNh1sK8eOZi1xzYOdc+0q9m
zFi/+H4NedFtfxvN45Gw2umDFq3or+h9YBPq2T+N6ZFacigSEHqRXvKyfLoXlMmFqyJLsWVtIU0k
fhPnTo+QrWLbtaaT8MUZI6eOxfQxIS4e1Z07bAAW78HRrKCKndIn7BPvVUIRJ8eZJFropbxz4pIm
JK8iLNG+/1f2yatGxmMJakhukRimPGJirSND/Wm0bdYacRrOiP3f+9KdnhDbfLtcmo/R9W0oHrlY
ADZxjl5W/JZeCm73eWjD4+2A8D+BkGE9DoGi0R9Lhwnp0BZb2azjkjZWRThKL+Z8yZGciglX4HQJ
cnLk/9gE2zZq484Q36rjjl0M0p88mo3Mzxaw/cmmiwu1lqzgtGaYlEWRAr7icxo/M5T8IC1MoRx4
I6rn6q9YwxAcpUn3J6phExp/BEYTZv0MIChhUF8j58gsiO5Ev5lPr0+U7WilcbO/4Q0j0i06siOt
4na0b1yT8zeTS8Iw3hrYXKO+UJp2tvz8INsAFDfBdgdZoGAxxK9kKOGuSxWV19eqv6lIYCWi+nGD
Xpvh6zQuxP4jVUpCJkezwRFrKrYR1X3XAgsl6f+jcxAOoQNCe0lioyKjY6MJIEGi/2ny/tCYaqUd
0qdU7UrSSadGq8vH0tENhDpWjWIfwhVjmHkL0OZY8k8zfYuy7YH5NNZUte6hAa1wOFCpfTUFoESj
pZYwnbAQlK3fdDCEYw0L/nyWyE4YrwGTYRo9XHYZ9yXdHHS4QVcxi3Nmi9zfIwZWj9Tlgd8YyaQf
ysiRUSwk0S91wvtJ9vPndc3sJkpWvfe3ifeH+DZnUyVHCZ4KWolRjhCS9WJyrrkqHOSL41l4YJ8T
HL7CI+hSucYHUpovJCQ5j0uKPsj3ujUVyM1XQT1bc/tgFmTzNsFVSaRDO4KuXMSemY0kFSbqicE+
I0YAAg/2ByIm69RFtyTldcqe8mB28QqvmffmCxRRP3Q+ngfOpFk8+CP7BwOlgW8Vuj++gV5iWJhp
JpvDXbLlKU7aPOfK2e4QlikIGCkxGGPLXOOWOuX8uMFO/SRvd0dMN3bZ0Wo7Pqayq5gB0P2UplcT
0Qt8HuUdRs3gqykk4vQsBbZw7/+vA5LIUsEd+9nKQmsou5AjtsPfRa3GRlBJ8I+lj9gj6H4cCC1B
FjSZXvggKlx32PW15pc7VEqj4qQT2pXiNqWRZRfb8kxNSHFUhZXRoVIXhVzr5YU8sCXLxsU93qPt
cl/6b+z9Gkp9oPA3rXxLDB0OldC3udBCjoIjQ3Qb0RO2JLSVqI3ikRC5HfwtFlPa3W+rJa27cPYs
4kB5bfgZ4Ct1RPvhKrQcFYDWL7HnWpYC18x0yqhYAjri05ted4r/dXAzRJfMsLmSl80Xj6LzBy0f
KVe9FBcY2GAOsw5FCeWoR9IDTZdkVn35I7Qbw9f1ei1/savRaekjObJOFbJ+bdWxEA2LhCcJIx9s
hHcX0jKv1LUZ1EGK+FUz5XTXLKoKUi+Chpn60bU00PwYI0KHHzLc1GsVot6vZAWm/zSbnt7P4A/K
e0sIT9+DwsOWGI41rNKCDnSPHCGd1LTqLhv0CAOfx7vgmq/NENSo9YYr5eK3/Q8npErq1b8vOaqk
yi/2mNplP5vFmv3tM51R8YUEWzQo8Pvg5kFDSoFb99B0hhLHEgM2GTEsiIs1AP255YS3B3ABU90h
zT5eTTenWBc6PdSicZLYizafZAQOlCqs2BlO9jcDvcOu6kvv0SSkk11t/OQvyi+zqYddNrcGpvo8
wM5ggnLzC6YItFQHqKe7sQViI2A9QNo1T6zXw/DLR3L+87ADDQsnkbj3BZjst1eaY4Wn3Gl1dSov
k2BiC6QiKrpmIbmkwHzfEN+OLrtG9SlmrQhYzyIe0slS6aB1serOsWo5XDfAw7jLmYm5ExCzc9Dv
Jf4Rt/60J9IHVZvyP+cwBW6F12Gc/D9CW2zn09gQIEB/7SkDvoow52WiE+yA+z5R16ETMrpTRTgj
5nabCW8JSb6BRjb9PZrceoxzc88li61+2Y1cAFus6F7XVqLnH85QxXOz9a+AXSCXfeXxSIcPKDiB
wZDv0dDJFxhmcW7Su1c4UO9oStgZizfcCSpVebnqCcw4Mf5C87XMxbK0XOv6DJWrtXLPUB9TaS5V
hUOHCh4i+X4Q4v0S3Qhb5B/up3vTWRzZAorTLcEvZgYUGnH1i/nUgK9GMIA12QrOXb9QoTrMIR4f
2MlD8rLR8PJ+EAMFN6L0Qd4pYPVfxDN+sPB7uq0azolAZIsQsrGQ5C+qpd5p2EmsPyFGLxRNvadG
+FCAX7cTVfcHNhmK3LP2Uoq6h1dFi+PJOt46LWnBNgmqVHm0hg0/IBIYH0aJS01njWy5LdnZk6U7
TrFpFsGxDa3BuW6KDIkBgTr2a0oJyV+LkX4sDfWY6UNjXInqgLSdGShSM9TqtFKzpgsi7DMezYwu
aUCKSshYaW/gTuPK8HAZDkSQ52l6QacJAP0pq7s6rLOEjnbhjpXHAfz+d+QLhb1MMuuH70isGCnw
AUynpN28dnE7pUcpsSEDjUmRke7XIiDdKEzNWUqwj1K8rqf9H+LTCjkbOB5OPaAekeNoBI98Yzkj
FmFjZBIY7ANZ49ekUX/YnJa+jFMsjLFrbgSDGWL+E2Dk2kXQtyz5vjvwzsyrpvxr8JgDBMM+jW5I
Jm2T2fdjlZej1MZ/omxX6UXfPIbhQOOz81kMU2Ba+x7vHH+mGMRulghC1d+JtZswAnKNIqC6QoTJ
3IjjD4e17IhLuEkAt20Q/+0LVF2oaImdJOCE9oOLJsd36kIzL7HfLI8Z4jc+gs1Nsf0FUOiKrDq8
iz/4a31GwFtuZBUhUNCuGWum01qVpVDE0RLKulYCKoRGV4yAgHnEGYxxlTD3Q0MR+NXB2/6crpgV
TWTp8EiZxr0k29BbQuGzsoMPQx2BQbQ565V1e0xXCcI0BklXzUtEVC9rHyo/KY6pD5ttoibfeKsg
SxwRoMsJT9gNBe0Li1yEoGkX58zuyGyzh4ZKr3HXSxf7g9+nYU7HluQVPb7MiTjFVzZ0zM1P5mFh
fYJFRg43Dh/ySBDFOEsHjZbVKm3BA1I2BViVIFJuOQzDRibkrQRJeMorRcr8kCUUNedkof77C+3t
vQF8e8bIE7lxM1olRlOvLVogQy8hRP+P9R1boTVrE0NnpCZEI/dHDPKfzgaU2YBFw9fJoQoEEZkx
glNUrDehC8cxiOsxH4aRVUoWKCQ0KMFb2VPyDEAeQ+aH6fWfWC7KBik86VJ+SMvGR0p7BaKUrWRs
Yfk3ySBnG99srzt2uMajyxoIHrEdzOYqWoRENSdMfwHaP4eZeQ0DUNqHLZXQTnTVO+16kRhp4RIA
wROAZ4CTVtCt0OF5grdBiNEu9soGW0shYx8URG7JpcV40MSdVIpx7z99OxiKJJgnbz3KKWy7Flyh
Ig6JvLySKoNwz0afvfpL3ZclJYzaNosTYTE6L9srbUI4yA8GPKfKGdrGRE4wrvIbSGIAFQQVDaL1
TR0OD2+a395MJyXVUwxs7zwpk7kW9VyP86hWLDjtFRWxfC3shOeubmwSoITAmknctlo5x6Z0XtG1
Dk95Je1WEFwE1j6He2sBAdhf9p2WibMhRl8YUe1UP7Rs9pROYvKieNIkRb2UfdK2el1hGhWJfldQ
nyCkNonKMVsn8e7SdYWUnIgfG8F6/IppY5YidJATAyEuMngtneBmXtfJw7tYPDzhdjitle3+pGWA
CqB5PR7lth4sJJvxA8EhVY68yhTF+Q+qVaMLCf6tVnjmF1NEnZrt5X416n8BV77qByiQtufDHYqi
TEzzWtgZYK1Hq+71yINk5xLfBUyfthS/CSVtZhOGD7fioc3Xi/f2gPWHJyPr2ITqt/1vO4QthKgN
e5EbLyAWLfS4KeiHn0vyUm9f0KxI82nf8X1LHDO8bPGynCFLmF/0GjKQv3jg3o3/9ol3lvEYLDyZ
6sw87UBcWHnFo51MJEh07kEJRJtQD6tiURMmWXnk6KBKTULorzRE/6nK5SDOKQbk8vmasK/Y0THz
iSPWvCI6PascwS5Q+Y40BTAgvTrCIZxVLeovWJbXDQ2pAT1twK2MuIFl+HX9R4Zu4ddxZh64fLZU
93UFSZ/EOtSo7RTIx0moI9cE/32qlN3IoOEhqgLzUgNiw7PQho1weZ7hAJb/Hg2lQEsSqUapynwp
xhZLhNTJgu61j1ITQh77fIu4f91zVWrId/MziQqdmJSYjGYtA5xX5UEK3a9p+VlRxN1d8ZaqcAjw
28iCtJXNPpPJ6Kw689ymBWZodVZxbuxkLryNOhL6avGXtE5n6TVXoGBytHjqLwvXV7PMNdVU5f1n
ngbrs3y9zF/YTymhN8Vz6jhQT91/l7MpP7ALsYsm1JNHKirzVCx5W/nL9VTHPEgUSzG9Lty6ZjqX
lFTRzow2OHiq3J2A2nSBkuI1UV+zwDIeRB2s9dGBRgGD3CoegTca/lWOacj6gADF32F5C3C9KYnF
Pd+gXUzlIGmEqemX0kjtansvb0Zmaq0n6nir1ssWFoPbewf0M3SWalNxhot30QaHQ1Jv986cWBkm
zFsVwOGjQRCBeFDwYTIw+BbSCUex7G/Zv1/qiy79H3Vl1IQMs+X0Axnl7whm6gmUMxEbDcpJKnD9
YTy0Euq4dJTizpPlM/6ZXA4ivTj8sgrX5Z/jEvcyIL3T2xxuTkFuwOwkVk/4w/OLvJIlHNKXH4ho
1YCuR7BM/8cG4J5Y+f24A1+MnJrCSKBXqt0UDfhJdVYpbAt73Q8C3/X00YzPoO+3I1J9T6vvNya0
WyrS72yil03kCDqLt8yhM4Uz4w2alYfTR2lGR1nQFITpeSE2i53y5im1cfnkWUDbuve/8w8kSMDo
rQql/yzLnIGt8U76B9WHF02w8vQfsi9KMtLAzoyE1PKYcQwJwCqramM87HUHiXVjc7NHscup1Z2M
2wcjreiK34d7nLOMWhIMHae0R0EYY6pHW8PD992IfU4tbzTWBf+IbzMTrzfG3yns0Egdqp7IJYCK
BJIrjl4xGCIeR515oaZuUdiPMskviC25pjZHDf2Mox37foyNOs91kYKVh+0HNpUCfheYd1B08T6G
xr2yrT8+SYTzUvuiGXMazUqoV4LWyHn3SWWwxeE9+jWqMc3UTR4NDNRoCNxjZ6hCRVgEcei1V3YS
R50jwGtJerY2kSdloeOlcqy5z/cxq0RH1n+6iF+XjpIIo48NGpZz1WLUTlN/1sgUFbXl+f4fPd/U
XWf+I+9CkoTzbHy966RrcDurgiOibhIcHVBhRMswg02bTUeoxNWjdZ30Oye9YWRdCFuAGD6OHLLR
01gndTR0m2tBE+T+XWnqKiFyi77kjnzC9dTyKoGEzBvRJNgQyi1AOCeA3163x8IEI5DVtrJzdOXH
9IKM5ZHJJyae5/YH4GMUnXjbXd44NWgF62e8fUs6NDA7+/Yf7tNpwEMOmJsV1wAqe6/+XxudWOHJ
4ZgXMFAjemfp5avN8pufhQ6psg89spfSgBGyiM83ZhGdo7E/pKjllCvc6vH/gLYumGZJ5wb/BEkj
LcyG7v6cZOEwMWHkZBQH102lTct/L21OAcpoc++tj66yex/bgdjjbylsGXQ1v7uMWuA3cqvd89Xw
A01tyNm7Q/QU+DaKmlIoixOwmDQ9dJ8lnAu8kdeo6HeH3Jp4vYnLwEWo2VgTayhcqO0/Ww7ybHJc
lG0YGVoJVGyTQSlQNh7K6N7OjPuzvcQxLRek0XieDlqf5c10KEf1W5VaSitdo3SHTqxQR1wnzQra
f8/TMyl07JX4gCVwNACW0VNGkX8RsfRCjOe8KqEiQuGliqZn1bjerEslwULQKL4pQB3rQSMCPjJ1
gqy4Z2HfacmtsFdVH5mbO3IlpjOPRZGfm1i6HyqkoXLe4wHiXoKgKqBfF4CIPBj5V8psICjK2zPj
/jQVU2hyrdCtM9GHu5JxJklwWZxMEPBpv53QHxIftjz+dz1OMIJOoGuWeuhpGLjE8DKz+BAHlAeR
Ezl2Vgv77RdaZo98lEUE07+mszxELY01pAReGchXiZwCCPgT3Yg4meInN73e0cMYnopOLc5DsVR1
HuzYGHkeBtFh/ZHJjuefce4MW8EimENO8bdEMCTpw5bn/8eblbmuRXLSoEwaAYJ6EhPAnRKyhdM+
LpinUc8RJpf09UwE1ZfYLci5ayEkqitDVq/ZkRlKe6/gGRhRfGCthm+LFnSSQvY8RIz7s7u5za7y
PPfdOYXZoVrPknK1aMNmVLKAzPq6oWyZ1L0QcPzarxHpVavWn2FTCHyb3vOMsa3B0kUXED7kdI13
v3hHwqOvYbn1y9/8jo8pdcfuZxHv1VBsJY2I3Bu19YMZ7fKi7UrhVgEiHNu7OG5ueuFXDgXpVL2Y
hlSHOI3eRwHZLwIDlkGz1aV6/2mHELmZVzcWnGaw7WanvrSAkYtFA4bgKWioabfWxv4q4f52Anpb
RhLAv6Y5pdVbdkOM159hNvyH9Nji/PhyxQPZpgvMoo5WkL3fL+KJwiyynSc793UZBwcH2RdTIVY4
QP1lclOBUlEzubPGg/SMn4wNpfpA6TdzQKg1b+HBBtdTEYJZCqaKbMddnn7ogwAbYFP9cgTOU4c+
g0r3mQ23IKJ/5nmpqxQZkKmp3artMl79eQPe+T9WP2ao8m/Ak2/IAeqlJ15DiHb6Zljc3aXkfYrc
010MqPbl1yW/SkrT4qWm0qCeb+EdmBup7SaTonrS9HawafgRe9yaE06jZs+m6R8+e2iSx6tbRSKU
yyh48RCZTW1OXXJLDFS5SgnRiuvGIA1BlAbrL1Ud91aWsPMQwo6+FW1LYi1ad0xvddi7t1odO7wx
1gTCNp0AFamndWxQ+WSdAdWoCy7NFTpTkQCpINT3kMVbkU8D/npRuPjJow/1Vx018FKfoyS33Uh+
7u8vR5ZB3zlvOHCiC9yHwwDKmIPBW+g/AWsOeFDdtLe7bfVaNlTjEf63y+KRloZ/o5wqvP2QSwdw
NUAUnAcIgyyesu1V8bkw/0LtC3KW3ZTL1cuqwXcegeZZ0tOP8U95gnC+YC16PzwRGWslB77dDwEh
jOqCLlKwVY+kzz8qtZssEpzv7RLh1rv6dmxQV5E6zrem7Hf3GYCh6vSGD4ZlFbAdkW4RAHTOaYF0
6XkaIeJekE0wot4Ghw8alWhBBKfNXMMx3stcgfHzNS1K+6BP+IGFcWUOHHaIrHmmGcnrFgLMCHS6
DCGhMXHURjqqydduUS/QPCipZvJ3i+EUU0PZiGnkZsQSLskCykjvFLfJkIm8Vpqm8A7Y8FJli0jU
hiY2Z0cnozrvLhz6UQqpblEQ0sos0Mjeqae+JLQ+HkI/+3po2yyXN9RqKDv8n21eKn+n4XY7KqCK
sodUdEmRCsSzMUOnMy0WXZ3QKua/Gkgxuj/6LtG51K2/VypwE/xjkIo0t68mwGgmAlkHF1b1gCE7
v7l9OwY5pg80j+YFj6egno9ByxSnd094uSGUJ+IiXgYRc2sus6ccqrxx/KbQXH0wjavDX1ZAJXgt
MZFGH6TJHEhn1x4HPXGK44yGR2N0GZZYsDS4jxtbkgUeCkklb8MliUu/eqSDzqqwgD/xcU/UMNL8
ZTm2D/UmOrmQWs70aoNddKnOkr0dYodUrYC9YKjGu4hyeVW6H2fghPLSgNu5xNXkMWF75CYZhM1o
FquvJNigo066JEoMTSn0gfkqInYYd70AdKydzqLzqgylFgcXuF1+NQcvOWdzI6Od2wC1KFQ2zSkJ
3Pja9qKZbU0fK3XMQU7AeDDubbx7LhtShWlEr9F/BbkMtEUUulP0VW5vc4U0QJfB0hzNxnX6Q5ms
aYHm11irYLKDWtIf+/t1KHUqQYf+shvjQBE2hyATvxp08SnZav9Lo6EqDowmF6qjo1tuDd62ydlk
0jyMJ0gky+OX18BymCjra8FInHCELZ1AdleqtEsq9I2q/Aruds0HFa8WbpUEk2n2M98xXr4LC6xn
e6nTW4V8B7SY/5Ep/rJuaNYMrCtAV6KK4R9B8UTP27ASLqHM1NYn9+606J6Q5ScvOLIFwemOQw/p
rDiJ4kSLuuQoGlVrp0IH1oUvWefpvc7b5h4mY8uoRLn6vFg6C7kprM2VCLGP1InUPkIXr5phi6xh
AKimGSEolNMqkGY1N2bNqFApspZ8Rzgped3xR0ftlL4lXC2XDy80QjrfYzdCpxXyv6MmVn72Lin+
DC8dKluZVjITAOIOptupNs43KSqQ+KE6jqhNGlUQrjachJK/c4lLeuEl1zvragFRKG0jXr41lMny
25kWRvptsmn3pGSyUyc8/wPI9fenZZVgDjE50OIPObMZX4tSk2ZQSXCP6gsZBO6WSr26b59PxLP4
RsaBXtqhy6Ums5vNpvRzRleVTC+PLC8Ddw+vtUuzJ/k/VJyQBJrc4FyKC7YkUIZKWYCX6iZMlZuF
KqaJ1zx66qx/Tvk1Z15rVlAFwbMtA++kkD3UYCp3gqGk46xq6JhNX44tdxg+3PoMgLPhPA5YCDgv
6vWT4P0TkNZpTx8ZeBAKtRz/qp5GMi56Y/MnOzMz4T7KzOSj4/ZzZJuG22Et8GPEv3jQoW4QyW1B
pI4reA7d+1JPtHw98aR8PqdxSC8QKR1ugjBc0sZSixCYrgnFrfby3ufTtF+ezU5TwPkBHvC3n2Kn
VeZMUfsMTV3bYZ09dSR/5F7AijInZiLWIFfBfraESc9HPk26oG/B7x1jIHOtyUd8CIUmXeVA5ed5
P2TRYdQw1VQRzG8SK/UYfwFnxluEsmELuOTC5UkBHZoyOQY/DMezahYpaCPqji1v5kKT7qb8sfwt
r6cxr0xEvkj/B5CLpbqvnwEbM/FSme4CSLHMNglFy8yXSF3EU9pPTypiaKlrailgCDlMFqDOVL7t
3iDkjm0D0al6rgTLc1E7TNJ/hq/0pCWdQSAQx+pZM6P1wbIY9d91RzxzZWV6BZYOH5nAYkJsTuU5
ltrN8W0NDDraXWg48r2CGrrohuFvtvStjlvT1hNLf14HF0djjeLVjmNZoa0UtAjgBQ9UFnNyeZgn
Lv4TBJAzASK3ImsBudazBJNfsqRn22UcQscGapW5Brszk9BWaudeI5PL745DXC5ZNNfS+754CyTg
iEOOBCLV8dCXsuM0ndLhwimr4HMfV8Xv8esyED73a7I8LjP4syFtSdErP7ryOsX7QwGJYLAKkDg6
XUmcywTSECsxmMslYv+my/+Im2JoOJBVHhN6S1KlMm84DITH4ErCromhIKRVgfbHrmYzLWt7JblH
vv84MlMfJRb6NZHkYha3lp7izddJGNffrG0en9N/d0VolHrMeKPbFmvYasrIqw6FRQkvgoYu7WjY
PWzvJgazFiDaAqnVVjai/Ud69HB3u++nLkxKN2Q8wGoY4VqVQ5Sj3QeJ6F1a6+vD4i8gl14Hrp/X
iY4x2lIsK3/HXquq+xJOLoIxRS7PsJOQaslYvEJDb9RpraK5vrEUAisQS354uUZvHraqclOnN9Vo
fFeG6xOEZHfDuhp8ScknEZc23o/WcwW3sH4zLHmiChzyEhQQ3+9ceNOhL39y7V0LeWVdkcGfl+0j
Az4UfGV3TA7qhT/GhYdtxmh732DBoEAAZs+sts8iVr6T8F2dnO0LsWqP2orf0xV+Ni5E9xM6RXAm
FyiJDIuVzhSi0nSDe0dAVqgfOGtnrEieU/QoV5RfZoWo0yHgElQepsUvbRc5PBoS426eRLbHef7h
P6BbQCWxRol1L+aEzLrFjaFgdIUesGJB9WlzMLQCCVST1VasGYYloEJEiSA/ioKNDZge3gGL3FCJ
bO9PrksKLVRoLITr+vbrh/MIyzFM1C+wYvNTQkaASsxO5nHeTgey4ZGFiEBsgFGceR3OegUZbkUy
Xvwr2qRZ7eAUKllvRG50XMqjXJreeC1npidG6FZ+k9D0NXpLk6zNiBghf70+VD64hnHHWbewtuZ3
/o6xbQJjuFVQuLRBit2AbdY14TDb+trchaeN1gSqFkRsFLFYn522pQ4FjzEBJDrVtBPq+GlqRQX/
LYAiLylNm8DVsLhweXgNmm+gaLFNWrpoasL8Yqlw0NQS2Lf8NOUbv7pgbM7LijmRMw0A/n+33EuB
HrSnU/OO712H2uM2eD1KEDKUfhTWXsdAsbG6lBskV2mn8t4nYcqrYxi1BMzzuaRQUfKZTqC2moFV
Low1tLFe0d9VzQU5R/tD75WR74MYwIEyUqpTSsPAyh5HAyKsac6QzpT32BHXygETvHtjbfmlWlG6
9yLWBVgstnyQKRYYu30vN4/TpigG59euWNzEIIEnugstljceJqQEP8iNoKr9bYH9jniJbqQFXy5/
gToSPQ9WFYrg4bUwK3u1PU2pCkD/RI4BtXbGde6sZbRHVebwvQDtRSmyGBZ24gyJyEMvnszIbeUU
Ngkx65o3aaU/7A0u3f+mRWR9nWdCsKWiOsjFGyxyy7v2wFto99naqkvvHj0j0XEDGyi3obu4XxMr
DI3ZQHU6y1koKPi76GRCsBqjtlwyA6Ts+cpYH8lzGTofiStZ4Mqtbyoyjzz4l4OilET+XpzHK78J
y6KmRA9b4sUh9X2RUfQSed+n7XRpY1igtRThArBQS/LZIrm72xpa5bm42/N6ADeoLWXUqmCIUlfm
3gZvZ+Mbrk7MOchl1PMcXue5KGaD56j8tlZPqm5x/nzRZ7lh+tFfiqEBNz+C6GE1N5CLY8Fms0lD
wu5VYmhRlHQdfhZMAYmz2iETzdJqHMMC+5RKlUtOZjNF2glHaui3LBHZMMw773zyq0vsUfFcoMeK
X7hxkVN20KAIxn48p9DLy/pfmzHoBxYPvTJvBoBrIHQIrmCZ9kPj6Y336aFQcWFy6rjyJu0PBWZP
wdS83A3BFWYAquNsWRh0Pb5Ctwd28xSK+mQrqec6TUBH+kq1i0P/12+RVwuWDGDWA3gOi6bFqhui
Nlb2t+J8OhYGMiMqzCUb9kpl0ABsjA4cX1RhMBrC6we5GvTGRgcYHVSHO8BMy1PiTvhlyBwksSdW
XRwg2R7FONZ0j26oo9N36GxbuoW2B70T2CnAp5DXP4L1kgHKwvwLbkarZjeJdqn8iLslTLR706it
ISh8SSuzbbBihbG7xuoMFRo31ffhnKrhyW6ZDjT4/XUHZioOgeDffG/Q5zeV0EQ3sN94Z0r1MoPw
qNu4BItM4BXJLAa3asffdISf/8xF7tTIivf2PtTnxj3awqQbVOqPvTMXYFm/PT3uLwbp4SdoHYBa
cdl7RzHsVMOyoIXHB7QV38auoKwX0XfSQRls/5+gePUT9rSrsotANsC7rjpWwJhbQCGcJVC7mGWk
KuLTBhqvM2lK0WKMO5m4B0tAh2WRrwOXrUIh3tyokhR0whQOFTlRC5/SdEXLmhlk6E7W3nJsrS2B
70DCZU/nVc4cag88aqZKHUHGGp7B/2FxCf/35bzdXzTCnTlUpSa0IhiqoK32hInj1fmgTECtZTp8
ahl1h9OWJqJabF1cOUynJ7zz5OyjbtSMl9bV4xtey0HLNXR+3UCBDaOmNKQGHPx8HA7mNOBhtFbq
6GYgTZPMmsx8HMgDWIGgD2pCKhd3BHOEP2UIfFbQbrOl81Ab20y5UcYawd6Cy9KEIlhhnCjkd4iW
JiLUlZ4iRPMNT+DAnCATYDNOpCZcpmDTtRB/x0e4inwOMmI9XO6g8RkdHiDgY/eVgKjvpk37V0gu
/sqXJ3dDUOEoTACJSFdlhB+f0ZSRQ//s45Ewhk5OUeS5CCprxyOzb07VNt5O9HQWBet5r2kM4Jmf
59I2y2U+o458EBCT9FT9jJ9hQvTg/omEDNUbwi7tTIw9a5ML8RvfJCLxjMpMytZRvHPU8U2WUsK6
kBlZV24OMmmZOfeveA+V/NeZxAk6qsXWt5gK7ZT4/ZdcTU+UKrvN3tSDXmnfPllisK4XZZmWasO0
47O3O8Q+TH8sDx6+KqYfphifkaJm2j7DjjXGDx2KkmrxbbVZoyV8XgSNGnQY/XBrx8p0+3zNhs/k
a5ORWsJZNdDEkky3PbdB328Dz0mVtigoiXMwS58l3wiZ87w6HjwBfYfkScU792YkuJrcQZzhIqoM
ZAXk7cRpDpPUPr9EhKdnapkeyoNBCz/P4f7zdD0FMbkb/EhS5bDrmB5LHCupuZ5WXE4Hi1C+svZn
iz2nJarBzqEB3CBuXia26FTzseVmnslu4OjPogGyAo5iuQZy0XT4hoMbK2gFFHdSVLWxtxxEQaJt
8bQZ8IdTL3SXlqMevdTgQRyK5PKQR3RgzKn/LCimkPtuGu/WMwqNnkkvJ+0myy75JAs14iJdF1TN
6X1L3t/0Wsx4iqP13rue3aY53JMKXgT/wdoMm4hAvLX1hOyEqDtJIYnFz3A5hdBx/nyNz09vKK6E
6/asz0Xz7SQPKDOOmz10Tc32VgnfUJb75CNr+nOBZVq5oF4LMzL1AFDAZDE0G8NUqZUCXN0uw26O
AkAWico1x0qKJ7y8xGPk9dndAL1zbJ+mHPkE7jdexs2GU7j039JJt/BtdS4YJAhHOyS2hSR612ds
Nz+7P3kp1VWTlNyk82YkZ9xrcFu3bJIIYpHee4U5O4eOQQiTsfJEh0cDlF24HPZdg22PYmc0yz+f
DhPbGhW68Ixk3QnlD7yJ9QuDTm/wcDYNn7nYpbaWJJ0AY3Vjov2KvvXLKJ/LTF1VtRGaMbaF/XKi
FjRyu1Rt2eoWrTABG3ElcKmZjkyTetO0CynIj54oFo3m+qVaM4IzYkrmO0T2nWc8bPqG/UTNg/YB
joePlCw6bo9bDN/EpK8LQrn0FmR7rASWhuYvtZjLDo0ZAfpTkrzzZ760i9mw15BUxb0Cwam3WH99
SYZOWipYSAtFJ88eEd5LN02lOeBJyCXiL4Rh3NOurL+xXLjZmXQ6sK2d2OBBLPNV6JZg/rDLJT2X
2pRH1E48BCJj2AMBF4Y2miY1bXHeO0wpX/LxoX+6SALZecvG3IYFI9z1DF8Yu5BMehFMvrAhmtHH
un3nEJLuF9dkCUNIi26b3jYo6qb73WuNw6cCnnFOy1zP73rUuBpm/u9vFkMHlk+KNrzlounUrH9K
Hi7zmstdjz5D3/7WDswZ2rfTznRfV2pR76i6TldGU4iIJgP9saPzXXvOFrvjCIMqKAqlF+mv6Ysz
qIbVLP7sO/XDT4VVqmGyxJx6qoaXb5puUbuBcg7UIhTaYEWc+qEdDtm0/ebdng/5Bg+zW3NwoXuD
pRCHLOLCmWDmqF4FxUStHpmmNmWpqmQTzqWlAbMD7B4E7r5XWCMS7XgnWJGUZyg73E6jf+xO0m7W
gSLDvs33+AJDJ4Y8Stv3nM4zYlujUbG7DmhC2olMejEHeSdjmMq9IcrsAGI4BsHySc8qdXiw1Ye/
J756UlvdQ7r/GgUf9pWTaPi9XDVTDnNjQW6YPFwXP12mzq3Z7+4QsmPcyBWEJGmlnJNKKaaT8K0P
omH2fGMT+IO5f6arP+HBd0Knp6aa7yt8Scf+jAP91ybb1qaGXuD/gp3a0PZwlr0KdIRCF6HvL2CP
me4qG0H2RJBkSPexg6KqNL3Ah/KMZ7Px26kY6prhCWQTaU60ML6Vcr2FXKJggS1lekR7OwfYZxU4
83CTJw22Zb3VmOFEoV4HRDkUCVuO+6XUx+mz02Yb8FqVKGsNIQ8Dm48FhaiTg8BlkPfbiziPMmTC
waIBXin1PY/JBUyZkpe2dju7Y/5oCWcaLwzZDYpv86dl0y6hHE5LH5io/C3j0WDdpy4QZXeVmCOL
rTQm+a0ySzGNG04s1DDVGFa63pVGXifPnDYqaC5LvMrNZXavuAPaDKPaUsjr0Fif5Bi3Q4E2H6S4
XsqrSnwNVVognLx3pjKHJF+XgniuAjzega4zCOg9jHacwfAzsTXeMydg4uxey0wcWhwm/rOC6tUw
irCgqV792M/ujNsth6LAuJEq/eRZ11ZBLVYIY9RYN7Vj/hsEWOZLkpWAp1h/Fj2+WywmI8lJ2hN8
nH+KMWitf2RYgZgyAlElrLuvzERk0A8iqjyYBkGc6UQyTCu60LsZxo8NykF8vdhkIwco6jX8uEUo
4FeiSi/Ia+5XFHVvv0/xvIm+o8AO6+bS/dVwHdPFMoZ7bjRub1qPIukbXJoMk3SFDDuWzwaIUZjW
2rpYZ7Tmsb3em1xfGZQkCioAlIoReZALeSIwGID+soAceC1+6/skSxTJ1fz41tReGj1ic5L1UuKC
fKfjSYL0pyx9I5tCw5Tg5Tjzx3+kAQdsEVJlxyjczb6s+pS+sKsNtYs+y1pCioIc8UQDEo5m2q8X
74cfPu8kdjrFrsqH0vVOK6y6nrOdWEbs1ne4+cW74MzmKwfwKsqkpdHY7WMrhNmu76WfwVOX0N66
Nf7slZWe224qKTUqLU9UNY69ld7jCPyDar+pJ9uhEGv5ASVE+EDFhlOUjfqSdNa3q5IYNJbm/5MB
CGSkvxLNO99Cxuopn+xPANikGGGpXXpr8afZg2J3cK0HaVwtxHb+AEAfwcgHE1okyKWKjuT/jq88
cp63Nrw0wqLHZF58OmOIsEe/v48JMWOB7M8j2z1ZOUJbLJ48Uj8v9yfLFZTQI5FRespltwqr4w4I
VtSuI7VGq5zCmSLVOZmeT0BgWWO9v22rHsXIjYsQ9gr1fccG7/yhjlKtu4Nv8hf3LqhTzq8YdJGK
NQ584d3OI1bxJy9KCi1I5nog7+sStXi6vhFtzmzEQT7wjwRNMGKxKecFNaAurGgwbpVch69+v3CG
ikB2G7mK45cVIECr6PCmClDeFM2Wjmgt6cWilQ041sP74kFpSszeG3Za/tJE204+n7vDDrWAwTuU
5BZ3Blo4J1BizFzwrA92PBtE2LY18xoXHXwzKpDncCisTyYx4xAYRfyBDZGxg1H3F7teD41C1zeO
/lSiWdX69elp33GRUg4hUe71IB0XL+RTyPof7pDoSdwFbB8t0dWcw50uAqUnqFgqW7adoPni117k
iv/NvgUW1K0yxu/ZG1QJ1l7GysTNz+TlFWJtCCR3/0amCYw4CklMuWUMKjJ3DZ7xdp2/2dQIalao
I7Lh3Z1c38q5X01fmxEFNC2ZMFxUlYmhEEJEt1mexxmD/JELci6BUBv5RFZ1jFu+femvp1Dje4dL
8XQ45NF4sIUkLoXUjTIa7ZdTMZ5dy+sNCpMIVjiV8Pz0Bl3K//LTn6L1P+5WQX0O3EWD5B/k4O0p
aKtOzvxLw+PnZ0UlAgvwu58oXdgPUHCs7So9YOT0kxXsLEcCH0jhZ8vm4p514mvypDnrQpOsKTTe
6qxpexAtD6JNvU244FSlM72zoUrO4emBKgijdYb7ALeYTUkA8DggcRKVla+N8X6/M3nfy7DINjTD
Esv5gYlIag5jO9/nlVuSdGZw2y365fRjOX2KlSMRJRlhJWlspHleEnWNOhJybsnaVnjbpvoqoFFR
eYNmMMVccbSfvnyqiAKa36VWuxA4ESXdE8LmHUOrlFI6qRJG0c2Tku1cA1s5BZLNAax3XCvlMEMl
O389ANGAh2a3ckG3hb6rW5SN5VmSj2ou8Gw8RSFCF/Yqf4LdmLfcdrqC0Kbrk9Qp2JuPZw75YsqC
lbpp9o64VFrOklF+GPyT9XclQZXyY98NgEvQSyYCSyL4clXumZ2qeGa7CXv08pRv+JOoPMnXxwIr
A/GEHCS8DLDnNxLtvUildUBdFWv5+2lQUBY9SpOIKGh+YfUVP2r+5GjcybZO7p8jfjhrPHR3caPk
lsF7fP9hwXCR1IpfCCn5TcwZMkPmynRVVVDJthIcwP3gobgb1X+ssBvrn0TjreXku/5yCJQX5478
QvOaiJYV8t8eJhp0maE2x3uZF0OWaTct7DPy5ibXc4ZFhe1WN5jRwtUnzPZdz7ate3Yk8cHHArlz
o8a9kNRbfK9sLMdOSaJBDjMfxpFtPYtwwULkQIY7Cw94RvxiwNv1hXK6pmYfg6HsYsbHMF368wPG
SmZV/CuqtrydHM431cGdNn5PW7Gt4SbSO6cObiD8hDaJmTs5XlRNCUxcB8el3LmTj5cWhzAyPdxr
np2eH1k2+qeIDbcQcNpi7iR2mP8xUmctjq/lGWs4JgfZK4wHlwHIV9SEgybv0jyn2hVYOJjLsUUe
PQ1Lo0BKZFP62f0IAEkk6LwCz4cpvb/YIB6GyZ/JeZeFGZsYTdbV+TraRVHmDMuRaOcR8TzoQkFx
CBCm/zFLIpWs0dWBiLNdDb3Ey6PJnJRb5xWJDFrkHEu51bEhjVUDLWr9Et8dMEUo1fP0Fb3vBYg5
FgC6JcvsF2odIM5emhCjNcd8jVj2+1cHGSIbXlD0+2CO7x27EOTv2efzJ1jg9jFQWG15C2Q4+NQo
p7/tTJv6BcomBcFTR/+TSZIPra8LOZx/rXU1vEBP2n6azhE5yfwM/GAGMIW9MId72SInHMwoJxWp
ANfwNCfv22ovWNNbGE40IjV0aCbN9pXNTHYBgYYGxJzTTrzXxbjD9gfqSvLPCppO8l23iCz8gbF8
2k0BaIgq49yYREYbHD4pw6L9c8gl8ndYaSnwLEbgXjy0/DDQO2GI2zY0wtSrt3xlm/fGdQplwLqW
rmX5sQ7/q5fe6wIFDHR86rCaSKTB6TSRGZo/SF/CRWuxH1g2GwAbrxV2oSa7byBZm+7tHFbHFbsP
fpRII8ZnjD0maQrF7hBwfpq9fxF1VYRBNjkuYCMYInoz2lhvPlxgSFeEepDnlRGkC7yFiTPIr2X8
1wU4QpHHXFXGa8qd6TDDk2+GgGfr/t7fyrgjIWs8cW/ZqXjxy7d0xL+GOq2gz7z34nH8kgg+REy9
XjHpZ5t68U/ggAmkTqrmwBaZAzzWDqOOEkxUsX2NIOhBDEup6K2BnlRXUO96dJwQu5g2+H1l+NBh
k1nGNYJLrJm4GHkaof1FejlcTTi0cXTWHQt6mqGF7LMrSQLW0L4or1hUaCJttEWAr4KCXu/7ei9j
uBCBoSSsnZ8sHCDVocHpx4rMJThjNUrnaTYTU3WDThsqRNPUryH0xHP+5578+GrEbQSVEo+eCtjB
ZeHxCNg446V9UT5REjJMP7oX1mtzmQB+ZUavCfQU8YCiTeKVSAqLj+YrZr7DHncHuh3PhDDr7Zmb
nT2amTnRa17KxZokUL46hylGbvp39Ex1vXMA2sztfyucnbUxLYpZpFb4qkDCRJ2newGw7oL2H9z6
PlydZKDcNnr+8/x0oIOPbwFv1u5Mhw81rXwKEkEAQQWkf47xgDYoiMfLp06pFIZEb7Es0SY0ylyF
iKkEs1bAAN8JAOZIuK81xBZ/9yWtPflXFOW7KnE7woQcFBCZ1O5hL/64LX9hc7zGxf79b1RWfwAA
0K+fS5lZYp7LmLhzRGa7RScT1YLg3eHDCyFJwOOjtfww+zJxkzSgeMb8kcCkwGYiaMUYJb5Gbh56
jDfuWm5dtJq8qaPkAfwlvGQj4EoN71dwyCTYe+DIfCylnw6zpIab2bTQPETqV7/+u1aOPLtzr6ZG
tAtRadzW7QPYbAzbBTmoNBJOeivbrOaehUJQBKpZZxbxOWBkJdLwZdD4EfyQNUiOVorKITnrnPtA
Zt99zXqm2Rt/usUV1MyKvDtnu2dxokey/3oP67v933jxS5UmbxRZG/mu1YFpIq4FppyVWLSrW3YM
rpenJXlgM158g+nSK/dXmh54pVWJ/Jez+z+SqswmW7AgBTN5MWyKzMiZAMb60iiofHc+nUftSu9I
1NGuxUDmi0iasROyaI5O4nUauig6wE/svYD/3xsEQz809OveaRzFOtzrRlc2CFmRe9ytkNgDW4No
HjL0a5FF3KC0dAwK48sEkEfe2HErv4egLrb3Uer9GSaStZAlU1J+mc2DbMxggJdCIStFuH+tBlqk
+VvlMITVXk2u069Sclw/Jux7eNIG47axlEpYHNXlNnOKACFP6Kc4FJXiCzLQq5lnSHvyQ4UkhSL/
6HOhKsZkexKH2WCRcokfAcU1OwwHzTnRPAgV4oM+jsooSn7iF6ItQIAumA1Z2Dd+0ZqqsiDCM4OP
i/75TQLQboNuKWIcyTYG8ZW8vIGCZtNyQ66xCiAEg/kz4K7+JrsX6x42uZXFuDSgtlw9QiCKr1FT
/0BZ7IgXTKPNRWCmcp0Ag414I6FhtN5mmxF+vxSTRpdTO+y4TZUqTrrgDRaSE6SBcxCf8fXJAMzK
OZTZTAAhWqSydljhOpDc/ZFLEKs/PxQWPmfy06hg7BAexlSDfH4Q0iQAQUYYQ6FD9mcRVAL6pDaw
KaMycQnAo39zNcunsZy2zQ0yxR4/bcUmLofuarVCw+I6RVxu/c/BGlzJZ85aINnY6FerNjxcMB5Y
iXGoUjADRvKIprT5IJH9rWD8J3kpa1oz3VgTukrpvsll9HHS1EVoitNUBOpjfvnaCRkJceAnF4+v
3InJko6fHdYAUfZvrPWMByAOxW/cDFNdCVJPhFi3U10wgXbEXfKe6nnscw5Ub3H9URh296jsF4nX
CL08H4sSAMBd6AYVLJowyDrNzr1BtfjMOdUuYI0I65DmOMljjM0hhDpD7gnz4daTOM93+KmTpLdR
O0K4xRG6urhcwV+zNzQbAioA1TXd8Wsd6cz6cnOOpeXeYNi00cBVHXNfc0cIaBBhq+Y4m2BGAggj
g1a7FCbmd072X1tAsdgP8RMJkhRE0dEF81d4Cql09+6L2DXlvgVcdF2vv5Yigu+xC15/59SJNi8/
3bDZQXWlvyNaoZD0Kb8EnCmrFlV0223hgu4Vf8MTXA1hdsyuiE/20e4Ryxj1KSTdaPUJ1QyXdKrL
lQMyLGu0FeDvWOyIv+t03oTVUAHKM+bCqrAvE0zZdsiNudQjNzoyOcT60TTvL/g0wWxXL+KNr+tY
8nLTMjNL37AtYwhezLbh6zTPr58t8dTt94PSWCeSg9pUEybAmC7U7fEs6hhqOHFPa+7JoFW6KD6A
oUMxEMr1aZTcoy+sDLXvigUolKeZJFEwZ5iqu1V4S2p8FpYqjycrYae3uOKD2cwghKY5nPXED4ke
0BPT47PXQBL2jzcasLTdXrVDaVC+NjZEhposT5oqjJUT7jGIOQYpndPJ8a8OyNfaDjOv+fw9eIn1
LcVQVkVVQGktb/8qMDt3YUTj/s4jP9XdXiWNsLk3WFvWPVd6ypP7fHqaW8l8t49sYhmMkzJRQVo6
CTVV3lLJOK5t4Z/b2ESRPoYMTZfllExE+BYZkM1FMNLYlAWtGsoKzWaCQ2azzAEeECztd72+sNK6
nTn8U4Q9RK3YdJD8A0T7Gv1/Hy8fcagYVhiBYErXZwsL1wiyty0lsyvMxUyJN5Ds+j23u5k9ozMr
RvJqeaept7adIc8KlCwUnJPFiyljeRijE3lbbm2CpvaY8UD1Mv9ZJap7iYrdXP/qkh+TvyZA/Ekf
jQjblfQA0BJnVxiZfE9JdBnV8Hmp7jAW/VbyXH0T1mLPunSg3m0yZ/J20oaK7zbnHJkJsqJFRw15
f6zAhd1pvIeVUZvtvZXBagY9BijSeH5tzPQTu9PdwNfnsPgSrhQtBSR1tUmjfjavacSuh2v1wC/j
hxSWyQx1gr6D7C5yCZZOp6L69gEYN8/7FhDnKTC5MxnSE/1Vd94oQQ2lFGlP4kRU/+OtqIt7oOI6
FI2zeC5Jlvi7COJFuFB3Nhg7NCrSek4fJ2+7QTV4wsP7mN6B9S+Kh9QvDJFT2TAKkW9cwViZLZ2A
QCwNbBS/cqpQwrAF/yf5rgAloL2jOKPH1+VAVp7GVGixZbshmXaJiZQSl9YjZlWqIvDunUgFMHSc
bwJY18qDucefknIAla2vmJCbDnm+jvldWUatvXj9bf34HZf3l9WR5EINb7VN62VuMRgsmtJxrjGA
TtccD1+svlOhSCW8GMJszZ/KzF4s4Ur10vNhxD9PseFKw76e/iCrSW8mMFYK/qx2VgXxsXn5q+YN
+9SthcE+usW74oKHOq3Vgi2Vu8otwAEtUPVF5YSbUMs9L3T3vwi3FU5wfWhV9G9N8kn7EW4USNpZ
uj2cO9nReOilOHwAMUKVL6nPGxXyGPC66zUnx4pH+8v5WUX9nbdxuais4DBS5OYrnWcn7RRGBx+h
L2YkptQS0AQJTMz1Lex1/8mI7SthOZq/tW9M0HRqRwPF3DOlmtAkWpc6tx6tFu3tAQdSy/t77fZd
8ylaWp8vt2+rhehi/LF0j3Dejqj5SCxy1HZsVpaiIR0rXuUElJAEIM6UMWltDUfKIGveGPn5jyES
Z8Iz7CjPQ8MpI6JP7CzRR/f7ehMuoyBaSu1RoAbo0FITvllFzVUunTDhWHPxXIHUduDNHbJEkxmJ
drsQx4WJNPVvhHVQoDceN1pqUKY3FwFL1RSLt/GgEM9wECZnEvVrgG8G+qv5REj8x+8pHmoZ7FeA
u/d9y/vvvsycPEpBLVWhkyLzBQIo42LRqwS14B+SK9ihmrYMvvmMAgv5F2Up4ccsUoNQlyydPxcK
hFl7XRx3AlasK3+/QSwzfu4JsbNzR24++cGt0TJS4o5fsLnZZJXhba9hqIKVJDTd2NCcpS6EnAvw
H2+WRCawo9MjUMFeArnKy+JItZt/Sm3fdBYpPErHS2+Y3GEF6v0GS1C/7LMeRtdUePUJ/V8U7PN3
0V3KO55GGbRvMhrkG3CNATpsKSuvjqlaJDKA9VIzr3GP2tVd7Wx4O0gHnGKcPLxyIcJXVRmd+68K
qmbXYDbwAcLTaoRuaI+cXijq7DkMGqeSYXJ+on9lruv2Bh/6JC6IuBsXLavGkVSrSUNAg0fQCcfr
lPI+Bnb+dFDc8LcAa/f7j+vjR9V2feS9H3dk8LdGOS+NavVPyoaDHyHdhreXAUFWBDtrxCU1PErH
MNIeIutLximOd31I0+MUBzwPJYUdcxEFKOUgdWC+jgOAxzfVFh5zbbLndBrLDojjs+7TYbVyklMV
hXQdMC7TX6UhlNv6eVd6wPRay3zrb8AZE0UVQQeFg2Z+pK9L637mBSIURFKwP+p5vNZVt4TLU2cF
jFkD7Vl96EfVI6pnRd7NtostK3rmoPnrBSwI8FI+4mGyLkbRBMR16kc8dZoqkX8ZkkWKa5rjXJ+w
d7NK12BJm7FCwDvogL89AEa+u3XaKFfWJ22l4xR+z6uZkPBWYLtpoLdyUGzyyMMg3EdanX2Ou3NE
pH53tn5pF4MdwnAbhF0rDWxSEw5uKGONRN5z6tGtEfg2ztrg/e0Ah0gJfku9uCLy7kXpa19Eo/nL
chmINREfCD10BT/5fCQzx+J1pBGeyxzABFkEeLU1t621AtTSqDLXXZ4RCi3KMR4coPU8mJ0ZHkcI
3ueJoXzP5tj76MVbIIqRQKZUHRTovm2GwbN/v/oVmT7Rp9RsLtrR6V2zJ05CJzudARjGLGHkQ5vP
+GrA49fgthR+LckjEOagWbwi1YXmdqe+JgkEukgRSr0891epEmSTzJu9LZ3KFUddyFyOG2AgFC9P
WAUu6Sinlf7/QBMPKvVCdnsluRMiZHqSB91XTshzRWO9LzIy1/drEdfZHBaJ0FBMJ1whoE/1q0XV
3OmvhAcDPscx5C71TlgeqxgxQRQhRokR6LtnBDAX3fzNS0hkZicQ5jJB9bhs5rdzq43d0topQOGq
+XEbWPuw0PGW5AoQ18djTAbLl0F79TT305dIzf1LrIWchvKpSoYvvU/IKGrGF2ThFXZNvO1PfGKk
WI/3om/PK5jEu2ff2NyKS5FqzrNtH5qyEBLLCxJEyIj1JKkrJCmA4uVy3NH/NBvg79kzYmia5CK6
1Te1YVQAogk7+drtzKpID5tNCi8ebuRBivHiet9sZ+ofrMDSVped2Bc8ir8CXUpNhhOAa1j5OETV
62FrMKpShP2l6wu9BFM5OB7qMr5VcndelFeppH9yQQyUcYzadUSdPt3tynFTIyHXKRvqLYvWtSAH
hYTq4uVw0nhFm+LaEgPiqsWpPRreq+IThaoweJmGCIFHYynu1d5MeuRcW0+Ul6jn903EYA0MHpfN
4TbopNqTRMiLgpJrOYjP+cJ7Eo7u1S9TGjqTZ3KRv4DkolU9kD/a3WAMk9SXJMx4gSICLHnSwuYt
g0SylpZGSyNpBWD4QvIPuCqssMYw4m3GC15rX8x+v9NGu9ug/0vVGQvwqg/lN3kwR/ZRR75AOeCE
2cRwUtOI0VO+WL8Hy1Lvfh9irEgBMXH9u60BeeVbVggVk7sdZckZnY7ASZQ+aWmT0c+uc0mXauaR
qt5HwA7PyyxSYcoZkMR9JGYdziYMDhvpPvemkmH5+xJ6kf7sKC3H+0VXCMlyrIhwNFyGldisAfpY
ayhKr53fJDClJOca4hotnaLTtzVxFfeO0QN906Q3SjeZ+NXU6MGlSygmFwMQv94zfHePZ9XYiz2O
tjFFd7BkJ1BWoz2gDrOf+vWikNbMos82nCAxIQX4qlRRB5gqR5lC1sjDeiQyLIoH3Z2iQ3/kwnPz
AKAWdhyix88ma9Pmh8jTBON0jljodp7S/tBH2oR/kOMrZDz89eGP2/yAIo5ox6K5l0V+65IgExsq
3vpmD77oclaT1l+KpBnz+es66pWFp6d+TfOkq3tQbKOLsDg4UA04NWEOkhE2j4KUtlVIB5nvBq23
Q9/tzcxbq88LcQN9PZQ9jOBNuCaR1ut889HEeTKJB023S+yfbkAgMPZVO/5slZkPMDF3aE5lJ0tk
PXtuc3qj+LQXikK8HvbcqJ4eZ1nOyrOJirzQf6A4b9Cq1GHjlSF9snM+hwQHNVPioEJLvbw/g8dm
Od2+KM7TqsnnVYDX6cLhQZJOL7AZ5ulTVzFuimDg03lXItE0LsLMhB1PLQVvHzE/Rx6bLv7PKOin
Q4nM2hy2D7GWb8zpZphS9Rl/kDWWg+Q1oHmrFbpzqocABgHag32fiELLlJrbiKFEDYkfwOv4gJvq
3v0JAVj6Od/DEuIQdDYMBVZ/+0QH4PkkM7v2VU3eM/nhpQUBkMKDe5bGtGpuGLotpgSM0SuQNCvV
FWMP+n5mxXRnx1CAJFdaqA99pU3QEiZRy8QSrsEb99CdH0iHEgocWQyAWbfBp+eirgazimwmjFG6
QZDO5Qdn8cL9ohgjEt0V4V36PVD9Yc7chTCkrSQnuezWtC89ahMYKxIh3iytrGFMzm+iycB7eyVg
/DIU40Kdlm0AG0QymyqwlgDi+b5IZdctNHcoV/27CSFGzm07njI8zTQ6JVEJH6IxBZFVUqC/BF0T
ky9uycp9IriR3n6Dr4Wo00U0qwTLvT3Q+1f+rdPvqsdNh3MAkhxybaP1SYFWtetT55yE38pAt15b
Bo1d65nzwD0oHjz52inuJCw9AP8GPIJmmBTcXWc7AK+ihzbs5ZUy7sjE6pOcnD8SjG/B9tl1a9Ya
WEDX0JVnHVUunnhthh9Yjmw7pxNnO2irjOiRsPGbVtx0kqFF6IAXqvfQXKCh4avNnNQ9B3SN9b2W
AR4MlCPBRYA54xSTA3a06JBK+a9Q2f7CMv1izSQPMz55C7SQsozH6w96yhUkO72pJ3Iw3T/jezFp
Dc4RqNkFP5+6WoAFdRIegvrYGENmI0uPENFET4DaoFnKY33ZKs9jF+mmVPhzkM+UUDT2QeQe0r2l
8SeiPaR3CJNv6AfXtZTXz4nLVpftPFS0RMG6M9n9ZI15Mnh9k1KLlt8gTWNF8oAayXOwdl3Blz7+
l+TF+/WJqaYRKFmT4XD73VMtopz6O306dXsc4nOX/dWVxB2e3q3+bjbABr1rZVS0VDyAGHREj1yH
p+tL22Yss5aTYmCRgUStpBOuBrZsmAVL9RZuzibq60yWe698tUs0dVmOVThGcASddbbSM3XDK2QU
ATbbBpnTlPYiMAzqInfgji4kgkm3JTvIgNBPQpD2IZVvFvnCVrUdGQsh/AevF4mCGD75ydmGlgPA
dTw2uoH3bNvwECjwtkMP78DS3Bg7qA+O69JbCCbojAzhcBqvZtjDl1a4E0G6ydSdMpMqj25DEkUu
kWqZtscl3bWDbHw3ALdb9OX3qhXoK5MtIJsUftZLqaScVLi5usyPKF5RnC+qMzNdGkRylRirSJne
TyPjgL/RIb6kQnFHCF8qFHbSPb4nN1IsmGFiFj9LVhBs3yfeqrUEHO3uNakPr9ocdLe4cPATWlDV
UhequMAdY2nCRUSTIW3ljKBNTXYcFlMSNwCjeMdkOPf8s+CCwSgzQw+oU3Q4I8EZ86SiNs5FbCJC
fUjF9G9nbg4H2KFl4ypfg3Vqisxyzc+sflJjUUvSYUm23C6pChaaQdVB5SqpzbU+ttIdB/sFACkj
FYnQuGGldtMRf2N6IpWsLJRG6rzkM/3rEGBakIKtKboJXHj2alt3VWVCLV8/mPauAEDLVABww5JY
vPhRf4VIZ9atY/Q2AnfXP8oKYp2qcZamvhX0tC7TcKNmAUWB428QUBMWIruO0dO/ywqotzdJuW3R
6d3nSPy4opoPssYBNd0C8m6H5LQkjqwSUlfPhw7x87dZTenVHoKjpJj/WgVh4/57in+GgC2hKlMI
w6pPyqZgr26HsL15NuKhWuiJm8dvo3hsKsYyaXtD6qJPAY3mN8tNwA9KlOrjdOPUbEWUZSwTZ5zN
lIGPm223mUT6jAl4BmPggYUgsqc0OPrXmlOKKiYxUsiWumWREQnV5RXuqQwsNPCMH8ejDUoCO9Yc
U/YcTaDlXTtmrD8eIadak2OOuYWDUAEjVorEJ5tQZcbnFnCIWbQlyq0S7qtwK5U9pNcjisK6ajbj
TPiplgN1PJa2lsRS1Qs2B57eqS+pgQGZfskIryaVVAeQTPH78n8/N5IriKwW+GDdqtJU2APtTtc6
Qp8kcvGvEVjHd/0pVcQFe81cChHAD2DZaipjO+CDlDfhagTKZLNBBWtPhy6oqg7UOZMwAdT1pGHW
RJo8jAv6orUiWWhpsM7Tu5yeCm9b+bEiQSUQrOS4o++VmXJZof8z7CwUamwYsbXMmeURWpv+gtgY
LGZAtU++ACZUMxqNNuaajs2UR7V0BQzBs/lo03Ty7dVnCqUvY32Sj33Vsf2bknexdAMBe5VE4kUZ
Hn4kD6WSgbzmevnWzXF4uEtzQLImE9uw6cYeMLGZp09UDkq7fCAPOFovzu0ZfdSpahYU49MwjeRL
rp5KkGvKj1MxkxeKmX9zL1Jmd/y6zjBZ+DEn4sAhzfaa2wYoTHZZgzEV9VW17Nyn8Nc+pxDkaFZr
vNGZbgV1T3xQ3n7ncTeh5UgQPj99StsB5Nijts50H2ZXcjSaSK2V5ODBO51S0Rnkx+YAAVYBFQoZ
0dtJ8FQ604ZhHmQhgMQwbnE6/ocT+LNB8Obd/5OZIpVeQeMtNa+YzM6Hlw+FtoiQppc6Ycso2SuK
iRBZ/Qk04EyRE9V1Xc2rlx8awUd4LGHy13Pmnymr2nNO9SncTUXuNmJr0PR2J1OWsx1qxJ7zZSWK
HJ0kkr4pC79aH/rLQNAzXR9ZXGnHqZjjkqmlq2TUsLIrLKe4qoLZEC+l/Tb8WC+L+I+ZbKRu3EV5
VuYt5rsSoZyfZqL2gjZrowVBjB58r2pbP7kEkeZEpDptm+aClA0k+xKUfnY91BOPsd9qvfzul7Vy
/UMvtrqye8zK7UkWlIEZoLnx0oxNeMK3XmuZcXBgPGUhmK/HpTfoKWgm6HN47Q3oSztS3mDxWV73
IDXD7c4if+KYVQVZ3tilPtv2E45X6hoPdQc96nfW1EUKHtPfAQ8N5lJYzYf58Czvv7M/nF3O5Kfz
ZQ69qFbgyNfh45J9xnbLF+vSYhrsaluJk4ytYtS0nJ+JHkawikkekT62LsdSa7BkVOlh0HjiG/+K
LBINksq41F8YmQeY6/rUNbjtmSSDsHRIRCGahK156Wl9B7aZ3TqEn4tgfMx1sscHrauD+dVmzd4y
BpuTlfRdGgnBu2T8mtE0io2Bt0161B1DPETNYHqgM5W/J8o7Nyv53lCWT9KjQcHifdPI89QDEniq
Idav69VmtqqMsuQ1GdxzloatipmDbkykL9phkiP5ve56FxlO7yLQRa5oqwwD6EMn/bc/6wHb28Sb
EQJ/b9qVe15rTPw9xbrM0xn0f0J+YazzCk69irf3FYuhZ+q/31uoUWFbLBrevGkbobOU6KFzEBoo
SwSwMY9gM8BRLSR60PI3aUTd3jDa+T0FVSJtamrsOwbVuSFl/rStax1IvSdoF0B8iDlLpp8w8nSd
dRM+jscBDaSLur4prm9XB3UdG9n5mEMCPize3t/RV6aFF9cuzjy0BNaPlFgY9EzJEfc4CFQGmEFi
1Had5hlUnVPQzXjhPAeoeh24SWAwTQhGL9EQSZckGFAK8d7xpPZqlWIK2D5VnqZExyVRHgeEu+gF
pXKvm+O2uim6DN4Xnsj1Hk49iAd4WH7rCrQhks9bzjTkvC7JIy5ay9JLm9eRNXWhaIlh6aWUG96E
GxQ3Lfdr3bGON9aXorOs66DLV0sVNlm740Msp8yOKMq5IjKqPS1Y/BfeN2Yv4paLela5VNATgpVm
m4Hl+4aJVRVaPER/MojOZD1hDqVeFAfGr61fvEOxe8fTnoRbs0v0GN929e5NVpZkznmtYbNelbqZ
4RCUMTk8N6r3hs9jjTEgHvM11tajUcLnn1zRbtvJBgJl2ePkoUSwSbqHk9QRw1ku9Q1zfcdo6Pzo
4s/Iv2+FXVtqY8NJSYk9SHXC3pPATAiRsSu0MtcY3ifBGOKi0dbD4auwNjWIhpWqmhA8ZtMTfThh
bbtf/9u7UcyzobSU4MAsK4utruPBu+Ovd74dXhoWTnF2uY1rxzCm7AaFUiv3tzj9Uf8c5da84HG6
TGHJh1yUun81YgX/2eGMkKOtyoAeX/75p8knIfdBCifiPAyKdbdXI680LT5oQdIF4gHHGdB7lTH4
MQ/E+nnCOaKO15LlGe1qorsYE8BuIYEHC1w1eInHFYzsaAh3bSX/yjVZdKDZTHweUhLR5ZII7k6T
SAK9Nqe/2hUIY/B/MdgJMM7meu76Sw1LAj5sgOIAgWCRpVl0I3kyFMDYcbUamelKiD7Ul2dno//V
wCUvzbOG0FkS/qC7BWrCk4/CtPOd2FASu0wvMsiy9MpxwrKRG8Cm9kCzbRd2GU8+cigeqsmAd9Kj
OcApJsrRTxWbr+QUX6QwkmIEhgnG4aEpu6uBlinEcIa/9qupeK/NBx6zTp+hIW0dQJjL2UmqzMwZ
jbYn3dtDxGKMGm+eMUk74BY8apP2gscj/S6+lFV+U5utzPKeLam+be7psGZa8Qa1ivO6nYeLZTB1
nTtZx2ZgoLIN/cw5pcdqYae6+KWdmVb2ErD1dh/GRN2BOWiXGAIE0n//6tQW9ohm/blNO6ujdgPS
jMToZLke+G5/LoGIbLmn7LM9HIttA43tV1gIsVNCNfV3CKnRqDpk2LV3lVAaRCt9BAnhT5zAMpx5
9dO53b0L/bZSPsnKXxcokWwFMfyzWuQ2wCsg0g8sO24lsX/kxBRmpRhHjOzL3sAqXF3NgKazTGuT
zeeJv/mlm0XewDU4Xlrthjzv+P7cSaB8g4Vd6NptOin2dh7SewNGnDwiBzQELAYrrFfUn1P/NJRz
qS8HJNkdgLY6bXnofPve2ySwcc5L3aPPcJkheisOwsingWQpJfdncbnShnv5NJrg+2gU3gJs/qjv
mQQdCXVoUBk2oqmuHqf0xgsK5x5AA6Jhkdpkf8NSCvzjcOX21ui+z5YTalcn7cBN3nRK7w5yCLQf
OjdRX7+wXPYZU4RjsuIl1XDhldEQd2InHVeoTn9PKW8bPgc/Vz086/Nw82d2+6xIowA8IVYr95VR
MovHNXxXqYuts4JZxiacFRgV6z+hqW8NlX2NQvjWbfeh22owBvbJLSymcem/V64/gYIKCMFElt39
6OyS054bEbjUp0C6No3KKW+aB+6Do6ufSCW2HLvBHJyB/zX1WhKTEWVe7yhPOpqEa7qJfp17U79V
1cNsNZ2vdlbqVp/Ht3dtV0JtNq1Ai44IPEM4z0/TQktsqfG3bzQ88WB42LdLfoxmX+UTPUw3x3x0
ko2RTJ8xKUhGBSvMX9gIxJyNmeBjTUGNe9k3qiE5XWE+Sq4pC9D7uWKEEEVkipyatIlScroaxw8p
Kl9Uvu2mWVtSOXKRxCbDBUllX6209DCcVLbg0pr3p+tUFqi/2QG+mUo3EvPiRQTPasGDsdbSllyQ
c23h3p/jouFnNLMxSFVxOXW2zphrRq2m7bNnDdBvxiPUXB11CRYNBd7lnwhzkmL9SvVkd+4tfchH
qEyEeWhHFvb28akXCizPGaoL5x6+8qypfVKNiDxkv8cp/MG0Whjfnbr9qSGHdUgzuSYzFst1QM5v
9QU/pLBzQ/uuxD5JPITgBh2SbEFrrWAE3EDwQoSKqOOaNJqajXP5aiu7ui9R85rQXzRKqfY005QT
OxmR2TU9K4k8ItqwT4WPy4m+L4/nmpeZnX0fMKnNSt18J2tn8L/PcIz3yCaMxAKCLrxeHuPA3aHE
bgPSM1h5Q8P3uyaS9cUPtUIDXHgmXuhXC+87VyMp7gCOX3YYqHbURaZDKQ3DB635SlFggM/2hGrY
5/1qD2uMIJN4+ZrMTgVXy4mVykUSZjlus0M+prAbIx+nHVAMoeEfpdCDUcpDwghApK2jY70blsxA
z46LZ4+/RQKgIR9cJRGdCqCVTIVkgjBkWMxUdd0paqgW7Oq8V6qrvAqSg0E4GMWyf1oq2+nukatt
AiFc/xQHX3IiByOXzOIk0V01odTPH7DAmgnl/E7C0QpDzof2X2DLSXWXprDIEaC03DXoWoMtf5SC
jtGCl1Vq9QQR0FLppbJRYTh0IrSiwxrcg6vGSls5rN7l1TzxUSlgBGXRwkQM2OQRyc9ThBGMqvqo
4yW7GlDMxtC3riwjxSdZPEXGXmUEUAxP9/bkMgkHVS7Abg/y5J+mZGxPo+WsYeZbXSRLBEp6pkN7
e9gmYpSuritxZXll1eN8CblZHf4Zfc/K9ATFpf90vLrNlf641ILDOR9aIIJSqxLJ0EuzsGuo/IKw
/htu221CW/pFX5klkLyajIa3DgqJcPMOjyUYqiw9JQqt3P9xe4MzRRexfikKR8sydu1EjigTT1um
y1eSsBQNGngF6B/vqgWFhu8cFam/WFpn8tTs1yzLlNwK+17N4PRuNAcQHjzYekaXhZc4ht9UP0WF
yN5KggIJLRUxrmd66LfxspFbzcPm1ydLwDaRatuVvJ7ToMa9sMJSjZ3icId9YnEI68/y/n7YIWYT
Fo49tydOeqc4vVYN2emo4nXT3ASoUD1u0nUK71HwmvPy8Uh1jAaR3fvhe5s+pgWFadmHU1tqK+wA
1m/uECaNJqtp0QTYX2sbJ3/UtcsEEc8xUyOu6i1u6+0seagDzgeAaSGBjElnISYqE89eci6/RtyZ
GNtzYeG+i3lwSKcA7n3N4cQsvsWK3teb1B1YsVxZLMFF3YI+HD6uOArciVOJD3LlR/JmALLuOdFl
O3C1lq0yGzYLoD3BhmCcvR8KAP5KFy9rHAMkw65z4n+Q5TfXAIRM9smfYo0rIHvns9mnqzIG/sGx
HUIPgbCBkUG6zV6xIFFDscDixakUc56x7xkFPoSkkc5waqnrZ9aRAWlXYLaiFlyRgaVDfREzm75l
1FHCjDNRWqJkeiPWd3t3M7NdOuTXEgfCWQ5XM4pEqUmmcqd6XjdShqaQuSepy2i79rPKhINMMpJp
ydvtUOVM04WXPHIX5i5gXfRyBCs4vU0gd2hBwmQt40t1DMhZcP96wTrKOAlGoV+MZWywGzxFhMUT
QW7i4VMXg+Rk7gD954n0LuAwGmulcFymb2l5p8pFKVluK58lrWSczdrFioDJiien7zJYEQgO0En8
6PBwRSdcoVLmqZS/C6OoKBeW6u0VxQ39NVOxvRp+l52DpwJTAYZSoX/EJIgGM3/MdUkEEgV6yh3a
z6MZIV8RlmUFsCeiQSeUkWazCUf7tGta/4QO/FVg4fkHobg2xlYLCPabfv8z8W4xmu3KHPO1ZCSj
96zzhJAK9edIxGGe3cRH0RCGusPx17/HhaeCi17cTBi1HjzwXxtkptPyM42aAyOfy7XTb8LJJUHk
XxrBKE+eoiDewoga7RXbCcpOdqBCYzHgg+BP9gaVgWXzDe93nKO+QRYn04aaBwJFKWLGiypn8zom
zRQQ8Sj9wSQQYZd/SDtEtsV6IkISrvTQQWnJloIn6jaiUdmZTcX03JrBYRuqGliE5RfgpLOHCRsj
KLoUQhEcXF7aOj5R39js7AyWE4Yi5swv09b95t4mKlloX5NQOsJOycjina0Asr5mUEO9PhHTp4RD
Td2BQOIhezODdO7mbSnwcoTV8ujKdRdPEBsHg0Fo/j3j4iuSF/3tdlCLfhS5qQjnbcZhN87XO6/K
RZABVB1mwxB6TifqFGRPCsGvfjjdBBgKgleoLIHHTIAyLFgklgBbcn9A2vnwtjUQRs8OEWn+z4+w
Gg+qzwQBBBf6qGj8T7AaHO5sZCI2Xpgpaxzx6gZCyphELgDikYby/9JWyJZWMeCiPcn2ljcXzRYh
Ba4CsCHhRV+UrgBQ3dClxDm2/9TpISyj3Ab9oHlSLHEJ7cOEQkja4XGkINL/a7m72/6PYcsN6u71
VIuSqcG4vc5N+cEoEJVm+9gWMWceuatxRpARPfoJjZGosseR+ds7loLq1esvlzaPzZ+isgjF2sKg
lJyTeo/5cvvloGtXnUvwJJWby2stKnMn5Y+9NbyenaP8Eg0XaKoD5sSym/f5ovRz4wAoKmyuPtAt
ugEEaan1nViQhTJPP8K1P0bi1mv6cGrDPN3LTnI+MIPA9jfuZcgW9YaYJrsL2QOdIZewe7h7FoZV
5/IYQPUjrG+T0K0MooL7+vIsMCsMmkQqkSp6aU95igOcUj/9h8lZxIlEj4dYds35fiq8lPkkXaPG
TyBADB0phEFWmYqQI84VMcA4HiLjNvBFCvgHMK6MWrccitNDs/7FleaJxm64NuSLWEVpcRWTnnqX
A4dqD5/oNoi4dOVJNjAFWcYrG75me7K0ca4cNp8uAeDBsnKVDf+A7lpl/b2GC/Hs4TT7aF0sAZlp
PlGjqS/tB0IkunhAc0zkNc0Kiz+9JcDr7r2lP7/LLgfJnX6nzm8gF3A/E5S6lCHlgSUbUz2XNUUv
i3DmvidH6pZZAlk92Y4SmSqucnSKsETESml9DTXajiBElnaDtc4xxjNRsdth/5ej3peH+FEv/HdC
cRPlkTp5tygMos4aS5E4l11BozCUPiHu8cGqoR2UpHb9vhXirL7fQDqx/7J9/tWydSYan39ctjsU
RDC3WxxzIwxJog59E1DB8nhdNeGzX3DuWhUDEQTQwBWBdlCwi7wwczZMsYGc2rlNvccQcKJWDjOm
k0KkmRMUU3oAS/d9oWTsOTUcQQBPZ7+c/dnJRV9Gh6Wt2aX1O15IGc9UZXjwI90kQYtn7abRZl4F
M1fXXUC9UMmSn9aJhufN1dtxa5IwbvHE+c6gr/EupDy5yrINtxp+JTBf8bW+NvOyi2wD5U6auBM5
GDl4VPj2UY+6lDuZomOK3KscnrbMix1nN02kcT4v5ys/h2GRu/B0pOFCQnwq88IfcTeGJtCq3cEg
H62YDBade9zup1JjPmRg6Y5DMs67iJTXbeH7bLzPLd9dOhfcPveLXmClcojlT/noy1iSY1swO4dm
YCa8Ls5H792NJWShJZg9AoKlsi50jYLNskQjZ2U3wAIFpaxZByq3EiIx2WlyRpg1XESyLHN8Grr0
7ey386irUBDm2meaS2QiXL71op1cviEiJsiWCliEgHAWQsa19lvSEqjRyIhd6OkJlXhKSjhqI8Jk
+Ot7zqbLNrC6rho2y4IGdVFXmrFbOkFksKX2IFSiXy/KEMeK9dinfdRbjnqbNJFcC1R1oBMaVI8R
1q1pUVOLg/FTEhV0sfqrBR+Jpb6RwNc2J6HK2ZSyTAKJcKspgKMlh3RROZDuCRo2VVLWTHcIpj8T
AEc/R3HrIXNaGa/6Y/WlVUSaDGfImk5Fuov8qRQJuWfBSUVxh7WHscau0UboBnljh2UlQrfFkPQ7
zZXkcHDEPoTxAOT083I29kqCKw0vt+lK3s/sNpJBWFHuhyH1s9yYw6p3ZEB6Ymgf6MfxWFPRrg23
/VD5T/YwEfI7+c2eTgPcQHZYIQLQ8ZI9we4mZwRSdKgsqg3f6GDDAN+aOtWJqwLwQAI4ZGwkPBsB
KVyLYl1RgJaNFs5p705XiBI14IUxZgqdjQf/Q5OW+XzZYLNzb+ND5wcMNbth8BWkMLtzqEnSqLMi
vziJueT5Ygs1rFawx79E0La99DxZzq5uItX+uwlL75954oTvLf3FOOZu9ipMm7AqmhYKCoXyoj58
oYx/Tso0968xPqNl2+JUL3tV7fGrW35TI6X2NNopPJ5aTl7uhl/UvLKBGzYKQTyiXyKxKJD7D5eP
znVW40cDe3kSd3UTnoRMXsXyWaDzBTSZVLNjJ6SoErPriKHNuVYkBzSVx+SoPPukLgjfdPCOcK6y
DgDOGVuz7BWJAFvU8fN6j+Hy1H+q/s+2/RGmweDkIAY3GNuGjXRDWKVhP0LVig1Jn2J+AhREbDeP
+SeqHlcGngDi7LUTGwTQy4zcDBIDvA30IzbtJbgdgGgPNuEbvrRkMISUZ1pGKUjVQ3nVN9+MaUYC
NTj6HelDghk57u0JAKPg41UsUnCe1RnvP7DcCqBZiHoernl7GgKYGw1Vq3/vuBEdy0rHDlfRR0mq
TqHVc2WIU6eSfhuiT3WCnGH+8Pw+rcturf/dHwdxBx0LwknuMpe2wiFd/RenblLy8RirAUkLh7lh
KvAPohMWASc3cyKkhAAjRrjZbhaP20BWjacD+7+en3nKZIb7ZtFGv0l0y+Itxn9jsWynwUPHZdSt
H1xDE1nFmcOsWZh4z2huo7Q9Fs4c1LB96KPXRu5bNa6CjgSOaZU5eEyd8rdzoUfm8EnEaO8+WSGL
D47D2OBW14ulTEfq8FiNoKJWONHbRHofGFmFYE25oZ0q7jKw285G0l6qs9QTeqMkvEw/xeyyrbNT
ebIv+KmGFLT7JcffeUYR4XeEEOoaU7+cN704McA7RHGtRFJu65EW6l5jBivqj6xw2tjm6dcR95aE
34UlhpGn8dJMSM2Fn6MvlkY0xPxbZCCkbhWjOvKWGPLM8HtWw+k8R8wPuZSuJsrGIB/Hn30oBtaE
ldeTW7ugOkMyrsXOnr5NOwi8nkunD4OnHunLC/nxYZfLldiClzDvU3Mhr9FE+oDPFD2xfXmiJ5/o
QMQ5/Zl6qEI1TpKQrb08cCNq2FGlziQgv+mvdMipe6ocxgLEpxJz6yzvH7Eb18NtwPr/E8wchr/V
bcHNg6YVxjTRb4CVpurLr/194NXCAZA7NrqSDnrp6BJpDPZzzKt/oMFbzZY0mPI8DDo091knhTmW
dkY77zzN2JsXw71N1gNI1IQPh4xSaFRiGmRhRvj4Pzi7sNoFGUgdEhbDpYqZEXm0smY4TjQtIcp/
2KouihnE+CqvDowt/bQyxe5lXeaCbwYF6uBQpldNkLZTOI2EUUv1J4Rksv+eJHqVkr4bG9OcmNk4
yTk7tKMOhRFheA2NrrdelD2Ew3sEuJKFNksfCqX7TqSNT8+WlpYpA9NHjSEsXFH9hUi/fD4fme6q
POuGP7Rpb9m1xDBWMy+75YXEOCB+wN8MiYqWSUrfyRa0e7mpFT/exoNR5saCuDj6omGkbKhsT1Jw
0gynDoBWzZNMl0Ea3PC+wMJV08w8IRD2igVOvGB4ADMQnYp2w4u+9FLDGF9T+beZ1i3ixZ7YFuSo
OOhMMXQi27brsRmAchXzcRUeBuE9kLHJfyOZh37xIZ3JP4Aycb5qf676mCshhx9V23KqRUecQMFj
1HejPlFy4W9Qkda8E/FEcF5HtOgM2/OsvOmjW64jqep+qUF/TqA/eLn4H2j9yq8oOz0936+7yBtw
u1BABzFIZPigJ9k7cQcHsWGZgEj0W/6S8PkPTA/jkS/1uJ5YlTU/H7FAcOMKEBp/eDXYcKywwdXU
rHj0zXN8DQjNVftoe4vsSh7+4MjOn1W2xrfqo0GtfuGnDjcDXur2m7+4i5iJ1GBJ6RVeU5S3llso
ENq9h7gOTs8jvGs2r16swBmV3gArirnz5+WaQ5w9yC54ZNFU48YBnYmnY/L91FV+7gfYZKQlcS6K
6DRBw2o3oVtqnipdtzfLuccaDH2DRySbCuSiOJ04dh5lTDB+nMREt229/qZHJNSFWlSoUlEItQpB
LWqZ7pe3o5F+w8b82l5cM+rDxRCmZgsw6qqx6sCMIBkZXmE4fSVTHD4WRCz+A8uem9+h8A+2xpPj
nx66JL5qX/MMfLuIyi56Z57a7rLKAcAsiefMBn+UJU6djCsqgX91B1djBQLw9OG0T6fqtqgehfRH
i54HLGQhSydZz2eJzy9/4YDgLSb4BfPeBzyk8bE45dyLXqHMmfrRtqmzN9lLrxPg6ijf57yndTet
lDbaYYCgpPGiQM+25MtPq18ThP89WLZCmCxENtw1oenpRoj/I4BI0Bzi5WMi0q2ytuEGogrHy7me
Bwy7MMsBnTVA0J7/7R2Lquy8oaCAleCkgVm3ohesxhFdAxPPvngndhNb/HzwfB2JDnUJpe0hTlWF
q7jxTUrNDAOYHuVBXsYlA70A7kphxmOcKyZXiHMNj3gVAnBWoo2N6Cn50InACDggUaeK6peOUCvN
QovEVDrJ7tHkvTCIkCVz/DZHUM8wG5z3LPFfiGJBvayWUfwFDNt3ViNMi1j0NqOFq+UX6qUqiC4a
Fn0sio96g3dJnQmo0qT61NmziHXkYHOoIZUb4oveU52FVLJ3tsJOnkbRPjTUReffLm4cIeUhTdOd
HlC7RF0qMsmggZJBsi8FR8JIEMY9deaxI0iSPhiq5VByvlrp/Bw7ZliRrxS/uM2xias7m1S/boJd
GWY5o2gOWMqpl5jUXML93JsEq0DYF4GJMIsCue+lBeOGP6Be0Iw2ri140M7iH763ur/rl6PepkcE
Pb4LoOeipM5EvHMKbaEJi8aolK12wU5I/9sL+XSje2ivz6JbvJ02PrDm2xv5xAUqhulLXerH3ZFs
EoAvO1aLvt3VWo+PrgN6V4n3YQfrqqUdj8mzM7DymkB9foByoUVRGu/DffZpIzZZVdRa4ayM5aIE
bazMbD/04BKPCRzg0aQl8k6VRz24igzaxzZkbVaHX11gCZGsAp3ChTigbaDS6PZ9zQll5KI44VXf
yjEypVnIYzPF3/Acx9061mf3WJMiqV0niuKbH2WWrz0Zjh/hPIVvCcm+ZMT+04KBeY8gAAcqH4n4
vIIC7iH6CSMCuHVV2UzxhG2se4BE+SoD6iJgH708f8zUcskAUeoKvzf0ZCKsVm4YhwwHt6J5Y/19
HRcaU75gJE/JEaq626CKBW5MIf8z2VMLQUwOPY6hKNXXroaEYlbAYNTNbh8lygF5KNOM9KAh4HaX
IaDetCtIJlOH92uOCuDpebncJ0lgrfk7ifbnx8/KX623UB6UkwygxdaE6gBYn5o5M5NTevejxEsm
2hxmaDPROJo28f+4hMap1A/GUhMk/l9C+WxOhUUz1lHLFSifqDlzcew9rdwMHoscyfkO9MLaCr0e
x/xvCehrR13psdsBaM+FKFmRMG3WXurmvjdqhBULlmM6s7dORtgla3VfMsybR3sqiGlfXfkcQLzo
GcNSmfX95ivT+7EU9ZUFhkvQJ7K84bWSkWLAeoGvtlHBplTVm0dW3hg0RfgNyO+6iltyoLzizhQw
n9H/F60f5ATG8RccNKaCmSFDVP2h8R0JuBpxQSIasTJ4r2GjF+HQCJpGYr2WKL0KdfwdGqDQwqvl
CGrx/q4tIw8jNEK8lxdrEf8QGl2Lzrekd1Aewnk9hp/DA+P63A06v1/4Fktojr3IdBXz8yb6Ss/b
XlUMVIQZnlezdJHg0mbGX4OjZVYG0zb+ISCwp6iBSGODqUeXQ5Pl24K/0n8dGgrXkkC4JDf/ioui
kKhPE4e7W8Dt3HHEPYCddt25ZNGlv6IX/XY0oZAFAgSX8k+KBdUdNd+Nu5FjHN4PiCYT7IFRcVrt
o5AES7soo3Ddy9EWVFrWM1EdwJyM82n+fzwFI8Ey3zu0rvY7v0Mfd2zPO4W5ETyRxnkIH7U/0ULt
2rXM1lF7TIFTdU1fF+3PeSaqviYXFUXsIWcFBAoGAl8eM11wCkGNexk51c7KZd1oYG+AKpXlvnfl
dPvObCA4tHSR1RkOpNDyfO+X4W/3A3BF3BCskEIgrret8ihvbyu1fd8kcMDISAbu8iM4r8O+U0zc
Uh1bcR0YtARR1TqJWUN89zZT/IJ8ufWU4m6ZT/GLITIW7WArGjAc21ICJwrOoL2s3CKTlwMffK7q
dme1Cjhs4xIU5RSNXtxmN0eGD/lt4amrQi0IKzS2Q1aHPxTg6i0M/RkUxrvt2fpOWWw0OCqDxr//
aXKh7gqPinzf8OiRLaShxGzKErHZF2mX77BLpypQHihneLbKBz++QWpJd2On9t/92SjDSLCzH9o7
F37+W64gyQKwfEO9GuiDl8WyRMc0Y7ckZdEOCXMj5c6sMOcAnFQqAnt5pvd56TsiOloqB/+Qfo/L
GplxGpSkMQY0goVUSpbCqnSUSaXGUKJadpgtmbf9HEw4tEqWcZE/AWGThKpdfL001fT4XRuXKc4N
Dcp57YO0b8QRjOKDoncxOzhqcMuJvBOQm0NBB/bTUfCpW2asYMAJxt31xnzSRW4s4usar8VCttgB
RU3zk7eSvw/M6SGt/+Urfo23Ge/T+JPWvsTCophyhVgjhzjkbXqnY9zDV1dJDfdsl4yPQQ+ZgwDO
w6rSCr60rYeGKQjx8101cXLRBeIqswikYrCOWLjyOqEDv9oO20ziPltT0easedeE0z53Ad7R21V7
uVSwsygbeuSsQVbE/LzK6pl+Gif+RkoSEyeghZXuHdstbzVh6CCrpovRWvULiMlhiS2p6enPXg//
vyEh570oaKj4hGVgSc2aolZ9VeFiKm8sRaSYJ+B0ZiEei+YDHOcdSTsJ8PYP3j1ONGG8xOpDCY/M
CWzlAABO3fFcx99GSzGpr5WqTTO02lBBo/PIsIvf0NwEn26bGEK2r/s0uuhvmMbcklRU9sFii6N6
D87yqwK8sGKnLKVRLC6HVAGOfIMB0kjuP7INunqgE9+2xD9sTKqHkPcEOvl/hWGE96Vkq5jbShX8
luaJX0w1vZTCDftDUEQhp+SUwVU/XokcAgpv4yJyHn9mn4yzG7Y1mzddJls56uAHMyjthhKPslPI
seaKk5VUj8uO+d81b/lItXYgQ3r4wCgl9zT6uTpmRHerEGtMABFfEHf7Kul+jekm4fyz2ypjWPN3
JBC9NQyMWN8mEDY5ZauMlvJIdQBLrRKR+b4MT3sgH2sCjA3+mhKl5rZu8oKn44TUcrG7iNYg70OV
95l8e2X+jO5mFztyGVd+T6yc08oZKD0yeg90ld+ed9k4Lbz3x+cd6inLzYVXnsqYf5ke9HpHkJyz
47m5ccHDrT3J5Y3XyC9d/0r1L29tzJOHnh5EDWLYD2X8qh+xOlXK+P1YjfLxmXzKxH3rilgIlAPF
BFtpAIlazu17Wt3eBEsGmWGgrqVQ6aJUHgoZ8dYOih6fCU+X9tIdCPzWUIsqXTvOY8AEz+MROVba
HSP3dRp27nExfxJhKoTYhmDeR/C3zt7rVHuKK4+ILpBmXDUaN7K7QTveBXguwhAmhfg6jaCx40zv
78TXnSNXSAH9b8icQ636h6Ss8ucNbsDO37Q5IVWiC2SpGZsZhRPrn5JAh9v/EBQjwiACRirw4eBC
b0NEh7gtIpNG7Y5dTPN+brqCiISi//MrbNx+jGSJQ/toKyc3Iw0tOJBgASGmrQVkGOjmEMCMFOvg
yKeQR4bbLWaWms5s3oYePIgsA+T6e/z1JCKXf8zPejavbiqCEYdiiK3e2KlmDqq3nXyPzW5NSgYA
URw9+K8ukp6qk2Ui5aUHbLYJsxa4H0r7Q5HQM+uLhDCDpk1J85a5+bqfzuP0Fm2YLa0petGQCh8/
u8c+OlRpg0v7ywRypD6YZisvaZ39B1LaVLf0IF9tMoWne++Zb1I8V66WCMzgLtV84QstbxsYQVpg
7kg0o2KBeLw+6yIfICX2kcVHmQQHy+OVtp03+nDbJ6jSdg1YbjKdA8kRY4PvjuZ00IycNEDj/UuR
3101lWlLfCDz7+xi0+mGzpcfpoU74WCWwyzZnOLLPw8//LHB5TQwZCKQKPkBLik+vc/1GdZ3Y0NC
e2b/JfeaYtABVQS8/mQVk2aFrULQwbB63/XmAQKvn1lGmNZTHxYO8KGoXz9Ap0QkpUNl5fUL/HaS
HtACuw9nXWMMxDIrIdbsnCtGP/768cM51YAw+YzOPRzZV/GLi939faEOf9J6jL7BDiUQgev6Cota
IvzLWVq+oHd7Oa6vxku05pqkLSohMC53NKmcgVlczbEHKMIJLsV94kAvDx2wpqeSRlFLaN/csvip
WldorED5hoNJmQeRiKn40GL6OazBC1zNsmhhzc6A5yRwf0FxuHmrJjB/e48wBarxDmKpPQg3B0xb
88ss0VBkd/k90VQ1l9DRu/EzWKMTtUK3GVBw0iWYSOm8DR1fobqA7WWE+uLNWDzU/wSuZrqYaSxT
OexE3uEEz9KJgOsk4h0il4ocgK2Q45pfINF0xf5XRL+lGLCMBLpLEojuWtkLIDLssy4Bz0Gy0ctG
KfZLEQiENEyMIMD7n2sA4rs0WlBlXS0J1m0Y5EBiQYD0nRRsxOq9RhbBz92RFv7H7YDzN7nJzOKH
2lfB8Z7cfFZ5We/fZBzKTyNceG2zz+ppK6Ga9bbwBIGQEW5YLq04V0RuPHv+FksFlYYyLv49aT15
dGa5JFUZLsGrkvK4mQ4+PlI5/tReRk8RsrGvxazSkEK5NqwscAGgP51EbthX+RHwm24/jKsR1SUB
fLGwayFx9aS5hNGAUHwZEV112eEFp7G7t0byuRLH+a9K7qYpHwZAXRaWRrTj1V9X27F5Psvb5dpo
GFDJeiJFybBCtljLSAYUTPYCPbiI1JusYTC4bs0BgxT/hyCqOfQko6eIFM6HnXFJnRb2S3097t3A
44rK+iX/6hZ+PTNAyYkxxtCdDG67iE4mplt67AMSz+LzrjVFPtRDE/KyxggLyqw0LPuYKGPkWW4W
I20Ghi+X90eqiGmtTEzduiHyq8rUCdbZWnpQo+XhH7YD8n5FTDAVykTduvcbXGTQkqUilQyNJurR
K1yewixbsO8n20FkJtgebBL/U7aiqavBp/w2drHg04QYb1jtLpviuxMrZDTNe3BgtVh9Brw2nGWm
Mk2Tr+mQFIIuWd9e81OeXYllJmUf+1TpylXH4E9r7A1fTRNieFdzJdz7+m4rHyge1qC0Q+LypkUk
Yc8FQVTdVj/yY0oEi3tliUN5I6AwPKeCO6PE1hy+3teiAIaqF54BFNMyeXU7pfABHVdZgn6TMAw8
oLokrdOAzp0cGlHY+FXr3Yz7fqYKat3OicNoOLEcDANgdFpF3h0yWxi+1wch3DWSF9OMc5pDf8rA
Xl9v9Ae1GK91IZJylJM/eW9tM/GTUPCH3/+7KTxm7Cob/epbMzMzKkvAsTPymG2TP6ZwIXyFIwEE
uxIWLVj8C1+hMs0eYRJIU1OF66CZu6pYe2mCl/ydi8UYdqsLodwmfG/6cpj/JTxSi2J0I0+8M3Z2
HeESFLshSq9z4SLYHWMydgCq12SHCeEkmp/AEJB4/LV+bv8dzGssITGhkryP92W/aUzgIPp7ZPLG
lgGYBifahq56ovRuaQ4Yx51yNAz5VeD6p1WRKqH4Ct/d0ZO/T/vrWJmvoJIY349gBzULwDC0mLqH
J4cIWRfYjw6p7QhpF8T2+4ALhwRlI8Kdec0kczIY6BN7WkRlnSMiZFXGCYzml7eivFMp6Am8UDP5
xijkCRvbkVgIBMQqrcj9pPolcGXlZ1rMfDGb/ESM90weWmuEB5GLPznp7mOIZwfhPcaRtGn44XNK
XTnOAwjkML6Yjz6nzSnKz/fCpxwJMsTU8hOjq0D+hGex9bkuXSnqgwjXjDDRMjLCRIqJpvxen32B
dUaRTPkU4XHgkugxSEMaU6uE8LUCaaBtTa/0qcDCDf/zyklRelZlEtzIcDxdzoVs1pySSU3lhkMF
/joKsi+1vbhWphsmAxardvqmvh5t6g2LtN0coLG454wTug2z1QzS87ZLgapsWAuPZsHcEjiNTb41
TMFEeIGbT/wJoxnz8r9iPQ53lg3Dy4btxanOWLGjUPTZLGSMwOVFaLYY9T8DVoeAJyBYyf+E12J1
g7hRt4i/8cuSOrBmcCOTOmZ6IQydS2TED9uRG5JmXWnRkzLnnekuMnbn0HzASHsUgxKjSI8unxxw
b3yw36VlzRO+1LaFMolS+2kdfef9iUfVo3Qa9Squ2r2YNBdkLmjZCMZE3ljPvCE3ps446o9CGwV4
qaLvZL1PiKwN6OQXAo1QWzb/9CY3z2Cgvv61WT9cR9AfCr0gOcUBRnAAolWdffe+Xp6rN43qWTv5
4WXEJ8xhA34BRW9zg3HNQQq8UGa0Z0f+usu8chvECqsnFoO6hau2evlzKyCYvagyEJxZUuEZALCR
ju0R9IhivvfRZdTvZYjuPKagQDsO9KjsaamnYNO+nmvv9Gie7PCToe6BI2bvmeYvAMvroAA/LfMc
CTe2Xs/4j89Zhk+HZwPpXgwvlKmPjYpeXz6uBaSf2WAuJyOkTB2c7Rgtf9gUY2vmlM6QHH+YRKye
KiRxu8A2xszNP9h3mxN4yKX9MRxVj8jWXqu9fmFZRskZ3iGL6O/pVJEZDbYvFjnT2GA2/2N+72Ye
YnHJxcYXaeW/wNCF99j9Weq3p06A284UYEjUrFl5dSAHaCot6Ymu2/KQbKjbyTlN5pWceXWhczJ7
IfGdxLHJqNs75v4kvhQl4XzSz5YFWA2sBg37/rCQ7f2yw34+WzvAw9T93fklp2eNoXx9MsesqYSP
o0YJeEyI/9ReOJu9eA4fxoLka4xBUXjZMkPGqiVri1NSW7NJbgfp3z1N+ztlqQ31ao42JbbiamrU
FfoUCwPXTccjEgthW5OUl8P8uSJ5M1zEEL9rOAABE8YCu9YyKFfosmZQSqWSs2+gDJN1hMdi0Jeh
L2CUa3UqWZH8t7jJ6GDkzYd6KMK6AvYK7hxItpQGkrtbpSkWumsTkMAZKMLoGJ6EQoE4uMy67yBn
XyAWwTo1wW17/tF16gAleAbBv1WQKXAsAF3fLkDCvXgNbsuI7mp3JqUYB5Uiip5aUyMtphyw1AEh
XSHVFFiyPHyfTLy1H/fPVyysC15PKL1d2CKZyetkDThkQ1+X6xbvPUPJvCmCoOlLSXpJoH3jTxUe
GMc5AfkuoStFpY/exYcMlO1yoJkJeDdPl6D5OlP5WFRpKsrbfFQlIOHv0tU5wFK0Zc9EQD9nIReN
ccaF0CQViGPVBzCWOqsRQydMIZIMlTkJcodp0SvTIfXjOmNk5en9GbscgFQflMMC7dP0ru3Lb3Rd
c/lUUpwKWjAI8Vmf5Dc8qcFUk9crHxghdrBa2LvyzA2QSUYhPXxhHFgSM4Gawe/ih0HLqL6u/DIS
B3kadmKFZ5NkZYIng5akqYqbj2xNT4Mmq/qh3ru7agkpB+J21sNTK8D9W+7IlJZw+aMJUpcddH4W
fZr78Q9A+lCYqElkJCAKjL7o8DxOh/8jSq9X3gVQvuw6i5OXRGHHFREm8ntOg5TQaC45KNofVFrh
umPGrQlN7aWJi8gIZNPgI3jaa4FYhoBACuE1+3cGYjR9lPLwVm4bxh1rXKLwEDSx0Yl987QJmsnn
t+iN0BBucWLHOSPeAJ6zKjnwqgLKs5CStyFjHasU5VFzHNeQby7KQTRSLHq+0kJxdhjsy0TITlTy
0g5SlKDYRsRqa+G630P/jDY9zQo0iXOfkNPHqBhQM3bILv5NYwmRMn9Gih9gMtVM9Uulh0mrCTnM
/2wxhcZPBWiq4PSlh/xrDtoRJ1jgl1aj8/anu4VJJdcoaHJZL0mEcuZ5zT+KVTvutqWoEVw8FoIp
miXcN3F4VHTguDREY1OkocyWDkZeI2vfAfT56Ae3AkbOIv0fRcFMvyd5DVPXGfrkj9W92i61ATkw
RiWjxsbDcP3sjG8lwQk1Hv6RqWoKajYD7zUS1ZHS0d447iiLPXemM79xdaBPIM7Jn5CNeV0l5aJD
xb10+be21MbC79D0r9zGgU14b3znhacU9FRMTPVK3HOO5V1+N3RpRlQ4Lt+SfYZ7DoTwzwJ+XQco
sBD3DuiryY7P5KQFL3Z1VjlgFQ+tI/hglTiwhoGgInXktTcKoRFCqxMXATSJ2+WUbypCIaa1VcbI
RkGZftmyRtSHGWXo7KOjG+ipDRSWJh818s9y3Dcnm+6HPgtKbrG1tOqB8zaj7U91xsu0Sa/vwFab
dLwkhlk8jbbC0qCGCbfa5NQCY/yVvf3denco/dTYU9SldptlpsEJn8v/70S4edO1qbhCqs0OO9qT
2uHjlqEPbdLW3/LHE8U5OkrtmreZ5D7sWH1A9C1NIZjt5nGS/cDvKy9e2yKp1yy7SWFsLpnib/e7
V8lBipEime3OSvSAbMgcZtfdeG3Ezon/p0FpQ/Kw62DQnhG5P5zy8vg7FTKIz3ueJfn+fHgulFZJ
N0vFB4yrs55yZ2HWND8Q73z65t2qTJIvWGWqaYN4oZN9eGG6wHCrzX1Qsum0OFUCVsrjXS3/EZWi
SkH36ur3PH64Trboh8crfDGueICax1FqyiBUpATS/7a4mlYyPwkPSasucQqIF2oR9OZS2HEANNVc
w7ZizGtZpfJ5e7mVzlFI1Me6CJLZFoV/wtYcpA2H02VSktxkWNQVLNxOUG2sGh4GZEZpb7FlnIFL
HM/hkYvgEeG6kfWp79T44bO09WIo0gjUgEn5Ua0SZtpKCawUmm61FbqZzz6LhW1bMMZIuMHuGTBP
zFFcmOjqUl/A5OL/VsCF7VMViz9Sk5emYptn90YVu1euDdLjHLJZ/w2bV/o0ZYX1kkyDrOjRB0X0
HZxCM7AU26Yl41wGzi5zy0ZqJ8m3FfxGv4p5+mNIWirXt9sC0VnHKSIbxQ2JmIAWAUMz7BPZi7sd
0ql1ODU0c6sS3hRib/SdnTw7j9EO2Os+E9kDZnj9jTmWZKKnshnMWwolqIsGBYgwsGNJu4G1gGwH
zOEhzizkptSy8nFRfV6Jx9yRk1utSSvbWMjaoZHzoaTXXQ3c8UXF0p+eLNx25/p4V5Ce1naJKsyy
3iMyc+qCN4O0KnqK/Ibp13dDoeG7Pbje2+J4+PQ87bj6FgLl34tq9Zd4rE3gqW6vHZ0hRdv+q0HE
2BDGsMyqZrMbFsWm7KEsRSedYM0USjDRlB+s2UWnpkdctvaYkzThNcwy8Kjxu+CGf1V/wYlt9MaU
S4GenlnLcrS1i3yFC/RqnFeX6Ef6PqOdx/Lqr5GYh8qmNd3mqWx7o81mhmfUBOAIrFZslB2bMgHb
J/by5AJeSVZy8h4WZKtkX8XADrt7jll1OpLSVo/iFFrp+mH9J+msrGwW69UeFwNIIDujgZWG6mx/
0Uec0EgRxcFEG0qGx4ppivJ+37LPA4fbNcUEyrkoH+UYoIPVJCqIAS9V9IIeVvc/QDdRfMZkU8ta
xSaLRZX8ovkROJnprLjBjL+RRhP9Hx+qsHXLOgS0dTDD+wHzv3GYXSySNGUX6MRTh+6efVZ1ZcPg
3EfFlJehcHs83eb0kQdMK2okVVOIBR54hMoGjma5H6h/BAtj86isohU9zY08UFUZOvRXuq4nAwD6
tXGHS7+7W5ZLiqpXjWV1hgFDH58d3wpgKdUItwdQej70jd1TyrQ0u+sS8P9+OXsYAyDXHvRKNkzu
hFE1j713TuNa667P0SVx3wledaW+LFQIsuTE0OpmUN4RXeKgAOV5YQO/6lGsh5IahJf3CGPgZkGQ
qAxEKLJXHrTZWewkQJICOFmnNwZzoty9eNPa5oaQiT2FF/CX/FIwPuhQ0FPggAs6ADydFviO1hwm
5n4Jts8a7vOU54YxccbN31t8WzMqa8lRp5eP/jzL12DwPXeUnf3SWUtNxkhx9tSBlvsWSKWqZ0vg
SwjdV9n0UzmiMasYu62oco6WgvpWOOXX8eE79/TMrvilc45ffD+LfcNPIZoD/H74N+CHIWYJt//C
IAHjlWw90EEdRVCQqG9BxWz43aBXSPn5z5D30Bvoxca8VAJ8mNYPXM+AwhuqRtf/ey+0905SnTnG
5hfgm04XeCAT84kgsfI0AL8QdDuCaRsj7eREZ9XTPo8WRd+G2znhwxDnQyRCFyJPdhw3qhTcLbJX
P+4NAw3Jck5oLWYRh79jlWsOf+5aKY9zZbHMAApe6EqxtCdfefSWA6BywbaPojSATJvw2HD3b4bm
c9Ui3QGLK0nMk2FP0YY3UsJLlMfJq+3LwCgWPeBGQOhoNy8Y0WRK4Ng7RHVVQQLSBdDLWWfSlAnY
YznGsLNqVgsFlQqj/RJ8P5j6A2oWNghrgfBm10BgQtMuklFH71dGCEMcXBikQFAf17ASbtmCo5aU
Ytmi0OCc4OikMnHRaLdmttsULUb0z3rAfp5If9retQlkNUpNpiDTymy3fQLxSrJyx3O7zPDv9YUw
VSuPoVwgwmYqIKnMZBM7RUymkaYVDCQDB2XUX2hl3fWOEK7DzfD2pdGBaEpSnxuZw+Lm6PfHKyTP
H+Ns419jnQTurLGtK000uMM4HzeGqEU8bhH9LgF+421XOJ7GndAfo+f+k0oESDk2gwCnE6EFZd3L
7kGo7Wx7n8be3q7UdwosAnBTwrVArLzy5mxbBYE56H4vXdagHPVgmVJMfJm6MLfvCAh1EOInGFBi
8rMhU0n1EZr1p33mOgNZ91Oni4rksZXK81sc8eWPxIQY1FSjbkkajcJGmI+NP1FLkq1sy27PmMqV
oRX00tpACN3SLFZRNM2WKPtO3aC+C8fULMa2/t3wzZ5/jufNXMj23Zuz+NJWRB0nvm1Y+4V3/1aV
wsrphPBWJbtRYbA3U+WdqDcL6uEUxgmMz8cespZQcSVXMyxFuXKrswGgl+r2NsngEi2BZOJ0F66S
gTdO2MMdObweclbsx9qk5SsJVj1RO0dbHz3T5tC9H3DErGQVyi3nafIXHeitNraLLJpRe2gzcHtx
9LodXY01g+mFmA2sQJB/LmlM6X+n1GB2WfW0uvx5DyT40VpGcDisH4LZpjPii+YThHIEa8jCsZ18
vVcpNOE74KpJdJxeWNmzNfQ2/fCdI1cps2sSy0LFsUsPWGzYBt4qm6bQ3IIOIHz7u+p3SaEeYvzm
oZwPDQJoOU9GkmCk8LBuxXRb5/GDBquT4PQDC/iQCPnhdc6z29zvZzyLYLCJHqndvlvNdPq2Cgxg
R0zC9oRq+66l6ewOuUGk20ofuxlu3Qm0UkcnOBv1674A258j/LQyU8+PsjA/7OeYyq1jM6gG71vC
y0x1LOHpOMPdk7X7mRWCEp4bTcMGx3+IHq9dBqK21Wxk8WzMHm50rLlBkaH48dwqe5ueo3FL/gCI
019c/OmmTteqsLza5KHQfgqq+sYHef9C/uAb33as/MHj8nYzywCyt2oBImPSEQShuXVypm8LxP/R
y3FqkQGHL9lzeajSOYQWsPOtoFaQUiBDO16jJL3+UApjbH4W/gF6PCPJ9dB3+xSVRhMDM2JRT42d
Mm9AO9xRjwNtYHSTa7e9jYtgjya8DWSXL7H9Uc2pWkBv/x/ErYsPeazZvtrn3lrpefNrnFZ9ic/h
G9spkfEXeEjvZdGeL1WAy+sKK77DnpZ56sfdAmPcBsx+zTbuPjNO8ra2xCl0VvU9OFx0lVwzf9Fd
rLO46mQ+/3xf30K+e59dcgIEmGwpP2TJwgvQ8I2gCLdIBsv37NR+Uf4NtO6nmBknExRNOkkSm0m2
6FadTQvnwC4eGZsgEWTlGnns6SjKYfGeStnarF/ut2Ozmt0T7ePVSibK54Kq+HhGxicMZyZWsfsd
Xfm48DhHUISjrIR5e5PApFstvtgt2L2c9ThjTtQh94IAUjn4nNgoyxI3EdSXZbYzQKc/1OLF6w1w
i3ioCbC9JMJ0+azNOZwVoahcMXA12P88UYsoTMZE/704gZPGixvje2Ea8qb3ATkMauJVtzeJbaHt
TOgPLYe1ekmOmu6Aft5QbneebzSIJTlxerpBUD8N72kNKZWcbcYhuCtA3AumbbwyzcOPFLhLbCEe
3Q28EpwzK6lQBqqbrF4bL/+17Nys9I9/gJnhytFLJ2SHVbgbqaisqDyOW+asUVCv7nYh6tontkA2
PHi/R8uCR/ACCDAXS2TGUAXHldX14KGgYLv/FpE9aXyC7Ts/Oa4xay36rn7MCf2MiZpERG/Mh5NH
88V7QXpmf2f/hK93qFWklX76BdBjeCJFRoNdm/j3jk/vZlGImVfJu68IFAduY78g57RDuKDiwsY9
jzs1JhJg9i/GfUoIKlWjT174jxIFewfWQ6aWK9jECHiPrUTf108OyVEBKQ2SRgoNltqGLO+TU20n
1PtQ8C2jpZ6NVuizLCdRNaHWfvDWu4Bm4s8har6895K32fa12FDfTY4/Y+5hfwgmjaC9wZdGGx1R
JnB23rXbhneFGylK5GQBxcb4mNATGudfhIaYOhAKqty4T2LUKba76ln85Mo7rD4xdH3HK5f6ZTJf
pNt8pgaTDRJmd54g3OIyrMbABYgAVbNBS1KWGilqPr0WzqIPQzU3lm/sRhRy9SaWIV+BR6KMY0yF
4Hqs0XeZOnn4lvS4NCSlXVGpejFpYeJ0cQdTkaC3bw7zlvVxvFyoQKVbZjgtqUCdJDP4yoOIcA+9
AwporvgKcMNPt9nH6nVt6xHZoIqLdx+Lzb2rrqbpWrEx/YCJz0aOzHI0BftFh4O3kdGdzhYR1IzR
vpdz6+E9SH9CFhCp55+u0a0PdljX5lZeug3NkPpjSivvX9ElVTeMZ0J9hwjw8I4lVn98oJx2FcUV
oocLlCrw5rZY57zJU24AMM3sxHuwGgkcVqOwa/4icdU+CXhoNv1cVT12QXiRSTgRZNLNe10Jp05E
w/YWJ8xiKx7M6jc5c7z/U6FpzDEZ9dDodlpjOJpvpd5UOaOX5c/ektk4t2qii1kZMzxnwY+bulhw
VaNXU2f7cAcCCcj7NJ5ST8BK/lo7TZUshZ56yhzBCtMense+HlpK84E0R0NWCTJ8+AspTZLgAvOn
7ufJ4QfuIu8F+Uj2zmJXtgy97f/hpXYZmAuDvXbPpreSe0Mi/x4pjhZjb1iZj2AmXlkeK7sn9VVd
pF9UsOLjmAbx2ybkXHnZVJAGYy4sMVsDEw3JQF1+vn6lW03IfYc3UzV3SQuwHvCEakIu78MIRuOg
nMWBjor5GEf88Gh2KtDYeBfk4zud2GKjU6MJ2WfcIDQCOcOPmTZkT2/WyxrgvLmbOQXaCtXaKvVU
O2sakvWe87IfLUvGlOLzs6ltrYqIuAMKFfg2nH2+Kvi+nTGuK3udcpg82/aYeiuJLj5P4o8+rJCp
TOlI9SIT6JIkm4c+KJ3ShCk9dd9mDqi/AbDKnTLe4HMnRiYghgTzJ8bHpAKToaU3CZOne4+T4NuI
/gLJap/MmTWJTCsJROExoo0n96GErkmaqXlpvqpKAx6e6zJUOooLopP5Rq+473yDmRbd4OdyoRzd
kAcP+iTH7Y1Q/2mk3tFzSiCmjkn5UdBP4l0e681ILpcyE20s3CEbSNEjppbLJl7M53xxY0XKATmA
GThg1TMXXiMyo2Z/CIvk7lOd0mlw3E1ul5BVjfQyI805laR80fNL1TFa6hcP+F7TvHUu8BwWbREl
kR2Pu4I9gztEDv8UmbPElLJrCz60xLvXbMA8WGR40JPuCRQ31/hIJNNCi9laqLO8yZwQtP3yHHOa
2D9fSQL7feGzR78X7uyuTDevmraSP4sYhwbHF5WzWawlNhaP6MyYqLNZNoNhnh25O2O7tZfo0qpO
+xzr4vhYmRiFiDzhI+tGCYMgNZjlCt75OJ3gwQois+0HFxSrvoZ4GoJIFrPbiW3N4cpZnilQHurM
5DavViYjchNlfs435nrWjeKfODaMlgGKM4N9qZeCxGdo2UZFPxbKG64AYUpbsf+CNyb/nYPsfREN
7CprjGOkB3sV7s3AYPB84hzMrRYgJao9xoLBJIQIN54gvLA29cLqF7/pklcegoqjcCIjt5ZiVJLW
7imX7+sTPrGVYig2p8KFQNJ89S/d0rTbETSjm5lgYlN5ZyumCwUhGDbWFiBZP9hJgBRbSffY/X8P
vel3XYpKWOIaIxJd3LW+9NbplIDk7Od64WIvQB4tESZeEqPrJpSvR8Npf5xKzovRCMKswEKiyRKD
a4E12Ny69s8R3Ax+Z8IU7LzAF8ckWmOt7EqvWLdtBeV2SznOhMNxcaCqNbjpMGQ5daN5ZfWS2XKb
QCBuKjJYNl446wB35oWgKHYjCUKrvfqMPfYDsacpYmlMrZfjuHs8p/B8iWp66dEFtsj/QC8xX8+L
h2UvONCnBFFdvAdMsapPEuO7kVHMF8h5f7Z6KrxRHK/ylXBMIrQoBoW6r768AeZ3Wey0o1Ah4I3T
N0nn0x5tM/CtChKgJ76V1+K4utbQGr5LGJwC2fpgzr+4blV7b05W8pfqFQaOp/Md+M1cPr5P0528
L8mVFSNDGvkUYzafH+1zafmG5uP8cKuDLzYG/ZlN8tNTyMWyJCWmlYw1h5F6QvGqyZUAjUlNDnwT
mFZDzEVsriEA6XmSRiXBP/WJ1MJNc3Uf2Z9frusZ5Vmig+D/+BvI0wEDGPPlwwszyY3St/s05i/k
9dSHXX29yDZqZTYD7XgEF49bXbphCUwUrN1/vBIyAsAv47vsjKyT+9e8KIMLMxGasNsrqRAQ3Xth
zcePnzlbjpTW5pXGut/Pi1oocKubZPqAk8/gsVPR6hWn/gx9klS2jEN2mA8BJ0P7P5v1da3Llsii
2jVd/S9FvKEvPdkozAfyCWA/Hmfmbvi1TupRGdT3fhU5uxYDFg2/uiWQAAxfW7BSxQVSog7Maj3t
CKkaBe/L9lUKvgqeQq310eUbn7xJjRKIP+jbdicIrtfeL01wXzHk/7AX5mT9CAbSRcUUUCxiXMfK
vRn3Xx/iJBumwt884WS3M7QeTh2FNACod1oQtl7NR4geF/z2F/Jbjo8rKzAGaU9H+0d596XyIQ1H
m/fOwj7Zd1WM2FvRZKjUfhYbwxGDSu+7Mjz6lcsZg5SJOKFltuzRL0vdw8NbBOpRpfmEa/gNEm8B
HTdKxg3DmyN0nq9R7ZU9VkHx4ERQncXjiLeW97rPCRcl4xWRNUWrMPpnfdTx7zU/QhfZlz5DRfOn
6z4FWDAg+AfIGedM8ZUPGXC7ZkNzU6SjSkimEonCOXsnQEyFjU/c0S2Jdhn+BjnAMuC70dU8iOZ0
idKQgvqW5/zp0XkzFlu9MnHdbBKrL/sfREnPUCq8jll8P9MhZulNKpmVmRjtt/V0MNwZElgfhckA
PH7wtm28tGGCBwGnLr1qRTrD+M4twMYA1svvaDYuCUhHN4y0S6Inj/ywYu8J4BfqfinETMfGwnvV
rgvzyFv7FNN8q9EcSBWjWcpYCU2M/Ht5/NlYVW/GRGJxjfDUZhctrif7AMC48BjbvSFwumvcdXie
OS07X0jeIhQX+NEKJbUct/D880C4erXHXDkDRSqDDloDDi3sZnSFxa52C0Q9PUx4dfgrrjx3Pl4V
MfnxDgAdCipA4xc5k1MExzV+pFl9k60fSrhlVux3JJOJaaSGW3iliL7HTgmnVuZznUMTozUeeHzN
SZEguWXAqNOWdc4VmAsNyNslqCJ4dDrKQcWnlDRBFOACVybDwzV3zETxTduDgpwojvblrWpDervD
SATdBgE1oO3+wy9CDcQ+ax7yaqtoTFHeS+i2kH3T4iDoo4X6nGUQperS4zyuhb3RMDW/dXExphPS
H/WMNE/C7nhIAtiOBJQ/++ooXh0ODXwBbfoyEgiPdGz6pGWzcfbRxv2nMN+7Efca+iLEiOJwKKR6
YfD38jdKssyXx+sAJtpa2isc/5S7s2TumAgiLhWjKVsimlufy0dN4AUlY9BNGTJEmbOx47HsHpqL
tRMGax2fJut/dLbyEhHGShMj8roJkxedKhsdIDPprVSCdh1RfVrIGsF7P0YLQJW0L092WDLxpGRK
yfk302QbyCBJ0uGpoVq9+vKa0qvYbNN3UUGLcoEyl4e89YqIoFxdIKz3fG5NB5GibQSE4hUYvG7c
harmMYwjVlfAUxktMVjwVPjtf0Ua/z6ZpnFR2ckK40tsvZ90yA35E3yx52ydP0AH5II+mOiAy4Y6
5mDXgSfY94beco2bJeyH/oGNejHQOjGoPrvxtOZHGKw0Mo6eQ9XCiZQl3lf2c153vJRFwRCXkYLp
fFxTTYz7LV7t3IOX8bufUG4dDaTAdOanEhB51lkX9FGsmm4wtT+NSn+KiKMNa4l/Rv0Q89MlzRb2
bA1Q8MtXxNz/xOKfByo9DuRbf0B3lL5dFSZZD8q4wcCtPtyjI6NT05rA/ytbXWAu+Uxdt5Og+Qhq
P9KBCdhJwUdF16YjLR/57gnb9tQ18kMbtX/BOr1zN8mQAl6/2qyhzUocvN6Zl4Trd4mx8xI8oKLr
yDkNrgCNVJpMAUSwnCOZV9JBaY+A3EvlPjEoRfaLwtGTCeeEq8VBLzDE9QtKu31FtplR+JVVBDEL
/WW7dGIuqc83+whxQvcf0SsJeKqhrdUuRo5dPikeCC9jCA9Ky0jvI/AgFoJi/4m8zc+RlzF+IETG
AaizKjyQpAMeRFUBEixGh2brMrRgIcmf2qi2mmo6lbNf6mpc+97zJUs1wGnm0LGEvyyUytk14kTW
Y5vl3A6zf1aJwAInHv/jF5JaGJan2cY34+11vnmtouBWLH118lLXcycaL4qpuyv98cyN5t+WPdSU
96PqogDzyMcNzqy8j7tCPeLbDuJJGv8nWtV5mp20cYsFhMjDe8t/95qbJgd0PRNbimxmFPKRtb6R
aXpmc8yPHvAZ6SlPbifuAOK0JR2V3QND8WV7jC8lhya5WbHwVS5IcCnXjdn5Fd+lhA8bEry9C/J2
RPa+vxw9o/SY+WqYFmzC0wJHqOJiKXVQXnZFLrAGl1cRO5CVzQSamM4rY+XQTTveegzF8652uMv0
do5EqhNJAF44wZUvybsy4EwAh6GPnflSZsXzP2U7xCdGdlX74SPLFv72VRMTXQIiXS6fJQRrhC3K
QSO1SB2a6P8AbRWPzG5Ohv9jkHqbcEemvbjeiHz2MbmVi683cqNt81XSe4yC565ywnDXvvNMzj1L
TUqz5NMuyHssIyDE+O0oEP+foGr5Gzev9/SMFeHn5iju/6M/+SRq9RHuNpAvijvdXAh2by0nchXT
eZvdPPrWRfhNRmvXpuzlmHdZnZCzad0KMczTXPwQ2z/2kpeXLD5z5GEX+yNEtSZjEYfBCxvHoRKh
d3icrGvE+/xJe6WmZUqM7u1nokxJZtUz7oGvQzi1W+jezAm9WMn39pEgxFJbiblsee7HfZ1Vtf/p
gX14z1wH91nJpobGHpnS7dMKT+6dVx1X0D2Ui1lUcvLM985UtTmwEBLC+tZPDuJbcXhBTdmSWqaa
rRr4Th7piA8dJdoO7+9z2f0fdhgyqf1NNMCk/jYO96iapIBukHgaUpCjDyMmBy6J7M7LuFqwJTwc
HiWPRujHtLVjQ/A84aSegga4+UnBnRp1rPe/GS42Sr3e/Zq6NiJD5fL9H2zM5uM5HvsEzvobFYjP
CEHesTjX+o+6PtubZaKooaffdeKzzkF2HLPy0txwsLbvOoBhFVpSR3x4ws0hdYx4Ac+00q9n7hUH
Iz+fYL5L1IT178aCUFzGS3yFssAq7uxyJ8MB0aiqHBqex1wVUHEYNU6pqzuJzKhHx6Ts9YKsawxN
Js4qvP/azxKOarxSmzHehzsXxZFxMj6dCmDi9JsX6x+Fr+guiYK/L2YC/DRPAKk9hknWO8qq97ey
2chr4OzsgOiLggJEZ9+PJLrXDz8yjswu47gJxtkoA4hRLdNvBVn7mgFqP9sq9psWp6BIanPrBtSd
SH3MkuRHTyvVsimfV51he7K/MwVkxdpmllKWz/b5W8Hrym+FND37tpJhRYNjh7dlkLJrtqtQrFO1
YiQWlUwVGc81/FR+22yMvhxeNeKUqSw2QlR3T1hC9fDMObkEBvqMPbswOuyLqfzBBNC8dcG98xSa
X+aZ+XEgdG2vJU1JZ5dF4fOq3Rx7Jq/ULwNmW5Hn0jNOD/V+aBmzI6cGyhXODDqPsvszXsHpxmcZ
B77vLEI2o+jknw8jJmzGcSR+AF2KkSzX9zsHNGeeLU5j/BlDxGz9dAVtkaNzRlQNWzNno3pshMmi
UkldCcHR67mjaylaKQQVY8npENPMi2KrtrZDJG9cftupGN9Ps1RbWBrckQwSQkGewS3YzJPp68Rf
7rrwSIL6k7Wts6IqagPs7nSJtBRNuqZzz+C+t1IuLB3AE36P5WjDAKVIeWqYrqZj6yARcanwoWLm
0MGiGiCXJBRyh/pIBF5P2jFUVaO/uwCoJnTBfNbCoGufdDRKVNZpr2m2bllMVgJzYOIrJXlFqjy3
Cx3TmtaveVhFWTVlHALMRZOS9aSf36z3FdZjFshKaEkNdifi4psmg1gl+XD+DrHuF4CaGBxfDWpH
q8nwyFypArDvFD8kYq3lTFE/kVuwkwhB9GgPAQ1CPO/R/MZ4bkkrqdKnbeKXn8NAd321XJStjsp9
KFKh21OIcJMiifiUL368KoInZDmFJpt5fUsnZpLWUTnU2F8SD9ibQHyeJPS5UFqk10iTXquDmtyA
F/mJIeXhOVMQfXadgMANxxebJBqlZngbin2GXKyNM+IWDLo7A3T5Hf5hf+YmrSohxJa9wKP4NNpi
M7kIODGB1B3NdShp4o7YAnLMfdy6vLE3R+MaR6RAuKEm1IZIJ97CltfxLS1/GGXguCZtmTMhfGTm
lW05ri64UVCUvTb/9+WJhrkvO0rNduuBqutQ0WLCAfBVNj6FGbIBzJD7F3gSQoLSG2PnisyPQmah
ZLX92obBi2TZymktRLbrTJI3U9YtUPzGYLHTe1bvYE5JKW5GeZ2TpvLXoD9hi/+6aRuIfKHTqGpt
FrPUoQFp6hQE3D+D7dIAc2TCCZbrZEQymmUk7k18Xxa0rNd5neaudO1NBmESB/DW3/8EnwRFuNAv
fermJP3RbzpDKFgAxa3ZwD0oaluQSEEJlGpgVt5Ix4zMTeLHMDJWPgsgZvtG8cVYwK/G1ie8FZQP
82CcBJvNPyMXnFSi/Ps5V3kyZsRdGMQdrgFmfK2Yw0tcjke7KRgpH4mLfqxhRcFo0rPp5X5ADOTO
ykNDvd8CbpJ6SRhhduqKLEYOvmI9SsZKkX3YRDn59M7w0jDiG0aLJ3lpasVBAB/nb9aQzF5RgE2e
z2FK86d9E1gwwNvPH694xPCOGuTvY9jykx2XCjbwh1nDq5PSfmYsXBBIeuYsuyK6UXPyECFkBKBL
VejyNJODYC2RvHQxKYy0rH9AiwGaiVska0DjrhS8rKqLKywiBeD0UFhBGARYVgNxoB5I5XzXoZS7
FRiEgIaoUJq/iqNHyb2zNIA2pJw55RZAvWRWocDe8Im4OT5J90x980/qCT/vDhudZnjmThxRI7gy
UxBlQVnw3szDM/CgVBlToSl4rt7JROXfbFqKCjfrQl6bOcO8lDMV8cImdHJl2PxbLzzBS34BlLAI
QnBqz7sbj4/7MYYl91gv6D2tCxzENNNFADRjL5CHyxAr6N1VvGnLiWjqjL/BmMs2GWhaxDppAOY9
nytzUB7Ag64DC723lov0ZNnq3N5KSTxv7ryOg3JTBt54ez48uYLsPMjhl4Upqlh1+jNRedx2X+gw
Il/XZWHkybIIX9wbvp2euZL0onXCFSuacQCQzaW4I0nMvDP8/LnRQ6EkvbKVO3D4CwMCEy8UxGio
cXJfNlHguoV/Qh/kxiXXYa/UPtL3Z7M8g/+3Kj8ozh3L2lJ/+SXvzSPcTIwL73DE7T/RSKHDaMHC
akDrcWD/Oh/1wmUJ1I+cMSa+LiX02qRFFNd5hIIBXb83NHpwaWVWVGIBWKhws2pzBXrdagji74o7
whwvdBD+uFk/daGk6F1Pm/GUj0b3uixb41AI7RGrTbpWOlqtWTH/vj8i2uZURHbosidHkaJJFDih
IQOQIhEnQTBPsACHTh9EhY638lMjBPRUcBSytwbmxwOX8PGFAivjlCLdzWnmy+DpDYNmlgCWq06e
zh05pvaQbOOgQXSzs1vEmurm3pDnXKn1b588QowzmRu/HniIAdyGrm0lOOfUSLhDKmKIN+okzR7L
HEwBCP2YtrsjrGX1huFZTaLJdfcrZZyO/1gmMex/0d0q36xaUh3s0kITuQznXy2G9OgVpO75xmdJ
Iacsglfit/pVfpuzfjVuTqXkKdgYjMfirWZiH7ig85ivfUlDxePnJPjtQLBDkf3vNx92e/Ne3tvD
tnXJifNcFhYiy2KKCeIY8CQQQ2moQ0OgTm35FTFvyYpfTbyjHaaUUFkLQuY9JxQhN+rdf1Cv7lfQ
A1V/2lBBlOvD277+1y1QqXy+ynKQVZmh7aIky9S93x0eW/Br0dl8TA2p+rEbqonGmvxn4ssQV6iR
TiXuycAV0dIfKx5RBgi2OaW74TtpU5uJx5PQywNElctU/7aLz3LQqwR+G0Jh0zhsi5Y98e3TV4CK
5JYBG2AKQzMU3uU6Fj2w7pnfJaI+jZD/eIT/sgW48iWBJzVZ2nExzlb5kdNgWm4nK//IbftNQXPf
Z0uUSuv6MuNusUY3TdbT0lKiZCRSmE3dppiIvWDaJidful6rt4928Owjp/XqE4S/KaDjPgGIY96B
ZyfLAuKC0tpyZz/2Bi06K+4WZ+gZVhVfSqA45mAosX6+V+CDnW+pELENbmGfO8yXOzB+ecQ+hyyG
4wVFghMs9n5aTQU0/QBLdi3Auw9ZgWd5r+v+9rrdkc0xS7MvNG+rKwXMYZY4DuihrKacNaRMMMJI
W8YJpIff4ypNzaD2ZlMBSdLngdonZ4jCRmlQIf1wQTcBApSwfTYRg/21QLruLRod7SPVgsjIAIjQ
LZrD6lY25Oa77/Hw0viZzq6thXAIHS2kZhpHmt8pitbNeggQlspUC9JscwIKfx5Lpum+o2atid8c
5xiBdQS957lY1CFYTPxnB66LsbwzjoG0ZcBmP1n/BLBGhREsHOvtDPtCYscC2GX9Slrz7heHvO1w
zTiVuz/Kf4SvhdEsYoD4hb0fREPdIDGxcasm/WbiRJaonwg5yg86ApNVTT8VUxXzuhWrAH2sxkul
tAvrQMxzrdBCP2Q6WdAhOGxqykVQWgtsLbKu1L5ZWyCpZ26PWog1jjS4MKh6G7zEpVs421UVBPiP
in2nGOEkwGPJ9dQewcBAoA2NhmYP+tEFrS2aOKNRktvsWWXYoop6Us6ln1V7M0XiV16gHYQkmTHO
7Ajr043UEwQ8p+csQQA68s19iOnQRwwMdcWicbi7BxIsfSwF2zbSGI6aCHcs/Ue32yPMK1wTBUwZ
xrqc1DTYO2lMNfeY+dU/THd28AfFSrk2SdQqywoPKLGWjBlHYH9mUS48BEoFwZhCOxlwKFsRY7YP
UeZCFWPV0luBrL+sX6Jd4NBbTDQNNoAzokPdzjeCgbbOOkKsbJ/CYKPY2zkXWk/4xQ0o5DX/NEc4
GXITW3jjVBJnkwqCAaQm2PEAp769ttyjSP8nGmWusdH4nyrp398JMDh/JH0cK0BeBwVaiF6p2Cyo
EtRK0FIopCjLFAAaBsvTD2SoNztscpQ0/UjVI56YuANaMncu7MAfLmUTosNDBWAlMVepqzPs+GO2
QwhZ4wG7zL0LwQcXimce3kinZaHadez0HnrF5hav0ikcGS7jQe3T1Vcrxcc+1/i+EvQsQC6zBvTa
MFNX9nAlqpZoSaRbt8/WI+nTbhGJFY3UAUk/155K0ILlPwTSfNBrdClXrA/XM5wU2YyUVyGyoosO
5K7VnFgMgf2dPxpRT15cCSXwfPh8ppDzYj5MrmLnyhxzaGEA0MSklU32sRpkmfsw72fuCHW0K/6h
vcyqlxDPJveeJQakDxhLNayMaEbVw17I8c7SARVT6vTt0+GfHEiI3lSvUCugjsABDvIa7qogskEZ
7tLM8tn8WV3p+6213MRQs8Zm3o6IsKng4NOjpJZktTTcQeCK73gU31nVYoo/0otJGjvyWZpqRrbV
yQklIi+wwTCp4a+y05bDsWg8pBfABH6stqO3FT/ad5RK3gBvCOnTl7KRVg9cp/LXM7pdMR33yJqt
CcstlG1iEStGbLiSruGVNzgEVnfVLP7DBcNQyjWN99UiE4DfsBzso5VVHVTNQmW4ixDX5r0N0xqJ
hCxrlof90EAh1xjL/j+WF/t+7+f6Yw/fNzCPKIMSrsTuCSO003wRJ5cyYu1TvFGERP4GguoDdgIH
J9FhOsNyUi423ZI9aJrkDH00CDvsHVSkLYs5JsUWkSirA6iWhAQTZNNroV+C58mtiHBLe4FvqNOL
pANWnHypeyH9e9WiR12rYq3LnVebiehUsSlHmK8k/S+pXjcv99Dpk3hYKfBp4nZbBlHY6lNCFg28
teCrVEsAFiPYE/o3p5bNMTmlcVTPbjmZ6rN8g2cdgwn3BUASdHBcliNjPJbZ1AleRAd4olhwOy6o
x0wAkPm7M4XkCYxVzE8aJaEcsPlECEAtNz0IkKOjcLT2ZGy+PSs9rn1cEyG+mLEDUaJ5W6CX0+Ch
8ZLFh6ILrsbxVwQteGsUBYIxqQng+exl8wjuMo9p/cKzzXs7x/odLnvVQNQ8M8HeEcE2d+Usds6x
MHIYIU89o1QlHexhOzH/IBJi37+Hl8Q9OhfjaX1swcvvVuWzr8jjokvzfX8HcyVZxYlfufhF4Opc
+nyRuUGULksQp5LSYtWJgQWXsJ9lLEMoU2qr8TZRB3OjTywVtmIScVJP4Hs5JNZ29+Fo8Z+9ZvSG
EJUzYn+SwwV4kdo9+zAGdPnHcEKR9CDc95LCTz+iNtmvJosNKYgk0Bld+3z3awBvB6DFBnX5EMjq
IC98LQb+Bf+jVgKAa0p4SvrL+P9UBdkvnUWzGLnOSIUAvq33TeVcNlyAFL4ivLFXyZ3zLLpE7GtG
9iMWs1BXOgB4GUPQzQ/+UbcyFich2gGs/ACXae0HwSXHv740+YM4PoYWKO4tXmwbdq35PYbrES6V
RXjXu5B94RVTmAZMSJyQ8BxT/sgyCpCA8x7eYa3Iuh0OKTN8WlphZdrifOAVKv5Sr/neDC3Efjen
3XL7o0iVIijA9jp4kycP6NfJsPC7e/Op+UmT3pMnj3bsS1aGflD8T5ve1XfmkDRIGriHILhTUUA8
YHi0mj8nWPO7hAn9Sc/TOLnslk17EKTZYdZfpWOyAyOUgt1kqLfQ53qRODwYrfiQrJVbADeTbRhL
R1aw1SR7FajLmONrUD6mvHr37g0Y89XEwvpAC2bZYp9W0KyL2x+CTlRzS83tDqhH/gONCWtNkQqd
hrSATA2TFuPfzoX1DEU+2wHQAEpzSoB6lWIb+atrsjghW5PLrwQK24ORxakR5HU9qFMvguykpaH9
Clx+AEYIc1K58MO1WSgJ2qD2MR1MFbRF1C+GMc5phENqNYOZUnY1FZIu+K+HGLHG5JnyX38YrLNa
SdOyR7J4NevmIs/2zP0zxa2WqHjMxFf7mqh941z5FK+DsuyvzTq0SURU9qzIeg/lvVifyjbUSsRV
ggkk/Z99AVizuAVykGI86TGault57pI+OHXKJYnnjy/OBprKyB8pmE4B5fNRxwLRkDK1gAYkkBL/
YueoK0V+FN0JSIv6uFROKGhnEb2FZwmyVFLTq/QoiuSAkHDuTKMi5qhR6JFQy6EqCxz/MSgkcpPc
n5Y0GNiyqFh7QmplCqMNLKMVmILSAlO2+HRv2r/uAwwiZjzWSearZp27JKk1Rt3H2/uj0G0aCl5Z
HWB5acLdiyM/EsjXqcpoBaSg0PMJmFFSTQMx0IBiM+DsidH/wYakzB/7UOhMdANh6cWCf1xIvnX4
njBzgBNf0h5zHqQ80F/arSnDkSXWkaNx+Y36SgZX3RcLueFm02Y7a486Q+T0xFV84IQqVomDv+aP
bTYHgLoULZlT5cQDv0qxDuyZBRWjGhPMKo8SQ8SA0qOBdzriyYgcFVIc/TYCRACfEL859J5QQjbU
0mDumTJutLBZLoBuY3BY1k4h8Os+HWTC7V67Yil9dRRizI+WUGgh0Fp5T6emAWBrEzM6uiOUDVib
7wHMjDKCHdgll8W3/pc2fFvip9oel3vwUyaFKT/jmet1nGRA3vbhpKwZHbVtPt9V36GvzStIuEN/
obTaIOrCY7PqJuy49QUuzuiZ+/BkeZU+sbihpZwRGzxp2O1LW1Ia0YhqKdJfS7w61shK0AnQIRlc
6IDSYc/+py07Rv+yZgFYGHy/xc+Wu6R7A2Yc0M0wg2Wu15RsYL1TDA9u3EO2x0OAs9pUGab0Z61S
xKOORBbFpF884ladWGKfEYQSH+Y1TMB1SFNBNHylN+rFOhgIKnfOhMzeYl2NJ5unjfQEp7miFumS
ZFEq2oxUwWhbfhglHZn5sjuBagnLj5cv8K2lK8DHSDz6jQ3MzgW5aR0xQ354yVivvCRiOZ0c5KhS
8PyaALZgTnk363kMOqBf3ixC8dYVqKsoVEcy2y91On/IWPER9ESm9tjf3gBlEX0QOQ3AE5foKRYT
2JCCeo4n1E2/sEtq7F2HMAGGmHMi3Iju6588uQ62dWsklKpnV/Y8ZDiiArM96X3T1RGfRsJyrHuM
SRN9tL8DsOwP+cZlR1cS8uSfjl/M+Jc3krrsvvEW4NbQ3G5ugy1v+R22kvkCa4dB0Wm2UEEVNMm+
Fiv8zN/gccVaKgNUmczKFLesyg0TXLEcDNA6KGzcE+of5y4GvibAwaX1twQS+HOCMONuljSsCZ7T
AbhegHAef42IN0YE9hADVx7nCjYxEMFBfyuYkFe5GKbJYKOBr1I51K7tqdOXqBE9PEpPmJRh9cDR
2ZQ97BYToa0My4WD4GIDTm2X+VB4NVHfRRRqybZLVYUpZQtkmIcd1EKyHQiTLDNNhWXFK1urhLC8
JzUubph3Xu01d2K1AR7C7Sa7muRTspZyFVrqg2ZrOOKZnia3DPjNYIWKlr9W5qVQQ1/LdTseNy6b
9+v3C+mMPiKCIqtvR3/wOQV5YbDiYwngglhRFhk3YJ92BMzy3yEHizB9633oqHjyxL+ReXAWhtjL
yuXvxylpSazIf83+T2J26foEV6IRDGHkctgBt/dZdo6EHM4cYLuMN2Yagu3baZWOGKiVlnsxsDow
/azxdWL0uZtYOxIkeBhHRDog2CHZ4eP1cPxHb7RPDcx0BL4nMBU1X5MMTmkzT0CUEqiIOdMQ9QO2
0Ux/5HQznhrKrkYdrea+ZG5fLuwAntR8UhqJpBOtnlM+6NcYnQ+QA427ckKfMKskKEduoCNzQ2hL
k/ah+bvKnTlJ3e+6AmHDow2QTi8XB9yU+qpk2szHkPTLaHMHZQs4ZJtEv575q5cIP9xC//3hI2Rf
JeZs9e8M5SKzd/xbjZkzqh2EmsB9wG9weqXXKcT93uQx1kTUj4t9il3Bxmy+/ITZ26CxmGocgNnU
Ea4W3NcQ+eQO12oArVozGeD+cYU/vnbnj1BKLf6jmC725yA/nS9K2bRLTglXqS2nwxLLrI6yB0AB
fDFt8yJ7CMiBfjJYnE+LzvlqU5XJEJJb16eB87/pU9doVgW/MIhU5SiamCUVgY0nt99RBBiZ+5kh
lJ5Rf1+vpchek6fw4tPgbnij2zU4zR5x66iGyTgp7m4ldqezvQlbpGhCaTPmUagMJa8kNwo33On6
H+J64laedYu6DSrRqfA/73WulGXKzj7riyjFzdE6AXXrxp0mQjZPoos31+3aCbbJ1DRC9CjwYzEj
0CYE9LLnYpKAqR+ZX7Qyml5dXWhB1T/Kmv1DsNiFlH6DCD3yeimB6Gr24BAtbk7mNHX/QMWGWs6P
f476mZuFK2pRt4ChMBHmf0wOis/6SoDE/w5TblNw/Bc3chx8pl+CTbF5xJgZBS+q9tn9W4tm38Fz
M91HEQEbKf2/KaLIDhoMJeUCp8dnzctnkm6PhEKkhKqiZCfi43qAT7aeRYcbfBxQGQCDt+1t2aUb
Bnfoc+AqywmZ2kfmq6pq+o3rglsuwvRGCg1LAc+maRGCv1E0bvK//+7v93K0dyy7C0hyLDuzkXty
Lmjo5scJKXbZB5kMIWP/fqqOhzNGkeOMFue2IdH0mjqEOZNmggSNFSgu2oKKwQ20Z07AYrCmFeCu
VUhgA8bUOLD1BPr2M30C7qWKdcj/KhyQrYVmjTYwmz2jlGhf+wMztM7eaIn0U5MiLjaeOqWF7zPF
HAq/gxqByZjn2ASn9pHIDiT+JS2cUOzX24TOBz59b6H7FXF1IuTjJF3WsOSJpMHO8SeJ4SvMuhRQ
kJ9rswQKYdYvLc386RrAXTnGbeY+v3t5qtO7wdgpc1/RTfdb6IXD12K+86hfmAPIqzN6KvuRdtLC
1eUb5efjvnPckOwu/VM7h2X7IFfeb2ofQGFJ7AKj7JNUiPzDk2/q7x2HzAd6Hogq0wgHUBKfmiEZ
11WEefnoozHw6EmZ1wFzwboU+5TESqzqrk62xoeYQoFnE7fIwKbKrVcjBcLJxw5oh4wZdrBOy2oI
5e2q4pZiUgbzt9gJecE3rsyaF0zwBXhgfoko2mnWnlS83FSI0EbWwzoGUv+xs6VHk3t01OxQjFMR
XHBA+Khss1iHDTxSErwgrsZsxKA9GmrmlqYYbcMInBFOjfGJNhmFhB5B804kolN0xEnAJts4u5P6
Setul3sXHTEtJbnD5EKItGg6znbQ0HIrql8MdOr/MJzjMydawjP/5ZvB/D/uB88rpIm6E6M9cbNl
FMHxKymGqwa1fzdeUe73nrysXxpWQbu+j/vgoR//yyIP/E+Vz7K88zV2OSKZMkOLd2EB9R8hDMN2
aYh57EEuOfa8oni05rgEpvuCicTiH+SR2bFSaX2S/Zv1O/pyo4WWVEddb9mMtgHQ50Fe42wAr/E0
N6fk8rVYfv43pE1t1/hTrOZhpD5eRlQWuj6vZtBNgMaKTBA+pVHJrzI4+OSVrL8Fm9O1Jtbt05W5
gMG/UM/YwC0mXp11dD1DkVQmADUZxdCPfIX27/5llYOx+J95MR5eXyLIm4QfQyKgkFOem9hDlpoK
22osC2u1fltyDIkptd/6PzC1V9ourF4ux+XlPABlnU17gHOchrP9Al5wQ/HiCPQneILlCxiF4ydd
bEpuInG8WzsnimeKF3MssA/5GOAd+IkiUI+X90Kp+PqrVLKi8y0XrVf6KY0Rp+07nIDM4w0Cv6wv
Bv3+VyDYF57ayIs5WfS8hAh32OyQU0wuFfX5vxnuQysqHRvMSFacbqAVMw/9XtcwEBQqwVSWKX4I
R11tv25/FGo5UUX/vk7K1yTvsSEIkFyOVRf48/xW/oY0syYkthcqlsRF8avOzNeIqQ6VGfGyOVxd
7Kbb+rtfWXWI1Lk3c7ASqrphJltVOZtUIeeF+1oqmtTd9hrFxhnNDyj23XZ2gWZnnROBBFXgxA34
nzT5LpA3erDrsr2DiT4qAhoOpRSOVrfstYRojhsTMu1Nfrvo01J78Vvpz8IgOV3LNCrdSv2y0dHs
frfBEsBqhLz+pqOzDeo8+ReysNvl2HownKpZcubpwuwESCMhHG8v0r2xV2jsK+9K9yIxdwGh6N39
ViEukl066w3n2axLtjPJtIbJJO2XyJPbpovadUOdpPFbBewRwG5mLAI4jlPc71oAXZBX9jpUqqMk
A8EkKCDA6cqZYUEr4Pa5VesBQjlvh9ypJR3ETojeCBj6pqX9tsfMmm56x4UeNH74E0m2eTMxy/12
2E6rPE/NsPPg+ylCWzrbOHjxphUKr1e8/3LGR7YPQUWXbx21Su66OQA0MMa45jLJ+tTFdFbKncfR
K3gjnD31XpOrPJdv7N34lVqSLB+9ZIB2EE/J6U03ioqIVkL1L/UTcof9mFP1O4BCtMWeb3A78BFk
dJIWUcogov24hDjTVx7BTu1u4rWkqOkV/kTfG/Bj1LfcAi/9g+6k22vj29aFqanHcyPG+6QGTgPa
MnzJzVRKtwLATlmfo3gUnL5P3P0DNlolOqpoqC5ZDhmufFNmgp7HxA14fC+jhEyNve5aj/lgXfEt
RhIdjeGuyp6F0HoB4F7gXtyp5jyB3+xU4tkaESSSmXqltqxAwzId2VOpOpbvrDon0c6j/+JiBHrv
ojYhWBqStrx8WVLtMU+h9jKGbVTm+oVp9lgRS49b+ZIJKjruZv8ThxtlWuffPsQ8tMJrQNF5Z5xM
0aVr7kw72kaw5Gd6mGzY7BFrjWT10Ufy0er6SOXfQF93aIuJ8dfQHAvKZIh6l4P5Uj97T7uOm4Db
gvTmvnsMtxbSwYLFXMP0AmN8HLuV8vAjLASb+AS6Yr/5g1Ps1ExrrDi7lSdVB3lzDM4dcpS8AYlD
ckhY10/u9sbGhEUJC6JzvumDIiclxe/qvHeszEaZreWP6LXgub1SqVYtnapa90fZmXPzW0X5A1+b
WjsLnDmU2LrdtnuX5BbNTOK8fNUK1Bcr4ay86VeaS0Ms1tvia5FvO9Y0P4Mt7HEoYSyh1cdgj0FM
sTGs6TJ0OxL2+1h+uiEiH84aXTAYZmmifx41UPZLQttabWqlfl26dc7DwZbIQkShmiYDtso/G2xY
RN7orEx5c9vt973u+wuIL/HOiVYgkoQgsAjxCqZR1o+WPRw1zviKdfQlcPUcttfIWy1xkax7uC2g
35F/F/F2RINEGSJf7qc7KwLz6nFwdwHdIvan5xdyuW4t8HndMLfLAKvbcjXrMo9/00yas3w7jW0E
4u1ETsmnAVBJZLLu58pUkejvpZneLTmUcA8X/SAfiuY7xjJ9SeoFVwo1FX64t+sPp6ovBk5KJXID
jxgEg5XOhQq8wXBfWbHkK6UojMOog9N/Bzp3KoAWQDKFkGOWwLIfUXnFIa+rMNPCaxJRuj6QVB4U
+L3EqYndrHOUzwqCbSW/SPjDpt17ezA3JduZWupkjggsjelohM/5Z+LsD2yK5QOwvJB98GDuEkNX
7R6CHaL+T/bhHQI/ZTf/JFAJGZg2N5XW4kNKRXLkRkoPHV6tmLNhiLeVTQwrlt5l1ND5+8dyE1GE
7h35JPIaSsHD2t0DGkiOxdWlDN2TUQwJX+eWEAQhnTTqD+Cv2eWbwtWwaR9hG432uoV0kZCixtKj
xMo6K0oPwa1p8Y1Y1Oqf1dmNcyvcWHERL+QmpV4FQqlMWf4t39IHUDepO+rRfEC1t/Pz4/cZi3A9
GrubxkwBAzYXZZ7Cd8/U58R2eDO8CEIgHpoFwWAU4N4285i1ncW/POGwjAhFq5DO5ad+/3ixE9OW
4d+DyegKKr3ezIqDYZdDLNpnl2eZQ7ZtPtTB6a1cKyEiORlxu43GQTC99yDpstrLvt/q+kT7h53i
TyGb6pkQRO0IGoKjmZ/6S5VFzEjfGeI9jUcJ/ucvHz4A34Zaq1y4tjbzFLWAfbxhEKJBdmEm7y5g
7cO2xDI8EY9epT1+bYyTWy90zvJa/Izhc/PYuMJPiPELlNXOMbZspdSyUfz0ZPtrXxJlWren2A9Y
1ZYbpHZ2pxW9RSt3Rr7jJw57/+rrXdzb7FDqVYpr9IHTQeliw78/94hMPZefoVNFbexlnLVkADI/
c9zkDckb9h9WSg+ii0x5AW2M9TIWrr1iH1fQNQu3Oj1DOJFMdZcbfeUHvTlN5l3ScleAQEoA1VQM
oJzBO+YYlsPkjT1ifsaUKpP4VE7rXeOy7lh5oZoTmNwDT2eFLESW4H8+B1RnWSSri0fILgGXHz6k
KlAKx9dST2dMOqFxjk2hEJpvG7K52Q5441od/M/W1YPLe9g3imV0RvVjgQP+GjpmkrOUmfreIpB9
ldgnGpqB3iCquiJamwIQkEvTFSycELtHR4hUyagPGxF+ivD86bGjhip8WgS8OE3v1/O4sxGAjNtK
+NyxbRXnMdhcCnzAaAegqICbEiiBJ1S0TxsCGbaMj1iM8kb6zsPG3ag747QISS7iOSH/j/PwkPKk
rwixnX5i683CLoCMAVfNsnqkgA+0NtBr+xHJXt/txSWOs4MbGnqOhFYOGIsrIpfMB3ERiSWNoioO
8WQIwVjYOAq8G25V7kykvrWyglb37WRJOR3OYXSpGrVWfjBDhO1I8vIGZJEEx+aK9GtTx/YZ9D6J
ivQRyv6KoW+If0gvIT9vFdc9jTvTMyGrB3cxsMyCCgCoq7OrHXfXzmTXTRxtWyh5aBPbdYCrhAkj
lxfDlU4WNKGIsERqVrQX58BPaMLjldiYu5QQgDdyQjHemQqdl7/8xRfWkkL1PGijcNZvKJfoOitG
hc1BTBkW7bqOtY3E7BInZk/1SImZccHMJDuNd3FE5MlMTCEQ86u6Zl6wH8YDGMhPfse02NgJuKCI
R3jCYNGAYkKvFJyqnHih2txJJcipmvnUH8PN24NXSKKxGvUsICzjOP3YuqEEmReV4Z5Q8SZm0ZRD
ZtcjZcJbnCM0+lDcfbwckaCqVO4WfalKQfdmEi8m82O1v1Eg2mLRZlgOx4NJqKToNHkdsZrvMATQ
qlXEWhkBqdOjWBauCJ4L0WQV7Y0tBSLq+u1GzN9lTmXo436S9cp2XrHkWGnpvmNr99nD99roSdvA
tP0z4SdxmSfTpR35RxlmxgDBqZ5BCr2OoY0/dFwYX2TUICkmXIm6xz2Wb39ReIQaoYs0KAnemzwq
CTrng7nmx/U43L1VnfQ0NNqJTKbrt0Mz4u1VaFhFjZAqFrxYu8SIAUyQ5F+4JaHBL5UTELdU2K7L
UMXpQrPSRR21xXPk4fJBWwfStY5eJO4D2ULP+ZOCX+PITX49gX3Lt70v5V1k1LwKLA+HsnzJqe4N
dHgNru0hnpCCzXpCoIeF0WX3XaOgelBoYLXhJxwKeR7KX4zaSM37C6RbvEcAptd5MNO3g7Dmz5bt
0sUWhXyH+bOb4TcRjmTm5xQc9ru7YXMZFMDSqqdRprkEgygwCPTAgciSFbqWikGX5NCTj73IIM/r
kXBHMt5AZ8m6xQbCy6qo+Ek1tP2HExmr0tmiLz+f3b3ZmdZvr7VpBeyRr0i3USvudwRYYjb8MPKQ
1HFnWCzj6yGwHUbmdqQtp8LerjrCLJgmhkmPxv66Fxb+h7Cz7+79C0KPIwzH8FMsreFd1yBA1sTc
BfuRz7+92O3QcKHDiHs03wFR/PmCASM3boSzbQ/L6qsPvguV+MRUmQH4joIt9V5JhkfF/PNLQgkI
1upVOx8hTVOi2aOUzHWfz0v/OQJMWkD+T4W1SrU1nndfOtUEq98oiJy/TEWuJBt8QijzxgIf0Rlg
/IcDKnz/SbQdqM5LI52KLz7gEtSV4J9uDnKwjEodEzZN5QyzuGPPW7tPDFsxNS8Il+L+ZwemT2IP
Laa1CtGBM1lsuY/c/4TvJESYfrsK0ZJeLFDpz+K1MdiTkZoBFf4UYTy9rFtW/ycEzBzwJSWzEMWk
qRhWmgj3aIjF1ovBiGhbKINBXAUP3bbMLg9q+XlMfLxcyy+PiyNnGaD0FSDtQO45IpRIZgmct6I1
BmAD4NDo0InlXdMZLLfAzELInrSEwOL/kvo8XytJNqvj9/f6+rm0Q3OF3CpVBo9hwiNmeao+BOa2
anyEUyQ5DEGygkaOghkVxAI1crwZAiA/qki/2JayHNWFKqZxHfS1gY8+RkobD1xuFDGPi6xEAAQk
WiC87afCWfOGPl2b3NzcJbojrrFD22o7mJvIHEfG4PrfT1/aTDTu1vQogr+q4S17j0Y0dex4sQoT
0xFBYmRzlHWwM1uhRX8uJn5kj5i3ZbB5aduNMBok7gL3ys+Oy8qEusp3jEvsPByNBmWGTmxS9aB3
/NgWx+lRL+Grvo6NrjFBYblqDIyiO6T8R0uzFhYq8bfN+d+4JTRXJxb1QP4HOxG4oJ8jBfIfP99R
bGjbWVnRn6zVcnipM6e57E4LwKSgyDGwKYawt8sb1RziCnrPLw/KrlhMPR4e4+XnXtDPfM64pDSz
6xFrzm4Wt1kpj/55eKBgXDjOSjOpey7SQRQyua5/H2A4AmYuxTfgQOgUu0W6AngFY+s7jTvCWrzc
YFjC8sgQRxTfCW2TobfL/8DWfQyOSNUaJQZ3EWzaDPQBrOTPh1FvV7eUmLOnDGCofGGSrnb61iJT
ef/28D6ChcMYn7uHelKMdDdQmpmR9rzKnfr2ApKzy8CNtun4nNYVxEnkocjM8bO1FyfwKygSkZZ7
Z44Vv7t1BQAmQZ/JpNfzO7Bh+oNwXhWgOq7VNqlx9GNtaVWCdRTXf5mcDDoIujLdc/Kr9nK/Bsem
2gVTxPRbbFny4PtCHGW72ULwTU8lnqzEr/1MZM5q1Q5d5WlvGTZ1/Gl8di4vSMqARUdwHHkRshn1
3+n80IFTaKvw2k/S2nDhsvTmnUOG2nhw65XBaAt++WXR/yg/MVrgKbnedvl4ovBdu26HuzZYJu8K
Fz3quunyxTELAv9Gzg+Go6saDR7jyUueFebl7SJCk9UP2mCd2H87WCvl5NhXCK2f6210z/fmW+VZ
mp2LhBcASsmOWxv1lLNxGR5axvmUDmh/YSVjGskEwqbXwnf/QD5PM1N2DqQxZtmdYC/Ikbi15w4c
qnS+J6Tn2SQPxWihTBDMANGIL3m9k+R1awtB/5XVgmmxcHvOMdBpg/+gW+pw2iSd5J7CzoZqjVzm
5jL+v4G1igXRKhbANr/TAOO5e52OAtMOyhjY4DCTdMnn/CrFLuCcbdf0c2IW3+hz4w8YHmNBiHDS
EC0agzpsTFHOkAiUihQ0oRapIhuIebIAeaGqacBMHZPOm/rqz6GAbGCm7/6+lTe6I2YOqaQMKp1t
01iBxyjYMBDGEEFSmqkm86BlKamIpJzoAoYQjW5HbAuhbi7mhjwOk8/5rxzpcecgGEgRqrmXV/Mj
sZ/40VHUGl6Pmu7vBfEf0GChcZxBMwxuUfigWzqu4voxnX8FjjIOWF+PC85b1zdkcj7qLwm+b/5n
i/wx9xs35ixT5RatvtjObjeKPegRcSHh1e/oKqP9e3nsJnAAqSQ/Sxor+3tadkPoebN13qrXX/Xl
BgSMEsYv6DcB+fx+3Gt8R1OOMJFLY0d5xHl5rX+LlBp7GojNcEFzu/wQu6AJKYQ9p7akFmtDAdyp
HO0f/W3TnFuaI7TVFc3oPRciZbraaa1B5H2446O6CytZxaZPtEMedn2/Mwxao0sLSiUcC6eAKemh
pwEnBfkbqpOuQvE7Pt8mz9AnfvMTA9fLPkc5yxPFau9TorZ2PbwQm0ODjmw2zUnQ4oBUU53FQwzM
N6TnF3Dnj1ApW2PFs/SeaGe81hT7bmTi1hLaUbXXQlI8jpRNf3hqfr99l8fXgWqCJYdEHDtF/xZU
+DGDgIx+ZtUi2pUYtIyTrBRAs7xDJfcyaPNAHoEmxqZpAxlRmuBzbQDmF7OTbB0nC7n6vOfzLOim
SzK+EzLDtcWrDyyLPkr20jH7sEcQrNCNhzdAIXsKPFLSOxnrMuFVi+4AD4wDRStReDuzEW24vCFe
THQHSDfIHLz3ucwyZsuRcWiDnu1BjBr4mzsO10qk67y2cRngGytKeXkzExJJWbo3I7hHM/aBKmAB
ArpoNzdKYaAdy867zE1zy9mJGKY21ebVv2fwQrPF08nu5UfuGzaDXyGwj8DPC9IFGSiu/n8gvxWs
Yc+o6sfdT8655RwfcYyqDMwqt4Ths9VAV+URvb0VhkBTuDmfOk8M8xr9akccGy6Q6DHFF2tCXE80
ixqZUxLOB8zee5AXzmhw+5YlQ6v1ism0v5sVg0TOtePoGK7dFB7Owh6Qqyc4HqONOgSzzn3CXd3L
lY9iuts+nYCd2+2XoLb6yRUNm1nKT0au/w/3UFiXD/b5JI0HuWmfCHz6Ffkc7u25+PanYGzx5azu
oWqBSUNK85akV5NCGKCy9V2qPiAZbJRcmxIt8WmoZXaxlblN+ahqYBvegNCPQN98PYwgWkZ7H3Mu
J8wLLw9PCbI5uSFTufZUsjlYn1AhxYSBJKJ8ys+O0n3S+JovQKUIa/mPkxicuy7d0jkc5Ag/dGRq
irCXnLDnu/E+wuMWaZuhpVnqeLQe3uwNVNyLVQz5rjozMxEcLHhwkj9YMJIYwUjvfiJggU1M2tWc
1W0bx4mZNKhFW1xAJZXJs5AJRtQQZ2RhRuOQPUxqc/5Eunz+TfkljuUxPrVqMyl2n+o4JqYvPmGm
ud67j2d286NcqQkj8bFW
`protect end_protected
