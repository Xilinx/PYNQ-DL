`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner="Xilinx"
`protect key_method="rsa"
`protect key_keyname="xilinxt_2017_05"
`protect key_block
L+hTHWNlnIBxA9rTkLcaQvt9rkblZSDzXS4wbClmlniXQQjWA5ouqw3CaI5c3PCu0+rKBDTc9BiC
MQe+45dHFW5H6DkVF462SAfw+CCJdYNGysEIyspa5vuVQkRlTr4Kqpc2/ZGR8PCxx7MSh1a/JYnZ
hYSiWEF4H/6x0FHxfOqBARvDPtKtPZVEX3rMHHmVy6k+4tIFnDMS04Q8YrqCj9VzGA4FYm0LjEEV
lkZ5EPqc9ytFyoaPpNBxYsGJE5Z3t2Jw3gUCxRz6vGTp+ibODMRW3jZLvoTtkER/ZZkCddaPZ574
dWkG0Tu+YtBqdQxSlkA0Xp86bPbwfGMRwNc3EA==

`protect control xilinx_enable_probing="false"
`protect control xilinx_enable_bitstream="true"
`protect control xilinx_enable_netlist_export="false"
`protect control xilinx_enable_modification="false"
`protect control xilinx_configuration_visible="false"
`protect rights_digest_method="sha256"
`protect end_toolblock="zPKEWNadNeQDv0NZ/nWvWBXPqMr5ymoa+G2YIQAttEg="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 206224)
`protect data_block
N/QfClz5CIxBYCh9hI2+iDsSv9r8JxjPQ1kVpVELL/h1mUamJooaX2L53STFLl8HiCJbLbDue9b0
4pqAkQKcm4XRwws36pzMEPuo+pAots8M627LXmSsKCROtnVOIGsQeOAWTpxwQ0q48ovaYGvGMskw
ELJWt5BL0Wri6PMXNi+3SRh9vbRYsIYbyst4UNdelWHTvUy0T+ejpFziCjSJQl7fu3Xpd83SQpz3
UnNN0x2BzzLbB+aZtPvY1+NJYRj6uX7NLcRzxW+RyQXN41kWomJ2WpEt84aw3ZiMfUyUUJfMKzzo
vDn+wcRQZSKlNHa3ZzWf42M0/XVvaE/JDY7uIqd5/5kVxyTDyZPhVQnioGqa0G/cZy3W3/xa48fO
tgAk9nyp79YLxHam1kM/Cs7z+lPKfyYvy93svD0dTFKB5vkYA0Xk0MHtvBTrnrCyZ+0sF8bFuSGH
/qoXQPai7uCNqV8+1Uo1QNYfVpAk6+M3csjSR/EGzFTNCAiH6v+YeLjJeU2QHQF3jDyO4shL4xQM
pzZ9YNjshgbZEUqyENKs7mZAm8ypPOmwzMlks4Cv92qyiL6UdZwGMdTzGvUR9oOYSy3hD2D+Uvok
PsXHQ3xQw8wqDHlK30tOBL3vUqTlbsyBGjvWnyHOcCCD8AfhOo4WqK3G/qfpDtBu6uTj6X9sZjsB
mG/KwcOqkG+SvOM6ZTRiS34CPpiAKxidQjDNaZhFW7mFHH/Yq7TiF4XBFF8tTDvjJbf0UFweNf2K
zwuhjo1nFTRkAdK1y1aPL7LOQ1pMr9o4jxmgTvvfcE9UTNRg6EirDrXPuhRtM3crYf4NIPoF44Dy
lmrqIHgPK5KSzT4zLwIxZ5czzytV2kMdz48M5N9li5eRvvUcZ64lgJZQBFpAozmJdUJgAgut/+Jy
IIv/WROsb2cOIFvly2qOmpzvqPS+0Xin/DARmXN5lD/0ra9pnXfGU/MP/lAxYvDa6W3BEuZk6Zzn
TIr/x9cf6OPm1va2emikxSVJ9iYzOGM3TBwVDWn562jQ1BzAfk1CayzihQMRCQi9rXbnZrDQvCYQ
t7lTSYJ3/owGPbXgxZpS9Xw0vXb5Whqr7g0NNDruy5AOF1xnmBkqoG/fN0Vm2XYhbBcZPLYJ45I/
2RgIjcRUNm4CHMykKie5B/HakQpaayriNcQhEUYJQ8GS6FwSgu2TVWM7vpThw8RwMUaDW4J9fctC
SrT1kp27qMzkoKYadUzzmU5l136J0hyX8uGZkVYHHA5knwuwNwEZShfIr8JuCmc1mw/llvNL6aRs
/S9OVpU3Zcuh3MrFH5xjn7wS3kCs79YxjMHaGykKvXV+TBHyZmBaJtkySBYyqowXIjfWe/TWglVw
OvIp8YVRKg0Lppo0R4RjySbAZrraO52LnYOo1Y/M5rSoHNRQg+iWY+izN9Gqaxb9tjQ/l5IviQZI
zQG7heNC1Hx4Vdw9Gow52QvRhF5diUn3Q1uOhizEnv7eDwix+jZPlMRLEWSg3XP96sGL62SRv0sL
HOSHapxW4/spWhP9BC9Uufj2dFSFpj1oECsWToavtQ8xB25EajgbqObYO2XIPCrYs2CxO0DfrHhV
ohvToxsv7pdP1TVVFUK9aIjz0iVcL7wYo1srnu05ktvSF9khRmh5ViZ/VTAeeQHWADn7lUMYVd6Z
CelzS0X3fFczwrlsdywmR+i0WKAFOOgQ3ANDbjLpi9KbjA76pU3Nf/P8R18tAbMRAO58gU0i6RSt
QWh0uhdHsjVRQG+KEKCp8/Cs8PAnrkHV/Tc+zF09WFkHB0jUBlfoswKEfioT/4R1/Anz20svsVHE
n5LxFInuDhtQ4J4IRxa/XfgYXltChsXYnghPV+WhP1JRG+QFDRkL1oFzs71xgX7hZsZK55ftZlnp
jzmwR4ca1jTV49NDZIuxZICRcmiGD1X6qU8YQmwzPnunHuFG6mz+X/vyJtCMCSwPQi5fFsnj0wiI
iZ5IhSuEA4/lGYu92+gv9UvCczEsI62Czd9mUiT7134I/ZO5BUnSeDTxalRWF6hZhCGFSHywtgIg
Pmh9pmvwcQjQ6ji9/LVrAYYLqmgvJ1qxulmuucISSK8CDSHWDqcKMj4e87urqJGJaGlA+AGyLlVM
OkwI1VSktoP0z7Ooi0Dt3UwQ5Piaqf79sbmgEel+7VPW/zupAiBAk0sZQPVfJTaIakWY1EurDTAY
7EVGO1SKWe8kjiSfqfYoW6ojSqmw9FTKMIRuhNJY70SnKjyAeW6sKUhqipoYR74R7beqYrK0tu5Y
8eLiFdhng5Rop5ICwkfa6kvvcod9kR+hHOnLMg3KjqgQkQFj7CaVvisQDft6/ezzHSnQ4Y73bcIQ
g7MAk3M7OqCWClRr3uq8jIMdFfGhU2QW3eFjWsvMZBqLrgNcXBc3kJU+x4U2ehg6ZxHEJRt83Ioh
NZd2u3g0K9CaiRjZ6pXodKcpfbcOPR0PS3vq89n30oaOoRQFNZV0KbeYkuHG2fVHUpCOU55FwIUM
PTmg081aone1aOd5V307MibCvjpQRvTOLSqgZeWtJbUMaM62oefWNZNC5kEXFNeviKM22M1cUr7g
+VqgAD1+qjk+Y8UWn2XpJGdb+pCWoGh73EmhkvCuO/0miKuG6loRpE94DAOzFg7mvTDtVSe0uXxJ
BOvDNm0nv+qvOPDdrLElMoNlMg9rUTcNYRYxjVgCP1AdbDdT6s9FzGrBlD4Gl2+hlEgQIY9y8Rub
KaWSxNnXxUyMFpic6PLsljLxrdDKE9ipaiO3zG2dlL1Sfge/sB+k2sx14AylinRcI4pBj26LsTo0
q+EfwELgfGnkG0SMJ+vYZnaUt+jq1fPNof6L0KAzUZyMeYd0k66W2Z1i0/nn02nQAi8nqHQYfi01
WgMjjkorN4kNrFLfFyLoDT0v8buP+pMvI5jBLloH3huCkBZI2i1bnK2/FVOC0cf7DowJLaUEI6fH
YJJcqxA8Nt8di+DcQp8SMLnRd0yNvd1/O3yEHSs5NRjwF4dWGlJRvDVAkBtRIZYYxll61BQLhquJ
yJnJ0dArh3FtOzggpYjj1EgY0utpT0mGn/IJrZBVEDCmazf4JFatIJkCch5q4dT8ZRoqZJg2AH5Z
P9EAWZFfPvxE3EMzFC6Uzq0SHptybzI1H/68MHjr53AS46wciBrIultyVDJ7loT5jaXiwQLya0Hw
wGgQpTuIFT88HNKWIZvt8hUc64prqulTaEvss+7mIMxrwqtDXLHYgiWGO6vWZBpaKs2er7p9bNSF
ERuq9g/1j5SUY19vZkPDVYY/Si30KpAC8VzVROoo9DN2nVs59rkyLldwdjQzgoFUU84qrv7nIPkg
QnU3m1/omJeWrAopANnJaqRmdB5SZuBry2FaIBOejX5OEUQKAlLQ+sKuaihosn6OSmpzb880vKPY
i1WYLxvZHhP+3uZ2uEnttIZrvN5qGJXC1fQLKa4/9sfZWRvn7eKS7CDYZ/a4Diwe/mtWIZH1zUFN
Y/ti7X6c1bvAHahNjp4ubGnaY6FO4vSqw/c/UYBEoI20oQFg3OS9tDQe4NL5Aw1SpAEAW80vDMut
mSADEU6tCjyiad/E+BIurwIs5NAY77wi6hhp2lhZcvCQj1V52nfWhIdd33q/K8l/jwh/94sJzFR8
+nm3OpiEBhzO8Kn1VmMdkpgullPMl5H72/3CC/9jBlkLB4ROg07HlgTrtNuCU8w6MPcwi+1pJRrt
zEeEY+ffmrOTRBAq8lDCMwS6wREzaIFfaT6xm8rTYLRboJwilrb4p3dy+hlQGzZouH1wbxMO26J4
1RBQ2TvBpdb90s9Kpp5R4csBeCRtSkmELen3lVJkOTfava6M1veGeM67NvALKrNPmZY0HeRvJVuS
UZrXElmhGTgBrIaEI1VzANinELD8FRhUuF5Xbmno6AxteaNc+hKqTNrghFHGWU5kn6U02aFsdK7Y
u/vH4OWMnJjq2m4+EPKP7mPUhOLPsaFlbP3WYYMX4o8G35zlZG6bipWtgZKOnYVYKM0otdQYVn48
4+1nOWs8hmrcxhWvk6TO0MGQOsiF5ij6iklS+s8Z8IVUi/0WJw97vFN7TvcN9AvVVnlX4x0ch5+2
1+YoxLnZiQQqbcTu8BQj+9Wep0Fm295uzRNj7x5hKe1zZhfwa1AiYdyNRfkRb3vFC/KNKyDoaLIA
9xq7cGhtDHSEzCPZJivqZeh7ZcoE2igpn3CCpt3SX3dVtjWGiXSE5HIBxGLI1LzuEACBUmu5s+EC
UYpySGE7hfLfWnKqDXyVSYD+WdacNJLD7SRmakjc9ZLvSlWB+VQKb9Jwpz/cqp3dkKvZ7UbmKADn
W2ZGW+zc8boaSGsL60VqWRyrjzISNDR50SEbML7AWCCTC40MMd/FIjmxgtbjdtyiZe7ovKelFGRE
MZS5arxwe0lVFFUCXgni5lSlnygoNndDw9TTFhJMpwTczCDXMHx5hk7wmSOIRlxxs7v7ueceMnYS
+DA/kXhYtg6q3KvrXwGPI7ls0s/EHK7gZxyw5nDmMM37fDM57P6t9HbVj392NPhsg/OHIriAp267
E8LUP6K26jW1sMCfaCxCZ7A8u+VjgBkjpy62Hkwtbq1gHQHAeCwSWElhjKsqgCD64lw8q3aAUI1J
YsLTw+wUUVoJznLfs6ZcB3gjH4v2dxRwrlvkAQyS3cbRX3/YdwaFVrCP6u2F7xsDy/KeM5nKDi2z
M4lltzjpMnuOl+FDnfeFTbaImJxIVqQD930A1iDshaaVN/39yRdj7uMtVHhtF0ZHUYgDcAGDGnV8
ds5fT1JOa5OjQ9OeCRq2smr/FVrkOWLLGiQi5U/Q6E7q70eDuRR4coQn2uVY9INngjC/LwSEhhDB
dE1RMyVgeDt5XfRkl0Jm1mbuFQw7FoP8BPmSPXSPlek4iWYMz93fBFgJQhir9vM6dmepVWPvKR68
+KNMTpLaqNwfbb8Z1MPM/jpXCTAkl438/zh6P9zS2yKZ/NIC8ZlfssTipp/2iYEA1WaqxuxIw/ML
15h2e4nlXpjsYg3tuv0iCSpV5AIfnMkF4JdIfjNfJC9e/t3TNcSh3TwpdxvZ9LYomwVwsKA0pfXI
5KlXAMLQf8jNRTbIqc/WT8uR4ZNubBnOjQl3ePQlRBEDzgr//O1MqBmvpCK6LupmIM9ecs9sqNvx
K53Et2izRdDQvUBVlQl753hiEZBv+YYXgX57ly89GPsNnsIVGwWA8R6msjeunDHFOK0Z2kN80FrG
VjpiAXSKOucfLkz3zB29llFU8ZUCwUYh5LKcWFPP5gaO7C8vFfb266zchGatERPQfbhUb7GQRz6W
1SHEwtmR5a7XLyvt4ngI+WiLPVA7aywQs2TblrbOd5KtZJSKAq/4eKW9x3rzjTPsZiwpS5nGITSq
1zWpnCzEgQd7o95F/0ITYkII737XFshVn/MQF+5saaVEsviOWrufINo94a3xwKNqI584NtUBzMBi
5KU6+gTsCNcIXrDwmoBwOsJg8fAMzXt+hN7qexdwNnFC+UXwgb06/EzSG1whYAu+yqSvBQYzcLEG
1wsgMYcLR9OH5PnIGzz1Uh/8IchN9WL8l2lICIL8MLzV+saOTykfbK2sKNizFcoXbh/chCr+SiC2
Nh+3qpDOyIo+FUB7jRTc/pPN3cSTkQw2rvCdZHXEyM3E3N0Voj52XhUqRM69JIi7q5zXQ5H9FTbd
0n07F+HDXh2EPUKsum8A5hN4StOABci1wqtcisouZoGEY777tW4r05YOTZ64KNn/lTzNHqL9BU2n
rE6LgI8lDNhm8ZyVFh3iL76aq7zmQVJzCljmc6RaZUupGhnTf996CQ4V1HC+jTakr0Cuql51uVF+
tDKNXV7EeY2DiD5mp0uO/NErdBbOkviIlpPtKTzPfNUCCaTWoMLYOWZBU7MpGjBkMi0AjkkfNWz4
nP3LpGeVLVA//US3UZwLYoY9lla+rtGae6pPkdoUj94A9CTuAn21uK91/Rphok91zTLs6QCFDvPL
VcPCLsr3FCCe+2Eo5Ng1fYdo7HO7kXAYi46jExOCBjW5FMXrMK7isq1NxI59VPKEoYA7haznEof8
R0SjH8ZL5sFMVvneL6+F5IvPj3rdHXp0D/uJwpLM7Oqwzw7zUxVxcyDzQKs6jQ5DPt/mLLDZcIGU
xwig872gkVksZpjGDchYy4u0SiqgBXsZOfpCAKHC3cO/xOV9bAxoOIVy+NgZ5nHhpyzd0n+hDmOP
nQ8O0ro341rZvOEHWzxkLb44TOUu6OO+wWX0HebLS9Co0F2XDtSo5NQqCrU0BPIexufXN5tuUrj2
UEHs0ZpSSfCrcddfdzp5m0okWoabboAo0+TplWqHza9yrNuwaM7uIgYaj/ii2GRrzXM7o1AnWZZa
3WgJ//cmfibEFGIej6iKEP84reOAW5lqKKPujJfHcBoF+Y2XaGYX+16oWMdX+0lHrNeQGvz62gGc
Qw3/Pg+TKugI1bIccmY+Evte0AsGbTDfuXMxIKxBR2Vipb/D2Dz4sGYoWzXqqvNhColKlYnEMjT2
tIcYI2oT+qdqxhGQSEoxtPCNdAPxRS/SpBlG3ZBu8sq7kal9DuuQNtMaN+ltwCWx8S6dOGggJQ4p
fCZFYYjo8wQAHqmt7cxN0i/qPdV5zW7twQek4N/xZmzPidWcu+tUTg1tZLcIhOFWzGGOx4B62Li5
Q1pcHAsFGCXgFEkdHUUCvDE0grtnYn7i7tspie8O1CKajlqq5g6Aep8sXxnQu2bpOZ/V/c3UCfgO
f3dTsEWk14V2yeqNj/gHz03fVKLQLw/o0FCHJTyEhADAZiYx1lPpxgkXL8Bs1nZoFifeQSVfhzsE
c4j68McLRhmFgrZ16Ogh0S788sDTTJ9+dpgR8rsMFZsT0gwRzsDrGxjXGztE9wVQnRwkwixtgfAB
Kh5fp8GFwBuQ1bV+18IrLB0qZP0KErBVJBaNidtdPpgHnps1YfeFGQ8/bsFciW0YWn/f6E3jr7K/
HMbuZTAZ4X1ScmxVqxUPwDqoUAqNVWZxxO8jwknIm2OBm9jrZiFvl5R8sXjzLecu90SzWNQfu+WC
t8AUmNLIpPBfV8ZbWMAwluevgKt1yPuimhOCp9V8uaUGMbV1zeMKM3WWFdGih6iOFm9DzMZwwuxy
iBvGJJgpUukeYjLQBnlC7cbeJQ/A+1FJ5D0R9YivdTqt8oEVMZyY43P+peAH37D/k1nrmlXhkOE9
kIKM3PGWqKXLBkrEdDvdRorNUJ9noe+EeVSXnHiK52ZhJy0nBxUT2r5wYhmKwstqz7xklekTEbn7
bSaY7l0EAUf5JP61Q2wcoL46S2nwT/0JHHH+N0pc9u+Ermg6j2B6VzzrbooPRYu6Mq3bfOWDAFoE
qpA+zp7b1uao6sd+UYiN/E96lE1jHUu151RLZe9l6kJSbuaDQ+lF6UgboT1GvYVvF8x7XZbGg1Il
rNWy1SPTejLhz5YpxqYcO1SPeXkNe5v8/3t1FI4xKC3STT4NsC0QWZXt8epcsA4Pz/cdh6nywGZo
NlYTKVCDoUbsBg5isvDEzisG7bbPfobthrLNPvC0c1s6FZrQQEuJYLanD6xbzgv4S0i9iK0xfr7C
HaLl5j63Tk4NA73JH0l1bxAROAAb3SxjnxwhEIu+RhNXjG2EhWy8hshcvPFatLX4MIcdAu0uBJaM
aOF02CVZVd5hOtkplPWLdK2Om1K0oxYB8ZnddHe+DJrwe6zsUq0nrYVkYFWznynvCXirdSP28Enl
vOvZjZur1YaY56UgAMsdgAMkYpfwgtLv4h7LMkO8RqMkj+P8xWtTV7mFjAp/4SXGdhATIVRnU1ui
yGorQ17Pyz/bT5MNvZWx2nPvMLolpGIiQWuqavcLBCGVvDBxAJ87bQa/mQLbtMy40uYR9mEOE5yJ
DshwLm4JNSzdWqp99EKpznOvsnzK/OoAThRf+MHlyi6W6zpDnqDhIWL9H7MrdcTeNXivTqhjTRHj
1UDFgdWwG8YEgY5/fYNa3UWa5aU2JXMWuqlbky896uRoIpilEusrw78kNV8gL924+v8I2ZMyq1nH
lOZjj3fU0EWfmBrb6RTTQ+y7f0++EVc0PQF/5ecfBjNBaVk+RZjFQM6roUHHES7NJmpixIWE1DFU
7wfPCK2O8ihRc01ja2vmLB5JDb7oQzbmMpPaPduG2PKBel1boRAiIiJbmZreiFbiFc7rFnyIIENs
DjOZptAoe6n9ZEgqAkArnqEZoJNMNzJKCgYpxcBdPSKw7s2q0EZSLL5B62PBSi+sevqDAHjNlC3o
/uM2LIUnSwrygH5W+DAkntdy5sROrnVmsL+REJkYIj92757oF5MbNxF1+nEHPOtORkCbQwowfHiT
pbYuq4+GwuPh6B0wO9RTXKGbufzeVMKxdCe6pZP1E7D6zgvzC6X0BQY6PjsM1jmjE7Y9UlWogFi0
t2cwGy61E/aTCI9PsR5uE1Vx6BOa6flf81CyJkaCrgbgvYHy6RZmIsZase8uo/+gXJgNm/jNwgho
AlJLh4hbsMFzJqMYlJF2ZU1wZ1I19Cqpgi1ZK1HyjWozkoJZ8EFS8AimJS8l93BRMP15TNB4G+T4
vHmIKUZfTL3YnHhbYZ9NrfsMqghd+uioI72YSsrPdXosbW8kKGAOMZ0+Nqt3zxOh8daf2hx92a5v
vb64XXNvKTvY7lzDG8l4MMUmZ+m75th/2pl4lRRm7nxUu3vBINXitHKYlHiMpwJff+t21dGzoX2e
09AV3whGIwdLUhBC20FCHsBLZPAd8DWfwm5FdjbiSk8HuzaUcwyUwhFvk+2dJmBePy7Fc2T/Dt8q
awulyH6YcgRxyNP96pRaRqkVwh9LrvOHjekSmiWh2mfvCJnTQUOFwTuAXn7BvOmDazSP6HV83yoI
ZhN2Pf4z4d2tt6y9zg+JYwx9awVAITY9miUa8j13sOM/PCD5ucCBvUBAFAklV9z7ghqaJ9Nme0VB
yM6WNyEfQ5tlY4J2M0+HM5WK7288cRGoSQauleLAQKB9zO3+xFWqeNV+uRD25WK4e/mLGJhYL+cN
XCoXKtTB658AnfgGdcgsUd9zyon2z0Rv3uDoJqTQApbDdEpZnf7kT4T8aTVEHICAqN31M/4wtQ27
KUPbNawluhSUWv8hK7SKHTsOD+tZZJERqnS0BcUs6X4eT97lBhNHVS7B6ctBRRLQgTl6+cTZg0qH
k8PTC15dbxiNa1s7eSKEg0+1WPp2BLqXf3w0Qm1+WyAROdFGlVBUS0vM8Q06GSxdFsbXx5GfydUK
PN05k7jIAcOOBmpBgy9rsRa0z7uL5zGsSyniUG5pH+rDddBM6QqWwMYxLfuk//tWE5Nl3jheUnnW
vTtaxfYaGq+N8Uxe38NhkrMcc465e2rhfAHx9TCpPkt6Y7sGx3rB4efAhyPXetJIOa8s7J99pRvw
5Pe5g1ddz88Rf/S5K83gU5cgKUrnUo33hVEA0gL/+qLVuXqOqThFzLtb2oFUoRYONqKqyFK0mu2n
VR507/GUd2vpjuUPG4rwyeZixNClsx8aoVZsYETTK34/7IQRYAQKqRdwAh1W1fXEuCTMVku6jhQe
WDe0oC2r8MktwpAKNIgFm27R7sopjXtOQAkBdm07XmrQ56HNh/UHmoWphkVZ1qJGKrMH0FDCXZLy
2hqteBKs3DPs00dFaKDCeoH8gQOymvs0HkyFpCDR3rAVoDkl3Yg+4CmnoYqnMndG6wZCWuexWw6S
1HMB88qoChdV+25KMFtuVzhGE6F12ugfUilf7Xtt+l3Vjr7dcVZUQAiUn+hH8C9ihXLCONQGHqKg
XzZnj+SHQrrto6CjMnp/bvXH3DyLsK08OOWWBShwpCRAsb1e8vrg2B8XyKm2i8sCdV4IPmCdYesf
IXbUuqmfOmtM0PLIESZbEAro83l3Xynf8mgnbeE/kxd9ns0QtsgpWyTElQURoNJSB4SSP1FgUSSF
PIIqO54g+sOtl9PgtcWOmPHS9JEBG73a/mecqusLTIBmmvkWuzmYJF1DYy0Z95mXjiFhhKBKuO1O
UnkYFtjFwnMppl8CM3V0d4sPqJQoE2TUKQ7DKvLUF/ARrinH+DqLxZJoeQ8py7UQr8TDzQEf7czu
GCC/bSiqFcO8DOlHV1IFMsB+VqPYYJvDZyjwLAFEyjXoW9MypP2nhjyNcbv+eaQqBofTcqL0zwTx
SPk359PdmtTIoxKfp4X3SZamZVTpitrIIifptXEUo2fCwQXlLL0ysvrNKRQzmKsj4fUPJpCOx/m8
BnRZzKC3CK7Mz5smqcnU0THZT2JORWvm3LRtQz0V9pAQM1KZheXCINfjwLu3IVB12Vj8edc5x2qV
Er/ddFimFPXSXmZHti5kHM7hul202J3iK5iXf4IVZ6zqwMyCGcB2re6t7vfAF3GgN4RM2+k3Hzj6
eCrWN3Yg+WwQJxSWrgEa6QkCYhiD5giGp/zHnOKorWFbB3V9SMTGFFuowI/+yPzVPcnqZKMcA6HB
i40RzfhN00CxOL9KCmNKnU7+WfXqS6B1gMnp2OLacTnXvcgmmJKn49crtnEmvLA1f7H0bC/6qdQF
LgFeoTuH42vYKM1zE4CdZGGaTFKsFYe+zKeEtBLVPDusgOcZbeJg+zkhsRdlTegK+6DxpgFUzh8x
bxXd1a5tMQEd4H6Ot6f+5D3YpVk2WLLNIDgvUAd0Tsv4ooAMlpkaqPYpqXjIxds7RY9DkU3PGaNv
oe/RZxcQpKDQR5QXHi2efWnCFTYLt5ks7Bo468/7uM/A7G4OrQWxjLuPIbh9wP/l16ErZzMaST2l
nBB+g/zPbLYycfRMh3p/cuNhPo8NqY98FkT7DTfySjBsiJIfDPGcwNvpHAt7NvKaoGmUG7TE3IeL
T43lPaKVuJMTUNnvVrC8WHdjRu92ioWzd2QODSxzo3Yom/T+2uOkcbsi5iSwqzil/cmGagGSojgY
Wuf4K716mw3mBlrV515guazG6a6CNl0Tkt8wX9vlk9m593bbi2BhrRAm4FC5ds1zryM4yGz6MNQc
VGDUvbCWxruTZl82b+4ou0CWTObgtfCDhCu3vsWFrTE62UIHwwQqzQ0oOv4W/BwN+cy9Sz5mXvbt
zse/o/0FSHchJr5WkmRaa92uOWf2jbCT0N2KWYscTSEPK+e1yk58hBPNcVuqyr3Xhkb7aKUH3z3o
g/smiu8cLiS4bg6jyDsmct9Fn7yDn1qpKpM9RO17ae1OyXRwU5l3dxdChkciKHynKzJbumzA1F9b
Wi3gccI0RVFGv1XbQdlVo9sJv+/gl5DiQBfJ0JFCRdLLT7ulIgcLOLDasDWohyMcuHpwWijJ4xFk
3qYRz+uP8HRvRTZ6pO6oN4qQMXeVxUzU6LopzXIhibl9+TFKjZ7+BXOdOjhNk91k2tecfD4cPEAZ
DRUQhx7ksE8dav7Zup9YJ9CLwMGgoqlnUgTYjsqSWTXjbnUrYp+WnHPdTiO0c8TtfxgM7Lg4fS5g
cTy5vRmmPOckMYr/DV8yOLLymfDHwSq+mBfzeB/wZEQT4Dv9l0GQkHEJddlJzYVunO8oD6hyTGtU
fzxiggkJIs+1s3DWac8Ef1kZbDCfnHkm/B3liTD5NyAdFOaFBp+e1V9YCOBdS0M9VF8x/UW1xVsA
Jpv8Tf8yyUajvYgMDI7/Q22u95OMbwcVgzrmOIBFLtCzBRWfdkrXdty3BJsIyc+I2j1LVgtZ4arF
gh2TbhoS2aHBM5Cx10YLLFbBeLMkHqq1uRCPYgifQ9BbHB+8TVh9lC7wdupHy8Z2g23KCQD1tRYu
C7zgQpHojdNasR6I/NlGrlxf1ZM+3z7n1bnm5NH6pOZKPPw88PnbsIXO7PGx9b6oOJGwylmTEh6n
EfmwcWfnkJL+9A5lj/xkEmf/xEqL0RQ2bMWVFfTktQ2M2BwqNv9NA5vqp0+nwPWs/MiaSOesz8H9
vQv+YX3x6Xz0qFqJD4bce+COn7hzQvZd1wqFK58DpO1AHuUhgb17ztWwNNLI96jWIrA8UCbfdVEe
tUBEeTNL9TyCD11JOAq39gjkWyHXvePnxRInFQ/ykwWevQ3uBLLvxHWzZUD9EghcoQipIRB9jNge
DM515ejeIZqnA1MDcaUx0fWnMYpALJ2ReKitlIsU5Ec3rgLkXi8DKuhIqwqlTMy3cyHdJURUZZ2D
6e1zPOnufb3BhtkbBQC6HHYn5Jss1ho1JaNIYMvDE6iQi76n/WTn/29sldEShyzHnbC9IEB3riit
IWevsk+D06hKxF777WDVRP/Av7eLPxP0PNvPtO+Kf5szmEgw+qzfRFr+7fhuCJ/f0efe/Mvj/qoF
w9VazydTCXd63e5n61Fn1YzaPTvUwRq2Xf6DAA1+CaLvYi0KBblxrqMERcPfI0iBbZB3j5NNX1DA
VU1GikBN876j0KIC0lYB7mvL/ZKSQRCX6F/pYVjAJjmxXxEOmlDUcgSY0UZkXMGPIWj0W29QfD6B
KRnL2Oxsp1Uf0VeKnEHqB6SXO0YtM6P7c5TZCUyFY8QWTy2DNpIR03A5NAPUCZni1vq0ZtyBmaL/
R/+U/QeS8SRMi0i8zB0jB3E4IJpHMLw8RJ70EDVSyAhalEdgVci+4NTRIKF2umpBje7awFQV8DqI
0qjE4XZ1vuNrR+cOERhl0fQiuD70Kd7K9KpD786Tw3w2JctCRTBXrhq47JMA7p+XDjOj3fSrUY4S
XTYd71sjYtl1J/o4D/F8uFJwT6Nxg7nWrorbVP2DGqzgmS6kjONEF9uqehgBP6ARbfLSjOHeZjFk
A0do7Z2tds23MGxulWN2iHCpRkQQeJ5HLGWLiUne+oCh6uCCtYPUCTpYtEzJT062JOqNkWekWwxR
buZF5S8TgV4jpehWHTq9HyWtq7d3bcIDSHms2rM8ngBePahJsiN4M5mwD5fHjZojCpzRi2THT4KL
Rx8vqujIsvXRdYWGip/IlBuV2tCfKF0SFFsfQajUB+cH66+lVMTlFYAePbsNRsXoPZtBJP02sb7E
5WyfOSEKXeG+p8OkYdBQn14VPuC6F5TcOj90pnw6pBSM05O4WmxycRGYEu4rrd2TaleNVdpswQh8
r1+guv4AMHmG1xKn7uvrYHw2r4EtADsiMOhEmYjVyM05rz2McJ3IOLhZfwpHAyJVobADk4SN6vOe
HaJobc6IkTkskqYHXXnLXn7TwKgVha6/FkClbkmp7YOBkGEyvjS516kUKxLfiiYZ9XtVOxv6J6v9
k9mPp6YWCzgpZZ7whJJSOxYygE6R0OfPZQCpdqWiGsCosWRq643owJkzUCO5yih7Tfqofr2K1n+j
+S9bu1hcwpwMpgjdq5iAh7WWWE+5bWXOn7uVBFzK801+3Ah0rNWgfWCxmBrgtWbcyXUOseQA8xnM
uNj2YNxcHjvwF83wLdfCaw9Q7dbxkBOnIfSe/zDrot8eeXcpXM3tuiASBmLslX7zDS7prw979XoD
vfq210ktcrJ4HE7AWbsmJkoqnr6Cypg+JgmxX9L/9Ux8gX20mwcWfAvAdZlG6QU7+Gc/ZVhcTPOy
6JaZA4DF2DcyzIDeuhQ5hBRR92PLjCQTXNKRoSlN/rstApLO1jEKx/S1vsUwmTOtRSKpBoA3myDg
rbbYUlvGGVSNkvjSthn/uDK4QfkNy2jzF8HiEdpj+k+gSni4XLxwnWVSbfReBZfE5EBcb3zmc3m3
dMdiOWG7roXp2hq7YrQ2Ii9QP9RxIfpW8UIVqVZvpunZX9ZlFPCCdYPyATGvw/8/iO5wL7Z1PP4e
A/FDAjnihjudESBrOepvkr5Rm+TbKpYPrJiGSIdpE0r8fltp8T5RuueSHMRt7tiX+Co2kwLLkEwc
jdKk5DFM3W1y9VrCpdxKHfiet0Px6ytyI3C8mxe25Rd8az7WnEjfsFGW9iploEQH5mztgMhadTRy
6mZU+YCkSeD5W7T7S9ZdwUK3SeAgkyTHr2d3oXBEQT467wLf0yyoyCLQmC1dejOpZxtPR9gsjCbo
VZpBSpfy8XSpmty6YRaYMkhuVMi2wTVPpyp+qV0CpUk/jBHllcebwygaB+pu+xVZY74M5DBHUkow
myiHWPt7bYF2Sd+e1/ytn1LO5X5Fx3jUEvhiIXDMMOC9ePyV7TSXTCmKaT80gQ0nXZJlS1t+6Ij3
S49bbwpSADjHVSV4P8iY8yAWTR6qjxoaIH36VH1NeIQvmcm+IdO2Eu4YmC12JlwhoLVT0Z9DY/cV
ZWcbhbpEfifCe63khHETShcR1L0Jc3/HF/VLirZke6PLBMBJUo2/l8Kj8MRChUpobBnwm7+fMt0u
Mq/zOL6OKMLn9rswWcL0pFYONpetXaqMh+Q/4TM7JBz6HM9QSAusAK48TeL0F2awbZvg2YdS05MT
MkP9OZ7fVe4yn3+iu/Vw6GBgb5RnHeHqkspvDDifkJ+W6qKA7kb+QrS88gWxlB321VmtGgMTkvYt
i01ga6PWuRxYLfru9YSTUWMgsxfAXiGqTdj0KYC+jQB+OuOYSlPUYLD4sUx3CSHFIAj9S79qL43e
u2qtiWCf4tlCBk2NI0yxx7nIjaWtIJpus/yIwLZbA0n8xF8X0PL17vGaEKCNB2jIHg+ItUpj3KKZ
xImQj8vw99++CSiQKWlWt+/Rpe0HMcyrIRRZKLjurZK8lsb38sE6Vj0u5x36YWmo8sOMSGG9AmHu
Fdj0JnHHs5QC9M2nOiZwo5+q0SbknOwrrzQQF5HewMUzU9k5qWdqxLpiU7UbOnDaYU7mPuXxy3L7
nNH1fLl373NRbs1HWnooz2CYOhd2EAyr3CgvGwzRzNwa9vVsz6Zg2GipvcYYc8G67+Iv2pDJJ5hV
mUStmTpqQtd9FJM4GhZaM+J3k6/j+ZCbtOc5PgN+SRpFCoEGEj5kGZTOzpAIht4cDabGLb+zJTbe
VRaaropnAKk3s378VvLxwk7sOgEPW3BuSUJMEzAX2mXt9+2jZvT3jZMTm1SSW6Va9fwLzi5a+v9a
Rz8j5COwLR/VGogDZ+L+V+uRPUpM6awmNl59HwPBqRbyLuOdhxSS389lXanJ2FXQ6Eb9j7TUNCYA
z/v7Un+CYv1PInVtTXu3/BpjA1ovpIv2IFw23QoWak9v7+JufeOlabxRksVeNQ895izbPwJMKmaA
PrS8bMdxnnDxHBYfeqrXJ09qqXINEnr4Jd6SvkPrCI1iQfr1d4EaPQuH11ksGFCVsAQ5/OHC6zAc
KJBj6qJojFUt4blSPmAHvAu5CF0XOcfZJ7QTnsudPjM5ssWgo5f5SaGuhDqVkG/7cpvA6c2sw77q
SvB7Z7OQ5SkggCuFyni96VeG78rKfDO1UtFVlSKqy0w5KLcBQ1QhfJTLf+a3iSrGOEhCdiTaX6N5
8N2Z8cE3hCRIMyaPQVAl35ZFaMbT7WRy3iouK3EbxoskmYneX52ZRh6RvnWSI5s3mWi6ThkKrIIc
fXwDxtTO/hLgT6pAE9q4TJynuVkUrCW1ABSt3a1a50RokmKlcUpN+pT+1m6kh0Y7v7tCjp+xV2Og
PJqX4/bE7/Q4k+w7dTjdtgqaJYY8L3UmiGd6CrVi0YMQTV3j3OZnyDwQB/o9f6lVH49ST/JR8yOC
FPzej05YKLWjbyUL/QqPA2v/C3ABhtpiutK/UrvtXY88IOxSLw2caJsuaYMnXZzylNyK2BwnhAFV
Vo+1SJIJpO6Zkn7epj6J7MEga8XAY5+4XZ2nby/ls+5vVhN8m70f+at1sSxDXzdjkptkJm4eVQ4c
kNppNKNgH1IlUHmOYMzi0wmcdHbdRC4HGB9/ef6Ep5UpJW8Ix020xE75OfdaiSm8/lUhiDLQNWXe
OuzVsWC4vb2KebIJywpow3ZVqdb2z3faXke8nZGa+6Hde6lVMA+BGdNZ4ntzDL4xJ4j9udVEJhTi
Rl3BJvvcRz3LJFi0gvXF550Ukt/ZjYgWzRJmwY93SZsXFZnVasXiOyZB+bCQv42qaSglTUSJpLCB
qSwy2QiAbo5LM5m3atnCC7+94jSw7bisiYvmoNXN/2Jz0ONn+fcJpQFCF+RkPRBVDL+C7ZHqZuuP
SrjFVS3KuwYPsPjYV9rcqh9gnrvgpWMRqG54IkrL0PE6FTE477nRzYdT4a0l4/J365mqiT2y4Q+5
ECgWWkMW8ciGQbDP4DzDrZHsyQCkjJwNaqMiCwGLt7MrKaU2KUHlHYAaH8vd4ioKIKAtVOKknT/k
T8Tatbur4CsdZIqsDSgIjM77EkvCeSeSSuDECP2eOSe6bCUcA6eOWOakq1bi2EJ5T78p3KY8gfva
2zgce8WQUcq/qYKvfX3zr8nDAQwhkW4PkMdI//80NKX8qusIGwhHirZvrhtRjCUeKBQVKfnVrruv
Y7YJjSFaTTJ6jNL4QnxV7ChK8zkVzCZ/INPFiaKPzy3Tpos+pThoUwgEpFr00JN7T8zHATGLkfDS
3I72apJETPgsmciSBTUlrmNfTkhZjfVV3iNRjzRQd8ZghnVxTyY/WZ9H31su+6wSY/0MwJeLLz3O
Tyb+R5qN9TnkNps+FglU1j9/VgwPZ07nFj/n8aOO+ofUll98q6DR6qC8UoLXSBU/iEML/cZhP4s3
xaJ7t4CZzTiMB+2dY3mvY6MRbqDUJK8hdm602a90PjtkUPvn+nEqL/juAONDu5dxjnR0qWse/95Q
WFK7KNzmgBtmIEUOjyd+RfIa40binEWVG9+XRYHRUwzuPQv/5KsJgv1z/Qk28kIub/1mcDmuU0eb
WBPk1OAKsH6ImWyy9dwQZEAL8UG+PJI47vTgtLCfW2zB0T1QJvImjagRoQzY/9InpxHlKi/pkgsG
0L8aAXE8Tb/BvqXCn5wCcPHgXe3rhDdNSz1BttSDYfU5EyUt+kJplTC/WgefbprONqyuO02V90Ch
eaXTdmC5BNCLBYGhjm7xQPObRBr86R1fBSVNN8CzjomkjzjzZ8/kZuCy/ySWfMxS2FgLjMU8E4g1
MF+PE5bkglW9F7pjYHRDdEnlJ/qvbrurCx+4zS7axqT1yqcuICAOs4a14rLN+BX5UccSx7niuBVB
0xGaOhNFIzwVI2wFxYy1MnAu+NPCaxxqOf7iLl3iYhKvaJ4qKhPWpWyWk73VhEk2CxSNBpcDFf+F
glRjg+p49usLZNUQ++9b4rxCQKfSI+Ro8Fk2vKtYE7ns0rbt7LrElk0fCkfiNm/IFPgJ+cgzIPdq
5pz9mZ8AE0ssnR/j3aMJNfP8I47BDAY/U2/+E6QqJ/4keVWBAWPTBfho5WiLxTMrTdetiZqshUJY
qyD2RirW6+Lur5vkwsADbVSHocyfsYqo5+ZQSj/NopeVnTB8x4HhNLo7XP/ZcAQ/qL/29hnd1JR6
B37SQLOAtxFdvSHmmlsWxdx8hokBpN1NWbjgQpXPb/8TSX4aPeoeMcSDDJHJnAwEKs0nwTf4Skxj
UC4q7A5TvVhlBDg+bhm4ohUlQmK7BBKoY+P6aLh4A41HS9MPOnxJeG0aZo6YaYVVxiGn5gyDra2+
SkLD53fw7N7nP7BIq66gumwr7wj/l6IYnuuJjw0nmFv5sOmb6pOUUSGlSpOdTj1u69lpsS8uM720
rGZ1Dv4gHlwPdyMtOI3SHKIiIPwgrNPdIw3vMcrC7BT9ut9AY0gVbXLRtib+mJRjY8jUzEHMzTz6
DF9CRZD2ASIq+ckTYT9gZjqAk+MTUHk9S9m30CElDCbV0GbIfNCPso0TL8Ufm9sTY7Uxsda9er74
n6tF/+fu8/8fvuDZ+YVGa/U0LwbhaU1aOrSeZTtV30GqiLoBkxOcee1/9Eo+qBlXjtMMp/8ycvBY
JqIuPygzcNbayYLjzdngvxLFmL1cQTC+/btYsU8suBUT19MJLRmoDj1IDtgjAkb3qzjAdCTrZUmm
DzdKa72lh3UqyOQsJAY+p3uy0Qd5bNqzS6Cajg9CBiAawHvNQL6YBlEkEOlnw2xNIesL6qlXzlG7
HLi0Le2TYuPM2J8jBzQZGitqcrYet+PzWVQzPhkCsoCK22casgvp6qY6MhuCREOPQejAMyrwg7Vw
2a3MZnNDVdU3H7xvuJA5YnNcz19v/KJpSnPORxPPYsjuAJ0g6Xv4sQdb6rOpsJIQShI6XEJ1Sm1i
rriEohSk01JCN0QRU0LN2WO8ps24VlVC+gv0t26625177tqNyNnf1hPgLMpzt7ciPjng3iAv5uiD
i6xQapliSBL7SO8UGTuoydfEKkUxdqYnLiwm8bWDvlFETBC1x2wnZC4ZLQKMPTG428tZ2epncyu3
X9BvUPEE5vSDm23G8Ruk418wEHHOGHj7lUiqnYAe+tykQvw5EX07pQ0p9sdwO9aTnUZ0dg23dcBe
HJyYxsu3BRTwf8jTUs+r5ExLXdsDfz1YmLPmHmyEFUs8jR4NnIWNU6oliNmSyR3FCxLswb4U/XlN
U1uD7uc6eQaGXhv3EKJn8H2gFGDsVq3ltZdBJzbOU2eD/k5AqXXQHR6iuywbXO3doe36Y4acS5RO
ZmHOCyBknEXmA4q1GFOrELGt/eCitDBDpU0fUX1HSH8iIazbnmcUk1DXoWGVQswYgOViGodD/ZoU
sCHUJ0e2SjL5ONI/M6KPzM8f4we5Gq4qnAtCgfeBEAL8xm/VF4I0OlL4XVC42Wudm9yLNF+YXdKM
2k7zj5fchyqDn82G30RrtMha9sluX/0aeAPt6yK6VFSN+ZApJe7qyPJhTrJ4fYhVcuO9iAeKsbSJ
mOdEgixz1K4K5+9eZmkJIemoRvEXHbBlROP7Hsk3YCaz+W3/zigwbVkcJi+uwxjvt6hGEzZWE1Gd
1pwbhwlWF0PPMGeAjWJtIUFIGWVajBIDkdWngwe4vep2F6p6nPC9RJer3NiB3a00ZTGiDxUKJ/vi
hudEa20+Ye82n+XOz8qwczmUiJJCFE4vZfPS0gaVL3QVpjnjDhrGfXWfo47ZJ4BCl4wTzv+xyHJA
6uvTf9+9PscGYBttL4D9KcZp9rnJ3GI5Eh9Wnu7lLd8q50K4tDIfUpGckWPzDIYiWDCyvonP/8q4
phC3G1RiuwvD6sGZU2gG+YxiSl1PuFwnDcoacFntSugpEUgR5lE6/Ap1YEmlMivFLw9I9ec7XvKH
pegmQPWEP8JSXLHh79O9A5aUqloIS1J40fDz5btGbCxqbr9w4Znj+f/zYHsObSD8qapO5/O2h8dP
eUl8A7g7FKFu8Suug5GJJx8ySNdxEn/c/n4XRWHQO5aXMzKRCRkNl3z2GN3zq+8wonz7yhkr6aVx
/k+vMpRUSjD4wfYiB/JaBJ7zla5zYWRKh1jfbBtjkn3QoP2wEj/cWAIzLq/JhHe1aMXnI2w2n6Jg
u/1Flv9Jm/lCwA22unxHj4wHusLWFRb0/bIB0IXt0mPgzRD+VlIs3MraKNapXTgkI6n+EzoGWXk5
+h8XgdfuZfb/hmUqSHAXXaWvO+R0739/awHSvPb4wnUCinqYI6B0XmFdeHvw2BZZS8pho8WgSeYP
//ke7QF5nZi2Zow54+e1Ebf36MH8rV35xraR40OlIr87u91RphoWwRbzolZhq90AYKKsqy1HJjJ8
KDijgmuPCm/M2m9E7wu5M5n1KNXDmm/fH2tjEPxdaXmoAqxgPDFG+ws7mc1Nk2gHObPBvswCJK15
0R/qqZ8WQgh18oQh5P+otMGWwdeMapJUFw0AM2qAyRAMxhj6AVTkVztPPLkteFTiapnmy+mhuD9+
Ca5yEvrQ5SaGPQESnEBdX3CFuFmFAVIQsXMGMXGnX1ruvV648XfPlAWdHpEFuEZWiUU6AROrlLxa
xUAQ/oIiDUfxCRqQaBZg2GmQITP7f5wLz/bJXuWeTDI9jznXtEHMaFLMRRWgjHXo8xlWhZO2bJkZ
/8kmvFjhmJUjxzIRijQG061rfipsWqRCbcAI3oqZ4nNpWA70jclbKQ3YCovCfTt1/YQToknWCN4+
/Ik+Jj/0GQvcLUytHpd0Ls5ByVjFCkiuwvxtWI5q/hS4Fao+i5sxO/eZAGbm1vZbR8B5QUMAObLN
cddGcIv1mSiVlEJZrmyPB6vH70clRY7DmDiYc+OYo6h9ek02xce2fkkBVszmiBqlfi5YLZ6kmMNH
wk4TpNdXUe1ZxFZrgK+MY5elBp0BljhKo3zPwd4gKsfStwTJFFHggAbc9VRmHFCMwSMMWbr+2apD
cUTTorMYvL7jEaDmYK8Mn7Oi0sKDHSgSB2YIUHBaYElUwIcwU0D49f5N4YGcvccnAt2sdTWD068q
cMzufQZBG/V0g+EYxr4xA6I/47OoPF2JAiYvgOcPNqVCTKvz7S29sC3jOTGhHrozJNRbQ47LRDik
BcdxcyW/AtM9FTgD4Qy6oQlc8obebeo0+TFXjoUAw7eEADRocOmrzF5X2+W5lqO7nNQOcQxpWmll
Oai5obWEi5jpQ0MStQt2QDbDGBvFLHM1DG4osFckjL4aWJM0a9SfsFsP9sVbn5ZUwtJCaCtqAdYt
LIe7H50Ahs5kpJquexBzsnS1Z7+fjKOQEz6boCJMTuGXbNQ8rz5RYDhf2JcmZ0gU/HPldGPSuyU/
wp1bDhWi95kkjnK9BubAzIe4Y1gysFm6uSPZthVSxWXPAQvvb7509ZvgwkCtnJoZvx/l6KBvX1AK
aVKOmZ4yGyHVif706OYPIrQ78h5Z5cS+bZgca4KWD2HUGt+2mDKulYtgInlfYbbrmndLOj3Mbhnn
9iAsm0QRlqCcMO26mBjkHqcY6vpfyrt4WXIPjW51ETtAMIhl235oN9ayA/PsbmeAO9Z3jmECqwz4
uGey4VdWaSEJXQubvv8Kd1AZpMi/3mvw4j1cOQsUxpSFCWC+I3lMYqutO4B9xoOwlJ8LsS2wTGAs
5uqLRMAOg1bsGlYHyx9VDRjn1DBqcKN0PgqyeOPSh45vQGMlUGDUFpn3OJUCZRWillId/yBR3jrj
WTzWFcH8N165ayX/yjBNM2Q5rity/anhImVJ52bsa83IXgeJUfLLmJfVkmScu1EZOR70m+93LtFz
lVrDVrLvEH7DZ8JVSMl1yMTlhHrsZ0+F9hLCEDhRu1o/qJo3BUx8tA91XhaTAW+VWNnwp5GaMoqj
p+NX+qe17Zp9K6BB8KpgEFTKZmPbHwZ7vSvFYxniwyrwzVRTVj9ZDt1vYnpNo1MXHs/6ga14SpMH
3LBlRTXttu8zlnJZdi+X3OgWh2xW8+A60ZjrLxqc5sza8RVL906v09Z64mWMIAi7KqRT+IYqYSEe
mZdVva1afv8OEbBh43IcuoL8m95ekiDfemVsRw9+xEtWVpLjSCh0ok8BfymotOHv3+EVnYxAmQHN
wGAZIKbg8BSiPYPvOk4v9Rc5F/B2PCjoxm3yaGinML6OjibFwYluU+muM+E8ab/4CUOO0B+NK8Wb
JAAhqX0g5+hjfsVpILeWkCkGIpGyOGJQo+sqnzs2ttAFDRdkbebTdVH0+cI2Yya/jZR12pjb4xSU
2zuEyg1rpxbnht+pidSNimwfD3bnp/SmqQW9NOucX2cLf8vUrI3wsvNB1ZtqgnV03M223yYoSg29
pcIzP+DlXUz7bOAw1iOtH6nYNeGqJan/WJUjlpVVOkSlFC0RrTD7Nmqg4iZjJ5oQNLffIIfUnXaJ
7AYG219tQEjxWH3eHhctOHqWxqRi1AtdoEPLpytkR4ugzUgIbH47WIyKgHFDvaCKnuDKgy9deyzN
7Xt1fVVEGD0cAJZm84Kz9LTLmzFYPn4Tw9Cs6rygNxel7TEW5jJ6gCJgqrsP8UkjFaDBaWwMJwYY
FOzUOo1kcHi9tlp5VyZIYr0ghE7fM4qgAM/QNe1g6jf+plNv87IMZnMSddCmxvO80LqfFgtgmsBB
9v3/MLyc86becwLBp3ynQxsfs/UkkToUoMNuHzKe9yf5OA46Operzo+lR8M8hF2nWlCjiG2IE9nI
p4ioq75Gavf3T6+Y66vYRrQC4PCFMw7AmrnA+Msdx69aAWWDITnOIPBHmBp8ifNKJDlTn8e+gZTp
i+82tfHhKbZtcQwBg42FFJlX9pq/+WvEP7H6Jf+yMu54XXp6GW48LoII7L/v8AgQc+2oWZawMP5g
5JxjqMxY5/kQgMnWhyhRv5Ra9K34PkSAyGenJOCb6U6CKI1uTkPTam/GGKCNew9G06ujcYenzNhz
APbVmV8yZNz7mxhn5LHV8lecmLheSwDFjRjp1VBe6RELiTTqz7ud/1jWmqmzzWsSRAHVmHSr/VyG
7/OWiw8PhvTBqECBlXvvHDLr7gEmEy0S1+BmzSN2oxSqQS8h2oyg5ZjQ5YOkEzQ3Nz8yQ4O/wBJi
QdB0RXTtMqTM0+Pm+cAgiD9gyXCgWsWEpM8/TWvW1SNpdzZy46cqSdd5KNyDjX2PAAy/8DlPiYPv
Ms0G+09cWcWrgBvuK+bHBx4sBdkrQA0bABUc/cJ5pdKWHzqC8QSR93Udv5yCXunCrgngXpo9J07p
jSjhln8rhgbTFbDu03IRPEFuwZ5gIOCecKhGmemoQeWvF05u5O70MPczkM7s8MkoeJPVCTkSTf8s
ppYNtbPdVU9O0KJzc2x9PmJPaZbyvVWkFKSEOvqUWkl1w2tANaaL7O5GNik0jZv9Wx4hEZycSODp
8nNHTftHzOQvThrkVcZ6vET51pFZaHGoMJPpYz13e1m/Cikda9tswdSajdaS8Q7hUk+EYgGAS14M
vrKiiWD2hzToSjG17vRHQib1nnlXzjrEFTQNdIzumtw9r8NC7u6ZyoubbEXvngpcaQcURbh0fIRq
p9w6qdPumu8yYIg4QNH8+YutTx8Kuy/Om3Wy9XrXxzhURAGbrylJ/R1BZLKvodktA4sg5Fxkh1sS
pijNSaa6fVgc6JR5jeg2ilMljPjZ0ZddR9wLfhDGypel9rObOG9VvtBVrK+dKHa2dSC8Zc79BwX7
zskZod2Zg7iKogg52gS46Lv18dF5pqsfHm5y2HonK1gegl0XM8U7b/bPdr2kReZMOs40cHl7z6pM
hjD5k4t8iHY143YYOICVNCTsdfC74tHvnS2M+02TTHq59FbD3QdBARHhho7dUW7vkczTfEqcuXNN
3dUQFFEstuXB5Q79tt+BIQX7LyH+2UEGXTqHAxzXHN/pZmlbyXNQ5cFuT4wUp/SPJY51p1h38Moj
rgTh1h7BgyKRgotJxwSYEUVP8lM1JJTikjgbTfEVtD7SMpdXSh8aqmhjfSI3M4ipblkoWzqyjfOl
HYp66/ZTUkXT/3EZCPaVNj1puXRPrzfi5OZ66Hl+6ASPAd2zpPedbipDneZU2hQtMzFBt3WrV7ik
L1G3S9Nntx3G0KM59UjW1gIrL9opdrlcGU3TPCohcVpJASqiGFmt0z8/8A5lrpXY+ncKoIflums8
whQm+7unCBTRQs1vBWI6T18+ZV40PvqShGtD6kr/x2yAb6KNInH+SIu1ugQEzMRGsc0M69VZzG0+
II+/QgdI+FY/YUpOXDNOaDtN6qQh9nAVH/fpzSKHGCJKeuAv2OyFICQOzaRAdPyCyhKKcEHYFR7x
fh3qZDyHR0ow2y1COwyaioyg7Khe+I30dfaLqPjCa0stppQaIM0utyz95rpBqpaBHjs01jkGdxvR
K6VZWB7+8yAlABBCGQmhweKBg9Im+iGWzzxq9s/EQL8qlhBRVM51axlUzdqgFPywXl14tbcgXmX7
zxdBAHyf85JNbpNSH3qyN941MR5gPecxNa0UEf7KI+hHcRNKU7+p3NSgV12l7iOpJzOH8LdvKU2N
uNmhvGno3R6TNiX64mZFhwyL1jyDFxtxI8fX3s7JWyy+CteFX9O2d0+NoMGXp/7ZBIoLVDoZQvFK
8pfA7U72eE50DE5Z62/PuM3fFl/z+zRtmNFVYS84tFhPaVoZfgA40xPiSPXwrtkaJVHKS1Bd33W4
R1PMsnMhoaZh1TYxCaqrCFWar8PYBp7KBPVrfZcMpqa+BITD39mO7+E+FGSSx/pKGE3pF/qbUer+
wv2Zv7JWUFybyTn7VH6lWe3nFPyC7dcVDv3W65T1z0j0zVxspyadXRaOAS47CquTRTT4hZRHZYNl
fSx5pY71INyS6COan7vGXZgaZt16c7kdQFd8QgMjNh7phgmZn2BSAoKyhW1hA36927/dv28toOWt
A75GOx7qPp9vGD9QzZX8PZ4hVSKTuZU6aoZGr1lfIuj+ojTnnQukUFhISV+ILBJsX8q0i4Bm/hy4
G1jZOo4acBc8SOFvk33RyRTl2K58P7hp210/I58xoGn0gXvG3lU3vbRMK0neESxDcr62tvwXkhAK
Zh16vauTlw7FHVTIXOjGtb6n06fJ1iy2CleIG6YG2hpNx+ocPV5x0159VtfpHe0wRbGijZbSlkKQ
lAJfh2kC2IdEEOSlhMMKgM2FSeNLeuPzluTNv8R4iMxlF7Bggb1sIJaHyjunpa5eEodCPJAqvt1+
6Vn4pzXWZThavyYSuBL3rgfcpLbVAVnPbRYHrmuJFdMRafsd7/tQvQe/fs5oY6EWL5SjkpJfC7My
vDlS2h6k0uSaXl5qHTGywwEAPmK1bYRYJP/pxyMxA15uTf4mnXoNcowLjg4IBhgwZ9B/utEQiVMM
uam5CpGAStW1D7CydB7pl9HHI+iEbIpPlCXVcGQpZ0wViEd/CxtUZTZ62OjTpH6Y8KYE7rKLYqfP
9Ut8qQUwfUos5JFuN98px4h8Edn+SqfShZ4Swv/GQxDn59WeswEmZtoA+ENMIwKwR9abZfhQ+5L+
VFBvqLpkjbSlZ+JkrqoJXr6te1Wjeswg4T5G4OG6PxuUyjUOPcJyqP3yn1AiPXpXwOMpz0ZwJkst
X5q9xUR6czIG1mrLOHTAAj+jZYQdFAzrbNShtx5OA0PaAd70vzpqSAugUQKrDg94GfmM3M5T7r8v
7qF53rJtypmi7B+HN/8hPECNz9C1FmPqoFoBU7DfC1I6GjVw1lx0A73VO04vb/q1GGPbg1H6RATu
0hit8oM+m+jfygcOVz5GwQq56mLCQjaQsRpSt9CyMjf6eqjyCK38p8W31fwi84gk1/4KAvZ46cL8
2CWD/fMK8/715ksWMe5O1JmRWUyG91yy1Of8xurCcMF1UcXpRIdOiF5cJIMctLkfPcUbMbo0xlR3
iuxLK1K9SNeh7Qlsu71+KayZ7zeAMu2J5UrjNhbZH5AxsQkDLZA3nl690PhR1tJZ7Y/tapZg9m2g
ZN5k81CKOK2H3YKCCfkDHlkD3CrQbpJ9ZufSrMjrvSWIMcN/W5r8Rf48C4UZYAMgK4WHQWjMqjrk
MWR72+yl1tAVXptJocTYBPVCrairn20J4Qg1J6TlPmnMN/Pzn9irj8vRaBOXC3F5rbi5FO3993pN
YLR1wXVJMk7Mnb4Ls8/NYf7Wa3LzZIjKhV/oFuxPb+z5iDnRY9jaDHFr/RhCjYd1mXCdd5tkC72R
+Z6gkc1rRMq1TDKV27BdtqnIvhLdeqxGo1SxqKfuOAShXrsP3j0aOrZgyDcdxHNcacN/BpKRI5mU
puPgjPmaGbMH3Kk2+koKt/A19StVBaMyEuRfjzBYDK6bu3z/b17TajPWK1MbxncYpvmj/QgHF9y+
tY1SNJoH/qcHgA4nqfzQL+q8WMU4xSGe2TD8+wQmWapy3+mkXR5g/+p1ibshhjx6QcIq4Jy5FHlc
zDrrH28QgbXRQtKdXUDpet7h+kzJ0iKQammpZgngtzH+CHfunxTuVP0CzTPQd1qCJbKF1ikodBU6
HnKvsSf1swRAo39ur/KAHHFwJobgKtxxFpnFuCWPuwLW+W8oLI4PPgtkis00mvY7PhzdZ/SY+o8E
a03fjjbr1EvhkhhA5Cj/q9t7jfpcuXJF5aYx6arK+b+xhQMB+dHaqtFk1TUFlxj0IlDIRwOpFkI+
P9IJz9UYbSd0A6gFmv9TXXl3ZnsrBrJUyKowVqiZy/VtNkbMDoGif8xOPe9NNqnBSFrql8d04xOw
ceujgp4X8rxQiJY2RmObeCco6ss3AJKuhsDLupHo6Ba+Xc3yFZh0D//TvEmNfmLwt44z/Bj5q36B
HRD5AgpFsR6q0ugjMr7DqeXeW7pOZ/m+IQd+Rkc2fGraqgd2yC4XTBg/Fp1YkCrlaXtvwnNh2qwe
Ckuw1DiFlC06eckK7t2CKZOuFTGaYZbop3o1aE4g+Wh3g4GaIUNYIXSDZ2DI8/7d3YyVXLESMUJH
ALcftpcgXt6597RjICTlWhIIUbxtfJslF2wNFLAWQVJ4m4lpJC9H0VNwTGAC0HrtcO3C01dqHzz/
Fx5AIMvQg+qdZmg46RC5lxObYnbFRe2Rb92dgr/4XIFUlzvWeLaXtpjXMGMr075t+U3K7cWK8Wpn
9j7sJnBGFY964Vmvk6yDC4gZSZ1p6hoBGrejL3ufU2uU4MP+FCWnMWn4+csRuzVhp5hPLuei7o/v
HX27WtPfzCma6yBkdEeqCMM57MHw4yZOI85QurFebKVs6Qd31gM/gDj9RHP1XsPfMf02IIepXqM2
Mfypped0w8a2ZVMOkepS/aGK9uW/YqP4AA9ZrvFK08fE8lRlrT2HBrHBQ5ZH6vks+MU7hCLQ0wN9
OlI/QjsR0C7/NIX0DH/JZj8UrwfxsCeVvqZ3dEYxpiw8zmw0BG8ACVfZjhu6aF2SowdCXvSvSYih
Pc0bwohl13Jdc1UmE8rQKVwGJevLdYPBlXs4UB4Fz20Bp5UwTmH7o0R3wV0Z9LWHUW6fv4H0iQDP
l+33nQWp+p6hr97wgWvaYeWGHajLxK/Ol07plVGoulHDgZWuktJt9nh3WGCb8ZW2pTSmU/s8ktNE
/mXnEnc9bPiXv9NLVxSpe8a49VNYv+VkI5S8P/OpOX64sMYF5ZdVdcGTZiRy2sD2C4IV7GaxYs+Q
zAexsm7c2ueURQkCLc0aup5fe0M7fBs/yqO//XGMjkgaN25Creyj9G7y/dtXEKU9nLKL0nPTBYWZ
ICRfhKx8Ftn+kOblKyvUU5/rwBxfnU4335FF0jlIl8N9gMgDigi+UCznIOFU+L5ahA7pD+2bxzS/
qNmObNoHw2xPayZ/TzjYLwyvQnj+lG/UK9SLM9o0Y/IpXKYPKaXcwYhJrV8KfVzuL2RkTZOHDR3p
vNMmD+LCMmoCzdQDej7nH2rcw3JOLSx9k6TkCThQwtX8JAOq93Hf6lxhPXToUhwh0H3WLf9Qva14
xRwr19sfaYA24AhamyL0puU3a4bzfQFKG7D0yepgVc5zvA1OUOjYiB2sH6bXWW9xcBSUPhEf3Yph
+B4yU7F4n7x3pf6XxnkmUX/KMjfof4AfH251L7yDZ0s0MqpqXfPG0+aJx8Rxgy5okUnGvl3leHyJ
I2ED0pF3EYTxfDWmNPpasl5LevsEO2UjONS4oRXihw4GnR8dyPBU6UMABs4LQDbPmjdgIGNSWP2U
iS7aEhvciMSRc9rraVnDsPAqXvnrOLHddIuclbH6w2NX2mynXwAWHky9Jm9G7KgzIWHUX0/wn5eh
OYqfNKfd8SwmbK3KAjVkG9HxbdkbXP213RNnNg5Tjuhj9gFANVwOCL6+nSD4zrkIlHeUBvuMwTww
m/swogUyqO3dO3cj+rVQXzZUgxHR9PMR3h76KAMjos76xCW0Pmaeqjlkdm1VygYALdnd70XRBNKh
ScZMGPql/egUlMUqGZtzB/bqbFJqHNVEKnofFoWkkjUuZRsC+d+RiCD3mvefOU4ksYz0p9Jakzoj
W/gy0BA6mfbvA/C3TbyAePjIzP1Su5gTIHXOeABP9WrsD5x/F6SZH3bzI1yq0mLFV7L8LlQ0N4pP
GkxjHaZy/3qHX/ZoXTsNWYJD2eJHqWkhfQ2dasutecwC2SzJDbvN/Pl5oQeqyHhDxWvlcjFUrJDF
ak+xRHFa44cUzAyzPYvw0MqQFaR+lhgjeQ+5uPlFSuwlBccKjOmrLaetfwA+HN8GsWprzaf+woHC
rKkojCBRBWg4HVcHeFTp2Fc2fIwbjU+pRNZR6bQQvOeMBbKljMFxdQ6UOuLH8EUQQ+aGmwEuplOm
/UK8h9recubvA4K5Mwij5nE8cV3mbhegxF9cxApCdV4RPhMTDzv/1s37d+z/6E7dia3ZPfuTlwMg
Khk1sRnpcbeMlP4Bc29kFpeGadF4fXAvq6etQGW6fRwBAoDSB/r7Kk2UTDBaKoos0mU/8K+ekHes
uL727n14QNsAv1WP5CamO4nay5e+Dli8lh7NgPqvTcrZk9s2KNIG6S4tjic40P07SFUXtCFt4+C2
EIeUkIPZrA85pWPnI9FFFYUZ27R0DUs8H6O5e/EO0rOEMrl7GhJ2KdRLKJExi9ggkN50K7sMMYgm
YTilGWzD0vxXctZ3aTlqa+zTS0Zk4pgbZRbmuaew1wybim03OYyXqhGBwq7oNONkxAB17WOq+lHt
7ZuuBS9uZ+A2iuBJOnFxJ3BtGGVQVfkhlEbvUPaPchQ0xhnRF7hdi6B2OjmpkPWw8HMoYkEm6uL2
z/sniIEntjsWQjZUS+rq9unI+uOVRBOtcKOdZ7JhY/GZVxiy3l3iryZKOjDH1ihNcD7O6vac3a/D
kKF6o7mKwtvJzr9ViIt9zlR9zSqHO2TL6+MPJL2CnnS3df9IMUGjR5YawaX8mNGGS5Ce5s6mxtul
5Z5TYs/NjnheX3VgNkoPPoNtXuD1Xn5L9uKFoDh2H5sastOOvL4lAQqyzp17kbatVvQuahk7pO+f
OjTAh1yK65QHHYyYvfN4OX2DppRFKtiTma2CcCRistyTrgWlec/pZKY51ARJ7B9QD0fLHZnxSCnn
Wg9bicDTq/d5BRqVjh1OHHBsb5EnCvns6s4XOsEpsFpIrWAT2eq92fVJFzddXvkJdTAuiH0e1M8v
EJnawYDvImmX7XyTJBKQbnydrmgdepuwqKr/mT0SyldNFLt0tKEQ9pnthvdXk0CNRH5+YSYGP/3s
6Tgg8Ni94Bcpla/8/yJAjcliJhE4pkWoZZCTTTd0g+vAo7ioz1l9gyfNt1kvqO8dYa2P1zzNEoSg
VvJx0kZZyZchoZ/wk2wQEaYOmZT6G8T5F6mkuLK2pJXI62oj2pJ14D3Pzf5v3VZL2v3VPy+XrKia
Y1gpxjpO6Xpz+ESe1qiNrYsSQWoBznlwYDlVQb5JY5xOTVK13FHjxNEEMu1QT7Fh5wxExYEbsFGq
+j/TNRrHFxzRNSti8Ai/uD95RH0zd7WAHRoUR8Ue/HjW1DxiT0s5twneoUZnwCTh0H7oUa9K+lZi
59Ppkeg9XhHWXc+xMuhtHzmlagYbuBrhdPFcexr5TmhrVdTB8P5G0a7PARPjbrRrgJ3mgAe67d8H
tqFMlidHJMLYu9VnUtnHFmigGPTghaYr6YWMpAMarIVNPjtZse4CP2JYauQYV72W0E/Kf55E7yL3
Gf3u0DYA2GkokmST/nV8K3Vz32Wvr2FkaBSKyNKT1+3AqJHl2NRxmHJkuOyqLUNjSnBijacFh1vS
MoH404uk5libzrbU6XmABzHGcKIqb9BAO/DLO4vCet8hR9tbqfUsODTlW+foVFuF/3koUj6U5tm8
j4RiGn0dclSkpb/cZsaDnVDPjQuWI1edlGv+DGlpcXK6vkWIwMQwBjiv76mor/Vzt9v73w4WilDb
o5jjSJsD0WethfpoLpKDqhJcJxnBZ/09gEqw6j+w8azmmyYJ2hW19YpVfTYxH6x6NHc+Yc/iUl5t
kSvBQszjUdXXJzz2FleCbQxD1Z5WpvV8BzBk0KvplCY0xUatAHXJ2xLEHHHNq6OLI1eFKfHAjqX3
SfQiHM+cf/q2ecr/PGFFvms+o1K8rVmWbj2q0KYpEI2TAbAvLSv2kGDUSY3OV1zzxagLvfD92U7U
GkT7eelod8F4MbBSqMK1GyZURH9EavYPnqqQRTGewQ68g+EletxE9t5I/V9bJE1KajFxCjIxPYZ7
YEsh9sg5Vx+E0nmwLsYgkDwVTNza8xkxVCrLVXsyLbsXi8inaQP6kRziJxb/anknfVYsJ53YxOPs
ElTfzJT8QBk7poR/G3olJ/oy77q9oQXRXgg8ZuhnR1ssfHjVGdYZ/Jg5+1nP2sgr8CC1A7VTmyhJ
/dsc8PB/YSjaySrDVkfpcNVoxlUjxAP8TMMu8lLoYe4C+qTicqzQpkrcSEWsxS/jrYPGnKgmpeM2
+pqIqONecMOMT1HUnL7UNWWAXH3BODIaBdAqPNJZGo3mQPiSw/tqZ7GwdebGQ/kRw2iv5yIOJ5ba
fkju4vik11Pfxqc3ii5nRz9Rq6hXMXjKN/tlTmuLOb8Igo47dvzBq9/Q2oSfwNoAe5Tt7dFYtrqI
FcxjNitaCV75eWAF/lsXD3HzzODPmKVVEQDpABu42K+MpWZ12R4Uc52GAsZpolkCDl+EjcbNUVOE
dpXQLBtcdFFLc/vmkb4S1qazPRl9v1OMfS3Y/RvgYixIzvmd502gMNwn0Ku+JDyp9JRHEvSES9E1
UjiXFkEAevBSvgOWHcajzFv9EnH6o/pX6F8bvKT65RQh3sSlghOiURQyqvZsyQk1szNXV9FIGLbp
m7Ti47xtz+Hi5Eo9aS/vNN7wMwqFaJaDKPakNuaxDe+PEZyRTHkwzvTNKGFxH6hxZtKbho9jsv/1
wfzSoDmQgfAkWo1xwMFmlZ7DPsNv9Qb2WNY20w0sSlEvgiKwLoKQciPWmr3hbcEbyDVhpbYRqGDw
VoHXKb2xfIdIMO2H8qT2aNWAif7ENziae34wlkYtBHV4zP20iECsXw7pCy/VhRXufvZiyh0c5tXd
C3KqPMg1gygyWb0K4sMPTxx9m2XdIQpA5n7FxmWL2q8bkppg/8epFWt/+brsyv4ODy3IRppNiqkN
LZd3UkWEikh0WyXKtWkJD+W15QSY1harhqyY+b3lpraFPla+kKefX90IVJ7YSveaFnJ0qiedrJhw
5rGV095e+UF8FNsZv9AuEOeZw+lPvB9MiKb+eMetExi390/sAStRM8rKSW6dsf4ozIXwQwRcYcOz
xO5eCs56Gr47mc+cvExoTyWoeo6fmoN6aCLCksQUMUadQLb+CbgsC6JyFY/3kuFAv28bZH4lWQ1n
TfQLmOhFA/ZO69m5RSegXIbnKs0YM8kyJldp5HhsODsVFXwUCT93+m3yrvhKszRSp+WGIQTUhMHh
ja/54VU/bqugnNokuqOODaqvgyBNAJhIbbdIooE3SPs+1OE8+m026PV7B9jIWbNnyzISy99FBkOb
skUyHUd6kIzUVkPKATMmDknfNNES3eLPB4z3jXKvSs69t8SHSFMEd+yM167Yp8o4rGaWCFEtzq+y
yULuRCLSlEvce0ICfcox+WPTm/eTdMG/UQjLAfm6pekb5ftikliLQlq7gHTPAHvRBNYaJFGj9KH7
bT0R+bHszbY6Ows0fSTWZ3bVomxZQ/XiKoHXdBhmibI33cHOglCpeGQ4GuCDthBHBhxqCLGBT4vN
Tw7V/sQIo45oByMqbQOkCq37RS9pYdhjg2aNLtjVwoZxHP0KxHw0mFZDge3ROPlU3qGnGsxfBU8O
TIYR+N0hY1Y1kiiw7tkI8/dG3R+RwQRmfY2Fs4X8u12tF6DaDJ0nzFDpagKVEGQR+tP7vXlBto1P
wBss1Coi5pjkfCWy39HvoCD6C4rz4ahwQ+RVDVTEVo8XbPcUPnBsw+Fgw6V3xUjcdPZvDDMSNZ1G
1DQmrK8HIX7q8q5JV+R56u8/Kx607v7qyvbIM3evIxIFg+8SXXnzt8jWm1akV/cpRMnWwbd6fRrX
OHvR8/ydiu9DsE9ue76HRsA6CWv6sbAAlyEQ2HLSp5M53EUyn30HkW4gCaP1COiKhAl51Vsedb9K
6gNEw6vd47e1k3qJ/gX0OQqJ8WwWvHeC5lhtFFY6XtJZYKHPuoLzeDu/BofZeTyTW/Gj1UZxGgs+
nJQ/SVu9ooxmLHJ7iHIU3f+yWtt4ECjnh6vSGNfDNhdcFVV6KycYhKip8GAbt28N2x+IHYsXLb/o
yQ79ULIfhSglQ+PwIPG7wpHkhY4T/tfSywhvHy7G08lyP9FvOQaPyPQU1wvZe69Ak6GLvYuG8rSx
PnzKTSEyLOfsVZ+c5EjCFWcev91WSiiNtMsQRdbsmdWUt5QafhcQp5wW3xctLbk6I/SaoxHWmfSE
+L6FpW2y9Ng00OJ/apjbAr1zAU1CLX1XH0dh6Kmd4DQf2DwLP7HXQ/Xj0W5UUf2QtarL+Wh79pm3
4dqdEdmzMPLsaYTUBOaxZRdFpLfAAUlfTj5tnLtLtZp2D7fFESeAQn4cRokHbWTIMlh3D0oQ+Hkq
L4PdNi6yWUtLeTUIBuxSVE2kF2BSrOQ46YaD/Ch32gPSPGGoAC1m+1H/A/6VtnAybOHvbn00rSFV
abBuO3bPUzzXBk1tKYsQVXYLeFz5/QuapVe15/uNYlCgu82czyND2um614KstHg3oCNaW1R1MFpW
hNpNhPlMD+o34X6fIT/m4lp2PSEthlahln9ZGFzU/voT4yF1ljt8mx6/0BXaSMq/w1ovleUMLydq
LnMPbcDDUelRkaY2t+EBJDIxaZmpvvesEEeypYOVMiJS6IDhdiE3myRc3/XvGG+4g3lPFnlR38Er
aJpf82REOT4GCViotz+kOmIdKl0PZPdzIWdXdIRJp3OD2YTY1l4W5VOTyXmBVWs9hStBFdgsLS9v
LintxfuZBGs3AZ5ktCH6Nsz2eb2Z2/2Ipt7vatJPW4HObp+2eEWfO+uFDMpbLUYYWHLUu/SXWwwc
NoxWdvgPBPDdwsAr8F6O71vFF3zjq42nQwBNG/xR8VyocF8jU3wWcgmHtCVVdui6Ijv0OuBhDA3+
bKKpMjV5FwAfkmVjNNpxlydrpnfb8JcFfS4ixbg/OXp9rbNUs4zoGa8kK9anc9VFlb44z69XO88H
F/pDF0GUeig90/Ikb2C26jFsFEp/xoWho/yjNee13ssYwN8C3i9c0vR9ezGwnyx7/NArQii1OCxE
M/4HOLo/VjcvcPr6GCtgGHo/Hk3ImU59q7f2MlFIx243CvBRqwRg0+6kM/fE1lI/S1Jr4XSNcYS3
1xBZIfRPKEVO8dzhMOpcjfEStVJc7i3Z3PM6KdYXI87FdCgZq6k1QHj+G14Fhv9BfDvzHJtq2i0p
wUe5K88UcX8Cs31cNo64dRBwuY9H3JDuOtrSJjcsdehR4WkVSKDZRWKikYneaj307EL5PodILLLs
x0eNIlR7mO1NRUw14Kf4tJWjFAvVSVVWkmBUMphCHbq6lbHSA1VrYKChKuuxzzlFXYqRT/vyN61X
Qpgb4lpFk4Fmdy1FC/5A2vHZlT84H5E2IJ463HWX2VUH5iO2X4H2DVEDH6eQEOVUHN+hvJmKda2U
DYtz0J3queXDIrc+zXyovcODh0xs7wEeOD8T5LNAEvKu6d+zF2pVyi7A8PhI5GQa7mQsp83qQ5Bi
AcAxu986vLGBnNuxgCtovIZaC8Jl+IhW7KsKnJAU+51plKWTves1mS5D6iTZh7sgyi00cuS1w/oV
yDafS60GcWKCFUjaMtDTvgYHL3mWxMe6g9ej6N1ETy4U+32Ad27OJj9+SD2Pq4Wt65TJ2Xpv/HXP
6pfhj7oVSY3hMPLrceaIU7qbODJDI0zzPBjdt7TCn7fDy29sAl5iObFRL56evQYhqsBHXuIS7Mlq
PLnSCzIehppm/zhSEGItTU85EszfwruoyTElGXSLY2rUHSnS3ghJQEZ14St4yB2UjVJ8vkz1QPjR
LLjAVsb9M8alTAXuO/rOy39rDzceAiDyPyaFP6hZZJFK/ILIgJysyhbFed8o3rl5vCKvTZGTWzmN
C7EXaCTY15aXn9xOazIicHDmAUNBwkosFeHkDIPk3LBhkbQy4LU+mU/jJuE7Yusz0JId4VfMoEyj
ISwgEP1TOKAUC99eQxVYJqhaaruv1688Mw1kdLEy2cdZvaYNJQ/dkK5Tx5Kf3icN8YuukZ6I5PHq
My3UsAr62GqES5glrJi2+GSwtYyqUTnPf3EUaiZaXJ7dw/gA94glyBBDYOHgdAsUO3ejZq3/Jzb2
nBX/ehqfeQhFS+3v6VYU0f+yBmatXS6Pf8Czkccl7zoZ08vJIFYL/sB++sKBRXkTE4q3PFC8pLHa
cnLUn7XYSeHAkleb29L07ivVrjHmY4a0ESFEwHNIW5no/2ynFZAGCr+hNttTk2nZJr6QY4BdCTug
3FTAX7br4z3jwN2b8vliw/fwEtDtPW5vUiMdCWs0TCB1sYB6EOpRD7Wn+H96CpmsJ211+My/pmDz
cKIE/QMcXgmKfNYNyU1e2WHZKNG+h252sKm8T4ulhpzzAyYNDdXcw9ieky9CtGJW6nzJltepjyC6
wocmm/5NtKo4G2hdtyfTytw1tFFOkGtPb9rxTfmitF6ma9bF7ktKnZI+lp5u8u+LmR4SpiyfO2hm
hDGbKZVps3Tma4zlZaZco01W4XCNbDoaQdH2T+fEZseGUr7LrQPEacMOwx78MpXJRxWZpRa6dumS
3U9Hqw/RZEK01qs0eWqvi+TRdSRpvr1R51IAwCHs9YGe8fEMP0PdLytOAXuETMKrZtXwVe5KF6S3
JKLL8Ssg1O2sgS87OhYGh9qW6kY+Z8XI1VpwqPq4bp9smq6oxJTOviYo7WlQlUlTKYZDK/GY2W72
9Ff2aBZ7R6WK44hjWdSiZn4cSJbQ9FBxx2h7CiMJL/4IzW6SWmF5zk0CBC2JjWw22EBSdxv9QDan
MYoaDv3psJKiXRvPbupkMTYJ72yBDsOIftboUxieqiU5bNLF94w5rju7CTUd4khqjgvnOKweypwc
M/DOK9CDyixn0uvBAwUsyy3G0De+x6uL7h1Y0/4FX54JfTD3muBTW4it1MB9zB52V9g3kpsOtALD
kQ3F+b+kueczePg+UIl/UndfMV0mbqQ2Mi9XfkfEtwYM/7Lafa5/Re/j61MKX/yapQmlTeeVPub0
EKrcVoBYa/d4VIRNqGpwzVXM77Kzl1fOiUJGvPRU6pzPXK6TCvv+eLGlNBO+e8Jm5l19R1Cfbm1L
FryMAcuy4NTOvPJRkB/eV4MZb8fvwphJbvjTxwY0OQcc+PL7QvChnxoz49UlpSg2Am1VN/IPXhOp
nEv9yBelZoMQs/xMD+df0gUm4W6U6N4T07UQ3c7e1eD+iyGjbn8VUTdbLZ5ndMHSie5JVEE/h4hV
zReF6cv2/ldZQ/pU3TwTuQQIp1dvNyQma3Vgz6gGH7PDaEUhrICgF6Qpzp85ickyD17ksKWfNqU+
Oe6I2MoAuxOX41N6QrNjfqQE0MNLiLOnLBzLFKC2w+MrLLXag2HhV6UrL4zLtzxcUj5744He3Swq
tjCWmT094vrzTXk+JTHSaBFpn3ceknyww+2y+pBamnfb0k/9rnwGPxprFeLnvOgV21RBTj6wZaMC
IwiwkoG9u96rBEwsG7wQAY/N+a9FfQzCkC2e89umILwHgGT738G700+2zPhFEvPKKTb+cm8WjHlq
mJ2UAb6M+nWIwB+h70k8tnkZ3uBqbPz2KISZ9hkoFabxnSbBn1Lr2xus8/+qHOe/ULuvzbqSFyeY
gU3r+/Ykl9tFwQZekH/ccBIacQbSUv2/EJFbCmzXukB6qX/MVTSOkbiRjPpsCn/PT+zNldzdPtTv
Savb7LUocUUBA+yNtUB951bv++GqXRUeaNVSOJ9CE9QxmgOHbv8h87DfMCt6vyN39KeIDM10r33T
F8A8hIqa+99qkoW7HG0wB04ClokxslUVO+6ALpAU44bgXMNPD2klmO8c0FHG70IYf1vfkM6PqRyf
FKhDoNq4S1sqAtX+QEhZDiDmWewffVNo5J+6NWz28ljyuWc29cHPrmdSusa8NP6DvNIABx7RqiDN
VN6N9A3Srfceyr0VL8YBuTm1KMAQ61qaHtncb0xKjra1QBqPqTPK5JZT1MVpKnEoSK12geQB5UE0
5ZIrbDvLuF2tDjYMMYU5z+rLFJHf6HUMLyjwZSDrwRl9bbgDbPqra3LxF0vG/d1XODXmZWFEY8oS
GA7deSjxWIMgaeaBX87RfM5esQyHZDAIpYsO/sSCSfmPsuEiPF7qqXPTahlxuqZBPALso53DN0fJ
LRTyUmi6gLlmUuYQzpcVGvVSsmVuSbDRGny3YOBneAe4AGsvwl83xt5XzGNSoFsJXe31MX+EBBFO
itvOiD7ByN+IlJ/6RQvK35UUsyu1BuuvJMMvxtWzTXoHcAGzC76ZYgUzZUwvl5gLLUaLQyB6C+VK
bmGch2kilJ1KUFzOBG5jD0LuZZtum3n4FGnzLW/wV6+EGJmjOxVmQbwP+tFK0pfPI6pke/JK4hk8
5ukfMtYeqUcTc8M5Opcp4sVCqa5QHNCRURFlbEEBCzNBVhiAcr+dOI/V05M3UFYzxbrzIC/5Ws5y
Gd7pjC8VpaKpuLo5+Jc3b1tzc9iy1a3CQ6NrvsWNSH1xZaMMBD7YsKJw5108gzSgK2VDPNTqiDFT
Kehhtaa4xt6jz3davtgpdWm9Lo8y1vAziC9QnzsR8p9UPyrz15BWROJbSf6RHodvx3p4jjypY1WV
RR4of1wxzmZ7/QH6qmQ3uID2lfyaG0nWImIk6umpAKbyACg5DEPqMdzytjYmLoyooIpvjetgFkYO
KdMeqi14MADgfdToCIfGf2i3JQmAFlTP4Scaxm90TV5lWHPRGjItwowwlo8WT2sary9ULLV9uQOL
7GuCijLn5voOtVFtksgwhe1V4mZvO7AFj1HfN26X/j8a8vAfnUrWLbnq0d++kOIlUHbtzjW6qX5f
bzKb7Ri3d0ZNDPKz4ke+yAJ/LsQNu/causEOaYUfzrBKCsa3EOrk7wxqsQxMUkgEGjQiqHaorw3+
bgMzFwp6jSif3U0KxdSwGRabfKiIO0m+gkgUIqg0RUwjSV/yQQOLVJs8wws6loRpUPggoUGk/wHZ
C+QYoI0jPYq0H0WOwHkGsfSYlpmZrmC9XNu3lwSID/9C2NYKBRVb8bM6GTVeb74ms4sX1KYkGLbV
TAuVVm5oNMihvc8JA+MlTdWqvdYwOjaSisyfZQJTMKdMiIuyAQxnmhxkIWvtzyqlhPRPqclLzWnM
hJoX7vDFIx+fN9FmuSEek2EhXhHc/4xURiOcMkyKUNgNN/lBEA2y9XIjs99IEWxlypU5b0MmTj9t
3tHpTLAa1hMsqPJPRGppWMvxmtSgNIlQCa+H491ezgHW9/DiVF9Bt4QiGcMHMRQ2ozMwxYTjfqx4
dLVjUyKR1+vJnVCR4nv3QpkOvokNIt87KgxEZe2DI/pyfLMZd7Ir6J+a57yaI1P7zQ4rwdbTTFyN
Kau3+TkdNw0cYZsrzCHsyB0dUxs5p37uybYdjcFo+4SlDgiiy97kl7HLdnl3vO/0vmSas1vMBxVh
h6/sqeeeaYnawtwH8ogdC4QyGyArc3CuuP250A+e0sY8VJWQ9clirZYEoJQnZoIzvrGLfbPjW32v
7RAp8npZN7ntLVXH4JzMF4nleh9SysCJtgoe/5Lr355ZLHJ/L+fZGQ/cgKp925uGnJDpgaVRoIcf
r6ZGS4860hchfWjbIWEuFCxQCXFGi9VuJfQ460n4aKH7x4FcVVupCER081P2QsR9+kCdGuGoduj2
bKSauugOWgTwV17sLDPTVwDn0c0PFp7rIIToFPpRHevhx3UY72juTQO0E8xMvWabZJ6p6FaEsxg1
J3+JN+SYrBp0vlLZiRuG3Ro989C67jWH3fldn6WPtMw4sDCqZlLK21jfpiHwxtUYpnQDoKrqZ7aB
GK24sSObIFjhwZ9qGSA98mRl20XLCTQcHk1lf4rREuNziga4Dyt70wumzAqCePU/Te1iFvH2rOwh
Xg4DuS7PSl/DFXATio4eZlc74HvCd8WqG401WSBQaPWn8lq22hvkP1FXZ0h4cw/BwKUf8FnTlQ2i
pr8dC+KUNmbrMO1VAZjockKwbNeUQ4bzRuIxPXAul0S176Lu8EGvDGwpkqJqfrmW5Ur51Op4qKrs
J3Gi3emopJHNpO13KQ0LavVqA+I+xZrL6TpGv5EKUyD1b6MBKAl8wcwqrougGonqN0/kLMwM27lX
HNYPsUN9HvtKW6lEl4gni8zw50q+lMfcc+lIuf7iVSkceGCTM7XkE2LcJiM8HrOum72sfV6n5NeV
oty/K0NxjFYm32AAWiVGnzS/wsPQb/d+pR+b1wN91XgTP9A2nTU1qiGCDHJ63ykTCpXRnlKmigLw
bD0HfDg+4CCS3JLejcmjZSrlWCVpNokK+kCmH1v67Ifbm4vdDLqXJ5JJvG7/qCRUIyAqAtB3CO3X
hOHNBQlg0cZPigcR/Bfs7PbZ/hlhuIC2JnMclH9QsMTU6VcYxWH4TDBVoKYl3EnpZfbiw2+KUZqy
hAQthiuD1wsqkOnLI7xTpcJnJiwn/0N+UuGiGJwuVbH45g/ibswXWus1sxmwfIj9f/4VxvX5OS/x
C5bhmfWY7fwL2E0mb0Ln1xVBG7mOBrEdgr0h3GvW7pfzFLvvXxR2FtMw0BlS7uyvxhe7Ow9sOfp2
k2mEbfULwfk23fTc+3M2AtoV5N5gYrYwE0OrF+opeZEg+OhrNlbrO4ZckE5PglJR7vzGr9cK8gjj
/iyoiU8nT1jMcGoa6T8Fc1/gbiVdhvS7hDkVKweblRIo3YuBYmvXsO2BmYHJTKJFjDPnrKwOwrHo
dxQ4IM+Bzrdp/XTz9l0Nke1xO3L3GKZZS4x7ZAkDRoXuSX812/2cJbVGodoC1yIcuaYgS6+71EI/
ErSoCuz9g5O3Kbd8BGGR0e0PeFl3XrNzonx8Jdmuzv0M6FS+2C3ySmH95sE7hvq+iOUkowPtjBsz
c6utx0WvJt4EUqWxngPJNqYQGORKetpybCOLnZXKhkUGZtqyVdFUKlIRfKHVrZEckcsS27Qi9lwI
ivxXHtr8dKbJY6FN6ghJHWHEZf9IwYcBblIuBTGeplI7Nr7z23xwoZAea2v1o7WI39s4EQH8+zuL
cvwsywt/yGtAmOwKLpOoIaK1P6Cl73mWuyFgmdCja8HH5OJoyAhKlB0o3qASNqKvfJmaGlGbHU3P
T4lcYqNjoWkB+iz3XCHGWS3AymvNsyKYFaALoZ+Ra4b5gGFqHN5SGCnouCYr3qEJk4N8i3Mhlqbh
QhLUOCooyN7aU5QMjO95WHmpOBnIKLQ/PIKGIIRipuNf6cqTPutAfXLyu3U/2qiGQkcMFgR1G35d
nMA5/7MsIfaACO49UitAUOPIJqU/60cHD/etdWK87T3nRVvw2hnSPQ8dm3/U2HcKi3nvzJkmmj4M
rAef3iZ1+lwt6O9JpHsfWG8VBSvXNNgNiVve5a6SQ9TZTYiL3y4zYVNQbZpf0CT3CWJMY3vTlpnJ
7bRUOq6T0HGDZWKnrxr8Wg+k4bSgKxGhRvrwNLSvyKzrlshPDlD1W6T/Sjj9ATnYL/ASNoK5C8om
0C/S+/+0epBH5B8OxWfRzqpNis5Uhp/kUMLoxpJqnPvXIsEECh3QpCM+Jo0UlgX5UTyrtnQmS1v3
IWnqUpQLo60TnF2J6g8kocqgGSILKG9IvdGjrERw4Ux2ISra+qKuSgZPiJiYG4GVynCMA/yCqIKj
kSiw7C7w496NeVwqRXuHFiDLISDOlz4re5+iu1vTvtnKEcg/coxvf9XbYtIG0I95xKXC2izwLaZM
AD9IZUcAYZObUi0g3mAHX5L7lgkjnCDXEtvjmKXAIx8ktOsSrCfSXNvUyKJ9jf4QNi9Js+JV7u5L
PvQF4kpXtpi5OyQg5RdZAuX1rfBeemXeqF4aUT4/gSCEWSwtB7X182jqs0sUbMjeDg0SZ+DJF4+j
01IEnkwXWlO4yBklECComslZmwGF0Rwgq78uJ3GtzDG6ELrW9YAYVpey2n+sJoo5sNBfeAIpdqW/
6dfyZK060J3/Eq+5JyDNEvjqW+HvbOaXhkIwvKf91zg2hm+3cix4UtuPvzRBuCDQ2q/hjAP9VdHQ
v1OuEKfbvUQkiByOeF57InWCG+CKVVHkSvdVBbiFgA4Q7npm1mQNamzDVcdfKzbtAqezV2jyr1Y1
wHvcdvYKTOmv44ZIzab3jUcxMMzWISSSNciSlO9aqFzTXP5MYShUciW6YljslQPmh5WsTlo70V0i
Z21sKWuvTRJmNdxRjJaXjX9AVuVVjHvYY1Iv6iS3QsUakBWUA3hiHnqDdLG+eJv5453Gg9tQlDvz
cKLkDhPfG3MHOQ7Q1oDqqQSo2pPi/Eb/+vS+p6XLyTLFjuvGyKXIy14IHGhNv2fVgS6h9Y4dVLVq
huR681MqA7em/tPM51OJnRfL0g0MAUOegprbYinrLYcOvkmCBRjzEIDZN7ATTeb6+Ce79aYRkmG9
RRudyR41b30Zn2YzNwKA4lLEE+LDrodF83mkvYgUD8/+tKuRAdrsT2EgBa0c7fcbm7ZWBTBx0Ddw
TagABmEEslm/ScznZOH3Pa5zLJdyycguTq2ZOwNx8n/ylOTlmVeRlkNwUrwItVobVF1watAHuly0
NUj0lyssGY3gAxftzIxACEPHrzWyZMCf7kT83MrATNGtBoDyy6KYOPZyryiceCeT8XoC6KOQMLQw
opGjEZKagYbQELqQlesm0C7DHwHVAbXMxKgsyOqbArkLi0SthI/lfL0ZbwV47MNO0yhmGaGJwEy6
qsBkkySnDDJ2e0pIaFei41jCnZs7oOMC/2nHThQjHNCuL9VXFjs0wjErwUOINE26hGUGWBGujB8n
bMRs1lxa5lfQZ7RRTuJNWXNOsOAHH8qTQGbjPmLjQyCR1DbUjN/1rbfb+6AQN1EPm40ZMuCYzXT4
FZhf68sbvvSNSLfyuYc4wMT2omKQohQxyvvz2u2cmD2kvXkJ8YzLY4sONMJJeoEofFQT2q75qCnE
a9lXP0c55yA/Xgso74ecnwGK7Vs4vvX3J8BsahHhZpSXzrKKnPsy+mV10NkM0Mex8/XgA8iVCJWx
FaMmRWpLflAc7Nxepwz0lHH4RQHFJPBQ1PyxyWimRwODmWL35nOkAma3oRA2dNKDSYo8wp94W80B
nsoaC6T4S5ioGXZjwOvG14apthG0UjMs5U+qzw1pNPIFBHw7vThEgNKlEQViqOxasdX9nXYRr014
hUBhKH7GWzUfQb1g/LdzxP0E94KG66ao+w4jh5fSif/d2TugIaBi0dVuD4Nr05TNIMrLlQq4+Nun
EEcsP9twGm3E9MXiVXhk13DDqg18O2euSqzguGru2HXmb4UE0VoNjh0nrXO7acO2OZJ8I4pR/NXt
RcQNWSCH5mRASXbU8n8oK5Kykwengr8HtrHdMUnkXetzJMFIkDT0S5ses1JTJibL2yxGNWwW6/yN
5ic8an5HGDzKSHTHtfPBBxCMhQAopZB7hFgB7novO7Ogjzp/BmtthIoFF5KsabZqI5oA0x9tFvSf
qEkqNphWAzxpCDoPfezaMV7tSfJllIy/aRxsSfD+cJGRI4NkcIMqxEv0HtDlIrvgzPNi5HKM/GWE
ix71ZnYCmjEDA7UpBpcJ84U52WJnPRHnsQIrYUKyDSGC/2PlONiiwLM4ZSkc6CrO0YTtYeu43QCA
HfCmPbdP1E/LPMe788iHIv2Oyx9X0djJtADs/aXBNkc3M8Ii1WKEoG+FtdGIJcoj/pVZNIaY9Ths
RoT4psFxltvdH3DmNXBrpMb3IJRq3npnIW47xmAgwXPKxVNcCUYhc2WDMZDO2Dx/hYAWMK2c3b4b
pVPsCytQn8Gl4TdKmjGk7VyXZ2A/unhERZeealBW6x8mag+2O3YcO07UIwG+iIHb0c4s2gU8RGyC
gpws2e5YofnFVGDK5T6kz/Y/E44viEIrtU72tW+yRYhlbrCBuwLd1Jy/vteE1IB0V9zST4xBOYKy
rKiLHyK0H3OQxTye/jLAcXQB17NVVQUKua3/hzEqrp55tiGHtJMBebyIRq7IupVAbAyX1FuT/rqV
PClmdu2joySMLb6yLACNBvURLNQ6qG5ol9noobIvpL3Tlg4ClGq5KAo8/uXe1jiBs1NO/NJlUq2u
ITxS3wMK8vWE9x20rNInWge8lZdwNuSYEVR/fG3LO27yT2nlqef+hMhy0CgSfikWiNk1b/IEpI2+
5hR+pHkUDWfnVLP0bYG88eewx+z8QW/Rot/pFbL4uQVwopMNSZ0moF56DJGvL0UGfE3D0URmUTuX
DeNDLCv5VsxaoI7La5QfBsb1dOW5hnyOUgvKu8hV0K2C8RsptZOvAOB8haHMTmAM8Enkd25RuFB+
CVC1WZe3BPWR43QD4iTKYc5tLZMATWXnwGEOyBsaYOrth7fZ/VExL2p/AYtMLcbOgrH+fXsNZ+iE
09PZQVIoKDiG6YvZqRUtYAEcYdIBrNaNukuIVgrGNaN/6512/6qwW8FF616p4RpHcegQZJ0XOj+T
WHIs93cViZwau4GL81SAz95ZXSW1dSkPVhsh0xjb95gYgjffxO+vcauDEGNglVFO3k5qKeqAWBEx
KWv5F+qOZ55TEpGHcgsRZqQlAEv0FlUUDAN3Fxvrx7s1/CGsYs43Tb+ahWambBwYO3KGDHyJnw9E
oKV8nDWpxCVu7IVj+WszB0lihNLwahIF0KNQ1NMWUSJCl5DpnFj7iwsOqz2baE5vkwHjB48u9gIr
RLNAGvwsY7oWnEPxY1z+R106+lRTmUUaEDvN4/zM5G9g8g0kRG1g+Gwgtj9sHktRSX9ywsYVoEXp
kQ6E2BMK8+uJzlaEnf/6fGe2/aLV4XRHKvzgAEGXIKTaCIyvSQ0i7WetUFcMZah2yHBL4ther5mk
qQFHuyX7ok0cY8CMH3pRDGZZj7yGGAAr5Z1vvOBWiYEQ8KlxEB1tIhMXlOz/NtvHGwbYTrVkgMmD
uazDlUxPVpvRc9NNputuoRmnNFow5MNZTCgEJDdjZDWy3Kw9vD7pl8ToxKHYlJF6/u1Y1JON7D2n
s99IbfKExMzZ5+Jrg4IUSpmFUdg6ZV4pG/wiDR2bHVDmLB22O91nnJiYYsbJmGBoipxK1qlDHzME
jh4fLz90hypMvmev6iDvYpuFMRN3/qW9ItnRmIK7/IPfrbWUxm59UCDWzk1PeeNcV+cQbVnF7qo6
7FjCi3S/bNWKFdzCMkWHzF2SKvjJTxCclvCoT8V6V9U+1aDrOomD2U34YndqazbVDfPoIEEnU8+w
p97kDvo6trbB3a6nL7Tf75hcoBnY9VI6o1mB2ynbBrdO9pOVF57pMJHq7Ud9vOCBCP0mwmlRgBV0
DxOG5mlH3uYWm+hN9LhNZIO65Gf0ixnjNRF+CyIjnOKDd7b0u2YHWTUGR08l9SiBUYKDcOn7EcYp
aMTxfGVVEJzWi6ssyop4TvAv7T0+qqi6tndCPAB3dB5r2CL9R+YciJl9WFo71K8Zo1YIj39ttOkB
gx6XLLxg1KI0EEQZYg/sEp1qI3YTNuaeVZOG/9z55uBHpuag58+S66XR5fC/X/Vch5SE/E4HxBIE
esCUBq3aDtpNN8zb5f7d/IYIG+p74aKYdimZSa9jY42nG1tJyyLsLyNjkenfy0etdYs0PRr693YL
Rs1V2fHBGZ/S+/lt0+nODC2Nt8s4yprUU/lT+3XG1MbxF8zZ2g//THs4sedpWn+iJ3/66QbXLgbw
i4he3OEUb8Wqt2NSxEVkirAPzFaTUUsjg6ag3EY1a8CwdEum4aK7j0Kp270CPvi7KmsBOu6nuAHX
AuxYBEPrLjf/27S862RsgkCyILyl5xkE/rGwj4RZHWPn/ncqr8jxMSGBA1pDnKT7eoIWKSq83eTL
vF1ljsyLFLHzhE4zMX7SsdMz+BrLh/49gcIMMC2XCqjF54ZGZgecTBfe/PdYZpgHziDVim/vruh8
nqepG9dsMF8QxYpkNuZdc+xafzhh9wlzszi+IWKK0Xzo3j1gcRwQN0823mb2rZhFB3WuoNbs6iqf
SnuWUAdiHJOuElZmn6cwIYDOj165K7SUI7Ta0K/tLBQ/qlaqN4cnpNSH78a36J/LRfONE6ZPai3z
H/PWIYuYOvPWUdGZLb2dqOA/D3puMCH05ZjmPuJx+v2P/XAmkTwNUuouA6xVNl70ZvGfhvzSHcU+
gDl3v5D7hNjYNGXp3J7RtBexC8mXGVZQTXug2NrkLzhWapcciwHeCErR/rCl71oO62uC1RpZnhPT
BU7tm/GvKnKUqHl1ajcYJI5kxKIwd2s9Jo1QjvuC+tauu473S5m20DBtnCUY83i2spzm0IFSLpO4
Gy9QO+9nuK5NT+i3IyQXntyfeQ+k4z5+sK6DAiTRxv9VBGEbp1gw36JQNYX7J4eejVQwMYrQxgSY
SczwK1Gxa/3+jblRNUlatmJt/GZvzddAhvNR2MOLzymo3CkGvWK5R4oWDD25czhe5e3/fSsT14QB
vWol7zFZP19+U04ghdaOd/dTbsv1uA40RoVt8Vj9mtx0omZERf0s3wZ3+DNu9GYoHhQdrkjQ4dyI
cgWdMNehfWd3VhSc1fr+VmA8mvHqpsJht80gDVwbvNhJ/gOrtppvCMV7+iYbeGkto421QZQkkIpA
XP+PnCUTc+zxVP5Oe8MWSFEmUi6qyj45EMZwG3/xxREVBhZu1nycZ6B+fZE0AG89YjxvWnot00Rn
UujoI0adY1dclw7L8QHKC3IbBpY8C/jDJPsUojn6z3ioyXLo07MWLIb0+rLN//QxnVw6EpbWnIJA
OXUPn05VTMcdjKixoZ0no/wuOMmu0rDcVS2ysUcErM5Lzzajl/naDFUFBj7k2Q9cHhq7BOXe/vK9
udV9Yq7cHQNm46A1dzNHPerntBne+eeAPuid0ZWDRUwlapvTx6k62jQdL4GTsY+mCFdaR6vzPhAg
lj1huzq11trnt0VDapO8Nq5TUTqGZ/XQ+jbUiSbfHWrmPGFm4T8Kh2+ErySwB8N36CGpCauZ9pgl
VOCtCBRLKzuzMJkRPYrFf4ykkwKPC8m3F3pFRx7XakEAW8J84bu5Z8qC63vmAXcFul6+6g6280ko
1BzY5q6Ab5pG3AAbkh3EMwOyjyQnJzOutf1vZGgCAdfLFcDtEIJl2uVbK9rrTUoVeV0sF0v1EwDI
Hs/CxekG2TCj3+n3TpgPk0VuIZhN6NOvHUqEyXsv5FMBMoJSj1F7p12CNNBy2Fg6BGU30WMZf+ms
4mGsShXw5KupfCl9e4B0++mfPrP4Ljuab7pY1lW2rm1qOrk4UoMdx5bx1gBJR5B0D8FwSJq8XyjI
HrWXjWzcU+WghcfYOAEkEWJ0Ax2R1RKUUFj2Er52xGS4aBreZMacwr19cQ1JrcAyFVH5sd5SsCDL
7aI5MFZrdSCtE3lq2g/2sUwtyLk4QoOXQc9yYcw0Kqk8hkaRimtVfVoMzkk5D2IweEB4kcRNp7B/
LYTWMTOBCp6DKpSfZV5efBp1YJuxjtRr6EdJOozpjCb5Ypqhb/7G+sSEJ46W+W8hIXeBxTcwKwsE
6sGceVS5nZrlsH1aZLwsfDsgf8lcvJRlH+sxMgr9MzU+oBtWKyuvgplFIYSIHpO5y7KiFLsYqnkp
mfN5mHCpz24gEavj7jb1/k8CRtIJJ2jJFSjYQiC8iz8eRW6s6+lHbPKdLclr0tfZ8525IrYk816K
z/nGjFrKN7YoCyKGErGw3F/DYn88mvJCT07e051wHqmQw5UFwRgTQ3CT2WpBXOinX8LANLvVE3ry
0324cQxGbRJVGwSFeMjlmUc9yzAiUaTVMYd9mk9VPid5gInOlE5pHq3cFio7hfLIg1wf0ZdUkqM2
tMcLKTkv0y65j+a/U27XssFhlMdC1Y8Q+FJp5gkQWRZCuL0Wj0k97DLiMxOaf23RKs2hzItv4qNB
8Lg8oqkSoiOQ+7fpJ7o/g6yH+CuqvmNF5hqvAc2Oo7VdQy/MB1sdtvqA8LgtFeCKJHKTTZV6yMNo
Up2Tky/JpB0Er5xU0HZ5R3dhIwg1Ngn6xbzjHQkuDvm1lR3Ia8m8TM/z9JhiEHfOL0s/GveiN8AQ
Kyc8HD48PZoOFFEpzzkrtebXLXpMQv+e4irhxqrYFX0SHj3Ac/1wXE634Clg8PEmX0y1MZNfYKG5
GWw3cw3YxfMYWC4SxiaQcUghbvegciBk/J161KtGEj7te8+vO30Q6zwA5onOM5F3JA3D2u0K/I/g
1gsgkRX6jdI+A5++3IpE8cKLsBgP1aDuxfy8xm2KuRDbzmj8MmyZoPq5At8EHJhxelTcgVanqoO+
RSnlRCOkh+nGA4YPRdACnEFGIWKHlOUysdM3TiAwhQTxk0r64yo4wfs1D5AfIXnO7/9MBagb8AN+
sictdkgKqZ5BwC+VBPLZBCdqBYnmngbQ2Foqc7hISAIlhdWgP3I+A/MVhEEjNURWTZWR2uBkkJD3
DZxBpSWi9U4VU77fpl1QVUgC0CoTON87iI7TEU6hR6n218Vg9SSl5LSyQlq+KU4+rxE7JCtkEd7e
agkvwgsK8TNL//311TSP7GsB2GwxlZ4V+xXp8ERswkut5xWUKrHttJl964omwPpY59NWwDoaJhzQ
mzW5Fry5SHeJpPMOBgGCjSgarGk2wBb5nNrYQ2QKsSk+KNaEYnSef/Opk/YIQb3uyhBonER3T8FS
N0+TkX9B1SglLFn+NozW5RZljtqc6zsqgsq2m8YTncuTBomFd8pMEzd9ajeOXpphGoJNtsBPQJIg
mVQohamnbVx/nrQ2tE6Ejz9Q0X4T2UJVjDOvW+63jPEIMX2HO/n3Z/RhF5wAJuWHU9FvyGNO5dnL
Z3J5BUQlezn+OSQuczrjS/dAoXCZLhxQzJiusVfxfEMWO/pIyEzS2ktghRWzxnAJfyiLEPd4SOwR
xfpGwj37/9/3q8zuDb6XfNl6fNkBo82iFk5vkt9HQgk5tLrSlyf1d53W5jhmL2T5dEH4Zo6QEbcf
20ilyThRGzxkPqSNXlllm1tvIrIfqERkz6J8oFycWYCh25FSqUk7HAhpFQfmKOFuhrXd+wEACoBA
/cfUVkcrdpKvIoo9LBn5aHRs6bS2fJxuoLyLC0YVMU+fyQsD55C15ZTPfeDTblrmB5Q31SMgrJYf
MntWm/QS8zVfKrynr/mlzVxgjUglaZ2hXJboFWTbKu/YLpcbG4xV7tkZQWoKl7aEDXQDXa+P1bGJ
NArZpbeJAScLwS1zxbrMQCr9gaK/9TyqLLrCJLV6+hJJSmqugYuvtjWvs9HQsFMgd6LdZoPe+v8J
M94i1zpRMBAibiT9pJnxXeiCNqygdEml5T1rjxdlmQpolIVy6w0b6FMVi4cEq+d5w4HPBHl2QhlR
oWYWNPbSmzqrZdNc85yB212qRtj+sQxmvn7xyQEd/nC+wzDuVB94567zsAZNmrNs+0JYqTc1g/bc
RAbMqE+v7KPhGId05At6jSz+O8eKTCgFjIAx3RMb+4IDyTnGY84Lw4DdUrQvHFXP1wMPG/A9SMl+
8PUc9GwoY+Oss/VVBlvA5uEV3iKL+Jhvj9Y6GjXHDuwmP43zloUDlngyeYXaN37ERuxC7bupHC7x
7SFWjtXTVEXtn21oTCRadiubOIMoZl1kjEjcAPB+goPKo35JwcSN46tHvToCZ5f+KPiupqDQuMDD
ceqzj14DpsUao3MK26Ts3knhcdoQW7U7aPodIPHpPhNWVUmHf1PAFHuZ9W/J8NCXaSUFHAoHp6o3
NaBZqLKyS7v2t2HbGimNzyvV5A5SJG/r0fnyGZl4B2XE+W/xdEyNI4xQ3ZR3eI5CcMLICglZQchB
r1s8HTl1wcPEV82XSHMh3JwrdHglZ+sLZZLZUaWVMvAW/H57cz7iKC+AMbd3kfm6GOIQqNZHBdeK
JE3VfMRF5OK1QJrU8NC+jyClA0kcfIMxN5n1Ygjx6z3SVaq1IKHkiSWUfn4Ud8NgjdPIDtFlOFhu
HZSA5Z/k0oOUEbNyUNzq0a4syWSrtTliOQyU39LNF/yaozYQum5Xtx4SPr7vFvRELxpY/NzyBuQa
FuNwO/PCLsKsc4tn+xDfbHnKCMf+ZwCtxbeFnCGphGZVci2XccLZhj6NZmgyqWBQLnDP4/+XXkZl
VzqUDLLSY3KwKAcb/6eD9LyZmx1tqVBTfGyaQATQWdFfYDKWENLaWuZ4p16mHEWDKkE0xg/kEbKe
k+z3SYwHJOcBtiU5//E+q+ZbytW1t75pfyamtOeB70uGeEE2Uk7lIGHBLcaNTG+DYSLbprJ0LjhV
utV3W7Ptx0WmOuckMrhlPjG94EcKl7eHAS6C6aQVllV5OdeQsnFbviyOoWxgqL2ennstbTUwkAKw
B8PuvV2QmczAr4sOpZPD9BJnkXpl7CKpd0IcBHwy5LFSmuSyUUC5PZxd1wE+DctcMNF62MXBdFSK
GawoddoHpRR249taEFHZPs3evPxhwJqc4+d0zpO6wGGeTZyRtFrCyvhCl58aoWL4WGnufNPle0Do
cWdyH6OOEbZtteDy7pMoilqGFp81XrV19htp9OW0QuMkfXjq93GKZYhd7OMckRvpDto5MiUKFH7H
9G5Qx/lY19Yclf25OCEFUhngBEDA8G32oilyN+NgZ0dNycbodQB5TnEXN9YohTMEuX0T6B6W5zBR
j/TG9r+1eO/rQe53P3m3IK9CoaMIFrBZJVxwSjPH8dpqMch5xuFSQZMFrSZNd6MuDxEEoztbuQ4c
M0S4raRbR0S9aTeQrFDfRmbaPVu0mnP8AdyR7ggwqUnvHz4og7EE8xfwLoMQPjYOYBM/v+w7ppR+
85NMZxac4B3lJ9pP1hDdIHyvTbKpmTyiUXbnii7NSnJC/B1evSrs6NC+oxZ/NXcMY8f5L804rKG2
sKw7hwi47n2AAApz0SLqQPh2qkiD00eNWKkcSgGcrCAa6PYSBG0a0eUAw5dL+jteL3K3K7cBK6xH
Tou2nGIbPAajCJKX8RT+Ylx/mML6ra00RbXZ38XGvKDqUppCHdip+CpZvHhquVmCj5WRZSh7LKkY
pfXqfPt3LIeKI1kl1Q5vE4VfUfB3UCYt0cvfUs3SHSEalJAg3GLWaw/FJrOYQGjib1zpvuRGlfRE
8XEUrnoRr0zvY7U9obT6tYGlePHEDaZj4GEipuSMPpEx64vJi6CIi1CYhnQ3ekJ4+Mc6TqIKmalz
VlNTKYoW+m4FIL7u94Bj7ejD+xniNSyvbdw8BGBzKzIPEKWTyCJ+vs7y9FM4JOR5R0FH3A17favK
higsFc1sg9rsRfWvjJ0KuQm4M3KLsamkL9RGhmNMOdybOF99BK38lKiNk8n1ZmoQTbS2YNEY2Img
gGgxLYVyk0wFurGsSGdyVOozpdzHVLWjYECxpYZNsP2Fcg/TqbNXRl+myrN9APeneIsLsfEgbFQk
yIlnGQggJioORQcOnXXNNKfPo/ggC7Y+MmjoA0LTLXV1FM6/iBKd57TZocvl6UM166AOu6hXZ7xt
LI8MLJdjkbdQPIHl96XpJqSsbKrM7pWq7bEyQymyDEp3b+Q43b/YYwp19yz0qFAOkBQ9/JJ2YaX9
JHtqaGpTwcSkpG40p4f9mHdkgGb4k6qBHA7lOWLP0WU3YQ753NY81HjyzK2QuVLoA79jBNTysJIV
9dJ07l9JRmjgWlIe7zl7d3f+zRce1BOOTjweyivz2wtjs9OZsmbSrbbVk2vdih4ieheSgZNzvCO8
jzuIzlCqdobgJpLusYqoTMubNJBcQLSOIPvlujBbTjr/dLwL9UYGUEFLNj/HgSk8TvOWmXNODmda
SXMPcXPhz12nK+XpK+89zZhC6+p8/DREzyIBidIUiqg86AqFWB2IaS62IW49OPpDKXiKy5kX2uKC
XQL1bVchnc+uwARejW+SPhwiIc4/Efu9Ad2gZT0vPWP0cDvEDxFxXeIKgOIuTJPwmHRrZiefGa0w
FTed53z9A8PWaklcwZNwswbt8IE+utV4pgcClP6VY4eOVeOSvcukg6gIW6opWbIlv3K7KbjnkOpS
YsRueyICaj5UH7eUFriB/r3OJYJi469nuzhvBjBUp6HJkWG2KsIZzX9T8bqa2AIeqr1ag6ziGd0P
VXtRmVbst+705fJQyvBBaNMeEbbS+iF5VUXsYmB3CrVHDl97hp2wZsnaDmbVj5BLCFojTRcDSpmk
SOuz+YULVNhNLRHgoJCAQ9knOt0VI2kSDMoNuibEfRV42d8pD4LlPnbvFSK58vs2SXjSwkp+mEYN
pviCC/I55KpxniDtzeQRJV6qqNBOsLDV3P41Hr+i/thP/JiWbLR+WSUvxaBp8CvdhBDYVk9jiKUY
6SoFfiqnmaCS3C8JS/UVvXoq4x2EAAxbcgxjID9Kq2DThUM2dnMG9EL39sUGKj1POYXEa2oxJ+r4
W0DbzM10lhLWoksc2Ou0ppRa5+/Z4jiUR6HHBML1fg7x+VmEWGVtCh2PnjfKcwwgjU06A/McTN/O
cLkDxJ+A86fPzVSAqErCT13SHH1xfZ7lIVGlIstkw7pxYIDGtS8pMPiplO1AltiRip0wJCmLurMb
W6efc7sladf2SZh7xydvyiE+yqlGsd+1bERs9F87YF9mUubrPczvitySfUo/uAp01jW8jwnrUnLW
pHexlulXfDKWdMzX5nr1a6Osal1I68YcQzBAunBEcwlfEdg1yf7GITtp1+b2b402YQ+thEk9vmRH
vibXz9Hk3N7WitZyKzMfAyySMcnXF9VXRbb/8zFUiW2aC/L8+KTCVXDw7fJHrjwnwhf9f8u3bmK0
OEwxr7GEY32D13CxSFu5PpxiTCKD9K96NhCb6pYK4qGJUS68Qfk8MBFp55+9A+6cCSzclnpa2+MO
20mxuqBiKynZx3hmZcR72++RWo8ne/FfTwaNPpGuPdKZuLhb8jrE1bEEnhi7R3L8bfxmkxQdZ5+m
Z6xDxT5uHI0foEx2wAMNR+xHwUT/i9bTlF1f2IWw4YgToYomIj45QDbpOVG8C+AUZ7h3w7quhbay
lb697azF0D+x1FytfeT1SQuAB3rQ3LY7Lk/XeLVaE3crgtM6suCHZkD/Ep6+Wl+D4m1AN+2+WER2
kXUbheM1YlanKL8fGUsg7BFcRTBhlrOK5hDDoZ27iwS4eHFWMs6PNnhP/8xwmT4pyxGs8VGpqGsK
tHq06NVBGmyeY6Lx2CV9gW8K3iDuelIf/RnA+wbcljE4N6M1ixBrAvXfq3eqlWTwDJcBYNbAmMN/
hE8rG6uldQ2hiqTLTcoe/aRmF88Hi6uoP3rYgwBOTAdhjzSJERIWHH8g+9XQfcDIVKTCHp61Hd0P
qg8d03jI8vvhVf1ofByhku6Z3Arj5iiCAj5nkmAsEUehl6OtDly71uG45Z8gCUPTBWnQpBXehY+3
E5tSDD9jgDDlEFBB0zfmFDSPvCsJgMagRrELDzRVOrjV3lRCOhsV0H27UY+aW4yJOLbSF+05xecd
o3XZK0uCq5rjFTlZ0TkYCw4ud+LgO4xJ2XCGVneos0eF5pP5EqDu1QxcoLm6ZBC3IitSc0VPU7He
WdW6QE7jTDbQVYdk6UXr9ATcJko0+uIAKKf3+wPAgQTPM/rV8s6i3WWDTQwAyHiZzxPOh6ezm5X6
cmIPqC6j0GM8aVXFsXiwmoy1ucGNRcebmbozl8FSWBdJ8cNr2lsNGnjCpwj2PARwEP95+9N4g1Ib
HzIa8BSnoMQFkQv6UHfd0t0CwH98V/WhXfh+D6vC9mYnSVGiHC7fPP9bdxy80a0J1Dlok34R5CFF
IZvrgMvfxyxOLB3QD4LKndlTjudgaaN8Mi7ja8YocyhV4wMKUn22+/QbdGg+6rcLQET02KQTOUCi
qLSPhx+FABYnNcNDF1nnkbUN90dUkMtoPkp9/9F3V/7KzJEYCgRdxXCJOHAuNujkYLFl9oBgn+2/
yeltR+nsbJ0m5iu1FSolYM8IjddAFFCNQ0aEFn10jrmTVYfBkLOoAjAwyRK6Wd3w3RUraaE0CO9y
lFyFD8p2hsAoqZFmlwEU2mxq7xdjfrOv3YjH6dn42RaThu/03TUEYf3kNYwoptl8uD4RsAHKgpTz
+8JUOkH4qm8l2XLnHp1sLRurjJfV/bf9/EASS/ypDQ0wIzsNiUm4GEXDi/O3xz5iF5OCF2GejxWw
w/Z2U2trM4c4II1522jIzDD9KY5O7DvHnFfKUgrYFjdk771NLsHIgmPp1SODBer/vY4oZY/8SMRh
CUKzVjks8BfDxs0W0335ezTpgoTMJG3R2JJO0r7aSlzFPKPrRFs6TDyJCVe8MnQaZCMVhEYjyg29
mubxP+OMX3YxlKY8ecfRyosiQvMR2WdQSdXyBqiDbs5DE2mEvHIMsbvW1JHFuVSri1PpGefTyKYJ
P6uDP2Dc/L9aqjwkjOe4N7lPF2bVaL+BNenJc1m13QICrrcG/QoQtLRX4dSgmDyYyUSbRvb8huTH
NQzWAUUH5DpMLrlF5djXpMO5Dws2F2io0DyOGjKzGXI5lP81HuU+nmVFk6mekWuxaCHb0P4if/At
nRO9klPGsTJDyMjTXIfrK2k/bfblHW8KLpWF+/EaJHodqeWbzPnO/zA/XbqESbCDowQaTPBy/TFM
BBlmQapjmzN84nJ0nwdYKBJ6uh1Clggmini8sWHWNDiAuOKeajDpxtsy7yFrwYryCLUtyLBH4whr
SqYZX5ctuNl9ML0IwB6t5SFzq9lNJFXV9iw71pmz27HbQqKbj1xXXQLfMlnyXIPnVUjiLjf4ObrM
b/39GvssIzgdeHivhv653VWjEj8I/YUaW3uq1AIjdVQqaq2OHW1eLhzMA6Y35YKgtJqyaaaf30Ir
YGfg7nmHdfe+aF5dFsagIafbuRs6tK35bVYvj7fRrU7DzzxGlsQjVL3ZGFMY4/V5DxbPpX5Qvosf
THX/StZwrE95ACmwg3rGt+BxpjLN5iHQm2TBmVcVQKXiAOns7y5bX3DiwoxhdZ89NuwD/pYQSRUi
Pz1QTPiUoxGek5dwcyuI/F7jzaKCy57I7f93YqXxSCyyVnKKHeGb2RHLOeHjqAEK3ClcZurkM6vU
oKFQ1DGIrcV0W9YqrFvux+YYRXL2EJAROcVVpaWEKbnbsRvKubzrXrKfVJlhOHs+OULbaYwIFvsq
/AVWCdrr6PNrvrGPC7dp7dikiU5n2yYbl14wiFZJKEuo/9gTCBszzd/qEErQB0dqhl3n5qLlpY9m
c5+blyL3eEtT1WS22tGgovNQ8o9Lg4V0r8vEZr65fuN+fl4zKDJUuBgHVj8Tv8P7sgpXfpO3moBF
P2FRW+XufZvtN1kQx2GzNqSJRGZ9YohntgNkN8mVUXUgNxT3KeeC+uYINner6/F90xBEmXMYGdoj
7kCrnuscADAyo5vb82+kg1zFjPeuhZ242JDa9vP7N/cIj+Q0U3UfcTnH0vV4WpG1TzCbEimMyOG8
Yghoxk1idSQWWfRmAi8wYd8EWLRgKncoLTcs4w31wmGCwTmehvMWWVV5e7qMfEx5hRM+BSNRYWbi
eXGWAAlqVpC5t6prEC2HrC3tm/rsqyqVaqD/BA4+vFSJBLdnZwx+Ch7n+vxZ3hGN2liWnFllh3IG
J7M5Wz+jN85wqdzc0z2Y8kmk9byWaZSIBRfenr4s27Dh04Hs5pQcBu6qyPA/w4c+bfkUXD8aw1lE
2U6Hqclyb4S50aOi1Vr7U6mLao3Bz+L6kZQdIP7LkBY5Q+Uh2cBdyvV3Jfyka2dB0SjeQpxNKTbW
7f1hb+1yZ4Kf8f9AaB3PICktt+etzXLNQjMZZjYKsmNRZdbE2/S/60FMXDia5Sgq3eGkRAuz2WSa
qqZrix0iwMgZBQYXH0RISl7kMIgIzv5Mw50iqPCHeOGP3wZOyfjSoBthbXLc4eAO1gvM++RYPxvO
ulWMAWAUxoASga94NGomtSmswV1zmdLFBA0NxNVKcj+to4QCYAbRPRsTDfP9vKApSEhqpJ/6yXfx
LuSyfrYUt7KkqWb2QB47+s3YQzrkjpj4YTeYwQcNrJK4Ak2Kc8BfHW12EmAR+THMHxoaAgrc1035
8Z4cc31iJtFaIeDizcqFjLx3oEBxubGgR96+U66voCX93Pppn0siCbgnTeTS+MRlbZ/rGBAb+5NB
h7c6kPsI4TUingGRT79eOoEyVkto+uDwRgR8F7jNTar9WQvV9SnkbViy7jXtLlrNwCOnM3bL3+i+
LMB7S3mOI1yZk8B3vx02shiL77F/93cxb6WGbLoPDukX2T7mEIYaBM6KzvsOOcWdZybHIoqOAOy3
rpPKDSZND3vt08JUjdJHJz/g8qmL9mA3qpHqdglgQA5JXeTmkepelr8jknPkM98esRYr/5DwkQNl
vOwuzm/9tfLQtyqrEVUlpgp7MeE42yiCd6cHIx1svCFYQi9pNeUbpF1rdmi7vYZwhflqBtaIMgmy
e+PqBdxDu5UhtXxtbXbfchBqfrwjLUsdrEhjZVbNmhS5xqeNG2GaCz3eKCkwYnMb85Z+2B/RlzZG
ly05SJ/K3eKFDF6Emcs+hNw7x0iz0usqUwr6M7FU0t8BrVxyw6WC1Fk368+fzgGFLDhgIjI4vT4U
ZyhpntEPRvD7R80hgv2Pc17T9AeMHEXE7cS2BFzWENenW8L8cFCOdGxknexiRhxvPQofeUDhtEwS
/onA8/Z7XgsyXAl+Pid3aWJZkw5lM9KNzbsDcTxNVMR3Yqyokua19CuQM/34fg2ZhHZ9YODnzcvF
tDDOt+evFSLrdO7vPB9ydGt8xOb3jtg/FtcmU8y44I9PST81+uwR9cbYbBiIzJnceUgabzwknuOZ
0VC3XMoI8B0ZufsqAnebdjL6W6O7i0QsYH1ij8FzMhcs/nwVlXxBl4JOzxSEI87aGuGacFo3aWpX
nevuaKmsh4NPIAwHy1onU1NSetZechrVwi82TZPUXEgUuvBaCmSVLDswy3fQgdvTcTwh21fr6aZW
+7JnX8NJJzeHhu25gmsUNOcArb1k3MC6BNGp86+fkp/nlSrbYqQWFxQp/53M1pleWX9i6RkPFkk9
wtYVd9YWvt+VC0m3prUkEgpf3XNdBVc/MJjtdZAUg2R/kqbMsb+0STSAJ1LQ9w/XpIO7lwNWlayB
RwFFKBCMhr/j0RisnkOkrgqQNgn+To4W9j7/cHRIuYDBSKTv+2dOKKVIi7rsktWhWBpiS5/ZxY4w
VG1XLGX64I6RPP075uVqdtcIBsBIDkBkEaKQvcNeFzH/YO2z1xIDNf3fPJ86x9q7TwtXLhJpdEwA
/rFZ57LY0Va/U6QGFWYH7t9rnYssiNdoSD61sz/VoHie87A0bSozsFe3qJDFu+vs7fwtfLljNwBq
yQ8IJ1lKKxg5xDPqStxFq5DSz7n92pIQxxVpWwgK7/8zoWt2BJwGSDQDJn10CM6XDTBwnIWzR/PT
bjoroQ/vPLFa2d7D2HQ/oQ/a3WVAKk2c6l+wBPxGo9/7g4enTYokGR4PRyO54NiHZ+IxNb6GIR6c
++QIgGEuqRLBhCnu1fqo0g0KPUJ3z0rOBOgxrVpoEigWWTQ2NUBjQRzgyDLkPAUUVGorVAHffCeo
qGc/mw86kl3GS3jfls97wTVupjip+r/QL2CixuDwKVBFljOR21E+5GhEQBZg9rej0w9WAkuNUJdR
0NcNgZpTPdQT/tr68w1wsmnqvobJfHFC1pwsefnZqcy8AzxoiiaIyT6TltTjEkFGzVpzmsTr4jKV
w85X4AXLxmXLdgC8P9Q1ofooPdU/bh/Su8YEQniCE0bVEUlJFa8md7p+rpuPQE+qpVJve+NiIHpi
+6l5f1NEAKo/ojmiby5lBur+S5SaQahkYPQ8sS/TiIIEaFgNDwsQ6RjNG5qQYNDnDw9SGfV6c58B
u5zMAttj1ECdKnBDBqm54QQQWBpmjgmxzO3s/iir+9d5MJ6+4rQzr1TprZUdTT+o3uijt0ITX4nk
LOU5903VsdhCxuJLMxGJkXTHblBkZZg9aewnB9Dsh+gdWoMtYIwOy9Hxea+/UTOTRBndLz5bv3sD
iKmYC2S4xykrGELxIRPlxxW5rMXRbNSbVbQC/NCeF196DzCytQUH+wGcah2w9vUd2khhkGpYsRFd
BMH3qgWlQD1mcBM5F7Lm8v8d18BjE04dMIPgVDF4l/bnkri9zvz8teL65v3gh3xa38JW8VrmJCBe
tehytg8wX9y+yKDzB5ycxrZiSEnzsSA+ifJ1WDNSt5AS1H2Uwbny/pHSZlZSAUybbaP84Or3knI+
2RpSfIcT1KtdSAJEyp+OTgR45BctZUGBTQxl2V1vsjWHXCVgLLBLk9COPWZwV6HUZyrgcaG+qnYL
nrNax1sdQdQDz8pE0ydIKX5pPU5k8OH1UkEchBeAtdtGGcLWCpjrtP95WSlADMwHLT0m8tFUxI8e
ja09czL3xunhFbp2zMGMpJnpSqdRZPTNhsz6iRajsrmgPbyKTu5iA/cFJeJxVCMGZdlNyUeW1A9f
I7XgyH7uKiE4yZAD6ig9KZZHYkn3LCJ8xA5BA45PJXkT5So1von/WDI8hWFvWm7x2pZluNj2KCOt
j683zqOpQpZBIP5fWLxtCzUZvewSRXxqDjz8pSpbmWe9Jw3bWx4qZbA0kRPAHv5zQE9sSRBQtFTf
WdNyYg8ttfU42G6B2miakUzzMkNw2AoG7iT2SHdEl0Jeej3t8aD5oVT+7/HQnOo+dK5YHPpVzZdU
3rJRSGx40BHfGzJiyaYiumIKaxYR8/UB/g7sg5qg77CS5HgdBTwojxYT1rWOf8XckDYBLUjLcmDy
PvfG/e9ZLx+s+Qr5Wd84SM+bRaS/wlllVNgVehgOAYydknSeOfxDuJMnFkCXSzIiaQf2Mm4bqQXp
YBJWE00K5k9uYEQ+opvsGppejI9ZscXBt5stdP+bomYRbAnRKgLBdEhmBENmkWAHgd9Ez1g1EDk9
9y0aWc2xOqaB7XA7vyUH2KsK6VOgxg9EZdxcg5MXZuMpBPmZemxri7IcNBU4MwOY8nAK1//lIwNM
ebDhjQjHvKsKjgCY88EWqN7EYYmdwkzqZLB62x655xg30Xp/DTefzfMDmKYyQNcT9+biocvgBj+S
P4AoOpgUqjeheDqRDItR2R2uVTtWXTU8mDF5gzBnxHunoKlIKjVib86ZyjxwDqOkxwiXI0c24ltz
23g1nTnbza+7m6i++Z/7A4qcdT8Bc4x4RtjVPkwoivoWdbEoX51EkR7ocF1Glc1b/pC6PvgBGFlg
Oo8TBK6e94c32X8+yi+u4N9Dd45bGCgrNc0BmfSmYPEmKvC+zRBwAwrRq62l3imUH85P294MMVzZ
mnS2H6Iez4UMYUjXNJVGdv52J1yw+rAF8lq+1IHBQbp02G/azF4wwJfxm7jsX5PyWMWkSgTAX98C
KcTSquUWMV7BJtTbx88TwJUnm/X2ug+C6Fmk1hCMpjt/KgmXs9e2PG16Oogf1H8pPbDfC8mYT4Ip
xV5ihdoNTW+D7Yji+9XSlIl5vUosM2TnHHv392Y4agtIgJzWE/GwLzho3q8LNZcEXCqrb8Bpk0t3
tM2ApEIVM9q+qu6CUEsX2gVKaDQAlhacHqNpMHpOD0qQ21tp+9/UE0hJuf7Jl5OtIT13urCLSc9M
eVjnJHPVQVTKJsJRlDKiIMmxN7vdwqY1rH+/3/yqWpm1sVbO55jLc0/JmVt1cQKsVJAwz+RL7roh
V9zmSaom9mokO+Ch3qEJHgHST8E6NDmtb82KA2/0jRbK17405IQJb0L7tFWw2CorzDeD5PzD5CEA
Thj5FuuW83XIRGQlCco0kt7RRKQ6lyn/9yZupZ/7KK4tVlTsfM9ymrcSZr90QXrBTlcyaEcRJtcA
E3SRTzRXSS1JidPziqLrZYr18/ieaLP1yxRrzy46EgAkwlOai+SmSzP4/0jklYMxSsH+4FXi1hAQ
ln/2KNOl2vilrmBeUhrAq0PB88jVYmIcpz1EFDQIvqGloTW8LJbZskd0v3OEmwPsmbRlckSlsL4F
Ua4nyMh1upbSVdCKpVpJ49w496/d6zqR61fS/K5d4X+jO/OvDB6NFgMLWqNeZNAwP3to3RmIhAry
FiwMjc3GtzJrYtv0DCqij/hAcG4r/1Bt1PLNSDYlCzQJg0wKLgC8p/+gIM/M6b7jZPCYCFTMTtA0
AN3Qn4vIv88IDUU8ykx38CdOzIBcvNdQRu9Dn8hRJrdIY+fM3KCChDGPzK78PSJ2n0OLhdxUFTGh
+amdUK6c5qKfAClQ+wEqG+YAHHhsox83FTQuSXiywH3LLmAAk/7OK3eyRYbRWcHBgbcovIAPuYYq
gwJWs7Q1VCXaE4ymMu4s1+T93C+FVs4k/vU+QAdVsDoqoyDINNx9MkimmW8IMtr1fWublVluG5CL
oK5eF3Wv49JE3ohAyYgRh2HRhMpKyoNYImHCTFgCIZpbNpBXxZ53sxy+a0BI+KfvUUOR7ixPqPhS
14W9OFHAUWV4NnUCg0c/KfPWfL5tqm7fQocB4e78Z4UhPnWUBRXUss85LL6nKOjHbpqPv3cEGNN3
yTNHJ/ZiohdpVJInc6PzU2zhSErAdU72ywTDToUSCNVtiAoYgmbs9P4t33wMgcpiqpTJdHNKHVR0
g2+JxzW3zZpT3jVYGYA/d1BbhYOPxOx5ts5zv0rRlQ9eJwL9Tnfcoxj/BEvbvkuaPGJNZ4KZDWtr
5Xh91NevpUDTIVmgKEaz8imE/Jv3l6TaD+FsHnI9ZkrOycnsNdPZl0PmexwI+hO3NKWUJ76vB47T
O6hW2htsvtqSE434cCCiW3EEunmtlTcY5dphnNEjPQTFW9G4gowwfk5wy7WyPN8dYIMFFT+22Btd
3Tu5gur2fAhh5OEFTK1h2eniJSwmxJ7lwN37pzK/VLpF8jzOPjhuJAtiukYRh3H6W2hfoSLxiJXC
Rh8MlrvZ5jT8IzPaZqSAbqL7H34gvF4l8t9uVy5lxKCemCc5UmmPWdn3Mgsiqq2SsTkHxBaqnOwu
RSS3+ewk/zcS2IJwPva/vuXe/3y+cFRc+zaafnF4slfZjkG+55mv6T3hUhCDrs3TT+CogCm5f1aL
fIsM2jE4sgrI5SRikCwc01GZyw7nAdRJAWtgukh6AwFtA9AbQ++sS0e+T2rD3bTI1gp6EzUts3Xi
HCl9G2SH3odsKqQih1ITExYn4GwG5AWO9K3LunLdb1pumQ2Sx3Dw4d20f77o3rOTEdsyJbhXsE7D
Pv7HtF9kn0kqwTPKZstDvyKKF0UUJvbTULgNrHBCGBDaJB6EWxEbMKTb7WDM3wbtpPDnNpO2iLlL
d9E+AIyRElKMXvo4MJ8T1QZjUSKR3GhNmdm5F1GngBK+fZA0qNiSH1ZKxnb8WH8+Nn/4C7pw6Byi
GN4jJCJYovH/KPL+YUSmsruszENbf8qRUro/c/wqB38xbIBZ5KcYdqMUhYmNVlsT1ZmjCKVobBVf
L+WJtg8/16TA40lt5ElSCFPVaevgWw4F1bSVErnPsH9gy9ZH9EZ0lB2RKg1Vc2AAixtsfNgi1F/J
eK6i5XKHSQYOCRP7eEliPxK1/s0F6SVkEGwVzk6KYvmMeBuvPL4AJnPKvJ98UCQxo0dTMiyOtdaQ
zor96k5JHF7kNNL+LcsOfFtVdvApfst+y1DNZ6/H0YW2n2LgLsuNKTu8/NEqtEKBT5whKU/D3kTF
82kk0g7uNFFeUeJfvIIs0JGaYINMoToBx44BsWepwNq3NnkmfH3qtKGvf51dLZTqbOjgm/ms1zbQ
G0ir8WLCTDoIRJKN/xjyxpFczLpZGeaHHeBQmkQoESNdB1hJf3iSRYsdd2JSOpMMIWE+WU03cpJ/
MYoF/aFy3dgAedRtKIjYIytSA2V9G7actI/15jqo2flNR/nWaFZ4wV7/3p8H71ioLKPW68Hcf7II
eKKPynxItuCHCFGUQ76kqqlo/9v+TCg2QBA36svfq7m8W8z63sNhEto0UIz4eOQLlpLuoFM+X43c
2nrhJ4dfj269GSHdxTM0Ugd+daASo9fQ8iLpMAj3vYuYD04HvrPBDkntNyIMzuHaa1WLP/Lg049S
1KzX7tCfzDGZMJD8J9D6WNSWa3T0nH9i8p7+oYN8pgyWd9jmah9vCikQEaJ7NiveFmM7Bt5ptmrI
jt/GGYtfcHFdgfX7gTOZ3iKm6vXsp21YCqGxmFOWFi6Dsu3sdjjhhpI6f+pe5T7SRHeChWuvYuux
+iN4aVrRvfEG3HH6UNml7zkM/MFiGjclOOPC/qetv4q5Lv/MhrBGPopYP5Tlu9agPgnx25Bp27ZL
yvaxvhxmjzh0tkgZ3E9QOZvTdIPYJc5d170ltUUUVpd9BMyj1YZxrUObcORCVj+iEjf/leezHDtQ
reziVmqgZWBTE8GRA1ZUNXvv2MFH86VZr9aWymy0m1s5+5ZqqVWHCoBlksPyU8qNC+t2puwf9GSx
MeAPtrAwCnLuw13ffw524uVeC7KXj/rC/HDwq2M9VFD8+Ho/EF6IFAWTxrtLsT5pXo7Yih+UTemx
NZqNnv3NUFYP3CYl4OQi8vyLjnj3z3rOreSnIQkf+82enM0MyctG7EFOADuP03pY/67NcNzow0lJ
IsO1V82Oonp+P5xJn3LdPdRtRCjvFKsYpVMkcuj3Pujssi138wwrYZTyOQ2fB7Q/uhsnHyRhPko8
TPbjy6ilXkXvIdXWtC4mOtqRBeUulZdVBTLV+jzDa+l39jLGwQvLDOuSMvQjhixM0BePCJ5HCKIv
XRBXLT+p59PVmEPfDqwvyly/IWYf3gXWQYu1eumZSLTJaOA7opEUU2dAkVavLZM+RI9xv9gro8yF
QDdDRSB+yEMtfUqJRGoW7Lsdlu6VBwOw3F0XwoKjfmLZA95DvaeJfhWZexItyed0OLF1E3HnzMT8
JNxJAYWzkeWRa2PGUHFy4CzEnuTqf8KmrJ1hlYTSTqNJdgghQnPt+tpiefdJwng33W+JEDwBZiHG
zqiZgR5LAUehwBUDD89ulpBcnp47YNkzMKpnbl7oHk41x75kMBFktr4nl81JZoMI6NizFL4p3oag
iPzTzZ1XELXfqOqxX/6EBVLO/PlSsqgQu64yEUwWWIbUjo7N0wok0fIPLBEUCpX/d5XHOOIWMPjE
emBwwVFSL5mQkMeAk6+z0gWPD4M+8AZDI6C858jT9Bdpr9SlrZQEn6ThcO7ztBwLVaf6xV/JPJbp
GC4tXj3U52hfobi/L0RmKF5vEB/rawSx9Y6ssQysok/cxTm8BTBmSRwMg+AVH8OI6xpTYuSDZvhZ
J+uDZX/f6CqP/O9z3VojaM9NdRtkE5ImNMjb+J14a0cT81mJBipFsCXrXxjFJJZaMYo7uugGjhO8
Q2vaS4nDbtF712SqRRu4D6U1zPLgcPraqJxH4jqEiNNeZNdnNejDfIO2+P+GSZGfrJfvbHsKdBKz
M0UT/XtFZtpEqb5Rs6CZEkvHaoXlF5VyABxYhaQbbYh/aCOhe7j3guCTJNHui2GX1AxZ+tGiCcyE
cHdYizW00M0UWfWqg3Ao0zo4GBPFRSZKCIY0jXsXtrOUmPqU+G/sJAc8AkJfrayv2PPePKDARQvW
uOEdYKh2HCHfgGVHLKjmfehyO2PKo/urHhpI1CLLsynDhTNr1pSNHCb2OoSL5drmmKpvl909KlBZ
LuUWOKGiGhFAUR2lemk5aVv0KR4hSc55XYFWFiPbg7xOIjEFh3dc0VjwI3mkY/XzR88qvOA715mx
AwvUltCYiroceAReOFb5B9cD3I4YbAgtGMbfoHlOqNPxMVDpNPPkCQH4ANejUPJvBcgOwaq27Fvm
7KH/ky2dMbz+pKhjMEtc/kZmvr/DqrhX8yGNfhfRPOmItDkbNHpuU8NDc74lbq4TarsjX0ukRePb
pp8KSWGtczh4Y/VNEkYlu64H0ZkRPj6UfdKaaWwHLOEhdYXzSf5xnuZKRYXvGJxpFAPmttSnwPV2
N7ZPkrBLUsNu8XwjtTVHMzDFNtMdhoLxYpRMRydc0ubReq/wIydCujC92u3e13F745ffCTn7ojCr
zHnBSIQJ8xCs4zdW5AJ6KyTOTcljuC7cF+9tLnndYemhzBCOgM9Ge3nNiHEBo5b5nGwlpgx1YZ0e
tK9GcLNCf+Q1tKwv45U2QzpmWxybLOmpZjOCW95bdkjXbDR+3XIY7fRDbhRLPt4y7MKtCcYnn4YX
HSg4EjWD+b5HfqOUNGKp822yphixbSSDNuuDkljLyuFq7Pr0oqIrIahm3W5VsDA5YNUY/rdWmewe
26wZ9rNYtYH5MkBHK5P1RFcJ9Q/nwfKDlQSu71kUJnpst00QzmUxJuuikyWKc2mAiNl5CRU+vbEA
6G8tXTc3cN2ZnLMz1qELQzbBbYnoD5RUqBxYrHtc9K7uuXJJhhKGb02SMJGJDYLQoLUkT3di3Wfe
j/juOs+Py4UKdvv+cku5qen9PyvcZclIWEq0fpEA3B8XvyiulJQMyrjVQ+XGW/3U9hsyJVRwCFOW
LVtWbDKO+qp2KiiFB666OAJxDouBRJzsKvuUZAKngEhfdaTLFZwRPodH8rH3Ve8BgEgeVaL7cj5q
UN4Gw5ph5tc91A2W8Mmpp9JUyrAK1bbDR0tB1u/aSq2Iq/981UAeV2nZ8tnYpLhvbkZRaZnyvqOb
P0eIlSyxxAWlJjwm7AaggD2MGCOMRDPwDiPY59e9cYH78RIvtCc/1gKFZCXzuJnjj56n/6ZnR8Pq
5LUPiV9X3OYKALi4NuAwstY/tPWc/ohqYl7hGbUjemdDjFpcTDEjTxVwNLmM+/L43yF3OLRvp6vK
hNNGAgnBDy8ITZMQdtA633i7fS1DeXnE6QGVHyJ7afYkGxi/bla8XfLsj0wV4NGke6SI94qqbBPd
rJnrW8LMxlkZ2v6VVtU4s53jyjDgmewByzJ5+1Z6Q0bw7z4FLceNP6LBMdgaDHR9S0Xn5zqfx+mw
IcyZTOj762CzY7xgIyoJfT4Ucm0APqQXa4jChshMp6LfV4pzQl0xjUmjKtpZ0d3/ecqYnZhv24gg
gx9aomBKeuKyCbIYliX7aLuAHczTu/lb4sdzx5CquKfH8slhUGytCvA5wc9yibRDU8it5ozYMOkr
ZOp2MjzbR6NrRntbXiYXrowMv0WLXT2Vu+fY8YphbSNl5/ZV6fZnhXoR2wKm+p3tfdOR8uPNYmNb
BXgX1+wUW5+ZFxV8jDp0Mplc5/sNXe4NYIK6VbwjwPtcRStdU6CH7y5oMaIMZf869oIVnwzI67c4
Sh+8vdvdRdSu7Aeua841Agkikxj8h7pwJggslO7fzSBRP4DSXEwtETItM2NOqQ17eGGBIsxQddBY
bIyCqDyS8MPhvjuSH3yIsjtKVvDldwVGtIRcN/ML8L56m518q1atXX5AmnUVpKtZhWlnb7ISLGgZ
Z5eyv79X5VoWpfOggN8oD0QGupZQEOP7vj4T1QZxqlBpXhRamWiw51ghNV/xieOh4S9lpoGn3rTp
FeYIhmEfNADWQ020sQEBg1hSeHC26pJ10Lxntm4shu9bw2IKZKn1Mh9fVzPyr2GBqQceo4zm7tSD
aWFTLTa7A5ZCzyqweZY1qSkOWw43WgOLTby2lJTfSK5yF0tzn4zZhWpXGviDVocDvaGvnh/SoWp9
8ShbONyuwFGNu+x4aC5+0iAookN1NApFVJs6jxxq2kob8NWtF/pLgk/dhfeAxHx2E76G+VTajKYI
J+UB91cL9cOicwVS6oj1SvuPThXXyM666brB6sdhtHfT6z8OffLBcRbPelMVKiwpJJ9HPJFsoxTi
yozN7kG0xkiuuxBZxmxSdsiNkf0BVKA8DgR4xP0+Imrv4y+I1Tqd3WehybQCyYlW73KPHNcuo7NO
EBIbP2CYHAUCed3sMMZPInP8jyYYDTSLQrZKVXdjryMDOaGs8xhD+aT2A1UQudk7XoJFEttePr6O
hmvGJUmJaFLorg5gcnWOMrQG6Zrx9QZR9Y/Hn+wGbv4az6+E7gPYPf8W01zoLSjZ5WdeigZyXSmS
X/68iwr+s7fdFqP4rR64wuyT84hHPUmRT+GGS5cngxAvAarho6UFxj7b1bX2arKiez8haW2Q/5wZ
dqT71b31vcdJKU5ASSHJ5ytuAAxbrrrdYnd3+vSVDZ3VJaDpnwIYejULOmh2vkRztvOQXHFTmgCq
jsiguDZ3YDFHpedPCxpVBK3gMqnfZgTM8iBksQPbegEs6O2SZDyoHf5JKGvBjtwW6DPy7NFv/LEs
K+8ejgdU8WlWmwkNax0fwJ7f1q4lyxE7n3R1c80iiQBoblHFkbdyDYxYCoIawfqSbYssKaq0D2e4
vjYQJYpBYv9FOifjby+wnuVBwtaDrbcXMPsbNQ1MdFrriGHNG+zvnDcfAB/j/FmNQ415aWOB2Jzd
9quOTShNvzi7cxn4o8U6UzOqqAM8TuORTBeFdLCF1wXlSe4cVQ5R1vo4W3N8ksnHMfRu8JWZbfrI
EfueBD9YMg8knN0MQCeNkjZRzFlOUTndQiMa2ws/iOXYrB8GECCx4/i6f8T8FkQSThY2Mjg+O0X2
39WCsjPwA6irN+6Z814LJuW0ccixCH18iloILq/VVyPIWhTBDWTcdObXVvOXgGU9QubtHUI8oyE/
u1lMLuqqyBjvJaKUaZrLZrk9XNydK3iMidQ1gZNk6IUoSdVCslfUjGtmHIfbaA4Dk8HLk5Mlog3y
r+C5jQe3WI42U73DJvH69xryIpig+TfsokQ5sL24WnOvPepN45TMfVddyf9z6B6rOFpoRG0M/5lG
VjIGxzgNW/izKLiRjTi+TZiLm/OShCFgqXcJcSHqJiiYBneVy9/szOTVKwzlVly6hdh4K7GZ5yz9
dIR+ebX5GscyBU6CmQvQfpe66c9mc3D4igPXcrORcJ78fOGw1lnHD+uuMUhCq+dbDgYthf22ZK3p
qlRu1KjMLYnBBwpnjiADR115I41Q7prpFtzbY+kq4tuZmt/sU8kKu8+Sk54dbqKzl8HajyYbmqCm
REOn2bL1AZNcKMD4AU8GO3bEqMOLL8DL7MDohGPZDXx/PSbM19A98u+zQiis2jQte+9SOFrvvqtX
Qx2J/WwSanRKb4Zqr7OZuuIWbVQecOuoidaajU8DSlx+ET79rkoygfxhEryLvJDwLN3TFRpzPmga
N4VKSAa5FYCv4v/zJNxXqU4FSfaqmRJcjWpbL6R7inr8UYlxewcyWAd9HEhDx6XBs+H74kijpGrW
GQyDxuzcyo6kgg6SOZW/5EQL0YwFkQjQdz98m2OtpNWd7SMXWTr70GGe1ncdMpuEwuyTYbM7QDZ6
P/vFIl0GWbrPB9n8iqyAIiv6MhpM8n31Kote1pdH98vdSE6Q1fQO1kH0HaYKNS1Of+Xw6RLs8Yox
6knGVt45XX/p7IWKPUKSSbn7QHl4bdqKVetZ/6FJpEBeajaXh50kg5G2Uo5tho/TAofoW/t+vpSj
enWCSADUKWrl9+KrsA0JRrT5ZnMEqdAnwpzSLS8ub6RxBRm583m52Kxq8h1tBloK5gmzdRPA2XfF
2Xtw4Ss3tAinOa1r2ILd8Dthnswag6l4I7X2t4kkGIf4tZpZWF3rcBmurfCEp++NIHM5z83EBf+m
BSMsbx5X0u2QUR4oM+SRjMh2WcIStb1rhOcGwslMV97Ec9bzkbR/DKhRggD0IA/myAjz9HbBKmvY
zqP9kfc8xz5rKOgtqpUm/43ylfaVKv9UjN1n64d8Vlqxlckf9alj7vlvxWrFbDipp0ZK4yUvKvnk
x+9jFzMfl7gu39RdP/f9+TS5PGKdsqLonHQMkzQTVRB9FZBouf39l7YS7RLJAIRaycUBASiTekj8
7FxAt/Z1hgOAqnUzZ0nfEHmK7X9Ld8pFEHEDyK0ud2A9uFXtFxW0xNQRMbdMGVPmB9UcIlOMvqHf
DePJO1Glu2pIwBP93ZFqlATLc/pPK30E2E2CmZGGsRtWG4+S97Oe2Ab+RZA8WNh05XLgAXNnA6jU
xK5JBxGw2fg0GJy72oqa2+6h3tF98Oq3v3azx8OHDZHewo2y3ec4bxhr3WhTl53QjRDYBCrEEs+O
nzRFZmvC7hhSKelvAeJEPhQC0ZNrn3W0VcoPyZwTjtw4fV2pij836ko6WqZN3T4DysMBgE7qp6OQ
wNgWP6LPk8omWt+ZsF8t51xxKvp51Ak8iqiX6hjLHExbCKdx+anvfl1grA5pBpV5tiNlc6+DuE6j
KkvfrEQ41eSu72t2y4PKZ4v9yueryGAuOpjWhUSNeKy2dUqTCxNTnkZIAl/2jkGUofKED2Yl7bzG
l/trReGFyNWOQrpzlraUK/XSMRiiNArfVLZ/wm+zyvc6EmAXHC+JRm/zQ9JnE8omeilWQYpHnGs1
JE547PGIeU8PKk1ON72N7Mvx9bD+SPWiIdoee5bZ5vEBnpeBcWvN7anjTjOaH7jUcOUg75ooUHex
3RAVT2Z+vuW95niaYcLF6sGdi1ULPU8J6KeNleyIBgV8a94X0EHTv+/j19lRpVTU4DsSeXS8lJfY
D0t0qZcDjZXIYlCFhvI9iayZJkf0Ke1CCz7CjaLa63cAReeBk3ILYcm9ajGE0Wh1G+oPtO+SbyEj
8+zCVgqI+WRXogsKUcDZKPpOVk3y9WWAl8HNYtaBU+V8vke5cA5yVJVg89JsxE/sqXxsYRgyajg7
8p9qxNoNeGYZeSab4rKB2KVAHCeV5jHDrs/MgHDlU998wlQm39fOSCZOhk0rcnn9+NO2E/ebgYRC
k9dT5ccFAuLdDAS54Lbc8Ee5QH9x205OaRwUfk/A5H3T4mZdluM2l23f1VqW6eoqj21BBCe1UN0U
l5snpLhs0RAlmPpgJfwtXvL41j1RtvDIaNwPli62lWoSjHc3P1mDZXzYEy3DYbDHjLIuMSaOU9Fo
iv6HV/e6qBHijONOAH2PQ1jj1I5AMOpx7qZ7KJ+W0p6RrEDf51wuHyP83IeOO8jE3oLyE+BXYqx/
uAA5mifLSNzT0es84HssSCgje2HBot6/Q1y5twh6H+aaskp6Fcjgfzov8ADP4yywAfH1pNnNhirl
NIkME6X88eqkDmUAfkUHYjAiy81L4sdLuxGrUFy6XpAoCJ2GF4D4j+CiXp3A+x6je9ExRB57AMAc
58EnzDfb4LzHyH28/YMwxq8AwzrKOINyDDvLK0v1Aab3pEInQap46HQOPyyg23DVde06caIpZpnD
h092zrObXO704fMxLHfrDUsVGhkqPFfc4RMq9lO6XfFdXrJsBHpKzNkjXvK+f8WvrgVAefRnJTcu
Hk2M7Szfdkbu1vNtYwNz+ZHEopwPPqQVMf9zDmLWhZk9zqCYlxquxuwvzC1wZUZMDIaUdwi1K6Rd
f87qvj73EVw977PBKMpSye0P/FppQqTdnTE9gK95EnqPxtq/Mmkf9VfAdoWb1Tc6yGUZYVvtGOl9
OttoUxGYMLVy0hjV89dlCdc3sPFPW/us4u3HcQvXmvbdY3v5FKtA2jAP7x6fS7NlveR1sIBATcN0
vJxzuqMMk/89IhL76eO3S3/t5hG9ON3dZoZhDwjpxz8coyi+1nUWekCaQZo7/Yli5Wsawo4T/ChO
aJXeGDmC8DJRrmkPPzjt0qjpbAEB1ZE/QVXN3hL6JbEVOpjEu2RIEIyMwEtS/DpMAwy1g0M2y/Oo
+Qhg0reheFSVGSPdeUvHTEpKS5JmFo4hDeOziBHGrzmsoqz6GrA5m2P3BgDiwKOah93cCmL9Eu1Z
A1JkM9rlWe1BXNHh3/8erm4ehKMCYKc3TlKuqRWP/w4E/h4Y1SEisIWvJ8w9RSHni1J4b7xnRVpt
Lk+OE+et4KL6eTJHMxHm8KvP6WByAiBUzzly3rghglbtStTkSRJqRmQvWR5qrqDGx1FjS5v4jtWv
YutbSKMaUebvxMkO+k7mKMQuwEnU+DPhEZqPMYLPuXO6VHYwisiAq+7m1BKeXgNuXB73sUuyGx39
U5BPWbC3iFVyJXgafGTTavQ2MEY/CzskdjsCCuoE5cx5eX2a0j2tCLbfqxk9gNSg/Le33kza6oaL
GSEs0gCS1Fck69FGtkgSiSqxXPGX8lZnVywo8+S+79t8nX1ZBTsAmrEshaoOsQOUdvBCN4RCuDcj
ba/V1AXriGyLx/0agADtDwXIriB4pmbMgV8coL0YZ/T97XCabSdhBwCEQA28bAU9soSyT85SBu0/
t/oQSDCi3htcVtt06iOo0JspjiQDPY3fxUzHQ3jx/qoK7LfO78p6bNkSnzb2n7EsVXYoSmYzzlju
4HsF1vQcICiVU1nyrmlheh/JGbOKCjROSbGRI1xcBRr5ZKVn2rweW7S9poWVJfMQhaWOUIu1dfog
7yG4wp60YhRe8+JeM9aPXn+e+Il+b4YdpAKwOg6HXKNzwjvOncFJ+JCL8krW0XFdZPiP7WIUFAAa
04iYg8E3SdAgFW+CiOL5y2LL03mFfpqv8l3iSl112MVNn4C+YkOlAsULeKXxImlF+Aj2YDP3vvi6
sKMiLF1JODpSl6CRVZwaON2m9bi9/bU6MqPyIhqX4tT3WwbLNGkH734nGtEUQefANrWlBY9TH79f
gnOQr9Msb1oJilX0xpp24TbN/qUAbUyFVrBX+ZkpX+/6XEFHIW1h/oUAt8/TiPelH7EBPbrv5Met
yXR52zCvwulPLSQs9SchxTaIVw9KnB7u4r29fW7Ld9QKaTolCql7dHa8YHB8utjdqjiLKfVBDw/5
FjULaC1m5qmwQeG9YcvgAzxvjVmxGZSCNaH7KygaALBMbdAxPMGa3VP4tfukFzlsY8XBMHCkQic7
9hvbOehSmWKrdYLTpnq788EqT0+mCqeEEyKrNVdPLZalXjAsS90mBH8Kf4VlABGwbZOCNyNb+3I1
sQuI+wsAQuVaZ/uq3n87Ut2IOuBvcF0vdY791YDR4u/36tB47hyg/Cvx17F3ADHs8j5Bvj48tt/1
oZJ2ddMtFbND+5t3l5AbG7OpP+nB/smYFqhjQFTufHRMN/4QC3TFU1xMyCkhTqR2wKWF6RiAjMeR
gIjK/eXwDW4tt5Mts8KVaEGvnJ2gQ7KrxRMRnJZadGkX1UAK+0/LxjNv5lKCtxhCRBI8VZ1HbKtf
ANxTgu68Dmp4kkzqipyu0fHoV+f9e4vwdGQqznmwCXwBgd3w71cuSDuvPHe/EzLISIKq/6bZ8w5H
ts2srcZEnYycCQpCsizvdG+AX9rNh3oBjT0gZho0UB7qC5PRgCo6v6HHmzWeoIYmgxkZW2AHniql
jwyCwaiizJtDcJJQRP/d/O8NkrQaCLaLKbmDUYY8OY1iS1nqmGPA6EEj2Tk/FFC3k+JtXvWPgkAU
HcMSUsgnwL5YT7FY7buFtxJQontGGNvc+X4GZkKvuR2LphaF8QoylPYCmWThHoKm2/l8hRGonw4t
jP6opo5hARAPWvaYmPRbaFHgupfqmsVrhFaC76G5CSxVdL3i6u8wYw6XgUCA5zocFHI0sVICBIae
EeU79qRMu76nasrq7GlUWN2fS+yKD0G+VMp+/nhyLYG4J9FQJRpxZ2TmkwnUHIT37JEHs2nqzOJz
NM4MA+2BnY8dJeCpw0IfE/qhA5IRmDW6CsyqFIrTabCM3Sv4NzIoCembV+ys3ugNT4h9peXwNg8U
3gXdhKAb6HQjK5XYBeeLzpwyey11KEyyOXTovGleLY03UueYHZD8dP8Yo3uc5FKC6WIGMBAXtf3c
x1akUs9gKaR7qV5u+5ypxw3vvQauH6Vvfhh+esxzYI6ArhJySyC5Lzaz3R40VxUx7FtSuupaziZv
m45uedE7e5TTj+Qb/NS4PnTVGxHQTeofm/5pXIrneq+V8KEJmwYCX358Z24WcKKvqZSY1XiCTAD/
nq2nRpIAhkMInpgo4Oh7FPzw5o0FgzhC9XSUMbRvt9AzntALFdSDYkNKoZLYJamGh94FsFXsXei2
XGtsDCBR+gCONjZ1O2+GuGdD/p/iWvx/uqD/fIidiNLmP3+Qk17p28m+8TAObPEsfuWXGBLaNZTf
2tvHVVf0Rx72q/3N1jxzNMw6PWsOk6FHRcpbM4+i1zUTEwOobAYYVae9HKfLMlNkhRI1pYwR8NZX
e5duCd9DDH3a0gr3uL47mpNMHz3mXfz849KKmQHu2/S5FCZ679dGEolfsXUlJssEIpagxYQJM/YO
AYyjopUTDgWbzH2kqnmoBOZykwys8cXEZB1SDkp0LCLNnzuMXoh8k72b0xEujr2mnRcSPEa8jGAu
GEGU2uDIjaGsB98XiZuMcVzjty83hgaiR1jR9OhQAquou8rE7MDgWJT0C4mTHAk8HCWYJHUWhwqD
FKHPxLYnO2OoLLVVRKDDmKHxxPtxQucgouM+7shcW+A+jXfZULmIj7QkFTCXWFBTUTKVXxBawZMO
9OIGj+OnJYBbscz5k4/oDHJfrNAWFayEELRvhSdpdmkZziBO/NDR4EfwznUVh3F1zTPFTbWsgYFW
D1ru6+H3ptajQLogxwrjO3I+LDsMaTAubrYvR47xpw58UbwsqCgU1DjlMeZQilxvnBRZOfQnxhMn
24X+X+xZ2wy726qrgdwbc+zRhziTs+2VzzivUeRr9ohOTKdpSuGYEHWhrt4Z8MMYp4NRseG7wG3Q
sbNpSXsAZhgUslEFFxVTLHuw4WhS8AK/vGJlsyHKQsaIGhMWbK8wy3oXmmW4ZEU4nFJGfK3W7Bb2
/1FvEFnxNQEzAJ1ZrFW6nzvJMacrJnxYMNqlwXFjiPpUXYBBx7Mx5xbqX0CpX+8THcr3IWtZTtiR
oSOP+0f/VW5koy2oJXBZ4pOhQ0KADRz1ogc9boSfXELCqzzzrYXb7eFDI1KIsoudcovn8cKxTR6v
3gAyPs5fMbY5d6JcsQl5wWXwhexvea73NV5rM9nue0zWW4ZvtziMxEfYL4b26Z25IX2yl6qm1MeN
ybkZj6KsdWvrtX90qCo8fzbHxrf4dlkM9PRrS0EWLeqsB4Y4rHuGUO23IA/yIm+044t2y+vBxhvV
71NcHKFzQ4DdVYIuGt/6elA3KCd+1pArRDk+LoxBQLfghfdk2dC0j1L8ES2j/IwkuuwVXZF8B3G6
2++YZcyAgaMpNEgJdfWCvCFRd0Y7YLUBwuA7cGP5YVLzKdJzTwfQm5yKFW+XWo/Y6W3abP+LvJdL
9j2NDnidnE7B/8dlZGE4+pd6Rlm7xhpsoJ6DThlpITfKARWbk3I5gFGC+FYKqebLhJ7jICKNYOL0
EIAuJfwfZLQCyXt9SNJnZBavTzJZ/hJ/MOOfMuEmFqmyrUzqkbw3nXvFV0ofO7Ep3+EZqcyfcNOR
H9hT+eOdwxStjcDV4VX4trqx/3kFwKgka9MZ+ABCV28f4o+ty42SKdRBcIpgEATLucPfDNn9bLIq
jwHo+NCTM/nCHBg4qSIp14N9ttFN1tg5eId70xh3JaKiSdopOUlIdVm2pYcnj9iv+/6b+M1kLaMr
VoOwxRnzHvZtxSFhF7lgtSrKxW0hvu7m3rGwfkVeMr6I5Mh3gbuu9asAWyUZEJukT5Npy+Weo3ih
OjZLhYnBGOLuqWU56Fg+ODfJoJT6FiXzvFfior8tH/ZFJL7L+qN6484NV7nI3UX6BMHHmIlR4EYP
CQ36GnwL9M3jbS7aZlg4KZdnwWO1oVFbGaWkeuRdrm2lhLvX2HfgPVkTbORkoGeIBnwnn7NUKw1w
a/ngKb8Ml+ZBbeu1AICF5g8bhQ1ffY50nimPYfM58jXU02VHu7SXL0/VqnbEflv3jIGstiy1cX7t
dQmtyripskVpzMzxrIbwLfRP80NoXtBjH35ChaQ2Hli7Lhh/kYyRIU+xdrVcseT6UDF4LlkqxHW6
0Z1EKKMh+WPg0JQKOsd/WGhFw3/IYJZ1/FR0B+aVLBrFETxFR+OvQyNogC+FSEDXqYWsQ3wFWiJj
OJCX2HfmVj215bu2XjOT0UdyY1bZZhzsRyYN8b4SHZM/vxFMzwoEWMwfJfYlNi9N1Dqu3VqS4Zjj
KrSdD8VtkH5pd/JDNYeAvs8nOm7hM5XYQJApNn/eSZGS70pe1pQXlRDzBj84d8fwvsapPMYdzLf6
6FYmky5TP9XjzyesliQ5NRhx5woVsn1o8n7+7x6QXrJm+TU7ryneEL27r/X68B6UmHZ/Lj4IXJoJ
Wv2uFSXBzP8DBd7jyTOb19Tkz6SHVYDC0lgUEMAql33/Zb5mvKijmKcPlMVfvjVfHGOrhm6xNKny
ZVEFFVZGxVVwxj+7Q8ZzMW39eRNlKZIkLFynIEjltH+pPMpDnqn3FoHrlbwYL05DsA7zUarD7V1k
/C8TWo5xuw+7zrdUJqC2vEbeRGSRGeJqCESSvtcy9zJhYhJZ+lDmmBF6zlA0keScuQ0ryMEGEdf/
1E1VuZedBcDzr/4S4F6AQvHOiQBVrg35ZDIHzPYFnL7OmJDk5HwGyFhbs0jB5zvHqf/b4AdAsAvV
cqo+pp/3wX+L1UUT0agMoSCx2UHZF6vcIrDetMJdrzupSCTyq14+W2nBsQwaKh+XrqrBBUj8Z9sU
RI3O+ZGiVVrOFITNLPpLG0r+NlbERj1fASPHxJeP58xdEz5KEoWP1j5d+7LdkfJ+yj8DoxZ3rrE7
6L53/XUVWl49esn+lc0sdiLvg911xKntSxmenPXCKTWRZjJteN0NrKso5M12xydhcITlfRYUhFDr
ehb4vRc0jBxJ5N6h6cxAxd+Dwk0tpODNnubHBZQy+lyv68xU4HkG07dCWTgNGhcjThMYNdCr4YrO
o+x1PxScq7ktpeQZupU5Vmr/Nx9zfx+iofp61B54ohqZzcxiVLo13e4JoX0eYFyZCl9dWNdWg5bF
+t5gEWpwpvBVf/8jWA7PXuT+OoQ0EzaA3FS8ciSlVYzt1L1T1BspFiWHeWxz7TK3B0Wqungqapwo
u4eNM+qKhZCSrz8wpAwqMneFSNxB8xbCGK1HW5mzPMt3aumO4Hu0G6Novo1SMBXlcp8BD3hY0dsm
R85TgpRQi759+PaKBEsGMpP0QiISf/EuM5aLJslNILmusjpG/7ubonC2LTILotI6bChOmAZOL8fN
K3oYhfbnh3x566BXM4El8+jgITutzIM/ZBShpIFAntLC7qAfQ5b6aWdo8i81UY0NwcBAwaQW7p49
fnFg3oylIz0f9McswJSj95mRdJAZDjeXgzqWaY5R4Ti/JrL0VSZw94B/wYEet7Qu1oOprarYlbxv
oJwZdfa1DdmuSF3ZRYQ10EHe1ZxGvATVarIYOcGqCrK8Jkr7LN3H7L7iHa3WmHAwWrogM3hHyFad
OVEvJMq4I5gDdvmc0GTzncyBGt+aOakknptEcgwMDJX3gD0qMzpjwaCJor8fX//DqkgUHd3nTJ7n
/AovpmF3D7/U/ZwGZs9FwfE1ivLuwpndR8JiU4xEU/BYbqF0BtZ2qKDofC1FiWm3WXubd+dbLHI4
h7o7tp6QqJlEWW4rkmvC2WA20c1lJAoOAGa1zTDxpMUN6kPXOODRUxBaOZtcEgb/CRRwLZqc4yhz
FMQQnINl2Cx/5K4ZpdS8ZxWuQeLtYLJ5i+NZvvp7bifO6ntH1ISTQmMK+pDV1qwstnzofaA+2NGa
GoJnpQQTLHxuUhBt1Tib+IeMC2usAyHamaE2ww4EgLB2Jz1yqYxVzuAfNVWX3gvp1pn3bs/z09lm
EWjNDVgX9J47YW9qUuxWtVC/H2gCT+eGUAB5IKYpVDuoC5JFlolXQobrAuA8evLoLzyyIZbztsy9
qI0XYDSQIsZKZLUtpjsnxaT1afOsmHWs1csFbmfGT2Vb+b+FtK4y9jG6h59jcqsCkcaTni2eMETI
arOvl+ED0GbbAi0ctcMOEwLP5lD/YExcHwVdoNwJv2sDlc2ryavAcEG6pqyFNmpByNXo/+yFTtlP
DLNBvYJ1DndrA6stxV+FRD4QifNVQix1zk1mBgGRJksvtNS3V8/1QPOzl7qJMvRo8/MgcEfqB1L2
HbBoFcas2BP9dNCvVNXwjNZXnIi8dqrefc7uO35DA0eR8BPlGCiC5fwukQkmZxmCTuZoqxGL5mGg
yu+sHjwMfhNsgsU697PunPvKDDvQFGfx2WRwSMfuiRGFu0XIh3VH/4yn2Slqwt0dm6hAuj9FEgH6
atF7Z9E7S5s8FxJkQ78coZ5fdigYlAkarPIK1pc3cM/1DtdM377JGWzgdNQ2x50++3Y180ivXpUA
ol5X7rErJTwsudohdb7jAhu2X1NMOs9ifoLdQPum7WldIA81zazsxap37SCC296jKuGFRMYblVRa
8QjCw9UYWGGKQfaifqgKaC4LyS9BB9oI30wkZVF+P+DrSG2Bcsfhv2ww6LczfrLU5im2Zxwxb6UV
kD9/8f8qPWiX+pXZ7dMvh4ey+K3FUuZYQ1eTNBFLu3i548wUu7NRquBLGIZBwHh+UeY0E91s6nvn
vw3XooRZjF2v6zpkuG6xbWXy7OtK4CjmmYRQcK2wSdl49zn4x35ePD567ibHo7Bl/31JPqAFqUB0
KXU51FB4wkUrYe1eYBn3EOcLFXHmn2Cs9vEcdpRUFd8R7ULkaQMoZxv9OolFcC68VWTMpTkAYLNu
l+BcfXolAUqHwp1FhHPQBYdAgnlEtwHhXI0tXrBKiCKTyNtvp6UgZkLcU4yB4mM+2K2I8S5W9bsI
JIqN11SaObVwtodlBPyPzAUY+0CUBZ9FiTTV+YpYrEOxDSJ97R+U1CeFBF7l01icIztYeue6Xxpu
w+cEXWXpw7a3xBhHf5fsmu2Np/TuxyJqmc+qQR+sAK7Tw2hT2yWLKbFfA28LohhoYC+vTPbD3PZ8
fYZ5Dse1s78qmuEf2jd6lHPjIY72Faftx7A1MmNF064cYk9qYvFkwtgjyGqzUemyUgEr3eOBaIXO
jfSOY5csN7PbXlcsNj4bl+aC3CBG0BtCy6N8p/BcmzSXPCIcg1nUOH0eQPh5vXoQLulDe0L25x5g
+WSpdm8PzfHTaS2P/fiAd5rIgETHoeAwNIo9DUfndJ45AZiqF4egjgwtmxjUdf1KoHzEyAMM2DBk
ZB8PMIGNgrajfvgxSoamE1+ywWWV5DZoZcS/q6G+69X9oHFPfeT2ZYvjsoLE4lqwcUpWiL6Mb/rX
M/BXNWRSJ2tebgcV2zignZah3VUBQs8+ZGQILrk0uxpi/SX3CdCNB7xlL0DqRPfOoE/rv2AH/qnH
IuZtF3A7xlGlLlcoj2nh73lyuSpk5D5aWFGJcWVqJ8KDgQoQ4BkqcWncX3nLsikRohse0tvLXfPr
aOhivSGiKeXlpQk+pITkRgKZzN39atXaDEqFZqzqgUqHeEsFC6gWz2KbWpqWlFmIYRl5ZCMNqV9r
TScc9vUV/19eKBHbYhNyhs+9xzZRS/ucoL+ROdl+tsBCeBp2//FHoWf9nT59HVhpdHoRU4xRVebb
3C68c1YMxEAoKm2BU75Wa6mRuN9VsY3WGhn8JEvSscUiOK0qh1HcduZAbgLDwTn0Xu7m2eRgtjwK
TcUsTVhkPAzaR9J6EcYE0eiNaiYIHF1Tx1U7r+hjSx8XXTJKVaezmJejnjVOByPGVMej4O+Wdsjr
9BPpTecv9UwuphANVSVy5QhwoXcTr6RLmgYLYkHCHGOEAmcSgcxmCg08qhQL3FJsYdA+pKxV6dUz
yC7fXXpU3QLLT7BVt9kYGa915qGWY02Pj3ivBmAKQC8sO5rxwWNxav4yHMyt1v/G3UKDz8aIE0gX
DJh9BUh+Qck/h/jZDs28kto9ZOEVEAb9tUiK/rLSh+7vId43NeSI/W/W7yuiAclgs7tiZeVNbOiq
fHMaVN7znPXH3wdrttTjLgLgK0HzcaRj/Cobp4fngyxbOMn3MVSF21OPz/1KRx/mPSdycMU1n13L
UwJo2igBiJsh7M6pR0LhL7Td5Ajlq4G/aKtap8/ABFMH4PCEy9BFRkD5nMpteRK80nueccEq9YQg
j5T+HkwzvIGxNKA1BmPiC4ZK+ON93g8cwfjZy0US96RkUGLa9VlGE1y3XcZkyE+qyMC1rEi7PvKW
K+Ldgr7iC43YvhtnJFNmPjjR9Flx0iFCGiDgnSbyV0vYNnZrluPLpb7tH5nvMKIW6yYLJJBY5lAH
ZPsdwO80ocxBZNHws5iXLufWgZzrTtQ2d0cdF0sS0cXw90PhmdGwRqYCuJjDFpFU8BcTAl++ccKP
W7fAdKIRdpsXVUgBQqSUv18teExUbCKELi+kuKiCYEmoKLL24w7y9lPI1QqFyVwN1QQaXqZyWU+/
pmAR8Aq2PrFSHkvyea45J5LQYUWmD1DYeN+9lfZbSgmnsBUt++DXdoUgSqn7aiTmReYYk1wvS3sc
z7zH5wLQ8XEbg2YZYPP5H5RaYdL7ivqFKmTYAyGghmeeS8KcG0FnTiMRXVsF/2nWG5e2XGWyp3ea
RenmOvNB7l9id5td9+v0Vfbu0ilOtxYu0BtKbaY5fJbWXLcwkigRv0M8PiG4kiYOTMwr/J8S6RYm
gnVKemwjTQeva4zlpOS44Y6IgnETM2/7bsjF4Nf33t1/aBxy2O5C5lAqANq326pfvGDD1liZBnOE
Z79fYwC39GtTFYkxGcrmCPm0vYWSJOq7YPGcrPWEsoKq2PjQkLfYnuT9n4CWkiIa/+UeRSx8afoK
nwqmozDcNyosaTp3mjsdGRNAxtSouBu2pS9OUzuCfQiHzFU8g25kp3FZHHIHG85/iCmynoSxnZk7
Gu/fMuwGXwr35YFWdqwsaY4+FtFXxJsgGzdMMDiQZbPhU//dcYw9wFTFo87I7mqrSblw3tkNqlVQ
sO7cYJ0g58dMfpZXNhwpElLmUR4pBxDMxGjLtLz8ycVy3RYXFTimWiXnF47nOWTZmYg/9uvRlCv+
npAMZ+3Our54ym/GmQTVBJnBwYFYiNv+etArYTB/9pGJ9cRibB8N+cMKTM4BvKjN3Ih1Nl0yAFe5
LH4KMi3zgdpU+nz1Fqtg4dKA4s7enY+O81+yTDeY9DlYWTAA1HF8fWjLySV/J6Vtt3XaStZTAvR2
P36GXzjdsSmz8C5fsl4HV0n7y6DjhMcqYWNWxPbtjES7k3kQIcTXAzX1TWs8odIMV229+RD6tBME
llK6L8Lk84C6e04A5HHTmLm0KcRLdIMf1GgEml9XHERDOHyTbOF2MRKNTjskfwY3SING44OHKYn/
9499S21m4JCo+KsT4vaPPeEJhjO3y6lIs0nNWdiFyRBXwlKLYaJjS+gbMMToC2nfsn9wTQEHG/m/
iZCR0EKpv6CHP4zM6WDViL4rbgmXS3XVvR2Vt5/uu+XvA337KNELOfWwNOl1DE8oEc8sFlsm2pzt
eJ1LQaeeihYZW1mEKmIBGZ0pV8QCGnVPbi0tscN70BYweNyYQte4IdkUSgrQ6HP7LC7nVP8Plql7
iThhBGDgXznH+dHX9eVV7q9B1DtypumP8uYDGAhlSb2gxAHYmdSrQqXqcn393VIv7IQkPFgM5zi6
d2TvX7E2iRdXo9CBkYSnFjPmDX3YOptPZH1f5gDsz8jsNR2UPj1GWIiKUsrPDPurA3Guu4TXLGlj
uec//a6BvzM6IioLuS38IqyBkZWkHx1UqvTr5Ksq6uxBhv99bitgOHOUmPBbcxYzdvO5n3xWFkDA
DFxqJsIOzMr+RasPVcOVHf8ZdtDjrFBx9vbsh8zC0G5H9NPEZdgBTjtO2gOSJjSQnoDfx8NXZL7U
u2dTeiyCmePi38EUCGGds1k6w+slWm78S1omUAxMWFMzs9PoA384qDXJ8WNnSLIxWZZe/t7Wip8g
bkip7GNaD0AU1USe72AMlYYNTUbwcut5b+VQxwN0ptZ8fIYNcfyWV4126nznMPiR2XMYPONElPN6
u2jMhsHucB4dyIamehuZ9Op2rKp9tI62dsLUH2s9Ti4VN6kQ55xlto+MHCtQ2mwyBnkvouKtgIUg
6HKVcss1n1DNtKMWLV7jBNcKgTdSCXInxzzCXVDz62bzqezTPDvjBcnZCmke/jxRJz6CfpDVbZB6
GHR61uYmJtx5lmaag/2TWVEbJd1egBncTtiWZbwKXYNLV56BdcfWopNVgapYQ26laI7LhJxSoMFg
ddjtpiIlNCWxH0Me0L98FeR2sRDoHn127EIxC+T+aJlItUL2Rgjm6kcmD4EDE3qG+rLIw3kLAwth
okWuQ7MXTo3gSSutGPNHRzh0TWra13KYhBWfwEB/ch9pKm+w0dYHRr8dW6Hhfl8X46oZiu4fl3wb
hQOoTVfHeIFexEzbJni1thG75o2ejjTfWRp60VHTciYcrUkkdGs0RqlSn97LNN7WoESjuprutUmc
wecwlPqYMAyekhan8qWNCGcvl6F9F9P1fe5XrKEjkJZJCusAwC3P3KaxVDit9Eva159D3Gc3udp7
FmZFGb9ILVSNJbNhZ87xAKlag3SRCT2xtdl/ZnsRZAiB15J1Emen8/mmjCyMC7IBEEIa+BIJ39jp
DX7B2hdLKmkxsfbwcJrl0pTN/BzQUkJ/qmGvQvKpjUZYcVdgCzuEix7RJdeY8RcZ5lgfuedcEQQP
9KpRyxA1MzAGx+7T/d4EAKVuB4baoZ191e0wk+VPeBkU+IUUN4mKNJhaQzBeug1DzckU0Yg+KOAU
u7G4owW4+0S3DuK7sGveTpmmcU3n7stbNwdwHbM98mMdQG58S/eLTRRohFltEZX8N07yOUm1jZKz
QVLKtUBg4IFdKm5+3STw9kIY4gKaiCbnhiHK2UH0QD7vL3CYqkM0EuDA/R6J2CkR4xZZ4gAoTRiO
EdJZ0p1/zKKc0jB8k3OYonDJLWRN/n1m7Tdks+v9WCvs6sxix1gVqTCJDndlh0b25l6vAkRMO2vy
xovJUt+lgA3d+F4xaP7YpfhrNt83Bh8yxX2NNiuKCIhUZpklVw1ATy96UUX2a8mDgHCgclFK4qwh
yOLthvZR59arswAxQ+b1Zh+THWsPzVeZt9GmKHYV3Ib9+T2rBYauh1HDVWxn3MHjFv2kbzIAxMxA
DRpcPoNebTAWjqRFJM2J6u/hPSa/ltZRN8g841x55iUm/b9x9vs8qmqiDeCmIiC0Jnn0KJrP62Cu
Qb41nglmiOjaTOKhNxGhpihb7EXPhEOYvOsGCkOoNH/1SrmvacSe69HVNrqukoUtuLladU5FW+gs
18Prg6N2nBGf9YOSpeN/LL2D7NYkKhCcAohjWXn18vXKg4FoFgXBzhmxj+vA2XjuFF32MapH8it/
zEhvV3LQbzYHXuYTxblcpt/ht8jJqvc5wUnXfFnk6dIjF2bEc080ZvNx+XRWtay/7fb0lFM6cKgJ
KEzhELVpBPELcsVlHYKRX4rUTIeuOy/WG9A28kWS0z2Dq3qNzJT9Vu7bSCpPagm0JKNB4BXZaSnX
b4nGpSBRolu28Al4p/wopke2UpL/j3XrGax9jVx7UyswZTVCmw6CPQWPAE9plvPYnYabBbIFyWKY
FdkxGaJld6EWzwRTo/y2P8f6YfqF7+g544e2SGgFTdC1oRCH6WAVanbdiyti92Gkl06Va1DAvtOx
IT6AOd3hsg9FotevRwLbiaHFnbcPrrTYLIDfnPDyBFrWVmaNMmQRtJQi8e4NEvC4J2y/Mweq8mDR
XZeDFQyqK+PXiTO+I0ZdCneOsm752MRxTN1x/QlITQal4o9MS+Zl42GDxjgQxKg/QVjG1e6rghlx
NPnnUud2uUpFY2BywVGWOq+yfpbNRPbcgKBEJwwNALcBKonETk2ZrkN/XUqCms49UvBUKQfAWK9c
/uU+DOhz7p9RWORYoqSDmbCckBK1cKCUR/DZeygOwnDPD6OiPwW4YJvqE0KaZH6SzOdUkW4sbwSB
tDz7RDqEJc06dnoARE7qG1YMvZMbsBBNm7OhSFN5YrelggvRc7JIjl++M6dq+ImA7Kv2swxgaRBN
H3/WnyhB6zog+hQmD3b6AE+JlOkRuM8seNbyUv/0otWHj4Yj30WzYVNaBY/A0sYsn+lpfLHaQ7Bq
dAFk+BabetrzanVeAzTmKtiVy+ayuEcirrqSwR0Q/kSvRpwWWluOYCyTBapPCfVAHrBK4BREZJpb
r75DpGXNhkqgHVQqPNICVBwWOQPFAahemllGZ0ueJ0mtWrJSY6ucaUIzhWsoUTzygA4F9+OA+VGH
A5fwS11vAXoB2YoteCyR4MlWYkK6jRVlONbnXpQiKRZUf4HiNC1QF3k+VNGQr1lsz+B+S/DYrdug
xPb2PxVDVxn80875U1+YhJAjaJGuTnvPw46v+lqeR4yGFkXZ9ZzWJIjcZKD5JmAlu/iT5qnNlTl2
1ejnAnUA5zvjq47D515EQhL0fIjzptwJlgYupY66p78Wb/BKEkJs6Bic0Q9qdi5bWJ9O86878jk5
P+Gld7pPe/XibtFA0jJWlIP7Skp8eniiAlvOeoBHvAzcMJV9dj3Vr6295toZadkVoP+seeFiLMsI
Oyg9Qxq8xvAWjIAmdayD32UHBq2v7lcwLPvdGMO9D2WOCgqPaz6DPmPcyqXTWOgNEMEMcv9u5iUC
4IeCfsjVhwbka07I01LdEqyOz4dbj3T8ARChabA105UfK+8xpHSyswP5iqWwl/LsGcs4GLNmCNuu
eVXO/6ZLuArp7wmKz5RPe0EFKdEXUUzONkkTbALMsW8nGrM8mmeA5J34YhQV5HfGIa0wQCXFu0Jt
UY2Q4Z1uaFNsm3imRYBOf9JVBoIBKJ3XoPcAub+pyQxWUDi+ghjVCfyyYU84Xh9KCXkO0iEfh524
8WuWNyPBOPKkWYALYnUS9JjKuLz9IOsFWi86tQokzPHsPA6X3nAlNo1N7B5uF6F4YeC8O/cMQ+M/
sKR+4JmyAKQvupwlLLOp4YddY8PddwzpoCzpycbxHOek36c73r+T9FVToCMf0eZ0GiFb2ePc4S7n
7LR04XfphbDg5CsSfOtn+Ng5MUP+d8xF6TjnoVVn+J9zfQhBfbP96rVkFTDJ+zZ5q8vTiFJuD6pm
W4DzySqTK2LybkQPgrQM+g6vUVXiq/tCZ6s4BVdfrHCE4kt7+/WSFKf6w2xOvGy+E4KSWgOTs1y0
V8Qq5Hv/GvRYOYr/cAAo0wH/Bn0loY9KPW1kD0NC+IvpOF5DMS/e3xaUrNjMzU1CClFhhsEdvFrg
oOEDblfabln9YT5sVmyxqMFjN7VUNh3NHORjdTD5wEexR+tn1gvSaBXqBoOjHj6z3+vjI6+xx246
1LJtXjzjAq7SWQPK6sfo2SoXO0mZgIG6m8RZF0shgkmig08Cv/YqCUnhAaBfSJr1282s8QPSIEWg
zNPOFWxgrAV2UWJi1aPJ1rFYauBguYXkGBeIOlek5bqMLTVoYjAy2KpSGGcdd5KAsPJFgp2ILRAn
ZQlFX1ZARu7qHa3dzObE3d5ZbO40TCdqqVxu3Vkl0egQI3aYM+X4QZOvL7aFvnxRHCr7Pxdc2ity
ZCLZ/2vIwGEsHh8OZug+ohA3O1Bav3Vd9pgHwUz4r+qa81jtflDkoSxe1gcAkjoqLFNFkLZx2z0x
NNALGWlEh9SztuYkExsxIgrUcqgrbJfyMDdq8l3w/M/1PWZFxXE22DI/NgAZyfuqwwqtIRqyrc8x
NsDFdF1UlEiM0SBTdn6apdxhWCw6Ct7T/cQ9Kz8JOuDCKGYQUtc/QYxY9vQmFQxCRiPBn3ufBx/B
L/9sVdJrzdQWje6DbV1aVJI16lFnmxfZSTPrqb+GM0FtNybGHDstTa0f9Bzu8TgFB+WL6W7Vh1+T
Zfvl6wNNz7PcXAs8hmQZ84/0og9BWkYKeBzcQMZojZOyHiDqsk5M8g+Y5BRHIMqJguDC1KGCWsyf
rLLGZSF8SARFxU0rPz47330ig875Bpqz5qVwI0dL+pCRXWD4N4I4KXIImu8iQtjXYsCvvNhL5Cjt
O3ixDxcl2OfVfslmsmhy30w78FZSxcLO+DVdEk+ugEt2dRA6PpRjIncAnO6n27BsRtYdKes1uUlD
D9hFe5RqBMveJjJt6OawD4jU1+93dy/74nIPvqb8HPXLfSmSE1Cyw0TESERlAmN2w6qt3WpINEFc
eXkB85T123nnf21uKaOVFAyI8hA/FYQd25GE18oHFivjcBvymQKS4Qdonwm5xcMbhPPImIb2iXKv
FW710/oRfIq3ghP10apl5B7tZaOHUuqzCoHM3HBPAn2zCgE713jr9DK3pzVQOe10+9h7/rkcd2Qa
RGo+DXvkeycdgwZKPbMcfV7WCqZEs/YyXGP4TiS2L4y/ZFLOWW5mT/zWsAo+2nP5qDuXqROxF5Yl
gDc6375obWbRC+XfSNxTvFuaIJVjhxASUy6vMw2kd+qmSNSIc5aGFaYX3vn0Huqso16kkka/C4mK
OJV9wn+0xqkq48zi11teGoQVs2gfM5TI2sh5iGYfYVE1kv2LlqzVli/wKucbDqPdTSW++CO+U8vR
6j9tyDl9vZT5nK0hG7e6zn+XuWDW5nDCWT1LZ5wkns7BP6Amj7Nhoater0JtL75c36UY33t2lfsD
nX8JhO0xS/2qsB3paoqAjzQSgRzYLVbjrG5cVtzb1y7KXjCzNGlYZH/TxoAJYbMFKw1Qum9NFrx3
HcCi2DgeZSzbtopAcVn09WcZ4bu0I+VUqQpfnhUkrUWhbF2+TIDZY+H91+8Fd01N/m2yOp2LKsmP
u1XITx0yewIMId0rQPzAU+0j7uSuZNnU906uGA5c7fR684PR5hLr37CDeRTBfI5DwyVZNhhzHCtE
hzo5MdmDBbG75wrfiBezlqb26ofGtatutKLSdgdUOufgxpgXDsfO7OlnG2JHtEnRYDWUKmvZpbtc
vad2421CNy7eYLFIB/UG4kKsQHV462LxpQcte9iIrKwxwmn/BoquD9O8B/FEkyz/KoTJROLfmgAm
zbBbfxkmO/OcM+4oFVimrG2QKQALKrvJbI+J/bB5l5ybBHAX9vSl0wUO6GmCq4H3mLfpIEbCAOAe
wdexbSRmdQ/3VaJOsxyny0PoKlncvd7z/1z0J+GPKXJORbP7md4WkPQX3Yhs+ttfdEGGShmWLz8T
mwFOo9AOwUjMQNcQa8MoKxcjljK37SMgL6/nw79vSL/5bMstMRvBkCtYKLZVetMaRaRLcwBrbdzI
9bqiVnBePFp9OGIXR0+h484Ua3uG6MXCwNvtUDHngC/lhivkNQx7Ah6PjNXXcIEOluqaAGIX3BBq
yT8wLAX7Fx+ghBGtOFkY6SYoLUol1wO/2HOsJ7Ztjwkqxrhe6sH2B/aTHtLvS3yxSi7WARK/LmbD
ISZEhqdQHfBeOv0Q9iozAaNcPN2OWHDhhhozh+aTWDRAb6+ogqRfG0J2BlvhAXIXWFn4tLHvFkNb
Q7vAmrFMASjM1ddJEdQ1SDVA3R/Q6Wo7neaCY8B8pUDmWtxBrGSIomlrovuCQxGYHnwyZCMYmRwK
Q7qxPlZx/Z5vubyn5bhjEWh4o71wOlICH0ZeCy5EhyIMURFInh44z3aDON5NOx5v91KOjdxvmY4F
e/CGuiXEWL1qP9qqfLMv19vcLCTO9m/KC1Tvjt2hOAPb/eJqcMPt4B5klBkrFKGnytPgWY6rXjAv
h0bix2r7H6sqBR/b+EotrGhxTtpCf7/WKfYwn8UhIJDZ5Zv/yEbsjsAYlDB4ztuULtR9Cikj2B6b
b4yauFO0thL1vTlZhi7jtXC20lcAxMawA5TDkv9NPBuipwSJNt4PTge/upWBZWEUW7r1EJDAy+aR
PkftIhswPrs3QhTMvzfZcCpj6OS7ETEyKkgafEK9oGbrTdmRetLYteGk+QkploRfpLcyPkyXNO+p
6HxJZUTCh398Q6t1hApMX/BCs2d6WXFRUb+uPj3WS5urL1dB0jdsQ4SW0c2aKxSRbGqXOLr6rP8g
As4zfJHXToQ+ktyxYDUWERvrZVsfy2tXMofFgLVgLKTmOQd3Id0GNYt8kHRUamslqWaNil9IoIG0
zmOB1B0dPL8SpJQ4cccbY16w/TbcWGfFjYmOhXT/GqFg6VXGGNdDFo/SAzEA/D0O6AsIJvhqZ4Xi
5glZzP70U3AQUQHvCw0+7gVgjGcMtowpJc8CimABEgQ5l8r2G6dhdIfmMS33RwVWYMmzxU0ms3eO
FGQRkSGnINy50Ehv4oeP+Xuv6DatO+wOA1M/+4+rS4W7kzk5uWTvuwcQ72V9/HOODQLvGEpg+GQZ
TXmZ20gMaG4gEG5HSb61iAv15twtzB3F4F7lTYx2mNJnBKz55ROWII3TvSBccHCPuAUPYjCdvYeo
OlXdJ/pO5DIxrqMD5IBcFiuCP4wYwYOv4XKSI8fgWlWeMYc1nsWzrK9lVSzGPyS+C6aud1ud+tQK
RE38x720wsuWJP2fy4dnzToUthBxXLTgWg/Ac2c6TDBsw5mFNIegMZQ1HkHA0GuZmsnSeh16rBIe
8m6Tg1HWLnZhlmrUcWivG/cAyR0XuKiITrif6p+hvax4P22uGyH2ZGJYshLArAPFAJ/pv6w5N8/b
Jw5lXCNA9L6EhoUPsX+OxI0pe6i0G7C2D8OcAWz8jAgQc/ryzD3/ojsMvEbN4nBSd96kAY9rxmzX
GZxNmNembSJhcJPJIvw+RMrUsVlucmavl7ZTT0xhyw3R/9tSKbSwjiQTPig8yJRSDlud2c6JszSv
ka4Hfe0xvi6JFTOPDRoTr5b0AyLtrVuRr5Wvucqa6/uAVRoGccP7oYJHt+HtXm+yuIeqguP2ZHoA
ypnDTTeQPVqhe3m5pKqDnNyzWPTxBWteObKbpkEyqY+bofsUBSE25n2BD2S1EuIx+CiokacBP6gh
32CD+1TeNi/glc/TD5/hPXH/MsL85gd3yRv6ayoJiKhC+Nb1xAiz0+odGe5k6TVR7ZyfwOmlw+B6
ZaK+Lsc4qNJq0mmpgl/0R/o7iybFnaN6nIAszpLqqcqzTwKO4s6mCN2BVBKq6J3Gp8nNEh/z5AGE
NrnY/+KZJPhLJq3zQxdVtP7CZKlmNeYrtLh4pJw2s1yvEgJ1LgEjY6g4L9buJDZAsOCpnwt21s2Q
AkgE/LJKRZU69J3scONomzT7jbRWv+8Nbm1ptFkwwGcuvEyY+OXXJNtN9T2bkFBCoK9g1W1fuh6k
SBNrCL1fBHeM5UUs3nY7CR+0ezNiJJ4gNOq1/PSGPSa8P4EAZazJRbJG3eGVTlwWvCk4V8jqr0EF
Lh/aTZnNNaLhS37B6KVmxwm5YPsIHUoM2F0f5irYGQijnv91rVjpkqMoNd8otsT5J6AS5hVzSyvs
1Mmyfq4Wvs3hH68cjVcv3xxMCPrRNWnT4SuazUr+uxcNVbWKeJ9NNdFeuoA3WVyYQCzyNrFvJSWK
BfeatxVaBVKp48MdfS4ApwMOri7QPHhV0s/oOj3Yebhe9VZd1GS25zpOe2naU7/5Een2ElDg+UH2
rPxr4afXxYC7WTzIHqaVfF9xPZln/ob4BRG5jB0R0Sci8G/0w+tJ+eH77+ZNgjrUz5jVEZCmiXzj
0wsH4n1Z2ixgxg/tvKNmYOTfcU29UdkrWG/iqGzsB8nHLmEZHLmRBknCHvbiZFGdTy1GdwXQyXnz
Ur7TBL2gSiT3mcewUGszA1XajPNPpAoKo7xSIYrhJZYUM4DzVLz7NXGEB0nOoDDstQ5fB4j4r32e
U+WzlqRCZUKlQQruR93gaqivkyWvetSSwHGY/0gG5cAkMu/W6EiD+02doSL+ObhC7vj1VOra8FVZ
rFRAqlBYFy4JDakPzRo8KqF5/WZSNoUhw7l4rKxLUZsnKwUncwKib5uWQurvOiqEWJfwY6U4PWhG
IWYbn7AcqymFlNM6CKrWWZ0LAZxcuEug3MekSFLgppfVUvOhy71knATrlDHYJAJ9vbvf8yZ8MZ/o
bdDhNNvhnxVWMQWjxoGmNyh7qZFltX8tz84fmyGCgDuk6B3RfiRDQw6jsOuizXMmUO+rSax9szZX
DcxcJ4TgU2M9iRgcfKicDZmbu6aPypN54m9uRq1VO6weS3AhFUa4vXevljs+74a4wx/T7IfTpRor
eGNLH5oK9Vk0JByWWmckGxPhysXdhuYTtpX0gzZcp0o4HOG4i462KNQGoDeNM+BlchpTteiwdf/3
DRTh9gzf9WoHlR8AvU34GIbYuyTaTK7IhReBbmLfcVRiK4wb5IcsbNe9UbM9H+ZJvh3ywUhJMejf
EUGHYENV6iDpf52xEyOCj7yHWTqChKn7MPz+ffTJ2Q69lGk1hoKbJaMCAoeFrN7FcyTp/b8ps2aw
DkBxZ+FME6lBLsg6ilNEwt9YpD3Fi6dTSUEcagiXd6+h32maq8SgP5j2/wLE4JhCs8ytNzmVFh/V
A5f4Ivs6vTtLcXcEbgt7BlXRjHM2TDE5sYyePhEKAinad6sLDZvZ2iTXtdpMLts70mVI0w4jOJ98
EQfqIbtg1sh/1847R06l268UjyhbbSueBnwUvs71ag2TYbnH1AzwA7hMMzAno0Jt24NMG20hTrWo
WrEgN2FUEq+kWS0oRYYzkPWH+1IsXATfUhOngd3q54BmUjG1dOYA8o6fQoqba9Ssbm/DfEUE+rFS
qHMnxdgHhfzfVWRk1ratUfx7+WPQExJnP82PoQY9vspjb9M4LzxQIYLqyNF9hoWeUv8+q2pH7Vm3
nH2W4Fhj2G16VUvjpmrEKTYwOkAU8BigmiaToNdXGLm6mEyt+CcTDrJLE759Wzm6ZjAjN9R4mqS5
KZlC7LzlaUZNg61+Poxv+9IqwZQ5d9hE2trMi7zG+FGIPD8otfG14XfNx1ZnjsIic17Xardesrqd
1B9GZ43y3KooIAqeca2uPNjmSuOVkKBSdLavAUWBVIn9LBnis0Ic4wCpisau+gIixw3d0pePIM/n
r3z6jSJzouv7OCZUgMvZfhcX9Yrm6T++kAZalUWuSKXyApXUz9gvH/OIjPJjYzD1i6tmDGnBN6dU
VDiCQWb/4NG72TooACSD+lzmOd1BtqMgFi1h+wmBftL/z6643yzjZThI0TppKRTXUiiCECtNMe/w
Diz1ebZ1nf+W1j2ESfQ3scsF1dh2aIL1+kRHXWQNv18GuIMhoUGhqX28hyxw/J5Wpgps8h0KsNZN
Pd9ZfKXBltiCpbLqmf6ozBHis0vFcV5L17fi3W7q+4n0cxXeJftSkQKMN9wGMM/Vhx90ampPCQ+G
Q/BmW+KFywqaAJ5k1l0Z+giudbROGzk5CR4EGuDPkdzdqQhNORnqWBVOPFUoIxRo5VXeq4fC7S4X
CI1QYKeGZMsOKRjD0sBx7mjrAauWvuDWg+ZEd8w3ASCRB04wstAVnvw7JOXKnc/0VV/vzbOmhAsB
kkaU2Le8PE9iR3gq3HhkjYi2fAMCJxdQFxkrBQcNGxMzxDqsB2tVdNuCWcrZnc3ZcgaNm3/bavvU
cxRJdVv2ukCssWbXD5997eTsya9OgZR42ph6nSM2KUCJeN4ow3JVk+7KtbwQ+4gsc2un1C0e+0Ro
4XC89od5G0vNbi/F06BZhhJ0f1jKZh8ajUD6ZTJUZWci9CNPN9ESKr9Ssmf03vllDLT2tAMQEx3m
d3dGX895VGGgeXK85pP5xL7/2iQ1xb4x4yY+pVhZe0zzCh0H/sZmBhkfXZlsZFSVQ4J65cfQEEcM
wUqOj7b1JEaWrreavoCxrcQgRoOaE69Bqo9U2AsaLnXtUVX6v7TTN4N7nKRcFq2ECj4KwUb9flcN
oFhdnq3Tqqg1LIu2589jUdWMTPplfb2f5OGT0JpPDVQQt3SWOEsYN/qoFd908Z8P2LdGdYh/hADv
9RV6UZ6lO8RUuhAiEDMLRW8/pXNCFQaE6Jm+ql4k2Mrjree3Mz65fp1oW9ylw/zFbkgb+l7FY8Zi
TL+QiVEnwV4pk1W8pjWmbDKuB5tmtjxeCEBgfeM/yyxzI4GKyMw/+Zdf/diCgqB3NqgfC93CZTmA
7ujp1HHPMcyD8tVlj7JfuOJ3jCr6KyHpJ7DbPo6jIpWoO0bpo+HSUsH38IcM7/b00b9XGGkWXfOC
KR7alx/ZuRlaMY0Z807+psVCAE5XkDNA86UG7vgt71poTL5z+NV7x8nh3a1yRQKRPKeQMrvfnPo6
z5UcqerN5meHlNpdyvjh5tqLv8g//fuFSL11j3AeZVSk/PbyAtQj9dJtTWGWYb90dyhrrnMtacR4
6hT6Bf0uMMPjIJVIuE5J0gsROPf/PdcE6K5bvMu1Oj8JEr9kjUk3K2IFjohfHm8qCaIePOPSW2nk
HGsQFgdPko0xbaANr/qwlvO5DPvZu3EGQdzDpTa92tiHsu+P6jkJCFCsLloAoDqIC7j2unDfuvNS
qYyXgJyPdaP5zwQDOoiZSTLdOJyAaZAWSsSUN1uzG257Spb7GPJkYKqLD2WY/eC1pbIlakCwGav/
9GML4pL6ezLS43DYwi23omQckImxdz+1TNohhg298svW9OMPtPJZry/4rLK8jqEUIxnHU1BPf2Wn
4sPNvBRuJS8H+Ds7KVMHisFcMqn5h7sPO+yz+8Fe+vNytuFoxFO61jExI0x0KvIAVjIXSmVjvnm+
W9DISAqc4UXn8vA0aJgQh/60xjnWAnj09pqPe8/m3OpySFXmdJXAK6nFGDdhx+rzIAqi9jY7kJJu
jCWi79FULbJxopJd2EYeC+r9ggzLcZTPD2zqaNSbyz/FieL1R7V1r2Z8NkZQkBnBQUiTDKIe2qzs
IkjGOsbrsErGc2ce3ERAJmGS914vWxUTMHwsWWVy8kcOGg/dhp5gqpxmKcD2xYdqcUjBTyQ5r5RE
kz12HV0iGbynxJZHgsVqHdn71X4dGnoZmsfhmmj+zDbGDCsi3/08lBtGxmKp2llJDnYFrmAp5kWc
EonM4eekYs5Rl0B5gxzuzT8oI3tiOja/vLrpmI8UM+Ea358MuXFzAGGgZDihhpCbKQ5EM94QVM0u
dIaKGuv7+06YsuG92zSvH2MJ7SvvJ/K90tPfpCLiW7M5CjP9ObCodWKmKcbGouua35bCKnZGWCZU
+pkHmGmZcWYeezwEDl5CJrK4cpSn90dz9DoIrDDkJ1yLJp7N8EX93FLVR2jVcSKsk7NroEaAlgwO
Z14R9VE1OWztPB68hvxg0jccsJ4wkAvcPCaSfvQzpGhFtGE/P1HFHbGjfolEDw7Bc6ZXkfwLHGh7
IA6ZPzCpL+U16sO5/I/GYUGOPqQ95xw97ObGpIDGFkv9y69KNZtguZ+UmHScvIVNbTvz9r14/ix6
Hc1Sjv4Zo4hppPOUUiDeZvv9CSNUMuZV6Hs5Zg/IJIRoeteHGUoChmdpCssoSjNGnYYP6qZWThX7
QekOwCIFe108RLVlTlZMb6pmgjqMPJNHmPD9JXV69ZAO3uNfHfS6hS4SvrUYNkp0jTcz6LGE8RgF
iQCrPAZ2bDGx8gCo0vmxlUkqYtKrAL0AlFMP+evL59yo3VQAv5ivoy7TI9Z2Uqm+kRYWEfeFtPIR
bO/mmTNexmqnHHJZeye/a79tR9jUdu7Sz2QrBGeOhyQmp7lggwJbO40FRUxRHz542GXoZLV84Dx8
3tGk7TkaysTNJVTfq/V37KEdk1YN2ZLDspI1ADBQLm8F5kHHxA/26bSRSLoPbmadaWd4Eaf2FNlf
micLdTuAQpisYz0Sx/kDdbWMQNh1NBpuCUokf9JP+tomAKpPUKUU0RyLcImZCmH6u3cwwBmkSfnP
FfKcULXXz29WESfoAI+tiW36KpwMpvK4fEdcfhfG6L77w5s0xf6pWd7wqGVvXLqEmzxNbYNs8d5V
VGveTpfVRw1hTloly2wdSKgzqkghw9VfsCu6HptL0FAW9IEkkJKy4MQ2CRQVHeaIixQFo86ng/Br
ma6e8fNfM7kEhnMkFOBbQy3CYOVmFPGWHnraKOM0/7/aTFTnYve3pGeLmOKouIHQkxQ9qLGD5G2U
oTuF6/jLTt6oC1qO1QlXLZc6Zp1dTXOhG3rswOKnW5Ghos6eOO892wFMXcNN3A9XZxLtxrkcqLth
pT0WuOQzb0DK+EtIFw7r/lt2CqCQFPkUYm7SvGG9pv5PT4FckLRohNkrS1/KlsMVz6S/2foH1u/g
uIMEZ7r3TE3xtfj55s500NNZlPuar03lFjsjIzfiFfr/w4GTnfeDYHt+Au7G01iXHclpNQ8nhWLA
MOBJMIXubbRS/8fhTx+rNnE9S8Xg1+kMdegYlsEq3fuYPIAJ+3Plo7fIan/DI+XBO5DqVmd3VfZy
HuPtxu39T9fRwpe/m0OskQwJi9K/CWoUGGPv8+xPKBYLAy1D5WhAbkxVFijSd8bSKO9uLTH/KESl
m0cKtWnsAvuQ99/i9oHE2cFIYLkRn4J2h2TINRhKcpX21aM+kLPCVZhVl98UiVO3sl6we02oKyuj
qYDwLv6KUxjYhkLkId7PNTKM3M/gHqVTb66rv5KCZK36I/SwTM48Q8EQwBBONOqXL07zkDhbJ8OX
A6drr6Fw3XvVv+tVO5DgGv1xj8//oA5teMnW4JMNn9VpjtJXHgNbw4ui8PvNwP6jX4wMK05aceXu
X5GlX68OuB2uQp46G1YcNCJksOAstBVYLW+UzOrwFiVkW1Sdp+stwWQs0OzWNqbtlPSCtZe33T4/
Y6kOjBnHDilskpUQ4VS/0Vz7rngz+QgHgXG6/YaR/xIdOGXFWNdAPhPQcsf5/uayu8jGKpq9yFvH
TsLaXQEpTopq00tbCEhR2gixkurrgGMoNf4m8vZC6ltCPK6BhQl+C+ePum3QvePHCEmt5N1vfbH4
taJ9MQopKluTjmfHD2XQNgGyJ531CtXywh5K2KpOg3sQiZo2FX3nWd9xeVsZ75L0TU8sKymKTPEg
4TCfCf90QhjLOVbshLJa7qOZTC7t8AxwmC4mnkZkMKJCYzFjpNvxHKmDlvARPfFW9ujDzXWBEbdw
ot2ukPyyuEk/3k1v17vWHuqdqXRwBLbSDbnJIa9n1Lfv2hSGUkJ1haJtxUWZjaJHwpsw7veCxVCs
/+g7bRmaCnp0lBBJoctH/mKodVeREEZH8o0oKTqJq9AuHshEBOTkd1RcX52HNAlK+16d0q63KfH0
p+ZQX6z9ih6zQEKcSrXlK4ve5/QmFV6fj+WthxZfnmXq1SZ+KcZAHkyGa5+JwwtfE40hq92gEaQc
TnBkN8y1BJBw2GLmHsYtKyAIfebVZ8C8AVNflkCKjvPSY6LxtdAl0dzG1yYS9aj5Pesn2Ll1dPbZ
8fOOYXYNleXApKqmqm+dIjptfFz7yhzZBgupRpEhl7FoFW+ufYwWp1mzra1/rvlijjL8QX/RkoMU
OpOliK5p5srCHK77LdVzlkwvQEQXoziwzjOi8wtY4U3sjL+87RfatGzuf2hWcrf7meMwwlEEVpjz
aO2NSrA+WZOBssXcSDj/L38Um3G6NEGGc77kWgXL47TDiQ0Ke8SkBd6VRwtxOPmfd7M3vkKbT0Ia
0MjbpbQhhy5AO4wwWM6cVSyOTQTVHK19hxg/C+Q464lHjutpTeiNyPGJPdxe/f22hr9KUKANWaEN
pfXDJPF+n06KXf7e5bbvCKLVBiehgf9WhBg5svnAKzCqCzhFbwmDXCt6UiXAWnHJC86FSaFt8yBu
7I1KkysdBmg+TMWi+HECN+44+G7T+92rj1nBr/JWEpt79ZU1B994UssfksLC0i24ikcFjxXbAyvP
7QdDh8yfsn39aEYsNiGvquCJC5NZlmFyxV7q++0PWyV6BZUq8VUJiUjeDhRw5zi7MuErjeWX5z56
ZA0jKiSoXQYDcEiBvPUfTDUggHw0upsRypO1c8XweARlx5zMBKuUqSdiBPByc2Z3125/x44qOJX3
/ELj+Szw6y2Qbbqy1muJSTS7lmaLQl+KFXgn7WwhnuWz0ZdRjCV7VIJ3MSQUkaMjc6vm1xeG0WZ6
XFJxTY4Mj3rxREOQZeOE95Eknhqez1ce/ZUaPe420SvHSMXuHsWSwe8nugFLths8hZtKiiaQ/1V7
jKqvAXiv/kVfcTcv+YJSVjliu/QgPzvTia++jtBZJFqAQ/rj2/QB0NX3eSRobA4iN8xE8VN+ac1G
SqQda8xVhitITjXO7j1Wv7bEVOr6u8XvsWu7YGZpze8Piqwuw+EEESvU8zGqz7TIie4vUyWGkP3s
nLxLXuKQCCM4GaWAtQtZ6UV9gONWHD9KJEjC+eUX4nZHCrDPjAeLnfbbhnh/ccMqJwav0aj/+JVn
C3UgrPhBeHPlLB0cCw0sSE/CW3Tib7iYQq8ZVIB/bJ+S6tm0/8Rn56S1Qr0zsIUAlAlPV8yPJ3BN
D9gq2Jsn4f0yn6un+0sLgj+0D69UDbP9O+89MdOEbTHWQoXgRK4E56RmzrN/Iegfzt6D8fYiM4Zl
Nq+6KgMjgOKVLHEvitj2A+d7Js5oaKDGZO8srkv13+J6lGQ8dYUBM8wT0aEuBtTOrusyoBdo8aOS
ftpn38MjasKTEmpWGojy8ql5JpBlzXthFwBT+tiM1JtDa4LLixPomqBuYOmhWwzYaMypwn6D6fRL
VV6IHd79hYOGR+pXxPaVfLjtFPrYHIzAHzUoNG/z0piFewA1SnsUZI9m5+I9mZe4SzMZpky8NgiK
X/2up5YXPLf/OneBd+22nrcpyYm1R410j2yPwkEnC9Uw4KudlIyVCHF9OP2Zxw6QsU09Zm6UxgoU
MJvYoMy0mQOx6dzMt8vcOVCMx6EWizx7mqF7JvKr57AkSZ2DsBiJs67gh34RgJkAVRTppIH9JWiL
Z4VRyKU5m6yqlgAI6yx/Uh7P40i1sUny8T8WoJEgTugpiG6mjHietsMdfd7rPI/tbM/17xNIT+/6
sGi9/GAv5KudeRVcNdDgdsHnC0vT9RqvRHZJyaNRiz05jLjfSleHYsTUCLkNRa5E9Q5MLLKOsi5j
qMQ0OaegvJJxlQyOZNtLvf+koJRBeqJ89v4M4GdfeFYLwSMXtBBt8Rin59pD72nQSwa01sAJrYfx
MVu4SZOthacIXMlFVaLh5mywFzpWvGj0Ybup8zXi3DNUWHWHrZ75A8q01qUYvgLGnTVq+TtZ9dUF
DPaFa3OhufVi3HIT45Y3Z+mkWTDvuu2/90wvCErGOgdzIYgabLptHOtGloChnuGk9XWGHz+5fRDJ
g8R4C7HAjoxfQ48Sw1IBuX/ZdXwF4W3Xugbc3bt9+Fy+njojNCaLe0wl6kvOdbjAsq/Pgk3Fa72b
MqJT3LNVYqv9wOey7NqUm0MFI3KEKlh6DwMpzKtmeOmJnWHHvH6eX3XRMsoIQFt7tD+XKv4wCggM
OmRtdPnDv60pdhhE5dxdDDJcEQysTqaFGtauL8MjT7NAOE0AYeWSVyNqmp/+s2702YG30wkQh1pG
Tmkr2F7HpITeFHTAFTL2kNTZ+IQlCXcOeOrKgCW3POB3FNlhJcVHnl29vk5tbB59Hiv+1fTov2KY
ZxtkK5p56Es5Krkm0uLdEHN9XW8sgvZ5CbeHu1ZebWXI/zLTXGlbsw2qjH4D8eJwcUP+zWG0xEXm
V8Rtz607qs+ISu6I4nrZDAwa4AWikCBtAg/AKwIByMC16mTsh2i2YPIs1LRV5EC7yxLBx5GjSFVd
IgLJdTgsiARuZ1HBrOSq4EVB0FsXO8ZJi961S7nNsVMkASvkNqYlv9Ndfs9QmGvE3o0KE+iArn+l
ZFrl0ZgnUI/8py2NV+SuyWTxLXl8Lw28YKn6Ta9anLLfZHxmzEqcrBLc9EgA+KljYNfKTEBJNwsW
23XDi3MwcSVCTfAzVMXb/fSRGFuRdJCASGylCHMMUShLMi1Vkg6qH6SoBLYZSJdhFpkOCaiDXhJ0
Sc4584Jz6GpTkzwQSUz6SaONFQB2SjlA8ToApJ4XmYrZnPsnhnskzv0vDzN4i4joQJbOHEa+2Cnz
7ELTiFo2t+hK8vHhjD/aQ2QqofaY6Z3KeY34qdNG1Cy/DgyVh48kZI+Eu1s6AleBn39f8tS9oaKF
7NVqlwJwOMlHF9Ziafzkg9jMBAtoriuKza85TGHr23UVOD5JWiI0SVDfK7lryyGxTViLbBniTEOE
a4uVfUQ++r2BmToE6r34HXxK1IoIksdu/OOhBvpMK7Y1jt16sgiLZ2oRCSF9B9sOOUHt0Y40iq9W
B60jvQfYBai7r00Gqv7Qk7zO1+wAW7GdKDqucZXDpREODuh9RonpoXO8xcsj/Q5bV2as2LpxS/YQ
nmalp3sekChlFWbA0VMhJha8rf7nlrUbwJhgDyTvHDpz0LrJ8ywSlL1yo4qbStnBHz8nT23KDxg1
ikcDISTK4gwPH+pgQzLJdJY+ZTxYH29M3YxElL2tHSeC7iqVXSLE6FgPvHjDBChvvSu/axv9GAqC
8Ua7jsdikC66WYMsC7dTnpTVWjFAzLahUABUQUNOtYRYOYGrs8LKoXB7/aZVDnOmr7bvqQfI3e9U
U11iM+TJdGp5kIFo/+P86+9Yf6k60aT7owTD9niPheGjBa93i7x6d8Mj31T+P4apoy3ZMyqIQdPo
iRmJXhIq3dozZWkmZ5opwtY9EeRhEXrQPl6PJQ0GhORUpFu2VLvsMkA5Hq08vFThxJHYAA98WiKT
H4ZYq4rQX8lpo1Rb8FiechMNAGbRfnqtae7J/+CB1UT7TjhGs/90pdZJLPz7juAWHIHA21Sdm69c
PR+okynqKruz7MuIczYDrWiBKyaT20YxDfosoxo5+bYrO1TIiMUkyR6kLF2Wtgcod8mO8T2m7hsC
XOS+WUCMycl+GBFGLYoUZvU7dYeh+SAYOhQRzW0geKUIZsh3G04qKT3+PmPXoAqofa5ZLXZ6Bt4Z
jMpy7ckzOZMGvkqCc0j6uBF9pwrJjlml68oSvQFp6vvZUUAGdaWurQ51laJ/5wlTk4hV/oTM3XGA
RcoPjSNRGHG3aFRptXW+UEWlPONLNAumfFgizqjyuDQFjE1KCARbna2Ypx+I+FU7M1V+jWzrZfdg
e4ozFN4SDXbTXPuTLliHOi407v0GlhP3C/PQvY6mEll+06BQfpT+yFeionne8TQO7Qo+8/axnr7K
Fcu64UyUft4y4YUFO5wxLhymJZ4Viw+3vrbsXcJbOoRPI5XM9yJ+LN1X5/0sGXGWBh4pugegsccP
zx1VuVCiEoiQwbm+0WTnwSXHAwVJHMhl4db2MZ172cJstkFVzFzINUewiEmrKMDTuvzdwxcya3td
BD15VOceYGO+J1IvkPRRvBG+sd8h2p32qzm6uwKXFwNPNM0s2p4kr3+sZWAqqR1RVWQeu4heRW44
x84PDAgmbz6ezCKvkClJmxC2RbcwTCnemLw0nUCw55O589IDBRZJiW99+z/QOf+6E8Em7Udi3Rsh
bEyfJIORfbkqn02zDzU2JlaVmhzjxuBrUR/ryYLFbfR5nZa1BI3b2p65ECvBlJ2LLpOpZDpl3W+S
WfxiN/o30E3nuUnvOGSsRyzmHIGogSKI/HjV59kOWq7DVeYnranM70Z7x04PWlqYe/L/CFnbNn21
VfsRW4/Hsxfehqpv8CqwLAmF+Pdz0ZDfErpulySkV/Yu3xTHIMTJ6lcclW9fZITBPLBDxmoID80l
qJsiZSK5rgs1n+PtWGrO8qe2jzDHmEwrqXGFUh8/Dr3EVWmkKzh7KcmQ+b4aUEp4om3yocrn5Lmr
AH6PmDjNGblxVnaqroxUR7oGlAH8r2L0iC/nCT0NVwNldVAPpvs/vp9m3sImRj4SXpVKnYZ42GIG
57BXIHTSghgIEe/kdhY/nars6KeUclP2S+OA8PJuAyXpKtnsdckzdkodkdtkmQc3mBy7XrbWPRdp
amPcDjeIwICCnLqH7//9svqElCnBNUMlbQ/EtGJWYlPG2gdALAw4wXnxM5iI/M07+ommyCFJOz85
veVEzK2CVwFnMh+nvd4OdF/8WpJOlVnkjnkTIhucelNlJvsCW3KSKFth2GeQRDdlLaLUHjMDNQuF
CYgrj4ij6unSzTczXGvYsGFTbGIBAOBzRgiBYyBF7bAFS1ANEquoJZnOQFjwAW/1q+NmOJrjpDTK
AX/8k3I2Ss6oU0VMmqWlhDRSRwrDV5g5J99rGyr6adkc4lUgVqxMGNZ/SZO498hGMsnQtSV06kbQ
d8osZ3OS15KnxUVEhYFpdO8mk2ra1f0cTRuKib+IoxiZYxjQq3waOiFg/11j+Lsz9plZxEX4adtp
15s8IKkhpwoeLXncZIJ/J2nWCCEOmwK/GzQuNRWz6/23pg5GGAZw6EiVUagJyOdYo66MzXrXdfhJ
spUKBQDGLUaMooCZ96UvuxgtrwR7OMD9bXaQCKKY+OH8l6grdiZWc7bhdyTfEu+GefbXlsGAzDuT
UcvDiCpVMGlUgidX5aUwB8M6gY2ZIsREy2rvCg6wlBMXd4kWNwDEuBxaFgRN30Ah/rLzwMXLkbKy
hSDzmvQsOC0k6X9oHyanBFwE1g8nMR9EATpawZUEhZvkI/hC353ThUa/y3AMAGqkG+oUTXIm9faP
2dDcv3xWXDLYN8Ha/vA4KsZKlUU2ezFW7b3x1fy6se0foNCy0R44tnUlaPgSVD90XxJ8ccYfxiJS
5988r7Z869WaXnJkZJD5OEfmI2cPkRssKVXeWYdzq2JqVE1gPS6qm6fMLdLpQHA4CLq10rNg2Yox
m/cggQG1PpuGU4OYdo8Fj5U8UPAOb+7A+Nj8aYIYpxcWaY1QQIOkWvVAGVKhP8FtfwcuQ/f/o9WP
+W8QpJ7UBENussfrcuzIs2Di3aV2+N78+JBgI2Se3YJK9aAa0hhi+pi1v1LRGCA6TqRCOM/tDpB0
gITW5/+pf9A5ULWwxp/hV+ciQb9hB/dM8Zdkn0vM/7GVNFAh8xuV4uVFgyiyJsMU+IHzcauXwfMd
fgLMLuJC4EeXBygEZGxTJsbgwkC92bv/UBGpYhmpntDkhtmFkXQItF2TFugDAAbxyVkm4ThgxaI9
DTX+VvO6t4XJLNG5mp4gFIWRN3ScnRaB7scRFqaWKjISiIhILF0M18YiCmYw5fmf9kaqRX2nx8dY
lynK9tk15Qj/PTiSrARKw1cePwKtKL6S2M9ZjQKNizZrrfmup8XGmsyNAsStZiBVLbDhXFRbMiwO
IF1W/hD3UWjHcATCvtGUrU2pn5V7NU4rT7qC2yO3w9utdxIIUEFK0y+I3BcRd8MdUrm54pqSFBAR
LKsYKpx0BL0wYrhsGA6ScgmEz0PuMourORYOIRuWuq2s/YzAxi6Jc0VA1TDzEJmpqCWB4aG7d4i7
CFp7OS0GAGdz7xWSezvw2b3LxBK+TeJ9BZ45TKtH836TjhsUC3OVugzAw2fOcJYqCK+ZBnWBWOsD
kYFz9QzNRiX6T324nihi604AtrD6nGWZAgiqS7MAKGIU7b4QFSiBmd2yZzcSVP7u9ISBZ0Y4DC9C
i5UqNUShV2G+rzAP3ghMgRhEBgemgw7layR8c6/yMVfpkx3085kXr5e0bq5+rmnAJsI1s5DtsWd1
6iOSzvWlJdnxNEWVoXItxW6S9lZ9S85Zj0gaINlekmVnhu/GLWHCKHTCeTouWMQbIC8Qr0HivDS0
T7U1yIuYF+XPrPvG2+SpMZuwKZO6MRbLx4z8SXXx3C4REE+hsj9xwNUsAMqk4PO7ggvNAiu8lIeK
6aXWcNfOp7ddKDgi5ldyg8l5UVzIm9Di1qDfMOY/tX/tR5Na763nYX6Py1/Wp9VGRioaCBxX/Jtb
LadoKoWe5YjzlWURm0Xq4y/lxhXYY+3Vh4a5Zvm3Yf3O0ovQ2iyBEROusjtecfoMWzVWMydAUkDd
3gQGgBbVYPkDoeNFq7dwNc8NljUN5xHulHCMiyuqj7m4YFUyHARKl3COg20eaMSBYtmbaZ+IKK9R
QwW2h3KLy1m9X7crDwGjjvUqywMSaV1M8EfN1X5m1cWbRvWuTpZQ/6crqZ5AXqr4EFsvAQa3RtrF
0+qTk0NbvErpBKh4U81sTQI8/5Cz41ie6wFbPEOeYe8wEaR1UNIh0P3NiPiQJ2/EbDAX8kOz0uKD
BQA9cgC/efZxb/ITduGW+tu6UAxXkUkPefeha34Hu3onNKyeX4bDyBXTA9aWZoZM4BmlD9Da9wGs
46TC9HPTMVKs9x4v4yipjIOM0K4UTqmzaarJ0m3il9jhxJmuvOrH431WlHK+tezw3qLDGXShplzZ
jgfTvrcD/VtZksZKNrxw1eJWLL/nLw+1qeAM0YxTiyZROIa9n5qaEQMTo/r4iGorivDWLbHiD3dT
dP3wS+IC8qgblPT5WANg7k7+w2v+iUMaP6LaXuGVHjqme9xFGh75m8iSaKMNUWb27hnZ8NIYGESY
RjTe4mpsFT+TJgSh6TmCqcWsTziPHBhcqIo9w8KWLfbcAuvha99QjuFAsmsgXRLYpzKASDrbIw7A
3sUsmZ7i6fKdRJvo5S8F6YizYxFUB+GaY58nRGUscGqB/22iiEo1heaq3ixiOxoShlx+Sf+7f2d0
saxJHH39QfDVvYDpdkb00+GcUQEBtSyWJ8Z/wR8EkUKiQRAMf30/AheeRFRJuqX+gbpaFEkSR8m1
GI4HDx07a5HZqCRI7ftBzKF+0R9UFUjWrTxJ1pT4dQMADT+N4JrqquHPIOxr+VNhjFSMRfuTIzNo
2Z7q91DPWTWhLo379MxqXBivUHI2nlSgYGv7ipHJfDszsrptcj1vj+Tls8yQLb83Hf+xwgXIHknp
YgTn4B/lLJMGdiNeLYX1bMnFYSPh7w/QGn0bUyjx5U0GOuk1Et0M2T3sC0nplvEXbtPjTRwDBIP6
QARv1JfxFgPlEnb7nF1hBVPhIgLNmNgQn+RCdK8qDauPCggOwjT3/QbLPBFX2ptdSynZbMOZJbpv
Rcpja1h6oVsaYP4DR3cNCcWhm8JDsNlIgUDeduTEo6YX0rEzoYFebdRKPObW/zfRa4TXS6KjT4+J
XXgwfDwpst5BCwEfpzkZNSiSHZnJLKwRs0flv9xQdq59UYke1LZPOJq5m9gs2viVSwqbhio7jlL5
1zk2kAtxgOhv/PfOWcd3ZcFpO5pi1GOL9uJLeIAHivDefcE+DLQMNL/nNThzEvC5l91XefZfJPsn
o4NPz7JpjvljYZe5Yo5M5xhBtXXlO6LtPppZgSHXIa87PZFTKOdFyG9opFPrQXcD0NoKOh6OX7n/
sVj0xgL5qxVx5I9f7hR5sB53GyJ8mGwFE6nEKR2AAKTmx+MmuNGkTfY8Ck9DSf2iUOoGn0KzfEg8
ZMFzGoaEWJ63Lu/zmVaoYs7cJeDOHSGlkdYZ8KkmxCRbeRwHJ3urcCJyGOlyVW1xzlDMdDVp5i52
ESV5YxfJSnVte2eFpY9IURBTqkCM98TMCsAmFmtnSPvmqU6k6tjApLAdqTDCAyB4KtHJ/+SYAsOC
RSM3a7dJjnf57ANC1peoP+rkEu1iZONUdk7WaedWx0tVAf4wiUP0nBtvMCg3RZ4pEn04o4Nw8IT+
v3gHRDthSIWg5XPaF/DRTwgcev2Tu1p11RwJRCfy4Ri1cigmVEVk1XqaV/zPcmSfHG1eSuz5gKHc
sSnqXQSfG8SWGGjdjjXR35JhDU1EOPISMAfNufjt6k23EogiNRxbfcp7ymZB0Ax8yd5qgv8qHr5L
c7f2TTc8e3DqqoYYSgSNn6/tmPoqDvd0i3O0PG6zXlTK5H1ZquJSxMlF9uFjCTcp8q+qDgjKnc/c
wFP4FeUmCGbz1xbBoLRvU/uR3UtyMWWz3dxtp8X7/qSyJj9tri1hoxwhTLx/49wl5eYVKmSTRH3P
0dSc+G7ZDMXE9bUQhHfqbRTo/x5RfuKSa0uW4oDQIZ1NyFpllRMuVACPdn3jyUHF4UW/2bF1eVdh
SZxAockX+0RjIHeX72vnKoH8dFePXbpy/U49NLycuqlZdvdMn7xkew44xUFQuyfRs+7fheqGSckS
U7mAhxQ9MaTPanxzGxulCav+0ygiy5pPS3dOjC4Voj8H16zC1iAFPmHP6q2LWd3mGF9f0rqAQbXG
XJ+v0aBMOA7YskUzcaJGB1z+fIbM/8KFhDLArIC3xiPsgTtyTlJFYlJ58Fbcz/JspoMo+2AQjuES
9mWN04sSRNzf6xxT501I2LBYvGNNvCCZ1bHcv0QuZX1NIoyewPcORX3oaRWwNie3xHKGBB8mEBIf
VmchFU+eNT4jyUwq+aHFbP+IFWQjiujRnosLG6gNGoUPv+zmBRb8070veWOPos8wxnybYeyJR4B9
5DkjDu8vJHoGP5auK6nU1T0s2n91dUGWLZi9qIUaZnxmpTVgvPQ7dAEzilaOmuZA8n6+iQCAsBC9
jDBAVpCsJUCK1Dac4YeNBJ7vFZ2GBSbnr5clNCbkBlzXy7+SI/by+a9i4PTJDop4PaKVGm9IIScz
YnN/7GX28/k0y+P46Jm8yK4wXNTvN0qFS3nWMJZNt6fkcwwcvCDuF8s4s5kbl7zewNxli099dgvk
B8WXSGhY/OlWlA0erzR+4+4MTLCVKni5qxpdhWuCYAG5zlt2/0IYWhvAjYL3stsljA/VFGOcry42
080zKM0PSw8id8on8WyP+yCLrms0zFVu1pVkzZW2skJl/PhHic0aq709xoOz8HSUVH3dpF7Tuvjh
8fliwck4UEBI6v0Bp+PBXVz/K5O0F+3mNyV56vALm5ybr5GOsW6UG1zki99YqIPcnmRSawoGAvkx
Od5S5GX5eWG3KPfdd87j5TLPHaBpd8oYdx1/v0MhZpOLHu7Xy6TpeeXe3PSDvcq73qxDXUWLzqTS
C0at9tiN/xi0RJIgx3q1rGBpqRKEd3BtSS9CkUhE6EvxDxv2wkWcsSX5lTBPwYuq3QYShGasPkUA
Nz7OpkAm8xKuZx6kEJquGSuVSVKKdviT7mislHKYladuo+9TovOWvmkY99BaB6GI9LsX44GkvJl6
CZ6gjeWsqkQWeb2o4sn7zJVWd6zf+Hmb2fjCzYNvkm/0NDdkcdsM2It8qhrxKD8pKyR/JasFe7mq
hYqyjfqlFUiuU+9nedsJ8ZgFwJZLY3jLnrRBbtshaGX2TqBjencK4z9fcz3yQUGrpmPRNpWoE/Uo
8ZjK9SjnErv74oOeiqn5EJAdbZyoiBzIwA/hEc+RefijjKFLMHb93gK7Sl/F4a86V+wy+DSRMtoB
Efd8SpuGnWQhoyW7cROu21l9/5vpV4zTyshc6Er/qV8mWbEuQScWAnKKQ0+bcynsTs/GwkouymtL
fxn3NbxbsoptPZyjoPLBBrOqq2QCkPf+QrkU4Obdiqzi3mbN7Vj8WdsA+CkL+FWH29D76Xh/K2nf
8545pZSCZInQMtyC7S9W5cV2+ftCs664gYAwo2LIRUJR9TrDtc4jEzN1xUV/8B0lVH/STosUYNLF
ce7/mA4QubKFIGD5kgzinGJDP5Dws3oy5vPrGApt+f0lMjA2dsc7q1E35u94qP1M+bHbb9BwB0m4
gEhNTajOJHVjir9zL7PLQkxu2lru54gZ7Rc1qA+sg1Sn8D4nivU0u9mMK7/VjdACBKvIktdIjjbx
VlJGeDAlLDqqIIq3ZYUtUKbNv4gtYWSyk8bqJp+13gAhXz+Y6SasPvlgFRX+yDaaKoJMFpVsxsHW
I47/Mxk8NCLh5jKrSR/UbtW3KughatP29+VFYkjtp0x8rP+Zvy+lj4yHf5mpUMocdYMlHP0sL7Qd
B8gQPWZyDYMJttFBx5aOVvhSbTMq/6OFAxwVEbGnHEzcV0Tm4eOkFOUj+y383Z9wqW44JEyXnVlZ
3eBMlJbSzNvM+aI5FXSId9/ODr2E3pxoBjCdqOJOFem1KMeU6S8yyyNRvhhiyRVhN9kvPgIHCJpj
EQ94LmrJ2Ikdj/5/rUdkzC0kraTie5p+uEOCSA2DIhME7QzB5laodZ2MGTv1K+pKeXpfjlHFMswQ
l9UJk5X65+zFe0pf3K6TNhxy3ZWQr9Vi9olLyTYZkGuVEeVT+wEhhviDzqNW6ghp1nDuExj9ojiX
CNCZJSUpk3/gWC11UO6VZK+kSuHXF/mBFl441wxEiRZtmN1jvP6TuiUy0UI1IUraLaZ1VtS+SgWP
x7yVCSizfiGQVzfUUj2OQ74CmP8r+k9j0bJW9ym3ur5MJk+XkzDi8jDWIdkBcjPLVZSC74X0JlmC
OJ3nf8E5WDDfNwwyDfnj2nu2eBem3VJRskHYDay+Et0PV200P7eixYn0QSab+nRUr1DXdEtAq6yd
GLoZJGUDlGt041NiGdviaJCbBs3oipylG54oFIiFxWJeoT5nu15e28GA1NCvHLkiFkfK5zOphgh3
ZiRaDhQWFrGw0CszHk5E+/arRF8vYB39zOnaPpT9Z8PSV3ZywJCZmZSA/g6ZwCvMKRw4KhzzTwcl
gr+WsYc+u/nGXoV/Q2GqoDQ3EjGD9GvgfvDo+oAaooyHqIWRBMV4m0galJ9ZT8JDVgBUlRdvIGiZ
+03DqNLlk+rVA6h8QfXt4MN/o5+xI80YyDc6wsnCHp4ThAUHM0KqZ+HSpd2BEoAsw8TIZTy4Lacq
ygZ4aOetSZ0OCkH0oVtcveEh0N+JFmmitwwvWV/VniLFqV1QPSNhAlgODF9w1inZn8ux48A9+IgU
bdD5hRQRPJxXvjj38aBiZfh33zcokzeo62aJIwHtj8v9V0m4U9pEwL79Sr0ruPKqiCEJHm2CDwv+
twzcsrodq1ezn0tQ7BYRiRhZX8szInSb5MxCYMQ/vy/PD9RwXBVm/+I9rg78eJaqIUb26XLyo46C
W9WbS5huzwTzfiyW2n5TtsbP0Jexwoz9C6ewiaYWCBygtlf8emzcj/ez3GSEo+Drh+ARsTTzP+3J
EDu8TY4K/nnmc+4YdC5U2dzp+qted/Gbyvhod0QSp+qsF7DFEZMFSPY1I50cq8H9JpgCr4pasv66
0T97ZqBZuvvIDmGseSXd+1JuwsOOuUqdV2+qbIRfJbtY8Cb9d8YjHLXbBEhsmxnebCelt7mWvkks
KgSul9XavypWTwMUY6wcYRTTzhnOh4D87Uy6UlowPybcgEzR3SjRIMB2ZMchveJ2Lw7i4Qm+Klmg
zZJExhRw7kBXCHlPAyhF5rurZvbKyOEbUrB5JhcubHDS7+d65Gr95k7A0fAXLTCYZZeU5xFZ2ESX
ocEaIvEOdulUrYcEZRDrFnVVOvSZPxh9jeBa+yIrD+wgmlKDxcQ5EYYQSm/lZQ5xephRHzSWQHBt
e5cT0FGkBXQL5tmsksypfwIx87fa6Q9W3v+tjkPh7Ltm+nT16o7pCK0Z/VT0Y1+MC2BsAgT+XZLl
Hs8+iw+/zWpb7FWSWHr+wH8LLVauPqAqEq15Vqjx7tUYmWUXYoUcNS4Id2olHemclOZvcrt3Nnip
vmmQ5+RhWuxI0tkpuGXc8bJgcit+USg971mrlLD+V3CEJucN3fvqP3tK+mCUqQutAd0lKBve6MuH
lbx3waHbqFmD2fgjTGIopLzgfSV0Jl7gz4iDdx31sr/DmpdmZGBRrVA3PieeACng028XlS4/6kzm
rkiQBTRnPx8gASk4/7HG34grmFaXi9cU2HAZVX/BX/EIhaZQZYKKAIlLV09uo4Bzw/siSACgPkiB
vOP9Pvxfahj0YY3hGN6obuVgIoEnmMuWFgTIZJqtTrLwdd+kEsHz5A232kM354wtdYQnTJx1odyY
0KUNK6dvl2+IArz+UXEhV38VEYExGwgfOkK/p/gsJzB/EIb9zPKKjoEB5TP+tKBt5AyOeydAAmHz
9KdN2V2Unb5EbDT8L+/VXwbVitpipjVP/gk24aL8mW5cAaOVFbF5WdMxoRKJ37RR8GWNXf6d1drg
ULxKB85baVemfbHgWk/sf+KqFfywPwzkiNGXe0AlS+ka8IwxdatkJpLjJblsmQhGI5BmZ58M2dwV
XSm6tAdwosBbT6E4Mi2Dv7eY1P1//gsFoVrc9zPI3IS3eZZYNJAGzqUO22DqjauOqxCzmO0shvVt
3cvHbpt4rnmeChQpqSXc5BoySXAMgRgaWVx9gTvI6oIeUy5VyZNqaeGDOnQPvSFpNXMT+KMehJp8
Vay7rg8RgmFS9tyAzS2CtnZ2HCuQ/RePREWcb31w3WoiUMATzo6xnBtLGDhyXc8pqSrAGfQj/IP+
8ARdlDre/yl1bj9DaZ4T2YEUBUl7pghirfHVZpVfIVLoMpVvdPVvi0hDpZbkfV0bGP5yRg/pDHt+
fQClfSexb/OInBq0DZGRvEfuPE/omVWZm7Mb/HGvBNQx1Bwpcwwfw0uhjYujOUDSwxlWEADof2In
XXuA96Hmp2EBjQIskrpBbG0swJ5fAv18MBykaO3wsKW+owNAu4PxFBG2QjXkzBM4fSLUsun7w+ft
tkhvNMjRBIDtrNqlDEETiZkogbzUr36Nqs8vA0WSpI9MYDPhzFAyTDiDUXvSzqT74eKb/cP15d2V
ARTnKLmSAeYgnWOE83hIbZO2V7/h4Yq9h+1CwY8DxhenZZj/oVjZX/MYMWNEA0WXjEypmARoO+YO
xERhAhjycHLcta614C1vFmdCyPSLXzuubKfzgMHoCBVOYmsjVsUIjzO2W4qnV8mOkvbcpjJ5eeFY
davxNyoi5vsbJi6LzsmZW0aWRd+Viif9xqA3X7h797RhunWFZrGU1lKMMYqZimmdeKRKX3OMrnoX
279O6y3CFmU99iJ1oo2GaY7BFBFrIhziDuVymQMGawUzUwz0P/BMc7pn17I34pjLEf5O8jXaPsR7
H9aG3v/z8DRvGikOEdcxYE9bnihCKBzdVHz7gvLN/YBzkknLnqKqPhPNkIf4Se8AASqYQ5FiGHDc
7Z1Kcu7wz/sz1pKNdvbSk2WSHFj6s7o23z77SYeuK15ldMr/zG2hkP9OwKX/ECg7WSzUSPjYz2Sn
Q0mrL4G2K5ETD2n2I6txl2C1bqEOwyaL0VwYDxFocSdlUD7jY7aBfhgG0fbf7mot+WjbR5KHf6R0
wfZHUpq7LvEEQ/g2+LpMRJrAbJlD5SjMniJISzSIC5UyQcUObXcqjeeuICdA2UvNCnfHaYXFUWX0
12Y2zopDLh8/UqIJ0qj4A1WyPrluz+W3A+gioF5CsOoFRivo7fm4Anll7Bb0vVDcybh5VcC3J9o4
L5kzgiA8hMI3Xb//JQHzOWNbug2VX+TlWbkqDY7wX/DyOD1clUcHSkp6vmMeLz0s8GA6Sld/7d5Y
kkTvlxGHy7Cr84xARZnEubUXR41oyYCkE+qYojJWkzTn3fZaVf6cTxcsxwLst+ojrHf/rKMPoSmA
NH5tDaS2h9a+0/QwYeGOMyVyHj4ca9yoVJb5LqpYYbl5k8PjDDE8/njf18DPvZy31xbEa+Rkk7Iw
9PRKUMnfe3jJ8NBg4fOKA+MR/GTldrIVl3ZQh6IEA34CLMseP8huWw3fyHNXjRYwoInNjuv08knZ
umFmavyYFnvUmS7xInZB/MBOVwykTd2aV9+QJsyk5K3V/7rRTndgDisE1I/8eRt/Q/5RQuBJGEOW
yFJENZNmBu5ew4cuTmqT1aeIJzxrR3ghto+12Jznvv9yD3QRdgMMExUxbkx4k92lUXy9irdkTi7U
ejyONblR4N0ihw1A1vP8iciQ39bkNcl/rLDat4wZuvjHSwK1F1L9Q2W2ADVBxdPpYn/w6uNSDz+y
kphiQye8NUwBL+Xp+cCSLgz7rWPxPCDTt2Jm5dbbcw9oEy94MSEMANJpK3r7QjQn39sMWqvvT3+b
2R8D0fz6bFSPzMpBZ+AqpktaaawZVjZhjaipw4B350AAEzzr82Z65bqP4mTpE7A+L7cC/G2CIp33
ns3Ec4YVCd/zWgK2DzCweXARWJjY9kF4uPEo5f8baXJg7QHnvptCgPIt8Y6upcjzbZq6WBwlEX3h
jbrmCwpl32eXa/wZ/jWPfx8/qiItPIDuDSTxcbvuC4hw8+SgK+Hrux/BM2vmZayj8UlBGv6+Ys3j
iH7fj6daMd6KwOdyRQARatnelltGl6xMr1k9zlf1/h7HAwruOy2b+g6lTllImlyGccE5qJRTCTPW
SoH6yb9cWmXlUppzgF2gFcdA4d7HUWv3a7NxP07T7ai0lM9d4N6YRyOiJaJoRpPofChMIyqTpFUs
w0reCp7CeS3rbN7uWkMhQWpcnoMFOu/l9ysuctv7ou09ilVwBGP3i4K9nGVAgPen3CHb90emGc1V
djQRqPgW6OtaDTeQ07DXCSuTOI7/AIrxhbJG3xTFVMKuQg+N8Cf7FRcjKGo0kZ3nE9muZEer+T67
d5HdTNEJ5p+l9gW2b+U6j0DGiJhMk3Rbq9yleGh3HVJ0vDaBV1Bpkj8iK3vEERmAyn//x9nh9YG1
Bk4GDTeOHfSCaJt3cy2LsVmgjYkOWdvYDJNG35ZZ2xOW3+q00T633UHOL3LRpqMPoXsKx1wW6dtr
VsUXsR7tOiFeWD/JpSv6/PTxLiuGxmDSY0KCKtmUrk+fNrHteWxwzy+MsAHVq1F7YTuuNo3gUE+y
GkqgKmK/vAtHn9ZBHG8IEBkXceD5l6pyOJ6Bjg3RrzEVUkkJJ+8UqGXx4qyqUN2mkAoknoTiz0QI
OfvyhubOqSHc+HnO+YRP19aH/KPUvgynjv3jltRt0C/wt7tysPVVshiYha6knA8X6gi6UawqZLYN
yab49XPHHAbhbjymJWaHs5z5kuuGJJoIBCPRpVruq27PIQUxU+6wHSP1kFdss/kixdreqO2rxXLW
CNJQBGw66zpGcl5QtdxQH26DlVKYQS2d2pKo9LrPctof9K8s4ywYrUaKwZOE8Vprsq6AbXV0kzbE
E22Noehgz+ZmqZvnbR2T3P4JE5oi112qE+6pI6/mvTiQ5q+/XU/4PS1c4sOkMq8Kw/L53tRGGwBH
GjAizVsOVMlK+f/sgAhUN/dnPAT23plVyeEqNhFnl49X6ctBzjFUTkRZcmPKiY5cVB8eBAAoUZuN
ObWPGLzD5zYgQIOMbM0B0c2+hC7BdSrDVN8Exlw67Qdj83UjkjStABKX24lrIisMdlqdtc2GMaHn
Cii/qQLCV97GxTsKDkK98phcxqiSDXWLhaWM40QyvcqM5v/chSHlfCELFhqMoUiCvtntraOqLqkZ
0u49UC0C61x4yb8HmPdWbGA+DaJD9Rq1Lx1XCjo3rLofvs6r+yrJZ/rB8OfNk0xtcEkFPJquo3ND
4kkguGCPBnOsOFLFK8xXKpxFiKq/ZEDWGvlbOV+U9h9FYZx7PiA/pbjfYCB3CKUbPJgftg01zGBf
CE5SZwPxBvdRIeLSBWtB5CbNCjnIYVBEs/xWP6DjL4PPCdVjzf6lW1WrYXnchqDeWU1NQWME19c7
kUPktT9m5Fm5iRm3QqaMa1ZcYSfKQO3/fki1bUgy3nJjuZ4e+9WAI4Hfriy4uhndil3oWqEeLJkA
87xpDK1vci/aEXW36iML0AFVClat1bEBngFqrDHMQ1dgj2tMPcOo37bcI91ztZPRLgKSO4kYvwpW
/rqQiwiLMpdeQnQWEz08A73HhqkPGTdg80vfmw5ZU6JtjM1xIYn9a6Lk7/DtK/EXum9z6iVeHubp
jBIaoK6587M5H5Ewbf8CHoSBpRfXAmMGebyS7M9eFw2iFIkxkKm2JgWBNYJYnIYrqqcaHyXl4E23
adFHDB37s5LMxnC9WSBcqYEIz8X2s/xWXUosgLA+E3sQLjjGg77r4ppqX8x4OmVrrMpvmhilt5Rf
Lix7d/ZoMLWnYo2icyB8a4gFbO2OuDuzBHeQf9INpKQV+xlc4NNgM0sNn5AkYqsM7sD/avgtb6VB
ETpgnCWxZIOUOiLNP/zAkI1sg6Vl+FdbbYbgVy/6A7SLND5uku1iFkpDyDhkrn03Ywv2zBKKaFOM
dQmvrOylmfdAQZfptYOb0vpA6GmSCiCUmQmxejnuvVe1E2eTqucVn6SSpqXqkpgudL/0qz46cBbJ
5BbEUSHaK10PqIptvAdeLJSNxtA1iUXuiupnYxhQjggmXreUTia/PYR7yoMMMffCPDkaKoHynOiE
QXyLE+QuGl3WvJAfXqb0L7oqGO1zrXCbjIN88r0cE3VaepCPY2V0LOT2e8L9OBfUMF4VkvsbaVsU
Eelt0eGx1uEs6uFJrNWKyKmy9xYBGNFnP/i9aitrgz8Vur5h9GWIHXSMATSbLHrDyIqADiNDbuah
RBOOaLspWupui0Pxs73p5N3QjZwUpufMO00Rl3wPJ4HZr+SuglyfwTRSZf+dTUIU97qhVZwwY8Nh
tNWi8D9GNRpuYp65xmspyZhdWWwE+ImmTv1EKes6r483QqvAXl20TTlMKhRKi52DLaBoWObhLumA
meduNbRyboxd//jqNthYPkhZDsqOlb2enetk2WTn9ACNrH3Sn17EUcE7MeqFUthKp9wSKTfxmPWf
8GOe4Vukt/R5nxr1HmwHCsgwx574c7S3/mLHbQiIm972BbyEuvjNGHthyvZ1/oosgPw1Mjn6qs1A
/IszqkQK3UpVtWKENF/4f/e5ds2bLDObpPLeNgvS4Pw1Xv178F9JzpdqlL0v2F8o8mJxM0//W4vF
DC5jQg4dEte4YfVGzvFMb/vMu0aH/seNfs3yzhTW8XdyFHzVN+6xYVBbi9jDccSacpzWKKtbqDVL
Rlr5jXLEaa8/rEAK3YVeB4Sv1UKBFpXtDDGuXIUEUTeKLTWmBytAyM73m6DdFIVEK2m4n67NJzfv
ohp05xvmNmyQwlqflN96l76IEKBk5Az4ug9s7NHms7vT5BjZBBN7ZluouxmM5zUSnfy4YtyIP3zg
dEO5+UTANcoS7DIYg0QvMfZBXJDtfrtI1YEnyHKmWVkFR3sSmNNm1sBLvHmGe5atrtW71F4Iqj6b
TeZMANFvJNc9B3qi2FQzG0NJKjENO7XVVogSj9jBNz3IobFtv51pS/KDh7H0oiM3AHjX1/lf8Kln
m3Nvcu2DeLi1waje6bbaZ2ycDnTAavpG6ZAOtaK9KM3myWPvS3Lx2XnwsAJqmlgxbiqEdBxqcNv6
Xnm1/v6+4EGoVOI1niIHELF2gz1ByPbJBrfk5xp7My/kCG1evU0Q/QWbW+cNztAPVAVoCCpk1pQL
6XCjrbj+MVyjNHkOok2pmYr7ALpRt0R2BHdNAZy7HZH4f9/SRZCyAqJ2uAJDsz9yJWeNV0dI6Puw
Hq7HM6FYBPdufH/c1+5yPtQ8PxCwlRBxFWXggs516TYGf7JPKRU5r9dqcPhR9v6YaZTbL7L2fUH6
5gY8muNS9o4hMp8JV3raVwKAQlwCj0CNUQGvYT/81Ct+G27iPVZ/uu3jYs94CWK2nrWUx9zZ6Z6W
kOpWco5eAiEICr1sLK5USeJYSjiCbVC75h30DrN3dNNDNoSMPzmCWLfpQnODDC3fx0lKQh+g6ntk
yLB2110ItHVVzBNnkIUHAlll+pvTzVqy5tXMKDj32HaLFAwtmn87QrOJ3abPdjiBfTHJMHeXGfzo
58jG4GBz3darDI05rVT+nvn2jmHFN/eOWNBEaYFcE4P9yb/3reH8vhXNyoHWkYM8eadE5vBgcBDV
x83Yzz/+gjWQy2GmVcX0CR0d4zEKLVoPhSX/1D75RQBwoQ1X0k6mhB5xpa9fAu3GQlKBKP5cYls+
fIxaOe5fW7JZii8jtLFJJ6I48aR/Qievb/r4Mhe4gz5KWL9XxvRDzYTg/uMKh8odmR5WsJZI76+f
Z6ZWsvCSgYXyN24JaSCpuxmN7LLCiCHWu3miaGZ+hCZUvTlcgthH1KX8e0VJCIorYy72GJSoNc9I
ty/j9oZYM89m8Oa3THfuuZ6svEWoiYb5Wg0sWikWHxZmIwzhPDHXSJS1VuT4NdAkt344ZISYhXSD
pn8JDWD0I+cvS3Zxm3v67TpX6nrR4cdgtJDYFDZDua9ZRLZIdXDeB6/t4wiHG4A0wjIcvJ2R2NFb
I38GFSL3TxQAT33Ya4TH5lorz6u0jitBS85ddNGJMTi1Nv7xZce6cecexdrBhikfKGwL0t2W30Kp
i6wKd9g3WP5lfYNwe2ACcI4MNYK/L8HDunKT4GZywvIHxDOSsttq6yhbYI4m+bvS13m302eYypI7
3C3inGA64+CMlyR4eXui5mYy1xPBwSHtaCFIy5utsCHt5QN6IjseTj4W/a3lYaJN5f3eYB/mZrOE
uzdmbtQwVvDBcy54FnuKQ2OtIOKwuD7qvwxByFo8ku/KFzPs2oyD7RBZf40a3Mj4RgylUFQWMRLp
YfCAN5b/gn7toLr1r3h5yQvZm5NBquKY9TSm1Qpiltfv/G9JRPYKdxq04ns08Jo+VcKY4iCoNZ5R
kFshYYY3S27oV0DGNtbh8RC4Y7SSS1Oyl9ewUBNkuCJ/abMeBiICLxDaJp6T1apHDKwOETRYfBtP
Oi+YhzkRl+w8sPwZtBN7xoRTH4NCx3xHtRwUJcDoRqkaWgnE90jaZXxswQl9BpoNLClVRO+/Ut4z
wdUGjoXzDxcAypuMQmFd5SUv7+Y7RMKp4C8FmZ8t3U3sAoCZQ0tmk0oSLaA6sNIqJ/qwetaHZjYq
q7/VoNh9TbvM9gBMGL3sjS67YWssSI/0PZ0VplyXUSGKrs52GnpuEh+ZARRggKgSeGkS9pSnuXva
uj7l3d/fqA+0ul/j2lWK+oWuMnfixE1//0ZZsQB9/Rmbaklj+sdHmLr1NjRUz7Xs9+YiGdF/pQKT
Cj5cyVVL4hCnjA9Iajt4Yg3qANxtY3UR3EcRm0EUtKd20lEk6ZARdQOZcBOrIpPj5xB6yXieT4rE
KjNVT24UuaRynMwa2DilakyhJOGxATYJE+l/WYXRYynWysYSTdPcOI7zo2MgJKJDXoNdauL3Zmd1
l9HkpiU3F05YM9M9bLmOOnY29lt0wph/xmsS6IobdrkAfKn7mdnWupijCzaBY2uneW8yffi/g0jr
DiTECpHbk7LPwyY+K9PxkIT5s5Tbp6/TgZysTZhQT0DjAgTE45/nzaz8WmSmZv7PedrKnuOo82Kk
YSnGVTNS1C5oqQGQqVYLuMe7x4Ysz1ZzEh4J8NJL8JL8vKb9VWC1EM1zYyNVDEOXe08+gOmkM+37
z+ZXjfzrvOzYzqFEYAhwGOLVN7xdijNnhQYVO5sXjQRk8/jqcY+P0TQbZvq0Bs4zjErKq/fB9Cfd
Nz6ewEo6LD6lOg0xchpEZ4/dvME7okS9UtxZ4iwR27o17RONguDEk/BCYDVXy+4iA0FHMYBVdzEd
+uLs5r8qqWdXE/PJ9HTu325TGj/Z+PP4laAy5O67YdRqHKH+PQ6wios5ndLJlFiqWqj6mJJkzfdh
kuiF6KMtpW8UlNTcd0jSgCvL9MY51vLfIYE4vujYIbRZdyPK5kzS3n3dgUusp/eot4Q1Tkfk3TA0
yfQNtfMeulPRjU8HiLMufPPsTI8ZcS7U52uEc0nKBlC5vTTvkScLAkMMnFU1IwLKyjwR1ecDxL4M
5sYOWtmwaUMbf40c8QKruqbkDuayvSR56c5iMcO0a4OgXbAWbTuTGprBYWSLqkF/olgbbsZzQw6H
4YPaZQTh3dS9CihYjbF0UeSNXO3xNskSAOIuG/CbNPa32BPMaMtz/0iVtdiER07JASu1foNwOxyy
AiZJ5wMDP/MJsunlmGq2gHqzxCQ/XdGP7VhuM694d/06pgUs8it+/oduu8dDiqQHoDkKE+e28AKf
l7A8zoYDJ51Bp97QQhYAWc22HvdAHD8jXSUaXtnkZkjitwTIbEifMP4RaxyrK70iSYOmpbpFtHxw
/xRk4DaYqPo1i1sbzzPQ0tPo2rULO1fXKp7naIyoWiKykoOP31V7VfFJE9ZD6CtJmPkM6vC6fPxU
yuisIOJQMXEE/xsgSLbmEC1q82BK5nz31Z9N2kPLXeRwvaBGylHDfpFznDazw7cHz2HWS2Wh/Z1V
Wx1GOuxX/klzB9diXVQhxY/wsnJlIj7xTCJLgH/mQk5OdQOM+c8yfXjcuSUmJUTdvFyWuJR8Nx5X
pNyBNOuOuOa7t6PE44kSyWmn0QCR/cUZ8vbZCcaEo77UQGEtdk7Y86QW/gXPL9gvJaNc0EIK9Lsu
6DBFTXlbm/aX6aP7tjk0CXWPvDIjxA0gIr8tHnomCQY9jIZuig9x5bQibcSNhTX1mthEXanuTXn8
UvVNGUU9zcczqRMOuiTPrin16zVORhzzzPrJ1wc+UQcXJ7h/aCV1+C+OZgAZME3Pu1iLYDHkMifM
VPSw3QJoqiqC/cPT9ubzMWruzJFDGNwg1kIxRQ2Az70SeIsr66jNB6Ca6f7xPj3aFXiFcwqkO72U
3/M0yZ10NDz9+Imwo+9J7zynUDnQEYT4qI3s2ZYaO3VhZog60yDi5pUpr4VocC1HLzlCYNAaB26s
DkIsLDMnruxfYYH0LRRmAJVCq3shhDxiPVexVC7LC5RlqhlXnMR9bGqvofZGgMlenlzqaxQH13wt
4fOc/crNkjHHZdRbVYGcri+xx01VnBX2RIJyYC8Y3rsmoGIKFQXHS7eot2f/Kx3QYJnntDGESGHK
2W7eDRCwgdUwmKPIX1X2nDKSrLkRzWzeMYBSUyewRBPAt83n1V11QFYvDThHpecwc25pq7NT58Es
IT3eyBKG0VbBj9AeiTfTbHsrFsC0bwxytSXtgDU6L3Rg7Dcxf3xCwSWIyyzUaE2/nqKmFERF/5Gb
Vwsjj6dAYUaAtpuEO/P8PUhUEazM1tkP+50rErMBBfOcxamjZjpgjOjZurU2iSIGZcQd0nI+4aWd
tJMEsv/vH+PUPe0H7NY3u1Gn3k0CkiqgL23M91c24fbuQjkhKmCJhj3tJFAtGwtVbq8ztAMbQoUx
p+1SMgWoBv0URpYughf8bmLISbpPZgYPksrilQHzz/eGv3V+emdabKKsmEGFsajDJY8n4Cf90pIS
7by3HlHbCfVKqyAeJHhhQLh/G2Z2IyXfO3o8AKGf6sKhWeLDKaLhwge+4AI7ZYLPGYqVDsxKT8O8
Qa4c4hLXeBj82wj4DdfK4zFvLcoK/7TI6oJTy1uxSSKXgvv1gIjh23HegqLHoNUSYyRUqqFheD6u
Xo4mXLvg+ZKHTeMTTTvxvbSQbEJ1O1MQEyTzFgnG0zYE6if8Q9wUWdXQtgknSAiRFlQCSFRL2vRE
Bt7LPufDlCBirxgu8a3xJY1Tsm0JmCxmBKjRl13v6kCkaAOSnF2jrVJZPOq5gmAl7vmG0DhqsGfV
ADE/AtJnYx7EtScV1K5bwY1yaUKNiXX0h3FDelB6lim2YHfLx4D5DB4AhDqpWCxQrAqM3ZAavX3e
NL6heaiZfIOePoAFGXzl+HMmo4kdAbX66c3+6FdZDR7oCGuYnufN8E+RW2K60geEkr2pGddV8frK
kzQLFX6hpBrB50QdlGrX9LHz5Oyuqqljm7ha+o7AOd9bUG5rlw9mHHbEBI9m42vaS+NIFsr0O6qL
fjXFKlee8JnYbeR82lDUtyXCLH1kM2J2tBMBCv57hB21yyXz/kzRNzR4x406443iKEz+AjMl5Dm3
hEGtQkHhJHyuPqGDKfmXXh2IWVUBsD+LISUNf2FKMpVf7b9+Y/pW+eTtRbuZyrzlUW8DttLvIXu5
Va/YQeZ9eKdEEPWhdfjCpxIYMQciCWcLkkrPPxoCbVkxKWDll66lDgvtwIncs9MmM7B/i/wm2Ran
oSQE/3+giLUFhQXDkstB7xNeEVBo8CPP6BurwxPUfw/K4S3jVj2a1ZfVAZazySZVcR2ZUYFsHuRC
HzbwJjRVgCgsHSH83KUkW6Kq0WuWlfVrzddInd9fYtaA38AefIPP8A1kHefy4/m6gcpeM9NDM2A1
wYxReejzDCRwsLwA2xb5ZlL3RFMdhCK91VbEW3riTRVtiWBqwmtad5Y1RPcR1FxFOn1F45kqHWeX
/wx4JcCoNzQIr1WRruv7Fqu28zdG++eFfc7QM3E1C7GwyP94cbDVyaJIWaNT4H4nQDV4L1JXTLe+
lFYBseaK4VzK/YDMgpU38Qk31i6hLxJL7xleUNaVBPFlsv8LIvVZpgN9VFtrYoGSZF1emavyz0Xn
pL655znl1SKIiFq3jBizxdamR3M+pqshomoQekP1nkD+/o9w7aJ85v/+49+T9M0tHqflNXZ9hO6r
dsxK98TeMU11IDWHCg6z9OWymp6FdmU4CnLcLbv6Utm96RZMcS8/rPKVavSB+syeVhhd4m43rVZm
eveKAz5Lc0d5fn0A9Sayj0P53bK4+hiubI/wxRr6a45VE1OMNJMiLF22/ReTuiq/eTFHY8mGQRc5
px1C4GtQdvaE0M0XwgnBacLIu0Ei4rMSfPm3OGrVXNN3FvDKLzLYiYOaQWtXsNSKxmHdK1WqKchm
m5Qjp+NAidCVI+sh0YQcIvCEg/aaKyJ8OXTrmsy9ovXrkwNHc8t9vCzbnmbOrY9epHG2DP8cLqtF
xrx1TW2uqFGghZlti0E+/4AqVqA29MNvpVOCttDW3pkDXr7b1iUqzDEgDJZsmzEJ2U7IBv93XiyK
Q2TsV2i7Ier6mpaKkPDq8UsZ1MVMR8HP21WiyGvY5k4aDOJkg3/0EFkcE6EiF4BBoWtGOjkgdlhC
vrLnVc6EoOeaVORRuoYpBCSwY56x/bMb/aJeJ9kJc72Y+anq8OXuE3rRahGJ1H4rr6ypQZTzSJeo
MW163SDkPwj8Sz2NbG+2foEjULuSPAVRN/yd/WbcTIL8G3V7f0b46Jh711MrMlhPUXg7BAZLhRqp
DOYhaS+xhr94xRO3dvhIJP14oYRe0mf0bX16Tr+jwjNG2ZeHWYT/OtPEQeL6YFOsS5MeKpzEbYKZ
hwXA7pZk5OcwH8p8cjGF0UQTQl5EU3zLQ68g9sbKKwLKnASfyVJw8MVZoK0mLKSAv6QDqG+cFjDE
wJl8XA4z9xrM3nkzcNlN+PCDHU+NpwdO7wpie/GIX6FuENlDyoy2qQVowPGDDyMdZyncMKdoG6ux
IU4hFm1iqZlSwhcCa6ugHBJZ/KbODHpGajREQFauVIpNomDCpmUnriciyFu0iSOdwpRevujcmEsL
f3wedJZto3opm8JxVXlE1dmnIVqFMnxJjB9rWTMl5liL2oxIiRSheYEwA8xPkAN1BpolI+utauRb
W6V1ga/eAFWjRMtPLLhdyyROTrh2N6K/o6E/O+c5F0Ssf2N18aQYur2qf0OD5qOP0rGCoH5O54yL
jwVjfGGuSvs3N07bc0zg/bhSxyO9e5PxQjDyT0bRzGlGd6AsI6ntrGUYzOffmy/ZHjIm4GnLjmjM
X+6ChjUiRs14Km5MZgbImCWqWKFd0M+szVaWM34K81psLoGjem6wL3BhqqyKaHoPKKwegUsS2+dy
yaejIpdP4hWX2A0FhM/c3jX6E1k+xZrn1WJF5ApHaEnW0AqVVhoXHtv3FTvT3klDUn6EerwZlJBd
dfxffm5hPYadWKgn5OJOHG2157Sw/F0fe/M6iZ1b6AI4zPH4ZY1Zp8NMfTPAos87nj9zqObyctaj
/NvEqX+Tvq5Db9EiPk6NG40woWAhS2UppW/gDOaX4UVdVIQL2sP4MSEUvLsjihD7jGlCD9LUDuzf
lAMOHjKKuZkqm7RpUMC4ddZ3eGTLUJI5LF7LduL05J8oPQtIPv7QmWy45LtlwkL8KYx0Ifkd5HeT
qQ1OcBiO8kGz+D0iA9WgbsOjqekSyYhaEbwcPSkJYKHzHaWzq9pgK6y4u5pHdUF9h+GABGNiCcju
KgPjDJHekG4aLBznVWEqZUqoxP9/ndkj0lbPu3/+OW56uHY0BI3p4y1nnks5m8vVoNdwg47bbE9b
jIDYO4VkIisl30P/nSGEeD6IvHwRRQYsQjIbooA26R8HY1AtnE1O+M1mqAINX7cb/9kPswG1ZRit
JqGNizEJ3Vj/n5iHRnVZdh+PrIv/q+6Pckf+cYMoc8smBCDh9OpObORj7r2cRfjzYQ3GUZGUV1Ro
y1FfTRwc+y8VoVfuiIP8AbvRcWYHIESX3vz1FdkwCiMxolntv58856AtGcZSjuzVJk4DmJdxrEoI
9gu36J8AqiH6meIeSolImctAhqGbnDmuRoQIWoAwMw5tSQzOhdjK8YTqXZSPyYda/HqgjHMCuITq
DddF4KwzTlKC4oATsZ3Ow6pxEWI7IwUFnOiiB0Wo0RRbC0evaSWshEOCIJ4Tv06Cz3FGpbdOHyVI
xjkatbpO6f4WxcNpVA65naY+2wzJ+/tX9QHsj52I1ZN8j8UijCufRzJg+0xwlPG0OgO9pS8GRB7l
sbLGrJF413q5cM1Y7i6tqJBgAro742NaFVoe99tkbaSj1WcRPNhFzaZk4GIBk4ha9g13ZnnDN5nQ
V7z9OvUWnJI2hILVUerEf5VTv4zBhtDhfKIpMnOE0O9yKpvGka0NgUBXu9rDCtBbmcDv/d6jKr8c
FlQLa0d+FGQp1ApJ2qiY4t1Mo2bXReAgEJruqqgm914yNvBFjbXZQ0RYIl8ra0l/mxcZMGmCjN5k
89zSLMNWB+m6mHbvNPjdHz96MumJ/R+g8Vj9lQR2TVoZ6Tvfy5u4ozZbPG84wfjn4H1KxUbt/pcs
4QSDaus4tPgDSfAsit4L2GWqTIMLtID49dmNypqoyu/qN7xso+WYhYnYar7k3pGdbZlTNhcZ4W0n
RKCkHk7E3RCJGUAjh5fECNLV6+775qi2GqsAgOd49cpJgsaT5Gthc542/8ijBljrPAE6Z+amG0L6
u3DyZ0u+KDgtoc7bgO3hC5LrAkR+nuPiUlj+kLC8k4htGK20cryqXoWIvCwuce1tNt83UDnThRca
lYkpZ9a5aVQb9rNQJgxOaeyQME4hJVVa0I1163BRmRGStusGAQCEu1/kpQnSDzZKHTVI6WG1dL6e
t4INJrGENHTA5VHDD6Jqe064x+iBBbqXNU5fn8EaxLcBnV4Uf54LwbGtN8eoyVhr7cTJSFaV+Uah
JKxWta5jwBY3r8FmoYt1yotghfMUb7H9BQ2SsMgXLv7BL+g9xd9gGQDILoHhnZmf93WstcicJHp5
AcpxPZyVrDR5xCG5MujWfPYBbkxbGkVrRI/DeJcxDx1RxOgNrXxF2mAUyzQTMCQYunORTYeWD3f4
tYdGajqgCmDVXM5NhWdIa3OQvbmEaHBi8i0XwR37Px59ClBhK2V0uoF9aBsDpCIDuEqdEyvIvoCp
+yoisqk9Fu7fRSmM+SbLAO045uaL+mes2cekwXR9oxWKvUGxYBPhyfcR8D7xcHmtNgQxhYJOhYjR
OyVibeW2lyK+L+4ESjbPgScoXtZKlRjPVgzx0yRxWxHrQ8ZLzCdpD/nHwm+E0Z5psbEYwh+HfI8p
B4FS7S/TBwpC6RnbHA4UpyZWfNYU2f8MTOvBXCUrRg4t8aEf8aog8qdX9jqRxDHKtu8UYsGeVHig
EGcUrHQY3UiQmqQq0gZp7VLfPumC18P8cZwPO9TzI/YQ2dNKDqGFKD4iUFiPseKKY29F2V+jDejn
T5w4y+uqM+FkDDVLrFhtOcBvNL117L8vOIULa9Eu/3k4uMxDOPHQ7VGQcT2Edj29Eq6V1SU8oUQe
zw7odbh0zm8/n2non4ebUcsRLkCpMA4p10GUJXSqCKvQVGDCTv814Kq4L7kdDs9SM+n0C2FLuY4p
KlPJgGDYQl426SISZmMEB6fdezRO/0AQPeks9q/EsYeYkygldQu/ZpVkOtwbY7KwAy+PkO/0FXyt
XfaoiNFurc4Lk0ZyrYaaymoW0dOL1hMNA/FvmcGYZYUG5kkLUNDQTnb6hGYxeSEdHgGCuc5+bm7r
OY0sVZWNqIHg8gAI4Nol1Z88rue9AfAOUJnPOOLgakx7j6Xd+knogWJkD5kIKF5P5I5XVw49v99g
ZmaCZdKLwwMnSNmklfFZ++huXw14Hn3FEePjPfpHZn+ca0Es9VwHdCSODRMGHTJVbyG5uXaUkumb
r9YbIWC8Qo+uXOq9tygQqCdNCGjGbobPvv3oODqsEzgVXnilYZbhORyEZfYsm69G96V6O/O4C6+/
m7jUx5vFn0Fn2NSGUN9PfO8FqzC5A99mBQV2Jgppg3reoegDzrkG5eymPY9A69O8C8BIbAiqEnXc
hZC56X+9fOahU5EsLfp9UxIgt2Pl7/wuRnZvRkFOIMHTJAiRP2q/VcZCwgxqUCHQGsi37/upQf8l
aSSFjok0xvoL4mh3+rs8t9ajPB0PZ7DAYmSTUUifDhHFiv6ZG//1/73qqBLydrFPmHZaJ2lxKS8I
3Y730xr5g1vHMVRWSMLeoinaTWbBLcIvKW1bWWNi17ldGZxxPaQuJC0ra8kxSbxDplzzBzS/KaIw
FH3OnAxdhXgu5Joy9m7/nQhAv7ltP250SIy4PYq3PNH44ryqGeP/1NFITENNml619+0QqzUiE0ds
KSd+4CXHbBp0hgX1nmLK7LSbGYuNwOh7H6uWwjuRtLMlLDJ+MPuNnfXlqryfJbm2YiT/UTSCfyio
wiarcrihUKLldYLSViI8ioX3p4jVJw4Y120byVuKJMQXeqOJLPp9ALY1xhZP7myCctvOZUZv2Rcj
oGn+yQbH8Wf86lgcfS1tRyZ1qCUX9nNMppqTOFQawtzLUKmdG2xTTs34DOanqfhKWzQUUSbkdVrs
2Iz+PKlsyu0D6mEoiDBaHapWmWhiFzP+cTlyxCK0tZJJFGyGDJr6BZ1JgjERuxW2sR/+OBuOwtFx
iCcSQw+lRQTJA3uO/7B9vHcEpFMWQkSwJ+wx9JMBLK3o5GnJEXT3tX1TVi8ovlm+fWnEBdXbBwyr
3NB3gNUGqH52tkYtXp3BTTYo350CgWeK80CO4gC4dto0skTfHXswYTVl7Al0wxm6yPOfQMk8zsSx
uC4DYGKWZmCbBhU9UG8Wix8NpzRjjMI4slGEV66pnHIjJJopX1WsAT0kU16p8vTh8AFRhr05GML7
IM11dcBAP3ha2o0vXA08C4Oy6kAqsS/N1DIIhdWeR3JpGC50E/uEsMMei+J7ZOar0xhQ04ma5xsK
Rzc2tXCohXuSC5zDEjwuWREO2kRu0eztOQ7Q4L02DHuuZpMij2AoApkd1Am2CE30GD0ju1+LNYS8
GasfrYAt2fx/QezbCNiYXlt30iUHU/J7ZE+HxmS/WeRDD7Z9WEvl/7IEjjwal0t21glQfhWNfvq1
o86bR4l/VGop14blgyTL9wQweDM/hK9XVviK7i4oK1IryhaqHbm0iyy23+LFJoBleDI4CoZpyB6I
p7/GkETwrEQczsCEe+J9nqL2t8c2N+4jdkLbM2xqnubr6qHpBdNfaGgvy6nWLRWtj/KoZKeKcb8d
jZujLmhSlaXJFN1cvfuvxqOEL1cwB7RPsMq0iNZE986OAcSGFnAS0IIOIkvbEPp6ROm/u5mrTFpG
N/f2iSC4r2F6vYwxViH21+Fwy6C4JuiS3b/dFE2feOv7V/Sf9fLYP5+JyeCBXoqLjqcpaQbIVYF5
MDcFVyGmgmT3zghqB7yjXpcufIb/TMoGRTkUwDNTqGkYhdXzJv/Suynq8MxHVngjPPq0fukubPJJ
mfTBawyDcn5nPeAeWH1QkgVKvlir374r2dob3gqGzRVKHMgqnXmsAeKA51bvFcXTrAmMHr90vFBt
O+CerhllHUzJL2Za0hU0qqHXDirHpFDCyrT6M3s3GqPZryFryK092wcDu0LzGP+TGpYGiR/OtzHE
O6HCZWMVqLN5pmCXTWKQ0cWp/SLVgYPK9UYjc0dQx3svgTnjxbPbbuRltvULP4q41N9zuaUAxolU
MrSF1RIatro1NxNbRybW4ieDz8kir22tZTqAqx1CQeZwj6vnjwMGe+Ghn2UxdCbyfR/r7C7M8z0+
vg6Pq6ctoVuvInGdbUafmTRZl35llLIcAp7QVefq5BWXNUhfgG/H7vMhbdZYqkca5mC7yxKmvGwx
YzSA5wNAtN7iEMntPjq+S6vu3eZQT24B/lsLaIqYIyQN5YRolFbbj4Zn0ZLhQYXpqh+nr60kvIXD
1lUiYEXYgXTO8VS1pPVWFyYl7gh7VBwgNoEk0fiLbP3pAOz9ooX6T/dyWI4uHFrxnixgFsDHq2ov
0Pw8qwzX4r+KpIWfK2B3nFgfPCj7viAjbGV5uHTleCQyMzMIBx0KfQf6xg35XJ1RYg/WNMM349kl
KUEKx6sS9xJnpwdWsugA9QKAtBXrEv3g6+FN76KfWfd/T2nPu7rc9kmyQ+3ywvFCVgH2xTHN2G9W
mVEbDYPNkMTpNEaLgdIDreP8EQ19h/kI3ZZuKlwtbPgG54L6ky36okzPbTF9up9E7ud8/PSJuOPL
VKdOdEtPVxB6JSlQm/l+b0+YrdufkDVoVqIVnvCwl9AkbNkTCSaJAxGoEWMC00FlbybMzvSDg5Ro
LltdSppXfmWEgwFYqONg3qoZHMx0tVlxSeDNMHIciEY17+SRzmOxsRWCT8DN2/yuMZYLwGdEGm3F
bSc4CVHOu5sT0vOuzRRYjf8yhiiBnlVmn9jeZQ6Bd8rxM4n8AcKJlrkhsRoQVJRceniehmCUCMi5
kjuW40M26Bb8CmhS/qSnxbhjbehG3vL8EaK+95icITt5Eb3mV0y0vb6P9Igua3lfI/lZVb1lIh4z
Vn3zfNlNB8qrBpoJ3f1be6vyPpDbSlO8B9Pgu5aJ6/20EYjf1QHY68LrUbZDM+Dc/3FifLklShM/
hhZsbaLlOK3oMQ80v8u3Cs/RepZ5LgqKfskbwB2VJALJMYcHdJ7srNmErBjVgspMwkAOAnAZytGz
zD4qbUFvnzxBnRwHOT3Eh5AYwdLErONhoGa6tcBdoEeknPHTlxsYoNEUWEs29sm3nbHnGXkQf1UG
EpkyRrUykOUaLOhh9lFg5+F7uH1Ef1byZbEid7Ocu/KQLX4MxYgMz6omKPDSqMAAeErQKUJ6TmHj
BDhJ9gWWvOmBiFut8JvqjryZYoRY3cUlN2KUdW9Itwg2Hl4iZPimtEIhJkXIeYTBqpFAc3x5+BBA
1vjQ1EFFZktWFVvMtNQlBhaa0EktytLykBv1MxaOhUI9z7oWZIxrHUNPqqD3dobp4qdimPh+v2Bz
Lkx5SQrK9SsT+oPg4NqCiEuawp8l+4xERZPfvT3orve2jFLhRwv5bezBHVlomQsYasqsI5i995Er
O7dewkkYnLiCsfNq9vsz6PSeUm8IOkmYpiVJX97cUWxs5wnJPxpThRrdJjFldoFlNm3p4Xh6jur9
Xf/oR2OUFM0s5vL/gYvdOVjwtFsR7wJzQlWbKxZyyccVxBUlvNuHAaxsYElrkRkuIsrjH9jLFq1E
56Km/Qd4pp3cCrGArJ4VrXZvxQ5oc6HS7s7eFb4ZKr30O3cvKKdXiTXk5h1Dc8AKGuVC3lnS33vu
VPRNzqYKzboLCJg/x/sHjANMY7NNaP2k04w1aLCz/UnMxHV20WlMa8Hyqh0FoVw3VQYuUwX7AyaJ
6iyhVGzp6D3XUmwV9KUgmugPGPYilsPh+J1ciCbLheP5KeJ/BbUany7E/GgrK1ezgia5aZVJQGNM
i4guZhmTZwKca7hFlv7S5UZuV2CNvAT+WU1jH1i94f4diDyk0LSAmAl1999QhbE4XSEN2At7o/qG
6+cHYCdqIPNpBmKUgxq0jnCdka5+WdLU0ym9DoxJf4VjFpIaUo737ppbZSg807IFnZLB+KohhyWV
0v8a8As3jQ4bcS16Jc26gHeN8whNtW37YzyjK/BqHvfk+3mCXVOG+oCKVZJWi1kVYXE39mR3FLCM
1aLMXhHA0wI9OSOyU+VP086Wx2hhA0/suH76h/tAvE5bdVuUjX9uj5HzF6t10J6RojCTt+F/22TW
6ccJXRrdzisYTZ01bS3puYsvvgR/NdLEAwsVHMlqxLeHbFepVzBnIa9eXmZ0vx/yG9zTsGy/hhYJ
ot2vZMZ8cVeJ52aEeKEJkEk5pEc5Xv7ODkl1Cqbzdzk8kNAgYntHTRMqO4/VNk0nNGBToyBPI474
wDlibe1bOv3bTRVguNORme5WOPtTbQz5wZMt5KaWboRQM0/URKojX0oyk7UMd/cjZ15+J9B0tDKY
HS/jtZ3aCfbkh4kjgonm1LzbyjTr90FMJHaa7oGb6HzMj41FURh04CCqjcrAju0/GYUTn7ZWSuEy
lXjGV2XIlgvWH0BlDwiR3l6uMtWeKkFog3nWvwG0Ga7bW7aAcTaKJKzBx6cBaAy9tr8Hq7ZME3Lo
fWhGkOB1FbYan3y5t2QFgjtLR2qCDICYEBWNyJb5A5NrCzhN/bB61KtFgHLbbPWST8SUNcOUEPe4
8yXS5OQJGe71UzalTVt7oBR61gZTcjFLDWwsYixKcSlJM8Zn9LS7nl3yhVDVBfAAYiNFOgL12cgp
UznxtcallaqfKx/i7dHVGMGASCwtHSRsBACUoM7TAvkqtR+W6pee0dF1hH8JCXOGYQi3sZHnksOn
/6LX1bT+fo5ZwPrG9UyniBEMiJctFWq2vytVk5HLXS/Mx6NCRyZGJ87x3pL6z0P5rY7AStVAS3oa
ScbmTW+xPygb0CTBnZjXE9wkGmLUWJ9gnVOVK0aaM7IrqnoFLQzKaVKwdulJWZPCulkDJE2Trdnq
nwJ6PF91lhQVVTS3PCk+FglZmD2SVNdgAaoUkoEDi0Qspg6k2IOMGt6zLvNFQiuW13f/LpXqbalp
2qxbqG+pNOiwW5OAIHXjdJ1957DZuR6u9lhJKOZ2BmYi1gK5BKt70T+iOrdvFX2/SiIBlHKxGNxu
3nvZ+dOPKp3ThUFFZ867zQHM48k/beFWxab3PGV9YzfCz4uni0VfBnm76QFlDJCklV+jyLsKBqX/
j3lTUnjz+WPep7c645tPD48OzwqRCd5O2QtPtFLY6DY1MtvtHqAQTFbvzc1k3P1c1IXZDZrIXIOD
akC1TluJZ79uWUJ6iUYTf0Am84ewHSVwzmdJAS6mheRAdHoB0LHZjNTgoKtWLvy+GxaEb8XWSyZv
Mn6PSudxlW+YH5Hr4CuC+6KC9pPGHKm8EoQqKZZhkmqNTppv+FUNyZTCbhprOiDwqL1/N3K9Y2NQ
r24Vs0xtG7l8uQcVu5shP6lr1UCFb0Nft1WChHoR0wMnjdmTuwdYvBnKTGXzldiBf6kMlfUrkssA
n70BUjJKnwWfZDRghy2nhS7MC/xRHIsHSakLkCoV2ykjLZP77hMEroSHstleUUs86Ff5vJuAeYjA
gPJI3X0iNFAxGk3I7FzCUqecT89ykE+9+6BscyjCGl0bwhIWTVOUN2vWK8wLcn1er5oMCK573xXd
dqKXrTwMeWOLlCA0tm4Qrt7hQ6acxZYIbyPor9RIhuEY1J2jGj3c2lLF5CtQhdcpd0nIevaP+EwD
hQgUARgvmMOnuaCI/HrD0i9akkNPkCjDN7hxYXAHFHyKYv9Rzh+NZR3vftIpNubDkwBvgm0P1eV7
ugISxUL9+Wu0aiOeyorZrY/nGRGlgxwPHoF8kdxLADUdHRmhyJXnTZWxnifw/6Yrlsy4z5HSNEFb
cvJQDoVbQ04PPY31tIP/2pN0ljMiLANb0GB6c43i2x6ewr9Etz4oBqrVleKYB8yGhudQKHytJ7Ii
XgF7iu79IC6ke5m3EonTVgkgCNuT944MKpA1l3sgwtvWcWpJFhKt8fHYBGF+gtgSEdykqBLvGUfV
76qMcwAD48YVIdv1t+z3iDInahNoPixlegQRNHGiUrdIK7paXWtQ7PAwK4O/lvssDZy6TJyzcCo9
5vIJ6TAMgnBzuMUZdyyLvYbobUECpC+TkFf5ixYeqh79Kzq1Z9/TtCpN49dFIMmU/1KQT50DH+m1
WM6zwKf71l+vuLxZWKV6ALUHU7GY5cxMWLJr8DuMkzzR/XArVzzNnljmuATxXtR41saSURDkc/xg
s743XhQk1J6x4UfEiyWqXklMeomCqwAzQ7YxrJaZxDqDzaAlKZYk8Xh6olpxRP0we793G2gHcgut
x5cQvGXV2je8IjrdesrnDeWIfeyQ/h9Iq2pq9+BvgXH+k9fTjfoOPN1vUxNk31HR3AkrT4ex9j72
c0TQtx4amiZLl5bt4Z7jxrLGzvl5sPgJQf6pajDSQ7cTEE8IDrniv6I0ppbFc1yQHU/LOzymZ3m9
fUwUHUlNIZyTLrplpY2L+qOSk7FgFKbM7p+kw0zNTMCwAlqlFQ3o+Z5iHCFYrdpQvuDZQdiZ+etn
7i+6L/8mHBDnXj54ikBtgT9gUqQZtotDXxuIB4JC401cSEU8jQyBdKVkS0pEydPBZJWDtirWlEOJ
kUzIDJshzDWLa6q43AcMBUzVkNnQQF2L7mddC3VamkIbIDFx11QXYYBfTAqB1OTNzq4wWnkUE6e3
FDGbVSULiuYCpvHE3LPFb6VXzw8DS34qjL9RdAMpxQMlga32v8eyNUBlxHIH4+wyDfy0cmGOu/q5
Xu9wf5k6PyJ2ICxvZl9l0n9/q6enP/C7aEpT5rfg1j12doMQKFUwSfhV5j6tnuFLiaGR2dyWvUF9
vgb2rLBKAfCYdQ8fAHbHjsJFcldSNPckAvzr0jGhz1rShjLJN/nhXDn7mfOAj2FybnHTR84LtdsQ
2Fxe6s6oL9xpTUEaht8xLRf+snXIuq7HmkZl50fTxZ8PLfWfb895htC3ulp1BL6bahVyKU5Rif85
ZWBIkNcn2Hp4RzuFjrFF2Rd2LTztmIcDNinPG5/LjUyj0vzSs6KhaCO5TRSVlOWd1Gl5kTVtr3qg
8KMANlzNn8O1jBjT0jPQtdedQfC33UfWfR2IjskfPj5Y+mld+Mk4w636PYsK5OkTFpz4LtS9fVr/
0WtJt5eXp3n0FMjSmayzaUoZTYxehxyi7d4GSl6esRUnfx/wXV8IjTbEPi6j3U2IPXSDE7DzYQ8d
ARfE6QX39LRRZETpPWfGv0ox58etWnYVR51fvWouRY/JuF7G4K6gx39f88GiirxlqEJJW0BCywWT
FbQLuwxWn04Z23dRl/Y65hDv2XC2iYlL3E1EQV2uzrAyVGbUWo4Qr0tRPoM+ZHANV2ZpEC8pwh4e
ewBLBJAtxpxXfnQvrOUdUQPieZi9ySkLiToDrRHoDHZ4aZuq1kQBr343FoLdtCVL/orQbIMcY96R
kG/FDYwyL58gMu0BSD4EdNUrZK+3E5ZTDVko6yW/mzft/uDlvn51UItPB0ffXnIasldzOnsonxhu
2D7Mm7yH7m6a8g/jV1/yLEqDw5dvowsGGTcr1fL6RY/SVf2hsFBu45CNUxr3X64WMDshfJsOY96A
iAP2dGU9ERXBDnM2dumsOfXQNVA/aTgQjFf02J8bwO7it9Z3PsvZcFJRA3lSvqdr+u5/aScnOqp9
K/xJPG1RFCLTcItqYXdImNWArRPWSE3GOTZPAw9gX5PnChowr3HdCrZamSifcp6IDJc2IOxz4z65
U8zukPkKRQJnu8Sv360CBQwW3NTVTXE5T4OGo/z+5dS3KB2drufiJhxZ2sylPJwQ+vv3LtEu6YVx
UjIg96D4j6voI1gxr0ubrZf4zKbzHHBehSe0B958Npl7FYVGL8ZH+N+qk7akkaUtkJ2zzmf2UY8l
oow5QDjoWacibP7zLg87rwowEARLaeJXHWAJ8PF4TtQ7Z/cFklc2CfKfmDYjhOtQrqfUz0C0hyU+
znhzSIGI792Fko7OtIuEkpR3R3tUwaTCXvQ5WSZDe0duFlzJ8qEQL4+CyECtCaB+PDltMSdPweUb
FdebUDHNjyku9mfKp2yYrU8dmFSAUpUjOuqE8qBS0wnTGkupgvWZGOJpvD2zzgXJ+Sux30QJr7ky
wOe1RRsTYDi/1dD4FYXAKFmlaqrcynNsiru04ypp+QJBPQUO4fModuq0bvc6ZN5OzLINtNrO/SsW
4J518042kDp3oGG+9IzppuWIph0GlA9nEcYbtFs23Soqt/OLbTtpWmmWGMguNqDc796f2cCFQOZo
fHS2h/FkHJ/j3NDphG8+9vxvAjHf+Q7bEwCB2DpFmaSjRvWAzEIkv44+vXimxkWcFiXO9sI3Sg0k
V0dKuAQ0/dk14phHKxmLIxCr/SNdj/i41clyXnjqJdANKfDXcLhv/Fc1CRRszj4GVJBKOiyBOZyf
i2m9M/xje0AHv4jrAQB3gXS9tBIOGbq/c84r7SQBo08xGvBjzF4KcKp31/Qmmo2f3cbM/P7UjbRR
MB5LxELuV+fgiZ0gKR9Tud463kQJpDS0PHLUicfPZf1jObG0dAZKQza4zD2JMFEs0shbzXBvebdZ
28bbUJIKpcebmixJzEvSnha+SjlpPjmBEYBLAXlMw4F5p80apVS5hFXfX0va6EMJ3NHzD7FPOd+h
UM5m0UqINAUOQfDjKMHNKkwjQNQjPBxOe8cqCrrdx972EMVNRfVis6JPt3nCA838TNZiR5t2Fw1/
9liLyJ3vjW2A+ppFK6Lnys2IVLU3Gr6vC8mSERTg2777qvF0WU0XZj9la5cq6uvlUNgYo+3+swlu
8D1aJdBMiUmlqDRl7/a5izxTAruPpj5U6T/I27LqnQxwWckQma20wEMrwnAcQrNdJuwDTqSsV7gj
69QmKQxiZgrvpL1e/JSwmB2zHYNoBdOhcWD1p6NLbWv3s8kvOp5Gq5ICt6aWvmtu3dl2InIj8fnP
pMCUKfnszdg17xafNIVyo1OBxX2TRYyixuG6rkNycSz1r5cupbZBW5hCKwkQywhvo8+HqAA64MAv
LTmlHoJ2rcliSoaVwKfoTXJM1c+e2zypM18Xk07YlNghaYvTAxivZvBO5pN0FTLrmkt8Vgf1a2j2
RJvQE9lDFO0g+shnXNwAZQfoV8eVZqWisK7BLqTwoCCUoM5yoKqzjmvzKg4Km0lMUh8MO0qLo2hK
fWMmbDZUnP6lRuMO+SI/uPSiNdvDi1xqAC/xJ3gOVj3MClJhgHdAJaPHVFKaXiphTpPZICQRcFph
MbXQ/BxVQTYzPBYzwZA4RT+MrXjLCZzvpfWSBTcfyMj7xZKL2i3EOKC3A+g8RclJMAbJEMUz7swy
JCl8Rewti7WtcykWGVNNGL0q2BWinGCSkSerWNOXAd59f3RBT0ZqwdThqbH3Y03dHJZIO6qE0Rhh
kEuRJCkmsrxN1fcKil3IavhqM3k/auWSrJdNCu36KzUAssCdOdjZ0dI6NBXShWdKLOJurI9RyVFP
nKiKgXvtcIE5c5N0n9cpnMedj3OeWh2O7dkcirRdl5IzvMNOJO7lp0gXussEGCMd9xrCkXWZh0IZ
7Lg97dXh8c2QhMKeadptnDugXkvRHoYv8m8BbWb9TXXiStNH2W0tZ4zqhtguQYDQHw/7akwCoxqd
bU8zKL4iYcgJjKhbCRtNWepgpkYL4kvUqXVle2FUT6MdOZ9ar0e3o79xIiLhO91AysSjiWjFi6Pi
X1JihO86VMBJ4wdno1K7J/Dz7t4QVSRffGAQ9pszQaE1vT8mmC8c4w2WtSisqs6EXXI4ZPsJi3Ih
aA7ERbz45fG6M45aOtE08QOfnK/3tK/B30nGhPse1XrW6va4d0czHcRRPU4MF7lL+MF9LOtDxXva
xT0EjaNRFgHKkvdeNUT3miD4awGv7g6TiM6ZW9Mj9FrmFyo6yGmFWKOlEINx/isyRtSz6PqNNwSK
TTaDN1G+pZAc6PqIx/IIZwb5+klae+j1/IkPKUvxo1PVXv9i6IAahz3eaKtGBV4TkLtZtVkZuOOp
P47JDMWYw6g1U0/rO5RTbMhZjsuMgTz1c5xdFVcg00+EvevURzBois1CMnO39GiWqgBPQj158RIG
hLt5yfzPKMPZH2X31tVmXwIEAtDrO93sZo+G+SQdtTNF3ijtDcN6Q/c0Ntdpa/PcNdfHEELmqykt
wWqDpkbIiqFAOK+tloy8MSuTkU2YhgeV0JOSeCz0YubmG5hbrEfx2KZw26HNuZTFLlWzLYVyjTrE
PTzu3VX2fbaPwM9ItwOTtqVXWkQ9J2MAV0IAgtF0Mf/YLIC0jLJHFJ+7Hc0HC11y7QD7HbrOnzQp
Cm0C/t9qIBDyzHJLhMUPMVA7nDbb3xDRxBXSqr8f7GhQGam4uTPqVJC5PaXu5frXHZpm9W7iKMp5
1nJwNFhGd0kORt9duQhVsqFuT0GZye4fszRL+DkNvLhe1mFuaMQmumKaH3JBBnWgtj+4qdV/ZWpA
K5N3pCAdtchc9Ikxhgt+xLjFCDM9hpNh5R6DnOjjgBwx5z+IdGhSDzPqddn30y4ZlbEZOWU/o/W6
I9ofBQKQEP0Hq3eabWEziUvVJiunPCUFZF+Gc7RubjCnucjE67ofDHyqVzxWeYyEgsYFPL+obn1v
vwDmIUlyMQ785ektfl1GJUhNjS3RjqBW+5AcP6J5bo3hNVKpa152rE9V+7WS6tROZjo3qZZbXG1G
Bby83CMX7E8wmclXyE8oMsNVu4kHOpl8kduC6ZR7Jx9+fF8Cj5wj6srjQhBaR/h3fKnKkXxBvjnV
cZVndpjfK94sh1yrquvEwkHj8GpVSDRVuNyNompV0rYeUTZetxeSeReADtFaG5UleD5MClmt4AIC
fq59uctHawCMuvfFBPaN+Do3u3QlUGSHmme9ytIheo8KDV0UVGILSDEn/hw2b0+kSgprpDrEvkyN
5yY4FhrOn/Ti7plvvEKU7mgXO1BmvjmgfWc/TNLQ+D9FPFhwMjCNkT1VMn1sV2BmfcshJoKXjejD
pkrc3sOJqzWavRm1ZZnd71rnpboTtL4SmcsSHZgqL9NocIjCutKWUYMe27Mys00s11mPGnqbH2fq
L+svHJ7v4oLnIL3hZp6X0x4XpTIqCWoVZc2g7EhQaJoNdCqtD06bktD1Zk167iAXeCDSJLFvb2Sj
8rFNKmJAuyFj0AOu+ZzFM2uXoqN9M7EQFJMCwMPYva7kTlvvRYrwNXmEZ7WsBsZORJPfPeQMS234
Uz2EtxIGNmufrmHY3oHHXjdE6GLyIwLXOwX8dGdiVph319J+8Y9zfYzs7pZcVg8kRpjvetNkXR5R
d7SMla0z19dg2Sds5JagryL2qwVh4lvNmf1Fg5rYEBGDvgh1+DjOX7xLaISrXDFhMFqLNNzJL37T
wxJrJ9nB7jgmC42Deo5k+aT8e/DUei5VMd531Ipr4NOL/iusEoceuaJg5PrByrHvXl8p1Hvpikv4
v1PB+V8YbaJnmr1EyZEmxMu5/wbmVCex3MV1qU8vaikVGD3+892ODL9TQfoLL7eO4IiEbKPzwT5i
f/EXFGFrxS36PdtddXv8bO6DjYZs8AtshUB2Dz5Rw8l9zNsb8aOdmESgky9QohOExYYZy+8xWDDm
Wlf60kl+d31/cQpVBghjc/OgwVI+oPWJ2yE9la5vTIwqZgF8/dUUkFq1IbzyIsh2ejUFQwrBj7vC
0Lvm61g9IjfeypfFo2RFAd0E/zo19BDq1Lcfffdo26++jdfM3dQdZFHY/8Nt1RwsOZP6LJqUm9yg
xmtPctYN0V7m3eGRbUTCbFk82C+RmAOw/Z5Fct8vhm1hr4zpZ+jGBZ3CJihD0sAm5+xoxrv9pSBK
kbysJchrfdMn9p4iVHsegd2EtmRuFwY5Ji5C9t9GWN0vLWx7cEni22pVgjCvcfr8eZaJMfCkAmYZ
swnXvNPLjy7Axxn4ZePorVMsyvFaDPpeKP0lvsLs9PZelaG9GVeVo/MV8z/Aj0Efvsy0b/Of6RFT
E+ytGnxxz0z90WZsA7PEF5XdfIl3mPLjMQDfz6Al7wjqLuur0+9O/AQuDtYl86WwtxK42TgtF3tr
IuTL+VTeUeEBclQMQpliUXJbYb3sKnHhDD0/4bWt4/fqMJkvws0bw3yjFPaRXBmU5xLhqwPt5YB3
zPKh2lyZfTzot1qCM9aocUWw+h+0nU+wTOFRnNfISgxtL7mnEsKJf4o7qheDIJKvvFTKPOFHB1Gf
ysf2KryKI52beEEsfRsDwjcMY4EBe0/HJEvSy0QG+4XcppQs2uyTPeS5GdnpC/CdRfMGJ4yLFjxO
Wlf2m71dwYkSn9tsktqntq0gNWmDffVJgcNpeVSsCfu5IxE4oAATwvgLLBO2HDMrSUtJ8jE+7uJF
LRHYTw1oyQFi0qrliIm/3FLWisppaCov/9Ic+gDTTmSDQYxdpeAZBmKM0zq4vE2vkIab1PqHM9j3
CBfM+OtSBmeIRRqqZRz15G2r52s5m1QeMv3s+L9xO/JFoz0hRuQislGvBz2qpqF5CBrw9Dx5Gpos
PNqvyvbfE6Ojo4JsiCi1SOoBY1s1QX4Vc+5xtISrFipBXnShHeFfW5BPuSYBFaZiNOq6i/gonQD0
SAlWd8mPeDUbtCYlugNhIDeY/yLOL8WvDGzmfE/rkvx1xh999n82gYXVMLl9SL+lLx5/4JmIlWcn
lT1x3kYA3XLS1G2p5gj/IHS+oZ9A51rfDoVWnP5r+AbUUOE0GnmKFWBa6MLlW33M81kJQ8+G1Jmz
hK7BX1z5nqJw8351bL7+nbibP7ot8XwgvwpJO5IVFZ1sCeSa6KsVC1U9vXWmVkluG7kDxKzEzFM6
STR5CjT38Lrz3EM4L3nXvt/59YffPATE85gCGZYMjOrBxmhOe59ZWV2xz+OzJETMKFTOPytusF3R
7XvyG0MECzJfKfqjU3QNMBY3hrv/3MAJndo5NB9cXTSXMVbUCBIN6RP6QpL+3S5iVvYiHIVRzg/V
mCHKJuPFN5kk9KLp9144Ll3GDaoT4v8xHWHJiU31tOfgxaTV0xlcZrqlN+2NJAJmMCr3SEOP9Trv
zXE5Z6g0NphViYxo1jK89pFgwzAEVP95X1xqjM4wLjIfJMRYxo91H6tbQNe44QRPaha7Vfmljwdb
h24TfwgQ4o2bXd1GrsnBK1bUceAXtXZLH+Pc9OE3SFKKonOb7l7YRGqeGYGXYVgPtqA/5/MNCBbD
ZSuN1kRSlgnIYRT16JRE9jxZVY22hMK/OwNjfOoM96QDaVQDAVpKdu/MKBNrMCpcdNkDer52JH4u
rwApcB/P4Zz7leNRLLg+c2yNSR1LUrn+czl59dg/+6ZBKUs/UPcm8RXdTAkVx8mxZPJIBENviRJy
jCbCQUd0PAw+N+NN20S4a5mOEQyJvgimOppUjMKV1qriDseg87ZEyzkjJ7m+Z4gWdDScpjtAI10x
9Isf0j6MmVCUDY3E4lurOrTzGKol9YDe+yghNjLIDF68XOcA48pwy1PhYv4xbGUFMECOk8nD6y+J
vfg3OVR2Qc52blcn4UpKmWFCu02B0t9LLx8HN2J+S+wpduXePCO0sAqjf4rLgyH/Q1F0F1nu8i3r
ALvDScg+97WpMuS2A6746dRzpbMfpcRYOObMdKNEPzl5RzYv9wYH85NKbOQ5rWeZlsi8vR18ZYYb
TfUgJM9n0a85l16xrMIs65ZuW8Dc1yXxti3L0X61fdLTgbBKP/sOH+w5GVZ/zYxhT5elW5CP00uB
O8gYH74XF2PRHxdvmEkpgcURR8YrqVESBMD/EHd+MmQdpI3tthB9LDfGmDeuepfVKxK6U9NUceIF
Tof4yBF2qsL/34SREzJlu5TA5iJ3Yp7Sm+4+pR2siJ1oXRDNbn/w/zUCxczHOsNjyuZR0wOjHZtE
FneWpfoh1Z1du3MTRa9FZ1abKBDyHtqrPWfi9KfRsakl6u2KlDcsLUJt3EZSHiJQQLZQIJm+kfpd
HR2svuOcN2truWfG4UGs29HUZWl6XkEMgQSJ3iznN47B2IrUc+7Ya0npe4MdJ+3bS1wZM/6X3xVo
xwXQr3cq4o1j/1W2t/Jt9nM9ZpMZjECbX9QdaRQNdcIWsUtN9Fo0uNE1wh3xy3OM2dPX9MEdQsx0
HIZzmwTTF5pWVREiWUR4Qu7Yb+EtNQw8aVyiloh8bfowBUEmR0N3xItqisiRrCHJu0lDw1FsF19i
Mqtjq+Qfsg8lU6xZtU1sbBhPkiBprbVwtGgMH6zoQAVIgFZ0Hdu9WbGumCbX6TZPKBNHnEIiFvzG
p/k2kZuof/V62bjmY6Ahs14I+x1uaMylbRBu4FTwzItrMrnotBXzzJGOFt5vcl7uskcIq72T6tz+
dD5UUpN9eCuiyCdlS4IBAGP1/FS571Kk2N11dttTWZErtbW35bEPzkqh0vp1TOU7OfLfAYjwBwt4
aFe60jrUl3wTKA2DIVlw/ErE/KC2jHp7Ob/cGW5t1XFi5tnya9cDIGwRrF+zfCwkoAfSCwYnPzAn
b2rplvIYMwE2iLMoeuZhCFhkgICV11GJPCglQ7GbAKQe3rAF1cHa/VjR4GzbmspGz6tjEL+KWcNP
s/tNbUpj8JWmL/kbUfxUKRv7W0XAEZ+ozYyaW0wXtFAek5/drHY0a6uY40ktNo+QhB109JcZM8g1
Lo22hpbO2M2KmUk3dVndSea8NEBVmPv7TykwvXBgw2FuUBcjzdx2Q6jtE7JnAEIOa+MoSX733UOB
A+77ZdH1jqLA3oDzW/EU5fkmtziDdNXjoLTiZ3XDZBHhkhHYYR4UZ4uB2hVvTFA6FHxLK+WU9K4/
0TmXFv9cEaxdGeG3JaktLI5AW+flxZNLWzDQouSq8d+9HuFh+Jz80dpSgjZWzFhotQmx0qhblPzi
1raX5m+7O1o1AtbJHdRC3sKfDvTIzk/GUN+k0RY49Gn+Bsk/QpmYnn4kEThDOlZnUCAILSXlDWFM
8aemHjjuBKCYo2oeqBxXsMSBzGb6AKRGldXdDN7cyOzzCtj8gKd9TbQwTEKxWXUuKvdrNql21edb
aq1iT8MAndTbCrVwgReI+Dj2byd1IzaHLqB3Ixms9AKSRIOHbC5TrWL4zYAo18jXrKjfsaiP+0wH
3afMGETXVf2mWAgFbfN/dvRizDDLFou3xPrM4+GD4tiOze5LFKy7Kir0lWsDR5xjH1q6C89QjIz9
TvMYMV1/LcDcxUBV6XbE9zrv0G6Ez5euPLtFIERbP6ec2roNFBX7v4GAlpiOYZkyQiL4OuGR5ZAB
4W9Ou+RE1J40JC6Z3iC8nnRE+OS3C+YAEc8NeFVlDpoQjG5Go7JuBWBxGI/jel+RE6MyYhg/pqjo
XI3ddt7xemkIp4JMDK8aR2MInQqvGIe04vfi6B7/BWbAXNym1Qedm6R1X/o5PE7uQ2ULzCOe+a4d
QoH4/ASwQxNOngvw+KmfppaD7PtVEpRie/UgLQTKmMAV2AtQWwZfSZj+yOAS0U8ZPXUoCceC9RSW
RkrwwlBM94ETj5iS1cc/ioRr7DGH17mC8/BtDg+UXkoXPdaJMnXnJTHbXhqQA6JBy8tIBjw1LmpY
tnyuD8cXK1aPu1IxtwOnqE4KbQA0HQv9Wn7QuwjB/WLsRIHfKrysSELbKMS+OOFx1OgNWCnwdAZL
O2wGOIqFRdj+wUdIf+/xJ9VACPg0gcmXeinE/cpEnU2Ch9iNqiPXcWOt0OAvdPAaxRnWpX1LCUl4
B2YxZF/cZuaCFcXI3yjJyHKxulabOoOgqfnob8hxrl4fAjtJ8RSrRc5ypyKnC0HMopGDFEsQp8JB
81iwTyoOioO3DaxsoQqtsFKwUlplOhbpVHTSnS9fa/K9DbbQYfTjOlzxs7++Lg+EmLlYPQjqDSOA
jTFUeWh9v7SMF9tVTvayv83eBdhAO+7PvyuRUrCQePGXstIzrRHvR+ESD5VOutCseQdPtbGuqcmN
uQDtG4DgZ9jsKA5cIOOJk6Ekq8ac1J+dnB1YH8x7cZq7QnHcoSYeWznOl3qDcTZxoq0guoaiLS4u
sRueaLOT1LYodHx6ndKqerucPZIcc5Lya0/LXwZkaCHF3zJWCmfnNPZL1l0A5SfpnHz8EtTQqfvA
ZiLpXFSXYG9ae6OGiroiIwynhhsvdquAFhJ74i7HaALpqKMQif34wiuvGpC2Tu9RqG/1TEu5zxmW
evtDF5Ur+GaPUqrINtUU56sTa6HbtJ080I/Canm5qouHDYCQB2mdojnFba6IUOnkpF9RV8GXBenc
YRAyFUpJ8y6ySlrjK+ndGwWEyg7PmNp/+wDzY3wr5WYAnWn68vqzbeHQYoNQmutaJofBTayBdiY6
NO0lbcvSy5ZMCactbL4cG6tVa32Tcad8DilRiXdmBZhlMV7V2+ad71Se0sbb1Tdd4D4llvhnPf8M
ytW0AUN736OUU7mev29eYOi4sP0mFDIfLUjPY0jBzEXFRgy3lCmdBNGjylRpzNDTHU4qp0/yftjv
rOv+PbdHfeLmWDoOqRwT+Xfuj+vOPtnlM0J97JwufOe/E05F8+DY73iIKHknZXPcRfjBcbb0qHG7
hSmYoGsGDDsA+HK++FKylRp7CeXMIVOjdt4hfP5qccJ5VTLPw7WcFAfMGNuwpUUQf9tgoOsTfT56
D9Ze+M5MixiHPNqUg1iCzKu4EDOu8JYAsIb2jbwZ2BF1M8+2X+0U2em2FCxf5zxLXCSyIHrMX09p
yUxl6Ia7udYWXJg33219rSRnDjo9xQrzfqSAUyQHbrpko+ue/LZRfp4HwJRLLP5lf0nBO8JAKe3o
ET6eMEp/YCGXy2H6/m70ejD2xH8pb8sBBR+xZQCtgf7oaRg5xtWoeF2kXzvDzIZ7NGXauNwUc8UE
1+eydS86qtjpr/hUW0xqEs6yBXgfaWWnpS3mNjGwN1ENqwXYqc7lTRRUs8+Y3aNfDo7WLxawYil2
XM7lvYaRrIY1D3OpykvCroSKrBimmJZQfgHpy2AjgrymDhfmiuu6lEP6RtmUN06lOt1AqLjBHrsj
n4f5dL1lAyaWIZz3vE40XOFXf+nXib3BBH1UuHFIm5AOvCMxHtP83kZ5gKqHfaA4gxwsaeVaR13y
NTc+0XWOgPK8fKeBm4ofACaiAN3QGsyum3dJSEoY+WFNfjTSinIjKGKtbCbqOOmQkl2yOS/ul2CU
gBHrJpBFbkMeTrXZ+O6DiNnlfWYu4IwHZwrGQs2N/4eBzwoWr0MtB2XZw/+TcYdZyD7ekDf+Ybmr
kDdgYrKtKA8dDlJYoq81Wy/MTUybhAZKvvyKwT+LYBf4U/DEnVXUCuUzkS3ru/8oBqmaqNf21sW7
41ohAYGwgJcMu6Wppg5lCZFA59KdS2VT9j2w+npeTeco44erqdV5JAJVwtk5MhEuuFSldgeE6OW1
/hs8nMr8Z2NNI7ndPqH40o/S0MWZ9OCxQOX7jyqdZd3fbs/RG8rGKGEHIbKpxKMJVfEvefQhYFoQ
+lmRJBg2En2by46FlLXHEsZcGbkZp/T5wCeVnvUN4TqHQ2C42hLJXyTADOtsuTqT9JCgGV1wilHa
N91t+XhYY4AtGtKkneXvUMrHWQyx7mBzFCPLdas8IebDrNgMhq/1dxD9R50fM+1maSlvByzBVxpX
SrPmGJvUHudsDPRaKa/icU2nrzLdV/dXmlVTBFCHX+Ijr/C4SUcVLGTf++J4kAxjCIUZy9AYqFcH
nBZZeKX+vsaEMYbohI9PwmBY4MKCULCKsyVaqbOpjcTTWv1KU5hE2C6aJ6zT83Sf43u6DVc9AeUP
Eg2SNwMmxFjs+QXICTHcdmEd573thEIJuDOYv5ErFtB6k2suS/7leqqPgazC8kZcmK0r7NCk+aIY
KEOVTazeIUikAjJByn2ZzdInBKUT5muyydYM4uqQNr7IwKtAPfyIDZSlYe1bAp4FdCy26QbB3OSw
f4i8wjA1UFl98LzP66Y2vyBCnGEg5Rd0EathvikxZpvKsWrmwdC3LUdr0ssBU0srUcu7IrTq/h5P
B9O2laRY1VzIQxmNAzLyXvTt6+YwyW4qA5gSiYdjzUMjLdGowgoYIA4WqjxLuirMdteX143y3syt
1eQBxJo0Ie8gjIql0waNH/koviFHCjybfZA7hhV3PjpuyuoRLU0nhwqy1CMpV4+M6P5i8pFd5qEm
BzIvmzu4EbCM6x73F7l+oR3N2JD9eC1YZWET88dAXlX1je1d/rnfxNwNohGWg9fPhGr5UxRoscI8
f2RJfC80GbLT32bJxtovNaP0KAkKQLkxXlm19mz9uCf+e1Lg5dkNaV44oMmPnltCnF8LxJS5KwFb
D4Av8A5jLb9kE6KA6ZdUyQKTyq0XnMn9o3Hfk/Tevje6zyGLwn7dnSaKjhJT4umkXnBVXfwCeHSE
ce4v+2qP/gARUBSAMbFxUFJz5E3BNoD+L+CuqWtcF5hKi5BqMCVLWZQZQ0qXc10GctWHOydtnCY/
jSM+MqzMgl5rYtBOacFK8DzadSCINq27jiEcl3BI+3iAmLnFfT0A7aJBxMrJqyPqpa4znWTbkx9X
K7r+l7EZcNdNInSMs50gHh06ymoA2X5LkrV1ywIgVGq6zKt3x7dmNDYsYyhWUF2mpesWWlmN2XJn
9TjaiWNZ6+W7Hf1BSm9Z5BbmyHJM2dROQ+0W4AsggcLH880TZZkoy+TZSq7NHgLZLgvEhQ6BD4MJ
CoryrqWuowQyAdA70ZPa0fmc2S2MEFjIJP9HTuSQgi0NRATIUVU9UOoVnzseLGTvAXzKEc0vPvSy
93VPagqQ1iq2TKGARZhh3pqxRW8QzR5QsUmYpoIwPrTY7L3jEmS1uKD0oEBtWHZe2TEJ1GixxiB/
+3XWwbK3CJdCmYGBB0bs0Hy2Aj1AXiB2Z7pqEluIFPSDKBqPhOEfNH0bc423hzIN/ce0gh67HD8Q
9Ix6adX/d6OIzt5G6kSaYBmOeQnJTjepSaXl8DtJgcTT+26FW+Cq6JljgqRNa93N8AcawV4mQfv3
km+/jX4WnOoQPWR6+uX4sWTFRsR5sDMCvY8paWUUB+4WdsxAyYm0n1zWmDvBfUAHxCRjIqBo7A17
ZhAILsycsT3LNUF8e4tDO9tJBN5YjkBDY/VYTvqA0wTVEJCXBFIn7mQQtGlgBaPHFHiIXhLVCW+7
YMKMFl4dItk7mA3DX6qpTNWOyEHS2nKi01YOi+DAxI8A9qISgtkSsp9FdemEX6hEk+okYqkMesn9
LYWG23IeOKtFXlirEOsIUBXCo6i8/60s20fT1zDq57Xtl/W8Bci/UDil1nrr8xejUQn7ZWz70YS5
8yoVBhwzSfSrwOxjYhLBf06OfsZwp+sxOIgiBwOOm3hBOY1H9C8/cpWwj5kTkGaPh9HHjEM1Nn+6
NoaUSwbb32RI1A/+N7u1E4xS6ae4nMNXwPebMP2BMsvP8oxsDNWIAXFqUNIgwolREKzJR8nMPs44
ai8oXj1CQ6cT62ErcYd90usEixBi2LLsTzA+ZzSBko4FZ0AxhTZtU2ttap59yHs6edBq/vsanQSG
sCg/49SkA6oMnhPWLFy7pcfCJRtKIr9rSxeSh72HARb02QgY5GoZzMS7ay2u1G7Ez/Jiu+QwhoH5
YBULPRiaSYVTaiWGpmGZAVpS3mitgTSzMuvOIp52oTOskKRCFVw+9ww7UqZd2Kpr2vFuSMg/Rm3y
PLvEQlgGBfhlT6pWQiJFqLZupbFjfVsfBnGhOw+VonXS7l3KOnUV12pG8XPAiLEK8ZBvMaVgFuuV
/pptdUKLB0c64pHcYmQ5FOzuvgXscvTxQAhCCwdebXzf4oebwXFUzFjEQHxinjANEDgT3JzzJbEC
SzNrY75CT0NmSz/WBrS+nt1wq928n3a7Yo6gg7NM/aICDEa16iPfZomc8M2NpuGIFChc6q2ykfHl
JE7aGQj8WkgaT8AR5sekYidb0NhNx4jIxLFk0CuTudPAQgJ5eSrR+cF04GJeuGbeOepI8IRRmr3k
a02QhQUgTkcXPJjn4A3E90//k77xUZnQwCStOGWjCMG3u2WJCawqJjScXiC/fmS9wQTchtri5Mfu
GRngbUhNX4qmxHMdfq05b4EnJj1rcrYQt4J2RHYuKBcXP/Qnr+72FH/LJ2uRFHaUw2NjD2HdjWqm
Ig5zuUaVMXI4lcjSXIPLQi3WE2kitD9yxwk9sao0q+0hYgdCALYqkQLisHp4YgD8hKNjoZAQupkc
BfeX9HEWyyj9g+5NHfRsbryjJtFbcw8r2BwSsOOaqZkAKMaKqZQt2iCnfsnigNUrfuMcPaMMuZJQ
swg+nKriADWZeKFRVXdrzZqwCqvTBsboqGMLTIPflNh7Cl3wAUF5w4bEdAqZa4DbM0DisihiWrTK
8h6UGDQ95PKefMb9Pa+MbQGymu1bF5utnHCgMvSklBE2z7O6xyQ5zi1ypqt0X3LFaUcrKohfRZj4
iuPxMZKNdZeErCr4OG+9iK/DL1kD9FSGmrVi1y3QXtF+ifGwy2ZDydY1D5b/D+R41LzqNmZrBBoO
u+Hli1wul4uWDmUvyQdXKMZCU+wbUFPgaluU4FA4XowvEWLdkeQpcqynBWhtzpa6YVeVnKbc2a9F
yGCEkeXvo3NWHp85jHj56yQ2vUi+sUM1go/x8By90JNlVv5aPXpO65r9DWQncQaHky+K3nsJGCmo
+/aogggbmqM0Z3i5THOai+ESqqNrxTjogZQ4MmNyyWtepmhvb+EGOkTmj0PheezRDipCKOU07Y0h
LBHsAiTAhjnYr63JuWRrQ7qLrfejus+LYKWE7qHQyc0FQxd9y/JAH0k5mLyJNleVBogTCuq5HIMH
2mdtaEv65UYNbQ8OTAM6hubuIk1Vfk5fObA7W3wgEvdeJf3eXaVqOpoZMyUkIKKS53/GbIV6H3M8
KFqWLA1qERl09ODtoMN/BuXdjNYbXBDQSXKO4cJDPlVQZRGpBIP/+tkQjeyGjxqWHdEoO5TLnab/
lut6MBGsCF6br7Cnc3RMiYOV0POyS/0ij5yq1f1eI7NWAZM40as/bPbefNn2qGDir1GZRy4AZW47
x/JDzzwgwY5O/xeT4guJjaXt4uASnJNa61oYrwXSOaHJH7rt/CAwej2GkptKZA11T7ftXoZ9WQx/
oHoxxi/B3INJGEYbTlnEINhtDwbp9G/Nw6mKiUOdvkHZFVRo/lN2SZEtgaGXCXh5Qpv7EL9lGR8w
pYOhWXxkif5i32RqwUWQpL4v10E0GC5L8JgAM/sZ+i0xbTHz6Onol1OPP2zG1uZXaihLD0f+KMJi
5XHNj/4XLUhaBX5JyAFvohC9VLsCCD50C3dwZpzbwkGWFYLR2c2gtqvmJIE4WVFUklk0tGpFWP7c
9vFoN+3d3IzvvqJ/y4fBF1NJ8yEeFqsEqRje3FAR4wLMDJ3/fc1l7rSDZnRas3ApEtTspawqKakm
gXgwoy+0anOYAOThRyOUe0FAf+UEroFb+KvYAehB9O14eG9kMsOW243KC7dXGlwZbFpZ9S1JGvVt
KGejHaoOPDcx6KmietlhIk7obVmBcObApUNcOlSd7r557n/2KxmVMvdTA8Cpsg8YxOETFDDd6g96
eDNqZIlNo+ILCZJ3zFlVES83s4ent3zNyhirWxcV+Jwwu05H7fxeklNzaYqrRXBSTJDWhpaBH4sO
mHLV82iSRBMi91F5dd41FZ9lNABB3Y67lZqRZnh3qCehRCfOO3m6FqdRlyYLdNWYv1uaslRmaIbV
qZGWNd2MQhrkKASw+gLOXiLGqpC4b9uhXXSrKy6qHSMCcp2it47jXo09arps4ec3X0tSb6Pk06rq
VsQqwwi0QgqKt2HE8qZJIMZ7yM5GxZDxI1WcmzpOCHlZBdw+xWRbBAMozXXJkj5wFqtKSEoO7QSa
IcHbZ7mRfjg7eVTxCJPzZVQYRV4hTXVK/1pyLjwCwcq0ld1fJwe/qV7mxURfG+xFqupjfxvrD3Ee
6t61fHp3MgBO2jDgBUYi2qYvPv2UFo2Awx8lYaLxKyV4aIbwU9jGBbW8MVYWkDWShKra4fvWVAiO
NPPSsgVKAF1Ft+92CqEQfPilgkj3bR6i2tSYQ9Aecjg3WBLPrnKYs4pCwp0/C0IrJLmZduNyKzX+
PgpJhUu4Djd37/+ocXqXQ2HiZmuTYLDV9ND+JxgqXVW1lLi5NjZIkQ8onU5QBEhyZL3agI8jVUY6
36Mwx+tslFpBWIJlnY44VNC+/YhArCKuXXF5dh3elURDaKu/EXeHb9ma7UAm76X941DlRe99emSH
JPdwFlwT8eHTc5Q+4keMCMm3T3EzM83LB9oGi5NCz6RIZiZz73ujNaBmeUCD9YLUMNRpCvT1DPbJ
Nzy2TlJMo4M7ho4/gZLYDees0n9RqaaSUUAXnjDOQbaxvViTfj+baLCzWh3+h+yyQYNDyi/8NOEc
smqUmeNeh9N44NcVzF25Znd1qGkZ8MP4WKIembTDqzb/xZzyoJZSZCFvt+VZAG1VtqltYzQPK2P5
YusWW3evStO++5T9NBIyROSjCBs5rESEYN5YLfeEE6ijFVFp5z6oavRM7rrALd2ohYrCFDh8Gy5A
4mxtEwKMGjbQDjn7K/ps2nyFY+WqJqXns0LZR3Q1X3GcbpU6hz5txLKOQ4GeELKkuBy0KXwC5qNd
2ZODXn/NcQTKymYPB6johaeJRP3ATV3KYPsfNxwfXwVbYL/hm6RY8DzqH2eseSxcBAcRl0GZjHpQ
pVb31FxDwQROzHGptgtKL+0I7SeuUh2jSuMy8spwtEujbR5VfPgbPbbS726PIff2Sy+flYqar8t3
+hZdAJHatPhnG8TrNgSxq8D1Dspw+9rfth1cx/ZGvA+e/s5PxCrwfHfdBAICwrq0HA9y85ujFoa1
ihvgZi/hm3rPcAA4UNkmK3kCm65HIXj2og/aQHK9ZNkjFp+JmOymlZJPKv4eemtRklF3YFrasvcj
iaFFlQ748vjlB8HFDvm60cRH5h0J5ox8aSmcq241BSBWZHyp4mrCkkgRoPqiMMhC9cd5bUxvCxtA
cjsJ2DSzMqWf8w6e1qC08n+VDESFlVSLpE10Ue6B6E0SmqbW0iklhUzXXLrAE3D5K/mUkeqb850f
/41LQ9Go6POotcyNDYtu5thFV56r5Gy81zwXfXTITR1TGv87dgIZBAKAYA56uf69CwyR8J3TtSBY
LcXS2yKPpPzWe4b4nv310hwXrCenUt60MA0ckwCWxCGYer1TswhoGliXHMqOkTNnsUE6b8dv1ZAz
tOQgMZ0+KQ1YZpvKBxmNQHpKffTjH8q8TGiJYwRjxJCYTndJ7Nx8EbzCbWe+BaI3N6EQ5PErJTmR
XuF3SJEBzy5QjzB1wX/ccj3JQHcxybEH+cdOjrJHcNVvHdMz/ksPhEmMOrqoknoW8QR6meijyYW2
pebPIqWK6SowI4ipbkbbih9px46qcdHjqCfxra9w7+C6JepDpz9P8XGBgb0PY1dS5NMgBzKA9RKX
rMLKSbjquCW2ZpxTFSM9OGDmhrsE+MyliMamSwbaDlUZAima1v/YRvgSIPEFIqmItn7n7ZbkEHdK
011iu0eTYpMkjATa3Ex7dm7MUIqiwa7kEgx0Q7Qsv4fEAxKtHY6D7N2d2uzeghhPQMqLPhrub9IY
rEtFaeIYAyWpRL4kIdJoQVZ+m8DRQ2uZQ2ZYBEkXXFw6tq/aM5BpvjzmJK725owfW5FM7Klfn2x0
1gIYCdFdAP7COEBCLdfN7D27ystk7uUhwHcH4vRNBGF11WguoL72rgqUelRvwgq4cuxjcKL1MZFN
KGv66gbvbMLCfLnHVFoIJql1nqA3hnFyZmiiDNy76Scs/x8SSx8rQlpmsCSo2yL+m/zfvoSH4rio
JTCgIrqSTOo8ggHQZOgZbK/aR88YyDHu9lnYE7D6OGwTHhJHdrkLmvKVBRGoQy0Bkenn63coxPhM
3Z4FuHoLaGEdZh+2xrtg8UK46Px8gUfpN0X95fyTz2HdUNzceTCaNNcekBFr8/jLO5fNLb5XLogC
WCOT0lF/JjbUasiPk2ZN61f8HLN7m6svGKwT2iUPAAPMt5ByQRlNrO4tJGmlOH5g6er/4NJXrweH
wcgbajvQrlC+YqQk8nmC8tTXzk99H+cvh7mHROaB+udrHcWu9RFGpcNlTybuUP10KUtQTH3cJqsD
iOiWf1KnSVuZe7Mhc9YKunjqKuC/YMADPJASekeQTxSJyfGGSYFNxMPjkM9d6h2mBttUqG+PTlWp
Fwid9vZkphblUHeDTLS3GYF1hgIUszAIxOAGDf0dacemWZhBD24VDtFzDbKJRervVbV3dNMhacbD
1Jtin5UKxM+R1ZSwEgk4wJKebN8nPtgckCf5eGfcbQV22N5YzssUJ06Owhclt8R/Cpo4gzpbhrJz
pxzfDy+OxyaMb3FizDlnzh04EHr+Aif9R/F/FYuDH7ntYb2jcJ6WdFqkX3rwlZrNgbDgMniSyZ9+
VvKRvLtB2weP+NVvUTfYwWSgbVg3l8Ok6Xq/WHb3BWBVb3q0grKKgpBEkyqIyHPAPWmmNcgIQCHo
K4+RwlaFkUrl9X0ziZkzyoosS7PC8OPOEUHpHS9P6eofQDP9KdppupBrVSGvnXAJ9EiRzVbb8XUj
rx6pBXt1WVttXR6V/pS1zV7XMJ7dfUr6OWqBbSfur+JQ6wqF/ntuXr022nmkYLUsEMJz/DfEqKtX
KQIvjqQtvcryq7pr40D+egi1kCCFJJ8PP9WwmPWiSekhNUU7nArtMki2yZdde9U6yGGG4S93/hF+
0+8hJbqFNU+Thjo/YTvFWDsyeus0XUelYTkG0G60nsPVU/FQbFXBYIg/unR9c68dEaAouKu7XVys
qbe2RHjxiNCPwKM1YZp/CmpBidPl+nXLVoFcFF7Q53Ayk38HLOU1WONRx2eIL2BTnKQ+Z0qbgOAR
+1xsPuVGanW5MVVw1cUKAMd9ihvQhiOXSjfYhnHjI3L2qHyML3Mwoxo21T0s8LBBxrslKYQ45IDn
sBoZ6fCxBGfL98ARP18ThR8flYCWXAcomW3AvKLLyrTnTbeZyABlDEYx0+nRcDSqyrATAvvIi0XG
GECldCuqSBW5tR1i2JzgFkYqNyQrdwdfeQHAnaB4b4Zuj+xys9BmM5KpSuWMzixp0OZA3Z9rqTwi
09W65PQbeO+MrPvXffZJuUQ46tzf0NAagI3gGUVLuMgijXzpuZvLa+l8Tx5VynvXfpJnOrF427ZU
LozpPIkJsEd738L1Aq2drfs8sADGiiLxs2vXzU7zDh7GnZfPEh8tslElsu5t1x05+bZDKwSwADVS
B7lEcz/U9e0owEDCDTNP2OETcjIju2ymFWI2VxTh7ig7hvd/aCjjo/Vf1MFzz8U2+9OXzJAn2aLp
9PYevXdHurR0txQ8pwnxXMb+kdfwCXmraKz6u4hpn1Ua8Cuk8PE8ois8c+68nJCq6pmhR8IOFUXk
ZI7IDsluByD8zRQqsHT1ib/vLwLnV7wQfDuA8ncn4U4B1Ebqon+eHojCNETeSuwUmqyQ/WSGERB7
QNmNp82KdzxPJeLH8kjdYDr8yZD5jIcEfL15kPLIhZZl5MI8TQtphuPtlbeVVALhP6pn8dOFXTzi
nFPyblcVts4URc2AuqwOuOeCRcvyjZxpTryJVmu5wy1YnUBE6NBW5J5Cjhhyz5NYgPUnTUK3UmTp
XZ0MfJLULehk9d8YF0t+M+D9RJGXnT4+0IcL38q5J3TBykthy0K4207wMT2qzGwDpRlzV97rhARQ
kCl+46XCAjM9fm8FeOqSdOpKbfYq2HgceNsE5qnYyrO7hBDS73WXa05XLYEpnBmec4h51Qpxv3az
h0ePNrVbQhFWz/75LMciBcECp6/9ZpGkPPGTUsTPMx3HwBr17dLXzKTdooxo54wHrXgLlTU1P2kR
0TFr+DovfN6u7ReoedBtjG6JeOdKyEz2TTy3qwUHMcmK6yI+t75cSd/+pIiOaX8qaFJq4RppykTf
MPtKdB33tqurXjGNbYfwYJEOq2u7PgUcwXZWEBmouJeXojIg7djJ0dKOBSKCbLBImNIADN2OOlLL
Ig2EvU0iMGSzzn5MlKaoOnIgo9DnOYsCcvnC8C4nTxqB0lZLxyTCNOp2XbofyfXRqLhi9VVwMaZp
7EAP2HhuHCGs5HZ8SL3PSH+xBpgCoPI1hisq1P2FlLXFpxFXgCU91gQJAU2+0ioTbX3cYYsoJGx5
hENAF95skay2AxiXzQQUD+ZslvuwdyL/RpPHSWZ2Mw5dlDLs7r8eq8V7mZLiaNovUm2iUGR8L3Tc
MigzFTRsGmaxnmxSqAy8C5Evb0O5R+0+OWJ6hl8Cqaa9ueTD3cEm5RPwvmlbrM6J/IXFqQPq47f+
RDGKSZwjAA58GkMxLu7O7EWHDbaN5OqALW4c0zmWEiJGUaV5YdxQBjxEDbD7awSdnhEyac8wQcEO
tsaNe25OKa4O1iNBCsObQ6Suf+3mEb7Xh52JICMPXDm+5jioMKGaj1QTV8W5f5uJ386My0dv37ef
HwVLNG6EKz3LwdBtDj/1mc5xe0V/vlHkpmyfWJGXikzERxukYiPeSgWdye/eDttTgCBOytI7v5iU
8wkwewtOl8aFSNVwtcow1lVBX+Ivqmd4tycYFHvY+TJw9dw21qgcQ4glawb4BVZx0TuUX0yA7xu2
RssMq4xJaqgQ/64IR53etSimtV5C6PXyVja4oKmYpSvPuLVMkACwv9CWqUG/TmR7+xce/5FCSK9H
IJCOClqD9O/35oBGF6IoZ8tmqJ1YUQ3coS5cTvfMG7cHYwP6kXyKivaS3UlJXSX0fbX1l9dN3yrK
1LR92uIPccoO0XppUv/a8kPjlEMg9IYDhKLrOSQwK+CnTlwLBuDjrL0o2CNi3b9aybYCbrZP6EmG
o0LV6RcTgHcuc+Hp1t9W3GvNR1wiTXG9VDtbNwLzb2k+42rFQ+O3TXAXnizanppQyCfLYfMI+IiI
jHQ6cbtzan1Hch5nQfv568REG/qlakoUVldJ1O2xgEi5HMWGjeHdlmyDz/GNlrYAz4X5ZYk90Jx9
YFW/18RIjdtgeJu8WNRDFXan0i8at4r3nwCPh3cGu2TOH7OybPqKFd7VmZOTjMKACWecEbwwVw/p
lcjpTr7CSQBg8kxguRxsuTI0VCJowZHOGJijfxXJpk07EwxLP3j3rTrZMukfTW0PQHtlV+8G/g8j
1L0Xcyu9nKCSb8MSeOIcLZCTAZ+K/vOLSteqJvcj5U1JkALgT15Sq2dOwPEBHpGckS8GNsMo1e2c
I/xQMqKfUTnluSmnttzMJ+mb7V1OfzYbSsGEvgjqNQmNidvXphCL3gJbKZX8bi0rEoKeW/WtiysA
JoOzxci7DfjmB/gbzGIfjQd2M8FVrS6J/+iy65WOuWOkxY4k/CVD7XWOSLtq4E/c1n5lA+dR+S+7
RgQsCbDaeOBRDDf2Nlimdyq0xGwZwdC5zGguLD4XSVMh8qro/Z+FOdICYSC0JT/2omjcRcdQmsvg
I7a0yvFSC8FKVs+a6oqQJgLTkmzgPOGj5ylAONTuErPhMg6Asnzvq9fQkPQm2eG1URyx6YDwHXWL
EbyD0f82TnOGigU2OPyDVDM46uksDtZOuwXSWkdr70PtpIBd64UX9uRd8FLOlQlkDuvlscj6cPY3
rZjfBlMHOTwGE8VwsuV94FvCikDGv55ca9n9HJ9Qgt7dns6bgcfaq3LpFWLUx905vY0kXxE+HE92
jH85vgYgLPC9a3XWxHjmqFLoYiASEjEolnUsNg35GvqYm3C3f4LuEeEOBII2yBBk6ouInTJlHGzF
3wlsIkQYtkrqM4A+mOez/jVHUgNw7EDnUUnGijAucdJCXKJHdy1kABpx6tkVCZepjLySp5e8hrHN
ORy69EE84f1CtK5lI8amSKNXFPBNX5ditk+dcLeGztvYWeDOkr4BU+CLPowx9wFVZYLAlf9Cpvkk
W2i0FMfzv0rox4mI9TCT6ID2H4Sm0wPCYrrwf5U6OE94UDTTRP5icY39sUEQSGR0NPwuVhN2YFi6
8SpmgjHmdYG8Tgsj80bYKNo8F6LP4z+f7Ur+1KvNs+BPQ5XwbzAZ2A8eTp/LEH1aK6alB2FFHir0
wsyULpvZF4WH1OUS/53D0UDjZsvRswmzceZWp8zC4SHypp0x9sgD7UzWpfs4PaDNEpZiKGa0pJRk
dpYW4MI6kR2cZ2lgymSfXmALijcwzE46r7Ddc6bxfExOOybxs0hrb080y6JALQD7uKEdAhEJyZR5
UpuNLgEN2ttxgiQdnOFOEFUrKg346nhqaEy9l/s7wlOHP/vrCnlzwO3Qzdn+SxUE0+9TEtjgKMAc
d71qBlsKEdIUw7p5Kj3lTylVyy3yezz4GgUW02pmPwPAG3/R1RCXdBlRKJxN1JNLCxRUFo8eIdRW
OTm87kccyYlCOVSe6l4kfJHe9GydkGKJiCLTSDBuQobbXr7EiBkvyw7+xSLiMsPqH0yhV2nr0gQp
JL+U4A5DVXJ+uA0ibWobrNQenOG6gNPri5xHBni8V9rkPeWwFO50IsLAB87XexIeTsyVwfHYVQDb
rps50DB62a5l8sWgKDtxuIGtDI9OkmlysaebHKNq4CpRGqv1Ou1tJ1YkT5scMaPoO0ptKAPEllwZ
Io9tyznpZPv4jP/+chUHn7xthgIObUzCxVsVIQQF+5Ovb0MnhoKK+GHWsHN71qogYboovsUTdcuz
8Rts/ADibRoTkWv+1gifHT8EZsEYqygU2YN8Krih4fUasRjKdUY6MHH/gd529kYgMr3jmQzT4RdF
ySpJ3tOOHe7SfKUB5o84SeCVu2W/or2Q8+j/YV+jF/w6rDYb2yx2mQMzFvxpQgQePWxvEawSDtVG
aCHrlNMG5aDdB0RZGN93i7cJkoceNb6I0k1A9QmdpoBb2P3u1F/Rxb5W0iRpVee9ud3brDKjJ1/d
8CDDx6IJaYjY/6zcwF/QkbtSfQg+mVmz0KxDOH6PyyAR+1dujWvZNaxaP2MWWX+HqQbgpfxbj/SO
wLiymy2/6le5t+Q4WZhysAQNb7YcneWT/dcmd0NNnf1em85tidqfR5vmR51e2EU7Wt0v+Dp3hMMi
TvOHwZyqictpm54Tm1u/pp1M3m1qTUjpTgwbWPa9yAN3yB5VY3Cktk0BusG+t5nWokyebKxhmSYt
08fz/7rsL9WvuXKEltTswBH6t0Ulruh9rBLvyngV+nDfGtk0VhuPISP5c1lQhIklmuE9EXGud8Rf
JMtLcEIeNgDSE4CFn6rsz9gFtDxkkL8nVRQPfZBhT7Tx4npXJSciFVgqfYnEnjFZl67fF8ZG1fHs
wzgtejF2emAFQBTRWZg3/OcNvP2ukU4B44G7qiiTnbk5HA4sLYScmGbBJ3glgx6zqrtl2CmJg/fP
BLp0cuKgJpKgda2UuCzGt5xw7+RWV8X8bc6TjpAiduC+0VVI0rskQE4LEKZ7awF6Vd/ZkhWGRFV0
q1HjavUasUFxhUftfA9focw1Kubj9YOPhpXl5ZD6Yx9cm+Dl5cd923rrsMRdYw8RbXJ6WiC2CihN
NLyfGzqNuz/NH72KlSnBKOL8d7NVrKJMdZEnNj73tkR4Livkc7X3dYHjafFU9pya8NyE1QnE8uNI
MpSgFoj1JjqbkGRqEq4cNpVCdPGeMSkJfHAWEnaWsDCPDDlSTiCUjr0TS8dqGHZrz900JcvWiTUE
6Tfn2xCyZaaF8/vF6ArIQOHhXrXDU4aMXNJInl3YMy+o5bXp2X0w/ggi/uvBmHnpTDF54hsdtbM+
tyUoykFumgH/x0FersW3+IFsBP5D1nJD/k1OzxJ9FRo2nWUQumDPXTL7hGIpUCM6JI+teSjULdsO
2ljRsiPWu2uJ8ngvIms5dcVZh6tPwYaF9pr7qdDxwA+OJRQf2Ibp0CY9UXVW4BRAq5z7+2IvLieW
Zu20Y+QEeA75llSlhROkHzDWTGnuHcNFr+WrT2jfOcmjjrAabXuND4/IWMw3reTwmYSSFWJxUF8T
KQaiAYtrCCNlCXNy+pFPguorRTvet/VJyGjxb48tNJZnDXROiz24EPlIVOrctrwZa2cFfqDeYK20
fKUpY7cx7U99KflWbL9Kcb6uWnrkK3BJUEBllmMufJOy67qgxXUryvj3ygqnc7Drhb0sdWjbzeJh
6AWQt3hjaRiMZf6xfEe7UzSMt9LpXY40QMxiwJ1kJZ3f5T178CUtGKO/AvafvJ8HHH9Y/AGs/YYy
PIXRvrKDJZH6rvTAuXZLrveKhwaHTsS9QdABo7PxihPiUBua9Q4NsqfLW44vbZoy39qDmyIpAECJ
/58cPbexp6qWoTCG1o5dTeTiLbgEX6RXxCS/NwfnHqY5ON02Jjt3MtAZqTKV8ls7OXoVSboTfOzt
bLWaVpIFW55FhxqVIdkcIq0S2PH6EZOfMsND65gHI2Vqua883epWu0EJgYYdhc/7oNShU8zP5zN0
fVDyhJdfulRM/WJKT4fIn8oD/Qwb4iZTVGmZ83y8noXSnfVS1TbnE+Jn7D0rj2PhKNLx/5CggmGP
Vu1Wim+OgJYXQ4cKaJsH6m/OcA/vzQ4gWAYXA+tFxAz6WojS9sEbkf5jLY/REP4DsXxlYdQzekN2
ZZV32aCes2p5ZIvxev/IsOLhF4sB5CsEfouj4/p6fbGfwzJBTAh1bh2W/hXrPnvTC4MJbRUPlGtk
avr7u3OsG52M6wlwdTqR4xGLCVsbECSQ9fM0otmsyjOicFgQLlbbMin6z858zstzC9nuDFJnhqzC
BM4Sz0Xqnd3lfrVGOlcdqZrve/UdFkyDuznFnUaCuCo3U2p3mGeVMqqc1ngea4Lm5V8yo48OeLZX
p1wHUFUEk4Z+VvTe1VCWSyKtSFFQxdDIl+/esXrIK+qk/iC8fk3Ra4teXOaQev+cRvWlVoZjr3X5
vqfK/OTdT2qocfrGk1bsY8WDJnFHeNh5/pFTFPc683qOWgnI0rdCZMhxuGhQc6ulcbIC2P9bAv0n
aB3KryxKfJ+MJOHFaGKDvk5QC2oCS4OeTfuyYansuuzlnbI33nK37D1r8qZSyK0C+RCnng8nOWZw
iFYXovnbxaG5bIqMGZdfGWhX+VfYasUZNTMT8aA3FggAPn3NiwXjhPOdtW89ra1EyJYyyGf1xI0V
+r/SMaRg4zq/8U5+czM6T7P0Py7Ig/NHq6mIXvDzPNDQvqk0FQ3aVJp7XJDWtRLSWxkIoWT/Mjds
i3fPqG4vj1Cqpw0ZO1slmtS01WkyoZB1MPdu30vip/qLuCI8FQetWXrS838vfDeWSoETXmbqjmkG
Z/JIIHB62MMWLAZ7cQTPveVnYY/xaiPKsVJRo018o22PdBEHy400+zR41CNDIlS1pQ+Mb4D1iSEo
jKbLL1Fbmce0/6fvELY4UUE1k90qiymuKvKpwLQOsHSOoI9aLfzxyc3YcDEIdUaCsk8BqiEGOxuD
gADhnZnuTJfUaRS5LVpAs2YsWXUgr5+kdILpXkomLBQUt1ZWY+7X9xOsKZYJmIEend+VJCqMMG/U
ZylAjF40xetBVUVXFufwJsfh3vNZNc269/a4ChUxSQzDR1CM672A/gVph+7CuQbI6zDocFR5EQka
WOsbSRY1xhnvpv5vN6kef45cxcNfW/S7FDOK+fx/cJg8pu7SJuUrmko99sjqSPeXTQecFgB/vglK
/DS9+PN8gp31GCXErXqjYfZIxbuxIg9giUlfQ+cpMTw4P9Yk32SxRRB6ctUTx8AfZjR0r8t9+zS1
QsV0GJeHSxZOQiS1iTfZdarBEW4cYDMSa+VDxNPNNk+ekuu2bXzaSszubIbLU6eMBeuKC6MSeZ29
KaTm+2H0LP8JvYhKxae65ZzVhqVb/WJpQ6NNecXEb/rT91VjHlGXxJoFQlBaUQykHR1gGOUH5Pgl
YgCEKJPDHdzX2qjBRncNa5ti6nsUm9NR7u2uEQhv6jwMYS0siEjSlrTvpkE9xGTCbDPMiXhEfORv
oZXqgcpAAXVBiFh4CqbR4mVcEP1EPxpGI96FsKrZtUfxqegCjZs4YEpDrIsEcZ1qlaksaoCI5MWW
TM1RQTWviaSnJKO7BnHzYjdQfalRZLIKvBt94WyBqRLWu0IfJJWMNlkYvQo0g1fZChVOK72aI25j
81sIeGlIhj7ce6kOX1MjOT8cZSR74+SCF7JAA7W3Jo7BZ7VKKprbT44A8jhOgt1ygBL6BQTuUzth
hdHkaPMzn45F0UdT9rf8CqBAklRRow20MHDRkmP0Wqnw90QuEYxoWR9uWwqPk8eBW04drDdzkfj2
3KZbPc4tZYUL5EwyBJSJt1ee4DRl5IYiCg1tj0PZqRhjWgvcdJSfTW+UIr85C7DamcKKwLpdfJi/
Ko6sbXCBVxJO8xhSiCmtXzy1gEu8FRcWEWr2JPGQT2x5l7yqvRP+S7LmZ8gLAWLXnz4xNlQhj8cK
E7Jug3spZiZavzSv0CquyDrFkxIKTJQPH2/02yv7B1341QrwjCgKNjyNgmdbh6RB2dlVQ69DUCwK
2rpq6NML0yfd1aNYWG/JYaEI3XMlnAaYdF41nUwClsydhZMMsyGUKWg0IlxMC2hEO93NiCXQJ14c
Wk8Elt4I3xd5eAH0haopmzYtN5PaLalw84UKu3SJN89Aaoa5Y3x0Cshuro1hZEZPjXl/rdxZpSgj
7Su2C/zc3gCUJXQqT2QNOnYJUaz6aTbkj5OYzI3DpuVuccSGmQ2iJJc3JohfIGjHB1zrcA/hV3rY
LhxK4kNApB7s/UvfatJRdRZW77n+B3XRdYZ7ea3GvpYsTQRyUhICHJUXrV/hn0lRH4zHmPD4l5N3
QLn5SRyqOrMBCTqoa3xcT0L01S2pyuTCNfeDke74H2WnZWU06T8U06L00/8/Akqtz3K8VBAuVOby
OlVaQQOirHgxkXNdyz/5pQfTPCiHFY9YllAJkkHCcwMqwqtQSpvBzWVo5gGoTKuWuI5sFBV0vUqC
3q+zQ07QqYXJu5ODEhMHxc8aT95TemLGAlemGzsg+AnlxznRleotfK6tpBfNotm/VrMNzBFeR/Ed
oDEEU6FU9xe9W3zMdsg8fmi47WePo/j+cM9gie/2ZJUt+OnkMtLJzNz9c4j9XwcbrPQB3wcMfvbK
3OlN2y0KKayWz7hZ0GGzUM3izexEdsrRP/BIgzk9AGAyIfPnqgZdw6mOPQZYmV/lkPxFiWxEQfHZ
wJR5KHHlcHav7ylQg1rfW/3Vt4aSzrSjM71kAMNiWuA7W/q4J0jmeHVbtiM8/5nXSeYf0ofXdbZ9
FH5YnkoAtqqLgxdsG5lfMzLu5i0gpygd7+KU9MVJIN2ZO9Q3OaiI+9/JD4369A8CfN/W8VkeybPO
5lRs9bIr2J1jYwZqsa7vUkPb2y+7od+f6OSWaU8RZSblQyqrCTb88PU3Uu2VQ7XNQ6Qk3ADDAaZF
EgRRwJuogHM41INotMt01QGcwW6hWEyXayNbCxy5nj50hQ+vo37CBg2waZu9Xuqh+4Ytkc8cB8k7
hg4JYWx6gr+sujbxM4ynJkBUMBmTT5qMDTVXccZOhiWHzptlj3qnYdF79flQ1jIlJNSj4GarqQOS
6zVunZmd8H0W2LzpMxbKn1xKkgrshHcMf1qdd4dLKBqXysZYTYMIiwjGqr8xv8lw2wZnb5XZAsck
YAC24IhlvH5+025WttB27CGs+JahEhAVxQi0vV/THE6SLuieyl53OeC8HIYQLdPp/TemUXvGl1Kq
hBAAuGE+HgWV3HPD8Y5V8sFhfS9X0UP2PFNncpxWP8+GwGqFmcDwYmI1+M3SGtf24mTLNH0HnuZ1
m74x/wScimMIb9c/ewGMeBQeyy03qdIYPPWAcruI5L0lNj22XRlxYevSiKpIDVHzZ+TmsxaTIhB/
BnntjT5ENwH09n9+p8AMsc+AhdQKiEnH9/ACieVdX5yYzqT2uhp5jJKv9E4B/PGhntk0se7YUuwv
iL9PMGsq+Nzix6P0+qJfWf+LQD47zwMFNHeJJMVNMpVl5huf7ylgbiSNKCtcJy9xA4y+7rCwbnCq
ellKN4S2axS5ho0rBR3tp9h9f1VA/5AXh7nlU1eOp4As547vWUq/s6dy/LleerWyKYZp19kQefaO
nV6XHRR6ZlTiTKz9eO9lbfUdaQ25AElxVRqShl2hVo9wOJCoftww9rDpn2MgckIjdPzXrvGMAVh8
IKJWoqgyrhiWFIwiwOuwH2ZcA2hBzQyN4hJ136/57ZRvW7qni5jk27Wr2lIblYSPsmKpYDdoRy75
xRxewSuUb3/T/JrbLLjeRz8RRxnzAUe9wMl5HBUiPmQ3AVp9s/t2Fm1lHQRNzFi/2UMJJeT9Xwgc
UIGAdEVLXNrxTlZTa+HtlD0vz59+LtZCbZKmWMML8IQt2ZI0yP8uLyXARY9wF4BWDnIPkY6Sy2ZP
eS6cYKsnIla1oxQZ2fK1Eh0E/NOGn8i0+0y0TVLlfkqHVw8XfwlOPmVbbXrd0ZhGWB7Ol7IXtSut
ODDOjHTvlefSKB07xsuMcb5FRZfq9NIMJWxwTZx33LWRMgKWF18yBP9RLGUJk3Gl9LMoBDscD3py
KpqOBYVmjoSDKwybFMKzFwxyPzYTujYzqcuNPteyDR42dTJ6XovGKk5DZinjoWfSoWfA784l6wiR
qZ6R0Nss/crb6CxkxlA5rTEPk23Pw/clYWamjNvA2uC0dDf4MhYNjGhNwjeh4z3zhj16P6FPcOrO
mktZ23vrYglgt5lYbHyx8KQyUTszTIrrEMbrIAWY5hDpV0Xj7mZDmCZ5p5UL4m4xcHPDRjywcNoi
l2HHdl7MBVY2R7cG0IZsrjr614RD8NQCpjoB/LH0DIUj4BrXs7nzLSmtlZOs6TxCpcUN1BwPyzVJ
VVve0888ZXhEwzqD61YCuHe0ky66sQGUdRf3bHlAbiEWytW8xfz1V9g7SUG4yjhJAH5GTh8WPwhD
+4jgbhI9n82n5Hi3sXYzVqjoT+1FqzSyABlTLLQGbF4vB/JDfJJnm/Xp7gcvtyMvtkE2TCb4HnhZ
lCNwvLxnlZ2oT+5OEXVShlGQso9FPDiBwfAVtCk2zF8sP8CrUHiE0vM1Prgg0mzs2szurOTQj6Qj
wvIeDhGYpD/WsXQoMEIs2eiY5NbeOP7W1DOwEVJzdY2Kxp4gNKxNoUSeu8vD7UQFQw555jqhl1M9
dEJCyzwRVFbju96MXOp4B47Pqbg5E/vxApW3Q4/5CpHoISordoOF2JHLk+KMn35niHVkBNrkafSN
xDjt0TF1ycCmDP8Az6O/42RrvvDvIFdWUAi2IacfWlO7Rhj15HoDB7fhis/6vFZJq+5ktAvs0dwz
8GW2BqNl1wMkLfe+JGCd4p17Zn6G1NFT1stHAqv6JujtTUBoYADoSGq1dnWllqQon0uD/cXisogV
W+n9y90gPQqraJy1ECny4SlERfJ6glKyQuVVHd/AJwC/9gh1y3JZl6t7aIXcxrIGi60MuFmFrEpb
bzMft5NnQvYEuUees4g4lENpJYmH+ZE+hIeLJVPvRk6pEW07ePN5KWzDxuw5+V8jGFWGDQfyYCou
lz94ltiiBOGOt9uLLU2BgN/gUOlWTY6+ZWzAIzpBJMHw3OSBY5KxHuaVv43WHj8r6No6qKTqvshJ
CfkpdR302g+yRT7gAHuI9gstoiW1Vk/BFak4r3MouzupvTI+rVR5USLagWMgcyO6wKjgpxOrUB0j
keKtx4XuGFZ96fHG0OtXdx4YsZULLLUh1DNmdhgd0vDet8Mfhht00Abg66EXO7oXlTzaqD855nXd
r2mrhjAnwrdDucxqck+OfLhYy86uXc/FU92mQpMaAGMkMLLKwPsnVSiQfnAM7hW9A6wKLeox05kH
4EUrUpTMOY64IhPEvsUxSLJRtjwpLvJ337JzRwLo4+koyPjIrIQQyOw8N/Wh366bI5DUnGL46oN6
cVTbM2XOpguJLyxfXrA445d0cWICRzBqEhm5la2OF8FDaUf82GHgQeLVXqvozcu2YC8dbLqlwee8
frSu4BdkXG2GAnPbH62LF1RLfdZcoxNfXeC/eAc+LeMFiZcyI6CjXbh7uB0wibP4FXQ+mIRJyAv6
LjJ933jT9wWoq4cHR0Lq2OzmNTJFptVNyCjHhK0W5Bs9LcRvL8QGpxlHZGPmC4iAuJPu7vDAtVmV
D1eO6e4u5i6H0rk4ISmv3GSoSoAAj0iR3xUj3qGSAnD0k6XehpmPYhtz9+SoTg/4oVmZansLN79m
7lCTd9DzQLtvvXLgpk8UW5ZEiq9ggi8zuWQxU1791B27HzDW7Fs2xYlj4ua9vdtK//cJuBjNF2sY
Deq43y9muEdPAzJ6ev+Brq9RpLiOndSKQNEBukKSKICYnbpIcbcuT9x4D83Y9m9rPIjxC74tTmoc
w+tZPcoSwLKinw/wMXlv3uDM/j3Xj+8JWBg+1F71rH2YqX1igMFNOH+OiGEo/JM2+uHuIzrthtQp
GDQDlyRWeq4PWL9ddMlUCfW3psBiRhhHNk0LQGHBQwRzUrhJ5ZMMgBQxFWNWUjKx9CWj5LPPCi5x
vhdOvJIm7HSGYN3WK3jqqQmgyB2YCj2l5dG/6dj6g2uDOEgY3x38TZvBK9K0uCSs+ADDVL+TQwrL
hjffaUe62q1h6qd39nRWbAxbRfhFHvIRM0c1fMvSfpGe/6aIBzD0FMzsN0RPk9iRMh0PCSqcVQ0n
F/9LjG32SaSK1bTp75GskIO2fM3dEQDLr9zGp4jT1lPtDnD73vt9Ily/0LdZiV0gibNHcxbIhrUF
GrKvjY/sUSujBywEgVvqTLcNVClDwRYNelEdEeRXwE9grBL8Fn5HuM/ce+RVvPQiiJHfzGfsuSYt
bwYlhkDGQIEP/Q1pPLdasQePNwxRTdVDqRCuFwojOnykwclQKIl3ojAbAclyfTYVts7CKjgjgAXF
HXzgLW2i3Zis27SI+iMY07OCS0kUAxD0aoiZuIeT/BAjOSytl8NrfwtTI6zOKread4FYdI93WBwt
gnMR8/EOsrFPtLzAZDZsNzwCGABuX7ROKDgdb083rD36KHthOHaUa+RF0/gy4by7y7ft5pXwxlxP
S9exTFVAKvJE59KWHjc8DdcLcZGFhcDsI8PZ4gvI+xMbZ6bGop4qO74z9vEBDYCvncnOW8f58tby
9kSPoBfxWe6RM75ygcVPiFebKHVFLCn7dO+xtgFu/XqJvvoTvx6A7Cma1S9VOB9qoiNPygVBiHvs
YN55KBxRaIp9HorG+kEW4nnAAvxtVjQIQQbI2yR9gyPMK/AaPjuNzbjGVfg6BBjI84Ngi/TNgP3U
9ZcWlzmpPuLTVcQ3z0PEMNuvCWJjyWzncLGjMo448WnMCqxFjQXkyYVbpCOyEqje1gtMpHXWb8UO
S4yL0QleO4LtsG8kbMWuGpymP5Nj/NO6buEM93GgJVPGo06LXiUhljAXY6eCviHXSfkHQTRVSP4b
uXcaCcuP0T8sNKL7RdxkZJWv6kVGBhqptb8sj4+VT9oIriYQP9AirbeB0yCak1qg21z4s7Q3QAbI
XtPo8VEz9A68gzYxhQoCaCJo/gkN50XU+sOghuVxPcyQWs6Nmi6qaWuDQ/3IjodBjcj/MiL7VVKC
MgNF35KKKAP9DUHwW7sthMU1bxRo2oFWHFwLoxBxj19Y2vgyuu3Y+/0rK0Z7Z9wXaUfaoYNPrt28
iDc7W42IBGj3x1YQTHsH2NWpvKRILLY/Tj/003sPk33QnGBZuQQFXFbuH8Wbm29zsS1YHQftewb9
Co2vBFSQiKpT7tqiyk+GIclrxYWwwnS/sSF6YUIiGBaEt7Lh43medi7NoCPCBSK5Z90dJxKKcN6j
/q2a8GySlJUFiyY4rbIUY0wzCQX8cDQghWPTvMTbWsI6QVX1bB15g2i8Ahl3hBh04MGLuVluTAPr
ufiGWlxVICpRV5l/r3BJZ0iseRuQo/PUhnQD4c1284lYbsE3n16xwROfFljF55CFrVDxsUYdCTEI
/kNBPsTjIATGrQZXt4X5wuuFLcTPcun4tB+ePHEPCbmZju+nh36E2C8EnOZJRK2W8eP+1DTPb98e
C8+8jXxQlekgWVL7gd06DJVqkNNRq7AacBBhWACwEFvYgU16BE4r45WCZlg/344BLZBoz+PmEtdA
d1S2YDtsxPYrxkuYYZYoWffWCEd1wfgmM5pYkn5KrTxx4TYh/94pfQNCabbkuYTwR6SvFTa9nPUj
iKjb30kXLuRRLTqBO0c2r1mj/QrWBvovxFJKXyD5anH2XKBeGmf/lJkph71tkCKu3qecRwa2SSRH
M9LiSUcTnvQzUO/fskSnuzia4X6IpzWN3nxbjF4V1YGxmFQrVp5C8TvNWFspB6Hc+kIQoSafscEE
vdCNRslWw1mKK4R8BGlgTe/QMhSk2n7VayDcqx02XmhUTi3ztGsOb4Xq8BGIote+Ssyp6CrbVOqq
gxhC2cnm9jOaIiQCZdyViFeDBnlphxkFqU5C/L57cJnxUAXCXRj5jFxkP5N4exKnVfvA4w6I52lX
39gvtwxMZ9o+wTMNF9KhmZj6KAXdLWggYXVdeDOQ8F99T0QCTIt6th+7V0XtcejHK86bGJVWfCrW
hg5Ib5hAGtFOdz8+5gdCVBJHu92gBdaBe1VVC3AhaYTIU1m8Fl9pOZr2f72TlZRM2bmOhFcMcBnN
rRqojfEvznW7cFdwGMu0CNpXnRO7Qru8ZsTawS8471NREimrkJumq+wxKSi8hUXT+pNZdJRuZNfK
+c0j7/VZkZ6KXjnYx+oveh5E18An4XrHE1VzQnHMqFgF9Ohj1R2CoGwTOPPT7Qf1GLQIg0t9qxJC
3CUY9WEeo8Q7fTqfPAnfDi5fMFK342vq7xlNaIC/SNG5HPaNu6zl1BHLUkRKYavqmvTUqOlmHdOZ
w1hlPHl+3JNtKyEv/clLjM+Q8aXlPijIR3YRdfgdE4uzsMytJ4aAEmSlmTG1u8G5HnCSjL3qcU8E
7L/9grRf/sWuZXH0ZXnr8HUphyveCPGkJfhWgP5hGCzn0O0Q3jhfrKQQzmzc2J4WdGz0QHdlfi87
eeUkVl22BaNVpyIvpdUgYh7U5IGs1f/maQ0uatnsboPcuGXafOJeSYK4+BRAfgdqNAnESdhTzLz5
0jmOxybjjYohOSEhlKLieEBkvpD3X5KJYdL8yCPgJW2b5/TTRfPq4EeYSzijIs5IiZUaKoCx+jcf
jBmz53zGgQg53/UEiJAyvQEkbmKOcEE3HFJWRD46Mdc00xunDOB5JEqO1l/HfdS9BA+8YIoL3zjE
X4RXI7fHcYnnIUyXrfkycaChH++u5LB4/waOvrVZ36m1P7g+Yz4zJdtFBVqF7uRjLX+Rysn7O2xM
6D9+5K62+6XRqD5xQauG37NgIf+BY7A/wuLQFx8GD45R54ewqkceHd4lhwyJlWFbnjolKSBX5Nke
QdeKrxi59Cn5ZsHPz5IVjoddUNiprUCUksTLkaftbvbZ+o+kDwMKb+qu4S7SLughfcUqSbFsAxlU
9lIiZBHbKlNvnfgH995M363dspX2sB9TlEAKTssrADQ4oK0FgEFu1qalSuwQnr9Sxt1M0fa5eq3O
F7Jor3N38z/vVmmYpVjViOHrQpJSfxOMrIlfemCQzU2BI/OlozFAh7XGHAlLgFpVzj093NcWPeqT
U0cfnWkIaZoI44KFBNEolCttcJBOn7HE+75G+h8XzABMlSrvbvEv89t0jz4V6diBSSjn1Sdlgq/y
FH1SwdxQ+WRGFiX2k5vWcgrelI+HLy0Qt0CS9BNbpxnEDRHi5q6WQMefF5R6XzCJd0lXVWoIfPOD
OVpvJLNMU+LjwI2rjyD4iRif+7+Ej6kSakJ9ZqjKUuYIr6nYUoczIwfZNlyN/JfrBQMkWksRFJnd
WM0f5HKRbxCgXGdsHeQcYts7bGNkURbLEL9TJZ0uNLdzd8tDqdXH11q4EgBj0D0Uw6BIQuDTS6r5
CAuLaH1tsBxv4c48ljdjhYM+1wH67NX3PlNOGl3UbqRcpJMI0S8SzN+2JMYGGgjmfZ+8uXU+jTh3
eYs4ODtru1YbNbB7F3YPUpRfXT2F/0KaxITwpprOGmmn6fLK+wje7iVWc+0Bt8+N6nyLjHFOsxkd
xwTo5ZV/vcGb4kWNx+wSPMN2hAO58rpijiAnugoykQd7hQND8RH6WOh9Vz1oWkvB9QdECn4oTn81
orQW1ns12xnFFywTBwSUtn7UG5cc90WnlVUwg4OCz6iVJ9T+eX1aGsdymCxQSIfuiyt+FsIl9cGl
afGkug1rQ/hun4fibacXvjpAUnl2w7k7uvbWUaqWSPssB1L/ophusn10V846+4RDnSpLbgY7wMAh
Meo20nbMDoGMdWeySVvwygegp4OdHX4tL8WafrWnNC1PL9USD6HDpyFKAAl6NfLFhrWK4J9rMDJQ
bsoWlDSduefXJPukOqb2bfDYGMwUA/OlptGEeB41bkNznqst1Xxlq7PWJsHIz2KvwgnqI7TR0qDZ
GENsFVv+nVMJDPUjmV5NEnHQIitZTGdiG8TloXbxe2oMEkGlELKC5mNaC9Vd5nC15jIealL6EupV
dsAfEnBPji1BQ14U0CAiCU3OLb2qIQpa54QpxRWgGdfkkZeGVv8kNnJLFDfS1i320U/TyZl7woKA
WJIWPItPo9qXXCFYx0fPakI93TtcyWo669+7B3qutxZR7nV2JcNVoc73rLrfrOOdcL4XSLN8DfB3
xefK45xfVUHdiYh3Q5aTAh74obeMa/zPgCI/mrkJ31UtqJXeRwwx8GBdwMRcccYviQQ3C2eLxhSU
o3aDgrQgP7isLEK1skVgH2e08yPl3Be7ILKd9L5BkLwU2byGHpv1F9eRmLfjFhnDexWMipT3jE31
/bpnGlzqFpofi9N7LLhFnsj2C3VkSNGz7oOk9zPClD2yktn/aVn9ui3fCV1ZA4paLuqiIkC/FdjX
9XQexjBgiCp1m7Vcr6xTLp2p/fn2/qq2jki6EY7vGqBc49fbohB6i7h7Mr60HSkH24nC4u+X1b0U
o7gSQB+Vh1mESYiS4jIF0nB1uXY2ZZR8uzOebb1Kjr0Wdtzk5XtYDBorZP2+IWB+yaqBecFB1B9O
ZHMdLvSOyYiLiqQVB+hRYF/VwwSyfAgcl8jvunloBCwc2TZsqrXd9nwvMDawLBqsqcx6mqS90dV2
zbASU+rZnri0ReTYSf0T7bgIQKeI+RPgtnhvo81/sikUSa3lCinAbOvKPF/FNE6kXW6MZh+AOzoV
Vb/NIUPBfB2G8hWiBLmiht8isTwRBXvGrMEThzVpfz66n/UF5yiSatX9Uy+HDM7pmTRc/YLzRM5Y
+iZYRsjC05exQUqAi1zta3hvkLHcR4cqB+SYrF5Wga4dHGVA1wm7/XjOcjKv7RsUkCq6qUROX2yj
7Ziiz9qLY+R1+54UVdtrPof0VlO573X1oHX9PxQPDhcjftc+zvhPaBhyCp07DRqvURf78iBQzmEK
5wD8+o1jyC+pea3voqt3g+ylci/o1de1/c0deMxP+eCQWwQ+qW9tWESO0KHsMUWQ2C/SNn8gt7nl
U/oKdZoF588PYAegBtubV2OxUqqJYAqSilZHnc+Cizx1bCMHtxT4hBVWcU7GsVHmFMGsTjZP5CD4
YBmioFVILdby1MIUYw9H+I6iwswrrMkJUYhJ26sEjLqjBwCFzWY2cGoVeUX4wi/XK7zJp12cbGiH
TLfW8E2VDwAnssWmyudA+QR/++9eJH+c4DVnMDt/x54HY7cVVKaPl+mY1tLKajK0X/Oyrzruzkyy
U9/HJUEyGG+jgRksC/0AbgblQ2H0yPaoCv0T/DH8R9Al46Xvsha6ob7+PQOsx5VVFTxVWrh860nI
vIAFE2HI/EvpCb8ZXwcvNe6pmKKwdwaGTddLeF45GgGmlxQcdNLxcta3mYJ+WVXcE4QPFLfyo+g/
vChPzqn35a0AS0+dG4IVMSMfF2qIqmIKur7cz9HB65vd+VyoYngiMsSwaHA56InbKWM0u6NhVeQr
Rf0Iavs11cbkmB9oi+RA1tzNpt45C5kkwoaodWaMW6FU+GH0I2uDsQwCN7Ul3alXyndrK0hI2zHB
5b466ymi7eEzBF/k3PM4Jae7KsYL9g1zvAG2tSj9tv5Kbh4RYjn6AyLgWtiQubyTnNiZxBhkRDhl
HbMAR3BWlMlx2IKgCDFWFKnAEhlsWznhlOuqRKnUCBUbIRNpBddJnydP2xhfQaCXl/eekjZxjh1O
orv5/R/e+x0LkupWtTo3tbpqCDEeHQ/AdoVrnac7x2fTBMF6dozn2wOjnYX7uCOvSPgGQ+aoha5+
Mo8cFuT0AEXuDSQL29VBf/K4atx13BvsHdsKcG16hXe7X5PaSUG1zZVuunagOYtHywxxw3YnElUP
2hMi9KeudAtrwaZj9nPbev1M6wIr3FXbfqkApZr395ZuKcsiLXheq8JGUdMiGxId6LHtg/9OmKcv
oVuCSBtAZKQVt5GCORnbrkx14gyDuwQzjjGCphKJii+ORdKTGV1w3z5BxvREvGOiyivoJqVVeeF9
rU4HlBvx6ew8OsfOPZBQlBlxLLuIheK/lSRsv260eWlY/e5zDuMnuhukbG6bhJjuLICMx1H4Gr+f
hnU0hmckWWEdqZSinG325eTw9lVjGR9eSEXfAQJbuHsUtyJhN08e88W87qOWNx4OJCVQAYVIsCoe
gFBMGlE3Ah6IHHjYd156IwBdz7GMxX0h+JqR5cBLQRyw045Em+n3Ploef5fYNPDHr3m2AH2eKcSO
ocNQ8HE4pUsV9qfKhWHgasbtVEItqtXvPpTlb9AKDyy//wPNTYrSU3f7fSz52zMY6v5oYaaG+cvG
YO/ItjZ+0Kwy9JVm4XkY25BR36o/eCBDgS54fHhgcHx04ILOSz2YMEyBjy6hj4vA06+oYhDKC/kF
2XEeN0Qp/nMlK7mu2bNMiXYl0aZfUBw8wGjjsoOorgaJkRk5BvlNvSnSPc01NvgediMskKVsk6dr
+EdJmnMSsJSeRmmF1VlneAQvfd4lZVWfT0tIIpYrEPGpPshDSWp9HozChB/cB4owSDNsLcOk/1zW
Gt/z9boMB5PC9/tOx1S9P35zlEEtKwfJmtBMiW1/a/tYRD7h9cSZxQ2WQol8ixOO+521AY9pIDnM
dHzmeUi2KIDwAkJ6GSvQCq43hhLB26a/cm8T2MFbqFbcBoMEEjaCc/JViTJ3YNlYbOjfxr5+fR++
NXOybxVqNqElyAiOdBKl546VC97VYDpbQTI8UwcqBR/+KXXiuxZTcNL2rKiFE4QYl0JQMZVSw+yw
q3TaF3XNy2pce/BggFU6SgffcJkKAvV2DAQTZQ1my7iJElVXwa6NSy5SW729FHZN+/APQ+/dhfOW
x8/wt3UdGGsskM5AR/Q9QeHhLEHRSmC37sI1xFsZDgaC5SVHIbSQPtEiFgi1tCAuyvoDy/JYogdI
ffu6cyfGsli1qICC1j1Eyj37ax0lcHMm7O0H1W7zNxkicGRqfiLgKarT/QQhSDMoLTJQZ78ZlzUY
2cSa/LRmP/2Ut/k4uKg6qGwlNbKntTPOEUefkzeNTwls4+OCYlhpw1VIoFZ5yAh64E0RIiQSAS5h
Tsjo45Z1Ye3J7iBIVzkRNahAyHOnXRzIrLWlCwyycMwclXBy2eYfVO/bLIebJvWOZDZYAuAUyseE
zbSgW9DcuA0IthkNxSXCCHw/31t/Kh6c8PysgO68fz8ZBgsZ/aTTDnr7Z9DLJxfocP5utWCuDArD
bT0hlw0swZHhljOeXYohJnKOixNQWYJjYw6p5u04jkKrR/JGF4k83yvGHqJ4H0DSmOpYKIUVi0gK
xYiaFv9uC6196k+Pc5o/u4eTzanuXZ9rbl3lcvFkQ0fPW5rwG7PTz4XaM0B30p1RxIXomLWSsm85
ojmPE3L9jg9ZIn4W2/xCrhM4qR/GkS2FUNlk38OH8VP+G1GbLBUlCbE6yOuhRwQJyGUZf40xqfCa
oYER671SRDhx2pVDiEWYaZfVGNggf5sMQQ25rr8pvb/Llce9EfvzwJw2w9cUVtlNM9v8sPo0e3oC
L6YLMd7Tm+5nmNL/PKKZ2+06eFIQoRuFLUmR2c1sObXDmGuNgBa0po6pz7XOvqq6jg5NIhOQ6e9z
75MPT6bJW5Ft38KPq2GHSF7gq25667jCpHLl24y3FRVQkXxHocLKZUNdbm/WWxdCScrTv8nKS6mA
pLxG4WHdHsntcxVwCS7Okx0hgDA41CftHCKV+eteytZxwjzYIeVwCti9Mrr2dt4MSnWgT7MEpu8k
qA38txDHQgff//E8p7pOjiHhlIeO8kwKsXXn05Q/yhxvKoBtR5RQUIZTeS18AjbzLsmmC5T5/RjS
GeVM61PuFbJj1Q11BoK8QTXWlU+vWwjDWCsbukOj97OSLEfo3j7con7s29rlKYt8ITt2Auf2fYCn
wK3gQ9cUx1XyLRkkQ8/dtbCim3r/tBi/I4RDxageBRmM1atbCIKNi/CenU1MnPjJ70vS2iwthOo4
soWITf1FNJFbc9KputT4UPEGaX2DVl0a6MGfCVobfw29QeVFmow+uc3aDkCtzqrUJJu4t4/diIs0
Ax8wlmBjwqKdLvLvSJjyN+uj7SxoCT9e6YGUTaeKIDT2wv1TAKFQmTs3Ujq3Eoaz6B2Paei1WT7W
rZXo+dHFXvAEQQLzwd8WzOOoe97Hsft7Gv2PV1cJhYrS2dqVaZybppix20w8vYV964RiNaNcNbzV
nZxTb4UrAcGtR3xJE7+AWnISLVckqlTxZIN6T/koqK/wTjpP43vdhpQYaAP8rK7i1hzSlgJRAJq5
Q5do4OhiUhVLO9B9k0INQ/LEno3wBLhHg4R756AhYDyH9VMaHOFDGu3h/CjSJSO3QPjsPfYpHwKe
mRRkcMiI6YYNyobg7n6A0MfVkX+S0YgFgro1PZEB4KflfjMAIvnX0g7JSSYvvHeCAPwWwT+CS91Z
rJLSGMRKineddOTwok1YNv5lO0ne1icG7Vcd0+fZkTUMIbFTYrq4qETaG1kPhMDMVCkaIr3bGIlv
TNj9a1GDNwB6amJ2FYvh0M3q7mOE1Yl+BT/UWoU28mXh/t7QLDweAZRq12Lgyi8iNo/2vAn6lbcH
vSqgiGscQJenoURAG+cJlsZ5YNHgfc95UC6/RGZXpbrM9X4tK9P03J5rgvLC69ZLQ8OS7aejjFdD
Ai/s4zG3Xg9bnh1o78g6FO6gDXt1vcxCM9xBOiHaHBfqk7GIyY75u7sjMuBRbq06qs8vMcgUfjP2
tfTF7fj+dFPTyLXpg4jmYNWyJ+/XicujX0mCV+djd0z1LzZ1Z+UJLgQaZADqORZkF6PU2y6mtcRV
31k8X/xzWbE1Pa/5AEtjSn8UQHfiypPBblJvDEdSwUuLO7WDWbxDu1v+8qPEEk44e3NaUkHPB6yy
os9NBCCYUbf99WSa18Z56kmmC3JwMfOXmtdo/exzJVZvJPuepvJBor1ZD/+DfKLsSBnhvteoymnt
5+r0kfghjd72GaLoh5bbGtbGJ5TnznACIkDUCqnalW58VzbCA8087bjSqKrlBK7sKFkxsX5Twf1b
VCf7Z3WWtcNsYSt76SWvxojEJ+tMJakYC/w/nfUnklKdIXCed7M3OsUUzREMHdrE4YcvLqYMK6wo
tRqPFjB0nv0ESCGRLV5XYVZTpxVKt/qTBPLO5ox8ZRZOO/i437Xk6fq9vhu80+NlVaaS+z97e4a2
a233udLkPz5ESCV2SMLx0+q2rOQtlQJHOBmqqh8T1J3CKAb7bFnIiENdidRF8HtMxuv79kHbV45W
N+C3OmRgZk/8CIk82G1kRM++teJfcUodzSo9LC6fEbBUgVWRETu0iC1RNXOLOPoR+0craUz3q/fU
xzMFWEOvMqtDfSgw+/hSi+rgDzcpm8p9pM0oNP5RxNxTBHfwWKF1eTxg81YHizpobRoo7i3dhaZ+
lVZBnPIHnW+WA7l+07rNUAMDhGGqjBvZfoqUB+q+31fIXWCUZm4rYKvUhPyL0zpxAPDIXii4MQf1
G3AutOQgAnPfJuVumZEEYg1hwPuGgNi8PeOYUr9E0YXsKNLtlLR2cIFT/etFaCYOQUGRUOH53NG7
9CXKQ4S6nLyvbTtRrSA0q5q0M0feDZv5U5qnKzLWm4oitXZsxljkSIXsDurP+qqt+mB4+yjjhyTY
hWdrq4GNG482Pvh82PB0BVD3806+va+AHRldcLFKsSa/yRLAlK4L2Jh0ktVLTX/SEbGW0z+8CbtC
H1ee9fG8s7kVnHyTSfnraCFkkmX82v6WvwNDH49tjcLT2P8Aeu1w3ls27MOhGlWCtebq5JA0u23p
+L+HeUZL8UwVFfcnL9LlN9D2zwCDcQOxwAywiAeRCf5OYZd+kQishvHjjcBYNIMI4y9t3zX58Cz9
/2j9TXJp54Tfi7U0SEjk0UwlD0LngTrW7yMHHnjHZ0GJEVqJ4olv8bodbv+Mhg3bmTWYhCJhGfhI
0dtCe1DABSaQR5V+0E5bs4/FXNHL3iinq+V8Z5bPC20yr06W9DTVEs3PNqmlh+tVXCNrmDPr0Sj4
lj6Ck7gjweIx8rQO9bTxHGQfWgGCoYevg09AaBkhnuLldWbq6fEtFJ146YVZAmy6ttxiSk3aHWhU
qxG8vem+9gmtNiqRYKh+lrVgFgvqo3APQe8OYLoo4Mlu+U6Cj/h8Oxu9OwGOAtthfDgpIntcu5e8
T7XcBgpjdroEleYHfQHGKHfNoxz0S8ZJXBJbAGYEFZUOEIWGoTl1OMzvHbWjknQVdUVQbFDIhltI
r0eLXcyhYDHfeTvLzoFcXFCZ9icrRwSc/GkpAGvI9c1cyXssU50xh9cJ+izZ1TZAQ/b4kuVsG12v
EH8ZQvRM/HHAwAMLszAcQ0EzFOK3MbvVCwQTbKWSWaqNkuWQC40Fc1vEMGTiNw3JE05bDu9vPhFw
8SF2QpiAKtHRnnE7D5NMfH4Yq6aBWk9N4k8qz4lcsBAGdNmpp7owAjUT4BK0u6OkDlBYp0g0OnXA
po2mUDMm0ISfY0aNMOPAPDfbks9RosgxlAu1ABjx/80dHD3yaI9lcUzglGh95hzhA7u3U+F5ETzg
zA030tfTu9Rlp41Lc8rGcMu787RFQ5cMYI/FI3i8YToCS7kRNr8M1kCLtm7V/lHdd30kf58teJxl
pvkOttQN4qhdQoVm5YxXMEpp8/kEl0sGZyNm+X+ljsYrHdDjpG4ITyrNLscrsgHlhNU99oxovTIX
YArLLpFEeYZ3n88VQGmI337yHGTfF4u+O4LrNg6aGYqQ/fsQcYPi+c5Bx4nTE7cP6CjjCeO2D6HJ
sNSvZ1jXtAAMH+YLucvCzo5+qavBui7ZqM0xJ1dXo0JiLDennNeVK7KX1Yx5ve4TyeOprUqq4LsW
0L7ErNROwBlzBWVF195hd6zVIyJmeGDhSpT2ElRG/GXxfaUAhr77lSSMGrPnVTRYCrLBOVynLb71
8UWO43XL03uyK3lxu3KvBqS+0yttR9gu55drpySUKiCI743Pvj6WSsbpgLt45ya2S7xKJQh7YS9G
q1I5OaoHFUxWUegqLJjztH5HWpEUk4lhjqp1ptRAj6mC+Rvm4gdzvxOkHQBOOL6sdOC1S2jBTc4U
6JmiMMAsdYwTPPsNZ1ToJy1R8uOO4w6yfl+GHoHKStQv7NgzAKdsGCYvgcCzgChe3Axe+wb9ICXo
iBbUTJSTPgX8VyOHWpKYN6S2opjdoZoGDhXk+THgvhMaWyti44U2rMu0qc4QZ611ErEnXQ5C9Zvb
MVfab+fWnR5ZVN+idFkzgZzSlvYx9eWK4UROX00Wav0X1UojWseK5Y0l8hqMp+l3jlkgKWZbGlVW
62tYK/mId0+fHOWw8pRLf5Bx9kQ1XUbh14aCWJQuh0z9w2AVAraOdAXNsDjfk4V+2JakwC0ynPQR
yOK+prbi8Gkmh2yN3BNECG81hh82jZmBsPaWog1d5Tx129IlV/PoWRH1b5mFFNjeozfNoM6C6vDb
YBBNo1gEvIPKGinFSksqBlzzO1DzYj5CcrJUJvGD8cdHR21l1opJcNCyKeFOvF9qKqMd0zX8i9Zv
ESrq6/sE0Quymrv+224X5+zJo4sE5bBurKPv6nv/F61oBU5BA36ySkzn2dvDsSZKhVhf9qiXaXpT
AiZHvuUQFPoO/1bGFPFPF7CwvuiOw0+3onQzspFa9A122h/dYfWbJJWeq6vQ92sIn8Icid/F9geZ
srsXAQCacQMVb7HCjXkxGH8vD79sxp29jEWVM5BaRpFEsMs2Ez6QnGGruymlpmiSlL57QhsYN+RN
rm3p2IHCcFYqHnp8WMPNZul1qBEKpg+cDIS9nNn9hoaqc5uWE72r59HKqNG+ON4ZYgN6+xKDWB+P
wjkjCU+BUnwswN2suUAW6OkNjoWIZMMESxP5O3pUzzp5lsYO8rLOxm673L/xR24iYlN1zNWMTql6
ywdBEgKYEpPXJeG8fDqs4E6dx+mp2C2fuIDVRMV19EHVmd0yroEcihmbTfrRdUku7x2vwVZwz2l1
1X8b9GjoBRiyvVTc/w2AC+dOs+qh4ThVTucHaC91uKfWlDhBP5f1ImjN5DX53dU1t1i1jbHu9CnF
ScvNbuEaL2R2GP4qauXnzLrdzazFA1EuKwrpKlFWrGdPkUdJ6EnFZzbO3k9Q1o63VhEg983VLRa0
UfKfTNrSu32UQjMOu9GAcHum7UfwAvtclcgqjWXKG+3etXjex/hrYop8a2+VtVZUJyI1vK8/nmTd
BCryQm9ihnMC7bbsClZ8mRnnh1/GYwVJ/lCV+AJyqVS4eulIH7j8kQUjgSSkwsjtISuOaiVY1ai7
AacuVdtBwPE0iT8NERoNGN7DDvZFPG2eRO4zLkJjOngEGUbM9NNwWRwbPlGyQ/6hOlk5m4kIDE/u
irJqEDxDSL38N6URmHWVRV23hiFHpQxTvWVC0pg4vQJxniz2Tpl7CKTrRx4nJuxN2IZa7ce/+Bcu
lL63WH5rSqQSvxanIG0BAYl4081E4DwqNpU5Lip5Saq9vwivTy8YMqOjI08iM9pyGFTITCrVK/k4
sGxYPmrtQ7VQtUo1G1+NultWhn12EYMafeKiclTTS/vYYZhNcCJ/SM25cku1ygqKgr5VUdDo+3/1
QVT1MrH8bIaNyi9TuHzWXGemGGEhLspi2Cc7U9Pbe/pG+FSZSCHlGAlrD9ajp5ibZDf59CISI0ge
9bsm8w9ZXucFIM5/SbKziXjBBpERA3QRw39TKTy8WYfI5lYveyerpdhDn1WYET4wLICpZh++705J
mt2eu7HpEBewRvk0CsLbRCd0w7v6xYh1p8mA4WDZcEx0CBn67Oq0zOSp9HNVXPj+rP9Tl9KuE5Ov
Dy6p5acXMAv2OOEG0YEMyCzvl1LKYkAbjETY+0P4I7OdNXZDlt3SiMRxfy+0hOeCR6xL/Sa+GMFR
rv7s9BAdmFsbjMr0RQA3RxFJgcHADKrgJfZZg+FmO81yWTpCPHsHPHGgYDdryiI3/KzftEglg0ml
DnnD7z6im5x7a4Nj83w+EYD22o1jTTcpMg32TiET6QubIQnGZ9pWn9ynamgXkPVSIMXpLyx9tRkU
S0hRMUG0NvjYuBsNbly9VFZxgpT6izS0Ns4Fz7a0ZN8xjkRUpDX229zKb5u+RjZRbGoFrgmHQsto
/1E1Bsq5BzbQnzjDa7+yVV+Ag5kG6OE06wFC3eW0j4N8JoHWl2VMilL6XeKYx98qrvsHqjYQ4fhJ
cH0XzEbc7v8okMAyz16O+9H7HPguIPpacH7ijO49RlByOuY9hQfmURS8IHMDCU6UX/Eeg/moOmYu
QKayH7LvzMKO365SnQ2Au15H63xxbgmwj6YNt/L2kEUNPWgcd1vjDXHQ62wGiviWhxw2qBLBIXQS
vIjdd/INMBAbqa9ua3a/gHC5NpANE30nrDoEydCnll07ykO3zWMEbwKS0NioRoMZPgqa1YYoAJ+4
ho87+G6xlVybhPyPWmt1VG0wWBbWrNFXDsQ36g2/MA9vWRb80OQbZYbK/EGthTJCu3CGUlk4xA4t
ecBc5ORiypPSJWjBa+AdJFe+7hMJS8w0x03dvhlUid2Z7JpJ8Jf5ymygcEVfPvNO46dG5aDajRnT
/6HE49dIp+AoY6WqJgGuNidLV66XfQeOcrCecJWS0fceCRnARuD6Nzc6W4K/zS6/NR3bbgiqAD6E
xek1HcHd8xBgcaUWNUg07TKwEjjy72f+TmNpzKdoYycjLWGclX4P7BUqqFZN0NhFz2Bf/hdCEInD
QVW6OMgC/6/S57e9kxqtIRbqiMd2ICW3nwu6PZ8w2SuR0VqdfMb4rW8skZJRB4XOSbGYJBLBecCj
T0FsEqalfSMeHF4me5xwy0v6y18G56NMCv3hBrXIF4lf6WJEmhe75OM755yx9nC7q5/b94Tg0krl
9o2MBgXmWn2l2sJGgHjSqrfzAxHwa/8WfuDLVUisbdzMwAwUE8EVPrhE8Y+DZ/wU2Xcg2MhMrqdw
QIbh/pXNvWkQyKs/94GNtWkJ4hvoa3bbItLggrHV0+TK5J4DnDwqw9XcJ2ffBo9ZPAwmWRqltcKW
lR1BoxO5686LsXnD0HGQuSamyG6vSCqGBp/W80VMthPWkam8GC4LVTNnKv38XBKYme8rwbuOdVSh
f0O8siJmLfnc7ULhA63PgC2GoSJPyoYGl7ssVqQ+LRsSmO7qlJ2vZfKvQJUJ+PUflyC8TRaYTHKP
Q8eHvlTzGNyj9LOIDVyNt5IRsEvY8qUX8OkMlZPnv9Y3C/sO/6gziHg5wedmHxQtS+6JsEiKJkJI
vt+SmCA2nyvxwNcy+KhnXHjmc79cgLvNqia8awAqDKCF6dsaTAQ4ur7xh4PSljgQxeIJHXt1qXRj
jLSzW5kIVzo5qjdaEwE5zJHYos3nmIDnJKvE+tshh5lRVIwttlxpLgkWMazExalNG6zauZwMdTBu
bDnel/lVxzepxV6Vo1BrAUZf1LZe9ZOj8CIz7DNSD//hzqMEyW6s38IeM1UB8bY0lBmh+AxnWxm+
Ieql1QsnGMrlv/JXhIqWPykX4s5jwL1Hx72AIe89BRkV3ImEjLzVIQf3o9P8oE8B61cD68hvVkWW
Ap5ZgdP/F19icKWiXG0rmCMkFv4GbF3XxjLEeuVH8hFA+Xvhc3TljTJU2MgdeeUFJTyZBTPtycHE
U/0hy0pV80zarK1y8BtuxmB5lkq42pVd9oXNpg/uu802i0d2cmc/J8XzPWO5/LMiXdb6An2bFVyc
Gl5wDiddpo8eliKnZxDkltjIJ4yM8zpgN5FYUOj1vL8s2GI04SxPaMe3ZHoOexPXuINVzMUIzsDt
xHEthA588Atu9kbVMl3+rCHU/9vRAPq8CaoKuOqnlPwppTYzMPBAw+kzdCoGebc4RQ3i9nvbCpgV
RrlPPFuKgy9IUp3Z0wPDl6bPg85WGVP4ayEfIuY0JhG8CTCSTMLOIAhLQmSKRLexOH0Vj1I6ksBT
vcBvg/A/sCeXXb46fakDQC1PoTwBdJ2Ysw1NzSwztClQ7wTqbmTHhHsWoGDWxlx6mU6Qxv+M/PoQ
8UIgOisiY5pVo7RX/m4TMZoKHdyekw/+ScUapnESb2xLNU+i/G+fAgL/3QGOkEBIYucGLdgwH70B
IkOcrsM6ATB0K1zVh/DJulEsRrsNTtdVUSbEnNc8HG+oB86eHD2P80dkI5+dhhBKKPH6hOBF5GQF
Me+sLVxwTEhwqWs/MWdkWFp3TCZP0/czSwJgdWycKP5UFKaXSfoolcaSiA5dd5/IvCY/o6mNat26
UiCWLGsy5xEAlqmb/y/95kY2md3B+/wV9ENdmSGyO2BmxsLbwEJOkxx15rD2dV6wDspcmJB4OZQZ
VongHki4eUV87wBm0d6nhr6Sf4pTFnCy+vep/2av1eZc91ZYpLneF90+iG+KVR1hjN4hXn3SFO+i
kb0g6oS9b7jYaJ+4BvR0HLYt/Itb8lTpYCBUyjkckgntE3Seg5m3kPOrwZoFE2uCzYADkTXerqTA
J5nv+zN89knC5K+cM5AIQ9uYaMMJf6b1kj521HR7AUzKi3JQEeIRO1QYt3plWtFRIcxYzhop2QKQ
1cH7g1oh7A8uSnBMoDWjTjCEXjLsmYQ+hA4ndR4zJcJwfWlkSsUl5cfWOtbqSnDS8RnhDbd9wctg
A63sgLpzWbow9JzRDGCPvaSiA2JAiNGsVvRi7ImD3dbO5m2aixYdlFTUAT9ZgYN3V1sdKYc72Srp
C8ZzlTGJO/ehYVskKyVaV7+DKijOawnv3q5ccRRiheZO9SAwdV0JIDkPruhgQCdWxhXXrKkkEKoA
ahMWUfcOtb+g45EYkt7vh2FrKySJ2ciJ6pnASn5BcscvPzV4rKYNg/u6mRVgfaS/eHsDGFiXq49S
wlszm2ZQZQB1ABRBXzcFlsmj+U4ULHjAvoDdRL7PDHSkZSCA4XbxdqiqBnSx2kCC+6nrki8hwFWp
vCVLgl/HlKM4Vukmp65MNG9C7Qxgypioq0kkZU295KhVKXM2qqpuSSmdmD/3oWd6PE4M6R9uVu7l
RInZqFNmZkye+rqvTqjVyJ+VdK0X3Os0YDvxQi0gzyVlM8rRrn4TtB3QK/CqzjZP0dCnlwhQ9o5w
+zjLIak7eVxq7IeuCjD0/qztZ1R/sJ25lFj5aU/SMzyDEvu6YZ7MzDGXVzCcBGrB6psFBs3pEMnn
GivKGILc1tubQVlIzzjAvNivwLC7owy5LaaylWqxo6YqhWATe8uRWEJvl9YU/fjV8nZzylR+KQLV
oeKiOl3rnSR361K7g5n13/5shUmnihbaw3v6Swllz5AoeVXrbP31S0f5ajZwx6fkhAw3JJJxV1/q
/9gEozHUim8By8IuD+HwsmDcqfow8Of+6wl4p8sHnLrd6UPrlGq06/Ha6v809Dcx7meonywM+Lsz
3YARxEvgQs4xKd/QxPHE+qXtPna65hIEByjpEINLX/7wFWwmkTr5EUe9lFYo5Asx2ydNHNws8FV9
VpBXwXTrJJF5ShwEYUOYx5GAWILaodued75NN4pmIcJqCdaFBUpBMziK4Z1r/b4pOjpVbKqM1eE0
upapCnVC+x5F5zBIG/xp2DQseUT7y5HBO/jdwUSdCbAtvnD2TVEBt/Jzd2S+bH4ilF9I0R6SI7Vv
bx/XP0jAr77I/7fvV/bSV2z7uDvSAiZTtLjNsBBM4uIxK6Ut80g7AuUx/Eqozgb9hfUsKHpT061N
JgHrhzaf2V0zNIqhWNBiTkxQP1kyOdQZCiFBZu4mJQfLpJ7zpwIr48b0zbmdI54L6SGeQr3xGBMQ
t3JC1eyDQXrr+m3IQcPc/QeW2s7VwZilK9gxzK+mYaeAkSX//1KFzX5gvvgHB7yV+jPyYw+QmNZf
PQW+aMJwP6nlXthP+sG3mMM8m0T36dXnF4PL3v8SDXL2bkzbAFt5LbCiLjoHTDZQcQokYtTZz8AP
7XMzpZL89VUBLpnQTDC3M5s+dFpQnPFOfdT3CcC+0ZhVsRmMwlSvzOnAyORDxFMgrIgiB6clknbS
HSaE8Xrxl4xlOSiDEz4jN7Qtc8TEwgEpG4xbGHgeN5luV7it2YTwUmHCk+Rsl+mjoZXTxOgRf31O
wN3e6HnjX6kYmgwpeDdgTN7gCaQ4GiYiZVaWaUjP0gqO2EqWE4LjIBngICi9/J4lItKsdtcfFDWx
3xsU2anenZIMTAbSvV7pe9qx4RfiXU6LnjTO0DlWRs1Ln7DEnGWZM5+sy5UU6dQN0er12eay04N3
Yx2bKBnPjehWGhIQiVdqcVOC9Ce1fiL5L1/HFh4Uy3aa7s3rrdcx6KF554yjkfyo1jHiDsUkE1kY
GEvfubmO+E0XVWFB+EezydIN81mMzjt6R3j8lyWacM9I8bsjoLbZ//Nvb7FdzTojgH13do0GhLUl
o++SLcaRcHh31f5Rhqhoc7VmqlFB8rRVHjGvjn6ns/Blm8JcE6XfWHDOlPIv9IG6xJv7d0X8BEPb
0bUChtCpKMEoesj1USB4eGKqvshK0YWozTb0VG+mzP56NsdeCCE1qAwfhvGHdsAFPD85CThAp60Z
VTiajPcoF/GSthhiPXC6lhJ7uQd3JeW5BLVJauYBNURb7WG1G6f9CVZ4utu0neHU1O5oXBwcagzt
Nnz8gFiWzA3/X4pwWl53+I/7Mksn+kHWIfT9nPK0a19GAdXY+UJ2a9oJnVelh5Y60uaSfop6h2qd
9NUL6Btpx+lzg3mLHT5kJZ8jPoxLJCfRfMcG+ulyocNilq8iE95xpA91OmyiojzK/h59zA9DKYWH
kL/6gySE2mMjWE+tgDxOvr4BVd33/xypcp1+7piTFDZMJcIexxAJ8jsnWAur9O8kYL16wAJhss4T
23cjMDhJn7GeZKqW5KimNEnmkStmd8jzVj+A9u5c96zHFXxwpRhQ1WuHH1BJCCjasLCECQCNRSGp
fWmkPqBC1+EsflrscWpgoM4h9BCM8yf8a7BU4ayuZylyDW162GFOIlpGd6ibi32JXVIUS8ze59x0
l8uHco8R0A+m/iLqF5il927HwDjsgde+eWxl2QFJeOMqWClFEVJs4QE/jCmkGm9gGN59qRExjoED
PIrknVcfBUt9EpvnTjs/v2p2BEbGy7BZQi+S13ZoAyPCltSiTGuRVM+QMBBGdD2IfB4tZBawrcKp
asDK/fnF/7Iu59grJ6CWy40qvt1onmJjxknnLk/52m32ztXl6F7vYHAhkGp++iRwC89ND7VmunWG
NVpuTvwvGpxmC0t1KhKZZTBt3SArQl9Y05qbssWreyxili8rAnpCTTvLVN/OTDdjLqR+L457g7MN
5dHaKwrkC7/v9knSKOhqKKRxBF0QrGF07hcoRWtMN8gxA3dr9dQpXLR7H5AvOL+ydGvPHPI0mfbR
T8P0i8dCPvHhMYjE/OXJ+JO1VCLWQhT606G8iNIZEU/gt7dSSrK3esqjU6gDp6znAOhz1UIvqyIk
wwRds48RuxQSTyS4QsGt7xilK5LjzYjbm/IS0yUIilP7xZtovEJFljEioWhraYBCwH8RL2NNx8eh
F4EkKcxFRPEJA9pHY+AyxJipxiFXo9FOZNyrqyDnHRqZysozKCA5n4tG4R2/ntWBY8mzdH7wQErl
xued/S8lKUqjVEpA/adIK1b8t6WIBVVLSPH/jvWjhcWomJbvL3O/MveVbPMqhvjN94R3idUgyE0B
ds3lMuYXPmVylk9eGrUWZ8cL3A8kcv+w3jeqPFrWe2LrZG37JOIfAB9geocHUVaw8bwaS6a/AEOj
uGo75Horq7bW67LfSsnwBsyPxYecOeDOQV/p8jf28tAj3B9gEBwBHMtKJowVsVzMU6q5WcGT9Pmu
5HoPLWT1VYOqZWkMGEMohljYAyv+sdPVVuVAmkE07cyDE6hFgactbY+P1DfCLiGo1FTeWR172P81
Gu5971odg0FnySjDqi+dx8UWlYtG8HdwZCqmn+9g/QrLDCx1tSaK2kXBvYZUXm5b5qJU4NMPbGKm
F9oOF5+OJLz7XxI/QpdwXkZUC0jiyzvBUDJ+4jPEKIEOwpM3njMv3UwGlG7dLMx91x3Lla50SS1d
Ia3Rckxg4jfPFPpOZr0wc8yhWjeCozPBjII6NiNiAtPvht4MAs1XRYrYxRSq+BUDVNb1+0ju6Tsu
cecMZuPuWSB8waAB0yK0OqVwapL1uiNKqeqWQOOoRm3LNRRrwbvn1HF60QSh3qguzYG0Shrjd+vX
oJPNbM4bO8LHaRTdwz+9AoE65A7CBkdHWIBUv6uzxl9GhQKIyZVP29fll4Pgk79wLwW/nlVIH/B6
UjxA+O+QlD1aVKKhbPCq/H+2kuL8m/NBRiggDKT25AWtWqlT0TafiMgnOpvr1brGy6YSwpxmibs+
d5ANEzZjEIBtodFSljHIoSzofYpsCDLAWQSwplMt9T8m9Nl1PJzQOMxY3W0n7slRW5N0pSvTEuPp
09ZjwcaLS/iSvMm8wlUG4tdy2O+EQNqn0weh2OpfCcN9d0YF62hYcMsmXCBasmWptMf+Q1BbvD1D
m1+9BWMWx6jh0pu4KUnQ333hiztfVPMl59jeYNWE+2ojGdyA/+y0Js8jPu0lvXgenVViQ8E6wpD7
O7jead6BFk3a/MJYFAXuz+Phcsmz3T+JNT0BrV0EyCNDlLB/88yPoDZrVOobtZagiaCqys29mrfJ
rkjxPyXsvzOjmy08C5zOqj7uqM2wwhtDc/fU6C8XZczAvyTGnmydiRH7o5AuKBwGGq6MAeV5x9Ou
CXGkWl0v5r+l1E4EFLCynh3QX5G5c6H1m6nmM1FPrWi9EktdHjHE/A8sfD9BRi/2ImYcy7w2DtBk
Qp/5rXBEaS7PuM2tC945CSjodPjVXyIy/B4w8geDPWAENJ1n55APAVFKKXd7EtYfzTI/KgmJa9aW
nTSxV0DvDC4hMoy5K5+N15YNmY6z1MrmoyGT7DuHU0H+dmxFjBV5SMyB4gx9BuNf92xrBEiJEUrx
r3g+0LPAlSrd9y7TyLDxgaVop6xBRDX1nrdWLw6sS+4/gHC/Syh3oNgVEljlRHGIxhs/nYuV3ZM5
vrfkB9j6zj7p0bw6xxFccZc5wMFEm8cYZ0cx9h7XeGXrzUfzHIj1nugmP2hGIUXnqCLHHdZP1yqn
mK5OkfFWgOi1CadlUqrDhpBCenoMyYZiqyglL7uP9wReUEumZT5E/WqDOYELjunoJSWgCJJKcbWw
R5AwEsZmThkOOn7OoSeWwZoPqT7rLNdeYbLSdzecagXZ0HKOT/Vp8lV6b9nrm1x4GLZxfeBg7oRp
01S409yrlXry23rsEjtmbrq2p7m42nODz2N3x+ccLCLCqtxoryWRcrfHX2SIlxUGi3IV7zDnPCeM
TvcNP6q6LOkZTeVlvAYSvEK2ZRn9xmE9z7JMolTkwpKvIMEEm53XE5Rx96U3qNnpxAQNwRkuZ+h9
FPa+qU6aGBQ6aMqS0DCJRjtwvr/5d1ImLgzSzZ1Cf1lSiwOop7stahczMIcL/gMNGWXLSywFxO61
fHPNZZGGAFcMol2Ms8fQZ2HyAy9+lOACWWXginu0gBSBonpj7zdLLhYOoDczsKRIQjXdKvkn+fl8
Ksv2vrXbbpZCseCSWE6YFJhL29lXW/KSH34wZl44VDAIJPwOVH4jBJKMfaT+3mnClM3vRu95vvxp
rjdTJ7/e03AP5IHu+wksHsT/lA7kdVEDpU5HXWe3b90mrqZLigpCf4nM490jQfmV4xN4cuno14n/
rmojEJpsdmPNeBCrxa8XaVBVQR2pstpHqMc/Ox+r2oK7z3fXPMQIib6VjYHRmytPa8BUxWmd2b7G
9WM60knx41EB57uVt0X/AAcWquKCfZ+uj5bqddz9Y0fPnIPNGqfhBh7+TNiA+Yk774rdBPGAWTRq
SAd6zWms7rRmnP8biTMvtk0KW/biZRCm6Y+A9O4f6s9Oj3W7/jQQfp2Ha5ZGuKI6ph1r62UaWBBG
pmxlQLVs6/moEGu95iOH8/FiHbO/xhVjLdGtWgREBM1QTEVVErOq6pkNmZpqkHzwbswEt12ADrWz
I1ambsE4obeLiVVEsCLzTWx9jN3ajhkUI07APWrsZJngx8dU1kZIC6D9EumdbbENPKu0NHIkiJjF
YGoUUEzDmwRseWZeARteJZzByx41kas88mpJ3FjdeMP+Pe22so/p4vEVatwrZUPnFJz3OA58H5ql
O6pYAzb2yMO1uTUUPdjGUBk1h4GuDlmg+yWkAUlVAK6re/n5TMqt+LNssBrugrT64+GGpUIRR+EI
ggtifjSZMFZiN99b2H3FVbTQTh3iBbmP23x6T0EbXCm1rW8FDcPyiyA5wVcJvOmVbeTZo14BM4V8
is9xav++8t+0HBitbaxzgOJYJZlCvFYlXwXwKkvLhdQDEGsihdsXnlPCgCyo/5ZP2nZfl2KQ/Awp
IfR/Lry+BQpbTWvd9nMi3hfieAktMzkv9U0pLj/Bc1GK3mLlfb8aO+p6NDwFj8Be7tDTNnyGIryY
2UQrXPXqGjzsmpJmzoE1HY1fkZqOcOgBKA+pCPuPcDckaknFpazs91PtUA6KD8Lc2QQOscURlgaz
XFdPiUaV/HiCADv4YvbXrjG8mqmLYwgNq8Z8GrPg81brCk/P4A5Zc3o2ZVB657rvODzFkvEwLP4c
ebxR2aoFDq9g1E/Ho622qbBA7ipYUZ1vSQhyi2mRcIl4oRUZXaSM/sG7uyQltdCDKmxvjHB13RDI
YpAFHsNuR8kosVdic3DcCSQueawgjdEaxnECmHLSL3gzAhUZTkiDW8ve1jTISSrKGL8xSvp1DKcn
wd008PTHAGbLwDkDAzGghmwa8nBK4nH56+ynP1l65B6Xm9FZrSIoyUjnFKu0gon43fMOA8X6Garp
mBmK99lBqtIanGaglyQMEC9EtDVz7czeY9ia7X9gCq062USKh0n+2yL+zWZO7uz+jl84xaEgB/Jk
KE6JZhDjCszpvH/XP3uYIhfYO6zVwvttOizhW8Gq87sDpVa6WeuZTylzXE+RP1hTrncGgPhBML0K
bOzpVhTGpXy+AMDmV5KlXO0vfedWoFhI/fa6yq4J6lAqkJ1Lmbmi5C+b9qRUzjVEd4X178S+0q+O
v9YRQ4Nwj6HDRqiqEczhnSWz1z2+vD7ZNkyTRdm2jmkmwQSzvCJwcK05OfRQD8q6F1c/kyf09G3t
1AYXq9JLwGExjEgOiARd8wrzZsSIeo76rGvAa/c9k1e1ZopA89xfw5I+/21FqeJGUOnHVU8xZtoK
xuH2qpk5jWGdEVr4AZeW/OWBnVxA31T8QWUy4jZShfKnvT8974GFmLwWFxT3tJcFlgll5B2EJ8qE
Yv4t9xtls/qsiyTzCOAinUTrukFw0iUFBi4xRwdLEPc1x4ZmuJ6h2Ag6mv2fvyKnW4ZXH2W2w1Ax
pIw/lXgaGJNcFzTl7K2zPQoGAi02/jUO4UDrr29lhRRvZXVoan+ExoOcxnEuQjYlCS0agJyNdI0v
sRcK9lIPYwvPS2Q//EkO0LZkMnWdA7+1EJASA1ZxZjcNdv2AXzjTGUPllGdD/ah9mUYbBEIlILXN
Ntl9dapiseHzW0oT5LxMKOTkUCvEV+cFxWz6oz3NQBMeizHzJazOpxWaXaRax+vIjgUsA453c4Hg
7tSxwxcNhWOUmsCk7Es0Sy2ag9FSe2KTJ31Ii1y+xMm8ZnVuJk2QHJsLg7JzmzXd6tR7V5WH90oU
HykC+J4o19O1xQMZZx6ecWLt2vEu1uI8nBZhfk/qRqPGglZa5Iyf0v1eoPq+umf8xQ19fqYT2sLJ
VnBEwv43XA5ATQftpZ19BaOynuURo75g7qUUMKI7Gs7EjHhhDj4m1hltv3oFtCFO2gAMQJ3PxNar
0Yx0Cl11rovsaWYRdDIdhorsMmtNSuGfuiZUwmIuGQpcEFKGfDjKb23qgSx+FQNavA1yNp/ls3QU
tEh2gNH0Of7JL587b7t7HC++wGeQp9kshK/5GW5J95bjdbQAWphpd8TJe3C6+alwJRIf19fQSRr+
dqr8dCbgI/1er321eRuvHodxeRPSR1z2y4uKHOy40h0rV4PN3Z3wJgkRShcQzXMV/AApFpiMl5rb
A8ol5cWFhT7UtpqwqlxrlD05JhSAnPM73St8lYuWrrWKWJT+aUOGYn0Uv73hRiaBpF5Kl53Ba+39
INW6Cchblt/KeC0sEj5PgTZj19HtSW9blAHMu7ZmYWILvaI4j/OjdLG4iZFmcJPJ+/RzQf1+Zd1y
9iPW8Fpx0q3ND7XBs8N5JUAERus/EelVD5MiZN3svyOhc/KkatcqwvhwdRCcL1GjCSlPMzM+VWqL
cFEuJZQdoXH2OYfiBJWe6wXJpq12KTZFVanReqPg+kuEJmIbz4ddmyhvVBrNYZK7FPpdVa2Ziwll
eOTjavypshz/i9tvn+8TtECgZyBBCaMc1hONbYKaSWqggE4jdsa0rGlxcEwelNu6wry7ml/ftXiJ
ovHgx+7lz4cV4H+Yo1KU2SH5KTtzRzqosO98nVwdT4QRDHHL4vp8EKSVrzul/316TERr+V83KoSb
OOy+E6GoIf0Pt31eDsdZAJ8KLP9/VPCLc4FHhJhobbuspkuPkrFb6Y4I7mgyyVp++xWANlD1S03Q
ICtsQAMB7LIE82ToAKuspmkVAU4orgeFN/WvgMMjdkbncM05MgkTxpQDXV4DWWMmn3iwHrBUhsA+
nSU9qu/blKcPdMHLevdeqQ48inbxcD2YxWU52Iw7+x7Brq2+ZEO8ZmAO9GpnwKvkVesrvfJ6XuXZ
4ty/t7/+zKgYLa+bIRGIcMPqa9/sM685D6ePB8SyfrAUrXUB0JK6eCa0BtLmaVuL61bJFleiIHLO
6FD2P8dvsyrjONxsxi/bdL+W95+IzWq+dUjTNX5132JHUQe6WdmCg7+cf5JZ7cMh6cDS61NxL721
LvvE7RbXPcGd5sveM/4v1s3GXm1UN2VXcnHwqqW7me2ANPWOOeJ5UUM6hjsVQ19PxE1J/aLO+qgP
emZpV4UGC4Q/OwsU4IeqYskbWdbrCkVil7doYqhiu/2+I7ZmCFkWbYRrQBe4H98d7Pf0lSajssMO
yGp76c+jipkwhptIpdBPM728sWMLtoVCNsz5VyKlIz42JQgGghsfkJQZo70kIHCYPfB6Z/GZCexM
8nnH1Cf1t2S2jTirwOdilkDXW9JUKmn1HasoeCkswsrkcY4CgsU/K6/uv/fALBgqKuYdpptLJnlw
Usk30IMDA8lt5q6U4WJAyTUslpl8CGWoFfcNtqYc9KqpVTCoAw+32iJPZ4R5QjtZf0QNOWU3j859
4AOFz/kVqT+C8p2g8kEDbw3qGIuQm/WvThv96ZkOexkD4dtMb5qGdeh0Uu70efOAeUP3gvui+fe3
IGWjyC0vRAqH3Srh3f61VxRWEka3NvYlU25u3OFKp80672pWhmFL7TOT991rH8VtMA93qOxxaPNP
sT7WNh+wDqKzahrVtFAfi91VIKkc/1oLlwXVnM5dbrBYjMvUBKuSZ5tm2kKOB4lKfPu/z7Cglf0X
hpU6ev7JTtvcokpWkFH3FaK+rK7sPHKpAWGj6df7QhMSDhZiwsjlzpAfybEJBvPyZkoGmlEEF3P8
cKW74/NXeRSHgGIGusVDHk+RaZcQLcnrTUnGDZVftHrBdsdfaeZ1hMj7HK/IKyvBh2rs0SSyD4RE
1hiLJ06wmjGMvL+h1gu4fd66FNtY+upt6GM0DW6w9jpgGOYlsLDI1liJBzdi/Z8S7rC+iUpT/OKY
asiCTPtpQhy+PRzM7tI7iQ3oDcZT2l6G1zhX7xg1yk8O61YsY3608Sl1LbozIXDJnuLBO7gJp9IL
uHJOpy6kK3s8mwfcT+y9mjQ1Z0jP/bD3nfx7oJPxQnBEOnCBwvelthxGW1KNB/I9AHDicSe60HKr
PKOejPtXT4HGLaCP3amz4WIoWxfdPuZwC5Fx0VpRJ3XR/YGIBfqIb80XCm62ZB/vrm4gVKcAobrb
2cIQ5AMGi2CADpSrTQwvTrzmOvS2kwHW12dxAANNPhDC486uEqlcmJ4z8ZF7jlGQqaAQiUq3R+wl
1Ygoqg+BV/Yj9Q8Pk0sATcR+CWyg3fUfh1CVxAaFol6m2Zdx1VpNL95LpSQHNTynKXUcaZlRo5HQ
02S2MWimNXR2/CSyzAWzgo4aAsBfKsF0A2rxrHXWfHEhT9dxFM4KqdvIOAT7lg6dJ1lLGWnfATUC
ey+9ffV7Tzs206prgbJ02WlH9FfYS4+Z0ypsZ8sLgZ8NiE4K47/TaAk9psgPlDYOxwNWfN4pb2gB
Ay0joEkCb2YGPQTj1VnY1gC+Sr3Z8vwiIkXf1j3oZgtIzteoKvTsHu98V7XkqJjmOkiqo3EuWj42
Nzo2spWzbMqVN5UvgJrk5zyo/sLCoJLqNY03ojUE//jFDJnQ9yrogMIqWLShZt/zlXxeOobT+J+b
aSH0YoH9bnAYdxfHmcIyTK9Zb/D76Z0UUtzfFLt97udBOG9cDSG6Cq3m0Rx7ojG2ftw/g0A8eliB
a6VdwQmdcgqEQSoiVxr1Do4X3n6rc1+N9drGaH9fsgvdaf64l932muxx7DEH/rldnk+Hstly3+9w
19fYgFQBJvx7ylkOgaGRlfWWo4+/Yo+Pnbpn/A8QJAopxRhNbXGetRvORdzCFeWdk5rFIvXH2nbx
v9UU+2O3hvMjsNwW9ZpAg00LwU5FR5ZUwaWzfJcSdj+XL8Idgslnh5hBcWy/SvnsUeMyVaPgujHa
x4N/mC73LyFEgO1C4KqDI1epjeBL+LFtM0PjHIeEw/1sPBN3zAKuJCcq67j6HSMFfD+JT8tmylrq
s3GCV9dwr3qR/J0WdxziFdWoO64tjBAqG2OBABrlfOUcQNT5sOtEmIbjSTE2vv03VBchJ4n62Ciy
JcO1dcoBelNsOh/lLC01cfzYg5IRtOTqS2q5Ln6vEmlp8goP/NzRlhCJeaBhVLufg11QlQjf3QOB
YSvx1Q4dYVfWcbmwRoH5EtHXzgybZRX7ND/LEEPqm+qcAyCQ55nDQrlfFpL21Q6uRX7zPBTrcGzK
agLSfPRNCuRnfUnJpc9ACEHjzlnZcvB3nNSlQouu6QymDOk/n4keqdC7R4ZVABaj6SNGm4QDwaMw
x1IAXlF67NcqJ474gey1AJQWfF03+y1x+HIOrxH9yK1s9+WJHdTnKoeUISXZc8G+Nu/Whe06yWl3
+2qXsUW5nFPIk8zLIZsdybBuaM2fApAOnV7C8LR6l+2A8demM9Jv97o2mq75fcCfoc1zF3V2ZLpb
Ha+aXhKvM86WX0QxELU4Xt07ELE9qESlMiK1Tn6q7/rmW+jqsPzbaYGOgt6CIuYOBQYKT8W2LvbO
JOAzpVZ8WmP9qee8Z45ZXh6QeVLSJZQDbiVJXCjB2qt7jEdkyO+LMZBnALeqWZBxedO4kAgtS2JY
/+CfqPJYEJF1MfxepycDlcfVrVdTQ+E6OxQkdfO++PWLMRllt/Q0/Rgohk2u9k6Kw+yU0xLFVOPh
ojBtssFxk9w5sVy7xKNBDZYJMhkQ01oo0QTe5YZghlO9ZXrORViZOCnhuIJn4eZ9rmGZrZ359/um
gmj44JSFvVC9qZY6jI3ZrSVOTubO9w9xxWq3qEE4l5ZzYX1YAqleKDBcW2J6bnCUoyB2Xub6oiW5
xlT7Zj8Sql0ERcUHoq9Jrbhvm3HoOkeIWbD9zznQqMlGdElmc0qUelgS+Vto3YnamyfF9JFBtjw5
v6ya2V/NKUQwmFFscw3ofpy6y+GziTfqGx1Wnp2PM1xRDrrvM7xOfvoF/6cU/WU/xd2x0NI40KIt
HrfRzVuCjPeQYZyWku8aqPD/Esn8T7yw72YDeZw9kWqKg7F1kK/4SS5gkiNkDAwyq8arfAnJAPaQ
8BonbOnR//93oP6TBY+BJVv6SbibtHVwCP8C4wTkhmWF+agOi6Ij3BG+wPN9Zmed31Ky78ezc2v6
HQa+jwDeye3CThzvcrbZXWYQ0alZnkuU3KCfDxRZOST7COuMUNHgcgRwDBCNPR5GOeO9YTHYaOUy
00B7RK3c4urJOQHOF3JJqS2FMPqMM5QvvGP+oJ+jLRz6hPvzBROMKO8LySsyR26J8U/tSEMC1Na8
T3+zhnZhMZ8Vb809sGlkdytYCkPV+0+Wu3493/sOqHpIwlpeht6Gokancp0R0yswTGL+xyIb0/A4
gPasDxREBxznwyJVpKDxFN0+64Ixfd1VFQAszFwUgMe1y0MCCzQzfOCeHC9Oo9/ndud65pV3xey/
58EmmuVVwDK02CciWZcNDUMo2ZLWMKZ38+CUe4FgMca1YU5/WqmUUHsCcOPKsxZof7o27W2/rKdw
ZfC8OycSAOFjjy+NqKljTjR9zPF+S9Qd+SfalovuIu7BshBuAs378gcN9d77iwS/v+06zVM7/TpR
lWTmNu8bjG1Z71zy57tIyQ6v8PBmise90kQPxN7WrybP5u8zTHqt3d0YAG/WVvxUwHXU0XCEZdWw
H2ZeJ/vvxhQJKOkvHXKmHHmh8iO1MfkLtbLAQWzsnTk8gaEsOX0e4tlrefIIlJ1pcnkoY8WWQPmv
KBN13WISFQULBuq2HJ4O+bzgPu6UxTvfp3ZZX5iD7G96xA+a8xx9woNgu/SJtaupEXCFSit4aCaA
ZFGzLvQj2Um3YpcDRcRIbr/YeBzk5LE+4Z430wNFJylcCh78DO825ZYWt9OcaYDQqSBrnQ5W7Fr5
GkQtaesJNX7eUXWy7lLULf+pIJWLXRAOmtq9RFSA9HDbEXkJif5I1AOaziNWzHh7vWeqkxCWaUrF
KHtSGnnXnZxxUsuWz5nb22BDzDvKyTyZBewGLn0qmr5Hrfd3KYpJIOEyWv7Dpe7q0+w/h8RpE3sB
0B+BjEvbTN81LPH0fIe51IMP85u5c6sVj3BHu92GBzYApAXprlQb4nH6jxi4mW9JOK5MeW0ydsxi
WLESBpZDf58TfQEOsssTbNmHuQpMv68/t8MMwXmlkRM8/bp4bBz1d4uSXfrC002oWk2lqKJJf5Db
m0b59OUTXq/8C6NqsJX8Wdtw/4Aj/goFm3F8EaKOwkFK+ElKHik2CWESToGEZJKmOEbzgvPljtmX
QDXBmNj685Y1DgI0PT7unVH4DShxX5lpYP+i5aIfCetalJiWPJDTMl8L+QuQhhmDgA0IK1m6sBf7
sfGCPDeVEn+IMyljL9wMWs1OGbbmoOnNg478tQCwmXyi9lSABsxNwvZgLGNObiDlMlH11NsI1ubJ
a4Y/qWoXjdRVFcBajzLKgSLIiXv9Fg10YOcErcIahBVaxiKhGr4rSPIV9b+1FQXyWVJd5RMGb7o9
O3EjR/sbkXKL/xrEve48RBwxi8+L9Xq9vXucjHSuzaKeE9fJ2GRu7xhpGjzCX6UTwXy6Wvm8DurQ
+JA+nA42XanVhQXKHZxXwo+EYwS+VFV5SyiA9dG4y1c8Hs4EmzO3ZuLxoWxYoUlneTHSyJ8JbjuZ
QFPrLa/FJ9rfJd4QOa1JfpB+00gSDKORJT9KE8ftVGl7z80k7C9cQIOHOXwnW0Wtbu77SUuIqcya
vJKbeJ+WFCSoauUjKvvqr2dHC0r3tlXoYmZaqfcUT7NdWv6Z+W2bIPPHrgJMszyZXMTLl4Z3GOWq
BUrD+En1T/DgOLtZ6Gs2zyT9gxfDcUiiJS/NqUXbqpw40WoejPJC7vEy2KCD16tZIX6ofoHFfi5U
mQor8b70k3iCnSZnHt+UXBNUHd9SnlTBuTGDrt0hyTqNZnkLeHYg0CO83K5ekTabISdbYi+i/YeO
AmLEt+fdFPjGRTxKAbhfp/jI2anAYfup9isYRNq/MWOhPYdn/NuZquYpJp7PIatlMVBmXA38gaCg
dN54m/KqWSyJacsnYNPZ8qnSzg3VMndHjKzJT4LwYcv24hqiQpfzZrOs03H3kObNR5WRTcu6BTY8
1cVuFtmdiunQnnopjRN2kC+TewbvowXsMgMipIk2pWmdojNRv5aZIxRPtyhaskLoBqJny0JtBivf
KHSLak0BLm6ZIBZSU6dL8UXQNPhiHbuLq35KCF8ENlv3U1srddS2vti17AIntyrqq+3OqS6+K512
SV9j7aCve9fHWlxX9dRsa+7Fmf1YahwvDv+T98p82tai8H7LIBSWtXxtvgFackbCeDWAokj/CYwi
+a6CritYutTOrHJ3LNRPgHi4gJY/kqz2kwS6ta+yYXUhisq2NnnkdJRY2xB0siXz5kWGG5jAq+Ew
2i2AuH7GgrEVnqj2tIvcMvsjCjhACS9U63lxvbDXqWrw2vfSRhnujO/OnPHfARxyqiLmn+fwlHdI
cMAXkMvdrJosBN0z5tCRagCHbIFIF8cPj87qef42OXofGSJ5ImTowhxOoIfmR11rigOv2ZAStih8
WPs/rYAuIblGs9MopUH5PxPdBVwW00UkGcX9ErdhdKj66R/pU1EG2qnvq6J+90JJBqQIcsiTsiV2
p444caugTtND/ZliUk2ImoMiz/E1X+AqGz4xLmU7LUGU34fksgqx2p60/avOfLFDZTQwkHMCgLHQ
Qa4GOc0b2JOpfE4onuCTt7K0XwWuqkjC6XGUJh6dmL8O9Z/5GjdqDi8VmC2yQWDBnEZuNFx2o2BY
hO1PsCf6PPtUmRBZpX9bBTJ+pyQoATyIzyCICsl6At3F8yF7gAAZLt3tdMH4BALcgxmtMIeBi6Fy
SZwq14s6vOLKa5JADDRI7rqOgndgroGjcRDM/ipNhIMrLhDmWxNhuRQ3mDzsVTEfzwMfwx8lVkMB
T3dI4SYdNc1CQUelpuDnmmBizNnVPAYs7opbJ1GPMMOYhyBez7MI5pPTHWJtX5vJ9HlA3/VFhDbI
GQy78dPclUgW2FvgJKHhlAgiBLZjk6YBKzT0apmK3jlTmakcwa4eAR+DSLRHUDGT5tvcvTa8rnvk
4HazDeFyfo1lqqkjI4MdNfpgjaUTxx0zHdlWr2q1IKC77109/KZ9MYlLCUvP/gocO5dKPCt5HWW0
TYIBOj87ugOCIzX7wciWAgzPH4AttucVJxLfdpXYnlIRSfrExjl5fWiAOdpDwZjhp2DUJXYm56z5
z4yjczuzPivqJV+w7YFG+kNxfS7mTXthm0U1WUg5wmd82BbD7xMXq51BZCBwMcJJuyBhMe+FR19d
ilmjUf+OEa4zqU6gmLxasBtYXfrYn6LFD34JzojzWz51CJQ1fIxTd+X2rGQVfpstRTv4TBn0KCVg
eHT6yU+PKgmIl0cboA7aPX3ppasUEcghDnCRk5S7VPxv1bQTxy7N8SkqTUI02LmwPuzL6dMWiHqs
o2lZfE9ajd589H/n7pOptJlDQTgTza/hAfBEkbfWxpmbw1EOTpYBp582MQux48F0mKOEpwOJyA8j
WUPru29XSurueVApzWTprj71a3s2BmfqhgVO/8JQn1v2fKb//zbM3XHR2WEWzNv+aVFkMmJJ9fR/
km3bV5dOh0xEmAEYYjFhgMkYpdB03Eo6szBtkYy9/NU025sLyilA0bJNmqZodLJ6etZabbGsiEnF
0nxB6oPv9Tiwv2N1oxC8ukBjyxkmtST+VG91wJGjeZE2dy/0w6e3BKYDq57iwiMQ4KiybSEvW40j
05Yg8NXAGmrdBRJdeYnHT35Y6zIF1avnxfChPGu95OtGpRJmyxByRVxIr/ZyN7PYwmrn9/fhAc0y
hB17x9BheglMG5oR9tzJ7dy18195Srt7tq2lSmxBiSSPu50BhYITMqJeKWYB5ZvnvHgmPo/HM3rs
Aey0VkWFEMnzmNvzaNq1VicpuBpNX4jmJQvodvNIVL83FJsM5kBzROA9msAsyIFQf6fildXlBWqC
7Xj2LRJKL2X+oYshciFpqwnSov8zUrkLzdJ6J9VfmegpvMVQW3qOZDvHEZucgj2KVTe0QnHwFW0I
BuLXkzH57jAFGPhRDA/OPTvaIOPESV05rkhXbkOIb6zfgOp2mfSQillR2DmbxzF9BJCAXkDgUKjs
NLuuSsMSlorDzIBBj20k53qoQgfO5O7g+rMc0Hue1JzLL5UbjGP6xhV8/vyUSnjtF8xiNwqy+Udl
Ekp9tL5JhGEiTMzaWVlPtqYuzGzPRxZsCi2WaLEOorIjNrg77vDqoJok9KREP5H1act9D+4XRy65
Z3ePhwZQsmCkMoOzzzFyMe5NSEKdey/S80998JcwVpxKURJe+xemqS8nfVR76JVXqJwFV+O55bP0
RfqyPM1/vg7trk6hsWb9eTjBdSao64nRANZZHFzTSYjNA93n3Ql9Wq0+2dVA2AejiR9mWjniMv5N
EXyRijrFgNoEFBdi5g25YIO20VbtlSPKosFBV3/Q3ZQxsFn14lshxrmO94+remYX0F/VF0uPJP2K
i8bgvrYrn5PHIXDggtqp7f4Tqoixganp2haW6U6I+wKhL1132FkGLjJfOHJ0CiczjIc4r9sAskNC
YcBhRyvPcZfxS3JbRJHBqqNtliURQOyyUfyUL8HwC0uVnhQ48dSdycGv4DtfLy4g74517nkYlnkN
u4JMyG/pUDIXr9Y+2sB0SK7EZutPV3p9hh5PO8dKa4LmAEjiXGAWfWU5dzNsONGJGNSFQ4mz2cT1
MhE+si+Vj8THWon/cHlqWzJZZN/rHuX2bKALTCaHFboKuaQ20GkhdjacodvecxA6yTbb01rxzgWn
czytGWI80O998Hw0n+x3ldtqJGWMLmlVaIs0rHL7DEyUgHydymeIYgkG2Kdg5Y1+Ur6PwRWiRaQh
+wxdyu+4Iin3PPBXD8neKvwzzeu/19diRzv9mW+ytgirP2Y23zo2/UaUriWWAfo8Fh9PNiSOa5UY
hlk/Ag8k4Ru5s+vhCMsoDqDCbQ9CDp0IHfxfkDjrLuHaY2p6wByv7wxfJmtfErmyDflEcucamL8E
PkwwxKsBthKGDRF1PCZtF26A+Hs2YDkloR66EuURHKIfFRmg9Gw25D4ubCdMRxfwSVTKwNAX1zA8
GNDdmZsGzB3YEEEkA0qLWBKBwLeULwAf9PasFFORW1fjUaQLR15VpP71eYYMuswzWGW0WHFIngHy
MpwbORMLnlofqX/ykUwjgtyIlnfX4RAxMno/P3B9wYjnKzeci23JPLf4ASE/oPvFROh+IeCff+xX
1l9x7vKieRebugEh44c3yb+D2gWGocynSlBG/74A5Yyj02VATJF0W3uOKK9U4MDQzi/LE9OtkIqj
BTweneaz8iAkUb/Ad/IiWPLtJlxKB/YKmLOX1xZM/UPnVt3mYMrWIS1WCClRBMuhW9ltP752ZF6W
KsDKw/xZn7H+G0FFuPfem58tzzq5up/Ji5NQAYxpXxrmgeGOiQEXqdMN2dktmaAwHSh/ntRNrEMQ
vMQE6LtebUDkC7UEgW6tm46bO82JxkDOoEnfYMT8ixfk3xzTX+fASEmb5bEO8MnG33V7hPpaNKcS
4vhF1E2gp0JxYZfDdJ41TBfSqU8Dinl+g92pSRR/xQqFLXS2jAJgeDOad5EYM9xb2oAQirtmWPtJ
SMpEgfjoifvdKTHCi4aZRgFxsdzx5cs6pKC0OD4R3emYceNc66K8lLzoyXdfwLL0jXYmQ0ho3yCc
tqryrj9sz7/0E22+Hf9IExOqVwB76TfGqxoIYmcfyZHvSQacVFfhSdTdYS7Tj6aPqh12OP2LD7mS
7To0x58x63PxBPkfMhaiv8EJ10k1ftLOpEarM2b+OYp0q4rdhtUMciFrETXGNJRgBVVIaVuIhPiF
36GklACood5dD3MWTZM7jtYQ420o7p703o8KBN1X4Ob3Sm5/claXb90876NyQQEBEcin6YW8dsJq
sP+Z0R+Lk6rxMDVOB3ewKWccIpTC8dUIbuA0cuWtR6JgifMiQkXzv62BZ/xxvwOUZOjLWU0Lq8yv
DMdtLLKAlxVet5i8adgx6q71mvhArnsXVGLVOFYG3wmr/1aHVcTGMobdWCmQNJqh8c+plEDom0nu
pb9soM2+XyD8s85Ejyy/kVnMHnrSLJ6zGog2kncec1I3BJxmgq6vuoVET3MmL5Z/PObEbzZvKQ/A
VQXCK/+xZWTkzkZyCyEPJ3R7OUu6FYHwaUEQm2Bgh666XDItjMk5MhBCUdxNW8CMUh8WWuFlXL09
wGKcpfThtiRpYbURaTMVDhzFRLKDXGOFDK9S3Sfp5TJrKU5Qn8rCt97BKCPSeY0EfHHe9VfBLtZX
XGibdoI3FCWPKK1GlGENJslQMifgCKSbGNxrOCGffHJfveP1Wgw98a+2vP5SXGhs6KOuvcCmkvrF
zj+VjRqwq7yn/6FDeARbxyZNmitwW3Mt6X4qdPi8rnlFR4YWxU1mJG6W2YRT10rOr0AAimmRLA2M
4gd7cBaynPdOiyXPyw7neEXblavXXDkAPK7HvalbF6WQMy/2f7skddqM1HGzn6YSP8mA7/Nj+ch8
sM6uUtCyJS1f0h3miRdAsVk1nYoX0ujwsOq4wBlE3BFuqUTPjd2gy19017/W9WZJSBsq9IotGtbd
6mbuwFBURk1YM/jk/geaJmnCKmw1gd7WayMl/embt9TwaDzpKF9fG0NM8OM0afTiAANMcNl5rbDE
BydJhHhRb9jzvxpOwsy/axc4+Pzp4F1D3slMS6t1vu54rKVgGLjmHuVRW1rKciRtuvfi9OIzSpDd
4talz5KhaXJTUYBFT7QpMZCIVaTiWCgbwOlRVcNs5yol+hBHJKoYQTdDx4AAl5P8JO2PdfxbnnCG
GqrepLVa940N8Ox560SiG5Opy02mrt4zmvQ69JJAbdaMU3QXMWxH9ubmgbm3G/sTdwHt6OvokfJN
5QU/uOPt2K8gPJyqAhOzWPY76umuuTGucXyL7ORyXsuyy/up17wYxaG/Y74iaqR5YqtV8pN1bFTY
zDiP5CQJF8QKcGUe5bTDPR64glxN18fMT0Xpi00VwNw+roJW6RDBbfGVl6Z7vThwAUrmFrSTtkKP
/q3iwH1rZjHQG0iU2XEXXDb6sqQfesFvfS557OckrEaZKZWz/G8XwUzkt6DX4Q9TSKusXDF3mw9P
x/ngd3K7KEFNVa5VEJGyaWEe7DjL89Q3kAM0ayxa4qiGWCxjDkXm4rr0bLx3ikzfFntfKcCnOl6p
Nz+qfPcTcE+Pz/oh9AnOByn3DDP264CT2vXF6TYnZTYAAr4eAD48MgU2s+n2z9KkLgnBlzzzHSVE
Z0Q00jbMFmb9KXCp5peo9y4vzEtsRBm+kioLgszU5R3ogf89RvibUEr9lPxb1Z7MVi/VbssdXOQM
BOtNW9MVFRnDbqBjJOg1+q0HXVCQvU1inCXrCeDjNfykMQVE5niz/swAVt3tEUqRBjrLnDo9pFJQ
zckJtoUL3fpzJaumrQegMB+Y3c3dz93YhD/0jmbMNs+E9uvqF/LHZO1v3v9CacGoNYJ54wFSzdk6
BL47Xr+x1NXGAt0QIOhTfWFdKJZdTRis00u/hGLeAVrNWWhdAn3yRsaWyW+6dAjpcXL9s1YVXN9B
P2JfUURCd4z2KMCoeqRLtXnWJCvNH9WASIsKsSgq1yVHfxB5kIgkmF3tCHsNNrD4Qaw4qz17w3nF
jcODcCIg5Pg9WPlN0zDf8QrnNQcNetJHg7NtXJ3rwoDeY+FNAQwNyANBAqVC3Sev4NFYl3n8NT7w
DrAlbMdkDsEEogwNS83Gp4BnVVDS1Vsg3LeeHh4f4aettsVkv4ieX0HyFZ35B3sYkrB2/yMdHZir
2DTzHEdquKorwr/v/SSZWPLikzB561/+BVew2yqwwxQRqMocAmmFs39BwD/D4l/0ktpmu0EossYf
tpjoQk7/E+Kbd47QfEhNG/DWddP6svoOQq2H3JCHhaC8RYkr3FflXvrYShNBiPIXQAfFCl/EGkUy
iKsq1fqf8yB8Uh+hqs5FOU0fMGK46fYLFJWUOdpVxf8xiKNjPwrHLfdRR9aYJVLVxvvQqLknVAob
qkJjac5nY7b1tDiIbLcOxgKyRGDIVGO5XkHr9sYJa8O0puC3+z6Nk0Zc+miSdNmh9ySzzElCbWc0
Qt5F9ZMaZrPeFrUlzOjYbjfxdRM/OfbsBiUh4qXoXA6J3VYEBzCrZj4bB05u1oz/c2hwSceB2vsX
ZksG4FaJKdnkBJWy1vqZ8D8EkOqkTSvz6WD7A3Oy3d4G1SFu2ZmjdguENJMzQyrv0QFmAp61mnyj
usPukvR05zy61XyhVRmW1Z6sjTTezXER2V9I2hATRwe6xW0SRN8bWPe/y00eC6zs2uB2KSJb5mCr
KYY9xRhxvMLyckHlpM6DEfMZYBC1ejiL9awj7HfWni2/tWNuGw5ERAuQs52gq7H+pgHQ+L+CoF84
Vp9aqt5TSm8KjdnoqLcTaUllwuGSXVQqtABTTzILU4VcMC/MqQ8gCeyF5YLBQmr2utXaeN2nJxKV
cf9xQbCF5m20cpmfLBZjlyZpw5tx+FgQXJ36Jh/XM6JQfCl1oNaKNqL6pLBjQHS/TtEe6ESISswt
8adzqTuqsNwAkrVw0hB7XXv98Ffy1lwME8zqS5Dalv2RPxCJFvMZo4ctOdZYg3gvhZLxax+aKQZm
CHj/X925pUxdP7Lglwsb1KdBVBAA7HfNELFGUhk86V1RpwuWRA8JNzr5Yd/PLVWVzlXsrX0GEoML
1RLoWPMlxA6LJl5BCjJBOSdpSjbZ71g5YBpzlb4RsXJVBbsye7BNLRRaAb2xcj25Gig9CQsJ2aqS
xnMnBFPUr2CEQ/ydUh64Uhgi/Rqaadbgyxj86Jho2ftQR148F0DLX9ipeVu4xzf8eE6tfOcoChjG
jM3xV3Y62l6HHlhuBRzRTOKZKio3PJ2lbt6xlsORAc8RJq6IFRcMEXaW+d1eyukZ8PzMoPtoXWtd
tHOYsGFRRTbrx8GDd6FNG+BiDSVWOx51KpL16owEEr+TW6PyeBLooextIfElwS+w+EN7EMI4IvL9
TiGOgN2oPgGe3G/R1xrz+Yfg4jzUwr5ww1ufwE7YOlgvhneTGSzdM2Y69rk/9iqmS9asP8EYYDgB
KhEWB0jwvwoB6NqNkhmhg5hLwoCTkJeLypEKP+DZJ27u6HYSwTcyUMbC9uh2wq+xFuqM6uCCymA7
eS1msh8sEzgFes6Fnjt7EKf/D3B7B5uyr0dIXFmy0QTO69jF24Q5gmPnz8rHnRCucSE3FpAESm9y
6Lr+sCzuz2goSoyqElKGj9OzbIz7WF/TxTkTT5veJ7LCSgmv6+CcMi9pCACmEeayCRxt0P7m4rSR
6MQwoec0+K8FONUQGIkayfRcpkWcdNT70xiM7BGHu92wznEGAEuPl6XiGwRwkdEdrK0iZoPlN/Qu
/0C/Pj5Gn6E7njo3CMfDZZjlcfqgOzXSPQSnpWp+ZOiOPzj1ypDjnwkq0ngi2+1cYcfc/9ocxnev
sl6FbmWtmL6gluAPP5l9S04+oe50xN5jDRTivy8Tjs1Gjq8bXOyULTbtRv5UIBvCnob3ENY5L3zQ
Mfe/hFNXgU5JgIKYn/nesou9JWwjqGkn5lP8SFKGIWd8e/1Y0OyAslSbI8G1rMfC69bvprhgWaGZ
kMkgad/J/1SKLNTuAfT+IVGBov4LCx/cJ9W5ViU/VW7ehzhvSH8eYctPYOimGi/oRgCwXych2ICE
yHa+z2dxue7OWiMwzLFBaIqVqtghtCUEFvA8HxyV0aQLH1DS/qQIhCHm3E5OiU2NcZcb4bgSO+Yq
/Kzv7fVQb0QFRfPwnF20C0LR8xqww3Brhhy2UPagvjRzHGyI9505B/8B/MAurEY5HNA97AlpZ8So
weSx2WHswgxiSSZRSzjfbAxyrrcVgzqCzp5PQScHa3F2b0yQAjhwVgo61bysgRnjs7wQy/GvPyf1
tr3VZUfTv3x32aqPUD/GL40jXtZBdj8a2hrfzCe3WIxckmMeL1kWB155V+RqC6dI0VP37M0t5uAb
kRqdmurvKGHk2SR0QGbb8L/GpsVhw8TjXilQbjC/3xpqiSQbMjZuz3/FNYFXDAdOTm6vDgpUs/2K
0rFbc+4v1Rkwomq7BgatwdZ3eedmpGPAMgN7Dlne4TdoFEm80tR9FtFGonQFRqFqO7lmKstxOJfx
g5T4zZ48hPPAmNl4+2sSy3mHYf6Ncz36ggkhHs/V8/1mMnn8n/4pK2lVMkEFpGq9D62Kl24HsMs/
0ld33El3HKKrjrNo+RnJ+fktR6r6bZke0y+D7EEiM/eiX+LOVYrXtJvqrTdPd8FnaAUXj/9q48wH
0NNvYX4es6zEvxb6Sn8i/r3dpdBGfXUBMoejsHv8nsytJmBB2S+XLAVyAj7jtBoCOxBkQ4dhtXXL
Yb+0995pc80YfwTADlnNGAa3z3nWlAwGiMbZstIHqvl6emJCEQsElkg6BnkA1fnks9h17CUkvswQ
yMMIphfqgdWwhW4v1tkGC20cvBK9b1UkgjNKxNx3qCgvkIG0hzPJSrwXDw+cOYWrTeIP9bPWzIZY
B/AgLAmz2lRcncEUJgiNKDwqxPRBKifpRapkDTSuellHtq41F649/yfjw2Lhz0YNK/T2KMelrToK
DOdc8/gymWnREV1e0omtLqupix6WBMI7CaxceAXPXBOuup3IibNRCSyoPLRApBsUlEJEpw5Xm5f2
6ICX8g2FHlFdHkGpwaoWjDcHqfDOwvYIG+AON+KXTxxKjS7s/A1GlBTo/71Q7K+xPef3uz46a7o+
5tI3AcMUapjX4zJbNS63H8k/jmob91mbFFDHkUxRWg7lk0Q3acm7+MaeAgmtXfJ5Q9miEqKjJhX/
0tE1eOH16HGjmsjB2h7RzRb9UoFLT8YgUttSJOTL498qey4bGQ6MfJvrV8XELRXnXRMCOi1PE60Y
AAYBMmyMROLsygnihTRjL8aLyaJrvy3+tJktw4T28FsnnLwC7rctf6aMSEXLYocIUHsBuYxcIGiO
tZjAYiTtdNT3z/vhfdTshTSuOC2zkUgWVluU78meQNnNadE00DchuIiMN0af9dAYLbEyuk3wH0uV
K0ZugNJJPyw1mZPBuq8fK5nRtqOsjnmeKIIeFfRxYQnW8/n0w1rX68O7O2Hz5O1EYmfBOsgLhqAJ
9S8yHfDuyzlCXnxKGHc4P3oCv1ONpHPJpZKh5GNdwMg0wHrwOf/Q1gnRSNwzv4ooozaUAw9tOoXR
J9rDEs30PZs/dc7xK26pSLmh//SXqk8FKhSZeoipwXEUqyWJ8WuuZn8PmqB5lduh+rW1i5mCasj0
3bB0dXJLxU2BMMRnE33QuCwy+ZKxyGY7u+OIjqtMNxgk/j8KTbz+ND73xDYVTn2iRv7wakTeUOof
9JkOE8xO5x0Jq5D75AffBC77lPZeUWUoWFDvXdTVGh9h/zpX2TN9DYfqGshuGnCFn8AGpeNfeJss
TRLC9D6yP7dRby4hkqZ+cWm4ZHfXP/MHXUopBhfbZpTfn3rHR+jCOD8uN0NyMDES1H/lDPazJ/07
greqWctA0ZIfTyE1CCWfl4ZkqXwGo7N96mlbjx5POq64cEALvJ21WMKK5sjdCk9zS4eUqX5Dmjmw
pu2jpxbsUyVkUHbkxafVsxbZHLi8g0FUGv6u0YEbfjKKOOwLP726FGEI8uvSNP9Kdp4spjQSNO+d
r7cwIHjktFdqd/ChWr7tGPgk6jacDPGvEEiaKsl8jNxKbvotN3RbeRYvGBsh+NavD3acJFWloIja
5vSarhXVxZhVNcF3oDQnwP5ABgrMW01h9JFyBvOxlK7tzZANYpVRAknAcDFx2u/I2PsOzFuWluIi
u27vS2uP8KLdLIeTlfO15aOkq15saPEFPpC4qlqUquwN++h15xMRytOMa9HMU35tLDGd05W+VL93
g+V5pjY92Qbq+Phg0nyQmmEy26/DA/a8DPzJLM8DqFDrSkTXfgrUlozwABR0SxK1O7DI+wfeMT+u
7rcw66T9z8ixESByxra/TUknUSuyjgJfHHDiBXsgxg+UkdDfHwY+Js8GDIo6IeoFardJf1iMT0XD
619ApB0zjoM2iymNGkKSMpbh7qNl01WhThnibReBuXPNqQJPw2Y5BqiqwRbGsAeMVBtZOlk0oYNO
16txh4iY7n2hZstoSOU4wvZnwlh+f07/KnQJfpiRIqHBVZTMSbHY8gDgYIvH+YRp+0xfDQ31I1CS
Np9Re4TokFfYOp41fAjiDsPuBh1ya8kH+k/F9ar5iIrHLM5vBnxF90K/WGaWDJP5BpkDh10AcN5W
C4cm4ovWrPV649fzOmyMQIZDuJ8ofrj+t8UU/b+JyAuBAdrpT1vaZwu11yPe2/b5KAVUzVnUhmD1
EJ1stZTvcDvF1pWX3FekGWpeb9MjMnYqEgUoMa5Sr2pUY15XAfRGPKSkhjr0KHFv/ql9d4UAp1Yh
0y+NF/qddJZOk1lcK2b8ldaVzmcs3HX1crvarldpmvEHWvA+IllccSfSWzuj4oBVYp8IerB+fwj5
+vD3HAzV3M2jHcSu4ptxQGR1aLgp6EqOB8lNebwFTK0UR7sideKOUIs3TVih0sCgQZL9y0ivW0Kv
JK3b7KzRsFy4JYWLH1rvjlWzw19P3RUtRyz27NdhVz9qW5s9s7fEr6xuaQV9Rt9wOejQC2WzitCd
XeCcufP1ndTEbOnZyJEsAvuINg86KgPlkT5AU7SZw64wf2rgvgxbzJE2X4nEIz6EoZsF3WDP1u45
VKmzu4vuHBm+/fxh8RHsSNCAA+c4fLMhGX12jvC2fwmTyB4fyEqsl53QVYHSHuMt7QWu2bqrR/U3
Szfp5xJpH6ZUaBeB+DJEuMEfS4jLeg+Ek1DSQi8maPUagervRbc9mHrSlWt/LDV0uXUvulP3N3Im
JVZw0z07Fn6aGlhXi28WYUqC8/hiMIyFdt0ilLvpEUXP41NoU9nSP4Mi98r3W+pNijP9DjoSSNvm
8O6qic6Z/76MfhlnncuN+HrBAQ2znqNIsrQZ4A2KxUJr84tyAN8gKosR/E5V8M7iayZ+0Q9T7/Hb
qU2w0g6PCNjUtAyAYeij6jXnE0XcqCzQW81+NCaNsz5jUfjTf/vCDFewgYsdqbVxkqP5VNNohd0D
BW9F7673LXUna/c/WQ7MXttlHK/FK+wkFpGwpCG/1B3LQ/thDFCEs/IQ73WxmcUSpZ9u/EgSyVsh
nHOX8fB0CKrUU0amuRGFt1yG5vPpJa+BZuCh2iYt22LpyrMVMGSZPUmaFol0YzUuwKJ41IrNSIqa
vdtzKGbwoUO51NWWegx08ehm2qDhBjfwxHhnoCIpVe6HbtCOgpuw4lrwEAvO720FRa13OzBF+6Ni
jgaT9aAXR9GJg5oDUFNaZ6jGcvMiAwpG0Z+rvFjEabOLyt/5u0m3u5waythZo2J7UCNFihTCbqat
YjpvDsKeS2+PyI2DzLBzRp04cGGNWWYMP8HygZtzGeLupnEwj5FyXWziqYEikKogi4ufLlWinA3R
TDljg/qEID9lcFATLvz+Km4fHZHVEpyKOLIfRaD7CSEQd7InCOjhTQjcrSWE3KqImCod/kBSsFsD
b8btplU5ngFePhPANtiMHLHuZ09WDHq2gX7HyY6sXCY04wsnk5zxJKeZjHJeUn9P5K3BYGLcQcoc
Kx0pNFOswYHiXxUiLsnvDRq+bTmreg/36N0zWpL7etQ/hnZc1aWvY1UZmCaJcUZIUpRPbViOxBYm
FXx+RCqqpesBeHsn3cMRDfBL7H+XskGVsodXFlZqEFZu0oo2awDshrprIf4Gn447IpP9Az16FKY2
ATh+qwc6cOC3j1hxblQ+dd60FVmXgBRM47XO65psm4+PIJFfD+rXMdoayXOPLJsSxPe5nA8wE1pJ
l/Ugx8XdrexahrHAlXQ6T0NdVI3UOOXq/xFQ/mnNqtg/eEsIjcOMdjrBYILM+ss5WXfnyAZGBQNW
vYLIXA224zlizm9xDtEp70jeIR/hhszUjpQiDVherbf6YWU7kcuKrGzszOvQartDV/JVA3tcTMzQ
XeBDovKpL4a/iosQMNausNFfWRmUdifz2oCs8K3bPqyuDzlbUOFxFBt2CHExUt81SMiJ6BRAM+Zq
MFTufiGHRTTbEifYbk5+8qZYhN3+1TEEpqVERl3/2/yIzsWDDeIc8ddROhjvYdg9vSQCEYk4Mfzx
4OWuXX7IeRPYc07nSw+Hibz7/gmuPqXtESRa2iLa33/U57aWaE/moq8mTul8PL/5e7RCn1tkuHv8
aIhAKEk9Fksf9vgMs7bT8/xUD303nq1hS6jx2S2zghyzn3DfSYrtMO8tM299OvhVZ1NHvK7N/Xuq
Gpzx/CiTC5wAaHt4Cq1wdo6TLqN7CcuHGEunf5zgPdAEit6Nj+8Y/2xodQu/Rrovoih4DJ2mNzz8
SHJKC1a+Ijo2R/6Jv3TagZW9cMWNZ8SFvQM8HBeq7Wrrn7A37etCyQ/ivtUfXJpkBjJpE5f6MtxC
tdQrG6cMePeGZdtxCCZWX6H3Pgs+X/6nLpKZQO2pWhfCcr0asYY7p3R/TZsESA+1pVL+o1+f+IHG
Fvexu1MHcAYXO2jnrKuhpyFmhrOkvujqKNnKITTsBW5voQmUugvkbbgUgfCLkh2JPbHzsJ/35p+I
wuMVLDhKeKQtFGO4NKUKg0qjqQOyFN1fNEpC8XoOG3bEv8PRfcX5YYzMYFp74AvDma+vUQUeZBFz
lAAJaFymxylrje+jr7Ijc+b/QyWXqUvPt46m5x669pd/bC5axxi+/1l5pg6dyzNCF3PVRdnkV/4x
HciIJqb1+JIakU1VcMZYZmkmUkUEyrRNMPlMo9PPaV+SZ4CtH99Y+tnkorgdXSAwu4iSKKgS+6Rv
97efVYeuyjj0DWkAaEAgbOXL6agxBb6k94jXnwyxFhfskkLp5lp/1YbEr8Y8a5vCEsBnuOltLUzh
y2i8bboraH/638jGXC2Wca4VrqGdTn3vE5BdTOCECDWA+lvi41kZWyNN8dVn83OEvgOjJ1J+GREA
QhAk9CTq/LyhqsLLUjlEZmNVkeudnWXd1ytqhLBFobytrD/HeugDAUUiKCToWUeA5wd/pEyhgbpv
r5NZtvjtwZ2QQQsmrhcAO2sx6ZXA2rWU1rnExLXueRvUGgrY8liY5UvMy9HlMFbK8oGwY/i+InxW
605idDhDzkPR83m/PJYWHcmKxBaNuZhnVP1k7oLhaDuRjmh9mtBr0gRu48qHCp7pJ3RRxj1SEv8z
CavWCW0ktggGGjNt4ixqVWOediPLOhd4kMn0DSH141Nw/w//WgG3E40zyxpxOFFP0HYDtCsq6KHO
UC7PO/5hVcoxc6xtpJNutZjvo2R7B4/hJNpV/T3GHHu8UfUIEuL/lrQyNOqNG6pDeJ3sp1kfrBdr
Lo2io/dL0mIO7QOrNbho9d8OJVVsC3p14u6q3UE96HGs7vObiJDvjTb/AJpn++iqONHk+AkhB/iA
9vyaHGqUBIJiS5G2N5uie10CMckIBZJBoQ+ogog7188MNozLDWd6bCHa5KArnXwJnaVWaMvk8Zka
hmzHZXQyaVZLUsbpj4rlwmqYRCTgBkTgNUD2NqG3i2caTOKlMlJ4mJIexk5TpDbKORSurDI8Yhpf
2TqKGm7ckchuPUhQ4RxYXKEHfaAI50JZ+Et2uZ41Jnqa/WtExvlIAH9C70gAMaQc25EOyDx5DSFo
Ny1L/OICeqmFXf8Tcf8XhWBO8D8mzIZdWjvR8mKtqEo2tf6z/2FFM88dXAZKO2D/RRyhv4jPnFED
fU5j1wjcu8RS4UzJm+VMQaQgmMzBO1Zov2+0Nd4nKKmxGBQ68P1N+xSDrRbvkwJxPd14A7DjwQib
8Yf8wX7rVfHnU8cuY8Zt0VWf7nOf+9UFE2mdG9pF3EyfcMH5jvEOznnk7MQHoxIBAxe8+UoVtFt/
vdx51N77HsPdH7vrKX47H9wAvUWFuAFSC8aUguJ5yMN41VrpPaGRDSPfmVwcg/XrNen97eEi5vRi
P5HIRn6WWwzIlfYmsBX+098oCFoRMBST9flw9BpVjcR1vds8BO2NQyMKPM/wAnHYX5q3GR425CZz
PEBMlOOy2TwB3UtUMtciTxpQkYstnu2b+9y0f+O7VlxeujZj4lGJ8TPz07sg7y8wnWWyp6iUKpwx
A9cWOLc86F3cc4vzkDI26ouhccNv0WKCLnlRlXXJ/YNHT6um2kKU29YMQqm0/frBuZl1KoESouXa
pIU6lU3vjSVJ2CUUBKwOvbk4v2nWFptdaEGsCXlFqbaPtuFYE5vnk69vOQbu0dzZUUVApmd8B3IG
rE6FCw214GLVoKsW8cfPzHXJyJmQh3cbikrGaIzRWENaNcw4fqoG1zGr91ktXke7jOWwi2eZ2ri4
jLFCrv+r+t337nC+absd15/B/MR8c1FHvwyuCM3CJj1w6ZQzBFWfuMJHb3KYio2aki7u6Ish8NMk
sZtnKOZflfTgurW5c6D8kzzBIg616zRRh5yzfNmxX3uLXi+u9AZj6aWoQf5S/pX2xcaC/nEO3Pxz
L30Q8dil6n9Uk6piSYEdb61a/P8P1IGlTzxvTgZyEddX1mp1JYmRK1njdNNGxgsCj/BRAH4cY94t
EdmmqUxldOeXZsd5cTUHSc9mRTD49wgjIc5qaSVpkttmvOZweqofD6/hoUQW0aE74+xSLLoCH5FW
7gXjMpNOtsAakahsCJMoU+jwMkt4x6bTcVC3PBmVv5ucltUXIbYtwcXo1dVBNMNxOfCRH6SJbe4K
+Uno00cB0CBVgb1Sl7ul8B+9ttPp9XY9bf/M/kIhPwlYztX4FsMYjftgKyzqfnniwrJcSDumSrPI
gZ29av8RV+h71gMED9hKBTH42AnogFcDz/1KUCQPWL8cyqR6nI6oZJpYdi939lEwgv+0iSpl9RE1
MqFj8hQEuiO49x8wakkDywDGgcj5841lSRXh0YDjjZRlNubuR5RqwlGDAdb+OFBqkJZNrB9tYeot
HH3XsmrW5KB54f+k3LappUeBIde/JPJCHmqJtt1Ok/sCx1IpQgpdNKwCGXH3+H+7MPPYIEGkYR0Z
ZmDmubfZuSvjL/slsg4fCeoP9V4UWtSMoR8GpP8EnlhXgHR5ale2dKu08brK/1pBoe665aNAJSbM
bC/r72B9sXfZ8Desjjgm4Orqc/SdEx6B+dN+QWd/fymOTh0eyRgXr0qLqiwlOuJbpiShMMgzAZPx
JSOPWCuUc1Y+/JNV0pB9qYesbQC1I0DvvjCi2+Q6n5fom98AhFHHTzVEkPBrUhkK7v0pUT/OQt/X
DpvnymJS8iUvhIVp6H1gYjHbLZ0TQu4bniAFQsGkcSVRlyT0wE3/I9tNh5t7rbQoBovTt7QFGXd8
I8Z49gdDbQ6oMPMP7mXpS0EI6GtimOTFBqKqpxkJxovCKBLEdZWDaIoTtC1Izx6T2Xv+pF7p7t7Y
ATaloeHwiJ2mt5n47D/xe6K94lkB+8YvgTLKU80dA/c7yLwf11TLBRJCtLhLw5w2uaE8oPfhWGPp
M5USG+fDUsGQSTVgFe7i/dlxMzGBLmSVBAC/TsfTibvE9VYrFf5OvUhLq9wpp1T5mRmKMdsv+gpP
yFVEFOQsi3u0aewCFX7nGfK4vBlgc+WMgJSs4G7WyIS8bip4EcxgzhngwPM0b0cHf0OVMxs3fxUL
MZE1JtcEMmGEizAHz+DaHyvSdCKsfOb8SUVp4sQlLCxtcCavzBmLdsUKJq8mveSmnFS1LVeZ3qSN
5nKgGq7+m9XjZBPIJNPz6Tjrv7+eoO+ugR1b8/KQ9Oxuo5fCLhj2qn81eqrskAJgIEtLQyrTed84
9TH4rHVUafn7SLKHe9utxxjGltysG7ZT3gLBCgo7fhgH+wmVtaG1hATHAUs7UXVj0DpgDTPgRJBJ
coQ9+FDR1pd9fdJfVrKF6dsqWMv+cnSnnf/138Ytc03Vwpx9S76DN87v1KTNdYm9/99Ip1Rb+/kI
TDTHu5hH9SteHl5CZLZpajgFK+Eaw7+YejSoHGcsiaWNUOWL0uVcgMfzqdalfOL64D58w7qIvD06
GzY580KCI9tqlHvfJnYLPcNnWeZ+HPDMJCp451WCIdwD1FZ0gbUnFa7unbmawEmwQpIHrCwmSyk3
tqmjc/S9FY1X141AeCxI4+OeQ6QHrRgyHGaTsWGrisw2AfiM+/rb/7mn0wYGClZfy/EYY8JWCegS
6h1MhXWoGY7l+6mlAJO5FJ2fKTqg3IXyawGX+FnOhmQ/deL6Nu+BGnGkiTq6VC7dQZvXnpfyiDAc
XlAo2irxWa8Ksic776T7PmkR/UemX0nUuZ3XXqW9A1IU8YMOnXlgcwGAWWkqcZsXHW6DlD/5qiBR
HJcFnUdNexP4JxXsJbkxojKwbWxb7e4IgwqWEVi9DFIN/GTQOeVSweiPOwYV5YRT5iEx0f+YyWVa
oJTqAVI5FgvkB0ZnNvdFmke7rJjEMRnA8t9y6s02i8ZIDT8dcWt6yhZTE7xtuQxQIKyYGdZYv47w
1jsU2Yh02rLBcOIcu2I1rUBtxPCmvGuaEMO+h4qL4wDM4SiqDSeiOtU2yfkt2d0ISqwJAn94Izoi
hdo4NekwPQLNGSgXkuLz1KoS4xbMAq0AFSYSSqW1f/zh7PN02iIVdYnjIupwEJQNMWEyN5fm4m9o
3KoqioTFNz8UAZU7QyYE+U4xq8JWXWnBscCYeSVieJfFOPnylYZDTtevv0QO6gyfZl/JoPQpxV/o
2Rj4HVST+t++YhSd/mEm63y6guPPl12rdcFxEtCkzCgYdrRo9duWLZ66YWGSYJIFRgSRvY7zHhPa
BvRWtqf2vErjt1REGnkDrf04lzIaMrKCJ4V33NNayYRSsarPEfRrA+0uF+D8HaBnbkM5TpTQ7tNp
l6vZ0wBcXnMWOvAFv5L0Jx4Z0G8KUSn9SLtQ/tcic/warlF9qI/4qI8cGWJE0BrVU40IHU6nLMmb
1SLXv6rM3EBYPrF9JCFrwBH4abuVjGy5PMX/OfWUKNUuMQv+1OxsTtlqrkQv7ugdTHjGcZIP15Rj
LERO404d9ybZ9eSnQXn150torclRvTj7PxQgRgWKiygcFwsg2GhtAMMiNfxNA4bAzz+Ehiq4wv9S
BaJZ4pbKwu20haDjFMkflfERMOK2QLtlxEomlA5h/+icEgmXgPsjxgrNX8LByKHO485WXQUT6zYU
VabDOf+Z7+WLFIhvoRwyUnRFgZiTf5Yw39uCkqt7qIfAGGJnNSpmRidJBLjMhPgbW521HlpTHFwq
+qe9rDCZmI1q5PDjbyPifK4uuDy8XIauSGAAhDnP1jj40JRnR7jdquGJCeV2AuGTg0c9re3lIwFb
2c1F7YbPUmoYS5e9KU1z71kgZ1K743N7kJ6r2GeWFR+BYzIL5kBjVYndyN4RYir2HJVrk4rg7vPG
yONWlEdCSo1vSsZRDPErhbNRqgYzD1Zw+hO4FzeGyVHFD+fcGA4B9M7+1T412uC6rhuw0EAabGY7
yvVsc0hG2BhsIqmzsNdMyJ03X2bW2povsvLxYZ/uF0JAJO23LpANTe1pWRGDxCQxZH/tpHRC7+R4
oDZ1e0Pjoww2xTMIYCI1Xu7KdvfmpgZbcQ13oYkbW7ld7WZH0MS1rLlxBvCFyHljhiNFrece9aTs
XzE7UTuq/0XrQLcWjaQxHVpN7/9L9RTplLn8itqdYkdHGVLXBLvl4ItanRd1OQCt6S47LUzwwoM0
BRXc/3nMvCuhICElXzkSTXztPTJWqfwUieUQgsQtHzDK7TRFAzgaLm89UcoKBfl0qtIo85PMjcVl
bZDc1Z2MfJHVkQO8dSfVVnCMIwGFBNsJXgONZ5R+3UWqp/mJO5c0b+x17EwM5dIhZ4OkOdYOLy9q
VtFw804QX2o6hY4q7N3aQ+JT+hQpbPeZ4mJ0Ozhbojuw+SmifAMaDrnAInD8mlyelC62hz6C/ciq
nVjfBaWgyVIIBGAHnYh0n6BEZ8e7ShRniKGlPsKvM/VIIx9xUHxn49czKnvbDdbeYoDPS/JO14/H
d4iC6j43SyKL3VGDCynKeQJY4D4E6cIdhYEA4biwJbmr19Dxk4p4Xzzu0FvGHdIzi8jqfZpF+32J
XS2gtnl67DIKagvi9ifyuSKsYXJdy0/rWg5GPadKHqiHcAVkP/C1JUXsqFr3dDG6ta9qogUNw07Y
fdWzVgn0wugTGp6eqNlUmoakSFFSwnXp9wdne+LSuUO9QOaOo681f4w4Gv+MH18fvfKeXGi2V7VI
g6zIviTuUcpf6vIn8fWfRSoFUVgoHBh5IThxntPRNCbE/pqE3VW5oR2wBW8+BxGzW6cGZ3RoXq6B
XRz7zz5yKeL1XmM96+13+x1eFNmfI7H13m1fZ84KvdQBBd9wbogMDvtW7hnPXcx89ysL9WmFtpsb
l9Xe5ZEy1qW7acPPqstZXrjsYMJiShuWfc3BRxcOUKkLTqOfxiqFhmt9mEK9Qe36Uu2euGqNPcOj
PDng7yHdWP0vviFtX+hnxfroY4UD/vhhdAeSS9s/p3TcYD1j+dDyOBntS+vTxJXbMY6sIDftHyBP
3AD0wFR+/FAbZKBFz4cQ+YortcaLDXSMw1jFmDNXr/VSnjZ4y0FU+tTj4q6W3qLCD0RHnq6teuyc
5aGdlC23DjMdoFyY95LofnCBRWPXC96W1J8t6vhmM7AiNf0jmB/K+pdW55yEhi4NH9Ao3cbU8jkS
gNaX5ALHETuM+tX55Fd7smjoMsl26fAkbCdDQnbVK7GM9zkNHx+rOy04g0aALZlmu7KiEF3e4yM9
VZ4UZTJo7Wx8Df3B0VaKrq+zHYxE9/fyBD0Q8szWiCq6n8B+ig3hbyy+XkoazZxuvQOrFWGVZOGf
4uVsMc2wSmG/vaQLOWa/aw7RBoWbUDGto+59ajruej9ZGE4NMzuaMYo7kz31394zWaN5GsVRyD7g
glJesKLnu9y+6V9b+7cnKCoEiVALkNm1F5bdgULFRr4kBzNjt+5y7IHf5nbl10c6jWgKlebO5CvO
siNWSzAAd1gVrg8d/XnsRciDA2kqJqDr5s1Lvw6it5Fl0+nKtxUqXRcjmghVv08hDMuobbq9pD4V
U0pY1TqX8OAG4ciLx369FzAD7DDQARzfqHt7y0MGy2SbCvgE4ZRugf1WHPTdUt7MUEjIQjU88myd
A4uVPqgTxRB2/NrHPCuz9ZCVDbAU4dDVbanceCmBAKPhz0ziHDHVk6V3KSuWWz4H1538+46owNU0
ISTKSldTsgMkkdcM61WG4ymzaWa/6cffiw4EJ5pi2SBZKZmt1SxcS1jqG4GThk2R8oCVMpwp6qIZ
ekPP+0TNvywcUS1TsmwZs+FXToADIM2ZPYPNyZAYp8I3sAfRJWXO+IUJpqm0wqF5eSYH+ewa3HB1
sMRU4VgH0qr8FHmd8iQ+OYL+VppNUZ00ZOAgWmtkWfILfHttOg9CCQr9w8YZJkM1BlItfKz1dmen
oebUdFxEGaKfNecSBuG8A+DHJPYr7HUk2TJFQoLrR1/uC6P2Z9aiI4PJn2kDqa+c1uqfv0kcJjG0
LpYstJki/0XPOxGt/fcPD6MU+kUZggFKqfQ9eT2Cn4UuXGFzs2GgZ93s9DnPeyN9Hxo4EEniv44z
6fnkU4R62cqwDiGxE3zAMS/kzGsnt6idDCqEGYvsWD3qWP1UbCnn5/NpabRPxZuyFTWoddOin6+T
170vRZLdqrfdUqPtZAOYv0T45becdJeisWYEValsQGEyfKC5ahzzk0ap4GImeNWZW8GBxosYHLoQ
sraAAkOWyDYsMqssWW+nA9Gn9MLJ5ILCYdWNZQUt691VQ9gXhYF7CwAHf2vYh3Hu6BFrgGXP0OdP
+vpWz4wgRTsBYl6PQbPxxDYVnyyFOu1o7nnzCOTKUcC5LxVQN6KsD/YDZxPxqLqPjhpXFrtjcxbi
M6Qxdkk34FPsEtKHStfZ6GrQ61uYpyjS2+jKW/6nUFFJmepoZIUkUCwV7hbxzb+BkTkOC10Vwwr7
T956lsvCJ3qtodap8KpGDxVJ409KiKn+APNYpxiEMVI0Sjb4EuitHEgIVMHAUokQ1HuPEfc7myU1
9ML3BvOvcwPx/7VsC20vhTfizP5vQSrhkXZwiIKUimwejjx31VB5J0ptvJ5wpKaBg9Ihlndvg9gs
3j2SYmvxicgLY/Huvxf2U1AXyoal4oLgFOUFjtFTlGMLGVHSEPRw5ZnleG7UvygqSLhENMxUuHNU
APT1EGF6dYCKXJm8ZZNiihichDGC8Of3e8/DQu4DFAx4/fojNcKPqVS5tvQnJc1/TD//Bb//8BGI
hjkD2sPcWSVlYEM+U84OS2J8ZUY98DopCSwhfrWn1uxX3pFj9LIikMRyKMePkwfFIQJllOpz5u8H
3OtXUos5aK/v+MplrK+iOpnNWqmdowU7eGzOnS5EhsO5EqKLz0Duaet5l9jZ9cdpKgQ2gFvw6JHj
QOIAXA5E7GH4K6imxvAxhBbl8TmGz3pxJenx+PjKLFQD0tExPEYPscnv8/WNXKilBemw9f6P5w+H
PjOt6+6Nrj3WVeQhAfMSv0KOgOhCrDzA08DH5l+BzlBlUVstOJoTqnS6e13aXTMd3jm+DlkZ8kpc
2bO0MZ0g4krkKOOtapeRdrba2KJ+RxeHfxJEOmDaea1jYqWMEK8DxHtdMltqRx+m5ZAY+I7DJvgA
H1/FAphrigfa6xL6zNX3GmBBE9CqJwjg+HujSmSFU06kUDYn7oA8ekn0D3DxhfzpreIhalmkceP5
2nhP6eqJDv9lnke91rc5sMqUEnv0nEKp8XDkUsE5UVatmecq2jBH79tiTPsQnpXDLv1u4Z1uZryr
qLS8HUd5aYcAm8g5yChk59b11CYgmjBVyir7RULT7GX0PqR2Ncf7Vx29ivlFzWHy+eqv7E9UyXYf
m5pKoLOB8a3ACX6IZAM/xc7H9NfBk1Jh2NP56/3LYvthZHJ/tUEQhIMRo+6kdDpZaUvZawmF1GL0
qXNv7df+JXlGOcVEM0Cr+RliN4X0IKi1IEiRUNuhSNow2o8br77ErO0X3tXhpNjE2GNHkCYHJqCB
e9vxJCNJQ2ACu/Ieg/JO2j+YtMpf5XDmykm2jJAHCRBbfDCboEnACa7YPC3+W55StIQCTM9WjOz8
F+vz2/uAeJrG1R4I89IGVqdKfc3oTobttLNZvr6IFqkQUhd9SlpRtFH5rIUeQFtW0SqSz2D4BbTf
IVukv/OPPfuCNhqgcvtcfO0Ci7UbgjgklO1/KBKZRmU3qL4NR5RsKLDJLhbLcY6qApoutK7hRYU/
v+16H+wGLX0xNiVGLNlxAqidBMcehRmBiGUsMNjaLbeFf4o51GRw7cuTvTgHy8EBK26OqsDAJrMk
tJELJj0hLS5ERj57plzvpGrlB9bzertD1PN0Bg1hi2s5Pw0bJ4QILQDZ7LaHaR4M4tqvsSzWZQq/
SzKwZjmV53+8dZUE3+OsLG8iZMoMabSfNjp+28VbYyz+b1H7F+AsouSNeGJExrRi0JcbSHr4hl1L
OGBsuRmPiF8dvUe4i3XmkyslCO1Y2mcLxGGPo/4ki501Csi/NlXNdBoiTK5GR/4HQM5ZxtEDdufN
72dCeZFLTo5D+xJWOpMYuRMfs8EAlwQXbD/9qB78vkdYo3A9PQbk704uqZMIKWjlWAnVQhtyT8dY
de4B/o006/OYDdOiNEW65FCf8oaE5OEGmuugNwubfZvy+52VYKTujjHUqkoDFvNXUCEEOcxvIqys
o1gExZ+850zqohJDEUv+IQvSlvTDBoHWyOYlC2Jrw/iH/RIAjEK0YbnNZySFpQ+PZ3OLTG/lVIZU
/iUxJp7x65/x6gx+6L6S2R0JVg0H508cZ/7obq8tK2IxlVObv2b0n98CzxQAfReXbyIALGpOR66U
TprrxLxun8ZJHxzYxDRCzRu3uhLTwG0PtXVCYM/Y9RjQ5otQyteI0HH7cogWNNZ3P6YpNFF7lj1l
6WW47Q1WM/TXRbANnkAY/b6rIJp3Tg3axvJB+vQTJgDRGQxtpxZTkqHWgoqc+Q3feZUqvvoBFp8u
Nkn+jCOUXpK121ZhtB8fy1UjT1qN6gtA/fi4Vc8N3AyDKg9VSjOJ8QVfmHsvxXKQcX78HR0CHI2W
u44z/PPAv3oaePZ5U12CkQEG+4/5nBybPRth2A9DnlSPVJ29KQs6r44PoMFK6EKNZkpXtAUvvVZ5
9fVifkElTqXjC6nCLiGW/+/0qYdv1BKgt1mBnn7PJvsyNuBrSfm/8e2dV0AfsUnXFiyQMhoLwRtY
pXPQdRkCBE+tlGyzg9QaFLO89sKWX++AwIx4pW7E5DxUTYGbsC8UIr7BItyUaw/XkFnUkgDKZQDZ
Rpp1+uu0zRfXay5JjG/DeUpAqIvLqw3MNOCAalOZ80dwcvxC+3yRkM7jw/Md04kncsno81VNmzsY
wIl2cDcpgokaopi3I5kHIH+3nGPq6iEomIHBVgNZm5GZQwEebXb2PSM6WCbuTMHfn1RRrtFuo52a
d44VTJFTJsjSE3VS2nYHkR2Zz07Gz3nHfOihGbNsnC55HgPgi/w+YMBFaNxT3+NPO6Y7yYVDnBV0
PxaVRLC4cD0UGLwpKMkFrWVOh8omqhUUnAdpFq2RtNfWif+9tuBumIQx4Oj8D5Y0WAPl8uQJmoru
tG2st4jm0zuF0K1v8nj+2l0R3dXl2jsmOAwD2LsglJYcbaM6e6mk1hpoHQsYOw1Hk8WVtmnqjcki
7MzYnlBahxZyKCkZmmhD02TdZTfzEIE35e75ItgrtR7cXIS+WRBOzbYqlbSzroV1+ZYl/Sf/WiW6
Czqr0s+kz+LtQD2ViKBhHttfOy6YRXms9Sc7S/AUouggnyBYHBaLLJ3mH4jRcLga4fqD2Go5iJ2B
5cxbHQW+IGHx4UAa29kYc0JKT1pKN0n0au6IbU6v3s0iHEiKC3U2DYkQEAd9qC66OHXMYAfBm6q3
jKSM4+GrBoKBuLFfQ0C5enlE0V1g5GXXnTuPDyS2rYL3vVfNTxOiKVQSxRiu/keK0BBszR26w7zQ
mMsYgO1c6TfMMFZiiGWX/p66PE7wlj0vHY1ub9mPrL51rPCrYB2VtEX7Jr6dJbgktR9hf7xiHtLg
M+tKIPYoVBOFwiipm93rOg7mHavRhY7AAvZrGuPHI2ocJp/WkGMsxi7Lw41Mr6l0Qo8YPAiel+6t
WhDz50tYjZDz9GqaeuZQvpVMnageXAr4KeVjeGb+yXBK7/EAL84+tqGWHPafdMwRPHAU1WJZu4e2
vhEb4heyFwK9w4iO1U9fhmmblpuYlfrNHyIq+wRxQQPSoqUZSYIhlP7pAAiOGH99ICHNejpCL0bC
ItweOlwn8G9BuF+Hx2MPSSK/ClffIxioi3qYPWEnluLjWd9Tm7zIiY1ODueJPOk2PYNmA64tA5nI
Q/AYZ2C5bmCiBGIXkVRVTqkV1HXwpcXqU9xIsGDkf31WR6NYB54dZLIFSVL7Y1KiaqF/WJaetXrA
jZPAWbJwcTEnapW5OdP6kRaABw4p7ll22LbhGCOg2o7zyIu07EbVlaewvTi4LmpqLZ5qIgtAn+GY
pv0T+wibD6/8r6cNGNQsIqlL1aHOZnpHdISVJI67lP3fFNiAGqlsi+fxPNq+BV4QFk7w55LTlkOR
8KNZ+3XMJ9rsh3LE031Ab4sNnwn9cQuyr2A89A9wzb4uQXr6ii13YGr8QoCSalApduJ2IOZGmQaH
lFVo7b2kt32hai7XJhvJrDxexr5NCvMu9+efw7ezdSlg5SDq4u6fOjGGrCwu+V+wpaF+ENhlTTxj
pH2LoforZAO0pNvd2uLuh3NQn4zBv0RsB2qnaL2tIc+tO5PR0P2nDdDPS27TexJuG4KY+RmxsZzy
WkMaLq1efcPuxg8C1MaxR1ckNVJnIdgE+34pWpRr1tF3blKLxhhnwhubS8nayKLaaXQ68KBotE48
MHsdPWwkiGsUR+tg37QFLuTrqOzxyzDpdBhBJMqHEpI+0oXhhnH3JAYOhX9EWdA3zfeb+GlSWpPc
AhT460BW17O8iO4s9sJ0v0GdEg9vNDkBHOL9k8rQ2NMcF+31KFW2ByiGmV74KsTrccLl8xwJETTt
n8pRAw5cNd8B1t7wnPYWa013vBQGak8qPcm0FmN30Zqs/PNYFa+Da4RIFyhyI5YGH8eHMfkiYu3O
UIVuCBGMDdpWAcBaKBD2c/MRLY9y3etQjeJJo1wbe6NKNtmuwrfN72K9z5o9AkgSL2n3stk4NXiz
I1uMIjw8riYczcs7WnFpo98qvOK7R1N74pDXo+J1TexYQWFEzemRIu+Ve+ITOuXkQPiawaA9htQ2
CCvQrxb5JukRVTIf5AY/tXT2XtyapYHSq1tgv9mpN+A5BNAO6HJdvjPBZv09w8izxMIxjeVXttCX
T1FEQCsHQ1Re7jXFHJb/fbstg7YvSVYklWZutRtSDySpY4q+cPO9N1w1UJGqvBFVxA1G2xdog9/r
LijI7j0tvNJ2mJe5lx/UrW8nFrsG5g4r4h/qxNwTle5DpWWWHyKO1RWji9qjlYbAxp8rbsA0A20e
5NjXLYhDy/cnGUL4JMuZfor7DoZlR/dzletrfc8IcKkq+dtiVNnEF/+4o5VkctThG0QQK6NRIwxl
Sezxt4kx00gi2YB9PDTU3Kpaz7ToK17f0+L3xVufyxlZSP2jCXo1Bn9i15yskxTTWQHyievc0mrI
9EWysDxpJXlDCOX+JPM2UfKo+r4NrL69OLfx8z9fcVXKcCUp9FCc/Y7kRzuGenNzMgK7+R5E25M1
tVGqQxdNiN+t08UL6DTmblqaHIn31ZOWA/7WuAmxrgkktSFzzz4rMU733XZc3GaxvRVfeykN8JTg
yP+WlU6DSSHfkC0nz2uzCMxguH6eSs6Yj+DDEnReF21zCCz0I/sHzNqfVER6mc9ZRbW8eP3FLvRM
RwS3675l2oj5V24kMsjHGg6B7v6wfGvnmNZGJdRCQa5fz76ez7MxtyhcFF+KtF8RZIQaq92rbpr/
XSMZHCHnu7LTautCUuEEsGKhxeVfWxU4mU1yuPrMFbRAfabB5ty2MKjNuEKrraYtQvcTqiH2EiWn
KXj+eE9gohfT2Xvxd2Bwy/YKDj7nYcYEFdFonb1aGplv8ow9UokAlj0PoC9gsSQ/uQ8anC3YWykq
JXSPEmnsZ3CpoRrxxCOdGSQqIL6/zYsgWlEtMs5ertc+50Y2cACjJ3mtS7vFLhXOA2crP41q0w/j
wiRVnDG2R9trnsKyp2tNpQOgE81b+LnTGNAEdUsPMfsesMBBvlgXQf4n06Kls3bapAfmpYPWs/+6
Ux4pKv5xre/DovRRb/ik0TJsRR1ac6GzW68eJTGioHEMB22GBdQOOJS7mlXlZGTgOKHvs+fRLdf6
nk1Fi+iBp+dtUSp4BXqW2TIbOZ4az3w1sQwjVimLRX3GMstLvL7QUChfSFSAGeVe6z3ukWvjy3/G
Np/v0j2brvRl/1tef1AVUwgf2apHJjSy5nFATJOdk2xcHMUtWX/pojpC07r+jgcSaZ2gM38NMH8f
YP5xjdjS4RMIwOgbtc3roH1ISOtQ1xxg8+vtNA0FBUcmCEDWmAg/TTcSxijFxdmW8cP84fT+dAvG
uInoKAORAi5Hxy8eD8+1DVB/dXDqtYSDnx8Ar1shoxuqoH5Tpq/EMXeSw0EdEvyMR1HCe1VFtG2M
hp/fveu10fJbHd14EPgh6UcXdqUR+/TDKyIHicgy949tuSqtKtnO/9ltUbIDuVlqy0gJqng5CWw8
FIRFJSZQa8znsUUwFMRwiy0NeoLMNtkA5ImQm/4Qacuow1KENnrJ1V48uLjYR+tNfkdgwCwXGSRc
tl2KD5hkQK/nHD7U50eUjK0jyL9p01fn5Uz9jj+MnFsYxNAroGavd7i908kn8hTa3pYj/AWymY7P
Y0vIxAdpeKYuh0nhKbHzOkmSL6e9puNPB4tqwbtVewPdWwN2w2vkpGppN82TY44HQm02417RD93x
ooN92dcNr2d21+k9dPnRBHYNYZlfTaam8wLAUFeqvX5x/wLHnW5s6m1Kf5qtI1+BlLCD2ToWZduY
wrmzkFU26MHcSNAZMiUKxZKPKZPt80RNsddm8psEcWrK8RQqIi9X8ELEMwfS4y2iE+zWAKf8tDs2
sgUOIs0IFm8O8nab2fJmTHjXYQnySB4BpVGgbFywzcwAfXb9VVKKbyHzdrg1xFmNpgE42mM1J4nr
I5QjZ1x3SqD1BuU+BPfx0S0HxFWc8H7+eyLWokHBb6Rb97EAN1r6aelBZmaik9bd/4/OCFCtJU/V
x0+lEM4AJN2m3r4MFmfw9ehKkALNgu3FBG6xi3oxXCCko73TB/o/Ka8BrBaM863sU9MYEMTeZ9V9
U4B04/msmc9n1p2rz9jf0EvX9VS3eS9Q4r/hx+KBj6BKsF9xpy3UK+qR1waXSX4cs1j7wnXurXQ4
ZMmcxU7ndHLrEMEziQ1xoq/5Ngp5uxd6LKYJuqKIRBd857mC+hljeXEJxnlI6LVbg6TM4GhEiEIA
VxTPpYTCGZPb/UEdHY9YB5MGfUInMhI+i3uwld6Eub2uubSe1lbt0sB3sC5s+C217n0ipIJTfsmn
AYCD2FKIUCTeRG/BVfZmqU0Mgwjiiddyj8IKzu58FA8PzxHM1rZFvSywe5CjMl4sGliEc5kRfoQT
mT11Yaal//i0Kepab0wa5XPHJcrg879rKHyZiwTbkHDMO+ZKUMaX2nSMw6VQtJAG8sdh8TcYAgC3
6XcTpIkQDJdr2cl3+7vYXCO0ULQRtPc2gwaFqrKEXKv/NHT6egPM/nDmcxzJVnBwx5/zESb+St3M
IL/viWZliABqoe6pszxKIjY4q9yK2Wwb2kQpAKlxw8iA7BIjzTWMbdBdKkpURwgW0vA4lT2RHCmz
3OtR9CaiWzfLYF5/uoc+MQjToopq4MRZo3cr1x3r23bzsG+3rpvQFVSFNDRDQqd53Vx5NZ5ATII/
gFmiuoDpz5+/rn8NmpCkO5wQK5HE1j3n5DvAmMVNkZFitGugeXR+Y+fM/j+VLj6lKG7SKE2f/unm
jn0buDFkOpeqztgd2uE/w+Jp28O1PK3spNPwzd25C129o0cAImuFiJ0Y6hZBVHUrylG0rpGEGiW2
4Yc501E9H6gwIR4gNPtrKfsR4QYHQbHkan4xG5o9CkjKwScXRkp1vY9lP74UU0Pm97h3oI0A4HY5
Oe8j2m3PhoqnQoGUufDHnLIfBjEN6uHY9KPFSYtrXX7PGoo1ag0sf2UFTNrBewrq3Ubx2oriMPWb
LQ2QoeuG/cwEbRgNkEW8ffPJqZELtIWLTQYOLEEFIftoLih5jMQKdLgdadJbxOsy5RoIJACWH1A8
2lBH/lfni8Jmi4x5kf79CBWrq1gRnQDdaUZ0M6ZVA657AsrpxnRljSALngmprQEbpFHql9ni+6DY
T7UQrxcmn2LSNUq3e9ZQjR02Jk6qiRJjKmmgHLMl/NPkbPMYpFvf2lD2j6AXNjl/we6HCUA3T0xX
oFyXqNN3AcIMjBXO4IIEfhHu6pxcbcD6vr9/jGGQw8ldsLGW9tz99/RxIak3svXZgx4JGz32ADyK
BN5GOxUHvTCrn4BB7QC12Kw1U+Rj+Si7E7sArn9Pgam1nLlusRigd97MErlC2YakKX4haCKqGGKI
Yeie+FKx9aKI2Kv8/l4NQtSWhq9tnPslRTTP+HDXjLEnspuV3+ErYH9A9BYIuMUx1jKh7m9yOC3u
UvBaHh+jwqDmh7Z4LnmLtBd2tqExWyJ6jXJXzpWyvmyU9CoV4FUoD3OpIPIh717LU9PmYDa09orJ
KzGkt4v9elPo8X0I3rkAHo4CTUlHdEhiHc+I1mTseM5TY6M9O1WKOekw0Q0JJmrCvw1cew14jC8v
J6qutelnH/6DhWOJMQ9EVjYjcRABCVV2+ZT99Iptw/vK0l1/smzfXqESamRXZsE+DyTx9/eqKLq/
zTz9qd8874fi2EOToU6AWb+V85pfiRwh9+SnmEaxe0i1fsPWIVWSGfqxtp6VR43CAe+baD5lAaum
7vyKO9CIz55KsPJVNs9FZyGgSqFMwBX6ohGNQBH9lOmFSrcj+n9rsoTLHL+qI9FdzCYDarHJCUzl
hU31wP2sOkj0LkR6m9zLWj/pHbp+pxwn/tMM7KORWE5wIh2KYJ9Wh1mQH+SMNtIBSfu0adkK5eWw
73FyF0mFmL5GHIMtYw/l8hiNx31i6o0PvV/SaR3UqX14PfzCjrSxX7Y137CGy5veBRWkMcsAnvIo
HVLygcSMYJN9uSup6k3BixM8ZHYlNvVh8A2SNtccgMNeqdQTrQOQNrNPObVl3J1fZ4YtnO/ZtEYy
3joRtlgIv5kGV7c9iijX6YAdDJCeBOx9WgtL1bIbBK/KUpShqg4Ut0Du8HMGUPo74Osm1KWCleDo
ADcPGMC6oBYrMxjNBsEDNzaNBPxVXIbrn4pJMaRwQOEWA/fbR8EJjXwuUt99hDiCZUW+yTlGY1a/
+LKGKbqhNHpUznAwvWOpkQajdw4ErE8pSXzjTDcQ6xCwWct4m+RgodKSdpCZVgX4R0cITp4xIsC3
A2Gs+BJuJ3NOJc92T4I2V792eYjUcOEcKmsgCkcKJGBLV6SIO6hrJyExUqxhRhbZDYJNu7DP0v+K
DdkV9z76slho+ZvF1lQjYoEJ2pWFoWp3kA62Xg6wDSG5WE89cMHPWVm73EMF4+dVvUR1JkSr40o5
W0JkCRxkOzNMEWqRV+/rxJZ7bOXiGE8EnWbO1Gc5gu8h2rU7F2+W+FODqLAjou8haFOyRjhclMiU
NtR8YVBkKv4FtDDE7d9sCvyCN/FAKvFszHaTdC+Oz31M/W4C01WxTegqt2lL7JnTa98CQNY9lhy1
8PZdT77AGMzbEvyERD4BX0Hxcq2gIzXQ/WMtmiy8fTOrvqxUrFvZikV2OagS9g3Ngr56675blMEU
8u1RZxpfQx00lr6hzkTnkPFzkAt4csjQqMm5OmaH+MYAR3y37dZSQKxqKgZ/ryV2BJG++HWuWpIJ
8d9wHwfr6fwLNRUACTDNBYWuWzLwWHCmebude/vBhoAUBFBXQ75o9A6AFnS6pd9YbG7IFwt9CinA
12g2ghiKAFbkVY78ylplpIut+3zVQjHlmVDi286AKjwP22tRDjd7nstzgXw+FfohxlWb99MTRv2V
eEQmrCIage7dL+DzkpvXHfmN9T7DrBwiL/4yguFQEBiA40mZwLp/hEQcoTtX4LxmX0+ahqP0OtN1
I8DQ3UTLp9obtWbf4XuCqHP4PBhtqOFNqjeK02/6tlf88jA0NBssWr4KGfqwTsJyNC8Qu0N54iwx
xzFvTnfQJivr1mq4VrTaYKe2BW80RtofRQOngqREGaQgO66S89uibeKtYGNdjh+6q0cJX/qtpHIO
hesaChvma/Y3BvHZnKI6ja0R6jSW6mVIc6hZXs6CRP2vfdx8xSQGrtgYBa2zMJsOIUsV/IJinAej
yGVN4BXnVj4h/N4SG2sr7bzTvssY8sIdqxFilveY5SMX7zHY3ya/tK11y2X0Mqp6NZksA1HXrlnk
Z6G76nSEJrdj0Dp/7PmSAPvNAzCG1T/U/tFBe/Ewg0MYy3Hszdpqk2yNAc6qDwWtHWuF+jhdWEsN
WQoSndCQxvlkyqgD3MyZS6U4PMr8jXofEAEFFFCK3YpodjFamKueLxlaWOBJu9UsZSTOsegOlR8v
ZGJP7eaG+SUddMDXAUQl/vCtNs+Rew9j9m4d3aZEqGyy0yl8fC4GYbwep4ZcAUJb5fSOqTyY76nY
z16B/dlY7AuDd9mtOQcIaqA/HPhXJF2c+QHxCWq/7TZZz1mADxoB9gO91wwq/k6CkuCX+nIlO7oB
2eRuFRjAkkJZBkfp12PXAPklmF9M/lSQ7Er55CjKrGd1LQ1Em/Z+9x9K9vi0QpFNjs/VAtbBsG+a
+cqt6pbsgxCWW/FO79ZMrsTKES5inBnG5IW0S0TJ62GXIifkfQ4MUu3Ks/KVtQvMivBA7NDN9DFD
JZ9q0QgOXqTu8Zoo3d2R48IPF/0s9Lbh0U8f5CQiVXhQE9+M7RAtsCf4xZgfzwFbraxH2TqeuP+Z
J46987n/kHexgEH1+H3Pqb1elPSQM4OiBAsVuDycJTpsymjXQcO+GTUarkvPRv8yeyLjZtclwOgU
SINxYQr7Iomz5qXR6N2kJH1Q2+7fIK7N4kQpLVu8ZaMpTiWntoK3QzDDKLkZTdaoQifV5dpN8XYE
ZpQ+gCwgmfnkpLvNQRUcObV/8F23ifzoQbnD9jvXbIdRG4vUy5Lr8EQCMqqDuwzdV3WdT6BqCJmd
PjFJeIO5XIwo8lAhRwveJhmNCjGzBFA0HsYvWGaHEpKmyZvacYpFsN3Lqb0ZzMd/IDTK9j8p8W4C
iudbZJMudcdAYgvV6gdVh6LGN3POUTNY3u6Xl1YSuiHRtHjoYF/mPjQbHDV3JJUYLfYcST9Wda7o
kJx5nJDqhyXBrLPJEnOcX3nm+ffSAJLl35yJtWDnCph8M3LM1p3L84wecLD1uyDpr8pw+OrMZnFL
97QYQrWuPfl9y45v8v9z+EZJJNSWcj0h6cyS+cdAbYAjef7DXM36eRrKXB72ph1Fx2VGEWOcfcbT
w5BPv8E65ycHUB+NyRRr5k5T/RHml5SLGDDta2u33nP7vuX7MFx6wfaT39WLiaC0/CGTBmJvp707
WC96Lb9yNYqRMwD0Pk4VPqInu0W+JKHE7a53Sq8oawMWIhJ2zuX/WDQMAR7/KgR+SBb3wU6g7zoz
oWBYCt71n9lyJ4Qf09dIJZ8aztfUlyA0LLWzDhfX3NEHBIB13P3RJdwU4OsySgxxb64BtS14NwXc
uCG+El98T8jL6cgU8akLXnuMm1L/QwD52mSsH/lcY9tcYGJa+EhArSLYWmZUy4t3qhWQ2rPeBygl
LJH7hki03JylUvcCpkWZii/YYEMqxI34Dp0ki+iHJ+DAyL+jeuaJc88nR4JbBLVX//PdduniAKZn
8vJrO7ltfXmD1zxrWGIreMlbhKUSQfCd+G7b6qBprGB2rmtkklC0hxoqDWvphneB2Yisar4b4lsp
O69Tt3IcEPBKLu71xMzhASswifsplTkffkZ8fGtkc3CNDuO/hMtjwJ4D72d4sW52vwpT7KcE3OXu
egxBJyPWMacbG1GaPakL6FROgXti7q2g3kyzCBraE9JRNKRfMCF6hVr3rhKg0k6VWSJgwV5WNgfN
+zvxFk4eRV3Li4lDaX/9iuJ7MXg+adtbq6iEvgYYVnZPUu2j1tPvu27HW6b3fVhSJ0Ue2Q7gEIsp
zJ9dR9EEKojpga2ybQKXGyfrc4DVlYxE11ntUk0LxLABJOrV0n5eFV3BLbr1St0wREq5AweusxQp
QPWXlQ6vwoVMqTLDDzVGebTVpJZdTnrbsozyBXi+zOxJX6mih4ffZw3kXvY4jRmVTtM4UGhr+UD7
jLDUZYXWTpNNgyQPtfeT5KFVY1btSd1Fk2S98xMYhvl0/joll9OnQepV/QbbM+/2Bl224nPgG5mc
ZcxiWA1P5UOkbaoN/PjeTEgpbBxtmkpKpCDeNqzGh2nzCDIa1va4DjcDCJrkOQ+jhNFD3iENEY7j
szWOhHUcZJRVw9clXNNyvB7Rws6KVwNPmBjQK7iaBjw0yonBgRW8Ak8QuzJr1xeTsodvW11ubtji
3LJtlMii7+P14SKxQDM35pnamlZY0nd2JOBAiTK/W9PJ3QQYmMQ46BeG3ZgkR+T8qB+btpvi2hOR
xNrv1h9NzG6ztUrIAb0UQZeDMEPaLNZn0hPRq6efQW/ghQKoLzglk7SFWocL8WHod9YxalpHoS8B
Fr9wntgv7k/8SHAUh+DCLjaXo5cuIfayIKk9kFZtHoYfa/+Towyef1tWpjzp+qkAtm7XnsHU2kwc
gU8qxJVx0DFBW8rIK6+6/oTAoyuhVEDbDa3/J/hMhwew1Ccl3xUOW+QB0xKBzJEhwgIGH0vgp6s5
92Zq25F06gqHDGgMQLliHt9YlM8DmXiTJVDsLNyyxy4Hr3m5JNW2+eo7Q+WrV9tFlTOfNnuOT8gs
HDt/1rtEKr4Y33UTxpCcfoiV+UaUFaexSnrPpgEsHy185fyrFtthImV3QSAHhAucqYY1uvTFszyr
od7wDsdMON317qkvqGv3X94tqj4wbyZtaBZK73B7d0Ca4RWrC8kNEJqTsBS/ebTdwHincJ7JutDB
7oopN6Lw8pQjqHlFTbIc8EhBHelmAIsI48TnEvw9NzOxPzgE6ALb/uhnngTRT5MV7dhS+cA19p96
15TS2cCPHaePQpBUiV65eqzD910sLgibazm2+lkaxQAyiFPSu0DAXQ074MJo4771PxJgAI+EaqkT
vbT8fMBcBDJlvsHncv+2SNTA80k8yThX86zeRPUEuXMugiYXnLdXUiRqy9qssD/v+tVzRA3QijjH
i7vRe8bevFSOKxK27oLaRH/Xm+A2h+Wycv50tgN9lvr3qB6fJTWkVO55Nlfg/j82OLf0vem1S3Ms
QtUk6vHGQswYVpmfafYviXepwyZMUvqwRkf0RMWMwR/ZUVhYS9AIJ9C3Q2/lXDPMDRdWFAI/vg3H
AOfWksv5mvGjMij7V1lVYdXgMvBM1op7j+SQzlldwops+xnmT9qRMw4Fj3nsvjw8AqhaDOVXde6C
0JZ14e3dow8N0MySDdxX9lX6vUziHTy2iT2R2SdM4eJ16168BSrbbyFZnVqieun/BpZfLgz6e2W6
g6B6Ar7uPG5W5r5VEPWaVxLEP8+izm754nIc/2niLLCKqYjpgQI/rjFk5i/JuDn3Dl0bAIhz5/Hf
pisuhmpOyHE4aPv0JUlwflCpodAzG167K+IedC5gWvmw/V5X8Y5cSsiMO0xAng8ZzCTtLTyhi0VP
NjsvMKBBFMVoPJeDEnlbO6/QNJqYz13rhjDhH8dkq74o6IzyrCeLnSNvkqjzGLgHAsRs1kX4bZZS
C48i2nYYk7oLBB05Gd+PKkvb8T9R7DUEqqSqSJ1FvnLa/dk30tSDyxm9VRLjiTEb7haDaXXA1j0t
5GsCpyVGCOYgjCyHpU4ef+q36Mg79dZW66mxOXLgM7ZV3ILrrFRCf5TyLHPFlvjtt8CqyHu2uCcq
4TsABjqxElPfMTu41CK+EjFEquya59JNQexGhlEw9wTVFxKblOMWkJEwU7WYOLH+5qV8ZYArwjNp
ik6Q5RJ8wmZGd90nrux5to6k+WcrrylBb4SpkMglSa7crCzIIT5OWmgW+D6jilAz8JovcCxblJvN
JoM9tbWVdt+B2Lgn88b16mwjreoQeskqKblfdshQv6BWjumXqkatcNq3O3DApLBYAgL85BgDenGS
+dHpJgpH3KJQxUclo3B5v+EJZiH2LiDwYs2OPi2VbfYFoYW3Piai8pwZkYvfRBDn1zcjr+HBJwXq
VOy/UDS8ut6V8zp0ODMEcwPPELz9xrMsSvbwafgLr+8SpPAm3onMIvY5DuzcCPnCi+IWzFBYT5CH
T8s0j0dNduSoSD5K+ZCwfIxJc1HkXPanbGUtxo5OqnBmlUa1EXFgdlKVx0oz16CzPYZ8OpF+3bED
r21wjtOJi6Z97OHBTKtFs95QZmxOJpbw3m+kpZXQAedyEJqJ1I1lCTAniJlgTHTQ147wJ/gixxdm
ZGtyUqN7mn+pl+UaKzBe0yZ0Cn/c0a7vxefLg9AV5NDF/+0kMA6JiL0lM02M2fZamVcLMbQ1e4la
BNQSbaqbAi9uIrDC6Dbz3zOUZIN+nQWWNe9B12k1olm1IvgbOqmj8Ao735FYNrlpZJQQf52MpWBb
ygFXpFvDKSDJ2AQdbDOwopOitMsxUxoxqFw+FPntlQlflNFJ8Ce/HReg4KdpBomMEgjrPLGHbKxf
06iUoHI33zrmXWbkrtEAsxz+xRJzLeR5wMwxFY1/P/uGhJCVvhwb6FshvNZPLh4FLmVd44sx4AVR
bQ3A+2KVZanwvN7ceLdKSmFzg/y1DI9f70Scqxy+3R5EHfoe1qbcFBE5F8fYAi+Kbu/MDpnncuOc
cW1BXeM+X4ZaQKPbOQNPnafey4sq4XAjN58OuTB7Mcix5oHoEjH4DBZe6SC0cd39GYxU5TUNPFJS
KW8RAgLHmjsWH2856OKQxAwymobILPUxn84X18JRZdpKElgUen6Ljy7wcuy6QvBwbgufTluNObZw
HMpF/KLOFd4+gpEc9oucRogUfljkV+ZgyUpWn/DdZsHXZiP2yche2HUfrUA5d/sMiCI4qZDJ7S/y
Oj+5x3nqOsWH39U50fYhzIZQxHgIu3RsiK5uNBy7h1jx/qfr5JIpiYa16Ua+ldo3DWdDzCEJBP1O
UM3NvjkhHQaLhRiA1tWYRaHFbFc0P629NWsrxItCM9K7gcggxfFOCCpQIx/Er45+yjkOkxJ1aKuL
jw8KOeILm3FEIb5piNDNc+nrKjPRGspU6ZtRE+3kocWTSmWMlmsEGYox3Iav1NOcCjxBEoEHdIpe
kZvYa95djFNw284NOK3K7QD8+2Q5AQ08tuy0ZF6FN8+NqE6Ol+sGxmD4tRErh7L3rp605Kcf9gMn
lvE95Gv+7xrUZ0gxZyKyFbvgH4T0e9I4sYPXRE6POhRlrJpY1XNLkIB/TqY6uP7iX4H1oBaBG8XR
VjadzFkJ9/lU5JU6575TlJkjQxDZ9IVAps8Wmh0XeGinoPrIFbkbTEgISNULV/u9oEemM0ELnNk/
M95b2Q/eN3CrgtNTdclba0POaaXKV+nPiu6DSrEc+yk1xWGqJG8aG9mNLG/wJe0619tMS2Fdl2vF
lF8uu7uVHis2T3wiIwNYccIbG9OQvPmAdzdJWmE3gHmYeI8DoZ36whiLWLBqKkYwJqNWrxXmtluI
CGGTjIe/SHzqgSD2NzDU9nJ5NcVmK8X9DxK1rA5X9eSUUIk/DCvgSB4Xudq+kb8fTpgqBCJnp4UO
Z5QrAg/I/DUh5eDcgDs8IxEaTWA0ujKO7HEIjoqRBdpjRNpmkf72gUh4d05xLCX7CVyhRgXOrdVt
q1MKYB5zc3zDwOK7Fih0hoIj+YtS4+2dcjSJwUIGxe4Zp+okjxMoKlcPDYHVHOB+Nt8nzhKVLWAV
GeSdGW++vunvgNIejATnpaJsvmI2GMMRZmzDyKlUKs5Dqu0ULcaNCz8dANPk1rj2FUjzp+PpsKph
XHl/kqUiRBDIclMQRsE9BzVeFsxNhcq6gJmRcy+fE7j5E5TVjOGOnt2XHrjtNTUs0BVP0ZZIMkda
dcycEe092TBE+ncwtusp4iYTtaqdh2kIPVIXa3KplpduWYBlrTTyYdoGeOSsXGvdxxwbip6iA0FI
8yDlFksuX4Mwh+ZlS74WPva2t+oHIWPC8W9Tt/JIRmUnOlrjARIJq8WZeQW0EztZdqmNeyeG0FDL
OHu4cEmRX2O4bE4pGfn6EkaJuFYS+I9tJ+fftf6djaq+N7vwM2re7FNc/nGZhadDY/XxVDbFw5SD
FS9MtavgtZYONM1X1NKMvFkSPwDKUX+huE8fxxQhCcB63eHfksWQfW5lRpv4dlHi6KpfDSZBBAw6
aB4jTbwuBANdXZ7YbYe34RYUVoV/YhgUMlDBeR2tpbAktl+pc25dREmOVEw8v/vg+Rfn/llKPdMU
MiTbAOfyVDDlgPN3zSdd+NDHEYs8ub//4QbwP7wm4XjemhxhAHf9DkBeMxNc0wxLHZ8vO2b4Ysnh
yBRGQs0FMYgy3MFQAKqCTOAuBXSKpclXTRpAzf3Pl9WfxwyDuEFjhtU4uWkpY9HN1dYS1hL4KOQ6
gDHX31tE0lyDPyqXMXBOZltyoeDx+sMCoxNCnDbfBqBh8vIMBJ5JJDnlWWjnU/Rb6gKSL8ezJf+A
O/1wk4OJJHZ6TMuOkYnkXxGX/15hP7MwBMtCQFeJ08KJM7vxhuiicPUzeHoCTJ8nlnj5PAZep0DN
tlDbjXc3uaNzF0KaL66XTxpuWS+XL88jcER9FmmGWG+k6VeZfGw+5ctencv/0rxNYOt5hQsfDyLf
UE/0SrPK6kJnqbqDM5mTZNeRfDzF693Wu6uwACKm7htXNiG1XKyVLkAFnmH4vSHXhUOUoxexoCkb
zd0q08BErag23waf7rAEYGda2BRoP+EQuIT22TPQ8n51DoHBdn/ypr+eKMk6UcQQnfvXnVWwfc9o
dzqLQ512ox2x9Mjm17Ve+vM/IzT+ZITrs58QnWNzBQtDEXKlZMi83q0FPcrrTbIuNWfYYmAE5ktF
H+1+gZKW3Bi1yETKXA2/argt8u5/HZGvJGwp0r5JfkpG5WZeUy7fRhoWgyDkY5UOXQlD+8iRUod9
QYGKIRbGU5aXfQSOIH2FIf34tbmSMruF+ZqOzNxOYO00AxfYwJnkttbFkhWTK74Fv7Ow87Qo6i7I
NWczFrASF+VX13haraJGxVQ+8pTH9I4OoHc8HronfEtQOStZBg8c7CvLM8N2f9drWOc3zCtc0FRm
9nRaMUrQFWx/1jRRYvM5tyWEDRapw9g2dXqtp4TtsRSfquLB4ONS4s1/j69tdEshpyP2XCqPif7w
VolYod4B7vLBVhG96EjSIGRQv5ZrHaMRPGjPUD2a2DrfjdP32UFkAjNGUWo11a/5r2lh/GPFJhu7
v6U5MFzhWi+EzsopBu6gok2D8yTjo4RLXn2vjOhRQQQvXWDzayXy2DUkKaqmlgd/Cnz2pufpQbE3
RGJNXzNEBEfCdHk49IvDqbg+F3yYeVdIl6ycWsR7Q/BdC8HqGk6Hj3LC+NxQ3vY0LesvRTaEueqI
ffp8foT6ucEpPTbVUp6yX+dvL4u884ZhGjyI0nLnVoyog5SshiuuR6JuIXoLhbYVaPwl6exPNZ96
yySIVPIPfIhoEClIsYVmUOGUEZIt3Njgfw4HZslWlYjZRIwdJXd8qNh3C/RmWs5t7MA40QtFCXeU
1MKf8LCp6E8Cuq/1JK6RXHxMpcil7vBWgwgE5+mPq3MfOi7XjtprjG3KyHN5XnBCMR/LRAMOIJT8
fvOs8SPBm2n1QCT4xha3Uk8huu2XtkgI5OBpMtpOECm9COSuIIoAWS5qhh06iM6a2WkMEt94n9Ia
w3NT2dZ69u13TgY8wWVZjQ2Ao5wazUIBwURMSVk5Ofhytp/ZBgNm3MwzpQn6gi8s87v4ABKxGGtG
ME2WNEhXGdc4QQW+aQOnV/eDAAahLNNBcad/K8icBnHC0QH1vbGrkodDPzEgb8lHh+rFBzd4YNC0
kfTaOTqL5bGHjmodeAJI+OuqvVhsRCeTSchr+J991aeTRJT72FOfbeLrRM0zkgj65RS39d2K3W6b
dVEevX24twp+Vn08UOzZB5dS59zhureFPNiWIbbjG+KXLq2VlY6bduYRh8GPpScrHS4L5XIxzvHm
M6MVvVSHvePqwTFFBv2qrlsS8Cx+oa9M8VeQymq6vXrJkUUoMIZIO4MPjmh0PkdWqcOGhk+0gBWp
P21CqXbWq5XdJp8LHuDATvk1+m3iL/xqA3AoOK0vcsHrwpIOB6W7MJmPTxPn3ZaWlR6+8lYaAhjQ
K8UnykYUaY+oypuGgyXjg849hTZ21iOEPIbNZHfHzMZr3MHOaw9GMzH6Xs5aTB274XFjrBuRPkQt
eelQ0dkeJHsuUaKu1uayjCxB2mv+kimUzwsD1Yo7JIbUP7KFxlKH5sVSy90BrrHGpdq+Zkfv/K+a
CL5bS1H7+uNv9NhSuUEkLAo4iE+NezCwoDilS6MBfS0scOO1yebhu/aK+at/nuhrsLw4BcWX/YeH
P4RPp4YZKVgGU1FDxKtLmrtafVdnx0Cno03uMIsDOeMDrvW/ZE9EvMHLZOwqcnt8lZpXEilMUF6B
vlwaGs//iSTfVZLny9TqCp8JLTvYar37i/WXCAKX3ynasv/egrWfI7aWHcQoIULhA82LXKyk5F6v
AnaXyQ9JU9gACx0mM7NaUB0btVDg01vYUiHkxbbVL/QJsfCIbTTYM5LFwP/Wi7P++UB16RQCUoaQ
D/Jrj2PMG/iQVlOjMBw7ufghBsAZnoCFBLN5Hd8iDziGTHZoz66Khp0QpsYDHJj5JIXHTdsXwrid
5UHvEfIJrLGsC1v+lfSKVyQjklbXr+thLxCFgKE1KaGsfDTyk1y9oYDxDE/Ww8hSgEoDcGZPPnYv
MHlDxWWZfZh4TJPUSI6liNIY4zk9bGoSR1dUvFQ5vvqyHmdn7TRJSt8OTiVep2v/pJbvFkDhxadd
SrJaweZ32/7tFaQviTpjTzL97hU63F8jNTA3nnZhNU8foMfLY9cHDLzxDVejjUan/5rZv9BR9sA0
LMIwhqVnuViBCrOBRE1HZUg72SCjOQtsmtqkcRMqLFGTkDK9RM56AEo7c62oMPkz0Zjrqdmz8BWO
b8SHJeKBBmPG5/AbLuTy6K8pP1e3h8YGQ3I+d/d9wVRp2GiGqTNWRYfPkM61QZYzsWZ04sT/beuS
RXLDh7O8y+/FiBXDNUuJGw01Zh/5XIelFylZR+XfBkB+F3LLV2yQzgs9LAkTdmBpimBucBrtIQvn
NyC39foybhZFpn6E/FT3ANNoIF0I1Y1lErBD0BigW8ml7FWCtvSShr0Z9hKJpd5CE57I5CY68BTN
aHrRJIs15EJitJl3RDY3gfVrSobGpdc8NtJJjHIA6RxLeCZtpt1B7ylX4Xc1Of3uXYVzQps6n8tg
vZ2CGK0isoXX9WDLV3dsaw9FU19fs8bFTgZdWWgvfQNHKuvxu0FskbqKL++IB7SSuB/RBxeGvcWZ
h8CJchYSyoYaol9pD+vpo2wYelxlCuvqtQvc1PX9XHqINMytjQUnphS/5xSPgZIJX870ODchLHow
15VRlGvgQ2CzMqjZ2hCYTs5kzjGc9xs+BKIRZTvjgB0sfzqQHMaxcrE3Yv5er53f+VbC5WPkhaAN
cekqOfUr4gNPKNlIOTPjn++D50oNHVwLl1TgcaXVFK9n7ALLQnVCHwWk6IGBYomx2G9DmVN/1dmE
GaRNnkQALCB7HxQi825B3uwdprGLDNL94rtU96KnXDNr2IzJy1szjCiz/DGpNio+qlb0p+rPGo3Z
8TFVfSlBystA9xsGtM7GM4h8V7/SJX4k3JQ+oILsxmHMvTe1UXKydBxRbY5TI7s2ewVrfrzLvX4S
Po6I3yeMmKPC213wip46ty4rFbBVhucr/Ixs6MIyAOPUACIn6bdOOaxu4bs2mdZJvljhKpaAAuHn
NHsgdE1Q9ZO18uxRVqKgIjHXNx1quHUkBVlXvwVDrXacgYE/ING1uw64768M0k6Mw9kz56ZVaKqt
SgImTnkn8wYxeZA9Vobe/grDh+3vcq4rXCsDa5bMQUnE5KZjNnqxYBZWnzAxxC7O3ZCqNv1vQixm
B/q3QFPgtqbdXgKx9R0OYFSMFJddJUdBN2zial6swPaTRTAJ4pbHqsHMcFzMJyPAEzcstYrF+/CX
SjxhblvS3WNKfjLZXjjji+3LDGB50oJypz1lntszQ8Z9RxI1wI0b6YClwQjeLkWarrwZNIgVOIgB
G8RqMRXhrnP9lN6BHWDQ5roxiWSzrqAl3uVPfl7HzFYeTr2LWRTbTBB16luOUjKlhHq93ecEleE/
RJ6/pHfez4a/Vd00ONAnxrNil2DMUS0bcRbUcvGqnz5QxLTGE3vIV1cmcfmNlhDJ/liO9mbNjTeK
JNokJnMNDdgFynjqHXcPSJN8H43zGMYKR7JAe/esTt8qw/pcAQ6A/Pe4UkFTQjbvouOo0Im3FJtJ
Jhco/R8Y7BeYYxI9sBvMeCQe/JMC2Zt79LrOs3yMGxZUBPY2NYGFxMqZD8tTkHENgWrNhHf/isbi
9w6KN4sh5h9EDjygzuXopCwTV6pAk2MH29Iuc2Ocgr0kdH3jLcbq5vGVJkx44QJjT9mgicKiFdG5
6PkzSJmvAGSQTvjYrZorvsb1yv9PqIa6oHSc014c6HOY0YSfz1Q9iFN8di4YpCFxQqW9XWw5Istf
SFKbypmcjqGnxVYtP4tJTGf2i2ntZC6nvq4NiaUGD6xYmol/q8TrbktjxjYRRUyw3OGLZA5Qgk3i
GA4ZmgPaTl28op+zJ74tM+9jyifeAgfOi6SpZvvim2l/VosbAAMK8bxxIc7XtUMif92LJKl7A+dl
h2UtTJsB6Zt5yWAOxcaV/GCF+xm3mH2D5bD/swq5gCaUi34ubvzXRmur2rt5olMNdhBy7F7dmZ54
wpd77AVhkBIu2W5zp4sAgtWs3hwzXD6kg4HM/PdVKfdgi5rJP59Ur8hFK/ifBJ9jpXjGQvWKwZtu
dQXkARQOrqsta6t+33baSqn+lGDK06GF/s15lSVJo04VOFFjzCpnmQ2OK/txL6v2+kpSbqPaXnku
N6sO0uT6vLCraR/Gy/lP2p1wDUfkbbUKopp2XI0giP7gBn3h3nvLw+lbqUEH/gZpAxX5qb9HPvbg
ix3NGVCJR2HhIy2gaxuvPm0LQE+pjXrZQyRRQrkbjLA4qFdFkIUREXGCKkh293ML7Q80g35+xJih
eQNVIDC+Yfbz6MeNCouge4CdU5NAp2PtA+/nCJ3Q+/PDxw/I2+ifxrltHamAG3IIUwqy/iCQT47g
LQLzFlAYcRxfIWyrSlXJiboGX3uxr6yhsfY6Z7MIBUkqcCSp+r826ITgXvyKSeNSKnGBkaNh+qud
r5K8EzeXMGHogwrwt8tHLhawvKwSUY61W8JiYkyoCqgOh9/zRxrPHCSb23LmuWMpAioYWpC6R3BU
uLtpv77p2gIb4X6lAsCycA8lHREoBo1ZmqksIrPrT/pDdqvhWrHrpBamrZZGGNtl+XC3e7LBD5/t
/CIMw2PzTRyktLUEXTMU8L53Ww6yBm51lL/xGOrc3KWgwofLXA1DbQyTdrUxHRjz5hp8UO/Var4H
wKKgs6GhGhBWJiPN4p76c5oAE0F26EWz4ZKavezhBscZ1jJxQrmw0544yVuQ9Pt9gyuYmAXDjIgE
i2kEUiVI9Co8i4sgbBGS91tkFbTHQcysthCOuT4iKjpAIvgHVzLrmWbb8fezdM2r5ZqZz4xAFNDH
xf55CVnMgMbhGjb3mUnk4wzrp6Zg10LYqnDFXIqg4gJ7ZPOPIYsdSwAtpVxJ0YYeDSJ+fh3EKUEZ
oOMAmuozXdk2FDcNNJoXDKBiucVBgG8K2IezojbxRiy9CYurej7dg2QuX/lgQhigYlCMWm3Ke/bc
QF81AywpVF4x7xKTBETjRgmGJKXlQIe8HJWXK+u2sbLVRswqzMn9ibJONh4roId91PAZi/G3zuhr
j/mU9wmsw5qw9IFypc9pYBN+LUXWI+iBu+IpxjNDN39z7gg04ZbWJct64ckgB2etKVYaRdy7j9Bf
NLtXytQyrJDSQ15UEUNpCORR2ZksBXs2fWmn2Dz15cJ5lOxiOddqUTiNJbpmtZFTV7+mNPbWBTLQ
Er4zSeo8xLvfvErhl1E5Ji3dRSi+AQl6J9dQ4ipl3KkTzgjJpKMYEwNDup8rd5Dm5WcH+oSHhQTe
oJMk05aPmiJFoLNB3DHEmMh9WrqWeTbnm//uvKC+YIrb5RT6MN1tpBlSjaNbOnnqzJ3A3SwSSIS1
DcaNyixioVSmlBhVsrZdvhCoffdoiWqiCc0SwJNVI96/NOUrPgYOKkmBwsmh5ECciYIyN06+5jGN
AdEuNSByl0AbQ/CGY+Umf6F/lTnipxT8JuZBMVRSejYJr+q06N7nWcj/JOxKw86tDbtFC9gwRFz2
tsBHdsq8DXot8M7gTQRKHrtODzfq/BF+vY/nHR7mWKYGiouBO2IvMHn82TuZ4B5zQpNx5qA2HVGU
8EMkDWbqrr9LNMSlDpfkvuN6NACQNa/5NQoJiKHOFttRFcxvlTbSOQr4+yhyfqWeYgcT4H/FLlbD
GjYvemElUpYPj/citmvJJkIHwXAGAjCKxDVJR66oIC5DjhqDkhYxki/X1IbEAeOVRL+0DsUXGizg
DaRSpYN1bAbkMB2SgZxj7BUTBYIhSwW14wA/6FVjTo/oslcXE8UVWACimVyArL8MUhayg08/G2Cu
xDNGo/fuJZWIeVsZYs1FXfE5xB99WfkTwmxcDYxd17ZHiO2jZIBsUduf8h6lcAUeJ+SzfZA5V4Qv
6rMMs2l2b5OQUsGgA/ffJqIuwAwihQcBOw99b7PlR05JGcmfPhv0qOzC7oLlWlby18aD+IzU5sfQ
NU8N2brV49ISQwuywS4976krhfR88jtaBu/uB7kxUmx0hY+gzm3XNyLeFET4oE46heGzJNS/fQKB
IO+stkkTLzUheDYquGHNSpTgOguLLarUr/aiLK+L2oaqhQ4we9HAibkTmoDVq1lXBRhUCQaqPWIi
7vEDLTzQrOdo6cfg5CMJD3qHQ+N2ISGafHwIbYgBQt4/lV+0GmQgQE5HsOvOOwa6O3HC1AbyYN9h
ZvhrSriyeFPikRq3EMY/SnwGtFXXBQyYeOihz77Rt7+RbPs9qMoiU1vpPzF2jXHUwjLtowG1yiW6
HY993I+NSULWJ5f5Q8T9ErFjcZVAT/glXnZZUrXUAN5EJWQcYgYEprZ1Vqw2kFw7oUBYUdv/ta4H
bypbL7FudKGfzu3EK7fCh7hbNe+f0GZLVTgTkhoNyH7Lx1CXgWjOMvtp6/M27I5DqDK20D8DCddi
smHlaGoa898Y7ExG5ub8mJaxiqS87xdaorRApcWm7XU4B9ThZyGHlDwdPkhnaWxjvLHt96gIRV8i
xQWoohh6vunk9enubqc++DcwFIFks0WQyiv6fRa/2EJnBmgefX45Cjop946YLOza4YcFnc0q1sdp
clxxZCtRftAJq/VRt0zddNCTJfVjP/lQAvhS/LYR8WNLthj1sA0hEuVvPhg4XCMzcxyea8yDDFTe
xzQ7QGLFnQ2TcxHbfa9g2kHxw3Jv0vo/p+oc6bLi9qYDGMQcml6AIig3wEr+fOLqI1nCXLHz+bX0
c7KbhNecpQE4Fuxkx9F1EybOIqj0CxXls8J+tOWh7LnBw9Q3SJEs6IsEKVgI/jsgnmVXhR+qcLxR
cc+sLWfd6ue+OrUKDOtR8vsdleIfiOEnE0nrmI06I/8QB/mMTt6mirnUHpHB0Q8WPIwJ/sADJlGn
5aVHpzpe5HwRdTNaLfHTE8asXYmdi1Yzg/d1zfpO5e+vM7CZVcSOc2aLrkJP8SDKi2zlK62E6Gi4
YUpTYqWmgoxtIOMD0t7Br1wjQShxNuJkrfpmKNw0MXvpQSSZagQ0g/Y6xl2I6OLJ6r4f3UGHr6Hu
x62VDTsMe0025k4z6G427XB6K0vF7WPXOiBGZuY8XTnu2VkIVEacwt2QhLYbqM7r+Bb5l/g0daO2
cXbUi01Ptwp12zwYsBVkWG3AA9pjkr5E76YgKom2enMy+PY8yBkfl9c3hbazd60Cw9LUQqxjf8VM
yhMa1rgN1SkGAP5JjKymKCu4T7/cIVwEWHhefkHN6lsbdi9NjK2+H+4DtmKA5uhtzBNXI5K4oUGt
/D9oQZqQlTae4GFpGHFlAGyERmYN/nS/kJAokMKwlr3RnNcukdVx7FeGgfP8HjaGs+wsbkT/0jHU
3m89JPwXGWif80TnfoqL79X4T0z0eGUlSDfENM1TIJJHAVe8u2CkxpVWKkpo8tUtuAyHgUvw7gae
PUFfRExUFEwdIFUwq8p+NIGZEg17fE1gTjshP4yT+urW1M9hTqWTf+T1Etv2A2PHSLv59O2VoCKZ
4aEmOnYyvjkdh8Poje0ptOZujC4hwQI0IqikbYQwcXp97kVsFPqkvv+7n8F98IY+d7qFk5Af/z7f
ubM4p45fTQ9FL0duOcsyYGbEHW3YLt7l+uEJOTv4G2Vo3jn+nP6Dve53w+9z86fgfIMVNiRXX2+9
295tTL9qkztEze9Pb/i0R3u3L4E7Q2rReuJovtdukxRqG2l4LPi/f8PIJJXVLz7/L+kbzSxjjI04
PCm3OaPFYA2C+yXa3NkoVoN0UkbDlZ4DKKwOtw9uKX3k1IaINbFqnMYTWkArU1dRzgIqsIGBk1SP
rujG0QG5GMIQMIG9dSpv3dMetymYLoPXR5LfwbydutmHQVYpNFkjSceHgexguZ4Qs9e1z0YJP6ai
hKdF2E6BZN5T+IQCTHZEabyM2Jqnf5zr0BHyCV9WnzglVGOncG+eBJbykA+D4efije4nszK+v5e/
yqpGdXkcTL+0R1L/GT2+7pAulYc2L+p0+UVp4azKCtNkpQB+cwOozT6B2QyecfESxMWeh2vvi5yN
0Vf25LCwl5DmrEwcAwOXN05hef+cO9viW0Xbcrdfj9sbTi831tWa90nUFJB3n5WeZgUVeUEoun+f
vZvrU3oruZfO4KEff+UrjiS/XnJd4foKEB6m2o2OrJns1CWIO59eAnP+xP3wyqWhuOqaaEqS80rg
kpR7NNaroIpmIoQK+9qeB92KGLFPMWbn5d9h4lBknyZbHavsREhhR55y/KikbLjhNkD2fqcwOoDB
uQS+BqlDcJYpdQ0/2Q5bJkRnpWjzdzb5YCDAymjNh6Fa7zjcEDKLcSs7dOL7DsBkpgjTfmWLhMoT
R3gG+kwndcpGjvMCExMACUT9JGKHoYz/bWWoHoFSmpVuV/+TcfrF0Ce/uPIOk9pz+vah/RYbthyn
B3SrYqK8xrXZs306I3naSyVCENaO63nWQ4zJjPsAeupWiSUayy6EfqLBaeDcBXYjJFnqHZLuAIQf
gvSX578Wmx4ryXF/BmlB17aCkP2nZkNu8CHTFvLqgbnaH8TD79fAzLmNgYr/RJJzDBkeIqytZy76
7dMDUcfytPdyAjbxcgswlSWl2QDXc5J4HUjXyUTY7+MXPKke/JxbIxT4tvAx22gr/VP74R6pUjYj
BbAnLVlMeNS2HdHKHZbaP0I4rw8VOIvS8IOG4+axG+/a8StInNOGd910mNQ8YyZT90J06PmurKUM
Wvrk4tpCWSaWxONg/Hs7GjeMZ6TUv2ttGWlCrm+SPzE33p+5cln8b+DdDblgH2AJx3lTJ/WGetxA
Yc70U/77WtQeIdF1gsmBMFHPJIZ63wPAg/ud98xA28Tsi6nvD4GpGrAWUzeyoe34ZhGlWvlG97Tp
OB5ETUolebIjcNUKC5EAtCWM03rOgTFmD2ZxFeqUULgDdM0CT0f0EkDMGVd8qEQSLpZgDVjAUqW5
R0soMEhy1ZRnc/FoFW2b1iGeya8jqRP2ukQX3kgBrrykEO7w4bai3EDSEL1dWkDlD97ulAI0DTUL
RxciVvnpfh0XUg48IiHHKOaan5NU2qtxteA44JWkMd9Wj1haePAfL/Au7u5w4BzAPmPlkqyd4Czy
ZPMsQozLVaU9iC1nAkUA/bn7YwA9+s86rVkJDf5KnpO8G/lnlMU0httsGqLToG9IXHzQImCLcPVl
bmTD19xzkjiCAOhZl33gmMqKRodAVxbfqtkj3u+jK3Mqr40MJD0689MMKR1tgFLeiUaai03gsrvq
dpHkHKpIrbKshLj0zop+khbzjZKBoxG2ZwsWRC+iK+TA5Lr0q7pDJN9qqvunUloKQyV4t+V6IfVZ
GRHLPrME1KBeysayd00esoK1/2MPRjaH1NOQEGUvdrYYEHbwkT/zFP/Z/a2JjxBbXzg4qEiYkxBo
0tr20Lo4OaiaT+7OXXuZkeaGW9RuVtCNgnpNi3AqObIsq9uINMlxGzjvQ9oWEd7OkWXIu+lJ1oYD
xQAnMKozWmz/rKOIBfkfwTrop0Fb2EEDf2ZrSbE0AJOXAE/v/6tRm75v8j5Us9FOY/bJOEXh3dPu
KsTafDwo0//ejxdMgDvhk1na5M0PFwqjCw656eKaLvvD0lohr+xCruMcNISQolvC18QM+TMDpS+5
/tOjhocBbR7DjGwBFl3Z3QkiDB6UYecAB+63tggp6xUVYw4mghM3HXI+UQ5JOEQBIN/dYaUdkqeI
5GamoosMXTnmhlirSlgH0QacCBYSeyDde3gIkeFYItU5wn6oWXy3Is2tfFz3zGcR8t8LZFn2XssP
HoaWhqputJQ7rXi2Nkl8YKDPIKtfYV2KtJ63aqxkskBbpY0mhn3iQnCNb6QBg53U2QWDxnRsmDwV
yMrOj+GZ08slxxRboIeqhRTD5gfPkjTjTPKcSgVLI4/CtpDW/5DMuOTD4l12pmpN4vVirFAUUWha
iI/TakAJwzAxXabNDyG7JrwqwBrasi6bK+N8IRLc/nlb6B8bmaOnw1dzKaCvhrSYWjBzTh3M68lG
zgLL8hkgCLVa47tdrYO2yoxrKfWWBDgyi0Ec8Q2dKcFFXV2m2fjKB93zqP0tj6J/31nBxktRll2K
zmJFvIVSQzBGKmxg7cfYjy+9G4pKPuvqTUUfTYEZAsWacznaILzU6jD5ohJ+4xXK/ykipVv6N/+T
2iYHMYmDbKY14fxTQVDOcPy+8rDAskOQ4Gs5l1xKXkB8NUE/DT4G9Y/IO4u2j20x6pTQIWU2fwHm
kV60J59rm4S82HO4ymLhSw5huTo+LW+DDyq2OiF793J0NnmFAN/NDVaUgZ8fBaXrzVr4orzPeObn
EBrIQKrLbjc7dwSX3fODUox4UhCUZ5iw0wicJWL9glhG9JhGt8e36rfO8HyIzBZcUPBqUT/2lolz
0mjlkGIKVBqEdZemph/zEHh25/NuwqPyTJkxLDWb5JVKuGnLwfUjIydWHbDYFljcVX8o8LsSv97s
161ow/pKN6JObwDarxZgE+9IpeYSG4cbkvF2nav2ef7LSVhM2LTLZRJGmTmPBjBIm1sKQGcSbO8k
mBQurhqVFDKFcCnHSKo6V3d4DgppIymAG4rp5UTQU5TwAr09S6/zqpes80WXza50FxZ77BkXTGPw
KdQaEe3S3j0Ki3/kztzsG+W3CjJaJowfuR2LmmSIR2DJ0aj5KYN89uQBv5XfhLZyWnfeyuP3FbEs
YUVl3bGlnSIF8LPqru4yIHutWXAgUHyocnxgLiAOr4triGvLAOeCM4adQha8n0yKqN+BiZAqK7wK
Bc6eclkHq6qniZTPiX3qTHq6Ad3xX/mLwwIMYJG9aCZzLu/3e8HbHWBt3QRtDyYk/OuCGPitM6WN
PMHR80G+GIRipLrehZ6aklmRnkJxxEXHRhVsMw8nWyhFKMmG022OPaP4eW30zXeLuzB7BXXA23Ok
VKen7eoSY1W/jR4irLCtSbj3LUCxmKD8rqgjuBI9exVgobQxtFIU98O7fsY3Cy0FVfjWVXeyrA5N
z0Raf4mBivABHlQdJgwu8nN54BLiEFOvK/zBujTRNRU9Bb9XXMM8hIlrpcvHwT+JVhfkI0X4k9My
Av1ySqm1a6V9+Dic6ZQ8w3Ao2Fyrs3M2pkCBXKdxu8AznUdEbn3DKibqvuufH/yWKzCvflYeSeOQ
H63MxwO3Wa8TDhsa6rznxD9iYBTw/IDYY6priQ1rq39Qy3QftH4Kp7ZHgIj4URr10FFWeqsfWkse
dY3ToupWhOdUvBlfugffk23Jfu7CZiksrX3vSe8/S1bAhVQhEE3k+IcDwt/uNuYXWvqUA2nH07vQ
UjoMyVreSy4ctJZ1i+N7xnrELT4L8epY+lnDMSp/AQ7NM+wi6nmaY1K9++ouQQGy8wZOOLGm92so
A+l/k4h2VFUWIJjYMc6zq1iDBqxZ2FSUZBpOmEMKFDbxJu7xz0b4FvNLRBlVtsqBDoww1y4ZxRyg
Gpc0bwB2AkKVh55FCFH9SF3XobupGImKO4njF4WAHqgf3TrhMiF6qMU29NvHtfvhiBuYQBQJ8f3u
/waH87IIxDccD0vAlwmHEX9m2Ivmy+36ZpSUcKJo/J/xbEbCK5paYAa1zhq5D9Qrokvp4x0ESWkv
nNWIrfN1TqTQ43yscXwO3ouisu8E+8Sz+oiqXHS4Te+EjBW8XuwfVM+s02vMk72W/6S+zQ8slCJR
rKxWzkVFwL0lLE/ZL1qKZejQ9AcDzZSjDTTnTvlW4ljF6bf+XUJJN3WSZp3fElOVnxhJZXdyGtua
dLdCqsrLEIHJ9l7VN2+QNvkFr8M/iWNmJCAfoazUvI54gUFlKjKiPA100ldIsflQJMsKWSVIDY3l
yc1ND/O86KDdTbCnkEpGJ4unAhHMHMO6sa/p+idXvlJFXCETYiaED+byet8paSFu/ECIKedZMXPM
fPEsXuZQxOcHotBD9UoOrlrqoLbW9R/FOZTSAfmnIr6JfaHbgH1C3gNBDc/jx1v8kZbXN5E6T7DK
OVlfutt+ZvxGMZsZF2t7cGmQXqc8a2apWoVJWw8pjpPp5K/Ab1K4YlzovANv6tJhxw6KFuMBquaY
7Rq+y/iXanryqr9xctujr3M07BJMLoNl/QgRJY/F7+NywOFIIbg3CcMYYIhxUgkdp9GeMjwByPrF
sBuI0zQOnkPJhy6spsi44d7xlu+EEx7Gx6C+5a6rgChTHZYB8ai1dbVwqEO52A3C/PwOwVMg5Tza
iuz3S5gcml5Gs4r8T6aoeNRCRze2LDXDU3Q1KGYMzfLxf3Bq3+kwewKKoUc4GcDMGHD2THC7TNMH
HZVJTPylJS7ficdwoUb0EGEwNLWuubBq02+fucPlnovLBJi5jY016xnqIrxbovsXqBM70iCnXsxN
nGXgVAYIhdMushW2uiqNjqdsdR41ceoT8/8YZPehhzo+MZMimBhMsxg+PUYzk0yolf1UkbGb5zRD
F7/oTvfxSqVRHQntgU87kuCvM0XK8sfiBNTi+KpMtZ5wqQGpSh+x+RVXbmmcDzfeLVAvQase7ah9
UO+qaEabijGtNQO5lJ1yFA+fEGGC9AlKiN0A07bnupp2yKoTYb/Ag7POpvI24zoAsoSqcC4DgnuC
OCgKda99dKw3Dhp/xycBFU6Ln7mMwyB78qpW5Wxym7oYDW67387JTF8LShsqyhFulEGJiRfvXhDw
Ep/mDc9LqoWRQW9o7Kmifi9Ay7YPnPWDciYsPwS7EQ5/WaZ/EMm3dZpAYlXMAWPo4D/qSyRI9h3M
X+NVi0oi9XkU0PMmfe0qGwmwoXCaNuLCVGbcracyGrjYheeVnmWwoCTn1Mce4v9dfNKo5JtOskZL
hic95JLBbXg1wjuZbsGBl/rRNMG7hil/D99/81MQnygVzGIJbohhbrf7Anh6vxxvzF7myoX2/VlU
0x4pPuDqIpCECAgrGAjqZgNUXK3y0uvHHqI7OD6V1CwFJGo9U/mKRH/ORzsg7oAEom+oDSZBah6Q
B27oi6S8IVhohBfy0Y3e7+RRAuNKLvWKMTl4WfNorKPkK4g6c9W4LRCNq66k4KEcBFRkxUJxhem1
scXl3kEAgc0iXUM4lFIw9EUrdYWffDN1yPQxaP9QP7dHtkD4OUF22mY5lL6xpNGZ8DHSurOOONh9
3KMYFlTE/iRffbrrM9LglH1omSTLVePegtzs4c6jmHn6o79ftPkOrxZh4AAOOJ01kGOIIbs90FcD
PL7lmMh4w9I82wDQ+GlEZgbTVE+2v6p9ZqCkjsHhRSGNkdXuPy66Bx9PPnir5pE085qZPRNRuyik
nj2wuYFuaxS4zLVSRcb5TCHu4sS8a392ebIU9x/XQFJHd+OqZ7F5OnbeJ6LkefLPyHnme/1YyMNv
UPb0IjsSnSs8vuBAlpHCuon9GIQffD+dnPrluxclfLkLEPGnZ2+CjrXXCWpcem1EYzjqLhdg2R99
9domTYxrXT0yVAlHcqZxfFcrsd87s6nJHAR1CZM6S4i87SbhQTtEJOnbIJ4qbB5cRCO9saxbWhFV
vZyri+AR0id2bYnG28F+5qIMxHisyZ1WKNhD5U95lllB1jc6AJ1P86gVCJ61dw77+ZNWEVJ86C5A
NbsJIzSEO4dL45iQDVloSbB8frQwJN5/Eiq7hVYa6hCZRwkGDJSIsl7GkWCl0HrX2ipXo/QsIMFE
T922f2bLi8oYTyDpx+Mgn7qgSmYJEGAiX9iJAIbdY6bfqrhzPw4OPeP1vYhs2dgtYwxvxZKWyH/2
ir1KvJYN4NNbgSarAKzN4WDqiFwC27LmhYDJLuVPuHisZsfJKpAoB4a0TVL0zoyMQMOxTcKZoDs+
g2Uod8h3JRS+aktL+jSjfhCXsztgG5p1dlNqg2jd9QfOt/p/1iN/nOPVtletTidODdteAXt+ntI9
/vnFXvmA03mTWPWIbGBfni4xGkqdvsgmFhiS/J1EuUXeL4xrFBCMsy5ozaLUrbo/OUSlrEtoBtsw
q18bip15nfqeQlcvlUqXArkh882uPqqD9bFR/N9Jq+OT//Tbq9O9AaVtah5GRfiJhvsYS5bgeImO
8kPTvrNZ3hgVCbAG6Y0jixjrAmsjXKzpgpOMOmH/CR2pCLAv3g+eT35Zunb1/SwKTPM+d604KCjW
IP8wWvd1kIB+VTg5Qu8JNmk2IcwzlqiKzLQeKR35YwSlVZu5LKIZf9DFxQKYzaEcbJxJAlviA0Cj
0g5z8QRtu+jE+mpcjzF6jeaZdFjZ6GEudow8A4/SGvy0TLvCyBVdWtr1cT9gRRDn9/yPmXbqIYIE
4SiVpytwreYIkWkTwLPMFBBTMRigxh3oWVTk+XF/oWR2do2dtehSZHUHsASA160Xx/RHHyRl41W8
5JEDoSdJrzIIS1TE6/xjXVDTbMU7whfS9BRtlWgMT3szW199cXSGBFoMu2h6sBe1qvsx6Y7i5O7m
vVwC+TgKbKy2UDg56HmrOrEBp9d1FHMnu182FUvlJ8tIYWEf0nRhSoIxdAr2x6YLaQPNenHChfoe
lFDXo3j5BVW27xv7U1ZgnUVUpHvAw3GzFsse8NH5vqx61EOvFrDyYitBH5bkUEzrege18O+0f/3q
FGsMlDYEu9GoRLQA+BmwWbqqm/Derlzkb1IYeYpg5qlvqYkdxxRZXqpp9GeUESq3okhmdmpP3zI4
UaCiriMIXui5j4WZmrvdiu/eDFhjlS5288VDpCCldAE7OZF2G9rHC8qseIjBUCo9q3cu7jqyP43n
RF3wX6WL50aBniRDmr6NfVYQReoNpDixcqFlzZcdJEx+oCj5ln2jpHclI4u5biKgAZHLdFqXjHX2
vGT+m36ojLYtQyeCr76qM0eQw7rzJuICrkh+1BDr9OiOtBWXAr+pkMXSi9omIuggNl/bReIkZBnO
WDhqPf5FUVffwKwtzPjcI3eq64nc8OKAlr1TDGXnlPhH+5BxNgwNxIt6dveNHM7M7g9Hm4VFhIhx
qw7hhsDH0hIuwZvzo81TwImzbawKifA7QDrE81URuyCw9mPM2zTdbt0dlDrCCcl8hCiouRLoZM0P
XBCUVIynIMOEBUEMCo/9X9uewvj39MrHKYvMi0wddnqAe3OZVvAcWFV+P/YkZPcgUilXSz30pNNr
s67gScuZjFrEbhRc0D0MyQ7S3jfHofZf6g97FK+JL/g/Hu0nZueNI5eHDFQ5M4t355k+/0qaa6FI
MWOOG804zzFCa5lEA2Ih49Jn/kzOgGp2YhUeIVc5vdGMYzbyddIYyAp5ZwIM4muyArErsR7Fx6N9
ZEHY8PKrR+KcRNxrc9hrg7rnuX+UxDAnhY/acvP4znvHj2LJ/B1XwI3fYsyIIBU4gpR8eArY6pLX
Hh5jtQqL/N67NW29PHwLnQaYsMqHHnOfcRS5YvQx5ZwLjBfcA3DzfzGs9YdDvyRTWPO+G8RvmT8f
zUKEcpQl3us6FpLPGIuUJrgWa16Xa4MypJOjhuve+Fk7OFHqwYRsB3zAncu8eKAnc5M+0LBN7yLc
A75D8CENgHwlndHi9IusvVnjv3REBGGnH/h++slX4nGpc/7MHSNoXDRtQKGDCU3SlD+Ggd1a5dMg
jiSg4jxTuihlaeNx6vtx5cmk89dmRT6AzjWnXKx6iEHjPbrnsGoPEVhCMw3Xr6gToWc47hTTeLGd
fPj9DHChlCtx9xnWShI+Fgs+0gFtunaX2/YeOn9R3l+Oor0+xJpJ6htfUKwdG/qxHDBSnE6SallW
b/P6bEMWeuVjIJ4mpChfKhH5zxgFtbreQ8F/u7EiwOz4HQGWEghx8umgp+kBVs8+Z/GjM0T2GoPm
Xu8OQXZTmGlIm4YJRvUrLa6bhgbd83YjzZeiea9NiboyJGG3KBwozvAxZNNdwdNylZ2l/LgpUnq9
AgvN8osD4uiH7GoXZYvsRzwCynEJLq88SGvBhgAU02C8XjeKd5zdsbZPev9mVMUZF+s0fHec4Wje
ffMjUDb0SFBJa1e6YWdASao5ESNVOIWpoNwv49eCpnPJiLVLNczNd5XsQJ6JyTsKqgqZf6/iMR+m
KhbZAr7pqs4EQ/9lwrLNSqd4wSIEE5cgdk1G+ZFyJwNT4wf3+vjqQvjDDgQvjZdS8S5xAz8pCDkz
8uJD4GVIVq7vTzKsvC2vxwPT+ht5XnkqyCIxditf5mcrYWhx7ve/rHogA4L2E009aeA7skyRprd3
qTUwqe/7dYpzix9U8oMjLO8cRECaSmk1quH6EH23ehuhkT1kDPjfT8JyN+2+a+wRdT0Htb/BUoGC
sANmqiNUGccMaIVhZDj+gMZt/PCHqRjAlY8f8LDjR+rYjwI1sQ9H5MnsUZ6NQzjv/Ob5HKGwhVgB
5MKkp/rxvOTLrTvqGbrWD+2IV/E3rww+pf7zhneWJ33XLuCafKTr17B7EtHa3ttRlWJ1k1cs+WRw
wDo5NuCHaD1jncDMud2l1kaPOI/BBXUGcI3DxhJzxXdC6y/BitGXR1L9WbTaC6bEV5VUPRE4+6G4
TipsPM+M/UOK7wKd/awBU2QC2elv98mqFCKkq53JjdwfJB041o8suoTpVHyT3aVGB3dkFhQ1d/uY
djafaU+FFwcQWQuCnoY3EJiaAwwGNonvQxLkva0GXg/4/z7bmbCZ6I+pgh0XeRTGlWI78N48PeNT
RCeFAE66WjNsGyNfwnTEc3iJlV1BpMcoi+aA2+BsEA8L2YwYEopKYW4NIjeyHPcncNBf76voPQgi
dJu/C+lWij0FEMQgkRAwe7jQLQniQZk71+6vtl+p+CMTlZZRK2R9X2OS1BL7jun5lrI7fmQFPgTT
u2cvyEI5HJLfRDRJCFkzpLaJ0/aHskK04FryOPYVsYF8T7CU0xP6ZAAhUWSQPlxABglVA34qkA9L
8lwmP72ifpcCQNmPkCk55XCeWNZO9fr0x9vLiY9q/+frmSbE4jDe6nD+gLklL0mexwrZYE06EPiG
munzaO6ANSGALlh9Q3ZAAQT6VfegoNSGrALy0ceqn/g4BQJo+VrttQ3iheLw5d8GToF07dIgkmrB
8dRtHm8aDh+c8t0IjR6ebvsEAYB4C7RbYLvHXySZGmwpr2CUUJxPYMkFrQJdsvo60rXua0ooIWmh
DeKTJMYG4JgbV/KTfumtlalbKRcCGFnseEKRiAXgst2qMci7habcJtnV2YB/X1YPXd4L98F7b4AZ
Dx/FbHXIZWVhEPFbQgiK/UKDgakrWla7nz+D2Pf/DfW2qgIUVlcUc/BUxHQ06XpNCiyMi0g5ffUT
aAQLF2PGI7RDESJqRAERHEbaD97Mi65fMjgX2eIx2d29TZUf7EDNHOTdj3bYZTYAECkjpZp6v3D6
UfbRuHbF38z9aTcptBPlpMBHJsSjlayOsa724L8ubncGVb0OUt7LSPrPsKK9R2vjqqXnT+j1z31C
Dc84mpbOb4KzbUH3biZgQrt22C7Oz9PiFzhPABUUJK1uVkHSxomnp39r4vBUkHLoiqabcGCQ2ZQG
vFWKufO1juUqehuyC+Gl2YBQ34k7x9mMwZXqQ8IEcPA56+vJT7OaS50Gk9wzBmLdipYaYVuy2SOi
RrB3cluWIMTdbLLaMoVkNH/lwIgpgBCO3KisHGh0gB7FHM9Uqxk656rGE9sovxUsUS4eineiSfCO
xX5gwgP8DpopqbcRYztDqtBEa7wNZKDWeVi8bMlxHNhImf41yOkaG0qkaqLS3LmZCKgJHU0Zvrif
4WYmTJ1MUX72HtnUZfexiNprXT+YKRBokROcFlnIwOf/jR2/GhtgIOkFMyV5/wv4VRBdAuk09BlX
lPhC98hU3YZsXb2flbGubUR2z4MFSEWDd4j3chH7EOL2ybcS2zxYyAiA+4vGXIrwU+UG/x5eD/5k
dBKSY2huyX/Hhzeg1Gw97wYBclczxqPfEinxIt9BUMOJrZUhl6Bd0yKf4fv0aKQHhLYngbn+1QUF
HUMXNDvJQfYKK0FZbhbZi/Pwl1Ufw6+6QzA5OFje9Z/3i7kW0DNcvaltVcORZay5lgqsq0ceDaup
mrxpgF326EkokpQFDZ3V9fHCPXoYuwksJZk1PZIESK/RIRVYWPiHqzmfeUcLQwzSIqxIcqlC+Bk4
yTxoh4hlyvBgkKL9zIIe1rAKTB6e96cM5r54Ea/bM1lBo8d2g2s6px+kaJRdxP0J/wiihqjBq9O+
549e8JDhLIHNWkQYIESfybNXQz6Ekpj+p/EIfmZxVMvYLGAKxldLoeuJ+c7xcwcs0XtGSVgVHJx3
QDjMY/hvxpdBlFWOC0It40kCdF7yyWSM4auQYOeoqmiizFawmF62DImyYXYtbNuCuH8t34nVBI3x
PR1qB5VmHM99JLkYrM5Mw6j0BfeRPw2Oc+etXEQRCmhJC/YJpXun2/KVIGzYh7zreB0JtnahIhUZ
4dmTrSHuvfZZHRd2pjiyLX/e5es3F7IhQSXRyfEKpN5ilOAmQOs1ck0BQHrM40rE+PI/xVE6Cqrf
FThQo6fRkXnLD1JCRTywmVWrNjCaw0r4R/rZEGR/bJn9h29EC/XLUltM1NhtlsCJPJ3f5Tiuu41b
mTBXhD2cm5Zcna46z6vDCIo4vIJbAkz/o79ZtWrQ/QqMJJ+ZlWWcOwFzP9X8e2Mtl2ErWPL16M/q
ZYaLw8WlLqeUG21FEMgwYdK/CMhFagkA12C8jtGfXxY6bAZQ79vNBUsQ72nngBQPdiZ/Oh4sUMFU
NcTgnD7BRvnna1m4viDZBdieUipcFF1YOR/2TmoV1Cy/h5on04PK++Al34ewhPhe3K78rTa5xw7U
EZNLDHXkuxt8ZWmn0xtr7Pe06z0qd03jMpCZgR/sdVTlT7VKolCjndEt5GNOtxsv9vM+yPnZbF8n
1j6RjBjdmPtnKa0AAqUbrD0HK+1B0LI8aMacHVTZRO69bFmhCkWpzH06lslns4itpkTAYx5O+svx
h1pbN0cWbC6XDxEx92ejQHm86mp27WChFZm2Yy+iHw5df6RkC/eEFqhIsvhKsDg4JubrlaoEY7bw
0eyY+Yjnjy3oz26lni9xPtJArwLDHwfduJU6QvdKxceT5BUdLmkPupnuGBMjkWYbHKNa7ZkwSLg/
HqQjTEkIltocNd4PwBM1kMK6hsgpuU9jgcNEarldxBFlcI/M4YBcMEnpbF+PbrBnNA3AbJxBIXOd
zC0b5Bzof2pzUqIqBGjAMkt5Y/WOlyemAoZhVnSp2AzQRkTUG4bpBggV5olqBVOD/e+ERGUpOy05
hIlDsHNjMWs+AgSekskkNCVwokzQwLubjszQmWr28I7x+EaVnIASqFQMcXiw+G4IAFklajSEr2F6
TYaP2/3amTM3Fz2D++ckGAw4DUbl5/v15Wew56bYYSZoih/+H5iY5vrvmE0rs9+eqVkZbmLv+zQm
BHp05KNsv+bAbWGiIW5aBRsFCsk86eqNRcTDBwDIWhR9f5psC45WZtUt/fNEd5mLuCf95PiMl9yT
XxeyejRHDtlq3bab3jQC85NM5ZP5lGg6teueIEqcC4TXOPt5FRA+MkKLeKHCDjTL2+xfcumPMHcm
EX10he+ODq0OAKTUcz23Cwmvewz7KR7EqTWGEKokjNbFfe3Dlj7/eLgY85QcBv6XWrehJEDzQ0TG
ZZoghD30nlIatpOGQTpmsadXnkRuBz8DuZE+j+P4mnXQf7+wQAp4o1H5JyPRjWfpyIOIpx+l2UoL
hdNDsWEVEJduAQ/4oVUUB6C7WF3/NITC2fEL/cHHAvEJHRXH7jvr5xaTRLxHYUYMrIuU5QIyIADg
fcUqG8kM6ueizJapK0XTht4eMJScjaltBznDSV+DgjNeKkxCehShMUnnkLkn/k9NjdwegRA0V3o0
e2v6t9EB3RJdm/qZsuIN/ym8WmEtYJWHm17M1La56yZGAt10KzJ1Pt9qgHBt301n9Tiygh4+MgEd
G9MR27yxL3lKtz/YcS85/nl+hVHkfkdTFBVkFgvwmaR+63FE8cclihmb9sWL3srDeiDI6wCcjKBs
AQsAmUsgQQDUUpIXLrWpf2kY+lNVHzigo5gw5njV25Dzvb6dhUF0ySzOq39Psgq4yAeEhrYPFKjV
nD6x/cymZHzpFCuPLOphKmEKgGtfkOLz+mYZA95g0MVpSEfXx0+9BA7jaDwEjJslHghs6H0ZJ7dR
kEPyGTXERnVBUfHnamk9pjuAqjnHrMIPv6zEoyErfE82gvK8pbtqljkNk9MXoVVRcq5EdbG40JWi
c0du4s98DW8Kos16UdlRqXxX1LvZdV3j9Y/gE7tPBSGTCuoWAfgUhwkZ3UTvjgj1sGEW3KNBB1sl
9KtkLDB5rdUkU+7DsItf9p43SMLBb0npgKX8EQU5ugQhL+FRmaPkEiH/Jv6j5SLwHvxGEhRbdeQs
DuXF//dw11sTCzmlm6Whi1nPrWp93cPU6+v0pkmBUdIc+iKyTokt2leNXxTPDbBjeIw3PKvFighl
oCfRKHWIo26YHrc8PtaiGyXlk/kQ4aqwQCk5uBHeVxDp0j6e/lL/naLtkUexMpPlP5cLLyy4YeyA
8x3e/s7ctJ/cF37A7YT/JMGniB8unUPVnq1iBNc6Jy1FpXzKQNB9CyI/1zHsHWijxU3TYEuBzJuH
Gjocu8uttgKBWt4mQWul2TvHeB5BJNLMXtXXwj862jP75HuMGYDy32nyh8gnJ/rjV6tGnfv00akH
/iy62Y22Ue2+wi9z18VcPgVunihN1ZJB8cJOT0p10pZ/TazCJQ0L2+wb5XSRzLqGcps0I7qQWPEo
TTq6XK8W/shsjKTjwJudj7e9IiL5iauzTcUamxDMSF8/H9/Pf5KetJtAhuS09YNC3dAcev3YzAXx
AfpYXzWeMtSdCHzersjZyhNE1ZJUHeKwPJ1ltloszu2rZhZathRnbNZM4SKpqv360LGEEQ5finPw
CIKnl2Y1d8RzVf+SGjodmP5DIUOfMJvZYyrzuFCq8JCsZW+F9YqmR1rNtWWXH5Pc8mbbXJNzYA5V
Mo+P/6i6Cex380nHDUt5ojZK0hj4KKzahYSZIcTKejrUv7A91NwRNXo1+YS3OP1RrfiXSjnyd6ye
xibLuQM7Isg/oiwHcDUV+F87PwzgThwH/jEYOBzqP7iAZdhaAoz+KFPGYclDCIm88x5UtAYncQ9f
0Lv3jAphfQ6hwRouqQNjrTMj/l0zyYq9zujUMVZ2X5oiq5owKHWyXZ4lqEypbOETJkkEGUqMOGMZ
ThEViS5+VwyOH+XB9ziTjQGL43pFv/F72UuI76RRn6HuwxrzmluXSLOZcxhDiANxKXxYEaZr4cxX
U4keh+Wz790r4NinHascLpPbIItEUzxt50zo+kxWlnUWq4qCea6PQ9IqNWHuBmTE/T2PdYUPkUrY
cATuK78XT+mSi0o9CAuO5sCefwArXpIV601u8gsJAu8g3RWlzNIKRDn03+VY7J2+bNpGkARjo9Tj
pP5Vxz9iNfib/tgFo/z74rkOWKaJYLokwLsB5zsWKO7uwXGcV6MKrG72xNUxOXrgyI6mpwt1seWR
GQLTqZxwo84BlwYkHns6XzFSD8DtIioUmc06u9C98UYVxzDcWRq1h+I3PdWT8JzCHG1i3t4uhQQH
X+ZDNLNLFMxls82AgBto0x2SDiN6kU3SpkI1SkOCENJUCkJdHb541Srb4rhqfC07vaSaefuqiE+y
D61pOrS0rwoVO6hRgUr1Al8B1oDEut3sddKpEgI74qLJUoZaFDSwr7wUNut1hfXLIE86lI35nJEz
9fAHOR/R7hTul8bO+RfgA6vZDWSJERoiRVn0y+grcltL3P8pZFDfvCvA3kUrWo+N3X4MWgk9Bw7s
TBEpXqnoIxfaD1064wkwr/vChBrxaz/Czw/HNQUCHxbC5gQxLgfbOZ3K7u372HcO8nNXMZaNRf/y
QOcw7K/bHqBewoGTjjeL4/g5h3tCRvgYVP2165JyYL5BPI+H9Jae2GX14h4dPmDGJ5EZSa1Dp3Xu
xqFh2Cyyq+8UZqpyaKCrXo484ROzyOuB/2AtYMk+IHLtjVeJjELJ2w0z9vM328fRcFrY6CqcLLKF
TIlVkHVjo2JuJJ5Wal9q/yvfPYF5E8ij+ZPQeX/qax1gM919EXa/gyQE1mZDUoD6zKaFM3n9vyWX
gCBx0sn9aHX4WfilQez8FI7VNruERwgnUblbkdI8D3/xNqByBUDV9/KRWvdDZJKXH8K9OGIXhDxm
Xc9o98ltDRVcIsZSPxIYqfpCOSV5i6vKo7IiY2i66f4ZbdrxLkk3kAWtoha+K64C626jZlkNujwZ
Dncah/0468X6EBINfjxSMuloIfFwRrtLDfqZpPhlkZYWBnR0kvu0iFuZVUhRAAfuHj+N32FaZZJo
CSTBvS+z8olprE6NYJMpuPt8F4dEivO8OhxCOMVFGgH8DHIt+NUkFeLUrSqndT4Lluj5crFd24G8
SiqLKivXCcCH4vaF6c2v0pwsSyVRr4DBiWlaP0rgAuxXCV6Vr4TDkPpEmBJKLuc03ZGd8KMmumFQ
XEja8AwTnUlLbCgEwVj/x75EBRcZC0gAeCgLEsy6tbMJBTGZjOwmw1XYsC6dtSLiFxuHVmrHnUdc
LwGF5MxpznPfIjbDrkQIf7A6evuwd3YUKffKg0OBnA1wrLF/sariPgwGk9u7L8yUV5QkUy6f2Lmo
LtfT/vnQnSuaRfDc+8z61MLhX8/5Fy2RHMIEKNB+zmZt8zdNshc1BMEoRYHrYN4+L4Xr6b2WjYSp
ga8I0RZau0lmzhtcahRfP57R0GchXxqANjOYyLi4Xjsw36i5QnSTXSsKsRN69qCYl/kEmqcWMw4Q
EJO/Fj02UZcM0I3lfjzfI40hc9tGosVu3zdOJ+fmoZP4zQgNrZzETwMqpiJwfkpFdeCrLT/PVcP3
Deh6xEsPVyhiyWbpRt+tr1p9jfsCylhm485TiQbols1iCDK3pUh2tbjvpLq56mOV+xOrg7ZwC+zj
D+Loo0Orcu7CZQztfIq4WJ32h5h0Ag0FMeboaJovM1FyFdch+0seDJZCafx0zON0SvQV7XwtnyoL
0NsbkckpJs71DHuAlAxFE1QY4UVrfZe5/jGJWhLzrqm2/M+hVIIQI6lj578j/Ll8WB7kqkQzW8XZ
XOGo/eNXW2l+eRQ1wjxXFBwmoo9kZQZilpS9evgr3pdBbHvomnLxn7yhmtnZYlCOkPOuTHTJ7ZWg
p1eGYEU7EYRcjJY9tu5faMV8RnUwujRRAnRJKguORU5oUV3W5/GQOn6FDNLz4Nag+/pyq87Y5W5G
+3yxYSpsHrQs+HK9idUfJaEyHFzmreXGx8/13WKI/mjfGg75Nzhof8RgMPhFw2fOT00QSdjMqrys
YSCewKH3S714cFi8pV0WBMi4Oz78mnBn1TXn9npzfeiknH4o5B/zY8BMvd1VAS7z/grnMIG7PtRI
ItlugAyeh7WfhcxCe1xnf6aRq9Hw2T+Lu11Vs92WsTqXefNIAgg8eI4ypBaToYEzknt8+4mOUD4E
cc9kvXzLTffHgN6NswQ/uD+3K+rR4kuE0nBiWXn8X1NCpo9DQHp7kbmznGIFJYkoTkmpNivRkVY2
Wr10t03exNlWzl8QKTw7xbNPtcbrKNT/n3X1Z+C644MhTKUn4b97f1Z6nlq+ou3qp9Z+BbmRuCIf
guky7Hdljm78EllzgV9bX4oTR1KJKvvNm94j19N8gzcQpd6zkYfxYz2W6gBmS9PRy9E7X2/hY6Du
Nqdy0UT935/L1QOif8sXSZRSokCvgEBJ0ii1QGG3misUPd3GA8/VrbKNu0xXY3GBgAf519bxv+hm
E+g345u5fjQdMlDz+vzQQZWXvntRva01po+po0GlVDu8BdqlG/DL44OdbIUSizTszw+VCAQOj197
nuGdKnVpVKO4i4ReiP6FQXg/ty6yvXuMOJmYO2XeyH1+1zEM/TZ2Xz20eTHJCKFtveSuDuZR3jPy
BpJXrK1k9yQv/Qc/n5Ev0i/OYJAGThMMsxgpGTBMBFhRSKJN9uZDFmktznTK9msAW1JZY+oHeYfB
B9q+kcSRHbm/mQD29U8Ubg/M8JwW0YrAuN0AEBjh8J15hiGsNpPaXvagZDHKqbemNu+IDBh8k0fk
k2p7Fsi7WBmAQRobzTAqA9qTA2Bhp8eaR6TeJpp4V/6nPQs5z6jwFVkn6UYvL9rgii3tsjer/nkv
+mWb3NBInWGhQw3bsxTnfcnLh2RP6M6wVqzG+f1AVdQgee016ZULfF13XflPEG6R2GFcJD6vm+u+
awoXAe4bCAvrNo9rcdhXjWleElA2wEFSeJpJFVU2/19yAowOUh3VYiLFaiQpnfB/CwP8LUPSiXm6
tGxSPI+sNYjzcMrOlBwZ3GDPhN4RLkbJIkvDn7h9+8FI3Y7iiSqzlYOS9nre12R1TIH1ZW0RclFp
CvOxtsXgseV+G5a1SIvf7nkPj5xL0Voxb8egxJBGRUpGJvao1090bgm/bXdCC7RdEN/v/CtZWG8k
o5f639+yWFujaXqkGAIG0BLpAXWXBD6fP+vxW7DtvaAOjm8Eo0+GZEFpG5GQCQgxC6Pcty81lb+3
TuL6w9rDN5Bs/8XFIczymBFx2/o8COCHRb7m5HTikpbrNreGE3Mqt4obVBBPSyLbp/em5ETCUSUG
xp66avLNqVNBL3Cmxm+kuZqRxymTWEYaPMZytP0GXOVFcbELMuWCcTlu6EZEAMj0GI0JUaxBUEej
KVArw0fyMFTZ5ZLs5WQIHLOoBZQvSGPGuAbMRmm713qJZAd5+MB4sQYnsCX97Mdj0pM35eFE+eCP
swh/YUrL/BXAHGCFrjUM1TiDKTDsy6Mkm4jQiGkAmHqhAVhXmGTsNth1CCzD7qcSfCgHXTHKdWKc
0ew2ZUCFXe1P6lZsk+WamUv6b9a9fuiEERzPpMlkKnyFUJNacoVPB4v36rq/v3gU22AIN0m/w34s
zI8BLIPtmOXGhZYKhqOcSbKajeBwAQdUhkfNCb7Q1kHjasmJy3pvfPseofzFCNtED3sOzPUvOfc8
rTwjp1fKbIRMvG8ypd5pCpSQWARk9FS9suPZEKJ8HFOVA9YJwBHgxnQbMDhd+BmMaCuQzcAVtW88
ITmODWC3Dv4lh/02b7ltDSG9lAP5s1dYJNKqBow+MsCnihKOQk7kWmSn9IekubuhxOf2hn63OAUN
xWAuW5lllQAyflrRHB/G+kDYapg2d0GeMoX9S0pIVxecPW32HT9Wax2azH4/jla/ji7FAbHXDTiB
eqs/9bPGVsP79VmJjez/A1kvbqZg4TapM89XhTpR6IXqm0US0GsT+AS19DnAX0NgRljMXdWvWDMF
c5YR03Zt5s8nHc247zEVuUf8LWn07rvz5pAUv/UMyKTZKpGAdW/qUBNjp0S3JCsYbofVCtu6wbzJ
vwGbRgmV5urqD0l/2gPMFrDE8JU9O72hp1FzLAo9A4Sr8fd/l+ehsKt8W0NFPgTASourcL8Y11jF
3/6UYrRs27IhquTzDv7pn1eRpeJFdH6rSMVuzOE6nikzWWHIp6goejLBTfTQM/S9b9qtQxEGVpzc
61fBm9h234awW6SjcjxI5FMN8Lb9FqZqrbWq7Yaju3oXhluSjvQ/p6zd/8osNZ6vjGfY7RBEtWaV
ue1kIYb46eHuCm7KrlRouPnb2n+4Mid29Rsmg6zQfu+3ZyJSs0/W23babGOgICmYwhoB3SNjkOVp
GcYseCJWv9/Utfn58xRV+l//6SjDFyH1bj/N/qrS/xDzEgLJYbquC+I36iyteSJMXNOWUdePbdvf
DVMo0/u2SQNox/fqtxwUJw/zfDUyaOjf+RpsuwURL7lhKihKgBaHngWMYrzjFwwoKq0RyIFuGU8o
quHfvjPYkvMvLLVZScxHvlPU9hOiSjjXjzsAjlCiVoom6Bj+cWW46ULzKtWDQd6EIYftap9GZSsy
zsDbjYDZ4WSpopF0vNsaaEZlyB3f0mZr5nxmXaaoWb0rarI1jC+/F+JF+KQAKow1UUUD5PN9NMlR
XK/8ArylX7W/31PsuZrmQvdfsMVIkh09BdD5cMMEJXCHgDgKk5RhLmflIoyhCv+En7AhPyHixMzX
ezJZcX+GeaBOK/eZQ9Rv1EzaDaBEqy0GetOCt8HBj7ne/3XpXRDbMCfErBMCgQNQCfYkJ//fPW2a
SDIRE61N3LTlVA4QB7RBV+8edx8OaQOpvCBhLNGkGJIj0uYPAKGoFz8xII/lZiAdGr0ieU4VUssN
d4hJpECsZOyT1iww6tVBOpyGtEtlPAr+mgI5lYGUAyh5i264BqXuz+ADy+gN1YIAIWEBK3IW3AK0
iHMMCjsfWoSZ41q3BBX3M3j7cLXSCaIWwNK+3hLlHfZBBAhKoffcYdkOoY1SXria2BjpISRhLC7H
Vj2PPWKFH3GrXp5jAnIHqkghwu1CrvAAPV5xHyNU8yjDAxcJpOvQgBrZpmxqLYsgtsV/v7MBll04
TcjIZSmHIY/XznPA3cOgToNXDj+qY9oqFb7gY0YRb4XFlLyijDN5J2KnCz1U47Vmc4zbtbHyAOW3
5i1gwsXKhrn8icr6PpO2ckWS0y/+zg+ilr0/NDL0quTdY6OuSUBASvkZkjdseaAankzoLTRL6Q+M
Hq4i5SeO6ZevoI0Qy/wYJOGB48zD6uKDCCcRA8qhu/5+ty5wgS/OYMbGq4BJV2V2HZSpPBSgSq2r
Uz9WQAa9Vv+5u5G+qHt7Utv5uTarvFJasCRggXSZEEeEdNsnN/TW5wMVqQ3fsyCs/gDnmfhfctL7
x/lq5D2RebjtHDH5OL2U4y+MySfxqYHgxqlAIPfE2hr+jR1BNmyeqbJF909tHSXzW3EgDsTUxise
VubERlSYb9V0N0tKVp2biupObDraUvNclcmRmEytCOHH4GskRZtUjhv+3Ff7fQgpuGY/ssLGKOO5
VorL6BI+chKol2GER2PYAZNLPkuQWt2hHRlaa0ni7C++YpoziW+oAT96slMH5pMEuDe28kkgO4mk
h9S2bIkWfyybuIMnL6FoiLYVOsSNhW4WH7X+e3ga1lcwHy5L2tRk8YQKiwrLXwZDRCpK4wtX7/XH
iXG/4s7kJcA++B23+H+xJ6jCIV68+fPRq3G+QkqnKsI/wXXlyKrNlsl2lLtyzUgMFwvzZqzZ2ag3
sYozu15YNGMrvW6dT77/mAznbNKim8Ry/rv756tNeTi8xxQW/M8smglxCPVUp/ElFBaIcTgiUIjv
Hq+vlTij4ocUgLYoGD23LDjaOtrNa+JkvXk7/VKrLtJfQ/bmEOs8X4zJzbIcSYP7ER4M9Tmr0nAn
o82/NDRS+DHzXB+5OJ0ibPwoeLnWDk2BPFCSV1jtnRrPSmDRbZ5mKafDa0RUK4Ur4sBHmp37HsqB
+w5bL3IioUEpKC/EHcM5hsYyoieQk0lSBqpaIVkqcHuuNDJS291Ie0nWWkailcgZDNcq8nD235XI
aOZaP5u+YGGMQGR5oC6VVkbNF7EAnhOOvsOGBmkeFeT3y+AS4lMyUetZ9p9m/LKHkMkQj74uRyDX
/Ekcp2BMhSXLuR8t7YfV0O3K13/cojUm+qhxgAzf4YFUg1mIELveM5oZq3nIaa8q0K/369oGqqt2
FJGCU6swFgkmdbNt2770c2QjTi9A4mM3X4Kf7EFBR+r7mDLVvJ0AwsoPTjen4d+Oz1Q2bFCV1UHE
WhpEy0xjD55bm21E5pX1PT2IW1Zt2KURaVpiGwKVCrFGm+V7Axo6MiFpsbPog33fbXCUc55Y+on8
g0qc+6UqTWIYKwX71Ak9Yirs4VTT3O0Ks7Iic9utDYAElfUQHe//eO9frsPL8u6Wv+GFloweqAR/
CAdgxfE8FKAtj1Ce0mBTY2SiVP/24n5h1faE49dJJ9HBkzu6kM2o8ppmbYbO//39ujFZWiUrC6iJ
w4Y2OU9FAuJRkdlBDZnWczhL3gGhJlio+q+2SZRol1ni4mO0Do4ys6jXeBzvvAISw4y6BOu76l+d
b3vcZgq4a5C/k8/var0qwl7ig6O+sW+0Y5U8qn84NZha3tEey/AJLUXeecvMP0ZRDbySK5DvlirU
/OT+qzq0905sLzN3b/mo5i4N569qpqkc5/RpU9tyXiV03m5KP0HMmfGs2kHVlNh1P913oWmPRTwz
TF//NV0t5gjM+Yj7FSx1mdTyZ0TKEQF1IjqNxtGxPX2fmYAv9aP5Yrm35zZVLXwQ7XmFE4qY7In9
pd8XenypqHVzTymJ8ocCVtd207/KdRNqJHdRWrOkLwqb70Gry6sitQ7mYexCE4tVnsDvNn6dvEsA
6zY1AzmV9s/rQBUHya4tBIfMvUp1kU/sSZLzSL8uLtpPTBkt7oUd3sMwLfdowPJxbQL2cwN4+5Jb
YWoamnpH7LonOcEcorRY77ATbhuoR7LYlMp5XbvmsHFkLkfFyXgHoC24aBkvUkwAgYQSWNcbS0b6
aqYUlz2TZseYHWNc8tDWKAzHfTEZZ6xxGopOovU8/0zcvxDgyb8CIj6xv9UWlkvZZ40GjZfoLTQb
lZz6coJZVM9DKNEOJNodSIbAhXIDLMMPbWeYJoiJPeSH5IyzfagLT2fME0PrH8SrFIHuwFb4q86S
UUA/Mxz4whNlBY8TOYffk702CzB2YA2zs0cA1j6MVty9Ji7pydbUnODnIxfsStjUIIlGeAq2OaNN
3MExruj2eVHJdVdcjuklL0LuW67ox8VmbEuRGnGDr1ImfINvT36wMZOfBNIVqF/M/qVBcCIKd9Sz
lguHd1SO9fi1cyJRtsjTEz1km1N8WBLB2rUdZh6QPDnfGvDZEUtHg/HyUAmGg6Qcervjjeq5Arvh
AoMj/I7f4QTUsmmfIWbbEW0q3idIDybh6qeiU1kAetpCqG6uH46CYVSH4XbZe4uEZVYAqFPnp+X3
s3XFSCO9B3pirBsFqDij7f4N4Yv7o1VZj8meIdBeUxTCHYynMccqDJkhhLz5Vu6MMr25iYiepj4p
6a0z0BWEaLX0c3Rc/dqYuigaQCE1b85jtASwUYGJVpdInTXkYVYCm3wWV1pjdaMSiAAfg8lDtNPO
t13NYgzL9n+9D5FXVbfT+i3kMSeTOQoeRiwxc1dcqjdu44dN9n77lvFC4vWlLaHQRn0J00CRIvfR
t2zU1mvgTImSxh00/5i5spcNu+zPJ5M7OhuxJh9+/cqTFuaekoJQGAG8ZLfYNpfnHPSLVYNGSw67
JPU47Qww3uOKAsVv7C7/rkSRW+Nkpm2FAf1aXEOrPpFHNLscxhG0jBu4kHU9JHzFjkbRdtJEWtp2
3dgmY18oNBS7ssxf0zEscq5RB/rVcbaEliYWmVjzhzjEwo//h/VuateEOlsEmhPiG9C5PjVUeGJF
KyVW2qRH4zMAZLxq3r9H+33D20UIT59hol/YpJU/YaTTswTZh2+Uf3kSKBQBXyW4TsJzGgl4mFhG
MHOMa5mhzXiknFM9keQv4x1Dle+0bFvky4fiwew3uKLBfSG2tIxuMU6BlgzqpnXXSsKVekO5/81j
GtPaMMpRlkWRrQBPSxuAi7nOcr/pVUW3rQRU3oav4FpBXkfKa0ATrEE8J3gY27ZZQ0aTAepbRwuM
V+Lj67hfkjXIRgGBt5mERBQxPN81YykGhGfVr8tSh1MBHuzYs0I5VYThaClX74pre4nIyVmyG5FQ
QSHONW6o+5SeXJx6Tqqb8hUThK3S9/r82dMmic/RbUfd8goBILombBceKHh0QgilRq2GSpyAN4Iy
pQBgzu9YbT57MUtmi8g+yo7BRV+vhlb/JhbfKheGzDUROeEDF7MN52ed6RKXKT5x8MgWjyzj1pQ3
YF8r1YD+YPAYmLnxT+h8SLjXtaglvdxJOGn9iQAo2gsf9fw9RM8mYxtmvXP4/Ul6H+qjcjSbDUsk
Dyf9MaW867Tzdt+kkFhtgaLvpEoB/ov3ckPJu8TyVC866/gi2olUqsryb6nrxbcFn2+OUllCfO0+
bByGHGrtXtA5YLQkT4yqOGP/ZnBBLoiCE2MhXtaPSgZaTPZ+wCdTt9h57U5FRIFar4gR5h8ViH+z
sf5s8frkyvLouTMyE8clU6u3+/uw1dzcsb07I6o1kQeAe+edMixen1xLrDPme0vC2C/ZtDBIh86k
4I7TIX/SiMz182ompeFwxzxGdcgUmpuCUar29kXFXC+2EsNSBECSYtCSXG+ZlymrrmDo+vhT1DgV
esFR502boPzbGKDPyLz/eGgDCr13RPL7KKLHf01OzbSsMyMhw6nk/pOEZ99YzKsM8kpBi1bB4H+C
DT7ZSoloK+UVg29GQG4/XoikStuLrhQ4vwcHV1UT76eEs12ZSUrvTy5s1k7iLODHNDTc33cUno79
UTnC2GdPR8kMEudDg/mVupqaaoJiWR8gcmLSNEdEGAsaNQ7n1n97vCnCpem/JRBJ0Q3Rl1RglNCp
gLBYvQP5xl5+sC5CW5aPF/RzHATMNs1xBgjmI+mmL5LjIDFu1HdGIaxD3BagKozKOWoZuMfh+JBr
AJWtpsEIS7feVAIluPkINTV2aFo37UuP4cadMm+mCoMZu9Gi7dz9PM9Wqib+wgWAViegylh+AIkX
KFAf/Swqm6y+jpo73qjOH713hDZPtlKtpQxVll5169NdgLw6HxfbxJqIGCbdMtbH+oSLR6gpWNce
J+qDEBhXkd6DVE1rLFzkLQ28OLQ+ViK4bBylrkt6bq3A/sihRCxAyyEeg6K7FjPzK/SCOswsmNm2
5t7HaW+DEXY8onDWPnARAsTaV7hplIEOHJCjDc4tY8SzngKCUhLl+Id/r+LcoGZ/a5v4C9oq1p6e
14gESoZhKNFsWtI3r1DJJ5ZPZr1qcDadiDR0i5+Vetetw9X5dgvkZC+KdB9xLP32D5BoSqx/UxCc
ArJm41TbYqcxir0CYXK9tb/jsQQZZgOEtg2jHHw0hgoR7Po1zk/H8+KXfsanpVEf6LpMLrZ9I368
oUro3sTJFlm48WJCOz+ORCJMAB53hMzEDyOsNhec4Tn1jO2g2GIh3YWZCCl2HRqpGLrSR1oF0ZxD
E8nLnZ/htoBFvVYigWFqRzAUFm6sQjPhHlnBk3O/QBjv5SZr2vSWzAHF9PbGMnqdPDInMz43C0G2
1sKPrOKi/f/t7aytyTpnajJjIKx/nefqZCuJxW6uQUaAp+Y4Ts5VUZAJHi85gIPa6j4KqKhch7uQ
UWYYrjUr6sfwezSwajP/RrUkdDJwTHtcOhg06iMneuIZasWnYvtPgyCpl0eQEmZJCd4tMY9+tSbP
zXsYiGTXrEgZT9GAVbtN/0F/Zv2U4Z3YdDv2LhkQrNrdaNq1AwWOTWlevLg69oV9uoOVx26p3jip
RJmJuZIET//Dm1FTEB4XHQ2wS9zElRZeafZbOFol9nl/dSQTBNJOHQ08LpaatWdtf8tk2ViGAFqk
kSF0jTuIOkpG2qUS1Fo1ZH2J8CRv0sj8/mf3MxUR594UJ9au1jTVxMfxQv1PLiZsx55sTCS8F5xN
XKblY+iaLTMBt2B9d738JHCzGjP1N7L9Lj6Ppd2iiLeOe9psOTc9XphjJMdrL8wUuETmQvcbkfYW
GwSrIiuQS6uk1S4nnLlMf2NYcg2VO0QJEz4NZ4Md/qbexExfMfWNUBnGQhi2UfBvFk1QXuUInYY/
rPqlZtcX4NpS4YMCNZgb/DZX3Pe0xM24F7p8pxw4QJGPocifLce5dDDyl538nQ8tTLGoFkKZTY2e
YD3PC6/uCmx1kTMoqwsbXBKhBowXWlqRqdFT6a5Lwik64+1WHiy6AKDj2XCGIaLCi8fJykDFsBKM
YTqOUd51NF3wpLhAvql9WS4ywHri2E0tcbCUtzVNtTfFZ+Hcn+0Xch073YAX1sV9mhzamuINCxAl
OK3un0k7wAYUGJqZ9ikJY8Up4fiKLQuXTuJya7f5HeHbrb+1by4lSeCOcXUY/eYxfM3xB5rU9e78
0RB4uMZ/ke55apacuHRp/EVrrYAbAB/Ix3aZeWiRGOSUykaoMCUTOkVDuV77D4p1Y68H638lRlxb
YjuLRKzujXsl8ksRINSvPqQAcldMeNCG4f6FRiaCwDiFxMkKfjDGGSDVjZWeuhGs76npCfBCGtLP
1zfB6irKMAxtI4nNSBmAxwRUC+n/STDES4XdIQL4ejDACcN+XFLE2ydA3/rGjI7VAwppKb/i7170
vzUj+ptTDzW+55wIkK173W+JQBQGSpWbX9EUg0tLwn2HHxJhsGQFjOzTl8BE/CpM3yG1eKnd1seA
Dph/H98gN0uYn3/ya3dNrHEwnn1y3k4DvQUqxdNQwELD037ZrwgTjB6Xx/IJQRdD0mVQN4pZrJEJ
yBp9l3KTFUfOUhb7k3m1nAq77iochyBv4m8kwABEGTkYLrsrJCFVS7VikBwna4awD9Kf5xwYDd9C
kClEybvNoxFkrHSuWhMLCU+3h3G65LwevJggn4iFeMPGZify91eziVwShayPVNTq3uiKqpl3UCh3
mbi35lw3tqfE6ndhEShRYPRB0k/1DQa94665ATWzvFwcSY/yT5YOgypufh13W2rw0z/4ynSzQE6N
jZvlYe269zEeScgk3ozR0q+UxNnmu+xpCbdM5uWphcPlXunu1uA32TSoNPJTABMH1LCw3Jc+hPBW
PdgybK2uu0MVROs/w9IX/Z08SGuoCuDabDHpUnc2eH0Caq6IO5hF6KV8BjnFs5cRcRm39Of7srlf
RV3BJLrkWaMGDxPJxPPHFLsMRGWCnFC5a8/CK904Us9Qicpn1gDMXEXhZag8qNMmLZhQdzUUTzgV
8zXmm0VP30MLkjTkuUJmXInIusuc0+MfwdVmmC8lRx4C6jSO6VgdWbj6Im0JwX/wm6uzEtdDJoWG
Qtk2bFVSv6sAo6DoaoScHSSjf2E5dnmRdIpezZHXodY5dZGwmnMyygc7d+XduWv2DC8qfKRD/ifm
0xW14suqthdiaICsqQhJnQmr1NwzchDDoi3/Weco9zj1QuLpX+hdeRFehXb26F/EPn/SP79CJW9v
B+I58ylj8ja6ZZ9KXoUoy2EqbuCv9WQ33LvnHWRto2VHf20OBEllYapnmSPZ4GQvEM4rSUJRXFoX
he3JUFmaQikgZvBaYhdvzLuatSKv2e5BObiKEmv8fxfL5skadXv9hzzMDurSm9rgU0pZ+1hQpeZY
fbfNccbfqQBuQVzaACcKjyTqcPquNBCF+Sct0wSF7opc3n2dYLnCnQJBkCrWGF/87rGQmSKiIviC
rSPALLhwz40wpT6gQRVzBXylPISyB05APR2DGwwSYnv0gs4lus+efpwTbeax2kOvQvWoNfnLqWWA
AxxXhpN/hg6cybuun+LGFfeVNKHD9yzZUrf8EJRlucUrtj6TCjxMY82bSVSe/zdOj5Z4xOu2HGhK
ChItTmlUudXD9HqrYpLfJ3ZB6cQ4rpJcl21smwDZirzNyt/scwS5IVV+7Dvj+dQ9ifM07niw0PPz
/IxQKGY7ojH5lewqC335jTUhK+N3TvULNQ+Dr2oJGv5HMCvpn4f5FKft33mmeiEGDfKMdjro3JtA
QKAm9kgKgn4SZy1ZZacvHsQ787K3PlJiA2zsvNRiJqUe/5GewIsFEI+SLhsJTf2dndmv91KgkQF6
620uR8Iu0m2lPeueYCKmddIpTwnKDU5+Qcu8W3B035+QWdq04hgeO7XjS/aH12HySLDnYGkMCzVk
L4a2z/VNNv7LRFmw4Fhw5DePDBbQNNn7ljcGiLtSGs8nnux9/8ZZhCQci3+3hwh1TBA1K/0l/1dA
KD8xM1KetHa9oMuLSDqiqfrLH4nKw9acZmAi9vJyYfjadCIIFP9rWEv1hbVncZ0uMMkzN3c6jd8n
PsTeH1mCnnDqNt8aAQqwkAv6v4ISbgxu5joJ6DpW+F0o9kscsF4jB5o+ZjW1MZoWCXXB0oOen9Oz
zTxIH2lUGDkV//nSOcgwrb/m7lLN06qmPJXEArO7vXnoH2xGtDE0eRvKg6vqe3m8x0wuFFSRSqeY
EHdVB9SSRO2hYiOD2T3yv9U+ZJeglXzyvZzL6Sg44EbgZjrzs2fUmXd2PE4knXXnN3z36655/9eY
EcVydT9Q/BRhuI0ox3KDfToEsWx5OMPrUALXqpmyXf4ymwG9dNqXgTU74ttx6Gf8QiSTq4xdwBKx
M3c0t2Jh52HVPB0jIOLVoEyHXQeebtQist3dlxqz0JrFFWyCmRMGJvAT9hJekuP62AyTfyPXDBxc
b6pqkBLegoDOyAuncGYvxpRg99G8PTuk9pkIeNtq9ocF5fNhQcjFPeXpwWHodBkGKOK8r1hg5k6U
mdvLWvSDUHeTENGAL3WWQ0dpMIj0TRhx+Z/9IfnSqVxtUr2lPM0JJbG4jr5OfaFYIrZ0lgV6eI5t
ZTedl4NBuiCD17K+70sfB4vJWyTQOq52zC17Bl57WaO+CXuee+Hp497Mds6MY9QP7ZLZvmGjRaC1
c5hW4Edxwz8UwaUm4bO4hOTt8HkE8otDImlSD8Lcr1D8lpE/6TzkpZYdFXyAi8NxSx2xNWC/ILTd
pAlwcAX4rljFCKjS5T+plFQkL0UIT3DFujEh44dqxwF08qFioStupS/nYBiXvtKxoRqn1cl2faRi
+WX9RIiWO5QCZIFqV/tW3PHKRYLwOtIdG3rPlZ2X5E8tUawKAlKq/mtUZ1Jic5ZL3XfJRcGBVRp/
N5DeaAn1kTTGZcDcePxHO1jlzeM3IsVsh+KhkedZMq/Jc3z1hLG5zovkAI83r6mbjSrdJtiGX871
89shY/6C8d90GvWkmIEnV9Hrd4mbLipEh7NXttNKoXEdgajBweQWp1jknsyJ0dFsyWRHjwfmJCT3
2mRUY9lkMpYuF+TBOpkmZBoRY4h0UeAAcOiP7wAE3VgjGKi9HBu7vFjjI5npIiZ2GbduqPyKMOQL
9ttE8Lal8ndqPFNFeQVry3Ztu1Ud3qi+bARKyygsQycr3u7wiP9X49/bA5T4ayrDIRaUMUZRCyiM
m0CPSzD9ge4YBIqoM2tRusQzxuLRERDivyjVq6M1kjsrxIv7/q3Un2tV7FxUp9WlS+Ck9Xght9q+
xFi3TvO59TU//8A3Qt7ADGFfSIy6GEqr8y52c9xWR+Ko/opG4vHMY9/1tO6mEPzY8mfF9fr0+PE0
HXk24otodDUEciRdXvVhJXM7dw2DYQRMZ8usVuZ/1+0mr/C9o4VGLU1dxHfApSGrF20vUv8/mWH0
XNt++aE0VynE+2eMciQHKl/Ec7/u8i9V2sUwObcHlflKFV8dwuD731pOOBvx4OdT5PfBWUz0CWL8
Tfm1C1ZAj2/l+n/PQOzNBaEmOWRatF0it3F6dEfa1e6zd5Id6gddV2IXiVGb1TpFPfTJvtoIOBAS
ZNjl3mgvzRNTV3OKMzj3PyPlFCtFGZbSpZi2yrkyZbWn2nE+1YvDTM/UNPjF8cm17O+jkZdKILMs
edhB76q0xGTG/5m7slg1TtGcdHgvJwBRjkMR5FOn6MeX90GB2PITz8By8i9kHOfZhFfVrRX9jjGS
YeKr/6+MJ7Mge9D1d3mtgFmlNB5BaGRMsXV+Fn5JsUh7nFsDMtYsA0xhAOMwzEeM7BIiWSAzDRS1
0Vpd2GcI3yZ0GMX0ccEAp/E4CkmeoiSTKqTLNVE6w5BTuKNWMySpucpal3LfWKjN7cDIQ8qlyOwS
DJd/HgkhM/vx1wszUIpVBu0OrYJgNYZ5qMvAK5lrwpf/G4LgLoyibt8tJBTDNQAVsqXl6XLk4lXT
NPxDPFtS7T7kzY/ibtfg9b+1XFY8xgPNmt2zHViAL15INuUK3UX1c8wZetI8F9y58XgxD4BHDxJW
YeVOdILSuwYtR2ZhQFBq6w7oZzXTSNCRGkHFuS1HruwtbSP/+Z5QCvVEZh9ziSSW0jfcoYS/l7hm
UEmFpY91S27bbw01pfr9jVce4dglRjxgILEa2Ewte96vnPBd9I4Ch/2++5fDyooFiaPn9nIZ4aO5
35cw8VNXVRSLkhFItbIPGogFHRSGdP1XMJcrN60gKoVQYR4l1Xw/JNgAbE1COMqr+RdnXdP7vDNi
QGRd0hDpyaoX/qbi97bXTCizA6HodumIqxGDm9kH0ZRLS1N0XKkmRm0lkPAyrD4ic3PJs5FpFxkS
bYH2CwbCzsNN+NaDZzf8SvEzWp/+d3k31Pyyr15myDftVEUYiPKzebDCoDq6cwKKGSAV2RQVW2ru
B4jRzoJVhxDu57OJBJFs3da5OlBEYVUMvdD6OFu0xt5pKwIMyJbVPyfJlBhQKNEGVFzyGXggT0DI
QvzDJ6H6udtf02HXAqvdND5J9N0yR1euIchaXptsJjsCYGrpM6vtDKJoG/sNGDHdHpa06aZM5bqa
5KFohJ32HoZCR+63z4Ls7mbc9KbJp0NaY1oT/7cbgxH2HzvPJtfNJvLU6PmMBV8GM/TAWJRZ2t3n
iPEEr+Etf31drg7ouwdT/HML19LGgomkN6Oib6CzxSHpmafDJCh6LvisSCnNlqJqpRkoClf+905r
96DRZQKtoNXyTcDYsWQt314wNFk4gbj7v9IxNBbkfjTgC9hU/QdjmbtK0CMq4T0Q7HrudFUrN6hD
D8k1XvaI2Tk66rl/C92TVYHyStGXcFv8LbP0Wkfry7eXdnhlc/5tUu8n9ogebO0+985QQbtLpF01
tR+BoVmOHkP53j7iClCmQgs3f1OdUKJF9wxlkfLHLt+lXwuTCOvronfS884sIfmQhc3VR1g2ZrSD
Fx8gv+3UhYr9YbloyjjrtCEEhV4DFR6jXyNk3O6dQ2V+YJxmXU36aMoDHl8f6vAsUAwwiAeiyoiH
zYrMIJizRdH7Rc2UD16WOnkm4yrSEgJgRNYdKX+GLm3ua3jT6Mk8x809xrWV5jA63pwcRUaqs0AF
MAb1mdtX/JnOh870bWjaZeSzQkZTLv4huidYdtqgN1V/a51z25HbXc1elJt7iJcPrGOpMrspT1mF
RCZPVbMW9rTUBbGJWhQoG4GE0ve/aBfxliFDvLeWGcZuNwUlxILff0WhNgYH9rr00RQSNEPyQKEB
C4C7K2CctwfUeL9gmbODpIVJUXdigaM8vFdoxXGd67MRdIU9rcade22kwPFx1FFbDKhQju/z5aNh
D0g8aLoCfbP3xP6ZoxZ8MF4QZ2wIUgSj/ZbOR7v/V2uCr1+rFgCUMoBha5gmHJkUywiZlAGaBKgY
7scP66tzZg4UqwPTDNeikSyQL4jYTLRmQagbVXLLavMMr6sdMxvCbjndRpey/owdgI4G+uT7F3nD
6sBv6MKU8DO13aJn9ayqnVHnH2DbBAHguZO4PGOqV0TrlY6I7QBrZWkZf0WNOUoImbx+B62Z3HIv
T0h12A7J4MpSFWj3whl1/Or0djm2CH9I5CsUitSKT5D33SfiIEAGu1TySBWWEenjGePQml5+owR/
gpVQ9PxLm7/RCWZVEIWnYosMVgb9nH0uYG15D1ho6leXKXJ7pfbtOf6rMPDWdGtp10cmK89NY5N6
ejVLdyba6QsvQraplmx954eiUKxV0QWJ2Q/pCaNGganZuDbJB/ukgWN5IEXayFRFc6nJrXxi0fkV
CCo7y62noNR001zBQWNIMA4Lsc1lD5aydf+3iw5af3J+P06UhJ4lvZ/Rh4SNZNAHL2hRCue1qYad
/JHu84kChSMqWDwKMtTm5F/qEKBP11V9jALc7MxYjGwCLqVV9NS8B1ZXG9+cFFd1Ejid0G0GaBb7
CtXbpNPAcjcpL9a6+JoDRZIP3fHNsZrVZVQmPMmf+cuArY2gXxZJ5ZUr6+ufGUso68FWVyVNENlu
hBVpe9A4f3EYyaTnppQyGp0kuPgu+NiU/Ag6zAlkK1nfnA7Pb8Osvtyn2BSqBR8RqrSFr1n4xex5
La6+UmMS37yZDpbbjobXkxpIe/ydgcJM3cFiIwxdMKVzaYm0NtdgeSPtP1/oPoisqSkO/jTeEogk
Lu0zwUvH5ZbTO5vJyitx4DIcETZuDv92vpuH1ZnoI453niStpNZtOWJ1WTwlBMtOm9W+0f1HtZSl
zn3RT9zGpeOFT66yKZx7nBd8HEtHZaH0Haw9Y3d6Z79QVWKKS9poJNue624XNorO2HM23qMA156j
UWW9d2kiMYjjcoCryvbyuGrsQESPtKPpAhkSS0YNPUTK4DfSjmVyLeairZ2zQnsgHry6eL01KNH1
GZvnIFIz/ENXXqdj8h9n0yKnL3z6JlDLdFXyEkm+0YujY52cPhKzIagMqihJSC76rEln7Xdm+Bmu
SDN4tvV+pqvslALHa4zeQ2qZw7mxC0y4dAiJqFOLS05GULfz+YlltsyXQKp09a1BarJGJ+lPeDjr
IJVsTlPwssvYpzgM3SODw7oaLqZPCMYuVzvyKJVoaWFFA4mPZERAErGh37Y0uVtntIZfC5b1tXe6
5SqZFussOdQBJrH7mcu2EZsZpeWU9MviZ4tDXfjQUz7mP4rrJPhGag2jIthwdxuG0wseaYzTzuA0
DRWE/eSXk2POx8W1hSom1iLXhtZnE4HFVl7FzMDInELVjhEk2SDchIoWsMUOG9qltUHaxeAXGVkM
PXf1MvHC3QYl5AggZHfQRcrRBVL791Hp3FamczSsNboeOdIlRsG5TUMQYv/mHApXhD/8igq4GWD+
I+/rqPqLSrfNnI0DOmsIuAJ162kEnhkgO4vMrSifh045c5xhThznoi/i15EQaxk6OnpMUPM1kflh
ttHWrHNhNJjBgxhHU6wRrxDZi5Eq8p9CvoH3hIVdgt7B17qC968gaIhErPVBMAZewFCQOGNQ5Uww
EZPhM1an4xv7pH/av+y4xjnM/9YcSbPErEUwhQZ21JhzyXU7A2ssv9Oo20vl9BdbO7IplFi3wwpR
gEh1rmTf2kArwzUtSAQy6HJCgBQpc4DkB+8wUNwAhgYKh147r9nnoqcD1BeAWztSCasdXVEyy6tt
GSs5otoO7n3wnBcHeCpI4FDBcCV1Zd9errHWFc2hXBwBxSOjJgh5xzDNGzWfP52nT+2FQZU8Syrd
offgvaJcZuneQTPtv+ln+eaUWW/B8czdHSrc3brJWejXOP7bvQjd7jPWYkLrmlXOt5q3B+s35/+j
UKE3a9f2zGDBXBP8UwIH5BwwZIetN1OCdyZ0VausN54orb1CrbUBEfzfW8zZ78IGYvXxf9el/zJo
hFDjoFA9+jw1PZzCQBPZd7ZybGx2d/MDHmYnnj/sAXjImlQYpGaZ822bDb3UuRdiTupKF0vUHkBs
bm6OnWwARcci4BHwU7yJLRkt9rSj4/3Vzk89+dhwviX36LMBNMrexpgLizegDNwoaK9WV+lHrROv
Uskmjf3Um6KTz7GknJsprVbpVijG4RfhnRN2hUFpXeXiPd6Ea8+AcfGE39DVW6/9Xevv7WnuoO5k
ujkPyaNBWVWfub3b7QXnzfTUJxYcxIkvshJl0WZ+jE62hXkd50wJuSqYXdnwFOuS0Y4IuzvVL4R5
MFBYAr5S6UIT4h0E4XuKJgRrGSykYwbnxXWKp+vxL02Px7Iez8UkOuWHIAAGz9317WHia6FY9WPH
vsyYYL8hjEGI160ugI7Km/2EVZnV1C/fowXAkV/Ts+sqCSJJsLf/ZBW5cc20vIYKKLQiwQiR9K3s
CPx8izT+hsE4Y7cpIRPmNjRwPKl3H6N5gn3TH1NpGQyp2VenaZKmapQIhn0LkBi0RT/aSY1skuiq
ZxcmjbGXyS/wTHNQeA8V+yTymsS3Nm6/Up08jG4ACZ2kfCq9vTjs4rkqIl7Itb0heWoG4bZWpk4K
SlQzyaOQJMivmEdWEhfV88JImnx6c9qXkyivK2RvTBciAY15mWpm8lKjGflJiGIB4RDhjizt/0Jy
x9AfTBZ+TIQSaUOxiz44Ncy+0Nf6jVF9lAeTxo1ow6MXHwU2CHrAH1h8XpPN1iLvC/fLwYmpyNLb
CiMNu4F3dCe+47IwuJurqfDrgdVxUHVBxJ94Mal5iZrLymKcfZ8AhTuK+89IQnotpPB5apyRCtKq
QqlHE5g9Ysqb1eupRiYWOlPQ/Qw6o3lKILSvUyUCZ/20d3wsEsMAf2TPUgZSreJ9kZaW9mhOju03
LIv+k+Y4bM/WxXQ87v/dOuiw3t/wsdPST3Ao+3HJgQwh7Rhil7AfYPlFlBqkd9Pk649EBvm3uirS
0MnKmK8odsYHrA8/ttxLjcggHrpVB7pLPh2p8KGldw7Eq4WrO680H95E/j4XHD6juYHw5WoQNOjI
phGvl8pZDPdgpF/BLwEur9+lWFDPee4HJ1Sqj8mZAczYdapEM9TzSfp9t09HUsPdx9k+vkBhH789
gWXgILnkqdGIHAPeroDxJLyJLVllM+TEAMXWRqs0uNJQBi3qvyHWBQjVI3fz3n9UUEzcGX64NDYl
Q/HdMNvX0/Q+pK2T0qT4wDAwk5X4+3D9TTg42WQlQR8yM0dyVEDn5a/QMw8K4zMSD/snU5PSDnfW
+lzWCB+H+BUhaiZ9QVrnSXCFDWkaDxDjEiSYoMO/ra3yYw5kVKP0hZh7U86PlIkJsUGxwfD8PLVN
9Nh8PtLBN31y3XOtXQghk+lmf02ESmUFBUTrWaFWpt0eGdINgYjxo4hKM8QBa0Ty9i5TZK+c5PLw
GoLf/q/oaFDOe/xFELlLdm92Li81x4TUELUYiqMqXhSzEzLQkoFYQw8/4yI+JmTJnk9l+pLCxxMY
XFtFla8mZULQIb31rdTGMaSnjc8KS9tYG9whd+9evDYifsDIIP6wWTMIr8Iy6oerSKBIOQvklCby
t8eeG3T8LRwjuCuMhEMa098Qy79yti/SPthhlkyddXdVSSMCfkz6bjorGp1rdXsB+nSlEy2fwr01
/55k9+pRVOI2RGRxRRqFELZyMooHmQnqwKnU/vHTs5xEO8pcUkyjx/XAtmZYQzKGjXMP+INHrh1Z
4e/KdqEipKn+KwJ5ELCziyERL6BiEDEahz+rkiJlbrvJGRlXPC4fL2Xn8ltUTpPHhFq4rlP5vjPr
T9OMrrNT2FdyO6S+eTZFIRs6RwJw/l0s+tHZbtEAutYFS6UkYxtQvzne6fj8A6BD2u+FQ0efhwZE
yy0zpbp9USIPAY0ed7F2YU6sQdpPHlUY8YMQjC6y/SgbPEUqvtr+3dyMiEu60PbvAPh4/845m6rN
jxu2CodEQlnVozkWx3B76SOVAsXff5MsoKGvo9hi8x2qz6AZPv77aFa9MciNgnhe6XC76CeKDTBf
XNBWU4lHjH05FkflSsVapFOm+oCJf6o1qGO2+L2iCYGbp3uEpfXDVm5dl0Og9bVwQkH+3Odnk6yz
mcrM7Zjj0rGU5SmuVC0mFO/sbVluVvasmOWp1X1GfZ932GoZHBfBbqK5V5lA7l5LnLebR0RbMwYA
As0adBUuYUvjW5yOnIFmiaX9MPL4YA8OP0ADNi6FgCD8Wrj1wUJM4N/ErfTgvfk0jbgh/N3BhSTF
gIxec9kMeFnk1XAhsRzAyyA8vwVXAHLSAZ5hwIEqn886mmN+4GDSjxaXT4+vNaaMBsm3V7qD7W1L
NeQFWeu2Mf4QcU0giBdeE7eJV7YvEtMekAMWNyir0byWMJlW3JjfQUg1+6BCFFxj0EhK7r8y0ezg
OV4Yk8AJhsZC3woxI5OEEeXuZ/ktL4ivlTx1uKs5yucxfVAEcZs4jIESPx9TVIPbmMMdtmFUset1
RFYC3MkXFHJiRxRcn1U686tNBTCldb77wZ7rPCHuBF6n5UZufCGa8BC9dMayb1fTBxt3oZRERf9q
w0EkQ2o78e1N7+xdQgnM4KsUWOgDrZAylUHiDZnfpdgyA3Yfllc+jUBHZmEeibPSU5MxDy5mgKwR
Gw+3Qnkrw3pQVNMeYiZ3Ysu/UUFDfSO/sJB9DA5ogO0qMnHIAIsV/9LHpQbL4wggdcISCGZqXmo2
H8WIpujB/CDfgBX78ntXeuLK6GdCVThuSR/a07Y2gwF7sSomJsOgw688xtRWv1xa7VAUyjjiG+FM
u5XGrHojqHmbuaUYUK97xC5usLoAOS4KefIStScNs9wEQuLzgUfmToUCiM2JeRIluOoQuo76ezno
Z5DauWzrSoS/p8L51qDcT1SnWhwYuth5JcHP1qEmmex4WhYM60J7XNs+jcYOiyuUObTClmaqhMn4
BnK5m+kPoKUOmjRFVf5Uu0wiH3XG3kvx/O9gD7aK8bDKh0AGT4T5Xkp4EJKbq7F71lxy3CTBGVSW
o10Y0PuJkvbSOexQdNd31YdVBkx2UyIhAWd85UN6m6fBcUVXsLvqQM0ORyYMtSgAoNv0ajIhLert
rP227/J/0lfGvymLDfqKkWSrCmG0UB3m3Y1Nw21rbrRa2m8uFxu8M3Tq2x5115pqhjv4vjhjj+FJ
ViNdWIPWWrMS/tz3gWGm70BBul8vevvZia8JW9kkBXTesCOQw6DGxQEwkU1PJdGiHoy1jGVrXTpk
Y+LA4h7tV4Gk+cMlLAgSVbkLwEXOhem01xUt0ETzQnoJtweQLaiJwYYn4yy5TFo/scuy8w6MPmJ6
JJULg8h1KMtoRKCXBxmULRFzFVdzcE83pE1YBjL1+tPK5N1xobjdDfwa5jnXUOMZX96twajLoyVn
mRk8Sj96leyTe9eg2HVTz0XuCREz5vzX4Yiszybok5Nk92cS55rl8+pSZq67jNxqY+AIsQwmI8Ce
lCkEJ/QVXXkvfpi0oY6jA2ukf/qb3slPkSjZU1LEep2mIBtWRBC+YTte2dA2rIY87urCpW8t4aw2
i09IJCNI16DGjOkSH2yG3rsAGzl2fPTynyNFrNQzeFWdua5BUZdAG4oPOY1GjODjnxizA7Y82aMh
BKxWNkAHwemzpN1WCedhddvyoeSH32cS4yNZPPG/36YrnNOkzVZ6Jia6h5DXm9SkzG+jYS/bNiTY
OCGspIiT496BUAVzaSqtJlI+fNSmdNm/t8PG3AArm0/O+HUtWbF2CzSMbr1KhxBwU+GU6blrek/S
759TVQpi1lfInWAVdQ1zEI9mURKy7lY39FEyQP5lOrFMLH2DM2KUn7gYwnRZ06LhkVND9E4Rvu4Q
cY3crH8RCfkZfcL+9SWxNnrnuMRte7XpY5qNAzA5Qa/YFJTB2XOFSHpg/0uCUgLAKBErFkpJMIH8
89q5W4rz2DeP1TKtCo4ZBjft7hmRhc/iZpfMtQ1RKPnl9Sac0zSIQTdxwPLe6t6L9GI2ng5fS+Kg
Scl+PxfdULag9Jyto+hjx9wCRv5xz8KB/epwUPREYRtrxNfqAgjJHfdrjHO/eUCEAGqUck+NWASw
c+GZBpcVFsuv/rmCoYXijg6tJE6rsykD1gmbNvB/AvvstuXa4NBUZP7hZnSbe7ylktYnsLAb2L9g
ULTxpEzhk+359Kt8WS0q6aeE1i5xJvvW+iRwWp5argTVXnvqquDPqj+rZjEQUt55sdrOMTYndJzZ
FQ0L5cioWYakkyOfJt9/1uJFYsfh5H1RZ38tHIFlazQuatf4ZfokLXPhAolSz1MhtliWcj3N9aoA
S7bT0s9fAqPQDAJr6ym5h20nDlnYzTtnmIQeDamItBfoUYk/GQeZBZDZDAkzKNJXB/UP7I2fkajd
YO6vcjL6M3X4HAUS+cZnC5hov3S+X31pQJxFMKwGWnVH94ZB7k1a3Y6HJogrtf18lMdrsdbeQpkh
/gZAomQF3huj17/4tbPV73yQjRap1GBr+2gcbOXfT88cFtIyfjNIZmtrp/To7SWkg34JPB7XmQZn
4Ds2UC5hXGC/Ti1CVTdlKzD4a4vffmg2NYa1675G8II6ZrPBLHzWe3kixb2ojtna7OFPO31sLSE8
L4ZsCzMmTsLhrb8SC8J5AWS9zxL7Iueog19Bqsk4ALE9nl0fzurileJck0buVLi+H8+twDJ/lM/R
FO99hnYtaSqQ1eMK5ItkMIZ8KRzxuempyVbYbDFycyGIhC+wlmht6Q4V3PgR3KPIbh5Ddn2gDBmF
Co5eM0YjZVms0fP6D2pc7lNqsL54Q4YSL4cPUWDOjaGx8owCFF+ilVc/nCfQaadZyCCpEdToBiYH
Cj+i2rkHsbuuKTxF51d/aFn0tq9vpTwKzqJCPaMtv+/dh2v1H7HuZLQsS0uXgx5gUvmZXGNBMqxu
aiTgiXacA2pQ79V6Ch+3JPKW1/c5FfJ0zwoLnrT6eyEUc0fZJxcEPZJRvnZjx5AYpx5/mHFPAHTg
pzwt19V1TtTZAD3pGulenlYEc1sHuJNoEWrVD/mSqCoRek++IajxNHgqFw1QYXqo96p2fEdKLMy+
LLP32QpiiEG4NxypRDo+QjPGZOKP0Fp1RT1nksvoFsbJz+uientyz8clPvh3ystN5KeB7PzBEXNu
gWCTbZQ5zAU2bCdbIp/8L2dAlgeToewVTMPr6jdpNQoALV9bxq/bErSZaoeLtXFgAZlIyU+/fKem
zkwZr/i/o/TchcB4UT3wOs/dulCWquFrUQKMb5FhueXxORaxuni3Qb/ihnismayDfJBvrojk7wjc
5NZYnVhASbn+RT6XnOpmJ4hygQ7D5qq8EBmEUiDkbrn3tPTSS9UQSLT6XRNenAHesdfxnOr8WiQQ
0ilDy5+P9HuGyiWGvKGC+eWlqevNFVkdhSLZAUkQrUspXBJtbWAcqK8e0XTZf+mGLvxQrU+Hxo8Z
6xBji7Yf8oEsOUU/qtQtfek7whu/svlMYNC80B0abl2tiwoqNTcTQgobUpAGuxlaggSJxvhGKaH+
glvSJVXORKSeQju4sxoWQZrAF8PNJIis08zMhH6UF095qW3Z/j9i78rlzzobU5VOlL+ULXmy0goR
POV/5Jgh8hgq3z+FK8F8x/5PUvmtfXDBs3go6R2TJ4/Od4akd+sAbepvsR3IGdmGBmR12zMgPsKc
7hxFBHhlWxo7f9lDdU/rCkjMD5/GlQfiy5AHHg5WQkXFAgaxJeIAuElXDZz/p4K3h/81bKSyTwd+
CiCUUqxtP76JoFm7Tfcwe+gIeCz/LmqRMP/fCWydZdYfY4GA9F0MDaYE5pO7mNwVr0YVU7uW9XdY
EloaX/4+uEmk/iAv7ehcE9o0XSRQuakw//2cXOAwDsBdIId7Qpf6j46Udww5vCRni/4KjKi74dv4
ByJU77n16q6zfM3u/JoLQpdb7cGQTjiArpHfrM6OB2sQ4GkRqoUimxGZI4CoqragWQbOzW568qki
14Qy2DfJYCpKTdN9cxskUlsCkKMjdwy+nCFVyl6M0TvWkyqBHgZQ83Isz8FZ+odRdYu5H/HAl3Vo
2G+EsEoZRo1JlZMNe2HSrXNuOosk+cARusVF8t5qCn0uy/WBM4CGp1+MFbEn7TTNgZEEqux2NYTP
wQPR17Kb8ushLEm8XFqwTa0x5eVZQHLeMPLRyXjQmIu7Vm92hSx50rRdr8+agJ9qHP768vfD5GL4
M3NWFPsCCRdaphLMwjnz3V7xCHouvpDs3fmRZglxiWvr30jn/y3Bczcp6ZZDAAWa69PYDEyD/hC4
8xbnuU+zdLUkpjFgtAU1r3teLHFwjTAhrZoAC2yaMKUSOuvRdj572mbFAWc+l3KOG8XvebFcPcf5
F7ucLfL/y2kf8Mgzqx18yNQh3ewEDnIVbxQ3yN5ORASkOIOsEr8L6OGgoBxTUtbEjJTKjWt9KUAs
GsGfCuY1HNe9S62eJO98iFFFiRb0ctF/3wuRElh8P0eU2+R0N9IIujD41Bn2y0L09HkSr2m3pOtc
m2/XpG40PhRhpXhrCJmz+ckc/lac4zYM5NFJFcnbEllgKroqeRme9oW/RSkYIhRb2DaqguNtJ+Qo
8fkzNuuxDd/lhyEgGkllzg663yeObBD+p1sdZw1a1pUxKaCOB7Ytrf4gZfsnAndUzSfpLIdLGsG4
hoCxRK/2KR7Hs8b4P2zDXBgnfjAT8NE7eX5igT688oSZwxva/B/nf+7kNsNmSdgSfQHvjrgJyywt
Ag6JI0fnlK2KAg0vAvYNNnqcTR0oYiwjOmZ5BrOfOOfa+lpvi5AyGMrh8OknEyo4ZOZZze6aUZ6U
OHiYwkgSHStQEdS9gm3iEmQoksgeqA7fmB+6vIub1zOVcSIFVQMmTQF3B5vOjbju+gq12tJ99u9l
mf73if/kYGCGsIxe/OgHEh6nA3gF1hxy9EY9GW9hEdWKG7j6cz8hDsYNnEiI597gq/y3ByBAF67w
4Msv+8+nEI2xMDs4+jo8F3ddPt7/bG8Ur46o9mdcPTAPSXJhA5sDV5GXn81oGMq7TtL9LUCu9GsB
rh81vZ8zvFiKTT57c89A9ay7ym3798nWNKjLMJwAXfMXr4cfK8nQtSQySjS3goft0ETxAUT9Djy0
xpRcJuzhtu4aQUAjJxP21CIQozMQHHwrWQvzrTRGy9lpu6gORfMaLyYge2unwd1r2+nAIl2TeQ7s
rnZmyteNagN5mbzaa/1o0AJFz1Dx0O2ASerDLwKRvHjSZnC6CmwMymRlre0CfCRyZq5dgsIWfI59
CXYgUMF/yuvKc8kP0cDLr+ptYaJpwCf0xNX140UWoxG122W7vQ7uuY3xTsOITeoCyN/WkfJ3JYhr
SlwHnh8JI1k7/emcMCoYbQIkTOWWeqCHYodKjdMHO6HBGp+DquEdYXxYfcVJd3PhEBhBVbfZjx7y
hGJq9NhWF92nJYQ+tKk2d/3QF781CRHj6L00zxnZURS7mJCHZPhdQ9qO3XkqhPHWvhE35s9wPblv
f1LcQ1yNARmNLrvGrkTWicLaTJg9ZCiChXtk42lutUqFVJ/fXnwPRVpB/ShrtMJLOPXSlpKQg6do
k6g4IFkgz3OnrMKWfHT7tPfV5cHMsAh2494R5zIe5v+ZwqD5UoZ2f/xCtLtm2E3CTduW7KLRc56q
boXF0HFoA9i653dDzhQv1d0uZogiIP6hyXcALtdFrjdijrbShi+cy2ddc3JEbY2wAzkNtRxPPgRn
7iTSHlaritMWO6JgDuEHH1VLqRDgDm7Gl/9P+P2+ReT41F550s/5WfHMRadhC6BP6wpuJRhYWOtj
m+Da5l43R7Ej4ibmSqgQ8jttMblJONtDsEYmYI3tpy5FjLp8JXySibOJpw86tYc4VTTVJmQ2Xagx
xKcdBqmUyK8xS7TOOFzjJZXjewXTBJcGk9XOX/Qiidc0OFQInmyvArpJuSKBbBFQ2qNc3YbNVDqA
3mWmLD4YCti0C4EJrxSei9HQnfirHZ/gvRoK5ow77BshcDJv+LasnDYXMCsocYdzv5COFn/5iw/w
cpAHq+NvS+0LS3F/VmEYedifvcz2Z5blmrqDtVDuOl1ld87ZJ3HHd6C9+FepSpHAoV1uxtyvMiez
vVfvwm5fluy+xHOpXTdaJy1XcyTS/HHAnaXibtzoJ77goKZu4xUyqR4WBJrXw/VupnkAgBtSPvZL
4Jhzo9R2+2Hpun3r73sraC+bMzY6EHxkpOPZM/9PjxvImu1FN4Qu9pELVxO8FoXTHOoXsNGgac5Z
GbhIpUpy+95NzPDTmXoPqI4EdNBItZqiCd3NthibMoEkZlD4BCr6p/JX+wXvQzflUMQ0d+UXbL1S
rkGkglvINmFO1oYjeus2sLsU4qLtBNAEJpj1wjDGjropmWlCOcjxVt15AiQ7OUMjN7Vowyk1IQFo
895SpIL9s1YtBrTNvd8r5XZg/YKUXxB4wamIWKN8jlFG3lr71eeGlc7ks4JKqxlA+o+zr7gzNr7o
wJBzyxiIbVMQ/HeViF0VmusJIx1tytkPhzyxLtLbAbk+7JhLydozPTKoUjRitahUlkxCgbShomwu
AWoD30JYSikl1qZvDoM7uorOG8eURQbSAnvKOrnpxcQonzWlqiVv6FE1Yeqt+QBbBVuaHrkIycpr
CXxT+4VZguw3h7HnXPcqMF8OcBz2rx62XnJD8MjvbTuScyp42sHZPL8o/dOdVbdhk8UjQQdgJP9G
Hp9I1UPztry0JWfH0HLzdIb7p8nBwDADYHGjhwQJ1oOfHYzeQUMd7nGvz6BFz8nc0xvgtpU+4+Lt
WClPFaDeN95pC9dS48CP9vx96otDI/UaH+3Zmr125R1ICql4wzWEoqh7uLTREoobGWqW3nGiOJ2s
SljAByS/2aBkQHZyF25j+6Ttg/adLbwArblcNcXi3MX8YOTZKN6tV5D33CAWpye19cZq364tGFjh
0jsZDWVGH5TOSLC+A5JqMOJpcdcf0JOonx6sPVHRbj04KXjbNkFOuyIKLjDmqisvMVHI07pKzTbA
5J3m3gw2ECLglgfrLqh06IYnkjsYVSF9sfuwQOtjh0lmpNjrhFvSQjPeRBMLghibZ5/BquIl0wVT
mSOCXpOVYDfa/9vvuYyQD93sVNnh1Fmm9E163rS/waMX9Dk0C70bYRsnVxw2oJ4macstSyNUDKNs
p5e5oWr3qQzv5Mcn9AE2xq8icSW6sl2HKnNM6/jcr74hGe5gLtfpecbDwv74gytsxj+m/rJwUNwF
v4FpBNvohWN+RShJWoUirMmNVDu3YtVfPv/MW57QoRwH0x3xzR/pUQJfhyZ/64ocjUW6BEojCTfc
bvQi6OuNw7kXAfyHoFAk/7NTzqnGgLUOtDevZ0vqKaKeDe9Z5lnn6+NB4pRuTzVWWTnOyfXo15Qm
txziwPpoY2ePseG5xYV05ObIgXaoMi5Pj6UMsgVM4qwnBADiHApVPCoJg8DJUxnj0DO5YqFenabP
yvZD4mwn7Fsv4H6yp5L8cKsyFKjYje08k543x4PRmf/m7qwau8P6q2Jf8XKyPH9TdBoh2USs00NW
KQGCKF+Ph4+bllZmC3NNDGIWyfVCv9PrMEmLmSmX6Vg+E38Rc7IJJXewwBYjY3mfkoeRj4k7K7Ly
tM8qekivCmpTteERGeDMvt5CqSNk6W375D26tDbawyle0ylApzyCPGSS5IqfCihAS2AQMZMMryc8
gBGpCiH6AUXhl6ltdLCRisp+OqBxqxtoTZfNHm8DXvlN7ZN2HPUjanecigLXA55mMLw90khBlv4m
QTmyHWxZPzg5pUIdF9246Q4nKc7Dw0BDiCsD+iJ6tuKOaqBOETvkiNnH8y0q08LYr3dy7DmnOvEl
TQxNDyMy0xyevveUGVQinglDyGofq3WL/2WNMY8J5dA91/9DdzMey7WIF2GR/r7sQXsQajZPgHPb
b9kECLCtt8f9TMb1+kwga9tsdofra0tcR45HQO4mZAQ2zth2kGDrtEKo6RhXizJS3dZHEXUaMU6S
PvfopCeIz0m0zm1RM65K6onerQ5bP+6z4gzkwu33mPuK/gzClGnCCaZo5AwbPCSv7lTgxLKRAzdC
w3Fd038WW5P2tRgasFTS6x1mELIjCZqt74O6rtmbOsR7uZTJAlV9vzbVU+t/jx8S547UsLa/rHsw
Kj8clBPJoWPOEeDNBRviNVx9UALTOLo0+SgwwsjwuCY+DO4MjkmLPDzOCOjK1AtNOHHv+zYmOf/C
uXu5Mi9i9Bt4//nqseB9uj1fYo51KujuFaI2qYNMkGUnEiGZZS76RbQSpT2uPrrHRIh0U2DOqrsm
X+TNw/wYJ8czL3At0AhZ8HA+TyFgjskK/d20zs3fUfk9mD8/3gU6yWgZqm0ZXCcc+l3pb9Wcyd0h
PhZGXigfehoiTt4LH7JSivBwC5Xlh6tbnGWC21TbIP11m/GyFWzZ6UT7QllHaoWrKUfF8fpyLzHs
6NuH0iZjZ31OMrIsg7AtlFP/BC1Yt9RqZVTXm21cX2hdFQ0aKQyhz1VJSE1hc/71384oRHTQWPj3
wfX8JWJZidxZ2m+XcgBrP3ejBx84z7XLFoqWI9lp5khXkAboLFsveQY48jH2nZhaZcwd6/5JQ2PB
Go38Mw9cPqQmEgddl3b5Z+tyhJcm6hPE1Jk1MabKChq7wGXCt3vJ0RwqUdqC4PSLYc3WNb73ntF7
FXTLXcxre0dHvnjZ/10sBtRqINqmJLY86bURyu+U3Jb1edFa44A8cmVPN01X+9jKKKNXUnBAJYMJ
U3REmuGGsI5k+J+02BWCzNtXCN5Bg3S2n60+Sg6wX2AU0dD4TB8qECXuVcSVuYOEbaB01JcM6yj0
UoBtspmjIX5GYUWTjFvzVC5ECYARF2OM9Skdh7SPmdtBaNr9VD9c1fEAedaTfpFXwac+kfb3ywP8
/Xcg+pHnT+aMVraP6QTIS1PPNMU06QwX2F0aL0Xs4oRb1mpT3biTVPOTegko2OkTraY01SsKX81J
sIv4tojaCJMZ2uiw9LOHEdSbF6BucAlnJbyN8V0atKQPnCZ4lafoTI3YTZVuWzfBCFpIIixEvB2C
IAyej/Mra9pPpfLaJ74iIJMSImHGgnYSdj643i+Y1WN9PBDC9a5bkHKEVh8Iz36P39ZbriVFfua9
rjd4LPN8SfRPZrYxB6V8kYLIuiFRoaqTNIjAfKP3XyiAsH3Rcl+q3/w1MgjiOgcTguuWlXTBpSFy
KuOq26tpXFsRQpPVUhZsKvZjYUdIIuIrgOB0gdkaqVrdTkGikavtLHA+aF4EWaWr9eyZNkPAQnKe
5S7Zkuc1OIQBXteL4Vh1Kgs+uwV6HPggOdgOJe/S9B4HJCooh2dr92UagUlS7SGATeB1RBpuACHY
qm5ZOTLm5yS4R9qNNAFLq61aNj07+EWX5R/rC17WkYnyhhy7RCPHvHwvVIkwxB/jUjOJ9WPHM3sM
pDmY4wOvoTDi+5tK/vdXIXgklZFYoyY1k/54flvzEzu6QT4roEqOcqiwkKoqYYSKYCppPPOg7Uhe
0eOF5W7EvCG631zkZQFhvVdgH8CXRn4PFFdpjgn2vmsvxaVJb77HjucniJqf63P2DGUiCYiXt7Zd
/TVd3p+0cEXKSKI50wpQCkQt0xm3xTz4e9OG4Mub4f738x9dZ2x92J6HtCBtHya6kKQIHdRi2L2+
iUsXl2t1rkivRDARLopZbAVg3k0tnghJ9pFrxUdh72yvOSvRi8dd5O2LcsMkAKY7FVMEZk0aaMRI
GBE5gzcDcVEsV5UW5AITrOtPK8bBlahFc47UhgQ4hukulVIyB3lSbwKmQDH3K29laieNSJhncivL
b2YAV/oncEZeZ6tQEdPW/uxG6FhH4peGTuCtEKwCG4GsE9S/McNtKrG+Hx22pw/gOmWzVUMEbqFE
8OFxpx/DTWmOfsVFIRPOQNAKsK23F5To/2zNjCKFf04p0KzaVGJ4WOdnXanpbjVPq6kpu1vv6MsY
yTjSMZwIxR+Drwl9cI3o25CzXgq6b7fRkeI7IyVmG8wo7V6ewjY1u5s1lolS8fr/HSbrfIoEqIt0
LB5B90XrTydB8uup/tAIs06hZeZFdK+i5+W0sj8axRFNkX7H3n01k+zLFHnZ06je54mWQhtzBWsu
7CrxOnCSLtKXQgV7xq/yM/XU2bYcMAME1vbdTHwCBKNti3ctFHWU/3SsAfsWNyUsNwi2aMhA1tAI
yAQx9m4rANlZ+MbZAQ/3EddmknAFwHx3rBIuA9hEw9yxKbPexcTX5hTF/XoN+uhhkFqLOsDgehLs
wWj0fg+wedLyJO1YhZZ5lAYgEij4YLueUVPkoa+yGFq+F+ic4ymoXFVUjiYpX5tZ8UKBpRYKk4YO
l+rYTkMd3TRDVknFBMaxPL668dunZEsNj2821BTPb+Qi/fa/3wYyqx82lAxxIVMGdV/GQug8QvBA
DNVjWSfSYLJ8CbxePo55K0k++6ML91rYyvhX/g1lsSFfQvqul8ZuP+BXSnEi/XbL8mNIDbQ68HqR
cknEu1g19ONE9850DHl41bI2HYMiyANGOR2DiObLMkmkyJ90lYvO6UxxCU3n6g/uhtBsg2qmeJHL
5GbP4t2iO3AfbB6v4OQ/eGzjFZcGm1CbHGFSgyW9TE/cB71TVzk6ltPSngOE5a/XqlhyVyhT1dry
wXXKaiICNgB0Y11ByrMEOJIiv4lnnwB854KzoVVkzMwtsfUE/DjChHVFPJaUvWkl9NvwAcOK+T29
Migw5N6OndEl8O+yFLf/d4WRzDqteCaJKSQIf3h4y8IULcZUW1PAM+wgrk/OTonRcESsouBGaXyO
Irs/ZIYJ86++/c53bTJ7iccg4jmB/2o7Ca2wzUih5ENgkB0Jc3LPYPj0kqqQyrypcPeBe+7+Pkjv
s9XurTwKMPyegNDkYzzvN1z/ZvvpSKlGwNBiJ8S4kfFxDgf4ZR4DHBsD9wxsFWuScb9X+h/l39H7
0rhBFiI1OLTWAGlAGe3B936J/wZb7V9pvHMbHEroj/9P34x+7Pk7o9VbKkFii7e1CDiDuENejoNg
GrfKWEysWBFIkIioHk8ns09U+QX4ezMJqM0r1zSNMhPFLDoQ5J3fmQ3R2O8PKPb8Al7aImrG4bHC
MaizU5jB6h3M/mGSysFj8nSoNTAS2XcigaXH9AU1YIZRkKRbLwvvAhVFjHrwEtLfbfQFswJAIbcE
xEk8MEvGfWwdeCs5i1t5kd3c9W2u/lEZKEKLsC0edlRqbpU1qosikfsnOnZJ2FRZ8ALl/VJE0fHz
MewBgU7RZiySCHgtvRAJE1m2ZUNzcwIJYbRgdoN3pVvY/LTvcr19fyUyLHUFM712Cx8UsX1j+U86
qEb9Z0b1cfltlAxt3QphOysKQ5NS6RU0yrffOjrdbEnXzmFONPYbFPNz+7hDuog9S3vOZV/pHMgl
dhASA6E11H5HEuELuK8pN3jASl6YSqy7NP/6NWJwo1Rmw4dwiWp/YGOIF/LVV3AS8yC3JGO7tTi2
wFl3uFSTBfkGHBKDTZhwnPIP8yJxPxhh7PO00WksxE5uHaaq48EtEC9VChtd2wWvfTR8X52gKMeI
Kwb725xlJ9FRUb3qwIF0QBxYXGHOKN8XFVMatoYnVMU0sJ7KcTw6m6tMinHpKZ6VeSpKAk6VFXMO
v2qVrhsve5zk+gEPveS71xxaep4KL70LGvCrvcwSq2wfYrbyStabWtD6T6yElKevoOq7O1dDTrQJ
MvkfNMsMRS+MfruC5ecg9zZRJpDKlzwJRafwNduU3Pjdrj2a0RXDkFthtzi+FHOrCtDYgLLRYjnZ
CJQMt7jgsYfwmlUEVvujthZKwCOCD5emChNCcRpcAyar38PnMEnIhd1Dinq7vvE9BzQtSaLwRl5+
B/PiNuafx3aJ33F5aycBjD+o3xE7zpOkRGMmw54Bgqm3xi0i9Y6KoNMr7TEKUgHMhkcFlu8Q0rgZ
AzB8dB1v8TIGxQ6HuWCpshXw5QuoMGYlZrCUHe4JsNPM+L6VRruycmtMf/3vZBnfeGYVSmVq+sZO
Vep0tktv/yjuOYyM+CtEML0a1QFDoZcVT/5ZLy/wz/uw0J9eF3WaelM1hO2wbY21E22mV+vuy1ZN
49FoqkEJpCLUJaglcvQavlu/bDXE+u3LDp3cST1SfGCrOGAXbT19t7TVbjpwba3FYi9lVvBrDXtI
HG3gqxmAGLDy38kzME9XkHbAjqVCPERvGeM7pV5y8k8ffS1LR96lwIuMK6anVfLKaBrYs07HXGaX
hueAiJ8uglOfye3aPzQ+NHEJU+sPQoLm19cHrXUr2Qgpb9BrcKe0OBNTlGgaZFtGKuoYaiezJVtU
Rh1fa9gFPJTsnfa4gjqK0pQ2JTwo7awf1MPo6LSCx5axoUbYnjxNPcnNZRgXo+twYr9Ivj41ld0U
163R3dF8+jOF9XdVuYYZJ031kJMPJShuoUn98wOizi82iNP2x+1P/mljYA8/yq1olNcysYzuVAHo
iXvebLsOG/SguiPhaKFz0JLuJaLB/otw50kEkxbAeV8zC1K9t6nk7rN0KHvA1M0bKNySHRfUTajB
nGSOkLAXa/Mb17ZGIcqlEKgzVrzTnHOIa7WWVrt6FwEzDTdgJBkbSSjrUdscn2qGvqKLpY2trX+w
vloqapWD8u2yJDv50dx6kd0YZ521Zb0almcZdiMli/Fdcg6dDjeWN37l0ell6CLKR6KpaPMfxIvF
qzQ9k9Pp31YfbUBUUU5r8fSCcas/SkBCPu3x6fmJ8v3koal+8gQjxatmyNvwUghg5sPmZo+4CDO2
b0ViTJESUEaWJM8+0FyYr3L4cbP1i8je5dRRgAGx01C9b8aIrJpXqGl1T9sVYsqy1IvjHVx26jGq
UOblJUzmkVnFi8BYnGrwnqUKoVUCJ9WKvq6Jx3gfu+rwJf+6vVuwjJKfjVpj8NFz7Fk2xyIlORlr
+NfpRf7iPzZvpxC5a0bzqhC5r4bXyttXTKgSzIaZ2icqJlYvIudHxqTLJ991c/MLVdI/O/yzN9/H
4eENwatuyyRp8xT1iLskVniL9mAOqcrPaejQgt6vHPvG6mQF/iO/O7MjurhrwtPzgCx3/t8cn9VM
2sMDb/hNsH1q3Kck8pdAbm4IiVoitxB0GIGJYh+Dnw2CZS30W0JOtHq1T0idCN2WlnEIjmzjqN8+
czKFayPY+0dhs+qpfQpsH/EUCZFuCCr5lYBnJ6RhLb+MwhyXkMSnJE+aV0e1OMW0mUOIYpUrTyP6
KWka5bmf/aH8nnf8uKepk2+wWgu7nPm+vjW6CaIvRxnFqxW7Ss7ymGi53FgPBEJTBPriNQ7r3HMx
F+1gRq/hPhdH0KxrRubtZfzxaVAScsVa8rKdnAR0CmIcrmyQxPpes07IezzeAzPDN110SKQcmj1H
2UGpcov0LkHJ3Ynfjm/KPKLT97jEl3PPil2+IZHRsjKJ3M8CI5+LzfR74V8CfIYKVw/vupis6KJu
CDeyBqPx+oY/LZGoY17h3doCY6mLilncCjK0KdxJqxZ0yrynu8wr/U2bZg7q/Mk4f1W3iJDKeOPL
OcvWGFMhDqjds4t2pBxq2b83NZYWV7FFVxIGjEScDKSe+CBhZocCZZ5q0VqcwIBXg8kpyRwucuvO
9OFPK0ck4b7gLY5vhEw+muXk0fEBJOnScOaq8hUpC4bKhBEyJIRyC4gAReJmZ5aXSKCnYw0IioS4
34UyCiR6dZKoCQLC9R4ifOi0AUn7EzkNmxx8g/ybmoPhQcouqB7pLk9iY4tNuAmdgJ5sZm70EM27
4DEVbV/2ogACRPsrM3NTblNAhKt8akvSRtaZPrylaTYR1HrWqxgiccd+P5iY8O8W9/h8LQtgREDA
pEj00xXxSfYyUMIADPryodxMcIckV252HMPQkRVqYH8W5Nw6NFu6OZeIOi7ZOy4NFKBul+LJKbyB
GojjpQy13T1UbgJmWE/ynP7w24lq7u0HG7pcrxUtdY6nXqWDxi9Nz8wjaoQXSWScaLTR0yja1UZk
eR5ldCnQWBp5Acgm4EvZKwDsJSVCUTui4aR3jBvdpsOy3E/G6T93gZnx17kYnBfel+dc9iV+pM26
eY/Kqb93/46XZ4ADaup0YB7Ema60GEFd5nwkp1osBJY3K+rbFC+SR6WcaaOdLjMeOKoCWMPQph1A
lpImG+HthCWjWYVEG0hcKMC/CEwbYek0TpFXkNXdn+dBQXUXZVibDI5sBGJxftyExEO4gDIpQTE1
Tr1G/W6K7o46hvfrW58Is+OG9LArbncfQL40M27sLbjlnmM65n6y9fFBoJCe6NwUwLCPQkLo581O
Iuq6Bs5HUkKFdu5xqjx8A9kMrLNVlzYbS6HPasNB9+xPjcRdf8kxG5Ce3QGg+4x2Bjgf9a8ayYlX
vB9FrNlMfQrpPYtP4neN9+h3k0bDgYuqU0azMNfed27HvY1B3rk/gVagnI8Aj7BiosqvKCAqt7rf
7a2CoZ6bkCk8U+PtH138YRFcYLWuGEl/OCggS6IeNMRwdw0D6/Fnl20RLo1SzzJMMk8OvsppXE0G
aQP8Rn8LY76stfmgwvzgwUny7WdIR5aJ+Oq9/UohTjfyQU338wYNVqwx+TpTQd7LJej8cl8cb/p2
TxKxkUcL27zJyuFHPdx5r/lxQAKr0H4uF/bSrldeppc84iCDA0ISoK8w/dt+EMxFxnhPraRfjNHY
RRJ/+KidDE3ZCsikj90xV5pzkagxgehML7RLRzSF0p4dnDVxd4bLd2LvEWiwHPltPpUbbjbH1dMD
NcprgH1TX30VDiwE1R0XLVlHiQeqUu4xD1EYSWGXJifOKrksH9J8nGsbjHTYOuc3NtkjLHp/cg==
`protect end_protected
