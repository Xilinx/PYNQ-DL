`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner="Xilinx"
`protect key_method="rsa"
`protect key_keyname="xilinxt_2017_05"
`protect key_block
DNTBN2yRu2sIJqe9wfMnsUORX47AqReIqzLkLKNVfjtioXHPdozxI/cS7zIGkAvqghsq61l0kF6c
kVTktHGV/ryyabraT+yb26sa5e+jwu6WhkZMByIgqhC2HM+F6H2fGFZpmV8/QQv+ARrVv2lTS0G3
niRA36fTaOmzW/PKIMG7hdIFri0d4elnY/ge8N6QTkzht1Vx/G5Y2WljWjRIu1kRwAY07zgtyssp
jS1vcEHZdIAyvBGmvN7Rd+CscUMgeJ1VtaM2zJLM82t25RrSY4lEo5PNdCbcuzriFgM/9XFe/fT+
cLQ3xpRVQ7nizXD/RENQA2qahLkzCH+zN1I0JA==

`protect control xilinx_enable_probing="false"
`protect control xilinx_enable_bitstream="true"
`protect control xilinx_enable_netlist_export="false"
`protect control xilinx_enable_modification="false"
`protect control xilinx_configuration_visible="false"
`protect rights_digest_method="sha256"
`protect end_toolblock="an2GZCy8s9TvJ/9c7oDoHkG4Wd1kHkLw+lkVL8mr71A="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 46768)
`protect data_block
vTOv9dmJOkIAdvr7PjKtuG/C1rH+gbk6bpmvlDOx0UEzfx7Hm/kVmLh0r/e8qjxPwlNqPBwzlhVM
2LN4AaEpkY7PeE0mpGxf48LBDjwnY7HH723xY6I/FCc3KdRjz0T/LZ/yuvS6kb0bt5cCbUhCSfGx
4dDPjCvaANF641CoMcxVdPbgpE2tQI/UCmqA74frFvRn8R/rtkEllSiavtgeO2mVz/BOfuKRMMkp
eLc+5T9e086byfuugKzqi5zwwiuar3I7zLuku0++iBqu8fTJBT4ZEKrF7iKuS5DHHEJQEI7+JL+K
IQQ62hRLEBG2SZ8cdSeMngkAivB48dtvd7XzLz9PiMOVOYYUOZlIss1+NlYqfFlolSBPfmx3BQZT
OVC1ydNsTuGATqisSAtfDeauuqguIdeLYcF3kGu3AHubC6Rz+91OCWdHwwTdwKvAXmwx8ZVJuVCw
Uk6UoD6gJYf2mD1B3vuzeQgqWDdaRY52P/TNYS8E807sN++R0/M+ofhZaGSbZV4b+zlqVF4nxDJ7
B5BYbw00ByIIQ4tPkiCYS0LRcd6kgm3TEWAjXD0JPAgAXxgREPJi2uBTKStGVUfIEeKDRKhzKkgg
/irY/kFcTluCpKG/5wRpzjbknXHxtu21wA3o2gsIn0itBygWI5U3hTj5F/ovmjM1M+ayPQP/vQKW
zir3qF9vM2m53h3bqmRy3dnTL5hB7UBjru7H6ylTM5WsJscyZhUgCmHRoN0e1ZZYUfp5wdtQXh3l
s0eaS/8rQ2LREDbdbcjUs71iSt00SjWv/FY8OF5400uylfKv4ktzYWoH55XVAfgiUfigAlU6PrLD
Dn4/X4sp71obdnB8PY2F+yHkWfXratwR9SK6+trBYV8VBkjdOTADjrs1S9i4+CKT/SLxXjUkpecH
wgUKyafG2koyzLLZrh1pbkolBEGA2s2aqZb1RDBw5FtQJuuh5B+ioTtGXpVEEj+47/hQq5lU0ZII
8/9czf38S75s0YT7cNh3Tu4irPSz4h+wO0Ls5swGIlx7ObvPVC0nZ/zjXWXoZeETVTspvKAJQVLN
8mxjrSJMkT90tKjeFEkNHsHS4HUjnhIOZVOQw7aFnMijRD+D5x/XlbStwIqcX9Fwh4U2p+zZx8xf
uKKNbT1RwuncKyhULiCDtWwjfiUf1pcu0iF5FUOZJSd6R6EI+7cEY0RrvrZ1HeI6MCzCQHEbgtwa
7mBuyR21cxECDGlvIVJ4BBBynkKcJxc+kHUSaOWFqQwYNfCNKhrs4CrBQ1dOFez3d7HaAj5zE38z
XP9weiP2mcIzivqPuYUJAiVSBUsrcksg8vCDZH4fpys+ldnDJF4O/Vk3BS9l06jpio/rHHi1a5le
JW1mudk0C+W0pEWlmIyVIeAW/qGXgnsu5YncPzauW1dRupNHccM8TblptADwMTPefCRoyuj6kVb8
xhmY0C6JWdnX6sVqNIcIlrpBjj8fGSWX6KOGj01TMKWyFE4IlklhQWotVNPxbvZSjcxzseW+XWlS
2CSbipi3XokH3YqLZS8E7YpAXWfGaZ4XeNl8kF5jFj+H0gCZKhjC+ybobcGnk5MM7WcZQ7ndsxta
lTf1/lHR/yX/1Kc5x1UiPxWUsPtb8yjI17KD8dKCGMm6qX64sJgcWGayh/Vx7DvxZPxEwb+J2jI+
C1Bk+ehol6NUbZjyKv1AifQI2EosPUJ/hmSLVnoMnLbQEDf4At+7+hhrb7rCXDpRGDTlRtMPBslW
Iv2dxgSewb2ICWcQ586XftOJS1eL8jlWiAlgP9JH2f3XLxAl+VopPFlZ3SOQ+Y8a7Zf+nNPgUelD
ZeGDHuLQdgKiXlA8flS4GQoDFe780BJ1uUS72BE+59HQV24Cu9hRvxyp0b9AjxmR05GE0covJNKY
X4wevM1QpsXAEFSRx6rdl93jn0NJtWA6rUYucqUc/fj9rYVUnpt16q4Qt9TureeuxZf3Z55qiMAJ
KIMSNJb9gPxx9Dh25ZDcV5+9fgLo63Nda2yt6IeJrAWx8W4OlncF8nCs09+7jPyIhbS0KELzramY
rVI+WTKr9ovQ1+RwQgTrTSsWTeOLgNb/1Q9jlht8gNodx8jbC+MM5NVxMAOjRpR4EsWILYU3aGmB
KaxVCarKSm6kEzF/5nUqRzSnudLnPtr4a3G27TAtOQ30e6WO5BIgCBI0ZRux+dfUpzVEoWtsTIJ6
XBMUbtLFy+lLeK/iw8KkE8I5MlFr4Pdbim3zWLOkG0Do16c92EhMQYFQrafOqUlViZVLrtsX4xUF
cdgccZ9JXto2JWalI8onRQoUJ9Dri56at7CpC8S+6jmMwYojBFY16mpMK35qU4u7zXvYg3I0FUGH
BKp+n4gHdu62r2OnlNB894SMW49pagYUZ3+mFZUhHb/PW3sd0O/RqtYdO5c/bmp8rQTH3hgEwVuE
NCWTVZ706wYK+vAGwDywXCaugeRU2AXqgrEBPb1ZNZDVvz/mkw60QyZKihlevG7gj6ib8nPjhtBt
rOR/DahIz/dDFMamJXanYurJMkFj0yNSS9Da8ebgz4ClXl4vUBzXJ2mfx5I0rHyMM51ujw5EzQpt
J60CDWY1U0c6wK/7qObrKeTKh/JCMCbSrm3f+6mkGRQVmE1LvEs2euz0fQcIz2JcTkYP3VdLMU99
O1/6ug00VSQNWr1rCioTG4KkhNtsopKyeHmfYWQDXtFt8cLWkOboQZBmvmN+RLTdLEdnGK3eSl43
2TyiF8iuJsvVe+HCEaN762TNhXe9Nu2TSAB8C0xf9FD+FoMOzMiqJqKXF6XiruEo3+xo8tS8yM3W
KI+wSfxxqjMuEYi6QfdCwqKfbOoyercUuaxSlnjr2349S43FLfZuVuBnIKcXa1xaJ1JEyjnnWBX/
e9Jr9LN2qi4gZF2ZgA9XIIG0ERdSjKQcOI2437jvSWBTrmpiEoXWv/b4UBmobX0+3bOdw488Nxzl
/XKsVyF9ZAXu/8deGv7Y6KnYXftv/3Ee7UwAyXewLBYI+gMLg6IHsECosdW8dYrF+dcVnYveUCeC
TFscbSAxOwSH2jpGU8Wz3/+wYpJOzO9aXYpFpELmYii2+BOBJbMR5sO4SPjQP0Vi14m7Scpx11wQ
S/cvTKGm0iyGDNlOJ6kcYL/Jm5abV2ew6D0mlXPICUwHanfRnJlEuT3oh2lmruVCGkgw3VFiaza0
I4E03HDNguzxfJ6gg+FpQUFTC4LdcqjAc9LF9sR3yq6iB/golnEmFm3F47r8J3WdkADUQ6TjKmi3
m1wP67vYDvW4AWTnxf0XxF5TB9u+UoMon8A08kdqvY+w2L/LxYKApapMkyZGqHz+QhYbPceVE4sh
vB2+4AYz8+1NupgKIDlDYMFPrWmSxh6KtoYhxRP2fCX4Gc8UsV+cg701kJJ584bJzyTO0vXUFKgq
TU84CIQpf/ZSHB+lBuMZOxB9B72PqrjQw6C2Rrtl3Wxtvb/uyFagnCc0gswD0OG1Tgit2fPDn/6/
qfN5iqC/2mSTnlmdQ7kSPelpYYtcwg2SKp/AtHWAkKIWmGnnl042iN3oY54E8X8cvCHB91UqbjlK
WraKQNQGBtNh1LX5OvLmfh2dNJa1YTqw3cpi2KMl+vxUEhIA4An8JfHCFNcW0g0NlDSmDjaq5NNB
6fQYZevbqfVhKPvCBg6wTa6Kx/pkP+w43up8qG+lIBX+tyLgQQqoDO2k6QJyrFwMk57FV88EZ4e+
3eDbwdh8Tejmpgubs7S9Mg+5d1Wl24M3aGypyFDkGqiKenw74CwXcG9x3FkWovU1ALkzhMqjVmCS
I28zZmPm29bGMYdT9CAXin13cqzI9koLTOQiLpYOdUWSWJLbz11I/Q4/RNDE6/6LsWt4k2QT/giE
ZruXvASn/sRhFT9spqw+5gh5gyVOJz0OPDIbU7rS9tB5H+03K9ac6HirWJl1IGnAn5AvDIqxyqPs
WTrjeG9KZIi+YBPKHweBKEsw7pPA8HSkJwKgcEdfHqcrFmMhyWBikogSHbCYfRjmpswuUZymEGAm
tNdbKej+9UW0AJoOl7fi5BjvMjUrH2a/nEK47SShVov5Reov+SzjSQqm1MoVJ24a6wz9vDGrwbvs
+DvszM8J9cPQLn2q0txjCK6uO5Yug57TGnELfo+GYTDzKjG7jLBHZxxDgtBI7z3objwrxQQyrF5p
Xw8jJn4+uWUa6ijs5fUJ3L1oYrbKXwh0XN8n3cgxQ8aY2Ctx5X86tBdWy5ZW0mJuKXuOgzRB0PLH
RE9iYXh7zh81jPvbXq94NetpM+xVeWrX4592unbcTCPuKE09LrNtKxZOzMfoUkgi5+jLFL7C4RbL
UJYbOU4tfip5sVEBy/n9qFeIdZd/OLgklBgskud2/MAGWF9tzYrmRnK75+nZNI43ww39iC5orQl1
PkllnSWJl9gYnhcjhvDxlB+tIR6+Gu9q2oFa6ajFOdEIxbXO5ix3+JY0CLspkWvgA6uzqU2oyHU6
EbWMh14T+WaYUUw2EBARQYG9MlfP9dOpPvsC8RZttMQtcJY/4kpYu61GfLoWkyFmDp4Py4UK75z8
S+O6+ZhvH3ZZadYJcu6uPmUm/Zvc3nlVxyg6p4pYoc9uqpLrisLFxTpxVb3wFIZ5bQf1xgxAGiXb
oLc9GzFnw1iIk+qEa99Hd7YfcEvtePp0PSswrWPd7LFz0oSidC3QoDMu7tfjmo2FgqDICkJY0ETV
dfdUDXsnZjUynIDLweDbV8ZQ9p5VW4UwyNTR6CR6mUsyD4W6JlRaP1bauMw2eqLOI4xHNWSPbPfn
MSKc9DS0WFxL5SXBMnWkVVy/cqfNq7ifHEw63MihDcxnXfVkUuxobm8FgE6QRI3Io/hy+gLYGYdZ
fieP8lpPcmOl9hsU94z1jCUoN0F5Jfm/AVABPCQ4qmly/k2FEVfVKgSABTZNi/ZanUTmVe8Uzpyz
/8Nnog0z1PlYyEz4wKFQNLC2qK9EK3rjpwaUbfm5CAZu7yftzKhKPVnJfJD3IxjpAZOZV/1ghoyc
sw/dQDJdvXXlRojlrtZ9f1xpSn972CGIhDtndhJKAMnoEOfsbPNfA/kEvu5gAmAXtLpo0PSkItv3
y3tpcq7pC4FGt/YuMeun1wX8qkSesozS9lTg5RvZu0F1jOwUewXaF/8Dfmggy8nwSCn+JmQ8zRMP
snHunwUp6mscGrTwgeNUaeT5lTg92iXEVlbpX0MkEtmcXgH7xJqg66w/mq17/q199pYZvPWagR+B
z8JXfLPGgSx+qY4UA0Q2ublVBWZ8eKYxPB+hxJMNE0IgiOV48DChMreqwDVOHa9jnl2J9ca9CpjP
QB8aXbnTmPpYNCIlT+XMZCYEBbxPdKU1tnvQqmLcIDpAm+SKT0HnNZT0GQtLOT6wQGFvftRMqLVa
VdXSyjDgu466EU+um8p35cXIorfZHEvN6STxlg5r08KlQ0os5U0rs0Vfrth324y2l4iRnl2im8af
UPrAk/ZK6RG/+jNLAoadY7PHdWkzUpOV6cVifBbNSsz72AxUFgqR7sbiuJuZpVj0yvLdO2zLPQp0
y9xW0d6UzKMy4iyxJJwUqkjoayCZAZHp5DNxDXry4DYQIq4RZJJgSqElisbpLp5KMjUpTB+RNBJ7
3rb0HLws/sxl39hRIl2XQMsEHKzhzu3swzRXIj/ZsbaEhKXfwRT5Xk6lOBviFYzCbMkvSlg9Nyom
/Jb3JsDP9kVfiwsx/cY18kqaO7ajA7UqcmdimACw9YAVjO6/jl+zlG8lmitmSFDnKRMYzo5qTa2S
Kn0raEEAtdQBnvUbJjdkTjNphQmSNgx9lKKUbcjqKikX1XnsP/U89UczhfgBJ9Hvvbiacz/3bSO8
nZtSxmrdll/QSlyu6A88tfjQ6Mnf74xfqc4n9ZKp7M4Pmd3aVjW+/RR3NFXRAkX4FnRecxmsXld3
Ldl2hkyHucGenoQuZcM7/zKHpQvNkPPnZH2varDkSZAnK9IGISLw4GqZw850QogutQNo+TcPAywR
enkn9unyb8FHNcfl/C/Uga8dCgpF72HQQn5d6VKbdGSuMjtppMxLqNaTnh908NPN8PSANOlkqD3Y
PvDZ4FU0rgvBVQ23KYlHZO5D9rHGEQN55BmvudIF0lgNg4OYeZ4mjg8VhzBwAdgXSXor3UuSdIl6
auIdSeULjDDxNiQLg5XJEzp8EMQV95P6q+65DLhnC3w4c4Rz6j0BS6ocZzFHUFxR9g75cRZ1lHUg
1FpB/ovTZGguJAtyQntFVc8M0vUzpUDaE9e2prCnFS9zbMdYVcLYv7kD6qEs6LI3eOZQpVTh0XXu
OZhGPW/YyUS9hx2qWmwDHMiPFChh/MngDiOjJWaUVDzYgOALKr/VX/405rUKMBHUIAykN06SRI1y
uuHRs5aG1KdOWCgH8ZM+cUsAeLWVNoWf25pNqenuFuw6ZcTGxJqgeXvcsm33T2WpaEwi3XsmVeyi
qg6nukext2VgSB4Bv31sgKowx+DGijrvEArGUKGwQRVTsmCPl5164hXAiIQotej/PKs8DUf33W9R
Q10qmqhyFHTCzyhpvVn3sUEO2lstO5jRc0r+1stmF9+EWoeH8F+IisgcEsAN5N/d0xsG7OvDV9uY
m3dJyNPJL9AKy49de9HEY9bodHeu+p57EpPeYeNrHf4tEYh2d58waXk4IlHE9C7oHtg0h3MogF8J
5Qg5XYJjGxCuN6BkM8UF+lLyFUeiXYEW9Vgt7lfbZEoTjvqorAUR/ODTLSnMrh7QokUgbDTz11ev
WIdekUAcmQF+QmpkVEPO5a6sMf1zghm11oV4G386+cyeLd7WsE7Ikc3mT4HWWruWs7sZgeyqpj1W
+zicUb/2mMePOksm7k4evgxiPipY9Wa1xr03QGDrKbQB4Ken5+oI+r1bKGN1nfcufI5HjhOskt3z
YHTUkHYj0AkPbzknX2+28gnJIc/zK9DWvTYN2a//qKqnn+QGlw3bqFKdZuNGmLnv5nOA/XnQTj1i
S06n3B8EzNdt0eOKYwwivGQ5K9E7LrhoAkaxXWiaPCvkmtrV81f+7STMoXE1suLl1CHLl897XE35
dEM7lP8n02nm79BBOBBPkIm0eKlN73ZRQn+cDC0rBoSi2PBZt9YLaHL8+iY2v3a2ELjlvQqCicRz
MwLUT3A4grSTxudkCBUcvBn/jKNTU0uStjdw7L3WKAbYaXyM9G3ldFIFdlznp6nDnkpxEjmR1zte
ur87Mm7DJtX0G80+bkvc4gTu7HClQT83MS8ZTOlf+nBbFQqeSTt/93N4ArhBQ9RSpOdZFyLIku27
MCjzPhQEFb+pt4AmQph5+ozBDDRKqFQ78X2v5FD1IRGpcrFcmgP/MkVsMUfsaqGBX1BIjXEl3CKV
Buv0f1MPnjG63nJctX+280puSRMS6NIncWw9svzX1q4kZEi2tHOQsTnfFemgC1FosPEArvaYlnbS
wTElZic0zQjRoui/EqOSxGGRynSQhEw4Ky4xKpH9iaMwzf/nhry8GSrg5mh1FgkNqQLHVpFfsyBD
MVC9aRzJjoP6dfmjbBDAp9ReRQLD6BFt60YwTy7Ae/RWQwRgUdjNH+Yf75yN+4G5ZX7dY9Mwe448
R9A2XhDa/yQEuQ33CnqsOuhFjfnYgS+40b/Hik6sOydj75K9Df0f3erlb5WMa6aMPwkMYEDGSG1U
5sXiy5dFI6So8iuNcUs90iAW6eGgzcjvIDxJK9lKD/0+wPVjcD8LZPZqLmSlMr2wgAd9JcXsNj8H
so+fI/S8LvL3Zg7wpZKJZJBBZmkFw5e3pTFiuNQ3zTuVa62NbUVbHcPPnbPGG5f3Q4EXGSd7J7Mg
agpc2eJguunbQmx0n/nzdJ4mBRCXj1QWRxliGQD0y0LbG1qkM1Gjzkjahs7tE60oJ8HtfcxP3feP
vaHAZpGzxh/Ttj3igYLYD9f0//P5iQTXSyfPevHuug3nIaOpnqyYIYcLN413ByhB2CRI3wNzxLSf
D/oqwMC0F1b7VqZP2ODxIFVLIxuv8AH4Df3SbHcCtCelogtt8ECKM1bsnq6ChoNgxVDRu0hqG1Eh
woPY7VI9w7kkbqtOXWY2pO2cDxgV0TOoHZHpBgRBRzbGauvtbtcCCWqnw5NsGY0cHFQMmiU/+/A+
3HoS8+bCfKDWMjz6nzT7B+1wvHAfsSo9UysmaVS0VW8zAghUl4V1j12CEeFWCfifHmciYjxLw7Rs
AqeM02WQ6+lc49IUECYTqOnlyCHcPRMPEZmz8S+xezV0dc/1PyCwUheFeL6XeKoz7y/XeLNr1hbP
csW6yOW7e7ZS1hmO0GnJ+/bIwUr57tyVfdP08Sdc9PLTQ/7I6ZQOkAguSaUt//a+LFF70iyR/yOs
nRvIPgqEdhvBANy4jCKSMJC0UrmFlJYArsWrUNk5CYWLtY5dJ8cnb7vZC06kfroxWdjXkhDmPd/D
98z0SnF/WODRMJrDJlraR+wqLVSFX/+VPvjh1EXrnNQG6gik+pxHubw6+tkLRkzWio7PqQ8eAUlU
OCP4UWIGZHGjJ1hG3LwsUpzu5ZEgEkX3hSJGvj0f28VtDyb7x9N4Zs2hh8vja3QyONGVxqZkKmex
uJPXdenPw5e9+3wnVfDyPvvAtS03/SARz3m/D07KJHBOnKXoZ8EmkgSps3kskALLWmo2Gh25/s+K
KXXoPLa38fhBtNNQNfRoTDQwoUBdakz8csAY1QBQ8xz/kgFTS4OcqKoeX7SuNjOpqNxHCreg0Lff
fF6wDcea9pT7lcd6nkbPUQVYnYNLzpenZReVYRZxVQ/3r9/5CtyVk8qBQl3aYpo8ebiuxIZOcS4o
dxjZz9FqQn+5DMmcXyVr9cVRdFPLgiPqWvXOKwWw03DuSs9jZvRPJOj0talGSAoFG4swR8h6Sg2K
m/elwChZKQnacPM8l/3pXeHFGdORQ4xwssC1fvTRu5dlv0tfbmI8R0KZkHq+CIVf+X/lF8O09QaS
VJHzaxVweH+148UIEea+/JMQ73JSQr3aVNLlYnVHbiadW69krXzlGQaK4hd5a4/WuMTXSRgFBDU+
oQGVvDjLOuKs3QzaRdzpIpZ8TIQy8LjIO/gk5LrHw45RC28+IgmB13U1raTn8eB55I9w5x3mceDQ
wUuTc0jV3I6bV4t312ciXOJDNVnar4GYyZkLn+BQ8ml1jzjd2YUYWvvaF6AHyQNCSY/0eJop5J52
bDW44CHOE7sFchgIG9AQdwkWg9fMYsg96X/L4PaE5cxfl7h80+zElbermkG0L+rU93yIWsXOAuRT
1JGog5BgMVmffs0H6JM6Y5j5Wq371TX2MAgq46EJSmaAefywpjZIu7wmGgmxp9hxo5aepTLp1JyF
T4JpAk8nOMOnSp+wRlOpA1ZMfEUzyktznDaNl4QQo2FJJc9f3aM1rYtLicHR+otdjuqlcGTzv3DL
GVCRlxm4BLiA+nT3NtOjs3uEzUCX6WmInjf8TINqe4jwAcI6LY5CSscWdRo0tg5coBn6aLih5yJF
vHcppEsbznOdRNZYzhJsd1oVh0QFeQI5ekk8xomcX4fS0EMa+Eaa8L4UtKHwFLz2wq/Lt1spdIC8
ppTtv3t4nWJFsGjNTIECeItRev6vKYj9ZzTjozapk6OmRo5pDQxm7UuXzpA8Ev4GvuTVswK/HaAc
inyNQeC7KHnX3nJuGS3gcKJhYnV/NQzWAvvkA+Icm+Z8NBQwIarXRXm+XscjEncyKyPxsg9tMrp4
CyLm/wcUZG06QV/JyyTH1eiWxDyMz+H9XIwIyjpO2Xfle6UneqJyvai/Lt9EbTKM83dBFUkO54Pk
Su1qQSdradaulATu1IksESp2HbcC+g8MZsseMyuJf6j2azxhTERgRJ4Bvxqlo57PpzhvOGhhKUNw
JEF++JAB2j/EMJlB79A3mpwpXkXebJt56L1i4/wZfdHoryZl4vKDlGM7rJ47c7Q+5S3F8jcdYO7m
sH5y8pV8IlL/l1ao94ykn/JL8oq4GJfcj3PrTicvNGrw2rie+ClKbvgWQ1aIoS8gyt1CXMgpPf2h
0nJ7Hx1lKMQ26ni53WM9g3dSXOEOzfrhxcQT2lZKpJYIARGpjskByPTneAtfVEFC5gPjgwx6ds6W
VjO/Czn5p95uudpT4iaczfsbXbZIunsr8FlRs4kBRqSyuwIZN+semRGfD8ZQ5PgQ3/FOjh9Bmvd5
B2YL60vfBehvyV8nMbmNCdo1op7mlrr25aOdxjsWEwDTYALbFBWeSgHX79m2VgTazUQQZLukVmCg
/15j8WcyebHR1UfmS4D2in4PN6hgD2+OQqvP2x8K6kcxxg53G3raMDWTafPMR3UI0lPEiMxCWUTt
OsRbPQ7EeN1xKib9QKSCJ1dfTyAdtgQ6sEEq0hViDJC86a19xUjtsYLxPw2UzxOhuD4TRhfs0BkP
rv2gveKsXfFjZqir9/edqAD6LH0nYHB0BpzR9lHCEN2OE9+JEVJny6+m1ZqMsI5/B3dG5yM96rqW
SrDDNchbacJxk7RGD2/Cd0yywVIsjMm59Ab4HB9OJSdi67JfZXxZhIb/J87GzsESC4zZoXv8aW+g
wz/9G3gAyHVJcBo76ILthbjsfV71LaC2MyIeDjW3DCMemjlvlHjWn6VTH6MaENACba6FJISO7/+f
m+ulWfwoGDSl6byy3W/1ivdW3FEXB7KzvmZgfr72TxiLOWcmdcfLJ6ei0wXabmgLg04oSMFU9fhr
C2/rwF4dGGz8YDlX+kveq5UrHwDskvGStHvkgwb5Chv92qMYfxN0J1mhvG1MF7kZYmXhySFUXs0y
X+DDzna/J9+eN2zj/rRXXVpKJFislEgtwIUutK3IYqpI8zZEo6fcmUOsS4UlQl7O2Z6Pld2thmtR
4dhTxc37WLPdnGgIzBpx0lnC+Q+Vrwt97z/hcGfL+N1dt81wNzLGyTdYzvMSXU49wWVmEHD39V1K
hcW+zWxB0tjuSEvYuCUd2GVw9KCYWQ9b0l7oq+Q7LdoWkpSvNaFc+w0x7V9Vm2FY28Bc39a0Qn1H
Cmrkv4nKmWPNBdJnXoi7sHWLI0pTYgxaSQS4O4QRGoBItUWZWTQUNklC+YqCtnhn1iSHOMqx7UWB
awOT2oL2RhwYpVbKjF+lhY3XWjAD1sop8D5S43g4eey+A3q4nSuN19zya7blJUWOr5Zptyz8JfwW
sGWbyd1BbELf5TRU3iaRqCzyGz5tuL0diNwAwjIYkpPSC+/AcJJn0tobhGLtXT5ejTRcS0/B1tSF
ONNX0Qzon2YeMcEFbhOJvULIk3kuoUKTtxAWx9oBQPHlM+atKvAVrtPLvlWSJN8Cf41J4OufBMPz
HZIfaLqcQ+kQO1Rn6o9Sz+cvdoRCR6eL5LFP9R90fNNbnxjho9XvFg9N/NuWPZjZoGGlLJ42h0lb
hyjwy7sKQUre3ET1ndXsdbZwx1WUqOCVbkUMXc6+WizjfRm6WfQ5ntxse35VOnWVsnIkJzqdVDx7
kzzv02/14OcuQYnIy5VWEt+QIj4SLDujn8MfwvTMFPuBJpeZB3w1+oKfR3XF2Bm2jHqM4Ecbfyh9
1G1W3T/TEMSW10wxVFNf+dfDC9Kj7ebl36+51EqvfEcwBgODJd+VKx6DF6CLW3Jk6WJ4WTMw0T19
fObuRM0OxFJPYS3Xv67KLWOgsWObSaGXEVOVuYL+kUpetXOSWmmMWjuf+KkIVxgUryJJBHUNMIsC
CPWEESDB7xLtg/LV19RZiYGndb2H5U3G6gI4YpxuDUrmFTs8VKFE+vKkcvMyPdcFdOOY/tvIZQbv
w0GK46N2wUOaU1rCi+/eL2qfNm9C/hI1GS6ES2tpCjILL+ZbTdiW/PxoKAkk6KW2YvzwkKmn3Jut
GWIAu8ASfZojOIHAM15J2QGxsXfrGONYPNQHw6WMtO5FbFiaN/+v7vlogj3wrra9skTPvZ95GbU9
MDpSVgAidR5z0kHKFC1SpwRHth2i9CnYtsvAQN5Dt4zcqPTAhKBF4GsNe9srlTMmVqAuH424bqc5
xbJvPdOcHG78Te3sVh2GUXEhHQwxvltkthDWkT+Qefu7QLVSAv1zNOaMj+2dn6AhDwkpx/t66OyB
SAdTwEAIqlf3+aKS6pJLsTeFdfntmQYwt9F1oie5LkTbuqCjEzjPmWOGMwHeP9t+5VrGo3oRIbdz
gKhPEtOsOa4oDIrHf1VRNvDGccDSkfVWLUQE++vfezWt+LBJc9886FohrD+zgr4/Hol1UzmWzfXm
jD2ktqw+51F9OkDyOs47YXnlqI+eJdTtuZTB7TjCpCfJyUMkNaC3sp1Tq0B/NBt6tchiXz0LyQbe
8AUeqMS+g3WTu66tcz9XMCfldXcuMJsk0U06CWy5oQ9JENfhNVLPEhn/sKbhhrCtX61pqtr0y0Lh
IgjoYMWcy9mG+B0+bgKV4pg1OhfsZey/3sHlgrIhZvZxXGK4Csd42kX0vEk1zD1qjk8M2TACaNAi
GYT7zGU5nbVnk1SZ+0c7YtTsE/367cGvlUwd+T30NfUpxzvb/Bc3wZu9WRR7H0oghqBHJmtyK8um
NhuIo1oCfbD/DO/1YuCLbZruh4QREB7a6vwjyLfekSDhWIACRZcmCfT3HMH2rLVMC/kLaG1MVSwY
/CdauwFVOvI7YSqx/OSsdwHjgfUL7YIs4qQY0jElAu01ghjBIOIO0IIvbffRTLsWb52+IiRYp4a0
0/pApw8nLxMsPCazqPlbXAQBU8NRh4cjAquH1grGF2IqztFiSp2VtJwQD1Q1vLLBqonK9RkFaKOE
M6VVAEiVmbdPO0js+xs4TLDA1PnoGazJhRb9O+AeO9c6Qv3z7nhzxBzbMqjp99MgHHRusLTnQM2q
L7z9IF01V1nDC3HTz03tyLB6DHVNSropanARAGLYAAy0aoHbv2qXABqWxu3rJvjbnREDR/SKTuko
cJas1qXbStJh04L+ausuibsV2C/HHRU+miZuN65qjjjxgod2FiC4J1G+9JH1EvhMKE9sjqX8Yxhp
5lXaKYZQig2GC1eWctV/c2FBZSTe10CFKeqAdXBgfnYT7okqyutklNUQs7Q5aZruq2oqRtYdP5Vc
gykXemaNzdVVwQdjSbYuQM5+pLXrHUflIFq/16Kuke/NVQT/t7mfgalq4eFS+XVNIo2XzeKnOSF6
7/2bLWEvNuFr7MpvE7RsBPsvV57GK1LrXVeSSgDvPN/slpnNpohVLHFz7Ewtn/YfOjDfEuKGhK/u
vfn7d7O/LvNTUZRfug2DUcXNow7K7/Sq/myQEi3sZH7UJrw+qjFrJvESyfnwAEWj2vgLEfFEYfMa
bivTAiLTdPPMlMHmwspndI1qmusV4TL37kC7Vx5IEZ4coAQ8YB2Mxbj9eUVw0QUPWkBiwFRP4DcM
QK86TaA4oNvsbL7GgcUU9kW2777IX5khZ5U+LQ4QDQgFThS9Ulwl4AlL+RldSxSYevOazGqUfkF3
eddWjaWD7gNK+/Tf+uUMG+6N7vLTXWJZfyVI+I+GHolS36dAjSZXyQGtJ3EWHAwi/FXEbHSC77Ww
IusnqniNXFPf+HM/F3UvPaEHMUacEMSGAHEtsojcL9NS3iTCbbNWpKuNV/wBnT95iwhQRoUZVYW3
Wb4lLR6zx1n2ZwdyA7kuHxcWVEC16IbjUesQNY+gMILO5om1HeKddm7uivPWgyOOJxz3+370VRJa
jBvzeDbb9G3Lay4IoBq5iGchcQaZwZV1y8bWQhDkf4KVBxVpO+GEs8N82cbC+558UGZGsJGBoSX1
45kubwrbKLDAimlE7hmX7ozZ0rJNsrM0l2B4HXtPTm3Y5hRdyA0vFrOLAAAHw2794DDvxhwYGwGy
hQu/qpBmHiPSskdxlvVNlrcbzPjEZ7ZyV2yMn11z6lF5VmvsOhyDu1iA5UFGplNbz1BbkGtlSTGK
XnevpFCOh3FmD3EpnbV2dCjxdQo0079iFNKyZUmWL8KnzM1jCEt6M+2gBXfi2809gQC08zRhTTfg
0cB9OWNqMEDS7yT0I47aKirvfFhBH5KZlPV0xDxNAutv0mrz+yAPts3Jnj4n+PAtVtqwruxCeASg
gKRpcqUAfBCZLwZVZulzZBj3IrKPKfXQlou8aGSe7X65DLZklrizvnzytdpoMoEOZiJdtkel9hek
ClZNGUKkDOGqSponYHYrGBLERkSxQMImm4MB1F1tQivSQpTZf6c6YX/PBZvDDfLmmDY9iF0j5UII
AE+hU93ayWDg6GrVQGBjjbPRu0yKv1wfqFILQeaMz9/CSVQeWcoufVfRwIks98JzdYXvLRthQdCP
0aX+vn6HBtjv81Ttoqb2o7qoOuqYhr+pOm0Nw+g9mLIPH/7oA0wTso4BRu+MCVsHbH9XP7xUu9UG
ZJTKffvdWchhKFUgitvFqq0N08u0q/hNmzgE4Lyvx3vhv7/rwhT2HTt2Y0uiDZiZl/+ykb+I8sPd
FKtIX+6m0Xfx1EUvbNKUX6WaJOfZDQsF4Ya7POe8DSsVGWYvI4Tk26iglP22kFQFQyp5dBrmgsIS
lDFmGjuw8iTdHtkifHHnPhMviH3zsGYhYrGGqlDT+OM3SB37JEk+g1EaeWorMeTDzcDn2RJ6gPJO
j5F3lIp0zFQs0XdRigeteuP7L9ab3UyxREqSdlTrKyVenx117RPBSi1nmBv1+c70ZRvWU8UjR7Bt
jFcvtmqF89J6sex8E1PYAKEBebsO1hBTeFT19svuCkl9v+IKAG0g3iSaIH4mDl34sybI8LnPwHLy
1fBFbzjVxKzw3rg4/5MMS8X/NV90Fp5X4IYdeLRc9ssZKSP7cmtB2+JJIiLjEKoQXTynQAkQd8OJ
oRcrrK2pqUN2S9HEJJ+Jn7WXHqzNpvzPHW8inCpfQKQITOgXPmy1Ohb1wOwU1phynmcHuujf5vqU
ifRZaj3jQfGed8yM27rM85nqBOLrIxHvi16zViOdf6Jqgkh6qztWvnJJQQat3CP9e1eWrJs83jBy
muHeUpNZiPRdDFYmGHcG7JbMs1Iub8Bw5m6T0aXoq/BP3YqFPebw1wxd/xskzmGYsLGc4Ab28zkl
4Vyb988+SaNjxU1NYVgw/s7U1mA+AW4VBcWpun/q94lE1uM6wb5DS0LSdNNuXmH/UOmb8NMXhjZ2
p+E++V6Waiwm9mFxocL3ceKr8ONAARzDDZL79ej3T0+iuZ6W87vl5E+7F6QprMjxMhGFN1L7UdVu
K5Ypk4ObdPxINRpiCdsBLUUjbCA+TkdQ/NuR7pRTUPBbvd6FOM3PxgPOUQv2hsHJP/vzliHWzMsd
a6GHZIRTAaWfU8Ik9zbU4HWctNPk54nUNCAaYuog2pnrMb3+37gxiap4DAE3Jk/ERn2MbNQqxA3w
M+vv7Toxr4NTdUtFi9P+PE3EULb6Xms8n0BejM4H9ysD22641Jkkdo3RN06m7raF6Q93UKoxeOq5
SqxtpD5AGqk5/vfph4RecLJOdSe/QRTsPbX6cZVbGSzDPuFUG42dh+fFemaukmWXmWd7HzhVZwJO
xShiReIJSkdwUD1AEwecvB7hlRuRQBuZ6O74GizPHCg89pimmx6RVpExilUQC1KKfIpXXg9Dyo2P
DEbQYUoPOeWjFuSidKuUzqQcPntImNf9X2R/LRqJuxZRLZ1yPGxQ9T+M9KpA07xr4l36IMoHUCh4
HU+qgY/a8ezgFS117PHQQTHlFMrlgWMguBebhr5D1W4JFUpcOHZ62V9YD1nTZDcB+qk6q7nRqz40
wqzb1Aaz4tIP2YcDcBnLrTu0P09xX9K6sIsPGiXyU/aKtcsi7/34DxVZR+YKLg3nN9AkWgLD0biV
p7fbYlFSujqSlMZWITMHjW7FGWHtClPCT5E/LZUzkjxwevEblbreBi91cJkLwh/W3dTgfieUOTB0
g8DTYoXslshaPiuE90hdTBkN5VmNxsg9vvABT2DAqN1HDzdpbu6ojMG9z4geZ5x0y6bAKLXnV6Xq
xbxYkxoKPv4eROTzPMGNj6svPUY7LVAJ1l49Gog8HjV+I5Gx6w3IgMszCNpEnVviCPAN1EneC7ko
zMO+1asrwbZqjU2jpMGGKFD4yv6MOwhKbefFadSLdBclO9aUhYr9WMIZ6vYY3MEXVMcdU3E0hmbg
MFtsBrjxZ1IP/YHUnlNW88RUcj+Msb1GO25fP2TezsSBgpBw9XR1XOe83/hw+Ga4Pbe+WfLZ5fM2
7nNcpNTb8qo2lGN45QiKFK5OxzlLZyjZKGarPrecuzQsYgNS6AONYngYJxMjorlHxOHZbKh+iva6
qiwUYIuytKGe8ojk8R/Rp+PfAHcM2fZP5EjB6orDkjNZWp4zd793nRsfN0fb8EidEjLhL4sxv5j5
9wDuvdRwZ6VcaMG/OOKQhmkJhTmeuR01ysB2DyGvNYhYzEn+vlfZTV/C3e13GkkRqmSlTy4/uCx1
azjxfnvaiYDVXB8xG7ZB9xvvSGswUeLasAwAXiPa68tlwVNn9LKF+MveKWoBW+5547w4YSvZpm0V
WANYZao4Vm/bbtWG2e/WLn+y/qWz9mJ4ApaA3Vm8mN3GBB3ObmnuxgjX5YKETtMW+p+T2im6K6MH
cKU0F3ZgmgtwRhlPTlM2gdFytl5PjMv66JnRdpcLTXpHuIdh17Bl8GX2li4oSJ/KvpLFzfTaPQJ6
ec7zdNZ3KG2RFY/3+JkiAfZ8f1lut7LviUa5vtflqj43bgewtuvGK8ASQYfiGjpYzbDYtxAMdCcw
OTiQKzfoDSUVweIgxNhTjeER7zw8v3tYAr5NxGeFZFY8nXdROb5gs2uB8R6+2FWM96YWI0NjvxDP
ylFhWzSQPmrku5Y3SgI9QTku2agJRB73YdX6L3to8g/O3beAn3Uz94tU60a7ae9ykehm19c+OOsb
736HRWeL8Snz53VdLUBncM3uwk0UWKC1lZ044fzLzjnxPZ157T/S6LH7jO7q+p+H6bRcowZvvQl3
/ebed5g85LCzqgV6+Xx+l3+0okq/mt0PAi0QGHhxuYTk0fSdzsmk0w6AMZw+Ws+OYt1P6Uv2slaf
VATXzPyZ8ogex3Jma33Qv9eC35/qTUVpxmFU4/3BEXPrGgRqFScteHj5j1nwGYScIEIS6Q5nD5ik
vzKbQ1Qg4do71Ev3rechbt0Q+ojMS9ymFAN7bNFliajAadw19rD6J1wiHJotfm5M3QuBrXgRp1FV
GSndPNhBxvZvOKHvEI+gGy0Xv35164QN+YJpbwj+zVVvV+C7zz7poYfR0SG7icSyIBMluOtWhqVD
bjzDGqb7p+SvIDNkvRbqh930ddHKdBRQfwbB+/Y6CuYnZAA/wJfaiAadCr2rd7h3GFevKj/iIEap
Zy3SnZkivOOC9z+SGd0Iu+1krs8y6TBgYRozOTVdGsks7C1dYASncaMvQs+79ZvsfPqnX6+8aiLG
mR53V8wkD7kKZFFmPD2Wcyw/V1zO4czsM4N/+i68axLsOk1YnmgPuvniaZ5JVEjJTlHblGGXiJPl
H76ZxW9KdEmF4G9hZD3EldAEY7c2OrportachaXyeIvenFAtnppE5jpuDig6QKeXr5wjA1V1P9Oj
WqURBFR7KQkzaW94Zd04ejeR4IPw1Qw0RXB9tK2bJf8s1Fwbz8fgnxFCwX4z2hSKMFhm9WZPJbCI
B81Vz5oTXIOkbJAeMks9DqXrLRAETUJMGL1Pv3PLujn8V+mXBl9uaLVD4E7N/8KiK7idjwuaZ2TG
2ilKOkQ6q3NS6GNP3D1AnPqfbphoV2T6Ur/1HKXpQ6zj82Qlva5RUpPnWPdvuOJjGxIa2jsxntpo
hufdbQBf/oju+Ewn6WNy+Et0DSYrRBXBWIpvSHIjDQ4W1pyO/tBRUXzy0jsZ0Ru1FZC23ED3wxyI
aO0e2wYCDfHq/PaIPbZuQZeaB3FuqfsnWu3ymrbphQXuk0WfWEl67FBx+ngOfo3891OiHch5dxRs
M89oiCGa2RVOPX2vdSErvtbRDUofdrHO/TPnUnaWof1wOPB5S/bVZ0f6SuS5b9hzpnZsTO4CwZ+z
xCWF1nIVQExvE/0oE1zckEjY3LfJTlMYNERczlbAfNvcMJjfoKmASIjxqBRK8Uh7f+tgfJP12+Di
ffFXGAMrFblUsoD2LLsZZfkJNcSNp4CgojZmQR3qeZ4aiXWPn1/sp78VLch9mY5vf6S/6kGbe6gA
cm5ROAc0/4oV/9J0mMZhBDrjt5YMLCYPibuEsRTKQRjNXb+53At/ISmaU/bYjtkKIyW02BXrSdnE
yBNcP9GKSYAlMiQtfDQOWLB1eiaZHcCW0OuQjROyOrw/2ncSIQxfJUaDaun3x+RNcn+2/R5q2EEh
GcKmNmPy+vENYKnI2oJ75kPGASJQTzRg5iVUerOIpq+9XSecsQQvnRIY0YiUMCb8UTiW6+KaKZfE
zkv9rntiPQBOpYXft4xj6V411pVUPKYn8d05fU0J3bD5P8Y0Is3XOP/Xx5K/y9R63J+tnFykROs+
SXfNW4DrXB14qYIUp3xIht0dAm7u0cB4zSOQBKLV3BLPGRDNUvpH2P1nZZ4BvQ+ULgo7uzH/EOy/
MGIPk33xjsKtRMNp7R5fYoO+Vib/vX4snjvg9sLLdpARO/EaI+kRjvCr9ErmsjBqyuuLDJQipbyr
J4u8/rfmr9qOlLWWq0Kiv37MV6m+0rW0Jsm1RXEyvUEzXjDAKblBvXJz8eUNaxocQk/dwQMW5FOO
+vqh9SClqqtwa14kxOKKnz7vpA9ovRfKIk05BUFKXJDRVGqTgUcNO2SjfbIzFttuOURJOctRVeQi
FEaj3pimD3Ory+VNYtkYloxQQxSjFLNnDprECjH9vVEyzO0J3QYfAKPflYP0wM81F2OGoUc8IWIN
mrL26ma3dY2D8X/qjQ0gKQeGkHTyPhYBH8HsonvcjFdTX+6at1LkGgjMdDOBdNt5HJI2rMJMdFPA
CINHX7HPFpmkDXWNlC9ONCpSr7DPo5GqQqCckxKuG7h47gum9fuPNQGC3m/iEtm08f0vMP1+OA1b
WDJWc1a3I+WHF//NcOfqHOaVSTdmtXAQBuQzHXAVWpfUNcVB77sxxDNmC2V7IrfUTkhC2JRJwlG1
8zyFY9urpnKoMZHtrTHHPMuIjILGCuGcEFGazxkiAqG26PpiAxclyLqhO/vihaVUN1DM+V68Xe9c
XcFs3qFKfgIglsxQZdnDWjLO4mW6EYprpoUUw5MswqhdKLbW3petCAxf7W8K0AGs3HRekejsXeVj
7WvcD4rNLlsEC7e59k5RlRlBgLNZ4sUgXGOerBkpln0FqBU4G+x9ZNWzkuFxkT3VkhCSX6OP15n1
UbIXiC6aRLnLa9mKBjgubVuW+u3c+vHGNhjkFDOpVPptWK4jNXRc73vgdmJLZcPq03sM/pfX5r5E
vsNwxqQYId1HokSLYW9aZlO975iKmUpAZ/zDhIef8b5jP3wpsttCveKD8hVUI7sOaER9yP48KVs5
BNXJH/PqJuzR5cGbNPDmlEvf1YvdnfkXi5GQurJ9JQ50StDfH6EhugiLvhjAfFUHrt5z1LWk+Iwc
98hgElKLlq0PZ2EqSP5GDgYGIm02R4iDbO5zXOQrvGI6sIyoupRekjXPyVFfwojS93rKyYBueaVu
QgdRcVE2OWmFeU3UzRFuvBvCq88cpVwz/yIKkwRrZed8rsNAhh1ao7SVqeE90KR1Rjh38rUxENDK
b2igupLI1YxQf0i0rW/xIw6i9OMW82jXcY+HigaoQDAq3HbDm+EUejRLjtfeNgBqHd1JqjLFdHkq
9BBQFjT33QECDBzDQw/cV8CVXaugn8yHyJB1uMp2FySOE7vuCB5sU0hjaa5gYVNy+OmdrujFCJ8x
T1keZezc+DLkPz06kXyDHBnudwLcIwKscY1UL6Uh/mYvwoGO6NhSGKtj6/yhdgYMbZzs6f8ZaZAE
32fhxC9+mDy/V+B+DH9ImbidHZqDN3oTGQ6XA+JPrVFMr0MFDKIYakwqv/iCyIuXn7o6v5xNpc79
XW7BaWibI1M8CfQv3vtyyifffpU+eNXn+1/PLjjUQ+6e5T8GWC4/CiNAEWmQ6v7kZP29JtzJrQ7T
c3s8DqSXTyzjnM4aexgizG40J/4jle93fLC+7927EuDXXHzaKmBIDkKRG+cJt0NG7kt74OykeA/3
X9sOyKqcSa83tecz+iKjXLGETJ5Zuu5TSfwkZi0R4lcBvsv0Z22t1IJ90mN7ocB+x3k45AEa7VU9
vCpgAAtidP5OqRoOgzh836emdlcgaiGMvEFePd48STUElmkL9DnEdR/EcPXis13P+JkIC59/03Cl
o7xQKy5h9XMrS2rFE8t2TfQriO5qkxleBs9wrt0P9pdOIUEKfyymT0vnLxoIlowZc7kloiip3ANv
3CXCyR1HwQ50eRNKuyJawKBmffA3vuSqMfyAWWU0YiAs7jmNezfCI0ey8mKYlB6M7xQNPROvO5tS
BKJqH99d8/UkLHl3vO7HEj9bubcwvGjH0rRECScXiMClAzt4yjV4lO8F0bK1lY9cG/4/17Rtz51d
MzN2hlXjf5kDLvGPkfH0utXxBK2GfbXnTVCkoo9sJ6ITisUZvYhrB+VwkXQ+gm7SmTstgOBHcl7/
xC4XgVTbuptlRUrtgdh3cLe9Kd9YtFnslg65DzNJrU9gbsSxH8/EQ+HqoJSTw7Zt0ymOyBQfu0iK
yBzfHvmbzswFBh6kRGkLWAdypNEax4NVSjRlmsm+WUjkKAuBxpahUGQBJQnrkLKP4ABa4MeItH+Z
mNNjT8gvsfstmZshygu5Tzemx+5XWgnYAYnsKzHjsnvXy4YX57fNKFPDTZ5zQQC0+ExwAEIWEtT8
X3GvjXtpFIUujWmWefiS5+zBoXf/gCgEgEL1JvNNh5oHFfM2IOaKZnKOYFwAdzDwzukCFpMcnsch
2aqzEGE+Sw06gLqIVuZ8434K51e370YCykv/5jMH97jBghAX7+IwdOAXU9SfrfDJ7GOfRwDngpcw
T4eM+BQmyJC6B4asiYBsccKgihakQY7U4SQIBInxWK3FEfWi0GaaZu5lEvX2RIRCoWZY8GE0V6vp
sc6GN+zBBAJewtEuA9Q3cDzqjPIR51YyFiqnIEKgk6ZjVH0ZniuXvrb2Bmp80rmywiRlPc1hPwq1
TX9zGk2Uy2MySASmXv0yN42VvJQ8+bfn7iComvdJAR2KCRiE130MocPd+Lfx6RA20sQpi+MB0Eyo
S8TFzbsKSOuF+NenVNEDBl+fPI2bwli/QBQOPWMsQDqGgS3MSk1MePX9+Ng2b5ZHW5wun50aj4cx
TpZfFcaD8AyWXLunbf+vPQ3JccngXUrA/yC8gPNUH4LbzgXoV/Wi3ugXoh9//zZ2+uNZsqnEtU2l
lFZfSnXtYHFahsm/imRjrvNO7GVLpyA0c0Z8Qg3ISf/YoPAW/jG8gUH1eiVdJw6QfYY4jB+DIW8v
8y8zRK47NJybyCISkIcjw+S7xudMrlu5QVZbxouL76iQl+m5I6TtGehfPJtiBeYMJXFk6y1b4fBV
ONm3giIzkf7G1w1nShWu/Zz2lO0+eOraDLLNUHyKAGJgiHeUGdaDeLaPCKU/C3ZnZBTpBcOaBgyq
xfTuKcdJhJpcBcE7LkY0lHgXRvONvA+oUFY2IguM8UlZ71RWyvOLhsog+OlHSHzmSozNPcb8U/6X
F9JQAPzcXF5RV0c3eMbGmrmOcmRgpYhGzHQquTSF99vrwbPNU+/vB4Nw2P6Tr741aaYKOJqmIc25
c3cnrHESBLbwOSEs3Dz45cBY2Fk4TANCQROhYA+EN3c6BLVkmqjGqYv1GBo50DVZItPqhxpFZQXE
N86pxbYTJYXDAaW1gvbGdOeAIB5a6DzkCsI1uCztYs1CXOBgaGTaUiV2Z146IPrAFLSIw24cwtI3
avgowdZ0wcCyPKNVw+mLKIPbuCeZnV1mfKfPcWYJ/MA9bTbFFIrVAanxBcpi6GXm6ybcr1UN6b36
SNRPIddTCimgRCIXWUEc93uzrQ/ftTJ8XIVOLo7OiJmQIH6JlCmiuqx+6BceEHTrkQKz1HP4HBVD
ZhJ/RAK498eweCGZ/1Z8EqSgPQdNN8LvY1G0c2VqHYDWineBXVhe6//0llKUv5ciiQvGnSdAz3+o
NQrBoz7SKT2J9C59HHUW1r8M38ZWylX+9ynN1PLPT4Kc7fIOup1+2Zbasxgqg+asBwmtmEsg9tTH
mMJYDx2Y7WfHNoC8vqJrxhEZkcDVZIf9MOe3D0v37tETPFrHoVxLHMBv7IKJUXg2J37Mn2NnE6zZ
IC5pff+c7GWlaXboEP9Cd+GawJOFhOeAvX3W6Sq7PZwo1j6aY4zOFAp60+tsS+RJhK/xSIV/kEnJ
0OZvOrKd9wK5iWipRBgxJE5zTodv2uftxT9A3y+m57FzDKax1a2dHXU9Hb63pKd0mxcz/4Fw/Qor
dkQjVdP8xpbyxbaCoEre9KStQjYtx/B95mvbS1FWkbWvp/32YTgRh2MupBfL+xL62Om3NmCA2rZO
NgIfaHrqzC7M7xN6cjZDdUH4g4i8HqdV0n3y/msd2+hRt8G1c8N5NAXG0k9KxzGRpIpwgeRpIjux
ygY1wHh1wgG00Q96pBS3PLT/73VjBr75+mIpEcsNcdtjVrihuJUe7Ot1PCfM1GRGE2X57d/+JCG0
Ptj675lDJntQWx6C/BIgVt6+I4rJoIzvKNARQjNNKOG/c/L0ooMP9Zax5IQUdBZEw8VQPyDPTIjx
a4F2rK7Uxn++uRDGt5feEw7K85JOk6/PjNuv9z/Owc1Gbv2a2C1FWcGM35X4oLeDMJFhmcuaVmo/
zpSyKqL6/xnKsEAfxx2YNQ3aE0o+wUWWF6Ou6dbcQ2agnwSGCI+810zpPtTqtxpPLLbX2lRX0Bdq
OqJERPTq9pdf44qQs2rHtIhbATGe1+Q5+mQS6kfkxGxByYZW3K4Z3p7e7vbg2JjXcxwW3502eCx5
YjZvYbWcto4axThiCVUoHwYIdn3iL5DDakiHvyIIkoX+SnKNP7NejwBAR7wWXLk8+rUxRN9rqF18
51P430dgiO+Or9QtIklKqLLjrfYy0GcS4yHUEUAxszYcurF63VVZXhJxUQMHSWPFGo7Dg8VjzMN+
32iU3P1q9dcHMEBRDOKX7iXHUOQfyuA0CC3+Urn0rDgdVhRGzMFDqJ1tt2Dhv2SL/NFCsbv+vu8n
+yQ9zgdYnsbWR4OL1b2c2fm9Kw5baKRmeTDD+Ihux7ZziwMtcjd0ZfH15MyyCGy6AvDB2TLfpu2K
hQiIDM6W96ha9KK86/ssK0CAIRroT3dO8QWQKWqzk60vFyTmNlSGGGe1atsgJRZv3RR9W9GMaGuE
YKxik2ZlIjmi/5Sc5ItbcvAgQsXyNsgpW6EdS6PcdJI7mDkD1W5nxDWkaSwdAI9iYJ+UiwI1V/Hw
Apw3f1B/BlBFWB5qAPzpT2Ls1FSDpK//6beEkJ0nB2EvSuydEva0PlwQMgTzvMxbiOZHBNx1Rpas
yRCD6lxmNKf+K8OHbzdTLu5YbZx4WjawDvQXDtvwO2ekHxqexAWmWK/SDXNHOtLOyKHU20M3qQB0
z0iHHTBG4nW3XFhl1vcWXhHX8hbUrbZwHQITkXtrWZcd+CNpn9B+HvyMNggOutpQ7PbS84/o9Cz6
H3dT0k4elqpHKyW43SkUnzuoPs/PEnMJnqYa06qjZgaXA/opgDXH/9uIoOv96VXV/HLgRU5WN2F0
gA7rx/J8xTLQuGRjsYcv6rv5d3tCK/ZGxc826K0dCBophBHsWQ4syy2z3km1fau13uqh+A4hv2Xj
Z97LkjhhMPUEtkf4BA4ZwrR1JagtDxk0Cekgv4WDdWlZg9/n0s7V/Vrubk+4I5O6u2p3hkj3VE8H
9afrs1/XKAABDZVO+NOMVD3XFVRRMvPBC4a6rLTNTpw8rg35YGjHFxJ7V48uMdTzpqic+3Djya7O
ee7uxDIkhUhQHLCrTDJX1G3GVgbHYiInpEskX5Vi5MRE8FEwTvSewu25ylmvbFsDSo0d+SK/9JiT
RiHAWUvoJaO95ueQ3AsOd0gl7ap+73u2Gqv+nkYASl1SbMotSZJVzbh7h96xW4VVuOKS3IK56oMT
Sel2EJPviLmRU7/clCAWI2Lud+dbKE3+X8YXO9ckeRl7aD5P+S7OcMttpBTbNq/xZj1tVTWfF4sd
iE3K/K/UK5AI1TWijcMPTluMucA0pZ5ku3bN2XaoEtBT7Z1mRLaHaaqT45rTqFCAqR4sN31KxeCA
YBx0ptsR6CtrXuigAV8IEFNFZJvsojyh4Pl/f7wsW3qhf/Q8pzOTsq/tKqOZb7uo3/lQDGIgmcN/
OAY5L5ead+cnmltgEVGU6zlKN3soxL8pXAwpFslADZmzjsip1dDKNTMlzZB8aZ/LY27hTdI9QlzQ
EBhpMUchdlQ3qv3umZfgOwaFomxeRsHncnThqUQ24+/G2u5mXEYl+A7VkroZqTXOeCg+MSWRl0Ob
jFQr/NHyZjuj0uVsjsa21yiaF063z2H5x0khSaS13MCZg1L941Dmr1dlIQpxQCqESy+q+C9rHaKJ
72o1yeEOArGAXGhUdlKYMr+HtvufBBNTvM+ZGlz1NajHcUrmnUg3gPWQIan0vFQsZeCW2SV19YcN
VBaxOLlo+8Q3G3SVU5lQXxMViLmU3iH1j4gUV4YZhheR4zZzEPTOtZTAkjwYftOWU9f4ZuKf3OEa
Q7vITQDzhp6/Vth4XfDIyn4rFpR6ORJ7zY6yAVOZkf5u124Ih1RntSBI3j1az799zLeG+vHt8CUe
P+Yvn+iQnlQkrSf6BnxFB83/ludKNpZoRwUh/gbsVEzuA1WoEFjUL9SVTDhGzUe2+47R/Qu27lce
MnrXY51uwGoPzo08NAG1Sf4vk5H7ljvsTXbolVB1CrArWUWnGvWPh+Q8bv9VYWxT9X1etv0t6sV/
XN2nCHV6Yhuet8nMs49kJktqUOnIvR1CEQ4G6PWXkOIyCuMAAUwejUXnqi9xorFx0YPbLU7fBefz
8vWd+Jvkh4wa+byLW36r78sTgy2jwUIcS7f4IZu3Icg9MVBI9Gy6BYyVvYRkMC8NKlIONswsqawj
Zed0bt8c3a641gMlwqxo/ugxQZKNkqaMymp9jX5cwY12d1OaCKpnF0ZLYftDvyO1oIwlrPLw6R2/
ppumsNXCM7SuPhX0eB6kOavz028Cg+dbnjTjylMxT4VVm9MAFdBJ0dB1GGyePBMbceShyMy+aGwq
q9xeaFP9KXDFPzWM5Mvt8SIh70SgftREbU6IA1zx/OVpFkWmCY0JjIMuw7Xh0G4aLgVX55DFPkkm
TboQsR8U5yL6njUb57rGRyN081gn/2OuTBGMAV2pcB9MlpPPeWpwtPVhCcQA24q/c/Q8vQ7V+rat
spSZtE6hYiZp4Jutd7oxNPlpgMQdLHcuJUiwRcFdBpz1TLiVUGcRhsBLDGRiDLYs5lYqSghgk2Uf
d5kRSAwW3fqKxFa+FbR+4hRgHT44TEfWd0Lnvqxx6VVikKZaug8qMCznkSIAPVsm1OUlmUQyieZt
pCSJnlqkukbzZG41Uaq0urDQH5xNtt1s/4sDi/ZZ8Be2+saQDIHMW8FpyvXDQ6tqM/O7kTQrDwEe
L3XfIDV+AwVkvWVgYAvBa4ATCaVrrxucX8XA0l5xxVXhV+Dy+n9BouvedV88kyX/iIQNzKyHkziv
IjLaJDgLVVLKfYHDJDgiJu61kEt6sU0NOJb7BQdfWb3IVa8j0XTgw3D2hGLzJI6tRqWgLlKns5g0
tkQWzdlaOgQpLQ7IEMRfXDMl5qbydn6LJkT170pARJju/fl9v831mctbOWo4t07DjmBDpp5s5EJI
CbTEaECCAcgcMn+89kyaT5i1OIXXxW7K6vphP6ZBpo/0AKbQtI4zOpw3ecT8Kvs91Pye90svlX8W
0pSZFX1BiBrYsB+VKiHahIxtiS/Ucml58NOAb+on++d3zqjluLhm1iazal51Q/65aPEmHKkYPNxP
kXCEgqtG5OwBwQl78nfzwk/GVNSTfTdbAz6s8NLLe2qG4RNa9J9cEA/N/ePnyoDRLPgNCNwq2VwN
cNzbycRVD84RQtw7rugR19yVTpYIjJX3F/qULI4mXJcWAXO0P8dZ+iwKVxZdv0AhGHddsRKm4ycE
o61/mHsFR+kzD6a04KH83TqNrpwI3cU/XFD1b1R1/VmGIqDeVfmmXSmrIm9Zth+d40ZduQSTy/QJ
LrSu5WrHpz2grKmVXeRcSwOqC48St54QtRtKTgZk+FsQYGSZyci0lh7l15Uv8KYazNGPsjihpT0o
NM2qipaQ4yJT4ecV173qfUaDNl64cQHaK/cU8veIGMAHdfjkMb01eM3jjrovOkPzRkKAZGU01uBH
mkrOSlfkx2GKfVU9fFlXZmk0Ufa3rQuQX8bgncN/dvugDDUEJfjDYDIjRmOiRM3ejsYGtNoB/z4F
xG8BylHrqJIK7sSjQL9XD6MdYzZ+jeN8ZdaoXrBEiQqyxJbnG1BjyWs7T6MIh45oFhg8CUT3+ohU
K5yqukRMnhMFG+v6gruCe31/SRUEZkmHHdkYtJIwQCI5tMWG2Y+PA8z/UmvlwEI06GkkVVEzqqGw
o36yvl04oZh0Mc+zTPwmIbO1lLfA5JPO3i8J0VXtMH2No5kz8Ei9DvzZggx92hOFObhDyUDf9BJd
dvP9I6JywtnHGEoy8gbCy0EHLY8N5MDe5irFMCfL16AEriMwEDRyhCUMg8f1aaVmKCz+l5yAjy3C
T99YG7UyYHZKueRw8gB7kk3vjRAnSWJINTA+nUXY531qRbDInMkY7iU9Y02n+rlvVK389QEH31SF
BEE5rGEIe06KT6O4rjAA4NeJhk4ji+Xif0bPxRQm9IL5W0Uhxd09Fi07EEgKf5rX5wx5q/RB5YZu
NfvgDCD0lU+pQIPcTzjCD0lzh1BJbvHqYt0D7fznuapZfZ9Gnjr+CjVbtxjzGhmvV4Uf4Fnp9FnX
A000WBtg5hL/gDv9fjEArbo2Z2K19k2v6UdBB4VK/9QTqvsUaGDyQAVpeU5yyyBJK59Od/ZZrgCa
+BuhBd4HVO5h0bZn11Iim4VWCIVriYbKhyfmnb4kH0nDx7H4ODcjy8/MAYUCkCefXPjxIflNYYAT
EqXR2qlEjn14q0lNNLoIeoBW85zVOXl0BJOSsrEzDiNoy7kHIfaC0VDTIJo8ePI7sBnBwnzWrZri
L8bqc2RkNAGBOFXiAciin7EDxz/iAfwxGpS+U9SsDH/Ml62ghleLpI09DOb5GX64HEx3OChEkCVC
N2NSVQg/NWxoCQ72VIkrJiH2lgNxkvQcsY6BT0N3HGpRRGaly2dMpQs+BDiOJB8FgyqmnF1AZZMh
81RxsWIyLxZXxVm4KxpDZZ+Si4ZNl1Zk9H1ARz6RvDHljiw7mVLcIclLL0fI+sYolQiErEyz8U+X
qZSSXDuZnB0aGjg7iJNd0VXCPgyHJfYh8xWjH7MFqzBK/baqI556Mp8IkJEQ1RRNTiAK1PuZHIe6
vkIWRG0q6xOHSbmUmyRLLIxixC190EEfN9cE6w8dnRgT98LNtZ8uxuNyqlJMLVFey8PVNbWLSXZM
QZ2iySC43zrHT+LiosIJ9q6/c5VTjZG63EHXtMt1GJl9CWkyHzWllzGylg5PEf8QKuFkX3mA1MNJ
t80qV/dXNila+ZTvI6tzG5diaxQVkxSEtIwM7OM0CxafKJciO5waJUTi2CVZByTPDVoNKn1qZTF6
bjtjuwVyKxHwmhtsc2HFHUFMYsF5maxZOU6QdTPHMvTVbN2UJz+fVor1iVwSI5u1Da6EMmdG6uDb
bXYxpxrq4ntw6WkPX7PVmHcQdLCgFjKQnC2O60py0ouXu8SKGYUfJF6iAidhxMqHdjy+t/m2mJFZ
vu5EnlXXKgBQ+LiJAcBV/TzeaURy0swQ8FQcPMc+J240Nx96wg6Aif3v3WO/knufwn/Uons+pWbV
Bu5YfhlhtlyhgXyxkFogT6YJngBlfjO+t5nfKpHNictTYXIIuiEcHQGJjsC3zu56lkcw1vaRnULA
Dt0JU4NN3pA6PDueHt4EwSDMzkK/1BnBUXSDaqJ3zU7mGZageUrx43CsK3BLMFbn6WHY8RqvZIaY
zpjy4u2ArAyZrxhZZU/kZpwQLsAa6DwGJbNPvQnSW2O4FMWtiwhLdAon8Od7nX6bVSIAxiO/1xAq
0jKXkvjhvvRFWqlHt/Q1u73Eri1ZiHawh4RdCndPIy4qXkkz9Q2zPOe8IKPDmgyf8jSBPIKgUcxx
2KreYd5DpchyGBbBgTGTk11FjJB6XkMlvDLbXPKym3EvOiul5ethJKJ+kRRkMJ4rO5XNooVjFk8E
3IByOleXsVB8DhtY/vQEAlX2bclTnvVu1/YhNkSGYig5O2RCltvF3nQO7e3iEbsQWUSFDUBCwlUd
rFvtT4IFXU00h95NO7ugyd/4BwdCY6dfC7tKAsEVfDGDkNIRmFokg14niwNphk67KobK87dFQTp7
k1o/iORUbuqZyfheprBmSQ7Nrhc5eYEmOh+5BzWNnsPmRrx5UN0FmKO9iG+IR0V9kwun3VSngZ8N
OqO85vrqag5z+FbKYZkUsomWiG5sZQHlySLLLVNLOfNxZmWF+twBf3ScgEYmplTfE08IJPejhSde
EILBmdi02BIyYAaIA40czifYKdqxRL+RvOs5xlb6njgfurQwjBwJ1ayqgnF23U3xOW/zNrLZF6ke
ZLRhRRrKPHwJdv/BFN30h5KPxUmJV2n4HKpDg+AoGQQc+PVyeK++yEgZZ3TzqVConlDFVF9T0RX9
sssaPV5zAe2smwvjTyvAlniSZDbY7IGqWB+Y4dwLAfYpzCmJHfOh565oEFbIk4Uv4rtgdVjSf1BM
q1tv9EVIEqE5DFmCGg9wYcuHW/Rlf+gRrwpHNxKl2CK8s1DKTHbzShoyJak7KBhuuf1WQigLjk93
B9v92jliO90iIUYYE/lSog5t0ZAeYB8Hxy8ZS2Xc+aK1r4acXUXr00mie4OqwOB6THdS80gssWsD
B7kKOO+aUM6/B/AyDPSFQ7e5HMnixUvMlDnCuGD3gMc9bKrnI/C68qfBjqpnTfc7MODuyNtlo/aU
W/UIXQUu419XXVVreLTVMS6XKle+rHJGau4EcQnUfEjlY0atMA5Q7DqBSZaUfI7ZpQRZrEHCtVlk
nllUwiWl5q4bA9RlpiXDrwB5l8XZOd9JLUtstPgcYlIYUKRAahZ97EyMqeKvJr8H5WhdKvw8nVOe
fXoQ3QOxZkaCu9aij8VZWi5Fy64BWj/VBttBzHKeWq32r2buirE6h66PQyd4ijYaxYNvQbw6LMBN
kJQO5OwQOKRAcu+h26eDmT1ZmjT0pR9eSdB2eK+JYMdf4rRq7jniibjwHbbuwJpg1o6fkcaRva/n
QRBMSNOQC0m3xzr/yXg8FHnI8b4SJCYulLaSVFeZfLf3XbcRZS2QtMFnpmBggxvuYa08e8ClsOk6
2RDrFE4D1BGpnQwZ2vwnK3vAiFeNkFtuYj1BI8myz8GmrAZjAyGfI8RlP72cwZNaQrJu8Izk29jN
yUCpwGO6OrJsV0BlXk/BkJJa2aQf5w3O68NNJD1bBAcQp8Z830796BWNpA8XB++yu8d8wCGokcNg
y3PefmRNdM//8v8aUAcuH9TEbRiIXCLTxRhezSYQHxCDkP3WW12Wzs4lr5xYhdRWH06rhl7IgYUL
ZVBxUEqOZCfZR7vuLq3XKkBquZKq1PxM0b7t31nYz4PCcMX55K6fjzndcoblK1LR10vr1nVLMs7Q
0+m3TQEGNZOt4eHGkYbG0e+n/vq+RlloXmhUXQZY8H66T46MsaW5PlMPh2snUn1LAfY4NbX0nzJC
+NG3wha7x/4qgqj6PksMrTrkc7a574p4AUx1dT6ou1DWkWy1UWrZNTHMYrSR4XmmRrRPK0xuIy27
p5zVj+EgX2br6SMEZkv+Dhnei1JOsnrigqff7NBx/RsuLPfVkLwm8xY9ZTeRCUzv/i7Fi80JErY7
SYPtXVCq8b3uxzp06gkI74aeQ3h5jOuhsGe1MndkbaVcKr4zQgjZ/Ws6TiVNcLgLqMaKJMsRSSLa
Gb2T68IibFc7TTfzLlP1NibsK20WVhegYxzl7c64fPcTwtAG1z2OpZWzOu0aPiP9G47CGxPgG4Q8
hf5vWOddtkqJUoG/56xlQSujoUkosGf7ECb7whPqWyYI+KSPG00iAltSk78kAu6254mnvNAonLIU
PouZF2JV9eBsbS06aPEmh2n/cbzgZRGhAIoIja/vA3Djw+uc1VarvuFJpeGEUp9X1FkS1BzuB3Pw
dbQhkpgbylH/DmJjW49clMOiHuwiw8MxFRmwoRiLoHC3xwON4RC9utri6Psn+RBRGmwS5CrYzZiZ
mjKqJudohzgHn/h0OW8sv5Hzxms90awa08Spdjufb6INXtOmRn2iAPF25ATzXIou4S+H4pEO5ZO9
CkZ47pIl0Uy/n/+Ph20wRlmJE5VsXsyYjuK0DSC/DvYkGOMGXEx47ocC5tISxHIJB3HWjXuPDhez
AGVTwRgEk7mIq22AqJdbWHRsL8jFGhFBCdt8aV9lpGUoqSR+lH98xs5bkZnRBSSqLbGCCksc+Ena
zjb+45LF+K4Dx+aPnWKrMGTpIz3Wwiy3Ebwq3ZVf6UrA/7urZkCb5zjgkV3XtB3cID/47v1L2RMe
L5QHK4ABCooo1/hodELKlwbSS6/0OTOr59CGwcOuUXBPYFsoMJsmYrNdxhkZZxuEmGceFF1bkyol
ELIctw5FhpnHv42mS1cWZ+cvLoyoztM+d7K1OnPKaHXskwPiMwj2ZTszUu8STpnAWON+WJ2vK5gU
tSXx+NsyhFdCjZ2NaY+dOAvMPC/+wdiuHT9Rm2RuusUI06Ggs6k+jMwHVyYu0A6024vFFhTHGQ0S
hE+QltPU9MOAaJqxVaRVjaJ+Y0tiWJ3d/FYuVMdXIGfORtp/sJGCK1uwocILRHTxPEGhOV63qYIO
ryhjDxrho7Q9AipCNHJprQ/Boi5wBnyyJqRe2gxz5yLRqUkSviT9ap1aPgiGfJVRJUkYFeT3Uw3D
lSbRAN939aLGWQrMRoD2u+S7loQ9/RV5HOHwxG2HInpZ+QWxRaw3p3glUq1v2lFLgNpCGdhtiyeh
1y7W4TqjhQDO9QA2aC4+IWbJsqjp5yerECGbYsypCZz2oc5UoPXXKMIpTs3FRNwGdkvAzpUTRpyZ
QYUSoiO3Y5AfDBrqE5GOfqTj7YLCFh1lWXfpYG4A2s+VGYIByKWtZZ911HCGdWZlsgM8PXVn0+kl
4bM3SE6ssCrPLUUEpVX3D/xtUpLgvDaQw/qSXDjyu3BFl/PTn0WkJwkh0geM07WMkPLHbzvivKSt
dLYDVDVfPmSTBT/6f2hV23Ozz1IU61eX6z+goXXTwem7SbLe6z01FVYzpGsfl7+7WZYKRjHhZJ3I
uLy9FLgDuGwCQ1e5hy/0vOOCpo8XUFRNe6OuURpOa5l4+1lCiO8Mwc6W8BeiEyNkBtdYEwt7au2Y
tnq9FyyzKdUYkDLX709aOUao7/VnnF3QXpxG6dffjYqAgET984U2Mz0uzHi1OP0Zr/eByFIZiKQB
3VMJoarrM8n2eyl1I/2VvbshuK9tI+al4gCz3iAOq3NYo7TflCM7L2iUBN4BdRFkM+eO4vNu/8oy
hIQSW69C2qUEJVWijeGC3ydP5y6Z2JT90pbMILi2YDEUYP4O61Enskv+Em7On/OXIJGY64rSMl+5
KcuNRoOTNhugOcyRNqXAABMsHtcY/DCQ8FphcHcEfgjh0fp/yKqWHdt8vA5Kaa5dhtCtE6vTDfbI
+JKH+y0xeaBQd6Hgdb/d6uMOQ6qq753S54bTkS0o6dxFudcHoqshvHHVp0onhZwSnhd78OAmJebK
19kSlZRkiCuk4uOLLoF4vl0xOPlJRgh39LFZsQ/LvLWecgZPc6gCqJXucjP5a1QjUMLOyNKrxQ33
HK1XkbE3bFkk7lgpJqJSStagiIPfFtGBj1/N+XE/ZIc92p3ytHCizWdW7ldDDVWnlgL5qLsbmkAJ
YL/VKLZGZRUFPRzAQklq9xmc+cF0/dClvzyzWVMDK2PJQhByo3zsLRAlH7Lna9CuvFyRcqBOdW/u
vf1UmexqgotMWwLOefKOhkIVAfq+JDl//AsI95wnOGARvylKQT7EntSgLy+FnoQlI8Ymi5x9pwco
Nx6MnwvU3aFW8KqdTy2GErEexFmADIzxO7/08x3OMclf2r9kJrDHRr1ROKAeUE0aznRZrsYzKc91
P1+mqfzoPtTn+7cLmDLjiA7fqWqDdpOdTd5O1F7HtwYgBH6Xa7zcqdzmN7s3g9vdi4b21Vr7PTFs
WAsEXXll1dvpEb8sYL//Wjs2lONoHIC0KJBCpQcbZF3JUw7cMzZsTXwjFNr63GMs1b6OMsPk0XhP
jqMmLxO8zNOrf+6ULn07dLvAjTExt0It2JrMjuVabKIqNYfN+piLgPjx9McUYyGI77hx06w0CyY0
TPblOakAdjovEQAYi+NACuIBWRZ6wvGwy1v9p5JGhVBV36wOz6AME3db3ju/WKSLsrm3O0hCtY3V
BDz9AOgBPL/oKAZLAaghVxcreF5SiFsWGp7Di9anW2nrV/9bDvjCRwCGgDpGd0AqeJtQft8GXH21
qqBwvrFTXOqDsKE6s9e4/5fKYuuvUBmaNuqjRvZUgW8n0zZirnkDJsWxYqbXDI/93ih52wfBLN41
egPnvKllg245slUEkTfPTNgaE6SVDAoBm8/MsbJk/u9wBho1r6RwxA3e5MIbAgHl08sN3FF0NJYV
O/KLfhPvkCoXjGAqvhw8x/PpwVDylzQSvREVANEvT0MmPs9LjfnxdECqofV84IIy6TtEOdkOxJap
ELO5t/xh6YDNQykF9Fy123wSD90n6DO14XnNJc5Z+1z8SY0/C6EkTdhIJGHdqOZRd32X9+/wh3ZJ
ybzQn8jDNL3bzBhMJG5EEEda2k02gNWsOr2rowt1Swm/toRIh+U+RA5H5DpSndG17YWzHdhcm/8e
IcX4cEqQe86gRBJVKJ3+xhL4NcHtOuKWvXOxXuHHcRba4bYrF3SMH0BiWrml0dbzAdTEYhVBd+pD
pBaXAIG8bzLnBFuwd+35wykfjObcGL56vjRxlnJwRfjDqoSUZ319d4spiRs3VFDkz8dvk156b9Cj
HitFTHhLVrVgbjJVSDx55wJ4SxeM57HhVo7FbGex4zG6gjH5ddPq4XgcCWhVaRIujSGjPJ+BQFWY
5nGp8mSDncu1Wlp/94Z0L78FnaaCEpakwrw9/LLIeOazy+xrTf2ed/YtkplRZD2MTLMr4NePlCEc
Bi0GIxC4o5XGhJ4FaO0kImiLilIsKI0XxA/ceWY2ShmcmiyxtKfnbFplJLSHBfkeePa1QltUXCOM
/Bp2Asx1Ki4JktHEx/P6Qs+BoSKgeWVKDe+R8td6PR9eWgDWejEEd1fuw7MHK+lPjkyg9IHB+07I
sAkHIlb0UWqC3qqz8NXrtpxnuLN6l3q3xX1VxuPUVmIi0aJJtenhJR/5BVIul42dnxA9R7DcJfn+
QnPtIDVBJ2MZ9yuEB/o9VVEoBC+hNfBOXw2nv6MjA/8VLx/VXUDP2G/Tp6KGB2v37Qf0b+f5FQF6
BewLXkTtOvQ2nn4pyDEfuuNp1Yu1Pur8jz40Uoobgjzur1BCd2+9E+uYw1IkUv9/COHBhGGyL5MA
uwZqkLVK7WdRu/K+5KGv9E+qg80BESChWMPxSmf8nXLIB/oZxCAuob8f/0eFQ9AKTDmSa8kN22wB
ThAjJS2oC81wsfpayJVkA7g15GlVh6BRN+hJDbtBMQ0b5VGyqW2E7AMQU/EunfSzNhC9AV7cDMqu
7tRnMESn2dC67cR611iyTQQOjP8eKAEkoSNKNbxNcm5V9nBgd0VOrOrUUvLfGNdqdsN2kiPw42KW
ywkkKzoLeS4H/Zp1yGM22uuR7rLqnEffjIPNNa4+fMoT7tvaEoR2AhTDpxfr0NHg8TGDIfUh4hmR
cXXN+eTRMnRiPzfRP8j+o68nqLqhI+Sw684wvGUcwVysVJt2tSbmm4zlXULOWuTqi5iPoZhi2b4o
2pEu1vaebsvDNxkTCk6ckosJCIN0aglVLACt5H5Nd2uyEekTKfuE1jvQxnHUaDIZncSK46PXKLpk
WJYAQxRMLDatlHjH1fZPSaRVgdQN3RUKxArhRa2KPy5sOwTj3Kon3CTVivzZWvcAUwnzFm6NS//U
nJ2ssaktei2GDL7AeadC3rbARg8+3cIXXQGDHcDBvO1CX5I/k1ZvYZzp7+zjkvs2G27VA78HvR40
ligsMqmhFvVaOFaEMVm5Je5oMJPXwMIeZNYWQQkKhcHvT8ILUmtb9SYqI2XT2uUedNu4nywnj9KP
v0maMmsi2qaGXoikBi1lDnrY+gSM7iS2JWjcWehDUKSncpEAKKDbGawRRrtmQiyuLz+DhxIw0aHd
yP6pS68As1El9w6BpOKmSSX2gYAiG2yrFt2wthasVIapU4d0V+GoIdNY+T4zuGdtokDt/VmuI2s4
Vadu+Rgif8cF+RUAQiLiaMbq0NlT+iEFLtJNXeCIugQ0KUyVGUm1MsWlHQBaA9J+ioPp3tUxntV5
BNTTbxz4Sw4zvhCIURX34+56qc41/PP6XNRSW+aM42NnxLT1CUvX7n7IzmI5Rv9QrjE2MoiAmE+g
v/CdoXxp+2TW8VXTJ7DmMWKSoVNeSW6A3NDW5IwJd34SDBFTGb+6GEF0zQHx7R269s7jn7mSzT6b
SH+4nRVQ+Pp1wlMVFUktKRJao6AKOxFEmIsMNntdF9rWDl5uNSZRgmLt5c4w+wfVs5cFOw7f/tuz
UMGYF+H7dKLRpebI0guDF7vT8ys8cmhsfH7xBV8wsguK6wrXYC6Ugqu/7o3BUhS4AIV20UmrmaGH
pp3E/G1LMrjHd0jiUBC4ahrk7iveeYj6mARlQNxFBmPrgAlQ0u4AlvJaAP6X6XOW6D4QXzMx8y2a
npqNqc0ug97FcUANlSU3NsAKlIiQasJO9bzIICGWNwc9f9/3w0IIll2DpO6Yi99VqUhwyvNgztxd
0GVBSKOuzJYxneVl5UPSFArYUrcat9eqJdd2x8ZUVUSl8TA/GocOR0CdKsm5cLtM3uuoa1OowjUR
vzD8MkXmknFB3xtspdDrIbSFrSiuQuJIuonkgnspDeLRFTYEliHmQd9HU5RfNOwDyYbN7qsmlbP1
qL5OLY9C4cljRB9bNlJKKSIaKU37AP4ob7ecGngWu8Bfwe35JlYkAlCdS1BoGmygWivn1J9dn+KJ
tFolf0xhkyZKnRiLAQMST+qE+ojrkG0MdW95ioAORGdRyQgdZhGya+hK5Kv6bqHpQGnurcW116Pw
XB1MeiF0zO04iLFUs3VwGxispCIRDnuroB7pKJ9aAdt3oOA+6PPuscYUbLJmnE+FrO7LwZL3w+97
crB5KhIZN/ZTidNcGIgrZ9MAXD8OlJEPz5BdjFurdBHtn3mLdJFKJDuH7jWo7Gz36nCgh0FwU+HA
NDn/F4I5+z/ol/FdZaz2C68jPRSzxaDGK/kOM7AlrhAM7x6uXd0iPOgxHa63jHlL3OHyzfhKqCF0
P70m1OU5FfWlW5rpLNjPv6JNb1FNFSmUTI6LFT5n1H1vaNUmZWdPKuO2g8LtXkmU+rVAu0FmN8EV
wV9ANQmHO5/6/5FubFL8mfugwnCWc1hhXL2lAtQqGXwWPLPdcQ4DlUmcQ58YG8EORoj32ki+MJMR
BFzfF/cF4ilE/xHTurJzj0+/z2M3Dr3BMDey2qrHW9gFAAvvhqHsh4SaAaTRpYeWdwlOQ5fnNxoH
+pB/u7F/MvwNs0oSXezmMH+IZousmiVblSbyJ0qbKr+cJ92nWEk6YgqNhcLL+gfFGcae0DzsvnP4
Ube90aMJQat6gxTPDiHPmQHttsEFJDRP0kNRHmLf/WwuYaCfYb5HL75DP+DY0Dy3bdotnouuXzGD
SLK64Ck02Yqjs9Ew5OGVJ+7nzhaY0vzeQvYM/ElYNQ3BZAbWNDy0HYTgn+9anP5UWY7Olvqhv2kR
KvxIU0fSHtgmNsGd1TGH8uB6GcjwOc4aygGEZxMF7xYqLgYk7YL9mx7nngHvQFWRR3j8zN1f7R9a
62bxfZmbjhMt7nVJmKcUMqSIPH7J+G8H8xtkS8Zn60s3tgZ0WCQktyNzcM7zSF7PtqR6QbN5qNGU
ungg5ix9LG9a1W/rPyJ3LrG414gMyNKNLb4tUjeVmNl2+htEOm4wNDMrrJHVUd5hXHSc0k0/WwBR
sNRKhvH+PyVb6GFqccbC5raurIqVrVyKt8LnlxNJSX+Z+pzGjwCR+1z4qVhkLi1SRaFg/zJ89U2Z
ArIAZNEjVGzjsY1Oea2wZ5a8tHda7UOTwkch05TVDtIpJBH9b7qqcgX8U4TPxslOfXRK6WGbw3mf
OcYfk2xY1yXQEwCFUgoBRdeBYMRqTRrKkh97VqWzPX9M4noowRSDvy7w9R1HQdAnAITBlCnSMPT4
FEKAOZ3X8pS7pM5oA0bmOiN7NbtiVoanZoNEZEl4WNOf+paaW58NyRR5e4Dtr3vdTkFAbfQHKX/6
1inUVFdFtFDrJZ1syqKBmGJnXHrb6aWSU+Z4CIDp/HftBlBmhCs1X1bf3eRZX4xNT1QHog/fs/+K
TfwoDXTi82G6rECrU8UatWYnU1HREGNIbJGNL7QO4g3O6/iwI6HT7LARz3Xf+hDkNWgUQpK2R86v
lxz6CGjc7gsRc/cY9A8do6/pjKNKNOsLJXEt2bCvXO9NEAAOQv6lH5SZE47w98n8vXfCM5DTUkXJ
wsmim+sr9IEsa5HxCO2lblH4+IS7yQAglprEzLnTRpk1l5CAt9VIBV6y2GHoLo1JlB284YLt8r7U
kMVczx1VeushpM6ETRma74Jermq3X/kKRqSrKu46ElsRxiFW3HA4bmThRFb31KA4xEn90Z+HadXo
3vqa8awL+CbfEFxL3cG9v1utfnytM3TCcAgAX0XRLwWriVRcChwBgX5Y6TppyNpce39PP/EQbaqC
bFWYaUwSwetbvegK3r+VjHVMHJcwK1zHCKSuH13kEo7uRjaisQG0laWZ4EsY4JbIJhu+jaLCrPv4
viWOwZiIOo0luA+2vyOPjTuersui4uyxJvAVGqkxpvtBjSeKnsQeV6Viis+c9tK3kNZylIK1tk+v
lpimi9Lb4Hxnj6ItTYwBSmZPTkhXvNXTtsm8ev6rlAgX9i3KUOgzOmjWfxJD61qH3d6zw2qw8Ip/
NjNvwzJEzzCNc97zCMvZiZCqS5DzI+lmOh7iEyl801lUnQzbI1F4lRv0Vm9ho2sx5pC/4NiL6lbB
I90phwW2WLxREFj59V6vsUzvH7nefVgoBMU2nFDv8A0GoRzElw2vL/FdVZNzSFyzZlPMT0z0LhS/
cH3b0mkfg6flm630AQthYtaN2ImNr9UICUmbOibnR3y1z/mAZ43ou6gVOBQzwdM/isui+PNLY0Qe
xGr3GMol/E1PzrJVHnZQYIWL7L+mi2I7Acv0McDR6Qs48iD5d1TWYx8i9HqCWublmqVhzrnEJZCh
qYsZrygET8o/3V849meGZVOWwML7A+rdiECtchWCvrPftjoku9pFdM4jUS8/UDQGDe65atfiyPZy
hmL2YIiqhTTvcBIzbmsE5d+LKviKUOuQMbVkiAaKP6+reNJW+6pyWcmBFIcCkm3CZTqK20Wo9/XB
frsNz1qOolUEmgXG57oKEO/nVciFjqc1IDsX3ydbVNIiroGbTu7CbZtYKX6BhWzhKDj9vtU6Mc9w
2WbcnXjd5nfJSUZEDmZSmWarGDRmiBgLj5czgvB1w2cBQ0hOlN19T0LM4BwY6Y7G7mWIMjwKNDJ7
NoLzrK9cj9szIfdtaGP8h5TQaIwkLDnGpeupecw3bQMchGigHWwHX8s+qhaT6GRVU1DHC6l+HOQ8
h77l5Jz6bkNQnnPSsL8vblrOrhvCoXq+R7uEuJMIaLdJsZYzXxCHin2B496c+C4Hq9JZGRlrr3jK
P2J6KQ3Nh+hXnQEGzLnE4tZzF6IYF96baf5vtcecZwDmHQlmcZKGgqZxLiyZlWf51aMpyj+68fLy
vpdtkaqfQgU9PW7rZXe3QwLRib9oynO0OuSnIMjJ8X4ozfTzSLhqfyenSUrGHtV9cdIOV110zYvX
1nVP160EyFpvac+Jj5msnQ7Jsrxkd4Fiqk2KRpj4DweNboRKBWckiVITt4K6YzbUcpcTSwQXaCYZ
egA0X3ZjQm/SltdWE4pKXlwOL9YVrtLGos47YA/fRGONIgpSPFuj5MbPBZiBbQCr9vgxK3Z9PWWK
czcd+fdf3LmvMf21kbEIpLV2Otxc5MrcH+7iwmGWiq5xQl0+bLER/5cZKeBHOWtpe7wUP/Vej7xS
+NsNxXdUGzrYjq1T89cBPnc1TYyryCiwO9IQngQm+GssrV0DzKpkIfnHudco1pYzh8dJv3Lgom0c
S4S3SxoYv3bs+Vi4RkxG6S3dlO9V7i/NsQweCvUa7xIJySOH0cS4Ys8EiBIEkLIf7KOaA/CYfV7J
D2NEe9ZYUlj62HHB3uCGtirobAR7ZEt7NPygrLdAwkVYSKGntpPr4J2YZNXjHzML6ye8cr+BS4k3
4DB1TLd4hJqj8RhlojrD4kvdfmTtRk1qZYSkX6EjqEnnLqq6UecbpntlJr+rCmMt76JtZJdiQoGH
dfpCw/1l2A7aQmMZn/H6YBMxXxRKOxvggRQmBNUTB6u9TTnpC4I0osgbpVCIwhf0cMmShrzZGqJm
+c9V+u9v8Udk8kGgn+dWmZ93SBQr8UQxlWUM6lTEkMeXicatiPys0sMzkN5GkO7wX4ehXcOJtQxW
UAquKQ83WZR2nJFkF2CXwZ/Cq53SprHFuqVYeS7S8IrY4BOoUfWfoEyB+ZDoY/pqD06JuIvHMkzO
AyjttVxQOz7G+BD234SQa4OtCG3biGinxTHHNn7eOGUQLFcKpxcZKpQypfxjTQgnOgs7PBcMJuZY
YazF0s5azi2LYOONKl/KDT+m760LMa+0N1MBwVD/WbkgV3cTyRZ688wC+dfxVNg69N015vXSe+gY
w8vAhxV2P9qOyg7J+BlWFX2YHbYXrNjrnnXZuyNPD1aJ3duanFA/Y4Oe6nVzqlhu8cEKqx5iqN3R
XBWDUOb3ZUbrY+kKD4y7k6EtA8W0GqqUNef70eX1SiHNoew4AgtgRRsLz1GMoBVIKhRSVNaGcdMc
HvudjA1pnW524XtRIVNabbv9p92sB/wVU3YP5iwYvoKm2Pu/Sw4U00zgM1PP1snMfar68E6feZ+z
cu3x/3x9LavV0ngsIOiLjIoBRytpxVbvFBPp3zeUjEnsd2r08RrdhqcdybEKd3bYrNJc2D1gHaqL
4UARyR2V/QKqqrRo8Kh0wJSQlWsn3k5Cbi8lWMaIdaH5oGBaDrbbOgj3wmUWEU3ym2ZL04ne9UjN
1Nam1jK0dLPw6a0QhHwDkTgSxbR946BXErzeTQgYIywZFLGlgVUWM2QHGM/lzlus21MKNOBZgbBA
9564Uhtrs0R043mezjS9XpM60MazrnRZu/GySuWQM5QSdwVI7umKbNkr3cdiBxzkZey46r8UAUgI
S3XgWxQve10MfsLVTipccZ0tOI87ylqB7J0SzlDvErdEcrUzH/V0EushJuCmpKaFs3bP7qUgr9B9
UayWnzZ+pGYnw3RZNQexckv0jjJdA9o2UgSolByxFZf5P2oNe5uAlnXRdhJfptTkQMOXNyjVrwUc
2dnOnnwBxJyzCFXWqBMVBnoLMLDj5kQTNhnw/Y2vycP0lPiU5kZRO5FifRU5Wjdbexv8EbNRKnao
QUWpZuGNDd5pHdtIest+fs1+WOTQvZZXhLHtWj9r07JyUOMbm17QiYt6UPa4CSg0LZO0xmJyVoFl
Sf90G4WyWd78aqeq3Vw1X4Yt9pgWzGATmgzejZwAFshXMgqj8hg4/AV6BnXEtSDxiIlc9fsJkjBN
wDVtbhLX4201Kj0s2N06jDQIiXAYmAVcLyeiE68BUU4/v9lKhS/jydjzd5FDhd4Iy4OytNryWzIX
SULTgzveAnRnvUJ+ktwpWk5EzTQFobF+PascixZl3eGfIGZZKY5TyaoZVINOPy/mo5vaX8RwtMAH
CO/GbXYVOuv0Nom1/wHKwzL51FH0UBaPT04mG9r8bdwPb1x29wRdB7/xfOqm6PF90sUY329CCxis
NiakQdv91ZuASsvJjpE7Ua63+Hco/ACBZL/1YQB2tboNRZyNprnZUfE2hpmBgcJt3PpichTpkTjw
i+uyMIXlTj3SqLTiT5WMzjO8298C4RGmZQZr+tBbslYjJ/iLVeClNhXrGbl1T+80PVuVGwiGjNIR
fTAt03G3A2AjP+0x1xtkCR62eDFtzV+CtPpPV3JDuovNv1cd7/fsRPrYmhOTBxUWgLAUId0gJVdA
A4+RaZJKIh/VUnAlJEsuOkhw1NUhGmUNnm1ljDvtj0VaEMa29zBI7t+yEK7MSdYqmChMIf5XykuB
cqu19eCsoMaN2WbzxYQMeaqazcKIsUFyrn+fTyW031KS8twOqWW3fCYWGF3Ryo0nNSw+8uYV4Z6O
vqOE9yVtb8KpqoT5sZcOtZt2W9gI62LbpaRB2Rcxj1L4sP+YfJ+A/CJOcfniMaZ6WQlFrAF9H0/X
Km1Fi1lv6jRq69VsMmurVEUkLMm3dGWCINoomEF1p37b5w3RBzV0s7aHM2/24qylzztF/T5CHnW8
whW/6sNxVDlizD8R2ufFo89sTHNnQd+Iuq0iyeh2mNxAndMcbLMBxyKMtyDwkJ2dKyK+QYvD3HU4
Siekbse2N4YfWXgfViBMUbdL89bxu+ybRx7V42UR40OpkjjtwJi8jKKaTnBiSAMdtITtUEfUEujN
lJyULfgHbicipFoKWpQjQ1jK4mAxb6hoO2c6YFmeI3p8jT2CJgKOmzBIekDSq/PhE97W32F5Kpft
p/gO/X0V+U2zg/pDIvLu+bsUMk9m0knJJOVc+PvGP+5L5+lsrzn1ioTsqyIK88xBexyNAvdjR4gc
3b8v9v4JICTGhS0DDbU9vlq/Jt/PpRSHtFb3gmEOvarqUZgTdE5M5vnlT/HoKryymm3JatQVniBd
0hIzIs3kQsfCHNhfeMCAfqOmYFW1mamBZKf/ZzDEhVfx5jPeb1Tr6RAmjqVApQkB+fJ8HfOZ+eNK
rKYx69DW0C6XEM+QewOEbZ4aQninSYS3p0voQx8W+cU7rqRnmHCqp4zgNzv6MtmV55nYNsHBbdUC
+ZMVqfU4ABEtPFvirUEayj6HxNsxZRdGePmBUlvei/rV96fgmd/pLPNjmO3II3oF/YonralNONJn
m/LiAqvq0zVy2GrgKCl1zus3LDKT6TkkpsCYBAXvnbzN+TlcVh/uEXN/fIXqv9dzujMkFoAKIan8
2LxWtGTcsy1GZEXvffJ9S4cpxVdQ03Jy2KKqgpMK29ao9/BY2C7w81h66FTz6CgZdEuYoXcTVYMV
VdUnP/yy9pHLrXfE22KbMay+eJqwU4tKsPeGKQgyPW0b02yHtsNf0cbI3jICqDqHow7WtVqEFPzP
OxWlcfjsUTe3yu96CA4JB/JYt8rMw5PuaXXnQi5sqTBViip4aln6B9TXqEKy2de6r9S8WSuCpHZt
NaLUGTUL7b1PFciplcImthRQW6wL41cgrmoXh+Pe48GZ9AdQlEpTDHtPHzAOUK+fRo2YsnLJbFY6
izB8gXZVqPh3mhz/X967z55BerXJfi7wsDsyGCMZQzwkeacNBnbtG7R07+NziOJJWIvCmaOwA7b0
q1roBuOzVmu4N4rgHilNAuHPF36KFY6bjRKiUJZ+10gtD0vIT2M3AYGAwmZ44HoeFNqy8NgqMW22
xbEocO3I64ZyrUpc8mJLc0kBg/DBX1ge2BcbSNyBzmYsMP+gAnlxTiApukzwtJRcCDn2dE5ly5zY
k4qu68GlQMXe4/O89xtGdBEUWHwZkEY31LunTFPiRl0UnofiiHPVvVVMRszJYVVf68gaJ+6ZQlKn
JCEGYGm83YflgLYhMiFn6xsAxDC+YCUyzBqlWokAYKAtaQjwFD1MfFWLdc5ULhfi/EA8w/eCDx0t
knBC4jhib3tVQGZAlLXMD42hr4mQfPZ+CRz7iaFFiOgHZ97iFlqNLe032yGNHPlmybApxNQrRyHR
9swHvAtl+nSOBlNyLxRYc5KEe1/54i+jNg3FmMsF/cDw2bzRlgYyyS2jVjnIkI0pWIgHdApPU7Hm
3/2cD+iX193qRIWUQFbmnUtSxjgHC3mURp7EnchjxNy2Dpg3UGJGcGVr+pCOlzgXxxPLn4jt/zBG
Hq8z+vJeiC9mkv6WJP9/YBbwWCOcSvGK2gOwEyTq0XfZxkFaoQKOQgl14S/TIoq/9iJJsiuvmLPg
RTYTN/styhA2UONiiGTBcRIOY6munBKsKefceOgX09Z6BNyIjWuZtoXXNSv27YO7RadmcnEySWSQ
2DBQyu57a53Sg0AA3Qz8DU/ya1VYg92po0hN7vy9rU79QJ4cxNvDSNy2vODREgBSaDJioKfhsVDD
y2pjpG2ndtF60nlitG1eJS/DtmsPdvGvODqta44IkbtPzs5GZj0z/PnRFuThEx2VFUh5Dm9aoBw8
UUV+Psik6qY9bLjKfm9cLLNsSdlMEerjNC5hbmdSYzdHlqt0GTbjlYq+1OprPAWJx46UtVncaQCT
Kma+PojFCEuqTSJzLMf8j92a0/C/JQp7bfkMOS83lNpjeW/3Hefl6dMYzyyjrfieAOcmhkzGOKMm
Ru0bMY64lhuxeVNLXJLTJ9dWp0hBjiQFlG/YVjceecrAq6qVZHuhqi5z6Qbw5qQgxpjuxkXA9DGM
Hw811ZY1xLE4TH69Hca/4BcDOfdPW6gmJGWPjv4h7Oc3QSDR95o4r9MBHphwqHiGPCTxLTJfc13P
JehyFBs4y44bYgQVhNcokmbmTF1w0qNCQ3vmDHlTgQEu0tA3ecznZe66l+XLmXF30Y7Rw7LDaCSP
FVR9BnfI18YnGAP+h6m7bvSLiKd7tlKlURC/tTXEDnWhpULThheInii4jei9nbliugXLI+LMW4Es
4s+2YHsg4O5GXsLvgXhNgC1GfGq2gFEule1FlnBH79yejTdY49vBDWXLYta4H5rU2jQnorlaRUsC
QBmdP3czsOaA6YvMHhTpXzGvTNpX61Q7uENyoAelJLrfAyM8aRprSHL0SXVh0F/FKomN1xueQ58v
4GcoF/98/HKlFB6+wC/Y7sRwTLYFe9lYU/lmVY9V8FVIeRz41v+RUGliQe2P7w78UIaCXS9+SpfN
zm4vH0R89CR6YRl1uVvhAWHFXLPzwWL5Ejst+k+BBxuTLXuKsjwdGE27vtOy6r3QrU9KaCB2P3Mt
FLGvxL155q2jsr3FSsXoAI1jWCAIYgTh3S2QTc4sw5umXXsIE72spFMbRAm3b3uHyy9KbaWcIPAC
iqb4hXW3MSl55KYmlD9ulasTHixNsoZqosveSaPDdXgin5EXiPmimzdvHAsMoA35YlYqFK67p5pv
giVBOALAsUer8ms2JsYGxpBTuu6gUK/c8Santw8NRXl9hMRBM2PQQD2LL4xlEEH32W2Djhb1CVqK
diyN4uQ38fnDSbSZO/39DUA9Y/s7N6jp3MG1h68sujBJOAUCj/n6gqEshS2npXig6BoUDOvd0FpQ
gXVcLQZX82JBiuQC6nIx7xvpKj9rnvYkP8UTx8GUHI/arA65C77ZOX5g7aKDVPa4HWnX6GpjLfh+
1P5NfGlesEC8l0MLLp7QxkLYeqI3+Snm0c1XgY6WFone8/+VEwcHi4WLjs38pvA0EODyG6esz7CU
noa13bAipbfHXo3O52hduRSPyw1PFrhv8AFLhwN901CzcU8xOLEgng5BC3bbeCWajDAj2K5der4+
3TJ2Pf3tKQWtF7j8YmD03wD0Aam7B0s0EKSstmVTvzLj22VgN7hxUhfTIRUBTvXViO9qeKSxpy7p
nMW1qg+93upfTpKvXkQStpn09HnACyIT3Rv0p+Zna6ZK3BXLfipqwxp9LeT+ZRlOXMEv3JoPrL/7
8bAF+LyZQLiiU646Xin8S75ntJeQdN7vH5tQP5daNXRobBC/zY5oDvNlZsNYyVvPf2IlwYtvEz4b
BxQd4skCO8KAeeJrVUg+VTPC3EuzysRv5vH/5nVhKdxeSlLcYb1Izd79UiAW+DLRGgGUsXKNEGOI
vKxNze/FSeUToB88PKXJP9a6iQK2qp7isbEtZiRoe6XfN08sPjxdq9zMkCDUImAwSOccLji2vWY4
xHmt6Bis0v0KnNRiEbIGiXML/L8XAHJ8YkbXKBLM05deFdSLexKEn8r6ojIT6W48Xfbv2rrFyWUr
p99EOZpysV38s/qFMeDVeWTwEgCb8OZ2963uNcGcmeG7kqPNbEqqAR/Qg/IK4XDKXNATeb7b8NLO
G3bX1mKX7kUBcrWtFihDh7Hu57+aOUu4KPIudfIi3Qb48jB35xIWHh44j+UPSZkam8vv0XUZgd3l
KaVWCG2qUFNH+ducXEZTjbDQeHM4ypb4JI0GHbKvXCBs3Euckt8x/edtXopNED++//3WSrZ/qwFA
LOi5ENAdtNAUkaZLerUs1w5vQ/Irg0213v7VuyPG9Iv7tvmxnTeppV9H8P4m3oBdCHvKVCLG2cX4
tgVZdJOYSXAGEcQdqGxNF21UvKfl+9OGemtbnrcVtq0QeSv34BxfCZN2GQ9Csje7xrAH1ncZ4yvO
ouJub3FWapF2VIEnAs0HbZo2wdGfBkrP58PEuh64oF9AfVwDQE/qPXW5nEO8joUoNFYCvLijdYRO
22aMSkQo3QbXcxrz91BGO4Zoj9cgx//a4WJzezAXSPdgxLeUqKL7sOPyWDcIL80cL7UHhj26WkkP
LU/1u2pgSCw1wC4PQxZJCmRn1FUpsxjKsAZIaEYa9OYl7lzHbkCnKJ1179KEntqZkUfUVvxGgMmD
oSwVgzZZ4QMavjERa9dmdfCQ4Y0TmpFgdQ+OAksJt5EtxBqKdIklLDzMF6iPI5OlfGkarTJhHnky
eq603bEwN2lO9q1STla+uIFIGVBgq3kjfEgtvsFrV3ZerrUGbUW9tLgw7a2V7LImklX+WScR3B9P
UidGq/wrlg6t0twyqccLyJss9k6+5TeK+z/dKlPQl6pbtwKtJciXU9OJo6ib6XRuff7PUuMJH2Hd
3Q7+dPu0zkxmxN/+6MG0NCBeuFsiDF9b/Kp0/rW1jH2lUFlFWBKUHRtd2n200eISqXVnYdfl0Wbn
3y9lxKQ53bl2w+WY0mFTBSZ7llYBwwUYUXVjLloZITGuBvNtm4hnOG20zHZ7E6j469Eri8FFWdnI
0ECa50rrH8J5y2M9JcCcSeC37uIqlDKtkZArRHLR/Y+qZE8w19ryyCgcfHxgvwI6fWQnDFZO9/Wt
zylUrNWHSLs0JIYcZLFvgUek82vOj7BKsMF8FED9Ukebvupeukzb1iM8TvNhCnvR8e53UyRR9R1k
wgObsbwoIHRpfrJKv2HWohJw0uirF/DaUaNo3Z0994twG8oxG3Pv7kzxuWXK5iUAGdDW7az2H0AO
8pjcW4k+aIGLUmkRhyzeOYilqajan/GCA0oOuaeryrLvk6LJ1lk+69BjaZvNB1Z4D/6MkwOvyieI
1a4idfutFXPTY1WIw9tHTJQ0XRE2qaTg4NHrVC2hN5nJlZcsu81jCgtTX0yXf9bSmRFhfRwNhp34
Tz45WNceZ34DhHbENLuIcpvLBvlnJJmqD7ukjpDGS7bz/f+ROuALmKSukrFPtrbkFPUYipR1n/yk
nUYqEHs6TxBhePnd+5Qpo+f3VsVMqZkC+cMhUy+//ehifbZ1AWNJvLWz7vg7lKt53HM3pmXoVhST
0AStjv7xCE/+KN0Yx8K4lmbk2xCHLHNg9XbOIO1kJdgb9cCoZepcMzQNHNHfWWfIfctccsGWej26
TKySOtY1PDuAzSG/lVxE+jEn8zSfbfoQd0A4t9a3IjWwUQiFG+CjPECYX4YCeaCUQK42F22WKhyN
C7X3XMciyv9+FvJhZtGQNVWXwaUHUEqlyBo+UmhtXR8Mv5fTJfOPGTsbdaypiySe5L2Zx4ZeHXP8
y51WtfDAIrwWEOzBfRDRCslqOeQuwW1BGDUWiOeieVUcchQVyb+SJ0tlKRXNZC7Oi7LhNIBfCAVm
rJ+FCWdc/oCvxnXw2pX5bnbDhjVZiSKlU9OP72HI16ho71c+aUDqJ24zPVaOZtXW8XWrVp7SaImE
28eQmfXw0GGkl1IB5KsuXpqiJdrz8LEHj9d+pD1Q3KrbK93bjrDC4yjhExuRndktmXoyDod4Ym0F
opwGeiriID8vzbtPSzL4wqS+4IacpJCqvyGbfZY5eM9GFmM4QTnhOVELPDpWQR3vSjKXUt80shBG
cPrXYYYlPwYgJeh4KiVJlDcqEkhuSbKjvOTNUckRfU3qzrkAVjepIM3Fltgh84ik4OTlVWGQfoyX
5GcIj522LFp1I3PFLFAs4RMU1yANW/Sfg1oCN2xg9/m7nmrj7f51RVxhffmAnRywPULDX4WJb83n
r7RYh/+PIZEanSljoFZd4pkN24452139R/hDPa9VDnVXi3hOg+LiWBu1qiFCTEnR2M081RSznxpk
EXZmjbWTA0lJAkw8vhwn5CamtYzRsIDJyYU5bENTE7Hn19b/Fw3E/gSweLQpDj+JqkR6PraV9dwK
wHeWkewIMjnLhEciPiCWsLZg2d8aqjntlC6oFT9Ax860XOiWHaa7JtkJ4rkCzPmkOD0Wm5okvaDf
IWbQj9Z0e9r8RUGLI8RyccskmLXEJyxYDXTrxdHA6HBusASgtWr4jcVuqWD+QA3im7ZEzlhy780r
5A4lIx4tW2GMj6jCLxatFyVzL80W8pBR5aU6GKvPF/zQjAERDpSWHnRTHGM5GoSb4TrtsHMGk+Ub
gtyO5Xy4H44SuOhgBogJ7psokbmQ0xHHJyiBgfjmcjgkvi+b27obK1Xr3xee3MP/k0fUBDm9iJvs
jDSEODyfs1+WynJ2FsP7e8uodu1XrKpXnUFdIu5cVoellfZAgG8DefKMv2DGouxdZq1V5LVCKbpL
sjp/Zn9b4+FEglwxkGAroap6I3asuCZ7prxiuzxCdPgi6Mme4gzw40VljdmxWCwhOvmjRfNhvh4a
/7AZAUuldevPaA9vGwEiJRgwAmNC2TTblmpr6SnVmXrRaWTumfEEduvPb0ySupneMWN7hikIPwhh
429mk5IZd00cap68zCb705hpaYlX/uwwzOPC2WRh5ZTiEA279hKtIdFwVaNe3oKSe23o/o/Solz4
nVJYRXXOtvsJyZ3lByzLom3BN51wStLa/fqbCQBwSRFYPotDNGl0Nmh8jERc8KP6IMhHT4AfsTuc
RBreSNtOQGrigoYj3HFt9QMK2nAhkwTCTVbxDJ5zI87j/Rk5Ai1k4P1WM9cpSxESIXHaRyj+Qh00
l8ERtgoeLb1EUFMmzvqNcn+qYYMAlhYatfnNLndbwsq6ycCWHG2zT+0zUW9N6YbYGFRR7UFgUfkV
QuULS9aI++qeoZkVhJ/2YOUL+neB9fJgM+bPBZYvgxpOvsulcia8Deko+/GYTMU5Do5Ie8cOo+Lw
Gv/HsgxBE9T0/ZgoCNLNdnqGLrQn6Yth2UTokN5Pmoi/0uEZMTtXTauaSHhchxj4CpvDp+RGS+kT
LbPpinwGpyT2zi5FFEka6fVYN7wGGgl1ui+iNIHfJxvI4rtGPnGCn2YH9TnBWeisKJhpjAf5X88d
ASkSXYtZUDPg/jVGHQRNRj/ZtzcPuxNFYZVbd30+4FEIxMJurBbiYI0b+i6Gw12V1mbV4dwyxhzB
ReR/w9laEZYUHSddM7j086uwHjB/7Vk0ARjj1xKkikP8zd3F6pQsYDScyHMABIquL1fucIo7LALL
DY5YTW4EaYjUNaK/eDPSikGmiDvIuuIpU5ZMuY7vbH7FIa+QRWk72Tr7QM0++Zy0XiR1MT48/rRh
9CEv/7pSosiQUCD4LvuG+gFv6ADzRQ3WVQpBnJIbfJl7nGWE2vyieZlVu3lMXP9t0tvpRkkXFlj2
GEmP0Rb2JZouJDyP6QG7DOaIq5Hp8wV9grQcg4Bk0q2pMY9PNAI1+UlzjNFGV3b8K1kkmdRtLC7p
SWTvLdIYktYdPoDRjuLgis+V96tnq6LNQ6o0JuoZpl/dN2kFo71uQsRwqmSqNDt5vZRjlZw981s5
DVWNncRjDIfa15X6UtAw5w2aSFewYXvHhsvu8mQu4Ycy+MIRFMbM6sbmh8LS2JtzHXfOOM32Bl2A
BLqGTNurLh7duBe+Y3o36rC0twTEWCFqHN5lwHN0zscbqjSc1XJxVR8LJNzdTHTALnGAxDnR8r9n
ym67ZlFscCABUWUyPzI21rcUV5f63vKwzH1+fcjX9P0ACE+yHNS2m95BF2kpqzf1QbrJItbAHtlh
4mf5wa8VlKF31qXc4Pa5sZGvQBQAVuqMUWyrgqIxUGR+IFlqWnlRPGGGFP1vS89DaL0nTE62dIkb
8A5+HeFpNUMhmMtLL8272BdmtLYQ9zoaw8IkOpwxxbY8oGo3A2sa/TwUz65Epi2ILzwfGI0PO5Qz
fHOWnx1lR9+pC3TWO7SjlQQ35cOq6OUvqkaP19jtx2+tn0KpSPgnhYHcbHlRDUfgvdvLUxbw4lqt
+c6Xk3aOK7gZD0f55h+6mD4AyFbF5S3u+rJqkOm0Uwaetl+9rRO8DCgS30XXaka372vWtKqzLpGP
7qUIQ1rXzzZBZDjSbwoVvP4Cw3luiUR/0RhXnpw4q2i3I4LCRpdgj++5NugrAPZZbPHB6NkEQlNL
qDAq/N7q0wBDlHr/vzgh67Makb+1w5ieTKZs4IkjsbwX9or8BEdVT5j2Qc+ammEOryjLk/PqdU4/
egjL8MBGhmcivjJDbB/dELzY+OqkcVMSaLIibJnACrhKV/AgnZGoKrABPFjVcujUTMvoDd+WerXB
2TBGw4iixwXdkADbJTf4lrk+/zP8vFwkhC5GNgbWc6fPKr+E9A5Ent2tpiTJljEZv7dlLtG2nNyR
0o8Y0sMf8didyVfg8UwWWBkx8y59V94lskhddjMUjcuC5n3lble8logRlTQZ/j/yd/kQoJn+UghX
rTLWSxFdU7LDpjKgZR4rQEbMmpFk359g29NHcih0NwYQ72SmNEhnNzVKv7XBoMcEFfO6r2Y9bFTe
QvswA0exQUKRDM32hCHZ5Ek+fB83BpixiQ9hPBBF5ZDS17scqmV0nRIzlElKr7woE6dpnSSR9FSr
lKS2y/Ka2cj8MgkxodA9ArRfwrtmmQ9Fqp0NTta5xwAb2MeaCX/vGisl3aKifOKTYKpfVY18EH+z
tjn4H29OTKabPdGJZpzVnIN1IBRDsHg9Qe4baLeVkh82CiTuKnsjMlr5frjERLHQWBLtPUkDxIe9
m2rw7Z4cuR2AXQk0kNbPNzBtD/JLLh3VnBOWz1O1Py9LoFA2niQyqYoFlEffutSghH+gMyTRK1vT
3AAv5Wh4oGs4HFPujxRBhI4CPjT91H/fE1EX/qPLgVN93xLyop9/hT2MPuvZ3PVrx8rww64CYeqh
UQx7hqvqgt0Iu9MnPYjvOV1eaqPx7FmeHZ2wZKvF42fvXfKlWajG5Wecp29hlJIFyiahn2E4MMns
OyPwpHkomQk8k8fLuBT4kLOIR09xM9wpQ5T2AAijYtZsR4hwG4ZbV1xYtduvo52EZzAKDMlr4zrU
hJ+OckZSHRc+r5B49qYENQmqkbk8AllRfE0tKnriFkhZb06FH2lFtTE0dXltGK/TshsELo7ymX4m
2oKX9bwBHQGaWO5omUt++X4ReTPTMAegn8Q/0lvJt5UfyRGkKqBVd3AOtNq72SL3UP4hEUr1UdBI
BbTdH5OvMhfYgR6+DGlx1pOCZ/Z/QjuP2r70NYt9XO0eQ9rHLtlr8qPNRcqCcVMALBU6I/m/fJM3
klVuZA7HD6iuVTu7Xifc90hU56G6Gbj6ov/Kp+BWMq+xuG8i8ADcgL/B5sbmxo/I9KQ57JTnJ7C0
w4WcGiGLOGK82Kg1OS9uFDdUXKQeLCu7o84kqkGXTllxk/+DtMss794E6dHblcRdtVB0K625G7CH
fgRhwaLkX2NvN9ZbwK3VoSelu7gz4tKRadi4S1bBluSkOXK+pchoaCiQbyZiucpXVM2T4oEL66Mf
5/PQtDopF6ICstxRNrJEUfTw6PPmQsF2YPH+iVeMb/sG7mio8CQ6IDg+O/7YBO9yb3ZyKR2PJuQj
asdjcKMpIVJW9Ww047m/f4oL9476+o5LN39OkHvw+ARRowjUtUExkNuPmkf3R8O3Dh+i2Y+Ojt5g
dUC2io3ftbP92GJzBqEKnogrj84TjQYh8zovm1R2JRsz6mmNK2ZDM0cE0HZ60UEyU11Rj5+qoIe1
7mCUjHSe3wEdp7utXRsKkNo5mbqoj85YFKKlwaIh5aaJyXXpkW9SMh2r4LRJrUEAWSaNT2+ndmjV
qUgdMjAf32QPIDVAVv8JDmsF0EU096I0caDOQO52ql4T24Ya3ktyUHNFYL5+X1hDLCIqkw4qVVW1
T6xQRrONUQ+eY0iCvEfv8As4P/cRXDp3HbVYICP94o6mw8ThCblTWYhoUS3vgFmxI98DcahU/+0k
ZqYBTpV5EGK+lcIMoSA51PyKPEd5/LwTo51nAqguNhEizMt59g7mLY2Xy25LvYBr21sr9Nw64mW7
1VP0QjR1wK150OghZ+xBU1qzph/tDaQGV3a1q79krxXLWN4Ih8NH1RSFVYHDkKj/aE7PSi25hQ4P
hmgsjFwtZKRWMhXhM53NkUId+HYMH4drHpbAd7sGhtjos3ZIhwqaJmGLFzETNiqLj06L+JXVLQrk
d4OgMKzKS7NJhxNskIOn4ic8GQ+5AlFhxdgk36fq1WlECKbR90KWxIwHbCqPEWI0f/AQK9E9BU/4
0GDTAkzxRYrFLyMkusG+g13fEtYC5OBFXP5s9NQYArRbSnUEZZrWp3SMFg5jLbM+cVQZyKjNbiSR
sg0QyJ9ucBxak5tpZ85Cafo4n+9aPTxxYiZN6zxTv6NWpoc7Hae11hlaLSu3OzeW/pTsleAUnh4X
JJhqyp7Awh1iZDgBcwH2NFbu2Uu8NLiZp/xROt7wKb0yB1IOPssYj6oDaY2FTU0/ek2YuCIIaRAU
EVIFvyU8ky456Nr853N4PTCli+DI54ikX1jfBkKPPd9FFnbzejnQb2wZw8E4281FdMGsSaE5A40L
r+4+iQbkyqPmES8qgfFZnZ/vwZ5pqXbI0MC/95Xx0iG7Ig4+NykRU09aI8HMZsi59t9k92QEDfQK
u7993twelLaaFAeaDh0KEMq6w6vykmEEWC5rSYq2yQxcpCamPtIO34PMAxURvOEjqO+DzmiAwZCo
LT5Y1YCjf3QD9XPj6KUSm9C8Mpijmm0y/0qLbzXCUcZKF+qoEVHceCL9rjBoNFjIRd9UsC7wWFLA
7zt2SlnEjnJ7GqNeHaM+0gPp2aze4xPBOm1jwc0WdmxHz4WlP6qNi8PUcuRaw7BI8kw1PEwqHccb
qESue4BsHxaH/5ILkjAf7UrfT83QN7FdLcTpbqXgsM9Tflqxumk4X8QBTUkm88VTczQ7aqXoYXiA
RQezQ/bK7vqrQjXKtN9/WuSghJIelUvdieTiSZY2LkIHoaijDJ3Kqy8IMML7uLZmqmgwv4ZaMXY9
gQWGS+IA3q6rY0RDW5rsoN2+NXFFSigjxGHnOg/pugV2laU8HVNwjEo0m5M3jA3ruzBzCZjdeA1m
d3yZxvRrVaFsQ3xF3g9TAjDKJuAx6fDTtQu6pR2Z7niFFwSx0amKpbj702/o1bqh1vO3kcsoTYf8
XmwMH4rBKeKIXfveLAdmcS5TLsgYYE7kQ31mr9U5sxJHwDMgoIepg/O8VYbYYB+pXU7ERmIAKKuD
Sz8d9qONvXRvC92dg9Y3h5lo3ZHXCcllfL8gsuAs/KyS4KqhW9meaQ4MjbMsp5s+f/+xOEzi10/I
E3OtJEC2XdBhz0kWT6BhUJ+34FyjyxNEs2AMvpg2JnfigTWRrZx93s7aTKSiCcRnNsY3r23Ogf8H
0NFcOWGkwO6j/SYSTq+W6t3Al/J5Qm3p75amHZJM0mx4SY6DAmdrErwciq5qyN1dAecsPcbXKS1V
LV+zglTktBZzwC5tI+U2NzPQ/uZwZBuLRb3dXuPeX9Ie7ivtfMbbTHMJpKUAr5eWjHKamcbtfQEJ
4ek7qoaI/IBmPDNzdxxo/NCI+zFx7X4c+TmQ43ZIE4rtRq5aZlXvUOwFyrrY2UT3wtGIip/lsez0
H9FOP0UsgZQ+YlpdlkWAJDreVPMRc8RiRnnwfLxa0rGyZLRFsq2LlRZ0J2+UJn4M5AL883PXyKA8
X8ChmVHR57XqG6Wd/8+/dY8u/dzJZ6OMx3sFMjguvePiG6Ku98lfVbfFqJ8uNMtqI3LXcYBJBO/t
ybaIGkFerOHjVuXSw2lw9sRyVOIuCd+fxHnx8XT1tRDvYXULEt6PgP4OSqU9vSA9dnWt+i1Biwz0
S7+qrlAK6uqUlF7cpWVrS46GqrWQPiKo9UD4cwUguH8qrZ1p6u5uJFICakChWbCgaMotwe7+l+n6
2JLwuCegamfxkIBFOChkmD6wG0rnI7wTYCSo5qKW+iWYfuQTNZAj1g/RgxJDZaWyYltWSOQysZdx
hoy7gH2bDjVFZpwg1LHNvyqwVVo56tmW4tJueEiumDGIl4s9bVZEVSTMZaMaeJ2h8ypCU2xbDyFn
2MKFOhKBhY8fAKbtCoAoXLTlJPG9XMSH5m0xsAXCWoD5jiVSr1wFYIvKzTgAmgTztItALtcLoVmi
gcSyVaykffQl42xnpZA2mp/RhMa3EaVgGIj+smUoCU8WYtjtChvZWCnbnokQHrOsggI6ww82kHoH
OTmnefJ9IGqTFzJfYKo2gQrMbU0xkqBLtUlfEfk8CXNtf+RmjWrz4u58gVk4AdJW9NRxhw1W0d//
XN6XnsbPIXTIUhBi94lOwCuzP4qUpupER65l3cypwajcDUgJwfjPGBXbmWUsGc0tdeRzL41CA6lF
ajKPPvfjv4MUr06W6FT/eK7g/x87lE+TuP1L+lk00h6p1Y/TuogZdzvGypLFKVxAj4h2BW+i5mIU
e8i9zkjKT2Mf0mIRxe+hxflbNTY0ym6Gn2AW5DiFcIS6ZAToKj5wEueMBVr4OFOJnnt61miE+mkX
V6esxgGE9R40fEYH60YWE/IrCBz+dnG+O5WkrSnuXZL6V/cXLc8Fz/1FXA+3awAsc1stmHd6bZ4E
UG9PDq000wEKlSRAs4s14T9VR2zHGLSyHh9/Uk3X3uO2ZuOXtM4IQrD74cmv7EYUvK9/H+bAoXft
gyA02lHKCziiW9+OsiAl/yF/4avZuackk1wVaYZnpVDhVjLhvmb8HViysVnr5ArlsFZ+KD4OB1ur
G+ITCkLjDFJwL5Vm4bzC2qkZWmn/TnHRhTDuRXs+mgxxdTG9B1vYKx0Y8jsvPIGHW4AHoTNqBPX7
LJA5lrbaSsxyTZRKvXvsugN4cRoY62RXUn9p3palt5L27tSHTwtcFAAswYHCDPQcNusxTf4SDfZm
IVq/DnRqv29nMsP+M5l2hBGQ8eAUnfYo0VQ8atqzkGuyUFA6CH3Xp2w9ybdIJbfTc41sBkhyi18h
ZzcisO7PgohSef0TIODJxFFxMoN0uOQU1j/rA8Ev3GYyRRaJss7fCNVHaw5YGoq9EHcr7TwLHb3Y
/33jVyVX9s43epl8+d/aJYoLFG2bUqDnpVFqCTeYH2xA48cgp/+aFNopKUEdcO+qFhoQ0baTFi+o
8hJPVZDoAdiFoSTLbW7rg8h+ATcV9/Qhe9iClf1YSX3/mNxlza6J7RU5RDViUVeR4832V7BoWRlU
VPwxLDw7hBgl2V0+vZTrv+dY5IpYKTUbrJ0RSTY4YMygGTWXFZ3IgZAFVCmREbM6YvdFul2EUp5k
xpMPGZA5tD2MK4JdIVegD7+uPvKuAizD81q3vj1oatXzeAmnBeJXpESe6wmQRlonAUy6g0mNdVpk
xMTm1rPJ4X3URqm9svpTa1C2NfmEagSzNMD003E8MnIZvAoGxtuIx2EHQ0UtCazbtJHid266YTQQ
HPQvQkwDhvfIibzC1T8OdKtjT9VEMkr1fDAvUEr0nYxSOlaQk2/C9akEc2eSctLm7rkezYbYkG+M
pMdPYBME0sd4Lejrerdsbq2a9yNhWxpuAcJCE88hOgeCy6+2RRhH085Y44bemy2H4Zd4NEGyvlz3
tnfXcwdUMvuLKAxBR7/J7gI4UCOPYAiAuhaMnZmq3PYdVq3byNr5Pu6IIWlysICrPmERUYBaUSLz
ll1K1qYCidezT3K0uQ1vkR4qXB3FrHYTfPPW4THNYEMTE3PXHEaYb/CtRACdDJM74X7GArsx5w9r
ewEoXsJZZkFkuJGicVVxJSZREzCkQITzi5vSJHvgWRX9WXBGgf7y3L98Xwd5GiBJrw0ZnSP1wLK9
ncESuP153Iow13O+m4WwF+tvKy53Y9y9XNiJ1m3oly0ezRlGqyOx52K157w/RJF+ThIKxhZNpgYM
gAA6nNznifyy83UrAkuiLioWbMlzVoRrvinhD9a8feL//OdqBLoMpiof1EiPQASF4iZqEDXfcv96
OoiwPA3s+rzXIwRmpszw3sD7G1AGomO4KvU+cuQHthCd2yNV6akx24G7XlhlO/LIBeaFEZiHUUuH
Jxru+pY9nmlUK06XWFcb+Y7uAf7XoCUyzvGYIBDDDx07YsNuCEIy7r6mG5q+bEvzLTzlAThh106K
bHg1da1li58zVe+firj/JqgFqbIKmZoPSAnYMa309e2t81w6ugtdCrsFrn1IbiuSYVOMXdcxx6hc
v9AWAxHjFIHTk6Kbv/EIRZkfoX64kIPGGxz48NmrbABsNBXNi2ROKuDHCmz32SJ6MvaKnEU57Smh
wOe8NWZZ4Nl4B6O0o/Jv5NJk5VA90upr81t5gV13VOFjQgt/AL5xs+KsNhgEHAY0FYZenc03hUCM
FVQj5OKhYD4l06WVAfTWejI6AEcKKLxN4R6vqnx5w5GluPHICSv90kZ+rDxw35pnmph2ewq6/Y8y
y1eYZnEhQ4pIYPH+EkjZTmnG3gDRqnCI1kij57iUje+1MbylVEyL0f3nk80sLeALBdaSauiWltnO
fTr1idRduZKWTk1mrjt+5LjH9FiN+dBp1q0HvdCpQaTeRzCuKFP20CIB3qXcakaDNavP7rehJpad
L9XRCgvp/e0ol5RoGPgQw9JVk9Glo2elGOj4BCp3i6e4JQFyu1Hzqj5E7IwFvFho5/r3w15Xobt7
abH06WbMMcBRUWtuGXnJTFyyQ+Y3qeGxDIsPT8ogVJmrgZc4lbVyZuQgGwyZ+G+8ZkLE1Bm03jeS
bm614Al+xMqcFsppua6iQhddMUT5qlVtWeA3z3kBygRBIYDj2WFpf3ZpRgeMjK55z8I3gYb6R/Tx
i/+XvcJl6rST8tucOHOp5aTvT6eugg+FNfJyNlAVN9ku8iifF17EO29mtTrj9BFW8Andn/uQeQqv
XgEYPTXmr/aXeka36K4HJUqG2nlSahYgqjuRLg9MWLOmugwRcapsFYyglpk3wkRRy7DiZFtk8tWU
WW4nqL38J4NGNK4XvKUamauTNQFRRfJy5fUUfRdcP0Hi9gPEup280T/SZkuq3AgOowNrq9MSC45Y
8cNR70ZV8juKxuIY7pPXjKwtaXXdX8sCMsoGuYpi5gu1w4OI3zrE6C/3GjhTw3nIJ1qP6ttSBoCi
E5AgqWsYhnq87az78PsLPQnLS24yLT28oW918uNYO8llx8IdE97ENOTkFWWHHigZXiY2u4XLNQZl
kLrAj3V5Q2rGjaf6v4dol1/ukW5jkLXH7OjJYsABRXUNC0WW3NUoDEmuBeio69joFkMAjwPFgx1q
+TGqB25o9NP7GxwMAQ9e1OAgkSuHJZruCJRbzpvtZEMWQBVJY9pGm90nkPPmPBD58xkI+1SLNN9j
lf9SqPc0iiKDX3UYxGo6aQLGCkU8uHPcpp4m+c8VKKmXJkCL9sxJGF3asmhPv9TMHD+k+LgW6x8P
rHmr+z8Anqu9bHEM0G/GNzXbBAchfyULjR+5eJxsyG06RzyzmCVKJ0kvzLuOoSbPg6CDGq0ZZys1
pvpkL3IRub4K1+KQxBIet9qd+Y2QhCmbANahiIxOcmz9MvmkVqKdGNybM/hYIwRsTyeR4Sc18GA3
NAUXshUbBXykwxFtzUlHmYxXTXvUFtTi4QilKOzQsnnW/iZLh3T7Jd0NSUMwyHIZ+s60Vr9BZHiL
O9IBHlugmZ6ZDPHLMtnqfkTrcjt9TrKzZyPkQ6OtoYNNV6bGHwh4yqYIJjB3/doxEZTiXhALj4hz
xaAHj1YefGt2kS5ZG5guRisBmgo+KBupAxiISlsBMpGuyZR0L032VB/ByA4Dhh3v3cLG/Q0C5aoX
jpXZuuvN+fxXXUpUx33YFmHSYD4CPhvRz6cit1oQ/imF8p4pVuyg4/hVB7B6mgSdqwODyBnE01ZY
fURPWnDE46ROldYUDJ3cCnqXF6eGa3KHcjii7Z9FVv3wVF5s43ZgSLM25k+nTjAxXLP6enlM+m6x
e4Ij2+2DlQSLnzQNUPMEGQ9Adfsb5E9oeajhqmEVUpAmgLuEs8ULTJdfF1ZAE+Nx3Bt3Zr1pNZCv
X1xEPl7u5lQgF/DtUdchEw9m0L/Vo1l694iO86Zfgqr0SI8t4+YnfRRkBmjPOQKEZgJeYeP1tk8t
uxrqsXGaHstAyGJIrKDGsGv/OhHdPi4GaOcwpzBYPmWPUWRKuN8Z0mj5eLvo262MYPvtdokMAUZc
AZOyKVD+O3DZwwAbieNtN0ha6181I6wHqLlLi5zah7CYOciowx2Hqq1VvHW+Ddg2D8KGUWBX5NYj
H5Iz5H4P4qZ0Z03IB0315EcaYxJDwuDQySKE7CcGdjcJ6MvByPWYWSeGJV8PSFspOuO6rbdm0Fpt
COjBRFouBdYa4KgJzW/5k1gJTt3RYYDCeqBK3BOrKGEIt4fYHC7ASt1bmLGxYpcE6qg0yn6JbLH3
C8o8BJxZfLoj0E+u5xWX1QXJawfloNaNFmc2hD70hMPyd1tTuhcyOmuKe7j4SdIgOQ0Z6tGHr8Ts
JOTlzvI69aowNKlJoGqPwtVQECeJ5RzMd7qkjglPEaku+p9HtUoNHqnX6dyl/ZeQwM7AaNHfGAeu
icrfo8m9lZMHuinZmfUFZuA8FlkWh7yA/jJI140ycZskGskTLeRO20aCGwKOQ8LOtuiMzz1VQnU/
gXYtADMR+L6/x0bY1gBneaEIkJ61LzQtWHinax4KU88eYrJiVTpWHbY6Q+nnUb5gIW8M/9HqLylM
h4+b8FHOM2D5PPEtgWRyOEgZSio576XJzdVW1M313pYaLbe1g/Rjvtj0IodBvZTrCz9p+KlaaXme
v3YsJ99S+cYwilowMdv/xVx46fMV0vdFjtv1KSuX7lg7q8OqI0kqbBq5QOzMMBuR51z/+Ngw0FAo
UjrGdVeBPF5iRbCBiXLzQzCOLdB9V5IBFYEDMWm3WDzfAAdhlMb2mQBJDc2CeIglCfoGoCIUTdfs
TdqcIbQD7RNRomA3q0HAY4bO/Wkaln6AqVVDUbPARieYtGq/tDjd++CuNWZcNYs7jhC43k4HiyKd
Q50C4kwpHLvysn2EZ7R0kO8ZQEOsMLCKhFxEF7p0RIF4aYyLXTFFlMHJlvL8rEksLQ9YxyetVGGg
Phm15yp1zNnNssfqJhFtBNsoB3VgAsAaXzv5rcYty+K0bpwyzzyE1egceZ//Bj/eQ5tcFERgjVzY
r4wHRTvIXYX2sjQh69yXADbU44e7Mmh6i95Jy+gx1RvSgikcoVsCzCKRkCgYXusLKU7echFV9e+x
AgLMk4E2uTqJsfhJBv/sdCiOIDlQ2b+yntxWQvKUrFyy+8I557hn0z8PZ4weuQg0NVKH3gV4g8iI
GOvWs2sZP2i5M6eBwM+MXAWTIChIXyH/RbPNl8hia6WvnKksyAWaAAVgtGFA288DRGa1ccDO2vJ/
BF/71ihW5Jr5CSm4blaHGwT2TI/0ZZHB9rbiRCsh/8fVXqYnEDciEv2yS7hBEMZCpokqHABCV/64
V2YDTHkO00sCfYhQt1vr4o7aU1Tar+GWoQsLn0IXW9e1Sx4p/0dpe5ejKg/50+imIRS0tGEsdLLj
TjShNjmyHkLwrQDmt+EU0txmyZ3FDWcCG5mVwYldORC5sjvk0HCRK+kfe3+ebvzkh/bwMbEHzX3x
xORuP6HHIkl0nkrAqnmxfM48oEhdMol7OcfhWSFoI4LYD2aVkU2XnX4ARKV/y/wt7LBIE+BEvEgu
Biv5rBc868aDOpeR+9BWY7e6MKwtKn/7LP54HEeCjmKvKsA1dVH1up/Fv5+m6Munx6NGUBfpmyz8
NN5GL+0s0xMYmZFKZblFcXudE+MWiWyCNus0WleO2DU45X3vEHNX2v0aIVFyFiZVV3aizZYWgKGn
wHhVka2M3FQEElLhlutGT/7yW4pnB6dCUrclOrOCsMDgav1r0XKRvhdb953bbVVCN5jXbYktLIo4
LwENyeGds3+lD3Rn67kbzgLNOAJL1ymwj37CFUwP3hjAEqBoRx1JaW4gvkayx9apTGIAsMZdQhEG
q8ceHKViwh/uyfpW/bb2JiOtB6/4EB3mDDOwJCINw3sWEGmSaQr1jn7OuiQ/oQcOvSkZYs207K/Q
5INlkC9twWdGD9iVdQlQHeuGADpqTHn30qSeuLx4poFlRPGg2+5Lo2Id7/zGnkkZGBRqt+gy4PTy
ywmsL57cqGA0K32cUoG6XQPlcZoYP4R/t9esKKDaFR7tLkyxWk3XiN4WxnCB76Oc2r96+g52TrvX
kLz9v11uUms9na5xp66aJa1lGKQ8XSBpABq3gNYBKpOsLWpr8es0I0TkZ7/81je338DNAERx3kw+
nh2cVgOlq1eK9/0Jx/VUHrDiehYrBILjt+Zrnrm3iiDjwxR/fGS8RVZdfswz4e4UXwQYmUNEFOK7
Rh5Cm+DZF32aYr+batfX0lTPDNd/Q+Ak9jQBmIjrrpLOtAAK9Hs+6VTmohZjf7sSm0Yj+1dd1siO
+OsvGxTPC+fDPv4BTndc+PYklRJ3/Nvc2xrpv4aRJNYYvazmEMPDZ/4YcqoYOmJm7zGzOXADNOFn
d4VLmNpuSbyBoNKJ7PPGMYqKJ6c6FgJajYH44mOwNiataNmTYgkQ5EkCLMB6Me6HS41Cg9thUdwX
Xab5HvsmjfYrXUS2yn6tx1rLkVXs7/njVGve+EH06tnjtL2ZJVDrmRvm0P1JngkUJZYmz5di4LGm
i1oJ7HrzHQaOsd9LgmUwti0Su76v33u6k19SuhpCWkAiv7uio3OiRsG/1aoePUid0qckd4fZ1NOe
xlHhr7RZLtGq1QIlFu5qx9L/MoVK5oldeMfUEqaJ/EcUL1Fo0qtEhcsp6JtX8uej13nC7SSSzIbH
qsUk0ngJVmKHieip3aJhzD6Q1CsAQTwT1veglBQ70kKV7VLpEoqMX4mkl5guSOt0Pmy8hZmDy4L1
rlTLq732hNqqvrp9HtA74xGqIaKwqOvdvA8NqIXI2NSpmuHHTB4l3zmtEEqGStoUG4MivP0aPgwf
vY/ueeEoRLP0zzaN66vGSbupe5goNArGTM+DxsCjgUVN0BXer4FTn3LG44J9mWtPHwzxZihp+GCM
2fdnLjp3tiU9QYCraWgKuZQLXp8QQ6CY3Gs99e5V8H6tnkdCda+nIYC2jHnFIk1kQDKnlwN9emra
+hDAdtPP+R+VR7vaTzsDEdQ/5RNeSwIwXW6PVVLhPGLc4W7eHJX9H8aYGco2SrA71IQKUCWGK7lL
h8Zlk4O29rTGJKL+ovbhZu9z1YjlSKZFs/p3WH/sFvQceGBBd8IpNOaMIG3fuqxTcvSOqtdX9Ai5
hvONejyvfCkxuOaIeIsRLh0nPv0ECUaKnWNTMMBlBl99LCXezk3hvFHl3UL05dELv6yCwlw6ffH3
2g1mwwNWxxEDXfJxhYo546bsTX8xeZ8agYJNYN2udYZmJG5MIoDZcW9G2EqnCud2mZ/2dilQBatx
oDLiYK2DssULK3WMP9C6/fsjaK3Uww7unApHtNG4kKbCLqGs7ZjyDBIkoNk/vYdIq8exjvbKoLeZ
8d9/L6waquY5nP1Q6+flSYzhzHJ9lctXIFeKOHyxxRQakxt0+VGAPKTc6ImbuyLY8bxTmw6s1Zde
PPMDhJGIW1OEVpV/P6gh5Ht9udW7UjBeCf+T/8tsFS7xHfogR7NczCBcnKZ6j0Sr/M+DDmB6cfq4
dWahvuy5asvFCY65946yvZhkq5ftRLqCwp52xXq/NhytaH4iLSkN9U70dw6NZDenM0L5R7F4tyKT
4f46eiwZBArbbNjf5VhndYLUNGQSDPLruL8gFFdeSxqo29LDs6WDQ3Kiepc8yjvMunYYUoHggaQf
9hBPamMP+a68v5EcPYYON+kDukyubPM1TzxtKjU7UDSBTCTG6KDLvRy6/OaLXVtqWxNg2AzHDQco
xSzPQduiI/bf55XikknDLNRWZWd3BSj41ITnaNY6/2Bz3NidDqbt6hbPfq79guOnpUHmML6AEXAd
5siQiFzuremNxvAqKo2afBIMA0pueClwCMfZjCY8fTnjOC1doHeFB3ysW7HBI6dhUD+nAtTG5ewz
E6/qCMdUHmGJ0+2d/fFPI18YVe0LQML6rMbY3r2v0kdjqAcexPoV9DvmBLw/lMUIHaCby5HQHH5C
sZJ2xdB1IxTUgyfX4EzF19O+Z6LCyB3C4KfgNkSdhiWTozC6pikTerKeTbHacLX0KkziZF6pXCdR
xQ9U6z+107+F0i0X6sKOXZIbyW/DULY8FWY+jmVuImIjESc86oAPP1byOd5sil8l2n/2zbG2TGEn
G+k5flFnvrjnuLayMJkpGmjDWW9+aDJFYz3M93o9qf4g/TrkOM3ckocYMIVvk15oLWmxkL/33NqU
BIfVUZk7RqU/WgpVvlv2RHmuwOVgpJf3x4l+X6hPCKc0iNzfjeolY6DpupvOoh1HkO1R/h2RX1sW
hg+s+QvW30TlH1BMrUm3y0T93TAsMxn96fwVMBugyM/0J8n0zvi/bdrP+PH3WxzZ63q9At60H6PA
r14hpJNFRZB2G3rPxQaQtTLLSoTp4pPord1oOhb9sxK+9Oc2cz2EY6kS5S9VprAz7jbBEn9HNvIF
MiXZjnjKaHg6DbSuaVdlKEtlHHpeNtfJF6KMrv15cnyMumI1Cqk+Sv/eK8AtCz93v49lJXMkYkJw
3QqYXImJsd6zX/1vjDNCcoteG0V8Xc3WmeojFNyjmWU79ET6EQdq/lNRTmVYqMky59tONOPKtrcs
aOd6NF9vU28HU46nkO3PrFzCPCbLwVoEXFKuF2MImb11QfrWSIkxHe7Sp6PCMLMlMA5XgzmkAaSN
QGNfcjoV5A0wU+GmtUifXAgO33KcLKs6A+vh2sMJpjMECcD79jaKzNQZAvSHTNQ5WTH/5LWq9DQI
RWZU1DwxqaNg5xTcCnrMJ7aTAU75ZGnT2bvueKsKK5hYFs0FtKX8E1MWHCPMiWkl8wAhGn1R3zfj
XoNwKMSN/FDhM83rLLPF/MblaOBYFeLrIeufb+/18/+QWYiGY/OOVKtdOLPX9Vt/by+426Gt1lwh
GvCTEQv7Bx49+5Ok7SRq5oKmqwhetmCZPZXDdQOVwt4QJr75H0o/8Y2osN8ZEnDKq/epNx5QZJkd
MBgdRHqmMCCO1DQHKwzajUM7NAo/zyw6fz9XGJ/86St8KmOTmfgpRKdTN1e6J9FBs2Ifq5QEaZi5
tz7ebKyFQ8UySZguXszrldZwhoJjPZutXd4lEewW38w/BYEpyvkAGvBAGtuAeiXLMbCGy9wedBrF
nx/Xa7ibXu5leFimvTJtFV8bZHKULsCoOSgTQOQMc1xc8i2DK3SvPiNSnutbnCZ4Z9xQi87n2OZH
HzvxiYQxB6WIh4itmt1sdxzy3wigjsNoJWch5jIlp0y8H0YRFUl+lJHvIys0yahSk8yIOdxBg1Ih
IYMvaCxJ8qBLFg+0JZFNS/6ZbWNQjPWm6E+tYN6zkV7Yizvpyy/XrNR7XiyJV5uQTdVw8rPv1RPz
HTMEJj+0aMThPEpZQIWvdPRVNNRBfB1q4nucJw==
`protect end_protected
