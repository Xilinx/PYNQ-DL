`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner="Xilinx"
`protect key_method="rsa"
`protect key_keyname="xilinxt_2017_05"
`protect key_block
EZkTjCqolmWiKCZwXpUwsylV01ZDbBLzMdTBGMEJLsWh07XphHJ91Gp0PysOcBqtZBPaUoaGenqi
9b6kUkGJ6e5GLsUEMH9n/ZtiE2cOvsngvzIuZbUqTEG9hzqET8aicR/48eYNL+8tembP2M69nhw7
4VZ5tGdz8nzwptnYfY/VGgCk4onZWB28CYzY68W4lV2arEmvhZz1RF5BRasJKepPfIHKPY6H4sEB
rgXlPSjZse29dgNREANEJzcYwFIJaxoJQHkIO6rFYfARiRgETRi25kdW8AkZJq3J3FNI05oiVfOV
gK6N9aRGBlkNpkGUMFiKJJLJt+P+57wL35IF+A==

`protect control xilinx_enable_probing="false"
`protect control xilinx_enable_bitstream="true"
`protect control xilinx_enable_netlist_export="false"
`protect control xilinx_enable_modification="false"
`protect control xilinx_configuration_visible="false"
`protect rights_digest_method="sha256"
`protect end_toolblock="UWZlu0ZsTZMc2EApb+oCzFElq2ZkNWcIrDEPFDASFeQ="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16384)
`protect data_block
mgC9zkgAtainguRWGRHKAQSKyoM3BZzPoNkz1VqlCxXXG3S7pXnaudp/v/JLruZLNKqbA3cniU5C
gjwpeqSFsfWWrjF8GNJRsFRDzx8mpowZTB1hZSGXmbXr6fqEt/izfhB1q4YZb0brANPYat7MuwQY
TLVkQvnh4C23Jos4hygq3XmigkaaMmo2KSmtG8VqJgZT7t9Wkb+kqpWvMMP/Z1svBG5MMqc7nZBQ
3iQ34HoP3F3R2czvJNA6eyWIUmKXhoIxfa6xXRTtrV3P2aoVconXIN6ZfB6PQ9HFaio6E1x7vnko
aAthdhUyNIyHeiG9TGNXCfYo+P0K+m82kujGo6lfFIZ62OER+OKNyvVzREVUH4eHjRjnujoVuZCP
lP+Wd9UVlPMO68fcfXuQ47IUlroLAQ3UQIJgsr3IosdXAuKpRCc7HuQ2cFzIUKBwZ5bEZ6PmM/Sz
ePZIIcH3B9u1WOWsOirHv8S/0fhI9TsqRHNhsaGB3YYCIJbHSBGVwnJ+mjG68sTIOhyEqpXKckve
vophZuFnMNupXwnZ2c+BAAT1zyE0FoTUM+AWKMmqbwyaXR5+4je2QkRAoQ3m8wOGy/5RjVLQURj9
abuWSIXJS9uQvfXyKLpt0BLGB2p3XfjAM9QIyTih3RrdYCbRe5aDQZZzW0JwcubX4CEuOM2aWUBm
zdW2TMFXLlzYbUFEPInPhxuAuYlk6p03CZbkaUD4Eoxufx1pyvxDlLUygBQflE9jCQTOhYmwfHLm
qEhWM8O7LukUpyFyGFMgRbSpATfbIG0N6i2Kx8PlBIdEtlbEHK43ddZLHCvooL8xtC2UmR4itOky
M00AtAx1c8lJoz/VlLjhZoPGjG5y9cgvXp7AkzybyIgyCBwQtfQjoKRzheibojk6Gul+XvIXtx6D
sPeowVxz1fz2zKsjv5gBlSvJtTnu+eXPXX5skmDOpL4OcocvFebnG4SZV625IluA2WQsOH8Uye6Y
y9ZlIOhSemxWVGhDnPlzVgIlysOD+5Etq/Z8ENBRnAVi6WjsiblSJbarixDtko5PjQDckT2VCIqj
jQy9DyxILqilCXRJimVI42yIBqkWnoL1yqcRwxNVvmlvYsNzwmWv0CobtAJhBu2a9rBC2BT7we/e
1xR7laTKr6mfZA3Mn4XiNVZTXUFuKemUW8f9eKKTbxyDMIZPXiD0yhDRg4xG6S7ESDhkxyYxdy6K
UQWImNreww3Ayvwydz5rbDBSo49RwbBs+NN+jZayzMlipriCOo52s5N08ZaOPUG+Eo4WLi42plXE
dYf+d7wy+EKubqTEGi4vRcsCPt01WYZV/dzVQI5KvR/f1osGc2X/kU7HTHYU3WTwWGb6IQ/nFTOA
vDAMe2BBdgQGwGI/nHQMN9k5f6SVjc3IRl2L0m7++1dMglY/km75PbAEbzzB+mrPy1/nD7fiY6AJ
aFGrw9adPtQzYrKJO/rhHAC9xcMjkN/Q1/q7qmpfgYZxqIq879gJP6VLq2nUB+Ag5eVXXpiveio/
axE753mTr0XLOrSpWr3yDTbaHlvZnPiPJc0hByW3b40TPh5ALrT2wBzIVF++0whjjDv2BTdLLmCS
HHJ8ZOeehSWui2pRRBAbXDfnWinGn8/TL5KSOruvxn/VkMQUDNeLVtBqQ7IUenmiPyQUfWBiaAWf
LfY02hrlNvTpZ6GenYBN6duVHuCb/DilJ27U6N7wgWtNfYjXMjqDD0amoClKCTfUydGiWIO5nwQZ
dJFaEU6cYMJgYHz9loJu7D+Hvpa+6wXNYpFQGIL1eW+fp9o9i8SkgdDAYcjl3oCMBHQAxTsMNpEh
mKL1thd3uteN3D4K1wcm9FM126FxrF03g70ZiW25CivQIKnK37Bb6MtJ3M/GC/WKWkNy8Zn90Sq9
qXcxbJZa4OMQ8noU7c6gdmDBIYnJExBqMdUitRhVcU3u0O17Ubty1dncIoL68PHugl1+R7Yyn3Im
LWBiYSVsYn/5CPEodquvo71XWExlSKSSCww+6gwxrE5qWWKOfS5Y+SSTjpKJbiRlcFhrWbqOA53S
8ylyZ23u78EDAX4K4JnO8bupWfgnCw7PAJ9u8ihHrFq7gfKVRzrf8uoPjGuKkkMPJA1ptt7jSKGM
K48ZQKUalRXw9PV/aM+f8oVWvl2WzrrDttAdk+eMDROlYOjbE0bljxIKGNwHGpL4EXSnP6zmVIrc
0JB73pDC3sQv5AGjp+H5JFgyEb8PxJ+6OVdMz+kvwqUhAvRuaOByJwSIOajCOWCuU996QMC37QeZ
601Tz/9nKQrOSyRbqYOlNbWGLZB27daLLg1cDqsMJQHy6K03rQbkRH4SGkxzBFwJTtk3EbA1dWBs
yhLd3YafYYA+gFC9M5rix/CzFuLQVJrR6qDAYx8DRBHi3OmB+9ijhS5c/iAjGDbXXVrSjPb2SDbe
pHqyox/w1lcnmmY0lasJAUxEGrj6r+F7mghJxu0LGRxY1bYNDLv7ixT7JH/+iTaJZ2bnv53yJB3U
ZAOsz5U+tJgrCOC3D+Q1pGU6OYj5K12fOKrZIt/tN2ey12R5xtxCo1qShpISTwP99JO6xBba7+cD
SJupfL0dhciiv7F+Tika9tJAbjC07J98521SikECAqkpdOUlc3kPjN7gz4KOH7KxEAp2+9QlFHLr
CFOY5Mi6tZZsROcwyeYud6ORuIAI+Z1ZRLtIYke0Q3LSwbZuTA5O9NRea/vodRGcuXpzIqPoxiK8
0m3DyxN2W5q1BGXbk89Qt2eEtkcGXpYiCru0+JT5nGWk/N0xWCr8TcUDD79aG5MMptkghvfqrBsP
CZsvhJEXHCVLdCwUpoONf8y/yeg8tpNHxc8VkhVC9WU7syJE6PC70nazhNGBU7+bCAQsCEye4wr3
M9B9E0xER9wpjNJwYuHxp4vtkot16fYvhjogGmdOsknD3hF8gwJ9tKGwyx53K034Y8g0f+hAc4vO
eeXK/r8Xhk92A/ktRINB7qvvmfmB/y2dzHBlZuZ4BIBdk6M+D0mHcMdSx2+jwv8fdBXg9aUo09Uo
4uJNF1jmmexX2hrduoUTYnQXkYU273PcudSekeIRwKTDIHVpP96CIrH5cHzjGw14gv4ZN/z5Nysf
pZ4dtyYIh0lCjsXPWYCKBvaa3RSi10SofKtBQto4x7KihmrFJmQh+gFdBAPOW3EcUQyNAnHQK/Sy
H8hVWi8oN3EKzwtRmZl3iGz1FuGrn59dH9BuXwwENko+mP0s5ieseunLkLX4QOsxbfsEyIdLzdm9
sEtWDsOE69Sh/AsLQbMEKVtVekHNlTxz3GS5w58DyRK7lf46kRxSk4oOvT6CMUBjwWaeq7P4nTym
pEbqe/MjqdMXZiUmRHW+AdCxXkoDiprgnNxyeKqbbMlnGx7uyfNc72ga5aTLbITDzocLbiqzk3aX
iuuIT8z9dgegvbtmKUZgFgilScNO/qrQKh8wuuQOVY3twrFm9ElJDJTHB8fDgbyHwDSspoQxDb+Q
a+B5GcdmfMJIf0puo0nAyy8sdlhRSbX/ktxVRIrqlNeAKtaU+QHwcxzSRwyAGK6UUcuW1YXFTnjN
GQezMSy14f98T6gwZJ5cUcSE1IZGDmUzXmZZvBSbMvAc4daO6duM2mtyye8VbmarIR0pTzNXhcuO
wevYwj73xkB5wHD5V+qK1Qo5JsR9HYWQ3yCjLyTreiyVYAJeZV1cx+3+o+vO8hsud2DK+XKXGFnt
6duh1FPJXAh+fKUC/vGlcAxzR8M+dxmxJ3qyzg+4wBXGb0S9/JDlZ5nmXOkx8CsdbQyiYYBTytYC
6L/TGBDdra1o6MkG1ht6OaYhGladRWz2qQW28nMdeY4/gNHRNNKyLV5XGjo7D2Y3PgE4SDYkfEgN
L6rUzQemE/WVNGSQL9V1IAx5nHf1cmjnCF4gCfoXbve97DuLDFn/NkItdFkkHGgrUiqKZcyQAvvd
PjRF79WLdv6Hcpb8dt+2TCuXWn+M+ljZIU8C6D9Oll7X+8hsOfMiRdMiv0hWWhlsGowbugY2LAak
QhWneawd9sPy2DO+7zSEWoXIeWKn61E8o35iyCcTctoVrFaJp+RFe06WDwIM3ciPZ4mvInoeuKiJ
hVq/Pv/sCFoqFoselZMJPe+84KngU1RidsUUD3TwBq5ymeuVh1tfTBxbTBtm3lqy05RJgyeJeSD6
bL4cf45fofbAuvHUi1hywogplQx2D0ThcPasRPubpMn9axSrRUiYKVjrkWywyePu0eB6EuxNJCj+
x9xj1BzbmwF1sM0m4SEPnFvDzKD41kaL+lcYaDpokNdn2plfJKpovVtYWKvD8/9yYtP+XmyrJvyr
ho3CVp6DJvcDwU/BavA7HXlcS865zk8qwUbkGtG+zhqkJxCm+0PGd34bEyK8dlYlMpZ0gU9wVKSq
PSofGy5cnKTUZMPwBS1gh8TCMX2jTvoxMwJfCLaxZCp0g97PmcTPS35j7kbx7tlgAkDh4WOSykvm
6up43+DRJwwwTo+QSaqZOHY9Q9qMbRuFaO9NGuBFN+fi+YkWoC1c3fV38F9rnj0S0NgBxygIHIWQ
5inEU/3nS9Zn+C3mWqVMLcKdxzmZuvxiu5oft2ngb4cplOQw07KJoyj3qFeqF2mgWSbjP4yHoBGy
lzjnG1kh1OwsOQtYq+XXfp3Y4AoF6Ua4VuHh0wiTro6AsHGhVevlRXaVhi36FrLi9N8hJnLl8S8q
XeQwtYFmdi265X95FjAmAHleUZFh02FH1pW7h7wZvhHWByN3zd0fYoExLszY07+3OCulZngvQdyt
NRk8Mc623aVGos7V+WYhcPBN8O4vA0YexvHstLVTDIHScUI108RoAp0u8aX2n56LA1wEcl9ZysIU
0ZSsmMtmURhpOQcybn9dhxgwZb/BG+o1aPJvWoQKeW3EjKZoEL2mo2LGUSb1gbLsgSKDiruQER/C
Cciz5w0FjF/btzPj21CMCgPfn3E2G5aQUDHX7X+1AW9Y9jcDdXPj774APbZ2RcFRJ7hTX0HFN6yf
l18GomaIeo8ESOjOv4GkVNJ93fJrDl1bkF7LAnIPQB+n1P9X3sz7JNGKuAf4YmQtwV1IfqdMk6hT
w/bn6KP76zypBpiD429UzjAct+wCHj4CUQe1oSSIanA681e+r6v6q+9QxK0RG6B7OHIWWEYG9fW4
N2UTAn77ikZgdfevTYFjVV+eFOCOd5apfEX6VY1J5RmsxcEwgANwTI9tFFkMC1KjpRWXGWEQAkil
peol3aY6Tf8e7Xj2JhrnrZiU4r/FmHm/oD+le/+mZQOCCoPGavCFMLdi2AF395Tpqdhl/atZuvNp
noNhayabvzz+XOq5BG/V+CY6NDMZ9bOxB9ARq/LShcIUc9pI8twH1MeHYizFcol5ePDuyjJYrmqX
atT3qNvdS+yuDGV+Ruc7aqQIHpL4hulLGL+WSw+kYb3l+W80MGTTDusgorTCmy/nAanBWKqBd39y
D0StKGOD1acbh+51vtyKRfft0Ej043A/9c+xHd3EP96iciY6alpwXTF7/bEjxmNK4aKMh2rJLiRm
569cJT/DBYcnUtgMhzVAvRODWEZpZefffy8UJSGKrhJl0Y9UA2/eGpbQ4d2BkmeNU5CfV64+7YNO
c4RHhgnOjpr03Amm/PLvruZMlqocJecqEWGChWF7MiTNgFY62mZ+LmewFO4JrpWvNjBYqgZy+vGA
Xu50oGvRbo0slhqAByah/a37VwR1ZI/xf6KLX5/AOMZ4cb25ngMLDCOMdVaH/deaVqHmW5XC3PQY
o9LNUHeI3llmCCEjzX+bQEmGY6r8uz6KX27T7a2Whx2do1Bt7KI8OMJIqcz6EKPP+kBYM4DedDsS
VcguzsAemNt/4ggnHiLiQc9fyk8Snx48MTiU7oQIpr+IN8UKsLu1jkEDaiiXoHqcK+3aa1xmPDLC
dZW7TxW8+9fdmOLRdZFwyBqn4txtvOH7zLzHSKP14H9Jju61sCdFZdonY1hhJx+FwiXaBYEn/UYS
JWZmHUt8CCNGvNjwCBPCUWhUn2ZuyTsLKNI/thP8M5Rqb/qzBLsv8UWdEe4/Daa/CpZddBXpc7GQ
9LDLc1rC1JPc9iPdEt7ULsWZv6uays30VGxLNhrkDAoTJNUiwdSdLBJPSReJMpStf9Y4O8vs38B3
ypyfSfPTBuU1wKLBz0S8nW5zL399xXdBBU3TZoHn7vqpC9bU3vqrsghu26IY9u/FLXYNYkexrG6z
3GWCAhEJbJMY4bg1odxpBr8KNYFHJvJ/IAV8WqOEZMGTxY9FC9x7CWkVtszwXVVNtiPdSwMJONOz
WOufZkbPmvVVjIkVpQfZGn3lhHMTeRaynfjaVEX+bbWeP/ZqM8F+DUwYCcyfpvP/l2hdjXoeSuyX
B4gK2bo+KS365emirRkrEQAJI/AhxAkTW4iorX1S7xRDWXzk7VeMUlB9112ww7wq4Pjk7UpKopp9
ySuOKOJQCSlSYfEF5mnjcIm/j6BeOaFfw+qDAKk0KJB50/SQrLY0kGZjo5VcaJGzcZOM8ciOhKzt
dpw6R7Jrz/ko3srLhXgo7+3G2gPywoHm3PP7maomKPp/kGWsX+gIbQ2rCFY5Dhxime19MM+Jb1CV
J8EYXBZ3UkwIsr57/cswThk1l2YPXug5fliR6MzHhloIQCtDsx1ItuortWCuP045czboT25riZy4
zkrtLybVGdcOuYvXcDOHTb1gdOlr3nC1PkWvzRzPSFaw54uUswfxouhFaoxda25366a8lnyu4jV2
ARm+69M+TwykPQswyfLNyAgbKkpy6rLrQjxWgg+MGrErpy5R8ySDrnB7WvrIS33bi79AEAm3EbGm
xjcRidI1oFjfU6+qTMn1gr5nQrmIN5S5puLe1hVfq5Ko44JS97cPhEc3hI/CRWUGz7gQRMrkIa5W
T3ANivF67XS/el835DIr7DdDEQRedmWfr0gHdhNh53cC2BeOB2K6Xl/w8sCxgEj0oSmc1U3lsGCI
Z7jM/V91wasVcGkqJMvezkT/ArKO6ybCkO0EML2N2PzofeS960d7c4lhcf7Xnh6aH5wzLrMSyLhw
fcXqJDcgRfxucw9g6u3D+tu2rc4rpNOPATSU0bg9NuLha/nu8np0hFLhl3k4Yv58AQTO1o0N7hkV
qvoPVNkAq0agIYiijTnItSi9X32TwMnKEH/BvzT28c+8Uu/G25jMI6dU1xAmvOC+pPVtqmf2cs3y
q782QoR3CYhEwGpbQ4fJzVifykC8+5gHJSLBtrOGZ5ATu1AOa10hpaCCzV+FvPSYGBiltW8FI7Zt
QbfkM88mRP4DAm9ZRqS6AqxpT7obTznwazvb9KGSrj+3qLZy7j86BJtWKdcdnUh8KOR8yD4Huqci
GvHaQxLs85gmyrg5CFoghhwtWic4vsbU5ymCKrc1fbN319A/JsSXk/frKsrgV9DTUVhJ5pMhmTsH
Hn/FSdEZGbGTvoSIGDTKiFzOsmmDXLxPf5xp0bXblgbUc7JLnTKp60IFMG3U6K2OhefCQcAmDc7Y
ndgakrhJnMKQuuk2hyFY0QwvOel8eOSbH4eJv+5WmZhCyxRfgGpKosiv1f343/T4eL86GQmrLg6D
z6yW2A5FyW0YVC14VOvyiZF8K+tqOUXWJvrl3ueRBhgql2qsk9brLCbL1xk9UCWbKq4sk/KbDxaQ
Y99Lop2fItzaAbLn8i1W7LBtcuPBS1jRFz4U6oMfom2GSXWcSprLYcCME/htjrYr1DBUF5orr/UO
04tly9pV8YylLW7VCdlh+wPwSzcHE1Z5oYiRwKjiRGJXihMp4PAckHc3yj4CBOljWuNYLiXpjXqt
m+FXLrTA9X9MpQuEk3o365ugSKio/F6jSjqKx5bWdlaXIGyLjGG25DR2kDLjAqBMtiABAjsD3Bxj
kzgROXMXkI7NPx6F5q5/pB2Q0I4WOPxYIJIWo6XmCBjINfBg807uAPRqfw7ENJH/eBrzZryIEeTs
ZG7z1rUJATG3Xs6dkC96eKwe95Q+3TKOck50sx5XtA4JArIwd5IIT6V8ehKsI4riG/6rB15V1EdA
03wUyhqWkhxlX+d3k2JPmsa1EX6roSVZ9ZfhetEu91LCTHqN+fUCi6piP9gCyxNepY2wZ8V3E6kz
AEwpH4VgSKnJ28hSGHArgPG029zb34Oe7pDz2WXiiozhxzivDDytmpRT/CsxLapgb0+v2/kn6MlQ
8f1A/E0An80Ozczntqwr6fk55BY+Azz8Glg6ZAFebjyuKsK+RG8fWh1OAxyFFNYjdtF+HYSy1g+H
9tc58D1JUTiRVDyNxhUc4RIYTK+t79Vi95DSKdxw+1klxMWd4tXvj+O9JnSZ/7TJN4odH1LxLjq6
80nikS0k0snk2jKg7h80upyAO0Di8CRbwEaFGcMMEGc3O4C+ys2L37KYRKhPUqVu5hGeGrX/Tn99
gk4ldA7Vq002151XEWb0VsQZcyr8MFBEESog/GhkhbYn9DRbOXcEMhS8EgvY6Ibdh7r2k3wCMBXB
SJav8qTZVTlVkZHqRVDaLztrI7fw5sDJoS/SXurAGvZxZhtzIOMMkuKDAyuH4bJFkGi1nxFZX28m
rSDWh0CyNZ0ymIcJk87pwO7U8bEZuBJiSjcW/b0GMM8ddSERUIHOTr4gSTh9dRbsAAFGbp8I/T/L
YoUQeohGniCotp/UMxLFU4crhU8F8Zz7UYfKzzERW4IH24r0CIouR0yif+b6M+iRdfOuWLsJw7Wd
ZfA0mnvep8eat72lEyqaw+u989ZbzEwsBKIT8dGgphCMsHCg9g+UfDWz+Mp2RX1EgRvt+ZheiYkC
e8ZGwApFdwzPDx0Sx1bGlShoOlS8TA/YRsSUWSfV3EtuWjPTLpQdEX3nh41mCq4MOIjt70MqMcZh
8J3xk3gCNhhMx8mEyHvBuG5bLX/WJ8LST9qVOdzZYKMhjLXt3n2qa3TP1+QRQJgzRoz1FJ0qA31R
lW8my6+cADbjWEtSqa8ikal1QMol5qQzKZA9cPwJDPhg3hBuC9iB9pKLXBkqdMgE4fTn1gX7XFdT
mZSgVs2kvdvOOnF3ZG/jcSHJVVEcFh2ZpHtaAWwODQQY/FhyUe/IgHziZZ1BH+jzSz56ndOqFsqP
MeNPPDjWxp/nF7TdOfm5nXC2OLVkxX1YfgWqIDRdU1cDqpA0IIsX5KStrDFYChF6k/p6rVk6GX9H
Q3xWnfnD4kkxCA9tZ2Vtcgoyz/BMr6qKKrAcTUWxgId7VLL38m8Z58vTg4JlwxEPaB/Fyf2D5IzO
oBcbHb6JXcO8dUsvQC7z7unW9DfjFECbGG5/kVfh6BRIcDjBVa0wYYAsM5B5fuAz5V44HeWrumIj
rvNJLz+q+v4nqpjAeOoLl1909sdJzIPyTx8ToHHje+MuAvcAmdkB7h9K+LultT9CP1HMrcML27Zb
B8ZEWi8jLLefeHCsFahE716oyUNc/9vNIZ3KHSMG7TvMi2ATIfpL+JsB5CIaTAle4C975iilbm/d
66f2n2mQxURg2XuLyiEsEE5MNzx37xbffyxoX+UKmfOXwu2BABvD0oEW9M5V0uHWRlCtqhRQuk4D
yz1LZfdpYdq5UWf74mRQ0tiRlFHH+EifeZN90p/HgQtbmYdSTJ7dCMebdrbdN4SfNB3LAsl9b7n5
4oaNExVbPt+RsteWs1tYPF3MNOxabrXAQpSsBJ7KsSJ1JKH48hAAeKncqj7V+ssYa5sb0x3NjcQR
UoPWkTwWRuy6eTyLs+07Pl55sr0qQupFOYmziH0lttwUG1FXLYo/eYg1gMDk2z4UlG1m5J9WPf2F
OoBuOzzUbuVeRFoQLXSyMGTx34eoPjya2eZ5iUVLVabCdywwaIwl2ZLwGnAJbcux6LqfrE7bDTOR
6RbiLUcuFmnOVASvjlPoYbivahf34fnuMhw6pVb6aP0RhcXYN46r42H5W5hvHOuuuG8G3Me04swO
DiDx5+pHxABshXcZd1jRVVW7leeDmBVoSI5qM/EQb+/ZXj9m3r726by/YumBdIU/ojqKS6LPodsR
amJWmbkh4VGEa34I8B8Q2AJoqrEntBvm95yJHg6o5sQSxa5rCp9FiYz0rYebdKz2/syB2WnQY1Rb
8bMbap2iKGnivmNk6B/MFAGxbpuRRT3NfUnP8MIadZSISV0pf8PNibUHa902v/MPd6oxlyU02UOv
iUDAM8yFjXrTHr90aL8ryk0mTjJpNaLe6dGT1Nh+ho65aFp+VkQud4WBuvLOcC+uh2F4zAUfsHKn
bwHRLRw19PTPjtOl8uewm3CcH/rYw4Q9y7A6zx8lExE4ScHwRfRQDjj7JZD75bIpDLPOYGJGPK6r
vUCYYK5xIj8BJ1rzNdr6uatDC0xwhGPSe1IdoTfb3EH9gxDs2o+l/lVmOJFTn2+xSw2H7iHNNY79
iJmb7vNb+jV/0raSRQ1rD9wIAeX4fjg1us3Urzo4eMzLkFqHtE+jSW5wAkfkYCd2RGjYwcr1KT79
og5UmARrH/uvLj2iBf4v9lUFxR7YiR58On0ugoNFb39eD/HTPiVnZi9DkBQin+fYeOJp9kWoZbVy
73ulorK8O3ErxqwFql+um0c77E837GAiPw7/S/bCJNJ9yzoGWYm7cTa0Njs/TGkUs4ZF5HK2AQ09
D9S5rKY22N/qFW6qwEmVJ4OwhsuLS0WAwoZ93CP/Gxy1S19gSSSPdZ5apDqzrMYxxuKNjYAGASpi
hGgehFm8svXjfsAkT0WZ2gcn1m67r2LuFLNVMorzfBzqu9UjbSGUF/aJecXjsXFINycick3EuL8O
NvGnTkRVgeINLbMdbYJq/FjykRVsPFeIMdlcNpXa1iysc4q/bkiPG183B5YMEazM9sjEsePpmtcN
XvOQGkcVpB6WU5fZN727QcZcuRhKxJQfK48UdW+BcXQ2jGEkB4x9c9Jg6mPq3b/mqEvdndyJFZ4a
6vW3erc8XL3L2zFjvVyYzi0FuvdKaBTU9qaRnhdM4ntAJzX1vYVxdqILO5ibOrxpI7UfA6FDjPr8
i7ewdd1JPvli7xSxpJh9EpC0SkDz6c/E/uhV7QwLT4IxJfkQteiHb3bkIXu/kYy9gVSuVjwvrjaD
CAK0PUdYdkQb7s6dCaKCa0t9LnDJNHAbt5BkeU14snB9DVJ93TBal87C3welxszPjGDXM2z95ah7
dvEmKz0aQS/bo4oPsdIX2Pf+T3KsMfyfl7bCNq3BMfh3yx1NdvvwPzBDa1jSxvRZFc0N0EWFij+L
DAvjlBiaGVG3LIP08SMGuGEcsCRL+mOBpOQsqSmCuuvyEGLjqat8dXnzwoz111nKfMRhDy4Wg83r
eJhUd3PHLREn9FGXG0o3tAr9r5YFWLNQ6exB91xkuhPnMKYwo6hVLt90ZcBE8W+DN+1KTNL+ibso
xVwpAPC46JmZojV5mmbnSaiMwxaykoqEHUcvN/9IyNedB9ozKEyqSiSwXv9wmTVpku52RqJuSIlc
DWdG+h9O1cmeXPDbPeqLTCwnX9wZ6oLtOmerSdiPTChPJPdhhRg2TFuGCx6EMiny/KcnAvvuHzwx
Vxl1Gh/8bmbzRAd58tzIRKs5WylqJg0suJa7o9r+nXRyEhb5X1tn0clzkXtNYa1DcPnB5btFwKAE
LjBxCekcxAEdVv/yx9Pa/vt6TPZXpv1ea5Dhtd+SwFbxfZli1sAxLbCThPtMTTIYiK6elx/0vbBl
6yXpHMjfzk7dDTLkhnbdCVOsQgyofdSpdT1hJZkBkLyHI0KzdclR5pVqcPoaXJ8LEz9Gv4Z2XVxl
V6nFIcJaFO/OKLtZFkfgULUL1TXJ+se7yQRezGdp4jWc+Ve/Acj0cBrvwfPv0kxDTP9ZQQmZO4Kq
XUJNWN1EzsXNtVvdFcpTios0RGsUZSP8xZXppJMbF2JAX8mApTy7ZGtPbN6oHjVFl2HU6dMF99BC
B82GJCtMq4BlfEfybgcCKBVErwlrn5BrLdwasli3ZYUUkiWSt7paOylOvqLh9vWHKPI7+Yhxf8T5
a2N3oFbXjaxdBhBwruEgB7OGfAWO/XJ0qNPC5pd4eSfYjzOFFxQLSQvawjKl4F/O8vWpzS+GH6jX
hd85ICMsFIwWRPMBu/XCRRheDd+P7KeYLFzf7FVXzHVKA52l+vs95f3dgRXla6qyLze8pIkgGO7X
QdDwOr5R5Sfc36xH+YmtqU4eMO3icjYEw0dNvea1oMrW7plY+p25aLkcSUqSFciZEgxbM4FI1kOJ
OPuHrHTcToUjVK6cBNz5SmM3F97D2t8vy6Mj+DT6Ln8o3Ox9duSoj2vVaJemla6PViKPWxGwEoDz
Lbak48vFmt/PWPX9EcPzBR4Ie301Wb+vxDV2VouW0dqdHtTBHE0OxaM4tJtusfTGnuHDUnVt2oxs
NGDBECWAEcJ5U8R8xqBtAmMGMyvN/vICBkyNp+RGtoH99/GYoXfPA2ZNX4w+14zLM/jLj9dBYIZn
ceeMro5F00+G2Y2liwmM0QjHZqI++6T3OPb9a1JVVBz2dtEppX7qMK0bkRFDfRRaB9YmMbrZ9uM3
YUCAFKYDAiOZ1NtebV+YGGJq9i6q7jWzGsuEw2/z1IifZz4mLhsonakuWi7IA1+KhEyPNXwhrsuT
lTsnAoNVE6FXfyxvVlKPB8ZvCJxeu5o1sYYmghgOPAJYmvmu+hl+VN8a9ZlSd3HNX8HWiQy9Hb9m
jVTgI5a9p8sYp1AZpYnHsJ3ADztuoKLGW8igLcqyZtE/gapAAOOjVZsapp9tEXxC2hb5wfjr5bZ2
GwI4KE8fyG2pd7OfyLkK0TovkHJ7jQB7ZkVjQU1de9adoin4/a/ABhUoSHGmF2ciO9FVCRdnzuPj
GKXACHKoxsy11/YBdG99nxK5YciG9LHlw4KF/f5MZEjbJswYDoNWwpG1uDGdIKWb0Z37L1h8FIWA
5QapRm47dPWrzHJm5N2bKiJLBAvXs6yplxEaJKFmFE/fn2J3b/dr60UYbkN1cWk5RfjgyagMb0Y3
sLoJ5GzRylAlGi6YA1CS8d+cWm/V9IGGAsbkxyp37PR5RYYbn6IUN9S1h4o2jvaUfORdftiKPgii
Er8yckGiTOX6VyDO2YquNJ8inr4kck1m/gazz3UYTSGnNnbc2aGkiczHvkMjx5MjMKyOfGxFzLcJ
uXtAA0saCtGwJ28y3Qzt4Ksy4qnMziCjUbPZQy2E+W+hduwuxagyEsW/J8PqadSECEL9OZ2J7Sbh
D2qSPP868vhELDRyh0jeYvFgXJ5kSnhOhOv4kIc5W0U7Qx9LII/e3OMRufW/SYw4bVpD9hxzztIT
62Idux3fUdz1yyPlGRuzRPu5uQUtYt0Z7Pb3ryxW8fXQcVHlmp+DTTt4JXQTfI/eHZEmLXuy9Nix
7vtFayjhLyqShHDXNZ5biulUekePbH/IUkSo9NicLxS/W7iYKWxCOb4JKCJL9duAiGBmzEl6G1eb
Xf3G1g2lUMFlvBgj0axixcNthAw8/ppIFhM97h8NB+6sddtZrlnt2hBp255yrVek6wgLk+tcNHJ1
DYia3mGkxKACJI6cr6y1hxKSrYXVvdSE07PUpei5HMeqklH9BGG9GssGiqqkxp72JecauHFgGtTW
yekIIjfoWnotPN5KdH2ArhqwJJl2pS7UXRZzkYjv4tc7E+aFY9dTBuUXcDmdxAx1AEFqC6F6KlJ2
D+9kk7aRPGZ1+xmhsQQbBiQ3dESJTj8Xo+qatUQvpNWIja6EKWrGkKbbRkg0sQfOCkPq9QRc92er
uPh6XPgP9JHkk3J21LOJKTowpac+E6XpXDizHIpTa3UaNStan7S6kAm5DTNRqvPHnDt0U95dANXc
2a1zknNVjjRg/Pv/JDSP2RYUtI162CCLQn4sovQ3AcYaR+LsfkK7uYw8LbJJl6xRa3ZtjUcOZRWT
sS34PdwYFuyMbtMTUtSIDjooBAb6IjDKS5oRCg127i4jEySXxvxzkiP+KkgBtkJIbd7e7zwnD81j
IqCxChPzU9FyQ8oaPfkybaH1GUW4IB75WXtf31iUrWyTZKs8PierFdumOxDU07nB8uY05JI3fRka
22BiVn71VmqcP+jNfytXQeA4KtvQ6Wix//BErPo4Y8aCBhiYEkK1iOp9Kl7d1Ubsd8u4y0zyyoga
oVKJyv8qRq9uz45wNf5Q2DgeQ6uq/q0t9PsWoqr/yQVj5uh1TJqfq4pqQpg+JeG0avKz00LWorTr
Ir6IErJE6qhJkizTzYpNHGqWlFvpug/XHzwr1tNlvWW4TjP+PDWN37uX/KJEfFcVXIIMgS1ls4RV
tAB034FUgJW4TQENK3DDH+996No84YYIYU0BOTDznderTntR6Gmo4Ljv8aeK9o1bacFIEoQnUyZm
Ud+gl+aNVVMn9Bzfj+cpSNfH9Grso5NY4I26J2+MY/BeSgdhLvyAtStjTYwmncNMIfmNeGHMZcX3
Z1ceMEMpjw4dTyHI1GNxJDQ/QEF2Oz3WU3wooVhkqzv+VYf9lfJZVCTMNb/AyDSl80tbkwrsl2YG
l52fhzUCKzfpfIwn0wRCyFJWml9/l33G5abm2AK5s5YMVl7O7YcaOsfUu/5jMJ8Nz1Ky+MhSt22+
e3IRFNaZzJ3KAt8JOZiIPpmyFba5VyCxDHPCrWRh0Arja+PiXSygGb3Ps1NZnoXqPZp+ueO9SZ2x
hbPKBjq3M/RoqD55FYIBjxKQ0AJj+iIvEYjnYcxKPscplXAMq8NBP/ROZ2MlO9gG0ctslbRAX1ID
KfRDq5xObvkCuxEZdHzEcOgI4dVRv8IETrIsVwvw7ltlggCYTPIdWxhn3NnVOu7Rv5f8ONDerVqk
LTNzHS1+3P9kHyC1wY6n4AF/XAcS6nP+1IGlCqmpR1FHYTJhY4mXesiRM5lkJeFSvL5SC235rLTv
guxevjN6Ive0XJMNfdGVMIeskNdp93uDAxyNpjeZmOBKuCat9Vjctt8FsJOTpy329UFMlVRqym6h
EnL6OOLeXMQbqyuKEv6Wuw3mR7sUWVJpYTkMAM3YSQV6N79ETNiDMvgTKQbBxBu0F44gYEi3h88J
dIXQ7NxElvcE4mYnaKkXY1PtLPHDtvqtGmBjwmGOu0oOLge4dsGV2Oikzdvtu7A5gl9TzkMhDkrl
sGxw00Y+DuT0XEnvAj9eVZvpGxv6YfaCxdlTlrZPfZ9kxhnapEJhFJgNSk49e76seHx+qE+6msZ8
4/tYurDqdUf1ANyRinVd1gSc/vwK6UVVn/W85qWOGpL0u0KtGR2lCvURHtfUtpuEVD52ZlC9aJ6K
UPJbqtIz2wk/6V+8U3h4sVjxD1cAz2Gt2IB0SwNzl23aKXMILjXJPHqUd6V1B76uhmUb3Upov5Fz
Dqc0tRUB5LryKfzK2cNsI6wf9/oy9Q7mj5j1MLfAv7kKsYtVs8CPjfpvJIA8V7ftqpRhJIr56r1b
XO8aQR2AGNQY+cs66s2wn5ZoPNBCKtUBzrpSf0Q3ZpuoFq6XBCWxrY6wiqv4AfS9W1aFF/O//eRf
H9RBFM0uDAFtMpazdopjxa8KKxt80LOEt+mnTFCWwVD2G9gBAA74y2Bfx8IRNmi64IOyILXnvb+4
t/VbuN4nZoCXN0/5Q3HNmEJG6BJOprQgrPy33c8sxHISnfaf21VvP1EgcOI5ml+tg5TWrqUN9Nm0
KNxb+z3v99EBkdQalIeWdU56+pxH5i59LwHb9iO2UXASBziSNGD8JzxZ2nC1EtJVgxxc4BuPD/Gt
X+aZEtc2HHojGqtYIVLLoNAOvKwXLV+RJvvkSi7zJGqcQPyG8OXMNJ8QCz7mp9g+1APNtnA9HaXK
5Ar3G8Ty+OyuEqEFt/x0gCK8+kk1gwspQBq3lA7tWQ9DfCfi7BMzbN+R4oYK2o78JoaAEtIex3jd
4qb6EMTg2dq0BKf8H9a6yRMqlZsWm3otrpZRgfRP7yNzb3lDHqj+gCaXL1AgJtEy0s+nbkyiuh7i
kMkgIJZorPPYs5+xcaGV5GIEPMHGm7sPtsHJAi9w7UyD2n7CdZfoEiGl9VfVRA15btz+liaDIZ98
pzfYlBUq7e1hVlt4j4Kofw4Vrg45cqpWH5rKLaminGq5OYem/EaDJMkXAbj0s5ZidHR7xWB+tLld
LoURPSYn/EKy4RTI039/kyufuClTj2EcUHdsSS0ThgOf+j6ltfh4jKXnVymKJRMRQRtHT0OSVi8w
iA+AZTgQ8a5o/8rOUX4RrFmNpELR+67R07uwJzAZBX+5SaGWkMEKDfZXSJkd9l8xN5WZNif1J//o
9fkBsjHUuftraAH1dohWY2cqTKAamoxS1FxrOc11koQ+2MJ5Nb9I6o2O0uGuOaMntrTGM99EWfcL
pqy5dzVZz3FUg07J8UCjthIdQH1s7iD+GSK/hGbqGrnKkCYiV719ix9qmfX1J9I3MWVx3O/2CzaD
ncD5AO/DvxokqyVjKQCMo1iwnmQnklXO01CF1CB7KWH8ypcFYjFAwhDGlsC1pYjKrBMQB9o1VTi4
922jF+fqUqqKidkcO00PQLJpCtd0DyT8FEb+0IX3CtJxPoeScHES0xuJols7JwcWgKvOqYuIhtts
syUxERS7m2dzpqzReBhL50eOlnEW4t4n3RhD9l60nOBPsfPfe2BhTHa3pZ0nqdhXYtfdr2iE8Pbh
3w3lB7qQCBxU0944ZRbT7ffaGw9VPJ9oFgu+i+1BN5+tZcInGdqMSLKFjVDdjNfcFzWpAqVcyhpj
VIMUQaYv5/wCImo0pGFF0Cqe4QXEwq7JpTsu2TKZ7skQIq+AjDgXXMliUisCjlmkvYCcOBqzh+mX
fsXevV8vMhDWM3RDWZds24WQrVAIK/gRo6WuUrypoD0Ngi3OqXY4YQm4ejrCjexTWlgbzZeXLjx4
u+OEfQss3hGvhLKEhrrrBDa7kcGN/BLu3TCYp+0skuX0JY/HAUN8r2/tMutTVuxFvLqb/2iWrwBX
seACvrKe3kWP4Sp2r9oGM/gXmppGC1QuxXa43tfMRN8+a+inSw6T50660nGtzoRWg7NF27dgOoA2
oFKPUPCE0YWSm0cY1rrhhwQT9kYGH1W88pb/inaWudFP1ZUm1B/OTZ4sZtRRmX+zRB13NHvX/s1Y
2mDyXuY6CALwVNJBGpJFHzae/KtMH/rV4Jg20SKD2Lp0aVCCYQGnsNJlC0VsTwk1Mp0uI9i/NEmH
LXA3shZfjRNTsDQlVYAx4JEwG441UxrwYZwhBhFgDbYIpQb/Yr/pLMekkp4AhloOlisarShKCstl
WxyAVnPB46rQhYs7F/+8hMUPh4jB1TD5wRfJBj4ZylC/TmN5hp/w7IF45ywVEo93gFvkzNo8ztCj
UDEjW3enmFFKH6kBkggdB3M5oLlQo8Cau7AVrV9Tx40cmPeSJgB8Hv4ev0nAgd+HaO0CUIpiFP2E
sOMW3aWBNr50SmiZIpjPx4N+RUVdK//G5/XprVtos5Vz7mbNbaBnoqxnoMMxCHDtlqAlu3o7TWUN
qv2a8HAeXBl5M06RCVC+iOqgPTmUE/q81NlPhZJ7Qy5XA6dOEvHNitgle77/4EZ7Ia2K1FYqBcAl
uiDJOaE14V0GNxJO1WlkDB0lYUvHACDQdUDfLxJoyAe9XiOlNd8ZHwh0tilV9AWxRmMkQZnj7Yz9
myjOvaC/BvYy9f3hCj/+KXyQhQsM+3mpypefPReRtTGNdT9fXz+LZ+jSzl5nDbENhcmZa7/w/zCn
kX/kk7bJfg2gxujZnTtiQyup7bbSaXl4vEP5FU9b9tpvYO4q/nKLdl+KbI9VMF+0ptb0iCs7+jjG
ed/iYLSCFTLnL7yx+6G1D25Ap0dDXEsjFAgMC4HsxhKyiiiq5QVoMUNhiYyMxVOfvrFyxiBnd0r4
5NKbt1JUayv3bWHZnu/P0AFxOKi5+jU4lHe5+2f0G49HLLtmfKfzziA/uWiWyXYlgU6KWJy509hZ
CafJ8g0cgEpYCbqoobG5zCPbi3AUk/zFctXPGNDjbSa5uH1LzpvOEbsh3RUsYyCkfmjKW2ezmiHV
klBlSeZjcUjDcq/PRBLpEdTKGBUQWKo19uxQSBvyN7EUPAlGGhb71fr9YDipNxb3/vkQ3sfnk82N
E7rQGiZGxtXVL6VkFpZKAuGg9CoghqudobIP2P/OkopRr4/Pdn4rwjlHn98ujf+OSF6idmzJYVHN
CprxZDBtr+iA2uv14/XRtI8wPK/GcjQ8wph1hCknfrbhzw4G32ANd7R9sNo+4isVr93z0LoY6y5P
2VA3LpDXLUhCF0Icd9On/SScnDCf5Pt6O38oPeZRFzvMNIpmCOVfzjDWlVk+MIGdFaedDlFauVAe
HsLv+XX54Qf9k7MiQJ1xoQpXWF/sAA8FN6UUoNG3kcRhwiPfygu9Vbt57b5EUuMn+x/6H78CxFfX
GQ1J3K6MoJWPjdU7dTHLX0ontwKLn/frFzdMyhYdCZVj+cl5OyvcQdeALGQoGfG1RgcOQPiDLOP/
jkJCLQvna1/mgJ/vDYJbC13gxyyqcN0S+8cAbgrdTtdx9DNQS12FZJ6FJuK+YQ9QROwTgMCoc610
KAIhvuLR3BYDPwIVeSgv/c7d6zNm1z1N8B2FM5L54ms0akblQLFzVdl9WUJiDOc7nT7iZnCsvZ8Q
hUQmn6Yb/3RrJZtCACAA3C7B5JbWPsnB4iXnBrpTYVATUVcuy1M208audQvrFE6Fez93/0WlSL/U
97pUpvC8y/Hk+yO1W7HHI3OimnigOoBLu8fo9nNahLyPJcOKjnSXbJDxbLudc2GUdI5HA+5xa/Fe
wxT6UXB6hUW2eS/3b0Ats9LmMEIrgjWsH5jXmYY3yBmdbtqupf7mtSexv/TfaD/ANLg4ASqA06R5
uOtYfhHL245WKUpN9DQaX3W0rtcXqduhVQ+TdMdlWLjQkvxKBp41P0RVg8VPz5BBbkcas/9oaesf
i0iGP9/YjHrBXIjB0SVO+of5pPcjdG4JJxqcoVR5F6l+UOYAZe8nl8h65oPnEvi734BLI1zgdBSR
UHjNZyyzY3YI1fxjpAL6Mf24XwclcFvIsWEEp7fU9q+fVNHc/LUfK/AThOMvlUomcqDB36CFk+YQ
SECvDkrKup3lzHSXWaH8NMnBVkxR6+njzthPF6hu3/odoHwu5N7znVGMd/IIHO3kbzcxrI6m9VQx
rLYyJzsEFJaV83RRCl2//5PfSdtta/yua8Rxf/M8aEsrynKUJDwMAC+yZ6wRbiQb5DUEPTzxQJSU
Qt5VnWH6mqDJ31pgCjJ2RCO1Do2AwwOw3qwEdR1qnyjEREB4DiZv5kOpFo6uHqZy08Et6kizCxTG
Kd+/ivCdJvae8ITLhY2tJczCsmnvaB4pY39P22M7arZ5eprcKj00dg5bnjBvQd+IvueYkGIgnFiv
dqKjA6DtDNBQeWCIu2ZsyWtRyynKYN1IKz8tFMVUoM2XrfpJzurjOfLu4+uBYJTf2NPIMsj1AmAE
FQVUysMfQ3UYF4+h9Zri8lxIrN/rTCzGvfR6W7214VBRhii8T3Gl2fAWCBpjMWFiMAb706tXSfsG
dzSQj7f74eoY5sBoqJIIXzobb5cNEWEJ3yVYmXveSHNpVFftl+xe6ZaqknlPnsWGCK4KWWNJoAcp
iHQTw2KKSfDCZZbhpG005oznRR9Xv6Mir9Wyw0fFAAol5nguC5eB0su/vpvms5+SXN6ctVO8DkQI
DCqo1zpcGPtTSPiBZRUm5JXz/sbgf0OKnx9IcWG5AXVA5730AEapYKZAsgitlz4imlrnOfGQJ44J
JdIpOWL51xStZEEbN7PR2bAzZ77gcPxr9TCfne9K0sQ3PA8Iu9vpiFh0fv02Y8hf1fr9CCEevne+
lxnYqfIc5uL1Ij8U+cv2qy34m8t0N5HzdMdrKzdIaSCDFEhJ2he3wTJFL57NWea23NcJB3oa7MeE
zizFJHXwRBE/euaGzSVAkemoHNWJlj1Vr1eDHeDMtAb5OT82C+eGzwMZvTLptrxbiNb+itKIfVUx
6313MUDYcxBQBUDTp655fNYVMxMVLwIRU5IAjNDdl0aDnIuGThWwSjBV4GRq+BNXNoQlszL0rbd6
tAxt0PexMNaF9QBH4X5QjORLnXlcK54thNRjvkLQCmHiq3qEQRiAwf8no6BX6IHd3ysj/UWWFaJL
xjskiJOREofcyZNSxt6GSS5KYi0r1gKkjD0oq5rVeWerK6azHMG1XrZfFfBT2zAG52Ladh4kAY8i
c+Lm/VbstWudCXQuUYH7XCtmQtIdlxMLyDIV0yRAO/BYv8ePQiy2iL8VvRqf6VoozkJpT7nQCl6C
o6T7/Q94oUIP035IoISLdYsTGlC2R0FufGgE+2oRvUoJ55qlmQchFP2G3LMkNy7D2/RNJgsnNTNX
UOxzrKreqgtt745gT1raE4f6/bwsVOM33MZ/Ro+S7hex0SWB7zvU5Zescydzz6tz7JuL9uPbeJrk
5YI31i3pY8FG1Zze5k/bgE00K7a/hYtlCS/UwP2uZjJCiN8Nt4D+6KgThdqgnCtoe0Ph/YXVjCgR
7qVdZEODtd7mfxs5zYGynTb2Ag+V3K+O+yDFrIsTfDloza+8ttXskzk6LOqb1a0C03940DqHes7G
aL5TiEmsn2n8NmPZrdDnMgdBkwllP3odazFYE+RkH3slSE42nGZyu+c1EXHpuNQXiSOiYdFpSziq
bsywftd0culTidfcjDXTyFPKaX/RJXVXvKORR8tMe/Xf0XFkaXv/fanpmvv9VcEIWzNT4nMKHKWm
Xv3ODi9EbxxObPC00Fi+yOAQQDdgvKK9yyYIP/j/uq2fu11B867ph8dLX+krUaPY51m/IE6kr/J7
OWUfu01/loxa4jyUE4W3B4hEKRnSP/hJ/Z5TCTGN94+TkYq0TaOMOBdvqpjxTzv/Rh45rtXIYrtA
DN1vQrcVlxqb1w0FIJO7SduB4Inv0zlFe8Vo88HLUSfziUPOou9X3N5fnPmN+DG5yAeLqBAi5B7z
v692X/Ln6in7hh3Sj6ZLVqU6/C11nDGfYxKzNU0L98tgunQm6BEBxlQau5Fi/AMO1kGOnWPMNJAd
LE4sJEkr3KKHLGWT/Vebl1PoFWpn4l2Nlz4vDDuhXJsSj266iI9/g/LluQlGiXhGgAZdAUciIttq
7FsfxWzUiiO/Jr/Ec2yTRyogrRGP4eo3Wl1jKUvgj9uR46JCUKQ0gIjT1zRax2MtYJR66xeikW1T
7pXPmKFNVtFzmYOJZimpMZqb1FgR64FSLRGzaZL/e9zD3BNwf5l7x8g73ztoEqme99Kqn7/GpciH
BjIZKwepIYNQgAFJUEWGDM4F9tWR8SIDr/uFl54CJTq5MCiZ504WMUWWnj8Y8NaVfhmGYg4YSPDm
PPx7DGYW9xx1pRQf0j6o5O2KD+L0J9XIsHxFqq3klIo/uXWkCp8d+G98dXYUvNZVG8BrDPPpZMKd
017HhN8m2jeDn2jMwYKc4+/mgIIe2Ouru7xnvATsLT/H2uFMQxOlllYd6mYTNNhjXbWWiCkHJEya
dMbT0xMMksN7AVX/UCZ7M74cV3eBkcbOscNJFRnq21CfOJTD/My1saDjddKV7VtFIMmdJUmj0QOd
0IlCL9UXbYbSvnajCeQfGxFU2TrfsBOHMeFnJSeZZ7+qFfhbPa8sIyz47js1wcADSKrbFTgESBVZ
uajMG/JFFwyoYQ4WDa9Yyr/e7ZRqVLykp8zNq9p53gvvrik3b6oxYHtSOBbiZC1P9Y1KJr0FCFZx
zWl7Umzql9wsOg6IBQ+rD2JkqkTRo7YHPd0zjo7NH10lZmRejnlY481EzqCZQdVBTH3uOODiJa15
1dJppd8NKKclsJ/L+WLDsk1JuDRIDWT4Dg==
`protect end_protected
