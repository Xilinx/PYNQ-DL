`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner="Xilinx"
`protect key_method="rsa"
`protect key_keyname="xilinxt_2017_05"
`protect key_block
g4Wfx6Gh4EiFMhn+WL3JYVc3RL3tUF5ErijOX1M9IDTf74/02aAlfpaMw9DJrhIK1b/o8Uz7LqKh
u0vYpqN+nUAkUQgGZLRFw8NNlzMI1uvuKDA7esMNJ7f1l5H95lZiNYeMFw4B3+mggR6y3jHJAU05
j2i0OJy9t1TYBq6lK2hXBOIKnL3LY1HddwQr/tktRS6bLVV17MCG5DSX2XXqMSaJR3Nxpa1KsF0H
3Sh/7EpsiGQaglDEQJ2mLt8EIo0akKotSMduzzTKw/2Ev2sK35GNPHkv4utp0KyLdfCZvpoEqQ/0
w6MDuNlgd34jbmvnxbEyNYUSbwAZwXI+RjIBGA==

`protect control xilinx_enable_probing="false"
`protect control xilinx_enable_bitstream="true"
`protect control xilinx_enable_netlist_export="false"
`protect control xilinx_enable_modification="false"
`protect control xilinx_configuration_visible="false"
`protect rights_digest_method="sha256"
`protect end_toolblock="uQMKD8xU9qCKoGHE5VHuB2ngMivjftLdda+IWxjQtl4="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 49968)
`protect data_block
usiyiO3cmNTnvnG+nvfWOBEc6OLtouECY+1PFUA0OZp3rxFGcbeWQVKZeeoIQfgvAM/i8gPxEPGT
s+mrJpyOM3aFTA53AOUF8EIAAsUT2Uy2bG1QLmkN9/7Cn8o9PjACKWu7LItfIwT+k0/qMjEc3Vl5
IWhn21kcQMYHcB9wKnRALsL1TZnKgo6UYqAXmH4moKhkPsieSvTguWybLeyHLv+3Ew1xyxUaGBCl
92+qjVdlk2w+V8hz4bHWt3DLZr3O1ABsDk3ufFMCvlJs2JbWEL92U943D7HxDX/0GjMlHfYYOaNo
hZuE40c4e78fCge8kTVlqvjY6fr0GCIDySSUwquNMAX0xszwLm26F/BiBhGy4dn2EbqppaO//TOS
D0o5uK2pido2CdBnpu6Bv3xilsDwdsxxEzlKo139ej/Tiuyq0nSqcpgvN6mU6RbZGz1+9uxVz4Yy
JrsSFtWzdtKMJZzdrwNgnCWNAB100BLV3+oxHEORBFBPZHiWTalLj+8+Yg/5nA85iuRTEU+ui24d
EjQr7i5LgC7TpsdUdx1SHHDPaKzuUTMskN/QmHq0CRORNSFqjeQd8PZkwQo7KpM70xHiRlYH7ihZ
MPWbjxEL1GVSDPTW72Qcvlx1FmOJ398jLD1fONYs2DC6nAOukFbzRouikK1aFdIimiTIyI8VOI5v
9zmbIFw3JY/Gtoi/rhdQjjCBgzUISWy1KUDxngf4B+kGCo4V41R25YfVfp4A2CQyEdQycuIrwOEC
Ee+NGeu1bh4+KlEIcIm0+1jUXNE8HHZ8MwWHNzlgOOoNd20BMo7H+XQ9+PeWeZ+CN99FMLJbeZ92
sHjdDyccCVq4bU0aXndvVPBUCPopgMlh1OmfJ1umgOlY4B5yzfcRF6Jd4ULBWc/Ow8JRDTTAZw6S
HvzcJRZuPTmjUfuVaeYDSbahZu09Zi5ZryzlQUaUzd9wkdATdqFFXm7iWlPoJ17BlU2/Nnq4phaS
CkPjv9U8kGxFyFFACdzRctXR1bVZ7yf3/sSgatzAvd+biBxufgdAJugE/WKhQ3kAKwIsDSfBb8L3
5dV43HakedDNmQ+2IIFlvwBQp5XX/z93Nj3KfP+UVDPF0YWsGISKyaXzeHOZmR9jSoHqlhuFBEKh
RHHkdSf3eoiMd4Bflnfgm4VgqL/W+fZIdSdXkN6mFz95Hf1XaU+8PJEaZXiURs7M3tVC7Pzgtful
b2rMKP2IziLsJ5TEuSLLWWKgUAFiVEApKUrsejRqdNWL1GgiXdNczh6iez8b+5EosDONtlIhFQ+l
q7BHmH/lwCs3MW7YLb4Z+Cjcv8W4Shj8DLyvuSXv8ojNI9/yObWd1OSW1zI2oxubg9pJTKabRLKb
nNystqKSbDmdl8OsKSEcEgTiS/jfon0iWC2Pr6O2cTuXANkdvQ6YDqYwnWGuB7hdFzzUTuEyrR3W
F4kldtC+xvOrdH6VzfUs1W+fb/53jRRsdmRd2qmi3pBH496V91pqQEXuul/+j4AjZLK6SsmMV51n
kvuv6wgfcxakfd8dRWt0GdajabXuFQESHHiJsWGK9Z4HmiQ40VVDtZrSsO+Zp5Z64MAVKv7gSI0t
Y86GpjztfPL3TDtkXeb8YErjx/wLKaQcLdcHkv+BcgtCTRT+DiCNI/D8zBmVfNjqp0dM7Ja/KPV7
hZ/sLn45UvPRsgW9Tc4nFQZRDOVCydHPbiTu59HiBpFCdLp7u0HcZlomukGAZAqkhzsLLcr1gUjA
FKFes5E4FfUrA0jpadwPyp87AeSJQ1xjCo1rIAzRtsLoMkEw7Fhix/Gla1ydqiDSmFlH0D8lRrBW
VvzdYo6i+hKfMj27BAzCLRaInOQ6exrthOwg3FoNMgTQzB9z+SDa82nm0h9Z8LFHwWD7P4yuHA5J
iPu7BNDsreFyo+60Y7VIkY4JcFqFg1OA5R253WdNoKP4VnOl8W3/miKTxEJlAeM7MWzoxRm43Sn6
RJcOAJp7WvWmO/u9v61a61XJ5NChmw8stdpeO+xRtqn3qQvuQS2I9rg49JZdERRRP/barLzTsyYW
6IRZiOT6yySr671VDxUpTK+N70RW/Ba8Hi7uVXf2L5ZqtmWLGzjrw3UrnK+3ACy5ssG9X+kKEuGU
/zQIFQXDu3sc4yK5MTSGMntIxHrXYiN5LSgDJgsa7K8pmmjbIsJDdbhCaD4P+616rrMiLDrVctxK
hjS6rFBkRdIQxpfvnWBJI8SQhrVtFt+AU3HRYSIVwq2+sYWuq8OeYqSlBTEm85a2v5MVRC/XUFDF
p1FFb0dKdnDT1VRbL3sbSZW2iF184P7Q8GOxs7QrV8QNAbDQh5MBfPPtl5KwNB24Rr7lyBZCgMyA
QLA7TXfOzepQeR9ZvXcO0szxjqrMTLGwjSPpJ/5/oY/brUCsNWv8bWthZIJXzjB1tiQDuPNA6Q7O
TAT3jsoN0x9ZBd9j72XaSbHOaVcaf17hdIaHlDV8r1kkjCo+beHJyG66S9+QMSbeTYdOAUSyQyCQ
/tFug+Pf9s18D5BG2JCnNTeu1pS4COKcTzqaoMIg2lWm5iaRdiHQ1RI3AVtznuEHdntTOM0DjDm6
XUuLvNYa2Zzrea5dQvI+Qx5iiTjyXfYTdd6uvyD1lFEYANPpqX/iRwQFOd0ortI1Rk9ac+h8iUpD
qJrS54Me95JOtNWA3s3SNUdmr5so7ZJGivLWqJpmC3OhsVzxk1TsrZctLijwtlPCopMhIPOr607V
K+xazaKizvf/oGj249GfZt5iQOZ8OLdoptl39R6P0qEsEm96ZVHDTekBDDipsyOvYc2Bvm4T7TAc
jGTezS9FiZMxFKlr+ILtfcbCmthlOJXSGWSnfjPxSXjJLS9cm9SYYaxbgTWKM/kuFN3q0Ot9ThyJ
fOoOCtj+PAzipluX35JUS8WHHHhfISREW5vGhHHV17+HzeUKizJB/aX6qVW+AQvwE0Agdfdg3jcG
UDnG2PixAILgEa81kGTYYqpDNCaoNQnFlGxgDn5HaCh8gje6aQX096iYY2usVvIj8h8ygd2vSzyJ
NbajIOciOL/r2hymLxZMxVyP84pE75opCxfWoEcr0vtZENhHBYRR+ESe2/4ekH79kJMYAXpLuqDE
ZTGl9/2mNgSWj6dPBAic1/eiuU9DNRMk3SCYjm/mzFz4s4gxCSCu/U+QELzyhZgT8XU+grpbc8lp
JCqDAOQRwkpnMaapxqhf9gfyYhgxUgSAk2PSsgJzX67NXYvbgapNEdhVS9XojVCp3mouOm+u6yod
L6tbZVG3LNo2sgwe/vYx2/Ft66uYpYqMe2RcfQ8nRimqH1VWnVnMPN6ryRAzjOfAS4ubu6nHIex+
gosL7kljtlKl+Nd9er5fmYNZ+O9b+idHPEsmFKc8uyWD7E38wc1ipilfgY8tjDmr2LF1mCXWNqRI
oD71K/rS8tNw95QZVeQHTKXmwEhXTSfMPPytCru5f0ol6L4rEE2A0V8eVZWTBq7Nkn93AVYPAomz
Yy/wRlNyOhzjbRSZj1HctZGdpWvyzmorpeZA7zGIPLWJhP0Q5J2uCA8v/p74vQ4/LYDgNhNHOyE0
Wrtc6dUVWnocuW6ziVSSvWDdWysR5zmTJe0zBD9sL9cge6Zulnl0d5DBZ5E9QjG3b05T0w6KfCK9
5swVNfE9GV5+MNZPjgWl5Md7pBO82NOmRu4t5c7JouXiK7T9rpsBjTK6L7PMlVVbxmWsl04qt5z7
b1tGy1AO3Je9EuwUC1rreA1gDmsop0WhTRbY/TCSwl1cKs5pUhjFZ9e2/qrT+kHJat+TpC2G9enl
6sAfdil6zr67nDehz6bmTo4TqKLlYB3Cu5Y8uSqfD/+1gRr5uIibT+bMimEpou4RI0xP0kmi8UhH
rqgmCRil72Ujpk4IG/jYukX/kJWoQFuZ0+b/jW/xdv5WSb+UlDaeM3QUacvD3fIfRDQo5rwQbQj1
Hh6O7fJFA2vlVUlpknza9/E583pEHVHMEZhbwNfJsDvcmeOebN7TrbSntWRaik/T+ml7V9j7Y/o7
D1OhdpaTPg4lbXeLYwv36N6zrChWSlcXq+5+BJgWmu30YKITTEEz1Ct5f0+gsJMtwdbnZ2h/pLuF
FSGcEuDohSHVrSuhUyxTWEdYbs+KCxPs9gisGWfLRb2iAEPv3AyL1sU8ob66V+9eyj0Sbd9W137S
MfheaS/OgdGL8vA/fRZe/K7XGygsl2I2KGMlN2aLd7iQPEmjDYvdsCZzBLejlmK9vU9ZWRuGrAsP
FjPhiIRRFIpKk/Adae/qgp69F3WDD019OYPf2T5NMqNuZMpRtiLE3/fEhHmur2CCyDXo46nIat4I
gX0mcAW7jHKIlKdj7cP+xvA1oH7kdr1rLPhVWs8IwFkN1ezysW9IE5G+A0npQsKUpjUz4FjgppIU
zNWxktHq/odSFgQTFj1wuGNPUap99bn+mC6EnE8OXU/c3D3KTXZ9CvIj7pUWfjTAxqMEjCb56rWs
fmxh3OXEcbGaIJTpz5+ZYQ1B3hQzNK+7pEMA5JNem3wdEMu6UUrVnS6kIiil6OrOEiwX1yudUfhd
vQKJZ9Q8IDHt1ptbHjkAEtOXcjI0aU+cHWVq3rRABZCe2BFYVL+53rJ5kcEWPENO9MN3p4indVki
nEMT8mXte5GZDCdRHbgr2pAKsYNbqq1tiIKoGN8Ldt5mXU8wDO9R+xRT6EM4F+iXY9Hu1hcXRvWe
a3YxMdK52mJoJdJzbqhNenjdCpP+ZDJ/EdTPEoKl0xUNFiNI4/UY2Y/YTQQaIJOyyPXWwozJwIsT
SCtSck4CEzqXC2RNryWRh73Bh4PzI2mhi9kaaSCQHG+H1G8VOwYIRGJPJscMl0qKESLtTAjVqiHp
p+D8YsqhUiL6wamvjJWZFWRPTKam39uDZszPQWaLZz1EEMApuAAWupITUc+VInydtRAVqkQlY5NF
3mwhpdokRJH/ZvNL7KXvLt+6RsuLDEkYETeNzKEibHPVzwE5w5Ijyge64abfEBxzPxXIumnxhKKv
V0hR8a81IYoBgGs27eliTsG9l57M544+IuGvsyB0C7YORa26bb+jDGuXOw6/HSQrJBmbQuRrKFJm
LfDerwNwVSxPD5Q5D4uze9SuXczB2LE2iTTC2X5dAl+TaJZtc6kEv+nVYLKAK9SGA4952PODPVk0
u2RACgB509BSChy7UIybYtDA1g8MusA3Ay0HeQ5HQM2bBh4nNz96Gyxmsbe4LpqAcfh1II0unMok
T7ZloEAs2nRW86VWeE6jcCITU/NCB5ksB+v0sLB93hhtTDtWLjWFxnbiJV5DWLswuTQ2Nx86BEJs
XvpqbCVPdgZiJ9eDUFPx1zc5lK/sHSubiDSn6DE92vXchWYiezqfNMu9lRyUfIWUIqU34vMixvY1
7Xsox13v9brpq4zrmZs9qftgNflW1Od42xuppSe8fhOUggbz+aHg7Wg5c9QxFzNcm39Q5fg6Q7Gi
xevI6rW2ot6Vh+AuSbheZ37goXKn1/B9ZBscAouhd35HjMwpSjyWj9pubxSw1dHjEQv7CvMpycK5
rf/OiURPvTAxsCwsuL2jw0pgLB/nzsrvPfhJCf21kxBQoAYQ4zpF4NYrll1eZDhVuGhPm6rNlxN1
MI0C9SZcpjnrPEXaWxsP15ruiGUfJrnxbZEwyZ859ASBTEkng2PE/vov8aS5FT8TdJ9DW6/HyBuq
A1Pt6JuLUwKbq1MK0hEGd69xEjD1rIhLsc1Nw7bcixulGnpMKmfuiICLBuoFvo7bjmih9yBO0uXm
GQPGOKycyV/zpZFSi9bO5kGEVosfyp040ZQ2JKY54DNuR5zTgDSqPIoV0M/aRYZnIs18pkW20lMQ
Nv5UXBpq/1wf1vx7lZfLtHKK4zdc4lTGKvVlMdSfbhkbs8Be5vKZ5XSIiQXNoLWVLVlZEVRb9q0Z
ijusiL3KSOXZBmQgzgDgcC8KQ8qWku7KK3Y50qS51K7X9EBhwQB4STPFSuzDRqZMhHSV9TbRr+FH
DjwjNRNJbLX1LEak9R6EBRVYTw6Q3SOOb3OJ8N8MVHuCAVXbhAzs9cpOJmYbQ6yl7LYyVZ2Pi2Nf
hOEFHkEMsmq1EDYzNo3rwPUHnkD7JsjsZAQpZbeMKQFlkyFKLvdD7Ffky4AQK2mT8LvmynYcPkeG
IEx4asJHWflNo8X/mXzZpMhvPC2m7EjRqV5EcCusBy06zSjqd6K0+iJB3DCuyLf1ypVPHUBOqT+O
xs26XsJe8dntUB4PhwuimSFT1odSR9YAa5PB2bkX5OqS1YRHW6e6HnGngBsM5kl/yejsAna7p3w+
MsWMmOCzheAcw7/tefZhM7qbuhhF1DGH6D99pz/iMIyDbsKMb7JjRxk1NBkqoKnThL31vskPU3cK
XUWaUwxzrhvCZCfCoDTq+9aSUhUvlKJoplj/RKoWD9UABsudDs9vStpoQcdJ16mTS7pLwqBzY7cp
ukxixGLwQ1UUMl0jpMseLXS+Euz/t6jPBgQkatKKDOQjAGMI+VxUR6LrYzaeJ8bzZRz+5mAL2w8i
hP2WAgBc4B20WoVvcL96m6Q8/o5qiuSRT8rexiIUxMVwUCUqKz1PSZja1uX908WHlgu6RcBd3gTb
wER4sM0hsugr7RGBR8cONP112Z7GO0OAhqHuZjVphKqYgS5Xw/Bdmnhz5mX48VEuNFqaMgsN0kAc
KLpzcldhDlkhtTg/o33Y8UIdwB8aHoFq+5ANjbnR28NdnWPbcr68rqhYvfF3geLa+1TCh1XiuIJ3
wJM+aw71MtfViv4oUFI6AnkxXoVkbKyPemT0oIDqBqvlfwohpDlam1faK3nFq81itUwoLbLD2tCT
4Fw+09p7mvssR+myf6FeBdJd5QPhkIryWVMJz7tdoBade9G0fk44Asyk8Tjm1uA+x2UKshPp//1e
cQzmhIpSfZsC9nS9ttLPl2WB0qVxzPJL2MtFqCjvqBW4ep9dS76XOAg+3GQXq42CjT2/wHJnFRqi
rr8hbd+5f1Np1AsdABGp4ZrzYMrMAiWIdFSe9kIdJJaECLsLlee9W4YAlziTftqA0TBXOK/vWnHH
SPSVzpCZkkiOZIgF0o9r4k690Xa38FKNLCU9o0CPQ24efJC7S3O+xwOFW07BIIcmi8AfNXbZRwsG
6LZPIG49ZIHjxEaym97dQffRdaY5R4oCIBrqt/0XLkVcYHYC8s+C4yxn8mT6K1l53VBhwVwbzul4
Yjllgd+hT+wjyh6i/gYyT4yjxAADjw6xi/pCJUMpyCpFtzGgEq10XXXLaqcWTCA82TokzHyc5e9/
Y76Q2CQTWTVmFpfvxZJe4bzxo1LjI2I7ELdwdm3zXF1LvvmY2U9s7k+BuOQN7g/sIK77c2SjxYjb
u5kTpIf/ODJOFqIboBLmuMBoa9EjzP84trkVICnfgrcDnSbAUpTtpu1SnnFp2PU9vtd/C2iwgQea
0uc6l6dhmCmVlgfvkvwop4QLUh+6gYdmD47mkOA8Ix2j0MWVOMgEg3rjeZd9WIpXX2+YCHtPx1Jj
04nwOn7x6IZVFMuGJdkZkOljnMDk5fdsD+iXVBTfCRuQ0TUTbkyFIGEEUF+SDf39GQ5eGTScWRnb
b53x6f5qn6YGCikx4OEZTgerhDiox7sL9k4wqlUi1SGB9IjN1+WP+v0IVdgYQcvHle2CnS9kLa4Z
yAXNnAv2pGG4xB4QcAGY3pTar9cit/MZ8aJr084mIvwHVSLzMkMI+NkkKk6gznJiG9rW2xEV22+9
rcAFfffoVdH6jZ+zYeIau8ZCq4LJlHkQ+J+KoGvXRYs3dIyxHewCQuVrC5bhSwxNWGRRbeCVHo+l
OnL8O9Qn60wsl+PtShlPW6sI6LedSfICcTnHgL0/WoHqDN9JyY3ssn+RlvjFCei1E1OMdWh57j2I
HA+nmQmxXLkFSHjwKcdo8eTfm1WQIoip6F/TCJTWtg2DEsDUj3fPM0uazUSXjPW1uAGZmmLIghG9
57uXj3okzj1TAvsIuimoPAsLDK+41JaLVXeP1GTKlu0P9Ey1zjrTQZmn02WsnuxC5kOz+Xeu905M
yjmh1bsnWynklxBGPJB0cM4LF121jvaw3J/nRxvUkOvocqgh0K+u+OzdGvG6gGJXSREsGo0f++sB
z9L1yBlIey+VM8XuiA7BWuqA2s7gWsMEswshlHE/gX/SF1wIp0Jxr8nyU3tvIbRkK9Njpgzj8WAt
CkSZB7Myd2qhYYUXJ4GPgVMNCXvUQcBOnqkZaKC/1MfVq3bfZStyxr8J01KpeWmnxYk2xpL6S3+S
kElPXHrirqsZD3pmN9mGqB8hRHp7zfUkQoO7So+fOE1Z68rpgz5rd4Zgd+PI8JJKSICS2CgEEpKX
FEJHM8DKAW779+8JT3GMsR8JglhDXAzUCmpZYP0IGPwiZOBBLz/gO4jqUqwohQhlbDJyTiNCVnV2
y/vgcMhMZjNmnn39mPhActFEIVa9ZWxR9IoYWBSpiKiqFZjAWvE/JuFtPJnP6fc+HTIRMQ37uvBC
z4F44koqW0iG73fN8SH9U7xmOpbytkf/y/pqVsV7P9XZk5/48ZcV/MxZZG7h8rojmq14N41FUmG1
VS4EnM9M0jjLiqlNaFoFO67fYC82zAZ5PAzdGRGGDfYEIuGc705NFQoukSE8TYXbqYgpgHe6qBYB
mHZ3kpvndhQmZ17nkTBwy4mmAQkRRsmJAFeBuARC8/x93cwFHeIBeHBdqyxM7NPx+qKp8ZzoAV3h
gOHmH+i+mEtVCExVq3c/HwxbcrMZ+8mBZH4rOXuIkc/XWOKEp8oNRxomDeqVouldUnyBRZNl+kbF
xRpuy0Yql7EwIAsNbgp2oGgLqkWi4xIGcuUGDESdWhs0cA2aOD8B4QDudXbFz1cl+KOZVtaX5uIx
WTUQ5uYyMXLQi+58TFpzpFfOw3qzParW//0X06Q0zfQXyzkKCmeG0ZmLOT1yfa0C0w4uTHaVxfN1
W3pFy7GnlTQFnm7TN5LX7tTM2AETYlCW1nj50gPltWpEvhRkrVGTjLD41fitwsNLTCpiqPlib5H8
4R7pJl9ng8lu72DoS/EC5tvKREaO4Zxjh2GOQYWIoUObruUeEWRU55DnOP2fgOPRFlQxQ4vW5Byd
2jqFiGg2n7TOGt8kpEZzHTvLs8pQHedt40VswYAeXw9NQ4zZ83vjTabaPrBLCfneI2P8TkjnbiMt
ujyq0MihM2QfYRYPlwhXdEWtVoQ4qQb/Dq04w74s77dN5QAnXMGzkOFU+CiWUIEW1uvlluyyjixn
NCGJgO4zgGoexQDodSob0WG8ujKJ6KS9j6ecWq2jqsn1CSH7le7mnPfib6Pwq+Ya+D1stvaZ4OSA
+ksna8VNxbuQ4JAjv+ipT8OKOIXgNmnzn3yjGgAWAHsoZHFy6LbqzTQNKwbZFbXPcBVDF6edC+N6
G1OI1QLjeN9SrvKJ63EoPeMIOaFNCIEPKabqQ5OFRGzJIm5TKmuN5qxcjla1mABXrw1NtYCeiqGv
Aa2Sm1LlS8R8FNSwoLh++KxPpS46Dkquvoso6qgo3R1uSfhrE2Q0tnezTDa3ro25illwZ6MVOVOE
L+ERjj3Eo6GWO/+FEZU9Y/GkSHL9+hsuZsKkzfqBDorzdajN6W6Lmk3QeTHZug5a69/sxEkKfxAH
iAnLYfJAvui3kxa1CgYnTw309GHZFsiNrHDmFaWFoODqwfNjQRMi6/blY/lAoghx/eewmkGgRRu7
kuyR5vwTnOcisJ3Zgmt5F+lSEx9UD0tpzBnJ2YvTPcRBqhR1KQaQh2oakBjmec/jrKeqtA3ovxul
512TFw4cyWv1euVUfXLZmFuRBVfmzCqaVBkv2Affwk7TcJHEqOrQrDnJPNzV6c0RYhjPVOGV0tgH
PtNC6HDYkpVZAtN3Fj22jcOFKNjBsHy4xXj40gPKzhhddus4FJ2SHDrTjX3YNzJ+i01FUSAhE6a4
3P6KBsxxm+e5xFDZWyn7pn3O4XW0IB7wtahHDQ7VQXCSWevNMTlJ9129+5Zo583l0Dpcb4O8/Rgu
zl14gsLuW/Ubnxi7Ts3tU3dHdToN5StcDLt9AqLNCX5yx8UwSgMB6MJuCwiuOkG8NXsX416VVzq9
P+2+J3cTZ6NpC8UGBbgD8jj0Ffsd9dYC2UzUeuhTDOICfntujWkZo1EYtYYEvtGQTB6DR8iJXHhR
lbQwGaGm23orepqQfLXsJe5IcXC20Ryz5K0l6mlkKHNqNCjU/NVwRKDVnOAxVN+9VjXXSwTNj5+I
XwNFd3DDR8lK3F3ldh76M9gZntqWI+W6hJ0zpy+z8Y9Vn4nvFeoN+FTfLeBhshzX1OIiWX0kqE+d
pPyxZJOHJ6L51zLqxGklPazcXDb0X0wFADWOa94uRYDCI9kqYSk9fa2eGokqZRTLZgwlHG2lLTeC
GI0tlRaR8xzCGGE6XX2/EeW9MXIYV3PzrDPO2+ooTZwK9B+rmnHeWVqftypEMNz/QImNJ6mjRF3R
bIMdBAtvQt7B3x0lmVvHu+Cw4qgmsyuqx2P32uoD7S5nWljp8LBS3Q+h3WLz9OkbFaumLr2GbKq7
CXCw/2S2nkJIznCvzjdjd9lT2vu10GDz2iiGLf5wqtQslhfFXTc4C6gz+UqtkTxsy9nI7phhE5p+
ABaLU1rF8U5df+LXu4wp2T5n+Bzb69B/yhmAs+kBTineRZKcul/jFmF7wjVdTW0xUm+6IzihEuLo
R2kY3Wpq7A4OL9guI83O4Hb1/YciiRhkVy4GucvfqxCFyeJ3DFJtGSM0MdscqD344DaFixVuZNHp
KneZ+9dRj8CTpRTs8LGqPHLqtv40zI9Kdk3hrwkU7zGUx+lJn24D0grNcGbFf7+KfYV8H2BRpSQA
NX/fCurUbMOF+Qkvwy0x9oVR9ptkPpP7V3Myp3Q5adWNk0FSl9kV3l3tIgSPBtD6jO5O1o6JiyBY
zejP17VSB1gltNFfpUZU2BMRagCfB07UYfjxC+QodXvF+OhlWhdD0qMbnzgxCi13+6mD6YTSjczC
BAOKZJGGy8ogw6qKGvA+NsZbqbxYrp4vri/P7rED9nnTVjlyWgjqGS2Yn2IcTZxqAh3Sx57ccWe/
vVqBAdYYx5NP9qCoRAo3giXbReMNQGnJGLsv39j0OxXD2tbF66IQulrqfa/VDJPlY0oPZaaODPkp
Q0SnQcu14HQDz0JCHCN4cAVs/wCBajOPlVo6XAtYZMxp68XFA1mHoeaZiTR5zg0X3tMghi2daNPV
v9FzVRspxTcSXlWIAK5ghZ9zKUOhOgSFfLp+yzdFmJV8mTtl7Wy+et2WnUnphxcv9JK2bkig2iFu
NWOwp+FmOiU+EWqyY7843HixrOfW2qN9pdugyGvjFBP1jNK2tkcqet0ZEkBtEwvj2SPI7JqU1DcL
iokjlGnSySk4LA+mIPrSKWNtYgUOtKZp5j2JLaBLngqKeQ06CnmYuRSSu4pTIkkRDV6xyWEEUPxJ
iH0bkYZTU5TiEiCEds/mgujf/mgnHAAoQZheT9Qw5/AFuJKx+tyi1N5tI9B8+c9mcQOujQcZS/+m
m8C0Smfhi6vqYaCJ9dYguxh7lHxSPlLl/MQ6U+WALQSRVk3hV/AVF2znhSe5G42Ky6efrpB/5Ouh
frSH7oWKlHw1i1JhvfQGXlPx+wK4UJJik0ekK3/IfeoWy99pWSrIcYY9x0xQMmc2lYb/5M6PCGwf
npe+YyyzWydbbmnqpFz3ClUsMnQlzJzHgRUo4XmBbgfWleUglQRdvXDeiseA7o0Hk3dp2oUrexnd
r0SjFUAf7yQ7XCYOSegh5MeEjWaQO5/qEe7XYV/JivvGINOeDArEFRbebV09zojpycFgHWESLZvB
45WwFVyAwpmtOj+A645Nd+pb6pK6ke5t1bs7KLKe7lIOYnLlbccAhqtCMXYJmveoQ2uTxaqI1OSE
ObJ+5HJFZpDJ5gPu482iEe0EbpFuIhNEbUJYWC9p1meZ5ECtGizzeY+wQd+cFlzKObb68LEDRHAF
RvTU+W9aWck7ShaBTWJBxdJteUJilZU53EVX1Hi4pFul4UGEJvD/rTI8n0HGJZ3UWto69lYUNYru
z/eVxzv2rcMsanvhuXVKkMCzRt2sI0HkwrdOUOmiMQPCm6RupryB/qqQo0bNyTQibgnsMm+dgHrc
XqOxid2WdvbI4gKm3953VHXCr3HreriO5ZFrSTQv1+w1L1YGtfS6TyojUrXY5kExKFW3LkcOURpg
BAX1EWfxAP3Xe/GiqufcX4Eyt0rM9ZVkifDgAgQ+MddqQfv0+sEFvWnqtQyY1hn4+qtmAOHHPndr
Y5K91Sf6+5eijHcZkygTYtYxLOfcRMpap00b4e32b9Ke9DPGGp9VNc9HaXV01mG39CNiLSBxQQ3G
AO86w/MJ6TR5oI5DTnmX/rSwS6ZDmuAzof+rCz0LCBvCTPyF6kqIrs9Nc4FGiMm7Yvkqt4Jr/YCe
bkMzJNqNJvgutr1PFAoTa9reUIlwBzzCtbU7O0PTWk/LC1822ZCk0OaoD/P6nXRWpCnpfVcoAKIO
kp7Mab7Wa9j7hy4MQ37SgjKJRFwBnAw0rihbcPHDFihfY/VGLyDmfkl2QgQGvF8asUsnwOC2HmVO
Lku4jBesLtGN0xMyOhNcQb/Ft5pjj1p5svan6lojHx4Y9s2AwAem/AlUAeQh4t0U2QB4dZhzLc+w
XjjJWyY8Bw1uERe4jhKPTba+n54ho6MAXSuxdLNTZg5aq3xvWwtUQDMp0hFeEq7r+l+7FUsP8gO4
VSB2j4Kma0mVWV4miXWi0m3JhhHO9VrSeu7OznpEe+pWKL0Sd65orPCv/QxOy6/3rYc6dkuPszBJ
5uq/pmkYBPJbjBkLaxeUbRK4jzXsuW9nlI9U1vsxZW2cNZZuUgxr5zwJXgcdbnrjtCbl2koPKzNp
Ajt3pU3qYzO+oqVUgHeyV62UopdV9E65lbw4Tzbr2l7WGqMiSAvDD9g63XpS/8ZQmxueGr8WRa0O
4wQCSnAHp6tN3FVu9SN7xNKwvaTFbxp1M0Z862CEvCy2I1XSS7FhOKI7W+Wvb7JMOzXf/xasz82z
OfjuWLPaPhcoJOZQKFUz3PdCc0t1Ksu6+27+7e6Dsz4yW2stsi1OtZ9TT+uF13RQ9kgbp7ogbwzK
GRK5CIgte5eZrVur8TqLCoX+p8Q8CBHbdZ8jtQSgSxKatk3SVWzCqa+QKOeAyVfjTweMwyhdYkGX
9c2hvsHepvyaK3TdZyTma8MuqGuxswAzJwANsYIsB13UKA6t2W5dqr9cbw6EFuzgR/VjjobcQpF0
pqg7BYgOQoc6PYZm9uaUqMgtuDp5w6dQSyrwicSfWZK1jxHglqoQW67gMGmxmf7E5X212B5nnj+D
CS2WVpyxFZnyHx477sG1FVvVOtlMG9FTVb2mWR9XZboCBA+CAk8wKtT4zqzPlp+asLCZme19RLh2
R0Vk7h6y4F/IY4rlVZrmoHevviphRkS6b34Ozlw7ErsxNuNh1vchi9JHI637sLuHy516F5lopPH2
6YVwRobl5obY137/6S01KYcYsTmBKjkjPzWsF+6UNGCM3AIBf72CF9f2SfMrj6do/m4o0wPOARpa
lmjW3DMqyN6NIk/uaWrWnvvMF2GgX1/XRVIIgvwQWqPonmv8zN6bWK/IN/oqvlJPxbVsVHk7E2wU
usDYuvgUiNuYv6wjYYSb/kTeBzB1mzYUJqFPoLTiqFe4VpxgjvkWjVuZcMMG+mh+NDOVyqPH/TaK
/zsgm9fnE2USm8DqQVKdD4V1m7vZe9ES/jFzgfDEEZXaNthHXAeuwINb7U0Lxj1lqU8qNQ8dn5XE
0GOMGYoyPedRPq17A+PqGh4D1b5I52CStjWiAQNV5/jWi4WGK/EjaSJSYQwqT768TeSXB7hzMnP2
LII9qRKsCqJn1qE+Hja0kwuFCJHvzpR1mnPCQgZQgvQH8pv4ZluHNmLUSAnqoa9jt7A79AVZ/Mb4
a/9HOINNrb/W/QVaS7g7XnhPeFR8UlR5iKbFxDeaSl/APiz4PmS9lJkOmsnqa3L9/pq8lWI2EgFn
KsLcHD3ZWx15f5qp4E4z4DOdh5gMRrxbHEcfbjPX5WjBkGjHt9Lo9YS5/p2j1qPLyki0HdG3+PsO
DWXLkpxMdTTQsoi2ZiQwcnnZp8zOkJ5m3GNnkQZZWkwt8UNVMSHbiICNmxfBsoHwDjMv1ghJ6Gk6
Ku8NUW0KxJKJDdOYywe2z8QZdE7LdlcyR1by1gFmjd4x/SjuiNQ0SD+KxC7WO8Xag1A4XiWCTPxY
EU/dn1WhJe8hzGByaymPdNSb+KBs05neQlaCJZXgr0AmMJrBqO3s8KszRDh0fVvs9TnHT0zflLHe
bH4omke4WY8CSAkG1mNMzZjsEkNDnPCrQgzhFRE1px740vikD+HkmVOgPP/dgBUNCMfEywKvnFvA
uHGe4cLxUQULNDEjRJL5H3q7Q9wKnJRw06MFFDy4d8WMTDZNeFKJLQq3r+PXolLE8nV2RfN3gRGJ
B6YS/3o9BYfOpZ/usI9wPvv8XKTKZxCJuZmsdph7WU6n32BntP16Bj/a7kai6lqiNK04Si3rheOj
qdzBbDHv5kAnVypXPzwyZl8NAm9Rb9SL40+hnNMVIWhxfxW9jKSFkC1E62GVmaC6AvDoaR6iU07S
L2wbCjaEWIWnjM7F+UprVFJo8YHc25gEDo0gfa+jMc2rd8rfLn9WQChUpO/RwxlDJAuDFa7FTeLb
9GpuzaaXAAkre2j9aygJXOPexKpLsVE3MPBEYW0apfcfBFcqwufWJ3a7LtmdVmrfw0yIcekKZkpX
6AMNk7IpL0F1AG7nWTb2buL07APxklzvZOklaGjhjXr8uxBYjyMSLP0CPeMKTnwpnm/V8jDASSP1
yVVmD9eZBSRFpu5WpLBKUjRi3kyQwyHEV8m61/DXzctpauSvoBQxxjZqWmi4ABwEmuTQ78LOuC1u
KM2eE7lI1kjVnnCmtCiRzu7y9ysuW3CiMbvIzkrEkTdiJgB0yzDEsTNMThxyjspLOS8CSDdh4+Ro
mdOXMHau9wnX49a4h+G4OZUJvGICyz/MfOwOYKVWE3mRZ0EAGfsVAQyNYwr1b9snSPWyMdaKxMZS
2+D3jdC7nY3vHTsgTF98AkeCVG+8K69CLh035nDnA6ncKfNjg3H1t66UP3zs5k7qSOGmV/CHurY6
O4Srjt0pYKgXRekA7h+W2Hd1YUBM8QEkjJcNjPHinUT7ftSaS4QwNZ5jBtd8HUYp4jF8Sa8IZ0Fl
BFY0A1I2eOrw4YpYqozYP3RTGIB7nwd6HpkhWCMKq65FMm29imC8RRiQeNrclKSjBCAl6eXOHwWK
5NdpR33GcjFFDMOkvCpCjLSHPgXih8DySi+nEWm4mKwplVfyBrA8SuyMBeARDN/MeEzMzyHzEdrU
QL+CkBq+Z7UVRhmPs0f5GWA9IHknB4VX8rZ91hmWg+ncnjQdhQDQknVIZf78OaZPD373mY5+va3G
/XIRpsqwDP3JXgCdYW63/5uIN2KkxqX/Y/pT/NIVHIz4bvRu3XfUHKthZsY5+jKQySh6fFMEGMCb
2uE2frSoM2k7lxaGtVEH7ILfDIl6wOMnLXTDQc7nTsCW5c8T2jwBTcg8i+Hpa7+B1RlEJREkkJ5i
H4156+VaMwJ/ab2NaCeqDryYyw84+gfNNtzECiE3VqwoL5KAOpvvwTbSPCYOL9mMKMjTM1En24LY
c/vQ/9gsiY9YnBZoCheaaqB4eNX/MToSr62wceLGPBiBLSrK1J0feyfVGu0y0kUpHKIZsMNaFONx
2/jC/Bw5R/l/ZcVfgJd8FqJW9dInoSzqthBXG39gXj33OLBqZjg65ts0PXhU3xnwFBJmFqLLL4T8
TpTRCWoO5fYoTaNmncKOwCw+EuHypkrj85FU+jYZyulmX6WQ4aOBgAPaeKWpwqqHXiq4g2KeKhhE
12gWBp9sqse3xev1gOFXWVVB5vy2azeGyfJgs/2NLzTFGMVTMVyqDYtkS10S3eMUvaye1WcaghZu
ED9opGob4jZsVJ+Ech4pFgCD2GMPGQeMV0TtqVQViDdLyWFmoQD9UIqNWv5Tn+1XtOLIj4GyJw1a
HEBhcbrmTvtyucfjh8M2v7h8JemeZ13MlF56mZaysalBUn6V0Q50Qmdjox7wOAjkhv2cl+KvE89g
m0i+kWime4LMe9LIccDpqC93e0bzRdZ+8wzbJjH37YECJ3TZqd1Da0TAOUDjdf+Eksn4CR86aDIQ
9voaGESJ0grD08cFWfhzSOw6Shsybl6/suwjayZGVtlAgHEh7afgnwIhouFhNZFIaSSps3vCa5OZ
SLbMHSsPJt5V00qtbUyyFU5WKiKQ5sUl0eK9lOzVN5YkU6y5S56iJKtTMKLclK5drhOuFjpR1erH
2vq48Exw25O9exyNndWHqghCMA+UQ+wwo+aGyG7alVY3/kzB9yRdQZisH+cyMX+l8r4nWiV7yad1
S65PkD6OAysmWxnyopNTOtFEqNQ/ObrUdxul3onlY7NQDmK3lV7HOMcbD+fd7xf27F8wFDDlUv9y
XSqG/vtD0zOSL3ELPXC+IsLeS/1mgUspE8LfDXxuldhYYKGhkZDSbSPvW2wZHsCweCecNzv4R+cQ
WaISAQZ2fKwEeFQGqh9YHHuBrGDdknsTzGYJuPo4d4fuLmGIPBj27HXpqWHv/Ya97ctKvyIAq7LP
pLJDl2yZEe3ELF53Vxu/b2p8XZc5kH2U31dLIhpOnbOEvFmRhd3L7ootTPJNWVMCMTnS+bui9p31
1Ct0383c6MAQDV8EM6JY+/XlfSRRddpxogKzXr75wEPO7qTH5sf7Ml/+P5JC7T+8FP9NETZCRpIQ
3gAG6CnSHPz2gHysG8LwNjBZiyWNIXwbDKV3FSM0/K2vr4vJjWM2/xOpy0mmz5NPOGqdXyoI9/N9
Pl1AJtbrv/7u5b2kQrRCg3xTIAqA9m+e2Ag7MiU7qhOAVCMWI3Xk3XRwT7uab2ZdGZ9qbRcEd4cv
5jjNZnX5poHx+hhEiuyQHHhlTe+uHjd4xiljXjWTg0qBp4gi0JDyV7FikrNq66UEtemxTIcS1EZv
dD+gvvbtjTZqdytqH2F8G84IN6odGZwvrC/f556yAgCrX1R79YgdD9AUyUvtNPQedHB1YKboQ+dy
1WKdpX7U6ruUuNtwnkrHUGCAylcNCSVFF2Cd+4m7TMcZhYNNmdOKD1m2nrft+tc+kNx6rsKvP0Ty
A2O1ZdCPEqZcJBDQlmNAO4s4We7sbbrTjfbgo9FFIyclgX/XeRmgqSAaiE6cdeuBaDWrfurxwfUH
uF3XqfrxXyP6xx1x8D5Y+K/5Zw3IlrY0XlRczCq8X3jY40wZNogMkfKHiJWXN9E2u25nPFZAxgFG
FCT+seKLOYvTehm4Va+HPIg/sDAQiWiadxWddph4U7Xl9GMvbb7vMuxHmNK0rWHNnVVNggM9wqhP
Xo0fh6ML/vpyrPL9W4AH9Vq8RjzW3G5chghLrYDFZ1sKOaqRPWsM9mtoMdFYBqx0wa1UpbSU0gwa
nwBEzTNjzkcps2NgYsI7NLjtDSrCXTWd/4aPpwPZdOLqdKi264pDLIzGOHNj33z8Ih6sEs56b701
03e4RYgb+C8r2VYgvKF46736I3f9x5ppo/y61E2J00gpHrL44RlhlWCcbigDydBk8xdM51AMvv5h
GXpycijGdfJex1WTFm6xUYxNyftnQ4EN/h/E8GKsrkD8jPMGQji0fRP5Ml+KRbFHN7f3PYtwCJGJ
6SVAJl77a3tdpZX2KAfg5tzoiCL9NXHEeDtRNnbkdTXsWWnhYYsJ8ScWkLNXaphu5rptR8c022xZ
H3pboxtCVDvHIZ7gQpCm+6qGJQw+DUU8bNVyMAkG46+OxFyyrQvG4H2EhvQvH5/JdOurd1jWFSk+
vwAzi0pAa1TlAPWMve5mlnkp/C/O4tu2ryt99+h/VbZANYNh/Z0Er9iawy87kVdAo0PWASNrJhgq
sN4Z7S+8KEKGpn0TfcUSogHOEjxpVzCIefxhFZEpZJFIRUbGTEAEZPHc1zTlT0lANlBENeqOXTmv
p25pBI5PySAZH5zE40mUJt7vLT6/Rmly5epTv/kfclp1Jlk6ZNPqGvktjs6TI9n2bv3DKwm/yW2/
z3KR+z7bK9ujHjUzJ7wdbplecvMvNXygBoF0ay9nSPEzqCjNXmucCxZSGv5oTl7UqwzP5XgE1wZN
Fu130i5rwGH+Te2Y+ic1WqygFDZihgrvKMyTIHQmdacA0cZcQ3kchZ/CbtEpF2YLYkRYO2TtuzaP
IBijHJL0ekOoHATKc5ObS+QWxEiv8PolXqrMcBn80npt2iEtodNx+ajBa6vz0eXd//lCYE2wVRHG
tj0bMAld4jZOJ7h0Rjppqu1qEgByiGXNxhK6Xtho4HQVi5Gf9Tilyp6Zu63OI9HPbTGNn3leAW8M
XM/RD4R3zesaIvTAaPqCWlPyXIdBee/rjlhw3rFKbQ1YNxM0GKCXpQH+1L4ybkvY1ZnIfcWpdULY
DdIMaXpkIIdoMKSwVrC/sLgtqLp0k7WHlaN94P0mw7ro8Ly8+7SmkUW/q5BXXB1xs+B8idr8uway
Temzr7qr2oTXz8YlyEPSEP69QOsopDrX4oDGmnk/OVqIZbbphxIJ76bfXHy8oRxVic73WqkzUNmz
9gP4+hFIQdRD1xQW7Kt5o5gIsgemVnvYTGqTgAYMcI4lBJIazwJKRu5A3fwyJgAZgkXcS0AHAnwR
Z+4445xTE9ROwq6oiK29Rn/83SXromDXpXvhBz+YZYlVb/WxSw1scQToyvNXeThm75hhgFwTiDoc
oMeguc2GIINlCRk0BTi/rL+uGrNjjstrAjaOi7zsPxSNuyP/c7XELL1ttgrbFoi8oepeuWTdud5E
40SfGcXZKTt1SL9udJNhClgYON4K+5WdRIbsdeNw58GrZVx3UiNZ2RGGDLZ3pIju9+b2vP5RM7qd
A921S7lBOA6IqXg0tHpOgWPn+Ce59m9SFWscE8GMjq3inoA4bRJx0/66oDghP8fs0SUoivxx42EL
ofa/rcOKM1Objo6M2D88hJkFOYs3g8F+8hyq9Wz9gPM3vs569xb8ir48wv3222jlcepSFA0ZUmOY
f6P3olz4yU6lDMHaWogDsGlcm1hUY6UZrWomNYdRCuXwjym1zyWF1uQ4yHu4ocIoFaRvAqc8z2r3
qhH1hUzXsYhMpjiFZeRApOcPYPmHlW2SUkQLVSZaDo3uzm6UTs+vofKO9Kb34gwoV53lBx2PX0W8
nTLSjPzI5SD8vMtT3wwzPhJTNgI9OLa5eyjMq/V/vDmhTGbguG1mkEBrvymy9sIIP4oUtjeyIkzE
64jT8gQbR1yC5HulXqYJQ90nwXjRKAoZpqfX3zH0CADSoSyOiK45cue/rBz3OUZKZabrxTOXdDFI
R6QAsKvETVYGBrSdQ4HNu3UQ8uwfLZqp1i+IpTP5cbFnpbi7YX4mOIR0QM2xgWMOw3RQz97fwVdT
+k5lvoDRH66HhJ4a/u5UJUD3kD9pUsS1PdQ/IE154Sjtje2qDYNDDmrYFlWfkBwH1fd36iN/GVs8
NSs4B4nqwBtowNTNTl3tlNtRBC/ddPuyUl3yYM5GjyEazOMBe6842n1RxmTBSXx0w7xOYCaxQOMP
GbvpcWNNKKnzbWV2yU5K8VW1ShzOPfyXsf3p3IamM7udiVw+0Xin680DmoM1B7YQaFm/vrRUNAci
CDYAJ8NI44AU+1Z+JahQOj0kM0MbXSAjujScisrw/nreBhvjFTAHSYX03taLCkKbjGPgIvvaWrOg
RmUrTAc3rbPE323rbPkbprTck+ik5ggwRqeigWKHz+3QuZzHlfQtxI2QaHvp9MNGxHloMiL/PIWu
zqRvxHzLApjLVI2txgn4m6cjycttNQR1o7Xrele8x4XALUL+RriK1VQN3qsRVgcDhNFju7IBYYil
z0QniUKZqDc2sBPN+eAegcWzv+T8aEzI3KESCkBAvuguuwuvgYHHunj0DClBtmN6u4pIWFqlKDf+
R3MSCnZKGmc8o7xQ0DXq92TE/BGrH9XJaElInVPlh0XaSk6dwRvSJn5nBlDveAsy6KkhW5eZjuLv
tr/Vk6sPZPmfIM5LAsfVVBJqUqQp8kmGqIHeBCcezWI68+ttJ8GmLYwrA+ViJixT8dyUu76x5/cL
IfR6JV5hbSAj4d9qK7RiaSEcis/F3eJI4FEFcF8TCYXNP0YHlDnvobW05VjsDMqNNX8UxMqML+ym
94K9jwMJYLaYaq7+32ucjf2oX5heZ5Gr1zW6FPpN/owEJYc2+nlWYB4s7Y17mg9RqdCwygQNHTIr
zrRB1RCBjUHGz+BFfwiGndKWyO9Tw4U86ofst1RmSI+F7mqY/ZdWhrkBgrQwxsn/gYYWNnb76QjP
Hvd+GNKtkBQXh0eM47eZLYSTfg5JIM6Lqby0kjUDCW17QmcvSMIpNcE2jtOykCTdg5GvlQJewCHF
/KjzkA9JveswHMEDDBMP/QY3lmCWaUDPf1zpagEgv6Db7w7Ahii3kge03eQeIPhSNzTJZfpGd5XT
tremLSctQCnsBJfB+YzC1OhhIfj06BPJcMLo+7E2BL+mTb7Peaxja9yFF9fC09yL1oV/8tHqyZ6W
yJQEhQAEVHorcwC8stqlKkT+E0o9Nz3Op9VpNG5UOu6tnP1KFVALVSKXnUhHk8sOfFhNBv2swG/0
3WuSOvFiZCfDm4600gSG4w6baxxHlh51tE2jxUBPaANHsys07A1CdW7RlSrqiqYgdXwxKjcYDzin
b7SiDPartS5AzxpTuUDgvp7CSnKUOh0wLeyuJS7PcLSqCwFgt6tSO8l0RuDq8oODjUEJjoEAD16D
FBNby5eBotsT7A12kRUoAjZW7QqiOEAZtXTxzLdfyFKNHARPfVP6gW7NB8sujAMhVCBZ1yickroH
eGRn5/yXyC1EUauDrgWNVHdcWHE3u8sjIyWbdkpio6C1TvW5DxNrE/3t1SHPs8S+sHxi7rLg43T1
Gttx+6uVFqRWFFUdx+w7AZukbT0tG0OCWHxp4OZGvR4NvWNAtz9Nl0RFdiwIbR9/M9Jqrmc6olhr
5/OhZCX6Kb6aifPFEIcowGzQTuD1eScKvtcwQ4dDVd0FKvt33DRrzpkSsTFEL8qAj9suQCb7qX54
pD1FlSRcZlalpnF2oG3auA/fqGKCyjM2FCk0o9JdlpNhtcuGQkKQ9DPTF7tqNo3F296HP1dydEkA
/+gY4fE3Qmk8/Ebf97uyCoEUw/SQWo8b9+PsmwV//DzIvfRhYgq3e5KNhrlLSZaJC6ZGmm5XFH4x
HsfWPfBIlXJJNyt0wF0ii/cWUWUQGJ99/GcXrb+QGLStc9tRlISrz08++CZp9ETH8ELTD8La8ywF
yPOv2etQa+/yxQuL/B9NPmLMVjqoaFuEtSbM2kcH4kFvFpGHYB9oUzkYiAbOvPar4v9pxKETvkBV
JFgM+zXDAMy7kM+jmlC1oe4OsZcO04fXJF+pjToKt74IHsj+G1JEMNvZoZrMjR60tjb79r3FqG9K
HDupU39Efb5z7ZOY37f5kVGeZu+VqUkZe2pcSMcipws5+f/Eke24GOWo+nPrb4DPfyDtWk1Pgr4h
mrA/g3HBrYL9WdHGSdPzUGOq53cMvK7oOIFb0povmETVctRsm5QZo+BamRLY+hnew0Z34hDAv2cN
kl/pPGcg1vaSPQC9E7PzUw5hW3nX/Tj9Ag+Gp9irt69Qbmim9G2PLkkncTSi1Yo5kHumxs90lr/W
rpDUn8NTnVPBPI3+ZM0IU8Ze8GW5mGK2iFFaJA6pctGH4TFA6U4hwz5Pe18wvsJbmXBEs3VbEzkM
hWSgsxeM5TvwWiKY3FFkxojzY2GaJR8XYZ+/emb9SkaSVGNKCDk6o/5eGboqR+KUJOxY710fZeD1
bFe99rwlMbzuE8TqlqhgJfJEAtAEWWs90rOqOPNX+sr+/0be22kXKmGkz5JibVUmo9iwhmN6jEd8
sNZblZrLb6Q7XsKBk7HyboFYuT/nzE+D+JO7Wg/qdW8A+26bPQssHfBS0FGhx7ukmOkN2wJwGXJk
LhIvfTl67kEnrYJrdLBTsFXB5ggKxjd0jOxGU/vrlqTglRyEpuQm5Ksr7pNsVMixkJ/UHFS0DLcZ
KAk4YHMcirQSt58aix+QQenjBTTpVFuy6ZTBzz325Qa+R9jdrBo7mstKBSg8+MIrzF7x/hghIloH
MLzc8LOynWQ3xzvVE+SWZobtYg7jzjDcj/3OdFUwu0LGauhscdgQZpLS34H7shy7u/NV3kBka1wp
l9OBy2OOANBYdslL7K0DYo7c8PZ+MQyDN+ErtFJ5T/HygQJkhoEAn1q5RYoj994B5t5GxEPTbRKK
96fF9f+nDufg2is48Tn3i+wJd0iQXv6Oi5O5F8v196knSIbRh2fvkFysKlXZXif66LXa2Gv1r+z4
Rc1yYwLrwlnBSq7Lq2e6n+xea8RSCYDSc+wL5vyG6ll0kA6HfZNlSft7QdcCSqBIosEuUF6wmovs
ztR0YvzLgLBASPWqZOyXP7LKWVYY2vZTW5fqCAqQ8gFYg2XT62Y5S5VnIOHYjqUTuuI9kYnxEam6
p7Z3H4uhRpfIOX30706GO9v/Rn50XmGp90vAsvA0bxvhZxmG9SXwZCNPRKx19Km3f1pNmU+2sUTz
NP14BKTAHpOMcbpLu8HBkI1VXYpDWAdZvP+6VsD/qAeUsTAB37SXAE5CrtLpvB9Ljz1J5lepM4/w
HP0EKZJrZBY/k+gwVF0Sw7yyUn9Wmb3KP2ODz2p2jR44LeUjQx5sepkVOLSmGsQS1kq+qcIxcRil
6MAYLsUK0ZZorSRKA/c09G6l832Zr26WNxCD5HGwAvDJb2+zRUlDpVA0vglUtt/rbUW+G1SH8Mdk
EnJWID6nFvJsunVK4garGBYd2xgbP9DsDaduJ/If6E4eQtIUom14wxry9MgTpu03Pe1HvX1Dy0uZ
jKKAwmYqNw3nypvXRagmEsrOqOqC8CPPu5vYjFjnPiEflLdEoe96dZHfZfR2ZpTeX0M1JKdIZ5OC
Fmzlj+KsmnvDplFYEPjHyozSejtQvxSzmaToY3S143yHygRus6EMxiVXas443SKq4EE4wMgibMKi
+flhKUZADZnMzlUM/khlbbpmY+x5nwe+fDzbu+gG1GD1yOOjnNwWcoUis+5wvJRkvLZwoYLm6V+O
CX8g5rtU6XVWD4jDnKuiuJVZU9wyo6QAFo91Ym8gK2kPTgnDVIaSzKmZWVQvypfYJtOP3JjPJYIG
uGj/pFGgals8QzK5GOxzzXs8ve2QSAWzfZR4EYimU8hbLiVi8eD1fH7s83pbH5YI0ETA+MLEkTrz
icLtOkiR7Y5fwunNGdROIVwggahSQaQIapwlK6BuFNtDGtkaJfwiuN+8y1biuC+xoZUBFT2rvopU
FScwKmGFnBycstcjIRK/CTyjfJIpof7NNz512J3iyaUYAXU+oujJ1uI4OsWDjWhObo7Ui+tRNgM5
NSXA8V1EXFR1ukk0OZTkC8J5i7uuMsl3PcpaAuArFTE0IJlge24KLrldnfKPbgaLRUW2R4wVG3KJ
WLFqoIDZ94fqSgSOIOqiQcenJ2AnSsQS0/MXcE+SV44hgq2y6I84G0daExU/dmRwYOAM21XVs8y1
BxUfn2BLQOwUvbzt5gbF0h4n/A3/5oesZcPGDidN+FGWdr9yLBKa75tKAbZ7O8HaSA6a4utQsZnr
u6p2+8qjLXIP0GFeKuNZOZ64s7PjqxbBKAQZsVoZD5uA5PaG9SreRfL6u0jHW6Z03+eR4VMuf+VK
aeICFTo2zbG5Wi70xn4OZPCGKL9owzhAMMuiAQXJtxH3N6r1FvPOzMr2jaRk1KV3MfQCzaH7JASU
HagxWY43AIYMBUiju8QX8oQpl2hAVxJQrXTaQFgjkgTQs+sfOAl0ilSxpxaGSqZ5tW9c9FA6CFti
vB17nJyDzZe5sFx0p6QQFPmBP9d/dkNIuMM9yUjJOKplZZ+UsKvq5yFX732GTFzmbZU/WzFIeCO4
PVpiEyykE3XARe+/+4ZoSYmed+ox2xEdYmePUoLMyLPxcwz7z5gnMosyKdDEsrsfG4iaqmZEKOPQ
EcPDz1oz+KoPnEkB5qNRaA0wo+qrEqWy5UtbI167I6VQ+nFqPCJcniS7fzSFcbuaXJKTxqREspCl
3jWRdglsve8tdzNE29mgGF2kGallC0nEvKFfFBor+kewppCnlowWOt0YWCohNo4pPw95PejQqKn+
lDzIt8ubDMohJexUnBJH6unH6MzJPDQTo3jykBwaO6GCnU8RQXL4B04EWSay1d305hiByDb/4/+W
nQJWm9q+srIuVn2MVh4LPstZnCpsUpDuJK5gSY+5GtzrUhqpHSu7ElcCOl6bzS3Hsut9V3KEJ/xu
Riz7UW9oaj9+BfnhCx07a5w3yvDa/R4yGM4cIw3eufDwsE6M0J5kedbv9PLi1wXT/5sVmCyGepOT
6pxQBkxk7sD/wkTqIiQyxhg09tta9D8v9/ZwzrosobJqrBTCBnhy4aITbGhLeAseAF87D02uzmpQ
QfY4iYZByAtlM2WoS/grWyUOJo3yNzfMdkfH+k9XTMnjLJDbwBJzbpWmztEb+kI5BhOFhXUs5FPj
IUVshTqeFjU10UhBGgdP10V0dw4lSghZJPnID85jinD5FZ8LLQm6vY2HKYRuRMwEmKfNn0dzmuoQ
NfehQiXbhPUO7MsgjQO+nMd/nGeWdV43q2epylB3GgLzXigK9j8Ii+g/vL6yFwf+QdDhcyG8WrFK
lDQmMajSRbAIGd8xxy4m9IakFKKU+QyCDzT8MM3Xe7XFD1jbEZy5sktPlw5O6ZveNR1K+xEdfWFo
ym3gZHbESBCi5J/NSsU5wjid8qF62P0/sJa3C/e2BhvfvjrZG7ue7vayEpZvM/1XI4PWXmTTqOT9
/PAOyj9GNWMmzMxhM0BB87BIi8pv+ylZ1A9IeQg1OAdM2m2Znno7UichoSC3Dmb0qqH2MPQMWQAN
t+e6CZreZw3yzNoxv2jAND3HWkBzi+/1PaspAZ5ZHwyK4ltj59UUB9RG/zgzQWx52v4PNchnN1VY
vHxp8bsXwVSToCgYRo6lxw7H27oqEeeldGsrye85EsQaz79VTulvgSiNrAb8b50vKG9lUPSEF2CO
qhB27x1l0NVeyY1ZbIMf0gP/CHXaXAuAN2JY12APYy7P4x5NxSBMtPpr4DJcxFadMK/jraGNAGaa
7X4G7ByjFSV08YVNJ3gcJe2ypLUR3NBQULZh4EPv1uejb/giaTOnvmedh0bjvXxaQ7ljPyZHG5XR
Sqc7uQJArDokiqZIhO9/WwcdiPLYqT/tZMKx1Izau79z0u4TtuYx9ICqO2+Nut88AjOanPhh8Mds
xir8CorakTgzMoJ3WvuywvGHQzMfwvTe6VZSyZt4NrAxLVmPZJs4JdZZ5mi8FwTd+PEDooynQBvH
exQzKRasWE1fQOOBC2c6tC4Zg+EhU2d1TUmTALPtkXqRgvZbR4XdtvLmXEAGrkwUqWAltof9jk+a
/unALFZ33HWgSJrwXuvWjzlZgkNx2OwiVsSc8RwVAx+8h06ANiI8yZ3ho4RPXwUf2RK0UZUEN33E
XLRQ1F2AfrJN9+I1ouyFRDzK5J8p7/Nj4ip57MOLPhd9fgLGvcsE3JcVUkQ7c5OGyGCi96g/67Cz
PdH7eoeb6XzkmNusMXG/SBlC1mIn0GeA//+8DW/y8sKYSxPG/QwnEaCIiNcxPgKPpbIb1W6sLtVq
5T66srez6QQOubaWOFQ0HPE+9YystWP53NfLyZDW9MAwCGxpnjZBbWwEUWWi2aR/DcnX+E98OMA3
mEP7dxXoM59xyqhVToBF7dLI2spTGnK4uCs4hroLalaeRCZkDQpnvRNLOAu+Ovkub+VF9Avl4a4F
6K2Cj0ghMmAA8u0L8fiDTTvoPb9Ugj1H1D6bWMqgTxpuIwrZmB29RPuK6isZA7Z1TkTtDCYOXfv3
ipw14XkUCRM7yQn6Il778OIC5dq4j2m0AfFvpJKNQBYExYjieNAZl99MIvTR/7e0yt0vq6JE+2R0
s7ipFXG0aX21OvYVnYGYIS+T6mF3gu5RvRAW9e0WZvhUjgN7moAul+TGQmcqpHIoKu28ORk1gCr7
TDargxWgpZ3oB74FYT+OL3PnkyCU4CW9U+R85/BrfPXjfhGG7FjqGQJMLUoLg7UxjXc7LcCFndt6
lIPqJDKlhkmX3gn8ZFzB3vUUUXfF77K0bX2abDcssnsbnB+6FLcelX2ZHoAWjtGkvAKiBSg+HAW2
pg5UAvznUXtNC96bSrv+sjnBkC0rdSDZdqh84mLG4HlsZzHrs5NXZxk1nCa65oKxlYmEYRHTLXDi
pj04n0/wmQEqunVn4PV9E0xl5DG/rZetVpsrHo2EvkHST7Inl8YmbDiYwy0Ts92F4h0m4Rx+SeqZ
jP+gxq8GB3S86CAYQW1U8m9wOWjquBX71z5pU417vCa4U0Mo4UT8kz1Pk19ch5YJn3T6CioshAHv
dl0ePaUw4cs4wwywsFjmXFpMYbdJE6CRZHNk0KjxWt+22tuDeEavzjcfobHPNwWdct+V/BzcBBeH
GauOZHKUNB9mqkfa6gY/EyB0diC9HbxBEWCLlBwmbPUV70Hq3R8FJ87MBkO5gG4eNvDqTiJw3i16
t23oLjIb7m7jV7Ww1WmJQdGw2X0trRilfe7hHEEq//K7UBzT+CUi72uWtVw6leGraneVbllB9v0x
gouyadEzU0plV1ZtEyhqhrYRj4wiUei6RWXgx2Ae7wye+eTpINY/ZcJwkeR02GA4ngh4pPYqaMe4
7wFb6LU0RpU8nK07MJqotdB763YcLBr5+V0Weosu5Ru4yQ1Se40dRYOtnYDuHqql0UQzTe5hsXRE
7odIlvHQLmVIE6/FzfP0OTE5MK68FjiII0BwhO9hpaR32+A5ucn5eBaSbIiPWNSARaUSFojiuy4n
5GwG41InK9FJz2hAX0RF/w4x89/SWe2z/1Dw+0NhOHNGdTJbMKu1L8iCbJz8gPN1ubpiQgunQYDr
/GG55dgd4TE5v+lACxjH+d1GtxC88YfBVNMX2thhZgqJRGAWdpOQFvR/6sf2ZMsUVfN/PmMHIZkZ
Sf7apYm2PfwYPuKVJmVqLeZd7kr1hfGtcXgd0Bg1VoP44JGdqkI+MDBmIr5NmfQUScRT2lDg5AtV
MdJpKrQsMNxkdENfnz0km0jE/BQBB9R1rEH5LXFSDOQBonKDYRegH9539pgNcP5fbwExLhsaP6iz
MXgnrJungta0rbkcusPmV5gPMZTvKXkiS2qt8/uPcGB3UYCIwbxPewl4Gz5r95ZolkoW+VbU3FIY
0B9pJerbC4tFlWZApkeocTNBERKgHciBONmCcOY54t8p6M7EYr+SS018wnMwYX9FEtIoUBXvxWd2
ucc7f8RkCx5lthYiNHXDRhRYvpI+ElhksbutaiSQZcOG+kDQZKfnKmzcZmX2GCniYBj2kK6FX7VU
hBBW5eAFAulGEEn1Jvo4fDGRfxoSk0qTIpQj7eynRNyBh52dsi6IubWdgIPoN/VvQ06tmKza608t
yGZMiclf+RJoTtDtYNAiZtaIaYv+Jr2hbNKXwljDzno/zcG4jbCV4luYH3PH1faco3G4hIxzdiEc
FwD8uIBAdGZ8GwVJr+07bk6Ai+0dZBETKlsL9HUdDRvgrsOA6YY8TI2UmkqKV9rAzOwTNfzm2Gqs
ZpiYBDaQ8XFL/EwlMLM5ffteDPj0GtaNmNFWWK0vbwAHfSBiuy0XvNAiqra/7K7xkC+Lx1qgU3pt
LbXowjL6R9TnIJALKeGyycYSFMvJzEr4YftRgSrnFIKfgoLaHAPbAE2Wt93XeT07H0lOb43xE35p
PvB2yRujQ+8BFlyTS504CQDrzE/5gwgBKxIfoHlw4k0/8vv+phGXsLKbd5WgAeeWFXmAz+oliVPZ
TxH6nQwyHKlANLgVQQVEqbsFURd3unJFLxPnMdTFhcMiBBbmxT2ctVSHCOxmaKVxP47MEZKe4sId
4TBMxEXIEKTyMGmml1ni0A954abuw1ciegh3/wDqM2swlK73RslIX7QKfxCngmTk9xixovfaYUpj
sJbWrVIci7bXfwDMILTyNbAap9rJ4cUuu9uPSeLG2s8XJ0RnIlhNqkvmx/bD/ACDUMPQynLUYrlh
skndwK6mUgFpWg/zBb9uEZnsORBK46phpIHAfTlvBFWL2ZUMT/YtFFNesCQDJ01Doil9CAlYEMPl
UapMWbyhXgBwqn/3kP1XBJ7a2Der67NeIvNCbwEVIG0cwJlxf+FsEj66Of2SJ1u6eDTtfPmrc5xS
gby02h3IZwztINfag0J4x7+o619WAi5l6IswxjzYvV5oGepySnQ+IEmwP5oisRm96P/DPrYq0tRE
vp6h3zojE0JnTs0E944nLQ/tye01WBcJkDsOf25ei43oqVctuBipy8pUPuFSjGpWET5Oh8J9eP7Z
DIJKX+uqsHhIReETnI0/zjCQh/f//oe+1T5DKTnN4550e8qKugXp+bkZcAFV990u3aeoIb4Rkas4
odPuAFUfU6XHXZF/hnUJA5f9VOONXQn5lSsyBh8zRtRDjJjDZM5NGxAamOibckEOv6O/Mqn33QaC
YyHK+DVnCTxFB7NJKW6/ug1ovpDQ2p0XUY81o74LHYV4DtO0/omxKlH9VMMVoyjL9MgzldeHEPr/
TSte/GUeh0btyFjuRUF8H3xOO/K86qNerLQ3f9rLniAaF2r/JbGAJye1yRCYoo5r0Qgmi5OxFiYH
bbFB/s/uW12SEqKaugtIYbeEPLQHFn4Y0v+mc2JZSV2AS0w2DZmoY8o3uafwY37L0Zi1GPB4jkZE
1Uh0xDlRh3x8QirAl2moGGAyqEiwAfV57D7UGpzzOoa4HBcVAqxbIEFVA+V7Uko8n4tqd8g9nODx
bEe+qRtJ+IJUSe86xLXrvCNpSRKQOwmsOfTC+LbWUzaPZNXFATWTfesFv2iXfL01mUptX8+bLpqT
xlKRB3dofANZYiad8Lb8ha9RNEYzFj89GS0eMfnGBQj+lc4zO3XQRutLEGoq4XqaqglhYZdhjBzd
ID71gsSOLF/njBc9tckn2J6Egk52v1aYDOhvJHayJeBeE3Upv32AN/Xbz2WzlH+127J41wSl2keK
EuvTZACB2PWQiQL84uqK3h1F6Z0kUJn+262AXt3d+f0TYsQg96HickdwnviFMMw+GbwpnfVDsTkf
qOTTAW1httH4iCe9iVU75xkVKnSzQ41Ag+bxRkR8WvjK4cSFMXTlI731ge0OMpmGKeTxSWeISJiv
LZhShr8m9cIFbUHPjkVHl3e7bHw/pf5iC8iZiertaVc4T88cjs12XrO9iRbZzWnMT6S3bHB9nzIa
C8WiixubCL4vtyLlyEhS1e/6JqgvkNNhh6Hprex5YW/lndBI25eD1mOsA0k6jh+GbYHLB43TbKBG
4sSIpqAg8BdkjZmI2aVnHBhjT03/bdcnbnUh7BgImElxa5THj3/BMM/XRMHHWFKqtbOAdOiXpjLu
CjEdv0YJfTgo4exIE81cL4xJ+Y3KenDNg4i6lHzuGYhDDsnYFeF4IQTMDvhaivHIJBEqYCd719lt
d9jpsu66hZDNDStQ7QABQI1SNg6aVJurJtNXgtXAKZ0unFucNwriVxkL8ZlBaw8BSQW2DXXSnzCa
8GS2ip8vBtEqKUyJlokMBVNIKdlnHG/wekVvPQpaVOtE0/Umet1/UTD71Ylq4gWcEUrUQt1t4RxN
/iAW631aLVDLfQyIDUcMcisfBjhe9nMqGFhyi9c4vdjM1qGY01dOjQJTrNhZoMPrzag3DfLXiufB
sNVTxWHO9yUw8EObbG1iXT/nXIQbzGH5Bzd22tAXmJxtyKHdpTGJH92nbwOppRVl9iKj4mBCud8W
PRDNWbztaRSB1dmRAFKt8wJEGbK8KMApq06evHR42Tqs5TgFMDMHmz2abZudlpVZ0svBpvqNWx5L
NNzjDqmyisosKjy2Emgh0RHzhU9zSxS/nc9q/j6n6f9cobVQJns24b+kd9ZBT+6g7K0KcKTIpMyL
+3ho8ELKK3bz/n8Sv9Wpz3t0lTPIbG+ipFqDjn2HbQaD6R/picKLVOM8kEGWHsy29BDwe3mO7zwD
VdB0FAQu4bPMwyBKNEjIVOk//3lTTrtP5f1CYeDOrX0JiHrfITlI1aYZ5WFd/uRCs4nZDXsUakWb
2N2SEVTZiGPahUkjB5qPFwSlQJXPfuUIaomICbZZFyeJkiLo/jac9ngjzTsJasKqYuCpgxv1xyki
+0sBWSVHdqjyR8e256zr6A/KzUWUxQgFNgHBwX2H5NqcPHihs33aSpYonjrzzTtTItyHSJO80gCe
1CovIG5F/thxduRE5UETdxFiZEZS/rNPg1bt6BPhyrCqAGzbDKlMHVDRfHzrKCz+XKLaBcVDNA3E
XtHygaZ8aN++DVCiTwrpv3Ovh7/M1oBic/xe50+hVKALr8LJQheWxP1d3KxP+afmU6f1Tr4ZVq9K
sH0LQQ63brB9C4mdBP09dRSyS34/KsYoAP12Syf8mS6sE2Y2ZVEWYrHy7XBRa8r0ZO9ypgHUKAYN
5fPqtlesziG3L0R8/NZjJrYbwOdcvIiwEczJ7/PTpPt0wDbKlOpf/rFrOhacn24dvsIwgeylweaS
aiRFXmyQpMgs9AMq62Xl5FcY40CeTF7srFOHUA+qGRZqamNqugGOiem8WHDslIVyWyopFelvVhvd
N+gMDWWFMcvFn3fSQJeqhZVJGA5g5mumwl/FNnqsiE6UC028YDLVyJkKxByNUZ78s783COGJlqPb
L21+h/F9+vVCTACKVrjV2+lcy2T7afwKBNnlxsGQ9khWPDTfNXNfP1jlhVm/9uQKA8e46eMgPb7N
yDyWhJwSamR7mMGyTqL+QFwB9gDSlv9VE79rM3/vRsi6UtNOFlHYr/VjbPNvc0FmVt2K3P51Zewf
aePj96mv1t1xuM5tLRt/H3qVMAVjoojfu/Vw5FTd8nykbMG+iDBltjlJnMLyMCJC4hDGKJi2qV4N
GBrP8EMJaY/2nsMONx5VXsCIKAWeetRo479oxfZzfOkep0k4hKgsy+mCfHAtyHgYI21nE0goxdtY
m9eSmVkMi77yiL5TOyejABPGYR1QXUkfx71VXQZHe83qrWchgawF4POFSWABFmaEIgFO+FMbCmk4
OtqFrIRxfQyPOGWqoacXiaUlwTFs4IgJYXCoOqoNkHUaHQuV4jgYxb86yB1sXnHOBqg3JLBIXzvF
ps+iOwoutU5TtVpZmCOBQKAVtcWvhiAHHJ9qJkACCBvtOw3ecAOvin92tr318/DZKEV33os1bZB9
z0Xf9hq8eP66/tMXfdel3iV+T0EJpCLC8VbC6vl9SLSTNSTzjltstGy4yuXbICdPOUsmzvCTKlth
supZnPcZqB9KCLDR4NwoOa1shBstHJA9FZu8lAKO/e3bdjv7oXI7Da7r9A0+R7hYC0F83ONqJo9g
kG/iyPo1HQIcsXDCbdCsy5bIxYO4bDFV/JwTYfuVH+seCn9+sLUPwGOPAy1whnqINb2u2QRdFlws
sXM2zWhfOMKAb67xER5Ee+hWAKfN+PxffNCxyVcR4vpel7WvcO2mlKobM3fGYvnyQbT7KGbRw45H
8ugSBD01kVjgDoSBkEPD/VZdApNgEB+/AmfzIRxklSgdTvY1SpBesiWPhbAyo6Rcrif42Iz1vuor
W1yTH/f0GFzbCHoKujzVGY9TtZF1NUaj0fl5+fH1NR4NaYjRAvZ5QYQlOn2zwWgy5zsZrbv3EgTK
DbvCOXSTF+ftBwfhIBGjA9QWbwHw9T48cCqKkKjaXYX/IPiLqXkpy4gWW+I8kTXAgBG02PL8wPR2
sSbgXn3s0/5pHITdoTDkaDztOXRB/rJRSwRLgQQxUdwwuOho6n9z8ppbaFq4UrVQmO+lnFrZG2xS
CWK2g2Rn/1D90N30+bM9w9yW7hXAnoQ0P7nKesE/fVA99VAMNCQGVYxmzz8KFkX32ovfhOIe5KFh
hfR1A67NndP1mV7kdW/aX5rjJPOMwpTWfpEhe3BmNnCTHCLJYq9XpaEfFwKifrrbXt/iRa1fIpDb
X9v+DCRqVVRwLw3FhsjalWiSA6A4ry7Vy2p0/lH1n1fy9m04P3mxRTlo34FAlQyWdAZnHW4mZIkp
j6KzvFrkZJ1Q5QnzLuL8OMFBacrcBRfUtUEMqmiZr3ghe6bMMjNa1XfNUJfyp9jqoQOnP0nOQrrE
Kho3i92c9A27HewyoeFEiPXvJnyCvBPTETcD1O7fK+cF7GpSzBgfer1TupJLIJIXjqStpKZKhTlF
d615qX2TYP1npFCgrNi5Lks7NewNkFajJIIll8ItpRV21NB9H4LhEnXZnBr1hNlv6tpUc6y4lDhv
1T6MEMdPKSSK7y+dgg9wMrNB/HfaEAEnotYY1O3xOx8r5wP/e/EtNLg7rgD0Vqul6dzHCAP5j7lx
Bi6urYXyHa1rBHu/wBKQo9WBnFIlUCl5TKcSrYNGgvsZqwGMj3i4DcKeE663QFxzQhr22r82rlpn
76HUTrkTZMNzJIVde4OpZ5f3LPqLc5wPQK00SkjH82hSUz1giuXmlJmCH70NcB0SfJjD450P8V86
pKHd0YrMuieNUA5qr0CVJIYOXLe/6imLIC3eeDVKOeM25qJwAjvYoaN1yox0HiJcYVuZVs4aAbud
3XvzArJziN0OQ4FmWo0rwe8QNh3geJM+N4KXVIrRGEO25qp8FifZsMa8GF5fsGdPp/xSwKdNGBYF
5HkQs88L8/X1WQN0bW5FCgGqaCYfT3Pb0/4m0qnOfh12LZ7leN65Xnaj54zjg4/UYoKCO09Fj3ti
kE+zzN/JiqaUi/ygM1YIXdHyKD0Mqv0QC9r97Jejl7iiT5WmAsQHhgNgFQqbVuSBm8yjfMIVUi9B
2Yp59qK5ARmdz2e8mVXRCmY5Hv2fcFngXWJOKD+Ezz3IrDT7AfL3vsotviI5dNu4abzy3EXrIyvo
cYXs3mryVngExSgpVYiqes7bfUz1leQK2rtY1OBqcn7nAzZC4ugJXDIuAJ66zvL6bvf2Nv27etua
MrkEQsG/RcBlWNcw/h6UNONuLsu87TOBT9exfQFU0AtOv37MhIfNZErsmvDLhowKgSaG4RdH7sUl
v1KZLftlbRIfeT124ZjtxqPJVxDnN0mHvCIEDX/WVpoQgQlguQSZll/NwqCNU9GDogp8+vZwMLhW
RqqdP0TsOiizN8aTWr+HEG3Bcngxs81TBs3Uvm51RPLfTafRJRYjxSa8luC2gDLnQFzGZvfbJEKa
3mWDKJ3hZRbsVkom/icS6QHiEo+Ke7rXqZJ7vy8QGoQ0SW/XbhgcEevnLdm6wfOs2ib+vCJMiFyF
bs3AJHCIZPZHt9GaJ4pbBNkaZZWhWcjF6Wj+NKct+1jmeAChiG/H2rFxy+/NG99dJp9XiDsaB0IU
4SZwpExRXD5IyJZTawq6Az3AUIMh/IeqDoeFEIyef44sYUN25d+ipGvG9PNG1NdV/x6US1sZtL37
b5wGH4/DBLv9bMpjFXfptTZ4xTNLR2r8wk4yk37vSf9JGoFQesTTEl4cqWd0zvDYGoYYIcc8WF0H
FfU96DUPwiV1jwGqRtkVbXaJL7YpejGVwRHaMjMjjw2KKJw3QyGu7E6Mip8sQQgkJIdm+agtLfDB
vkDazMjag8zgkjduNObE6eFv0+JIiaaeIhSwJ9J6SOAMVGeoXYTqt4GH17aS6rnOSu0tmpHVZa6/
dUAwXaUtgiGTOtUduSj1K1cpQoDUl717qyTtwTMyKgNGmG+ApNa5mPZEUNvPqFF1CG3vmapxDH28
CsNfh4p8MYEke9yVS1jq7fKzYoi7JklvUYo6zpMKo9kVPJwkkyC1fLo1CsVW0pnfTr5GCutATOwj
62pbxUq2a8HiSX0McYJodRFXyld+N/6m4Eml4T7sxWAe9osHpnzsTAFYGq3d7rTVaqIgWym7rbG7
qwlOBx5quGcEnfCM7AWVPHUJgfKLwF1MweqG/l6ZPchXw4W0VwMgsujXj6TGiuWMEBKn5SXmDtiP
zQ5mq+2uJyO24CnzDcuWjhpkKnvdbQDIWnv1DT+r0WADgXGwEzfu263nqd4r6n/S/RbPc804TlAS
wv7clx1jv+BeRsKe57yBCIQEXpZUz/XMRxCgYuG5opQyiUaPBu8Oj/XKluuukOkcNRETLrzSwPd/
wS8wiAC3Di44DprgAlFNL98iiUpNfl5oKXMxFbvCPXJCg6ebEaMv62LG6AGRxOxoLpfBJb3ZPtNP
86GI47F+eTeuYyoJ2tvxDyq8yg1YSuaC0W4eJO2YmN8kp6YC+TH2trLCoi6/un+32yY3k7PWTHxF
6Vsbmxy6PuIMkSI+BMnRu4cvOQkz94yGB5yDMAzoaoI2jAScxHJe7o36KExKfcfyNidWO12q5zBS
Yh8RBjk+o9rsUpWkfixD+9MwgpRZXxMPSqpJkA83aaWibKREcnqBBDtc+nTzLdTVrNdPBsVGxYzt
wqgwlBJ+GusK5/7Fo8wSACE/tx1VuHkdsk9tcK3PPV5S0a7vrSBBh4aCH7BoHuF4m4OEoARPVPRq
prLkk8W0z8eJAPi9HmBT/SZ4kRPP6GfUb0NDJJrIyJr2IwmVKXqkWQYnoLKD2A6xnEK/qCBgW5lk
j9XjFVXO83eDNI31DtZ6RdTvPN6H9P513iBcVXM32MgLz5H8rQtKfmxx83trtRNnX8r2E9qmJESU
ixSZTVojSMN4CPWgvuR//irmGKArrUA+VHn5kU+qbp9Ypu20rtYp83Ps0mEs5c0+GVlrQqhy8p/A
o2oiWyXhvDNiIqW2LZCHsmVxh4yOngd3nTbsk1CPfPEvjplL+wqorQjzfszr5rpMw5PmJfMssJHL
Fx1GLzbhqwBwnSXvGqe/FjPj9GuMxzAwqJWJmBxR3TaeBX8In1iL7pZsgilz98oIzCnxigK9397W
780Gq2JehnmAHBS8DwnNhusQpOZUXCAmAS+84319JhueQouCofZC0s8lw0HA7lFBCXWY647kcLBF
F4nGrcIuJd4t1lXGIvwLsrPSuvF6rZqP3P1hi0HjkrFLi9+ETf4GMYlwpGyZu32JoXNbLBUPm/g4
LVoabvJs9RdbQrptqHYQU1DnviY64CF86M8xRqgcUqmU4QbpbO1lOBwSI5fLtUNGbqqZSrUkxBf8
vBvDkvZoxy5Ti69LOqnMlSZNcI6Sz9PUdziFKklow63iOrF6yS5ibU9+MK09QJlsIDCPw6j6b5Vg
ITwcv8/dALJvEPn8AJIQPIpDZvWwGO8dEGRYYmTvLuyfpkszUEpupEx6xqpR/HjcM/QvFzpgQy4t
ixG/85J9S9HkGI0e1g6Yu66xCVFtckO77qQKdzMu6aQirsAk9WJ0eOSO18gUaXij7ns3d2CFG5RV
M5cnRNRPAR/aAOA87W8UMujyUuHbVOzx7FzaIJw4Y8NlW1JlCqmWRTC4JfJZj7b9KbEjVXd3f3B7
rF5VbTSCniNH2R7/FAgDUTwl7gUtlswADC3hyWK6fJnL2QVqeibP1P17/c3JyOgIrZEGu1g0dkkj
AP2yHHpULxAWCoaVIvCrc9IvgAvZXVpwd5XWxO1nG7QED3iYjkuLektVDFOk4Yqo7H8ek52SUzZd
NFg5r/1lt6zMLkt4AKKSClWC7lSzYCVSiWSCfp0ErAYmKZIPMwL6Qcpu7lNfoFVlJKJKj6i/NXnA
ptkUh/saCcsxyQNGHpquPgoPNnzh/BkHhZDisV8xp99LpnhvM3mI7NGk5JU3Sw54UK0C1xwyoKGY
R7eqq+yayznU0sEW/xBaYSH33AQH2djtdoHDiEaIgvDMm5RtkriUe2Imvm+tHmgZN4bJ8fLk4vK3
diGtCZSDm8tCYU5g+cJjBsVe2f2ky7K/yXT7Zl/2dd/04I8fl55FlncTPyZJhGBZATGg+kPVKpeP
dZ4mqkDo5MsQCzI9gpZNL6XXKHDGvhmfJtnDmJczDlxkXoUKJE5Ks/XqJ+97UMT3qGTv/W356yiO
GietpJRnzI0NAGYacFLKnadPdjmt2Ctin2RatvCS7bltf0woN1Axc4jwjXzhXcOx7vW9R4Sd+5n7
EfDrOjqbVlFFNjwRq3qM4GINWSjyV5wXmCxJyew0mVXFnm1aLxURDd+5ACRuvyjQsSbQYawAIn9o
Z+aENyj5mRwullnzqdUfIaK/GnXA0hw/tzYUQ1QNo/eEjxj69EA686Psy3PyakwWJUhInxtZyxrz
7jPSMNP4FgEiAvChafqu05ykvYNiZq5nEf5xSt7msszz02AqVbXO6EyQG+LALEML8nN8Z+BvMwUC
XM9pSW2EcM7ZwNe1uVmyznamr5ZheWaiDrpISNtcR5EMWaxG+egpg0CVDAwDELA+ct3kDh17uFy7
7b3de/O3RyhCjhiIGOl4jZjjt99jCWZnPsV0ADfsl5Tbm5eAhEQ1GOw7TcAetX16smS1a7+3fEP2
0JfDH8wLEhPYocyNZ7hP7HygGHDofajjEc7hNNLEVKw9erWhbTzTNtvDX9znOqYx2nLZ1zdWZaTO
PYnN0SUlXaPaTdzuCJmaED2SgIIxCN6VUtVKdjo2ARBNZZjXxGxMWRY11o71gAdNOzX4lpgaj2V2
rj7WpvhlwRfI65+NgJgUKFtj3eorYJCdqY5txX0F5LtaTZbe6Z/6ec5kBjoONNWBsjHxa2bzoq0R
DUS058BLxKdkf74STyNTXMaEOFidzsQJlTm32Q3FnoH7oZ0u//epRkghNtUFnItVPFHZI64z2Qy4
e0Cbd2KSrBxk4pxbXp+b3jVtkCQ8EqK7GzutMOrEK1HyyKCs0+3Hdz9uvNxi5QAkQ3E0Knxv3i54
e986fxvSPfehWmZOxaqCWQy42irqdTPDkGxl1VT4laFNZUg3ShKtMqqWI2lB4B0FO8BJ/lAWJh05
0cI3WVL/Vd1zSXjVyGnsOIns6si/ydBPJthRLiTcOfRkZwVh3k7oT7hEFSIzwibOdZ6/zP5Ez65v
ZRLjFL/sqafiowOk05fNVV9jHOTw9+sQyeNd5y42jUhUQEnNKHO04CqqwF//V3FFL26PzgM6C5C5
aoU5sIZFmyJiXvL4VrV+wTD+BClrleGaClp+JjAKEo4ljainaRRrL+3d6RXoa+ugQGQXyB5QFQ9Y
I9dcN6KCPg/G3yYha9A41/9zUpGJRL+j1iA54hyJEo4zILYLQ6oQqZx8VZmZNy6ztvyNr8NsbZU/
eolPMG6a3Vp8qwwCTmR5tigvhEpK8zkGj55yKYwP2OL5uzYE+wD18QLR+mly0EGLRQW/QDOI3Y0W
PTDPdQ7j5LwqVMeZ67iRdmz/5fGrvsDZaR3EAHT8HBeA1iX8lvSuJWmyQIjtCPw3fKNoqqj1/zvk
wXJLSGbgutH0UNMmp7k86iG0vusPsmQ0z8WohNyMbjfDq2q4NsaRvc80hyYwQf0Enh11IEpoKqJQ
yB2oeKgzHCuSpxb6PquGNrJTTqBlQAHUsAfEhHNI3PHbjXtIoImSIs3nO7HhjCF/lYFa0jEUgNQo
ECVRSpyA01QzTmdX73qjb+0B8oufSuEyoNUehlAOl8EcOKRhDF85nR/51yR4tpn38kZu6PFTPMu6
vlvMdXuE5YGEVljxSqIeG2QebJu6sVkD493Cf4kUcjHm3X+xPDXZvC9m42t+qBVUm3FjlvpLfbZm
R7ZUGQzTjtByaChvG0JseAiyhDSHxkHjt4xfhL1Moxh3iA0pvQIW5jC8jX80z5sZsZkltBu12mzr
wAxLEIRsVya6TYkc0QOoYrOEAfRbuPEH8wBfrYTyiVMOo7tp1Qa85HZbOIGZqGeCfAP7IEGPQjZs
XngDab0BcMM0KX/LB7f2GQIdqdq1HJ0T6Uvppe918QMWiHML0/fhN1jxY1Ba0ZLYGAXGcGGDBPiy
YjqjyRzJ12v9PaAK2ZE7qB/sIaq6m2BIObz1nIIEECADEIT7W3fVnQHYqXpI89xot9qKsq3py/cg
ddY85vcorjwh8k9BWYahrG9rCdOKBfb3HTq1STAmnUp7wQMcIQdaMlOOZat6myDa8IyiF1SWHpp3
9BA8cZU6O6igzSFYtgUvPZcVlHpIxGVlRUZTL9ItjLfnls41vmrZGICHwxtzCO+88kiHyxuxKv6W
Je2b4DcZBLZ1DPo5xR8FuMzHY5IdLpXR5ZXcU0hnhaiig9x67rQV9VkFrETZ76iaW5Pi8jxEJ74r
3LpHBfs1WOG8WZOhvolpwB/uLcqQHVSH4GRfN+Oh3LHXOvN8mI6Ho0jrXbiCrPR6l++k4bxoUnep
mFWbUQpcduEQHdqKHKLCEiBL2YfzGZprBpkooQOlZBVw0YjnEOnlUNOV30R26yyX8YX1O0ojORyY
k1IcS1pRqptCebTLo95mqv4beegGXxHcWmAsdwvbTcuDpmFZ+ZWPS6TmOuNSXyktv0wnC5bEsujs
6Y7UyBFtBo9H52BfABflHuR+tXA0ZWcgYCuCZlh+qLXSGUktkY7VjOFPGRysH32D2zsWp+PtfVgY
OxY4B/2ckpYSTOyJud18UxXFUjx361+QUlLAg3As8u84rtKUSakyqn6BNeHuJ/4rhflsVvvbmQXR
PIfHp8ARoAgOBjwGYC0oY6u+KHh955drWBA3nSKTupK2kQFX8E9iYcdDWMD+HHDHXd7BlBKO93js
bIlRFzBgb6ZhNOYVpNk7kZzMJ4oOyqIo/oWDw0EznYu7VGO5rlLJUVX2wuNd+5zNzhUmFYKNVJxX
tWGSzT+7waFUYrrIOc9NdsikErRkJOdvN6sqniCrFtOcYrpwOF36BRpbBcBeBipY92KAgiN9RcTa
Eq02SqdKzw3xZuik/BDzqKh1jHn2G29BVg6n/XXvErTv19ovYoAJx7N2WjcePGEnStR+Ht4DMHk1
r4T3kn4vMH1MxfFwse+ea1vKOmbNpjIHIdu8yvqri8wY0dBU6SGY7g7jI8b5QsJyjbzZYHsNPSDR
svV1jGxI9ioRtWZw3VuDER3OLnODXxFPU5Z/2AQXScIwo051ZfVznko2vIQLDotHBsfgDsCnrM8L
zyLZ0KxJukO9iIjISKEFeKCuTZo2jCo8sF+mc6VdDcb3kkMGpwboPe2XbhERnltPjM8uJD2XNftU
OOE0unyUKrublHAoO3iUY6kz5lozoBnDpxjxA3wRBGwx6v3HovakeWIrEfu8HWMhMJ6FEZXQr4HO
gIomED268jeskC7wMSbnanzZyMBSEXKBxoqVIVD8ia8/82xI+Ym0DqOfo99LVi4yV2xmbPINGhUv
rxRjirBG/9VHOPno4Bu35kN8w4W/NLsnh/EyAJWhBeBXDghYO1eCc7KOs0paF0BKNdPyouPRaiVC
WUDPCbXqnjOgqIqB3k5is2raRjGnvYtC0KB2tIpYOSIkEv+UGIFSmXxmjeKzC6Ypoz8kijixK7rF
VkkPnYCKnGEuqJXUYpIJD7mhYan2qLlxqcnQD0kw0gUQIwj2zUQcBYHOqS4HHAO1QyAtw/1n8hrn
JrICKpS7JxCwT+1eT1wB7vngY5TQYLGxH/z/bxnW42ZNB9y6o3Pz526wnnZHYXcsTak+cSbmOm5j
DxFIcWgQSFrIBfO0cHDsHhIf5a3Lxd02aRA/F/XhBup+6oT4iGOrehvCu5b3Nji1qGHxaZQpfE7d
lr6/JVtTwpsIlf93PbsZxhs1fqzIBQmc+bMRNUs5qLRN0JkN9f5A8F8uoZ42zy3DRR0sunc8kQCJ
XxwIJ8eW9YjFoX83TKDc8gvDOb5OJ6xjrVwBp3Ovs78hZqduHn5BnQAm3AWe166xZZukt16OXFV0
sxEZFJgyNVpa71NwS4ccUfBIBUyOGX6d1O5nna0125WPsNks/WAR++jj8sXS5EW0RZQqjXSLtthd
thFTRebnkto9yk73KmbiNctu6lK1dTeFCn6aPnIAeYtsiJhUgOf+iix442uedeIf1hYJIzsZkuxx
JkB7w7fYPsvGs7/ttH4pksS3papg14EsuKNA8i5gvxNQZDRKcJAe0VA8l1QAYk1g7K3N6iP0wgPL
oLIj+6bxjEXmsadRDHICwjNWMuvOW7CtRQKiZe0xh4Kl5X6CEEkDWFVRc3rwvaSJk2PDn8vKVm+s
wDup4hTwlypGZADaxLS27jIF73GKbBYDq0GfDy9Km+OCliSy4jDxbHlVnqKU/z8YRQM8HGovj3JL
aaFq7URmzNfIRr/yrs5wzLuGEO1Yyg3pNSPjPkLqqEmp/X2ijOy5yHuWMenvxAX7wdTqrtz0wop5
zIpyT1L3yZbTm4j395iWSrwj42R2HDIEn5PtTxaBzFlApE/fLZjTKKQvDbJ9o9kxo8MdCdGr1pfN
krGnwzV7nNw2Tbc69jrjxkptb8NKzEyR3J8KDxRygk7WgEToAdYUR+Fpig76KCvcWdwVIWh750Zb
5GWic5n5OspFKUPCladzB6nvPz7swuUxivSbyjCIpqDpbS9uYK75o9Yx3pavtpONajcMOZc2CNeI
KSDeUSUrOTyrhxsdr5njWxLIdrltLIPLASi88T+Uxpx9xBaVimiAj/cqfQPndRwicDcUZYfhRH3X
9T5TZ0ltZtXicX4As9HeiEBN2bIW/LyLWK1YHSB6Qb1NgEDOuY5gOCQW7CdZ0qGZr060Gp0RnYTH
xTM3MxOhdC7qUBGde7hMl8Ox+R+qzvJNpc9y33zbvLQ9mHDLqimo8+YrEejLkcse1xbsNfvveStG
XR4w0VbUBCHZHzV90mB88L3vBUJSENPsD81jbXPlPAy/HAaNFB8g4y6SELYSxFbW33qK5xmn7kJ3
Z6nIBNE5t1uYYbgVG1EPhwp3sKUN2fKrFz3zOkFuwVgUcSm4w7F2g7/aWGNxqWSk50PJzsC6cn5f
aYpA8FkgxVecFMl/y7mXmW7R5bnKyn1miHhcq5WlEFslQwE/IkM6mOOqLTJHcYYU2ifTC89F6Fte
bct/TUI3XBfxsRpNf9kOoWoNkyGUvIC8YTvsW3zJHckxeEf+iycUF18lMbGZ4dJbUaZOG4UxiQ9U
ANu5QpmXrV2L5Wji3PB5ivaKzCCZALu7pq41neXdno7f8bVinaIH+LcjmMpqcAA5R45NpagvbsWx
QSy9jBvk+Y09pxoXCKD3GUPQLKUx3vLUYCvzIUyv6B0mkExGZ0LPRPfQCVIHI8dzp7WtSk/sDhFg
YoYvGErm1COpT1D0hLjWM/5qeIslfyhTHuv6CKHk56at2kh75Jme1oe2yhy2e6oDahxDeL31p0q4
eTlAjPOAKUnt5aY4vsNkvrX1HZKH0udRfUtQJIe7cWyG8khHng58lymiokjL3zUF5sYo1SLLHRss
BNv5e9sgaBd00Iu36YvfRL5d48M7u1kMwQRjq+WeHKgdBVbq9sns/UJxywHSyjw1bRGtNq9Eq5Wz
Fi5kWNBbL+Sb6o1VTpWJPbU5sjvbjjR6V8q8a8vvHOw1bsRwLLL517uwEFfg14kYVHrs/dTirSLD
sxgjgYtpbleb1SnjaH6JRBDUow/WpSmg7JaAMWii6gWbQKXgKHhTIvMK6oAT0xO3ze2tOB84lmah
PvD0Lu9Tehbs9HkJFHIiBFmXXgSWFDrGjubBZWfZX/CAvCRUjJZqaV+txb2h+2UAFZPiFIuOk8BJ
L6Vz2pR9X0oA/CRIkc+fVQ+Vq7SXujVRAyjQr25y+NqhrPay5rUaHoSSv4pJkk2X+yBEyHhjTmrf
jF/vF6XLUgCW8/R8EfIaj3+OEMuOB2NKA+IgkL3/Mwd+cDJQIYE6yT0RKmdoBEKSC1XFbdQ/DlqN
rb+lsnIwwLV/zvSblxwWfdfxJTG8jjgDDWfyqJsrVAy6GGTvtQ5wO810dA/524HGxtWXmX46jjzq
ZV4eh3QeHdpHeHYZ2fLVGsh286TUGw61xYkXzIO9UWDIEmSORJLIzAd1eIibsqYDHs/p2/MheJvH
07u4FTme+UQJxNokEP2Dqpwrrptdu+Z2QHeHfO6CqUDLAez0Oq7luVuJGjXC5RKcFhTt4YrmkQ+9
roPAuyeNE9jgbNYFo5cZdvoWygNUpqPjwslADPJ7oz2Xu+w8Y+7Pxb9CUS2yaUeLXJhsaISTjHX0
phXm9lVX2fqSXkOxr0ksSLf7T/yT2ZAmeDJq2VdPFVo67XQmnXEkJFHPgsnanvVpz5t+ooxELdUn
aXquYe1j1PxtqKxxdTcsQvc/2qfyVY59AdCBpOYMH1XP6+ZBvIsYZG39KbJmeiBXrK3mRbK0ZnDW
GXlq2DAOaEGRcT2QSFzRRCSFeV5glxhAZViMGYWhjR6/jibsK+ydXDZbSqlwGWoomdlvahRNVtWb
5i6bdnaONuOZpp5X0IdkMoo9FsvLAe8amH2mhrMdZr/2PL93YRvZq8oi50QFFyC6K2Zya4MoVj9/
63755kaVTUAdUD7KG7I7c1dejroQas0sWpYXUKOnHTJ+1YdsuKxGQ3aLMhqVRZeE6r4pKhR1scbo
N8Rt/KjSOr0AYCEFrJ7LBgYQouIH9iZ9mTDQ363dH5TsLnrlus+f0W1bvIdYE4jo3jtoc7bA/vmf
c7j/+fPBDaPBodVJxlh9v6ugmBCr1OQDQacLALOc098BClAWLHioLpWvAcAPICaSr0z9yyeOXuTS
dXYthWspeScozVFfC1cVW3zx53ZPUbhsWdpjTNaMMBgAvs9hXECpGTzOiRzUH5lvTUgQqSFQFrMX
VQB1m5P0ky9Kp6CDyneJ8s+EmV0xj7VOZ2M+wyfhVnq90pz55vn7TNhzJX3EmiocmjjJkNyktRYH
53Boq9b8YeYLQueFOSGxSQ4laC50SwC6fu0/lSmplKuO8XrM+BOp6RRNE+f5615+yTe2m/8oFcLf
KXx1zrf5oxIMC8DrUC1/k3knnAql97aFJFktIS4uOEPLCEYwPAbYj1dQXxKPq36IlqjRFuuFrvO9
VbK3ogBihgm4eUNl+tA9MJ3H1JumX7RNd+cewlLsl7EBblIbxdsNGay5lGTWBCU+3F2pwz3GumsV
ccSeYMGUk/Aa48sXY/MAtm2Zoqv5mXuQNfgDV5KInakW6w3eavL5v0n3w+k07oIRsMw0Hlx9ArQk
wZyorT+P0gsn8EAOlUUidiNoUZq/l6uFegMQMEVPFeGm9IUuRjqeO9sBq9MLrq11o3wNZLV0eyXf
VG7pH4p4ekkawjWeFPlCoYO2Aw7N5dQx7ynrUj5XAca76M24aKpzsyfQTjC8S9yvBWS4lhCe3WQM
tHGDHKLws9sj80HCH7sDXAABDFH9eyseajLEVMWwmajs0mzqIA/B/vRTOSSzh7+KvewyJEpPdBo6
uU153UCTwgdmbrhtG3kiTLCfXQxF6BowD/BVp14QO9ZRk/JEN+mrmtwBSpMKkOzA/Vk5omitYKnr
MVvhS3L4YFML7hyO1/8Og+uxrArXTFPtWPKjF1Q8fP736huNqLJUmu89EYpxGglJFk+LfzKLQl4a
BO4/PTuY/0ydxalyjNKe5xPfQssfUNcktX+vdEI6PUp99qxLa0AtWeqELM/bqUJQYfnuCof69oOf
2Wi8to8yJBA+Fx4rfXAhB550dre8fS7+4WN2P00198dxttvD36b4b17Qgj49cmNYYEF0Iwfj1ytj
dJJk8HNPlQmlzp4Ghy/KN2noPWqcjP0RuuP7BxnQw9B2Ay0h91l2K3zUiuaQ0+mex2cs5Ir3TJWh
wz4JD/59IZj0IpU4DwuFGW2+0B6BhVR875dEUJWvmOwFPsD4UYUf9fqZSfNuQ2g7iPJAMU0bRn7i
VYASFErTJJbJ/Wo6eb3X6HlnYzyeWgW/4iRuIlvA4GSJpTixto4YN50/jw3LT5iXCiac3GSxbmET
Gq5RV1pimLx5ApGxqmQpC6Nu3ZqjsUqYEVmZ/idEFqdN1tNh2a11Kmx3Q3eBO0BLeTxPW7bvEcK6
3oojRtCwP1DEa0Po8FwABCXNVZN1l8N8LWTh+OZtGu+QBi0qkGAtJxkQyib6Sx/6db1L9g8+2uV4
GE9Aq2XnkL0OZ72eLjoEaopsCAGsHbv3dO7YE9m/W1hLy2Tj3MK67k/aCjkkg8nOjTPx+uXP52FQ
HNB2BVtGz/J2q+ymv7hfWZlAlBuZhAHbmFl/gjlTLYNufLjMTCNvr/lfR4FYtNPWP+KrKb1MiHjB
x+F4BDIT8MLRsLdFs2rPgi5ReuL+AtrvJpnXmZ33kbdpaM8ckrX0NVuYupkbgcIIMH8rJV8kS7To
Kbewk0YoSQZLXzA+hHoEnQD2cf0S2mCHKxvUTuvRmqNRP0fAFhkNZiOHxtelN+jrMZWoy+HaHuAK
spKerMUdv+KaaDMXAptQhIFu4E3FJmT1V/hRS+L+Jqo3utkVzvPqxm1lUHuyVse97FUnUrqfZyr9
diZ+FI6pYuVkjFIV3fvfLlCTEskSmlzRbfs/CYhX4GkpQLmLbtjPe3BigpATxhOHzpcLqRrdO7Vj
WPaRcO0XO+3m6fz/Y7ZvSaEp7d9K3exemJ5JArJHkJHv3v/skElbNmVUXer7x4XyBPqG9UsUHEhT
pG6u4JQ/ERe6ci9Kpf3bV/IsQvTJkpjixknz3ThVep/ljUnlYG46Wpu4xo/llc8ak++afGinDyqJ
GoSDYcfbiTrLSNMJv4wmXYqlTyc2XSdBd65XUoI0Vfig8vsMshAxStZcPKITaXmH+22UAQzzVH2E
zWbH8pFawK3fuC5pZlhAQLwDKhLhzZnVEQZTcoWaQOjz9f+NUvNTiGEck1+pIu4TuJRAr/WbxBFU
XcBClVPm2XXyP5tpN3K4JXw+FDVeF0YpaPG6HYS6cV6arQMQaEYHWUxfeVYtJLj3E+SEPePt9DYu
34+M66ioVdCqgYnoiuYkPjHRuu+7+yg7uwJXP7aE+WR8rm0wgZ+Inrw79aOGsDiKJCFH7u2FSdZC
w5lXEIuebbuJ4C6F7Rjqsr8D17J6Ags+4jvwy7WYwxRvUqw89cv9J+CYL7lmF4hoJN9Eh8+d1UCH
UF0/sx/0lM0JJcCaPdQZdwGs6TB3JQvPuz5mNFiLbVtQKfJw5E3uK+YJ2mjnVmTUbAlQxYZEje5k
YYBOXiLeKWWiX9/fIdIqO8zHVhY6ZVwf/EpCWGps1nSxLyxYxB7++q7zX1+u6ZJ5ocTxe1B2xvao
Ya7IlMB8aLmW6ZW61hOtV/iBjnz6kJy3cnysUrXeeDaJXP9Bp3M+vAWq3LqghQOZq5i88aX9tG67
TDzEruqHiqtGGqMv4EEib1ISe3pdT4xH/WKVEhSN1AaB5nBg4lqHRbPY63Ubu26nc2qSTWnQM3je
JYlaWaz3nu+6MaKXUkX16YFjwghaG7LNs+GdHZafhC6U4SvZOEFZIX0fMyUMNwmNpKJMgEbsjVK1
ctMy2V57sGGb3nm9dPwYnaZlBaD/5g2sQxVXkU4Cm+YmbTo41jfleL0atkQLuY/jk+D2LIec25qb
jR9sLDZizQvHKhE6/Qyr9p9+3fhpDklSm2VapNsyffYqURzdIyMi5KPAaLjpnBU94fVrhP7hvRzU
/9sPc3yRzpe7B3+MQAUIjKqbiRPRrTM046lU1NP7i6S/QcZRrxHgq6s8bx7wzk7lU/d+WB6mQodr
nf+VOv6Ay2p7VIrBQErbIGdaa2Zr7LtIQs+hEjXpk/ZmXpwP+4EBL6gI3UXFOFM+IEI9c43i6T8I
UklBQrZi635wmRqDHKCNa20zBHmxpIfZj5aEt2sSds7BdNkWBvyWFlKiYUYNayrFRdC1C7rzh8xS
WdiABIw7Jed1Bf26vOnbPl5AbPnUglPGajPKayBw4k0M0C6betbEMV0qsJ+EactVB89bkYVHXVCD
msvHsBobJVBETQK/z5sboiuoyOu+3MY5tQC42IL+rRGyEhFbM5eIMzsEYawkMLDm3hAQfIWEX7Qp
Mnuiu2j4beM4vJVmdSGC/W5nXXuWbtjHc6W3jEBG46jKgBoMuqOEGO1qpJixAizAOQokfHhZHkOc
er5o3OumhUSbniiHYEUKo7IFLm+XAspdjM0UbByiuZ1zHGRYpuF5wzK5a9UbZYaxYw/axFMh/V2/
he/H4VnHIw/hHa1wZBJ+b+O0rjSpyoNLeCRkfba9i61Aj0ruk83w4l2Gk0Hxw6H+jJlkDAP+Slxh
rNK8ezL5r0+8pJXtFRPS+kx54Fk3rpjYXq0p7tE/Iwd8UXe2ntvmtYU0GZSzSvjySICKb7I6FkvR
kwHUnTyQAsuOmuyWXUDwDcVIty7aTbRD3vH+YM/YehA8VGUHsdhqQ1fcJX/MUJxHh7MOkpkjWwxd
tAO21eugdD5vT4ELo836gch3m1Ur2gYq1tzfLheRo5rbPr+HWaZG18RKo0NnmDpfU4UJLr+R9izx
1PH7ciy2L9Lv3l22OZ5IvDAS/G2CCeLZChwvlHtwsPT6/B7lxWFAHzp/zh+2ma7mut3TuGM5rz/M
yuTFc7iCbWsL0DaZyOLZWGbQ5TESBXnI7JwoYdsr2pCYoM2en04Q5M9ty+GYX5r5+rkENHT/Edh6
Tdxc9NM7Lu36fyeEwkZBpjJAr7u7SQ2AIDY7rNVxPDq6czMjZsBKdVWfM5JqSThUaPsLFh5E4Z2w
eyEeYv0CH5jXmM8LRfWMVZOUJMB9LgkQwdz2WdXu4Zt6EAetYieTWtrgyc5gQdYpJ5ftc0YC1F2Z
VLpv1ovsoNdchVhv4ocSlaPKNi7KRlmfTde1MYt97llREgI66L36Rn8xuV9VdP43DTyvH0kEN1wI
g/y+MbV568UVbLfx5Uff7mq7dSy4VUV0gS7owF5dxN/6WNTfQ0JQ6LvXzscm2hU8w81H6v1m4M3k
tkaUdMMNnss/2cLRDLX5Ex4FttSZ/N25EVAbepqOEPQGSLdBqXdyDnFDuYGvgDeUzQbGZ1PqFRr0
xQoaNm0yiMmKs8lGmotzTGZ9PocZWx03tVuTGDtS8BVSqNux6G3dMVaGHqED6HyGaeeUaW/KUkx1
joRds3hSTvkLgv1uOV7DXHF9vwkOEWkyanhaPNz94IRPEtMabewchg0ODHJzL4NCg6rF3nPR4fwb
TKjtM88bEc5UC1yWlyZwoIBzReY3MHd+t/2o9lnM0vQrZldplzZ+5v8r/wq7w69b01CCTKTvsOa8
X8QsZnBtzLWsubfs9QZ8oj8H0nIN1p9xuRuYf8lTgGXqDebZ5qVQgGL0O7S6/C/eJxLC7HsxKLJt
eBt4slFi7jiHSLU6suzvICcFV3FeVuUHTGR3OcaqxUWRKsJ/s64iU2qL70mJMQTi683nIZTpBt9u
rZY381YgiqevElKBcZhGgQ2CiMS12K61/4GSSgP/S3mCqc34I/SgFjB4BkGeMdBYiJDwIzBYk5QL
L5q353PIbrukSP4EHYzMaU8Zf/ePbTZqrNUb2NvJLF2qKtHdX4ZModyDgmhbf4Nh20BcH2jTOuTx
yYsXvAnh8r2HBLea/NaYSqawV20SbJO5rugngqyY5uEvz+EtaxDDO/vt/Xcy1YHYIsQRRAiIzjTw
/iN05M8CjAtUzKRDcf6kmL1NHVV9M8WwGEKMT1Udpjr0Mfay3erMjwDK9JQY362jEufclVL1N+k8
PWaG3AFjE0C0Dn17F4548NhsbBNieFZLKEjBEzSOgdU3CtMBDyQVSYn2+//3f85X/LK2fmNaJWhM
8iI1s4tG30vhXgUp9z6DAbgZAfgZXmzi4ZqFlaJxte3N6V73/eTbi4PphbI1Af06HQvsDfTgYExt
9k+o/FveNnJYlkwQf5iFgmkPlAIOVra98MynMLHR5u87JlSMOzskPrk8mUnHBIoe6yt/ygDOXKfU
8CzN3sA47DJnVIF7dMLoHluSsy2VWS2vN6D0AiWJ3RT29Xu/bb53/wknR04mtaCSE6SAH9O/1HHW
XZutxDh/Qqa56hXnUu1fYeYjupF2qGkBYQ6Ym3nsXsnhNJBctNL3U3hEtr6F+1Fz9t5zmdGCtvVU
d01B3kyZnl2JqU56wHkYeHC1N/U/1G2ccSvQs/I8TsiNroFnA3rnghHh48tM8U4mnXk7fizgpDnB
2c3OqHIP2b06vTyOaEUjDWgmXbhpIE5rMOQf7d1BiXsWcSsqQfdvEsVebvDA3Rc+uWQQbetHJtD/
8UCOGUCND443ZN/nFJ3K/quu0wQnS4rk712/Rc36J7QGdNzKqtSYJd5ymUqVEbN2UIynm4LGu0hi
6VbBNN6UKpGyffBYPtak2gVPioyJZMqyKNGkuYPRiTTTHsZgCWol6ucFDmDPAe1aB/PmoiiNVhMB
H41S17JnxnVi6q2HIEfSrlxcr6lNQd8UIh4hKTcTODGVO25tr7e3ZlKuuXJsgs507R5uR2N1iWEw
n314vDeQZjQ9/w8iGUfdgF+eksOzicuTKxTiv7K0ZO00AhibFj9ye5+stvBd82AfWq96nFgXq7l+
OuE6vRQvwi4IKrQPM93M/DXQkaGtxQ16MlKdb9PHhgayZxdc4OwCz8prF8wOt3o+i0HjOdlfnjPt
RgUzaWvaG4BYtlrNXjmuVR0z94lF4j2syceVKL6m55K7XHhRVosqE1pXva6JaDR7m0JOdA/wfKwK
X2merBvbWD/LfbCi0SlJ4UXZG5nnJJxy6UeUkztbNNlQCDTp/V+3YRAFdACLnF2EzL0NmGUDKB/8
v1qwOC6x+4TN+HAiPzWdn8EbHsz9cidtuJ6kmn+Qx8mf9SysDxlpcaIA4aJVnV67n053uIB2YsqA
o3cwhcOL3TzKp+rBHCcX/KfZtwMxI0JpG6K5F9kwbTojL3563gAQ8XHoJYmbr7dFVYySH9l9DCXi
FxwspD4IFMjgQZe3UVlcrlKjkPUhOrz4WDgJPqleb2VF2C9fJlAaxvrCUxZdqkSUENxZuWYG3Tj7
zavFpp22RJsA97rgOoKczCU73x+9moctlAOiTSs3D8hy1ddv35bEW+5AesEQQW50whNy/Syykq9X
W8ck2QA++qr9GvLdllzaTmz+55prifCdi4vzkbFQYykVfDyxvQaBpDMQwOhVkqizQ/OrKpTrsgHw
7ZhIc9LtWUAHlEMmckbsQnnf9SV+hR/K/MHBQBkvBQ6kQzwhTBqN1H2/hd8uSg/4CfaVaQRLOa3/
YF0fctQwBtVYIi09mYrSvMB5NKko7xc4f7ugpQCM4JTkaAhLDrP+SJJi75hF+NRbc3+lzth3BoVq
eq3eAk9o6PVyx61x9GYB5VzuWJ00bX15ZYzR4ftu0EA9yPYmq3a2hvrjfm0MAoYywxQgDqvgGIYL
r0nOrqS5CuRsMS72AyLqtGcA4l7VaydHGv421oIilzGrB3EqWMbqx47D8ivnqlQ6mKpKOyYFqAWH
o5VjM53uPc7BovxCNnqDt7OzuCWmqCnlw1Nj5z1n3bZTBgdlNgErDwnpQfB1tnt2rR4SOoEAS3gs
wpJhXNUlDFXMwtj81ky4IYFJhXXxs+kcbZcW3w7ar8HpRiGqilV2sAOAZFVP+FdQ+B+sXouvp5bM
dzrqK7KuWH5bIJp9O9j3Z8TDD2VoYC0V2zTj7M/ojBP9BpvBouDNFBcOWD4mAPPKpZApUuFSS8ZI
lMbQSk+2scTRbdj8B74w/Hx95QwGlAgsFk1OtHMX31hllCWSHClTUy92fwI3NL+93AwZUJdq880L
BkvVgj1+DPYkkhiA/NawaUEqVZFCAy5WXDEYTLkIFXXfss/5eFXOvoKJCp5lN34vf7a1fGQ1Mm68
tSWwpEOiaymG+pp0DZWKi2jmQd2BOgxBgpG1jzPvdmIuWmtSw/oQiKFcDo4QtQaASx2OzDLIz8Z+
EeKAFB6u/DdpXECYHILbvVGFgdvsuPMFMDG3Wsm7ZsPyNGgaxzt2MzQ8rGzkzyc5dXetn2Aa6rKr
6fS7d6yYPgDM/6MKLiy6raHBU3MqoRro55voWB5sraHkNv7OXttb46bBtEoDB0e/U8CUtwD0NIwJ
V//BP8K2V6KSdKEMmiYbTWlqrRJP5wTg6ClQEW20adDU8mfl4Vmg0qSuhx/9ynv/8dSdznyQY8Ea
wEtljNxbENjCnWJYTD4s3SNnD0ZkkwW75OiqaYK/VJjyVM0k/TABKhrPyzKW99rMwSJzl/NmJxud
yK8cUrdbD1vALVDiTDX4tki+tQXB859tIxfi3ys9+QR50j3+1tQ/hJ5Ptjl6cVQw49nhXdp6PPWe
B+0CIixXZNYtD2baeh/Fy/jEc7l6XJ+nfvMGszDZQgRy49lBTvHpl2rpVgSWEnSZv9NwEza+toOL
3iWasaTfSTA1cr0VVF67+Ys+/WwCVGRKlwWMPQm9u9egeGCLVjxJUGTuW2E2twQsbLtgrSYJp3JY
Q+lKjfo/5owYRNUuntYV4oIZl9ozAErtOsfRBpylXHHGqWqExsOVKCELLxSvjUewxpk6ld8ta46P
lLe2sq7el24nOB8DizEnxaB31YQU3jYiSAfcbfbBZLsa5o+o+OXaQr4O9DJv1xey5cg0oanI9Utf
ch5H8ofFETYFl9jzv16VROUbymVZl5DmP74vCeOKj96/gYSXkizIc34y8N9TOcW36BtblpeW5HF9
1AlZvh/ji31B9ULLQNgIAP8CwfCpYWX4YldpVA2vmIvG0uJOGPJBUJJPVWmUV5/KwkFLrAs1T1vD
GdterCdrWjY+7KXl6Cw8VjcrAfmlyjKSQEWiBlNLc7xUVFIxT/T4bcowL38bFbBnEyxAUugyeiJN
7Ynwnx+L1KoNOnTs8kjjBCaW62vfEz5WGXF9BFRSvn3kBfBfFUXBCWJNk0SZXOBRqqjoI/ZmgKgg
ixlP0F58cKIa+1HK+9m5vE5rWzGkXzXAhJmm1FR+a7bTh8P5i1wd/DZiwLAky3tnq05qInGEeO3+
mdALDPAqqUpgtot3AMxnFKuT+HC4py1fW+l1EFobM+oVhXrMZKm3zn+EfYOFm2uF3A//wKwITOCP
stwGjH4L0kUguP6WhdJ8sIHnax5OjeJe7rZKIUUMhjhRbt9MpHM//skWg7+TL6ysZUXPkk5Sd8kp
hjyogJ77ePkNFuroQLN2qaHHFIhC0+dSEEfMP7EqfoDzxko3jg3MCykcK3duaI+OeTvQqA1Dki98
oCux9qdI+DMUlXZ8aDqBj0/Ycd+2EtpEfoN8ZPcPRxTgbDM+ctR331FdEqixhhhGRD70zmaeytCv
dny3Kmc1P/MOE3qmdn5eZ7KkmwE0oxobEal6JElWc8IzU7rEiPtNk38gTAFyv3h8rX3od3zSoSEG
Zwy50Upv19g97b030NIdmM3bI+4KNyoQHZr64c7wSeIlykSNzQk28WGkVR8ShShQZSOXt+UoYLSi
r31TL0wh8cnQH7LbpStI+5KNdDA/AvkaTSO9vNZG4FEoGqmRhynua/i/34MkIlkV+yyy/xxwGcid
jBTDO8YFd8DzhTAZNew8n+T22rRe8QKzh8OriKMS5mB1NVR0uKYDCnhcsTiYrZqv1Ja7kqClZ3kr
lM/WdHS96A7kuoK+djfqCWcKzsHCg/FHp5PZXCLLGrb6xKm7KGC61qf0B+zrc3FmdPigUcczqrWx
n5wSRJ3h+EE0mubBQB2am3NWrfOhD3r5DQplwxHBpV1zEzarwjScwu/wu0BzRDClKrjaiAaGNZn0
FCalWnJTdXVk602D3jNzmlBhVg3RUdLV/aE6BrInYBk0/1a5+ojhuoUch+IB1KbNrP2S4Xi/48LA
byuIo3kE55w8mGWYoM42Xtav5vylXCP9mGP+9HP8L3uPcHe94yZTrqcB7DBVf85tKgn04RC7dW/E
2JOFfLC+AmZhNpOXcDZjTEdfu63dTjB6LlexJx9QipShVFniynjsMDm46sSlObddUlxSGHeKhFWn
fwuIjUsf6UdIDCC5XlwzoizAcp8OP5t0EP+AO9uiwLUDPMI65hBBqNpOWqPd9I3qnn1q9AbbmILb
08949tvOvuLvrhQz5mXk4B6/FSi4+KF//Q7VwVsylNSVPRHQn8uA8Ooakwpyj9Wuy+s4aVqQ+qif
lyDOqylQj0r4cd5dE0EVPblJzz6rUthmx4qK1UepoCzqNRfuMTddEZYA++1FZBXxHPW2lRqDrNRx
WTMYQwQNrwDEyW0O6pfK1jOosRmCPuDqJ/MMnwCl2HYQFovW3OFkANnqsTGrdFiEP8/h4Jj1BUq+
Au3DVfEpq25VTPCTMzVM+BhGWj1n5y5YtqAYfV4sc11A4bnPWCDEwlArdtkfPcb6oX5rULaZOFr+
t6n73NiV53wjjwTJgd4bhkGw7QZPDuHcEC1lS3DDT0wmiDp9cWZ3QjIkJ7J/A7/zNHuM3je69n66
ZpvZL5+CmthKSL9JIojy0oMFHipaxNda4j5bgc2nPrK6sWQYjJrakfFnhGwQq5oWjYAZtEzMAG3n
nyaH0Hli9UoFK7a2enJBcc3/TGxMywHDDrJV+RhS+zgXorkYhiZxXEpfg3d6uD+9vwcJU1qmMrCZ
XZmoFTGdiyd35fhBdChzYlruA4ypWiH6G9mJUOrwJ+cFQCTqD48U/Y8PU4ACapiW6bLquJuXIRrE
tahFpHvCSE298WbV4Q8xLJ427MhWWN9d5fCleAqvsHqpCzAi67+KbnjCNgBZ6C58qwAG+N1l0c2r
IVbIzfbtHGvfBQXTGJm+aIeB+tc1bwXUQ1fWA64EuZMeAET/WEKfqib3bXhdQ9/bPbTqyPYFpv3g
XziEqs9P7o4wMD9/iVEQHpFY3Rolz52C0QzuOaj7mxfYHgfX9VMssHkS/0MRRqpzEWQ+dYlx3CYw
YfQo9ewu1AuzzUyPFzoSOpCHSxoJT6sQs9E74rXxYFGCENCqSjgfjNEhhgS35dzjBOjy8pc8qUkn
zeD4234hSviB/exx0GV4BczCrK7yvf+eSnzGi749FYIGg6xZl0EVKN7L3MH5/muai00OzIzWiHFK
HQogZCnCknIqECE5hh+g9GB40Yvmtno68nLhORA5/Y6Xmos0l2rvpjkAimtmuTaCiPoEt2VcCJOo
R31jtYp+BoMlUdQiCYrHpc6poaya00fAJVHOp6tpScl9xdUlE1zLNtHPQ+m4c3Bz3HDItYcaBD3C
n6ggQKAhnDN/a01fFvQ8JQM+t4RoJpLSHOpktxjt4IDND3z6b8qPvcYnqZbzsqQlmTqcy5XFWcsp
n2jRQYGNzd5mmBsKp3IJLBCbDA9T7YxDyXYM/H3qyjv8oUZFieobqGoDYShenPmPtXSwUK95WqMq
dBr/IruVN/nEJOVFuZKIE8ezV2+I3yiDmmfZJc0jdCa3HPleEL3osd4J/s7t8qVOEP/ET3DoBqQY
EJWthEtqxij4eJfB5r+8eAWYote9N+XDy36J+CJflWRdN6x3S8UsdCs3IidDYdhM2mqTypWzCFko
F+w4MdTm+oln2w2Zf8ONACehbIdtN4VgqptbBbm99wqwEqOv8WcHeYzFdYizHWNoSorS3u/9sBgY
c1gCxdyE+529lCpOLB2euAETBPvvOLk8muCrt9P4bHPe9HGi3fPSl11CHP7whal/eqTG3DKuS6DW
SJishmjYBill0b8KnecnmsCb+26nWWZkFSNGDkBz6Fl183L97zWd1IUsueUJrWLGVcgBbVTlzHp+
v4v8m7G91sr/ujG6JVXoPr9lkoDas4jl2uvpr/jZMd1wMn62uimqfDWTHbaXy2H/J0aYXt2A+ybX
wr+V72PmV/M2NORfUfP4AwGBN6QGHtvw42btAe0fcFAgmBNUPZpsmT67DmjnDRQ/gWmkizY5OsK0
X8cB7BKf6N5REaxHKIYOBpEdiiXzrlDUgizo2dYs+jTDCLY3VxQdsw2nmEZghgjLDCrXCPcyKxVy
gK2YQ4cOdgR1/jgsv1i0cUhQH44nfE1DIqxPLHXKJAbeAhSAjOIy9R97dxXrX/ZMTaZoI6lGwdpf
6fT0FcpOcc0kTONyfmelHV/Bo7rOBx7NKGrbAfWGRPcy6io/soMWvGpbZ4DMYIuDyljhUdsG3VAE
+z+ciRxWdJv9pZJYyddnX1fvy9/sY7xi2iN3qt1xs1CdH/DhUejcPHzEPsLIvJQzNBJ8Crw+oFH7
qButhDNaP69UY3We0XruD573J78MNhkZ4V45Qqc338WDDBlinvhwgd5wSeshbhGNq3TBWUyNSIvH
lqy+UjBIrvaPiEFuOTxGaQAosBfO7Boo03qTjYkeGV6uZL1jeC0L5+XzESprDPY4KfG2rZcBn4TM
NgXzpVclIb3FUrNUv1uBhlMhDjKH4o6M/oLj+C6KqLWiZyCiaIfZ35P31nY6K/oagih0rGyI/HjV
3Vv1CTrKC9jdsGV2ETvP1rH/aSdBZCNfNUj5xwwXxgPcjNVdfqLi6J5MMImvILrUqRRkoDKO6vUh
OZDo2UHebOuHBC1Lt7nYE3BbrVvvnQs6TBo4Jp5Qs36QFtmOj2MfdLYd1yksVszYXaSHuLdPHtol
9f7IYAep2v1xkGS6KqxISlnFckQeFpLFWtTJi0ZNG6X/OFCL1y43H1h4o40sTIzXFz/7/+fEmuCk
T7j0Od5SabWFQI8wlV7+T4NHEng1BoZwoQ0JSyhMV2k6upaEugm1RfrZ9rb5+ARyZHng46seUonA
H7UyOrMGpvTrMp2CA1wEJALIG0OqViQ6diCi2fpAT5Pm/BLdQEQTLQgPNetxbGo2zfEpPrXdCBmb
6iPBE23bFlN0q067g9qZpJ/x6RVZpp1MMWUp7H10j3qfoYyYppswmeoe0gdWtmakEYprGRTTGxRf
kTq/069Oo/V0KiksU+S3nXzUv2Omd6dNufEhUC/rbCXJ5K4KZR18o9mNADAhXEmGzw1YgvGd0k73
f9RudtNfx+O/aZ1sneZ+YsuAwFdDyX7k+1UnJ8BE2dNn1eGZoqq1SlYLv0C4TlLdIfuX6MCMrhsc
ZOqH1OQ04xcT9sGTrNSKP2lVngRrl6TnMfDqo+FdbkXhiRDxwhPVLjV4meCAIUNzdg5/wM4XGlAu
uJEnqEiWZbVLjLWKOfJNiehQ8pzc6e0k7X3Re2Pwx6H1bnoboMXF+/0GzjOTvua+dXGEtb0ZbDmz
VQJWhCmDPYBnLPVs+hv1QV1q2PjwWoYTV0MosebQGdg7kLnHirySnmrYIz1IrGFmFUryBHyrN04p
E+A/cLVBjyEOMpJZH6XsIrfBnSKprPMnmr8zjX9WMftsUSp+iEZp1Jj8+ROnnTm7VWhlttAHdKIv
8rsqs1G6/soatgdB7LeH4V3Ov84UVmmVYpSFBQLRR46ETKSiIwWYahEZNK5mrhnaAHkOfBXHTmsU
5WYDMbNNt1+amq0T7Ddk4Z7BjiLn4vy4FjaDrJ5yCZb3HxMgSo+q8N03+PHbVHKhDQ+ab9V99QKP
bliZWkGBt9ZHuIedeoZH2JMqhjs/5/G5PQifw6g5lad8l7VmjeCxlyrUP42REoxzMv4the3OYaRF
ajxWY+fBl9pFLk4bEG/ksOsRp/UzVp9otLjpY9WDFnhcbSo9p+SfRVtKt3XMs+0cFBWQyjJwJAYb
mdzRLX+uopTzwGKCOW/tP6r4tXs4GeMOe2I/lhEEZvZaZ8r3J7IGw1THsrefNcHclWlzy+zdtbb/
Z9J52oo3hAQJkr/ZjhGtadlyCZL6xxCWAgS5ElytJnA5EZPibqjyBVpZtv5OoFJsRq6L2Umio6Om
pURH3kzk0vRcT5x/whaFOvVHaf4V1KP80sAsznZZBdnx6AAwT4r6KWAI4yxpUvgYk6rixR9E0+oY
wJ7bkflNqEvgwFtiEcveZ+qiTmJCvZOiLYplKbSH8uvopH4CP899hPVd3aedRp0+hKhydb72Qega
PfTuCWtNYItj5qXjR1fnneqWnSDbg8GSyWt6D88Yt8jWkHamcM8gZEShbpPrMZ/iHjlMY6I1K8jI
VpML5ZqF6UALbxHEYp8p+jvHcIduh2if1Pc/DEIgIU+rKnEOQTk/SyLUZhvAH5D+u+jQzh9x4zI5
IR2YO33X0pryy3hHNp2uUXBpVt2H9NdTAN6dVoqoDLyYMz92iBVK2U0Zmdih1QdnIazv+R3XgwQA
pPJiMMhIw/s47iTTUef7vRgeFTjxvKNb8x/HUmQiJzQxAWuRFNQbgH1xexDyXf0i+xYdEiACSfNe
9w4h7DYcik20XyXFJcfo3NdZNgFu7QeKnCpdyA36JM3Q135IQLJbx0/QC7DS1oNsK5Hn+OgfTr6r
LdAOq2/5KKc7FnM3UijnOenVB5JkkVFBgTd1RYNSIV3YBlBVwJ9z6QPL9KSJnGSSfNAXao8GZwNZ
WbA5dPF8re0Yfijef9RHYk3r30XKoVjuSGqFcffUSzQmSKbQKzLZdfrnzxwvrsQYDcKmWGNB4Pqb
mGTul0xSqKRwzysQ/UsOIcBHsNf0KvHCNo0n0mlu9aVnc11+2xsjuaR68rGXdrJhHhapQi2P5Wx8
1xQkWjgEM27T4YjaurahMIFnwVi9Bqa9RHodUD+JzaCoQ6Yar8viH2QPUJnlG8I5nWQxN27F7MBG
fL1HbICo1yHGqTAimg5TLQe6C8Gk1ORzDKWNcVLZiixIeR3QNAqu7DXaqXa8KT/N/k3pZ3sOynxz
0EgknulMMZ+6HJO6/dzYrcL+PZZV3CsdzsMs4LwGpdDqzhnIbW1SHHCS7GhPgPPyzktO1+ZYLvmL
RmWUnEefqzlytxyH5iNK4o9tbljjPdSwNj2w9CNdiDWP4QK1sCpy0DpC6TB+mqkwuH6Xo4BeVPFY
MnDXF1vx1YWKLdrpCpaI6bolyjQbOxXjz9bjpKoR9x56MNAfa9OWgzOAiOZ6zyyaQruVxWJq6Idn
ny5AHzHT8gEjl5VmUG4fnwqnSr63iqji/hBmplauiKTebj6M797YWbd8gWY5khROi3896MFnnowB
PuVZc86Dlm4t4UtiQp4/E2DXXZXq7ZHtn1NtYXHRQLhfxcDumfetyG8TcTcV6OHqdWSQTlccAb8W
PNBr/OBOU3Pgh9N7t9fcl3orR5MRAxAMN5ZayYqwuabGYkWSwt1c0NOhB65AJk/huI9LdhLBrR+l
ZtYU0WCz1TDegO9ERMibnrMO8gjooor2OiCHRFdC45KLk4fOn5SipdiTvePb3JhCglE7+bciOZIB
q7aVvXejlnFASJU4IhiyC+/L10AxUSYCwxP+Djh3LDjqTxZbHLxUFk1tmisekrqefmob3+uIYzkE
8Loa8Q0wNjc/gstr3oQ/RPrWxJQ9gesdgytbQP9/mcx3trsCEDIp7cxdC5iHBrTAujQt0229eV2R
yIS2W72fV9O21oKFgG+NUTPC3LvL0DxGpYISAhUXOrCDWxYOmRFbVrC1pJHWOAbEL/5oaoshObY1
7IggPeeG9vDJ5972mmhprzV9XbcR+G6J8IkgGUrYZO9kcrLRnumLWWYgwa/ih0sTJewV4QSIWHxn
asHloD07g1flQp1DWP6uqAwckAol9r2BGNZ+onnw3QTaWwHcojCcq2maDqJ9Cz5w2J3uTM60n8Lf
TPpT/IdHbtJHDJB+uz1CxByu4VyWVr2MLGFjHdHAyjm9GKRAbAJRTtiufdwv7XaQVTso0bmO+Y9G
Cp2Qy8gYKIRcUt0Gx0PK+tgNx+2VvI/vyL7xdD4n2loL8nZ/zfkfgBDbwzO9z1bFLEKy3ifBQNk8
HW+ZP1wIrhqcgjzp8ZLqAA47sh10ugsWEF9ds2TNVwEpBHVGIQOaBziexWjvz+4LOW+AS33sfb0a
0D9ieNHBI/RDXuUF8hAc6POJZmQf8W99jOGHVcjWr/Zz3ceceHE0P4XSuLPmRoRN+ajhTWpo39i4
750DspJg8idpGKvIAbu0pKt5Es6Lr4V5hSgVKOiu5sD3KieSIubIQY+ZTBbW42ezO3OJ9+XCb8F9
xQkxXfkXcpXvtHW0ico5GVtPe3TjsHUWRHi0o1iR38AOUWLm/LI85GpJ0VF2uz1LHHTXvmmRDw2q
ZWUVAdMo7d9fB2rL0GY3/FsFUhl+/XPbEAKLXay4nc6EX0rcQoT6FG5cv2H9/tYttlJ0scMDLEvR
j85u6tgnPnTFUfHfXrxKLBTvjjLRhKx3JOtVecD/clnnp2ZoOIUTHsYCSUe36Cp9KsXOxRJOVWL2
IPbs2ixeAVqFLas5R9aKbkCYlrbOKfzMmbMQSxgJmRsq8gaXE1Ev3Dw52fgkd+Lh5pJSofw6QnKt
d7nXOJe+SsMEwZEqiXa+IMC15XBvEIRWq/EaPwUIdQYazi4Q0CAqnuJJoIdslTibdofiam6zsGxT
wMXq77WTKrQIQowIpdF7ROIc+c9xX13ZpKhre+JbU9c11tV2oz+hbymvCQZ0UMVP4j6R5MUpYX/Y
nUdVSw7S46pIQl119SzXNbTFhX6Ui4wUz8u6RS9JRyGQ+q/FHIXwKjdjGB0OQFbhtZOPiKqQe1r1
DWko3yTZtg5eWilZ7NG7MCFJ5PNHbOzvH1rX5UHyYlQyGxfHhqDAxcfvJl/O+vgo4EjETH8S2Mgs
dyEmSYP9kaxga9grd/uXGKroz2nQLaOxwF54QWGHU+jnS4lUYo/EpnRW1yeSJHUXnM3t7VoUgW4w
fqIHLz4uiv9NJMjAi+EW/wcxB0oSh+bIY3xN9fLoA3XrTV6992KCdEAM0jSMdai7CfIF+zyRIlCU
FR7zNI99w2YTPdwElUuBQtKKRnF3Yr+4hRnz4igaI6IL3EYkUvVrHibE3F8thW8c4acNwsctG8oR
5GM3tgehH97MU0xBKidAYcy9nnBGw5jEC0/n3Vg0277kM5CI8DbjB3VUZX2bBUtROHWIgnXZDmYc
iNAZQ5aoSpSuBTFQLCQWTTIsGlimBjNGvKMEP0R6eWcs5hB8yRJSa2aX0HXK8DoGtVPgEw3qYM9v
RpypWee95L47LCjrSstiq5j9cVu0ta+yGyiCAqfol+HfEkJsrKEMoCUhgH+rdFKpX3f2GWTOLxYD
M3FPHohkRh+hArSdKCMh3qXe76dazhX12TnRTO2AzPO62M/sd2/pfXFfM2hcdhIg25tRMljlfExQ
NpmiVbGKaPMkZ5nC1h19oMVXvB7fCVN5L6pDUfb5grW2vD/wY9KPinxCQTaLElkJMwe/QGQoQMqp
x5uz6mxTL7xLsgbvjAGdWDRTKvkSQ6eT19X3y3GkByxcrl7CJyO3fYDFu+Sgo1X+agT3p06LvZTi
bobx6813O33p+wLPkJ0xMAfZ7FDDmbD9b9jaS412leB/vJnTcd79OkKwbcVqTnapmfk/K/8hBBOp
ZVlTo5DwQrw41xxLvSc/ODOhFMXwoXje5CwJitj6dGIuFXM1lWa55fFG7wC7A1I0S2doGhFOlcTR
ylSTWxkx9d84Mm7QsSSOCIOS+xqp10zLb8ic8wPZvWvjoRdblpIrYUfW534vG9gD8yT2ATkMxw25
QSGayv2IOg9RC4nZ1j2z48NSt9h0t/9wKLx47VH3hDfV6TMAKlHt5d10DqU5YP3MLW/ib9RhVGmf
hPb/553jbQF8a/I1fHCinEjXomrKvZRY7e6fyWHSTgATO/XPGDDqtJMjzwhFy6q/NoK4+JFC9O8m
Cd07U8UEWhzYkkAJHn9vmKQjVqsH2eIOAEi8431wmn+3DwkuDwhTJHWWvoAVme6QbV0dWQ0ysfxF
f8AWURiRj9hyhtEwyBIUt/6nX2M4KRpXk8UOWRbboZa1zPPUcBpzD80Nb4QM2bRs8H+bB31isf3U
oiRUhHAPh1a68YiD8CwfE8hVM/Onb+KHjsLAjJD5QIjgAAEVok8vVVoxdACqKkVrffSaoNhz7YjC
WgDh6+c/0srkvd1E1OxXfRv7YkbmDrr5A8X7R27hN5LgBmkSiZmOD8Ex2xG/ezf3NHNeDG9YKCNE
xDD+REZZ7T5T9maPJkwLOGRzVI168SO/aUtnVaSBHZvbjUVuZEXZSqdYyTxx7P1V/GZwmF+LzlVh
Z0JmgiqjrU9h+6H9qz+87gYttCPQrjIwaDugzqx367j/IMzuxWbsGDZ/iX6HCHPMG6zD7zDaeuaq
NZoFpZ/K606PhJF/ATSDe0oO/Tk9BjlBO9222RgE/GK2wyR3m9BPG4DG9irtwIVgaVZck7QWwi9Z
AgnvipiFr3nojabvUAfWJ/Pj4+QcWrH9eNueG1CHvLK2xwq9mvTg1p22G5c8MGUB1ELZFZT3NxHN
pXrb2hHFPPzZKC3estYRNFulvwe4zjKSxMLXyGIW1/CEkAwj41u/QHgQDcCAGakoj+FYNNTSf2MQ
fT/ipWBkYa0XlX7d+n9wy6ja1pd7uf1GWTwl3r7DJzsWUCYaiIGEJkpl3HYc99rrJVPHT/am4Z1N
2eJrMpv63ZfIIYMsMVMcjjhNA4pP/NjIzR9qyZJBGFbyHVfVy5GVijsH9siu9727nuIS5hwPGg06
BAeB7fJVU4Su75VO+l7EClM/ufRC0OFhoy0ka/kQNzpm0njPWYp7VIwxD1Q0BWhnckE3F0rQ4l9J
jzZ4ZgHlDvWks6nXX+BJlOxypCMqijnaPuJTunHEZ1AzB085qiO7M4LoA3+EBaYxmGW33lu14jsM
qkecYDiqG3aTErItEf1nVoYYSjC2QPLJbFc/sJrGzP/oyP59W3nkUKi68eW0sJMVU0e7VsaegTVn
iiEMgBiiAbph5h3MPHu1NH+6Q1ZxQOgcekZfOAGZpBbqYMxNi8c9FBftI05mMTPWTY9GX4K51oBS
A0QuCrOqNcXYsrQGcU3ih/q2+dIank4P5L4ajXPPRnAGK5H2uXHhHGDJ4vL7HjsjfJEXI+9kHuZY
WYf0ciJ8i8XWI+G0p0luNDxg+oCv8nhu2VxwnabmnR498EhGXpnzO4riPc8P/KDL2v3j1sxpSRvw
Y5BAw7qHbtjsXcUDB0rP7NpwiEtnlo5pkUJwNT6bwaUa37nWGRyD+9miJLZl5g0d9f1ihJuF8id0
TVOLw8zjGrt/raK+Anjdeh2r4XuCYhNXdlL9Kn/MqiU6IfPDVx/m4SUH5eVwlQQPal73DvAtclh0
5FhYYHzASQF8YkzJ7QvYpidJrP9GLi2wOy9igoq+/efmmf2kbPGyCSKI0ehNWTnCieMFz9iFeOFV
T1d3FacFzT/ZePHQyx3WD16M0kPFPaPSC2O6JGIo9m+u4UQ+Rb2QXICCHGoQAYeCHQk43cnG3a6r
We7y0clcvg1zc4C9I0AHXMOVXJI2u6f0puv6hamci1cFDEw4/Eqd4Sus+EqfUsqMH5B7yTjg+wgU
Pe4vN2d9PFewFnhXn4RMaVX5YBso9Zq8JgcyB9gFf5hBghDHXi5+nzvRjpzbX0nh9vnoepIW4Kno
GOgVE2U/zDzaR9U5fRHbugbvnGExBS+0gssqGLM+RzUa3IT/LCJikjqczoRQWdeadH4cQkWmOmWU
F4kzfpwBc+6JfHUW0glhngBP6mUFWQSDc2BvJEUCR4+roEkvpQ6mt8IRkgyhOIpb5OnZQrJeC9dh
uSD6dNULen8RS+o/E/hdDTbJkdeOfuTyjeCLJTyIX/NAPsZb0it6zDjIxNeyXXB5Gjcop7gt0Opu
9JMfN9xv++00yK7pPoe+H6lLN9fUmsquGO1XwIfdBqfs1lVxuHdJPqhDyckJ/PawQz7IzfYXV6h1
haNfeSYvvx7aKHkeO7iTYiLmLUYPQTEUoqm+PjMZ+DK4ta3uvPp1rBVdKjnVulqc1PCz8B/Kk9tK
3BvkGQF1p5XE/KzbGbD9iYAPU5ZuJGr6naxBksfcLiXgtyz2DvbtO6Rv0mqgLOseWXee9zmhXn1l
oc8uoV0lWf62XVtrz8aNrfcIDSvclMpPO4UFakDIXB06L1sGYayqYwx6GfFjXmI3eKNVJAqlvi8m
fBxOdGq/kzHfcMx91kBFBe9wr0pOGEJmtr1F3umJEDOXedLrzafpVuskqjKDjZ0hXn00AEkgpGiR
tEcgoZxcuww/qtiXglqPBtVlZ9SY1W59fF1uhopKF/sLVjG5W+7jhFvIb/CM4nzLluproXr03Puf
Xa8IamfbbSOXu80xkAYDBz2ghLCneh3es2S8PFYNDOyq96VlLRVoHlamaSee5Y8giDSU1SlZzXgO
jLAiR1MZ7I94KY+Jw3K3FuFYvNQtXas9XksPjKe7T+othuqWs0yAmiP7hPyi+FMLK4dNmcWsDXLY
bmyh1EHQSDkaWyWgTXHQXmTtzwxRsrH5o6gX3scIrGRfDr2j8e4x6nnQFz9OT+HN4nFenKxJ15Ue
U6brEfkTRbsNf6TEIJMr5hiIoS6Tz6Yy7u9mc3F5LhM0x2xhsudNsw/x7ClKTDOdHEBhFhQ1VuAa
uKqX5KFVYSxzUl+JRvH/sxqoqZUJ6H5Bb1Pc5SJPwUv7oSrDLsYYSqY8KAPNL9Mj9JzDSPbDkiAv
5hh8QDicTq7zbiscp1Q/futEMH+UpWTytE5vFBSd6JoNEUNZ+mSHrauzt/QjpjLmwJKzPxlhPrKA
91HH5iF9NklfbVjStKStRt+Ln4CsXKhM+SPSYF8rLlpqI2/jP7McdBtnf5NieJJRAz/ZwSecVls5
0PZnlnmEBWKbXX+Rp3ARXovyhZy+MmoqRiCeSRCGXejCeh6O8cnhXG4bh5uEhYsc3xqLTnoRjB1G
Z/t2XFcAoGaTabD/DAvmJVHx3YGh4WjXBmEwCxuEe3zqErr9EHSG/rH70TWyBPEm7lA6zxeiFPzP
YCaWooQNtOJ5XnCdyY22xjza2+g3riQOh7buE8CzEsmXGr5Zgvfvn3UYwRjQhrVF5VNjQWz7NviQ
XTrd46iOjHVCKiny1TXl0Y7dkNm/XuwWUe1L4F50hUMLuS3fy0ZTyjcKye/5KGsiTEXbPl5eGZy6
fpeBky00Dsc9RZiOUTRmUZKfakJqAemYFkR7c1HLzU0hcm8tuEZZLRvxaU6JO0K+h13q1xOJWSrT
mK/W2n3J84pjjIwyLCgc6hu/ekh1FXfPZkl4YsAzmpXtcJzkpt5Qdq0qhSJl4tGMz8MLU6ysakBw
qnAzceQ6vFyDWzgogo9yqDMrkgMYJ9Q3ofU1PvsuxM6Rb8MFv7gtlnj6xfmO52gAa5VfTpeV0WXE
TzB3RYrpmAWUD1JNhBNP/LJL6T3NDL+2hSD5ru2SAmmPy0upcvLRHzTXI3StQvQzt3a19ckgmym8
WUQ6m8gFOLu9TxSKfDbIRTW5ASFeglbBQIdpjAvNrw9QmS+xAEITqKAwSYt/CCYedwlhI174PX1i
NW4hBvDu+q0lbizolVmEQaBIWQjRfbpcBeTjbgNLwToKorsTDZbZUo1P7NreLqWDTd1XxKbleJnL
Ve6YXcf4xZS61GH9MwAQqQtyTEVm5b+EyKd6VThsWwrdcbQqaiyUZtI0Yx4Cuf8z+AvGYByEekxp
QTZ4feLskfsX1KWNtTxPDHkzS6zgwgoigzNKXI5SVLrgsvPL3IrzkYZcbbNYtYcHw4635quq3ms8
ati8PKvBRjarK3yEvPfxVab5j72SQZwGhXjQWcV2gn0/umEoWupChaLsrwcr2seKxuYj4XBpRrg/
dMGrteA56Wy36/clX5y5UJSrF1BHwXjAJr9csGz4Se7r1cl7w3xU4clKDk6oFpFH47FNiCExc3qa
kiPWD61f0NtUFPHytQB8j5gxufZkz6kdOpNCoT4YYMQJK9TrwfXmbldBXiQA0aLNFYq3nJd8jDlv
hqrNjkDfdKryIC/Slc0IFBa2Yq/7aY0MflmcqGAfJtENmk2KIX2dxeeqwdrm2WfNVcHT4W9kBF4y
Q9kTDJp5kZUn0lFzgYhTEOgiIfvS50keBlwKfr8nBrGOWJ4ihR78AklC1C+KVMvy3WSerRH+qa6v
4wLuX2kvOOuckecG98NVazRlM8AdbBMH6H/bW8M8E4qbx0MUajJl6MN+zsU+Aq9+kzh8B9TXiMed
8o9JsAKrPZCjIR3LuwgVXER7+TmntoQA1laf8GPJgcJNci94hfSlkVoJGqvN3ZAKjps6Phjy0yqL
p18hSc3tsfuD9S1/Q6ZNdyMjY1z25gOeMsoY97qV1gZ7vCQMAw2c/jFEiXTi728sJispcy6qGSNx
AhjcsbNELt78VHfwn63IDYbCuBQZ2UrFXpgvD++gzm1Y26ex280e4fdUC+OoQVmX9BNq2F0T1g6a
XfveHo4HewDxn6fnsBlkbV/vQ7HuYaVx4THMy22pj8OHE6aVLcrdN3/xCaqL3XX01vP5m+AXOF/5
mvkPxXUdKCiyE4mZUmx1LVJ7VqGXCm3AOVSGfesqkEB1YIkN6oHjHifgVLA53/4e1kPsW2jCGis6
pCA/KQ+dky9w07vAC6o3qO4o3z4ccEdAcidfzRYPhtCvsHnyZY7Dvx+lvHV3jxsZ3gkVh9Tr4ssR
Ql80aeAhzH/69QsvYjFnlpgW+MhGn3RW90eMYu/FFcz1Nu1AnY78QlH32XPOshrAfvXnY/c0ySVW
QKFe9D+ELkT4zoR3VSCgHxzl6DD0YGE3n3w2YxwUUvSe3TBdgZW5F8W54gFRHFMLHymc0hDr2KHZ
BII/eMSNxPFGGR/UF9XhMe7dodOsdU40c5NZtB9zHaaoZAgZOXXXZSg+Hn/YYHXEA/kMvRdVZ0E8
mGEofEVf3i5uHgJF8Kk6kv+ovX60ZBXg51IzLChmaEkLwbe0Qev5VaF9rFetoNRPObWa3DJxLxnx
uyGjXX9pajFIHcfaPcOPNWl03f5VR7zyzLc0OwXlzDyJ2quSb5wMNwBw6uUJ+JGFth7FJ77UXiNE
4tPRHeL6SPNYsFb+MxhiuraszvTLtd7hrbBlGBpJ1FEdhXn3Xa7nlUCZXehusa4atHrZgfqUyFEY
N55h48CsRCa9/qa1DYrIQgrFWb1Y9S1QCFR7CG58Ht3xAJK7UoxWS+irKOtaHr0+dUfOMVVUh2t2
jOhGBMaRYlpBg19uezNdu1mggtzoBxSQLkb0N3JWPb5jHRPR+uJ9DMbeQFXZauzK2qov1Drr7u45
ePLuQaB8Dn5tIYW1vwl5UbNC4Wv0/S8T72KumVj42m+dj9zJfv9N9OfVs163YvHHzlG13uAxkM+6
+XW47if59SVD+WFSeuuVWnWPIfBnKzj2fmCWdB1MRbMOH4Iln9TprCr3rKms1TdbuBFagyJaIYiL
caUPyhOY5a16odaveQ+5idXSv4rgaCgW/0lkrQXkVoj1cznv1KswAL1Z7m+EVMRXn6UgKZGe59AQ
7TlJQFg9EZE/R9jN5EHLbn26XcQ3R8lUV0bPMM6Sn85j1gI2RNFQbx6IOu0bggyj5yyB0Mab6/E7
1tykBWfyLi4kN4QnPctet7vlY8ZZUy5fS4bKlkDfTpdbMLyHsLbcR0QXY5DUvsOMYPemw6iX4H87
yrkrL3RRJ/3/Ad60Zf2D/JPjWCRfPkR28BM9ImQmG+PDPPJm1/gzhGY0XI8Ado1FVBRfPCe6Ko/y
v2bZyjN5VDFalLaJPuuEwNtEVGkzGN0hXCTH44t0smIdjq5ZR4SGZzQ/IWzR49bjG+or1/fQl1xG
q5PrKFJo7tTy9RiheDHKQsAEZREtcFloIfseLTaYcTYvjj+ASjjXZy8rRJzgcK5QIeE83pL9G7w0
VFRcAP8tx7X3Bg6DPlB6kVhVAUoLxZ6WBMrlCTXazdUYJbBquBpkUYRboFV/SGMZqltGIlgkQBj3
H7+49+hdBBKXAj/o7Xo7cXR2ABl0ucVmqcEpzokC9O4FFVa/kMvJaMU2P6J5a6nE3e7PMCnTiPxa
nKNe+Tr/jhP0LbZ4WxuQwJga3A3Qo5QzmjKCLuC/FXbrktyrUJSC9sfEs8rzWuCaH1LvY3ihR1y7
WHYkKXPDfxLvs1Kzc9E3z4gYnlmwFG6O+DAQeOgB0aO/R1mkjhle9yrOtdJwlQeafiwEyjtFD7wP
hHaRCqV7M8u5yAW82GjLABgyO6Mf16Z3l3xrNf+ZoF0k/l3U+vKqaHrbiBTz9y4uwNfX+bott/kh
iW3wdalZOjXLLTlGu5l5CjPgYDKfzwZaAXw2kidjod5lO07uVW8KWKOz0aG10TEHo/mIBfouqUFK
JojW+UQwt0ibmVOyNPLkx9nSN7RUp3T/eb1eDaOBwc93vf5Z36v4IMRZiGCU6Mt5rAnc5GdmxOK4
98IGlm+BA6BkobqdrEaEFFBQw7xgkKC3Z4AGIUStq1plELzwnv2gTAb+hyCTT+T6dyHvylbPMhU1
FFu2z31PTrgSwjWZswyT7GflPtgKJTW5TDkqB4aYsu9cYm/4AZYoKU9a/2yn0OYzt1Urw+ccdfQm
gJWZs4Rjf98mJ0CGYQjJRHN6i9P8Z4hLPX6emJ0QkIoevSkjKn6056C2lnZseHvzWkFzu6erfdVi
8UFEyufEsr97WQfjEUYA2/sVe+0kiTdXrm7JJH7XnysAE5jcws6pdFzi9M4ltcjwsl1KLk9xIkuK
a2y+y7b2jBeW4NbEOmek8Dm8m3gE3cOr7aB5c88rRdb0t3Ix1QEh0vpoSmiC6tf/PjnnCRkVI0QB
UG2g8PHDlcFVu28cQ4HUILJR5kOl3x9b/6VEpwI3erOVj9bH
`protect end_protected
